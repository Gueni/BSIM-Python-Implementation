*** static buffer - modified ***
*
* ngSPICE compensed buffer
*
*
* Author: Jan Belohoubek, 01/2020
* jan.belohoubek@fit.cvut.cz
*
* https://users.fit.cvut.cz/~belohja4/
*
*
* **************************************

.subckt BUFF A O VSS VDD

*** Compensation Inverter Chain ***
XpmosCINV O1 A VDD VDD VSS LaserTrig SUBCKT_PMOS beamDistance = beamDistanceTop ch_w=4u ch_l=0.2u mos_ad=0.6p mos_pd=2.6u mos_as=1p mos_ps=5u
XnmosCINV O1 A VSS VSS psubIn LaserTrig SUBCKT_NMOS beamDistance = beamDistanceBot ch_w=1u ch_l=0.2u mos_ad=0.8p mos_pd=4.8u mos_as=0.5p mos_ps=2.5u

* common NMOS substarte virtual node
XpsubIn psubIn VSS PSUB_IN

XpmosCINV2 O O1 VDD VDD VSS LaserTrig SUBCKT_PMOS beamDistance = beamDistanceTop ch_w=3.5u ch_l=0.2u mos_ad=0.6p mos_pd=2.6u mos_as=1p mos_ps=5u
XnmosCINV2 O O1 VSS VSS psubIn LaserTrig SUBCKT_NMOS beamDistance = beamDistanceBot ch_w=1.5u ch_l=0.2u mos_ad=0.8p mos_pd=4.8u mos_as=0.5p mos_ps=2.5u

.ends
