VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO PNAND2X1
  CLASS BLOCK ;
  FOREIGN PNAND2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.400 BY 10.700 ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.880000 ;
    PORT
      LAYER metal1 ;
        RECT 2.800 4.600 5.500 5.000 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.880000 ;
    PORT
      LAYER metal1 ;
        RECT 2.300 3.900 5.000 4.300 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.400 5.900 9.800 9.600 ;
        RECT 9.400 5.600 9.900 5.900 ;
        RECT 9.500 2.900 9.900 5.600 ;
        RECT 9.400 2.600 9.900 2.900 ;
        RECT 9.400 0.900 9.800 2.600 ;
    END
  END Y
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.200 9.900 10.200 10.500 ;
        RECT 2.200 7.200 2.600 9.900 ;
        RECT 5.400 7.200 5.800 9.900 ;
        RECT 8.600 5.600 9.000 9.900 ;
    END
  END VDD!
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 2.600 6.100 3.000 6.900 ;
        RECT 5.000 6.100 5.400 6.900 ;
        RECT 3.800 0.600 4.200 2.000 ;
        RECT 8.600 0.600 9.000 2.900 ;
        RECT 0.600 0.000 9.900 0.600 ;
      LAYER via1 ;
        RECT 3.800 0.100 4.200 0.500 ;
      LAYER metal2 ;
        RECT 2.600 6.100 5.400 6.500 ;
        RECT 3.800 0.000 4.200 6.100 ;
    END
  END GND!
  OBS
      LAYER metal1 ;
        RECT 0.600 7.600 1.000 9.600 ;
        RECT 1.400 7.600 1.800 9.600 ;
        RECT 0.600 5.800 1.000 7.300 ;
        RECT 3.000 7.200 3.400 9.600 ;
        RECT 3.800 7.200 4.200 9.600 ;
        RECT 4.600 7.200 5.000 9.600 ;
        RECT 6.200 7.600 6.600 9.600 ;
        RECT 7.000 7.600 7.400 9.600 ;
        RECT 7.000 5.800 7.400 7.300 ;
        RECT 7.800 5.800 8.200 9.600 ;
        RECT 0.600 5.400 8.200 5.800 ;
        RECT 1.400 2.300 6.600 2.700 ;
        RECT 2.000 1.000 2.400 2.300 ;
        RECT 5.600 1.000 6.000 2.300 ;
        RECT 7.800 0.900 8.200 5.400 ;
        RECT 8.700 3.600 9.200 4.000 ;
      LAYER via1 ;
        RECT 1.400 9.200 1.800 9.600 ;
        RECT 3.000 9.200 3.400 9.600 ;
        RECT 3.800 7.600 4.200 8.000 ;
        RECT 4.600 9.200 5.000 9.600 ;
        RECT 6.200 9.200 6.600 9.600 ;
        RECT 6.200 2.300 6.600 2.700 ;
        RECT 8.800 3.600 9.200 4.000 ;
      LAYER metal2 ;
        RECT 1.400 9.200 6.600 9.600 ;
        RECT 0.600 7.600 7.400 8.000 ;
        RECT 1.400 2.300 1.800 7.600 ;
        RECT 6.200 4.000 6.600 7.600 ;
        RECT 6.200 3.600 9.200 4.000 ;
        RECT 6.200 2.300 6.600 3.600 ;
  END
END PNAND2X1
END LIBRARY

