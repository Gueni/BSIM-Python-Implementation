magic
tech scmos
timestamp 1600391712
<< nwell >>
rect 12 48 142 105
<< ntransistor >>
rect 31 7 33 21
rect 36 7 38 21
rect 44 7 46 21
rect 49 7 51 21
rect 97 7 99 26
rect 105 7 107 26
rect 121 7 123 26
rect 129 7 131 21
<< ptransistor >>
rect 31 79 33 93
rect 36 79 38 93
rect 44 79 46 93
rect 49 79 51 93
rect 57 79 59 93
rect 73 68 75 93
rect 81 68 83 93
rect 97 54 99 93
rect 105 54 107 93
rect 121 89 123 93
rect 129 66 131 93
<< ndiffusion >>
rect 30 7 31 21
rect 33 7 36 21
rect 38 7 39 21
rect 43 7 44 21
rect 46 7 49 21
rect 51 7 52 21
rect 96 7 97 26
rect 99 7 100 26
rect 104 7 105 26
rect 107 7 108 26
rect 120 7 121 26
rect 123 7 124 26
rect 128 7 129 21
rect 131 7 132 21
<< pdiffusion >>
rect 30 79 31 93
rect 33 79 36 93
rect 38 79 39 93
rect 43 79 44 93
rect 46 79 49 93
rect 51 79 52 93
rect 56 79 57 93
rect 59 79 60 93
rect 72 68 73 93
rect 75 68 76 93
rect 80 68 81 93
rect 83 68 84 93
rect 96 54 97 93
rect 99 54 100 93
rect 104 54 105 93
rect 107 54 108 93
rect 120 89 121 93
rect 123 89 124 93
rect 128 66 129 93
rect 131 66 132 93
<< ndcontact >>
rect 26 7 30 21
rect 39 7 43 21
rect 52 7 56 21
rect 92 7 96 26
rect 100 7 104 26
rect 108 7 112 26
rect 116 7 120 26
rect 124 7 128 26
rect 132 7 136 21
<< pdcontact >>
rect 26 79 30 93
rect 39 79 43 93
rect 52 79 56 93
rect 60 79 64 93
rect 68 68 72 93
rect 76 68 80 93
rect 84 68 88 93
rect 92 54 96 93
rect 100 54 104 93
rect 108 54 112 93
rect 116 89 120 93
rect 124 66 128 93
rect 132 66 136 93
<< psubstratepcontact >>
rect 33 -2 37 2
<< nsubstratencontact >>
rect 60 98 64 102
rect 124 98 128 102
<< polysilicon >>
rect 31 93 33 95
rect 36 93 38 95
rect 44 93 46 95
rect 49 93 51 95
rect 57 93 59 95
rect 73 93 75 95
rect 81 93 83 95
rect 97 93 99 95
rect 105 93 107 95
rect 121 93 123 95
rect 129 93 131 95
rect 31 50 33 79
rect 31 21 33 46
rect 36 42 38 79
rect 44 50 46 79
rect 49 42 51 79
rect 36 24 39 26
rect 43 24 46 26
rect 36 21 38 24
rect 44 21 46 24
rect 49 21 51 38
rect 31 5 33 7
rect 36 5 38 7
rect 44 5 46 7
rect 49 5 51 7
rect 57 2 59 79
rect 73 28 75 68
rect 81 28 83 68
rect 97 43 99 54
rect 105 43 107 54
rect 97 39 98 43
rect 105 39 114 43
rect 97 26 99 39
rect 105 26 107 39
rect 121 26 123 89
rect 129 35 131 66
rect 130 31 131 35
rect 129 21 131 31
rect 97 5 99 7
rect 105 5 107 7
rect 121 2 123 7
rect 129 5 131 7
<< polycontact >>
rect 29 46 33 50
rect 42 46 46 50
rect 36 38 40 42
rect 49 38 53 42
rect 39 24 43 28
rect 71 24 75 28
rect 79 24 83 28
rect 98 39 102 43
rect 114 39 118 43
rect 126 31 130 35
rect 56 -2 60 2
rect 120 -2 124 2
<< metal1 >>
rect 14 102 140 103
rect 14 98 60 102
rect 64 98 124 102
rect 128 98 140 102
rect 14 97 140 98
rect 60 93 64 97
rect 100 93 104 97
rect 124 93 128 97
rect 39 57 43 79
rect 68 57 72 68
rect 39 53 72 57
rect 33 46 42 50
rect 40 38 49 42
rect 68 35 72 53
rect 84 35 88 68
rect 26 31 84 35
rect 26 21 30 31
rect 91 28 95 54
rect 107 43 111 54
rect 116 43 120 89
rect 102 39 111 43
rect 118 39 120 43
rect 43 24 71 28
rect 75 24 79 28
rect 83 26 95 28
rect 107 26 111 39
rect 116 26 120 39
rect 133 57 136 66
rect 125 31 126 35
rect 83 24 92 26
rect 56 17 84 21
rect 133 21 137 57
rect 136 17 137 21
rect 39 3 43 7
rect 100 3 104 7
rect 124 3 128 7
rect 14 2 140 3
rect 14 -2 33 2
rect 37 -2 56 2
rect 60 -2 120 2
rect 124 -2 140 2
rect 14 -3 140 -2
<< m2contact >>
rect 26 81 30 85
rect 52 81 56 85
rect 76 81 80 85
rect 84 31 88 35
rect 126 31 130 35
rect 84 17 88 21
<< metal2 >>
rect 30 81 52 85
rect 56 81 76 85
rect 88 31 126 35
rect 84 21 88 31
<< metal4 >>
rect 59 2 65 3
rect 56 -1 65 2
rect 56 -2 60 -1
<< labels >>
rlabel space 1 -3 105 104 1 vdd
rlabel space 1 -3 105 104 1 gnd
rlabel metal1 35 100 35 100 1 VDD!
port 1 n power bidirectional
rlabel ptransistor 31 85 31 85 1 S$
rlabel ptransistor 33 85 33 85 1 D$
rlabel ptransistor 49 85 49 85 1 D$
rlabel ptransistor 51 85 51 85 1 S$
rlabel ptransistor 44 85 44 85 1 D$
rlabel ptransistor 38 85 38 85 1 D$
rlabel ptransistor 36 85 36 85 1 S$
rlabel ptransistor 46 85 46 85 1 S$
rlabel ptransistor 57 85 57 85 1 D$
rlabel ptransistor 59 85 59 85 1 S$
rlabel metal1 29 -1 29 -1 1 GND!
port 2 n power bidirectional
rlabel polycontact 29 46 29 50 1 B
port 3 n signal input
rlabel space -4 -3 110 105 1 vdd
rlabel space -4 -3 110 105 1 gnd
rlabel polycontact 36 38 36 42 1 A
port 4 n signal input
rlabel ptransistor 75 86 75 86 1 S$
rlabel ptransistor 73 85 73 85 1 D$
rlabel ntransistor 51 9 51 9 1 D$
rlabel ntransistor 49 9 49 9 1 S$
rlabel ntransistor 31 9 31 9 1 D$
rlabel ntransistor 33 9 33 9 1 S$
rlabel pdcontact 54 86 54 86 1 VVDD
rlabel ntransistor 131 19 131 19 1 D$
rlabel ntransistor 129 19 129 19 1 S$
rlabel metal1 137 53 137 57 1 Y
port 5 n signal output
rlabel ntransistor 121 16 121 16 1 D$
rlabel ntransistor 123 16 123 16 1 S$
rlabel ptransistor 123 92 123 92 1 S$
rlabel ptransistor 121 92 121 92 1 D$
rlabel ptransistor 131 92 131 92 1 D$
rlabel ptransistor 129 92 129 92 1 S$
rlabel m2contact 86 33 86 33 1 O
rlabel space -4 -3 142 105 1 vdd
rlabel space -4 -3 142 105 1 gnd
<< end >>
