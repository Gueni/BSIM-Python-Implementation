VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX1
  CLASS BLOCK ;
  FOREIGN INVX1 ;
  ORIGIN 0.900 0.300 ;
  SIZE 3.500 BY 10.800 ;
  OBS
      LAYER metal1 ;
        RECT -0.200 9.700 1.800 10.300 ;
        RECT 0.200 7.400 0.600 9.700 ;
        RECT 0.200 1.900 0.600 2.700 ;
        RECT 0.200 0.300 0.600 1.600 ;
        RECT 1.000 0.600 1.400 9.400 ;
        RECT -0.200 -0.300 1.800 0.300 ;
  END
END INVX1
MACRO NOR3X1
  CLASS BLOCK ;
  FOREIGN NOR3X1 ;
  ORIGIN 0.700 0.300 ;
  SIZE 7.500 BY 10.800 ;
  OBS
      LAYER metal1 ;
        RECT -0.200 9.700 6.600 10.300 ;
        RECT 0.200 6.400 0.600 9.400 ;
        RECT 1.000 6.400 1.400 9.700 ;
        RECT 1.800 9.100 3.800 9.400 ;
        RECT 1.800 6.400 2.200 9.100 ;
        RECT 2.600 6.400 3.000 8.800 ;
        RECT 3.400 6.500 3.800 9.100 ;
        RECT 4.300 9.100 6.100 9.400 ;
        RECT 4.300 9.000 4.600 9.100 ;
        RECT 0.300 6.100 0.600 6.400 ;
        RECT 1.800 6.100 2.100 6.400 ;
        RECT 0.300 5.800 2.100 6.100 ;
        RECT 2.700 6.200 3.000 6.400 ;
        RECT 4.200 6.200 4.600 9.000 ;
        RECT 5.800 9.000 6.100 9.100 ;
        RECT 2.700 6.000 4.600 6.200 ;
        RECT 5.000 6.000 5.400 8.800 ;
        RECT 5.800 6.000 6.200 9.000 ;
        RECT 2.700 5.900 4.500 6.000 ;
        RECT 5.000 5.700 5.300 6.000 ;
        RECT 5.000 5.600 5.400 5.700 ;
        RECT 3.700 5.300 5.400 5.600 ;
        RECT 2.600 4.300 3.400 4.700 ;
        RECT 1.800 3.300 2.600 3.700 ;
        RECT 1.000 2.300 1.900 2.700 ;
        RECT 3.700 2.000 4.000 5.300 ;
        RECT 2.000 1.700 4.000 2.000 ;
        RECT 2.000 1.600 2.300 1.700 ;
        RECT 1.000 0.300 1.400 1.600 ;
        RECT 1.800 1.300 2.300 1.600 ;
        RECT 3.400 1.600 4.000 1.700 ;
        RECT 1.800 0.600 2.200 1.300 ;
        RECT 2.600 0.300 3.000 1.400 ;
        RECT 3.400 0.600 3.800 1.600 ;
        RECT -0.200 -0.300 6.600 0.300 ;
  END
END NOR3X1
MACRO CELM2X1
  CLASS BLOCK ;
  FOREIGN CELM2X1 ;
  ORIGIN 0.800 0.300 ;
  SIZE 4.500 BY 10.800 ;
  OBS
      LAYER metal1 ;
        RECT -0.200 9.700 3.100 10.300 ;
        RECT 0.200 7.400 0.600 9.400 ;
        RECT 1.500 7.400 1.900 9.700 ;
        RECT 2.300 7.700 2.700 9.400 ;
        RECT 2.300 7.400 2.800 7.700 ;
        RECT 0.300 7.100 1.200 7.400 ;
        RECT 0.900 6.800 1.200 7.100 ;
        RECT 0.900 6.500 2.200 6.800 ;
        RECT 0.700 5.300 1.600 5.700 ;
        RECT 1.200 4.900 1.600 5.300 ;
        RECT 0.200 3.300 0.600 4.100 ;
        RECT 1.900 3.500 2.200 6.500 ;
        RECT 0.900 3.200 2.200 3.500 ;
        RECT 0.900 2.900 1.200 3.200 ;
        RECT 1.800 3.100 2.200 3.200 ;
        RECT 2.500 6.700 2.800 7.400 ;
        RECT 2.500 6.300 3.000 6.700 ;
        RECT 0.300 2.600 1.200 2.900 ;
        RECT 0.200 0.600 0.600 2.600 ;
        RECT 1.500 0.300 1.900 2.600 ;
        RECT 2.500 1.900 2.800 6.300 ;
        RECT 2.300 1.600 2.800 1.900 ;
        RECT 2.300 0.600 2.700 1.600 ;
        RECT -0.200 -0.300 3.100 0.300 ;
  END
END CELM2X1
MACRO SECLIBAND_opt
  CLASS BLOCK ;
  FOREIGN SECLIBAND_opt ;
  ORIGIN 0.800 0.300 ;
  SIZE 32.500 BY 10.800 ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.600000 ;
    PORT
      LAYER metal1 ;
        RECT 3.600 5.300 4.500 5.700 ;
        RECT 9.400 5.300 10.300 5.700 ;
        RECT 4.100 4.900 4.500 5.300 ;
        RECT 9.900 4.900 10.300 5.300 ;
      LAYER metal2 ;
        RECT 4.100 4.900 10.300 5.300 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.000000 ;
    PORT
      LAYER metal1 ;
        RECT 3.100 7.400 3.500 9.400 ;
        RECT 3.200 7.100 4.100 7.400 ;
        RECT 3.800 6.800 4.100 7.100 ;
        RECT 3.800 6.500 5.100 6.800 ;
        RECT 0.200 3.300 0.600 4.100 ;
        RECT 3.100 2.900 3.500 4.100 ;
        RECT 4.800 3.500 5.100 6.500 ;
        RECT 3.800 3.200 5.100 3.500 ;
        RECT 6.000 3.300 6.400 4.100 ;
        RECT 3.800 2.900 4.100 3.200 ;
        RECT 4.700 3.100 5.100 3.200 ;
        RECT 3.200 2.600 4.100 2.900 ;
        RECT 3.100 0.600 3.500 2.600 ;
      LAYER via1 ;
        RECT 3.100 3.300 3.500 3.700 ;
      LAYER metal2 ;
        RECT 0.200 3.300 6.400 3.700 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.600000 ;
    PORT
      LAYER metal1 ;
        RECT 6.500 5.700 6.900 6.100 ;
        RECT 12.300 5.700 12.700 6.100 ;
        RECT 6.500 5.300 7.400 5.700 ;
        RECT 12.300 5.300 13.200 5.700 ;
        RECT 7.000 4.900 7.400 5.300 ;
        RECT 12.800 4.500 13.200 5.300 ;
      LAYER metal2 ;
        RECT 6.500 5.700 12.700 6.100 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.400000 ;
    PORT
      LAYER metal1 ;
        RECT 0.700 5.300 1.600 5.700 ;
        RECT 1.200 4.900 1.600 5.300 ;
        RECT 8.900 3.300 9.300 4.500 ;
        RECT 11.800 3.300 12.200 4.500 ;
      LAYER via1 ;
        RECT 8.900 4.100 9.300 4.500 ;
        RECT 11.800 4.100 12.200 4.500 ;
      LAYER metal2 ;
        RECT 1.200 4.500 1.600 5.300 ;
        RECT 1.200 4.100 12.200 4.500 ;
    END
  END A1
  PIN Y0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 28.500 0.600 28.900 9.400 ;
    END
  END Y0
  PIN Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 30.100 0.600 30.500 9.400 ;
    END
  END Y1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -0.200 9.700 30.900 10.300 ;
        RECT 1.500 7.400 1.900 9.700 ;
        RECT 4.400 7.400 4.800 9.700 ;
        RECT 7.300 7.400 7.700 9.700 ;
        RECT 10.200 7.400 10.600 9.700 ;
        RECT 13.100 7.400 13.500 9.700 ;
        RECT 15.700 6.400 16.100 9.700 ;
        RECT 22.100 6.400 22.500 9.700 ;
        RECT 27.700 7.400 28.100 9.700 ;
        RECT 29.300 7.400 29.700 9.700 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 1.500 0.300 1.900 2.600 ;
        RECT 4.400 0.300 4.800 2.600 ;
        RECT 7.300 0.300 7.700 2.600 ;
        RECT 10.200 0.300 10.600 2.600 ;
        RECT 13.100 0.300 13.500 2.600 ;
        RECT 15.700 0.300 16.100 1.600 ;
        RECT 17.300 0.300 17.700 1.400 ;
        RECT 22.100 0.300 22.500 1.600 ;
        RECT 23.700 0.300 24.100 1.400 ;
        RECT 27.700 0.300 28.100 1.600 ;
        RECT 29.300 0.300 29.700 1.600 ;
        RECT -0.200 -0.300 30.900 0.300 ;
    END
  END GND
  OBS
      LAYER metal1 ;
        RECT 0.200 7.400 0.600 9.400 ;
        RECT 2.300 7.700 2.700 9.400 ;
        RECT 5.200 7.700 5.600 9.400 ;
        RECT 2.300 7.400 2.800 7.700 ;
        RECT 5.200 7.400 5.700 7.700 ;
        RECT 6.000 7.400 6.400 9.400 ;
        RECT 8.100 7.700 8.500 9.400 ;
        RECT 8.100 7.400 8.600 7.700 ;
        RECT 8.900 7.400 9.300 9.400 ;
        RECT 11.000 7.700 11.400 9.400 ;
        RECT 11.000 7.400 11.500 7.700 ;
        RECT 11.800 7.400 12.200 9.400 ;
        RECT 13.900 7.700 14.300 9.400 ;
        RECT 13.900 7.400 14.400 7.700 ;
        RECT 0.300 7.100 1.200 7.400 ;
        RECT 0.900 6.800 1.200 7.100 ;
        RECT 0.900 6.500 2.200 6.800 ;
        RECT 1.900 3.500 2.200 6.500 ;
        RECT 0.900 3.200 2.200 3.500 ;
        RECT 0.900 2.900 1.200 3.200 ;
        RECT 1.800 3.100 2.200 3.200 ;
        RECT 2.500 6.700 2.800 7.400 ;
        RECT 5.400 6.800 5.700 7.400 ;
        RECT 6.100 7.100 7.000 7.400 ;
        RECT 6.700 6.800 7.000 7.100 ;
        RECT 5.400 6.700 5.800 6.800 ;
        RECT 2.500 6.300 3.000 6.700 ;
        RECT 5.400 6.300 5.900 6.700 ;
        RECT 6.700 6.500 8.000 6.800 ;
        RECT 0.300 2.600 1.200 2.900 ;
        RECT 0.200 0.600 0.600 2.600 ;
        RECT 2.500 2.000 2.800 6.300 ;
        RECT 2.400 1.900 2.800 2.000 ;
        RECT 5.400 1.900 5.700 6.300 ;
        RECT 7.700 3.500 8.000 6.500 ;
        RECT 6.700 3.200 8.000 3.500 ;
        RECT 6.700 2.900 7.000 3.200 ;
        RECT 7.600 3.100 8.000 3.200 ;
        RECT 8.300 6.700 8.600 7.400 ;
        RECT 9.000 7.100 9.900 7.400 ;
        RECT 9.600 6.800 9.900 7.100 ;
        RECT 8.300 6.300 8.800 6.700 ;
        RECT 9.600 6.500 10.900 6.800 ;
        RECT 6.100 2.600 7.000 2.900 ;
        RECT 8.300 2.700 8.600 6.300 ;
        RECT 10.600 3.500 10.900 6.500 ;
        RECT 9.600 3.200 10.900 3.500 ;
        RECT 9.600 2.900 9.900 3.200 ;
        RECT 10.500 3.100 10.900 3.200 ;
        RECT 11.200 6.700 11.500 7.400 ;
        RECT 11.900 7.100 12.800 7.400 ;
        RECT 12.500 6.800 12.800 7.100 ;
        RECT 11.200 6.300 11.700 6.700 ;
        RECT 12.500 6.500 13.800 6.800 ;
        RECT 11.200 5.300 11.500 6.300 ;
        RECT 11.200 4.900 11.600 5.300 ;
        RECT 2.300 1.600 2.800 1.900 ;
        RECT 5.200 1.600 5.700 1.900 ;
        RECT 2.300 0.600 2.700 1.600 ;
        RECT 5.200 0.600 5.600 1.600 ;
        RECT 6.000 0.600 6.400 2.600 ;
        RECT 8.200 2.300 8.600 2.700 ;
        RECT 9.000 2.600 9.900 2.900 ;
        RECT 8.300 1.900 8.600 2.300 ;
        RECT 8.100 1.600 8.600 1.900 ;
        RECT 8.100 0.600 8.500 1.600 ;
        RECT 8.900 0.600 9.300 2.600 ;
        RECT 11.200 1.900 11.500 4.900 ;
        RECT 13.500 3.500 13.800 6.500 ;
        RECT 12.500 3.200 13.800 3.500 ;
        RECT 12.500 2.900 12.800 3.200 ;
        RECT 13.400 3.100 13.800 3.200 ;
        RECT 14.100 6.700 14.400 7.400 ;
        RECT 14.100 6.300 14.600 6.700 ;
        RECT 14.900 6.400 15.300 9.400 ;
        RECT 14.100 3.500 14.400 6.300 ;
        RECT 15.000 6.100 15.300 6.400 ;
        RECT 16.500 9.100 18.500 9.400 ;
        RECT 16.500 6.400 16.900 9.100 ;
        RECT 17.300 6.400 17.700 8.800 ;
        RECT 18.100 6.500 18.500 9.100 ;
        RECT 19.000 9.100 20.800 9.400 ;
        RECT 19.000 9.000 19.300 9.100 ;
        RECT 16.500 6.100 16.800 6.400 ;
        RECT 15.000 5.800 16.800 6.100 ;
        RECT 17.400 6.200 17.700 6.400 ;
        RECT 18.900 6.200 19.300 9.000 ;
        RECT 20.500 9.000 20.800 9.100 ;
        RECT 17.400 6.000 19.300 6.200 ;
        RECT 19.700 6.000 20.100 8.800 ;
        RECT 20.500 6.000 20.900 9.000 ;
        RECT 21.300 6.400 21.700 9.400 ;
        RECT 21.400 6.100 21.700 6.400 ;
        RECT 22.900 9.100 24.900 9.400 ;
        RECT 22.900 6.400 23.300 9.100 ;
        RECT 23.700 6.400 24.100 8.800 ;
        RECT 24.500 6.500 24.900 9.100 ;
        RECT 25.400 9.100 27.200 9.400 ;
        RECT 25.400 9.000 25.700 9.100 ;
        RECT 22.900 6.100 23.200 6.400 ;
        RECT 17.400 5.900 19.200 6.000 ;
        RECT 19.700 5.700 20.000 6.000 ;
        RECT 21.400 5.800 23.200 6.100 ;
        RECT 23.800 6.200 24.100 6.400 ;
        RECT 25.300 6.200 25.700 9.000 ;
        RECT 26.900 9.000 27.200 9.100 ;
        RECT 23.800 6.000 25.700 6.200 ;
        RECT 26.100 6.000 26.500 8.800 ;
        RECT 26.900 6.000 27.300 9.000 ;
        RECT 23.800 5.900 25.600 6.000 ;
        RECT 26.100 5.700 26.400 6.000 ;
        RECT 19.700 5.600 20.100 5.700 ;
        RECT 26.100 5.600 26.500 5.700 ;
        RECT 18.400 5.300 20.100 5.600 ;
        RECT 24.800 5.300 26.500 5.600 ;
        RECT 29.200 5.300 29.700 5.700 ;
        RECT 16.500 3.700 16.900 5.000 ;
        RECT 17.300 4.300 18.100 4.700 ;
        RECT 14.100 3.100 14.500 3.500 ;
        RECT 16.500 3.300 17.300 3.700 ;
        RECT 11.900 2.600 12.800 2.900 ;
        RECT 11.000 1.600 11.500 1.900 ;
        RECT 11.000 0.600 11.400 1.600 ;
        RECT 11.800 0.600 12.200 2.600 ;
        RECT 14.100 1.900 14.400 3.100 ;
        RECT 15.700 2.300 16.600 2.700 ;
        RECT 18.400 2.000 18.700 5.300 ;
        RECT 22.100 4.300 24.500 4.700 ;
        RECT 22.100 2.700 22.500 4.300 ;
        RECT 22.900 3.300 23.700 3.700 ;
        RECT 22.900 3.100 23.300 3.300 ;
        RECT 22.100 2.300 23.000 2.700 ;
        RECT 24.800 2.000 25.100 5.300 ;
        RECT 27.700 2.300 28.100 2.700 ;
        RECT 13.900 1.600 14.400 1.900 ;
        RECT 16.700 1.700 18.700 2.000 ;
        RECT 16.700 1.600 17.000 1.700 ;
        RECT 13.900 0.600 14.300 1.600 ;
        RECT 16.500 1.300 17.000 1.600 ;
        RECT 18.100 1.600 18.700 1.700 ;
        RECT 23.100 1.700 25.100 2.000 ;
        RECT 23.100 1.600 23.400 1.700 ;
        RECT 16.500 0.600 16.900 1.300 ;
        RECT 18.100 1.100 18.500 1.600 ;
        RECT 22.900 1.300 23.400 1.600 ;
        RECT 24.500 1.600 25.100 1.700 ;
        RECT 26.700 1.900 28.100 2.300 ;
        RECT 29.300 1.900 29.700 5.300 ;
        RECT 18.100 0.700 18.900 1.100 ;
        RECT 18.100 0.600 18.500 0.700 ;
        RECT 22.900 0.600 23.300 1.300 ;
        RECT 24.500 0.600 24.900 1.600 ;
        RECT 26.700 0.700 27.100 1.900 ;
      LAYER via1 ;
        RECT 5.400 6.400 5.800 6.800 ;
        RECT 2.400 1.600 2.800 2.000 ;
        RECT 26.100 5.300 26.500 5.700 ;
        RECT 16.500 4.600 16.900 5.000 ;
        RECT 18.500 0.700 18.900 1.100 ;
      LAYER metal2 ;
        RECT 5.400 6.400 17.700 6.800 ;
        RECT 11.200 4.900 16.900 5.300 ;
        RECT 16.500 4.600 16.900 4.900 ;
        RECT 17.300 4.300 17.700 6.400 ;
        RECT 26.100 5.300 29.600 5.700 ;
        RECT 14.100 3.100 23.300 3.500 ;
        RECT 8.200 2.300 16.100 2.700 ;
        RECT 22.100 2.000 22.500 2.700 ;
        RECT 2.300 1.600 22.500 2.000 ;
        RECT 18.500 0.700 27.100 1.100 ;
  END
END SECLIBAND_opt
END LIBRARY

