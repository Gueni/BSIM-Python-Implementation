VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO PNOR2X1
  CLASS BLOCK ;
  FOREIGN PNOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.400 BY 10.700 ;
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.200 9.900 11.200 10.500 ;
        RECT 2.200 7.200 2.600 9.900 ;
        RECT 6.400 7.200 6.800 9.900 ;
        RECT 9.600 5.600 10.000 9.900 ;
    END
  END VDD!
  PIN GND!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 2.500 6.100 2.900 6.900 ;
        RECT 6.100 6.100 6.500 6.900 ;
        RECT 4.300 0.600 4.700 2.000 ;
        RECT 9.600 0.600 10.000 2.900 ;
        RECT 0.600 0.000 10.900 0.600 ;
      LAYER via1 ;
        RECT 4.300 0.100 4.700 0.500 ;
      LAYER metal2 ;
        RECT 2.500 6.100 6.500 6.500 ;
        RECT 4.300 0.000 4.700 6.100 ;
    END
  END GND!
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.160000 ;
    PORT
      LAYER metal1 ;
        RECT 3.100 4.600 5.300 5.000 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.160000 ;
    PORT
      LAYER metal1 ;
        RECT 3.700 3.900 5.900 4.300 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 10.400 5.900 10.800 9.600 ;
        RECT 10.400 5.600 10.900 5.900 ;
        RECT 10.500 2.900 10.900 5.600 ;
        RECT 10.400 2.600 10.900 2.900 ;
        RECT 10.400 0.900 10.800 2.600 ;
    END
  END Y
  OBS
      LAYER metal1 ;
        RECT 0.600 7.600 1.000 9.600 ;
        RECT 1.400 7.600 1.800 9.600 ;
        RECT 0.600 5.800 1.000 7.300 ;
        RECT 3.000 7.200 3.400 9.600 ;
        RECT 4.300 7.200 4.700 9.600 ;
        RECT 5.600 7.200 6.000 9.600 ;
        RECT 7.200 7.600 7.600 9.600 ;
        RECT 8.000 7.600 8.400 9.600 ;
        RECT 8.000 5.800 8.400 7.300 ;
        RECT 8.800 5.800 9.200 9.600 ;
        RECT 0.600 5.400 9.200 5.800 ;
        RECT 1.400 2.300 7.600 2.700 ;
        RECT 3.000 1.000 3.400 2.300 ;
        RECT 5.600 1.000 6.000 2.300 ;
        RECT 8.800 0.900 9.200 5.400 ;
        RECT 9.700 3.600 10.200 4.000 ;
      LAYER via1 ;
        RECT 1.400 9.200 1.800 9.600 ;
        RECT 3.000 9.200 3.400 9.600 ;
        RECT 4.300 7.600 4.700 8.000 ;
        RECT 5.600 9.200 6.000 9.600 ;
        RECT 7.200 9.200 7.600 9.600 ;
        RECT 7.200 2.300 7.600 2.700 ;
        RECT 9.800 3.600 10.200 4.000 ;
      LAYER metal2 ;
        RECT 1.400 9.200 7.600 9.600 ;
        RECT 0.600 7.600 8.400 8.000 ;
        RECT 1.400 2.300 1.800 7.600 ;
        RECT 7.200 4.000 7.600 7.600 ;
        RECT 7.200 3.600 10.200 4.000 ;
        RECT 7.200 2.300 7.600 3.600 ;
  END
END PNOR2X1
END LIBRARY

