magic
tech scmos
magscale 1 2
timestamp 1598350919
<< error_s >>
rect 2300 3616 2308 3624
rect 1068 3576 1076 3584
rect 764 3556 772 3564
rect 2060 3556 2068 3564
rect 316 3536 324 3544
rect 2460 3536 2468 3544
rect 2524 3536 2532 3544
rect 332 3516 340 3524
rect 1948 3516 1956 3524
rect 2012 3516 2020 3524
rect 2108 3516 2116 3524
rect 2156 3516 2164 3524
rect 2220 3516 2228 3524
rect 2668 3516 2676 3524
rect 2780 3516 2788 3524
rect 2924 3516 2932 3524
rect 3404 3516 3412 3524
rect 3468 3516 3476 3524
rect 4380 3516 4388 3524
rect 4412 3516 4420 3524
rect 4460 3516 4468 3524
rect 1212 3496 1220 3504
rect 1244 3496 1252 3504
rect 1260 3496 1268 3504
rect 1436 3496 1444 3504
rect 4572 3496 4580 3504
rect 4716 3496 4724 3504
rect 4812 3496 4820 3504
rect 4828 3496 4836 3504
rect 156 3476 164 3484
rect 348 3476 356 3484
rect 508 3476 516 3484
rect 716 3476 724 3484
rect 1340 3476 1348 3484
rect 1388 3476 1396 3484
rect 1852 3476 1860 3484
rect 3452 3476 3460 3484
rect 3804 3476 3812 3484
rect 3948 3476 3956 3484
rect 3964 3476 3972 3484
rect 3980 3476 3988 3484
rect 4300 3476 4308 3484
rect 5004 3476 5012 3484
rect 5132 3476 5140 3484
rect 236 3456 244 3464
rect 828 3456 836 3464
rect 924 3456 932 3464
rect 1196 3456 1204 3464
rect 1628 3456 1636 3464
rect 1708 3456 1716 3464
rect 2492 3456 2500 3464
rect 3436 3456 3444 3464
rect 3516 3456 3524 3464
rect 3532 3456 3540 3464
rect 4236 3456 4244 3464
rect 4556 3456 4564 3464
rect 4668 3456 4676 3464
rect 4700 3456 4708 3464
rect 4956 3456 4964 3464
rect 124 3436 132 3444
rect 636 3436 644 3444
rect 1164 3436 1172 3444
rect 1724 3436 1732 3444
rect 1916 3436 1924 3444
rect 2076 3436 2084 3444
rect 3276 3436 3284 3444
rect 3324 3436 3332 3444
rect 3340 3436 3348 3444
rect 4044 3436 4052 3444
rect 4156 3436 4164 3444
rect 4396 3436 4404 3444
rect 4444 3436 4452 3444
rect 4492 3436 4500 3444
rect 4604 3436 4612 3444
rect 4684 3436 4692 3444
rect 4732 3436 4740 3444
rect 4940 3436 4948 3444
rect 716 3416 724 3424
rect 1036 3416 1044 3424
rect 1084 3416 1092 3424
rect 2300 3416 2308 3424
rect 2316 3416 2324 3424
rect 2796 3416 2804 3424
rect 2972 3416 2980 3424
rect 3900 3416 3908 3424
rect 4092 3416 4100 3424
rect 1116 3396 1124 3404
rect 1292 3396 1300 3404
rect 2236 3396 2244 3404
rect 2908 3396 2916 3404
rect 3004 3396 3012 3404
rect 3020 3396 3028 3404
rect 3244 3396 3252 3404
rect 3388 3396 3396 3404
rect 3724 3396 3732 3404
rect 3804 3396 3812 3404
rect 4108 3396 4116 3404
rect 156 3376 164 3384
rect 348 3376 356 3384
rect 588 3376 596 3384
rect 636 3376 644 3384
rect 3148 3376 3156 3384
rect 3484 3376 3492 3384
rect 4460 3376 4468 3384
rect 4476 3376 4484 3384
rect 4764 3376 4772 3384
rect 5052 3376 5060 3384
rect 12 3356 20 3364
rect 60 3356 68 3364
rect 300 3356 308 3364
rect 972 3356 980 3364
rect 1020 3356 1028 3364
rect 1116 3356 1124 3364
rect 1292 3356 1300 3364
rect 1308 3356 1316 3364
rect 1324 3356 1332 3364
rect 1388 3356 1396 3364
rect 1612 3356 1620 3364
rect 2124 3356 2132 3364
rect 2156 3356 2164 3364
rect 2396 3356 2404 3364
rect 2444 3356 2452 3364
rect 2476 3356 2484 3364
rect 2572 3356 2580 3364
rect 2700 3356 2708 3364
rect 2844 3356 2852 3364
rect 3052 3356 3060 3364
rect 3340 3356 3348 3364
rect 3388 3356 3396 3364
rect 3500 3356 3508 3364
rect 3708 3356 3716 3364
rect 3788 3356 3796 3364
rect 3996 3356 4004 3364
rect 4380 3356 4388 3364
rect 4396 3356 4404 3364
rect 4508 3356 4516 3364
rect 4844 3356 4852 3364
rect 5132 3356 5140 3364
rect 284 3336 292 3344
rect 364 3336 372 3344
rect 572 3336 580 3344
rect 764 3336 772 3344
rect 796 3336 804 3344
rect 812 3336 820 3344
rect 1020 3336 1028 3344
rect 1148 3336 1156 3344
rect 1164 3336 1172 3344
rect 1276 3336 1284 3344
rect 1788 3336 1796 3344
rect 3372 3336 3380 3344
rect 3404 3336 3412 3344
rect 3436 3336 3444 3344
rect 3452 3336 3460 3344
rect 3964 3336 3972 3344
rect 3996 3336 4004 3344
rect 4076 3336 4084 3344
rect 4188 3336 4196 3344
rect 4284 3336 4292 3344
rect 4396 3336 4404 3344
rect 5116 3336 5124 3344
rect 5164 3336 5172 3344
rect 2796 3316 2804 3324
rect 2828 3316 2836 3324
rect 2876 3316 2884 3324
rect 3084 3316 3092 3324
rect 3564 3316 3572 3324
rect 3740 3316 3748 3324
rect 3900 3316 3908 3324
rect 4316 3316 4324 3324
rect 4364 3316 4372 3324
rect 4732 3316 4740 3324
rect 4796 3316 4804 3324
rect 4908 3316 4916 3324
rect 5020 3316 5028 3324
rect 92 3296 100 3304
rect 108 3296 116 3304
rect 348 3296 356 3304
rect 364 3296 372 3304
rect 396 3296 404 3304
rect 1068 3296 1076 3304
rect 1132 3296 1140 3304
rect 2620 3296 2628 3304
rect 3804 3296 3812 3304
rect 3980 3296 3988 3304
rect 5180 3296 5188 3304
rect 284 3276 292 3284
rect 1372 3276 1380 3284
rect 1596 3276 1604 3284
rect 1660 3276 1668 3284
rect 1692 3276 1700 3284
rect 2108 3276 2116 3284
rect 2492 3276 2500 3284
rect 5052 3276 5060 3284
rect 844 3256 852 3264
rect 1564 3256 1572 3264
rect 2044 3256 2052 3264
rect 2124 3256 2132 3264
rect 2988 3256 2996 3264
rect 3484 3256 3492 3264
rect 780 3236 788 3244
rect 4604 3236 4612 3244
rect 4636 3236 4644 3244
rect 4876 3236 4884 3244
rect 332 3216 340 3224
rect 1868 3216 1876 3224
rect 1980 3216 1988 3224
rect 2508 3216 2516 3224
rect 460 3196 468 3204
rect 3116 3196 3124 3204
rect 3132 3196 3140 3204
rect 3772 3196 3780 3204
rect 4732 3196 4740 3204
rect 2076 3176 2084 3184
rect 3836 3176 3844 3184
rect 3852 3176 3860 3184
rect 4556 3176 4564 3184
rect 956 3156 964 3164
rect 2316 3156 2324 3164
rect 2924 3156 2932 3164
rect 1084 3136 1092 3144
rect 1308 3136 1316 3144
rect 3020 3136 3028 3144
rect 3452 3136 3460 3144
rect 4316 3136 4324 3144
rect 4364 3136 4372 3144
rect 4764 3136 4772 3144
rect 1388 3116 1396 3124
rect 1484 3116 1492 3124
rect 1660 3116 1668 3124
rect 3580 3116 3588 3124
rect 3740 3116 3748 3124
rect 4044 3116 4052 3124
rect 4300 3116 4308 3124
rect 12 3096 20 3104
rect 156 3096 164 3104
rect 172 3096 180 3104
rect 316 3096 324 3104
rect 364 3096 372 3104
rect 396 3096 404 3104
rect 764 3096 772 3104
rect 780 3096 788 3104
rect 876 3096 884 3104
rect 908 3096 916 3104
rect 1100 3096 1108 3104
rect 1148 3096 1156 3104
rect 1196 3096 1204 3104
rect 1964 3096 1972 3104
rect 2012 3096 2020 3104
rect 2028 3096 2036 3104
rect 2332 3096 2340 3104
rect 2412 3096 2420 3104
rect 2636 3096 2644 3104
rect 3356 3096 3364 3104
rect 3388 3096 3396 3104
rect 4060 3096 4068 3104
rect 4076 3096 4084 3104
rect 4140 3096 4148 3104
rect 4396 3096 4404 3104
rect 4444 3096 4452 3104
rect 4508 3096 4516 3104
rect 4636 3096 4644 3104
rect 4940 3096 4948 3104
rect 268 3076 276 3084
rect 588 3076 596 3084
rect 940 3076 948 3084
rect 1196 3076 1204 3084
rect 1260 3076 1268 3084
rect 2716 3076 2724 3084
rect 2748 3076 2756 3084
rect 2764 3076 2772 3084
rect 2956 3076 2964 3084
rect 3356 3076 3364 3084
rect 828 3056 836 3064
rect 1644 3056 1652 3064
rect 3276 3056 3284 3064
rect 3340 3056 3348 3064
rect 3420 3056 3428 3064
rect 3564 3056 3572 3064
rect 3996 3056 4004 3064
rect 4476 3056 4484 3064
rect 4892 3056 4900 3064
rect 4940 3056 4948 3064
rect 5084 3056 5092 3064
rect 1068 3036 1076 3044
rect 1084 3036 1092 3044
rect 2492 3036 2500 3044
rect 2588 3036 2596 3044
rect 3084 3036 3092 3044
rect 3228 3036 3236 3044
rect 3980 3036 3988 3044
rect 4172 3036 4180 3044
rect 4300 3036 4308 3044
rect 4604 3036 4612 3044
rect 540 3016 548 3024
rect 2924 3016 2932 3024
rect 3100 3016 3108 3024
rect 4172 3016 4180 3024
rect 4652 3016 4660 3024
rect 4892 3016 4900 3024
rect 940 2996 948 3004
rect 2140 2996 2148 3004
rect 2156 2996 2164 3004
rect 2908 2996 2916 3004
rect 2956 2996 2964 3004
rect 3532 2996 3540 3004
rect 3612 2996 3620 3004
rect 4572 2996 4580 3004
rect 284 2976 292 2984
rect 668 2976 676 2984
rect 1132 2976 1140 2984
rect 172 2956 180 2964
rect 316 2956 324 2964
rect 444 2956 452 2964
rect 2252 2956 2260 2964
rect 2524 2956 2532 2964
rect 2620 2956 2628 2964
rect 2668 2956 2676 2964
rect 2716 2956 2724 2964
rect 2764 2956 2772 2964
rect 2780 2956 2788 2964
rect 2844 2956 2852 2964
rect 3900 2956 3908 2964
rect 4908 2956 4916 2964
rect 5052 2956 5060 2964
rect 140 2936 148 2944
rect 252 2936 260 2944
rect 700 2936 708 2944
rect 1628 2936 1636 2944
rect 2092 2936 2100 2944
rect 2508 2936 2516 2944
rect 2572 2936 2580 2944
rect 2620 2936 2628 2944
rect 2668 2936 2676 2944
rect 3324 2936 3332 2944
rect 3708 2936 3716 2944
rect 4092 2936 4100 2944
rect 4220 2936 4228 2944
rect 4732 2936 4740 2944
rect 4764 2936 4772 2944
rect 4860 2936 4868 2944
rect 236 2916 244 2924
rect 540 2916 548 2924
rect 700 2916 708 2924
rect 812 2916 820 2924
rect 2204 2916 2212 2924
rect 2284 2916 2292 2924
rect 3148 2916 3156 2924
rect 3532 2916 3540 2924
rect 3692 2916 3700 2924
rect 3708 2916 3716 2924
rect 4252 2916 4260 2924
rect 4348 2916 4356 2924
rect 4364 2916 4372 2924
rect 4556 2916 4564 2924
rect 5084 2916 5092 2924
rect 476 2896 484 2904
rect 668 2896 676 2904
rect 796 2896 804 2904
rect 860 2896 868 2904
rect 1132 2896 1140 2904
rect 1452 2896 1460 2904
rect 1580 2896 1588 2904
rect 1596 2896 1604 2904
rect 1644 2896 1652 2904
rect 1868 2896 1876 2904
rect 2316 2896 2324 2904
rect 3148 2896 3156 2904
rect 3228 2896 3236 2904
rect 3324 2896 3332 2904
rect 3372 2896 3380 2904
rect 4124 2896 4132 2904
rect 4156 2896 4164 2904
rect 4300 2896 4308 2904
rect 4732 2896 4740 2904
rect 5132 2896 5140 2904
rect 1340 2876 1348 2884
rect 1404 2876 1412 2884
rect 1532 2876 1540 2884
rect 1628 2876 1636 2884
rect 1772 2876 1780 2884
rect 1804 2876 1812 2884
rect 1916 2876 1924 2884
rect 1996 2876 2004 2884
rect 2060 2876 2068 2884
rect 2428 2876 2436 2884
rect 3004 2876 3012 2884
rect 4444 2876 4452 2884
rect 4652 2876 4660 2884
rect 716 2856 724 2864
rect 780 2856 788 2864
rect 1276 2856 1284 2864
rect 1628 2856 1636 2864
rect 1756 2856 1764 2864
rect 1900 2856 1908 2864
rect 1180 2836 1188 2844
rect 2684 2836 2692 2844
rect 2828 2836 2836 2844
rect 1612 2816 1620 2824
rect 2764 2816 2772 2824
rect 4668 2816 4676 2824
rect 3036 2796 3044 2804
rect 5180 2796 5188 2804
rect 812 2776 820 2784
rect 1836 2776 1844 2784
rect 3276 2776 3284 2784
rect 4156 2756 4164 2764
rect 4188 2756 4196 2764
rect 1788 2736 1796 2744
rect 2092 2736 2100 2744
rect 2188 2736 2196 2744
rect 2316 2736 2324 2744
rect 2940 2736 2948 2744
rect 2956 2736 2964 2744
rect 3020 2736 3028 2744
rect 4764 2736 4772 2744
rect 4908 2736 4916 2744
rect 5148 2736 5156 2744
rect 12 2716 20 2724
rect 236 2716 244 2724
rect 908 2716 916 2724
rect 988 2716 996 2724
rect 1084 2716 1092 2724
rect 1292 2716 1300 2724
rect 1356 2716 1364 2724
rect 2508 2716 2516 2724
rect 3100 2716 3108 2724
rect 3212 2716 3220 2724
rect 3308 2716 3316 2724
rect 3356 2716 3364 2724
rect 3388 2716 3396 2724
rect 3436 2716 3444 2724
rect 3548 2716 3556 2724
rect 3564 2716 3572 2724
rect 3916 2716 3924 2724
rect 4060 2716 4068 2724
rect 4092 2716 4100 2724
rect 5100 2716 5108 2724
rect 1196 2696 1204 2704
rect 1500 2696 1508 2704
rect 1516 2696 1524 2704
rect 1612 2696 1620 2704
rect 3868 2696 3876 2704
rect 3884 2696 3892 2704
rect 4540 2696 4548 2704
rect 4668 2696 4676 2704
rect 4716 2696 4724 2704
rect 4908 2696 4916 2704
rect 108 2676 116 2684
rect 508 2676 516 2684
rect 700 2676 708 2684
rect 812 2676 820 2684
rect 940 2676 948 2684
rect 1036 2676 1044 2684
rect 1148 2676 1156 2684
rect 1516 2676 1524 2684
rect 2380 2676 2388 2684
rect 2620 2676 2628 2684
rect 2844 2676 2852 2684
rect 2940 2676 2948 2684
rect 4156 2676 4164 2684
rect 4252 2676 4260 2684
rect 4300 2676 4308 2684
rect 4364 2676 4372 2684
rect 4380 2676 4388 2684
rect 4604 2676 4612 2684
rect 4972 2676 4980 2684
rect 5052 2676 5060 2684
rect 5084 2676 5092 2684
rect 5100 2676 5108 2684
rect 156 2656 164 2664
rect 172 2656 180 2664
rect 204 2656 212 2664
rect 300 2656 308 2664
rect 348 2656 356 2664
rect 876 2656 884 2664
rect 1148 2656 1156 2664
rect 1244 2656 1252 2664
rect 1308 2656 1316 2664
rect 2684 2656 2692 2664
rect 2908 2656 2916 2664
rect 3212 2656 3220 2664
rect 3324 2656 3332 2664
rect 3628 2656 3636 2664
rect 3660 2656 3668 2664
rect 3740 2656 3748 2664
rect 4876 2656 4884 2664
rect 5004 2656 5012 2664
rect 396 2636 404 2644
rect 572 2636 580 2644
rect 700 2636 708 2644
rect 1356 2636 1364 2644
rect 1708 2636 1716 2644
rect 1772 2636 1780 2644
rect 2044 2636 2052 2644
rect 2524 2636 2532 2644
rect 3100 2636 3108 2644
rect 3132 2636 3140 2644
rect 3660 2636 3668 2644
rect 3852 2636 3860 2644
rect 4892 2636 4900 2644
rect 4956 2636 4964 2644
rect 5100 2636 5108 2644
rect 1308 2616 1316 2624
rect 1468 2616 1476 2624
rect 1580 2616 1588 2624
rect 1628 2616 1636 2624
rect 1932 2616 1940 2624
rect 1996 2616 2004 2624
rect 2188 2616 2196 2624
rect 2428 2616 2436 2624
rect 3996 2616 4004 2624
rect 4428 2616 4436 2624
rect 4444 2616 4452 2624
rect 4460 2616 4468 2624
rect 748 2596 756 2604
rect 956 2596 964 2604
rect 1788 2596 1796 2604
rect 2236 2596 2244 2604
rect 2540 2596 2548 2604
rect 3180 2596 3188 2604
rect 4028 2596 4036 2604
rect 4140 2596 4148 2604
rect 4572 2596 4580 2604
rect 4892 2596 4900 2604
rect 140 2576 148 2584
rect 364 2576 372 2584
rect 508 2576 516 2584
rect 556 2576 564 2584
rect 764 2576 772 2584
rect 956 2576 964 2584
rect 2508 2576 2516 2584
rect 3612 2576 3620 2584
rect 3644 2576 3652 2584
rect 3740 2576 3748 2584
rect 4732 2576 4740 2584
rect 2124 2556 2132 2564
rect 2316 2556 2324 2564
rect 2876 2556 2884 2564
rect 2908 2556 2916 2564
rect 2924 2556 2932 2564
rect 2940 2556 2948 2564
rect 3020 2556 3028 2564
rect 3788 2556 3796 2564
rect 4796 2556 4804 2564
rect 5084 2556 5092 2564
rect 108 2536 116 2544
rect 828 2536 836 2544
rect 924 2536 932 2544
rect 1164 2536 1172 2544
rect 1196 2536 1204 2544
rect 1276 2536 1284 2544
rect 1308 2536 1316 2544
rect 1340 2536 1348 2544
rect 1436 2536 1444 2544
rect 2364 2536 2372 2544
rect 2444 2536 2452 2544
rect 2636 2536 2644 2544
rect 2668 2536 2676 2544
rect 4204 2536 4212 2544
rect 156 2516 164 2524
rect 748 2516 756 2524
rect 780 2516 788 2524
rect 828 2516 836 2524
rect 1212 2516 1220 2524
rect 1308 2516 1316 2524
rect 3484 2516 3492 2524
rect 3532 2516 3540 2524
rect 3548 2516 3556 2524
rect 3628 2516 3636 2524
rect 3660 2516 3668 2524
rect 3948 2516 3956 2524
rect 4156 2516 4164 2524
rect 4236 2516 4244 2524
rect 4524 2516 4532 2524
rect 4588 2516 4596 2524
rect 5036 2516 5044 2524
rect 444 2496 452 2504
rect 508 2496 516 2504
rect 1020 2496 1028 2504
rect 1036 2496 1044 2504
rect 1068 2496 1076 2504
rect 1388 2496 1396 2504
rect 1628 2496 1636 2504
rect 1708 2496 1716 2504
rect 1900 2496 1908 2504
rect 1916 2496 1924 2504
rect 1980 2496 1988 2504
rect 1996 2496 2004 2504
rect 2124 2496 2132 2504
rect 2188 2496 2196 2504
rect 2668 2496 2676 2504
rect 2748 2496 2756 2504
rect 3180 2496 3188 2504
rect 3196 2496 3204 2504
rect 3404 2496 3412 2504
rect 3468 2496 3476 2504
rect 4012 2496 4020 2504
rect 4236 2496 4244 2504
rect 4476 2496 4484 2504
rect 4508 2496 4516 2504
rect 4700 2496 4708 2504
rect 4748 2496 4756 2504
rect 4796 2496 4804 2504
rect 4876 2496 4884 2504
rect 828 2476 836 2484
rect 860 2476 868 2484
rect 876 2476 884 2484
rect 1692 2476 1700 2484
rect 2540 2476 2548 2484
rect 2860 2476 2868 2484
rect 2876 2476 2884 2484
rect 3052 2476 3060 2484
rect 3100 2476 3108 2484
rect 3772 2476 3780 2484
rect 3868 2476 3876 2484
rect 3884 2476 3892 2484
rect 4140 2476 4148 2484
rect 4396 2476 4404 2484
rect 4556 2476 4564 2484
rect 4812 2476 4820 2484
rect 2428 2456 2436 2464
rect 2428 2436 2436 2444
rect 2604 2436 2612 2444
rect 4828 2436 4836 2444
rect 972 2416 980 2424
rect 2604 2416 2612 2424
rect 4012 2416 4020 2424
rect 4332 2416 4340 2424
rect 92 2396 100 2404
rect 588 2396 596 2404
rect 2428 2396 2436 2404
rect 364 2376 372 2384
rect 4060 2376 4068 2384
rect 2316 2356 2324 2364
rect 3932 2356 3940 2364
rect 4700 2356 4708 2364
rect 572 2336 580 2344
rect 604 2336 612 2344
rect 620 2336 628 2344
rect 764 2336 772 2344
rect 1500 2336 1508 2344
rect 1532 2336 1540 2344
rect 1548 2336 1556 2344
rect 2412 2336 2420 2344
rect 2684 2336 2692 2344
rect 3100 2336 3108 2344
rect 3500 2336 3508 2344
rect 3580 2336 3588 2344
rect 3996 2336 4004 2344
rect 4316 2336 4324 2344
rect 4428 2336 4436 2344
rect 4732 2336 4740 2344
rect 1036 2316 1044 2324
rect 1228 2316 1236 2324
rect 1580 2316 1588 2324
rect 1628 2316 1636 2324
rect 1836 2316 1844 2324
rect 1916 2316 1924 2324
rect 2060 2316 2068 2324
rect 2972 2316 2980 2324
rect 3020 2316 3028 2324
rect 3628 2316 3636 2324
rect 3660 2316 3668 2324
rect 3916 2316 3924 2324
rect 4124 2316 4132 2324
rect 4796 2316 4804 2324
rect 5180 2316 5188 2324
rect 428 2296 436 2304
rect 508 2296 516 2304
rect 572 2296 580 2304
rect 780 2296 788 2304
rect 908 2296 916 2304
rect 1052 2296 1060 2304
rect 1212 2296 1220 2304
rect 1404 2296 1412 2304
rect 1532 2296 1540 2304
rect 1596 2296 1604 2304
rect 1756 2296 1764 2304
rect 2076 2296 2084 2304
rect 2236 2296 2244 2304
rect 2476 2296 2484 2304
rect 2780 2296 2788 2304
rect 3020 2296 3028 2304
rect 3148 2296 3156 2304
rect 3228 2296 3236 2304
rect 3548 2296 3556 2304
rect 4844 2296 4852 2304
rect 5052 2296 5060 2304
rect 796 2276 804 2284
rect 924 2276 932 2284
rect 988 2276 996 2284
rect 1244 2276 1252 2284
rect 1308 2276 1316 2284
rect 1996 2276 2004 2284
rect 2396 2276 2404 2284
rect 2412 2276 2420 2284
rect 2604 2276 2612 2284
rect 2764 2276 2772 2284
rect 2988 2276 2996 2284
rect 3740 2276 3748 2284
rect 3772 2276 3780 2284
rect 3836 2276 3844 2284
rect 3932 2276 3940 2284
rect 4156 2276 4164 2284
rect 4220 2276 4228 2284
rect 4268 2276 4276 2284
rect 4412 2276 4420 2284
rect 4428 2276 4436 2284
rect 4588 2276 4596 2284
rect 4732 2276 4740 2284
rect 4828 2276 4836 2284
rect 4892 2276 4900 2284
rect 5084 2276 5092 2284
rect 28 2256 36 2264
rect 60 2256 68 2264
rect 172 2256 180 2264
rect 188 2256 196 2264
rect 220 2256 228 2264
rect 300 2256 308 2264
rect 332 2256 340 2264
rect 348 2256 356 2264
rect 524 2256 532 2264
rect 540 2256 548 2264
rect 668 2256 676 2264
rect 844 2256 852 2264
rect 1804 2256 1812 2264
rect 1852 2256 1860 2264
rect 3868 2256 3876 2264
rect 3948 2256 3956 2264
rect 3980 2256 3988 2264
rect 4268 2256 4276 2264
rect 4860 2256 4868 2264
rect 4924 2256 4932 2264
rect 332 2236 340 2244
rect 828 2236 836 2244
rect 1836 2236 1844 2244
rect 1900 2236 1908 2244
rect 2012 2236 2020 2244
rect 2028 2236 2036 2244
rect 2588 2236 2596 2244
rect 4364 2236 4372 2244
rect 4972 2236 4980 2244
rect 1852 2216 1860 2224
rect 1932 2216 1940 2224
rect 2284 2216 2292 2224
rect 2412 2216 2420 2224
rect 3020 2216 3028 2224
rect 3644 2216 3652 2224
rect 3772 2216 3780 2224
rect 4188 2216 4196 2224
rect 4396 2216 4404 2224
rect 1388 2196 1396 2204
rect 2188 2196 2196 2204
rect 2556 2196 2564 2204
rect 2908 2196 2916 2204
rect 348 2176 356 2184
rect 684 2176 692 2184
rect 700 2176 708 2184
rect 716 2176 724 2184
rect 3148 2176 3156 2184
rect 3356 2176 3364 2184
rect 380 2156 388 2164
rect 460 2156 468 2164
rect 796 2156 804 2164
rect 1292 2156 1300 2164
rect 1324 2156 1332 2164
rect 1628 2156 1636 2164
rect 1660 2156 1668 2164
rect 1692 2156 1700 2164
rect 3356 2156 3364 2164
rect 3708 2156 3716 2164
rect 4108 2156 4116 2164
rect 4124 2156 4132 2164
rect 4236 2156 4244 2164
rect 4300 2156 4308 2164
rect 4700 2156 4708 2164
rect 4748 2156 4756 2164
rect 5100 2156 5108 2164
rect 12 2136 20 2144
rect 316 2136 324 2144
rect 1308 2136 1316 2144
rect 2204 2136 2212 2144
rect 3228 2136 3236 2144
rect 4748 2136 4756 2144
rect 4860 2136 4868 2144
rect 92 2116 100 2124
rect 332 2116 340 2124
rect 364 2116 372 2124
rect 412 2116 420 2124
rect 444 2116 452 2124
rect 892 2116 900 2124
rect 1052 2116 1060 2124
rect 1100 2116 1108 2124
rect 2188 2116 2196 2124
rect 2524 2116 2532 2124
rect 2668 2116 2676 2124
rect 2812 2116 2820 2124
rect 3004 2116 3012 2124
rect 3100 2116 3108 2124
rect 3148 2116 3156 2124
rect 3596 2116 3604 2124
rect 4252 2116 4260 2124
rect 4348 2116 4356 2124
rect 4428 2116 4436 2124
rect 4444 2116 4452 2124
rect 4508 2116 4516 2124
rect 4988 2116 4996 2124
rect 5116 2116 5124 2124
rect 284 2096 292 2104
rect 476 2096 484 2104
rect 588 2096 596 2104
rect 1500 2096 1508 2104
rect 3388 2096 3396 2104
rect 4444 2096 4452 2104
rect 4700 2096 4708 2104
rect 5164 2096 5172 2104
rect 1820 2076 1828 2084
rect 1948 2076 1956 2084
rect 1980 2076 1988 2084
rect 2060 2076 2068 2084
rect 2668 2076 2676 2084
rect 4844 2076 4852 2084
rect 4892 2076 4900 2084
rect 5116 2076 5124 2084
rect 1564 2056 1572 2064
rect 3980 2056 3988 2064
rect 3996 2056 4004 2064
rect 2140 2036 2148 2044
rect 3724 2036 3732 2044
rect 3772 2036 3780 2044
rect 4060 2036 4068 2044
rect 4780 2036 4788 2044
rect 2300 2016 2308 2024
rect 2668 2016 2676 2024
rect 2684 2016 2692 2024
rect 3308 2016 3316 2024
rect 3468 2016 3476 2024
rect 844 1976 852 1984
rect 3404 1976 3412 1984
rect 3612 1976 3620 1984
rect 4444 1976 4452 1984
rect 4588 1976 4596 1984
rect 4764 1976 4772 1984
rect 5084 1976 5092 1984
rect 1228 1956 1236 1964
rect 1356 1956 1364 1964
rect 2444 1956 2452 1964
rect 2476 1956 2484 1964
rect 2684 1956 2692 1964
rect 2876 1956 2884 1964
rect 3052 1956 3060 1964
rect 4076 1956 4084 1964
rect 4556 1956 4564 1964
rect 2220 1936 2228 1944
rect 556 1916 564 1924
rect 668 1916 676 1924
rect 684 1916 692 1924
rect 1052 1916 1060 1924
rect 1164 1916 1172 1924
rect 1212 1916 1220 1924
rect 1804 1916 1812 1924
rect 1884 1916 1892 1924
rect 2044 1916 2052 1924
rect 2588 1916 2596 1924
rect 2716 1916 2724 1924
rect 2940 1916 2948 1924
rect 2972 1916 2980 1924
rect 3996 1916 4004 1924
rect 4620 1916 4628 1924
rect 4732 1916 4740 1924
rect 188 1896 196 1904
rect 652 1896 660 1904
rect 860 1896 868 1904
rect 924 1896 932 1904
rect 988 1896 996 1904
rect 1036 1896 1044 1904
rect 1116 1896 1124 1904
rect 1500 1896 1508 1904
rect 1532 1896 1540 1904
rect 1628 1896 1636 1904
rect 1724 1896 1732 1904
rect 2108 1896 2116 1904
rect 2188 1896 2196 1904
rect 2300 1896 2308 1904
rect 2508 1896 2516 1904
rect 2748 1896 2756 1904
rect 2764 1896 2772 1904
rect 2796 1896 2804 1904
rect 2956 1896 2964 1904
rect 3052 1896 3060 1904
rect 3180 1896 3188 1904
rect 3228 1896 3236 1904
rect 3484 1896 3492 1904
rect 3628 1896 3636 1904
rect 3644 1896 3652 1904
rect 4300 1896 4308 1904
rect 4972 1896 4980 1904
rect 348 1876 356 1884
rect 684 1876 692 1884
rect 988 1876 996 1884
rect 2556 1876 2564 1884
rect 4828 1876 4836 1884
rect 300 1856 308 1864
rect 316 1856 324 1864
rect 444 1856 452 1864
rect 700 1856 708 1864
rect 796 1856 804 1864
rect 844 1856 852 1864
rect 908 1856 916 1864
rect 1244 1856 1252 1864
rect 3676 1856 3684 1864
rect 3836 1856 3844 1864
rect 4316 1856 4324 1864
rect 4940 1856 4948 1864
rect 4988 1856 4996 1864
rect 60 1836 68 1844
rect 1100 1836 1108 1844
rect 1548 1836 1556 1844
rect 3260 1836 3268 1844
rect 3468 1836 3476 1844
rect 3516 1836 3524 1844
rect 1372 1816 1380 1824
rect 1484 1816 1492 1824
rect 1500 1816 1508 1824
rect 1932 1816 1940 1824
rect 1996 1816 2004 1824
rect 2140 1816 2148 1824
rect 2700 1816 2708 1824
rect 2732 1816 2740 1824
rect 3020 1816 3028 1824
rect 748 1796 756 1804
rect 1036 1796 1044 1804
rect 2604 1796 2612 1804
rect 2972 1796 2980 1804
rect 3324 1796 3332 1804
rect 3340 1796 3348 1804
rect 4348 1796 4356 1804
rect 220 1776 228 1784
rect 524 1776 532 1784
rect 892 1776 900 1784
rect 924 1776 932 1784
rect 1004 1776 1012 1784
rect 1644 1776 1652 1784
rect 2380 1776 2388 1784
rect 2396 1776 2404 1784
rect 3004 1776 3012 1784
rect 3084 1776 3092 1784
rect 3500 1776 3508 1784
rect 3756 1776 3764 1784
rect 4492 1776 4500 1784
rect 4684 1776 4692 1784
rect 5100 1776 5108 1784
rect 140 1756 148 1764
rect 844 1756 852 1764
rect 1676 1756 1684 1764
rect 1692 1756 1700 1764
rect 1740 1756 1748 1764
rect 1756 1756 1764 1764
rect 1884 1756 1892 1764
rect 1964 1756 1972 1764
rect 2140 1756 2148 1764
rect 2172 1756 2180 1764
rect 2284 1756 2292 1764
rect 3452 1756 3460 1764
rect 3484 1756 3492 1764
rect 3580 1756 3588 1764
rect 3628 1756 3636 1764
rect 4076 1756 4084 1764
rect 4124 1756 4132 1764
rect 5020 1756 5028 1764
rect 5116 1756 5124 1764
rect 252 1736 260 1744
rect 492 1736 500 1744
rect 1500 1736 1508 1744
rect 1740 1736 1748 1744
rect 1756 1736 1764 1744
rect 1868 1736 1876 1744
rect 1916 1736 1924 1744
rect 2028 1736 2036 1744
rect 2092 1736 2100 1744
rect 2108 1736 2116 1744
rect 2588 1736 2596 1744
rect 3068 1736 3076 1744
rect 3180 1736 3188 1744
rect 3660 1736 3668 1744
rect 3836 1736 3844 1744
rect 3980 1736 3988 1744
rect 4028 1736 4036 1744
rect 4060 1736 4068 1744
rect 4172 1736 4180 1744
rect 4460 1736 4468 1744
rect 4668 1736 4676 1744
rect 4700 1736 4708 1744
rect 5020 1736 5028 1744
rect 60 1716 68 1724
rect 668 1716 676 1724
rect 796 1716 804 1724
rect 1356 1716 1364 1724
rect 1996 1716 2004 1724
rect 2540 1716 2548 1724
rect 2588 1716 2596 1724
rect 2684 1716 2692 1724
rect 3004 1716 3012 1724
rect 3164 1716 3172 1724
rect 3692 1716 3700 1724
rect 3740 1716 3748 1724
rect 4348 1716 4356 1724
rect 4652 1716 4660 1724
rect 5068 1716 5076 1724
rect 5084 1716 5092 1724
rect 284 1696 292 1704
rect 572 1696 580 1704
rect 700 1696 708 1704
rect 844 1696 852 1704
rect 1116 1696 1124 1704
rect 1164 1696 1172 1704
rect 1228 1696 1236 1704
rect 1436 1696 1444 1704
rect 1788 1696 1796 1704
rect 1836 1696 1844 1704
rect 2380 1696 2388 1704
rect 2988 1696 2996 1704
rect 3020 1696 3028 1704
rect 3052 1696 3060 1704
rect 3212 1696 3220 1704
rect 3228 1696 3236 1704
rect 3324 1696 3332 1704
rect 3436 1696 3444 1704
rect 3916 1696 3924 1704
rect 3980 1696 3988 1704
rect 4220 1696 4228 1704
rect 4492 1696 4500 1704
rect 5020 1696 5028 1704
rect 5164 1696 5172 1704
rect 4380 1676 4388 1684
rect 2236 1656 2244 1664
rect 3996 1656 4004 1664
rect 4956 1656 4964 1664
rect 5004 1656 5012 1664
rect 860 1636 868 1644
rect 956 1636 964 1644
rect 1644 1636 1652 1644
rect 1676 1636 1684 1644
rect 3084 1636 3092 1644
rect 4044 1636 4052 1644
rect 4188 1636 4196 1644
rect 4284 1636 4292 1644
rect 2284 1616 2292 1624
rect 3388 1616 3396 1624
rect 3516 1616 3524 1624
rect 684 1596 692 1604
rect 2748 1596 2756 1604
rect 3484 1596 3492 1604
rect 4140 1596 4148 1604
rect 4188 1596 4196 1604
rect 4764 1596 4772 1604
rect 444 1576 452 1584
rect 2748 1576 2756 1584
rect 2924 1576 2932 1584
rect 3148 1576 3156 1584
rect 4764 1576 4772 1584
rect 4812 1576 4820 1584
rect 4828 1576 4836 1584
rect 1244 1556 1252 1564
rect 2188 1556 2196 1564
rect 2444 1556 2452 1564
rect 1212 1536 1220 1544
rect 1788 1536 1796 1544
rect 2316 1536 2324 1544
rect 3132 1536 3140 1544
rect 3340 1536 3348 1544
rect 3356 1536 3364 1544
rect 3500 1536 3508 1544
rect 3660 1536 3668 1544
rect 4268 1536 4276 1544
rect 4316 1536 4324 1544
rect 4396 1536 4404 1544
rect 4476 1536 4484 1544
rect 4876 1536 4884 1544
rect 92 1516 100 1524
rect 108 1516 116 1524
rect 332 1516 340 1524
rect 588 1516 596 1524
rect 1196 1516 1204 1524
rect 1708 1516 1716 1524
rect 2300 1516 2308 1524
rect 2332 1516 2340 1524
rect 3340 1516 3348 1524
rect 3404 1516 3412 1524
rect 3484 1516 3492 1524
rect 3932 1516 3940 1524
rect 4012 1516 4020 1524
rect 5036 1516 5044 1524
rect 5116 1516 5124 1524
rect 860 1496 868 1504
rect 908 1496 916 1504
rect 1660 1496 1668 1504
rect 1740 1496 1748 1504
rect 1964 1496 1972 1504
rect 2060 1496 2068 1504
rect 2508 1496 2516 1504
rect 2556 1496 2564 1504
rect 2780 1496 2788 1504
rect 3020 1496 3028 1504
rect 4188 1496 4196 1504
rect 4540 1496 4548 1504
rect 5132 1496 5140 1504
rect 12 1476 20 1484
rect 204 1476 212 1484
rect 1756 1476 1764 1484
rect 1804 1476 1812 1484
rect 1868 1476 1876 1484
rect 2028 1476 2036 1484
rect 2092 1476 2100 1484
rect 2236 1476 2244 1484
rect 4156 1476 4164 1484
rect 4604 1476 4612 1484
rect 4652 1476 4660 1484
rect 4828 1476 4836 1484
rect 4988 1476 4996 1484
rect 156 1456 164 1464
rect 220 1456 228 1464
rect 348 1456 356 1464
rect 380 1456 388 1464
rect 876 1456 884 1464
rect 1372 1456 1380 1464
rect 1612 1456 1620 1464
rect 2188 1456 2196 1464
rect 2332 1456 2340 1464
rect 3628 1456 3636 1464
rect 4220 1456 4228 1464
rect 4236 1456 4244 1464
rect 4700 1456 4708 1464
rect 4716 1456 4724 1464
rect 4956 1456 4964 1464
rect 5148 1456 5156 1464
rect 940 1436 948 1444
rect 2396 1436 2404 1444
rect 3452 1436 3460 1444
rect 4876 1436 4884 1444
rect 1228 1416 1236 1424
rect 2140 1416 2148 1424
rect 2652 1416 2660 1424
rect 2892 1416 2900 1424
rect 3212 1416 3220 1424
rect 4252 1416 4260 1424
rect 4524 1416 4532 1424
rect 4668 1416 4676 1424
rect 4876 1416 4884 1424
rect 1244 1396 1252 1404
rect 1404 1396 1412 1404
rect 1516 1396 1524 1404
rect 1628 1396 1636 1404
rect 1676 1396 1684 1404
rect 1692 1396 1700 1404
rect 1836 1396 1844 1404
rect 1852 1396 1860 1404
rect 2412 1396 2420 1404
rect 12 1376 20 1384
rect 380 1376 388 1384
rect 1548 1376 1556 1384
rect 1580 1376 1588 1384
rect 2572 1376 2580 1384
rect 2604 1376 2612 1384
rect 3660 1376 3668 1384
rect 3740 1376 3748 1384
rect 524 1356 532 1364
rect 636 1356 644 1364
rect 876 1356 884 1364
rect 972 1356 980 1364
rect 1900 1356 1908 1364
rect 2044 1356 2052 1364
rect 2332 1356 2340 1364
rect 2364 1356 2372 1364
rect 2668 1356 2676 1364
rect 2876 1356 2884 1364
rect 2908 1356 2916 1364
rect 3356 1356 3364 1364
rect 3724 1356 3732 1364
rect 3884 1356 3892 1364
rect 3932 1356 3940 1364
rect 4268 1356 4276 1364
rect 4300 1356 4308 1364
rect 4364 1356 4372 1364
rect 4444 1356 4452 1364
rect 4604 1356 4612 1364
rect 4828 1356 4836 1364
rect 4972 1356 4980 1364
rect 76 1336 84 1344
rect 428 1336 436 1344
rect 732 1336 740 1344
rect 972 1336 980 1344
rect 1244 1336 1252 1344
rect 1292 1336 1300 1344
rect 2396 1336 2404 1344
rect 2412 1336 2420 1344
rect 2492 1336 2500 1344
rect 2604 1336 2612 1344
rect 2668 1336 2676 1344
rect 2764 1336 2772 1344
rect 2796 1336 2804 1344
rect 2972 1336 2980 1344
rect 2988 1336 2996 1344
rect 3228 1336 3236 1344
rect 3964 1336 3972 1344
rect 4380 1336 4388 1344
rect 5196 1336 5204 1344
rect 92 1316 100 1324
rect 156 1316 164 1324
rect 332 1316 340 1324
rect 444 1316 452 1324
rect 588 1316 596 1324
rect 668 1316 676 1324
rect 1468 1316 1476 1324
rect 1916 1316 1924 1324
rect 2268 1316 2276 1324
rect 3884 1316 3892 1324
rect 4028 1316 4036 1324
rect 4140 1316 4148 1324
rect 4860 1316 4868 1324
rect 5100 1316 5108 1324
rect 5116 1316 5124 1324
rect 284 1296 292 1304
rect 1340 1296 1348 1304
rect 1388 1296 1396 1304
rect 1484 1296 1492 1304
rect 2444 1296 2452 1304
rect 2604 1296 2612 1304
rect 2988 1296 2996 1304
rect 3004 1296 3012 1304
rect 3212 1296 3220 1304
rect 3324 1296 3332 1304
rect 3372 1296 3380 1304
rect 3388 1296 3396 1304
rect 3436 1296 3444 1304
rect 3548 1296 3556 1304
rect 3980 1296 3988 1304
rect 4572 1296 4580 1304
rect 4700 1296 4708 1304
rect 4796 1296 4804 1304
rect 4876 1296 4884 1304
rect 5068 1296 5076 1304
rect 5100 1296 5108 1304
rect 4044 1276 4052 1284
rect 4076 1276 4084 1284
rect 4300 1276 4308 1284
rect 4460 1276 4468 1284
rect 4556 1276 4564 1284
rect 4812 1276 4820 1284
rect 4876 1276 4884 1284
rect 524 1256 532 1264
rect 780 1256 788 1264
rect 1068 1256 1076 1264
rect 1132 1256 1140 1264
rect 2060 1256 2068 1264
rect 2876 1256 2884 1264
rect 4060 1256 4068 1264
rect 2396 1236 2404 1244
rect 2748 1236 2756 1244
rect 3036 1236 3044 1244
rect 3372 1236 3380 1244
rect 3516 1236 3524 1244
rect 3628 1236 3636 1244
rect 3868 1236 3876 1244
rect 4860 1236 4868 1244
rect 5004 1236 5012 1244
rect 860 1216 868 1224
rect 1948 1216 1956 1224
rect 1964 1216 1972 1224
rect 2140 1216 2148 1224
rect 2172 1216 2180 1224
rect 2300 1216 2308 1224
rect 2396 1216 2404 1224
rect 2748 1216 2756 1224
rect 2796 1216 2804 1224
rect 3708 1216 3716 1224
rect 3788 1216 3796 1224
rect 3836 1196 3844 1204
rect 700 1176 708 1184
rect 908 1176 916 1184
rect 1036 1176 1044 1184
rect 1820 1176 1828 1184
rect 3036 1176 3044 1184
rect 4540 1176 4548 1184
rect 5100 1176 5108 1184
rect 28 1156 36 1164
rect 1260 1156 1268 1164
rect 1868 1156 1876 1164
rect 3788 1156 3796 1164
rect 3980 1156 3988 1164
rect 3996 1156 4004 1164
rect 4220 1156 4228 1164
rect 4444 1156 4452 1164
rect 1260 1136 1268 1144
rect 1516 1136 1524 1144
rect 1916 1136 1924 1144
rect 3436 1136 3444 1144
rect 3628 1136 3636 1144
rect 4604 1136 4612 1144
rect 4732 1136 4740 1144
rect 5116 1136 5124 1144
rect 460 1116 468 1124
rect 476 1116 484 1124
rect 572 1116 580 1124
rect 764 1116 772 1124
rect 1116 1116 1124 1124
rect 1164 1116 1172 1124
rect 1356 1116 1364 1124
rect 1756 1116 1764 1124
rect 2108 1116 2116 1124
rect 2124 1116 2132 1124
rect 2588 1116 2596 1124
rect 2860 1116 2868 1124
rect 3212 1116 3220 1124
rect 4300 1116 4308 1124
rect 4796 1116 4804 1124
rect 620 1096 628 1104
rect 716 1096 724 1104
rect 796 1096 804 1104
rect 1740 1096 1748 1104
rect 2076 1096 2084 1104
rect 2172 1096 2180 1104
rect 2220 1096 2228 1104
rect 2236 1096 2244 1104
rect 2348 1096 2356 1104
rect 2396 1096 2404 1104
rect 2732 1096 2740 1104
rect 3084 1096 3092 1104
rect 3260 1096 3268 1104
rect 3532 1096 3540 1104
rect 3772 1096 3780 1104
rect 4012 1096 4020 1104
rect 4204 1096 4212 1104
rect 4364 1096 4372 1104
rect 4444 1096 4452 1104
rect 4508 1096 4516 1104
rect 4988 1096 4996 1104
rect 5148 1096 5156 1104
rect 76 1076 84 1084
rect 620 1076 628 1084
rect 1148 1076 1156 1084
rect 1180 1076 1188 1084
rect 1452 1076 1460 1084
rect 1676 1076 1684 1084
rect 2460 1076 2468 1084
rect 3148 1076 3156 1084
rect 4604 1076 4612 1084
rect 4636 1076 4644 1084
rect 4764 1076 4772 1084
rect 284 1056 292 1064
rect 380 1056 388 1064
rect 1388 1056 1396 1064
rect 1980 1056 1988 1064
rect 2252 1056 2260 1064
rect 2860 1056 2868 1064
rect 2956 1056 2964 1064
rect 3084 1056 3092 1064
rect 3132 1056 3140 1064
rect 3180 1056 3188 1064
rect 3612 1056 3620 1064
rect 3756 1056 3764 1064
rect 3804 1056 3812 1064
rect 5036 1056 5044 1064
rect 2700 1036 2708 1044
rect 2876 1036 2884 1044
rect 3324 1036 3332 1044
rect 3868 1036 3876 1044
rect 1148 1016 1156 1024
rect 1932 1016 1940 1024
rect 2876 1016 2884 1024
rect 3004 1016 3012 1024
rect 3484 1016 3492 1024
rect 4636 1016 4644 1024
rect 5052 1016 5060 1024
rect 1308 996 1316 1004
rect 3180 996 3188 1004
rect 4300 996 4308 1004
rect 732 976 740 984
rect 1212 976 1220 984
rect 1308 976 1316 984
rect 1500 976 1508 984
rect 1852 976 1860 984
rect 2908 976 2916 984
rect 3372 976 3380 984
rect 4332 976 4340 984
rect 4732 976 4740 984
rect 4780 976 4788 984
rect 4892 976 4900 984
rect 5132 976 5140 984
rect 5196 976 5204 984
rect 140 956 148 964
rect 364 956 372 964
rect 396 956 404 964
rect 1964 956 1972 964
rect 2684 956 2692 964
rect 2700 956 2708 964
rect 2732 956 2740 964
rect 3276 956 3284 964
rect 3340 956 3348 964
rect 3484 956 3492 964
rect 3628 956 3636 964
rect 3772 956 3780 964
rect 3804 956 3812 964
rect 3868 956 3876 964
rect 4108 956 4116 964
rect 4140 956 4148 964
rect 4956 956 4964 964
rect 5020 956 5028 964
rect 5148 956 5156 964
rect 300 936 308 944
rect 316 936 324 944
rect 348 936 356 944
rect 1196 936 1204 944
rect 1244 936 1252 944
rect 1276 936 1284 944
rect 1484 936 1492 944
rect 1996 936 2004 944
rect 2076 936 2084 944
rect 2124 936 2132 944
rect 2492 936 2500 944
rect 2572 936 2580 944
rect 2716 936 2724 944
rect 2940 936 2948 944
rect 2956 936 2964 944
rect 3164 936 3172 944
rect 3372 936 3380 944
rect 3436 936 3444 944
rect 3564 936 3572 944
rect 4076 936 4084 944
rect 4236 936 4244 944
rect 4460 936 4468 944
rect 4524 936 4532 944
rect 4604 936 4612 944
rect 4700 936 4708 944
rect 716 916 724 924
rect 764 916 772 924
rect 1692 916 1700 924
rect 2748 916 2756 924
rect 3916 916 3924 924
rect 3980 916 3988 924
rect 4604 916 4612 924
rect 5164 916 5172 924
rect 108 896 116 904
rect 956 896 964 904
rect 1468 896 1476 904
rect 1980 896 1988 904
rect 2092 896 2100 904
rect 2188 896 2196 904
rect 2252 896 2260 904
rect 2988 896 2996 904
rect 3068 896 3076 904
rect 3180 896 3188 904
rect 3212 896 3220 904
rect 3756 896 3764 904
rect 3804 896 3812 904
rect 3948 896 3956 904
rect 5004 896 5012 904
rect 5068 896 5076 904
rect 5180 896 5188 904
rect 5196 896 5204 904
rect 828 876 836 884
rect 876 876 884 884
rect 1228 876 1236 884
rect 1388 876 1396 884
rect 1804 876 1812 884
rect 1884 876 1892 884
rect 1932 876 1940 884
rect 2892 876 2900 884
rect 3308 876 3316 884
rect 4604 876 4612 884
rect 5020 876 5028 884
rect 764 856 772 864
rect 1404 856 1412 864
rect 3724 856 3732 864
rect 3884 856 3892 864
rect 1708 836 1716 844
rect 4300 836 4308 844
rect 1420 816 1428 824
rect 3020 816 3028 824
rect 3036 816 3044 824
rect 4700 816 4708 824
rect 5052 816 5060 824
rect 1740 796 1748 804
rect 1916 796 1924 804
rect 3564 776 3572 784
rect 3660 776 3668 784
rect 4812 776 4820 784
rect 1116 756 1124 764
rect 1500 756 1508 764
rect 3196 756 3204 764
rect 3436 756 3444 764
rect 4044 756 4052 764
rect 4652 756 4660 764
rect 4892 756 4900 764
rect 540 736 548 744
rect 764 736 772 744
rect 812 736 820 744
rect 1084 736 1092 744
rect 1324 736 1332 744
rect 1788 736 1796 744
rect 2428 736 2436 744
rect 2476 736 2484 744
rect 2508 736 2516 744
rect 2556 736 2564 744
rect 4012 736 4020 744
rect 4220 736 4228 744
rect 4396 736 4404 744
rect 4492 736 4500 744
rect 4732 736 4740 744
rect 4796 736 4804 744
rect 4828 736 4836 744
rect 4876 736 4884 744
rect 4956 736 4964 744
rect 604 716 612 724
rect 1628 716 1636 724
rect 2028 716 2036 724
rect 2412 716 2420 724
rect 2716 716 2724 724
rect 3052 716 3060 724
rect 3964 716 3972 724
rect 4060 716 4068 724
rect 4076 716 4084 724
rect 4156 716 4164 724
rect 860 696 868 704
rect 1084 696 1092 704
rect 1148 696 1156 704
rect 1356 696 1364 704
rect 2764 696 2772 704
rect 3180 696 3188 704
rect 3708 696 3716 704
rect 3724 696 3732 704
rect 3740 696 3748 704
rect 5084 696 5092 704
rect 220 676 228 684
rect 332 676 340 684
rect 1452 676 1460 684
rect 2268 676 2276 684
rect 2332 676 2340 684
rect 2412 676 2420 684
rect 2860 676 2868 684
rect 2956 676 2964 684
rect 3052 676 3060 684
rect 3564 676 3572 684
rect 4636 676 4644 684
rect 60 656 68 664
rect 332 656 340 664
rect 1196 656 1204 664
rect 1212 656 1220 664
rect 2812 656 2820 664
rect 3132 656 3140 664
rect 4124 656 4132 664
rect 4684 656 4692 664
rect 4716 656 4724 664
rect 5004 656 5012 664
rect 5036 656 5044 664
rect 5148 656 5156 664
rect 1004 636 1012 644
rect 1324 636 1332 644
rect 1596 636 1604 644
rect 1628 636 1636 644
rect 1660 636 1668 644
rect 3228 636 3236 644
rect 4108 636 4116 644
rect 1196 616 1204 624
rect 1676 616 1684 624
rect 1836 616 1844 624
rect 1916 616 1924 624
rect 1980 616 1988 624
rect 2268 616 2276 624
rect 2316 616 2324 624
rect 2988 616 2996 624
rect 1100 596 1108 604
rect 2076 596 2084 604
rect 2156 596 2164 604
rect 2476 596 2484 604
rect 3436 596 3444 604
rect 4108 596 4116 604
rect 4220 596 4228 604
rect 4252 596 4260 604
rect 4332 596 4340 604
rect 4492 596 4500 604
rect 4924 596 4932 604
rect 764 576 772 584
rect 828 576 836 584
rect 1932 576 1940 584
rect 2476 576 2484 584
rect 2908 576 2916 584
rect 3052 576 3060 584
rect 3196 576 3204 584
rect 3340 576 3348 584
rect 3436 576 3444 584
rect 4060 576 4068 584
rect 4716 576 4724 584
rect 44 556 52 564
rect 156 556 164 564
rect 412 556 420 564
rect 572 556 580 564
rect 1068 556 1076 564
rect 1100 556 1108 564
rect 1708 556 1716 564
rect 1724 556 1732 564
rect 1788 556 1796 564
rect 1804 556 1812 564
rect 1884 556 1892 564
rect 1932 556 1940 564
rect 1948 556 1956 564
rect 1964 556 1972 564
rect 2044 556 2052 564
rect 2524 556 2532 564
rect 2684 556 2692 564
rect 2764 556 2772 564
rect 2940 556 2948 564
rect 3020 556 3028 564
rect 3260 556 3268 564
rect 3788 556 3796 564
rect 4076 556 4084 564
rect 4140 556 4148 564
rect 4588 556 4596 564
rect 5052 556 5060 564
rect 5068 556 5076 564
rect 92 536 100 544
rect 156 536 164 544
rect 172 536 180 544
rect 364 536 372 544
rect 1372 536 1380 544
rect 1580 536 1588 544
rect 1596 536 1604 544
rect 1612 536 1620 544
rect 1868 536 1876 544
rect 3660 536 3668 544
rect 3756 536 3764 544
rect 4284 536 4292 544
rect 4652 536 4660 544
rect 4796 536 4804 544
rect 492 516 500 524
rect 508 516 516 524
rect 780 516 788 524
rect 876 516 884 524
rect 892 516 900 524
rect 1036 516 1044 524
rect 1100 516 1108 524
rect 1228 516 1236 524
rect 1356 516 1364 524
rect 1372 516 1380 524
rect 1500 516 1508 524
rect 2796 516 2804 524
rect 2956 516 2964 524
rect 3084 516 3092 524
rect 3276 516 3284 524
rect 3884 516 3892 524
rect 60 496 68 504
rect 332 496 340 504
rect 588 496 596 504
rect 652 496 660 504
rect 2028 496 2036 504
rect 2092 496 2100 504
rect 2108 496 2116 504
rect 2124 496 2132 504
rect 2860 496 2868 504
rect 3932 496 3940 504
rect 3948 496 3956 504
rect 4428 496 4436 504
rect 4540 496 4548 504
rect 5084 496 5092 504
rect 316 476 324 484
rect 636 476 644 484
rect 3452 476 3460 484
rect 3692 476 3700 484
rect 3724 476 3732 484
rect 4684 476 4692 484
rect 4716 476 4724 484
rect 748 456 756 464
rect 1644 456 1652 464
rect 1660 456 1668 464
rect 1692 456 1700 464
rect 2316 456 2324 464
rect 2460 456 2468 464
rect 2636 456 2644 464
rect 4492 456 4500 464
rect 1868 436 1876 444
rect 2044 436 2052 444
rect 3292 436 3300 444
rect 4188 436 4196 444
rect 5164 416 5172 424
rect 2716 396 2724 404
rect 1836 376 1844 384
rect 2380 376 2388 384
rect 3180 376 3188 384
rect 3580 376 3588 384
rect 3852 376 3860 384
rect 4332 376 4340 384
rect 828 356 836 364
rect 1132 356 1140 364
rect 3116 356 3124 364
rect 540 336 548 344
rect 604 336 612 344
rect 668 336 676 344
rect 1244 336 1252 344
rect 2140 336 2148 344
rect 4316 336 4324 344
rect 4604 336 4612 344
rect 4636 336 4644 344
rect 4668 336 4676 344
rect 5020 336 5028 344
rect 12 316 20 324
rect 44 316 52 324
rect 268 316 276 324
rect 428 316 436 324
rect 460 316 468 324
rect 812 316 820 324
rect 860 316 868 324
rect 940 316 948 324
rect 1036 316 1044 324
rect 1068 316 1076 324
rect 1100 316 1108 324
rect 1340 316 1348 324
rect 1916 316 1924 324
rect 2188 316 2196 324
rect 2204 316 2212 324
rect 2572 316 2580 324
rect 2604 316 2612 324
rect 2636 316 2644 324
rect 2668 316 2676 324
rect 2716 316 2724 324
rect 2940 316 2948 324
rect 3004 316 3012 324
rect 3500 316 3508 324
rect 3692 316 3700 324
rect 3836 316 3844 324
rect 3964 316 3972 324
rect 4076 316 4084 324
rect 4412 316 4420 324
rect 5100 316 5108 324
rect 92 296 100 304
rect 172 296 180 304
rect 332 296 340 304
rect 364 296 372 304
rect 3100 296 3108 304
rect 3548 296 3556 304
rect 3612 296 3620 304
rect 3660 296 3668 304
rect 3868 296 3876 304
rect 3980 296 3988 304
rect 4332 296 4340 304
rect 4508 296 4516 304
rect 4748 296 4756 304
rect 5004 296 5012 304
rect 44 276 52 284
rect 236 276 244 284
rect 1356 276 1364 284
rect 1436 276 1444 284
rect 1468 276 1476 284
rect 2108 276 2116 284
rect 2380 276 2388 284
rect 2588 276 2596 284
rect 2860 276 2868 284
rect 3260 276 3268 284
rect 4172 276 4180 284
rect 4380 276 4388 284
rect 4412 276 4420 284
rect 4524 276 4532 284
rect 4556 276 4564 284
rect 5020 276 5028 284
rect 5052 276 5060 284
rect 188 256 196 264
rect 332 256 340 264
rect 844 256 852 264
rect 2252 256 2260 264
rect 2540 256 2548 264
rect 2604 256 2612 264
rect 2860 256 2868 264
rect 2892 256 2900 264
rect 3020 256 3028 264
rect 3340 256 3348 264
rect 3468 256 3476 264
rect 4300 256 4308 264
rect 4348 256 4356 264
rect 4476 256 4484 264
rect 4604 256 4612 264
rect 4844 256 4852 264
rect 284 236 292 244
rect 476 236 484 244
rect 796 236 804 244
rect 1452 236 1460 244
rect 3916 236 3924 244
rect 956 216 964 224
rect 972 216 980 224
rect 1724 216 1732 224
rect 1772 216 1780 224
rect 1804 216 1812 224
rect 2396 216 2404 224
rect 2444 216 2452 224
rect 2732 216 2740 224
rect 2892 216 2900 224
rect 2924 216 2932 224
rect 3004 216 3012 224
rect 3036 216 3044 224
rect 3692 216 3700 224
rect 3788 216 3796 224
rect 3804 216 3812 224
rect 3900 216 3908 224
rect 988 196 996 204
rect 1196 196 1204 204
rect 2476 196 2484 204
rect 2572 196 2580 204
rect 2876 196 2884 204
rect 2924 196 2932 204
rect 3276 196 3284 204
rect 4108 196 4116 204
rect 4412 196 4420 204
rect 4860 196 4868 204
rect 300 176 308 184
rect 604 176 612 184
rect 748 176 756 184
rect 972 176 980 184
rect 1196 176 1204 184
rect 1260 176 1268 184
rect 1612 176 1620 184
rect 1772 176 1780 184
rect 2412 176 2420 184
rect 3356 176 3364 184
rect 3596 176 3604 184
rect 4140 176 4148 184
rect 268 156 276 164
rect 428 156 436 164
rect 556 156 564 164
rect 1052 156 1060 164
rect 1084 156 1092 164
rect 1212 156 1220 164
rect 1228 156 1236 164
rect 1340 156 1348 164
rect 1564 156 1572 164
rect 2204 156 2212 164
rect 2652 156 2660 164
rect 2780 156 2788 164
rect 3740 156 3748 164
rect 3868 156 3876 164
rect 4764 156 4772 164
rect 4844 156 4852 164
rect 124 136 132 144
rect 188 136 196 144
rect 1452 136 1460 144
rect 1548 136 1556 144
rect 1868 136 1876 144
rect 3420 136 3428 144
rect 3900 136 3908 144
rect 4700 136 4708 144
rect 4908 136 4916 144
rect 188 116 196 124
rect 220 116 228 124
rect 1660 116 1668 124
rect 2556 116 2564 124
rect 2732 116 2740 124
rect 3900 116 3908 124
rect 4044 116 4052 124
rect 4076 116 4084 124
rect 4652 116 4660 124
rect 4732 116 4740 124
rect 4892 116 4900 124
rect 5148 116 5156 124
rect 220 96 228 104
rect 380 96 388 104
rect 1452 96 1460 104
rect 1564 96 1572 104
rect 1804 96 1812 104
rect 2204 96 2212 104
rect 3532 96 3540 104
rect 3596 96 3604 104
rect 3644 96 3652 104
rect 4476 96 4484 104
rect 4508 96 4516 104
rect 4556 96 4564 104
rect 4588 96 4596 104
rect 476 76 484 84
rect 780 76 788 84
rect 812 76 820 84
rect 2540 76 2548 84
rect 2908 76 2916 84
rect 3196 76 3204 84
rect 3260 76 3268 84
rect 3772 76 3780 84
rect 4028 76 4036 84
rect 3148 56 3156 64
<< metal1 >>
rect -408 3616 -308 3684
rect -408 3604 8 3616
rect -408 3216 -308 3604
rect 2196 3576 2198 3584
rect 3165 3537 3188 3543
rect 604 3532 612 3536
rect 2524 3532 2532 3536
rect 3180 3532 3188 3537
rect 3316 3537 3332 3543
rect 3324 3532 3332 3537
rect 4172 3532 4180 3536
rect 317 3497 332 3503
rect 372 3497 403 3503
rect 653 3497 691 3503
rect 804 3497 819 3503
rect 1229 3497 1260 3503
rect 1293 3503 1299 3523
rect 1293 3497 1331 3503
rect 1501 3503 1507 3523
rect 1629 3503 1635 3523
rect 1469 3497 1507 3503
rect 1549 3497 1587 3503
rect 1597 3497 1635 3503
rect 1764 3497 1779 3503
rect 1901 3497 1916 3503
rect 1933 3497 1971 3503
rect 1981 3497 2012 3503
rect 2084 3497 2099 3503
rect 2205 3497 2220 3503
rect 2237 3497 2259 3503
rect 29 3477 44 3483
rect 189 3477 211 3483
rect 724 3477 739 3483
rect 788 3477 803 3483
rect 45 3457 76 3463
rect 244 3456 252 3464
rect 436 3457 451 3463
rect 484 3456 492 3464
rect 596 3457 627 3463
rect 797 3457 803 3477
rect 1252 3477 1267 3483
rect 1396 3477 1427 3483
rect 1661 3477 1699 3483
rect 1757 3477 1772 3483
rect 1789 3477 1820 3483
rect 2461 3483 2467 3503
rect 2829 3503 2835 3523
rect 3220 3517 3228 3523
rect 3453 3517 3468 3523
rect 3501 3517 3516 3523
rect 2589 3497 2627 3503
rect 2829 3497 2867 3503
rect 3565 3484 3571 3523
rect 3652 3517 3667 3523
rect 3677 3517 3715 3523
rect 3748 3517 3763 3523
rect 3837 3503 3843 3523
rect 4084 3517 4099 3523
rect 4173 3517 4195 3523
rect 4228 3517 4243 3523
rect 4349 3517 4380 3523
rect 5037 3504 5043 3523
rect 3837 3497 3875 3503
rect 4125 3497 4188 3503
rect 2260 3477 2275 3483
rect 2461 3477 2499 3483
rect 2637 3477 2668 3483
rect 2788 3477 2803 3483
rect 2877 3477 2892 3483
rect 2932 3477 2947 3483
rect 3021 3477 3036 3483
rect 3053 3477 3091 3483
rect 3261 3477 3276 3483
rect 3309 3477 3347 3483
rect 3412 3477 3427 3483
rect 3460 3477 3468 3483
rect 3981 3477 3987 3496
rect 4077 3477 4092 3483
rect 4125 3477 4131 3497
rect 4205 3497 4236 3503
rect 4276 3497 4291 3503
rect 4221 3477 4236 3483
rect 4285 3477 4291 3497
rect 4580 3497 4595 3503
rect 4605 3484 4611 3503
rect 4756 3497 4771 3503
rect 4909 3483 4915 3503
rect 5044 3497 5075 3503
rect 4612 3477 4643 3483
rect 4877 3477 4915 3483
rect 836 3457 867 3463
rect 877 3457 915 3463
rect 996 3457 1020 3463
rect 1636 3456 1644 3464
rect 1805 3457 1836 3463
rect 1997 3457 2028 3463
rect 2125 3457 2147 3463
rect 2285 3457 2307 3463
rect 2397 3457 2435 3463
rect 2653 3457 2684 3463
rect 4244 3456 4252 3464
rect 4541 3457 4556 3463
rect 4756 3457 4787 3463
rect 4964 3456 4972 3464
rect 170 3436 172 3444
rect 548 3436 550 3444
rect 1380 3436 1382 3444
rect 2820 3436 2822 3444
rect 2916 3436 2918 3444
rect 3002 3436 3004 3444
rect 3194 3436 3196 3444
rect 3242 3436 3244 3444
rect 3338 3436 3340 3444
rect 3396 3436 3398 3444
rect 3530 3436 3532 3444
rect 3722 3436 3724 3444
rect 4106 3436 4108 3444
rect 4164 3436 4166 3444
rect 4404 3436 4406 3444
rect 4452 3436 4454 3444
rect 5028 3436 5030 3444
rect 5124 3436 5126 3444
rect 5526 3416 5626 3740
rect 5206 3404 5626 3416
rect 1060 3376 1062 3384
rect 1754 3376 1756 3384
rect 3108 3376 3110 3384
rect 3146 3376 3148 3384
rect 3236 3376 3238 3384
rect 4164 3376 4166 3384
rect 237 3357 268 3363
rect 308 3356 316 3364
rect 1060 3357 1091 3363
rect 1101 3357 1116 3363
rect 1684 3357 1715 3363
rect 1812 3357 1843 3363
rect 1933 3357 1964 3363
rect 2061 3357 2092 3363
rect 525 3337 540 3343
rect 580 3337 611 3343
rect 669 3337 707 3343
rect 980 3337 1011 3343
rect 1261 3337 1276 3343
rect 1309 3337 1347 3343
rect 1652 3337 1667 3343
rect 1981 3337 2019 3343
rect 2109 3337 2124 3343
rect 2205 3337 2227 3343
rect 2221 3324 2227 3337
rect 2333 3343 2339 3363
rect 2333 3337 2371 3343
rect 2557 3343 2563 3363
rect 2708 3356 2716 3364
rect 3380 3356 3388 3364
rect 3604 3357 3635 3363
rect 3645 3357 3683 3363
rect 3716 3356 3724 3364
rect 3885 3357 3923 3363
rect 4349 3357 4364 3363
rect 4516 3357 4531 3363
rect 4541 3357 4556 3363
rect 4788 3357 4803 3363
rect 2388 3337 2419 3343
rect 2429 3337 2467 3343
rect 2557 3337 2572 3343
rect 45 3317 83 3323
rect 413 3317 428 3323
rect 509 3317 547 3323
rect 557 3317 595 3323
rect 724 3317 755 3323
rect 829 3317 860 3323
rect 900 3317 915 3323
rect 1357 3317 1372 3323
rect 1460 3317 1491 3323
rect 1549 3317 1564 3323
rect 1645 3317 1660 3323
rect 1988 3317 2003 3323
rect 2116 3317 2131 3323
rect 2253 3317 2268 3323
rect 2381 3317 2396 3323
rect 2429 3317 2435 3337
rect 2589 3337 2620 3343
rect 2781 3337 2819 3343
rect 2884 3337 2915 3343
rect 2957 3337 2995 3343
rect 3181 3337 3219 3343
rect 3492 3337 3507 3343
rect 3572 3337 3587 3343
rect 3837 3337 3852 3343
rect 3940 3337 3955 3343
rect 4084 3337 4147 3343
rect 4196 3337 4211 3343
rect 4404 3337 4435 3343
rect 2836 3317 2867 3323
rect 3021 3317 3059 3323
rect 3293 3317 3331 3323
rect 1268 3297 1283 3303
rect 3021 3297 3027 3317
rect 3661 3317 3676 3323
rect 3844 3317 3859 3323
rect 4356 3317 4371 3323
rect 4589 3317 4604 3323
rect 4804 3317 4819 3323
rect 1692 3284 1700 3288
rect 1437 3277 1452 3283
rect 1948 3284 1956 3288
rect 2076 3284 2084 3288
rect 2172 3284 2180 3288
rect 2700 3283 2708 3288
rect 2685 3277 2708 3283
rect 2972 3283 2980 3288
rect 3116 3284 3124 3288
rect 2972 3277 2988 3283
rect 3708 3283 3716 3288
rect 4892 3284 4900 3288
rect 3693 3277 3716 3283
rect 5060 3277 5075 3283
rect 3770 3236 3772 3244
rect -408 3204 4 3216
rect -408 2816 -308 3204
rect 794 3176 796 3184
rect 522 3156 524 3164
rect 2932 3156 2934 3164
rect 1508 3137 1523 3143
rect 2628 3137 2643 3143
rect 2588 3132 2596 3136
rect 2988 3132 2996 3136
rect 3244 3132 3252 3136
rect 3596 3132 3604 3136
rect 4372 3136 4374 3144
rect 4637 3137 4660 3143
rect 3772 3132 3780 3136
rect 4652 3132 4660 3137
rect 125 3097 156 3103
rect 269 3097 291 3103
rect 381 3097 396 3103
rect 429 3097 467 3103
rect 477 3097 515 3103
rect 589 3097 604 3103
rect 637 3097 675 3103
rect 685 3097 707 3103
rect 1108 3097 1139 3103
rect 1181 3097 1219 3103
rect 1533 3103 1539 3123
rect 1533 3097 1571 3103
rect 1636 3097 1644 3103
rect 1821 3097 1836 3103
rect 1885 3097 1907 3103
rect 1949 3097 1964 3103
rect 2020 3097 2035 3103
rect 2189 3103 2195 3123
rect 2285 3117 2300 3123
rect 2573 3117 2595 3123
rect 2189 3097 2227 3103
rect 2269 3097 2284 3103
rect 2340 3097 2355 3103
rect 2893 3097 2908 3103
rect 3028 3097 3043 3103
rect 3396 3097 3404 3103
rect 3901 3097 3923 3103
rect 4157 3097 4195 3103
rect 4205 3097 4220 3103
rect 4381 3097 4396 3103
rect 4948 3097 4963 3103
rect 5028 3097 5043 3103
rect 5117 3097 5132 3103
rect 221 3077 236 3083
rect 253 3077 268 3083
rect 333 3077 364 3083
rect 596 3077 627 3083
rect 1229 3077 1244 3083
rect 1741 3077 1772 3083
rect 1997 3077 2028 3083
rect 2125 3077 2163 3083
rect 2333 3077 2371 3083
rect 2436 3077 2467 3083
rect 3021 3077 3036 3083
rect 3364 3077 3379 3083
rect 3661 3077 3692 3083
rect 3853 3077 3891 3083
rect 4093 3077 4131 3083
rect 4237 3077 4275 3083
rect 20 3057 35 3063
rect 77 3057 99 3063
rect 445 3057 460 3063
rect 740 3056 748 3064
rect 845 3057 867 3063
rect 1245 3057 1276 3063
rect 1709 3057 1724 3063
rect 1789 3057 1804 3063
rect 1869 3057 1884 3063
rect 2013 3057 2051 3063
rect 2429 3057 2444 3063
rect 2788 3056 2796 3064
rect 2829 3057 2867 3063
rect 2877 3057 2915 3063
rect 3149 3057 3180 3063
rect 3524 3056 3532 3064
rect 3853 3057 3859 3077
rect 3933 3057 3971 3063
rect 4125 3057 4131 3077
rect 4541 3057 4556 3063
rect 4740 3057 4771 3063
rect 4836 3057 4867 3063
rect 5005 3057 5020 3063
rect 5124 3057 5139 3063
rect 5149 3057 5196 3063
rect 202 3036 204 3044
rect 922 3036 924 3044
rect 3236 3036 3238 3044
rect 3322 3036 3324 3044
rect 4410 3036 4412 3044
rect 5526 3016 5626 3404
rect 5206 3004 5626 3016
rect 1706 2976 1708 2984
rect 2564 2976 2566 2984
rect 3220 2976 3222 2984
rect 3460 2976 3462 2984
rect 4458 2976 4460 2984
rect 93 2957 124 2963
rect 573 2943 579 2963
rect 1037 2957 1075 2963
rect 1213 2957 1251 2963
rect 1332 2957 1347 2963
rect 1860 2957 1884 2963
rect 541 2937 579 2943
rect 589 2937 627 2943
rect 52 2917 67 2923
rect 189 2917 227 2923
rect 292 2917 307 2923
rect 621 2917 627 2937
rect 749 2937 764 2943
rect 909 2937 940 2943
rect 1332 2937 1363 2943
rect 1581 2937 1619 2943
rect 1780 2937 1811 2943
rect 1981 2943 1987 2963
rect 2100 2957 2131 2963
rect 2141 2957 2179 2963
rect 2189 2957 2204 2963
rect 1949 2937 1987 2943
rect 2221 2937 2252 2943
rect 708 2917 739 2923
rect 932 2917 940 2923
rect 1053 2917 1068 2923
rect 1101 2917 1123 2923
rect 1229 2917 1244 2923
rect 1277 2917 1292 2923
rect 1325 2917 1340 2923
rect 1380 2917 1395 2923
rect 1476 2917 1491 2923
rect 1565 2917 1596 2923
rect 1661 2917 1699 2923
rect 484 2897 499 2903
rect 1693 2897 1699 2917
rect 2333 2923 2339 2963
rect 2388 2957 2403 2963
rect 2612 2956 2620 2964
rect 2381 2937 2396 2943
rect 2333 2917 2348 2923
rect 2381 2917 2387 2937
rect 2532 2937 2547 2943
rect 2580 2937 2595 2943
rect 2628 2937 2659 2943
rect 2829 2943 2835 2963
rect 3908 2956 3916 2964
rect 2797 2937 2835 2943
rect 3085 2937 3123 2943
rect 3188 2937 3203 2943
rect 3236 2937 3267 2943
rect 3277 2937 3315 2943
rect 2404 2917 2419 2923
rect 2525 2917 2540 2923
rect 2676 2917 2691 2923
rect 2861 2917 2883 2923
rect 2900 2917 2915 2923
rect 3044 2917 3084 2923
rect 3117 2917 3148 2923
rect 3645 2923 3651 2943
rect 3725 2937 3763 2943
rect 4029 2937 4044 2943
rect 4205 2943 4211 2963
rect 4205 2937 4243 2943
rect 4477 2937 4492 2943
rect 4605 2937 4620 2943
rect 3645 2917 3683 2923
rect 3981 2917 3996 2923
rect 4660 2917 4691 2923
rect 4845 2923 4851 2943
rect 4845 2917 4883 2923
rect 4893 2917 4931 2923
rect 4013 2897 4051 2903
rect 4893 2897 4899 2917
rect 4964 2917 4979 2923
rect 4989 2917 5004 2923
rect 380 2884 388 2888
rect 716 2884 724 2888
rect 1402 2876 1404 2884
rect 1548 2883 1556 2888
rect 1772 2884 1780 2888
rect 1517 2877 1556 2883
rect 1788 2884 1796 2888
rect 3004 2884 3012 2888
rect 2004 2876 2006 2884
rect 3900 2884 3908 2888
rect 3996 2883 4004 2888
rect 3981 2877 4004 2883
rect 4396 2884 4404 2888
rect 4444 2884 4452 2888
rect 4572 2883 4580 2888
rect 4557 2877 4580 2883
rect 4620 2884 4628 2888
rect 5148 2884 5156 2888
rect 4637 2877 4652 2883
rect 634 2836 636 2844
rect 4778 2836 4780 2844
rect -408 2804 6 2816
rect -408 2416 -308 2804
rect 1722 2776 1724 2784
rect 3034 2776 3036 2784
rect 572 2732 580 2736
rect 1245 2737 1260 2743
rect 2100 2737 2131 2743
rect 764 2732 772 2736
rect 2140 2732 2148 2736
rect 2236 2737 2259 2743
rect 2236 2732 2244 2737
rect 2324 2737 2340 2743
rect 2332 2732 2340 2737
rect 2724 2737 2739 2743
rect 3725 2737 3748 2743
rect 2588 2732 2596 2736
rect 2796 2732 2804 2736
rect 3740 2732 3748 2737
rect 5172 2737 5187 2743
rect 4348 2732 4356 2736
rect 4812 2732 4820 2736
rect 5148 2732 5156 2736
rect 93 2717 108 2723
rect 164 2697 179 2703
rect 381 2697 396 2703
rect 429 2697 467 2703
rect 749 2703 755 2723
rect 749 2697 787 2703
rect 829 2697 867 2703
rect 1037 2697 1075 2703
rect 1181 2697 1196 2703
rect 1293 2697 1324 2703
rect 1453 2697 1491 2703
rect 1661 2703 1667 2723
rect 2276 2717 2291 2723
rect 3396 2717 3411 2723
rect 1629 2697 1667 2703
rect 1748 2697 1795 2703
rect 1997 2703 2003 2716
rect 1965 2697 2003 2703
rect 2125 2697 2156 2703
rect 2221 2697 2236 2703
rect 2349 2697 2387 2703
rect 2445 2697 2467 2703
rect 2877 2697 2892 2703
rect 2989 2697 3027 2703
rect 3325 2697 3356 2703
rect 3469 2697 3484 2703
rect 3821 2703 3827 2723
rect 3773 2697 3811 2703
rect 3821 2697 3859 2703
rect 3869 2697 3884 2703
rect 52 2677 67 2683
rect 605 2677 643 2683
rect 660 2677 675 2683
rect 708 2677 723 2683
rect 1021 2677 1036 2683
rect 1117 2677 1148 2683
rect 2029 2677 2051 2683
rect 2365 2677 2380 2683
rect 2477 2677 2492 2683
rect 2637 2677 2675 2683
rect 228 2657 252 2663
rect 308 2657 323 2663
rect 365 2657 403 2663
rect 436 2657 451 2663
rect 900 2657 924 2663
rect 980 2657 1011 2663
rect 1188 2657 1203 2663
rect 1389 2657 1427 2663
rect 2525 2657 2563 2663
rect 2573 2657 2604 2663
rect 2669 2657 2675 2677
rect 2708 2677 2723 2683
rect 2804 2677 2835 2683
rect 3341 2677 3379 2683
rect 3421 2677 3459 2683
rect 2788 2657 2819 2663
rect 3220 2656 3228 2664
rect 3421 2657 3427 2677
rect 3476 2677 3491 2683
rect 3597 2677 3628 2683
rect 3693 2677 3708 2683
rect 3773 2677 3779 2697
rect 4068 2697 4083 2703
rect 4388 2697 4403 2703
rect 4621 2703 4627 2723
rect 4621 2697 4659 2703
rect 5021 2703 5027 2723
rect 4989 2697 5027 2703
rect 3876 2677 3891 2683
rect 4221 2677 4252 2683
rect 4333 2677 4371 2683
rect 4525 2677 4595 2683
rect 4941 2677 4972 2683
rect 5108 2677 5123 2683
rect 3572 2657 3587 2663
rect 3748 2656 3756 2664
rect 3956 2657 3987 2663
rect 3997 2657 4012 2663
rect 4109 2657 4140 2663
rect 4701 2657 4716 2663
rect 4804 2657 4835 2663
rect 5140 2657 5171 2663
rect 84 2636 86 2644
rect 132 2636 134 2644
rect 836 2636 838 2644
rect 1588 2636 1590 2644
rect 1674 2636 1676 2644
rect 3130 2636 3132 2644
rect 3188 2636 3190 2644
rect 3508 2636 3510 2644
rect 4052 2636 4054 2644
rect 4314 2636 4316 2644
rect 5526 2616 5626 3004
rect 5206 2604 5626 2616
rect 1636 2576 1638 2584
rect 1946 2576 1948 2584
rect 2426 2576 2428 2584
rect 2474 2576 2476 2584
rect 2986 2576 2988 2584
rect 3716 2576 3718 2584
rect 4004 2576 4006 2584
rect 4042 2576 4044 2584
rect 4180 2576 4182 2584
rect 4324 2576 4326 2584
rect 4730 2576 4732 2584
rect 36 2557 67 2563
rect 301 2543 307 2563
rect 413 2557 428 2563
rect 269 2537 307 2543
rect 317 2537 332 2543
rect 717 2537 748 2543
rect 797 2543 803 2563
rect 1044 2557 1059 2563
rect 1124 2557 1139 2563
rect 1572 2557 1587 2563
rect 1725 2557 1747 2563
rect 2132 2556 2140 2564
rect 2356 2557 2380 2563
rect 2701 2557 2716 2563
rect 2845 2557 2876 2563
rect 788 2537 803 2543
rect 1149 2537 1164 2543
rect 1373 2537 1404 2543
rect 1597 2537 1619 2543
rect 1853 2537 1891 2543
rect 2157 2537 2195 2543
rect 2333 2537 2364 2543
rect 2493 2537 2508 2543
rect 2573 2537 2588 2543
rect 2724 2537 2755 2543
rect 2868 2537 2899 2543
rect 3005 2537 3020 2543
rect 173 2517 211 2523
rect 372 2517 387 2523
rect 445 2517 460 2523
rect 573 2517 611 2523
rect 605 2497 611 2517
rect 788 2517 819 2523
rect 1293 2517 1308 2523
rect 1444 2517 1459 2523
rect 1565 2517 1580 2523
rect 1773 2517 1788 2523
rect 1821 2517 1836 2523
rect 1901 2517 1939 2523
rect 1181 2497 1196 2503
rect 1933 2497 1939 2517
rect 2205 2517 2220 2523
rect 2717 2517 2732 2523
rect 3165 2523 3171 2563
rect 3245 2557 3267 2563
rect 3277 2557 3308 2563
rect 3181 2537 3219 2543
rect 3149 2517 3171 2523
rect 3149 2504 3155 2517
rect 3213 2517 3219 2537
rect 3357 2543 3363 2563
rect 3412 2557 3436 2563
rect 3357 2537 3395 2543
rect 3965 2543 3971 2563
rect 4548 2557 4579 2563
rect 4612 2557 4627 2563
rect 4788 2556 4796 2564
rect 3773 2537 3843 2543
rect 3965 2537 3980 2543
rect 4660 2537 4675 2543
rect 3492 2517 3523 2523
rect 3540 2517 3571 2523
rect 3677 2517 3692 2523
rect 4244 2517 4275 2523
rect 4493 2517 4508 2523
rect 4909 2523 4915 2543
rect 4948 2537 4979 2543
rect 4628 2517 4643 2523
rect 4653 2517 4691 2523
rect 4877 2517 4915 2523
rect 4397 2497 4435 2503
rect 4445 2497 4476 2503
rect 4756 2497 4787 2503
rect 164 2477 179 2483
rect 868 2476 870 2484
rect 2460 2483 2468 2488
rect 3420 2484 3428 2488
rect 2452 2477 2468 2483
rect 2644 2477 2659 2483
rect 3868 2484 3876 2488
rect 4188 2484 4196 2488
rect 4380 2483 4388 2488
rect 4556 2484 4564 2488
rect 4365 2477 4388 2483
rect 4812 2484 4820 2488
rect 676 2436 678 2444
rect 1098 2436 1100 2444
rect 1332 2436 1334 2444
rect 1764 2436 1766 2444
rect -408 2404 6 2416
rect -408 2016 -308 2404
rect 1588 2376 1590 2384
rect 2666 2376 2668 2384
rect 4068 2376 4070 2384
rect 762 2336 764 2344
rect 1498 2336 1500 2344
rect 2125 2337 2148 2343
rect 1260 2332 1268 2336
rect 2140 2332 2148 2337
rect 3037 2337 3060 2343
rect 3052 2332 3060 2337
rect 3124 2337 3139 2343
rect 3500 2332 3508 2336
rect 4316 2332 4324 2336
rect 4364 2337 4387 2343
rect 4364 2332 4372 2337
rect 4461 2337 4484 2343
rect 4541 2337 4564 2343
rect 4476 2332 4484 2337
rect 4556 2332 4564 2337
rect 4732 2332 4740 2336
rect 4940 2332 4948 2336
rect 2596 2317 2627 2323
rect 2893 2317 2931 2323
rect 93 2297 131 2303
rect 237 2297 275 2303
rect 717 2297 755 2303
rect 788 2297 819 2303
rect 1060 2297 1075 2303
rect 1085 2297 1123 2303
rect 1469 2303 1475 2316
rect 1469 2297 1491 2303
rect 1684 2297 1699 2303
rect 1709 2297 1724 2303
rect 1757 2297 1788 2303
rect 1821 2297 1836 2303
rect 2804 2297 2819 2303
rect 2829 2297 2844 2303
rect 3181 2303 3187 2323
rect 3156 2297 3187 2303
rect 3277 2303 3283 2323
rect 3245 2297 3283 2303
rect 3428 2297 3443 2303
rect 3485 2297 3500 2303
rect 3517 2297 3532 2303
rect 3677 2297 3715 2303
rect 3789 2303 3795 2323
rect 5133 2317 5171 2323
rect 3757 2297 3795 2303
rect 4125 2297 4140 2303
rect 45 2277 60 2283
rect 45 2257 51 2277
rect 173 2277 211 2283
rect 77 2257 92 2263
rect 205 2257 211 2277
rect 468 2277 499 2283
rect 516 2277 531 2283
rect 877 2277 892 2283
rect 877 2264 883 2277
rect 941 2277 979 2283
rect 244 2257 259 2263
rect 308 2257 323 2263
rect 413 2257 451 2263
rect 733 2257 748 2263
rect 973 2257 979 2277
rect 1108 2277 1139 2283
rect 1252 2277 1283 2283
rect 1293 2277 1308 2283
rect 1373 2277 1404 2283
rect 2228 2277 2259 2283
rect 2564 2277 2579 2283
rect 2717 2277 2732 2283
rect 1053 2257 1068 2263
rect 1149 2257 1187 2263
rect 1389 2257 1427 2263
rect 1437 2257 1459 2263
rect 2132 2257 2156 2263
rect 2685 2257 2707 2263
rect 2717 2257 2723 2277
rect 3213 2277 3251 2283
rect 3533 2277 3571 2283
rect 3821 2277 3836 2283
rect 3853 2277 3891 2283
rect 4276 2277 4291 2283
rect 4301 2277 4339 2283
rect 4717 2277 4732 2283
rect 3044 2257 3068 2263
rect 3620 2257 3651 2263
rect 3796 2256 3804 2264
rect 4484 2256 4492 2264
rect 4564 2256 4572 2264
rect 4717 2257 4723 2277
rect 4900 2277 4908 2283
rect 4868 2257 4883 2263
rect 676 2236 678 2244
rect 1908 2236 1910 2244
rect 1978 2236 1980 2244
rect 2378 2236 2380 2244
rect 4202 2236 4204 2244
rect 4676 2236 4678 2244
rect 4970 2236 4972 2244
rect 5066 2236 5068 2244
rect 5526 2216 5626 2604
rect 5206 2204 5626 2216
rect 356 2176 358 2184
rect 548 2176 550 2184
rect 922 2176 924 2184
rect 1018 2176 1020 2184
rect 1530 2176 1532 2184
rect 2228 2176 2230 2184
rect 2372 2176 2374 2184
rect 2410 2176 2412 2184
rect 2900 2176 2902 2184
rect 3482 2176 3484 2184
rect 4218 2176 4220 2184
rect 4298 2176 4300 2184
rect 4484 2176 4486 2184
rect 4628 2176 4630 2184
rect 5060 2176 5062 2184
rect 116 2157 131 2163
rect 141 2157 163 2163
rect 388 2156 396 2164
rect 644 2157 675 2163
rect 820 2157 835 2163
rect 1085 2157 1116 2163
rect 20 2137 35 2143
rect 205 2137 243 2143
rect 237 2117 243 2137
rect 756 2137 771 2143
rect 765 2117 771 2137
rect 1405 2143 1411 2163
rect 1645 2157 1660 2163
rect 1700 2157 1724 2163
rect 1764 2157 1779 2163
rect 1869 2157 1884 2163
rect 2292 2157 2316 2163
rect 3261 2157 3276 2163
rect 3837 2157 3852 2163
rect 3892 2156 3900 2164
rect 1364 2137 1379 2143
rect 1405 2137 1443 2143
rect 804 2117 819 2123
rect 852 2117 867 2123
rect 877 2117 915 2123
rect 909 2097 915 2117
rect 1069 2117 1100 2123
rect 1220 2117 1251 2123
rect 1373 2117 1379 2137
rect 1581 2137 1612 2143
rect 1652 2137 1683 2143
rect 2557 2143 2563 2156
rect 4125 2144 4131 2163
rect 4708 2156 4716 2164
rect 4900 2156 4908 2164
rect 2429 2137 2467 2143
rect 2557 2137 2595 2143
rect 2916 2137 2947 2143
rect 2957 2137 2972 2143
rect 2989 2137 3020 2143
rect 3821 2137 3836 2143
rect 3949 2137 3980 2143
rect 4548 2137 4563 2143
rect 4733 2137 4748 2143
rect 5124 2137 5139 2143
rect 1453 2117 1491 2123
rect 1604 2117 1619 2123
rect 1652 2117 1667 2123
rect 1748 2117 1763 2123
rect 1885 2117 1923 2123
rect 2036 2117 2051 2123
rect 2068 2117 2083 2123
rect 2116 2117 2131 2123
rect 3165 2117 3203 2123
rect 3357 2117 3379 2123
rect 3428 2117 3443 2123
rect 3796 2117 3811 2123
rect 3652 2097 3683 2103
rect 1948 2084 1956 2088
rect 2300 2084 2308 2088
rect 925 2077 940 2083
rect 1988 2077 2003 2083
rect 2396 2084 2404 2088
rect 2620 2084 2628 2088
rect 2828 2083 2836 2088
rect 2724 2077 2739 2083
rect 2797 2077 2836 2083
rect 2924 2084 2932 2088
rect 3108 2077 3123 2083
rect 3756 2083 3764 2088
rect 3748 2077 3764 2083
rect 4141 2077 4156 2083
rect 4412 2083 4420 2088
rect 4892 2084 4900 2088
rect 4397 2077 4420 2083
rect 4829 2077 4844 2083
rect 5116 2084 5124 2088
rect 2138 2036 2140 2044
rect -408 2004 4 2016
rect -408 1616 -308 2004
rect 1146 1976 1148 1984
rect 1274 1976 1276 1984
rect 3316 1976 3318 1984
rect 3658 1976 3660 1984
rect 2474 1956 2476 1964
rect 1677 1937 1700 1943
rect 748 1932 756 1936
rect 1692 1932 1700 1937
rect 1908 1937 1923 1943
rect 2205 1937 2220 1943
rect 2381 1937 2412 1943
rect 2812 1932 2820 1936
rect 2988 1937 3004 1943
rect 2988 1932 2996 1937
rect 3132 1932 3140 1936
rect 3980 1932 3988 1936
rect 4156 1932 4164 1936
rect 4381 1937 4404 1943
rect 4204 1932 4212 1936
rect 4396 1932 4404 1937
rect 4524 1937 4540 1943
rect 4524 1932 4532 1937
rect 4924 1932 4932 1936
rect 125 1883 131 1903
rect 205 1897 220 1903
rect 228 1897 243 1903
rect 253 1897 291 1903
rect 477 1897 515 1903
rect 669 1897 707 1903
rect 868 1897 883 1903
rect 957 1897 988 1903
rect 1076 1897 1091 1903
rect 1124 1897 1139 1903
rect 1300 1897 1331 1903
rect 1485 1903 1491 1923
rect 1453 1897 1491 1903
rect 1732 1897 1747 1903
rect 2029 1903 2035 1923
rect 2829 1917 2844 1923
rect 2029 1897 2067 1903
rect 2173 1897 2188 1903
rect 2269 1897 2300 1903
rect 2845 1897 2883 1903
rect 2925 1897 2956 1903
rect 125 1877 163 1883
rect 301 1877 339 1883
rect 333 1857 339 1877
rect 525 1877 540 1883
rect 692 1877 723 1883
rect 1517 1877 1539 1883
rect 1556 1877 1587 1883
rect 1732 1877 1740 1883
rect 1917 1877 1948 1883
rect 2397 1877 2419 1883
rect 2397 1864 2403 1877
rect 2724 1877 2739 1883
rect 2845 1877 2851 1897
rect 3533 1897 3571 1903
rect 3725 1903 3731 1923
rect 3725 1897 3763 1903
rect 3965 1903 3971 1923
rect 4685 1917 4723 1923
rect 4877 1917 4915 1923
rect 3965 1897 3980 1903
rect 4013 1897 4051 1903
rect 541 1857 572 1863
rect 676 1857 700 1863
rect 1012 1857 1036 1863
rect 2644 1856 2652 1864
rect 2733 1857 2739 1877
rect 3389 1877 3427 1883
rect 2772 1857 2787 1863
rect 3421 1857 3427 1877
rect 3629 1877 3667 1883
rect 3684 1877 3699 1883
rect 3805 1877 3843 1883
rect 3853 1877 3891 1883
rect 4013 1877 4019 1897
rect 4116 1897 4131 1903
rect 4125 1877 4131 1897
rect 4781 1897 4819 1903
rect 4164 1877 4179 1883
rect 4644 1877 4659 1883
rect 4781 1877 4787 1897
rect 5005 1897 5027 1903
rect 4836 1877 4851 1883
rect 4884 1877 4892 1883
rect 5037 1877 5075 1883
rect 5085 1877 5107 1883
rect 5181 1877 5196 1883
rect 3716 1856 3724 1864
rect 4244 1857 4275 1863
rect 5069 1857 5075 1877
rect 1498 1836 1500 1844
rect 1962 1836 1964 1844
rect 2436 1836 2438 1844
rect 3028 1836 3030 1844
rect 3268 1836 3270 1844
rect 3466 1836 3468 1844
rect 4148 1836 4150 1844
rect 4410 1836 4412 1844
rect 4868 1836 4870 1844
rect 5162 1836 5164 1844
rect 5526 1816 5626 2204
rect 5206 1804 5626 1816
rect 1012 1776 1014 1784
rect 1482 1776 1484 1784
rect 1850 1776 1852 1784
rect 3946 1776 3948 1784
rect 4196 1776 4198 1784
rect 4340 1776 4342 1784
rect 5156 1776 5158 1784
rect 45 1757 83 1763
rect 93 1757 131 1763
rect 445 1743 451 1763
rect 548 1757 563 1763
rect 628 1757 659 1763
rect 852 1756 860 1764
rect 1053 1757 1091 1763
rect 1124 1757 1139 1763
rect 1533 1757 1571 1763
rect 445 1737 460 1743
rect 1076 1737 1107 1743
rect 1124 1737 1155 1743
rect 1316 1737 1347 1743
rect 1581 1724 1587 1763
rect 1613 1757 1651 1763
rect 1748 1757 1763 1763
rect 2036 1757 2067 1763
rect 2077 1757 2108 1763
rect 2349 1757 2364 1763
rect 2397 1757 2428 1763
rect 2628 1757 2659 1763
rect 2772 1757 2796 1763
rect 3101 1744 3107 1763
rect 3117 1757 3155 1763
rect 3373 1757 3388 1763
rect 5012 1756 5020 1764
rect 1636 1737 1667 1743
rect 1725 1737 1740 1743
rect 100 1717 115 1723
rect 589 1717 604 1723
rect 685 1717 748 1723
rect 1069 1717 1084 1723
rect 1629 1717 1644 1723
rect 1725 1717 1731 1737
rect 1924 1737 1939 1743
rect 2260 1737 2275 1743
rect 2381 1737 2396 1743
rect 2788 1737 2819 1743
rect 3277 1737 3315 1743
rect 3533 1737 3571 1743
rect 3613 1737 3651 1743
rect 4013 1737 4028 1743
rect 4068 1737 4099 1743
rect 4253 1737 4268 1743
rect 4836 1737 4851 1743
rect 5028 1737 5043 1743
rect 1997 1717 2003 1736
rect 2356 1717 2371 1723
rect 3389 1717 3427 1723
rect 3709 1717 3740 1723
rect 4109 1717 4124 1723
rect 4157 1717 4172 1723
rect 4372 1717 4387 1723
rect 4525 1717 4563 1723
rect 4621 1717 4652 1723
rect 4717 1717 4748 1723
rect 4877 1717 4915 1723
rect 909 1697 947 1703
rect 1796 1697 1811 1703
rect 2573 1697 2588 1703
rect 2733 1697 2748 1703
rect 3924 1697 3939 1703
rect 4877 1697 4883 1717
rect 5076 1717 5091 1723
rect 4932 1697 4947 1703
rect 1020 1684 1028 1688
rect 2044 1684 2052 1688
rect 2780 1684 2788 1688
rect 189 1677 204 1683
rect 1508 1677 1523 1683
rect 2685 1677 2700 1683
rect 2890 1676 2892 1684
rect 3500 1683 3508 1688
rect 3485 1677 3508 1683
rect 3676 1683 3684 1688
rect 4828 1684 4836 1688
rect 3676 1677 3699 1683
rect 5068 1684 5076 1688
rect 2234 1656 2236 1664
rect 2330 1636 2332 1644
rect 3802 1636 3804 1644
rect 4042 1636 4044 1644
rect -408 1604 6 1616
rect -408 1216 -308 1604
rect 2541 1577 2563 1583
rect 2557 1564 2563 1577
rect 4810 1576 4812 1584
rect 2541 1557 2556 1563
rect 1092 1537 1123 1543
rect 1380 1537 1395 1543
rect 1661 1537 1676 1543
rect 1484 1532 1492 1536
rect 1772 1532 1780 1536
rect 1996 1532 2004 1536
rect 2268 1532 2276 1536
rect 2541 1537 2556 1543
rect 4324 1537 4340 1543
rect 2316 1532 2324 1536
rect 3500 1532 3508 1536
rect 4332 1532 4340 1537
rect 5020 1537 5043 1543
rect 5020 1532 5028 1537
rect 1812 1517 1827 1523
rect 381 1497 396 1503
rect 637 1497 652 1503
rect 685 1497 707 1503
rect 973 1497 1011 1503
rect 1693 1497 1731 1503
rect 1901 1503 1907 1523
rect 3412 1517 3427 1523
rect 1901 1497 1939 1503
rect 1949 1497 1964 1503
rect 2132 1497 2147 1503
rect 2180 1497 2195 1503
rect 2276 1497 2307 1503
rect 2605 1497 2620 1503
rect 2653 1497 2668 1503
rect 2788 1497 2803 1503
rect 3501 1503 3507 1523
rect 3501 1497 3539 1503
rect 3853 1503 3859 1523
rect 3725 1497 3747 1503
rect 3821 1497 3859 1503
rect 3997 1497 4012 1503
rect 4420 1497 4435 1503
rect 4445 1497 4460 1503
rect 4685 1503 4691 1523
rect 4685 1497 4723 1503
rect 20 1477 35 1483
rect 141 1477 156 1483
rect 596 1477 627 1483
rect 1325 1477 1347 1483
rect 1437 1477 1459 1483
rect 1933 1477 1971 1483
rect 2077 1477 2092 1483
rect 2157 1477 2188 1483
rect 2445 1477 2476 1483
rect 3885 1477 3907 1483
rect 4045 1477 4060 1483
rect 173 1457 188 1463
rect 324 1457 348 1463
rect 388 1457 403 1463
rect 413 1457 428 1463
rect 509 1457 531 1463
rect 580 1457 611 1463
rect 717 1457 755 1463
rect 788 1457 803 1463
rect 893 1457 931 1463
rect 1037 1457 1068 1463
rect 2093 1457 2115 1463
rect 2173 1457 2211 1463
rect 2340 1456 2348 1464
rect 2660 1457 2675 1463
rect 2708 1456 2716 1464
rect 2781 1457 2819 1463
rect 3053 1457 3075 1463
rect 3917 1457 3948 1463
rect 4045 1457 4051 1477
rect 4317 1477 4332 1483
rect 4365 1477 4380 1483
rect 4500 1477 4515 1483
rect 4573 1477 4604 1483
rect 4276 1457 4300 1463
rect 4340 1456 4348 1464
rect 4509 1457 4515 1477
rect 4829 1457 4860 1463
rect 84 1436 86 1444
rect 1306 1436 1308 1444
rect 1476 1436 1478 1444
rect 1786 1436 1788 1444
rect 1988 1436 1990 1444
rect 2858 1436 2860 1444
rect 3162 1436 3164 1444
rect 3434 1436 3436 1444
rect 4676 1436 4678 1444
rect 4858 1436 4860 1444
rect 4906 1436 4908 1444
rect 5526 1416 5626 1804
rect 5206 1404 5626 1416
rect 458 1376 460 1384
rect 1364 1376 1366 1384
rect 1498 1376 1500 1384
rect 1604 1376 1606 1384
rect 1684 1376 1686 1384
rect 2004 1376 2006 1384
rect 2340 1376 2342 1384
rect 3156 1376 3158 1384
rect 3620 1376 3622 1384
rect 3668 1376 3670 1384
rect 125 1357 163 1363
rect 276 1357 307 1363
rect 317 1357 355 1363
rect 532 1356 540 1364
rect 676 1357 700 1363
rect 868 1356 876 1364
rect 980 1357 995 1363
rect 1149 1357 1187 1363
rect 45 1337 60 1343
rect 244 1337 259 1343
rect 740 1337 755 1343
rect 980 1337 1011 1343
rect 1252 1337 1283 1343
rect 1325 1343 1331 1363
rect 1428 1357 1443 1363
rect 1748 1357 1772 1363
rect 1844 1357 1859 1363
rect 1885 1344 1891 1363
rect 2669 1357 2707 1363
rect 2836 1356 2844 1364
rect 2893 1357 2931 1363
rect 1325 1337 1340 1343
rect 2109 1343 2115 1356
rect 2068 1337 2099 1343
rect 2109 1337 2147 1343
rect 2493 1324 2499 1343
rect 3117 1337 3139 1343
rect 3172 1337 3187 1343
rect 3245 1324 3251 1363
rect 3821 1357 3836 1363
rect 3277 1337 3315 1343
rect 3780 1337 3811 1343
rect 3876 1337 3891 1343
rect 3949 1337 3964 1343
rect 4452 1337 4467 1343
rect 4724 1337 4755 1343
rect 5037 1337 5075 1343
rect 164 1317 179 1323
rect 189 1317 227 1323
rect 237 1317 252 1323
rect 925 1317 963 1323
rect 973 1317 988 1323
rect 1021 1317 1059 1323
rect 1165 1317 1180 1323
rect 1373 1317 1411 1323
rect 1421 1317 1436 1323
rect 1373 1297 1379 1317
rect 1565 1317 1580 1323
rect 1693 1317 1731 1323
rect 1693 1297 1699 1317
rect 1876 1317 1907 1323
rect 2189 1317 2227 1323
rect 1940 1297 1955 1303
rect 2221 1297 2227 1317
rect 2372 1317 2387 1323
rect 2621 1317 2652 1323
rect 2685 1317 2700 1323
rect 2733 1317 2748 1323
rect 2797 1317 2812 1323
rect 2852 1317 2867 1323
rect 2900 1317 2915 1323
rect 3341 1317 3379 1323
rect 3341 1297 3347 1317
rect 3533 1317 3571 1323
rect 3421 1297 3436 1303
rect 3533 1297 3539 1317
rect 3869 1317 3884 1323
rect 4109 1317 4140 1323
rect 4237 1317 4268 1323
rect 4644 1317 4659 1323
rect 5085 1317 5116 1323
rect 5181 1317 5212 1323
rect 3629 1297 3644 1303
rect 684 1283 692 1288
rect 564 1277 579 1283
rect 669 1277 692 1283
rect 1484 1283 1492 1288
rect 1300 1277 1315 1283
rect 1469 1277 1492 1283
rect 1612 1284 1620 1288
rect 2060 1284 2068 1288
rect 3164 1284 3172 1288
rect 2260 1277 2275 1283
rect 2420 1277 2435 1283
rect 3740 1284 3748 1288
rect 4076 1284 4084 1288
rect 4029 1277 4044 1283
rect 4492 1283 4500 1288
rect 4812 1284 4820 1288
rect 4468 1277 4483 1283
rect 4492 1277 4508 1283
rect 5116 1284 5124 1288
rect 1108 1236 1110 1244
rect 3066 1236 3068 1244
rect 3284 1236 3286 1244
rect 3380 1236 3382 1244
rect 3706 1236 3708 1244
rect -408 1204 6 1216
rect -408 816 -308 1204
rect 170 1176 172 1184
rect 538 1176 540 1184
rect 3757 1177 3772 1183
rect 26 1156 28 1164
rect 1732 1163 1734 1164
rect 1732 1157 1740 1163
rect 1732 1156 1734 1157
rect 3757 1157 3772 1163
rect 1524 1137 1555 1143
rect 2525 1137 2548 1143
rect 1260 1132 1268 1136
rect 1804 1132 1812 1136
rect 2540 1132 2548 1137
rect 2620 1137 2636 1143
rect 2620 1132 2628 1137
rect 3316 1137 3332 1143
rect 3324 1132 3332 1137
rect 3757 1137 3772 1143
rect 3564 1132 3572 1136
rect 3884 1132 3892 1136
rect 3964 1132 3972 1136
rect 4060 1137 4076 1143
rect 4060 1132 4068 1137
rect 4108 1132 4116 1136
rect 4300 1137 4323 1143
rect 4300 1132 4308 1137
rect 4596 1137 4612 1143
rect 4604 1132 4612 1137
rect 4740 1137 4756 1143
rect 4748 1132 4756 1137
rect 5116 1132 5124 1136
rect 333 1097 355 1103
rect 589 1097 620 1103
rect 1405 1103 1411 1123
rect 1565 1117 1580 1123
rect 2445 1117 2460 1123
rect 2557 1117 2588 1123
rect 3453 1117 3468 1123
rect 3924 1117 3955 1123
rect 1373 1097 1411 1103
rect 1773 1097 1804 1103
rect 2989 1097 3027 1103
rect 3341 1097 3379 1103
rect 269 1077 307 1083
rect 189 1057 220 1063
rect 301 1057 307 1077
rect 605 1077 620 1083
rect 909 1077 947 1083
rect 980 1077 1011 1083
rect 1197 1083 1203 1096
rect 1197 1077 1219 1083
rect 1437 1077 1452 1083
rect 1469 1077 1484 1083
rect 1517 1083 1523 1096
rect 1517 1077 1539 1083
rect 1693 1077 1708 1083
rect 388 1056 396 1064
rect 557 1057 588 1063
rect 644 1057 675 1063
rect 749 1057 780 1063
rect 1693 1057 1699 1077
rect 2045 1077 2067 1083
rect 2084 1077 2099 1083
rect 2381 1077 2419 1083
rect 2628 1077 2643 1083
rect 2724 1077 2755 1083
rect 2941 1077 2979 1083
rect 2340 1056 2348 1064
rect 2484 1057 2515 1063
rect 2852 1056 2860 1064
rect 2941 1057 2947 1077
rect 3117 1077 3148 1083
rect 3245 1077 3276 1083
rect 3309 1077 3324 1083
rect 3373 1077 3379 1097
rect 3725 1097 3740 1103
rect 3917 1097 3932 1103
rect 3460 1077 3475 1083
rect 3677 1077 3692 1083
rect 3780 1077 3811 1083
rect 3917 1077 3923 1097
rect 4125 1103 4131 1123
rect 4093 1097 4131 1103
rect 4429 1097 4444 1103
rect 4493 1097 4508 1103
rect 4845 1103 4851 1123
rect 5165 1117 5180 1123
rect 4813 1097 4851 1103
rect 4932 1097 4947 1103
rect 3997 1077 4035 1083
rect 4068 1077 4083 1083
rect 4116 1077 4147 1083
rect 4157 1077 4172 1083
rect 4237 1077 4275 1083
rect 4589 1077 4604 1083
rect 4644 1077 4675 1083
rect 4733 1077 4748 1083
rect 4781 1077 4796 1083
rect 4877 1077 4915 1083
rect 5053 1077 5091 1083
rect 3069 1057 3084 1063
rect 3732 1057 3747 1063
rect 4852 1056 4860 1064
rect 964 1036 966 1044
rect 1130 1036 1132 1044
rect 1274 1036 1276 1044
rect 1636 1036 1638 1044
rect 2026 1036 2028 1044
rect 2436 1036 2438 1044
rect 2612 1036 2614 1044
rect 2804 1036 2806 1044
rect 3396 1036 3398 1044
rect 4570 1036 4572 1044
rect 5108 1036 5110 1044
rect 5526 1016 5626 1404
rect 5206 1004 5626 1016
rect 36 976 38 984
rect 122 976 124 984
rect 506 976 508 984
rect 698 976 700 984
rect 1044 976 1046 984
rect 1220 976 1222 984
rect 1354 976 1356 984
rect 1508 976 1510 984
rect 1770 976 1772 984
rect 2154 976 2156 984
rect 2346 976 2348 984
rect 3380 976 3382 984
rect 3700 976 3702 984
rect 4292 976 4294 984
rect 5044 976 5046 984
rect 260 956 268 964
rect 548 956 556 964
rect 669 957 700 963
rect 93 937 108 943
rect 381 937 396 943
rect 189 917 227 923
rect 189 897 195 917
rect 436 917 444 923
rect 461 917 499 923
rect 605 917 643 923
rect 493 897 499 917
rect 532 897 547 903
rect 557 897 595 903
rect 749 903 755 963
rect 788 957 812 963
rect 941 957 972 963
rect 1076 957 1091 963
rect 964 937 979 943
rect 909 917 924 923
rect 973 917 979 937
rect 1101 943 1107 963
rect 1101 937 1116 943
rect 1293 943 1299 963
rect 1428 957 1443 963
rect 1556 957 1587 963
rect 1597 957 1635 963
rect 1892 956 1900 964
rect 2196 956 2204 964
rect 2253 957 2268 963
rect 2317 957 2348 963
rect 2388 956 2396 964
rect 2596 957 2627 963
rect 2637 957 2652 963
rect 2900 957 2915 963
rect 3037 957 3059 963
rect 3069 957 3100 963
rect 3252 956 3260 964
rect 3332 956 3340 964
rect 3741 957 3772 963
rect 4020 956 4028 964
rect 4212 957 4227 963
rect 4637 957 4659 963
rect 1261 937 1299 943
rect 1501 937 1539 943
rect 1789 937 1827 943
rect 1917 937 1932 943
rect 3117 937 3155 943
rect 3172 937 3187 943
rect 3220 937 3235 943
rect 3421 937 3436 943
rect 1236 917 1251 923
rect 1380 917 1395 923
rect 2013 917 2051 923
rect 2733 917 2748 923
rect 2845 917 2860 923
rect 2996 917 3011 923
rect 3165 917 3180 923
rect 3197 917 3228 923
rect 3517 923 3523 943
rect 3645 937 3676 943
rect 3812 937 3827 943
rect 4356 937 4387 943
rect 4861 937 4876 943
rect 4941 937 4979 943
rect 5165 924 5171 943
rect 3421 917 3443 923
rect 3517 917 3555 923
rect 3812 917 3843 923
rect 3956 917 3971 923
rect 4052 917 4067 923
rect 4157 917 4172 923
rect 4260 917 4268 923
rect 4356 917 4371 923
rect 4452 917 4483 923
rect 4541 917 4579 923
rect 749 897 764 903
rect 1517 897 1532 903
rect 1988 897 2019 903
rect 3076 897 3091 903
rect 4301 897 4316 903
rect 4541 897 4547 917
rect 4893 917 4908 923
rect 4989 917 5020 923
rect 5053 917 5091 923
rect 4676 897 4691 903
rect 4820 897 4835 903
rect 5053 897 5059 917
rect 476 884 484 888
rect 1756 884 1764 888
rect 1804 884 1812 888
rect 826 876 828 884
rect 1773 877 1788 883
rect 2748 883 2756 888
rect 3580 884 3588 888
rect 2548 877 2563 883
rect 2748 877 2771 883
rect 2941 877 2956 883
rect 3708 884 3716 888
rect 3852 884 3860 888
rect 4348 884 4356 888
rect 3901 877 3916 883
rect 4493 877 4508 883
rect 986 836 988 844
rect -408 804 4 816
rect -408 416 -308 804
rect 442 776 444 784
rect 1124 756 1126 764
rect 548 736 550 744
rect 796 737 812 743
rect 796 732 804 737
rect 1044 737 1075 743
rect 2212 737 2227 743
rect 2461 737 2476 743
rect 2909 737 2932 743
rect 956 732 964 736
rect 1084 732 1092 736
rect 2140 732 2148 736
rect 2508 732 2516 736
rect 2924 732 2932 737
rect 3340 732 3348 736
rect 3388 732 3396 736
rect 3740 732 3748 736
rect 3916 737 3932 743
rect 3916 732 3924 737
rect 4324 737 4339 743
rect 4781 737 4796 743
rect 4012 732 4020 736
rect 4396 732 4404 736
rect 4828 732 4836 736
rect 4876 732 4884 736
rect 5132 732 5140 736
rect 1261 717 1299 723
rect 1309 717 1331 723
rect 1613 717 1628 723
rect 93 697 115 703
rect 301 677 332 683
rect 669 683 675 703
rect 877 697 915 703
rect 1133 697 1148 703
rect 1469 697 1507 703
rect 1741 697 1779 703
rect 1901 697 1939 703
rect 1956 697 1971 703
rect 2212 697 2227 703
rect 2317 697 2332 703
rect 2461 697 2476 703
rect 2637 703 2643 723
rect 2820 717 2835 723
rect 2637 697 2675 703
rect 2733 697 2748 703
rect 3133 697 3148 703
rect 3485 697 3500 703
rect 3780 697 3795 703
rect 4157 697 4172 703
rect 4557 703 4563 723
rect 4525 697 4563 703
rect 564 677 579 683
rect 637 677 675 683
rect 708 677 739 683
rect 989 677 1004 683
rect 1812 677 1827 683
rect 1949 677 1964 683
rect 2429 683 2435 696
rect 2420 677 2435 683
rect 2685 677 2700 683
rect 2740 677 2771 683
rect 3037 677 3052 683
rect 3277 677 3315 683
rect 3348 677 3363 683
rect 3492 677 3507 683
rect 3613 677 3651 683
rect 3773 677 3788 683
rect 3821 683 3827 696
rect 3821 677 3836 683
rect 3853 677 3891 683
rect 4020 677 4051 683
rect 4164 677 4179 683
rect 4404 677 4435 683
rect 4452 677 4467 683
rect 4589 677 4604 683
rect 4861 677 4899 683
rect 4989 677 5011 683
rect 5044 677 5075 683
rect 1140 657 1155 663
rect 2397 657 2412 663
rect 2788 657 2803 663
rect 3085 657 3100 663
rect 3117 657 3132 663
rect 3572 657 3596 663
rect 4388 657 4412 663
rect 4724 657 4755 663
rect 4836 656 4844 664
rect 36 636 38 644
rect 788 636 790 644
rect 836 636 838 644
rect 970 636 972 644
rect 1252 636 1254 644
rect 1658 636 1660 644
rect 1844 636 1846 644
rect 2500 636 2502 644
rect 2996 636 2998 644
rect 3332 636 3334 644
rect 3524 636 3526 644
rect 3754 636 3756 644
rect 3908 636 3910 644
rect 4570 636 4572 644
rect 4628 636 4630 644
rect 5124 636 5126 644
rect 5526 616 5626 1004
rect 5206 604 5626 616
rect 346 576 348 584
rect 2084 576 2086 584
rect 2916 576 2918 584
rect 3482 576 3484 584
rect 29 557 44 563
rect 125 537 156 543
rect 285 543 291 563
rect 253 537 291 543
rect 429 543 435 563
rect 964 557 988 563
rect 1172 557 1203 563
rect 1213 557 1251 563
rect 1261 557 1299 563
rect 1309 557 1340 563
rect 397 537 435 543
rect 788 537 803 543
rect 820 537 851 543
rect 1389 543 1395 563
rect 1485 557 1523 563
rect 2365 557 2380 563
rect 1357 537 1395 543
rect 1540 537 1555 543
rect 1684 537 1699 543
rect 2317 537 2348 543
rect 2413 537 2444 543
rect 2541 543 2547 563
rect 3101 557 3116 563
rect 3172 557 3187 563
rect 3533 557 3564 563
rect 3613 557 3644 563
rect 3796 557 3811 563
rect 4413 557 4444 563
rect 4532 556 4540 564
rect 2509 537 2547 543
rect 2637 537 2668 543
rect 3245 537 3276 543
rect 3389 537 3427 543
rect 3501 537 3523 543
rect 3661 537 3692 543
rect 4749 543 4755 563
rect 4909 543 4915 563
rect 5149 557 5196 563
rect 4749 537 4787 543
rect 4909 537 4947 543
rect 45 517 83 523
rect 100 517 115 523
rect 148 517 179 523
rect 317 517 332 523
rect 461 517 492 523
rect 637 517 675 523
rect 733 517 748 523
rect 861 517 876 523
rect 957 517 972 523
rect 1053 517 1068 523
rect 1277 517 1292 523
rect 1332 517 1347 523
rect 1380 517 1411 523
rect 1629 517 1644 523
rect 1789 517 1804 523
rect 2381 517 2396 523
rect 2436 517 2451 523
rect 2484 517 2499 523
rect 2612 517 2627 523
rect 2749 517 2787 523
rect 2749 497 2755 517
rect 3092 517 3107 523
rect 3316 517 3324 523
rect 3437 517 3475 523
rect 3469 497 3475 517
rect 3780 517 3795 523
rect 3901 517 3932 523
rect 4061 517 4099 523
rect 4061 497 4067 517
rect 4349 517 4387 523
rect 1180 484 1188 488
rect 948 476 950 484
rect 1852 484 1860 488
rect 1996 484 2004 488
rect 1949 477 1964 483
rect 2332 484 2340 488
rect 2029 477 2051 483
rect 2045 463 2051 477
rect 2428 484 2436 488
rect 2572 483 2580 488
rect 3452 484 3460 488
rect 2557 477 2580 483
rect 3692 484 3700 488
rect 3916 484 3924 488
rect 4716 484 4724 488
rect 3869 477 3884 483
rect 4669 477 4684 483
rect 5021 477 5036 483
rect 2029 457 2051 463
rect 2045 444 2051 457
rect 2458 456 2460 464
rect 2029 437 2044 443
rect 2132 436 2134 444
rect 2634 436 2636 444
rect 3156 443 3158 444
rect 3156 437 3164 443
rect 3156 436 3158 437
rect 3290 436 3292 444
rect 4394 436 4396 444
rect -408 404 4 416
rect -408 16 -308 404
rect 3588 376 3590 384
rect 852 337 867 343
rect 2893 337 2908 343
rect 3405 337 3428 343
rect 604 332 612 336
rect 1388 332 1396 336
rect 2060 332 2068 336
rect 3420 332 3428 337
rect 4004 336 4006 344
rect 4604 332 4612 336
rect 4836 337 4852 343
rect 4668 332 4676 336
rect 4844 332 4852 337
rect 5020 332 5028 336
rect 52 317 67 323
rect 180 297 211 303
rect 340 297 355 303
rect 589 297 604 303
rect 909 303 915 323
rect 877 297 915 303
rect 1021 297 1059 303
rect 1693 297 1708 303
rect 1741 297 1756 303
rect 1837 297 1852 303
rect 2013 297 2051 303
rect 2125 297 2163 303
rect 2317 303 2323 323
rect 2557 317 2572 323
rect 2925 317 2940 323
rect 2317 297 2355 303
rect 2372 297 2387 303
rect 2445 297 2460 303
rect 2605 303 2611 316
rect 2605 297 2643 303
rect 3053 303 3059 323
rect 3917 317 3955 323
rect 4237 317 4252 323
rect 4285 317 4300 323
rect 3053 297 3091 303
rect 173 277 188 283
rect 637 277 652 283
rect 1140 277 1171 283
rect 1533 277 1571 283
rect 1748 277 1763 283
rect 1844 277 1859 283
rect 2365 277 2380 283
rect 2461 277 2499 283
rect 100 257 115 263
rect 493 257 531 263
rect 717 257 748 263
rect 1700 257 1715 263
rect 2189 257 2227 263
rect 2237 257 2259 263
rect 2308 256 2316 264
rect 2461 257 2467 277
rect 2845 277 2883 283
rect 2893 277 2908 283
rect 2596 256 2604 264
rect 2845 257 2851 277
rect 2893 264 2899 277
rect 3012 277 3027 283
rect 3037 277 3068 283
rect 3117 283 3123 303
rect 3204 297 3219 303
rect 3252 297 3267 303
rect 3485 297 3516 303
rect 3613 303 3619 316
rect 3597 297 3619 303
rect 3629 297 3660 303
rect 3700 297 3715 303
rect 4756 297 4787 303
rect 4925 297 4963 303
rect 3085 277 3123 283
rect 3229 277 3260 283
rect 3748 277 3763 283
rect 4189 277 4204 283
rect 3293 257 3315 263
rect 3380 257 3395 263
rect 3476 256 3484 264
rect 3533 257 3571 263
rect 4068 257 4099 263
rect 4189 257 4195 277
rect 4420 277 4451 283
rect 4493 277 4524 283
rect 4564 277 4579 283
rect 4877 277 4915 283
rect 4989 277 5020 283
rect 4516 257 4531 263
rect 4541 257 4556 263
rect 4596 256 4604 264
rect 4644 256 4652 264
rect 4852 256 4860 264
rect 260 236 262 244
rect 804 236 806 244
rect 922 236 924 244
rect 1306 236 1308 244
rect 1588 236 1590 244
rect 2682 236 2684 244
rect 3908 236 3910 244
rect 4228 236 4230 244
rect 4404 236 4406 244
rect 5526 216 5626 604
rect 5206 204 5626 216
rect 36 176 38 184
rect 298 176 300 184
rect 612 176 614 184
rect 698 176 700 184
rect 1194 176 1196 184
rect 1732 176 1734 184
rect 1780 176 1782 184
rect 1876 176 1878 184
rect 2138 176 2140 184
rect 2346 176 2348 184
rect 2442 176 2444 184
rect 2490 176 2492 184
rect 3044 176 3046 184
rect 3492 176 3494 184
rect 77 157 115 163
rect 212 157 243 163
rect 253 157 268 163
rect 804 157 835 163
rect 845 157 883 163
rect 1069 157 1084 163
rect 1293 157 1331 163
rect 1364 157 1379 163
rect 1572 156 1580 164
rect 2196 156 2204 164
rect 2269 157 2307 163
rect 2676 157 2707 163
rect 3092 157 3123 163
rect 3236 157 3267 163
rect 3373 157 3404 163
rect 3636 157 3667 163
rect 3885 157 3923 163
rect 4180 157 4211 163
rect 132 137 163 143
rect 996 137 1011 143
rect 1092 137 1107 143
rect 1645 137 1683 143
rect 1837 137 1852 143
rect 1965 137 1996 143
rect 2077 137 2092 143
rect 2157 137 2172 143
rect 2365 137 2403 143
rect 2557 137 2572 143
rect 2605 137 2627 143
rect 2717 137 2748 143
rect 2909 137 2924 143
rect 3060 137 3075 143
rect 3204 137 3219 143
rect 3453 137 3475 143
rect 3508 137 3523 143
rect 3556 137 3571 143
rect 3604 137 3619 143
rect 3908 137 3939 143
rect 3981 137 4003 143
rect 173 117 188 123
rect 228 117 259 123
rect 365 117 403 123
rect 509 117 547 123
rect 861 117 876 123
rect 989 117 1027 123
rect 1037 117 1075 123
rect 893 97 908 103
rect 1037 97 1043 117
rect 1357 117 1395 123
rect 1405 117 1443 123
rect 1789 117 1827 123
rect 1460 97 1475 103
rect 1604 97 1619 103
rect 1789 97 1795 117
rect 1940 117 1955 123
rect 2749 117 2755 136
rect 4269 124 4275 163
rect 4388 156 4396 164
rect 4580 157 4611 163
rect 4621 157 4643 163
rect 4925 157 4956 163
rect 4349 137 4371 143
rect 4717 137 4755 143
rect 3309 117 3347 123
rect 3677 117 3699 123
rect 3709 117 3724 123
rect 3821 117 3843 123
rect 4013 117 4044 123
rect 4221 117 4243 123
rect 4717 117 4723 137
rect 4788 117 4803 123
rect 5005 117 5027 123
rect 5108 117 5123 123
rect 2564 97 2579 103
rect 3549 97 3564 103
rect 4461 97 4476 103
rect 4541 97 4556 103
rect 44 83 52 88
rect 812 84 820 88
rect 44 77 67 83
rect 765 77 780 83
rect 1132 83 1140 88
rect 1932 84 1940 88
rect 1132 77 1155 83
rect 1533 77 1548 83
rect 2332 83 2340 88
rect 2004 77 2019 83
rect 2317 77 2340 83
rect 2524 84 2532 88
rect 2924 83 2932 88
rect 2916 77 2932 83
rect 3052 84 3060 88
rect 3244 83 3252 88
rect 3500 84 3508 88
rect 4028 84 4036 88
rect 3244 77 3260 83
rect 5100 83 5108 88
rect 5085 77 5108 83
rect 2004 57 2019 63
rect 2004 37 2019 43
rect 3812 36 3814 44
rect 5526 16 5626 204
rect -408 4 4 16
rect -408 -40 -308 4
<< m2contact >>
rect 1068 3576 1076 3584
rect 1180 3576 1188 3584
rect 2188 3576 2196 3584
rect 3676 3576 3684 3584
rect 764 3556 772 3564
rect 956 3556 964 3564
rect 2060 3556 2068 3564
rect 2956 3556 2964 3564
rect 316 3536 324 3544
rect 604 3536 612 3544
rect 2460 3536 2468 3544
rect 2524 3536 2532 3544
rect 3308 3536 3316 3544
rect 4172 3536 4180 3544
rect 60 3516 68 3524
rect 156 3516 164 3524
rect 236 3516 244 3524
rect 332 3516 340 3524
rect 476 3516 484 3524
rect 556 3516 564 3524
rect 668 3516 676 3524
rect 1004 3516 1012 3524
rect 12 3496 20 3504
rect 140 3496 148 3504
rect 332 3496 340 3504
rect 364 3496 372 3504
rect 412 3496 420 3504
rect 428 3496 436 3504
rect 748 3496 756 3504
rect 796 3496 804 3504
rect 828 3496 836 3504
rect 844 3496 852 3504
rect 892 3496 900 3504
rect 1052 3496 1060 3504
rect 1132 3496 1140 3504
rect 1212 3496 1220 3504
rect 1260 3496 1268 3504
rect 1308 3516 1316 3524
rect 1388 3516 1396 3524
rect 1436 3496 1444 3504
rect 1452 3496 1460 3504
rect 1724 3516 1732 3524
rect 1820 3516 1828 3524
rect 1948 3516 1956 3524
rect 2012 3516 2020 3524
rect 2108 3516 2116 3524
rect 2604 3516 2612 3524
rect 2668 3516 2676 3524
rect 2732 3516 2740 3524
rect 2780 3516 2788 3524
rect 1708 3496 1716 3504
rect 1756 3496 1764 3504
rect 1916 3496 1924 3504
rect 2012 3496 2020 3504
rect 2076 3496 2084 3504
rect 2220 3496 2228 3504
rect 2332 3496 2340 3504
rect 2412 3496 2420 3504
rect 44 3476 52 3484
rect 92 3476 100 3484
rect 268 3476 276 3484
rect 348 3476 356 3484
rect 364 3476 372 3484
rect 508 3476 516 3484
rect 524 3476 532 3484
rect 572 3476 580 3484
rect 700 3476 708 3484
rect 716 3476 724 3484
rect 780 3476 788 3484
rect 108 3456 116 3464
rect 220 3456 228 3464
rect 236 3456 244 3464
rect 284 3456 292 3464
rect 380 3456 388 3464
rect 428 3456 436 3464
rect 460 3456 468 3464
rect 476 3456 484 3464
rect 716 3456 724 3464
rect 780 3456 788 3464
rect 972 3476 980 3484
rect 1244 3476 1252 3484
rect 1340 3476 1348 3484
rect 1356 3476 1364 3484
rect 1388 3476 1396 3484
rect 1532 3476 1540 3484
rect 1772 3476 1780 3484
rect 1820 3476 1828 3484
rect 1852 3476 1860 3484
rect 1916 3476 1924 3484
rect 2044 3476 2052 3484
rect 2252 3476 2260 3484
rect 2476 3496 2484 3504
rect 2844 3516 2852 3524
rect 2924 3516 2932 3524
rect 2972 3516 2980 3524
rect 2988 3516 2996 3524
rect 3116 3516 3124 3524
rect 3212 3516 3220 3524
rect 3228 3516 3236 3524
rect 3276 3516 3284 3524
rect 3404 3516 3412 3524
rect 3468 3516 3476 3524
rect 3516 3516 3524 3524
rect 3068 3496 3076 3504
rect 3164 3496 3172 3504
rect 3612 3516 3620 3524
rect 3644 3516 3652 3524
rect 3740 3516 3748 3524
rect 3852 3516 3860 3524
rect 3900 3516 3908 3524
rect 3948 3516 3956 3524
rect 3996 3516 4004 3524
rect 4044 3516 4052 3524
rect 4076 3516 4084 3524
rect 4220 3516 4228 3524
rect 4316 3516 4324 3524
rect 4332 3516 4340 3524
rect 4380 3516 4388 3524
rect 4412 3516 4420 3524
rect 4460 3516 4468 3524
rect 4956 3516 4964 3524
rect 5052 3516 5060 3524
rect 5132 3516 5140 3524
rect 3980 3496 3988 3504
rect 2556 3476 2564 3484
rect 2572 3476 2580 3484
rect 2668 3476 2676 3484
rect 2700 3476 2708 3484
rect 2748 3476 2756 3484
rect 2780 3476 2788 3484
rect 2892 3476 2900 3484
rect 2924 3476 2932 3484
rect 3036 3476 3044 3484
rect 3212 3476 3220 3484
rect 3276 3476 3284 3484
rect 3356 3476 3364 3484
rect 3372 3476 3380 3484
rect 3404 3476 3412 3484
rect 3452 3476 3460 3484
rect 3468 3476 3476 3484
rect 3548 3476 3556 3484
rect 3564 3476 3572 3484
rect 3596 3476 3604 3484
rect 3644 3476 3652 3484
rect 3692 3476 3700 3484
rect 3740 3476 3748 3484
rect 3788 3476 3796 3484
rect 3804 3476 3812 3484
rect 3884 3476 3892 3484
rect 3932 3476 3940 3484
rect 4028 3476 4036 3484
rect 4092 3476 4100 3484
rect 4188 3496 4196 3504
rect 4236 3496 4244 3504
rect 4268 3496 4276 3504
rect 4140 3476 4148 3484
rect 4236 3476 4244 3484
rect 4268 3476 4276 3484
rect 4476 3496 4484 3504
rect 4556 3496 4564 3504
rect 4572 3496 4580 3504
rect 4620 3496 4628 3504
rect 4700 3496 4708 3504
rect 4716 3496 4724 3504
rect 4748 3496 4756 3504
rect 4812 3496 4820 3504
rect 4828 3496 4836 3504
rect 4892 3496 4900 3504
rect 4300 3476 4308 3484
rect 4364 3476 4372 3484
rect 4380 3476 4388 3484
rect 4428 3476 4436 3484
rect 4604 3476 4612 3484
rect 5036 3496 5044 3504
rect 4988 3476 4996 3484
rect 5004 3476 5012 3484
rect 5084 3476 5092 3484
rect 5100 3476 5108 3484
rect 828 3456 836 3464
rect 924 3456 932 3464
rect 940 3456 948 3464
rect 1020 3456 1028 3464
rect 1084 3456 1092 3464
rect 1100 3456 1108 3464
rect 1148 3456 1156 3464
rect 1196 3456 1204 3464
rect 1244 3456 1252 3464
rect 1404 3456 1412 3464
rect 1484 3456 1492 3464
rect 1564 3456 1572 3464
rect 1612 3456 1620 3464
rect 1628 3456 1636 3464
rect 1676 3456 1684 3464
rect 1868 3456 1876 3464
rect 2076 3456 2084 3464
rect 2156 3456 2164 3464
rect 2172 3456 2180 3464
rect 2220 3456 2228 3464
rect 2316 3456 2324 3464
rect 2364 3456 2372 3464
rect 2380 3456 2388 3464
rect 2508 3456 2516 3464
rect 2716 3456 2724 3464
rect 2764 3456 2772 3464
rect 3036 3456 3044 3464
rect 3132 3456 3140 3464
rect 3436 3456 3444 3464
rect 4236 3456 4244 3464
rect 4508 3456 4516 3464
rect 4524 3456 4532 3464
rect 4556 3456 4564 3464
rect 4572 3456 4580 3464
rect 4652 3456 4660 3464
rect 4668 3456 4676 3464
rect 4748 3456 4756 3464
rect 4796 3456 4804 3464
rect 4844 3456 4852 3464
rect 4860 3456 4868 3464
rect 4940 3456 4948 3464
rect 4956 3456 4964 3464
rect 5164 3456 5172 3464
rect 124 3436 132 3444
rect 172 3436 180 3444
rect 540 3436 548 3444
rect 636 3436 644 3444
rect 1036 3436 1044 3444
rect 1116 3436 1124 3444
rect 1164 3436 1172 3444
rect 1292 3436 1300 3444
rect 1372 3436 1380 3444
rect 1500 3436 1508 3444
rect 1724 3436 1732 3444
rect 1884 3436 1892 3444
rect 2348 3436 2356 3444
rect 2524 3436 2532 3444
rect 2812 3436 2820 3444
rect 2908 3436 2916 3444
rect 3004 3436 3012 3444
rect 3052 3436 3060 3444
rect 3116 3436 3124 3444
rect 3196 3436 3204 3444
rect 3244 3436 3252 3444
rect 3276 3436 3284 3444
rect 3340 3436 3348 3444
rect 3388 3436 3396 3444
rect 3500 3436 3508 3444
rect 3532 3436 3540 3444
rect 3564 3436 3572 3444
rect 3612 3436 3620 3444
rect 3724 3436 3732 3444
rect 3756 3436 3764 3444
rect 3836 3436 3844 3444
rect 3900 3436 3908 3444
rect 3948 3436 3956 3444
rect 3996 3436 4004 3444
rect 4044 3436 4052 3444
rect 4108 3436 4116 3444
rect 4156 3436 4164 3444
rect 4188 3436 4196 3444
rect 4332 3436 4340 3444
rect 4396 3436 4404 3444
rect 4444 3436 4452 3444
rect 4492 3436 4500 3444
rect 4684 3436 4692 3444
rect 4732 3436 4740 3444
rect 4876 3436 4884 3444
rect 4924 3436 4932 3444
rect 5020 3436 5028 3444
rect 5116 3436 5124 3444
rect 5148 3436 5156 3444
rect 108 3376 116 3384
rect 156 3376 164 3384
rect 348 3376 356 3384
rect 636 3376 644 3384
rect 892 3376 900 3384
rect 924 3376 932 3384
rect 956 3376 964 3384
rect 1052 3376 1060 3384
rect 1132 3376 1140 3384
rect 1228 3376 1236 3384
rect 1532 3376 1540 3384
rect 1628 3376 1636 3384
rect 1756 3376 1764 3384
rect 1916 3376 1924 3384
rect 2172 3376 2180 3384
rect 2236 3376 2244 3384
rect 2300 3376 2308 3384
rect 2316 3376 2324 3384
rect 2620 3376 2628 3384
rect 3020 3376 3028 3384
rect 3100 3376 3108 3384
rect 3148 3376 3156 3384
rect 3228 3376 3236 3384
rect 3484 3376 3492 3384
rect 3548 3376 3556 3384
rect 3804 3376 3812 3384
rect 4156 3376 4164 3384
rect 4476 3376 4484 3384
rect 4764 3376 4772 3384
rect 12 3356 20 3364
rect 60 3356 68 3364
rect 300 3356 308 3364
rect 428 3356 436 3364
rect 572 3356 580 3364
rect 620 3356 628 3364
rect 716 3356 724 3364
rect 732 3356 740 3364
rect 796 3356 804 3364
rect 940 3356 948 3364
rect 972 3356 980 3364
rect 1116 3356 1124 3364
rect 1292 3356 1300 3364
rect 1324 3356 1332 3364
rect 1372 3356 1380 3364
rect 1388 3356 1396 3364
rect 1420 3356 1428 3364
rect 1452 3356 1460 3364
rect 1516 3356 1524 3364
rect 1564 3356 1572 3364
rect 1612 3356 1620 3364
rect 1724 3356 1732 3364
rect 1884 3356 1892 3364
rect 2028 3356 2036 3364
rect 2156 3356 2164 3364
rect 2220 3356 2228 3364
rect 140 3336 148 3344
rect 188 3336 196 3344
rect 284 3336 292 3344
rect 332 3336 340 3344
rect 380 3336 388 3344
rect 476 3336 484 3344
rect 540 3336 548 3344
rect 572 3336 580 3344
rect 812 3336 820 3344
rect 860 3336 868 3344
rect 972 3336 980 3344
rect 1020 3336 1028 3344
rect 1036 3336 1044 3344
rect 1164 3336 1172 3344
rect 1212 3336 1220 3344
rect 1276 3336 1284 3344
rect 1468 3336 1476 3344
rect 1644 3336 1652 3344
rect 1772 3336 1780 3344
rect 1788 3336 1796 3344
rect 2124 3336 2132 3344
rect 2268 3336 2276 3344
rect 2348 3356 2356 3364
rect 2396 3356 2404 3364
rect 2476 3356 2484 3364
rect 2508 3356 2516 3364
rect 2380 3336 2388 3344
rect 2572 3356 2580 3364
rect 2668 3356 2676 3364
rect 2700 3356 2708 3364
rect 2828 3356 2836 3364
rect 2844 3356 2852 3364
rect 2892 3356 2900 3364
rect 3196 3356 3204 3364
rect 3260 3356 3268 3364
rect 3388 3356 3396 3364
rect 3404 3356 3412 3364
rect 3564 3356 3572 3364
rect 3708 3356 3716 3364
rect 3788 3356 3796 3364
rect 3932 3356 3940 3364
rect 4012 3356 4020 3364
rect 4060 3356 4068 3364
rect 4076 3356 4084 3364
rect 4092 3356 4100 3364
rect 4220 3356 4228 3364
rect 4252 3356 4260 3364
rect 4364 3356 4372 3364
rect 4380 3356 4388 3364
rect 4396 3356 4404 3364
rect 4412 3356 4420 3364
rect 4492 3356 4500 3364
rect 4508 3356 4516 3364
rect 4556 3356 4564 3364
rect 4636 3356 4644 3364
rect 4684 3356 4692 3364
rect 4700 3356 4708 3364
rect 4748 3356 4756 3364
rect 4780 3356 4788 3364
rect 4844 3356 4852 3364
rect 4940 3356 4948 3364
rect 4988 3356 4996 3364
rect 5052 3356 5060 3364
rect 5100 3356 5108 3364
rect 5132 3356 5140 3364
rect 92 3316 100 3324
rect 204 3316 212 3324
rect 396 3316 404 3324
rect 428 3316 436 3324
rect 684 3316 692 3324
rect 716 3316 724 3324
rect 764 3316 772 3324
rect 860 3316 868 3324
rect 892 3316 900 3324
rect 1116 3316 1124 3324
rect 1372 3316 1380 3324
rect 1452 3316 1460 3324
rect 1564 3316 1572 3324
rect 1596 3316 1604 3324
rect 1660 3316 1668 3324
rect 1868 3316 1876 3324
rect 1980 3316 1988 3324
rect 2108 3316 2116 3324
rect 2220 3316 2228 3324
rect 2268 3316 2276 3324
rect 2396 3316 2404 3324
rect 2572 3336 2580 3344
rect 2620 3336 2628 3344
rect 2652 3336 2660 3344
rect 2732 3336 2740 3344
rect 2876 3336 2884 3344
rect 2940 3336 2948 3344
rect 3068 3336 3076 3344
rect 3084 3336 3092 3344
rect 3164 3336 3172 3344
rect 3340 3336 3348 3344
rect 3356 3336 3364 3344
rect 3452 3336 3460 3344
rect 3484 3336 3492 3344
rect 3564 3336 3572 3344
rect 3740 3336 3748 3344
rect 3852 3336 3860 3344
rect 3932 3336 3940 3344
rect 3964 3336 3972 3344
rect 3996 3336 4004 3344
rect 4076 3336 4084 3344
rect 4188 3336 4196 3344
rect 4268 3336 4276 3344
rect 4284 3336 4292 3344
rect 4396 3336 4404 3344
rect 4924 3336 4932 3344
rect 5148 3336 5156 3344
rect 5164 3336 5172 3344
rect 2444 3316 2452 3324
rect 2524 3316 2532 3324
rect 2604 3316 2612 3324
rect 2764 3316 2772 3324
rect 2796 3316 2804 3324
rect 2828 3316 2836 3324
rect 2876 3316 2884 3324
rect 2924 3316 2932 3324
rect 108 3296 116 3304
rect 156 3296 164 3304
rect 252 3296 260 3304
rect 300 3296 308 3304
rect 348 3296 356 3304
rect 444 3296 452 3304
rect 492 3296 500 3304
rect 636 3296 644 3304
rect 844 3296 852 3304
rect 892 3296 900 3304
rect 988 3296 996 3304
rect 1068 3296 1076 3304
rect 1132 3296 1140 3304
rect 1180 3296 1188 3304
rect 1228 3296 1236 3304
rect 1260 3296 1268 3304
rect 1500 3296 1508 3304
rect 1740 3296 1748 3304
rect 1820 3296 1828 3304
rect 2300 3296 2308 3304
rect 2620 3296 2628 3304
rect 2748 3296 2756 3304
rect 3436 3316 3444 3324
rect 3676 3316 3684 3324
rect 3756 3316 3764 3324
rect 3836 3316 3844 3324
rect 3900 3316 3908 3324
rect 4044 3316 4052 3324
rect 4124 3316 4132 3324
rect 4188 3316 4196 3324
rect 4316 3316 4324 3324
rect 4348 3316 4356 3324
rect 4444 3316 4452 3324
rect 4460 3316 4468 3324
rect 4508 3316 4516 3324
rect 4604 3316 4612 3324
rect 4652 3316 4660 3324
rect 4732 3316 4740 3324
rect 4780 3316 4788 3324
rect 4796 3316 4804 3324
rect 4828 3316 4836 3324
rect 4876 3316 4884 3324
rect 4972 3316 4980 3324
rect 5020 3316 5028 3324
rect 5068 3316 5076 3324
rect 3036 3296 3044 3304
rect 3132 3296 3140 3304
rect 3244 3296 3252 3304
rect 3308 3296 3316 3304
rect 3388 3296 3396 3304
rect 3484 3296 3492 3304
rect 3532 3296 3540 3304
rect 3612 3296 3620 3304
rect 3804 3296 3812 3304
rect 3980 3296 3988 3304
rect 4028 3296 4036 3304
rect 4172 3296 4180 3304
rect 4300 3296 4308 3304
rect 4668 3296 4676 3304
rect 5180 3296 5188 3304
rect 1452 3276 1460 3284
rect 1596 3276 1604 3284
rect 1692 3276 1700 3284
rect 1948 3276 1956 3284
rect 2076 3276 2084 3284
rect 2172 3276 2180 3284
rect 2492 3276 2500 3284
rect 2524 3276 2532 3284
rect 2988 3276 2996 3284
rect 3116 3276 3124 3284
rect 3852 3276 3860 3284
rect 4316 3276 4324 3284
rect 4652 3276 4660 3284
rect 4892 3276 4900 3284
rect 5052 3276 5060 3284
rect 1196 3256 1204 3264
rect 2044 3256 2052 3264
rect 2124 3256 2132 3264
rect 3292 3256 3300 3264
rect 4652 3256 4660 3264
rect 44 3236 52 3244
rect 204 3236 212 3244
rect 460 3236 468 3244
rect 780 3236 788 3244
rect 828 3236 836 3244
rect 1404 3236 1412 3244
rect 1868 3236 1876 3244
rect 1900 3236 1908 3244
rect 3436 3236 3444 3244
rect 3516 3236 3524 3244
rect 3772 3236 3780 3244
rect 4236 3236 4244 3244
rect 4588 3236 4596 3244
rect 4604 3236 4612 3244
rect 4652 3236 4660 3244
rect 4732 3236 4740 3244
rect 4828 3236 4836 3244
rect 4876 3236 4884 3244
rect 4908 3236 4916 3244
rect 4972 3236 4980 3244
rect 5020 3236 5028 3244
rect 5036 3236 5044 3244
rect 5116 3236 5124 3244
rect 796 3176 804 3184
rect 1308 3176 1316 3184
rect 1356 3176 1364 3184
rect 2076 3176 2084 3184
rect 2732 3176 2740 3184
rect 3036 3176 3044 3184
rect 3132 3176 3140 3184
rect 3836 3176 3844 3184
rect 4524 3176 4532 3184
rect 4556 3176 4564 3184
rect 524 3156 532 3164
rect 956 3156 964 3164
rect 2316 3156 2324 3164
rect 2924 3156 2932 3164
rect 3788 3156 3796 3164
rect 1084 3136 1092 3144
rect 1500 3136 1508 3144
rect 2588 3136 2596 3144
rect 2620 3136 2628 3144
rect 2988 3136 2996 3144
rect 3244 3136 3252 3144
rect 3452 3136 3460 3144
rect 3596 3136 3604 3144
rect 3772 3136 3780 3144
rect 4012 3136 4020 3144
rect 4316 3136 4324 3144
rect 4364 3136 4372 3144
rect 188 3116 196 3124
rect 732 3116 740 3124
rect 908 3116 916 3124
rect 1020 3116 1028 3124
rect 1068 3116 1076 3124
rect 1164 3116 1172 3124
rect 1260 3116 1268 3124
rect 12 3096 20 3104
rect 156 3096 164 3104
rect 172 3096 180 3104
rect 348 3096 356 3104
rect 364 3096 372 3104
rect 396 3096 404 3104
rect 412 3096 420 3104
rect 604 3096 612 3104
rect 780 3096 788 3104
rect 876 3096 884 3104
rect 892 3096 900 3104
rect 1100 3096 1108 3104
rect 1148 3096 1156 3104
rect 1308 3096 1316 3104
rect 1356 3096 1364 3104
rect 1436 3096 1444 3104
rect 1452 3096 1460 3104
rect 1660 3116 1668 3124
rect 1580 3096 1588 3104
rect 1628 3096 1636 3104
rect 1644 3096 1652 3104
rect 1676 3096 1684 3104
rect 1724 3096 1732 3104
rect 1804 3096 1812 3104
rect 1836 3096 1844 3104
rect 1932 3096 1940 3104
rect 1964 3096 1972 3104
rect 1980 3096 1988 3104
rect 2012 3096 2020 3104
rect 2108 3096 2116 3104
rect 2172 3096 2180 3104
rect 2300 3116 2308 3124
rect 2492 3116 2500 3124
rect 2716 3116 2724 3124
rect 2796 3116 2804 3124
rect 3084 3116 3092 3124
rect 3164 3116 3172 3124
rect 3308 3116 3316 3124
rect 3532 3116 3540 3124
rect 3692 3116 3700 3124
rect 4044 3116 4052 3124
rect 4300 3116 4308 3124
rect 4396 3116 4404 3124
rect 2236 3096 2244 3104
rect 2284 3096 2292 3104
rect 2332 3096 2340 3104
rect 2396 3096 2404 3104
rect 2412 3096 2420 3104
rect 2476 3096 2484 3104
rect 2636 3096 2644 3104
rect 2844 3096 2852 3104
rect 2908 3096 2916 3104
rect 2940 3096 2948 3104
rect 3020 3096 3028 3104
rect 3292 3096 3300 3104
rect 3356 3096 3364 3104
rect 3388 3096 3396 3104
rect 3404 3096 3412 3104
rect 3452 3096 3460 3104
rect 3580 3096 3588 3104
rect 3644 3096 3652 3104
rect 3788 3096 3796 3104
rect 3948 3096 3956 3104
rect 4028 3096 4036 3104
rect 4076 3096 4084 3104
rect 4140 3096 4148 3104
rect 4220 3096 4228 3104
rect 4252 3096 4260 3104
rect 4396 3096 4404 3104
rect 4444 3096 4452 3104
rect 4508 3096 4516 3104
rect 4556 3096 4564 3104
rect 4636 3096 4644 3104
rect 4732 3096 4740 3104
rect 4748 3096 4756 3104
rect 4796 3096 4804 3104
rect 4844 3096 4852 3104
rect 4924 3096 4932 3104
rect 4940 3096 4948 3104
rect 4972 3096 4980 3104
rect 5020 3096 5028 3104
rect 5132 3096 5140 3104
rect 5164 3096 5172 3104
rect 236 3076 244 3084
rect 268 3076 276 3084
rect 364 3076 372 3084
rect 588 3076 596 3084
rect 764 3076 772 3084
rect 940 3076 948 3084
rect 988 3076 996 3084
rect 1036 3076 1044 3084
rect 1196 3076 1204 3084
rect 1244 3076 1252 3084
rect 1292 3076 1300 3084
rect 1500 3076 1508 3084
rect 1772 3076 1780 3084
rect 2028 3076 2036 3084
rect 2252 3076 2260 3084
rect 2428 3076 2436 3084
rect 2524 3076 2532 3084
rect 2540 3076 2548 3084
rect 2620 3076 2628 3084
rect 2684 3076 2692 3084
rect 2764 3076 2772 3084
rect 2956 3076 2964 3084
rect 3036 3076 3044 3084
rect 3116 3076 3124 3084
rect 3196 3076 3204 3084
rect 3212 3076 3220 3084
rect 3340 3076 3348 3084
rect 3356 3076 3364 3084
rect 3500 3076 3508 3084
rect 3628 3076 3636 3084
rect 3692 3076 3700 3084
rect 3724 3076 3732 3084
rect 3740 3076 3748 3084
rect 12 3056 20 3064
rect 44 3056 52 3064
rect 60 3056 68 3064
rect 140 3056 148 3064
rect 236 3056 244 3064
rect 300 3056 308 3064
rect 316 3056 324 3064
rect 396 3056 404 3064
rect 460 3056 468 3064
rect 492 3056 500 3064
rect 540 3056 548 3064
rect 556 3056 564 3064
rect 604 3056 612 3064
rect 652 3056 660 3064
rect 716 3056 724 3064
rect 732 3056 740 3064
rect 812 3056 820 3064
rect 828 3056 836 3064
rect 972 3056 980 3064
rect 1100 3056 1108 3064
rect 1116 3056 1124 3064
rect 1340 3056 1348 3064
rect 1388 3056 1396 3064
rect 1404 3056 1412 3064
rect 1484 3056 1492 3064
rect 1548 3056 1556 3064
rect 1596 3056 1604 3064
rect 1644 3056 1652 3064
rect 1692 3056 1700 3064
rect 1724 3056 1732 3064
rect 1756 3056 1764 3064
rect 1772 3056 1780 3064
rect 1804 3056 1812 3064
rect 1836 3056 1844 3064
rect 1852 3056 1860 3064
rect 1884 3056 1892 3064
rect 1916 3056 1924 3064
rect 1964 3056 1972 3064
rect 2060 3056 2068 3064
rect 2092 3056 2100 3064
rect 2140 3056 2148 3064
rect 2204 3056 2212 3064
rect 2380 3056 2388 3064
rect 2444 3056 2452 3064
rect 2668 3056 2676 3064
rect 2748 3056 2756 3064
rect 2796 3056 2804 3064
rect 2812 3056 2820 3064
rect 2972 3056 2980 3064
rect 3068 3056 3076 3064
rect 3260 3056 3268 3064
rect 3276 3056 3284 3064
rect 3388 3056 3396 3064
rect 3420 3056 3428 3064
rect 3436 3056 3444 3064
rect 3484 3056 3492 3064
rect 3532 3056 3540 3064
rect 3548 3056 3556 3064
rect 3564 3056 3572 3064
rect 3676 3056 3684 3064
rect 3820 3056 3828 3064
rect 3868 3056 3876 3064
rect 3980 3056 3988 3064
rect 3996 3056 4004 3064
rect 4060 3056 4068 3064
rect 4108 3056 4116 3064
rect 4428 3076 4436 3084
rect 4684 3076 4692 3084
rect 4172 3056 4180 3064
rect 4220 3056 4228 3064
rect 4332 3056 4340 3064
rect 4348 3056 4356 3064
rect 4460 3056 4468 3064
rect 4476 3056 4484 3064
rect 4556 3056 4564 3064
rect 4588 3056 4596 3064
rect 4604 3056 4612 3064
rect 4700 3056 4708 3064
rect 4732 3056 4740 3064
rect 4780 3056 4788 3064
rect 4828 3056 4836 3064
rect 4876 3056 4884 3064
rect 4892 3056 4900 3064
rect 4940 3056 4948 3064
rect 4988 3056 4996 3064
rect 5020 3056 5028 3064
rect 5068 3056 5076 3064
rect 5084 3056 5092 3064
rect 5116 3056 5124 3064
rect 5196 3056 5204 3064
rect 108 3036 116 3044
rect 204 3036 212 3044
rect 572 3036 580 3044
rect 668 3036 676 3044
rect 924 3036 932 3044
rect 1020 3036 1028 3044
rect 1068 3036 1076 3044
rect 1420 3036 1428 3044
rect 1468 3036 1476 3044
rect 1612 3036 1620 3044
rect 2492 3036 2500 3044
rect 2572 3036 2580 3044
rect 2588 3036 2596 3044
rect 2716 3036 2724 3044
rect 2988 3036 2996 3044
rect 3084 3036 3092 3044
rect 3228 3036 3236 3044
rect 3324 3036 3332 3044
rect 3596 3036 3604 3044
rect 3692 3036 3700 3044
rect 3772 3036 3780 3044
rect 4300 3036 4308 3044
rect 4412 3036 4420 3044
rect 4492 3036 4500 3044
rect 4652 3036 4660 3044
rect 4716 3036 4724 3044
rect 4812 3036 4820 3044
rect 4908 3036 4916 3044
rect 5052 3036 5060 3044
rect 5100 3036 5108 3044
rect 76 2976 84 2984
rect 284 2976 292 2984
rect 380 2976 388 2984
rect 508 2976 516 2984
rect 668 2976 676 2984
rect 1004 2976 1012 2984
rect 1084 2976 1092 2984
rect 1452 2976 1460 2984
rect 1708 2976 1716 2984
rect 2268 2976 2276 2984
rect 2508 2976 2516 2984
rect 2556 2976 2564 2984
rect 2748 2976 2756 2984
rect 2924 2976 2932 2984
rect 3212 2976 3220 2984
rect 3452 2976 3460 2984
rect 3484 2976 3492 2984
rect 3564 2976 3572 2984
rect 3788 2976 3796 2984
rect 4044 2976 4052 2984
rect 4124 2976 4132 2984
rect 4188 2976 4196 2984
rect 4284 2976 4292 2984
rect 4396 2976 4404 2984
rect 4460 2976 4468 2984
rect 4572 2976 4580 2984
rect 44 2956 52 2964
rect 156 2956 164 2964
rect 172 2956 180 2964
rect 204 2956 212 2964
rect 316 2956 324 2964
rect 332 2956 340 2964
rect 396 2956 404 2964
rect 444 2956 452 2964
rect 556 2956 564 2964
rect 140 2936 148 2944
rect 252 2936 260 2944
rect 348 2936 356 2944
rect 476 2936 484 2944
rect 652 2956 660 2964
rect 764 2956 772 2964
rect 844 2956 852 2964
rect 892 2956 900 2964
rect 940 2956 948 2964
rect 988 2956 996 2964
rect 1020 2956 1028 2964
rect 1132 2956 1140 2964
rect 1148 2956 1156 2964
rect 1196 2956 1204 2964
rect 1292 2956 1300 2964
rect 1324 2956 1332 2964
rect 1420 2956 1428 2964
rect 1436 2956 1444 2964
rect 1468 2956 1476 2964
rect 1532 2956 1540 2964
rect 1596 2956 1604 2964
rect 1676 2956 1684 2964
rect 1884 2956 1892 2964
rect 1964 2956 1972 2964
rect 12 2916 20 2924
rect 44 2916 52 2924
rect 236 2916 244 2924
rect 284 2916 292 2924
rect 428 2916 436 2924
rect 524 2916 532 2924
rect 604 2916 612 2924
rect 700 2936 708 2944
rect 764 2936 772 2944
rect 828 2936 836 2944
rect 940 2936 948 2944
rect 1324 2936 1332 2944
rect 1724 2936 1732 2944
rect 1740 2936 1748 2944
rect 1772 2936 1780 2944
rect 1820 2936 1828 2944
rect 1836 2936 1844 2944
rect 2028 2956 2036 2964
rect 2204 2956 2212 2964
rect 2236 2956 2244 2964
rect 2252 2956 2260 2964
rect 2316 2956 2324 2964
rect 2076 2936 2084 2944
rect 2252 2936 2260 2944
rect 700 2916 708 2924
rect 812 2916 820 2924
rect 876 2916 884 2924
rect 924 2916 932 2924
rect 940 2916 948 2924
rect 972 2916 980 2924
rect 1068 2916 1076 2924
rect 1180 2916 1188 2924
rect 1244 2916 1252 2924
rect 1292 2916 1300 2924
rect 1340 2916 1348 2924
rect 1372 2916 1380 2924
rect 1468 2916 1476 2924
rect 1500 2916 1508 2924
rect 1596 2916 1604 2924
rect 1628 2916 1636 2924
rect 1644 2916 1652 2924
rect 108 2896 116 2904
rect 284 2896 292 2904
rect 412 2896 420 2904
rect 476 2896 484 2904
rect 508 2896 516 2904
rect 668 2896 676 2904
rect 796 2896 804 2904
rect 860 2896 868 2904
rect 1916 2916 1924 2924
rect 1932 2916 1940 2924
rect 2012 2916 2020 2924
rect 2060 2916 2068 2924
rect 2156 2916 2164 2924
rect 2204 2916 2212 2924
rect 2284 2916 2292 2924
rect 2300 2916 2308 2924
rect 2348 2956 2356 2964
rect 2380 2956 2388 2964
rect 2476 2956 2484 2964
rect 2492 2956 2500 2964
rect 2620 2956 2628 2964
rect 2716 2956 2724 2964
rect 2732 2956 2740 2964
rect 2812 2956 2820 2964
rect 2348 2916 2356 2924
rect 2396 2936 2404 2944
rect 2524 2936 2532 2944
rect 2572 2936 2580 2944
rect 2620 2936 2628 2944
rect 2668 2936 2676 2944
rect 2844 2956 2852 2964
rect 2892 2956 2900 2964
rect 2940 2956 2948 2964
rect 2956 2956 2964 2964
rect 3132 2956 3140 2964
rect 3292 2956 3300 2964
rect 3388 2956 3396 2964
rect 3500 2956 3508 2964
rect 3516 2956 3524 2964
rect 3804 2956 3812 2964
rect 3884 2956 3892 2964
rect 3900 2956 3908 2964
rect 3948 2956 3956 2964
rect 4172 2956 4180 2964
rect 3036 2936 3044 2944
rect 3148 2936 3156 2944
rect 3180 2936 3188 2944
rect 3228 2936 3236 2944
rect 3340 2936 3348 2944
rect 3436 2936 3444 2944
rect 3596 2936 3604 2944
rect 2396 2916 2404 2924
rect 2428 2916 2436 2924
rect 2444 2916 2452 2924
rect 2540 2916 2548 2924
rect 2668 2916 2676 2924
rect 2764 2916 2772 2924
rect 2780 2916 2788 2924
rect 2892 2916 2900 2924
rect 2988 2916 2996 2924
rect 3036 2916 3044 2924
rect 3084 2916 3092 2924
rect 3100 2916 3108 2924
rect 3148 2916 3156 2924
rect 3324 2916 3332 2924
rect 3420 2916 3428 2924
rect 3532 2916 3540 2924
rect 3548 2916 3556 2924
rect 3628 2916 3636 2924
rect 3660 2936 3668 2944
rect 3708 2936 3716 2944
rect 3932 2936 3940 2944
rect 4044 2936 4052 2944
rect 4076 2936 4084 2944
rect 4092 2936 4100 2944
rect 4220 2956 4228 2964
rect 4268 2956 4276 2964
rect 4332 2956 4340 2964
rect 4348 2956 4356 2964
rect 4492 2956 4500 2964
rect 4524 2956 4532 2964
rect 4668 2956 4676 2964
rect 4716 2956 4724 2964
rect 4796 2956 4804 2964
rect 4908 2956 4916 2964
rect 4956 2956 4964 2964
rect 5036 2956 5044 2964
rect 5052 2956 5060 2964
rect 4428 2936 4436 2944
rect 4492 2936 4500 2944
rect 4620 2936 4628 2944
rect 4652 2936 4660 2944
rect 3836 2916 3844 2924
rect 3852 2916 3860 2924
rect 3868 2916 3876 2924
rect 3996 2916 4004 2924
rect 4140 2916 4148 2924
rect 4252 2916 4260 2924
rect 4300 2916 4308 2924
rect 4364 2916 4372 2924
rect 4380 2916 4388 2924
rect 4556 2916 4564 2924
rect 4652 2916 4660 2924
rect 4700 2916 4708 2924
rect 4748 2916 4756 2924
rect 4764 2916 4772 2924
rect 4860 2936 4868 2944
rect 5100 2936 5108 2944
rect 5180 2936 5188 2944
rect 1868 2896 1876 2904
rect 2108 2896 2116 2904
rect 2572 2896 2580 2904
rect 2620 2896 2628 2904
rect 2636 2896 2644 2904
rect 3020 2896 3028 2904
rect 3052 2896 3060 2904
rect 3180 2896 3188 2904
rect 3228 2896 3236 2904
rect 3244 2896 3252 2904
rect 3372 2896 3380 2904
rect 3468 2896 3476 2904
rect 3564 2896 3572 2904
rect 3612 2896 3620 2904
rect 3692 2896 3700 2904
rect 3740 2896 3748 2904
rect 3788 2896 3796 2904
rect 4124 2896 4132 2904
rect 4156 2896 4164 2904
rect 4732 2896 4740 2904
rect 4812 2896 4820 2904
rect 4940 2916 4948 2924
rect 4956 2916 4964 2924
rect 5004 2916 5012 2924
rect 5084 2916 5092 2924
rect 5068 2896 5076 2904
rect 5132 2896 5140 2904
rect 380 2876 388 2884
rect 716 2876 724 2884
rect 972 2876 980 2884
rect 1404 2876 1412 2884
rect 1628 2876 1636 2884
rect 1772 2876 1780 2884
rect 1788 2876 1796 2884
rect 1916 2876 1924 2884
rect 1996 2876 2004 2884
rect 2060 2876 2068 2884
rect 2380 2876 2388 2884
rect 3004 2876 3012 2884
rect 3900 2876 3908 2884
rect 4396 2876 4404 2884
rect 4444 2876 4452 2884
rect 4620 2876 4628 2884
rect 4652 2876 4660 2884
rect 5148 2876 5156 2884
rect 780 2856 788 2864
rect 1276 2856 1284 2864
rect 1756 2856 1764 2864
rect 3420 2856 3428 2864
rect 12 2836 20 2844
rect 268 2836 276 2844
rect 300 2836 308 2844
rect 460 2836 468 2844
rect 636 2836 644 2844
rect 684 2836 692 2844
rect 1004 2836 1012 2844
rect 1180 2836 1188 2844
rect 1324 2836 1332 2844
rect 2444 2836 2452 2844
rect 2684 2836 2692 2844
rect 2988 2836 2996 2844
rect 3164 2836 3172 2844
rect 3356 2836 3364 2844
rect 3836 2836 3844 2844
rect 4316 2836 4324 2844
rect 4508 2836 4516 2844
rect 4780 2836 4788 2844
rect 4828 2836 4836 2844
rect 5004 2836 5012 2844
rect 5116 2836 5124 2844
rect 5164 2836 5172 2844
rect 28 2776 36 2784
rect 556 2776 564 2784
rect 1228 2776 1236 2784
rect 1516 2776 1524 2784
rect 1724 2776 1732 2784
rect 1836 2776 1844 2784
rect 1916 2776 1924 2784
rect 2076 2776 2084 2784
rect 2300 2776 2308 2784
rect 2956 2776 2964 2784
rect 3036 2776 3044 2784
rect 3084 2776 3092 2784
rect 3276 2776 3284 2784
rect 3644 2776 3652 2784
rect 4188 2756 4196 2764
rect 4396 2756 4404 2764
rect 492 2736 500 2744
rect 572 2736 580 2744
rect 764 2736 772 2744
rect 1260 2736 1268 2744
rect 1452 2736 1460 2744
rect 1788 2736 1796 2744
rect 1900 2736 1908 2744
rect 2092 2736 2100 2744
rect 2140 2736 2148 2744
rect 2316 2736 2324 2744
rect 2588 2736 2596 2744
rect 2716 2736 2724 2744
rect 2796 2736 2804 2744
rect 2940 2736 2948 2744
rect 4348 2736 4356 2744
rect 4764 2736 4772 2744
rect 4812 2736 4820 2744
rect 4908 2736 4916 2744
rect 5148 2736 5156 2744
rect 5164 2736 5172 2744
rect 44 2716 52 2724
rect 108 2716 116 2724
rect 140 2716 148 2724
rect 236 2716 244 2724
rect 700 2716 708 2724
rect 156 2696 164 2704
rect 188 2696 196 2704
rect 284 2696 292 2704
rect 300 2696 308 2704
rect 396 2696 404 2704
rect 476 2696 484 2704
rect 556 2696 564 2704
rect 652 2696 660 2704
rect 844 2716 852 2724
rect 908 2716 916 2724
rect 988 2716 996 2724
rect 1084 2716 1092 2724
rect 1356 2716 1364 2724
rect 1596 2716 1604 2724
rect 1132 2696 1140 2704
rect 1196 2696 1204 2704
rect 1228 2696 1236 2704
rect 1276 2696 1284 2704
rect 1324 2696 1332 2704
rect 1404 2696 1412 2704
rect 1500 2696 1508 2704
rect 1516 2696 1524 2704
rect 1612 2696 1620 2704
rect 1996 2716 2004 2724
rect 2188 2716 2196 2724
rect 2268 2716 2276 2724
rect 2508 2716 2516 2724
rect 2748 2716 2756 2724
rect 3100 2716 3108 2724
rect 3116 2716 3124 2724
rect 3196 2716 3204 2724
rect 3212 2716 3220 2724
rect 3260 2716 3268 2724
rect 3308 2716 3316 2724
rect 3356 2716 3364 2724
rect 3388 2716 3396 2724
rect 3516 2716 3524 2724
rect 3548 2716 3556 2724
rect 3660 2716 3668 2724
rect 1708 2696 1716 2704
rect 1740 2696 1748 2704
rect 1900 2696 1908 2704
rect 1948 2696 1956 2704
rect 2156 2696 2164 2704
rect 2236 2696 2244 2704
rect 2540 2696 2548 2704
rect 2700 2696 2708 2704
rect 2844 2696 2852 2704
rect 2860 2696 2868 2704
rect 2892 2696 2900 2704
rect 2940 2696 2948 2704
rect 3356 2696 3364 2704
rect 3484 2696 3492 2704
rect 3532 2696 3540 2704
rect 3612 2696 3620 2704
rect 3916 2716 3924 2724
rect 3964 2716 3972 2724
rect 4060 2716 4068 2724
rect 4092 2716 4100 2724
rect 4124 2716 4132 2724
rect 4300 2716 4308 2724
rect 4444 2716 4452 2724
rect 4492 2716 4500 2724
rect 12 2676 20 2684
rect 44 2676 52 2684
rect 108 2676 116 2684
rect 204 2676 212 2684
rect 652 2676 660 2684
rect 700 2676 708 2684
rect 796 2676 804 2684
rect 812 2676 820 2684
rect 940 2676 948 2684
rect 956 2676 964 2684
rect 1036 2676 1044 2684
rect 1052 2676 1060 2684
rect 1148 2676 1156 2684
rect 1324 2676 1332 2684
rect 1564 2676 1572 2684
rect 1692 2676 1700 2684
rect 2108 2676 2116 2684
rect 2156 2676 2164 2684
rect 2204 2676 2212 2684
rect 2316 2676 2324 2684
rect 2380 2676 2388 2684
rect 2492 2676 2500 2684
rect 2620 2676 2628 2684
rect 156 2656 164 2664
rect 252 2656 260 2664
rect 300 2656 308 2664
rect 332 2656 340 2664
rect 348 2656 356 2664
rect 428 2656 436 2664
rect 508 2656 516 2664
rect 524 2656 532 2664
rect 620 2656 628 2664
rect 876 2656 884 2664
rect 892 2656 900 2664
rect 1100 2656 1108 2664
rect 1148 2656 1156 2664
rect 1180 2656 1188 2664
rect 1260 2656 1268 2664
rect 1308 2656 1316 2664
rect 1372 2656 1380 2664
rect 1468 2656 1476 2664
rect 1548 2656 1556 2664
rect 1644 2656 1652 2664
rect 1740 2656 1748 2664
rect 1772 2656 1780 2664
rect 1820 2656 1828 2664
rect 1852 2656 1860 2664
rect 1868 2656 1876 2664
rect 1932 2656 1940 2664
rect 1980 2656 1988 2664
rect 2060 2656 2068 2664
rect 2092 2656 2100 2664
rect 2268 2656 2276 2664
rect 2412 2656 2420 2664
rect 2428 2656 2436 2664
rect 2492 2656 2500 2664
rect 2652 2656 2660 2664
rect 2700 2676 2708 2684
rect 2764 2676 2772 2684
rect 2796 2676 2804 2684
rect 3068 2676 3076 2684
rect 3148 2676 3156 2684
rect 3164 2676 3172 2684
rect 3244 2676 3252 2684
rect 3292 2676 3300 2684
rect 3388 2676 3396 2684
rect 2684 2656 2692 2664
rect 2892 2656 2900 2664
rect 2908 2656 2916 2664
rect 2972 2656 2980 2664
rect 3004 2656 3012 2664
rect 3052 2656 3060 2664
rect 3212 2656 3220 2664
rect 3468 2676 3476 2684
rect 3628 2676 3636 2684
rect 3708 2676 3716 2684
rect 3884 2696 3892 2704
rect 4012 2696 4020 2704
rect 4060 2696 4068 2704
rect 4204 2696 4212 2704
rect 4284 2696 4292 2704
rect 4380 2696 4388 2704
rect 4540 2696 4548 2704
rect 4668 2696 4676 2704
rect 4716 2696 4724 2704
rect 4764 2696 4772 2704
rect 4860 2696 4868 2704
rect 4908 2696 4916 2704
rect 4924 2696 4932 2704
rect 4972 2696 4980 2704
rect 5100 2716 5108 2724
rect 3788 2676 3796 2684
rect 3868 2676 3876 2684
rect 3932 2676 3940 2684
rect 4028 2676 4036 2684
rect 4156 2676 4164 2684
rect 4252 2676 4260 2684
rect 4380 2676 4388 2684
rect 4476 2676 4484 2684
rect 4604 2676 4612 2684
rect 4780 2676 4788 2684
rect 4972 2676 4980 2684
rect 5052 2676 5060 2684
rect 5068 2676 5076 2684
rect 5100 2676 5108 2684
rect 3436 2656 3444 2664
rect 3564 2656 3572 2664
rect 3628 2656 3636 2664
rect 3708 2656 3716 2664
rect 3740 2656 3748 2664
rect 3836 2656 3844 2664
rect 4012 2656 4020 2664
rect 4172 2656 4180 2664
rect 4236 2656 4244 2664
rect 4252 2656 4260 2664
rect 4428 2656 4436 2664
rect 4572 2656 4580 2664
rect 4636 2656 4644 2664
rect 4684 2656 4692 2664
rect 4716 2656 4724 2664
rect 4732 2656 4740 2664
rect 4876 2656 4884 2664
rect 4956 2656 4964 2664
rect 5004 2656 5012 2664
rect 76 2636 84 2644
rect 124 2636 132 2644
rect 268 2636 276 2644
rect 412 2636 420 2644
rect 572 2636 580 2644
rect 700 2636 708 2644
rect 748 2636 756 2644
rect 828 2636 836 2644
rect 1084 2636 1092 2644
rect 1164 2636 1172 2644
rect 1356 2636 1364 2644
rect 1580 2636 1588 2644
rect 1676 2636 1684 2644
rect 1996 2636 2004 2644
rect 2188 2636 2196 2644
rect 2396 2636 2404 2644
rect 3132 2636 3140 2644
rect 3180 2636 3188 2644
rect 3500 2636 3508 2644
rect 3660 2636 3668 2644
rect 3916 2636 3924 2644
rect 4044 2636 4052 2644
rect 4268 2636 4276 2644
rect 4316 2636 4324 2644
rect 4348 2636 4356 2644
rect 4444 2636 4452 2644
rect 4492 2636 4500 2644
rect 4844 2636 4852 2644
rect 5020 2636 5028 2644
rect 5100 2636 5108 2644
rect 140 2576 148 2584
rect 220 2576 228 2584
rect 396 2576 404 2584
rect 476 2576 484 2584
rect 508 2576 516 2584
rect 572 2576 580 2584
rect 956 2576 964 2584
rect 1228 2576 1236 2584
rect 1404 2576 1412 2584
rect 1468 2576 1476 2584
rect 1628 2576 1636 2584
rect 1948 2576 1956 2584
rect 2076 2576 2084 2584
rect 2236 2576 2244 2584
rect 2428 2576 2436 2584
rect 2476 2576 2484 2584
rect 2668 2576 2676 2584
rect 2988 2576 2996 2584
rect 3612 2576 3620 2584
rect 3708 2576 3716 2584
rect 3740 2576 3748 2584
rect 3868 2576 3876 2584
rect 3996 2576 4004 2584
rect 4044 2576 4052 2584
rect 4172 2576 4180 2584
rect 4236 2576 4244 2584
rect 4316 2576 4324 2584
rect 4732 2576 4740 2584
rect 5164 2576 5172 2584
rect 236 2556 244 2564
rect 284 2556 292 2564
rect 12 2536 20 2544
rect 108 2536 116 2544
rect 156 2536 164 2544
rect 364 2556 372 2564
rect 428 2556 436 2564
rect 460 2556 468 2564
rect 492 2556 500 2564
rect 588 2556 596 2564
rect 652 2556 660 2564
rect 732 2556 740 2564
rect 780 2556 788 2564
rect 332 2536 340 2544
rect 540 2536 548 2544
rect 636 2536 644 2544
rect 748 2536 756 2544
rect 780 2536 788 2544
rect 844 2556 852 2564
rect 908 2556 916 2564
rect 988 2556 996 2564
rect 1004 2556 1012 2564
rect 1036 2556 1044 2564
rect 1116 2556 1124 2564
rect 1244 2556 1252 2564
rect 1260 2556 1268 2564
rect 1308 2556 1316 2564
rect 1484 2556 1492 2564
rect 1500 2556 1508 2564
rect 1532 2556 1540 2564
rect 1564 2556 1572 2564
rect 1660 2556 1668 2564
rect 1708 2556 1716 2564
rect 1788 2556 1796 2564
rect 1836 2556 1844 2564
rect 2012 2556 2020 2564
rect 2028 2556 2036 2564
rect 2044 2556 2052 2564
rect 2124 2556 2132 2564
rect 2172 2556 2180 2564
rect 2252 2556 2260 2564
rect 2268 2556 2276 2564
rect 2316 2556 2324 2564
rect 2348 2556 2356 2564
rect 2508 2556 2516 2564
rect 2588 2556 2596 2564
rect 2620 2556 2628 2564
rect 2684 2556 2692 2564
rect 2716 2556 2724 2564
rect 2732 2556 2740 2564
rect 2780 2556 2788 2564
rect 2796 2556 2804 2564
rect 2828 2556 2836 2564
rect 2876 2556 2884 2564
rect 2908 2556 2916 2564
rect 2940 2556 2948 2564
rect 2956 2556 2964 2564
rect 3020 2556 3028 2564
rect 3068 2556 3076 2564
rect 924 2536 932 2544
rect 1164 2536 1172 2544
rect 1196 2536 1204 2544
rect 1276 2536 1284 2544
rect 1356 2536 1364 2544
rect 1404 2536 1412 2544
rect 1436 2536 1444 2544
rect 1964 2536 1972 2544
rect 2108 2536 2116 2544
rect 2364 2536 2372 2544
rect 2396 2536 2404 2544
rect 2444 2536 2452 2544
rect 2508 2536 2516 2544
rect 2588 2536 2596 2544
rect 2636 2536 2644 2544
rect 2716 2536 2724 2544
rect 2860 2536 2868 2544
rect 3020 2536 3028 2544
rect 3148 2536 3156 2544
rect 92 2516 100 2524
rect 252 2516 260 2524
rect 332 2516 340 2524
rect 364 2516 372 2524
rect 428 2516 436 2524
rect 460 2516 468 2524
rect 556 2516 564 2524
rect 44 2496 52 2504
rect 140 2496 148 2504
rect 188 2496 196 2504
rect 508 2496 516 2504
rect 684 2516 692 2524
rect 700 2516 708 2524
rect 748 2516 756 2524
rect 780 2516 788 2524
rect 828 2516 836 2524
rect 876 2516 884 2524
rect 1036 2516 1044 2524
rect 1084 2516 1092 2524
rect 1212 2516 1220 2524
rect 1308 2516 1316 2524
rect 1340 2516 1348 2524
rect 1436 2516 1444 2524
rect 1580 2516 1588 2524
rect 1692 2516 1700 2524
rect 1788 2516 1796 2524
rect 1836 2516 1844 2524
rect 1868 2516 1876 2524
rect 956 2496 964 2504
rect 1020 2496 1028 2504
rect 1068 2496 1076 2504
rect 1164 2496 1172 2504
rect 1196 2496 1204 2504
rect 1388 2496 1396 2504
rect 1404 2496 1412 2504
rect 1644 2496 1652 2504
rect 1916 2496 1924 2504
rect 1980 2516 1988 2524
rect 2060 2516 2068 2524
rect 2220 2516 2228 2524
rect 2300 2516 2308 2524
rect 2348 2516 2356 2524
rect 2540 2516 2548 2524
rect 2556 2516 2564 2524
rect 2732 2516 2740 2524
rect 2764 2516 2772 2524
rect 2812 2516 2820 2524
rect 2860 2516 2868 2524
rect 2876 2516 2884 2524
rect 2924 2516 2932 2524
rect 3052 2516 3060 2524
rect 3100 2516 3108 2524
rect 3196 2516 3204 2524
rect 3324 2536 3332 2544
rect 3372 2556 3380 2564
rect 3404 2556 3412 2564
rect 3484 2556 3492 2564
rect 3548 2556 3556 2564
rect 3628 2556 3636 2564
rect 3644 2556 3652 2564
rect 3788 2556 3796 2564
rect 3916 2556 3924 2564
rect 3452 2536 3460 2544
rect 3532 2536 3540 2544
rect 3692 2536 3700 2544
rect 4124 2556 4132 2564
rect 4252 2556 4260 2564
rect 4348 2556 4356 2564
rect 4604 2556 4612 2564
rect 4796 2556 4804 2564
rect 4988 2556 4996 2564
rect 5004 2556 5012 2564
rect 5084 2556 5092 2564
rect 5148 2556 5156 2564
rect 3980 2536 3988 2544
rect 4060 2536 4068 2544
rect 4108 2536 4116 2544
rect 4156 2536 4164 2544
rect 4204 2536 4212 2544
rect 4300 2536 4308 2544
rect 4412 2536 4420 2544
rect 4460 2536 4468 2544
rect 4476 2536 4484 2544
rect 4524 2536 4532 2544
rect 4652 2536 4660 2544
rect 4748 2536 4756 2544
rect 4764 2536 4772 2544
rect 4844 2536 4852 2544
rect 4892 2536 4900 2544
rect 3404 2516 3412 2524
rect 3484 2516 3492 2524
rect 3532 2516 3540 2524
rect 3580 2516 3588 2524
rect 3596 2516 3604 2524
rect 3660 2516 3668 2524
rect 3692 2516 3700 2524
rect 3820 2516 3828 2524
rect 3884 2516 3892 2524
rect 3932 2516 3940 2524
rect 3948 2516 3956 2524
rect 4236 2516 4244 2524
rect 4284 2516 4292 2524
rect 4508 2516 4516 2524
rect 4588 2516 4596 2524
rect 4604 2516 4612 2524
rect 4620 2516 4628 2524
rect 4940 2536 4948 2544
rect 5132 2536 5140 2544
rect 4956 2516 4964 2524
rect 5036 2516 5044 2524
rect 5052 2516 5060 2524
rect 5180 2516 5188 2524
rect 1996 2496 2004 2504
rect 2076 2496 2084 2504
rect 2124 2496 2132 2504
rect 2284 2496 2292 2504
rect 2364 2496 2372 2504
rect 2412 2496 2420 2504
rect 2668 2496 2676 2504
rect 2972 2496 2980 2504
rect 3084 2496 3092 2504
rect 3116 2496 3124 2504
rect 3148 2496 3156 2504
rect 3228 2496 3236 2504
rect 3292 2496 3300 2504
rect 3468 2496 3476 2504
rect 3500 2496 3508 2504
rect 3724 2496 3732 2504
rect 3740 2496 3748 2504
rect 4012 2496 4020 2504
rect 4028 2496 4036 2504
rect 4076 2496 4084 2504
rect 4140 2496 4148 2504
rect 4236 2496 4244 2504
rect 4332 2496 4340 2504
rect 4476 2496 4484 2504
rect 4508 2496 4516 2504
rect 4700 2496 4708 2504
rect 4716 2496 4724 2504
rect 4748 2496 4756 2504
rect 4796 2496 4804 2504
rect 4860 2496 4868 2504
rect 4940 2496 4948 2504
rect 5100 2496 5108 2504
rect 156 2476 164 2484
rect 748 2476 756 2484
rect 860 2476 868 2484
rect 1692 2476 1700 2484
rect 1820 2476 1828 2484
rect 2444 2476 2452 2484
rect 2540 2476 2548 2484
rect 2636 2476 2644 2484
rect 3052 2476 3060 2484
rect 3420 2476 3428 2484
rect 3868 2476 3876 2484
rect 4188 2476 4196 2484
rect 4396 2476 4404 2484
rect 4556 2476 4564 2484
rect 4812 2476 4820 2484
rect 5052 2476 5060 2484
rect 1564 2456 1572 2464
rect 92 2436 100 2444
rect 348 2436 356 2444
rect 620 2436 628 2444
rect 668 2436 676 2444
rect 892 2436 900 2444
rect 972 2436 980 2444
rect 1100 2436 1108 2444
rect 1324 2436 1332 2444
rect 1516 2436 1524 2444
rect 1756 2436 1764 2444
rect 2428 2436 2436 2444
rect 2604 2436 2612 2444
rect 3132 2436 3140 2444
rect 3340 2436 3348 2444
rect 3884 2436 3892 2444
rect 4092 2436 4100 2444
rect 4828 2436 4836 2444
rect 4924 2436 4932 2444
rect 5036 2436 5044 2444
rect 5116 2436 5124 2444
rect 364 2376 372 2384
rect 1580 2376 1588 2384
rect 1660 2376 1668 2384
rect 1948 2376 1956 2384
rect 2332 2376 2340 2384
rect 2540 2376 2548 2384
rect 2668 2376 2676 2384
rect 2748 2376 2756 2384
rect 3196 2376 3204 2384
rect 3292 2376 3300 2384
rect 4012 2376 4020 2384
rect 4060 2376 4068 2384
rect 4748 2376 4756 2384
rect 2316 2356 2324 2364
rect 4700 2356 4708 2364
rect 572 2336 580 2344
rect 620 2336 628 2344
rect 764 2336 772 2344
rect 1260 2336 1268 2344
rect 1340 2336 1348 2344
rect 1500 2336 1508 2344
rect 1548 2336 1556 2344
rect 2412 2336 2420 2344
rect 3100 2336 3108 2344
rect 3116 2336 3124 2344
rect 3500 2336 3508 2344
rect 3996 2336 4004 2344
rect 4124 2336 4132 2344
rect 4316 2336 4324 2344
rect 4428 2336 4436 2344
rect 4732 2336 4740 2344
rect 4940 2336 4948 2344
rect 556 2316 564 2324
rect 684 2316 692 2324
rect 828 2316 836 2324
rect 1036 2316 1044 2324
rect 1228 2316 1236 2324
rect 1468 2316 1476 2324
rect 1628 2316 1636 2324
rect 1740 2316 1748 2324
rect 1836 2316 1844 2324
rect 1916 2316 1924 2324
rect 1964 2316 1972 2324
rect 2060 2316 2068 2324
rect 2076 2316 2084 2324
rect 2364 2316 2372 2324
rect 2476 2316 2484 2324
rect 2588 2316 2596 2324
rect 2636 2316 2644 2324
rect 2796 2316 2804 2324
rect 2940 2316 2948 2324
rect 2972 2316 2980 2324
rect 12 2296 20 2304
rect 140 2296 148 2304
rect 156 2296 164 2304
rect 284 2296 292 2304
rect 300 2296 308 2304
rect 380 2296 388 2304
rect 428 2296 436 2304
rect 508 2296 516 2304
rect 572 2296 580 2304
rect 700 2296 708 2304
rect 780 2296 788 2304
rect 876 2296 884 2304
rect 908 2296 916 2304
rect 924 2296 932 2304
rect 1004 2296 1012 2304
rect 1020 2296 1028 2304
rect 1052 2296 1060 2304
rect 1164 2296 1172 2304
rect 1212 2296 1220 2304
rect 1340 2296 1348 2304
rect 1356 2296 1364 2304
rect 1404 2296 1412 2304
rect 1596 2296 1604 2304
rect 1612 2296 1620 2304
rect 1676 2296 1684 2304
rect 1724 2296 1732 2304
rect 1788 2296 1796 2304
rect 1836 2296 1844 2304
rect 2124 2296 2132 2304
rect 2188 2296 2196 2304
rect 2236 2296 2244 2304
rect 2316 2296 2324 2304
rect 2412 2296 2420 2304
rect 2460 2296 2468 2304
rect 2652 2296 2660 2304
rect 2780 2296 2788 2304
rect 2796 2296 2804 2304
rect 2844 2296 2852 2304
rect 2876 2296 2884 2304
rect 2988 2296 2996 2304
rect 3020 2296 3028 2304
rect 3036 2296 3044 2304
rect 3132 2296 3140 2304
rect 3148 2296 3156 2304
rect 3228 2296 3236 2304
rect 3356 2316 3364 2324
rect 3404 2316 3412 2324
rect 3628 2316 3636 2324
rect 3724 2316 3732 2324
rect 3420 2296 3428 2304
rect 3452 2296 3460 2304
rect 3500 2296 3508 2304
rect 3532 2296 3540 2304
rect 3548 2296 3556 2304
rect 3740 2296 3748 2304
rect 3916 2316 3924 2324
rect 3964 2316 3972 2324
rect 4188 2316 4196 2324
rect 4252 2316 4260 2324
rect 4636 2316 4644 2324
rect 4684 2316 4692 2324
rect 4796 2316 4804 2324
rect 4956 2316 4964 2324
rect 5036 2316 5044 2324
rect 5052 2316 5060 2324
rect 5180 2316 5188 2324
rect 3868 2296 3876 2304
rect 4076 2296 4084 2304
rect 4140 2296 4148 2304
rect 4236 2296 4244 2304
rect 4844 2296 4852 2304
rect 4860 2296 4868 2304
rect 28 2256 36 2264
rect 60 2276 68 2284
rect 60 2256 68 2264
rect 92 2256 100 2264
rect 108 2256 116 2264
rect 188 2256 196 2264
rect 460 2276 468 2284
rect 508 2276 516 2284
rect 652 2276 660 2284
rect 796 2276 804 2284
rect 860 2276 868 2284
rect 892 2276 900 2284
rect 236 2256 244 2264
rect 300 2256 308 2264
rect 332 2256 340 2264
rect 348 2256 356 2264
rect 460 2256 468 2264
rect 476 2256 484 2264
rect 604 2256 612 2264
rect 636 2256 644 2264
rect 748 2256 756 2264
rect 780 2256 788 2264
rect 844 2256 852 2264
rect 876 2256 884 2264
rect 892 2256 900 2264
rect 956 2256 964 2264
rect 988 2276 996 2284
rect 1100 2276 1108 2284
rect 1244 2276 1252 2284
rect 1308 2276 1316 2284
rect 1404 2276 1412 2284
rect 1772 2276 1780 2284
rect 1868 2276 1876 2284
rect 1884 2276 1892 2284
rect 1996 2276 2004 2284
rect 2044 2276 2052 2284
rect 2172 2276 2180 2284
rect 2220 2276 2228 2284
rect 2396 2276 2404 2284
rect 2524 2276 2532 2284
rect 2556 2276 2564 2284
rect 2604 2276 2612 2284
rect 1068 2256 1076 2264
rect 1100 2256 1108 2264
rect 1196 2256 1204 2264
rect 1244 2256 1252 2264
rect 1308 2256 1316 2264
rect 1468 2256 1476 2264
rect 1516 2256 1524 2264
rect 1532 2256 1540 2264
rect 1564 2256 1572 2264
rect 1644 2256 1652 2264
rect 1676 2256 1684 2264
rect 1724 2256 1732 2264
rect 1788 2256 1796 2264
rect 1804 2256 1812 2264
rect 1932 2256 1940 2264
rect 2028 2256 2036 2264
rect 2092 2256 2100 2264
rect 2124 2256 2132 2264
rect 2220 2256 2228 2264
rect 2268 2256 2276 2264
rect 2284 2256 2292 2264
rect 2348 2256 2356 2264
rect 2444 2256 2452 2264
rect 2492 2256 2500 2264
rect 2508 2256 2516 2264
rect 2556 2256 2564 2264
rect 2588 2256 2596 2264
rect 2732 2276 2740 2284
rect 2764 2276 2772 2284
rect 2860 2276 2868 2284
rect 2908 2276 2916 2284
rect 3084 2276 3092 2284
rect 3308 2276 3316 2284
rect 3324 2276 3332 2284
rect 3372 2276 3380 2284
rect 3596 2276 3604 2284
rect 3692 2276 3700 2284
rect 3836 2276 3844 2284
rect 3932 2276 3940 2284
rect 4156 2276 4164 2284
rect 4220 2276 4228 2284
rect 4268 2276 4276 2284
rect 4508 2276 4516 2284
rect 4588 2276 4596 2284
rect 4604 2276 4612 2284
rect 4652 2276 4660 2284
rect 2732 2256 2740 2264
rect 2844 2256 2852 2264
rect 2956 2256 2964 2264
rect 3004 2256 3012 2264
rect 3036 2256 3044 2264
rect 3116 2256 3124 2264
rect 3164 2256 3172 2264
rect 3260 2256 3268 2264
rect 3420 2256 3428 2264
rect 3468 2256 3476 2264
rect 3580 2256 3588 2264
rect 3772 2256 3780 2264
rect 3788 2256 3796 2264
rect 3836 2256 3844 2264
rect 3948 2256 3956 2264
rect 3980 2256 3988 2264
rect 4028 2256 4036 2264
rect 4044 2256 4052 2264
rect 4092 2256 4100 2264
rect 4172 2256 4180 2264
rect 4268 2256 4276 2264
rect 4396 2256 4404 2264
rect 4412 2256 4420 2264
rect 4444 2256 4452 2264
rect 4476 2256 4484 2264
rect 4524 2256 4532 2264
rect 4556 2256 4564 2264
rect 4732 2276 4740 2284
rect 4764 2276 4772 2284
rect 4828 2276 4836 2284
rect 4892 2276 4900 2284
rect 4908 2276 4916 2284
rect 4988 2276 4996 2284
rect 5004 2276 5012 2284
rect 5084 2276 5092 2284
rect 5100 2276 5108 2284
rect 5148 2276 5156 2284
rect 4780 2256 4788 2264
rect 4812 2256 4820 2264
rect 4860 2256 4868 2264
rect 4892 2256 4900 2264
rect 4924 2256 4932 2264
rect 220 2236 228 2244
rect 396 2236 404 2244
rect 556 2236 564 2244
rect 668 2236 676 2244
rect 828 2236 836 2244
rect 1836 2236 1844 2244
rect 1900 2236 1908 2244
rect 1980 2236 1988 2244
rect 2012 2236 2020 2244
rect 2204 2236 2212 2244
rect 2380 2236 2388 2244
rect 3356 2236 3364 2244
rect 3404 2236 3412 2244
rect 3660 2236 3668 2244
rect 3916 2236 3924 2244
rect 4204 2236 4212 2244
rect 4364 2236 4372 2244
rect 4636 2236 4644 2244
rect 4668 2236 4676 2244
rect 4972 2236 4980 2244
rect 5036 2236 5044 2244
rect 5068 2236 5076 2244
rect 5132 2236 5140 2244
rect 284 2176 292 2184
rect 348 2176 356 2184
rect 540 2176 548 2184
rect 684 2176 692 2184
rect 780 2176 788 2184
rect 924 2176 932 2184
rect 972 2176 980 2184
rect 1020 2176 1028 2184
rect 1148 2176 1156 2184
rect 1388 2176 1396 2184
rect 1532 2176 1540 2184
rect 1948 2176 1956 2184
rect 2220 2176 2228 2184
rect 2364 2176 2372 2184
rect 2412 2176 2420 2184
rect 2492 2176 2500 2184
rect 2620 2176 2628 2184
rect 2828 2176 2836 2184
rect 2892 2176 2900 2184
rect 3068 2176 3076 2184
rect 3148 2176 3156 2184
rect 3212 2176 3220 2184
rect 3324 2176 3332 2184
rect 3356 2176 3364 2184
rect 3436 2176 3444 2184
rect 3484 2176 3492 2184
rect 3756 2176 3764 2184
rect 4092 2176 4100 2184
rect 4188 2176 4196 2184
rect 4220 2176 4228 2184
rect 4300 2176 4308 2184
rect 4476 2176 4484 2184
rect 4588 2176 4596 2184
rect 4620 2176 4628 2184
rect 4876 2176 4884 2184
rect 5052 2176 5060 2184
rect 44 2156 52 2164
rect 60 2156 68 2164
rect 108 2156 116 2164
rect 172 2156 180 2164
rect 188 2156 196 2164
rect 268 2156 276 2164
rect 380 2156 388 2164
rect 460 2156 468 2164
rect 604 2156 612 2164
rect 716 2156 724 2164
rect 796 2156 804 2164
rect 812 2156 820 2164
rect 844 2156 852 2164
rect 892 2156 900 2164
rect 956 2156 964 2164
rect 1164 2156 1172 2164
rect 1228 2156 1236 2164
rect 1292 2156 1300 2164
rect 1324 2156 1332 2164
rect 1340 2156 1348 2164
rect 12 2136 20 2144
rect 12 2116 20 2124
rect 92 2116 100 2124
rect 108 2116 116 2124
rect 220 2116 228 2124
rect 316 2136 324 2144
rect 332 2136 340 2144
rect 412 2136 420 2144
rect 508 2136 516 2144
rect 524 2136 532 2144
rect 620 2136 628 2144
rect 748 2136 756 2144
rect 428 2116 436 2124
rect 444 2116 452 2124
rect 572 2116 580 2124
rect 700 2116 708 2124
rect 748 2116 756 2124
rect 940 2136 948 2144
rect 1036 2136 1044 2144
rect 1132 2136 1140 2144
rect 1212 2136 1220 2144
rect 1308 2136 1316 2144
rect 1356 2136 1364 2144
rect 1420 2156 1428 2164
rect 1596 2156 1604 2164
rect 1660 2156 1668 2164
rect 1692 2156 1700 2164
rect 1756 2156 1764 2164
rect 1788 2156 1796 2164
rect 1852 2156 1860 2164
rect 1884 2156 1892 2164
rect 2028 2156 2036 2164
rect 2060 2156 2068 2164
rect 2108 2156 2116 2164
rect 2156 2156 2164 2164
rect 2172 2156 2180 2164
rect 2284 2156 2292 2164
rect 2444 2156 2452 2164
rect 2508 2156 2516 2164
rect 2556 2156 2564 2164
rect 2572 2156 2580 2164
rect 2700 2156 2708 2164
rect 2716 2156 2724 2164
rect 2812 2156 2820 2164
rect 2972 2156 2980 2164
rect 3132 2156 3140 2164
rect 3228 2156 3236 2164
rect 3244 2156 3252 2164
rect 3276 2156 3284 2164
rect 3340 2156 3348 2164
rect 3404 2156 3412 2164
rect 3420 2156 3428 2164
rect 3564 2156 3572 2164
rect 3852 2156 3860 2164
rect 3884 2156 3892 2164
rect 4028 2156 4036 2164
rect 4108 2156 4116 2164
rect 796 2116 804 2124
rect 844 2116 852 2124
rect 284 2096 292 2104
rect 364 2096 372 2104
rect 380 2096 388 2104
rect 476 2096 484 2104
rect 556 2096 564 2104
rect 588 2096 596 2104
rect 652 2096 660 2104
rect 988 2116 996 2124
rect 1052 2116 1060 2124
rect 1100 2116 1108 2124
rect 1212 2116 1220 2124
rect 1260 2116 1268 2124
rect 1356 2116 1364 2124
rect 1468 2136 1476 2144
rect 1548 2136 1556 2144
rect 1612 2136 1620 2144
rect 1644 2136 1652 2144
rect 1740 2136 1748 2144
rect 1804 2136 1812 2144
rect 1932 2136 1940 2144
rect 1980 2136 1988 2144
rect 2204 2136 2212 2144
rect 2332 2136 2340 2144
rect 2348 2136 2356 2144
rect 4252 2156 4260 2164
rect 4364 2156 4372 2164
rect 4380 2156 4388 2164
rect 4540 2156 4548 2164
rect 4700 2156 4708 2164
rect 4748 2156 4756 2164
rect 4796 2156 4804 2164
rect 4892 2156 4900 2164
rect 4972 2156 4980 2164
rect 5020 2156 5028 2164
rect 5100 2156 5108 2164
rect 2652 2136 2660 2144
rect 2748 2136 2756 2144
rect 2860 2136 2868 2144
rect 2876 2136 2884 2144
rect 2908 2136 2916 2144
rect 2972 2136 2980 2144
rect 3020 2136 3028 2144
rect 3100 2136 3108 2144
rect 3180 2136 3188 2144
rect 3292 2136 3300 2144
rect 3500 2136 3508 2144
rect 3516 2136 3524 2144
rect 3644 2136 3652 2144
rect 3660 2136 3668 2144
rect 3740 2136 3748 2144
rect 3788 2136 3796 2144
rect 3836 2136 3844 2144
rect 3916 2136 3924 2144
rect 3932 2136 3940 2144
rect 3980 2136 3988 2144
rect 4012 2136 4020 2144
rect 4124 2136 4132 2144
rect 4156 2136 4164 2144
rect 4236 2136 4244 2144
rect 4316 2136 4324 2144
rect 4444 2136 4452 2144
rect 4460 2136 4468 2144
rect 4540 2136 4548 2144
rect 4604 2136 4612 2144
rect 4652 2136 4660 2144
rect 4748 2136 4756 2144
rect 4844 2136 4852 2144
rect 4924 2136 4932 2144
rect 5036 2136 5044 2144
rect 5084 2136 5092 2144
rect 5116 2136 5124 2144
rect 1564 2116 1572 2124
rect 1596 2116 1604 2124
rect 1644 2116 1652 2124
rect 1740 2116 1748 2124
rect 1996 2116 2004 2124
rect 2028 2116 2036 2124
rect 2060 2116 2068 2124
rect 2108 2116 2116 2124
rect 2188 2116 2196 2124
rect 2252 2116 2260 2124
rect 2476 2116 2484 2124
rect 2524 2116 2532 2124
rect 2604 2116 2612 2124
rect 2668 2116 2676 2124
rect 3004 2116 3012 2124
rect 3276 2116 3284 2124
rect 3420 2116 3428 2124
rect 3452 2116 3460 2124
rect 3596 2116 3604 2124
rect 3788 2116 3796 2124
rect 4060 2116 4068 2124
rect 4076 2116 4084 2124
rect 4332 2116 4340 2124
rect 4348 2116 4356 2124
rect 4428 2116 4436 2124
rect 4508 2116 4516 2124
rect 4780 2116 4788 2124
rect 4828 2116 4836 2124
rect 4940 2116 4948 2124
rect 4988 2116 4996 2124
rect 1004 2096 1012 2104
rect 1100 2096 1108 2104
rect 1180 2096 1188 2104
rect 1276 2096 1284 2104
rect 1500 2096 1508 2104
rect 1516 2096 1524 2104
rect 1708 2096 1716 2104
rect 1836 2096 1844 2104
rect 1900 2096 1908 2104
rect 2236 2096 2244 2104
rect 2268 2096 2276 2104
rect 2380 2096 2388 2104
rect 2780 2096 2788 2104
rect 2908 2096 2916 2104
rect 3052 2096 3060 2104
rect 3068 2096 3076 2104
rect 3148 2096 3156 2104
rect 3324 2096 3332 2104
rect 3388 2096 3396 2104
rect 3468 2096 3476 2104
rect 3548 2096 3556 2104
rect 3612 2096 3620 2104
rect 3644 2096 3652 2104
rect 3692 2096 3700 2104
rect 3708 2096 3716 2104
rect 3884 2096 3892 2104
rect 3964 2096 3972 2104
rect 3980 2096 3988 2104
rect 4188 2096 4196 2104
rect 4204 2096 4212 2104
rect 4284 2096 4292 2104
rect 4492 2096 4500 2104
rect 4588 2096 4596 2104
rect 4636 2096 4644 2104
rect 4684 2096 4692 2104
rect 4700 2096 4708 2104
rect 4876 2096 4884 2104
rect 5004 2096 5012 2104
rect 5068 2096 5076 2104
rect 5164 2096 5172 2104
rect 940 2076 948 2084
rect 1820 2076 1828 2084
rect 1948 2076 1956 2084
rect 1980 2076 1988 2084
rect 2300 2076 2308 2084
rect 2396 2076 2404 2084
rect 2620 2076 2628 2084
rect 2668 2076 2676 2084
rect 2716 2076 2724 2084
rect 2924 2076 2932 2084
rect 3100 2076 3108 2084
rect 3740 2076 3748 2084
rect 4156 2076 4164 2084
rect 4844 2076 4852 2084
rect 4892 2076 4900 2084
rect 5116 2076 5124 2084
rect 1612 2056 1620 2064
rect 3996 2056 4004 2064
rect 92 2036 100 2044
rect 236 2036 244 2044
rect 492 2036 500 2044
rect 748 2036 756 2044
rect 1196 2036 1204 2044
rect 2076 2036 2084 2044
rect 2140 2036 2148 2044
rect 2524 2036 2532 2044
rect 2764 2036 2772 2044
rect 3036 2036 3044 2044
rect 3532 2036 3540 2044
rect 3596 2036 3604 2044
rect 3628 2036 3636 2044
rect 3724 2036 3732 2044
rect 3868 2036 3876 2044
rect 4060 2036 4068 2044
rect 4268 2036 4276 2044
rect 4508 2036 4516 2044
rect 4668 2036 4676 2044
rect 4780 2036 4788 2044
rect 4940 2036 4948 2044
rect 5148 2036 5156 2044
rect 12 1976 20 1984
rect 428 1976 436 1984
rect 572 1976 580 1984
rect 812 1976 820 1984
rect 844 1976 852 1984
rect 1004 1976 1012 1984
rect 1148 1976 1156 1984
rect 1196 1976 1204 1984
rect 1276 1976 1284 1984
rect 1836 1976 1844 1984
rect 2012 1976 2020 1984
rect 2124 1976 2132 1984
rect 2620 1976 2628 1984
rect 2700 1976 2708 1984
rect 3308 1976 3316 1984
rect 3436 1976 3444 1984
rect 3612 1976 3620 1984
rect 3660 1976 3668 1984
rect 4444 1976 4452 1984
rect 4588 1976 4596 1984
rect 4764 1976 4772 1984
rect 4972 1976 4980 1984
rect 5084 1976 5092 1984
rect 924 1956 932 1964
rect 1228 1956 1236 1964
rect 1356 1956 1364 1964
rect 2476 1956 2484 1964
rect 2572 1956 2580 1964
rect 2748 1956 2756 1964
rect 2876 1956 2884 1964
rect 3052 1956 3060 1964
rect 3196 1956 3204 1964
rect 4300 1956 4308 1964
rect 4556 1956 4564 1964
rect 636 1936 644 1944
rect 748 1936 756 1944
rect 1900 1936 1908 1944
rect 2220 1936 2228 1944
rect 2412 1936 2420 1944
rect 2812 1936 2820 1944
rect 3004 1936 3012 1944
rect 3132 1936 3140 1944
rect 3980 1936 3988 1944
rect 4156 1936 4164 1944
rect 4204 1936 4212 1944
rect 4540 1936 4548 1944
rect 4924 1936 4932 1944
rect 412 1916 420 1924
rect 492 1916 500 1924
rect 556 1916 564 1924
rect 684 1916 692 1924
rect 860 1916 868 1924
rect 1020 1916 1028 1924
rect 1052 1916 1060 1924
rect 1212 1916 1220 1924
rect 1340 1916 1348 1924
rect 1388 1916 1396 1924
rect 12 1896 20 1904
rect 140 1896 148 1904
rect 188 1896 196 1904
rect 220 1896 228 1904
rect 364 1896 372 1904
rect 636 1896 644 1904
rect 860 1896 868 1904
rect 940 1896 948 1904
rect 988 1896 996 1904
rect 1036 1896 1044 1904
rect 1068 1896 1076 1904
rect 1116 1896 1124 1904
rect 1260 1896 1268 1904
rect 1292 1896 1300 1904
rect 1436 1896 1444 1904
rect 1804 1916 1812 1924
rect 1868 1916 1876 1924
rect 1884 1916 1892 1924
rect 1948 1916 1956 1924
rect 1532 1896 1540 1904
rect 1564 1896 1572 1904
rect 1612 1896 1620 1904
rect 1676 1896 1684 1904
rect 1724 1896 1732 1904
rect 1820 1896 1828 1904
rect 2044 1916 2052 1924
rect 2188 1916 2196 1924
rect 2284 1916 2292 1924
rect 2444 1916 2452 1924
rect 2588 1916 2596 1924
rect 2636 1916 2644 1924
rect 2716 1916 2724 1924
rect 2844 1916 2852 1924
rect 2892 1916 2900 1924
rect 2940 1916 2948 1924
rect 3036 1916 3044 1924
rect 3276 1916 3284 1924
rect 3452 1916 3460 1924
rect 3580 1916 3588 1924
rect 3596 1916 3604 1924
rect 2188 1896 2196 1904
rect 2300 1896 2308 1904
rect 2332 1896 2340 1904
rect 2460 1896 2468 1904
rect 2508 1896 2516 1904
rect 2764 1896 2772 1904
rect 44 1856 52 1864
rect 76 1856 84 1864
rect 92 1856 100 1864
rect 172 1856 180 1864
rect 220 1856 228 1864
rect 268 1856 276 1864
rect 316 1856 324 1864
rect 348 1876 356 1884
rect 380 1876 388 1884
rect 460 1876 468 1884
rect 540 1876 548 1884
rect 588 1876 596 1884
rect 652 1876 660 1884
rect 684 1876 692 1884
rect 780 1876 788 1884
rect 828 1876 836 1884
rect 988 1876 996 1884
rect 1180 1876 1188 1884
rect 1308 1876 1316 1884
rect 1420 1876 1428 1884
rect 1548 1876 1556 1884
rect 1724 1876 1732 1884
rect 1740 1876 1748 1884
rect 1900 1876 1908 1884
rect 1948 1876 1956 1884
rect 1980 1876 1988 1884
rect 1996 1876 2004 1884
rect 2076 1876 2084 1884
rect 2156 1876 2164 1884
rect 2316 1876 2324 1884
rect 2556 1876 2564 1884
rect 2668 1876 2676 1884
rect 2684 1876 2692 1884
rect 2716 1876 2724 1884
rect 2956 1896 2964 1904
rect 3052 1896 3060 1904
rect 3180 1896 3188 1904
rect 3196 1896 3204 1904
rect 3324 1896 3332 1904
rect 3372 1896 3380 1904
rect 3644 1896 3652 1904
rect 3820 1916 3828 1924
rect 3868 1916 3876 1924
rect 3916 1916 3924 1924
rect 3772 1896 3780 1904
rect 4060 1916 4068 1924
rect 4076 1916 4084 1924
rect 4252 1916 4260 1924
rect 4348 1916 4356 1924
rect 4620 1916 4628 1924
rect 4732 1916 4740 1924
rect 4748 1916 4756 1924
rect 4828 1916 4836 1924
rect 5132 1916 5140 1924
rect 5148 1916 5156 1924
rect 3980 1896 3988 1904
rect 444 1856 452 1864
rect 604 1856 612 1864
rect 700 1856 708 1864
rect 732 1856 740 1864
rect 796 1856 804 1864
rect 892 1856 900 1864
rect 908 1856 916 1864
rect 972 1856 980 1864
rect 1036 1856 1044 1864
rect 1068 1856 1076 1864
rect 1116 1856 1124 1864
rect 1164 1856 1172 1864
rect 1244 1856 1252 1864
rect 1292 1856 1300 1864
rect 1372 1856 1380 1864
rect 1404 1856 1412 1864
rect 1468 1856 1476 1864
rect 1548 1856 1556 1864
rect 1596 1856 1604 1864
rect 1628 1856 1636 1864
rect 1644 1856 1652 1864
rect 1772 1856 1780 1864
rect 1788 1856 1796 1864
rect 1852 1856 1860 1864
rect 1932 1856 1940 1864
rect 2108 1856 2116 1864
rect 2140 1856 2148 1864
rect 2220 1856 2228 1864
rect 2236 1856 2244 1864
rect 2364 1856 2372 1864
rect 2396 1856 2404 1864
rect 2492 1856 2500 1864
rect 2540 1856 2548 1864
rect 2604 1856 2612 1864
rect 2636 1856 2644 1864
rect 2860 1876 2868 1884
rect 2908 1876 2916 1884
rect 2956 1876 2964 1884
rect 3004 1876 3012 1884
rect 3100 1876 3108 1884
rect 3244 1876 3252 1884
rect 2764 1856 2772 1864
rect 2796 1856 2804 1864
rect 3084 1856 3092 1864
rect 3148 1856 3156 1864
rect 3228 1856 3236 1864
rect 3292 1856 3300 1864
rect 3340 1856 3348 1864
rect 3404 1856 3412 1864
rect 3484 1876 3492 1884
rect 3548 1876 3556 1884
rect 3676 1876 3684 1884
rect 3788 1876 3796 1884
rect 3932 1876 3940 1884
rect 4108 1896 4116 1904
rect 4028 1876 4036 1884
rect 4108 1876 4116 1884
rect 4300 1896 4308 1904
rect 4444 1896 4452 1904
rect 4604 1896 4612 1904
rect 4156 1876 4164 1884
rect 4220 1876 4228 1884
rect 4316 1876 4324 1884
rect 4428 1876 4436 1884
rect 4492 1876 4500 1884
rect 4636 1876 4644 1884
rect 4700 1876 4708 1884
rect 4972 1896 4980 1904
rect 4796 1876 4804 1884
rect 4828 1876 4836 1884
rect 4876 1876 4884 1884
rect 4892 1876 4900 1884
rect 3500 1856 3508 1864
rect 3676 1856 3684 1864
rect 3724 1856 3732 1864
rect 3740 1856 3748 1864
rect 4364 1856 4372 1864
rect 4476 1856 4484 1864
rect 4540 1856 4548 1864
rect 4572 1856 4580 1864
rect 4636 1856 4644 1864
rect 4940 1856 4948 1864
rect 4988 1856 4996 1864
rect 5052 1856 5060 1864
rect 5196 1876 5204 1884
rect 60 1836 68 1844
rect 108 1836 116 1844
rect 412 1836 420 1844
rect 748 1836 756 1844
rect 1100 1836 1108 1844
rect 1500 1836 1508 1844
rect 1692 1836 1700 1844
rect 1756 1836 1764 1844
rect 1964 1836 1972 1844
rect 2092 1836 2100 1844
rect 2252 1836 2260 1844
rect 2348 1836 2356 1844
rect 2428 1836 2436 1844
rect 2524 1836 2532 1844
rect 2988 1836 2996 1844
rect 3020 1836 3028 1844
rect 3132 1836 3140 1844
rect 3164 1836 3172 1844
rect 3260 1836 3268 1844
rect 3356 1836 3364 1844
rect 3468 1836 3476 1844
rect 3516 1836 3524 1844
rect 3916 1836 3924 1844
rect 3964 1836 3972 1844
rect 3980 1836 3988 1844
rect 4076 1836 4084 1844
rect 4140 1836 4148 1844
rect 4204 1836 4212 1844
rect 4348 1836 4356 1844
rect 4412 1836 4420 1844
rect 4524 1836 4532 1844
rect 4684 1836 4692 1844
rect 4860 1836 4868 1844
rect 5132 1836 5140 1844
rect 5164 1836 5172 1844
rect 332 1776 340 1784
rect 380 1776 388 1784
rect 428 1776 436 1784
rect 524 1776 532 1784
rect 764 1776 772 1784
rect 892 1776 900 1784
rect 1004 1776 1012 1784
rect 1196 1776 1204 1784
rect 1260 1776 1268 1784
rect 1484 1776 1492 1784
rect 1852 1776 1860 1784
rect 2124 1776 2132 1784
rect 2476 1776 2484 1784
rect 2732 1776 2740 1784
rect 2924 1776 2932 1784
rect 3004 1776 3012 1784
rect 3212 1776 3220 1784
rect 3500 1776 3508 1784
rect 3756 1776 3764 1784
rect 3948 1776 3956 1784
rect 4188 1776 4196 1784
rect 4220 1776 4228 1784
rect 4332 1776 4340 1784
rect 4492 1776 4500 1784
rect 4572 1776 4580 1784
rect 4684 1776 4692 1784
rect 4828 1776 4836 1784
rect 5068 1776 5076 1784
rect 5100 1776 5108 1784
rect 5148 1776 5156 1784
rect 140 1756 148 1764
rect 172 1756 180 1764
rect 204 1756 212 1764
rect 316 1756 324 1764
rect 396 1756 404 1764
rect 252 1736 260 1744
rect 300 1736 308 1744
rect 476 1756 484 1764
rect 508 1756 516 1764
rect 540 1756 548 1764
rect 748 1756 756 1764
rect 828 1756 836 1764
rect 844 1756 852 1764
rect 1036 1756 1044 1764
rect 1116 1756 1124 1764
rect 1180 1756 1188 1764
rect 1276 1756 1284 1764
rect 1324 1756 1332 1764
rect 1420 1756 1428 1764
rect 460 1736 468 1744
rect 492 1736 500 1744
rect 604 1736 612 1744
rect 732 1736 740 1744
rect 876 1736 884 1744
rect 924 1736 932 1744
rect 972 1736 980 1744
rect 988 1736 996 1744
rect 1068 1736 1076 1744
rect 1116 1736 1124 1744
rect 1228 1736 1236 1744
rect 1308 1736 1316 1744
rect 1388 1736 1396 1744
rect 1404 1736 1412 1744
rect 1500 1736 1508 1744
rect 1596 1756 1604 1764
rect 1692 1756 1700 1764
rect 1740 1756 1748 1764
rect 1772 1756 1780 1764
rect 1884 1756 1892 1764
rect 1948 1756 1956 1764
rect 1964 1756 1972 1764
rect 2108 1756 2116 1764
rect 2140 1756 2148 1764
rect 2156 1756 2164 1764
rect 2172 1756 2180 1764
rect 2188 1756 2196 1764
rect 2252 1756 2260 1764
rect 2284 1756 2292 1764
rect 2364 1756 2372 1764
rect 2460 1756 2468 1764
rect 2508 1756 2516 1764
rect 2796 1756 2804 1764
rect 2828 1756 2836 1764
rect 2860 1756 2868 1764
rect 2908 1756 2916 1764
rect 2940 1756 2948 1764
rect 3228 1756 3236 1764
rect 3356 1756 3364 1764
rect 3388 1756 3396 1764
rect 3452 1756 3460 1764
rect 3548 1756 3556 1764
rect 3628 1756 3636 1764
rect 3724 1756 3732 1764
rect 3740 1756 3748 1764
rect 3820 1756 3828 1764
rect 3836 1756 3844 1764
rect 4060 1756 4068 1764
rect 4076 1756 4084 1764
rect 4124 1756 4132 1764
rect 4364 1756 4372 1764
rect 4444 1756 4452 1764
rect 4588 1756 4596 1764
rect 4860 1756 4868 1764
rect 5020 1756 5028 1764
rect 5116 1756 5124 1764
rect 1628 1736 1636 1744
rect 12 1716 20 1724
rect 60 1716 68 1724
rect 92 1716 100 1724
rect 348 1716 356 1724
rect 364 1716 372 1724
rect 412 1716 420 1724
rect 540 1716 548 1724
rect 604 1716 612 1724
rect 668 1716 676 1724
rect 748 1716 756 1724
rect 780 1716 788 1724
rect 796 1716 804 1724
rect 1084 1716 1092 1724
rect 1116 1716 1124 1724
rect 1164 1716 1172 1724
rect 1212 1716 1220 1724
rect 1292 1716 1300 1724
rect 1308 1716 1316 1724
rect 1356 1716 1364 1724
rect 1452 1716 1460 1724
rect 1548 1716 1556 1724
rect 1580 1716 1588 1724
rect 1644 1716 1652 1724
rect 1676 1716 1684 1724
rect 1740 1736 1748 1744
rect 1788 1736 1796 1744
rect 1868 1736 1876 1744
rect 1916 1736 1924 1744
rect 1996 1736 2004 1744
rect 2012 1736 2020 1744
rect 2028 1736 2036 1744
rect 2252 1736 2260 1744
rect 2396 1736 2404 1744
rect 2444 1736 2452 1744
rect 2588 1736 2596 1744
rect 2604 1736 2612 1744
rect 2700 1736 2708 1744
rect 2748 1736 2756 1744
rect 2780 1736 2788 1744
rect 2988 1736 2996 1744
rect 3036 1736 3044 1744
rect 3084 1736 3092 1744
rect 3100 1736 3108 1744
rect 3180 1736 3188 1744
rect 3260 1736 3268 1744
rect 3404 1736 3412 1744
rect 3660 1736 3668 1744
rect 3852 1736 3860 1744
rect 3884 1736 3892 1744
rect 3964 1736 3972 1744
rect 4028 1736 4036 1744
rect 4060 1736 4068 1744
rect 4172 1736 4180 1744
rect 4268 1736 4276 1744
rect 4300 1736 4308 1744
rect 4316 1736 4324 1744
rect 4460 1736 4468 1744
rect 4540 1736 4548 1744
rect 4604 1736 4612 1744
rect 4652 1736 4660 1744
rect 4700 1736 4708 1744
rect 4780 1736 4788 1744
rect 4796 1736 4804 1744
rect 4828 1736 4836 1744
rect 4924 1736 4932 1744
rect 4972 1736 4980 1744
rect 4988 1736 4996 1744
rect 5020 1736 5028 1744
rect 5132 1736 5140 1744
rect 1740 1716 1748 1724
rect 1916 1716 1924 1724
rect 2092 1716 2100 1724
rect 2108 1716 2116 1724
rect 2220 1716 2228 1724
rect 2316 1716 2324 1724
rect 2348 1716 2356 1724
rect 2492 1716 2500 1724
rect 2524 1716 2532 1724
rect 2540 1716 2548 1724
rect 2684 1716 2692 1724
rect 2796 1716 2804 1724
rect 2876 1716 2884 1724
rect 3132 1716 3140 1724
rect 3164 1716 3172 1724
rect 3484 1716 3492 1724
rect 3580 1716 3588 1724
rect 3596 1716 3604 1724
rect 3692 1716 3700 1724
rect 3740 1716 3748 1724
rect 3772 1716 3780 1724
rect 3788 1716 3796 1724
rect 3868 1716 3876 1724
rect 4028 1716 4036 1724
rect 4124 1716 4132 1724
rect 4172 1716 4180 1724
rect 4364 1716 4372 1724
rect 4396 1716 4404 1724
rect 4412 1716 4420 1724
rect 4652 1716 4660 1724
rect 4748 1716 4756 1724
rect 220 1696 228 1704
rect 268 1696 276 1704
rect 284 1696 292 1704
rect 460 1696 468 1704
rect 572 1696 580 1704
rect 636 1696 644 1704
rect 700 1696 708 1704
rect 844 1696 852 1704
rect 892 1696 900 1704
rect 1260 1696 1268 1704
rect 1372 1696 1380 1704
rect 1436 1696 1444 1704
rect 1468 1696 1476 1704
rect 1788 1696 1796 1704
rect 1820 1696 1828 1704
rect 1836 1696 1844 1704
rect 2300 1696 2308 1704
rect 2412 1696 2420 1704
rect 2556 1696 2564 1704
rect 2588 1696 2596 1704
rect 2636 1696 2644 1704
rect 2748 1696 2756 1704
rect 2956 1696 2964 1704
rect 3004 1696 3012 1704
rect 3052 1696 3060 1704
rect 3212 1696 3220 1704
rect 3292 1696 3300 1704
rect 3324 1696 3332 1704
rect 3340 1696 3348 1704
rect 3436 1696 3444 1704
rect 3916 1696 3924 1704
rect 3980 1696 3988 1704
rect 4204 1696 4212 1704
rect 4220 1696 4228 1704
rect 4268 1696 4276 1704
rect 4348 1696 4356 1704
rect 4428 1696 4436 1704
rect 4492 1696 4500 1704
rect 4508 1696 4516 1704
rect 4636 1696 4644 1704
rect 4684 1696 4692 1704
rect 4732 1696 4740 1704
rect 4748 1696 4756 1704
rect 5068 1716 5076 1724
rect 4892 1696 4900 1704
rect 4924 1696 4932 1704
rect 5020 1696 5028 1704
rect 5164 1696 5172 1704
rect 204 1676 212 1684
rect 1020 1676 1028 1684
rect 1500 1676 1508 1684
rect 1724 1676 1732 1684
rect 2044 1676 2052 1684
rect 2700 1676 2708 1684
rect 2780 1676 2788 1684
rect 2892 1676 2900 1684
rect 4156 1676 4164 1684
rect 4412 1676 4420 1684
rect 4828 1676 4836 1684
rect 5068 1676 5076 1684
rect 2236 1656 2244 1664
rect 3996 1656 4004 1664
rect 4412 1656 4420 1664
rect 4956 1656 4964 1664
rect 12 1636 20 1644
rect 156 1636 164 1644
rect 236 1636 244 1644
rect 796 1636 804 1644
rect 860 1636 868 1644
rect 956 1636 964 1644
rect 1900 1636 1908 1644
rect 1996 1636 2004 1644
rect 2204 1636 2212 1644
rect 2332 1636 2340 1644
rect 2844 1636 2852 1644
rect 2924 1636 2932 1644
rect 2972 1636 2980 1644
rect 3068 1636 3076 1644
rect 3244 1636 3252 1644
rect 3804 1636 3812 1644
rect 3900 1636 3908 1644
rect 4044 1636 4052 1644
rect 4284 1636 4292 1644
rect 4412 1636 4420 1644
rect 4764 1636 4772 1644
rect 444 1576 452 1584
rect 476 1576 484 1584
rect 684 1576 692 1584
rect 844 1576 852 1584
rect 1148 1576 1156 1584
rect 1532 1576 1540 1584
rect 1564 1576 1572 1584
rect 2044 1576 2052 1584
rect 2476 1576 2484 1584
rect 2748 1576 2756 1584
rect 2924 1576 2932 1584
rect 3004 1576 3012 1584
rect 3324 1576 3332 1584
rect 3388 1576 3396 1584
rect 3484 1576 3492 1584
rect 3788 1576 3796 1584
rect 3868 1576 3876 1584
rect 4028 1576 4036 1584
rect 4204 1576 4212 1584
rect 4620 1576 4628 1584
rect 4764 1576 4772 1584
rect 4812 1576 4820 1584
rect 5100 1576 5108 1584
rect 1244 1556 1252 1564
rect 2188 1556 2196 1564
rect 2556 1556 2564 1564
rect 1084 1536 1092 1544
rect 1212 1536 1220 1544
rect 1372 1536 1380 1544
rect 1484 1536 1492 1544
rect 1676 1536 1684 1544
rect 1772 1536 1780 1544
rect 1884 1536 1892 1544
rect 1996 1536 2004 1544
rect 2268 1536 2276 1544
rect 2316 1536 2324 1544
rect 2556 1536 2564 1544
rect 3020 1536 3028 1544
rect 3244 1536 3252 1544
rect 3356 1536 3364 1544
rect 3500 1536 3508 1544
rect 3660 1536 3668 1544
rect 4268 1536 4276 1544
rect 4316 1536 4324 1544
rect 4396 1536 4404 1544
rect 4476 1536 4484 1544
rect 4540 1536 4548 1544
rect 92 1516 100 1524
rect 108 1516 116 1524
rect 236 1516 244 1524
rect 284 1516 292 1524
rect 332 1516 340 1524
rect 588 1516 596 1524
rect 828 1516 836 1524
rect 988 1516 996 1524
rect 1052 1516 1060 1524
rect 1132 1516 1140 1524
rect 1196 1516 1204 1524
rect 1292 1516 1300 1524
rect 1404 1516 1412 1524
rect 1708 1516 1716 1524
rect 1804 1516 1812 1524
rect 12 1496 20 1504
rect 188 1496 196 1504
rect 396 1496 404 1504
rect 428 1496 436 1504
rect 476 1496 484 1504
rect 652 1496 660 1504
rect 732 1496 740 1504
rect 780 1496 788 1504
rect 908 1496 916 1504
rect 1148 1496 1156 1504
rect 1244 1496 1252 1504
rect 1532 1496 1540 1504
rect 1580 1496 1588 1504
rect 1596 1496 1604 1504
rect 1660 1496 1668 1504
rect 1740 1496 1748 1504
rect 2332 1516 2340 1524
rect 2540 1516 2548 1524
rect 2700 1516 2708 1524
rect 2844 1516 2852 1524
rect 2908 1516 2916 1524
rect 3100 1516 3108 1524
rect 3148 1516 3156 1524
rect 3292 1516 3300 1524
rect 3404 1516 3412 1524
rect 1964 1496 1972 1504
rect 2044 1496 2052 1504
rect 2060 1496 2068 1504
rect 2124 1496 2132 1504
rect 2172 1496 2180 1504
rect 2268 1496 2276 1504
rect 2412 1496 2420 1504
rect 2428 1496 2436 1504
rect 2476 1496 2484 1504
rect 2556 1496 2564 1504
rect 2620 1496 2628 1504
rect 2668 1496 2676 1504
rect 2748 1496 2756 1504
rect 2780 1496 2788 1504
rect 2924 1496 2932 1504
rect 3004 1496 3012 1504
rect 3020 1496 3028 1504
rect 3228 1496 3236 1504
rect 3308 1496 3316 1504
rect 3644 1516 3652 1524
rect 3836 1516 3844 1524
rect 3548 1496 3556 1504
rect 3564 1496 3572 1504
rect 3932 1516 3940 1524
rect 4012 1516 4020 1524
rect 4076 1516 4084 1524
rect 4108 1516 4116 1524
rect 4188 1516 4196 1524
rect 4284 1516 4292 1524
rect 4492 1516 4500 1524
rect 4604 1516 4612 1524
rect 4012 1496 4020 1504
rect 4092 1496 4100 1504
rect 4268 1496 4276 1504
rect 4412 1496 4420 1504
rect 4460 1496 4468 1504
rect 4540 1496 4548 1504
rect 4588 1496 4596 1504
rect 4780 1516 4788 1524
rect 4844 1516 4852 1524
rect 4892 1516 4900 1524
rect 5116 1516 5124 1524
rect 4732 1496 4740 1504
rect 4796 1496 4804 1504
rect 4940 1496 4948 1504
rect 5036 1496 5044 1504
rect 5132 1496 5140 1504
rect 12 1476 20 1484
rect 60 1476 68 1484
rect 156 1476 164 1484
rect 204 1476 212 1484
rect 252 1476 260 1484
rect 300 1476 308 1484
rect 556 1476 564 1484
rect 588 1476 596 1484
rect 860 1476 868 1484
rect 956 1476 964 1484
rect 1084 1476 1092 1484
rect 1100 1476 1108 1484
rect 1228 1476 1236 1484
rect 1372 1476 1380 1484
rect 1676 1476 1684 1484
rect 1804 1476 1812 1484
rect 1852 1476 1860 1484
rect 1868 1476 1876 1484
rect 2092 1476 2100 1484
rect 2188 1476 2196 1484
rect 2236 1476 2244 1484
rect 2284 1476 2292 1484
rect 2364 1476 2372 1484
rect 2476 1476 2484 1484
rect 2732 1476 2740 1484
rect 2876 1476 2884 1484
rect 3132 1476 3140 1484
rect 3180 1476 3188 1484
rect 3452 1476 3460 1484
rect 3468 1476 3476 1484
rect 3676 1476 3684 1484
rect 3804 1476 3812 1484
rect 3964 1476 3972 1484
rect 3980 1476 3988 1484
rect 44 1456 52 1464
rect 156 1456 164 1464
rect 188 1456 196 1464
rect 220 1456 228 1464
rect 348 1456 356 1464
rect 380 1456 388 1464
rect 428 1456 436 1464
rect 460 1456 468 1464
rect 540 1456 548 1464
rect 652 1456 660 1464
rect 764 1456 772 1464
rect 780 1456 788 1464
rect 812 1456 820 1464
rect 876 1456 884 1464
rect 1180 1456 1188 1464
rect 1276 1456 1284 1464
rect 1356 1456 1364 1464
rect 1420 1456 1428 1464
rect 1500 1456 1508 1464
rect 1548 1456 1556 1464
rect 1612 1456 1620 1464
rect 1628 1456 1636 1464
rect 1756 1456 1764 1464
rect 1916 1456 1924 1464
rect 2012 1456 2020 1464
rect 2124 1456 2132 1464
rect 2220 1456 2228 1464
rect 2332 1456 2340 1464
rect 2380 1456 2388 1464
rect 2396 1456 2404 1464
rect 2460 1456 2468 1464
rect 2508 1456 2516 1464
rect 2524 1456 2532 1464
rect 2572 1456 2580 1464
rect 2620 1456 2628 1464
rect 2652 1456 2660 1464
rect 2700 1456 2708 1464
rect 2828 1456 2836 1464
rect 2892 1456 2900 1464
rect 2956 1456 2964 1464
rect 2972 1456 2980 1464
rect 3084 1456 3092 1464
rect 3196 1456 3204 1464
rect 3260 1456 3268 1464
rect 3276 1456 3284 1464
rect 3340 1456 3348 1464
rect 3372 1456 3380 1464
rect 3404 1456 3412 1464
rect 3516 1456 3524 1464
rect 3596 1456 3604 1464
rect 3628 1456 3636 1464
rect 3692 1456 3700 1464
rect 3756 1456 3764 1464
rect 3772 1456 3780 1464
rect 4060 1476 4068 1484
rect 4140 1476 4148 1484
rect 4156 1476 4164 1484
rect 4332 1476 4340 1484
rect 4380 1476 4388 1484
rect 4460 1476 4468 1484
rect 4492 1476 4500 1484
rect 4060 1456 4068 1464
rect 4124 1456 4132 1464
rect 4220 1456 4228 1464
rect 4236 1456 4244 1464
rect 4268 1456 4276 1464
rect 4332 1456 4340 1464
rect 4380 1456 4388 1464
rect 4412 1456 4420 1464
rect 4604 1476 4612 1484
rect 4636 1476 4644 1484
rect 4652 1476 4660 1484
rect 4748 1476 4756 1484
rect 4876 1476 4884 1484
rect 4924 1476 4932 1484
rect 4988 1476 4996 1484
rect 5084 1476 5092 1484
rect 4556 1456 4564 1464
rect 4700 1456 4708 1464
rect 4956 1456 4964 1464
rect 4972 1456 4980 1464
rect 5004 1456 5012 1464
rect 5068 1456 5076 1464
rect 5148 1456 5156 1464
rect 5164 1456 5172 1464
rect 76 1436 84 1444
rect 108 1436 116 1444
rect 284 1436 292 1444
rect 364 1436 372 1444
rect 828 1436 836 1444
rect 940 1436 948 1444
rect 1020 1436 1028 1444
rect 1132 1436 1140 1444
rect 1308 1436 1316 1444
rect 1404 1436 1412 1444
rect 1468 1436 1476 1444
rect 1788 1436 1796 1444
rect 1820 1436 1828 1444
rect 1980 1436 1988 1444
rect 2268 1436 2276 1444
rect 2588 1436 2596 1444
rect 2636 1436 2644 1444
rect 2684 1436 2692 1444
rect 2860 1436 2868 1444
rect 3100 1436 3108 1444
rect 3164 1436 3172 1444
rect 3212 1436 3220 1444
rect 3436 1436 3444 1444
rect 3580 1436 3588 1444
rect 3612 1436 3620 1444
rect 3708 1436 3716 1444
rect 4188 1436 4196 1444
rect 4668 1436 4676 1444
rect 4860 1436 4868 1444
rect 4908 1436 4916 1444
rect 12 1376 20 1384
rect 364 1376 372 1384
rect 412 1376 420 1384
rect 460 1376 468 1384
rect 604 1376 612 1384
rect 908 1376 916 1384
rect 1356 1376 1364 1384
rect 1500 1376 1508 1384
rect 1548 1376 1556 1384
rect 1596 1376 1604 1384
rect 1644 1376 1652 1384
rect 1676 1376 1684 1384
rect 1996 1376 2004 1384
rect 2220 1376 2228 1384
rect 2332 1376 2340 1384
rect 2460 1376 2468 1384
rect 2572 1376 2580 1384
rect 2716 1376 2724 1384
rect 3148 1376 3156 1384
rect 3404 1376 3412 1384
rect 3452 1376 3460 1384
rect 3612 1376 3620 1384
rect 3660 1376 3668 1384
rect 3740 1376 3748 1384
rect 3916 1376 3924 1384
rect 4172 1376 4180 1384
rect 4876 1376 4884 1384
rect 4924 1376 4932 1384
rect 108 1356 116 1364
rect 204 1356 212 1364
rect 428 1356 436 1364
rect 508 1356 516 1364
rect 524 1356 532 1364
rect 588 1356 596 1364
rect 620 1356 628 1364
rect 636 1356 644 1364
rect 668 1356 676 1364
rect 764 1356 772 1364
rect 796 1356 804 1364
rect 828 1356 836 1364
rect 876 1356 884 1364
rect 892 1356 900 1364
rect 940 1356 948 1364
rect 972 1356 980 1364
rect 1084 1356 1092 1364
rect 1132 1356 1140 1364
rect 1244 1356 1252 1364
rect 60 1336 68 1344
rect 76 1336 84 1344
rect 92 1336 100 1344
rect 236 1336 244 1344
rect 476 1336 484 1344
rect 492 1336 500 1344
rect 556 1336 564 1344
rect 716 1336 724 1344
rect 732 1336 740 1344
rect 844 1336 852 1344
rect 972 1336 980 1344
rect 1036 1336 1044 1344
rect 1244 1336 1252 1344
rect 1292 1336 1300 1344
rect 1388 1356 1396 1364
rect 1420 1356 1428 1364
rect 1532 1356 1540 1364
rect 1628 1356 1636 1364
rect 1708 1356 1716 1364
rect 1740 1356 1748 1364
rect 1820 1356 1828 1364
rect 1836 1356 1844 1364
rect 1868 1356 1876 1364
rect 2044 1356 2052 1364
rect 2108 1356 2116 1364
rect 2124 1356 2132 1364
rect 2204 1356 2212 1364
rect 2300 1356 2308 1364
rect 2364 1356 2372 1364
rect 2540 1356 2548 1364
rect 2556 1356 2564 1364
rect 2636 1356 2644 1364
rect 2652 1356 2660 1364
rect 2748 1356 2756 1364
rect 2780 1356 2788 1364
rect 2844 1356 2852 1364
rect 2876 1356 2884 1364
rect 2940 1356 2948 1364
rect 3004 1356 3012 1364
rect 3084 1356 3092 1364
rect 3100 1356 3108 1364
rect 3196 1356 3204 1364
rect 1340 1336 1348 1344
rect 1516 1336 1524 1344
rect 1580 1336 1588 1344
rect 1660 1336 1668 1344
rect 1788 1336 1796 1344
rect 1884 1336 1892 1344
rect 1932 1336 1940 1344
rect 1980 1336 1988 1344
rect 2028 1336 2036 1344
rect 2060 1336 2068 1344
rect 2252 1336 2260 1344
rect 2316 1336 2324 1344
rect 2412 1336 2420 1344
rect 2668 1336 2676 1344
rect 2764 1336 2772 1344
rect 2812 1336 2820 1344
rect 2956 1336 2964 1344
rect 2972 1336 2980 1344
rect 3164 1336 3172 1344
rect 3228 1336 3236 1344
rect 3260 1356 3268 1364
rect 3356 1356 3364 1364
rect 3724 1356 3732 1364
rect 3836 1356 3844 1364
rect 3932 1356 3940 1364
rect 3964 1356 3972 1364
rect 3996 1356 4004 1364
rect 4140 1356 4148 1364
rect 4268 1356 4276 1364
rect 4364 1356 4372 1364
rect 4412 1356 4420 1364
rect 4508 1356 4516 1364
rect 4604 1356 4612 1364
rect 4684 1356 4692 1364
rect 4732 1356 4740 1364
rect 4828 1356 4836 1364
rect 4972 1356 4980 1364
rect 5020 1356 5028 1364
rect 3436 1336 3444 1344
rect 3484 1336 3492 1344
rect 3500 1336 3508 1344
rect 3580 1336 3588 1344
rect 3596 1336 3604 1344
rect 3644 1336 3652 1344
rect 3772 1336 3780 1344
rect 3868 1336 3876 1344
rect 3964 1336 3972 1344
rect 4044 1336 4052 1344
rect 4092 1336 4100 1344
rect 4204 1336 4212 1344
rect 4220 1336 4228 1344
rect 4316 1336 4324 1344
rect 4380 1336 4388 1344
rect 4444 1336 4452 1344
rect 4540 1336 4548 1344
rect 4588 1336 4596 1344
rect 4636 1336 4644 1344
rect 4716 1336 4724 1344
rect 4780 1336 4788 1344
rect 4908 1336 4916 1344
rect 4956 1336 4964 1344
rect 5148 1336 5156 1344
rect 5164 1336 5172 1344
rect 140 1316 148 1324
rect 156 1316 164 1324
rect 252 1316 260 1324
rect 332 1316 340 1324
rect 380 1316 388 1324
rect 396 1316 404 1324
rect 668 1316 676 1324
rect 732 1316 740 1324
rect 988 1316 996 1324
rect 1116 1316 1124 1324
rect 1180 1316 1188 1324
rect 1212 1316 1220 1324
rect 12 1296 20 1304
rect 60 1296 68 1304
rect 284 1296 292 1304
rect 444 1296 452 1304
rect 524 1296 532 1304
rect 876 1296 884 1304
rect 1068 1296 1076 1304
rect 1260 1296 1268 1304
rect 1436 1316 1444 1324
rect 1468 1316 1476 1324
rect 1580 1316 1588 1324
rect 1484 1296 1492 1304
rect 1740 1316 1748 1324
rect 1836 1316 1844 1324
rect 1868 1316 1876 1324
rect 1916 1316 1924 1324
rect 2076 1316 2084 1324
rect 2156 1316 2164 1324
rect 2172 1316 2180 1324
rect 1756 1296 1764 1304
rect 1932 1296 1940 1304
rect 1964 1296 1972 1304
rect 2012 1296 2020 1304
rect 2268 1316 2276 1324
rect 2364 1316 2372 1324
rect 2396 1316 2404 1324
rect 2492 1316 2500 1324
rect 2508 1316 2516 1324
rect 2588 1316 2596 1324
rect 2604 1316 2612 1324
rect 2652 1316 2660 1324
rect 2700 1316 2708 1324
rect 2748 1316 2756 1324
rect 2812 1316 2820 1324
rect 2844 1316 2852 1324
rect 2892 1316 2900 1324
rect 3036 1316 3044 1324
rect 3052 1316 3060 1324
rect 3212 1316 3220 1324
rect 3244 1316 3252 1324
rect 3292 1316 3300 1324
rect 2348 1296 2356 1304
rect 2444 1296 2452 1304
rect 2460 1296 2468 1304
rect 2844 1296 2852 1304
rect 2988 1296 2996 1304
rect 3324 1296 3332 1304
rect 3388 1316 3396 1324
rect 3404 1296 3412 1304
rect 3436 1296 3444 1304
rect 3452 1296 3460 1304
rect 3692 1316 3700 1324
rect 3788 1316 3796 1324
rect 3884 1316 3892 1324
rect 4028 1316 4036 1324
rect 4140 1316 4148 1324
rect 4268 1316 4276 1324
rect 4300 1316 4308 1324
rect 4396 1316 4404 1324
rect 4444 1316 4452 1324
rect 4636 1316 4644 1324
rect 4716 1316 4724 1324
rect 4764 1316 4772 1324
rect 4860 1316 4868 1324
rect 5004 1316 5012 1324
rect 5052 1316 5060 1324
rect 5116 1316 5124 1324
rect 5212 1316 5220 1324
rect 3548 1296 3556 1304
rect 3644 1296 3652 1304
rect 3676 1296 3684 1304
rect 3916 1296 3924 1304
rect 3980 1296 3988 1304
rect 4124 1296 4132 1304
rect 4172 1296 4180 1304
rect 4252 1296 4260 1304
rect 4348 1296 4356 1304
rect 4572 1296 4580 1304
rect 4620 1296 4628 1304
rect 4668 1296 4676 1304
rect 4700 1296 4708 1304
rect 4796 1296 4804 1304
rect 4876 1296 4884 1304
rect 4924 1296 4932 1304
rect 5100 1296 5108 1304
rect 5196 1296 5204 1304
rect 556 1276 564 1284
rect 1212 1276 1220 1284
rect 1292 1276 1300 1284
rect 1612 1276 1620 1284
rect 2060 1276 2068 1284
rect 2252 1276 2260 1284
rect 2412 1276 2420 1284
rect 3164 1276 3172 1284
rect 3740 1276 3748 1284
rect 4044 1276 4052 1284
rect 4076 1276 4084 1284
rect 4300 1276 4308 1284
rect 4460 1276 4468 1284
rect 4508 1276 4516 1284
rect 4556 1276 4564 1284
rect 4812 1276 4820 1284
rect 5116 1276 5124 1284
rect 780 1256 788 1264
rect 4060 1256 4068 1264
rect 460 1236 468 1244
rect 812 1236 820 1244
rect 1100 1236 1108 1244
rect 1196 1236 1204 1244
rect 1804 1236 1812 1244
rect 2508 1236 2516 1244
rect 3036 1236 3044 1244
rect 3068 1236 3076 1244
rect 3276 1236 3284 1244
rect 3372 1236 3380 1244
rect 3516 1236 3524 1244
rect 3708 1236 3716 1244
rect 3868 1236 3876 1244
rect 4156 1236 4164 1244
rect 4332 1236 4340 1244
rect 4444 1236 4452 1244
rect 4524 1236 4532 1244
rect 4860 1236 4868 1244
rect 5004 1236 5012 1244
rect 5132 1236 5140 1244
rect 172 1176 180 1184
rect 332 1176 340 1184
rect 540 1176 548 1184
rect 700 1176 708 1184
rect 908 1176 916 1184
rect 1036 1176 1044 1184
rect 1500 1176 1508 1184
rect 1740 1176 1748 1184
rect 1820 1176 1828 1184
rect 1900 1176 1908 1184
rect 2172 1176 2180 1184
rect 2652 1176 2660 1184
rect 3164 1176 3172 1184
rect 3628 1176 3636 1184
rect 3772 1176 3780 1184
rect 3836 1176 3844 1184
rect 4540 1176 4548 1184
rect 28 1156 36 1164
rect 1724 1156 1732 1164
rect 1740 1156 1748 1164
rect 1868 1156 1876 1164
rect 3772 1156 3780 1164
rect 3788 1156 3796 1164
rect 4204 1156 4212 1164
rect 4220 1156 4228 1164
rect 1100 1136 1108 1144
rect 1260 1136 1268 1144
rect 1420 1136 1428 1144
rect 1516 1136 1524 1144
rect 1740 1136 1748 1144
rect 1804 1136 1812 1144
rect 2636 1136 2644 1144
rect 2924 1136 2932 1144
rect 3308 1136 3316 1144
rect 3436 1136 3444 1144
rect 3564 1136 3572 1144
rect 3772 1136 3780 1144
rect 3884 1136 3892 1144
rect 3964 1136 3972 1144
rect 4076 1136 4084 1144
rect 4108 1136 4116 1144
rect 4492 1136 4500 1144
rect 4588 1136 4596 1144
rect 4732 1136 4740 1144
rect 5116 1136 5124 1144
rect 92 1116 100 1124
rect 140 1116 148 1124
rect 204 1116 212 1124
rect 380 1116 388 1124
rect 428 1116 436 1124
rect 476 1116 484 1124
rect 572 1116 580 1124
rect 652 1116 660 1124
rect 764 1116 772 1124
rect 844 1116 852 1124
rect 892 1116 900 1124
rect 972 1116 980 1124
rect 1116 1116 1124 1124
rect 1244 1116 1252 1124
rect 1308 1116 1316 1124
rect 12 1096 20 1104
rect 156 1096 164 1104
rect 252 1096 260 1104
rect 524 1096 532 1104
rect 620 1096 628 1104
rect 700 1096 708 1104
rect 716 1096 724 1104
rect 988 1096 996 1104
rect 1100 1096 1108 1104
rect 1164 1096 1172 1104
rect 1196 1096 1204 1104
rect 1356 1096 1364 1104
rect 1580 1116 1588 1124
rect 1644 1116 1652 1124
rect 1724 1116 1732 1124
rect 1756 1116 1764 1124
rect 1916 1116 1924 1124
rect 1964 1116 1972 1124
rect 2012 1116 2020 1124
rect 2124 1116 2132 1124
rect 2236 1116 2244 1124
rect 2284 1116 2292 1124
rect 2348 1116 2356 1124
rect 2460 1116 2468 1124
rect 2492 1116 2500 1124
rect 2588 1116 2596 1124
rect 2668 1116 2676 1124
rect 2812 1116 2820 1124
rect 2860 1116 2868 1124
rect 2876 1116 2884 1124
rect 3004 1116 3012 1124
rect 3212 1116 3220 1124
rect 3276 1116 3284 1124
rect 3404 1116 3412 1124
rect 3468 1116 3476 1124
rect 3500 1116 3508 1124
rect 3644 1116 3652 1124
rect 3916 1116 3924 1124
rect 1484 1096 1492 1104
rect 1516 1096 1524 1104
rect 1660 1096 1668 1104
rect 1740 1096 1748 1104
rect 1804 1096 1812 1104
rect 2172 1096 2180 1104
rect 2220 1096 2228 1104
rect 2268 1096 2276 1104
rect 2396 1096 2404 1104
rect 2684 1096 2692 1104
rect 2732 1096 2740 1104
rect 3084 1096 3092 1104
rect 3100 1096 3108 1104
rect 3260 1096 3268 1104
rect 60 1076 68 1084
rect 76 1076 84 1084
rect 108 1076 116 1084
rect 236 1076 244 1084
rect 44 1056 52 1064
rect 284 1056 292 1064
rect 412 1076 420 1084
rect 460 1076 468 1084
rect 508 1076 516 1084
rect 620 1076 628 1084
rect 796 1076 804 1084
rect 812 1076 820 1084
rect 860 1076 868 1084
rect 972 1076 980 1084
rect 1148 1076 1156 1084
rect 1180 1076 1188 1084
rect 1292 1076 1300 1084
rect 1340 1076 1348 1084
rect 1452 1076 1460 1084
rect 1484 1076 1492 1084
rect 1612 1076 1620 1084
rect 1676 1076 1684 1084
rect 364 1056 372 1064
rect 380 1056 388 1064
rect 924 1056 932 1064
rect 1020 1056 1028 1064
rect 1052 1056 1060 1064
rect 1068 1056 1076 1064
rect 1196 1056 1204 1064
rect 1388 1056 1396 1064
rect 1452 1056 1460 1064
rect 1516 1056 1524 1064
rect 1580 1056 1588 1064
rect 1708 1076 1716 1084
rect 1788 1076 1796 1084
rect 1836 1076 1844 1084
rect 1948 1076 1956 1084
rect 1996 1076 2004 1084
rect 2076 1076 2084 1084
rect 2316 1076 2324 1084
rect 2460 1076 2468 1084
rect 2572 1076 2580 1084
rect 2588 1076 2596 1084
rect 2620 1076 2628 1084
rect 2716 1076 2724 1084
rect 2780 1076 2788 1084
rect 2828 1076 2836 1084
rect 2908 1076 2916 1084
rect 1708 1056 1716 1064
rect 1852 1056 1860 1064
rect 1884 1056 1892 1064
rect 1980 1056 1988 1064
rect 2076 1056 2084 1064
rect 2140 1056 2148 1064
rect 2188 1056 2196 1064
rect 2252 1056 2260 1064
rect 2300 1056 2308 1064
rect 2348 1056 2356 1064
rect 2364 1056 2372 1064
rect 2716 1056 2724 1064
rect 2764 1056 2772 1064
rect 2860 1056 2868 1064
rect 3036 1076 3044 1084
rect 3148 1076 3156 1084
rect 3180 1076 3188 1084
rect 3276 1076 3284 1084
rect 3324 1076 3332 1084
rect 3356 1076 3364 1084
rect 3532 1096 3540 1104
rect 3548 1096 3556 1104
rect 3740 1096 3748 1104
rect 3772 1096 3780 1104
rect 3788 1096 3796 1104
rect 3836 1096 3844 1104
rect 3420 1076 3428 1084
rect 3452 1076 3460 1084
rect 3596 1076 3604 1084
rect 3692 1076 3700 1084
rect 3772 1076 3780 1084
rect 3932 1096 3940 1104
rect 4012 1096 4020 1104
rect 4396 1116 4404 1124
rect 4556 1116 4564 1124
rect 4700 1116 4708 1124
rect 4204 1096 4212 1104
rect 4220 1096 4228 1104
rect 4316 1096 4324 1104
rect 4412 1096 4420 1104
rect 4444 1096 4452 1104
rect 4508 1096 4516 1104
rect 4540 1096 4548 1104
rect 4652 1096 4660 1104
rect 4796 1096 4804 1104
rect 5004 1116 5012 1124
rect 5180 1116 5188 1124
rect 4924 1096 4932 1104
rect 4988 1096 4996 1104
rect 5068 1096 5076 1104
rect 5148 1096 5156 1104
rect 3932 1076 3940 1084
rect 4060 1076 4068 1084
rect 4108 1076 4116 1084
rect 4172 1076 4180 1084
rect 4364 1076 4372 1084
rect 4604 1076 4612 1084
rect 4636 1076 4644 1084
rect 4748 1076 4756 1084
rect 4764 1076 4772 1084
rect 4796 1076 4804 1084
rect 5132 1076 5140 1084
rect 2956 1056 2964 1064
rect 3052 1056 3060 1064
rect 3084 1056 3092 1064
rect 3132 1056 3140 1064
rect 3148 1056 3156 1064
rect 3228 1056 3236 1064
rect 3516 1056 3524 1064
rect 3612 1056 3620 1064
rect 3692 1056 3700 1064
rect 3724 1056 3732 1064
rect 3756 1056 3764 1064
rect 3820 1056 3828 1064
rect 3868 1056 3876 1064
rect 3980 1056 3988 1064
rect 4172 1056 4180 1064
rect 4252 1056 4260 1064
rect 4348 1056 4356 1064
rect 4444 1056 4452 1064
rect 4460 1056 4468 1064
rect 4508 1056 4516 1064
rect 4684 1056 4692 1064
rect 4828 1056 4836 1064
rect 4844 1056 4852 1064
rect 4892 1056 4900 1064
rect 4972 1056 4980 1064
rect 5020 1056 5028 1064
rect 5036 1056 5044 1064
rect 5180 1056 5188 1064
rect 140 1036 148 1044
rect 428 1036 436 1044
rect 476 1036 484 1044
rect 732 1036 740 1044
rect 844 1036 852 1044
rect 892 1036 900 1044
rect 956 1036 964 1044
rect 1132 1036 1140 1044
rect 1244 1036 1252 1044
rect 1276 1036 1284 1044
rect 1308 1036 1316 1044
rect 1596 1036 1604 1044
rect 1628 1036 1636 1044
rect 1916 1036 1924 1044
rect 2028 1036 2036 1044
rect 2124 1036 2132 1044
rect 2204 1036 2212 1044
rect 2428 1036 2436 1044
rect 2604 1036 2612 1044
rect 2700 1036 2708 1044
rect 2796 1036 2804 1044
rect 2876 1036 2884 1044
rect 3212 1036 3220 1044
rect 3276 1036 3284 1044
rect 3388 1036 3396 1044
rect 3500 1036 3508 1044
rect 3564 1036 3572 1044
rect 3644 1036 3652 1044
rect 3708 1036 3716 1044
rect 3884 1036 3892 1044
rect 4060 1036 4068 1044
rect 4300 1036 4308 1044
rect 4396 1036 4404 1044
rect 4572 1036 4580 1044
rect 4604 1036 4612 1044
rect 4700 1036 4708 1044
rect 4812 1036 4820 1044
rect 4956 1036 4964 1044
rect 5100 1036 5108 1044
rect 5196 1036 5204 1044
rect 28 976 36 984
rect 60 976 68 984
rect 124 976 132 984
rect 188 976 196 984
rect 412 976 420 984
rect 508 976 516 984
rect 652 976 660 984
rect 700 976 708 984
rect 732 976 740 984
rect 1036 976 1044 984
rect 1132 976 1140 984
rect 1180 976 1188 984
rect 1212 976 1220 984
rect 1308 976 1316 984
rect 1356 976 1364 984
rect 1452 976 1460 984
rect 1500 976 1508 984
rect 1644 976 1652 984
rect 1676 976 1684 984
rect 1772 976 1780 984
rect 1852 976 1860 984
rect 1948 976 1956 984
rect 2092 976 2100 984
rect 2156 976 2164 984
rect 2348 976 2356 984
rect 2476 976 2484 984
rect 2508 976 2516 984
rect 2876 976 2884 984
rect 2988 976 2996 984
rect 3020 976 3028 984
rect 3372 976 3380 984
rect 3452 976 3460 984
rect 3484 976 3492 984
rect 3692 976 3700 984
rect 4124 976 4132 984
rect 4284 976 4292 984
rect 4764 976 4772 984
rect 4780 976 4788 984
rect 4828 976 4836 984
rect 5036 976 5044 984
rect 5132 976 5140 984
rect 5196 976 5204 984
rect 204 956 212 964
rect 252 956 260 964
rect 364 956 372 964
rect 396 956 404 964
rect 540 956 548 964
rect 12 936 20 944
rect 108 936 116 944
rect 140 936 148 944
rect 156 936 164 944
rect 284 936 292 944
rect 300 936 308 944
rect 316 936 324 944
rect 396 936 404 944
rect 444 936 452 944
rect 524 936 532 944
rect 572 936 580 944
rect 620 936 628 944
rect 716 936 724 944
rect 44 896 52 904
rect 60 896 68 904
rect 108 896 116 904
rect 236 916 244 924
rect 428 916 436 924
rect 444 916 452 924
rect 252 896 260 904
rect 332 896 340 904
rect 348 896 356 904
rect 524 896 532 904
rect 684 896 692 904
rect 812 956 820 964
rect 844 956 852 964
rect 860 956 868 964
rect 892 956 900 964
rect 924 956 932 964
rect 972 956 980 964
rect 1004 956 1012 964
rect 1068 956 1076 964
rect 764 936 772 944
rect 956 936 964 944
rect 812 916 820 924
rect 924 916 932 924
rect 956 916 964 924
rect 1020 936 1028 944
rect 1116 956 1124 964
rect 1276 956 1284 964
rect 1116 936 1124 944
rect 1148 936 1156 944
rect 1196 936 1204 944
rect 1420 956 1428 964
rect 1660 956 1668 964
rect 1868 956 1876 964
rect 1884 956 1892 964
rect 1932 956 1940 964
rect 1964 956 1972 964
rect 1980 956 1988 964
rect 2076 956 2084 964
rect 2188 956 2196 964
rect 2236 956 2244 964
rect 2268 956 2276 964
rect 2380 956 2388 964
rect 2444 956 2452 964
rect 2460 956 2468 964
rect 2524 956 2532 964
rect 2540 956 2548 964
rect 2652 956 2660 964
rect 2684 956 2692 964
rect 2700 956 2708 964
rect 2796 956 2804 964
rect 2812 956 2820 964
rect 2860 956 2868 964
rect 2892 956 2900 964
rect 3132 956 3140 964
rect 3260 956 3268 964
rect 3276 956 3284 964
rect 3340 956 3348 964
rect 3404 956 3412 964
rect 3468 956 3476 964
rect 3628 956 3636 964
rect 3724 956 3732 964
rect 3772 956 3780 964
rect 3804 956 3812 964
rect 3868 956 3876 964
rect 3996 956 4004 964
rect 4012 956 4020 964
rect 4092 956 4100 964
rect 4108 956 4116 964
rect 4140 956 4148 964
rect 4172 956 4180 964
rect 4204 956 4212 964
rect 4396 956 4404 964
rect 4460 956 4468 964
rect 4668 956 4676 964
rect 4908 956 4916 964
rect 4956 956 4964 964
rect 5148 956 5156 964
rect 1372 936 1380 944
rect 1484 936 1492 944
rect 1740 936 1748 944
rect 1836 936 1844 944
rect 1932 936 1940 944
rect 1996 936 2004 944
rect 2124 936 2132 944
rect 2172 936 2180 944
rect 2220 936 2228 944
rect 2364 936 2372 944
rect 2412 936 2420 944
rect 2572 936 2580 944
rect 2716 936 2724 944
rect 2956 936 2964 944
rect 3164 936 3172 944
rect 3212 936 3220 944
rect 3308 936 3316 944
rect 3356 936 3364 944
rect 3436 936 3444 944
rect 1068 916 1076 924
rect 1228 916 1236 924
rect 1324 916 1332 924
rect 1372 916 1380 924
rect 1468 916 1476 924
rect 1612 916 1620 924
rect 1692 916 1700 924
rect 2268 916 2276 924
rect 2284 916 2292 924
rect 2300 916 2308 924
rect 2428 916 2436 924
rect 2492 916 2500 924
rect 2652 916 2660 924
rect 2668 916 2676 924
rect 2748 916 2756 924
rect 2764 916 2772 924
rect 2828 916 2836 924
rect 2860 916 2868 924
rect 2892 916 2900 924
rect 2940 916 2948 924
rect 2988 916 2996 924
rect 3180 916 3188 924
rect 3228 916 3236 924
rect 3532 936 3540 944
rect 3612 936 3620 944
rect 3676 936 3684 944
rect 3804 936 3812 944
rect 3916 936 3924 944
rect 4044 936 4052 944
rect 4076 936 4084 944
rect 4236 936 4244 944
rect 4268 936 4276 944
rect 4316 936 4324 944
rect 4348 936 4356 944
rect 4412 936 4420 944
rect 4508 936 4516 944
rect 4588 936 4596 944
rect 4700 936 4708 944
rect 4716 936 4724 944
rect 4732 936 4740 944
rect 4812 936 4820 944
rect 4876 936 4884 944
rect 5020 936 5028 944
rect 5100 936 5108 944
rect 3660 916 3668 924
rect 3756 916 3764 924
rect 3772 916 3780 924
rect 3804 916 3812 924
rect 3900 916 3908 924
rect 3948 916 3956 924
rect 3980 916 3988 924
rect 4044 916 4052 924
rect 4172 916 4180 924
rect 4204 916 4212 924
rect 4252 916 4260 924
rect 4268 916 4276 924
rect 4348 916 4356 924
rect 4444 916 4452 924
rect 4492 916 4500 924
rect 764 896 772 904
rect 796 896 804 904
rect 1052 896 1060 904
rect 1180 896 1188 904
rect 1228 896 1236 904
rect 1340 896 1348 904
rect 1532 896 1540 904
rect 1564 896 1572 904
rect 1708 896 1716 904
rect 1884 896 1892 904
rect 1980 896 1988 904
rect 2028 896 2036 904
rect 2092 896 2100 904
rect 2140 896 2148 904
rect 2188 896 2196 904
rect 2252 896 2260 904
rect 2332 896 2340 904
rect 2380 896 2388 904
rect 2604 896 2612 904
rect 2988 896 2996 904
rect 3068 896 3076 904
rect 3212 896 3220 904
rect 3260 896 3268 904
rect 3340 896 3348 904
rect 3388 896 3396 904
rect 3484 896 3492 904
rect 3564 896 3572 904
rect 3948 896 3956 904
rect 4012 896 4020 904
rect 4316 896 4324 904
rect 4444 896 4452 904
rect 4604 916 4612 924
rect 4876 916 4884 924
rect 4908 916 4916 924
rect 4924 916 4932 924
rect 5020 916 5028 924
rect 4556 896 4564 904
rect 4668 896 4676 904
rect 4764 896 4772 904
rect 4780 896 4788 904
rect 4812 896 4820 904
rect 5004 896 5012 904
rect 5116 916 5124 924
rect 5164 916 5172 924
rect 5068 896 5076 904
rect 5196 896 5204 904
rect 476 876 484 884
rect 828 876 836 884
rect 876 876 884 884
rect 1388 876 1396 884
rect 1756 876 1764 884
rect 1788 876 1796 884
rect 1804 876 1812 884
rect 2540 876 2548 884
rect 2956 876 2964 884
rect 3292 876 3300 884
rect 3580 876 3588 884
rect 3708 876 3716 884
rect 3852 876 3860 884
rect 3916 876 3924 884
rect 4348 876 4356 884
rect 4508 876 4516 884
rect 4524 876 4532 884
rect 4604 876 4612 884
rect 1948 856 1956 864
rect 3932 856 3940 864
rect 364 836 372 844
rect 988 836 996 844
rect 1724 836 1732 844
rect 2044 836 2052 844
rect 2972 836 2980 844
rect 3596 836 3604 844
rect 3772 836 3780 844
rect 4204 836 4212 844
rect 4332 836 4340 844
rect 4428 836 4436 844
rect 444 776 452 784
rect 1164 776 1172 784
rect 1356 776 1364 784
rect 1708 776 1716 784
rect 1772 776 1780 784
rect 1900 776 1908 784
rect 2124 776 2132 784
rect 2188 776 2196 784
rect 3020 776 3028 784
rect 3180 776 3188 784
rect 3228 776 3236 784
rect 3372 776 3380 784
rect 3564 776 3572 784
rect 3660 776 3668 784
rect 3788 776 3796 784
rect 3948 776 3956 784
rect 4812 776 4820 784
rect 5020 776 5028 784
rect 5164 776 5172 784
rect 1116 756 1124 764
rect 1500 756 1508 764
rect 3196 756 3204 764
rect 3996 756 4004 764
rect 4076 756 4084 764
rect 4652 756 4660 764
rect 4892 756 4900 764
rect 540 736 548 744
rect 812 736 820 744
rect 956 736 964 744
rect 1036 736 1044 744
rect 1084 736 1092 744
rect 1324 736 1332 744
rect 2140 736 2148 744
rect 2204 736 2212 744
rect 2476 736 2484 744
rect 2508 736 2516 744
rect 2588 736 2596 744
rect 3340 736 3348 744
rect 3388 736 3396 744
rect 3740 736 3748 744
rect 3932 736 3940 744
rect 4012 736 4020 744
rect 4316 736 4324 744
rect 4396 736 4404 744
rect 4796 736 4804 744
rect 4828 736 4836 744
rect 4876 736 4884 744
rect 4956 736 4964 744
rect 5132 736 5140 744
rect 44 716 52 724
rect 140 716 148 724
rect 188 716 196 724
rect 268 716 276 724
rect 316 716 324 724
rect 380 716 388 724
rect 476 716 484 724
rect 604 716 612 724
rect 844 716 852 724
rect 892 716 900 724
rect 1004 716 1012 724
rect 1484 716 1492 724
rect 1564 716 1572 724
rect 1596 716 1604 724
rect 1628 716 1636 724
rect 1644 716 1652 724
rect 1692 716 1700 724
rect 1852 716 1860 724
rect 1916 716 1924 724
rect 2028 716 2036 724
rect 2060 716 2068 724
rect 2364 716 2372 724
rect 364 696 372 704
rect 428 696 436 704
rect 556 696 564 704
rect 652 696 660 704
rect 12 676 20 684
rect 172 676 180 684
rect 220 676 228 684
rect 236 676 244 684
rect 284 676 292 684
rect 332 676 340 684
rect 412 676 420 684
rect 508 676 516 684
rect 556 676 564 684
rect 748 696 756 704
rect 1148 696 1156 704
rect 1180 696 1188 704
rect 1356 696 1364 704
rect 1436 696 1444 704
rect 1580 696 1588 704
rect 1948 696 1956 704
rect 2012 696 2020 704
rect 2204 696 2212 704
rect 2332 696 2340 704
rect 2412 696 2420 704
rect 2428 696 2436 704
rect 2476 696 2484 704
rect 2524 696 2532 704
rect 2652 716 2660 724
rect 2716 716 2724 724
rect 2812 716 2820 724
rect 3004 716 3012 724
rect 3436 716 3444 724
rect 3532 716 3540 724
rect 3580 716 3588 724
rect 3676 716 3684 724
rect 3964 716 3972 724
rect 4204 716 4212 724
rect 4220 716 4228 724
rect 4284 716 4292 724
rect 4348 716 4356 724
rect 4492 716 4500 724
rect 2748 696 2756 704
rect 2764 696 2772 704
rect 2780 696 2788 704
rect 2908 696 2916 704
rect 3020 696 3028 704
rect 3148 696 3156 704
rect 3180 696 3188 704
rect 3292 696 3300 704
rect 3500 696 3508 704
rect 3596 696 3604 704
rect 3692 696 3700 704
rect 3708 696 3716 704
rect 3772 696 3780 704
rect 3820 696 3828 704
rect 3836 696 3844 704
rect 4060 696 4068 704
rect 4076 696 4084 704
rect 4172 696 4180 704
rect 4268 696 4276 704
rect 4412 696 4420 704
rect 4508 696 4516 704
rect 4636 716 4644 724
rect 4732 716 4740 724
rect 5036 716 5044 724
rect 4652 696 4660 704
rect 4780 696 4788 704
rect 4956 696 4964 704
rect 5052 696 5060 704
rect 700 676 708 684
rect 764 676 772 684
rect 812 676 820 684
rect 860 676 868 684
rect 1004 676 1012 684
rect 1036 676 1044 684
rect 1052 676 1060 684
rect 1228 676 1236 684
rect 1276 676 1284 684
rect 1452 676 1460 684
rect 1628 676 1636 684
rect 1676 676 1684 684
rect 1724 676 1732 684
rect 1804 676 1812 684
rect 1964 676 1972 684
rect 2092 676 2100 684
rect 2172 676 2180 684
rect 2268 676 2276 684
rect 2332 676 2340 684
rect 2412 676 2420 684
rect 2476 676 2484 684
rect 2604 676 2612 684
rect 2700 676 2708 684
rect 2732 676 2740 684
rect 2860 676 2868 684
rect 2956 676 2964 684
rect 2972 676 2980 684
rect 3052 676 3060 684
rect 3340 676 3348 684
rect 3404 676 3412 684
rect 3484 676 3492 684
rect 3548 676 3556 684
rect 3788 676 3796 684
rect 3836 676 3844 684
rect 3932 676 3940 684
rect 3980 676 3988 684
rect 4012 676 4020 684
rect 4156 676 4164 684
rect 4252 676 4260 684
rect 4316 676 4324 684
rect 4364 676 4372 684
rect 4396 676 4404 684
rect 4444 676 4452 684
rect 4604 676 4612 684
rect 4700 676 4708 684
rect 4908 676 4916 684
rect 5036 676 5044 684
rect 5100 676 5108 684
rect 60 656 68 664
rect 124 656 132 664
rect 332 656 340 664
rect 460 656 468 664
rect 524 656 532 664
rect 620 656 628 664
rect 700 656 708 664
rect 716 656 724 664
rect 940 656 948 664
rect 1100 656 1108 664
rect 1132 656 1140 664
rect 1196 656 1204 664
rect 1212 656 1220 664
rect 1340 656 1348 664
rect 1388 656 1396 664
rect 1404 656 1412 664
rect 1532 656 1540 664
rect 1548 656 1556 664
rect 1756 656 1764 664
rect 1804 656 1812 664
rect 1868 656 1876 664
rect 1996 656 2004 664
rect 2044 656 2052 664
rect 2108 656 2116 664
rect 2204 656 2212 664
rect 2252 656 2260 664
rect 2284 656 2292 664
rect 2300 656 2308 664
rect 2380 656 2388 664
rect 2412 656 2420 664
rect 2428 656 2436 664
rect 2556 656 2564 664
rect 2572 656 2580 664
rect 2700 656 2708 664
rect 2748 656 2756 664
rect 2780 656 2788 664
rect 2812 656 2820 664
rect 2876 656 2884 664
rect 3052 656 3060 664
rect 3068 656 3076 664
rect 3100 656 3108 664
rect 3132 656 3140 664
rect 3148 656 3156 664
rect 3212 656 3220 664
rect 3244 656 3252 664
rect 3260 656 3268 664
rect 3452 656 3460 664
rect 3596 656 3604 664
rect 3628 656 3636 664
rect 3724 656 3732 664
rect 3820 656 3828 664
rect 3868 656 3876 664
rect 4028 656 4036 664
rect 4108 656 4116 664
rect 4124 656 4132 664
rect 4300 656 4308 664
rect 4412 656 4420 664
rect 4444 656 4452 664
rect 4540 656 4548 664
rect 4684 656 4692 664
rect 4716 656 4724 664
rect 4796 656 4804 664
rect 4828 656 4836 664
rect 4924 656 4932 664
rect 4972 656 4980 664
rect 5084 656 5092 664
rect 5148 656 5156 664
rect 28 636 36 644
rect 76 636 84 644
rect 140 636 148 644
rect 188 636 196 644
rect 268 636 276 644
rect 348 636 356 644
rect 380 636 388 644
rect 476 636 484 644
rect 604 636 612 644
rect 684 636 692 644
rect 780 636 788 644
rect 828 636 836 644
rect 924 636 932 644
rect 972 636 980 644
rect 1004 636 1012 644
rect 1244 636 1252 644
rect 1308 636 1316 644
rect 1420 636 1428 644
rect 1596 636 1604 644
rect 1660 636 1668 644
rect 1836 636 1844 644
rect 1980 636 1988 644
rect 2060 636 2068 644
rect 2140 636 2148 644
rect 2364 636 2372 644
rect 2492 636 2500 644
rect 2540 636 2548 644
rect 2636 636 2644 644
rect 2828 636 2836 644
rect 2924 636 2932 644
rect 2988 636 2996 644
rect 3324 636 3332 644
rect 3436 636 3444 644
rect 3468 636 3476 644
rect 3516 636 3524 644
rect 3756 636 3764 644
rect 3900 636 3908 644
rect 4140 636 4148 644
rect 4204 636 4212 644
rect 4220 636 4228 644
rect 4492 636 4500 644
rect 4572 636 4580 644
rect 4620 636 4628 644
rect 5116 636 5124 644
rect 204 576 212 584
rect 348 576 356 584
rect 444 576 452 584
rect 524 576 532 584
rect 620 576 628 584
rect 716 576 724 584
rect 1084 576 1092 584
rect 1468 576 1476 584
rect 1724 576 1732 584
rect 1852 576 1860 584
rect 2076 576 2084 584
rect 2188 576 2196 584
rect 2204 576 2212 584
rect 2572 576 2580 584
rect 2860 576 2868 584
rect 2908 576 2916 584
rect 3004 576 3012 584
rect 3052 576 3060 584
rect 3196 576 3204 584
rect 3340 576 3348 584
rect 3484 576 3492 584
rect 3692 576 3700 584
rect 3932 576 3940 584
rect 4012 576 4020 584
rect 4060 576 4068 584
rect 4124 576 4132 584
rect 4268 576 4276 584
rect 4716 576 4724 584
rect 4732 576 4740 584
rect 4892 576 4900 584
rect 12 556 20 564
rect 44 556 52 564
rect 140 556 148 564
rect 156 556 164 564
rect 220 556 228 564
rect 268 556 276 564
rect 92 536 100 544
rect 156 536 164 544
rect 412 556 420 564
rect 364 536 372 544
rect 476 556 484 564
rect 540 556 548 564
rect 572 556 580 564
rect 604 556 612 564
rect 700 556 708 564
rect 748 556 756 564
rect 764 556 772 564
rect 812 556 820 564
rect 828 556 836 564
rect 924 556 932 564
rect 956 556 964 564
rect 1020 556 1028 564
rect 1068 556 1076 564
rect 1132 556 1140 564
rect 1340 556 1348 564
rect 1372 556 1380 564
rect 556 536 564 544
rect 684 536 692 544
rect 780 536 788 544
rect 812 536 820 544
rect 876 536 884 544
rect 1004 536 1012 544
rect 1148 536 1156 544
rect 1436 556 1444 564
rect 1532 556 1540 564
rect 1564 556 1572 564
rect 1596 556 1604 564
rect 1708 556 1716 564
rect 1804 556 1812 564
rect 1884 556 1892 564
rect 1916 556 1924 564
rect 2012 556 2020 564
rect 2108 556 2116 564
rect 2252 556 2260 564
rect 2348 556 2356 564
rect 2380 556 2388 564
rect 2476 556 2484 564
rect 2524 556 2532 564
rect 1532 536 1540 544
rect 1612 536 1620 544
rect 1644 536 1652 544
rect 1676 536 1684 544
rect 1756 536 1764 544
rect 1820 536 1828 544
rect 1868 536 1876 544
rect 1964 536 1972 544
rect 2060 536 2068 544
rect 2156 536 2164 544
rect 2236 536 2244 544
rect 2300 536 2308 544
rect 2348 536 2356 544
rect 2396 536 2404 544
rect 2444 536 2452 544
rect 2652 556 2660 564
rect 2684 556 2692 564
rect 2764 556 2772 564
rect 2812 556 2820 564
rect 2876 556 2884 564
rect 2940 556 2948 564
rect 3020 556 3028 564
rect 3068 556 3076 564
rect 3084 556 3092 564
rect 3116 556 3124 564
rect 3132 556 3140 564
rect 3164 556 3172 564
rect 3260 556 3268 564
rect 3308 556 3316 564
rect 3356 556 3364 564
rect 3404 556 3412 564
rect 3596 556 3604 564
rect 3644 556 3652 564
rect 3676 556 3684 564
rect 3772 556 3780 564
rect 3788 556 3796 564
rect 3820 556 3828 564
rect 3836 556 3844 564
rect 4076 556 4084 564
rect 4172 556 4180 564
rect 4204 556 4212 564
rect 4252 556 4260 564
rect 4316 556 4324 564
rect 4476 556 4484 564
rect 4540 556 4548 564
rect 4588 556 4596 564
rect 4652 556 4660 564
rect 2604 536 2612 544
rect 2668 536 2676 544
rect 2700 536 2708 544
rect 2716 536 2724 544
rect 2892 536 2900 544
rect 3276 536 3284 544
rect 3580 536 3588 544
rect 3692 536 3700 544
rect 3724 536 3732 544
rect 3756 536 3764 544
rect 3884 536 3892 544
rect 3964 536 3972 544
rect 3980 536 3988 544
rect 4028 536 4036 544
rect 4156 536 4164 544
rect 4332 536 4340 544
rect 4460 536 4468 544
rect 4508 536 4516 544
rect 4604 536 4612 544
rect 4684 536 4692 544
rect 4764 556 4772 564
rect 4844 556 4852 564
rect 4876 556 4884 564
rect 4924 556 4932 564
rect 5004 556 5012 564
rect 5036 556 5044 564
rect 5052 556 5060 564
rect 5068 556 5076 564
rect 5132 556 5140 564
rect 5196 556 5204 564
rect 5116 536 5124 544
rect 92 516 100 524
rect 140 516 148 524
rect 188 516 196 524
rect 236 516 244 524
rect 332 516 340 524
rect 380 516 388 524
rect 492 516 500 524
rect 508 516 516 524
rect 748 516 756 524
rect 780 516 788 524
rect 876 516 884 524
rect 972 516 980 524
rect 1036 516 1044 524
rect 1068 516 1076 524
rect 1100 516 1108 524
rect 1228 516 1236 524
rect 1292 516 1300 524
rect 1324 516 1332 524
rect 1372 516 1380 524
rect 1420 516 1428 524
rect 1452 516 1460 524
rect 1500 516 1508 524
rect 1644 516 1652 524
rect 1772 516 1780 524
rect 1804 516 1812 524
rect 1948 516 1956 524
rect 2044 516 2052 524
rect 2140 516 2148 524
rect 2284 516 2292 524
rect 2396 516 2404 524
rect 2428 516 2436 524
rect 2476 516 2484 524
rect 2604 516 2612 524
rect 60 496 68 504
rect 332 496 340 504
rect 588 496 596 504
rect 652 496 660 504
rect 908 496 916 504
rect 972 496 980 504
rect 1580 496 1588 504
rect 1676 496 1684 504
rect 1724 496 1732 504
rect 1900 496 1908 504
rect 2028 496 2036 504
rect 2092 496 2100 504
rect 2188 496 2196 504
rect 2204 496 2212 504
rect 2668 496 2676 504
rect 2796 516 2804 524
rect 2844 516 2852 524
rect 2956 516 2964 524
rect 2972 516 2980 524
rect 2988 516 2996 524
rect 3036 516 3044 524
rect 3084 516 3092 524
rect 3116 516 3124 524
rect 3164 516 3172 524
rect 3212 516 3220 524
rect 3228 516 3236 524
rect 3276 516 3284 524
rect 3308 516 3316 524
rect 3324 516 3332 524
rect 3372 516 3380 524
rect 2924 496 2932 504
rect 3148 496 3156 504
rect 3628 516 3636 524
rect 3644 516 3652 524
rect 3740 516 3748 524
rect 3772 516 3780 524
rect 3868 516 3876 524
rect 3932 516 3940 524
rect 3548 496 3556 504
rect 3932 496 3940 504
rect 4012 496 4020 504
rect 4108 516 4116 524
rect 4236 516 4244 524
rect 4284 516 4292 524
rect 4556 516 4564 524
rect 4796 516 4804 524
rect 4812 516 4820 524
rect 4956 516 4964 524
rect 4972 516 4980 524
rect 5164 516 5172 524
rect 4124 496 4132 504
rect 4364 496 4372 504
rect 4428 496 4436 504
rect 4540 496 4548 504
rect 4572 496 4580 504
rect 4620 496 4628 504
rect 4636 496 4644 504
rect 4828 496 4836 504
rect 5084 496 5092 504
rect 316 476 324 484
rect 940 476 948 484
rect 1180 476 1188 484
rect 1852 476 1860 484
rect 1964 476 1972 484
rect 1996 476 2004 484
rect 892 456 900 464
rect 1692 456 1700 464
rect 2332 476 2340 484
rect 2428 476 2436 484
rect 3164 476 3172 484
rect 3452 476 3460 484
rect 3692 476 3700 484
rect 3884 476 3892 484
rect 3916 476 3924 484
rect 4684 476 4692 484
rect 4716 476 4724 484
rect 5036 476 5044 484
rect 2460 456 2468 464
rect 3164 456 3172 464
rect 4492 456 4500 464
rect 204 436 212 444
rect 1116 436 1124 444
rect 1660 436 1668 444
rect 1980 436 1988 444
rect 2044 436 2052 444
rect 2124 436 2132 444
rect 2284 436 2292 444
rect 2636 436 2644 444
rect 2732 436 2740 444
rect 2828 436 2836 444
rect 3148 436 3156 444
rect 3164 436 3172 444
rect 3292 436 3300 444
rect 4188 436 4196 444
rect 4236 436 4244 444
rect 4300 436 4308 444
rect 4396 436 4404 444
rect 4860 436 4868 444
rect 4972 436 4980 444
rect 5100 436 5108 444
rect 1404 376 1412 384
rect 2044 376 2052 384
rect 2956 376 2964 384
rect 3116 376 3124 384
rect 3180 376 3188 384
rect 3372 376 3380 384
rect 3580 376 3588 384
rect 3852 376 3860 384
rect 4172 376 4180 384
rect 4732 376 4740 384
rect 5116 376 5124 384
rect 5164 376 5172 384
rect 828 356 836 364
rect 3372 356 3380 364
rect 540 336 548 344
rect 604 336 612 344
rect 620 336 628 344
rect 668 336 676 344
rect 844 336 852 344
rect 988 336 996 344
rect 1388 336 1396 344
rect 1692 336 1700 344
rect 1740 336 1748 344
rect 2060 336 2068 344
rect 2812 336 2820 344
rect 2908 336 2916 344
rect 3372 336 3380 344
rect 3996 336 4004 344
rect 4316 336 4324 344
rect 4604 336 4612 344
rect 4668 336 4676 344
rect 4828 336 4836 344
rect 5020 336 5028 344
rect 12 316 20 324
rect 44 316 52 324
rect 140 316 148 324
rect 268 316 276 324
rect 284 316 292 324
rect 460 316 468 324
rect 732 316 740 324
rect 812 316 820 324
rect 92 296 100 304
rect 172 296 180 304
rect 220 296 228 304
rect 332 296 340 304
rect 364 296 372 304
rect 380 296 388 304
rect 508 296 516 304
rect 604 296 612 304
rect 684 296 692 304
rect 860 296 868 304
rect 1036 316 1044 324
rect 1068 316 1076 324
rect 1132 316 1140 324
rect 1196 316 1204 324
rect 1276 316 1284 324
rect 1292 316 1300 324
rect 1548 316 1556 324
rect 1596 316 1604 324
rect 1644 316 1652 324
rect 1788 316 1796 324
rect 1884 316 1892 324
rect 1916 316 1924 324
rect 1932 316 1940 324
rect 2140 316 2148 324
rect 988 296 996 304
rect 1148 296 1156 304
rect 1340 296 1348 304
rect 1356 296 1364 304
rect 1436 296 1444 304
rect 1708 296 1716 304
rect 1756 296 1764 304
rect 1852 296 1860 304
rect 2172 296 2180 304
rect 2204 296 2212 304
rect 2332 316 2340 324
rect 2572 316 2580 324
rect 2604 316 2612 324
rect 2620 316 2628 324
rect 2668 316 2676 324
rect 2940 316 2948 324
rect 3004 316 3012 324
rect 2364 296 2372 304
rect 2428 296 2436 304
rect 2460 296 2468 304
rect 2508 296 2516 304
rect 2716 296 2724 304
rect 2796 296 2804 304
rect 2812 296 2820 304
rect 2892 296 2900 304
rect 3084 316 3092 324
rect 3164 316 3172 324
rect 3356 316 3364 324
rect 3468 316 3476 324
rect 3612 316 3620 324
rect 3644 316 3652 324
rect 3692 316 3700 324
rect 3788 316 3796 324
rect 3836 316 3844 324
rect 3964 316 3972 324
rect 4124 316 4132 324
rect 4252 316 4260 324
rect 4300 316 4308 324
rect 4412 316 4420 324
rect 4652 316 4660 324
rect 4716 316 4724 324
rect 5100 316 5108 324
rect 5180 316 5188 324
rect 3100 296 3108 304
rect 44 276 52 284
rect 188 276 196 284
rect 236 276 244 284
rect 316 276 324 284
rect 428 276 436 284
rect 652 276 660 284
rect 764 276 772 284
rect 780 276 788 284
rect 940 276 948 284
rect 1004 276 1012 284
rect 1100 276 1108 284
rect 1132 276 1140 284
rect 1228 276 1236 284
rect 1244 276 1252 284
rect 1324 276 1332 284
rect 1420 276 1428 284
rect 1516 276 1524 284
rect 1612 276 1620 284
rect 1740 276 1748 284
rect 1836 276 1844 284
rect 1900 276 1908 284
rect 1996 276 2004 284
rect 2092 276 2100 284
rect 2108 276 2116 284
rect 2284 276 2292 284
rect 2380 276 2388 284
rect 76 256 84 264
rect 92 256 100 264
rect 124 256 132 264
rect 188 256 196 264
rect 332 256 340 264
rect 412 256 420 264
rect 444 256 452 264
rect 476 256 484 264
rect 556 256 564 264
rect 652 256 660 264
rect 844 256 852 264
rect 892 256 900 264
rect 956 256 964 264
rect 1084 256 1092 264
rect 1116 256 1124 264
rect 1180 256 1188 264
rect 1372 256 1380 264
rect 1468 256 1476 264
rect 1484 256 1492 264
rect 1660 256 1668 264
rect 1692 256 1700 264
rect 1804 256 1812 264
rect 1964 256 1972 264
rect 1980 256 1988 264
rect 2028 256 2036 264
rect 2268 256 2276 264
rect 2316 256 2324 264
rect 2412 256 2420 264
rect 2524 276 2532 284
rect 2572 276 2580 284
rect 2652 276 2660 284
rect 2700 276 2708 284
rect 2476 256 2484 264
rect 2540 256 2548 264
rect 2604 256 2612 264
rect 2748 256 2756 264
rect 2764 256 2772 264
rect 2908 276 2916 284
rect 2972 276 2980 284
rect 3004 276 3012 284
rect 3068 276 3076 284
rect 3196 296 3204 304
rect 3244 296 3252 304
rect 3372 296 3380 304
rect 3516 296 3524 304
rect 3548 296 3556 304
rect 3660 296 3668 304
rect 3692 296 3700 304
rect 3820 296 3828 304
rect 4012 296 4020 304
rect 4060 296 4068 304
rect 4076 296 4084 304
rect 4332 296 4340 304
rect 4428 296 4436 304
rect 4508 296 4516 304
rect 4556 296 4564 304
rect 4748 296 4756 304
rect 4796 296 4804 304
rect 5004 296 5012 304
rect 3196 276 3204 284
rect 3260 276 3268 284
rect 3452 276 3460 284
rect 3500 276 3508 284
rect 3612 276 3620 284
rect 3660 276 3668 284
rect 3740 276 3748 284
rect 3804 276 3812 284
rect 3884 276 3892 284
rect 3932 276 3940 284
rect 4156 276 4164 284
rect 2860 256 2868 264
rect 2892 256 2900 264
rect 2908 256 2916 264
rect 2940 256 2948 264
rect 3068 256 3076 264
rect 3148 256 3156 264
rect 3244 256 3252 264
rect 3324 256 3332 264
rect 3340 256 3348 264
rect 3372 256 3380 264
rect 3468 256 3476 264
rect 3516 256 3524 264
rect 3740 256 3748 264
rect 3868 256 3876 264
rect 3980 256 3988 264
rect 4028 256 4036 264
rect 4060 256 4068 264
rect 4108 256 4116 264
rect 4204 276 4212 284
rect 4252 276 4260 284
rect 4380 276 4388 284
rect 4412 276 4420 284
rect 4524 276 4532 284
rect 4556 276 4564 284
rect 4620 276 4628 284
rect 4700 276 4708 284
rect 4748 276 4756 284
rect 5020 276 5028 284
rect 5052 276 5060 284
rect 5132 276 5140 284
rect 5148 276 5156 284
rect 4268 256 4276 264
rect 4300 256 4308 264
rect 4348 256 4356 264
rect 4364 256 4372 264
rect 4460 256 4468 264
rect 4476 256 4484 264
rect 4508 256 4516 264
rect 4556 256 4564 264
rect 4604 256 4612 264
rect 4652 256 4660 264
rect 4764 256 4772 264
rect 4828 256 4836 264
rect 4844 256 4852 264
rect 4892 256 4900 264
rect 4940 256 4948 264
rect 4972 256 4980 264
rect 5068 256 5076 264
rect 12 236 20 244
rect 140 236 148 244
rect 252 236 260 244
rect 284 236 292 244
rect 396 236 404 244
rect 572 236 580 244
rect 700 236 708 244
rect 796 236 804 244
rect 924 236 932 244
rect 1196 236 1204 244
rect 1276 236 1284 244
rect 1308 236 1316 244
rect 1452 236 1460 244
rect 1500 236 1508 244
rect 1580 236 1588 244
rect 1644 236 1652 244
rect 1788 236 1796 244
rect 1820 236 1828 244
rect 1884 236 1892 244
rect 1948 236 1956 244
rect 2060 236 2068 244
rect 2252 236 2260 244
rect 2396 236 2404 244
rect 2684 236 2692 244
rect 2732 236 2740 244
rect 2780 236 2788 244
rect 3004 236 3012 244
rect 3276 236 3284 244
rect 3420 236 3428 244
rect 3692 236 3700 244
rect 3724 236 3732 244
rect 3788 236 3796 244
rect 3900 236 3908 244
rect 4044 236 4052 244
rect 4124 236 4132 244
rect 4220 236 4228 244
rect 4396 236 4404 244
rect 4668 236 4676 244
rect 4812 236 4820 244
rect 5020 236 5028 244
rect 5084 236 5092 244
rect 28 176 36 184
rect 300 176 308 184
rect 348 176 356 184
rect 604 176 612 184
rect 668 176 676 184
rect 700 176 708 184
rect 972 176 980 184
rect 1132 176 1140 184
rect 1196 176 1204 184
rect 1260 176 1268 184
rect 1468 176 1476 184
rect 1612 176 1620 184
rect 1724 176 1732 184
rect 1772 176 1780 184
rect 1868 176 1876 184
rect 1932 176 1940 184
rect 2012 176 2020 184
rect 2044 176 2052 184
rect 2108 176 2116 184
rect 2140 176 2148 184
rect 2236 176 2244 184
rect 2348 176 2356 184
rect 2444 176 2452 184
rect 2492 176 2500 184
rect 2572 176 2580 184
rect 2764 176 2772 184
rect 2876 176 2884 184
rect 2924 176 2932 184
rect 2972 176 2980 184
rect 3036 176 3044 184
rect 3196 176 3204 184
rect 3276 176 3284 184
rect 3356 176 3364 184
rect 3484 176 3492 184
rect 3596 176 3604 184
rect 4092 176 4100 184
rect 4140 176 4148 184
rect 4284 176 4292 184
rect 4412 176 4420 184
rect 4508 176 4516 184
rect 4876 176 4884 184
rect 124 156 132 164
rect 140 156 148 164
rect 268 156 276 164
rect 332 156 340 164
rect 428 156 436 164
rect 444 156 452 164
rect 460 156 468 164
rect 556 156 564 164
rect 572 156 580 164
rect 732 156 740 164
rect 956 156 964 164
rect 1052 156 1060 164
rect 1084 156 1092 164
rect 1164 156 1172 164
rect 1276 156 1284 164
rect 1340 156 1348 164
rect 1356 156 1364 164
rect 1564 156 1572 164
rect 1980 156 1988 164
rect 2028 156 2036 164
rect 2092 156 2100 164
rect 2204 156 2212 164
rect 2220 156 2228 164
rect 2252 156 2260 164
rect 2380 156 2388 164
rect 2636 156 2644 164
rect 2780 156 2788 164
rect 2844 156 2852 164
rect 3436 156 3444 164
rect 3724 156 3732 164
rect 3740 156 3748 164
rect 3788 156 3796 164
rect 3852 156 3860 164
rect 3868 156 3876 164
rect 3964 156 3972 164
rect 4044 156 4052 164
rect 4108 156 4116 164
rect 4124 156 4132 164
rect 12 136 20 144
rect 124 136 132 144
rect 188 136 196 144
rect 316 136 324 144
rect 412 136 420 144
rect 492 136 500 144
rect 588 136 596 144
rect 636 136 644 144
rect 716 136 724 144
rect 780 136 788 144
rect 908 136 916 144
rect 988 136 996 144
rect 1084 136 1092 144
rect 1212 136 1220 144
rect 1228 136 1236 144
rect 1452 136 1460 144
rect 1500 136 1508 144
rect 1548 136 1556 144
rect 1596 136 1604 144
rect 1692 136 1700 144
rect 1708 136 1716 144
rect 1756 136 1764 144
rect 1852 136 1860 144
rect 1900 136 1908 144
rect 1996 136 2004 144
rect 2092 136 2100 144
rect 2172 136 2180 144
rect 2460 136 2468 144
rect 2508 136 2516 144
rect 2572 136 2580 144
rect 2652 136 2660 144
rect 2748 136 2756 144
rect 2828 136 2836 144
rect 2924 136 2932 144
rect 2956 136 2964 144
rect 3004 136 3012 144
rect 3020 136 3028 144
rect 3052 136 3060 144
rect 3164 136 3172 144
rect 3196 136 3204 144
rect 3292 136 3300 144
rect 3420 136 3428 144
rect 3500 136 3508 144
rect 3548 136 3556 144
rect 3596 136 3604 144
rect 3900 136 3908 144
rect 4156 136 4164 144
rect 92 116 100 124
rect 188 116 196 124
rect 220 116 228 124
rect 268 116 276 124
rect 764 116 772 124
rect 876 116 884 124
rect 220 96 228 104
rect 284 96 292 104
rect 380 96 388 104
rect 524 96 532 104
rect 620 96 628 104
rect 668 96 676 104
rect 684 96 692 104
rect 908 96 916 104
rect 940 96 948 104
rect 1084 116 1092 124
rect 1308 116 1316 124
rect 1180 96 1188 104
rect 1260 96 1268 104
rect 1420 96 1428 104
rect 1452 96 1460 104
rect 1516 96 1524 104
rect 1564 96 1572 104
rect 1596 96 1604 104
rect 1660 96 1668 104
rect 1740 96 1748 104
rect 1932 116 1940 124
rect 1996 116 2004 124
rect 2284 116 2292 124
rect 2412 116 2420 124
rect 2732 116 2740 124
rect 4332 156 4340 164
rect 4396 156 4404 164
rect 4428 156 4436 164
rect 4444 156 4452 164
rect 4524 156 4532 164
rect 4684 156 4692 164
rect 4764 156 4772 164
rect 4780 156 4788 164
rect 4828 156 4836 164
rect 4844 156 4852 164
rect 4860 156 4868 164
rect 4988 156 4996 164
rect 5052 156 5060 164
rect 5068 156 5076 164
rect 5164 156 5172 164
rect 5180 156 5188 164
rect 4316 136 4324 144
rect 4476 136 4484 144
rect 4556 136 4564 144
rect 4700 136 4708 144
rect 3148 116 3156 124
rect 3724 116 3732 124
rect 3772 116 3780 124
rect 3900 116 3908 124
rect 3948 116 3956 124
rect 4044 116 4052 124
rect 4076 116 4084 124
rect 4268 116 4276 124
rect 4652 116 4660 124
rect 4668 116 4676 124
rect 4908 136 4916 144
rect 4972 136 4980 144
rect 5132 136 5140 144
rect 4732 116 4740 124
rect 4780 116 4788 124
rect 4812 116 4820 124
rect 4892 116 4900 124
rect 5100 116 5108 124
rect 5148 116 5156 124
rect 1804 96 1812 104
rect 1884 96 1892 104
rect 2044 96 2052 104
rect 2124 96 2132 104
rect 2204 96 2212 104
rect 2428 96 2436 104
rect 2476 96 2484 104
rect 2556 96 2564 104
rect 2684 96 2692 104
rect 2796 96 2804 104
rect 2876 96 2884 104
rect 2972 96 2980 104
rect 3100 96 3108 104
rect 3196 96 3204 104
rect 3324 96 3332 104
rect 3388 96 3396 104
rect 3532 96 3540 104
rect 3564 96 3572 104
rect 3596 96 3604 104
rect 3644 96 3652 104
rect 4060 96 4068 104
rect 4188 96 4196 104
rect 4284 96 4292 104
rect 4396 96 4404 104
rect 4476 96 4484 104
rect 4508 96 4516 104
rect 4556 96 4564 104
rect 4588 96 4596 104
rect 4940 96 4948 104
rect 476 76 484 84
rect 780 76 788 84
rect 812 76 820 84
rect 1548 76 1556 84
rect 1932 76 1940 84
rect 1996 76 2004 84
rect 2524 76 2532 84
rect 2540 76 2548 84
rect 2860 76 2868 84
rect 2908 76 2916 84
rect 3052 76 3060 84
rect 3260 76 3268 84
rect 3500 76 3508 84
rect 3772 76 3780 84
rect 4028 76 4036 84
rect 4236 76 4244 84
rect 924 56 932 64
rect 1996 56 2004 64
rect 3148 56 3156 64
rect 1996 36 2004 44
rect 2812 36 2820 44
rect 3804 36 3812 44
rect 5020 36 5028 44
<< metal2 >>
rect 605 3544 611 3576
rect 61 3504 67 3516
rect 13 3384 19 3496
rect 45 3364 51 3476
rect 93 3344 99 3476
rect 141 3464 147 3496
rect 157 3484 163 3516
rect 237 3484 243 3516
rect 429 3504 435 3536
rect 477 3524 483 3536
rect 557 3524 563 3536
rect 340 3497 364 3503
rect 413 3484 419 3496
rect 669 3484 675 3516
rect 701 3484 707 3556
rect 749 3484 755 3496
rect 765 3477 780 3483
rect 269 3464 275 3476
rect 109 3384 115 3456
rect 109 3364 115 3376
rect 141 3324 147 3336
rect 93 3304 99 3316
rect 157 3284 163 3296
rect 45 3104 51 3236
rect 173 3124 179 3436
rect 221 3384 227 3456
rect 285 3444 291 3456
rect 365 3444 371 3476
rect 381 3464 387 3476
rect 477 3464 483 3476
rect 429 3364 435 3456
rect 461 3444 467 3456
rect 189 3224 195 3336
rect 205 3324 211 3356
rect 477 3344 483 3356
rect 388 3337 396 3343
rect 244 3297 252 3303
rect 61 3064 67 3116
rect 189 3104 195 3116
rect 173 3084 179 3096
rect 205 3063 211 3236
rect 221 3084 227 3216
rect 301 3104 307 3296
rect 333 3224 339 3336
rect 397 3304 403 3316
rect 381 3117 419 3123
rect 349 3084 355 3096
rect 228 3077 236 3083
rect 381 3083 387 3117
rect 413 3104 419 3117
rect 372 3077 387 3083
rect 317 3064 323 3076
rect 397 3064 403 3076
rect 205 3057 236 3063
rect 13 2924 19 3056
rect 45 2983 51 3056
rect 77 2984 83 2996
rect 45 2977 67 2983
rect 61 2964 67 2977
rect 45 2944 51 2956
rect 109 2944 115 3036
rect 141 3004 147 3056
rect 205 2964 211 3036
rect 13 2724 19 2836
rect 45 2803 51 2916
rect 109 2904 115 2916
rect 29 2797 51 2803
rect 29 2784 35 2797
rect 141 2724 147 2736
rect 52 2717 60 2723
rect 100 2717 108 2723
rect 157 2704 163 2956
rect 301 2924 307 3056
rect 397 3023 403 3056
rect 429 3043 435 3316
rect 445 3284 451 3296
rect 493 3284 499 3296
rect 525 3284 531 3476
rect 573 3444 579 3476
rect 541 3384 547 3436
rect 717 3424 723 3456
rect 765 3444 771 3477
rect 781 3444 787 3456
rect 573 3364 579 3376
rect 621 3364 627 3396
rect 733 3364 739 3376
rect 797 3364 803 3496
rect 813 3444 819 3683
rect 829 3504 835 3596
rect 1181 3584 1187 3596
rect 2189 3584 2195 3683
rect 2301 3624 2307 3683
rect 3261 3624 3267 3683
rect 3389 3624 3395 3683
rect 964 3557 972 3563
rect 2964 3557 3123 3563
rect 1005 3524 1011 3536
rect 1396 3517 1404 3523
rect 1309 3504 1315 3516
rect 845 3464 851 3496
rect 893 3384 899 3496
rect 973 3464 979 3476
rect 941 3443 947 3456
rect 1021 3444 1027 3456
rect 925 3437 947 3443
rect 925 3384 931 3437
rect 1037 3424 1043 3436
rect 957 3384 963 3396
rect 1053 3384 1059 3496
rect 1085 3424 1091 3456
rect 1101 3444 1107 3456
rect 1117 3404 1123 3436
rect 1133 3384 1139 3496
rect 1149 3464 1155 3496
rect 1245 3484 1251 3496
rect 1357 3484 1363 3516
rect 1453 3504 1459 3556
rect 1812 3517 1820 3523
rect 1453 3484 1459 3496
rect 1405 3464 1411 3476
rect 1485 3464 1491 3476
rect 1149 3404 1155 3456
rect 1245 3444 1251 3456
rect 1229 3384 1235 3416
rect 1293 3404 1299 3436
rect 1373 3364 1379 3436
rect 1421 3364 1427 3416
rect 1485 3384 1491 3456
rect 1501 3424 1507 3436
rect 1533 3384 1539 3476
rect 1709 3464 1715 3496
rect 1725 3484 1731 3516
rect 1917 3504 1923 3556
rect 2020 3497 2076 3503
rect 1517 3364 1523 3376
rect 1565 3364 1571 3456
rect 1613 3443 1619 3456
rect 1677 3444 1683 3456
rect 1613 3437 1635 3443
rect 1629 3384 1635 3437
rect 541 3344 547 3356
rect 717 3344 723 3356
rect 852 3337 860 3343
rect 941 3343 947 3356
rect 1037 3344 1043 3356
rect 941 3337 972 3343
rect 1220 3337 1228 3343
rect 637 3304 643 3336
rect 701 3323 707 3336
rect 765 3324 771 3336
rect 701 3317 716 3323
rect 685 3304 691 3316
rect 461 3204 467 3236
rect 797 3184 803 3336
rect 1117 3324 1123 3336
rect 868 3317 892 3323
rect 1261 3304 1267 3336
rect 1453 3324 1459 3356
rect 1469 3344 1475 3356
rect 1645 3344 1651 3416
rect 1757 3384 1763 3496
rect 1773 3424 1779 3476
rect 1821 3463 1827 3476
rect 1821 3457 1868 3463
rect 1917 3444 1923 3476
rect 2045 3464 2051 3476
rect 2173 3464 2179 3516
rect 2333 3504 2339 3516
rect 2221 3483 2227 3496
rect 2221 3477 2252 3483
rect 2381 3464 2387 3536
rect 2724 3517 2732 3523
rect 2413 3504 2419 3516
rect 2077 3444 2083 3456
rect 2157 3443 2163 3456
rect 2221 3444 2227 3456
rect 2317 3444 2323 3456
rect 2365 3444 2371 3456
rect 2413 3444 2419 3496
rect 2477 3444 2483 3496
rect 2557 3464 2563 3476
rect 2573 3464 2579 3476
rect 2509 3444 2515 3456
rect 2605 3444 2611 3516
rect 2749 3484 2755 3556
rect 3021 3537 3107 3543
rect 2845 3524 2851 3536
rect 2893 3484 2899 3536
rect 3021 3523 3027 3537
rect 2996 3517 3027 3523
rect 3037 3517 3091 3523
rect 2909 3503 2915 3516
rect 2909 3497 2931 3503
rect 2925 3484 2931 3497
rect 2772 3477 2780 3483
rect 2157 3437 2179 3443
rect 1885 3364 1891 3436
rect 1917 3384 1923 3396
rect 1732 3357 1740 3363
rect 1773 3344 1779 3356
rect 1597 3324 1603 3336
rect 900 3297 908 3303
rect 845 3264 851 3296
rect 516 3157 524 3163
rect 605 3084 611 3096
rect 461 3064 467 3076
rect 493 3043 499 3056
rect 429 3037 499 3043
rect 541 3024 547 3056
rect 557 3044 563 3056
rect 605 3044 611 3056
rect 573 3024 579 3036
rect 653 3024 659 3056
rect 669 3024 675 3036
rect 381 3017 403 3023
rect 381 2984 387 3017
rect 701 3003 707 3156
rect 733 3104 739 3116
rect 829 3084 835 3236
rect 989 3224 995 3296
rect 1181 3284 1187 3296
rect 1229 3284 1235 3296
rect 1373 3284 1379 3316
rect 1197 3244 1203 3256
rect 1316 3177 1324 3183
rect 893 3104 899 3116
rect 909 3104 915 3116
rect 989 3084 995 3096
rect 1021 3084 1027 3116
rect 1069 3104 1075 3116
rect 1165 3084 1171 3116
rect 1261 3084 1267 3116
rect 1309 3104 1315 3136
rect 1293 3084 1299 3096
rect 772 3077 780 3083
rect 733 3064 739 3076
rect 717 3044 723 3056
rect 813 3044 819 3056
rect 973 3044 979 3056
rect 685 2997 707 3003
rect 509 2984 515 2996
rect 397 2964 403 2976
rect 285 2904 291 2916
rect 285 2884 291 2896
rect 269 2803 275 2836
rect 269 2797 291 2803
rect 285 2704 291 2797
rect 301 2704 307 2836
rect 333 2764 339 2956
rect 477 2944 483 2956
rect 349 2924 355 2936
rect 525 2924 531 2976
rect 557 2964 563 2976
rect 653 2944 659 2956
rect 685 2944 691 2997
rect 429 2904 435 2916
rect 404 2897 412 2903
rect 509 2884 515 2896
rect 381 2864 387 2876
rect 461 2824 467 2836
rect 397 2704 403 2796
rect 557 2784 563 2936
rect 717 2924 723 3036
rect 765 2964 771 2976
rect 845 2964 851 2976
rect 893 2964 899 2996
rect 772 2937 787 2943
rect 605 2904 611 2916
rect 717 2864 723 2876
rect 573 2744 579 2776
rect 500 2737 508 2743
rect 13 2684 19 2696
rect 13 2524 19 2536
rect 45 2504 51 2676
rect 189 2644 195 2696
rect 205 2664 211 2676
rect 244 2657 252 2663
rect 436 2657 444 2663
rect 77 2604 83 2636
rect 125 2604 131 2636
rect 93 2524 99 2596
rect 221 2584 227 2616
rect 269 2604 275 2636
rect 333 2604 339 2656
rect 413 2644 419 2656
rect 477 2644 483 2696
rect 557 2684 563 2696
rect 509 2664 515 2676
rect 525 2664 531 2676
rect 237 2564 243 2576
rect 157 2524 163 2536
rect 237 2504 243 2556
rect 253 2524 259 2596
rect 365 2564 371 2576
rect 196 2497 204 2503
rect 13 2304 19 2316
rect 45 2284 51 2496
rect 141 2484 147 2496
rect 93 2404 99 2436
rect 157 2304 163 2476
rect 285 2404 291 2556
rect 340 2537 371 2543
rect 365 2524 371 2537
rect 324 2517 332 2523
rect 381 2464 387 2636
rect 397 2584 403 2636
rect 621 2604 627 2656
rect 429 2597 483 2603
rect 429 2564 435 2597
rect 477 2584 483 2597
rect 573 2584 579 2596
rect 461 2564 467 2576
rect 429 2504 435 2516
rect 349 2324 355 2436
rect 461 2324 467 2516
rect 493 2503 499 2556
rect 541 2524 547 2536
rect 557 2524 563 2576
rect 637 2563 643 2836
rect 653 2704 659 2816
rect 685 2804 691 2836
rect 765 2744 771 2916
rect 781 2883 787 2937
rect 829 2924 835 2936
rect 925 2924 931 3036
rect 941 2997 956 3003
rect 941 2964 947 2997
rect 1005 2984 1011 2996
rect 1021 2964 1027 3036
rect 1037 3004 1043 3076
rect 1245 3063 1251 3076
rect 1341 3064 1347 3196
rect 1364 3177 1372 3183
rect 1405 3124 1411 3236
rect 1357 3104 1363 3116
rect 1389 3064 1395 3116
rect 1437 3104 1443 3176
rect 1453 3104 1459 3276
rect 1501 3144 1507 3296
rect 1565 3264 1571 3316
rect 1661 3284 1667 3316
rect 1741 3284 1747 3296
rect 1485 3064 1491 3116
rect 1501 3084 1507 3116
rect 1245 3057 1299 3063
rect 1101 3023 1107 3056
rect 1117 3044 1123 3056
rect 1293 3043 1299 3057
rect 1405 3043 1411 3056
rect 1293 3037 1411 3043
rect 1101 3017 1123 3023
rect 1085 2984 1091 2996
rect 1117 2983 1123 3017
rect 1117 2977 1148 2983
rect 1165 2963 1171 2996
rect 1197 2964 1203 3016
rect 1277 2983 1283 3016
rect 1421 2984 1427 3036
rect 1469 3004 1475 3036
rect 1236 2977 1283 2983
rect 1444 2977 1452 2983
rect 1325 2964 1331 2976
rect 1156 2957 1171 2963
rect 957 2943 963 2956
rect 948 2937 963 2943
rect 948 2917 972 2923
rect 877 2904 883 2916
rect 989 2904 995 2956
rect 1069 2904 1075 2916
rect 1133 2904 1139 2956
rect 1293 2943 1299 2956
rect 1293 2937 1324 2943
rect 1373 2924 1379 2976
rect 1469 2964 1475 2976
rect 1181 2904 1187 2916
rect 1245 2903 1251 2916
rect 1245 2897 1260 2903
rect 813 2883 819 2896
rect 1293 2884 1299 2916
rect 1341 2884 1347 2916
rect 1421 2904 1427 2956
rect 781 2877 819 2883
rect 964 2877 972 2883
rect 708 2717 716 2723
rect 653 2664 659 2676
rect 797 2664 803 2676
rect 845 2664 851 2716
rect 749 2604 755 2636
rect 637 2557 652 2563
rect 484 2497 499 2503
rect 557 2324 563 2416
rect 589 2404 595 2556
rect 621 2424 627 2436
rect 637 2404 643 2536
rect 685 2524 691 2576
rect 717 2543 723 2576
rect 733 2564 739 2576
rect 788 2557 803 2563
rect 717 2537 739 2543
rect 708 2517 716 2523
rect 733 2503 739 2537
rect 756 2537 780 2543
rect 733 2497 755 2503
rect 749 2484 755 2497
rect 301 2304 307 2316
rect 61 2284 67 2296
rect 141 2264 147 2296
rect 61 2164 67 2176
rect 45 2144 51 2156
rect 93 2144 99 2256
rect 109 2164 115 2256
rect 173 2164 179 2176
rect 221 2164 227 2236
rect 237 2184 243 2256
rect 269 2164 275 2196
rect 285 2184 291 2296
rect 333 2244 339 2256
rect 381 2224 387 2296
rect 413 2283 419 2296
rect 413 2277 460 2283
rect 452 2257 460 2263
rect 477 2244 483 2256
rect 509 2244 515 2276
rect 653 2264 659 2276
rect 669 2264 675 2436
rect 797 2424 803 2557
rect 829 2544 835 2636
rect 893 2603 899 2656
rect 877 2597 899 2603
rect 845 2564 851 2576
rect 877 2524 883 2597
rect 925 2563 931 2776
rect 1005 2684 1011 2836
rect 1245 2803 1251 2876
rect 1325 2824 1331 2836
rect 1229 2797 1251 2803
rect 1229 2784 1235 2797
rect 1261 2744 1267 2816
rect 1053 2684 1059 2736
rect 1277 2704 1283 2716
rect 1325 2704 1331 2716
rect 957 2604 963 2676
rect 1101 2664 1107 2676
rect 1117 2643 1123 2676
rect 1133 2664 1139 2696
rect 1229 2684 1235 2696
rect 1261 2664 1267 2676
rect 1117 2637 1164 2643
rect 989 2564 995 2636
rect 1005 2564 1011 2616
rect 916 2557 931 2563
rect 1037 2524 1043 2556
rect 1085 2524 1091 2636
rect 1117 2564 1123 2576
rect 1037 2504 1043 2516
rect 1140 2497 1164 2503
rect 957 2484 963 2496
rect 685 2284 691 2316
rect 701 2304 707 2316
rect 13 1984 19 2116
rect 13 1844 19 1896
rect 45 1864 51 1876
rect 93 1864 99 2036
rect 109 2003 115 2116
rect 109 1997 131 2003
rect 13 1724 19 1836
rect 77 1824 83 1856
rect 109 1724 115 1836
rect 125 1804 131 1997
rect 189 1924 195 2156
rect 333 2124 339 2136
rect 141 1904 147 1916
rect 221 1904 227 2116
rect 365 2104 371 2116
rect 381 2064 387 2096
rect 180 1857 188 1863
rect 173 1764 179 1796
rect 221 1784 227 1856
rect 205 1744 211 1756
rect 13 1504 19 1636
rect 93 1624 99 1716
rect 221 1704 227 1756
rect 237 1744 243 2036
rect 397 1924 403 2236
rect 525 2144 531 2256
rect 541 2184 547 2256
rect 605 2244 611 2256
rect 557 2224 563 2236
rect 605 2164 611 2236
rect 637 2204 643 2256
rect 669 2224 675 2236
rect 749 2204 755 2256
rect 781 2184 787 2256
rect 621 2144 627 2156
rect 413 2124 419 2136
rect 509 2124 515 2136
rect 413 1924 419 1996
rect 429 1984 435 2116
rect 365 1904 371 1916
rect 381 1884 387 1896
rect 269 1844 275 1856
rect 333 1784 339 1836
rect 269 1704 275 1716
rect 301 1684 307 1736
rect 61 1484 67 1496
rect 45 1364 51 1456
rect 77 1403 83 1436
rect 61 1397 83 1403
rect 61 1344 67 1397
rect 109 1384 115 1436
rect 93 1344 99 1356
rect 13 1304 19 1336
rect 52 1297 60 1303
rect 93 1124 99 1316
rect 109 1164 115 1356
rect 125 1324 131 1616
rect 157 1484 163 1636
rect 189 1504 195 1516
rect 205 1504 211 1676
rect 237 1564 243 1636
rect 285 1524 291 1536
rect 237 1504 243 1516
rect 189 1344 195 1456
rect 141 1324 147 1336
rect 141 1124 147 1236
rect 205 1204 211 1356
rect 237 1344 243 1496
rect 253 1484 259 1516
rect 301 1464 307 1476
rect 317 1444 323 1756
rect 365 1744 371 1856
rect 381 1784 387 1796
rect 397 1764 403 1776
rect 413 1744 419 1836
rect 429 1784 435 1896
rect 461 1884 467 2076
rect 493 1964 499 2036
rect 525 2023 531 2136
rect 701 2124 707 2176
rect 813 2164 819 2396
rect 836 2317 844 2323
rect 877 2304 883 2476
rect 957 2437 972 2443
rect 861 2284 867 2296
rect 893 2284 899 2436
rect 909 2263 915 2276
rect 900 2257 915 2263
rect 845 2164 851 2176
rect 557 2064 563 2096
rect 525 2017 547 2023
rect 493 1924 499 1936
rect 541 1904 547 2017
rect 573 1984 579 2116
rect 653 2064 659 2096
rect 717 2023 723 2156
rect 733 2137 748 2143
rect 733 2104 739 2137
rect 749 2104 755 2116
rect 749 2044 755 2056
rect 717 2017 739 2023
rect 733 1944 739 2017
rect 749 1944 755 2036
rect 797 1984 803 2116
rect 813 1984 819 2016
rect 845 2004 851 2116
rect 637 1924 643 1936
rect 861 1924 867 2056
rect 589 1884 595 1896
rect 637 1884 643 1896
rect 653 1884 659 1896
rect 781 1884 787 1896
rect 829 1884 835 1896
rect 877 1883 883 2256
rect 925 2184 931 2296
rect 957 2264 963 2437
rect 1005 2304 1011 2416
rect 1021 2304 1027 2336
rect 1101 2304 1107 2436
rect 1165 2304 1171 2316
rect 1085 2277 1100 2283
rect 893 2164 899 2176
rect 941 2164 947 2196
rect 957 2164 963 2216
rect 973 2184 979 2196
rect 1021 2184 1027 2276
rect 1085 2263 1091 2277
rect 1076 2257 1091 2263
rect 1101 2224 1107 2256
rect 1117 2177 1148 2183
rect 1117 2164 1123 2177
rect 1165 2164 1171 2216
rect 1181 2163 1187 2656
rect 1325 2624 1331 2676
rect 1229 2597 1283 2603
rect 1229 2584 1235 2597
rect 1261 2564 1267 2576
rect 1277 2563 1283 2597
rect 1309 2564 1315 2616
rect 1373 2604 1379 2656
rect 1277 2557 1299 2563
rect 1229 2503 1235 2516
rect 1204 2497 1235 2503
rect 1245 2303 1251 2556
rect 1293 2543 1299 2557
rect 1357 2544 1363 2556
rect 1389 2544 1395 2816
rect 1437 2784 1443 2956
rect 1469 2904 1475 2916
rect 1501 2904 1507 2916
rect 1517 2784 1523 3216
rect 1581 3084 1587 3096
rect 1597 3064 1603 3236
rect 1677 3104 1683 3116
rect 1773 3104 1779 3336
rect 1821 3304 1827 3336
rect 1869 3324 1875 3336
rect 1981 3324 1987 3416
rect 2173 3384 2179 3437
rect 2669 3443 2675 3476
rect 2701 3464 2707 3476
rect 2733 3457 2764 3463
rect 2717 3443 2723 3456
rect 2733 3444 2739 3457
rect 2669 3437 2723 3443
rect 2237 3384 2243 3396
rect 2029 3284 2035 3356
rect 2125 3344 2131 3356
rect 2221 3344 2227 3356
rect 2269 3344 2275 3396
rect 2301 3384 2307 3416
rect 2349 3404 2355 3436
rect 2317 3384 2323 3396
rect 2525 3364 2531 3436
rect 2621 3384 2627 3396
rect 2356 3357 2387 3363
rect 2381 3344 2387 3357
rect 2621 3357 2668 3363
rect 2445 3324 2451 3356
rect 2109 3284 2115 3316
rect 2180 3277 2188 3283
rect 1860 3237 1868 3243
rect 1901 3224 1907 3236
rect 1949 3204 1955 3276
rect 2077 3264 2083 3276
rect 1837 3117 1939 3123
rect 1837 3104 1843 3117
rect 1933 3104 1939 3117
rect 1981 3104 1987 3216
rect 2109 3104 2115 3116
rect 1693 3097 1724 3103
rect 1629 3064 1635 3096
rect 1645 3083 1651 3096
rect 1693 3083 1699 3097
rect 2180 3097 2188 3103
rect 1645 3077 1699 3083
rect 1805 3083 1811 3096
rect 1780 3077 1811 3083
rect 1853 3064 1859 3096
rect 1917 3064 1923 3096
rect 2029 3084 2035 3096
rect 2061 3064 2067 3096
rect 2205 3064 2211 3276
rect 2221 3184 2227 3316
rect 2269 3284 2275 3316
rect 2301 3264 2307 3296
rect 2397 3284 2403 3316
rect 2509 3224 2515 3356
rect 2525 3324 2531 3356
rect 2573 3304 2579 3336
rect 2605 3324 2611 3356
rect 2621 3344 2627 3357
rect 2733 3344 2739 3396
rect 2532 3277 2540 3283
rect 2237 3104 2243 3116
rect 2221 3064 2227 3096
rect 2253 3084 2259 3176
rect 2285 3137 2355 3143
rect 2285 3104 2291 3137
rect 2301 3084 2307 3116
rect 2349 3104 2355 3137
rect 2381 3137 2499 3143
rect 2381 3104 2387 3137
rect 2493 3124 2499 3137
rect 2477 3104 2483 3116
rect 1732 3057 1756 3063
rect 1812 3057 1836 3063
rect 1933 3057 1964 3063
rect 1549 3044 1555 3056
rect 1533 2884 1539 2956
rect 1597 2944 1603 2956
rect 1597 2904 1603 2916
rect 1453 2724 1459 2736
rect 1597 2724 1603 2836
rect 1613 2824 1619 3036
rect 1629 2924 1635 2936
rect 1645 2904 1651 2916
rect 1677 2904 1683 2956
rect 1693 2923 1699 3056
rect 1709 2984 1715 3016
rect 1773 2944 1779 3056
rect 1885 3043 1891 3056
rect 1933 3043 1939 3057
rect 1885 3037 1939 3043
rect 2093 3004 2099 3056
rect 2141 3004 2147 3056
rect 1869 2977 1955 2983
rect 1869 2963 1875 2977
rect 1805 2957 1875 2963
rect 1693 2917 1715 2923
rect 1709 2844 1715 2917
rect 1725 2864 1731 2936
rect 1725 2784 1731 2816
rect 1517 2704 1523 2716
rect 1405 2584 1411 2696
rect 1693 2684 1699 2776
rect 1741 2704 1747 2936
rect 1805 2904 1811 2957
rect 1892 2957 1939 2963
rect 1933 2944 1939 2957
rect 1949 2943 1955 2977
rect 1965 2964 1971 2996
rect 2029 2964 2035 2996
rect 2045 2957 2099 2963
rect 1949 2937 1964 2943
rect 2045 2943 2051 2957
rect 2093 2944 2099 2957
rect 2036 2937 2051 2943
rect 1821 2884 1827 2936
rect 1837 2904 1843 2936
rect 1917 2924 1923 2936
rect 2061 2924 2067 2936
rect 2077 2924 2083 2936
rect 2157 2924 2163 3036
rect 2253 2983 2259 3076
rect 2381 3064 2387 3076
rect 2356 3057 2371 3063
rect 2365 3043 2371 3057
rect 2397 3044 2403 3096
rect 2541 3084 2547 3196
rect 2596 3137 2620 3143
rect 2621 3084 2627 3096
rect 2429 3064 2435 3076
rect 2525 3063 2531 3076
rect 2525 3057 2547 3063
rect 2445 3044 2451 3056
rect 2541 3044 2547 3057
rect 2621 3044 2627 3076
rect 2365 3037 2387 3043
rect 2381 3023 2387 3037
rect 2461 3023 2467 3036
rect 2381 3017 2467 3023
rect 2397 2997 2515 3003
rect 2253 2977 2268 2983
rect 2212 2957 2236 2963
rect 2324 2957 2348 2963
rect 2381 2943 2387 2956
rect 2397 2944 2403 2997
rect 2509 2984 2515 2997
rect 2525 2983 2531 3036
rect 2573 3004 2579 3036
rect 2525 2977 2556 2983
rect 2477 2944 2483 2956
rect 2260 2937 2387 2943
rect 2445 2924 2451 2936
rect 2356 2917 2396 2923
rect 1853 2883 1859 2916
rect 1837 2877 1859 2883
rect 1789 2824 1795 2876
rect 1805 2863 1811 2876
rect 1837 2863 1843 2877
rect 1805 2857 1843 2863
rect 1885 2863 1891 2916
rect 1917 2904 1923 2916
rect 1933 2884 1939 2916
rect 2013 2884 2019 2916
rect 2109 2904 2115 2916
rect 2301 2884 2307 2916
rect 2429 2884 2435 2916
rect 2445 2904 2451 2916
rect 2372 2877 2380 2883
rect 1885 2857 1948 2863
rect 1469 2624 1475 2656
rect 1549 2624 1555 2656
rect 1565 2644 1571 2676
rect 1645 2644 1651 2656
rect 1581 2624 1587 2636
rect 1629 2584 1635 2616
rect 1677 2603 1683 2636
rect 1709 2604 1715 2696
rect 1821 2664 1827 2816
rect 1917 2784 1923 2816
rect 2068 2777 2076 2783
rect 1892 2737 1900 2743
rect 1997 2724 2003 2736
rect 1933 2717 1987 2723
rect 1901 2704 1907 2716
rect 1933 2683 1939 2717
rect 1981 2703 1987 2717
rect 2045 2723 2051 2736
rect 2029 2717 2051 2723
rect 2029 2703 2035 2717
rect 1981 2697 2035 2703
rect 1949 2684 1955 2696
rect 1869 2677 1939 2683
rect 1869 2664 1875 2677
rect 1677 2597 1699 2603
rect 1476 2577 1571 2583
rect 1565 2564 1571 2577
rect 1405 2557 1484 2563
rect 1405 2544 1411 2557
rect 1293 2537 1308 2543
rect 1332 2537 1347 2543
rect 1341 2524 1347 2537
rect 1357 2517 1427 2523
rect 1277 2503 1283 2516
rect 1357 2503 1363 2517
rect 1421 2504 1427 2517
rect 1277 2497 1363 2503
rect 1405 2464 1411 2496
rect 1261 2344 1267 2416
rect 1325 2404 1331 2436
rect 1437 2384 1443 2516
rect 1501 2484 1507 2556
rect 1533 2484 1539 2556
rect 1556 2457 1564 2463
rect 1517 2424 1523 2436
rect 1581 2384 1587 2516
rect 1645 2484 1651 2496
rect 1661 2444 1667 2556
rect 1693 2524 1699 2597
rect 1709 2504 1715 2556
rect 1661 2384 1667 2396
rect 1277 2304 1283 2336
rect 1341 2324 1347 2336
rect 1357 2304 1363 2336
rect 1453 2317 1468 2323
rect 1453 2304 1459 2317
rect 1645 2304 1651 2336
rect 1677 2304 1683 2316
rect 1725 2304 1731 2576
rect 1741 2504 1747 2656
rect 1773 2644 1779 2656
rect 1853 2644 1859 2656
rect 1933 2624 1939 2656
rect 1949 2584 1955 2616
rect 1981 2564 1987 2656
rect 2061 2644 2067 2656
rect 1997 2624 2003 2636
rect 2093 2604 2099 2656
rect 2109 2624 2115 2676
rect 2125 2603 2131 2856
rect 2269 2824 2275 2876
rect 2301 2784 2307 2816
rect 2148 2737 2156 2743
rect 2189 2703 2195 2716
rect 2164 2697 2195 2703
rect 2269 2703 2275 2716
rect 2244 2697 2275 2703
rect 2157 2624 2163 2676
rect 2109 2597 2131 2603
rect 2077 2584 2083 2596
rect 2029 2564 2035 2576
rect 1796 2557 1804 2563
rect 1828 2557 1836 2563
rect 2052 2557 2060 2563
rect 1789 2484 1795 2516
rect 1821 2484 1827 2496
rect 1837 2464 1843 2516
rect 1869 2444 1875 2516
rect 1741 2304 1747 2316
rect 1757 2304 1763 2436
rect 1869 2363 1875 2396
rect 1965 2383 1971 2536
rect 1981 2504 1987 2516
rect 2013 2444 2019 2556
rect 2061 2504 2067 2516
rect 2077 2504 2083 2556
rect 2109 2544 2115 2597
rect 2189 2564 2195 2636
rect 2205 2624 2211 2676
rect 2269 2624 2275 2656
rect 2317 2644 2323 2676
rect 2381 2624 2387 2676
rect 2413 2664 2419 2716
rect 2397 2604 2403 2636
rect 2237 2584 2243 2596
rect 2429 2584 2435 2656
rect 2445 2624 2451 2836
rect 2493 2744 2499 2956
rect 2525 2944 2531 2956
rect 2541 2924 2547 2956
rect 2637 2904 2643 2996
rect 2653 2964 2659 3336
rect 2749 3324 2755 3436
rect 2813 3424 2819 3436
rect 2909 3404 2915 3436
rect 2973 3424 2979 3516
rect 3037 3484 3043 3517
rect 3085 3504 3091 3517
rect 3101 3503 3107 3537
rect 3117 3524 3123 3557
rect 3341 3557 3539 3563
rect 3309 3544 3315 3556
rect 3261 3537 3299 3543
rect 3133 3517 3212 3523
rect 3133 3503 3139 3517
rect 3261 3523 3267 3537
rect 3236 3517 3267 3523
rect 3293 3523 3299 3537
rect 3341 3523 3347 3557
rect 3293 3517 3347 3523
rect 3277 3504 3283 3516
rect 3101 3497 3139 3503
rect 3069 3484 3075 3496
rect 3021 3457 3036 3463
rect 3005 3404 3011 3436
rect 3021 3384 3027 3457
rect 3053 3463 3059 3476
rect 3101 3463 3107 3476
rect 3053 3457 3107 3463
rect 3053 3424 3059 3436
rect 3101 3384 3107 3396
rect 2884 3357 2892 3363
rect 2829 3343 2835 3356
rect 3069 3344 3075 3376
rect 3085 3344 3091 3356
rect 2829 3337 2876 3343
rect 2941 3324 2947 3336
rect 2749 3304 2755 3316
rect 2765 3304 2771 3316
rect 2925 3304 2931 3316
rect 3037 3304 3043 3336
rect 2989 3264 2995 3276
rect 2733 3184 2739 3236
rect 2797 3124 2803 3136
rect 2717 3084 2723 3116
rect 2685 3064 2691 3076
rect 2749 3064 2755 3076
rect 2797 3064 2803 3076
rect 2669 2964 2675 3056
rect 2813 3043 2819 3056
rect 2724 3037 2819 3043
rect 2749 2984 2755 2996
rect 2573 2864 2579 2896
rect 2589 2744 2595 2876
rect 2621 2864 2627 2896
rect 2669 2884 2675 2916
rect 2500 2677 2515 2683
rect 2493 2644 2499 2656
rect 2477 2584 2483 2616
rect 2509 2603 2515 2677
rect 2541 2604 2547 2696
rect 2605 2663 2611 2716
rect 2605 2657 2627 2663
rect 2509 2597 2531 2603
rect 2301 2577 2355 2583
rect 2164 2557 2172 2563
rect 2301 2563 2307 2577
rect 2349 2564 2355 2577
rect 2525 2583 2531 2597
rect 2557 2597 2595 2603
rect 2557 2583 2563 2597
rect 2525 2577 2563 2583
rect 2397 2564 2403 2576
rect 2276 2557 2307 2563
rect 2221 2504 2227 2516
rect 2253 2464 2259 2556
rect 2381 2523 2387 2556
rect 2397 2544 2403 2556
rect 2413 2523 2419 2576
rect 2381 2517 2419 2523
rect 2461 2523 2467 2576
rect 2509 2564 2515 2576
rect 2589 2564 2595 2597
rect 2541 2557 2579 2563
rect 2500 2537 2508 2543
rect 2541 2543 2547 2557
rect 2525 2537 2547 2543
rect 2525 2523 2531 2537
rect 2557 2524 2563 2536
rect 2461 2517 2531 2523
rect 2573 2523 2579 2557
rect 2605 2543 2611 2636
rect 2621 2564 2627 2657
rect 2637 2644 2643 2876
rect 2653 2664 2659 2816
rect 2669 2744 2675 2856
rect 2717 2744 2723 2816
rect 2701 2704 2707 2736
rect 2733 2683 2739 2956
rect 2765 2924 2771 2956
rect 2781 2924 2787 2956
rect 2717 2677 2739 2683
rect 2701 2644 2707 2676
rect 2669 2584 2675 2636
rect 2717 2564 2723 2677
rect 2749 2663 2755 2716
rect 2765 2684 2771 2816
rect 2797 2744 2803 2816
rect 2813 2744 2819 2956
rect 2829 2744 2835 3176
rect 2845 3084 2851 3096
rect 2909 3084 2915 3096
rect 2893 2964 2899 2996
rect 2925 2984 2931 3136
rect 2957 3123 2963 3216
rect 2989 3144 2995 3236
rect 3021 3164 3027 3256
rect 3037 3184 3043 3196
rect 3069 3144 3075 3336
rect 2941 3117 2963 3123
rect 2941 3104 2947 3117
rect 3021 3104 3027 3136
rect 3037 3084 3043 3136
rect 3085 3124 3091 3316
rect 3117 3303 3123 3436
rect 3133 3404 3139 3456
rect 3165 3364 3171 3496
rect 3357 3484 3363 3536
rect 3389 3497 3459 3503
rect 3284 3477 3331 3483
rect 3197 3424 3203 3436
rect 3213 3404 3219 3476
rect 3325 3444 3331 3477
rect 3389 3483 3395 3497
rect 3453 3484 3459 3497
rect 3380 3477 3395 3483
rect 3485 3483 3491 3496
rect 3476 3477 3491 3483
rect 3405 3444 3411 3476
rect 3517 3464 3523 3516
rect 3533 3464 3539 3557
rect 3645 3524 3651 3596
rect 3668 3577 3676 3583
rect 3620 3517 3635 3523
rect 3572 3497 3619 3503
rect 3549 3444 3555 3476
rect 3565 3463 3571 3476
rect 3597 3464 3603 3476
rect 3613 3464 3619 3497
rect 3565 3457 3587 3463
rect 3581 3443 3587 3457
rect 3629 3463 3635 3517
rect 3645 3484 3651 3516
rect 3693 3484 3699 3576
rect 3741 3484 3747 3516
rect 3789 3484 3795 3576
rect 3853 3484 3859 3516
rect 3885 3484 3891 3576
rect 3901 3484 3907 3516
rect 3949 3484 3955 3516
rect 3981 3484 3987 3496
rect 3997 3484 4003 3516
rect 4029 3484 4035 3596
rect 4061 3517 4076 3523
rect 4045 3484 4051 3516
rect 3924 3477 3932 3483
rect 3629 3457 3644 3463
rect 3581 3437 3612 3443
rect 3133 3304 3139 3316
rect 3101 3297 3123 3303
rect 2973 3064 2979 3076
rect 3069 3064 3075 3096
rect 2989 3024 2995 3036
rect 3101 3024 3107 3297
rect 3149 3303 3155 3356
rect 3165 3324 3171 3336
rect 3181 3303 3187 3396
rect 3229 3384 3235 3416
rect 3245 3404 3251 3436
rect 3389 3404 3395 3436
rect 3261 3364 3267 3376
rect 3149 3297 3187 3303
rect 3117 3204 3123 3276
rect 3197 3264 3203 3356
rect 3309 3304 3315 3356
rect 3341 3344 3347 3356
rect 3357 3344 3363 3376
rect 3501 3364 3507 3436
rect 3405 3344 3411 3356
rect 3485 3344 3491 3356
rect 3437 3324 3443 3336
rect 3533 3324 3539 3436
rect 3549 3384 3555 3396
rect 3565 3364 3571 3436
rect 3725 3404 3731 3436
rect 3709 3383 3715 3396
rect 3741 3384 3747 3476
rect 3965 3463 3971 3476
rect 4061 3463 4067 3517
rect 4141 3484 4147 3576
rect 4173 3544 4179 3683
rect 4333 3604 4339 3683
rect 3965 3457 4067 3463
rect 3757 3424 3763 3436
rect 3805 3384 3811 3396
rect 3709 3377 3731 3383
rect 3245 3264 3251 3296
rect 3389 3264 3395 3296
rect 3485 3264 3491 3296
rect 3284 3257 3292 3263
rect 3437 3224 3443 3236
rect 3133 3184 3139 3216
rect 3117 3084 3123 3176
rect 3245 3144 3251 3216
rect 3165 3044 3171 3116
rect 3293 3084 3299 3096
rect 3309 3084 3315 3116
rect 3453 3104 3459 3116
rect 2957 2964 2963 2996
rect 2893 2704 2899 2916
rect 2941 2884 2947 2956
rect 2989 2924 2995 2996
rect 3117 2977 3155 2983
rect 3117 2963 3123 2977
rect 3085 2957 3123 2963
rect 3044 2937 3052 2943
rect 3021 2923 3027 2936
rect 3085 2924 3091 2957
rect 3133 2924 3139 2956
rect 3149 2944 3155 2977
rect 3197 2963 3203 3076
rect 3213 3064 3219 3076
rect 3213 2984 3219 3016
rect 3261 2984 3267 3056
rect 3293 3044 3299 3076
rect 3341 3064 3347 3076
rect 3389 3064 3395 3076
rect 3197 2957 3235 2963
rect 3229 2944 3235 2957
rect 3293 2944 3299 2956
rect 3325 2944 3331 3036
rect 3405 3003 3411 3096
rect 3453 3064 3459 3096
rect 3501 3084 3507 3316
rect 3549 3303 3555 3356
rect 3565 3324 3571 3336
rect 3668 3317 3676 3323
rect 3540 3297 3555 3303
rect 3725 3303 3731 3377
rect 3837 3364 3843 3436
rect 3901 3424 3907 3436
rect 3949 3364 3955 3436
rect 3997 3364 4003 3436
rect 4093 3424 4099 3476
rect 4109 3404 4115 3436
rect 4173 3424 4179 3536
rect 4333 3524 4339 3596
rect 4509 3584 4515 3683
rect 4797 3624 4803 3683
rect 4189 3517 4220 3523
rect 4189 3504 4195 3517
rect 4244 3497 4268 3503
rect 4317 3484 4323 3516
rect 4429 3484 4435 3536
rect 4477 3484 4483 3496
rect 4509 3484 4515 3576
rect 4557 3484 4563 3496
rect 4605 3484 4611 3496
rect 4621 3484 4627 3496
rect 4653 3484 4659 3596
rect 4749 3544 4755 3616
rect 4877 3604 4883 3683
rect 4749 3504 4755 3536
rect 4244 3477 4259 3483
rect 4253 3464 4259 3477
rect 4388 3477 4396 3483
rect 4196 3437 4204 3443
rect 4077 3364 4083 3396
rect 4157 3384 4163 3396
rect 4269 3384 4275 3476
rect 4365 3464 4371 3476
rect 4333 3404 4339 3436
rect 3917 3357 3932 3363
rect 3741 3324 3747 3336
rect 3757 3324 3763 3356
rect 3853 3344 3859 3356
rect 3917 3344 3923 3357
rect 4020 3357 4028 3363
rect 4052 3357 4060 3363
rect 4093 3344 4099 3356
rect 3789 3317 3827 3323
rect 3789 3303 3795 3317
rect 3821 3304 3827 3317
rect 3725 3297 3795 3303
rect 3613 3284 3619 3296
rect 3517 3164 3523 3236
rect 3773 3204 3779 3236
rect 3837 3204 3843 3316
rect 3853 3284 3859 3296
rect 3565 3137 3596 3143
rect 3533 3124 3539 3136
rect 3565 3124 3571 3137
rect 3693 3124 3699 3156
rect 3581 3104 3587 3116
rect 3645 3104 3651 3116
rect 3524 3057 3532 3063
rect 3437 3044 3443 3056
rect 3485 3044 3491 3056
rect 3549 3044 3555 3056
rect 3533 3017 3571 3023
rect 3533 3004 3539 3017
rect 3389 2997 3411 3003
rect 3389 2964 3395 2997
rect 3485 2984 3491 2996
rect 3460 2977 3468 2983
rect 3501 2964 3507 2976
rect 3341 2944 3347 2956
rect 3181 2924 3187 2936
rect 3021 2917 3036 2923
rect 3101 2904 3107 2916
rect 3245 2904 3251 2916
rect 3028 2897 3036 2903
rect 3188 2897 3196 2903
rect 2957 2784 2963 2816
rect 2989 2804 2995 2836
rect 3037 2784 3043 2796
rect 3053 2744 3059 2896
rect 3085 2784 3091 2796
rect 2845 2684 2851 2696
rect 2781 2677 2796 2683
rect 2781 2663 2787 2677
rect 2861 2664 2867 2696
rect 2749 2657 2787 2663
rect 2893 2644 2899 2656
rect 2733 2564 2739 2576
rect 2749 2564 2755 2636
rect 2829 2564 2835 2576
rect 2653 2557 2684 2563
rect 2596 2537 2611 2543
rect 2653 2523 2659 2557
rect 2804 2557 2812 2563
rect 2573 2517 2659 2523
rect 2301 2504 2307 2516
rect 2349 2504 2355 2516
rect 2541 2504 2547 2516
rect 2276 2497 2284 2503
rect 2365 2484 2371 2496
rect 2413 2484 2419 2496
rect 1956 2377 1971 2383
rect 1981 2417 2051 2423
rect 1981 2363 1987 2417
rect 2045 2383 2051 2417
rect 2301 2417 2355 2423
rect 2045 2377 2067 2383
rect 1869 2357 1987 2363
rect 2061 2363 2067 2377
rect 2301 2364 2307 2417
rect 2349 2404 2355 2417
rect 2333 2384 2339 2396
rect 2061 2357 2236 2363
rect 1245 2297 1267 2303
rect 1229 2263 1235 2296
rect 1204 2257 1235 2263
rect 1245 2204 1251 2256
rect 1229 2164 1235 2196
rect 1181 2157 1203 2163
rect 1133 2144 1139 2156
rect 941 2124 947 2136
rect 893 1904 899 2116
rect 989 2083 995 2116
rect 1005 2104 1011 2116
rect 989 2077 1011 2083
rect 916 1957 924 1963
rect 941 1904 947 2076
rect 1005 1984 1011 2077
rect 1037 2064 1043 2136
rect 1197 2123 1203 2157
rect 1213 2144 1219 2156
rect 1261 2143 1267 2297
rect 1293 2263 1299 2296
rect 1293 2257 1308 2263
rect 1341 2244 1347 2296
rect 1405 2263 1411 2276
rect 1469 2264 1475 2296
rect 1533 2264 1539 2296
rect 1613 2264 1619 2296
rect 1645 2264 1651 2296
rect 1405 2257 1443 2263
rect 1437 2244 1443 2257
rect 1517 2244 1523 2256
rect 1565 2244 1571 2256
rect 1229 2137 1267 2143
rect 1277 2143 1283 2196
rect 1389 2184 1395 2196
rect 1421 2164 1427 2236
rect 1629 2223 1635 2236
rect 1565 2217 1603 2223
rect 1629 2217 1651 2223
rect 1533 2184 1539 2196
rect 1565 2164 1571 2217
rect 1597 2203 1603 2217
rect 1597 2197 1628 2203
rect 1348 2157 1356 2163
rect 1469 2144 1475 2156
rect 1277 2137 1299 2143
rect 1197 2117 1212 2123
rect 1181 2104 1187 2116
rect 1092 2097 1100 2103
rect 1197 2024 1203 2036
rect 861 1877 883 1883
rect 461 1804 467 1876
rect 541 1764 547 1876
rect 484 1757 508 1763
rect 589 1744 595 1876
rect 605 1864 611 1876
rect 653 1784 659 1876
rect 733 1784 739 1856
rect 749 1804 755 1836
rect 765 1784 771 1796
rect 861 1783 867 1877
rect 893 1864 899 1896
rect 973 1864 979 1956
rect 1021 1924 1027 1996
rect 1149 1984 1155 2016
rect 1229 2003 1235 2137
rect 1197 1997 1235 2003
rect 1197 1984 1203 1997
rect 1261 1964 1267 2116
rect 1277 2004 1283 2096
rect 1293 1983 1299 2137
rect 1341 2137 1356 2143
rect 1284 1977 1299 1983
rect 1261 1904 1267 1916
rect 1021 1877 1059 1883
rect 877 1843 883 1856
rect 1021 1843 1027 1877
rect 877 1837 1027 1843
rect 829 1777 867 1783
rect 605 1764 611 1776
rect 829 1764 835 1777
rect 1037 1764 1043 1856
rect 1053 1844 1059 1877
rect 1069 1864 1075 1896
rect 1149 1857 1164 1863
rect 605 1744 611 1756
rect 733 1744 739 1756
rect 349 1704 355 1716
rect 365 1684 371 1716
rect 397 1504 403 1736
rect 413 1704 419 1716
rect 445 1603 451 1736
rect 461 1704 467 1736
rect 749 1724 755 1756
rect 781 1724 787 1756
rect 925 1744 931 1756
rect 1069 1744 1075 1856
rect 1117 1844 1123 1856
rect 1117 1764 1123 1776
rect 1101 1737 1116 1743
rect 429 1597 451 1603
rect 429 1504 435 1597
rect 461 1483 467 1696
rect 541 1684 547 1716
rect 477 1584 483 1676
rect 605 1664 611 1716
rect 637 1684 643 1696
rect 829 1683 835 1716
rect 829 1677 851 1683
rect 484 1497 499 1503
rect 461 1477 483 1483
rect 445 1457 460 1463
rect 253 1324 259 1376
rect 285 1324 291 1436
rect 365 1424 371 1436
rect 365 1384 371 1396
rect 381 1324 387 1396
rect 413 1384 419 1416
rect 429 1364 435 1456
rect 445 1384 451 1457
rect 477 1443 483 1477
rect 461 1437 483 1443
rect 461 1384 467 1437
rect 493 1424 499 1497
rect 557 1484 563 1516
rect 653 1504 659 1636
rect 797 1624 803 1636
rect 685 1584 691 1596
rect 845 1584 851 1677
rect 733 1504 739 1536
rect 877 1524 883 1736
rect 893 1704 899 1736
rect 781 1504 787 1516
rect 829 1504 835 1516
rect 861 1484 867 1496
rect 557 1464 563 1476
rect 541 1444 547 1456
rect 173 1184 179 1196
rect 333 1184 339 1256
rect 205 1124 211 1136
rect 13 1084 19 1096
rect 109 1084 115 1096
rect 61 1064 67 1076
rect 36 1057 44 1063
rect 29 984 35 996
rect 13 924 19 936
rect 45 904 51 1036
rect 61 984 67 1016
rect 109 944 115 1076
rect 125 984 131 996
rect 141 964 147 1036
rect 157 1004 163 1096
rect 237 1084 243 1136
rect 381 1124 387 1216
rect 253 1004 259 1096
rect 397 1063 403 1316
rect 413 1084 419 1196
rect 429 1124 435 1336
rect 445 1304 451 1316
rect 477 1244 483 1336
rect 493 1324 499 1336
rect 509 1324 515 1356
rect 557 1344 563 1416
rect 589 1364 595 1476
rect 765 1464 771 1476
rect 653 1444 659 1456
rect 605 1384 611 1396
rect 621 1324 627 1356
rect 653 1324 659 1356
rect 669 1344 675 1356
rect 525 1264 531 1296
rect 461 1224 467 1236
rect 541 1184 547 1216
rect 557 1124 563 1276
rect 685 1224 691 1436
rect 765 1364 771 1376
rect 781 1364 787 1456
rect 717 1224 723 1336
rect 733 1264 739 1316
rect 765 1184 771 1336
rect 797 1184 803 1356
rect 813 1344 819 1456
rect 829 1364 835 1436
rect 909 1384 915 1456
rect 893 1344 899 1356
rect 845 1324 851 1336
rect 877 1304 883 1316
rect 653 1124 659 1136
rect 461 1084 467 1116
rect 509 1084 515 1116
rect 525 1084 531 1096
rect 397 1057 419 1063
rect 189 984 195 996
rect 365 983 371 1056
rect 413 984 419 1057
rect 429 1044 435 1076
rect 365 977 387 983
rect 205 964 211 976
rect 260 957 268 963
rect 285 944 291 956
rect 141 924 147 936
rect 61 764 67 896
rect 157 804 163 936
rect 237 904 243 916
rect 45 724 51 756
rect 141 724 147 736
rect 13 684 19 696
rect 173 684 179 856
rect 253 764 259 896
rect 301 864 307 936
rect 349 904 355 936
rect 333 884 339 896
rect 349 804 355 896
rect 381 844 387 977
rect 189 724 195 736
rect 269 724 275 736
rect 317 724 323 796
rect 237 684 243 716
rect 285 684 291 716
rect 365 704 371 836
rect 397 823 403 936
rect 429 924 435 1036
rect 477 964 483 1036
rect 509 984 515 1056
rect 653 984 659 996
rect 701 984 707 1096
rect 797 1084 803 1096
rect 813 1084 819 1236
rect 845 1184 851 1216
rect 733 1024 739 1036
rect 445 944 451 956
rect 525 944 531 976
rect 541 944 547 956
rect 621 944 627 956
rect 573 924 579 936
rect 717 924 723 936
rect 397 817 419 823
rect 381 724 387 736
rect 413 684 419 817
rect 445 803 451 916
rect 525 904 531 916
rect 685 884 691 896
rect 445 797 467 803
rect 436 777 444 783
rect 429 664 435 696
rect 461 664 467 797
rect 477 763 483 876
rect 477 757 499 763
rect 477 724 483 736
rect 125 644 131 656
rect 381 644 387 656
rect 333 637 348 643
rect 29 603 35 636
rect 13 597 35 603
rect 13 564 19 597
rect 77 523 83 636
rect 141 583 147 636
rect 125 577 147 583
rect 77 517 92 523
rect 13 144 19 236
rect 29 184 35 416
rect 125 304 131 577
rect 141 524 147 556
rect 189 544 195 636
rect 205 584 211 616
rect 221 564 227 576
rect 269 564 275 636
rect 237 524 243 536
rect 333 524 339 637
rect 349 584 355 616
rect 381 524 387 636
rect 445 584 451 596
rect 477 564 483 636
rect 493 604 499 757
rect 749 723 755 976
rect 829 963 835 1156
rect 845 1064 851 1116
rect 861 1084 867 1216
rect 893 1104 899 1116
rect 925 1064 931 1656
rect 973 1584 979 1736
rect 989 1704 995 1736
rect 941 1484 947 1536
rect 1021 1524 1027 1676
rect 1085 1544 1091 1716
rect 1101 1704 1107 1737
rect 1117 1704 1123 1716
rect 1149 1584 1155 1857
rect 1181 1843 1187 1876
rect 1165 1837 1187 1843
rect 1165 1724 1171 1837
rect 1197 1784 1203 1796
rect 1261 1784 1267 1896
rect 1293 1864 1299 1896
rect 1309 1884 1315 2116
rect 1341 2104 1347 2137
rect 1357 2104 1363 2116
rect 1517 2064 1523 2096
rect 1549 2044 1555 2136
rect 1565 2064 1571 2116
rect 1389 1924 1395 1996
rect 1341 1904 1347 1916
rect 1357 1883 1363 1896
rect 1421 1884 1427 2036
rect 1437 1904 1443 1916
rect 1325 1877 1363 1883
rect 1325 1864 1331 1877
rect 1469 1864 1475 1956
rect 1508 1897 1523 1903
rect 1517 1883 1523 1897
rect 1517 1877 1548 1883
rect 1412 1857 1427 1863
rect 1293 1844 1299 1856
rect 1373 1824 1379 1856
rect 1213 1777 1251 1783
rect 1213 1763 1219 1777
rect 1245 1764 1251 1777
rect 1277 1764 1283 1796
rect 1188 1757 1219 1763
rect 1229 1744 1235 1756
rect 1165 1704 1171 1716
rect 1213 1704 1219 1716
rect 1197 1543 1203 1556
rect 1117 1537 1203 1543
rect 1053 1524 1059 1536
rect 1117 1524 1123 1537
rect 996 1517 1004 1523
rect 1133 1504 1139 1516
rect 1229 1504 1235 1736
rect 1293 1724 1299 1756
rect 1309 1744 1315 1776
rect 1325 1764 1331 1776
rect 1341 1724 1347 1776
rect 1389 1744 1395 1756
rect 1405 1744 1411 1836
rect 1421 1764 1427 1857
rect 1549 1844 1555 1856
rect 1485 1784 1491 1816
rect 1501 1764 1507 1836
rect 1565 1824 1571 1896
rect 1261 1704 1267 1716
rect 1309 1703 1315 1716
rect 1453 1704 1459 1716
rect 1293 1697 1315 1703
rect 1293 1684 1299 1697
rect 1517 1703 1523 1816
rect 1581 1783 1587 2196
rect 1645 2183 1651 2217
rect 1613 2177 1651 2183
rect 1597 2124 1603 2156
rect 1613 2144 1619 2177
rect 1645 2144 1651 2156
rect 1645 2084 1651 2116
rect 1677 2064 1683 2256
rect 1709 2123 1715 2156
rect 1693 2117 1715 2123
rect 1620 2057 1628 2063
rect 1693 2003 1699 2117
rect 1709 2024 1715 2096
rect 1725 2023 1731 2256
rect 1757 2164 1763 2196
rect 1773 2184 1779 2276
rect 1789 2264 1795 2296
rect 1837 2283 1843 2296
rect 1837 2277 1859 2283
rect 1853 2244 1859 2277
rect 1837 2203 1843 2216
rect 1837 2197 1859 2203
rect 1789 2164 1795 2196
rect 1853 2164 1859 2197
rect 1741 2144 1747 2156
rect 1805 2144 1811 2156
rect 1869 2143 1875 2276
rect 1885 2264 1891 2276
rect 1885 2164 1891 2216
rect 1853 2137 1875 2143
rect 1741 2064 1747 2116
rect 1837 2084 1843 2096
rect 1725 2017 1795 2023
rect 1693 1997 1779 2003
rect 1773 1984 1779 1997
rect 1789 1983 1795 2017
rect 1789 1977 1836 1983
rect 1853 1964 1859 2137
rect 1901 2084 1907 2096
rect 1869 1997 1907 2003
rect 1869 1984 1875 1997
rect 1901 1944 1907 1997
rect 1860 1917 1868 1923
rect 1917 1923 1923 2296
rect 1965 2284 1971 2316
rect 2045 2284 2051 2356
rect 2157 2317 2195 2323
rect 2077 2304 2083 2316
rect 2157 2304 2163 2317
rect 2189 2304 2195 2317
rect 2317 2304 2323 2316
rect 2125 2284 2131 2296
rect 2173 2284 2179 2296
rect 2221 2284 2227 2296
rect 2365 2284 2371 2316
rect 2397 2284 2403 2416
rect 2429 2404 2435 2436
rect 2445 2424 2451 2476
rect 2413 2383 2419 2396
rect 2445 2383 2451 2396
rect 2541 2384 2547 2396
rect 2413 2377 2451 2383
rect 2413 2304 2419 2316
rect 2477 2304 2483 2316
rect 2452 2297 2460 2303
rect 1933 2243 1939 2256
rect 2029 2244 2035 2256
rect 1933 2237 1955 2243
rect 1933 2144 1939 2216
rect 1949 2184 1955 2237
rect 1981 2224 1987 2236
rect 2077 2204 2083 2276
rect 2093 2224 2099 2256
rect 2109 2164 2115 2196
rect 2029 2144 2035 2156
rect 2061 2144 2067 2156
rect 1981 2124 1987 2136
rect 2004 2117 2028 2123
rect 2077 2117 2108 2123
rect 2061 2064 2067 2116
rect 2077 2084 2083 2117
rect 2125 2103 2131 2256
rect 2205 2224 2211 2236
rect 2221 2224 2227 2256
rect 2269 2203 2275 2256
rect 2285 2224 2291 2256
rect 2349 2244 2355 2256
rect 2381 2224 2387 2236
rect 2269 2197 2291 2203
rect 2157 2177 2220 2183
rect 2157 2164 2163 2177
rect 2109 2097 2131 2103
rect 2013 1984 2019 2056
rect 2045 2043 2051 2056
rect 2045 2037 2076 2043
rect 2109 1943 2115 2097
rect 2141 2024 2147 2036
rect 2125 1984 2131 2016
rect 2093 1937 2115 1943
rect 1901 1917 1923 1923
rect 1677 1904 1683 1916
rect 1604 1897 1612 1903
rect 1741 1884 1747 1916
rect 1821 1904 1827 1916
rect 1597 1844 1603 1856
rect 1629 1784 1635 1856
rect 1645 1844 1651 1856
rect 1693 1824 1699 1836
rect 1565 1777 1587 1783
rect 1565 1764 1571 1777
rect 1597 1764 1603 1776
rect 1549 1737 1628 1743
rect 1549 1724 1555 1737
rect 1725 1743 1731 1876
rect 1773 1864 1779 1896
rect 1901 1884 1907 1917
rect 1940 1917 1948 1923
rect 2093 1923 2099 1937
rect 2084 1917 2099 1923
rect 1956 1877 1980 1883
rect 1860 1857 1891 1863
rect 1789 1843 1795 1856
rect 1789 1837 1875 1843
rect 1709 1737 1731 1743
rect 1581 1703 1587 1716
rect 1517 1697 1587 1703
rect 1373 1544 1379 1696
rect 1469 1623 1475 1696
rect 1453 1617 1475 1623
rect 1245 1504 1251 1516
rect 957 1484 963 1496
rect 1085 1464 1091 1476
rect 1021 1424 1027 1436
rect 1101 1423 1107 1476
rect 1101 1417 1123 1423
rect 1085 1364 1091 1416
rect 941 1344 947 1356
rect 1117 1344 1123 1417
rect 1133 1364 1139 1436
rect 1149 1424 1155 1496
rect 1261 1483 1267 1536
rect 1293 1524 1299 1536
rect 1405 1524 1411 1536
rect 1405 1504 1411 1516
rect 1453 1504 1459 1617
rect 1501 1543 1507 1676
rect 1645 1644 1651 1716
rect 1677 1644 1683 1716
rect 1709 1644 1715 1737
rect 1757 1743 1763 1836
rect 1869 1824 1875 1837
rect 1773 1764 1779 1816
rect 1885 1803 1891 1857
rect 1933 1844 1939 1856
rect 1965 1824 1971 1836
rect 1997 1824 2003 1876
rect 1853 1797 1891 1803
rect 1853 1784 1859 1797
rect 1789 1744 1795 1756
rect 1757 1737 1779 1743
rect 1725 1717 1740 1723
rect 1725 1684 1731 1717
rect 1533 1584 1539 1636
rect 1565 1597 1603 1603
rect 1565 1584 1571 1597
rect 1597 1584 1603 1597
rect 1492 1537 1507 1543
rect 1533 1504 1539 1516
rect 1581 1504 1587 1576
rect 1773 1544 1779 1737
rect 1821 1584 1827 1696
rect 1885 1684 1891 1756
rect 1917 1704 1923 1716
rect 1901 1564 1907 1636
rect 1933 1604 1939 1816
rect 2013 1764 2019 1816
rect 2077 1803 2083 1876
rect 2109 1864 2115 1896
rect 2157 1884 2163 2116
rect 2173 2064 2179 2156
rect 2253 2124 2259 2196
rect 2285 2183 2291 2197
rect 2413 2184 2419 2276
rect 2445 2264 2451 2276
rect 2461 2203 2467 2296
rect 2493 2284 2499 2336
rect 2493 2264 2499 2276
rect 2509 2264 2515 2376
rect 2573 2317 2588 2323
rect 2573 2304 2579 2317
rect 2605 2303 2611 2416
rect 2637 2324 2643 2476
rect 2669 2384 2675 2436
rect 2701 2363 2707 2556
rect 2717 2504 2723 2536
rect 2733 2484 2739 2516
rect 2765 2504 2771 2516
rect 2781 2504 2787 2556
rect 2845 2537 2860 2543
rect 2813 2444 2819 2516
rect 2845 2484 2851 2537
rect 2925 2524 2931 2736
rect 3117 2724 3123 2756
rect 2941 2684 2947 2696
rect 3069 2684 3075 2696
rect 3149 2684 3155 2896
rect 3165 2764 3171 2836
rect 3293 2784 3299 2936
rect 3325 2904 3331 2916
rect 3357 2764 3363 2836
rect 3389 2824 3395 2956
rect 3421 2904 3427 2916
rect 3412 2857 3420 2863
rect 3165 2684 3171 2736
rect 3197 2724 3203 2736
rect 3437 2724 3443 2936
rect 3469 2904 3475 2916
rect 3517 2804 3523 2956
rect 3549 2924 3555 2996
rect 3565 2984 3571 3017
rect 3581 3004 3587 3096
rect 3725 3084 3731 3196
rect 3773 3144 3779 3176
rect 3796 3157 3804 3163
rect 3933 3144 3939 3336
rect 4221 3324 4227 3356
rect 4180 3317 4188 3323
rect 4029 3304 4035 3316
rect 4045 3304 4051 3316
rect 4020 3137 4028 3143
rect 3741 3084 3747 3116
rect 4029 3104 4035 3116
rect 3940 3097 3948 3103
rect 3629 3064 3635 3076
rect 3693 3064 3699 3076
rect 3677 3044 3683 3056
rect 3597 3024 3603 3036
rect 3693 2964 3699 3036
rect 3597 2924 3603 2936
rect 3613 2904 3619 2956
rect 3661 2924 3667 2936
rect 3629 2904 3635 2916
rect 3556 2897 3564 2903
rect 3645 2784 3651 2836
rect 3485 2724 3491 2756
rect 3517 2724 3523 2776
rect 3661 2724 3667 2736
rect 3245 2664 3251 2676
rect 3060 2657 3075 2663
rect 2957 2564 2963 2576
rect 2973 2564 2979 2656
rect 3005 2644 3011 2656
rect 2989 2584 2995 2636
rect 3069 2623 3075 2657
rect 3101 2623 3107 2636
rect 3069 2617 3107 2623
rect 3181 2604 3187 2636
rect 3261 2624 3267 2716
rect 3485 2704 3491 2716
rect 3533 2704 3539 2716
rect 3364 2697 3443 2703
rect 3437 2683 3443 2697
rect 3437 2677 3468 2683
rect 3293 2664 3299 2676
rect 3389 2664 3395 2676
rect 3437 2624 3443 2656
rect 3565 2644 3571 2656
rect 3613 2644 3619 2696
rect 3636 2677 3651 2683
rect 3645 2663 3651 2677
rect 3645 2657 3683 2663
rect 3677 2644 3683 2657
rect 3693 2643 3699 2896
rect 3709 2704 3715 2916
rect 3748 2897 3756 2903
rect 3709 2684 3715 2696
rect 3716 2657 3731 2663
rect 3725 2644 3731 2657
rect 3693 2637 3715 2643
rect 3501 2624 3507 2636
rect 3261 2604 3267 2616
rect 3277 2597 3427 2603
rect 3245 2583 3251 2596
rect 3277 2583 3283 2597
rect 3005 2577 3219 2583
rect 3245 2577 3283 2583
rect 3325 2577 3411 2583
rect 3005 2564 3011 2577
rect 3076 2557 3139 2563
rect 2861 2484 2867 2516
rect 2877 2484 2883 2516
rect 2685 2357 2707 2363
rect 2653 2304 2659 2356
rect 2605 2297 2627 2303
rect 2525 2284 2531 2296
rect 2541 2277 2556 2283
rect 2445 2197 2467 2203
rect 2285 2177 2364 2183
rect 2445 2164 2451 2197
rect 2493 2184 2499 2196
rect 2509 2164 2515 2176
rect 2461 2157 2499 2163
rect 2285 2124 2291 2156
rect 2461 2144 2467 2157
rect 2493 2144 2499 2157
rect 2244 2097 2252 2103
rect 2093 1804 2099 1836
rect 2141 1824 2147 1856
rect 2157 1824 2163 1876
rect 2173 1863 2179 2016
rect 2189 1924 2195 1936
rect 2237 1864 2243 1896
rect 2173 1857 2220 1863
rect 2061 1797 2083 1803
rect 1949 1744 1955 1756
rect 1892 1537 1900 1543
rect 1604 1497 1612 1503
rect 1677 1503 1683 1536
rect 1805 1524 1811 1536
rect 1677 1497 1699 1503
rect 1373 1484 1379 1496
rect 1245 1477 1267 1483
rect 1181 1404 1187 1456
rect 1229 1424 1235 1476
rect 1245 1364 1251 1477
rect 1373 1464 1379 1476
rect 1549 1464 1555 1496
rect 1412 1457 1420 1463
rect 1485 1457 1500 1463
rect 1277 1424 1283 1456
rect 1309 1403 1315 1436
rect 1357 1424 1363 1456
rect 1405 1424 1411 1436
rect 1341 1403 1347 1416
rect 1309 1397 1331 1403
rect 1341 1397 1363 1403
rect 1028 1337 1036 1343
rect 1181 1324 1187 1336
rect 1213 1324 1219 1336
rect 973 1124 979 1216
rect 989 1184 995 1316
rect 1117 1304 1123 1316
rect 1069 1264 1075 1296
rect 1213 1284 1219 1296
rect 1053 1163 1059 1176
rect 1101 1164 1107 1236
rect 1037 1157 1059 1163
rect 973 1084 979 1096
rect 989 1084 995 1096
rect 1021 1044 1027 1056
rect 845 984 851 1036
rect 861 964 867 996
rect 893 964 899 1036
rect 829 957 844 963
rect 909 957 924 963
rect 813 943 819 956
rect 909 943 915 957
rect 957 944 963 1036
rect 1037 984 1043 1157
rect 1108 1137 1180 1143
rect 1101 1104 1107 1116
rect 1165 1104 1171 1116
rect 1197 1104 1203 1236
rect 1261 1164 1267 1296
rect 1245 1084 1251 1116
rect 1293 1084 1299 1276
rect 1325 1264 1331 1397
rect 1357 1384 1363 1397
rect 1341 1344 1347 1376
rect 1389 1364 1395 1416
rect 1405 1404 1411 1416
rect 1389 1304 1395 1356
rect 1309 1124 1315 1136
rect 1341 1084 1347 1216
rect 1357 1104 1363 1116
rect 1069 1064 1075 1076
rect 1197 1064 1203 1076
rect 1117 1057 1187 1063
rect 1053 1043 1059 1056
rect 1053 1037 1075 1043
rect 1005 964 1011 976
rect 980 957 1004 963
rect 813 937 915 943
rect 765 924 771 936
rect 797 904 803 916
rect 765 884 771 896
rect 813 883 819 916
rect 797 877 819 883
rect 653 717 755 723
rect 557 704 563 716
rect 653 704 659 717
rect 669 697 748 703
rect 628 677 643 683
rect 509 664 515 676
rect 525 664 531 676
rect 525 584 531 596
rect 541 564 547 596
rect 509 524 515 556
rect 557 544 563 676
rect 637 663 643 677
rect 669 683 675 697
rect 765 684 771 736
rect 660 677 675 683
rect 685 677 700 683
rect 685 663 691 677
rect 637 657 691 663
rect 605 564 611 636
rect 621 604 627 656
rect 621 584 627 596
rect 685 583 691 636
rect 701 624 707 656
rect 717 584 723 656
rect 781 584 787 636
rect 685 577 707 583
rect 701 564 707 577
rect 765 564 771 576
rect 685 544 691 556
rect 749 543 755 556
rect 749 537 780 543
rect 797 543 803 877
rect 845 724 851 816
rect 925 743 931 916
rect 957 904 963 916
rect 1021 844 1027 936
rect 1053 904 1059 996
rect 1069 964 1075 1037
rect 1117 1024 1123 1057
rect 1140 1037 1171 1043
rect 1133 984 1139 996
rect 1117 964 1123 976
rect 1149 944 1155 1016
rect 1165 963 1171 1037
rect 1181 1024 1187 1057
rect 1181 984 1187 996
rect 1165 957 1219 963
rect 1124 937 1139 943
rect 1069 904 1075 916
rect 1133 864 1139 937
rect 925 737 956 743
rect 893 704 899 716
rect 861 684 867 696
rect 813 644 819 676
rect 829 584 835 636
rect 813 564 819 576
rect 797 537 812 543
rect 557 524 563 536
rect 829 524 835 556
rect 861 544 867 676
rect 925 624 931 636
rect 941 623 947 656
rect 973 624 979 636
rect 941 617 963 623
rect 925 564 931 576
rect 957 564 963 617
rect 957 544 963 556
rect 884 537 899 543
rect 893 524 899 537
rect 973 524 979 596
rect 989 584 995 836
rect 1149 804 1155 936
rect 1213 923 1219 957
rect 1245 944 1251 1036
rect 1277 964 1283 1036
rect 1309 1004 1315 1036
rect 1357 984 1363 1056
rect 1405 984 1411 1376
rect 1421 1284 1427 1356
rect 1469 1343 1475 1436
rect 1485 1384 1491 1457
rect 1549 1404 1555 1456
rect 1501 1384 1507 1396
rect 1453 1337 1475 1343
rect 1437 1204 1443 1316
rect 1453 1164 1459 1337
rect 1517 1224 1523 1336
rect 1533 1304 1539 1356
rect 1501 1184 1507 1216
rect 1421 1144 1427 1156
rect 1565 1144 1571 1476
rect 1581 1384 1587 1496
rect 1693 1484 1699 1497
rect 1629 1404 1635 1456
rect 1597 1384 1603 1396
rect 1645 1384 1651 1396
rect 1661 1383 1667 1476
rect 1677 1404 1683 1476
rect 1757 1404 1763 1456
rect 1661 1377 1676 1383
rect 1581 1344 1587 1376
rect 1629 1364 1635 1376
rect 1581 1264 1587 1316
rect 1581 1244 1587 1256
rect 1437 1084 1443 1136
rect 1485 1104 1491 1116
rect 1501 1097 1516 1103
rect 1501 1083 1507 1097
rect 1492 1077 1507 1083
rect 1533 1063 1539 1136
rect 1613 1124 1619 1276
rect 1661 1164 1667 1336
rect 1693 1323 1699 1396
rect 1709 1364 1715 1376
rect 1741 1343 1747 1356
rect 1725 1337 1747 1343
rect 1725 1324 1731 1337
rect 1693 1317 1715 1323
rect 1645 1124 1651 1136
rect 1572 1117 1580 1123
rect 1613 1084 1619 1096
rect 1524 1057 1539 1063
rect 1453 1044 1459 1056
rect 1581 1024 1587 1056
rect 1453 984 1459 996
rect 1213 917 1228 923
rect 1165 784 1171 836
rect 1181 784 1187 896
rect 1229 884 1235 896
rect 1037 744 1043 776
rect 1005 724 1011 736
rect 1037 717 1107 723
rect 1005 704 1011 716
rect 1037 703 1043 717
rect 1101 704 1107 717
rect 1149 704 1155 756
rect 1021 697 1043 703
rect 1021 683 1027 697
rect 1053 684 1059 696
rect 1012 677 1027 683
rect 1037 644 1043 676
rect 1005 624 1011 636
rect 1085 584 1091 696
rect 1101 624 1107 656
rect 1133 623 1139 656
rect 1117 617 1139 623
rect 1117 604 1123 617
rect 1021 564 1027 576
rect 1133 564 1139 596
rect 196 517 204 523
rect 788 517 796 523
rect 205 423 211 436
rect 189 417 211 423
rect 141 304 147 316
rect 189 284 195 417
rect 285 304 291 316
rect 228 297 236 303
rect 317 284 323 356
rect 628 337 636 343
rect 381 304 387 316
rect 429 284 435 316
rect 420 257 444 263
rect 77 224 83 256
rect 93 124 99 256
rect 125 244 131 256
rect 125 164 131 176
rect 141 164 147 236
rect 253 123 259 236
rect 317 144 323 256
rect 477 244 483 256
rect 509 244 515 296
rect 397 224 403 236
rect 356 177 364 183
rect 333 164 339 176
rect 413 144 419 236
rect 557 224 563 256
rect 573 204 579 236
rect 445 164 451 176
rect 573 164 579 176
rect 468 157 476 163
rect 589 144 595 276
rect 605 224 611 296
rect 653 284 659 476
rect 749 464 755 516
rect 909 504 915 516
rect 989 503 995 516
rect 980 497 995 503
rect 948 477 956 483
rect 893 464 899 476
rect 1005 464 1011 536
rect 1021 504 1027 556
rect 1149 544 1155 616
rect 1181 604 1187 696
rect 1277 684 1283 936
rect 1373 924 1379 936
rect 1325 764 1331 916
rect 1341 904 1347 916
rect 1373 864 1379 916
rect 1229 644 1235 676
rect 1245 624 1251 636
rect 1229 543 1235 596
rect 1277 544 1283 676
rect 1325 643 1331 696
rect 1341 664 1347 836
rect 1421 824 1427 956
rect 1469 904 1475 916
rect 1533 904 1539 916
rect 1364 777 1372 783
rect 1389 664 1395 736
rect 1437 704 1443 776
rect 1485 724 1491 896
rect 1565 884 1571 896
rect 1517 683 1523 716
rect 1501 677 1523 683
rect 1501 663 1507 677
rect 1549 664 1555 836
rect 1597 764 1603 1036
rect 1629 983 1635 1036
rect 1645 984 1651 996
rect 1661 984 1667 1096
rect 1693 1063 1699 1116
rect 1709 1084 1715 1317
rect 1748 1317 1756 1323
rect 1773 1323 1779 1496
rect 1853 1484 1859 1496
rect 1789 1363 1795 1436
rect 1821 1404 1827 1436
rect 1837 1364 1843 1396
rect 1853 1364 1859 1476
rect 1901 1443 1907 1476
rect 1917 1464 1923 1476
rect 1901 1437 1923 1443
rect 1917 1364 1923 1437
rect 1789 1357 1820 1363
rect 1876 1357 1884 1363
rect 1796 1337 1811 1343
rect 1773 1317 1795 1323
rect 1741 1184 1747 1256
rect 1757 1184 1763 1296
rect 1741 1164 1747 1176
rect 1725 1124 1731 1156
rect 1741 1144 1747 1156
rect 1725 1064 1731 1116
rect 1789 1103 1795 1317
rect 1805 1304 1811 1337
rect 1901 1343 1907 1356
rect 1933 1344 1939 1396
rect 1892 1337 1907 1343
rect 1844 1317 1852 1323
rect 1876 1317 1884 1323
rect 1924 1297 1932 1303
rect 1949 1264 1955 1596
rect 1981 1563 1987 1756
rect 1997 1724 2003 1736
rect 2013 1724 2019 1736
rect 1997 1584 2003 1636
rect 2045 1604 2051 1676
rect 2061 1583 2067 1797
rect 2125 1784 2131 1796
rect 2253 1764 2259 1836
rect 2116 1757 2131 1763
rect 2125 1744 2131 1757
rect 2093 1724 2099 1736
rect 2109 1724 2115 1736
rect 2157 1664 2163 1756
rect 2189 1744 2195 1756
rect 2237 1743 2243 1756
rect 2237 1737 2252 1743
rect 2221 1724 2227 1736
rect 2052 1577 2067 1583
rect 1981 1557 2003 1563
rect 1997 1544 2003 1557
rect 2125 1504 2131 1616
rect 2141 1504 2147 1616
rect 2205 1584 2211 1636
rect 2164 1497 2172 1503
rect 2045 1484 2051 1496
rect 2189 1484 2195 1516
rect 2013 1464 2019 1476
rect 2221 1464 2227 1596
rect 2269 1544 2275 2096
rect 2333 2084 2339 2136
rect 2301 2024 2307 2076
rect 2349 2023 2355 2136
rect 2477 2124 2483 2136
rect 2381 2104 2387 2116
rect 2509 2104 2515 2156
rect 2541 2143 2547 2277
rect 2573 2263 2579 2276
rect 2589 2264 2595 2296
rect 2564 2257 2579 2263
rect 2621 2263 2627 2297
rect 2605 2257 2627 2263
rect 2573 2223 2579 2236
rect 2573 2217 2588 2223
rect 2557 2164 2563 2196
rect 2605 2164 2611 2257
rect 2621 2184 2627 2216
rect 2685 2183 2691 2357
rect 2701 2224 2707 2336
rect 2637 2177 2691 2183
rect 2573 2143 2579 2156
rect 2541 2137 2579 2143
rect 2637 2143 2643 2177
rect 2701 2164 2707 2176
rect 2717 2164 2723 2396
rect 2749 2384 2755 2416
rect 2749 2323 2755 2336
rect 2781 2323 2787 2336
rect 2797 2324 2803 2396
rect 2749 2317 2787 2323
rect 2836 2297 2844 2303
rect 2797 2284 2803 2296
rect 2861 2284 2867 2336
rect 2877 2284 2883 2296
rect 2740 2277 2755 2283
rect 2749 2263 2755 2277
rect 2813 2263 2819 2276
rect 2749 2257 2819 2263
rect 2733 2224 2739 2256
rect 2797 2183 2803 2216
rect 2845 2204 2851 2256
rect 2893 2204 2899 2216
rect 2909 2204 2915 2276
rect 2829 2184 2835 2196
rect 2893 2184 2899 2196
rect 2749 2177 2803 2183
rect 2660 2157 2675 2163
rect 2637 2137 2652 2143
rect 2669 2143 2675 2157
rect 2749 2163 2755 2177
rect 2733 2157 2755 2163
rect 2733 2143 2739 2157
rect 2820 2157 2915 2163
rect 2909 2144 2915 2157
rect 2669 2137 2739 2143
rect 2797 2137 2835 2143
rect 2397 2044 2403 2076
rect 2493 2063 2499 2096
rect 2493 2057 2547 2063
rect 2541 2043 2547 2057
rect 2541 2037 2579 2043
rect 2349 2017 2371 2023
rect 2285 1924 2291 1996
rect 2317 1884 2323 1936
rect 2317 1864 2323 1876
rect 2333 1844 2339 1896
rect 2365 1864 2371 2017
rect 2413 1944 2419 2036
rect 2445 1924 2451 1956
rect 2461 1904 2467 2036
rect 2525 2024 2531 2036
rect 2557 1964 2563 2016
rect 2573 1983 2579 2037
rect 2605 2024 2611 2116
rect 2628 2077 2636 2083
rect 2653 2037 2691 2043
rect 2653 2024 2659 2037
rect 2685 2024 2691 2037
rect 2717 2024 2723 2076
rect 2749 2064 2755 2136
rect 2797 2103 2803 2137
rect 2829 2124 2835 2137
rect 2861 2124 2867 2136
rect 2788 2097 2803 2103
rect 2733 2043 2739 2056
rect 2733 2037 2764 2043
rect 2621 1984 2627 2016
rect 2573 1977 2611 1983
rect 2605 1964 2611 1977
rect 2580 1957 2588 1963
rect 2637 1904 2643 1916
rect 2525 1883 2531 1896
rect 2461 1877 2531 1883
rect 2397 1843 2403 1856
rect 2356 1837 2403 1843
rect 2285 1664 2291 1696
rect 2301 1624 2307 1696
rect 1981 1363 1987 1436
rect 2125 1424 2131 1456
rect 1997 1384 2003 1396
rect 1965 1357 1987 1363
rect 1965 1304 1971 1357
rect 1965 1243 1971 1256
rect 1949 1237 1971 1243
rect 1805 1144 1811 1236
rect 1949 1183 1955 1237
rect 1908 1177 1955 1183
rect 1965 1163 1971 1216
rect 1949 1157 1971 1163
rect 1917 1124 1923 1136
rect 1773 1097 1795 1103
rect 1693 1057 1708 1063
rect 1613 977 1635 983
rect 1613 924 1619 977
rect 1684 977 1692 983
rect 1709 963 1715 996
rect 1773 984 1779 1097
rect 1812 1097 1859 1103
rect 1853 1083 1859 1097
rect 1949 1084 1955 1157
rect 1965 1124 1971 1136
rect 1981 1103 1987 1336
rect 2013 1304 2019 1416
rect 2077 1377 2147 1383
rect 2077 1364 2083 1377
rect 2100 1357 2108 1363
rect 2036 1337 2060 1343
rect 2077 1304 2083 1316
rect 2061 1264 2067 1276
rect 2077 1224 2083 1256
rect 2013 1124 2019 1216
rect 2125 1144 2131 1356
rect 2141 1303 2147 1377
rect 2157 1324 2163 1396
rect 2205 1364 2211 1396
rect 2221 1384 2227 1416
rect 2253 1404 2259 1516
rect 2269 1464 2275 1496
rect 2285 1484 2291 1616
rect 2317 1584 2323 1716
rect 2333 1584 2339 1636
rect 2349 1604 2355 1716
rect 2365 1704 2371 1756
rect 2397 1744 2403 1776
rect 2404 1697 2412 1703
rect 2381 1484 2387 1696
rect 2429 1584 2435 1836
rect 2461 1823 2467 1877
rect 2589 1877 2643 1883
rect 2589 1863 2595 1877
rect 2637 1864 2643 1877
rect 2548 1857 2595 1863
rect 2452 1817 2467 1823
rect 2477 1784 2483 1816
rect 2493 1803 2499 1856
rect 2605 1843 2611 1856
rect 2541 1837 2611 1843
rect 2525 1803 2531 1836
rect 2541 1824 2547 1837
rect 2557 1804 2563 1816
rect 2493 1797 2531 1803
rect 2445 1744 2451 1776
rect 2461 1564 2467 1756
rect 2493 1704 2499 1716
rect 2477 1584 2483 1696
rect 2509 1564 2515 1756
rect 2525 1564 2531 1716
rect 2557 1704 2563 1796
rect 2605 1744 2611 1796
rect 2580 1697 2588 1703
rect 2436 1557 2451 1563
rect 2445 1524 2451 1557
rect 2477 1543 2483 1556
rect 2541 1543 2547 1696
rect 2605 1603 2611 1736
rect 2637 1704 2643 1796
rect 2557 1597 2595 1603
rect 2605 1597 2627 1603
rect 2557 1584 2563 1597
rect 2589 1583 2595 1597
rect 2589 1577 2604 1583
rect 2557 1544 2563 1556
rect 2461 1537 2483 1543
rect 2525 1537 2547 1543
rect 2429 1504 2435 1516
rect 2461 1503 2467 1537
rect 2445 1497 2467 1503
rect 2173 1324 2179 1356
rect 2253 1344 2259 1356
rect 2269 1343 2275 1436
rect 2365 1423 2371 1476
rect 2349 1417 2371 1423
rect 2381 1423 2387 1456
rect 2397 1444 2403 1456
rect 2381 1417 2403 1423
rect 2333 1384 2339 1416
rect 2308 1357 2339 1363
rect 2333 1344 2339 1357
rect 2269 1337 2291 1343
rect 2205 1317 2259 1323
rect 2205 1303 2211 1317
rect 2141 1297 2211 1303
rect 2253 1284 2259 1317
rect 2221 1224 2227 1256
rect 2285 1224 2291 1337
rect 1965 1097 1987 1103
rect 1853 1077 1891 1083
rect 1789 984 1795 1076
rect 1837 1004 1843 1076
rect 1885 1064 1891 1077
rect 1853 1023 1859 1056
rect 1917 1024 1923 1036
rect 1853 1017 1907 1023
rect 1901 1003 1907 1017
rect 1901 997 1923 1003
rect 1869 964 1875 976
rect 1668 957 1715 963
rect 1892 957 1900 963
rect 1741 944 1747 956
rect 1837 944 1843 956
rect 1917 943 1923 997
rect 1933 964 1939 1016
rect 1965 1003 1971 1097
rect 2077 1084 2083 1096
rect 1997 1024 2003 1076
rect 2077 1044 2083 1056
rect 2029 1024 2035 1036
rect 1949 997 1971 1003
rect 1949 984 1955 997
rect 2093 984 2099 1116
rect 2141 1064 2147 1216
rect 2173 1184 2179 1216
rect 2237 1104 2243 1116
rect 2285 1104 2291 1116
rect 2189 1083 2195 1096
rect 2173 1077 2195 1083
rect 2109 983 2115 1036
rect 2125 1024 2131 1036
rect 2173 1023 2179 1077
rect 2189 1024 2195 1056
rect 2221 1037 2236 1043
rect 2205 1024 2211 1036
rect 2157 1017 2179 1023
rect 2157 984 2163 1017
rect 2221 1003 2227 1037
rect 2205 997 2227 1003
rect 2109 977 2147 983
rect 2141 963 2147 977
rect 2141 957 2188 963
rect 1981 944 1987 956
rect 1901 937 1923 943
rect 1709 904 1715 916
rect 1645 744 1651 856
rect 1709 844 1715 896
rect 1725 844 1731 856
rect 1709 784 1715 816
rect 1741 804 1747 936
rect 1885 884 1891 896
rect 1757 864 1763 876
rect 1773 784 1779 796
rect 1597 724 1603 736
rect 1645 724 1651 736
rect 1572 717 1580 723
rect 1581 684 1587 696
rect 1661 684 1667 776
rect 1693 724 1699 776
rect 1789 744 1795 876
rect 1805 684 1811 836
rect 1901 784 1907 937
rect 2077 943 2083 956
rect 2077 937 2092 943
rect 1933 884 1939 936
rect 1981 923 1987 936
rect 2173 924 2179 936
rect 1981 917 2003 923
rect 1997 884 2003 917
rect 1940 857 1948 863
rect 1853 724 1859 736
rect 1917 724 1923 796
rect 1949 704 1955 836
rect 2029 784 2035 896
rect 2045 824 2051 836
rect 1741 677 1779 683
rect 1412 657 1507 663
rect 1325 637 1420 643
rect 1309 624 1315 636
rect 1229 537 1251 543
rect 733 324 739 336
rect 637 144 643 256
rect 653 204 659 256
rect 685 223 691 296
rect 781 284 787 356
rect 845 324 851 336
rect 909 324 915 356
rect 989 324 995 336
rect 765 264 771 276
rect 701 224 707 236
rect 669 217 691 223
rect 669 184 675 217
rect 692 177 700 183
rect 717 144 723 216
rect 733 164 739 176
rect 781 144 787 156
rect 861 144 867 296
rect 941 284 947 316
rect 893 244 899 256
rect 925 204 931 236
rect 957 224 963 256
rect 989 244 995 296
rect 1005 284 1011 456
rect 1069 404 1075 516
rect 1117 424 1123 436
rect 1101 284 1107 316
rect 1117 303 1123 356
rect 1133 324 1139 356
rect 1181 323 1187 476
rect 1181 317 1196 323
rect 1149 304 1155 316
rect 1117 297 1139 303
rect 1133 284 1139 297
rect 1213 283 1219 356
rect 1229 284 1235 456
rect 1245 323 1251 537
rect 1293 524 1299 596
rect 1341 564 1347 616
rect 1533 604 1539 656
rect 1581 623 1587 676
rect 1629 644 1635 676
rect 1677 624 1683 676
rect 1725 624 1731 676
rect 1741 664 1747 677
rect 1773 663 1779 677
rect 1773 657 1804 663
rect 1853 657 1868 663
rect 1757 624 1763 656
rect 1581 617 1603 623
rect 1469 584 1475 596
rect 1597 564 1603 617
rect 1693 577 1724 583
rect 1540 557 1564 563
rect 1373 544 1379 556
rect 1437 544 1443 556
rect 1540 537 1548 543
rect 1325 524 1331 536
rect 1444 517 1452 523
rect 1421 504 1427 516
rect 1581 504 1587 536
rect 1293 324 1299 336
rect 1245 317 1276 323
rect 1341 304 1347 316
rect 1325 284 1331 296
rect 1341 284 1347 296
rect 1357 284 1363 296
rect 1181 277 1219 283
rect 1181 264 1187 277
rect 1092 257 1116 263
rect 1197 204 1203 236
rect 1245 224 1251 276
rect 1373 264 1379 436
rect 1389 344 1395 476
rect 1437 403 1443 496
rect 1597 483 1603 556
rect 1677 544 1683 556
rect 1693 544 1699 577
rect 1636 537 1644 543
rect 1421 397 1443 403
rect 1581 477 1603 483
rect 1405 384 1411 396
rect 1421 284 1427 397
rect 1549 324 1555 376
rect 1581 303 1587 477
rect 1645 464 1651 516
rect 1677 464 1683 496
rect 1645 364 1651 396
rect 1661 384 1667 436
rect 1684 337 1692 343
rect 1597 324 1603 336
rect 1469 297 1523 303
rect 1581 297 1603 303
rect 1437 284 1443 296
rect 1469 284 1475 297
rect 1517 284 1523 297
rect 1485 264 1491 276
rect 1277 224 1283 236
rect 957 164 963 196
rect 989 164 995 196
rect 1133 184 1139 196
rect 1165 164 1171 176
rect 1245 163 1251 176
rect 1245 157 1276 163
rect 989 144 995 156
rect 1213 144 1219 156
rect 1229 144 1235 156
rect 916 137 924 143
rect 1028 137 1084 143
rect 493 124 499 136
rect 765 124 771 136
rect 877 124 883 136
rect 1309 124 1315 236
rect 1469 184 1475 256
rect 1357 164 1363 176
rect 253 117 268 123
rect 653 117 691 123
rect 285 104 291 116
rect 532 97 540 103
rect 628 97 636 103
rect 653 84 659 117
rect 685 104 691 117
rect 1085 104 1091 116
rect 1181 104 1187 116
rect 1421 104 1427 156
rect 1501 144 1507 236
rect 1517 104 1523 176
rect 916 97 940 103
rect 1581 103 1587 236
rect 1597 144 1603 297
rect 1613 284 1619 336
rect 1645 324 1651 336
rect 1661 283 1667 336
rect 1709 304 1715 536
rect 1725 504 1731 556
rect 1757 544 1763 556
rect 1773 524 1779 636
rect 1837 624 1843 636
rect 1853 584 1859 657
rect 1917 564 1923 616
rect 1965 564 1971 676
rect 1997 664 2003 776
rect 2061 724 2067 776
rect 2013 704 2019 716
rect 2093 684 2099 856
rect 2109 743 2115 816
rect 2125 784 2131 796
rect 2141 784 2147 896
rect 2157 764 2163 816
rect 2173 744 2179 916
rect 2189 784 2195 796
rect 2205 744 2211 997
rect 2237 964 2243 976
rect 2269 964 2275 1096
rect 2301 1064 2307 1336
rect 2317 1224 2323 1336
rect 2349 1304 2355 1417
rect 2381 1344 2387 1376
rect 2397 1344 2403 1417
rect 2413 1404 2419 1496
rect 2445 1404 2451 1497
rect 2484 1497 2508 1503
rect 2477 1463 2483 1476
rect 2525 1464 2531 1537
rect 2564 1537 2595 1543
rect 2557 1523 2563 1536
rect 2548 1517 2563 1523
rect 2573 1464 2579 1516
rect 2589 1504 2595 1537
rect 2621 1524 2627 1597
rect 2621 1504 2627 1516
rect 2653 1504 2659 1956
rect 2669 1884 2675 2016
rect 2708 1977 2787 1983
rect 2756 1957 2764 1963
rect 2685 1924 2691 1956
rect 2717 1884 2723 1896
rect 2685 1823 2691 1876
rect 2765 1824 2771 1856
rect 2685 1817 2723 1823
rect 2717 1804 2723 1817
rect 2733 1784 2739 1816
rect 2781 1804 2787 1977
rect 2797 1923 2803 2056
rect 2813 1964 2819 2116
rect 2877 2064 2883 2136
rect 2925 2123 2931 2496
rect 2941 2444 2947 2496
rect 2957 2484 2963 2556
rect 2973 2444 2979 2496
rect 2941 2304 2947 2316
rect 2909 2117 2931 2123
rect 2909 2104 2915 2117
rect 2829 1943 2835 2056
rect 2925 2024 2931 2076
rect 2941 2064 2947 2276
rect 2957 2264 2963 2316
rect 2989 2304 2995 2336
rect 2957 2064 2963 2256
rect 2973 2164 2979 2216
rect 2973 2124 2979 2136
rect 2973 2084 2979 2116
rect 2941 1984 2947 2056
rect 2989 1963 2995 2276
rect 3005 2264 3011 2476
rect 3021 2404 3027 2536
rect 3133 2523 3139 2557
rect 3213 2563 3219 2577
rect 3213 2557 3228 2563
rect 3325 2563 3331 2577
rect 3405 2564 3411 2577
rect 3300 2557 3331 2563
rect 3149 2544 3155 2556
rect 3165 2537 3251 2543
rect 3165 2523 3171 2537
rect 3133 2517 3171 2523
rect 3053 2504 3059 2516
rect 3085 2484 3091 2496
rect 3101 2484 3107 2516
rect 3197 2504 3203 2516
rect 3245 2504 3251 2537
rect 3325 2504 3331 2536
rect 3133 2497 3148 2503
rect 3117 2344 3123 2496
rect 3133 2484 3139 2497
rect 3220 2497 3228 2503
rect 3293 2444 3299 2496
rect 3373 2444 3379 2556
rect 3405 2504 3411 2516
rect 3421 2504 3427 2597
rect 3517 2597 3571 2603
rect 3517 2563 3523 2597
rect 3492 2557 3523 2563
rect 3533 2577 3548 2583
rect 3533 2544 3539 2577
rect 3453 2524 3459 2536
rect 3549 2524 3555 2556
rect 3565 2524 3571 2597
rect 3597 2524 3603 2616
rect 3645 2564 3651 2576
rect 3629 2524 3635 2556
rect 3693 2544 3699 2596
rect 3709 2584 3715 2637
rect 3501 2504 3507 2516
rect 3581 2504 3587 2516
rect 3140 2437 3148 2443
rect 3332 2437 3340 2443
rect 3197 2384 3203 2436
rect 3245 2384 3251 2416
rect 3037 2304 3043 2316
rect 3085 2284 3091 2296
rect 3133 2284 3139 2296
rect 3037 2264 3043 2276
rect 3165 2264 3171 2356
rect 3005 2224 3011 2256
rect 3117 2244 3123 2256
rect 3069 2184 3075 2216
rect 3213 2184 3219 2256
rect 3261 2244 3267 2256
rect 3277 2164 3283 2416
rect 3293 2384 3299 2396
rect 3357 2304 3363 2316
rect 3325 2284 3331 2296
rect 3373 2284 3379 2336
rect 3309 2224 3315 2276
rect 3405 2264 3411 2316
rect 3421 2304 3427 2476
rect 3396 2237 3404 2243
rect 3325 2184 3331 2236
rect 3357 2224 3363 2236
rect 3421 2223 3427 2256
rect 3405 2217 3427 2223
rect 3108 2137 3123 2143
rect 3021 2124 3027 2136
rect 3117 2124 3123 2137
rect 3069 2104 3075 2116
rect 3037 2024 3043 2036
rect 3053 2024 3059 2096
rect 3101 2084 3107 2116
rect 2973 1957 2995 1963
rect 2820 1937 2835 1943
rect 2797 1917 2819 1923
rect 2797 1864 2803 1896
rect 2813 1803 2819 1917
rect 2797 1797 2819 1803
rect 2797 1764 2803 1797
rect 2845 1803 2851 1916
rect 2861 1884 2867 1896
rect 2893 1824 2899 1916
rect 2909 1884 2915 1896
rect 2957 1824 2963 1876
rect 2868 1817 2883 1823
rect 2877 1803 2883 1817
rect 2909 1803 2915 1816
rect 2973 1804 2979 1957
rect 3005 1944 3011 1956
rect 3005 1884 3011 1916
rect 3037 1883 3043 1916
rect 3101 1884 3107 2076
rect 3133 2024 3139 2156
rect 3229 2144 3235 2156
rect 3245 2144 3251 2156
rect 3293 2144 3299 2176
rect 3341 2164 3347 2176
rect 3389 2163 3395 2216
rect 3405 2184 3411 2217
rect 3421 2164 3427 2196
rect 3437 2184 3443 2376
rect 3517 2303 3523 2336
rect 3508 2297 3523 2303
rect 3453 2164 3459 2296
rect 3469 2244 3475 2256
rect 3485 2184 3491 2236
rect 3389 2157 3404 2163
rect 3517 2144 3523 2156
rect 3188 2137 3196 2143
rect 3437 2137 3491 2143
rect 3293 2124 3299 2136
rect 3437 2124 3443 2137
rect 3485 2124 3491 2137
rect 3460 2117 3468 2123
rect 3149 2104 3155 2116
rect 3277 2104 3283 2116
rect 3133 1944 3139 1956
rect 3037 1877 3059 1883
rect 2989 1824 2995 1836
rect 3021 1824 3027 1836
rect 2845 1797 2867 1803
rect 2877 1797 2915 1803
rect 2829 1764 2835 1796
rect 2861 1783 2867 1797
rect 2925 1784 2931 1796
rect 2861 1777 2883 1783
rect 2756 1737 2780 1743
rect 2701 1724 2707 1736
rect 2788 1717 2796 1723
rect 2749 1704 2755 1716
rect 2708 1677 2780 1683
rect 2845 1604 2851 1636
rect 2861 1604 2867 1756
rect 2877 1743 2883 1777
rect 2957 1783 2963 1796
rect 2989 1783 2995 1796
rect 2957 1777 2995 1783
rect 2941 1764 2947 1776
rect 2957 1757 3011 1763
rect 2877 1737 2899 1743
rect 2877 1704 2883 1716
rect 2893 1704 2899 1737
rect 2909 1724 2915 1756
rect 2957 1743 2963 1757
rect 2925 1737 2963 1743
rect 2973 1737 2988 1743
rect 2925 1703 2931 1737
rect 2957 1704 2963 1716
rect 2909 1697 2931 1703
rect 2909 1683 2915 1697
rect 2900 1677 2915 1683
rect 2973 1663 2979 1737
rect 3005 1743 3011 1757
rect 3037 1744 3043 1816
rect 3053 1783 3059 1877
rect 3149 1864 3155 1976
rect 3245 1964 3251 2096
rect 3204 1957 3212 1963
rect 3204 1897 3228 1903
rect 3245 1884 3251 1956
rect 3277 1924 3283 2016
rect 3309 1984 3315 2016
rect 3325 1984 3331 2096
rect 3085 1784 3091 1856
rect 3053 1777 3075 1783
rect 3069 1763 3075 1777
rect 3101 1763 3107 1776
rect 3069 1757 3107 1763
rect 3005 1737 3027 1743
rect 3021 1724 3027 1737
rect 3108 1737 3123 1743
rect 3005 1704 3011 1716
rect 2989 1683 2995 1696
rect 2989 1677 3043 1683
rect 3037 1664 3043 1677
rect 2973 1657 2995 1663
rect 2925 1624 2931 1636
rect 2973 1624 2979 1636
rect 2989 1624 2995 1657
rect 3069 1624 3075 1636
rect 3085 1604 3091 1736
rect 2669 1597 2723 1603
rect 2669 1584 2675 1597
rect 2701 1524 2707 1576
rect 2653 1464 2659 1496
rect 2477 1457 2508 1463
rect 2669 1463 2675 1496
rect 2669 1457 2700 1463
rect 2461 1384 2467 1456
rect 2525 1444 2531 1456
rect 2397 1324 2403 1336
rect 2349 1244 2355 1296
rect 2317 1084 2323 1216
rect 2349 1104 2355 1116
rect 2365 1064 2371 1316
rect 2477 1304 2483 1436
rect 2589 1424 2595 1436
rect 2621 1424 2627 1456
rect 2717 1443 2723 1597
rect 2749 1584 2755 1596
rect 2996 1577 3004 1583
rect 2733 1484 2739 1496
rect 2701 1437 2723 1443
rect 2637 1423 2643 1436
rect 2637 1417 2659 1423
rect 2516 1397 2531 1403
rect 2525 1344 2531 1397
rect 2541 1364 2547 1416
rect 2653 1403 2659 1417
rect 2589 1397 2643 1403
rect 2653 1397 2675 1403
rect 2589 1384 2595 1397
rect 2493 1324 2499 1336
rect 2516 1317 2531 1323
rect 2525 1304 2531 1317
rect 2413 1224 2419 1276
rect 2461 1224 2467 1296
rect 2493 1257 2531 1263
rect 2493 1243 2499 1257
rect 2525 1244 2531 1257
rect 2484 1237 2499 1243
rect 2493 1124 2499 1216
rect 2509 1164 2515 1236
rect 2557 1184 2563 1356
rect 2589 1324 2595 1336
rect 2605 1324 2611 1376
rect 2637 1364 2643 1397
rect 2653 1364 2659 1376
rect 2669 1364 2675 1397
rect 2685 1364 2691 1436
rect 2701 1424 2707 1437
rect 2749 1424 2755 1496
rect 2717 1384 2723 1416
rect 2765 1363 2771 1576
rect 2893 1537 2963 1543
rect 2893 1523 2899 1537
rect 2861 1517 2899 1523
rect 2829 1464 2835 1496
rect 2813 1403 2819 1416
rect 2781 1397 2819 1403
rect 2781 1364 2787 1397
rect 2845 1383 2851 1516
rect 2861 1504 2867 1517
rect 2957 1523 2963 1537
rect 3021 1523 3027 1536
rect 3101 1524 3107 1536
rect 2916 1517 2947 1523
rect 2957 1517 3027 1523
rect 2941 1504 2947 1517
rect 2877 1484 2883 1496
rect 2861 1424 2867 1436
rect 2893 1424 2899 1456
rect 2925 1384 2931 1496
rect 2957 1444 2963 1456
rect 2973 1384 2979 1456
rect 3005 1404 3011 1496
rect 2845 1377 2867 1383
rect 2756 1357 2771 1363
rect 2813 1344 2819 1356
rect 2845 1344 2851 1356
rect 2685 1323 2691 1336
rect 2660 1317 2691 1323
rect 2820 1317 2844 1323
rect 2589 1184 2595 1316
rect 2637 1144 2643 1216
rect 2653 1184 2659 1296
rect 2701 1204 2707 1316
rect 2749 1224 2755 1316
rect 2845 1284 2851 1296
rect 2861 1264 2867 1377
rect 3005 1364 3011 1396
rect 3085 1384 3091 1456
rect 3101 1424 3107 1436
rect 2941 1344 2947 1356
rect 3021 1343 3027 1376
rect 2996 1337 3027 1343
rect 2893 1324 2899 1336
rect 2957 1244 2963 1336
rect 3053 1324 3059 1336
rect 3069 1323 3075 1376
rect 3085 1344 3091 1356
rect 3101 1323 3107 1356
rect 3069 1317 3107 1323
rect 3037 1304 3043 1316
rect 2669 1163 2675 1176
rect 2653 1157 2675 1163
rect 2461 1103 2467 1116
rect 2557 1103 2563 1136
rect 2461 1097 2563 1103
rect 2573 1084 2579 1116
rect 2621 1084 2627 1096
rect 2596 1077 2620 1083
rect 2340 1057 2348 1063
rect 2461 1057 2563 1063
rect 2333 1037 2371 1043
rect 2333 1024 2339 1037
rect 2365 1023 2371 1037
rect 2365 1017 2380 1023
rect 2349 984 2355 1016
rect 2388 957 2396 963
rect 2221 904 2227 936
rect 2237 804 2243 956
rect 2365 944 2371 956
rect 2429 944 2435 1036
rect 2461 1004 2467 1057
rect 2525 1037 2540 1043
rect 2477 984 2483 996
rect 2509 984 2515 1036
rect 2525 1024 2531 1037
rect 2557 1043 2563 1057
rect 2557 1037 2588 1043
rect 2461 964 2467 976
rect 2541 964 2547 1016
rect 2445 944 2451 956
rect 2525 944 2531 956
rect 2308 917 2316 923
rect 2269 904 2275 916
rect 2285 904 2291 916
rect 2253 764 2259 896
rect 2109 737 2140 743
rect 2157 697 2204 703
rect 2045 644 2051 656
rect 2109 644 2115 656
rect 2157 644 2163 697
rect 2221 683 2227 756
rect 2253 684 2259 756
rect 2269 744 2275 816
rect 2333 784 2339 896
rect 2381 884 2387 896
rect 2413 804 2419 936
rect 2493 924 2499 936
rect 2436 917 2444 923
rect 2589 903 2595 956
rect 2605 923 2611 1036
rect 2653 964 2659 1157
rect 2669 1104 2675 1116
rect 2685 1104 2691 1116
rect 2708 1097 2723 1103
rect 2717 1084 2723 1097
rect 2717 1044 2723 1056
rect 2765 1003 2771 1056
rect 2781 1024 2787 1076
rect 2797 1004 2803 1036
rect 2813 1024 2819 1116
rect 2829 1084 2835 1236
rect 3021 1184 3027 1216
rect 2925 1124 2931 1136
rect 3005 1124 3011 1156
rect 2877 1104 2883 1116
rect 3037 1084 3043 1176
rect 2829 1064 2835 1076
rect 2765 997 2787 1003
rect 2653 924 2659 936
rect 2669 924 2675 936
rect 2765 924 2771 936
rect 2605 917 2627 923
rect 2589 897 2604 903
rect 2397 744 2403 796
rect 2365 724 2371 736
rect 2541 724 2547 876
rect 2621 803 2627 917
rect 2765 904 2771 916
rect 2781 904 2787 997
rect 2877 984 2883 1016
rect 2861 964 2867 976
rect 2893 964 2899 996
rect 2909 984 2915 1076
rect 2989 984 2995 1076
rect 3021 984 3027 1056
rect 3053 1044 3059 1056
rect 2925 963 2931 976
rect 2916 957 2931 963
rect 2797 944 2803 956
rect 2813 864 2819 956
rect 2861 924 2867 956
rect 2964 937 2972 943
rect 2836 917 2844 923
rect 2861 904 2867 916
rect 2605 797 2627 803
rect 2580 737 2588 743
rect 2413 704 2419 716
rect 2477 704 2483 716
rect 2340 697 2403 703
rect 2180 677 2227 683
rect 2397 683 2403 697
rect 2436 697 2451 703
rect 2397 677 2412 683
rect 2429 664 2435 676
rect 2445 663 2451 697
rect 2525 684 2531 696
rect 2468 677 2476 683
rect 2557 664 2563 736
rect 2605 684 2611 797
rect 2653 724 2659 736
rect 2573 664 2579 676
rect 2445 657 2515 663
rect 2173 637 2188 643
rect 1981 624 1987 636
rect 2061 584 2067 636
rect 2077 584 2083 596
rect 1805 443 1811 516
rect 1821 464 1827 536
rect 1853 443 1859 476
rect 1805 437 1859 443
rect 1901 344 1907 496
rect 1933 483 1939 556
rect 1949 524 1955 556
rect 1981 543 1987 576
rect 2013 564 2019 576
rect 2029 543 2035 556
rect 1972 537 1987 543
rect 2013 537 2035 543
rect 1933 477 1955 483
rect 1949 463 1955 477
rect 1972 477 1996 483
rect 2013 483 2019 537
rect 2045 524 2051 556
rect 2061 544 2067 556
rect 2093 523 2099 596
rect 2077 517 2099 523
rect 2077 483 2083 517
rect 2109 503 2115 556
rect 2141 524 2147 636
rect 2157 544 2163 596
rect 2173 523 2179 637
rect 2189 584 2195 616
rect 2205 584 2211 656
rect 2221 603 2227 636
rect 2253 624 2259 656
rect 2285 644 2291 656
rect 2301 624 2307 656
rect 2365 624 2371 636
rect 2317 603 2323 616
rect 2221 597 2323 603
rect 2253 564 2259 576
rect 2381 564 2387 656
rect 2340 557 2348 563
rect 2157 517 2179 523
rect 2109 497 2124 503
rect 2157 503 2163 517
rect 2141 497 2163 503
rect 2141 483 2147 497
rect 2013 477 2083 483
rect 2093 477 2147 483
rect 2093 463 2099 477
rect 1949 457 2099 463
rect 2189 444 2195 496
rect 2205 444 2211 496
rect 2237 464 2243 536
rect 2285 524 2291 556
rect 2365 543 2371 556
rect 2397 544 2403 616
rect 2413 604 2419 656
rect 2477 564 2483 616
rect 2356 537 2371 543
rect 2301 464 2307 536
rect 2413 523 2419 556
rect 2452 537 2483 543
rect 2477 524 2483 537
rect 2493 524 2499 636
rect 2509 624 2515 657
rect 2541 604 2547 636
rect 2573 584 2579 596
rect 2509 543 2515 556
rect 2573 543 2579 556
rect 2605 544 2611 556
rect 2509 537 2579 543
rect 2413 517 2428 523
rect 2548 517 2604 523
rect 1988 437 1996 443
rect 2276 437 2284 443
rect 2045 384 2051 396
rect 2029 363 2035 376
rect 2061 363 2067 396
rect 2029 357 2067 363
rect 1732 337 1740 343
rect 2068 337 2076 343
rect 1789 324 1795 336
rect 1853 304 1859 336
rect 1885 324 1891 336
rect 1933 324 1939 336
rect 1661 277 1740 283
rect 1661 244 1667 256
rect 1645 164 1651 236
rect 1693 224 1699 256
rect 1693 144 1699 156
rect 1709 144 1715 236
rect 1757 224 1763 296
rect 1725 184 1731 216
rect 1789 184 1795 236
rect 1805 224 1811 256
rect 1837 244 1843 276
rect 1901 244 1907 276
rect 1876 237 1884 243
rect 1757 144 1763 156
rect 1709 124 1715 136
rect 1661 104 1667 116
rect 1581 97 1596 103
rect 669 84 675 96
rect 1261 84 1267 96
rect 1741 84 1747 96
rect 925 64 931 76
rect 1549 -43 1555 76
rect 1821 44 1827 236
rect 1869 184 1875 216
rect 1933 184 1939 316
rect 2125 284 2131 436
rect 2189 384 2195 436
rect 2333 384 2339 476
rect 2397 444 2403 516
rect 2429 464 2435 476
rect 2637 464 2643 636
rect 2669 563 2675 756
rect 2749 704 2755 736
rect 2813 724 2819 816
rect 2781 704 2787 716
rect 2708 677 2732 683
rect 2845 664 2851 896
rect 2893 884 2899 916
rect 2925 903 2931 936
rect 2941 924 2947 936
rect 2957 917 2988 923
rect 2957 903 2963 917
rect 3069 923 3075 1236
rect 3117 1224 3123 1737
rect 3133 1724 3139 1836
rect 3149 1804 3155 1856
rect 3229 1844 3235 1856
rect 3293 1844 3299 1856
rect 3165 1824 3171 1836
rect 3325 1804 3331 1896
rect 3341 1864 3347 2036
rect 3373 1844 3379 1896
rect 3405 1844 3411 1856
rect 3357 1824 3363 1836
rect 3421 1804 3427 2116
rect 3501 2104 3507 2136
rect 3533 2104 3539 2296
rect 3565 2244 3571 2496
rect 3581 2324 3587 2496
rect 3693 2324 3699 2516
rect 3741 2504 3747 2516
rect 3725 2484 3731 2496
rect 3725 2324 3731 2336
rect 3741 2304 3747 2316
rect 3741 2284 3747 2296
rect 3773 2284 3779 3036
rect 3789 2984 3795 3096
rect 4109 3064 4115 3136
rect 4125 3084 4131 3316
rect 4253 3304 4259 3356
rect 4269 3344 4275 3376
rect 4301 3304 4307 3396
rect 4365 3324 4371 3356
rect 4180 3297 4188 3303
rect 4221 3237 4236 3243
rect 4221 3104 4227 3237
rect 4301 3164 4307 3296
rect 4317 3284 4323 3296
rect 3821 3023 3827 3056
rect 3869 3044 3875 3056
rect 3981 3044 3987 3056
rect 4061 3044 4067 3056
rect 4173 3024 4179 3056
rect 3821 3017 3843 3023
rect 3805 2964 3811 2976
rect 3789 2904 3795 2956
rect 3837 2924 3843 3017
rect 4045 2984 4051 2996
rect 4061 2963 4067 2996
rect 3956 2957 4067 2963
rect 4109 2963 4115 2996
rect 4125 2984 4131 2996
rect 4141 2977 4188 2983
rect 4141 2963 4147 2977
rect 4109 2957 4147 2963
rect 3837 2904 3843 2916
rect 3853 2884 3859 2916
rect 3869 2904 3875 2916
rect 3885 2904 3891 2956
rect 4052 2937 4060 2943
rect 3933 2924 3939 2936
rect 4004 2917 4012 2923
rect 3837 2784 3843 2836
rect 3901 2804 3907 2876
rect 3965 2724 3971 2736
rect 3869 2684 3875 2696
rect 3981 2683 3987 2776
rect 4013 2704 4019 2756
rect 4029 2684 4035 2916
rect 4045 2703 4051 2756
rect 4045 2697 4060 2703
rect 3965 2677 3987 2683
rect 3789 2623 3795 2676
rect 3837 2644 3843 2656
rect 3789 2617 3811 2623
rect 3805 2484 3811 2617
rect 3869 2584 3875 2596
rect 3917 2564 3923 2636
rect 3933 2564 3939 2676
rect 3924 2517 3932 2523
rect 3821 2504 3827 2516
rect 3885 2484 3891 2516
rect 3805 2424 3811 2476
rect 3869 2304 3875 2416
rect 3885 2284 3891 2436
rect 3965 2324 3971 2677
rect 3997 2584 4003 2616
rect 4013 2584 4019 2656
rect 4029 2604 4035 2676
rect 4045 2624 4051 2636
rect 4045 2584 4051 2596
rect 4061 2564 4067 2616
rect 4077 2584 4083 2936
rect 4141 2884 4147 2916
rect 4173 2864 4179 2956
rect 4109 2703 4115 2756
rect 4125 2724 4131 2736
rect 4141 2724 4147 2836
rect 4109 2697 4131 2703
rect 4125 2604 4131 2697
rect 4173 2664 4179 2756
rect 4205 2723 4211 3096
rect 4253 3084 4259 3096
rect 4349 3084 4355 3316
rect 4413 3284 4419 3356
rect 4445 3324 4451 3416
rect 4461 3324 4467 3456
rect 4509 3444 4515 3456
rect 4525 3424 4531 3456
rect 4573 3444 4579 3456
rect 4493 3284 4499 3356
rect 4509 3324 4515 3336
rect 4557 3304 4563 3356
rect 4605 3324 4611 3476
rect 4653 3464 4659 3476
rect 4701 3364 4707 3496
rect 4797 3464 4803 3556
rect 4957 3524 4963 3683
rect 4845 3464 4851 3516
rect 4989 3504 4995 3683
rect 5053 3564 5059 3683
rect 5053 3524 5059 3556
rect 4893 3484 4899 3496
rect 4989 3484 4995 3496
rect 5037 3484 5043 3496
rect 5085 3484 5091 3496
rect 5133 3484 5139 3516
rect 4861 3464 4867 3476
rect 4749 3364 4755 3456
rect 4893 3444 4899 3476
rect 4941 3444 4947 3456
rect 4781 3364 4787 3416
rect 4637 3284 4643 3356
rect 4685 3324 4691 3356
rect 4781 3324 4787 3356
rect 4829 3344 4835 3436
rect 4877 3364 4883 3436
rect 4925 3424 4931 3436
rect 4989 3364 4995 3376
rect 5021 3364 5027 3436
rect 5085 3403 5091 3476
rect 5069 3397 5091 3403
rect 5053 3364 5059 3376
rect 4829 3324 4835 3336
rect 4877 3324 4883 3356
rect 4925 3324 4931 3336
rect 4653 3304 4659 3316
rect 4653 3264 4659 3276
rect 4653 3244 4659 3256
rect 4669 3244 4675 3296
rect 4589 3224 4595 3236
rect 4733 3204 4739 3236
rect 4525 3184 4531 3196
rect 4829 3184 4835 3236
rect 4397 3124 4403 3156
rect 4893 3144 4899 3276
rect 4429 3084 4435 3116
rect 4557 3104 4563 3116
rect 4221 3044 4227 3056
rect 4221 2944 4227 2956
rect 4253 2944 4259 3076
rect 4589 3064 4595 3096
rect 4685 3084 4691 3116
rect 4605 3064 4611 3076
rect 4701 3064 4707 3136
rect 4717 3063 4723 3116
rect 4749 3104 4755 3116
rect 4797 3104 4803 3136
rect 4909 3124 4915 3236
rect 4941 3164 4947 3356
rect 5069 3324 5075 3397
rect 5101 3384 5107 3476
rect 5165 3444 5171 3456
rect 5117 3404 5123 3436
rect 5101 3344 5107 3356
rect 5149 3344 5155 3436
rect 4973 3304 4979 3316
rect 4973 3284 4979 3296
rect 4964 3237 4972 3243
rect 4989 3183 4995 3276
rect 4973 3177 4995 3183
rect 4845 3104 4851 3116
rect 4925 3104 4931 3116
rect 4973 3104 4979 3177
rect 4733 3084 4739 3096
rect 4989 3064 4995 3156
rect 4717 3057 4732 3063
rect 4333 3044 4339 3056
rect 4349 3024 4355 3056
rect 4269 2964 4275 2996
rect 4285 2984 4291 3016
rect 4413 3004 4419 3036
rect 4461 2984 4467 3056
rect 4557 3044 4563 3056
rect 4605 3044 4611 3056
rect 4781 3044 4787 3056
rect 4477 3037 4492 3043
rect 4333 2977 4396 2983
rect 4333 2964 4339 2977
rect 4349 2924 4355 2956
rect 4381 2924 4387 2956
rect 4301 2904 4307 2916
rect 4429 2904 4435 2936
rect 4317 2824 4323 2836
rect 4189 2717 4211 2723
rect 4173 2584 4179 2596
rect 4061 2544 4067 2556
rect 3981 2464 3987 2536
rect 4077 2523 4083 2556
rect 4109 2544 4115 2556
rect 4125 2524 4131 2556
rect 4157 2544 4163 2556
rect 4189 2543 4195 2717
rect 4205 2624 4211 2696
rect 4237 2664 4243 2816
rect 4397 2804 4403 2876
rect 4404 2757 4412 2763
rect 4349 2744 4355 2756
rect 4429 2723 4435 2896
rect 4477 2884 4483 3037
rect 4660 3037 4668 3043
rect 4717 3024 4723 3036
rect 4493 2964 4499 2996
rect 4573 2984 4579 2996
rect 4653 2977 4691 2983
rect 4493 2924 4499 2936
rect 4525 2924 4531 2956
rect 4653 2944 4659 2977
rect 4621 2923 4627 2936
rect 4621 2917 4652 2923
rect 4493 2724 4499 2916
rect 4509 2764 4515 2836
rect 4621 2784 4627 2876
rect 4669 2824 4675 2956
rect 4685 2904 4691 2977
rect 4797 2964 4803 3056
rect 4829 3044 4835 3056
rect 4877 3044 4883 3056
rect 4717 2944 4723 2956
rect 4813 2944 4819 3036
rect 4701 2924 4707 2936
rect 4765 2924 4771 2936
rect 4749 2904 4755 2916
rect 4813 2884 4819 2896
rect 4429 2717 4444 2723
rect 4781 2723 4787 2836
rect 4813 2744 4819 2856
rect 4829 2744 4835 2836
rect 4765 2717 4787 2723
rect 4285 2663 4291 2696
rect 4301 2684 4307 2716
rect 4765 2704 4771 2717
rect 4365 2697 4380 2703
rect 4365 2684 4371 2697
rect 4868 2697 4876 2703
rect 4781 2684 4787 2696
rect 4484 2677 4492 2683
rect 4317 2663 4323 2676
rect 4637 2664 4643 2676
rect 4285 2657 4323 2663
rect 4740 2657 4755 2663
rect 4237 2584 4243 2656
rect 4253 2624 4259 2656
rect 4173 2537 4195 2543
rect 4173 2524 4179 2537
rect 4068 2517 4083 2523
rect 4084 2497 4092 2503
rect 4132 2497 4140 2503
rect 3981 2303 3987 2456
rect 4029 2424 4035 2496
rect 4189 2484 4195 2516
rect 4077 2424 4083 2436
rect 3997 2383 4003 2416
rect 3997 2377 4012 2383
rect 4077 2304 4083 2416
rect 4093 2324 4099 2436
rect 4125 2324 4131 2336
rect 4141 2304 4147 2336
rect 4189 2324 4195 2476
rect 4253 2404 4259 2556
rect 4269 2424 4275 2636
rect 4317 2623 4323 2636
rect 4317 2617 4339 2623
rect 4317 2584 4323 2596
rect 4301 2544 4307 2576
rect 4333 2524 4339 2617
rect 4349 2584 4355 2636
rect 4429 2624 4435 2656
rect 4445 2624 4451 2636
rect 4493 2604 4499 2636
rect 4573 2604 4579 2656
rect 4685 2644 4691 2656
rect 4365 2563 4371 2576
rect 4605 2564 4611 2576
rect 4356 2557 4371 2563
rect 4445 2557 4483 2563
rect 4285 2504 4291 2516
rect 4333 2424 4339 2496
rect 4253 2324 4259 2336
rect 3965 2297 3987 2303
rect 3588 2277 3596 2283
rect 3684 2277 3692 2283
rect 3796 2257 3804 2263
rect 3581 2244 3587 2256
rect 3773 2244 3779 2256
rect 3661 2224 3667 2236
rect 3565 2164 3571 2216
rect 3549 2124 3555 2156
rect 3645 2144 3651 2216
rect 3725 2177 3756 2183
rect 3725 2143 3731 2177
rect 3741 2144 3747 2156
rect 3693 2137 3731 2143
rect 3661 2104 3667 2136
rect 3693 2104 3699 2137
rect 3757 2123 3763 2156
rect 3716 2117 3763 2123
rect 3620 2097 3644 2103
rect 3469 2044 3475 2096
rect 3533 2024 3539 2036
rect 3437 1984 3443 2016
rect 3453 1924 3459 1936
rect 3469 1904 3475 1976
rect 3549 1943 3555 2096
rect 3709 2044 3715 2096
rect 3636 2037 3644 2043
rect 3597 2024 3603 2036
rect 3661 1984 3667 2036
rect 3741 2024 3747 2076
rect 3572 1977 3603 1983
rect 3597 1963 3603 1977
rect 3629 1963 3635 1976
rect 3597 1957 3635 1963
rect 3549 1937 3571 1943
rect 3485 1884 3491 1896
rect 3549 1884 3555 1916
rect 3565 1884 3571 1937
rect 3581 1904 3587 1916
rect 3597 1904 3603 1916
rect 3677 1884 3683 1976
rect 3773 1943 3779 2216
rect 3789 2144 3795 2216
rect 3837 2144 3843 2256
rect 3924 2237 3939 2243
rect 3933 2223 3939 2237
rect 3933 2217 3948 2223
rect 3860 2157 3884 2163
rect 3917 2144 3923 2216
rect 3789 1964 3795 2116
rect 3885 2064 3891 2096
rect 3869 2024 3875 2036
rect 3933 2024 3939 2136
rect 3965 2104 3971 2297
rect 4029 2264 4035 2276
rect 4084 2257 4092 2263
rect 4045 2224 4051 2256
rect 4173 2244 4179 2256
rect 3981 2177 4051 2183
rect 3981 2144 3987 2177
rect 4045 2164 4051 2177
rect 4013 2144 4019 2156
rect 3981 2064 3987 2096
rect 3933 1964 3939 2016
rect 4029 1984 4035 2156
rect 4061 2124 4067 2176
rect 4077 2163 4083 2236
rect 4093 2184 4099 2196
rect 4189 2184 4195 2216
rect 4205 2164 4211 2236
rect 4221 2184 4227 2196
rect 4237 2164 4243 2296
rect 4413 2284 4419 2536
rect 4445 2524 4451 2557
rect 4477 2544 4483 2557
rect 4653 2544 4659 2556
rect 4461 2524 4467 2536
rect 4525 2524 4531 2536
rect 4717 2524 4723 2656
rect 4749 2544 4755 2657
rect 4845 2544 4851 2636
rect 4893 2604 4899 3016
rect 4909 3004 4915 3036
rect 4941 2964 4947 2976
rect 4957 2964 4963 3056
rect 4989 3044 4995 3056
rect 4941 2924 4947 2956
rect 5005 2924 5011 3256
rect 5124 3237 5132 3243
rect 5021 3104 5027 3236
rect 5037 3224 5043 3236
rect 5021 3084 5027 3096
rect 5021 2924 5027 3056
rect 5037 2964 5043 3176
rect 5069 3064 5075 3176
rect 5165 3104 5171 3116
rect 5117 3044 5123 3056
rect 5053 2984 5059 3036
rect 5101 2964 5107 3036
rect 5101 2924 5107 2936
rect 5133 2923 5139 3096
rect 5117 2917 5139 2923
rect 4925 2644 4931 2696
rect 4957 2684 4963 2916
rect 5005 2824 5011 2836
rect 5069 2744 5075 2896
rect 5117 2864 5123 2917
rect 4973 2704 4979 2716
rect 5069 2664 5075 2676
rect 4957 2644 4963 2656
rect 5021 2624 5027 2636
rect 5117 2604 5123 2836
rect 5005 2564 5011 2596
rect 5133 2563 5139 2876
rect 5149 2764 5155 2876
rect 5165 2824 5171 2836
rect 5181 2804 5187 2936
rect 5165 2744 5171 2796
rect 5197 2624 5203 3056
rect 5156 2577 5164 2583
rect 5133 2557 5148 2563
rect 4733 2537 4748 2543
rect 4500 2517 4508 2523
rect 4605 2504 4611 2516
rect 4509 2284 4515 2436
rect 4477 2264 4483 2276
rect 4525 2264 4531 2316
rect 4621 2284 4627 2516
rect 4701 2423 4707 2476
rect 4717 2464 4723 2496
rect 4733 2424 4739 2537
rect 4765 2524 4771 2536
rect 4893 2524 4899 2536
rect 4941 2524 4947 2536
rect 4957 2504 4963 2516
rect 4916 2497 4940 2503
rect 4989 2503 4995 2556
rect 5053 2524 5059 2536
rect 5101 2504 5107 2556
rect 5133 2504 5139 2536
rect 5181 2504 5187 2516
rect 4973 2497 4995 2503
rect 4861 2424 4867 2496
rect 4973 2484 4979 2497
rect 5060 2477 5068 2483
rect 4701 2417 4723 2423
rect 4644 2317 4652 2323
rect 4644 2277 4652 2283
rect 4557 2264 4563 2276
rect 4381 2257 4396 2263
rect 4381 2224 4387 2257
rect 4413 2224 4419 2256
rect 4445 2204 4451 2256
rect 4605 2223 4611 2276
rect 4685 2264 4691 2316
rect 4637 2224 4643 2236
rect 4605 2217 4627 2223
rect 4301 2197 4355 2203
rect 4301 2184 4307 2197
rect 4077 2157 4099 2163
rect 4077 2104 4083 2116
rect 4093 2064 4099 2157
rect 4260 2157 4268 2163
rect 4125 2144 4131 2156
rect 4317 2144 4323 2156
rect 4157 2104 4163 2136
rect 4237 2124 4243 2136
rect 4205 2104 4211 2116
rect 4285 2104 4291 2136
rect 4333 2124 4339 2176
rect 4349 2163 4355 2197
rect 4381 2164 4387 2196
rect 4349 2157 4364 2163
rect 4180 2097 4188 2103
rect 3981 1944 3987 1976
rect 3773 1937 3891 1943
rect 3757 1917 3820 1923
rect 3757 1903 3763 1917
rect 3885 1923 3891 1937
rect 4061 1924 4067 1996
rect 4077 1924 4083 1956
rect 3885 1917 3916 1923
rect 3997 1917 4012 1923
rect 3725 1897 3763 1903
rect 3213 1784 3219 1796
rect 3357 1764 3363 1796
rect 3396 1757 3427 1763
rect 3229 1704 3235 1756
rect 3261 1724 3267 1736
rect 3341 1704 3347 1716
rect 3300 1697 3308 1703
rect 3405 1684 3411 1736
rect 3421 1683 3427 1757
rect 3485 1724 3491 1856
rect 3501 1844 3507 1856
rect 3533 1764 3539 1876
rect 3725 1864 3731 1897
rect 3741 1844 3747 1856
rect 3773 1824 3779 1896
rect 3789 1864 3795 1876
rect 3869 1864 3875 1916
rect 3997 1903 4003 1917
rect 4093 1923 4099 2036
rect 4157 1944 4163 2076
rect 4205 1944 4211 1956
rect 4253 1924 4259 1936
rect 4093 1917 4131 1923
rect 3988 1897 4003 1903
rect 4077 1897 4108 1903
rect 3549 1764 3555 1776
rect 3485 1704 3491 1716
rect 3501 1704 3507 1756
rect 3581 1724 3587 1756
rect 3597 1724 3603 1816
rect 3917 1764 3923 1836
rect 3933 1784 3939 1876
rect 4029 1863 4035 1876
rect 4077 1864 4083 1897
rect 4125 1903 4131 1917
rect 4125 1897 4163 1903
rect 4157 1884 4163 1897
rect 4269 1903 4275 2036
rect 4413 1984 4419 2196
rect 4477 2184 4483 2216
rect 4525 2183 4531 2196
rect 4589 2184 4595 2196
rect 4621 2184 4627 2217
rect 4525 2177 4547 2183
rect 4541 2164 4547 2177
rect 4605 2144 4611 2156
rect 4653 2144 4659 2256
rect 4445 2044 4451 2136
rect 4461 2124 4467 2136
rect 4541 2124 4547 2136
rect 4669 2123 4675 2236
rect 4653 2117 4675 2123
rect 4589 2104 4595 2116
rect 4637 2104 4643 2116
rect 4493 2084 4499 2096
rect 4445 2003 4451 2036
rect 4509 2024 4515 2036
rect 4429 1997 4451 2003
rect 4292 1957 4300 1963
rect 4349 1924 4355 1956
rect 4253 1897 4275 1903
rect 4221 1884 4227 1896
rect 4109 1864 4115 1876
rect 4013 1857 4035 1863
rect 3949 1784 3955 1796
rect 3965 1784 3971 1836
rect 3805 1757 3820 1763
rect 3725 1744 3731 1756
rect 3741 1744 3747 1756
rect 3677 1723 3683 1736
rect 3613 1717 3683 1723
rect 3613 1703 3619 1717
rect 3565 1697 3619 1703
rect 3709 1703 3715 1736
rect 3757 1703 3763 1736
rect 3789 1724 3795 1736
rect 3773 1704 3779 1716
rect 3709 1697 3763 1703
rect 3565 1683 3571 1697
rect 3421 1677 3571 1683
rect 3805 1683 3811 1757
rect 3837 1724 3843 1756
rect 3885 1744 3891 1756
rect 3981 1744 3987 1836
rect 3853 1704 3859 1736
rect 3869 1724 3875 1736
rect 3805 1677 3827 1683
rect 3821 1644 3827 1677
rect 3245 1624 3251 1636
rect 3149 1597 3267 1603
rect 3149 1584 3155 1597
rect 3261 1583 3267 1597
rect 3389 1584 3395 1616
rect 3485 1584 3491 1596
rect 3261 1577 3324 1583
rect 3252 1537 3260 1543
rect 3149 1524 3155 1536
rect 3133 1384 3139 1476
rect 3149 1384 3155 1516
rect 3229 1504 3235 1536
rect 3277 1503 3283 1536
rect 3300 1517 3308 1523
rect 3277 1497 3299 1503
rect 3165 1424 3171 1436
rect 3181 1404 3187 1476
rect 3197 1424 3203 1456
rect 3213 1424 3219 1436
rect 3261 1423 3267 1456
rect 3277 1444 3283 1456
rect 3293 1423 3299 1497
rect 3309 1444 3315 1496
rect 3373 1464 3379 1536
rect 3469 1484 3475 1516
rect 3453 1463 3459 1476
rect 3517 1464 3523 1616
rect 3453 1457 3475 1463
rect 3341 1444 3347 1456
rect 3405 1444 3411 1456
rect 3469 1444 3475 1457
rect 3261 1417 3283 1423
rect 3293 1417 3315 1423
rect 3165 1344 3171 1396
rect 3277 1383 3283 1417
rect 3277 1377 3292 1383
rect 3309 1383 3315 1417
rect 3405 1384 3411 1396
rect 3309 1377 3356 1383
rect 3261 1364 3267 1376
rect 3165 1184 3171 1276
rect 3197 1224 3203 1356
rect 3437 1344 3443 1436
rect 3453 1384 3459 1436
rect 3485 1344 3491 1376
rect 3501 1344 3507 1356
rect 3293 1324 3299 1336
rect 3213 1304 3219 1316
rect 3245 1244 3251 1316
rect 3389 1304 3395 1316
rect 3412 1297 3427 1303
rect 3277 1224 3283 1236
rect 3277 1144 3283 1176
rect 3316 1137 3324 1143
rect 3277 1124 3283 1136
rect 3405 1124 3411 1196
rect 3421 1144 3427 1297
rect 3453 1284 3459 1296
rect 3501 1124 3507 1276
rect 3533 1224 3539 1596
rect 3549 1504 3555 1536
rect 3549 1444 3555 1496
rect 3565 1484 3571 1496
rect 3597 1464 3603 1576
rect 3581 1424 3587 1436
rect 3613 1404 3619 1436
rect 3645 1424 3651 1516
rect 3677 1484 3683 1536
rect 3693 1464 3699 1596
rect 3757 1464 3763 1596
rect 3773 1464 3779 1616
rect 3789 1584 3795 1616
rect 3805 1503 3811 1636
rect 3869 1604 3875 1616
rect 3869 1584 3875 1596
rect 3805 1497 3827 1503
rect 3805 1464 3811 1476
rect 3709 1424 3715 1436
rect 3597 1383 3603 1396
rect 3597 1377 3612 1383
rect 3581 1344 3587 1356
rect 3645 1344 3651 1416
rect 3725 1397 3763 1403
rect 3725 1383 3731 1397
rect 3757 1384 3763 1397
rect 3709 1377 3731 1383
rect 3709 1343 3715 1377
rect 3661 1337 3715 1343
rect 3581 1223 3587 1296
rect 3597 1264 3603 1336
rect 3661 1303 3667 1337
rect 3741 1324 3747 1356
rect 3773 1344 3779 1356
rect 3780 1317 3788 1323
rect 3677 1304 3683 1316
rect 3652 1297 3667 1303
rect 3565 1217 3587 1223
rect 3565 1144 3571 1217
rect 3629 1184 3635 1196
rect 3645 1124 3651 1236
rect 3677 1143 3683 1196
rect 3693 1164 3699 1316
rect 3741 1244 3747 1276
rect 3709 1224 3715 1236
rect 3821 1224 3827 1497
rect 3837 1484 3843 1516
rect 3837 1344 3843 1356
rect 3885 1344 3891 1416
rect 3901 1384 3907 1636
rect 3965 1544 3971 1736
rect 4013 1643 4019 1857
rect 4036 1797 4067 1803
rect 4061 1764 4067 1797
rect 4077 1784 4083 1836
rect 3997 1637 4019 1643
rect 3965 1484 3971 1496
rect 3981 1424 3987 1476
rect 3997 1424 4003 1637
rect 4029 1584 4035 1716
rect 4029 1503 4035 1516
rect 4020 1497 4035 1503
rect 4045 1424 4051 1596
rect 4077 1524 4083 1736
rect 4125 1704 4131 1716
rect 4141 1604 4147 1836
rect 4180 1797 4195 1803
rect 4189 1784 4195 1797
rect 4205 1724 4211 1836
rect 4221 1784 4227 1796
rect 4157 1684 4163 1696
rect 4173 1604 4179 1716
rect 4205 1644 4211 1696
rect 4205 1584 4211 1596
rect 4100 1517 4108 1523
rect 4061 1484 4067 1516
rect 4189 1504 4195 1516
rect 4093 1484 4099 1496
rect 4141 1484 4147 1496
rect 4068 1457 4076 1463
rect 4116 1457 4124 1463
rect 3949 1403 3955 1416
rect 3917 1397 3955 1403
rect 4029 1403 4035 1416
rect 4029 1397 4083 1403
rect 3917 1384 3923 1397
rect 4029 1377 4067 1383
rect 4029 1364 4035 1377
rect 4061 1364 4067 1377
rect 3949 1357 3964 1363
rect 3869 1324 3875 1336
rect 3949 1304 3955 1357
rect 3997 1344 4003 1356
rect 4045 1344 4051 1356
rect 4077 1344 4083 1397
rect 4141 1364 4147 1456
rect 4173 1384 4179 1416
rect 4189 1383 4195 1436
rect 4253 1424 4259 1897
rect 4429 1884 4435 1997
rect 4541 1944 4547 1976
rect 4653 1944 4659 2117
rect 4685 2084 4691 2096
rect 4717 2083 4723 2417
rect 4749 2384 4755 2416
rect 4765 2244 4771 2276
rect 4813 2264 4819 2376
rect 4925 2344 4931 2436
rect 5037 2364 5043 2436
rect 4941 2344 4947 2356
rect 5037 2324 5043 2336
rect 4861 2304 4867 2316
rect 4765 2204 4771 2236
rect 4781 2224 4787 2256
rect 4797 2224 4803 2256
rect 4781 2124 4787 2176
rect 4797 2144 4803 2156
rect 4845 2144 4851 2196
rect 4829 2124 4835 2136
rect 4701 2077 4723 2083
rect 4605 1904 4611 1916
rect 4317 1864 4323 1876
rect 4445 1864 4451 1896
rect 4493 1884 4499 1896
rect 4637 1884 4643 1936
rect 4669 1884 4675 2036
rect 4701 1884 4707 2077
rect 4749 1924 4755 1936
rect 4829 1924 4835 2056
rect 4861 1884 4867 2256
rect 4877 2184 4883 2216
rect 4893 2204 4899 2256
rect 4909 2203 4915 2276
rect 4957 2224 4963 2316
rect 5053 2304 5059 2316
rect 4989 2264 4995 2276
rect 4909 2197 4931 2203
rect 4893 2144 4899 2156
rect 4925 2144 4931 2197
rect 4973 2164 4979 2216
rect 5005 2204 5011 2276
rect 5021 2144 5027 2156
rect 5037 2144 5043 2236
rect 5053 2184 5059 2196
rect 4941 2124 4947 2136
rect 4877 2063 4883 2096
rect 5005 2084 5011 2096
rect 4877 2057 4899 2063
rect 4893 1884 4899 2057
rect 4941 1943 4947 2036
rect 4973 1984 4979 1996
rect 4932 1937 4947 1943
rect 5053 1884 5059 2136
rect 5069 2124 5075 2236
rect 5101 2184 5107 2276
rect 5117 2224 5123 2436
rect 5133 2264 5139 2296
rect 5149 2264 5155 2276
rect 5069 2024 5075 2096
rect 5085 2004 5091 2136
rect 5117 2124 5123 2136
rect 5101 1924 5107 1956
rect 4541 1864 4547 1876
rect 4644 1857 4652 1863
rect 4365 1844 4371 1856
rect 4477 1844 4483 1856
rect 4404 1837 4412 1843
rect 4349 1804 4355 1836
rect 4301 1777 4332 1783
rect 4301 1763 4307 1777
rect 4365 1764 4371 1776
rect 4285 1757 4307 1763
rect 4269 1724 4275 1736
rect 4285 1703 4291 1757
rect 4317 1744 4323 1756
rect 4301 1704 4307 1736
rect 4413 1724 4419 1816
rect 4445 1764 4451 1776
rect 4365 1704 4371 1716
rect 4276 1697 4291 1703
rect 4349 1684 4355 1696
rect 4397 1664 4403 1716
rect 4509 1704 4515 1716
rect 4429 1684 4435 1696
rect 4413 1664 4419 1676
rect 4413 1644 4419 1656
rect 4269 1504 4275 1516
rect 4285 1483 4291 1516
rect 4333 1484 4339 1596
rect 4461 1504 4467 1556
rect 4381 1497 4412 1503
rect 4381 1484 4387 1497
rect 4493 1484 4499 1516
rect 4285 1477 4323 1483
rect 4276 1457 4284 1463
rect 4317 1463 4323 1477
rect 4317 1457 4332 1463
rect 4381 1424 4387 1456
rect 4413 1444 4419 1456
rect 4461 1404 4467 1476
rect 4525 1424 4531 1836
rect 4541 1744 4547 1856
rect 4573 1844 4579 1856
rect 4573 1784 4579 1836
rect 4685 1804 4691 1836
rect 4589 1764 4595 1776
rect 4781 1744 4787 1836
rect 4797 1823 4803 1876
rect 4852 1837 4860 1843
rect 4877 1824 4883 1876
rect 4797 1817 4819 1823
rect 4797 1744 4803 1776
rect 4813 1763 4819 1817
rect 4829 1784 4835 1816
rect 4813 1757 4860 1763
rect 4596 1737 4604 1743
rect 4644 1737 4652 1743
rect 4813 1737 4828 1743
rect 4813 1723 4819 1737
rect 4893 1723 4899 1836
rect 4925 1744 4931 1796
rect 4989 1744 4995 1756
rect 4964 1737 4972 1743
rect 4756 1717 4819 1723
rect 4877 1717 4899 1723
rect 4685 1704 4691 1716
rect 4621 1584 4627 1596
rect 4548 1537 4563 1543
rect 4557 1504 4563 1537
rect 4589 1504 4595 1516
rect 4605 1504 4611 1516
rect 4637 1504 4643 1696
rect 4733 1584 4739 1696
rect 4749 1644 4755 1696
rect 4765 1604 4771 1636
rect 4557 1464 4563 1476
rect 4189 1377 4227 1383
rect 4205 1344 4211 1356
rect 4221 1344 4227 1377
rect 4637 1364 4643 1476
rect 4669 1424 4675 1436
rect 4733 1423 4739 1496
rect 4749 1464 4755 1476
rect 4781 1444 4787 1516
rect 4797 1504 4803 1656
rect 4829 1464 4835 1676
rect 4877 1563 4883 1717
rect 4925 1704 4931 1736
rect 4893 1624 4899 1696
rect 4861 1557 4883 1563
rect 4845 1524 4851 1536
rect 4861 1463 4867 1557
rect 4877 1484 4883 1536
rect 4893 1524 4899 1576
rect 5037 1543 5043 1716
rect 5053 1664 5059 1856
rect 5069 1784 5075 1796
rect 5085 1704 5091 1876
rect 5117 1784 5123 2056
rect 5133 1964 5139 2236
rect 5149 2064 5155 2236
rect 5149 1964 5155 2036
rect 5133 1863 5139 1916
rect 5149 1884 5155 1916
rect 5133 1857 5155 1863
rect 5133 1764 5139 1836
rect 5149 1784 5155 1857
rect 5165 1803 5171 1836
rect 5165 1797 5187 1803
rect 5069 1604 5075 1676
rect 5101 1584 5107 1736
rect 5117 1543 5123 1736
rect 5133 1724 5139 1736
rect 5149 1544 5155 1756
rect 5037 1537 5059 1543
rect 5037 1504 5043 1516
rect 4941 1484 4947 1496
rect 4861 1457 4883 1463
rect 4717 1417 4739 1423
rect 4685 1364 4691 1396
rect 4717 1364 4723 1417
rect 4733 1364 4739 1376
rect 4861 1364 4867 1436
rect 4877 1424 4883 1457
rect 4877 1384 4883 1396
rect 4404 1357 4412 1363
rect 4500 1357 4508 1363
rect 4132 1337 4195 1343
rect 4045 1303 4051 1316
rect 4036 1297 4051 1303
rect 3917 1224 3923 1296
rect 3773 1184 3779 1196
rect 3837 1184 3843 1196
rect 3725 1177 3763 1183
rect 3725 1143 3731 1177
rect 3677 1137 3731 1143
rect 3101 1004 3107 1096
rect 3165 1063 3171 1096
rect 3181 1084 3187 1116
rect 3293 1097 3459 1103
rect 3293 1083 3299 1097
rect 3453 1084 3459 1097
rect 3284 1077 3299 1083
rect 3156 1057 3171 1063
rect 3188 1057 3228 1063
rect 3325 1044 3331 1076
rect 3357 1044 3363 1076
rect 3421 1044 3427 1076
rect 3284 1037 3292 1043
rect 3053 917 3075 923
rect 2925 897 2963 903
rect 3005 883 3011 896
rect 2964 877 3011 883
rect 2973 823 2979 836
rect 2973 817 2995 823
rect 2861 684 2867 816
rect 2989 803 2995 817
rect 2989 797 3011 803
rect 3005 724 3011 797
rect 3021 784 3027 816
rect 3053 764 3059 917
rect 3133 904 3139 956
rect 3181 904 3187 916
rect 2909 684 2915 696
rect 2973 684 2979 696
rect 3021 684 3027 696
rect 2877 664 2883 676
rect 3069 664 3075 776
rect 3117 704 3123 856
rect 3197 844 3203 1036
rect 3213 944 3219 1036
rect 3261 944 3267 956
rect 3309 944 3315 1016
rect 3229 903 3235 916
rect 3229 897 3260 903
rect 3293 844 3299 876
rect 3181 784 3187 836
rect 3229 784 3235 796
rect 3181 724 3187 776
rect 3156 697 3171 703
rect 2756 657 2780 663
rect 2701 624 2707 656
rect 3053 644 3059 656
rect 3101 644 3107 656
rect 2829 624 2835 636
rect 2660 557 2675 563
rect 2717 544 2723 616
rect 2813 564 2819 596
rect 2861 584 2867 616
rect 2877 564 2883 596
rect 2676 537 2691 543
rect 2685 524 2691 537
rect 2669 504 2675 516
rect 2701 484 2707 536
rect 2797 504 2803 516
rect 2845 504 2851 516
rect 2701 444 2707 476
rect 2141 324 2147 336
rect 2205 304 2211 316
rect 2180 297 2188 303
rect 1988 277 1996 283
rect 1965 264 1971 276
rect 1981 244 1987 256
rect 2029 244 2035 256
rect 2093 244 2099 276
rect 2068 237 2076 243
rect 1949 204 1955 236
rect 1869 157 1907 163
rect 1869 144 1875 157
rect 1901 144 1907 157
rect 1860 137 1868 143
rect 1885 104 1891 136
rect 1901 123 1907 136
rect 1901 117 1932 123
rect 1885 -43 1891 96
rect 1933 64 1939 76
rect 1981 64 1987 156
rect 1997 144 2003 236
rect 2013 184 2019 216
rect 2052 177 2060 183
rect 2029 164 2035 176
rect 2093 164 2099 196
rect 2109 184 2115 196
rect 2141 184 2147 296
rect 2205 264 2211 296
rect 2269 264 2275 336
rect 2333 324 2339 336
rect 2621 324 2627 336
rect 2509 304 2515 316
rect 2420 297 2428 303
rect 2285 264 2291 276
rect 2317 264 2323 276
rect 2237 184 2243 196
rect 2125 144 2131 176
rect 2221 164 2227 176
rect 2253 164 2259 236
rect 2365 203 2371 296
rect 2349 197 2371 203
rect 2004 117 2019 123
rect 1997 64 2003 76
rect 1997 44 2003 56
rect 1997 24 2003 36
rect 2013 24 2019 117
rect 2045 104 2051 136
rect 2093 124 2099 136
rect 2125 104 2131 136
rect 2173 104 2179 136
rect 2285 124 2291 196
rect 2349 184 2355 197
rect 2381 164 2387 276
rect 2404 257 2412 263
rect 2397 224 2403 236
rect 2429 184 2435 276
rect 2461 224 2467 296
rect 2525 284 2531 296
rect 2477 264 2483 276
rect 2445 184 2451 216
rect 2381 144 2387 156
rect 2413 104 2419 116
rect 2429 104 2435 176
rect 2429 84 2435 96
rect 2461 84 2467 136
rect 2477 104 2483 196
rect 2493 184 2499 196
rect 2509 144 2515 276
rect 2573 244 2579 276
rect 2525 124 2531 236
rect 2573 184 2579 196
rect 2637 164 2643 436
rect 2733 404 2739 436
rect 2829 404 2835 436
rect 2893 404 2899 536
rect 2925 523 2931 636
rect 2989 524 2995 636
rect 3005 584 3011 616
rect 3117 564 3123 696
rect 3149 644 3155 656
rect 3165 624 3171 697
rect 3261 664 3267 836
rect 3341 744 3347 896
rect 3357 864 3363 936
rect 3373 903 3379 956
rect 3389 923 3395 1036
rect 3453 984 3459 1016
rect 3469 1003 3475 1116
rect 3741 1104 3747 1156
rect 3757 1123 3763 1177
rect 3917 1177 3971 1183
rect 3773 1164 3779 1176
rect 3917 1163 3923 1177
rect 3908 1157 3923 1163
rect 3773 1144 3779 1156
rect 3965 1144 3971 1177
rect 3805 1137 3884 1143
rect 3757 1117 3795 1123
rect 3789 1104 3795 1117
rect 3517 1064 3523 1096
rect 3549 1084 3555 1096
rect 3597 1084 3603 1096
rect 3700 1077 3772 1083
rect 3805 1064 3811 1137
rect 3869 1117 3916 1123
rect 3684 1057 3692 1063
rect 3732 1057 3740 1063
rect 3517 1044 3523 1056
rect 3613 1037 3644 1043
rect 3469 997 3491 1003
rect 3485 984 3491 997
rect 3405 964 3411 976
rect 3469 964 3475 976
rect 3501 964 3507 1036
rect 3565 1004 3571 1036
rect 3613 1024 3619 1037
rect 3629 964 3635 1016
rect 3661 1003 3667 1056
rect 3821 1044 3827 1056
rect 3661 997 3699 1003
rect 3693 984 3699 997
rect 3389 917 3411 923
rect 3373 897 3388 903
rect 3373 784 3379 796
rect 3389 744 3395 756
rect 3293 704 3299 716
rect 3405 684 3411 917
rect 3469 803 3475 956
rect 3485 904 3491 956
rect 3533 944 3539 956
rect 3613 944 3619 956
rect 3565 904 3571 936
rect 3453 797 3475 803
rect 3437 724 3443 756
rect 3213 644 3219 656
rect 3245 624 3251 656
rect 3261 644 3267 656
rect 3133 584 3139 616
rect 3133 564 3139 576
rect 2909 517 2931 523
rect 2909 424 2915 517
rect 2973 504 2979 516
rect 3037 504 3043 516
rect 2925 484 2931 496
rect 2925 403 2931 416
rect 3037 404 3043 496
rect 2909 397 2931 403
rect 2653 284 2659 356
rect 2909 344 2915 397
rect 2957 384 2963 396
rect 3069 364 3075 556
rect 3085 544 3091 556
rect 3117 504 3123 516
rect 2685 303 2691 336
rect 2813 324 2819 336
rect 2717 304 2723 316
rect 2669 297 2691 303
rect 2669 224 2675 297
rect 2708 277 2716 283
rect 2685 263 2691 276
rect 2733 263 2739 276
rect 2765 264 2771 276
rect 2797 264 2803 296
rect 2685 257 2739 263
rect 2685 204 2691 236
rect 2733 224 2739 236
rect 2653 144 2659 156
rect 2749 144 2755 256
rect 2781 224 2787 236
rect 2813 223 2819 296
rect 2845 284 2851 316
rect 2893 284 2899 296
rect 2916 277 2972 283
rect 3005 264 3011 276
rect 2925 257 2940 263
rect 2829 243 2835 256
rect 2909 243 2915 256
rect 2829 237 2915 243
rect 2925 224 2931 257
rect 2813 217 2835 223
rect 2765 184 2771 196
rect 2829 144 2835 217
rect 2845 164 2851 196
rect 2877 184 2883 196
rect 2893 163 2899 216
rect 2925 184 2931 196
rect 2877 157 2899 163
rect 2573 124 2579 136
rect 2829 124 2835 136
rect 2525 84 2531 116
rect 2557 104 2563 116
rect 2029 -43 2035 16
rect 2525 -43 2531 76
rect 2605 -43 2611 116
rect 2685 104 2691 116
rect 2797 104 2803 116
rect 2877 104 2883 157
rect 2957 144 2963 216
rect 2973 184 2979 256
rect 3005 224 3011 236
rect 3005 144 3011 196
rect 3021 144 3027 256
rect 3037 184 3043 216
rect 3053 144 3059 356
rect 3085 324 3091 436
rect 3117 384 3123 476
rect 3133 464 3139 516
rect 3149 504 3155 596
rect 3165 564 3171 616
rect 3165 524 3171 536
rect 3229 524 3235 616
rect 3277 544 3283 556
rect 3309 544 3315 556
rect 3325 543 3331 636
rect 3341 604 3347 676
rect 3453 664 3459 797
rect 3501 704 3507 836
rect 3581 824 3587 876
rect 3597 804 3603 836
rect 3533 724 3539 796
rect 3629 744 3635 956
rect 3661 924 3667 956
rect 3677 944 3683 956
rect 3709 943 3715 1036
rect 3837 1024 3843 1096
rect 3869 1083 3875 1117
rect 3940 1097 3955 1103
rect 3853 1077 3875 1083
rect 3725 964 3731 1016
rect 3741 977 3827 983
rect 3709 937 3731 943
rect 3725 904 3731 937
rect 3741 883 3747 977
rect 3757 943 3763 956
rect 3757 937 3804 943
rect 3757 904 3763 916
rect 3773 904 3779 916
rect 3805 904 3811 916
rect 3821 904 3827 977
rect 3853 904 3859 1077
rect 3933 1064 3939 1076
rect 3949 1064 3955 1097
rect 3981 1064 3987 1156
rect 4061 1084 4067 1156
rect 4077 1144 4083 1216
rect 4093 1184 4099 1336
rect 4189 1324 4195 1337
rect 4301 1324 4307 1356
rect 4445 1344 4451 1356
rect 4637 1344 4643 1356
rect 4701 1343 4707 1356
rect 4909 1344 4915 1436
rect 4925 1384 4931 1476
rect 4980 1457 4988 1463
rect 5012 1457 5020 1463
rect 5021 1364 5027 1376
rect 4701 1337 4716 1343
rect 4173 1304 4179 1316
rect 4125 1284 4131 1296
rect 4109 1144 4115 1156
rect 3869 1044 3875 1056
rect 3885 1044 3891 1056
rect 3885 903 3891 1016
rect 3901 924 3907 1036
rect 3924 977 3971 983
rect 3965 944 3971 977
rect 3924 937 3939 943
rect 3933 924 3939 937
rect 3949 924 3955 936
rect 3997 924 4003 956
rect 4013 944 4019 956
rect 4045 944 4051 1016
rect 3885 897 3907 903
rect 3716 877 3747 883
rect 3709 857 3740 863
rect 3709 784 3715 857
rect 3853 844 3859 876
rect 3901 863 3907 897
rect 3917 884 3923 916
rect 3901 857 3932 863
rect 3773 743 3779 836
rect 3853 804 3859 836
rect 4013 824 4019 896
rect 3789 784 3795 796
rect 3949 764 3955 776
rect 3997 764 4003 776
rect 3933 744 3939 756
rect 3748 737 3779 743
rect 3581 704 3587 716
rect 3597 704 3603 736
rect 3540 677 3548 683
rect 3437 584 3443 636
rect 3469 624 3475 636
rect 3485 584 3491 676
rect 3629 664 3635 696
rect 3677 663 3683 716
rect 3837 704 3843 716
rect 3725 697 3740 703
rect 3693 684 3699 696
rect 3725 664 3731 697
rect 3748 697 3772 703
rect 3789 697 3820 703
rect 3789 684 3795 697
rect 3901 697 3971 703
rect 3901 683 3907 697
rect 3844 677 3907 683
rect 3677 657 3715 663
rect 3517 624 3523 636
rect 3597 564 3603 656
rect 3709 624 3715 657
rect 3677 564 3683 616
rect 3693 584 3699 596
rect 3652 557 3667 563
rect 3325 537 3347 543
rect 3309 524 3315 536
rect 3213 504 3219 516
rect 3149 444 3155 496
rect 3165 464 3171 476
rect 3165 444 3171 456
rect 3165 424 3171 436
rect 3076 277 3084 283
rect 3149 264 3155 416
rect 3325 404 3331 516
rect 3165 284 3171 316
rect 3197 304 3203 356
rect 3245 304 3251 396
rect 3309 303 3315 376
rect 3309 297 3331 303
rect 3204 277 3212 283
rect 3268 277 3315 283
rect 3245 264 3251 276
rect 3069 244 3075 256
rect 3309 243 3315 277
rect 3325 264 3331 297
rect 3341 283 3347 537
rect 3357 524 3363 556
rect 3405 544 3411 556
rect 3581 544 3587 556
rect 3613 543 3619 556
rect 3597 537 3619 543
rect 3389 523 3395 536
rect 3597 523 3603 537
rect 3645 524 3651 536
rect 3661 524 3667 557
rect 3741 544 3747 676
rect 3821 664 3827 676
rect 3853 657 3868 663
rect 3853 644 3859 657
rect 3757 624 3763 636
rect 3821 564 3827 636
rect 3700 537 3724 543
rect 3741 524 3747 536
rect 3773 524 3779 556
rect 3389 517 3603 523
rect 3373 504 3379 516
rect 3549 484 3555 496
rect 3357 324 3363 396
rect 3373 384 3379 396
rect 3373 364 3379 376
rect 3373 344 3379 356
rect 3613 324 3619 376
rect 3460 317 3468 323
rect 3373 304 3379 316
rect 3341 277 3452 283
rect 3501 264 3507 276
rect 3517 264 3523 296
rect 3613 284 3619 296
rect 3357 257 3372 263
rect 3357 243 3363 257
rect 3309 237 3363 243
rect 3277 204 3283 236
rect 3421 224 3427 236
rect 3188 177 3196 183
rect 3293 183 3299 196
rect 3485 184 3491 196
rect 3284 177 3299 183
rect 2925 123 2931 136
rect 3005 124 3011 136
rect 3021 124 3027 136
rect 3149 124 3155 176
rect 3437 164 3443 176
rect 3501 144 3507 256
rect 3556 137 3564 143
rect 3588 137 3596 143
rect 2925 117 2956 123
rect 2868 77 2908 83
rect 2973 64 2979 96
rect 2813 24 2819 36
rect 2973 -43 2979 56
rect 3005 -43 3011 116
rect 3101 84 3107 96
rect 3053 -43 3059 76
rect 3117 -37 3123 116
rect 3165 84 3171 136
rect 3197 104 3203 136
rect 3293 124 3299 136
rect 3629 124 3635 516
rect 3837 444 3843 556
rect 3869 524 3875 636
rect 3901 624 3907 636
rect 3933 584 3939 676
rect 3965 663 3971 697
rect 3981 684 3987 716
rect 3997 677 4012 683
rect 3997 663 4003 677
rect 4029 664 4035 816
rect 4045 804 4051 916
rect 4061 864 4067 1036
rect 4109 1024 4115 1076
rect 4157 1064 4163 1236
rect 4205 1164 4211 1196
rect 4237 1143 4243 1216
rect 4253 1184 4259 1296
rect 4269 1283 4275 1316
rect 4301 1304 4307 1316
rect 4317 1304 4323 1336
rect 4397 1324 4403 1336
rect 4541 1324 4547 1336
rect 4445 1304 4451 1316
rect 4349 1284 4355 1296
rect 4269 1277 4291 1283
rect 4285 1263 4291 1277
rect 4317 1263 4323 1276
rect 4285 1257 4323 1263
rect 4205 1137 4243 1143
rect 4205 1123 4211 1137
rect 4189 1117 4211 1123
rect 4189 1103 4195 1117
rect 4221 1104 4227 1116
rect 4317 1104 4323 1116
rect 4173 1097 4195 1103
rect 4173 1084 4179 1097
rect 4253 1064 4259 1096
rect 4173 1024 4179 1056
rect 4125 984 4131 1016
rect 4141 964 4147 976
rect 4093 924 4099 956
rect 4157 944 4163 976
rect 4173 964 4179 1016
rect 4301 1004 4307 1036
rect 4205 964 4211 996
rect 4285 984 4291 996
rect 4333 984 4339 1236
rect 4349 1124 4355 1236
rect 4445 1164 4451 1236
rect 4509 1184 4515 1276
rect 4525 1224 4531 1236
rect 4589 1144 4595 1336
rect 4644 1317 4652 1323
rect 4717 1304 4723 1316
rect 4765 1304 4771 1316
rect 4500 1137 4515 1143
rect 4397 1124 4403 1136
rect 4349 1064 4355 1116
rect 4404 1097 4412 1103
rect 4365 1084 4371 1096
rect 4445 1064 4451 1076
rect 4461 1064 4467 1136
rect 4509 1123 4515 1137
rect 4509 1117 4556 1123
rect 4349 984 4355 1056
rect 4397 1024 4403 1036
rect 4509 1024 4515 1056
rect 4541 1044 4547 1096
rect 4269 944 4275 976
rect 4397 964 4403 1016
rect 4573 1004 4579 1036
rect 4461 964 4467 976
rect 4589 944 4595 1016
rect 4605 944 4611 1036
rect 4621 1024 4627 1296
rect 4669 1204 4675 1296
rect 4781 1284 4787 1336
rect 4925 1284 4931 1296
rect 4957 1264 4963 1336
rect 4653 1104 4659 1116
rect 4701 1084 4707 1116
rect 4797 1104 4803 1116
rect 4813 1083 4819 1236
rect 4925 1104 4931 1116
rect 4804 1077 4819 1083
rect 4685 1064 4691 1076
rect 4701 984 4707 1036
rect 4669 964 4675 976
rect 4717 944 4723 996
rect 4749 984 4755 1076
rect 4829 1064 4835 1076
rect 4973 1064 4979 1336
rect 5005 1324 5011 1336
rect 5053 1324 5059 1537
rect 5101 1537 5123 1543
rect 5076 1477 5084 1483
rect 5069 1444 5075 1456
rect 5005 1124 5011 1136
rect 5021 1064 5027 1076
rect 4852 1057 4860 1063
rect 4893 1044 4899 1056
rect 4765 984 4771 996
rect 4733 944 4739 976
rect 4813 944 4819 1036
rect 4829 984 4835 1016
rect 4877 944 4883 1016
rect 4909 964 4915 976
rect 4324 937 4348 943
rect 4404 937 4412 943
rect 4516 937 4524 943
rect 4205 924 4211 936
rect 4493 924 4499 936
rect 4925 924 4931 1056
rect 4957 1024 4963 1036
rect 5053 1024 5059 1316
rect 5069 1104 5075 1116
rect 5044 977 5052 983
rect 5021 944 5027 956
rect 4221 917 4252 923
rect 4077 823 4083 916
rect 4173 903 4179 916
rect 4221 903 4227 917
rect 4276 917 4348 923
rect 4413 917 4444 923
rect 4173 897 4227 903
rect 4413 903 4419 917
rect 4509 917 4563 923
rect 4324 897 4419 903
rect 4301 877 4348 883
rect 4301 844 4307 877
rect 4061 817 4083 823
rect 4061 743 4067 817
rect 4077 744 4083 756
rect 4045 737 4067 743
rect 3965 657 4003 663
rect 4029 644 4035 656
rect 3885 544 3891 576
rect 3965 544 3971 596
rect 3981 523 3987 536
rect 3940 517 3987 523
rect 3869 504 3875 516
rect 3885 484 3891 496
rect 3997 483 4003 616
rect 4013 584 4019 616
rect 4029 563 4035 596
rect 4045 584 4051 737
rect 4061 704 4067 716
rect 4077 704 4083 716
rect 4093 683 4099 756
rect 4205 743 4211 836
rect 4317 744 4323 836
rect 4189 737 4211 743
rect 4157 684 4163 716
rect 4173 704 4179 716
rect 4077 677 4099 683
rect 4077 644 4083 677
rect 4093 657 4108 663
rect 4093 624 4099 657
rect 4013 557 4035 563
rect 4013 504 4019 557
rect 4029 504 4035 536
rect 4109 524 4115 636
rect 4141 624 4147 636
rect 4125 584 4131 616
rect 4173 564 4179 596
rect 4157 544 4163 556
rect 4189 543 4195 737
rect 4221 724 4227 736
rect 4285 724 4291 736
rect 4205 704 4211 716
rect 4260 697 4268 703
rect 4205 624 4211 636
rect 4221 604 4227 636
rect 4253 604 4259 676
rect 4301 644 4307 656
rect 4317 604 4323 676
rect 4333 604 4339 836
rect 4349 704 4355 716
rect 4365 684 4371 856
rect 4445 844 4451 896
rect 4509 884 4515 917
rect 4557 904 4563 917
rect 4749 917 4787 923
rect 4573 897 4668 903
rect 4573 883 4579 897
rect 4749 884 4755 917
rect 4781 904 4787 917
rect 4877 904 4883 916
rect 4909 904 4915 916
rect 5021 904 5027 916
rect 4788 897 4812 903
rect 4765 884 4771 896
rect 4532 877 4579 883
rect 4429 784 4435 836
rect 4493 724 4499 736
rect 4637 724 4643 736
rect 4653 704 4659 716
rect 4404 697 4412 703
rect 4500 697 4508 703
rect 4381 683 4387 696
rect 4605 684 4611 696
rect 4701 684 4707 816
rect 5021 784 5027 876
rect 4733 724 4739 736
rect 5037 724 5043 736
rect 4957 704 4963 716
rect 5053 704 5059 816
rect 5085 704 5091 1336
rect 5101 1324 5107 1537
rect 5133 1284 5139 1476
rect 5165 1464 5171 1556
rect 5149 1344 5155 1356
rect 5165 1304 5171 1336
rect 5101 1063 5107 1176
rect 5117 1164 5123 1276
rect 5133 1084 5139 1236
rect 5101 1057 5123 1063
rect 5101 944 5107 1036
rect 5117 963 5123 1057
rect 5117 957 5139 963
rect 5117 924 5123 936
rect 5133 924 5139 957
rect 5165 943 5171 1276
rect 5181 1124 5187 1797
rect 5197 1344 5203 1876
rect 5197 1304 5203 1316
rect 5149 937 5171 943
rect 5133 744 5139 756
rect 5149 744 5155 937
rect 5181 883 5187 1056
rect 5197 1024 5203 1036
rect 5181 877 5203 883
rect 5172 777 5180 783
rect 4788 697 4796 703
rect 4909 684 4915 696
rect 5037 684 5043 696
rect 4381 677 4396 683
rect 4413 677 4444 683
rect 4413 664 4419 677
rect 4829 664 4835 676
rect 4925 664 4931 676
rect 4532 657 4540 663
rect 4788 657 4796 663
rect 4445 644 4451 656
rect 4493 604 4499 636
rect 4205 564 4211 596
rect 4269 584 4275 596
rect 4253 564 4259 576
rect 4317 564 4323 576
rect 4532 557 4540 563
rect 4333 544 4339 556
rect 4189 537 4211 543
rect 4116 497 4124 503
rect 4045 483 4051 496
rect 3997 477 4051 483
rect 3917 464 3923 476
rect 3645 324 3651 336
rect 3677 297 3692 303
rect 3661 264 3667 276
rect 3677 224 3683 297
rect 3741 284 3747 356
rect 3693 224 3699 236
rect 3725 164 3731 236
rect 3741 224 3747 256
rect 3773 224 3779 336
rect 3796 317 3804 323
rect 3821 304 3827 316
rect 3789 224 3795 236
rect 3805 224 3811 276
rect 3869 264 3875 296
rect 3885 284 3891 336
rect 3933 284 3939 296
rect 3981 264 3987 436
rect 4004 337 4012 343
rect 4061 304 4067 396
rect 4116 317 4124 323
rect 4077 304 4083 316
rect 3853 164 3859 236
rect 3901 224 3907 236
rect 4013 204 4019 296
rect 4157 284 4163 496
rect 4180 377 4188 383
rect 4205 324 4211 537
rect 4237 524 4243 536
rect 4285 524 4291 536
rect 4365 504 4371 536
rect 4461 524 4467 536
rect 4477 464 4483 556
rect 4509 484 4515 536
rect 4557 524 4563 536
rect 4573 523 4579 636
rect 4605 544 4611 596
rect 4621 544 4627 636
rect 4973 624 4979 656
rect 4733 584 4739 596
rect 4653 564 4659 576
rect 4692 537 4700 543
rect 4573 517 4595 523
rect 4237 344 4243 436
rect 4253 324 4259 436
rect 4301 404 4307 436
rect 4397 404 4403 436
rect 4333 323 4339 376
rect 4308 317 4339 323
rect 4429 304 4435 336
rect 4212 277 4243 283
rect 4036 257 4060 263
rect 4237 263 4243 277
rect 4260 277 4291 283
rect 4237 257 4268 263
rect 4045 224 4051 236
rect 4109 204 4115 256
rect 3965 164 3971 176
rect 4045 164 4051 196
rect 4093 184 4099 196
rect 3757 157 3772 163
rect 3757 144 3763 157
rect 4077 163 4083 176
rect 4125 164 4131 236
rect 4141 184 4147 196
rect 4077 157 4099 163
rect 3789 144 3795 156
rect 3773 124 3779 136
rect 4093 123 4099 157
rect 4173 163 4179 196
rect 4141 157 4179 163
rect 4109 144 4115 156
rect 4141 123 4147 157
rect 4164 137 4172 143
rect 4093 117 4147 123
rect 3389 104 3395 116
rect 3565 104 3571 116
rect 3332 97 3340 103
rect 3197 84 3203 96
rect 3501 64 3507 76
rect 3117 -43 3139 -37
rect 3725 -43 3731 116
rect 3949 104 3955 116
rect 4189 104 4195 216
rect 4221 204 4227 236
rect 4253 123 4259 196
rect 4285 184 4291 277
rect 4365 264 4371 276
rect 4461 264 4467 416
rect 4573 344 4579 496
rect 4589 484 4595 517
rect 4621 444 4627 496
rect 4637 484 4643 496
rect 4653 324 4659 536
rect 4733 384 4739 416
rect 4765 404 4771 556
rect 4797 524 4803 596
rect 4893 584 4899 596
rect 4829 544 4835 576
rect 4845 564 4851 576
rect 4925 564 4931 596
rect 5005 564 5011 656
rect 5037 564 5043 596
rect 5053 584 5059 696
rect 5092 677 5100 683
rect 5085 644 5091 656
rect 5069 564 5075 616
rect 5117 604 5123 636
rect 5133 564 5139 596
rect 5197 564 5203 877
rect 5213 624 5219 1316
rect 4877 544 4883 556
rect 4813 524 4819 536
rect 4957 524 4963 536
rect 4973 524 4979 556
rect 5117 544 5123 556
rect 4829 344 4835 496
rect 4557 304 4563 316
rect 4621 284 4627 296
rect 4701 284 4707 296
rect 4717 284 4723 316
rect 4861 304 4867 436
rect 4925 403 4931 516
rect 4925 397 4947 403
rect 4765 277 4780 283
rect 4653 264 4659 276
rect 4749 264 4755 276
rect 4765 264 4771 277
rect 4461 244 4467 256
rect 4333 164 4339 196
rect 4397 183 4403 236
rect 4413 184 4419 196
rect 4509 184 4515 256
rect 4381 177 4403 183
rect 4269 157 4323 163
rect 4269 144 4275 157
rect 4317 144 4323 157
rect 4381 144 4387 177
rect 4445 164 4451 176
rect 4516 157 4524 163
rect 4397 144 4403 156
rect 4429 144 4435 156
rect 4477 144 4483 156
rect 4557 144 4563 256
rect 4797 244 4803 296
rect 4829 264 4835 276
rect 4941 264 4947 397
rect 4973 344 4979 436
rect 4884 257 4892 263
rect 4973 244 4979 256
rect 4669 224 4675 236
rect 4813 224 4819 236
rect 4253 117 4268 123
rect 4285 104 4291 136
rect 4669 124 4675 196
rect 4781 164 4787 216
rect 4861 164 4867 196
rect 4877 184 4883 196
rect 4820 157 4828 163
rect 4996 157 5004 163
rect 4685 144 4691 156
rect 4973 144 4979 156
rect 5021 144 5027 236
rect 5037 183 5043 476
rect 5101 344 5107 436
rect 5117 384 5123 516
rect 5165 504 5171 516
rect 5165 384 5171 416
rect 5133 284 5139 296
rect 5149 284 5155 356
rect 5181 324 5187 336
rect 5060 257 5068 263
rect 5037 177 5059 183
rect 5053 164 5059 177
rect 5085 164 5091 236
rect 5181 164 5187 176
rect 5156 157 5164 163
rect 5069 144 5075 156
rect 5133 144 5139 156
rect 4813 124 4819 136
rect 4788 117 4796 123
rect 4941 104 4947 136
rect 4061 84 4067 96
rect 4237 84 4243 96
rect 4397 84 4403 96
rect 3805 -43 3811 36
rect 5021 -37 5027 36
rect 5101 -37 5107 116
rect 5005 -43 5027 -37
rect 5085 -43 5107 -37
<< m3contact >>
rect 604 3576 612 3584
rect 700 3556 708 3564
rect 764 3556 772 3564
rect 316 3536 324 3544
rect 428 3536 436 3544
rect 476 3536 484 3544
rect 556 3536 564 3544
rect 332 3516 340 3524
rect 60 3496 68 3504
rect 12 3376 20 3384
rect 12 3356 20 3364
rect 44 3356 52 3364
rect 60 3356 68 3364
rect 156 3476 164 3484
rect 236 3476 244 3484
rect 348 3476 356 3484
rect 380 3476 388 3484
rect 412 3476 420 3484
rect 476 3476 484 3484
rect 508 3476 516 3484
rect 668 3476 676 3484
rect 716 3476 724 3484
rect 748 3476 756 3484
rect 140 3456 148 3464
rect 236 3456 244 3464
rect 268 3456 276 3464
rect 124 3436 132 3444
rect 156 3376 164 3384
rect 108 3356 116 3364
rect 92 3336 100 3344
rect 140 3316 148 3324
rect 92 3296 100 3304
rect 108 3296 116 3304
rect 156 3276 164 3284
rect 284 3436 292 3444
rect 364 3436 372 3444
rect 220 3376 228 3384
rect 348 3376 356 3384
rect 460 3436 468 3444
rect 204 3356 212 3364
rect 300 3356 308 3364
rect 476 3356 484 3364
rect 284 3336 292 3344
rect 396 3336 404 3344
rect 236 3296 244 3304
rect 188 3216 196 3224
rect 60 3116 68 3124
rect 172 3116 180 3124
rect 12 3096 20 3104
rect 44 3096 52 3104
rect 156 3096 164 3104
rect 188 3096 196 3104
rect 172 3076 180 3084
rect 220 3216 228 3224
rect 348 3296 356 3304
rect 396 3296 404 3304
rect 332 3216 340 3224
rect 300 3096 308 3104
rect 364 3096 372 3104
rect 220 3076 228 3084
rect 268 3076 276 3084
rect 316 3076 324 3084
rect 348 3076 356 3084
rect 396 3096 404 3104
rect 396 3076 404 3084
rect 76 2996 84 3004
rect 60 2956 68 2964
rect 204 3036 212 3044
rect 140 2996 148 3004
rect 284 2976 292 2984
rect 172 2956 180 2964
rect 44 2936 52 2944
rect 108 2936 116 2944
rect 140 2936 148 2944
rect 108 2916 116 2924
rect 140 2736 148 2744
rect 12 2716 20 2724
rect 60 2716 68 2724
rect 92 2716 100 2724
rect 252 2936 260 2944
rect 716 3456 724 3464
rect 572 3436 580 3444
rect 636 3436 644 3444
rect 764 3436 772 3444
rect 780 3436 788 3444
rect 716 3416 724 3424
rect 620 3396 628 3404
rect 540 3376 548 3384
rect 572 3376 580 3384
rect 636 3376 644 3384
rect 732 3376 740 3384
rect 828 3596 836 3604
rect 1180 3596 1188 3604
rect 2300 3616 2308 3624
rect 3260 3616 3268 3624
rect 3388 3616 3396 3624
rect 3644 3596 3652 3604
rect 4028 3596 4036 3604
rect 1068 3576 1076 3584
rect 972 3556 980 3564
rect 1452 3556 1460 3564
rect 1916 3556 1924 3564
rect 2060 3556 2068 3564
rect 2748 3556 2756 3564
rect 1004 3536 1012 3544
rect 1356 3516 1364 3524
rect 1404 3516 1412 3524
rect 1148 3496 1156 3504
rect 1212 3496 1220 3504
rect 1244 3496 1252 3504
rect 1260 3496 1268 3504
rect 1308 3496 1316 3504
rect 828 3456 836 3464
rect 844 3456 852 3464
rect 812 3436 820 3444
rect 924 3456 932 3464
rect 972 3456 980 3464
rect 1020 3436 1028 3444
rect 1036 3416 1044 3424
rect 956 3396 964 3404
rect 1100 3436 1108 3444
rect 1084 3416 1092 3424
rect 1116 3396 1124 3404
rect 1804 3516 1812 3524
rect 1436 3496 1444 3504
rect 1340 3476 1348 3484
rect 1388 3476 1396 3484
rect 1404 3476 1412 3484
rect 1452 3476 1460 3484
rect 1484 3476 1492 3484
rect 1196 3456 1204 3464
rect 1164 3436 1172 3444
rect 1244 3436 1252 3444
rect 1228 3416 1236 3424
rect 1148 3396 1156 3404
rect 1292 3396 1300 3404
rect 1420 3416 1428 3424
rect 1500 3416 1508 3424
rect 2380 3536 2388 3544
rect 2460 3536 2468 3544
rect 2524 3536 2532 3544
rect 1948 3516 1956 3524
rect 2012 3516 2020 3524
rect 2108 3516 2116 3524
rect 2172 3516 2180 3524
rect 2332 3516 2340 3524
rect 1724 3476 1732 3484
rect 1628 3456 1636 3464
rect 1708 3456 1716 3464
rect 1484 3376 1492 3384
rect 1516 3376 1524 3384
rect 1676 3436 1684 3444
rect 1724 3436 1732 3444
rect 1644 3416 1652 3424
rect 540 3356 548 3364
rect 972 3356 980 3364
rect 1036 3356 1044 3364
rect 1116 3356 1124 3364
rect 1292 3356 1300 3364
rect 1324 3356 1332 3364
rect 1388 3356 1396 3364
rect 1468 3356 1476 3364
rect 1564 3356 1572 3364
rect 1612 3356 1620 3364
rect 572 3336 580 3344
rect 636 3336 644 3344
rect 700 3336 708 3344
rect 716 3336 724 3344
rect 764 3336 772 3344
rect 796 3336 804 3344
rect 812 3336 820 3344
rect 844 3336 852 3344
rect 1020 3336 1028 3344
rect 1116 3336 1124 3344
rect 1164 3336 1172 3344
rect 1228 3336 1236 3344
rect 1260 3336 1268 3344
rect 1276 3336 1284 3344
rect 684 3296 692 3304
rect 444 3276 452 3284
rect 492 3276 500 3284
rect 524 3276 532 3284
rect 780 3236 788 3244
rect 460 3196 468 3204
rect 1852 3476 1860 3484
rect 2412 3516 2420 3524
rect 2668 3516 2676 3524
rect 2716 3516 2724 3524
rect 2044 3456 2052 3464
rect 1916 3436 1924 3444
rect 2076 3436 2084 3444
rect 2556 3456 2564 3464
rect 2572 3456 2580 3464
rect 2844 3536 2852 3544
rect 2892 3536 2900 3544
rect 2780 3516 2788 3524
rect 2908 3516 2916 3524
rect 2924 3516 2932 3524
rect 2764 3476 2772 3484
rect 1772 3416 1780 3424
rect 1980 3416 1988 3424
rect 1916 3396 1924 3404
rect 1740 3356 1748 3364
rect 1772 3356 1780 3364
rect 1596 3336 1604 3344
rect 1788 3336 1796 3344
rect 1820 3336 1828 3344
rect 1868 3336 1876 3344
rect 908 3296 916 3304
rect 1068 3296 1076 3304
rect 1132 3296 1140 3304
rect 844 3256 852 3264
rect 508 3156 516 3164
rect 700 3156 708 3164
rect 460 3076 468 3084
rect 588 3076 596 3084
rect 604 3076 612 3084
rect 556 3036 564 3044
rect 604 3036 612 3044
rect 540 3016 548 3024
rect 572 3016 580 3024
rect 652 3016 660 3024
rect 668 3016 676 3024
rect 508 2996 516 3004
rect 732 3096 740 3104
rect 780 3096 788 3104
rect 1180 3276 1188 3284
rect 1228 3276 1236 3284
rect 1372 3276 1380 3284
rect 1196 3236 1204 3244
rect 988 3216 996 3224
rect 1340 3196 1348 3204
rect 1324 3176 1332 3184
rect 956 3156 964 3164
rect 1084 3136 1092 3144
rect 1308 3136 1316 3144
rect 892 3116 900 3124
rect 876 3096 884 3104
rect 908 3096 916 3104
rect 988 3096 996 3104
rect 1068 3096 1076 3104
rect 1100 3096 1108 3104
rect 1148 3096 1156 3104
rect 1292 3096 1300 3104
rect 732 3076 740 3084
rect 780 3076 788 3084
rect 828 3076 836 3084
rect 940 3076 948 3084
rect 1020 3076 1028 3084
rect 1164 3076 1172 3084
rect 1196 3076 1204 3084
rect 1260 3076 1268 3084
rect 828 3056 836 3064
rect 716 3036 724 3044
rect 812 3036 820 3044
rect 972 3036 980 3044
rect 396 2976 404 2984
rect 524 2976 532 2984
rect 556 2976 564 2984
rect 668 2976 676 2984
rect 316 2956 324 2964
rect 444 2956 452 2964
rect 476 2956 484 2964
rect 236 2916 244 2924
rect 300 2916 308 2924
rect 284 2876 292 2884
rect 236 2716 244 2724
rect 556 2936 564 2944
rect 652 2936 660 2944
rect 684 2936 692 2944
rect 700 2936 708 2944
rect 348 2916 356 2924
rect 396 2896 404 2904
rect 428 2896 436 2904
rect 476 2896 484 2904
rect 508 2876 516 2884
rect 380 2856 388 2864
rect 460 2816 468 2824
rect 396 2796 404 2804
rect 332 2756 340 2764
rect 892 2996 900 3004
rect 764 2976 772 2984
rect 844 2976 852 2984
rect 700 2916 708 2924
rect 716 2916 724 2924
rect 764 2916 772 2924
rect 604 2896 612 2904
rect 668 2896 676 2904
rect 716 2856 724 2864
rect 572 2776 580 2784
rect 508 2736 516 2744
rect 12 2696 20 2704
rect 108 2676 116 2684
rect 12 2516 20 2524
rect 156 2656 164 2664
rect 204 2656 212 2664
rect 236 2656 244 2664
rect 300 2656 308 2664
rect 348 2656 356 2664
rect 412 2656 420 2664
rect 444 2656 452 2664
rect 188 2636 196 2644
rect 220 2616 228 2624
rect 76 2596 84 2604
rect 92 2596 100 2604
rect 124 2596 132 2604
rect 508 2676 516 2684
rect 524 2676 532 2684
rect 556 2676 564 2684
rect 380 2636 388 2644
rect 396 2636 404 2644
rect 476 2636 484 2644
rect 572 2636 580 2644
rect 252 2596 260 2604
rect 268 2596 276 2604
rect 332 2596 340 2604
rect 140 2576 148 2584
rect 236 2576 244 2584
rect 108 2536 116 2544
rect 156 2516 164 2524
rect 364 2576 372 2584
rect 204 2496 212 2504
rect 236 2496 244 2504
rect 12 2316 20 2324
rect 140 2476 148 2484
rect 92 2396 100 2404
rect 316 2516 324 2524
rect 572 2596 580 2604
rect 620 2596 628 2604
rect 460 2576 468 2584
rect 508 2576 516 2584
rect 556 2576 564 2584
rect 428 2496 436 2504
rect 380 2456 388 2464
rect 284 2396 292 2404
rect 364 2376 372 2384
rect 476 2496 484 2504
rect 652 2816 660 2824
rect 684 2796 692 2804
rect 956 2996 964 3004
rect 1004 2996 1012 3004
rect 1372 3176 1380 3184
rect 1436 3176 1444 3184
rect 1356 3116 1364 3124
rect 1388 3116 1396 3124
rect 1404 3116 1412 3124
rect 1596 3276 1604 3284
rect 1660 3276 1668 3284
rect 1692 3276 1700 3284
rect 1740 3276 1748 3284
rect 1564 3256 1572 3264
rect 1596 3236 1604 3244
rect 1516 3216 1524 3224
rect 1484 3116 1492 3124
rect 1500 3116 1508 3124
rect 1068 3036 1076 3044
rect 1116 3036 1124 3044
rect 1036 2996 1044 3004
rect 1084 2996 1092 3004
rect 1196 3016 1204 3024
rect 1276 3016 1284 3024
rect 1164 2996 1172 3004
rect 1148 2976 1156 2984
rect 956 2956 964 2964
rect 988 2956 996 2964
rect 1228 2976 1236 2984
rect 1468 2996 1476 3004
rect 1324 2976 1332 2984
rect 1372 2976 1380 2984
rect 1420 2976 1428 2984
rect 1436 2976 1444 2984
rect 1468 2976 1476 2984
rect 812 2916 820 2924
rect 828 2916 836 2924
rect 796 2896 804 2904
rect 812 2896 820 2904
rect 860 2896 868 2904
rect 876 2896 884 2904
rect 988 2896 996 2904
rect 1068 2896 1076 2904
rect 1132 2896 1140 2904
rect 1180 2896 1188 2904
rect 1260 2896 1268 2904
rect 1420 2896 1428 2904
rect 956 2876 964 2884
rect 1244 2876 1252 2884
rect 1292 2876 1300 2884
rect 1340 2876 1348 2884
rect 1404 2876 1412 2884
rect 780 2856 788 2864
rect 1180 2836 1188 2844
rect 924 2776 932 2784
rect 716 2716 724 2724
rect 908 2716 916 2724
rect 700 2676 708 2684
rect 812 2676 820 2684
rect 652 2656 660 2664
rect 796 2656 804 2664
rect 844 2656 852 2664
rect 876 2656 884 2664
rect 700 2636 708 2644
rect 748 2596 756 2604
rect 684 2576 692 2584
rect 716 2576 724 2584
rect 732 2576 740 2584
rect 540 2516 548 2524
rect 508 2496 516 2504
rect 556 2416 564 2424
rect 620 2436 628 2444
rect 620 2416 628 2424
rect 716 2516 724 2524
rect 748 2516 756 2524
rect 780 2516 788 2524
rect 588 2396 596 2404
rect 636 2396 644 2404
rect 572 2336 580 2344
rect 620 2336 628 2344
rect 300 2316 308 2324
rect 348 2316 356 2324
rect 460 2316 468 2324
rect 60 2296 68 2304
rect 412 2296 420 2304
rect 428 2296 436 2304
rect 508 2296 516 2304
rect 572 2296 580 2304
rect 44 2276 52 2284
rect 28 2256 36 2264
rect 60 2256 68 2264
rect 140 2256 148 2264
rect 188 2256 196 2264
rect 60 2176 68 2184
rect 172 2176 180 2184
rect 268 2196 276 2204
rect 236 2176 244 2184
rect 300 2256 308 2264
rect 348 2256 356 2264
rect 332 2236 340 2244
rect 444 2256 452 2264
rect 844 2576 852 2584
rect 828 2536 836 2544
rect 988 2716 996 2724
rect 1276 2856 1284 2864
rect 1260 2816 1268 2824
rect 1324 2816 1332 2824
rect 1388 2816 1396 2824
rect 1052 2736 1060 2744
rect 1084 2716 1092 2724
rect 1276 2716 1284 2724
rect 1324 2716 1332 2724
rect 1356 2716 1364 2724
rect 1196 2696 1204 2704
rect 940 2676 948 2684
rect 1004 2676 1012 2684
rect 1036 2676 1044 2684
rect 1100 2676 1108 2684
rect 1116 2676 1124 2684
rect 988 2636 996 2644
rect 1148 2676 1156 2684
rect 1228 2676 1236 2684
rect 1260 2676 1268 2684
rect 1132 2656 1140 2664
rect 1148 2656 1156 2664
rect 1308 2656 1316 2664
rect 956 2596 964 2604
rect 956 2576 964 2584
rect 1004 2616 1012 2624
rect 924 2536 932 2544
rect 1116 2576 1124 2584
rect 1164 2536 1172 2544
rect 828 2516 836 2524
rect 1036 2516 1044 2524
rect 1020 2496 1028 2504
rect 1036 2496 1044 2504
rect 1068 2496 1076 2504
rect 1132 2496 1140 2504
rect 860 2476 868 2484
rect 876 2476 884 2484
rect 956 2476 964 2484
rect 796 2416 804 2424
rect 812 2396 820 2404
rect 764 2336 772 2344
rect 700 2316 708 2324
rect 780 2296 788 2304
rect 684 2276 692 2284
rect 796 2276 804 2284
rect 524 2256 532 2264
rect 540 2256 548 2264
rect 652 2256 660 2264
rect 668 2256 676 2264
rect 476 2236 484 2244
rect 508 2236 516 2244
rect 380 2216 388 2224
rect 348 2176 356 2184
rect 188 2156 196 2164
rect 220 2156 228 2164
rect 380 2156 388 2164
rect 12 2136 20 2144
rect 44 2136 52 2144
rect 92 2136 100 2144
rect 92 2116 100 2124
rect 44 1876 52 1884
rect 12 1836 20 1844
rect 60 1836 68 1844
rect 76 1816 84 1824
rect 316 2136 324 2144
rect 332 2116 340 2124
rect 364 2116 372 2124
rect 140 1916 148 1924
rect 188 1916 196 1924
rect 284 2096 292 2104
rect 380 2056 388 2064
rect 188 1896 196 1904
rect 188 1856 196 1864
rect 124 1796 132 1804
rect 172 1796 180 1804
rect 220 1776 228 1784
rect 140 1756 148 1764
rect 220 1756 228 1764
rect 204 1736 212 1744
rect 60 1716 68 1724
rect 108 1716 116 1724
rect 460 2156 468 2164
rect 604 2236 612 2244
rect 556 2216 564 2224
rect 668 2236 676 2244
rect 668 2216 676 2224
rect 636 2196 644 2204
rect 748 2196 756 2204
rect 684 2176 692 2184
rect 700 2176 708 2184
rect 620 2156 628 2164
rect 412 2116 420 2124
rect 444 2116 452 2124
rect 508 2116 516 2124
rect 412 1996 420 2004
rect 476 2096 484 2104
rect 460 2076 468 2084
rect 364 1916 372 1924
rect 396 1916 404 1924
rect 380 1896 388 1904
rect 428 1896 436 1904
rect 348 1876 356 1884
rect 316 1856 324 1864
rect 364 1856 372 1864
rect 268 1836 276 1844
rect 332 1836 340 1844
rect 236 1736 244 1744
rect 252 1736 260 1744
rect 268 1716 276 1724
rect 284 1696 292 1704
rect 300 1676 308 1684
rect 92 1616 100 1624
rect 124 1616 132 1624
rect 92 1516 100 1524
rect 108 1516 116 1524
rect 60 1496 68 1504
rect 12 1476 20 1484
rect 12 1376 20 1384
rect 44 1356 52 1364
rect 108 1376 116 1384
rect 92 1356 100 1364
rect 12 1336 20 1344
rect 76 1336 84 1344
rect 92 1316 100 1324
rect 44 1296 52 1304
rect 28 1156 36 1164
rect 188 1516 196 1524
rect 236 1556 244 1564
rect 284 1536 292 1544
rect 252 1516 260 1524
rect 204 1496 212 1504
rect 236 1496 244 1504
rect 204 1476 212 1484
rect 156 1456 164 1464
rect 220 1456 228 1464
rect 140 1336 148 1344
rect 188 1336 196 1344
rect 124 1316 132 1324
rect 156 1316 164 1324
rect 140 1236 148 1244
rect 108 1156 116 1164
rect 300 1456 308 1464
rect 412 1836 420 1844
rect 380 1796 388 1804
rect 396 1776 404 1784
rect 844 2316 852 2324
rect 860 2296 868 2304
rect 908 2296 916 2304
rect 908 2276 916 2284
rect 844 2256 852 2264
rect 828 2236 836 2244
rect 844 2176 852 2184
rect 796 2156 804 2164
rect 556 2056 564 2064
rect 492 1956 500 1964
rect 492 1936 500 1944
rect 588 2096 596 2104
rect 652 2056 660 2064
rect 732 2096 740 2104
rect 748 2096 756 2104
rect 748 2056 756 2064
rect 812 2016 820 2024
rect 860 2056 868 2064
rect 844 1996 852 2004
rect 796 1976 804 1984
rect 844 1976 852 1984
rect 732 1936 740 1944
rect 556 1916 564 1924
rect 636 1916 644 1924
rect 684 1916 692 1924
rect 540 1896 548 1904
rect 588 1896 596 1904
rect 652 1896 660 1904
rect 780 1896 788 1904
rect 828 1896 836 1904
rect 860 1896 868 1904
rect 604 1876 612 1884
rect 636 1876 644 1884
rect 684 1876 692 1884
rect 1004 2416 1012 2424
rect 1020 2336 1028 2344
rect 1036 2316 1044 2324
rect 1164 2316 1172 2324
rect 1052 2296 1060 2304
rect 1100 2296 1108 2304
rect 988 2276 996 2284
rect 1020 2276 1028 2284
rect 956 2216 964 2224
rect 940 2196 948 2204
rect 892 2176 900 2184
rect 972 2196 980 2204
rect 1100 2216 1108 2224
rect 1164 2216 1172 2224
rect 940 2156 948 2164
rect 1116 2156 1124 2164
rect 1132 2156 1140 2164
rect 1356 2636 1364 2644
rect 1308 2616 1316 2624
rect 1324 2616 1332 2624
rect 1260 2576 1268 2584
rect 1372 2596 1380 2604
rect 1196 2536 1204 2544
rect 1212 2516 1220 2524
rect 1228 2516 1236 2524
rect 1228 2316 1236 2324
rect 1212 2296 1220 2304
rect 1228 2296 1236 2304
rect 1276 2536 1284 2544
rect 1356 2556 1364 2564
rect 1468 2896 1476 2904
rect 1500 2896 1508 2904
rect 1580 3076 1588 3084
rect 1660 3116 1668 3124
rect 1676 3116 1684 3124
rect 2220 3436 2228 3444
rect 2316 3436 2324 3444
rect 2364 3436 2372 3444
rect 2412 3436 2420 3444
rect 2476 3436 2484 3444
rect 2508 3436 2516 3444
rect 2604 3436 2612 3444
rect 2700 3456 2708 3464
rect 2732 3436 2740 3444
rect 2748 3436 2756 3444
rect 2300 3416 2308 3424
rect 2236 3396 2244 3404
rect 2268 3396 2276 3404
rect 2124 3356 2132 3364
rect 2156 3356 2164 3364
rect 2316 3396 2324 3404
rect 2348 3396 2356 3404
rect 2620 3396 2628 3404
rect 2732 3396 2740 3404
rect 2396 3356 2404 3364
rect 2444 3356 2452 3364
rect 2476 3356 2484 3364
rect 2524 3356 2532 3364
rect 2572 3356 2580 3364
rect 2604 3356 2612 3364
rect 2220 3336 2228 3344
rect 2028 3276 2036 3284
rect 2108 3276 2116 3284
rect 2188 3276 2196 3284
rect 2204 3276 2212 3284
rect 1852 3236 1860 3244
rect 1900 3216 1908 3224
rect 2044 3256 2052 3264
rect 2076 3256 2084 3264
rect 2124 3256 2132 3264
rect 1980 3216 1988 3224
rect 1948 3196 1956 3204
rect 2076 3176 2084 3184
rect 2108 3116 2116 3124
rect 1772 3096 1780 3104
rect 1852 3096 1860 3104
rect 1916 3096 1924 3104
rect 1964 3096 1972 3104
rect 2012 3096 2020 3104
rect 2028 3096 2036 3104
rect 2060 3096 2068 3104
rect 2188 3096 2196 3104
rect 2268 3276 2276 3284
rect 2396 3276 2404 3284
rect 2492 3276 2500 3284
rect 2300 3256 2308 3264
rect 2700 3356 2708 3364
rect 2572 3296 2580 3304
rect 2620 3296 2628 3304
rect 2540 3276 2548 3284
rect 2508 3216 2516 3224
rect 2540 3196 2548 3204
rect 2220 3176 2228 3184
rect 2252 3176 2260 3184
rect 2236 3116 2244 3124
rect 2220 3096 2228 3104
rect 2316 3156 2324 3164
rect 2476 3116 2484 3124
rect 2332 3096 2340 3104
rect 2348 3096 2356 3104
rect 2380 3096 2388 3104
rect 2412 3096 2420 3104
rect 2300 3076 2308 3084
rect 2380 3076 2388 3084
rect 1628 3056 1636 3064
rect 1644 3056 1652 3064
rect 1548 3036 1556 3044
rect 1596 2936 1604 2944
rect 1596 2896 1604 2904
rect 1532 2876 1540 2884
rect 1596 2836 1604 2844
rect 1436 2776 1444 2784
rect 1628 2936 1636 2944
rect 1708 3016 1716 3024
rect 2204 3056 2212 3064
rect 2220 3056 2228 3064
rect 2156 3036 2164 3044
rect 1964 2996 1972 3004
rect 2028 2996 2036 3004
rect 2092 2996 2100 3004
rect 2140 2996 2148 3004
rect 1644 2896 1652 2904
rect 1676 2896 1684 2904
rect 1628 2876 1636 2884
rect 1724 2856 1732 2864
rect 1708 2836 1716 2844
rect 1612 2816 1620 2824
rect 1724 2816 1732 2824
rect 1692 2776 1700 2784
rect 1452 2716 1460 2724
rect 1516 2716 1524 2724
rect 1500 2696 1508 2704
rect 1612 2696 1620 2704
rect 1916 2936 1924 2944
rect 1932 2936 1940 2944
rect 1964 2936 1972 2944
rect 2028 2936 2036 2944
rect 2060 2936 2068 2944
rect 2092 2936 2100 2944
rect 1804 2896 1812 2904
rect 2348 3056 2356 3064
rect 2620 3096 2628 3104
rect 2636 3096 2644 3104
rect 2428 3056 2436 3064
rect 2396 3036 2404 3044
rect 2444 3036 2452 3044
rect 2460 3036 2468 3044
rect 2492 3036 2500 3044
rect 2524 3036 2532 3044
rect 2540 3036 2548 3044
rect 2588 3036 2596 3044
rect 2620 3036 2628 3044
rect 2252 2956 2260 2964
rect 2572 2996 2580 3004
rect 2636 2996 2644 3004
rect 2524 2956 2532 2964
rect 2540 2956 2548 2964
rect 2620 2956 2628 2964
rect 2444 2936 2452 2944
rect 2476 2936 2484 2944
rect 1852 2916 1860 2924
rect 1884 2916 1892 2924
rect 2076 2916 2084 2924
rect 2108 2916 2116 2924
rect 2204 2916 2212 2924
rect 2284 2916 2292 2924
rect 1836 2896 1844 2904
rect 1772 2876 1780 2884
rect 1804 2876 1812 2884
rect 1820 2876 1828 2884
rect 1868 2896 1876 2904
rect 1756 2856 1764 2864
rect 1916 2896 1924 2904
rect 2444 2896 2452 2904
rect 1916 2876 1924 2884
rect 1932 2876 1940 2884
rect 1996 2876 2004 2884
rect 2012 2876 2020 2884
rect 2060 2876 2068 2884
rect 2268 2876 2276 2884
rect 2300 2876 2308 2884
rect 2364 2876 2372 2884
rect 2428 2876 2436 2884
rect 1948 2856 1956 2864
rect 2124 2856 2132 2864
rect 1788 2816 1796 2824
rect 1820 2816 1828 2824
rect 1916 2816 1924 2824
rect 1788 2736 1796 2744
rect 1564 2636 1572 2644
rect 1644 2636 1652 2644
rect 1468 2616 1476 2624
rect 1548 2616 1556 2624
rect 1580 2616 1588 2624
rect 1628 2616 1636 2624
rect 1836 2776 1844 2784
rect 2060 2776 2068 2784
rect 1884 2736 1892 2744
rect 1996 2736 2004 2744
rect 2044 2736 2052 2744
rect 2092 2736 2100 2744
rect 1900 2716 1908 2724
rect 1948 2676 1956 2684
rect 1308 2536 1316 2544
rect 1324 2536 1332 2544
rect 1388 2536 1396 2544
rect 1436 2536 1444 2544
rect 1276 2516 1284 2524
rect 1308 2516 1316 2524
rect 1388 2496 1396 2504
rect 1420 2496 1428 2504
rect 1404 2456 1412 2464
rect 1260 2416 1268 2424
rect 1324 2396 1332 2404
rect 1500 2476 1508 2484
rect 1532 2476 1540 2484
rect 1548 2456 1556 2464
rect 1516 2416 1524 2424
rect 1644 2476 1652 2484
rect 1708 2596 1716 2604
rect 1724 2576 1732 2584
rect 1708 2496 1716 2504
rect 1692 2476 1700 2484
rect 1660 2436 1668 2444
rect 1660 2396 1668 2404
rect 1436 2376 1444 2384
rect 1276 2336 1284 2344
rect 1356 2336 1364 2344
rect 1500 2336 1508 2344
rect 1548 2336 1556 2344
rect 1644 2336 1652 2344
rect 1340 2316 1348 2324
rect 1628 2316 1636 2324
rect 1676 2316 1684 2324
rect 1772 2636 1780 2644
rect 1852 2636 1860 2644
rect 1932 2616 1940 2624
rect 1948 2616 1956 2624
rect 2060 2636 2068 2644
rect 1996 2616 2004 2624
rect 2108 2616 2116 2624
rect 2076 2596 2084 2604
rect 2092 2596 2100 2604
rect 2268 2816 2276 2824
rect 2300 2816 2308 2824
rect 2156 2736 2164 2744
rect 2316 2736 2324 2744
rect 2412 2716 2420 2724
rect 2156 2616 2164 2624
rect 2028 2576 2036 2584
rect 1804 2556 1812 2564
rect 1820 2556 1828 2564
rect 1980 2556 1988 2564
rect 2060 2556 2068 2564
rect 2076 2556 2084 2564
rect 1740 2496 1748 2504
rect 1820 2496 1828 2504
rect 1788 2476 1796 2484
rect 1836 2456 1844 2464
rect 1916 2496 1924 2504
rect 1868 2436 1876 2444
rect 1868 2396 1876 2404
rect 1980 2496 1988 2504
rect 1996 2496 2004 2504
rect 2316 2636 2324 2644
rect 2204 2616 2212 2624
rect 2268 2616 2276 2624
rect 2380 2616 2388 2624
rect 2236 2596 2244 2604
rect 2396 2596 2404 2604
rect 2572 2936 2580 2944
rect 2620 2936 2628 2944
rect 2812 3416 2820 3424
rect 3084 3496 3092 3504
rect 3308 3556 3316 3564
rect 3356 3536 3364 3544
rect 3276 3496 3284 3504
rect 3052 3476 3060 3484
rect 3068 3476 3076 3484
rect 3100 3476 3108 3484
rect 2972 3416 2980 3424
rect 2908 3396 2916 3404
rect 3004 3396 3012 3404
rect 3052 3416 3060 3424
rect 3100 3396 3108 3404
rect 3068 3376 3076 3384
rect 2844 3356 2852 3364
rect 2876 3356 2884 3364
rect 3084 3356 3092 3364
rect 3036 3336 3044 3344
rect 2748 3316 2756 3324
rect 2796 3316 2804 3324
rect 2828 3316 2836 3324
rect 2876 3316 2884 3324
rect 2940 3316 2948 3324
rect 2764 3296 2772 3304
rect 2924 3296 2932 3304
rect 2988 3256 2996 3264
rect 3020 3256 3028 3264
rect 2732 3236 2740 3244
rect 2988 3236 2996 3244
rect 2956 3216 2964 3224
rect 2828 3176 2836 3184
rect 2796 3136 2804 3144
rect 2716 3076 2724 3084
rect 2748 3076 2756 3084
rect 2764 3076 2772 3084
rect 2796 3076 2804 3084
rect 2684 3056 2692 3064
rect 2748 2996 2756 3004
rect 2652 2956 2660 2964
rect 2668 2956 2676 2964
rect 2716 2956 2724 2964
rect 2764 2956 2772 2964
rect 2780 2956 2788 2964
rect 2668 2936 2676 2944
rect 2588 2876 2596 2884
rect 2572 2856 2580 2864
rect 2636 2876 2644 2884
rect 2668 2876 2676 2884
rect 2620 2856 2628 2864
rect 2492 2736 2500 2744
rect 2508 2716 2516 2724
rect 2604 2716 2612 2724
rect 2492 2636 2500 2644
rect 2444 2616 2452 2624
rect 2476 2616 2484 2624
rect 2620 2676 2628 2684
rect 2604 2636 2612 2644
rect 2124 2556 2132 2564
rect 2156 2556 2164 2564
rect 2188 2556 2196 2564
rect 2396 2576 2404 2584
rect 2412 2576 2420 2584
rect 2460 2576 2468 2584
rect 2508 2576 2516 2584
rect 2540 2596 2548 2604
rect 2316 2556 2324 2564
rect 2380 2556 2388 2564
rect 2396 2556 2404 2564
rect 2060 2496 2068 2504
rect 2124 2496 2132 2504
rect 2220 2496 2228 2504
rect 2364 2536 2372 2544
rect 2444 2536 2452 2544
rect 2492 2536 2500 2544
rect 2556 2536 2564 2544
rect 2668 2856 2676 2864
rect 2652 2816 2660 2824
rect 2684 2836 2692 2844
rect 2716 2816 2724 2824
rect 2668 2736 2676 2744
rect 2700 2736 2708 2744
rect 2764 2816 2772 2824
rect 2796 2816 2804 2824
rect 2684 2656 2692 2664
rect 2636 2636 2644 2644
rect 2668 2636 2676 2644
rect 2700 2636 2708 2644
rect 2924 3156 2932 3164
rect 2924 3136 2932 3144
rect 2844 3076 2852 3084
rect 2908 3076 2916 3084
rect 2892 2996 2900 3004
rect 3036 3196 3044 3204
rect 3020 3156 3028 3164
rect 3084 3316 3092 3324
rect 3020 3136 3028 3144
rect 3036 3136 3044 3144
rect 3068 3136 3076 3144
rect 3132 3396 3140 3404
rect 3148 3376 3156 3384
rect 3404 3516 3412 3524
rect 3468 3516 3476 3524
rect 3196 3416 3204 3424
rect 3484 3496 3492 3504
rect 3660 3576 3668 3584
rect 3692 3576 3700 3584
rect 3788 3576 3796 3584
rect 3884 3576 3892 3584
rect 3564 3496 3572 3504
rect 3436 3456 3444 3464
rect 3516 3456 3524 3464
rect 3532 3456 3540 3464
rect 3276 3436 3284 3444
rect 3324 3436 3332 3444
rect 3340 3436 3348 3444
rect 3404 3436 3412 3444
rect 3548 3436 3556 3444
rect 3596 3456 3604 3464
rect 3612 3456 3620 3464
rect 4140 3576 4148 3584
rect 3804 3476 3812 3484
rect 3852 3476 3860 3484
rect 3900 3476 3908 3484
rect 3916 3476 3924 3484
rect 3948 3476 3956 3484
rect 3964 3476 3972 3484
rect 3980 3476 3988 3484
rect 3996 3476 4004 3484
rect 4044 3476 4052 3484
rect 3644 3456 3652 3464
rect 3228 3416 3236 3424
rect 3180 3396 3188 3404
rect 3212 3396 3220 3404
rect 3148 3356 3156 3364
rect 3164 3356 3172 3364
rect 3132 3316 3140 3324
rect 3068 3096 3076 3104
rect 2956 3076 2964 3084
rect 2972 3076 2980 3084
rect 3068 3056 3076 3064
rect 3084 3036 3092 3044
rect 3164 3316 3172 3324
rect 3244 3396 3252 3404
rect 3388 3396 3396 3404
rect 3260 3376 3268 3384
rect 3356 3376 3364 3384
rect 3484 3376 3492 3384
rect 3308 3356 3316 3364
rect 3340 3356 3348 3364
rect 3388 3356 3396 3364
rect 3484 3356 3492 3364
rect 3500 3356 3508 3364
rect 3404 3336 3412 3344
rect 3436 3336 3444 3344
rect 3452 3336 3460 3344
rect 3548 3396 3556 3404
rect 3708 3396 3716 3404
rect 3724 3396 3732 3404
rect 4332 3596 4340 3604
rect 4044 3436 4052 3444
rect 3756 3416 3764 3424
rect 3804 3396 3812 3404
rect 3548 3356 3556 3364
rect 3708 3356 3716 3364
rect 3500 3316 3508 3324
rect 3532 3316 3540 3324
rect 3196 3256 3204 3264
rect 3244 3256 3252 3264
rect 3276 3256 3284 3264
rect 3388 3256 3396 3264
rect 3484 3256 3492 3264
rect 3132 3216 3140 3224
rect 3244 3216 3252 3224
rect 3436 3216 3444 3224
rect 3116 3196 3124 3204
rect 3116 3176 3124 3184
rect 3452 3136 3460 3144
rect 3452 3116 3460 3124
rect 3356 3096 3364 3104
rect 3388 3096 3396 3104
rect 3292 3076 3300 3084
rect 3308 3076 3316 3084
rect 3356 3076 3364 3084
rect 3388 3076 3396 3084
rect 3164 3036 3172 3044
rect 2988 3016 2996 3024
rect 3100 3016 3108 3024
rect 2956 2996 2964 3004
rect 2988 2996 2996 3004
rect 2844 2956 2852 2964
rect 2812 2736 2820 2744
rect 2828 2736 2836 2744
rect 3020 2936 3028 2944
rect 3052 2936 3060 2944
rect 3212 3056 3220 3064
rect 3276 3056 3284 3064
rect 3228 3036 3236 3044
rect 3212 3016 3220 3024
rect 3340 3056 3348 3064
rect 3388 3056 3396 3064
rect 3292 3036 3300 3044
rect 3260 2976 3268 2984
rect 3564 3316 3572 3324
rect 3660 3316 3668 3324
rect 3740 3376 3748 3384
rect 3900 3416 3908 3424
rect 4156 3436 4164 3444
rect 4092 3416 4100 3424
rect 4748 3616 4756 3624
rect 4796 3616 4804 3624
rect 4652 3596 4660 3604
rect 4508 3576 4516 3584
rect 4428 3536 4436 3544
rect 4380 3516 4388 3524
rect 4412 3516 4420 3524
rect 4460 3516 4468 3524
rect 4572 3496 4580 3504
rect 4604 3496 4612 3504
rect 4876 3596 4884 3604
rect 4796 3556 4804 3564
rect 4748 3536 4756 3544
rect 4716 3496 4724 3504
rect 4748 3496 4756 3504
rect 4300 3476 4308 3484
rect 4316 3476 4324 3484
rect 4396 3476 4404 3484
rect 4476 3476 4484 3484
rect 4508 3476 4516 3484
rect 4556 3476 4564 3484
rect 4620 3476 4628 3484
rect 4652 3476 4660 3484
rect 4236 3456 4244 3464
rect 4252 3456 4260 3464
rect 4204 3436 4212 3444
rect 4172 3416 4180 3424
rect 4076 3396 4084 3404
rect 4108 3396 4116 3404
rect 4156 3396 4164 3404
rect 4364 3456 4372 3464
rect 4460 3456 4468 3464
rect 4556 3456 4564 3464
rect 4396 3436 4404 3444
rect 4444 3436 4452 3444
rect 4444 3416 4452 3424
rect 4300 3396 4308 3404
rect 4332 3396 4340 3404
rect 4268 3376 4276 3384
rect 3756 3356 3764 3364
rect 3788 3356 3796 3364
rect 3836 3356 3844 3364
rect 3852 3356 3860 3364
rect 3948 3356 3956 3364
rect 3996 3356 4004 3364
rect 4028 3356 4036 3364
rect 4044 3356 4052 3364
rect 3852 3336 3860 3344
rect 3916 3336 3924 3344
rect 3964 3336 3972 3344
rect 3996 3336 4004 3344
rect 4076 3336 4084 3344
rect 4092 3336 4100 3344
rect 4188 3336 4196 3344
rect 3740 3316 3748 3324
rect 3756 3316 3764 3324
rect 3900 3316 3908 3324
rect 3804 3296 3812 3304
rect 3820 3296 3828 3304
rect 3612 3276 3620 3284
rect 3852 3296 3860 3304
rect 3724 3196 3732 3204
rect 3772 3196 3780 3204
rect 3836 3196 3844 3204
rect 3516 3156 3524 3164
rect 3692 3156 3700 3164
rect 3532 3136 3540 3144
rect 3532 3116 3540 3124
rect 3564 3116 3572 3124
rect 3580 3116 3588 3124
rect 3644 3116 3652 3124
rect 3420 3056 3428 3064
rect 3452 3056 3460 3064
rect 3516 3056 3524 3064
rect 3564 3056 3572 3064
rect 3436 3036 3444 3044
rect 3484 3036 3492 3044
rect 3548 3036 3556 3044
rect 3484 2996 3492 3004
rect 3532 2996 3540 3004
rect 3548 2996 3556 3004
rect 3468 2976 3476 2984
rect 3500 2976 3508 2984
rect 3340 2956 3348 2964
rect 3292 2936 3300 2944
rect 3324 2936 3332 2944
rect 3132 2916 3140 2924
rect 3148 2916 3156 2924
rect 3180 2916 3188 2924
rect 3244 2916 3252 2924
rect 3036 2896 3044 2904
rect 3100 2896 3108 2904
rect 3148 2896 3156 2904
rect 3196 2896 3204 2904
rect 3228 2896 3236 2904
rect 2940 2876 2948 2884
rect 3004 2876 3012 2884
rect 2956 2816 2964 2824
rect 2988 2796 2996 2804
rect 3036 2796 3044 2804
rect 3084 2796 3092 2804
rect 3116 2756 3124 2764
rect 2924 2736 2932 2744
rect 2940 2736 2948 2744
rect 3052 2736 3060 2744
rect 2844 2676 2852 2684
rect 2860 2656 2868 2664
rect 2908 2656 2916 2664
rect 2748 2636 2756 2644
rect 2892 2636 2900 2644
rect 2732 2576 2740 2584
rect 2828 2576 2836 2584
rect 2636 2536 2644 2544
rect 2700 2556 2708 2564
rect 2748 2556 2756 2564
rect 2812 2556 2820 2564
rect 2876 2556 2884 2564
rect 2908 2556 2916 2564
rect 2268 2496 2276 2504
rect 2300 2496 2308 2504
rect 2348 2496 2356 2504
rect 2540 2496 2548 2504
rect 2668 2496 2676 2504
rect 2364 2476 2372 2484
rect 2412 2476 2420 2484
rect 2540 2476 2548 2484
rect 2252 2456 2260 2464
rect 2012 2436 2020 2444
rect 2044 2356 2052 2364
rect 2396 2416 2404 2424
rect 2332 2396 2340 2404
rect 2348 2396 2356 2404
rect 2236 2356 2244 2364
rect 2300 2356 2308 2364
rect 2316 2356 2324 2364
rect 1836 2316 1844 2324
rect 1916 2316 1924 2324
rect 1244 2276 1252 2284
rect 1228 2196 1236 2204
rect 1244 2196 1252 2204
rect 892 2116 900 2124
rect 940 2116 948 2124
rect 1004 2116 1012 2124
rect 908 1956 916 1964
rect 1052 2116 1060 2124
rect 1100 2116 1108 2124
rect 1180 2116 1188 2124
rect 1212 2156 1220 2164
rect 1276 2296 1284 2304
rect 1292 2296 1300 2304
rect 1404 2296 1412 2304
rect 1452 2296 1460 2304
rect 1468 2296 1476 2304
rect 1532 2296 1540 2304
rect 1596 2296 1604 2304
rect 1644 2296 1652 2304
rect 1740 2296 1748 2304
rect 1756 2296 1764 2304
rect 1916 2296 1924 2304
rect 1308 2276 1316 2284
rect 1612 2256 1620 2264
rect 1340 2236 1348 2244
rect 1420 2236 1428 2244
rect 1436 2236 1444 2244
rect 1516 2236 1524 2244
rect 1564 2236 1572 2244
rect 1628 2236 1636 2244
rect 1276 2196 1284 2204
rect 1388 2196 1396 2204
rect 1532 2196 1540 2204
rect 1580 2196 1588 2204
rect 1628 2196 1636 2204
rect 1292 2156 1300 2164
rect 1324 2156 1332 2164
rect 1356 2156 1364 2164
rect 1468 2156 1476 2164
rect 1564 2156 1572 2164
rect 1084 2096 1092 2104
rect 1036 2056 1044 2064
rect 1148 2016 1156 2024
rect 1196 2016 1204 2024
rect 1020 1996 1028 2004
rect 972 1956 980 1964
rect 892 1896 900 1904
rect 444 1856 452 1864
rect 460 1796 468 1804
rect 524 1776 532 1784
rect 700 1856 708 1864
rect 796 1856 804 1864
rect 748 1796 756 1804
rect 764 1796 772 1804
rect 604 1776 612 1784
rect 652 1776 660 1784
rect 732 1776 740 1784
rect 1276 1996 1284 2004
rect 1308 2136 1316 2144
rect 1308 2116 1316 2124
rect 1228 1956 1236 1964
rect 1260 1956 1268 1964
rect 1052 1916 1060 1924
rect 1212 1916 1220 1924
rect 1260 1916 1268 1924
rect 988 1896 996 1904
rect 1036 1896 1044 1904
rect 1116 1896 1124 1904
rect 988 1876 996 1884
rect 876 1856 884 1864
rect 908 1856 916 1864
rect 892 1776 900 1784
rect 1004 1776 1012 1784
rect 1052 1836 1060 1844
rect 604 1756 612 1764
rect 732 1756 740 1764
rect 780 1756 788 1764
rect 844 1756 852 1764
rect 924 1756 932 1764
rect 364 1736 372 1744
rect 396 1736 404 1744
rect 412 1736 420 1744
rect 444 1736 452 1744
rect 492 1736 500 1744
rect 588 1736 596 1744
rect 348 1696 356 1704
rect 364 1676 372 1684
rect 332 1516 340 1524
rect 412 1696 420 1704
rect 1100 1836 1108 1844
rect 1116 1836 1124 1844
rect 1116 1776 1124 1784
rect 892 1736 900 1744
rect 668 1716 676 1724
rect 796 1716 804 1724
rect 828 1716 836 1724
rect 444 1576 452 1584
rect 572 1696 580 1704
rect 476 1676 484 1684
rect 540 1676 548 1684
rect 700 1696 708 1704
rect 636 1676 644 1684
rect 844 1696 852 1704
rect 604 1656 612 1664
rect 652 1636 660 1644
rect 556 1516 564 1524
rect 588 1516 596 1524
rect 348 1456 356 1464
rect 380 1456 388 1464
rect 316 1436 324 1444
rect 252 1376 260 1384
rect 364 1416 372 1424
rect 412 1416 420 1424
rect 364 1396 372 1404
rect 380 1396 388 1404
rect 796 1616 804 1624
rect 684 1596 692 1604
rect 860 1636 868 1644
rect 732 1536 740 1544
rect 924 1656 932 1664
rect 780 1516 788 1524
rect 876 1516 884 1524
rect 828 1496 836 1504
rect 860 1496 868 1504
rect 908 1496 916 1504
rect 764 1476 772 1484
rect 556 1456 564 1464
rect 540 1436 548 1444
rect 492 1416 500 1424
rect 556 1416 564 1424
rect 444 1376 452 1384
rect 524 1356 532 1364
rect 428 1336 436 1344
rect 284 1316 292 1324
rect 332 1316 340 1324
rect 284 1296 292 1304
rect 332 1256 340 1264
rect 172 1196 180 1204
rect 204 1196 212 1204
rect 380 1216 388 1224
rect 204 1136 212 1144
rect 236 1136 244 1144
rect 108 1096 116 1104
rect 12 1076 20 1084
rect 76 1076 84 1084
rect 28 1056 36 1064
rect 60 1056 68 1064
rect 44 1036 52 1044
rect 28 996 36 1004
rect 12 916 20 924
rect 60 1016 68 1024
rect 124 996 132 1004
rect 284 1056 292 1064
rect 380 1056 388 1064
rect 412 1196 420 1204
rect 444 1316 452 1324
rect 876 1456 884 1464
rect 908 1456 916 1464
rect 652 1436 660 1444
rect 684 1436 692 1444
rect 604 1396 612 1404
rect 636 1356 644 1364
rect 652 1356 660 1364
rect 668 1336 676 1344
rect 492 1316 500 1324
rect 508 1316 516 1324
rect 620 1316 628 1324
rect 652 1316 660 1324
rect 668 1316 676 1324
rect 524 1256 532 1264
rect 476 1236 484 1244
rect 460 1216 468 1224
rect 540 1216 548 1224
rect 764 1376 772 1384
rect 780 1356 788 1364
rect 732 1336 740 1344
rect 764 1336 772 1344
rect 732 1256 740 1264
rect 684 1216 692 1224
rect 716 1216 724 1224
rect 780 1256 788 1264
rect 876 1356 884 1364
rect 812 1336 820 1344
rect 892 1336 900 1344
rect 844 1316 852 1324
rect 876 1316 884 1324
rect 700 1176 708 1184
rect 764 1176 772 1184
rect 796 1176 804 1184
rect 652 1136 660 1144
rect 460 1116 468 1124
rect 476 1116 484 1124
rect 508 1116 516 1124
rect 556 1116 564 1124
rect 572 1116 580 1124
rect 764 1116 772 1124
rect 620 1096 628 1104
rect 716 1096 724 1104
rect 796 1096 804 1104
rect 428 1076 436 1084
rect 524 1076 532 1084
rect 620 1076 628 1084
rect 156 996 164 1004
rect 188 996 196 1004
rect 252 996 260 1004
rect 204 976 212 984
rect 508 1056 516 1064
rect 140 956 148 964
rect 268 956 276 964
rect 284 956 292 964
rect 364 956 372 964
rect 316 936 324 944
rect 348 936 356 944
rect 140 916 148 924
rect 108 896 116 904
rect 236 896 244 904
rect 172 856 180 864
rect 156 796 164 804
rect 44 756 52 764
rect 60 756 68 764
rect 140 736 148 744
rect 12 696 20 704
rect 332 876 340 884
rect 300 856 308 864
rect 396 956 404 964
rect 380 836 388 844
rect 316 796 324 804
rect 348 796 356 804
rect 252 756 260 764
rect 188 736 196 744
rect 268 736 276 744
rect 236 716 244 724
rect 284 716 292 724
rect 652 996 660 1004
rect 844 1216 852 1224
rect 860 1216 868 1224
rect 844 1176 852 1184
rect 828 1156 836 1164
rect 732 1016 740 1024
rect 524 976 532 984
rect 732 976 740 984
rect 748 976 756 984
rect 444 956 452 964
rect 476 956 484 964
rect 620 956 628 964
rect 540 936 548 944
rect 524 916 532 924
rect 572 916 580 924
rect 716 916 724 924
rect 380 736 388 744
rect 684 876 692 884
rect 428 776 436 784
rect 220 676 228 684
rect 332 676 340 684
rect 412 676 420 684
rect 476 736 484 744
rect 60 656 68 664
rect 332 656 340 664
rect 380 656 388 664
rect 428 656 436 664
rect 124 636 132 644
rect 44 556 52 564
rect 92 536 100 544
rect 60 496 68 504
rect 28 416 36 424
rect 12 316 20 324
rect 44 316 52 324
rect 156 556 164 564
rect 204 616 212 624
rect 220 576 228 584
rect 268 556 276 564
rect 156 536 164 544
rect 188 536 196 544
rect 236 536 244 544
rect 348 616 356 624
rect 364 536 372 544
rect 444 596 452 604
rect 540 736 548 744
rect 556 716 564 724
rect 604 716 612 724
rect 908 1176 916 1184
rect 892 1096 900 1104
rect 956 1636 964 1644
rect 988 1696 996 1704
rect 972 1576 980 1584
rect 940 1536 948 1544
rect 1100 1696 1108 1704
rect 1116 1696 1124 1704
rect 1244 1856 1252 1864
rect 1196 1796 1204 1804
rect 1340 2096 1348 2104
rect 1356 2096 1364 2104
rect 1500 2096 1508 2104
rect 1516 2056 1524 2064
rect 1564 2056 1572 2064
rect 1420 2036 1428 2044
rect 1548 2036 1556 2044
rect 1388 1996 1396 2004
rect 1356 1956 1364 1964
rect 1340 1896 1348 1904
rect 1356 1896 1364 1904
rect 1468 1956 1476 1964
rect 1436 1916 1444 1924
rect 1500 1896 1508 1904
rect 1532 1896 1540 1904
rect 1564 1896 1572 1904
rect 1324 1856 1332 1864
rect 1292 1836 1300 1844
rect 1404 1836 1412 1844
rect 1372 1816 1380 1824
rect 1276 1796 1284 1804
rect 1308 1776 1316 1784
rect 1324 1776 1332 1784
rect 1340 1776 1348 1784
rect 1228 1756 1236 1764
rect 1244 1756 1252 1764
rect 1292 1756 1300 1764
rect 1164 1696 1172 1704
rect 1212 1696 1220 1704
rect 1196 1556 1204 1564
rect 1052 1536 1060 1544
rect 1212 1536 1220 1544
rect 1004 1516 1012 1524
rect 1020 1516 1028 1524
rect 1116 1516 1124 1524
rect 1196 1516 1204 1524
rect 1388 1756 1396 1764
rect 1548 1836 1556 1844
rect 1484 1816 1492 1824
rect 1516 1816 1524 1824
rect 1564 1816 1572 1824
rect 1500 1756 1508 1764
rect 1500 1736 1508 1744
rect 1260 1716 1268 1724
rect 1292 1716 1300 1724
rect 1340 1716 1348 1724
rect 1356 1716 1364 1724
rect 1436 1696 1444 1704
rect 1452 1696 1460 1704
rect 1596 2156 1604 2164
rect 1644 2156 1652 2164
rect 1660 2156 1668 2164
rect 1644 2076 1652 2084
rect 1692 2156 1700 2164
rect 1708 2156 1716 2164
rect 1628 2056 1636 2064
rect 1676 2056 1684 2064
rect 1708 2016 1716 2024
rect 1756 2196 1764 2204
rect 1804 2256 1812 2264
rect 1836 2236 1844 2244
rect 1852 2236 1860 2244
rect 1836 2216 1844 2224
rect 1788 2196 1796 2204
rect 1772 2176 1780 2184
rect 1740 2156 1748 2164
rect 1804 2156 1812 2164
rect 1884 2256 1892 2264
rect 1900 2236 1908 2244
rect 1884 2216 1892 2224
rect 1820 2076 1828 2084
rect 1836 2076 1844 2084
rect 1740 2056 1748 2064
rect 1772 1976 1780 1984
rect 1900 2076 1908 2084
rect 1868 1976 1876 1984
rect 1852 1956 1860 1964
rect 1676 1916 1684 1924
rect 1740 1916 1748 1924
rect 1804 1916 1812 1924
rect 1820 1916 1828 1924
rect 1852 1916 1860 1924
rect 1884 1916 1892 1924
rect 2060 2316 2068 2324
rect 2316 2316 2324 2324
rect 2076 2296 2084 2304
rect 2156 2296 2164 2304
rect 2172 2296 2180 2304
rect 2220 2296 2228 2304
rect 2236 2296 2244 2304
rect 2604 2436 2612 2444
rect 2444 2416 2452 2424
rect 2604 2416 2612 2424
rect 2412 2396 2420 2404
rect 2428 2396 2436 2404
rect 2444 2396 2452 2404
rect 2540 2396 2548 2404
rect 2508 2376 2516 2384
rect 2412 2336 2420 2344
rect 2492 2336 2500 2344
rect 2412 2316 2420 2324
rect 2444 2296 2452 2304
rect 2476 2296 2484 2304
rect 1964 2276 1972 2284
rect 1996 2276 2004 2284
rect 2076 2276 2084 2284
rect 2124 2276 2132 2284
rect 2364 2276 2372 2284
rect 2412 2276 2420 2284
rect 2444 2276 2452 2284
rect 1932 2216 1940 2224
rect 2012 2236 2020 2244
rect 2028 2236 2036 2244
rect 1980 2216 1988 2224
rect 2092 2216 2100 2224
rect 2076 2196 2084 2204
rect 2108 2196 2116 2204
rect 2028 2136 2036 2144
rect 2060 2136 2068 2144
rect 1980 2116 1988 2124
rect 1948 2076 1956 2084
rect 1980 2076 1988 2084
rect 2204 2216 2212 2224
rect 2220 2216 2228 2224
rect 2252 2196 2260 2204
rect 2348 2236 2356 2244
rect 2284 2216 2292 2224
rect 2380 2216 2388 2224
rect 2156 2116 2164 2124
rect 2076 2076 2084 2084
rect 2012 2056 2020 2064
rect 2044 2056 2052 2064
rect 2060 2056 2068 2064
rect 2124 2016 2132 2024
rect 2140 2016 2148 2024
rect 1596 1896 1604 1904
rect 1724 1896 1732 1904
rect 1772 1896 1780 1904
rect 1596 1836 1604 1844
rect 1644 1836 1652 1844
rect 1692 1816 1700 1824
rect 1596 1776 1604 1784
rect 1628 1776 1636 1784
rect 1564 1756 1572 1764
rect 1692 1756 1700 1764
rect 1932 1916 1940 1924
rect 2044 1916 2052 1924
rect 2076 1916 2084 1924
rect 2108 1896 2116 1904
rect 1740 1756 1748 1764
rect 1292 1676 1300 1684
rect 1244 1556 1252 1564
rect 1260 1536 1268 1544
rect 1292 1536 1300 1544
rect 1404 1536 1412 1544
rect 1244 1516 1252 1524
rect 956 1496 964 1504
rect 1132 1496 1140 1504
rect 1228 1496 1236 1504
rect 940 1476 948 1484
rect 1084 1456 1092 1464
rect 940 1436 948 1444
rect 1020 1416 1028 1424
rect 1084 1416 1092 1424
rect 972 1356 980 1364
rect 1740 1736 1748 1744
rect 1772 1816 1780 1824
rect 1868 1816 1876 1824
rect 1932 1836 1940 1844
rect 1932 1816 1940 1824
rect 1964 1816 1972 1824
rect 1996 1816 2004 1824
rect 2012 1816 2020 1824
rect 1788 1756 1796 1764
rect 1532 1636 1540 1644
rect 1644 1636 1652 1644
rect 1676 1636 1684 1644
rect 1708 1636 1716 1644
rect 1580 1576 1588 1584
rect 1596 1576 1604 1584
rect 1532 1516 1540 1524
rect 1868 1736 1876 1744
rect 1788 1696 1796 1704
rect 1836 1696 1844 1704
rect 1916 1736 1924 1744
rect 1916 1696 1924 1704
rect 1884 1676 1892 1684
rect 1820 1576 1828 1584
rect 2204 2136 2212 2144
rect 2492 2276 2500 2284
rect 2524 2296 2532 2304
rect 2572 2296 2580 2304
rect 2588 2296 2596 2304
rect 2668 2436 2676 2444
rect 2652 2356 2660 2364
rect 2716 2496 2724 2504
rect 2764 2496 2772 2504
rect 2780 2496 2788 2504
rect 2732 2476 2740 2484
rect 3100 2716 3108 2724
rect 3068 2696 3076 2704
rect 3324 2896 3332 2904
rect 3372 2896 3380 2904
rect 3276 2776 3284 2784
rect 3292 2776 3300 2784
rect 3420 2896 3428 2904
rect 3404 2856 3412 2864
rect 3388 2816 3396 2824
rect 3164 2756 3172 2764
rect 3356 2756 3364 2764
rect 3164 2736 3172 2744
rect 3196 2736 3204 2744
rect 3468 2916 3476 2924
rect 3772 3176 3780 3184
rect 3836 3176 3844 3184
rect 3804 3156 3812 3164
rect 4028 3316 4036 3324
rect 4172 3316 4180 3324
rect 4220 3316 4228 3324
rect 3980 3296 3988 3304
rect 4044 3296 4052 3304
rect 3932 3136 3940 3144
rect 4028 3136 4036 3144
rect 4108 3136 4116 3144
rect 3740 3116 3748 3124
rect 4028 3116 4036 3124
rect 4044 3116 4052 3124
rect 3932 3096 3940 3104
rect 4076 3096 4084 3104
rect 3628 3056 3636 3064
rect 3692 3056 3700 3064
rect 3676 3036 3684 3044
rect 3596 3016 3604 3024
rect 3580 2996 3588 3004
rect 3612 2956 3620 2964
rect 3692 2956 3700 2964
rect 3532 2916 3540 2924
rect 3596 2916 3604 2924
rect 3708 2936 3716 2944
rect 3660 2916 3668 2924
rect 3708 2916 3716 2924
rect 3548 2896 3556 2904
rect 3628 2896 3636 2904
rect 3644 2836 3652 2844
rect 3516 2796 3524 2804
rect 3516 2776 3524 2784
rect 3484 2756 3492 2764
rect 3660 2736 3668 2744
rect 3212 2716 3220 2724
rect 3308 2716 3316 2724
rect 3356 2716 3364 2724
rect 3388 2716 3396 2724
rect 3436 2716 3444 2724
rect 3484 2716 3492 2724
rect 3532 2716 3540 2724
rect 3548 2716 3556 2724
rect 2940 2676 2948 2684
rect 3148 2676 3156 2684
rect 2956 2576 2964 2584
rect 2988 2636 2996 2644
rect 3004 2636 3012 2644
rect 3212 2656 3220 2664
rect 3244 2656 3252 2664
rect 3100 2636 3108 2644
rect 3132 2636 3140 2644
rect 3292 2656 3300 2664
rect 3388 2656 3396 2664
rect 3628 2656 3636 2664
rect 3564 2636 3572 2644
rect 3612 2636 3620 2644
rect 3660 2636 3668 2644
rect 3676 2636 3684 2644
rect 3756 2896 3764 2904
rect 3708 2696 3716 2704
rect 3740 2656 3748 2664
rect 3260 2616 3268 2624
rect 3436 2616 3444 2624
rect 3500 2616 3508 2624
rect 3596 2616 3604 2624
rect 3180 2596 3188 2604
rect 3244 2596 3252 2604
rect 3260 2596 3268 2604
rect 2940 2556 2948 2564
rect 2972 2556 2980 2564
rect 3004 2556 3012 2564
rect 3020 2556 3028 2564
rect 2924 2516 2932 2524
rect 2924 2496 2932 2504
rect 2940 2496 2948 2504
rect 2844 2476 2852 2484
rect 2860 2476 2868 2484
rect 2876 2476 2884 2484
rect 2812 2436 2820 2444
rect 2748 2416 2756 2424
rect 2716 2396 2724 2404
rect 2492 2196 2500 2204
rect 2508 2176 2516 2184
rect 2460 2136 2468 2144
rect 2476 2136 2484 2144
rect 2492 2136 2500 2144
rect 2188 2116 2196 2124
rect 2284 2116 2292 2124
rect 2252 2096 2260 2104
rect 2172 2056 2180 2064
rect 2172 2016 2180 2024
rect 2188 1936 2196 1944
rect 2220 1936 2228 1944
rect 2188 1896 2196 1904
rect 2236 1896 2244 1904
rect 2140 1816 2148 1824
rect 2156 1816 2164 1824
rect 1964 1756 1972 1764
rect 1980 1756 1988 1764
rect 2012 1756 2020 1764
rect 1948 1736 1956 1744
rect 1932 1596 1940 1604
rect 1948 1596 1956 1604
rect 1900 1556 1908 1564
rect 1804 1536 1812 1544
rect 1900 1536 1908 1544
rect 1372 1496 1380 1504
rect 1404 1496 1412 1504
rect 1452 1496 1460 1504
rect 1548 1496 1556 1504
rect 1612 1496 1620 1504
rect 1660 1496 1668 1504
rect 1708 1516 1716 1524
rect 1148 1416 1156 1424
rect 1228 1416 1236 1424
rect 1180 1396 1188 1404
rect 1564 1476 1572 1484
rect 1372 1456 1380 1464
rect 1404 1456 1412 1464
rect 1276 1416 1284 1424
rect 1340 1416 1348 1424
rect 1356 1416 1364 1424
rect 1388 1416 1396 1424
rect 1404 1416 1412 1424
rect 940 1336 948 1344
rect 972 1336 980 1344
rect 1020 1336 1028 1344
rect 1116 1336 1124 1344
rect 1180 1336 1188 1344
rect 1212 1336 1220 1344
rect 1244 1336 1252 1344
rect 1292 1336 1300 1344
rect 972 1216 980 1224
rect 1116 1296 1124 1304
rect 1212 1296 1220 1304
rect 1068 1256 1076 1264
rect 988 1176 996 1184
rect 1036 1176 1044 1184
rect 1052 1176 1060 1184
rect 972 1096 980 1104
rect 988 1076 996 1084
rect 844 1056 852 1064
rect 1020 1036 1028 1044
rect 860 996 868 1004
rect 844 976 852 984
rect 1100 1156 1108 1164
rect 1180 1136 1188 1144
rect 1100 1116 1108 1124
rect 1116 1116 1124 1124
rect 1164 1116 1172 1124
rect 1260 1156 1268 1164
rect 1260 1136 1268 1144
rect 1340 1376 1348 1384
rect 1404 1396 1412 1404
rect 1404 1376 1412 1384
rect 1388 1296 1396 1304
rect 1324 1256 1332 1264
rect 1340 1216 1348 1224
rect 1308 1136 1316 1144
rect 1356 1116 1364 1124
rect 1068 1076 1076 1084
rect 1148 1076 1156 1084
rect 1180 1076 1188 1084
rect 1196 1076 1204 1084
rect 1244 1076 1252 1084
rect 1052 996 1060 1004
rect 1004 976 1012 984
rect 764 916 772 924
rect 796 916 804 924
rect 764 876 772 884
rect 764 736 772 744
rect 524 676 532 684
rect 620 676 628 684
rect 508 656 516 664
rect 492 596 500 604
rect 524 596 532 604
rect 540 596 548 604
rect 412 556 420 564
rect 508 556 516 564
rect 652 676 660 684
rect 620 596 628 604
rect 700 616 708 624
rect 764 576 772 584
rect 780 576 788 584
rect 572 556 580 564
rect 684 556 692 564
rect 828 876 836 884
rect 876 876 884 884
rect 844 816 852 824
rect 812 736 820 744
rect 956 896 964 904
rect 1116 1016 1124 1024
rect 1148 1016 1156 1024
rect 1132 996 1140 1004
rect 1116 976 1124 984
rect 1356 1056 1364 1064
rect 1388 1056 1396 1064
rect 1180 1016 1188 1024
rect 1180 996 1188 1004
rect 1212 976 1220 984
rect 1068 896 1076 904
rect 1196 936 1204 944
rect 1132 856 1140 864
rect 1020 836 1028 844
rect 860 696 868 704
rect 892 696 900 704
rect 812 636 820 644
rect 812 576 820 584
rect 828 576 836 584
rect 924 616 932 624
rect 924 576 932 584
rect 972 616 980 624
rect 972 596 980 604
rect 860 536 868 544
rect 956 536 964 544
rect 1308 996 1316 1004
rect 1500 1396 1508 1404
rect 1548 1396 1556 1404
rect 1484 1376 1492 1384
rect 1548 1376 1556 1384
rect 1420 1276 1428 1284
rect 1436 1196 1444 1204
rect 1468 1316 1476 1324
rect 1484 1296 1492 1304
rect 1532 1296 1540 1304
rect 1500 1216 1508 1224
rect 1516 1216 1524 1224
rect 1420 1156 1428 1164
rect 1452 1156 1460 1164
rect 1740 1496 1748 1504
rect 1772 1496 1780 1504
rect 1852 1496 1860 1504
rect 1660 1476 1668 1484
rect 1692 1476 1700 1484
rect 1612 1456 1620 1464
rect 1596 1396 1604 1404
rect 1628 1396 1636 1404
rect 1644 1396 1652 1404
rect 1580 1376 1588 1384
rect 1628 1376 1636 1384
rect 1676 1396 1684 1404
rect 1692 1396 1700 1404
rect 1756 1396 1764 1404
rect 1580 1256 1588 1264
rect 1580 1236 1588 1244
rect 1436 1136 1444 1144
rect 1516 1136 1524 1144
rect 1532 1136 1540 1144
rect 1564 1136 1572 1144
rect 1484 1116 1492 1124
rect 1436 1076 1444 1084
rect 1452 1076 1460 1084
rect 1708 1376 1716 1384
rect 1660 1156 1668 1164
rect 1644 1136 1652 1144
rect 1564 1116 1572 1124
rect 1612 1116 1620 1124
rect 1692 1116 1700 1124
rect 1612 1096 1620 1104
rect 1452 1036 1460 1044
rect 1580 1016 1588 1024
rect 1452 996 1460 1004
rect 1308 976 1316 984
rect 1404 976 1412 984
rect 1500 976 1508 984
rect 1244 936 1252 944
rect 1276 936 1284 944
rect 1164 836 1172 844
rect 1148 796 1156 804
rect 1228 876 1236 884
rect 1036 776 1044 784
rect 1180 776 1188 784
rect 1116 756 1124 764
rect 1148 756 1156 764
rect 1004 736 1012 744
rect 1036 736 1044 744
rect 1084 736 1092 744
rect 1004 696 1012 704
rect 1052 696 1060 704
rect 1084 696 1092 704
rect 1100 696 1108 704
rect 1180 696 1188 704
rect 1036 636 1044 644
rect 1004 616 1012 624
rect 1100 616 1108 624
rect 1148 616 1156 624
rect 1116 596 1124 604
rect 1132 596 1140 604
rect 988 576 996 584
rect 1020 576 1028 584
rect 1068 556 1076 564
rect 204 516 212 524
rect 332 516 340 524
rect 492 516 500 524
rect 556 516 564 524
rect 796 516 804 524
rect 828 516 836 524
rect 876 516 884 524
rect 892 516 900 524
rect 908 516 916 524
rect 988 516 996 524
rect 332 496 340 504
rect 588 496 596 504
rect 652 496 660 504
rect 316 476 324 484
rect 652 476 660 484
rect 92 296 100 304
rect 124 296 132 304
rect 140 296 148 304
rect 172 296 180 304
rect 316 356 324 364
rect 268 316 276 324
rect 236 296 244 304
rect 284 296 292 304
rect 540 336 548 344
rect 604 336 612 344
rect 636 336 644 344
rect 380 316 388 324
rect 428 316 436 324
rect 460 316 468 324
rect 332 296 340 304
rect 364 296 372 304
rect 44 276 52 284
rect 236 276 244 284
rect 188 256 196 264
rect 316 256 324 264
rect 332 256 340 264
rect 76 216 84 224
rect 124 236 132 244
rect 284 236 292 244
rect 124 176 132 184
rect 124 136 132 144
rect 188 136 196 144
rect 188 116 196 124
rect 220 116 228 124
rect 300 176 308 184
rect 268 156 276 164
rect 588 276 596 284
rect 412 236 420 244
rect 476 236 484 244
rect 508 236 516 244
rect 396 216 404 224
rect 332 176 340 184
rect 364 176 372 184
rect 556 216 564 224
rect 572 196 580 204
rect 444 176 452 184
rect 572 176 580 184
rect 428 156 436 164
rect 476 156 484 164
rect 556 156 564 164
rect 892 476 900 484
rect 956 476 964 484
rect 1340 916 1348 924
rect 1388 876 1396 884
rect 1372 856 1380 864
rect 1340 836 1348 844
rect 1324 756 1332 764
rect 1324 736 1332 744
rect 1324 696 1332 704
rect 1196 656 1204 664
rect 1212 656 1220 664
rect 1228 636 1236 644
rect 1244 616 1252 624
rect 1180 596 1188 604
rect 1228 596 1236 604
rect 1484 936 1492 944
rect 1532 916 1540 924
rect 1468 896 1476 904
rect 1484 896 1492 904
rect 1420 816 1428 824
rect 1372 776 1380 784
rect 1436 776 1444 784
rect 1388 736 1396 744
rect 1356 696 1364 704
rect 1564 876 1572 884
rect 1548 836 1556 844
rect 1500 756 1508 764
rect 1484 716 1492 724
rect 1516 716 1524 724
rect 1452 676 1460 684
rect 1644 996 1652 1004
rect 1676 1076 1684 1084
rect 1724 1316 1732 1324
rect 1756 1316 1764 1324
rect 1804 1476 1812 1484
rect 1868 1476 1876 1484
rect 1900 1476 1908 1484
rect 1916 1476 1924 1484
rect 1820 1396 1828 1404
rect 1836 1396 1844 1404
rect 1932 1396 1940 1404
rect 1852 1356 1860 1364
rect 1884 1356 1892 1364
rect 1900 1356 1908 1364
rect 1916 1356 1924 1364
rect 1740 1256 1748 1264
rect 1756 1176 1764 1184
rect 1756 1116 1764 1124
rect 1740 1096 1748 1104
rect 1852 1316 1860 1324
rect 1884 1316 1892 1324
rect 1916 1316 1924 1324
rect 1804 1296 1812 1304
rect 1916 1296 1924 1304
rect 2028 1736 2036 1744
rect 1996 1716 2004 1724
rect 2012 1716 2020 1724
rect 2044 1596 2052 1604
rect 1996 1576 2004 1584
rect 2092 1796 2100 1804
rect 2124 1796 2132 1804
rect 2140 1756 2148 1764
rect 2172 1756 2180 1764
rect 2236 1756 2244 1764
rect 2092 1736 2100 1744
rect 2108 1736 2116 1744
rect 2124 1736 2132 1744
rect 2188 1736 2196 1744
rect 2220 1736 2228 1744
rect 2156 1656 2164 1664
rect 2236 1656 2244 1664
rect 2124 1616 2132 1624
rect 2140 1616 2148 1624
rect 2220 1596 2228 1604
rect 2204 1576 2212 1584
rect 2188 1556 2196 1564
rect 2188 1516 2196 1524
rect 1964 1496 1972 1504
rect 2060 1496 2068 1504
rect 2140 1496 2148 1504
rect 2156 1496 2164 1504
rect 2012 1476 2020 1484
rect 2044 1476 2052 1484
rect 2092 1476 2100 1484
rect 2332 2076 2340 2084
rect 2300 2016 2308 2024
rect 2380 2116 2388 2124
rect 2572 2276 2580 2284
rect 2604 2276 2612 2284
rect 2572 2236 2580 2244
rect 2588 2216 2596 2224
rect 2556 2196 2564 2204
rect 2620 2216 2628 2224
rect 2700 2336 2708 2344
rect 2700 2216 2708 2224
rect 2604 2156 2612 2164
rect 2700 2176 2708 2184
rect 2796 2396 2804 2404
rect 2748 2336 2756 2344
rect 2780 2336 2788 2344
rect 2860 2336 2868 2344
rect 2780 2296 2788 2304
rect 2828 2296 2836 2304
rect 2764 2276 2772 2284
rect 2796 2276 2804 2284
rect 2812 2276 2820 2284
rect 2876 2276 2884 2284
rect 2732 2216 2740 2224
rect 2796 2216 2804 2224
rect 2892 2216 2900 2224
rect 2828 2196 2836 2204
rect 2844 2196 2852 2204
rect 2892 2196 2900 2204
rect 2908 2196 2916 2204
rect 2652 2156 2660 2164
rect 2524 2116 2532 2124
rect 2668 2116 2676 2124
rect 2492 2096 2500 2104
rect 2508 2096 2516 2104
rect 2396 2036 2404 2044
rect 2412 2036 2420 2044
rect 2460 2036 2468 2044
rect 2284 1996 2292 2004
rect 2316 1936 2324 1944
rect 2300 1896 2308 1904
rect 2316 1856 2324 1864
rect 2444 1956 2452 1964
rect 2524 2016 2532 2024
rect 2556 2016 2564 2024
rect 2636 2076 2644 2084
rect 2668 2076 2676 2084
rect 2812 2116 2820 2124
rect 2828 2116 2836 2124
rect 2860 2116 2868 2124
rect 2732 2056 2740 2064
rect 2748 2056 2756 2064
rect 2796 2056 2804 2064
rect 2604 2016 2612 2024
rect 2620 2016 2628 2024
rect 2652 2016 2660 2024
rect 2668 2016 2676 2024
rect 2684 2016 2692 2024
rect 2716 2016 2724 2024
rect 2476 1956 2484 1964
rect 2556 1956 2564 1964
rect 2588 1956 2596 1964
rect 2604 1956 2612 1964
rect 2652 1956 2660 1964
rect 2588 1916 2596 1924
rect 2508 1896 2516 1904
rect 2524 1896 2532 1904
rect 2636 1896 2644 1904
rect 2364 1856 2372 1864
rect 2332 1836 2340 1844
rect 2396 1776 2404 1784
rect 2284 1756 2292 1764
rect 2284 1696 2292 1704
rect 2284 1656 2292 1664
rect 2284 1616 2292 1624
rect 2300 1616 2308 1624
rect 2252 1516 2260 1524
rect 2236 1476 2244 1484
rect 2012 1416 2020 1424
rect 2124 1416 2132 1424
rect 2220 1416 2228 1424
rect 1996 1396 2004 1404
rect 1948 1256 1956 1264
rect 1964 1256 1972 1264
rect 1820 1176 1828 1184
rect 1964 1216 1972 1224
rect 1868 1156 1876 1164
rect 1916 1136 1924 1144
rect 1724 1056 1732 1064
rect 1708 996 1716 1004
rect 1660 976 1668 984
rect 1692 976 1700 984
rect 1964 1136 1972 1144
rect 2156 1396 2164 1404
rect 2204 1396 2212 1404
rect 2044 1356 2052 1364
rect 2076 1356 2084 1364
rect 2092 1356 2100 1364
rect 2076 1296 2084 1304
rect 2060 1256 2068 1264
rect 2076 1256 2084 1264
rect 2012 1216 2020 1224
rect 2076 1216 2084 1224
rect 2364 1696 2372 1704
rect 2380 1696 2388 1704
rect 2396 1696 2404 1704
rect 2348 1596 2356 1604
rect 2316 1576 2324 1584
rect 2332 1576 2340 1584
rect 2316 1536 2324 1544
rect 2332 1516 2340 1524
rect 2444 1816 2452 1824
rect 2556 1876 2564 1884
rect 2476 1816 2484 1824
rect 2540 1816 2548 1824
rect 2556 1816 2564 1824
rect 2556 1796 2564 1804
rect 2604 1796 2612 1804
rect 2636 1796 2644 1804
rect 2444 1776 2452 1784
rect 2428 1576 2436 1584
rect 2476 1696 2484 1704
rect 2492 1696 2500 1704
rect 2524 1716 2532 1724
rect 2540 1716 2548 1724
rect 2588 1736 2596 1744
rect 2540 1696 2548 1704
rect 2572 1696 2580 1704
rect 2428 1556 2436 1564
rect 2460 1556 2468 1564
rect 2476 1556 2484 1564
rect 2508 1556 2516 1564
rect 2524 1556 2532 1564
rect 2636 1696 2644 1704
rect 2556 1576 2564 1584
rect 2604 1576 2612 1584
rect 2428 1516 2436 1524
rect 2444 1516 2452 1524
rect 2380 1476 2388 1484
rect 2268 1456 2276 1464
rect 2332 1456 2340 1464
rect 2252 1396 2260 1404
rect 2172 1356 2180 1364
rect 2252 1356 2260 1364
rect 2332 1416 2340 1424
rect 2396 1436 2404 1444
rect 2268 1316 2276 1324
rect 2220 1256 2228 1264
rect 2300 1336 2308 1344
rect 2332 1336 2340 1344
rect 2140 1216 2148 1224
rect 2172 1216 2180 1224
rect 2220 1216 2228 1224
rect 2284 1216 2292 1224
rect 2124 1136 2132 1144
rect 2092 1116 2100 1124
rect 2124 1116 2132 1124
rect 1836 996 1844 1004
rect 1916 1016 1924 1024
rect 1932 1016 1940 1024
rect 1788 976 1796 984
rect 1852 976 1860 984
rect 1868 976 1876 984
rect 1740 956 1748 964
rect 1836 956 1844 964
rect 1900 956 1908 964
rect 2076 1096 2084 1104
rect 1980 1056 1988 1064
rect 2076 1036 2084 1044
rect 1996 1016 2004 1024
rect 2028 1016 2036 1024
rect 2172 1096 2180 1104
rect 2188 1096 2196 1104
rect 2220 1096 2228 1104
rect 2236 1096 2244 1104
rect 2284 1096 2292 1104
rect 2108 1036 2116 1044
rect 2124 1016 2132 1024
rect 2252 1056 2260 1064
rect 2188 1016 2196 1024
rect 2204 1016 2212 1024
rect 2236 1036 2244 1044
rect 1964 956 1972 964
rect 1692 916 1700 924
rect 1708 916 1716 924
rect 1644 856 1652 864
rect 1596 756 1604 764
rect 1724 856 1732 864
rect 1708 836 1716 844
rect 1724 836 1732 844
rect 1708 816 1716 824
rect 1804 876 1812 884
rect 1884 876 1892 884
rect 1756 856 1764 864
rect 1740 796 1748 804
rect 1772 796 1780 804
rect 1660 776 1668 784
rect 1692 776 1700 784
rect 1596 736 1604 744
rect 1644 736 1652 744
rect 1580 716 1588 724
rect 1628 716 1636 724
rect 1804 836 1812 844
rect 1788 736 1796 744
rect 1980 936 1988 944
rect 1996 936 2004 944
rect 2092 936 2100 944
rect 2124 936 2132 944
rect 1980 896 1988 904
rect 2172 916 2180 924
rect 2092 896 2100 904
rect 1932 876 1940 884
rect 1996 876 2004 884
rect 1932 856 1940 864
rect 1948 836 1956 844
rect 1916 796 1924 804
rect 1852 736 1860 744
rect 2092 856 2100 864
rect 2044 816 2052 824
rect 1996 776 2004 784
rect 2028 776 2036 784
rect 2060 776 2068 784
rect 1580 676 1588 684
rect 1660 676 1668 684
rect 1308 616 1316 624
rect 1340 616 1348 624
rect 1292 596 1300 604
rect 1036 516 1044 524
rect 1100 516 1108 524
rect 1228 516 1236 524
rect 1020 496 1028 504
rect 748 456 756 464
rect 1004 456 1012 464
rect 780 356 788 364
rect 828 356 836 364
rect 908 356 916 364
rect 668 336 676 344
rect 732 336 740 344
rect 636 256 644 264
rect 604 216 612 224
rect 604 176 612 184
rect 812 316 820 324
rect 844 316 852 324
rect 908 316 916 324
rect 940 316 948 324
rect 988 316 996 324
rect 764 256 772 264
rect 844 256 852 264
rect 796 236 804 244
rect 652 196 660 204
rect 700 216 708 224
rect 716 216 724 224
rect 684 176 692 184
rect 732 176 740 184
rect 780 156 788 164
rect 892 236 900 244
rect 1116 416 1124 424
rect 1068 396 1076 404
rect 1116 356 1124 364
rect 1132 356 1140 364
rect 1036 316 1044 324
rect 1068 316 1076 324
rect 1100 316 1108 324
rect 1148 316 1156 324
rect 1228 456 1236 464
rect 1212 356 1220 364
rect 1196 316 1204 324
rect 1276 536 1284 544
rect 1596 636 1604 644
rect 1628 636 1636 644
rect 1660 636 1668 644
rect 1740 656 1748 664
rect 1772 636 1780 644
rect 1468 596 1476 604
rect 1532 596 1540 604
rect 1676 616 1684 624
rect 1724 616 1732 624
rect 1756 616 1764 624
rect 1676 556 1684 564
rect 1324 536 1332 544
rect 1372 536 1380 544
rect 1436 536 1444 544
rect 1548 536 1556 544
rect 1580 536 1588 544
rect 1372 516 1380 524
rect 1436 516 1444 524
rect 1500 516 1508 524
rect 1420 496 1428 504
rect 1436 496 1444 504
rect 1388 476 1396 484
rect 1372 436 1380 444
rect 1292 336 1300 344
rect 1340 316 1348 324
rect 1324 296 1332 304
rect 1340 276 1348 284
rect 1356 276 1364 284
rect 988 236 996 244
rect 956 216 964 224
rect 1404 396 1412 404
rect 1708 556 1716 564
rect 1724 556 1732 564
rect 1756 556 1764 564
rect 1612 536 1620 544
rect 1628 536 1636 544
rect 1692 536 1700 544
rect 1708 536 1716 544
rect 1548 376 1556 384
rect 1644 456 1652 464
rect 1676 456 1684 464
rect 1692 456 1700 464
rect 1644 396 1652 404
rect 1660 376 1668 384
rect 1644 356 1652 364
rect 1596 336 1604 344
rect 1612 336 1620 344
rect 1644 336 1652 344
rect 1660 336 1668 344
rect 1676 336 1684 344
rect 1436 276 1444 284
rect 1468 276 1476 284
rect 1484 276 1492 284
rect 1452 236 1460 244
rect 1244 216 1252 224
rect 1276 216 1284 224
rect 924 196 932 204
rect 956 196 964 204
rect 988 196 996 204
rect 1132 196 1140 204
rect 1196 196 1204 204
rect 972 176 980 184
rect 1164 176 1172 184
rect 1196 176 1204 184
rect 1244 176 1252 184
rect 1260 176 1268 184
rect 988 156 996 164
rect 1052 156 1060 164
rect 1084 156 1092 164
rect 1212 156 1220 164
rect 1228 156 1236 164
rect 764 136 772 144
rect 860 136 868 144
rect 876 136 884 144
rect 924 136 932 144
rect 1020 136 1028 144
rect 1356 176 1364 184
rect 1340 156 1348 164
rect 1420 156 1428 164
rect 284 116 292 124
rect 492 116 500 124
rect 220 96 228 104
rect 380 96 388 104
rect 540 96 548 104
rect 636 96 644 104
rect 1180 116 1188 124
rect 1516 176 1524 184
rect 1452 136 1460 144
rect 1564 156 1572 164
rect 1548 136 1556 144
rect 1084 96 1092 104
rect 1452 96 1460 104
rect 1564 96 1572 104
rect 1836 616 1844 624
rect 1916 616 1924 624
rect 2012 716 2020 724
rect 2028 716 2036 724
rect 2108 816 2116 824
rect 2124 796 2132 804
rect 2156 816 2164 824
rect 2140 776 2148 784
rect 2156 756 2164 764
rect 2188 896 2196 904
rect 2188 796 2196 804
rect 2236 976 2244 984
rect 2380 1376 2388 1384
rect 2364 1356 2372 1364
rect 2508 1496 2516 1504
rect 2572 1516 2580 1524
rect 2556 1496 2564 1504
rect 2620 1516 2628 1524
rect 2684 1956 2692 1964
rect 2764 1956 2772 1964
rect 2684 1916 2692 1924
rect 2716 1916 2724 1924
rect 2716 1896 2724 1904
rect 2764 1896 2772 1904
rect 2732 1816 2740 1824
rect 2764 1816 2772 1824
rect 2716 1796 2724 1804
rect 2956 2476 2964 2484
rect 3004 2476 3012 2484
rect 2940 2436 2948 2444
rect 2972 2436 2980 2444
rect 2988 2336 2996 2344
rect 2956 2316 2964 2324
rect 2972 2316 2980 2324
rect 2940 2296 2948 2304
rect 2940 2276 2948 2284
rect 2828 2056 2836 2064
rect 2876 2056 2884 2064
rect 2812 1956 2820 1964
rect 2988 2276 2996 2284
rect 2972 2216 2980 2224
rect 2972 2116 2980 2124
rect 2972 2076 2980 2084
rect 2940 2056 2948 2064
rect 2956 2056 2964 2064
rect 2924 2016 2932 2024
rect 2940 1976 2948 1984
rect 2876 1956 2884 1964
rect 3148 2556 3156 2564
rect 3228 2556 3236 2564
rect 3292 2556 3300 2564
rect 3052 2496 3060 2504
rect 3052 2476 3060 2484
rect 3084 2476 3092 2484
rect 3100 2476 3108 2484
rect 3020 2396 3028 2404
rect 3196 2496 3204 2504
rect 3212 2496 3220 2504
rect 3244 2496 3252 2504
rect 3324 2496 3332 2504
rect 3132 2476 3140 2484
rect 3548 2576 3556 2584
rect 3692 2596 3700 2604
rect 3612 2576 3620 2584
rect 3644 2576 3652 2584
rect 3724 2636 3732 2644
rect 3740 2576 3748 2584
rect 3452 2516 3460 2524
rect 3484 2516 3492 2524
rect 3500 2516 3508 2524
rect 3532 2516 3540 2524
rect 3548 2516 3556 2524
rect 3564 2516 3572 2524
rect 3628 2516 3636 2524
rect 3660 2516 3668 2524
rect 3740 2516 3748 2524
rect 3404 2496 3412 2504
rect 3420 2496 3428 2504
rect 3468 2496 3476 2504
rect 3564 2496 3572 2504
rect 3580 2496 3588 2504
rect 3148 2436 3156 2444
rect 3196 2436 3204 2444
rect 3292 2436 3300 2444
rect 3324 2436 3332 2444
rect 3372 2436 3380 2444
rect 3244 2416 3252 2424
rect 3276 2416 3284 2424
rect 3244 2376 3252 2384
rect 3164 2356 3172 2364
rect 3100 2336 3108 2344
rect 3036 2316 3044 2324
rect 3020 2296 3028 2304
rect 3084 2296 3092 2304
rect 3148 2296 3156 2304
rect 3036 2276 3044 2284
rect 3132 2276 3140 2284
rect 3228 2296 3236 2304
rect 3212 2256 3220 2264
rect 3116 2236 3124 2244
rect 3004 2216 3012 2224
rect 3068 2216 3076 2224
rect 3260 2236 3268 2244
rect 3148 2176 3156 2184
rect 3292 2396 3300 2404
rect 3372 2336 3380 2344
rect 3324 2296 3332 2304
rect 3356 2296 3364 2304
rect 3436 2376 3444 2384
rect 3404 2256 3412 2264
rect 3324 2236 3332 2244
rect 3388 2236 3396 2244
rect 3308 2216 3316 2224
rect 3356 2216 3364 2224
rect 3388 2216 3396 2224
rect 3292 2176 3300 2184
rect 3340 2176 3348 2184
rect 3356 2176 3364 2184
rect 3004 2116 3012 2124
rect 3020 2116 3028 2124
rect 3068 2116 3076 2124
rect 3100 2116 3108 2124
rect 3116 2116 3124 2124
rect 3036 2016 3044 2024
rect 3052 2016 3060 2024
rect 2796 1896 2804 1904
rect 2780 1796 2788 1804
rect 2940 1916 2948 1924
rect 2828 1796 2836 1804
rect 2860 1896 2868 1904
rect 2908 1896 2916 1904
rect 2956 1896 2964 1904
rect 2860 1816 2868 1824
rect 2892 1816 2900 1824
rect 2908 1816 2916 1824
rect 2956 1816 2964 1824
rect 3004 1956 3012 1964
rect 3052 1956 3060 1964
rect 3004 1916 3012 1924
rect 3052 1896 3060 1904
rect 3420 2196 3428 2204
rect 3404 2176 3412 2184
rect 3500 2336 3508 2344
rect 3516 2336 3524 2344
rect 3548 2296 3556 2304
rect 3468 2236 3476 2244
rect 3484 2236 3492 2244
rect 3452 2156 3460 2164
rect 3516 2156 3524 2164
rect 3196 2136 3204 2144
rect 3228 2136 3236 2144
rect 3244 2136 3252 2144
rect 3148 2116 3156 2124
rect 3292 2116 3300 2124
rect 3436 2116 3444 2124
rect 3468 2116 3476 2124
rect 3484 2116 3492 2124
rect 3244 2096 3252 2104
rect 3276 2096 3284 2104
rect 3388 2096 3396 2104
rect 3132 2016 3140 2024
rect 3148 1976 3156 1984
rect 3132 1956 3140 1964
rect 2988 1816 2996 1824
rect 3020 1816 3028 1824
rect 3036 1816 3044 1824
rect 2924 1796 2932 1804
rect 2956 1796 2964 1804
rect 2972 1796 2980 1804
rect 2988 1796 2996 1804
rect 2684 1716 2692 1724
rect 2700 1716 2708 1724
rect 2748 1716 2756 1724
rect 2780 1716 2788 1724
rect 2940 1776 2948 1784
rect 3004 1776 3012 1784
rect 2908 1716 2916 1724
rect 2876 1696 2884 1704
rect 2892 1696 2900 1704
rect 2956 1716 2964 1724
rect 3276 2016 3284 2024
rect 3308 2016 3316 2024
rect 3212 1956 3220 1964
rect 3244 1956 3252 1964
rect 3180 1896 3188 1904
rect 3228 1896 3236 1904
rect 3340 2036 3348 2044
rect 3324 1976 3332 1984
rect 3084 1776 3092 1784
rect 3100 1776 3108 1784
rect 3004 1716 3012 1724
rect 3020 1716 3028 1724
rect 2988 1696 2996 1704
rect 3052 1696 3060 1704
rect 3036 1656 3044 1664
rect 2924 1616 2932 1624
rect 2972 1616 2980 1624
rect 2988 1616 2996 1624
rect 3068 1616 3076 1624
rect 2668 1576 2676 1584
rect 2700 1576 2708 1584
rect 2588 1496 2596 1504
rect 2652 1496 2660 1504
rect 2412 1396 2420 1404
rect 2444 1396 2452 1404
rect 2476 1436 2484 1444
rect 2524 1436 2532 1444
rect 2380 1336 2388 1344
rect 2396 1336 2404 1344
rect 2412 1336 2420 1344
rect 2348 1236 2356 1244
rect 2316 1216 2324 1224
rect 2348 1096 2356 1104
rect 2748 1596 2756 1604
rect 2844 1596 2852 1604
rect 2860 1596 2868 1604
rect 3084 1596 3092 1604
rect 2764 1576 2772 1584
rect 2924 1576 2932 1584
rect 2988 1576 2996 1584
rect 2732 1496 2740 1504
rect 2540 1416 2548 1424
rect 2588 1416 2596 1424
rect 2620 1416 2628 1424
rect 2508 1396 2516 1404
rect 2572 1376 2580 1384
rect 2588 1376 2596 1384
rect 2604 1376 2612 1384
rect 2492 1336 2500 1344
rect 2524 1336 2532 1344
rect 2444 1296 2452 1304
rect 2476 1296 2484 1304
rect 2524 1296 2532 1304
rect 2476 1236 2484 1244
rect 2524 1236 2532 1244
rect 2412 1216 2420 1224
rect 2460 1216 2468 1224
rect 2492 1216 2500 1224
rect 2588 1336 2596 1344
rect 2652 1376 2660 1384
rect 2700 1416 2708 1424
rect 2716 1416 2724 1424
rect 2748 1416 2756 1424
rect 2652 1356 2660 1364
rect 2668 1356 2676 1364
rect 2684 1356 2692 1364
rect 2780 1496 2788 1504
rect 2828 1496 2836 1504
rect 2812 1416 2820 1424
rect 3100 1536 3108 1544
rect 2860 1496 2868 1504
rect 2876 1496 2884 1504
rect 2940 1496 2948 1504
rect 3020 1496 3028 1504
rect 2860 1416 2868 1424
rect 2892 1416 2900 1424
rect 2956 1436 2964 1444
rect 3004 1396 3012 1404
rect 2812 1356 2820 1364
rect 2668 1336 2676 1344
rect 2684 1336 2692 1344
rect 2764 1336 2772 1344
rect 2844 1336 2852 1344
rect 2652 1296 2660 1304
rect 2636 1216 2644 1224
rect 2556 1176 2564 1184
rect 2588 1176 2596 1184
rect 2508 1156 2516 1164
rect 2844 1276 2852 1284
rect 2924 1376 2932 1384
rect 2972 1376 2980 1384
rect 3100 1416 3108 1424
rect 3020 1376 3028 1384
rect 3068 1376 3076 1384
rect 3084 1376 3092 1384
rect 2876 1356 2884 1364
rect 2892 1336 2900 1344
rect 2940 1336 2948 1344
rect 2972 1336 2980 1344
rect 2988 1336 2996 1344
rect 3052 1336 3060 1344
rect 2860 1256 2868 1264
rect 3084 1336 3092 1344
rect 2988 1296 2996 1304
rect 3036 1296 3044 1304
rect 2828 1236 2836 1244
rect 2956 1236 2964 1244
rect 3036 1236 3044 1244
rect 2748 1216 2756 1224
rect 2700 1196 2708 1204
rect 2668 1176 2676 1184
rect 2556 1136 2564 1144
rect 2396 1096 2404 1104
rect 2572 1116 2580 1124
rect 2588 1116 2596 1124
rect 2620 1096 2628 1104
rect 2460 1076 2468 1084
rect 2332 1056 2340 1064
rect 2364 1056 2372 1064
rect 2332 1016 2340 1024
rect 2348 1016 2356 1024
rect 2380 1016 2388 1024
rect 2364 956 2372 964
rect 2396 956 2404 964
rect 2220 896 2228 904
rect 2508 1036 2516 1044
rect 2460 996 2468 1004
rect 2476 996 2484 1004
rect 2540 1036 2548 1044
rect 2588 1036 2596 1044
rect 2524 1016 2532 1024
rect 2540 1016 2548 1024
rect 2460 976 2468 984
rect 2588 956 2596 964
rect 2412 936 2420 944
rect 2428 936 2436 944
rect 2444 936 2452 944
rect 2492 936 2500 944
rect 2524 936 2532 944
rect 2572 936 2580 944
rect 2316 916 2324 924
rect 2268 896 2276 904
rect 2284 896 2292 904
rect 2236 796 2244 804
rect 2268 816 2276 824
rect 2220 756 2228 764
rect 2252 756 2260 764
rect 2172 736 2180 744
rect 2380 876 2388 884
rect 2444 916 2452 924
rect 2684 1116 2692 1124
rect 2668 1096 2676 1104
rect 2700 1096 2708 1104
rect 2732 1096 2740 1104
rect 2700 1036 2708 1044
rect 2716 1036 2724 1044
rect 2780 1016 2788 1024
rect 3020 1216 3028 1224
rect 3020 1176 3028 1184
rect 3036 1176 3044 1184
rect 3004 1156 3012 1164
rect 2924 1136 2932 1144
rect 2860 1116 2868 1124
rect 2924 1116 2932 1124
rect 2876 1096 2884 1104
rect 2988 1076 2996 1084
rect 2828 1056 2836 1064
rect 2860 1056 2868 1064
rect 2876 1036 2884 1044
rect 2812 1016 2820 1024
rect 2876 1016 2884 1024
rect 2684 956 2692 964
rect 2700 956 2708 964
rect 2652 936 2660 944
rect 2668 936 2676 944
rect 2716 936 2724 944
rect 2764 936 2772 944
rect 2396 796 2404 804
rect 2412 796 2420 804
rect 2332 776 2340 784
rect 2268 736 2276 744
rect 2364 736 2372 744
rect 2396 736 2404 744
rect 2476 736 2484 744
rect 2508 736 2516 744
rect 2748 916 2756 924
rect 2796 996 2804 1004
rect 2892 996 2900 1004
rect 2860 976 2868 984
rect 2956 1056 2964 1064
rect 3020 1056 3028 1064
rect 3052 1036 3060 1044
rect 2908 976 2916 984
rect 2924 976 2932 984
rect 2908 956 2916 964
rect 2796 936 2804 944
rect 2764 896 2772 904
rect 2780 896 2788 904
rect 2924 936 2932 944
rect 2940 936 2948 944
rect 2972 936 2980 944
rect 2844 916 2852 924
rect 2844 896 2852 904
rect 2860 896 2868 904
rect 2812 856 2820 864
rect 2812 816 2820 824
rect 2556 736 2564 744
rect 2572 736 2580 744
rect 2412 716 2420 724
rect 2476 716 2484 724
rect 2540 716 2548 724
rect 2252 676 2260 684
rect 2268 676 2276 684
rect 2332 676 2340 684
rect 2428 676 2436 684
rect 2460 676 2468 684
rect 2524 676 2532 684
rect 2668 756 2676 764
rect 2652 736 2660 744
rect 2572 676 2580 684
rect 2044 636 2052 644
rect 2108 636 2116 644
rect 2156 636 2164 644
rect 1980 616 1988 624
rect 2076 596 2084 604
rect 2092 596 2100 604
rect 1980 576 1988 584
rect 2012 576 2020 584
rect 2060 576 2068 584
rect 1804 556 1812 564
rect 1884 556 1892 564
rect 1932 556 1940 564
rect 1948 556 1956 564
rect 1964 556 1972 564
rect 1868 536 1876 544
rect 1900 496 1908 504
rect 1820 456 1828 464
rect 2028 556 2036 564
rect 2044 556 2052 564
rect 2060 556 2068 564
rect 2028 496 2036 504
rect 2092 496 2100 504
rect 2156 596 2164 604
rect 2188 636 2196 644
rect 2188 616 2196 624
rect 2220 636 2228 644
rect 2284 636 2292 644
rect 2252 616 2260 624
rect 2300 616 2308 624
rect 2316 616 2324 624
rect 2364 616 2372 624
rect 2252 576 2260 584
rect 2396 616 2404 624
rect 2284 556 2292 564
rect 2332 556 2340 564
rect 2364 556 2372 564
rect 2124 496 2132 504
rect 2476 616 2484 624
rect 2412 596 2420 604
rect 2412 556 2420 564
rect 2508 616 2516 624
rect 2540 596 2548 604
rect 2572 596 2580 604
rect 2508 556 2516 564
rect 2524 556 2532 564
rect 2572 556 2580 564
rect 2604 556 2612 564
rect 2492 516 2500 524
rect 2540 516 2548 524
rect 2236 456 2244 464
rect 2300 456 2308 464
rect 1996 436 2004 444
rect 2044 436 2052 444
rect 2188 436 2196 444
rect 2204 436 2212 444
rect 2268 436 2276 444
rect 2044 396 2052 404
rect 2060 396 2068 404
rect 2028 376 2036 384
rect 1724 336 1732 344
rect 1788 336 1796 344
rect 1852 336 1860 344
rect 1884 336 1892 344
rect 1900 336 1908 344
rect 1932 336 1940 344
rect 2076 336 2084 344
rect 1916 316 1924 324
rect 1660 236 1668 244
rect 1612 176 1620 184
rect 1708 236 1716 244
rect 1692 216 1700 224
rect 1644 156 1652 164
rect 1692 156 1700 164
rect 1724 216 1732 224
rect 1756 216 1764 224
rect 1836 236 1844 244
rect 1868 236 1876 244
rect 1900 236 1908 244
rect 1804 216 1812 224
rect 1772 176 1780 184
rect 1788 176 1796 184
rect 1756 156 1764 164
rect 1596 136 1604 144
rect 1660 116 1668 124
rect 1708 116 1716 124
rect 1804 96 1812 104
rect 476 76 484 84
rect 652 76 660 84
rect 668 76 676 84
rect 780 76 788 84
rect 812 76 820 84
rect 924 76 932 84
rect 1260 76 1268 84
rect 1740 76 1748 84
rect 1868 216 1876 224
rect 2748 736 2756 744
rect 2716 716 2724 724
rect 2780 716 2788 724
rect 2764 696 2772 704
rect 3228 1836 3236 1844
rect 3260 1836 3268 1844
rect 3292 1836 3300 1844
rect 3164 1816 3172 1824
rect 3372 1836 3380 1844
rect 3404 1836 3412 1844
rect 3356 1816 3364 1824
rect 3724 2476 3732 2484
rect 3724 2336 3732 2344
rect 3580 2316 3588 2324
rect 3628 2316 3636 2324
rect 3692 2316 3700 2324
rect 3740 2316 3748 2324
rect 4284 3336 4292 3344
rect 4380 3356 4388 3364
rect 4396 3356 4404 3364
rect 4396 3336 4404 3344
rect 4316 3316 4324 3324
rect 4364 3316 4372 3324
rect 4188 3296 4196 3304
rect 4252 3296 4260 3304
rect 4316 3296 4324 3304
rect 4300 3156 4308 3164
rect 4316 3136 4324 3144
rect 4300 3116 4308 3124
rect 4140 3096 4148 3104
rect 4204 3096 4212 3104
rect 4124 3076 4132 3084
rect 3996 3056 4004 3064
rect 3868 3036 3876 3044
rect 3980 3036 3988 3044
rect 4060 3036 4068 3044
rect 3804 2976 3812 2984
rect 3788 2956 3796 2964
rect 4172 3016 4180 3024
rect 4044 2996 4052 3004
rect 4060 2996 4068 3004
rect 4108 2996 4116 3004
rect 4124 2996 4132 3004
rect 3900 2956 3908 2964
rect 3836 2896 3844 2904
rect 4060 2936 4068 2944
rect 4092 2936 4100 2944
rect 3932 2916 3940 2924
rect 4012 2916 4020 2924
rect 4028 2916 4036 2924
rect 3868 2896 3876 2904
rect 3884 2896 3892 2904
rect 3852 2876 3860 2884
rect 3900 2796 3908 2804
rect 3836 2776 3844 2784
rect 3980 2776 3988 2784
rect 3964 2736 3972 2744
rect 3916 2716 3924 2724
rect 3868 2696 3876 2704
rect 3884 2696 3892 2704
rect 4012 2756 4020 2764
rect 4044 2756 4052 2764
rect 4060 2716 4068 2724
rect 3836 2636 3844 2644
rect 3788 2556 3796 2564
rect 3868 2596 3876 2604
rect 3932 2556 3940 2564
rect 3916 2516 3924 2524
rect 3948 2516 3956 2524
rect 3820 2496 3828 2504
rect 3804 2476 3812 2484
rect 3868 2476 3876 2484
rect 3884 2476 3892 2484
rect 3804 2416 3812 2424
rect 3868 2416 3876 2424
rect 3996 2616 4004 2624
rect 4044 2616 4052 2624
rect 4060 2616 4068 2624
rect 4028 2596 4036 2604
rect 4044 2596 4052 2604
rect 4012 2576 4020 2584
rect 4124 2896 4132 2904
rect 4156 2896 4164 2904
rect 4140 2876 4148 2884
rect 4172 2856 4180 2864
rect 4140 2836 4148 2844
rect 4108 2756 4116 2764
rect 4092 2716 4100 2724
rect 4124 2736 4132 2744
rect 4172 2756 4180 2764
rect 4188 2756 4196 2764
rect 4140 2716 4148 2724
rect 4156 2676 4164 2684
rect 4492 3436 4500 3444
rect 4508 3436 4516 3444
rect 4572 3436 4580 3444
rect 4524 3416 4532 3424
rect 4476 3376 4484 3384
rect 4508 3356 4516 3364
rect 4460 3316 4468 3324
rect 4508 3336 4516 3344
rect 4508 3316 4516 3324
rect 4668 3456 4676 3464
rect 4684 3436 4692 3444
rect 4844 3516 4852 3524
rect 4956 3516 4964 3524
rect 4812 3496 4820 3504
rect 4828 3496 4836 3504
rect 5052 3556 5060 3564
rect 4988 3496 4996 3504
rect 5084 3496 5092 3504
rect 4860 3476 4868 3484
rect 4892 3476 4900 3484
rect 5004 3476 5012 3484
rect 5036 3476 5044 3484
rect 5132 3476 5140 3484
rect 4732 3436 4740 3444
rect 4956 3456 4964 3464
rect 4828 3436 4836 3444
rect 4892 3436 4900 3444
rect 4940 3436 4948 3444
rect 4780 3416 4788 3424
rect 4764 3376 4772 3384
rect 4700 3356 4708 3364
rect 4748 3356 4756 3364
rect 4556 3296 4564 3304
rect 4924 3416 4932 3424
rect 4988 3376 4996 3384
rect 5052 3376 5060 3384
rect 4844 3356 4852 3364
rect 4876 3356 4884 3364
rect 4940 3356 4948 3364
rect 5020 3356 5028 3364
rect 4828 3336 4836 3344
rect 4684 3316 4692 3324
rect 4732 3316 4740 3324
rect 4796 3316 4804 3324
rect 4924 3316 4932 3324
rect 4652 3296 4660 3304
rect 4412 3276 4420 3284
rect 4492 3276 4500 3284
rect 4636 3276 4644 3284
rect 4604 3236 4612 3244
rect 4652 3236 4660 3244
rect 4668 3236 4676 3244
rect 4876 3236 4884 3244
rect 4588 3216 4596 3224
rect 4524 3196 4532 3204
rect 4732 3196 4740 3204
rect 4556 3176 4564 3184
rect 4828 3176 4836 3184
rect 4396 3156 4404 3164
rect 4364 3136 4372 3144
rect 4700 3136 4708 3144
rect 4796 3136 4804 3144
rect 4892 3136 4900 3144
rect 4428 3116 4436 3124
rect 4556 3116 4564 3124
rect 4684 3116 4692 3124
rect 4396 3096 4404 3104
rect 4444 3096 4452 3104
rect 4508 3096 4516 3104
rect 4588 3096 4596 3104
rect 4636 3096 4644 3104
rect 4252 3076 4260 3084
rect 4348 3076 4356 3084
rect 4220 3036 4228 3044
rect 4604 3076 4612 3084
rect 4716 3116 4724 3124
rect 4748 3116 4756 3124
rect 4476 3056 4484 3064
rect 4700 3056 4708 3064
rect 5164 3436 5172 3444
rect 5116 3396 5124 3404
rect 5100 3376 5108 3384
rect 5132 3356 5140 3364
rect 5100 3336 5108 3344
rect 5164 3336 5172 3344
rect 5020 3316 5028 3324
rect 5068 3316 5076 3324
rect 4972 3296 4980 3304
rect 5180 3296 5188 3304
rect 4972 3276 4980 3284
rect 4988 3276 4996 3284
rect 5052 3276 5060 3284
rect 4956 3236 4964 3244
rect 5004 3256 5012 3264
rect 4940 3156 4948 3164
rect 4844 3116 4852 3124
rect 4908 3116 4916 3124
rect 4924 3116 4932 3124
rect 4988 3156 4996 3164
rect 4940 3096 4948 3104
rect 4732 3076 4740 3084
rect 4796 3056 4804 3064
rect 4892 3056 4900 3064
rect 4940 3056 4948 3064
rect 4956 3056 4964 3064
rect 4300 3036 4308 3044
rect 4332 3036 4340 3044
rect 4284 3016 4292 3024
rect 4348 3016 4356 3024
rect 4268 2996 4276 3004
rect 4412 2996 4420 3004
rect 4380 2956 4388 2964
rect 4220 2936 4228 2944
rect 4252 2936 4260 2944
rect 4252 2916 4260 2924
rect 4348 2916 4356 2924
rect 4364 2916 4372 2924
rect 4300 2896 4308 2904
rect 4428 2896 4436 2904
rect 4236 2816 4244 2824
rect 4316 2816 4324 2824
rect 4124 2596 4132 2604
rect 4172 2596 4180 2604
rect 4076 2576 4084 2584
rect 4060 2556 4068 2564
rect 4076 2556 4084 2564
rect 4108 2556 4116 2564
rect 4156 2556 4164 2564
rect 4060 2516 4068 2524
rect 4396 2796 4404 2804
rect 4348 2756 4356 2764
rect 4412 2756 4420 2764
rect 4556 3036 4564 3044
rect 4604 3036 4612 3044
rect 4668 3036 4676 3044
rect 4780 3036 4788 3044
rect 4716 3016 4724 3024
rect 4492 2996 4500 3004
rect 4572 2996 4580 3004
rect 4492 2916 4500 2924
rect 4524 2916 4532 2924
rect 4556 2916 4564 2924
rect 4444 2876 4452 2884
rect 4476 2876 4484 2884
rect 4652 2876 4660 2884
rect 4828 3036 4836 3044
rect 4876 3036 4884 3044
rect 4892 3016 4900 3024
rect 4700 2936 4708 2944
rect 4716 2936 4724 2944
rect 4764 2936 4772 2944
rect 4812 2936 4820 2944
rect 4860 2936 4868 2944
rect 4684 2896 4692 2904
rect 4732 2896 4740 2904
rect 4748 2896 4756 2904
rect 4812 2876 4820 2884
rect 4812 2856 4820 2864
rect 4668 2816 4676 2824
rect 4620 2776 4628 2784
rect 4508 2756 4516 2764
rect 4764 2736 4772 2744
rect 4828 2736 4836 2744
rect 4252 2676 4260 2684
rect 4540 2696 4548 2704
rect 4668 2696 4676 2704
rect 4716 2696 4724 2704
rect 4764 2696 4772 2704
rect 4780 2696 4788 2704
rect 4876 2696 4884 2704
rect 4300 2676 4308 2684
rect 4316 2676 4324 2684
rect 4364 2676 4372 2684
rect 4380 2676 4388 2684
rect 4492 2676 4500 2684
rect 4604 2676 4612 2684
rect 4636 2676 4644 2684
rect 4204 2616 4212 2624
rect 4252 2616 4260 2624
rect 4252 2556 4260 2564
rect 4204 2536 4212 2544
rect 4124 2516 4132 2524
rect 4172 2516 4180 2524
rect 4188 2516 4196 2524
rect 4236 2516 4244 2524
rect 4012 2496 4020 2504
rect 4092 2496 4100 2504
rect 4124 2496 4132 2504
rect 3980 2456 3988 2464
rect 3916 2316 3924 2324
rect 4236 2496 4244 2504
rect 4076 2436 4084 2444
rect 3996 2416 4004 2424
rect 4028 2416 4036 2424
rect 4076 2416 4084 2424
rect 4060 2376 4068 2384
rect 3996 2336 4004 2344
rect 4140 2336 4148 2344
rect 4092 2316 4100 2324
rect 4124 2316 4132 2324
rect 4316 2596 4324 2604
rect 4300 2576 4308 2584
rect 4428 2616 4436 2624
rect 4444 2616 4452 2624
rect 4684 2636 4692 2644
rect 4492 2596 4500 2604
rect 4572 2596 4580 2604
rect 4348 2576 4356 2584
rect 4364 2576 4372 2584
rect 4604 2576 4612 2584
rect 4332 2516 4340 2524
rect 4284 2496 4292 2504
rect 4396 2476 4404 2484
rect 4268 2416 4276 2424
rect 4332 2416 4340 2424
rect 4252 2396 4260 2404
rect 4252 2336 4260 2344
rect 4316 2336 4324 2344
rect 3580 2276 3588 2284
rect 3676 2276 3684 2284
rect 3740 2276 3748 2284
rect 3772 2276 3780 2284
rect 3836 2276 3844 2284
rect 3884 2276 3892 2284
rect 3932 2276 3940 2284
rect 3804 2256 3812 2264
rect 3948 2256 3956 2264
rect 3564 2236 3572 2244
rect 3580 2236 3588 2244
rect 3772 2236 3780 2244
rect 3564 2216 3572 2224
rect 3644 2216 3652 2224
rect 3660 2216 3668 2224
rect 3772 2216 3780 2224
rect 3788 2216 3796 2224
rect 3548 2156 3556 2164
rect 3740 2156 3748 2164
rect 3756 2156 3764 2164
rect 3548 2116 3556 2124
rect 3596 2116 3604 2124
rect 3708 2116 3716 2124
rect 3500 2096 3508 2104
rect 3532 2096 3540 2104
rect 3660 2096 3668 2104
rect 3468 2036 3476 2044
rect 3436 2016 3444 2024
rect 3532 2016 3540 2024
rect 3468 1976 3476 1984
rect 3452 1936 3460 1944
rect 3644 2036 3652 2044
rect 3660 2036 3668 2044
rect 3708 2036 3716 2044
rect 3724 2036 3732 2044
rect 3596 2016 3604 2024
rect 3740 2016 3748 2024
rect 3564 1976 3572 1984
rect 3612 1976 3620 1984
rect 3628 1976 3636 1984
rect 3676 1976 3684 1984
rect 3548 1916 3556 1924
rect 3468 1896 3476 1904
rect 3484 1896 3492 1904
rect 3580 1896 3588 1904
rect 3596 1896 3604 1904
rect 3644 1896 3652 1904
rect 3916 2216 3924 2224
rect 3948 2216 3956 2224
rect 3884 2056 3892 2064
rect 4236 2296 4244 2304
rect 4028 2276 4036 2284
rect 4156 2276 4164 2284
rect 4220 2276 4228 2284
rect 3980 2256 3988 2264
rect 4076 2256 4084 2264
rect 4076 2236 4084 2244
rect 4172 2236 4180 2244
rect 4044 2216 4052 2224
rect 4060 2176 4068 2184
rect 4012 2156 4020 2164
rect 4044 2156 4052 2164
rect 3980 2056 3988 2064
rect 3996 2056 4004 2064
rect 3868 2016 3876 2024
rect 3932 2016 3940 2024
rect 4188 2216 4196 2224
rect 4092 2196 4100 2204
rect 4220 2196 4228 2204
rect 4652 2556 4660 2564
rect 4732 2576 4740 2584
rect 4876 2656 4884 2664
rect 4796 2556 4804 2564
rect 4908 2996 4916 3004
rect 4940 2976 4948 2984
rect 4988 3036 4996 3044
rect 4908 2956 4916 2964
rect 4940 2956 4948 2964
rect 5132 3236 5140 3244
rect 5036 3216 5044 3224
rect 5036 3176 5044 3184
rect 5068 3176 5076 3184
rect 5020 3076 5028 3084
rect 5164 3116 5172 3124
rect 5084 3056 5092 3064
rect 5116 3036 5124 3044
rect 5052 2976 5060 2984
rect 5052 2956 5060 2964
rect 5100 2956 5108 2964
rect 5020 2916 5028 2924
rect 5084 2916 5092 2924
rect 5100 2916 5108 2924
rect 4908 2736 4916 2744
rect 4908 2696 4916 2704
rect 5004 2816 5012 2824
rect 5132 2896 5140 2904
rect 5132 2876 5140 2884
rect 5116 2856 5124 2864
rect 5068 2736 5076 2744
rect 4972 2716 4980 2724
rect 5100 2716 5108 2724
rect 4956 2676 4964 2684
rect 4972 2676 4980 2684
rect 5052 2676 5060 2684
rect 5100 2676 5108 2684
rect 5004 2656 5012 2664
rect 5068 2656 5076 2664
rect 4924 2636 4932 2644
rect 4956 2636 4964 2644
rect 5100 2636 5108 2644
rect 5020 2616 5028 2624
rect 4892 2596 4900 2604
rect 5004 2596 5012 2604
rect 5116 2596 5124 2604
rect 5084 2556 5092 2564
rect 5100 2556 5108 2564
rect 5164 2816 5172 2824
rect 5164 2796 5172 2804
rect 5180 2796 5188 2804
rect 5148 2756 5156 2764
rect 5148 2736 5156 2744
rect 5196 2616 5204 2624
rect 5148 2576 5156 2584
rect 4444 2516 4452 2524
rect 4460 2516 4468 2524
rect 4492 2516 4500 2524
rect 4524 2516 4532 2524
rect 4588 2516 4596 2524
rect 4716 2516 4724 2524
rect 4476 2496 4484 2504
rect 4508 2496 4516 2504
rect 4604 2496 4612 2504
rect 4556 2476 4564 2484
rect 4508 2436 4516 2444
rect 4428 2336 4436 2344
rect 4524 2316 4532 2324
rect 4268 2276 4276 2284
rect 4412 2276 4420 2284
rect 4476 2276 4484 2284
rect 4700 2496 4708 2504
rect 4700 2476 4708 2484
rect 4716 2456 4724 2464
rect 4764 2516 4772 2524
rect 4892 2516 4900 2524
rect 4940 2516 4948 2524
rect 4748 2496 4756 2504
rect 4796 2496 4804 2504
rect 4908 2496 4916 2504
rect 4956 2496 4964 2504
rect 5052 2536 5060 2544
rect 5036 2516 5044 2524
rect 4812 2476 4820 2484
rect 4828 2436 4836 2444
rect 5132 2496 5140 2504
rect 5180 2496 5188 2504
rect 4972 2476 4980 2484
rect 5068 2476 5076 2484
rect 4700 2356 4708 2364
rect 4652 2316 4660 2324
rect 4556 2276 4564 2284
rect 4588 2276 4596 2284
rect 4620 2276 4628 2284
rect 4636 2276 4644 2284
rect 4268 2256 4276 2264
rect 4364 2236 4372 2244
rect 4380 2216 4388 2224
rect 4412 2216 4420 2224
rect 4476 2216 4484 2224
rect 4652 2256 4660 2264
rect 4684 2256 4692 2264
rect 4332 2176 4340 2184
rect 4076 2096 4084 2104
rect 4108 2156 4116 2164
rect 4124 2156 4132 2164
rect 4204 2156 4212 2164
rect 4236 2156 4244 2164
rect 4268 2156 4276 2164
rect 4316 2156 4324 2164
rect 4284 2136 4292 2144
rect 4204 2116 4212 2124
rect 4236 2116 4244 2124
rect 4380 2196 4388 2204
rect 4412 2196 4420 2204
rect 4444 2196 4452 2204
rect 4348 2116 4356 2124
rect 4156 2096 4164 2104
rect 4172 2096 4180 2104
rect 4092 2056 4100 2064
rect 4060 2036 4068 2044
rect 4092 2036 4100 2044
rect 4060 1996 4068 2004
rect 3980 1976 3988 1984
rect 4028 1976 4036 1984
rect 3788 1956 3796 1964
rect 3932 1956 3940 1964
rect 4076 1956 4084 1964
rect 3532 1876 3540 1884
rect 3564 1876 3572 1884
rect 3484 1856 3492 1864
rect 3468 1836 3476 1844
rect 3148 1796 3156 1804
rect 3212 1796 3220 1804
rect 3324 1796 3332 1804
rect 3356 1796 3364 1804
rect 3420 1796 3428 1804
rect 3180 1736 3188 1744
rect 3164 1716 3172 1724
rect 3260 1716 3268 1724
rect 3340 1716 3348 1724
rect 3212 1696 3220 1704
rect 3228 1696 3236 1704
rect 3308 1696 3316 1704
rect 3324 1696 3332 1704
rect 3404 1676 3412 1684
rect 3452 1756 3460 1764
rect 3500 1836 3508 1844
rect 3516 1836 3524 1844
rect 3500 1776 3508 1784
rect 3676 1856 3684 1864
rect 3740 1836 3748 1844
rect 4012 1916 4020 1924
rect 4204 1956 4212 1964
rect 4252 1936 4260 1944
rect 3788 1856 3796 1864
rect 3868 1856 3876 1864
rect 3596 1816 3604 1824
rect 3772 1816 3780 1824
rect 3548 1776 3556 1784
rect 3500 1756 3508 1764
rect 3532 1756 3540 1764
rect 3580 1756 3588 1764
rect 3756 1776 3764 1784
rect 4220 1896 4228 1904
rect 4524 2196 4532 2204
rect 4588 2196 4596 2204
rect 4636 2216 4644 2224
rect 4604 2156 4612 2164
rect 4428 2116 4436 2124
rect 4460 2116 4468 2124
rect 4508 2116 4516 2124
rect 4540 2116 4548 2124
rect 4588 2116 4596 2124
rect 4636 2116 4644 2124
rect 4700 2156 4708 2164
rect 4492 2076 4500 2084
rect 4444 2036 4452 2044
rect 4508 2016 4516 2024
rect 4412 1976 4420 1984
rect 4284 1956 4292 1964
rect 4348 1956 4356 1964
rect 3948 1796 3956 1804
rect 3932 1776 3940 1784
rect 3964 1776 3972 1784
rect 3628 1756 3636 1764
rect 3660 1736 3668 1744
rect 3676 1736 3684 1744
rect 3708 1736 3716 1744
rect 3724 1736 3732 1744
rect 3740 1736 3748 1744
rect 3756 1736 3764 1744
rect 3788 1736 3796 1744
rect 3436 1696 3444 1704
rect 3484 1696 3492 1704
rect 3500 1696 3508 1704
rect 3692 1716 3700 1724
rect 3740 1716 3748 1724
rect 3772 1696 3780 1704
rect 3884 1756 3892 1764
rect 3916 1756 3924 1764
rect 3852 1736 3860 1744
rect 3868 1736 3876 1744
rect 3980 1736 3988 1744
rect 3836 1716 3844 1724
rect 3852 1696 3860 1704
rect 3916 1696 3924 1704
rect 3820 1636 3828 1644
rect 3244 1616 3252 1624
rect 3388 1616 3396 1624
rect 3516 1616 3524 1624
rect 3772 1616 3780 1624
rect 3788 1616 3796 1624
rect 3148 1576 3156 1584
rect 3484 1596 3492 1604
rect 3148 1536 3156 1544
rect 3228 1536 3236 1544
rect 3260 1536 3268 1544
rect 3276 1536 3284 1544
rect 3356 1536 3364 1544
rect 3372 1536 3380 1544
rect 3500 1536 3508 1544
rect 3308 1516 3316 1524
rect 3164 1416 3172 1424
rect 3196 1416 3204 1424
rect 3212 1416 3220 1424
rect 3276 1436 3284 1444
rect 3404 1516 3412 1524
rect 3468 1516 3476 1524
rect 3532 1596 3540 1604
rect 3692 1596 3700 1604
rect 3756 1596 3764 1604
rect 3308 1436 3316 1444
rect 3340 1436 3348 1444
rect 3404 1436 3412 1444
rect 3452 1436 3460 1444
rect 3468 1436 3476 1444
rect 3164 1396 3172 1404
rect 3180 1396 3188 1404
rect 3132 1376 3140 1384
rect 3260 1376 3268 1384
rect 3292 1376 3300 1384
rect 3404 1396 3412 1404
rect 3356 1376 3364 1384
rect 3356 1356 3364 1364
rect 3116 1216 3124 1224
rect 3484 1376 3492 1384
rect 3500 1356 3508 1364
rect 3228 1336 3236 1344
rect 3292 1336 3300 1344
rect 3212 1296 3220 1304
rect 3324 1296 3332 1304
rect 3388 1296 3396 1304
rect 3244 1236 3252 1244
rect 3372 1236 3380 1244
rect 3196 1216 3204 1224
rect 3276 1216 3284 1224
rect 3404 1196 3412 1204
rect 3276 1176 3284 1184
rect 3276 1136 3284 1144
rect 3324 1136 3332 1144
rect 3436 1296 3444 1304
rect 3452 1276 3460 1284
rect 3500 1276 3508 1284
rect 3420 1136 3428 1144
rect 3436 1136 3444 1144
rect 3516 1236 3524 1244
rect 3596 1576 3604 1584
rect 3548 1536 3556 1544
rect 3564 1476 3572 1484
rect 3660 1536 3668 1544
rect 3676 1536 3684 1544
rect 3628 1456 3636 1464
rect 3548 1436 3556 1444
rect 3580 1416 3588 1424
rect 3868 1616 3876 1624
rect 3868 1596 3876 1604
rect 3804 1456 3812 1464
rect 3644 1416 3652 1424
rect 3708 1416 3716 1424
rect 3596 1396 3604 1404
rect 3612 1396 3620 1404
rect 3580 1356 3588 1364
rect 3660 1376 3668 1384
rect 3740 1376 3748 1384
rect 3756 1376 3764 1384
rect 3724 1356 3732 1364
rect 3740 1356 3748 1364
rect 3772 1356 3780 1364
rect 3548 1296 3556 1304
rect 3580 1296 3588 1304
rect 3532 1216 3540 1224
rect 3676 1316 3684 1324
rect 3740 1316 3748 1324
rect 3772 1316 3780 1324
rect 3596 1256 3604 1264
rect 3644 1236 3652 1244
rect 3628 1196 3636 1204
rect 3676 1196 3684 1204
rect 3740 1236 3748 1244
rect 3836 1476 3844 1484
rect 3884 1416 3892 1424
rect 3836 1356 3844 1364
rect 3980 1696 3988 1704
rect 3996 1656 4004 1664
rect 4076 1856 4084 1864
rect 4108 1856 4116 1864
rect 4028 1796 4036 1804
rect 4076 1776 4084 1784
rect 4076 1756 4084 1764
rect 4124 1756 4132 1764
rect 4028 1736 4036 1744
rect 4060 1736 4068 1744
rect 4076 1736 4084 1744
rect 3964 1536 3972 1544
rect 3932 1516 3940 1524
rect 3964 1496 3972 1504
rect 4044 1636 4052 1644
rect 4044 1596 4052 1604
rect 4012 1516 4020 1524
rect 4028 1516 4036 1524
rect 4124 1696 4132 1704
rect 4172 1796 4180 1804
rect 4172 1736 4180 1744
rect 4220 1796 4228 1804
rect 4204 1716 4212 1724
rect 4156 1696 4164 1704
rect 4220 1696 4228 1704
rect 4204 1636 4212 1644
rect 4140 1596 4148 1604
rect 4172 1596 4180 1604
rect 4204 1596 4212 1604
rect 4060 1516 4068 1524
rect 4092 1516 4100 1524
rect 4140 1496 4148 1504
rect 4188 1496 4196 1504
rect 4092 1476 4100 1484
rect 4156 1476 4164 1484
rect 4076 1456 4084 1464
rect 4108 1456 4116 1464
rect 4140 1456 4148 1464
rect 4220 1456 4228 1464
rect 4236 1456 4244 1464
rect 3948 1416 3956 1424
rect 3980 1416 3988 1424
rect 3996 1416 4004 1424
rect 4028 1416 4036 1424
rect 4044 1416 4052 1424
rect 3900 1376 3908 1384
rect 3932 1356 3940 1364
rect 3836 1336 3844 1344
rect 3884 1336 3892 1344
rect 3868 1316 3876 1324
rect 3884 1316 3892 1324
rect 4028 1356 4036 1364
rect 4044 1356 4052 1364
rect 4060 1356 4068 1364
rect 4172 1416 4180 1424
rect 4300 1896 4308 1904
rect 4444 1976 4452 1984
rect 4540 1976 4548 1984
rect 4588 1976 4596 1984
rect 4556 1956 4564 1964
rect 4700 2096 4708 2104
rect 4684 2076 4692 2084
rect 4732 2416 4740 2424
rect 4748 2416 4756 2424
rect 4860 2416 4868 2424
rect 4812 2376 4820 2384
rect 4732 2336 4740 2344
rect 4796 2316 4804 2324
rect 4732 2276 4740 2284
rect 4940 2356 4948 2364
rect 5036 2356 5044 2364
rect 4924 2336 4932 2344
rect 5036 2336 5044 2344
rect 4860 2316 4868 2324
rect 4844 2296 4852 2304
rect 4828 2276 4836 2284
rect 4892 2276 4900 2284
rect 4796 2256 4804 2264
rect 4764 2236 4772 2244
rect 4780 2216 4788 2224
rect 4796 2216 4804 2224
rect 4764 2196 4772 2204
rect 4844 2196 4852 2204
rect 4780 2176 4788 2184
rect 4748 2156 4756 2164
rect 4748 2136 4756 2144
rect 4796 2136 4804 2144
rect 4828 2136 4836 2144
rect 4636 1936 4644 1944
rect 4652 1936 4660 1944
rect 4604 1916 4612 1924
rect 4620 1916 4628 1924
rect 4492 1896 4500 1904
rect 4844 2076 4852 2084
rect 4828 2056 4836 2064
rect 4780 2036 4788 2044
rect 4764 1976 4772 1984
rect 4748 1936 4756 1944
rect 4732 1916 4740 1924
rect 4876 2216 4884 2224
rect 4892 2196 4900 2204
rect 4924 2256 4932 2264
rect 5052 2296 5060 2304
rect 5084 2276 5092 2284
rect 4988 2256 4996 2264
rect 4972 2236 4980 2244
rect 4956 2216 4964 2224
rect 4972 2216 4980 2224
rect 5004 2196 5012 2204
rect 5052 2196 5060 2204
rect 4892 2136 4900 2144
rect 4940 2136 4948 2144
rect 5020 2136 5028 2144
rect 5052 2136 5060 2144
rect 4988 2116 4996 2124
rect 4892 2076 4900 2084
rect 5004 2076 5012 2084
rect 4972 1996 4980 2004
rect 4972 1896 4980 1904
rect 5180 2316 5188 2324
rect 5132 2296 5140 2304
rect 5132 2256 5140 2264
rect 5148 2256 5156 2264
rect 5148 2236 5156 2244
rect 5116 2216 5124 2224
rect 5100 2176 5108 2184
rect 5100 2156 5108 2164
rect 5068 2116 5076 2124
rect 5068 2016 5076 2024
rect 5116 2116 5124 2124
rect 5116 2076 5124 2084
rect 5116 2056 5124 2064
rect 5084 1996 5092 2004
rect 5084 1976 5092 1984
rect 5100 1956 5108 1964
rect 5100 1916 5108 1924
rect 4540 1876 4548 1884
rect 4668 1876 4676 1884
rect 4828 1876 4836 1884
rect 4860 1876 4868 1884
rect 5052 1876 5060 1884
rect 5084 1876 5092 1884
rect 4316 1856 4324 1864
rect 4444 1856 4452 1864
rect 4652 1856 4660 1864
rect 4364 1836 4372 1844
rect 4396 1836 4404 1844
rect 4476 1836 4484 1844
rect 4412 1816 4420 1824
rect 4348 1796 4356 1804
rect 4364 1776 4372 1784
rect 4268 1716 4276 1724
rect 4316 1756 4324 1764
rect 4444 1776 4452 1784
rect 4492 1776 4500 1784
rect 4460 1736 4468 1744
rect 4508 1716 4516 1724
rect 4300 1696 4308 1704
rect 4364 1696 4372 1704
rect 4348 1676 4356 1684
rect 4492 1696 4500 1704
rect 4412 1676 4420 1684
rect 4428 1676 4436 1684
rect 4396 1656 4404 1664
rect 4284 1636 4292 1644
rect 4332 1596 4340 1604
rect 4268 1536 4276 1544
rect 4316 1536 4324 1544
rect 4268 1516 4276 1524
rect 4460 1556 4468 1564
rect 4396 1536 4404 1544
rect 4476 1536 4484 1544
rect 4284 1456 4292 1464
rect 4492 1476 4500 1484
rect 4412 1436 4420 1444
rect 4252 1416 4260 1424
rect 4380 1416 4388 1424
rect 4572 1836 4580 1844
rect 4780 1836 4788 1844
rect 4684 1796 4692 1804
rect 4588 1776 4596 1784
rect 4684 1776 4692 1784
rect 4844 1836 4852 1844
rect 4940 1856 4948 1864
rect 4988 1856 4996 1864
rect 4892 1836 4900 1844
rect 4796 1776 4804 1784
rect 4828 1816 4836 1824
rect 4876 1816 4884 1824
rect 4588 1736 4596 1744
rect 4636 1736 4644 1744
rect 4700 1736 4708 1744
rect 4780 1736 4788 1744
rect 4652 1716 4660 1724
rect 4684 1716 4692 1724
rect 4924 1796 4932 1804
rect 4988 1756 4996 1764
rect 5020 1756 5028 1764
rect 4956 1736 4964 1744
rect 5020 1736 5028 1744
rect 4620 1596 4628 1604
rect 4588 1516 4596 1524
rect 4796 1656 4804 1664
rect 4748 1636 4756 1644
rect 4764 1596 4772 1604
rect 4732 1576 4740 1584
rect 4764 1576 4772 1584
rect 4540 1496 4548 1504
rect 4556 1496 4564 1504
rect 4604 1496 4612 1504
rect 4636 1496 4644 1504
rect 4556 1476 4564 1484
rect 4604 1476 4612 1484
rect 4652 1476 4660 1484
rect 4524 1416 4532 1424
rect 4460 1396 4468 1404
rect 4204 1356 4212 1364
rect 4700 1456 4708 1464
rect 4668 1416 4676 1424
rect 4748 1456 4756 1464
rect 4812 1576 4820 1584
rect 5036 1716 5044 1724
rect 5020 1696 5028 1704
rect 4956 1656 4964 1664
rect 4892 1616 4900 1624
rect 4892 1576 4900 1584
rect 4844 1536 4852 1544
rect 4828 1456 4836 1464
rect 4876 1536 4884 1544
rect 5068 1796 5076 1804
rect 5068 1716 5076 1724
rect 5164 2096 5172 2104
rect 5148 2056 5156 2064
rect 5132 1956 5140 1964
rect 5148 1956 5156 1964
rect 5148 1876 5156 1884
rect 5100 1776 5108 1784
rect 5116 1776 5124 1784
rect 5116 1756 5124 1764
rect 5132 1756 5140 1764
rect 5148 1756 5156 1764
rect 5100 1736 5108 1744
rect 5116 1736 5124 1744
rect 5084 1696 5092 1704
rect 5052 1656 5060 1664
rect 5068 1596 5076 1604
rect 5132 1716 5140 1724
rect 5164 1696 5172 1704
rect 5164 1556 5172 1564
rect 5036 1516 5044 1524
rect 4940 1476 4948 1484
rect 4988 1476 4996 1484
rect 4780 1436 4788 1444
rect 4684 1396 4692 1404
rect 4732 1376 4740 1384
rect 4876 1416 4884 1424
rect 4876 1396 4884 1404
rect 4268 1356 4276 1364
rect 4300 1356 4308 1364
rect 4364 1356 4372 1364
rect 4396 1356 4404 1364
rect 4444 1356 4452 1364
rect 4492 1356 4500 1364
rect 4604 1356 4612 1364
rect 4636 1356 4644 1364
rect 4700 1356 4708 1364
rect 4716 1356 4724 1364
rect 4828 1356 4836 1364
rect 4860 1356 4868 1364
rect 3964 1336 3972 1344
rect 3996 1336 4004 1344
rect 4076 1336 4084 1344
rect 4124 1336 4132 1344
rect 4028 1316 4036 1324
rect 4044 1316 4052 1324
rect 3948 1296 3956 1304
rect 3980 1296 3988 1304
rect 4028 1296 4036 1304
rect 3868 1236 3876 1244
rect 4044 1276 4052 1284
rect 4076 1276 4084 1284
rect 4060 1256 4068 1264
rect 3708 1216 3716 1224
rect 3820 1216 3828 1224
rect 3916 1216 3924 1224
rect 4076 1216 4084 1224
rect 3772 1196 3780 1204
rect 3836 1196 3844 1204
rect 3692 1156 3700 1164
rect 3740 1156 3748 1164
rect 3180 1116 3188 1124
rect 3212 1116 3220 1124
rect 3084 1096 3092 1104
rect 3164 1096 3172 1104
rect 3084 1056 3092 1064
rect 3148 1076 3156 1084
rect 3132 1056 3140 1064
rect 3260 1096 3268 1104
rect 3180 1056 3188 1064
rect 3196 1036 3204 1044
rect 3292 1036 3300 1044
rect 3324 1036 3332 1044
rect 3356 1036 3364 1044
rect 3420 1036 3428 1044
rect 3100 996 3108 1004
rect 2988 896 2996 904
rect 3004 896 3012 904
rect 2892 876 2900 884
rect 2860 816 2868 824
rect 3020 816 3028 824
rect 3164 936 3172 944
rect 3068 896 3076 904
rect 3132 896 3140 904
rect 3180 896 3188 904
rect 3116 856 3124 864
rect 3068 776 3076 784
rect 3052 756 3060 764
rect 2972 696 2980 704
rect 2876 676 2884 684
rect 2908 676 2916 684
rect 2956 676 2964 684
rect 3020 676 3028 684
rect 3052 676 3060 684
rect 3308 1016 3316 1024
rect 3276 956 3284 964
rect 3372 976 3380 984
rect 3340 956 3348 964
rect 3372 956 3380 964
rect 3260 936 3268 944
rect 3212 896 3220 904
rect 3340 896 3348 904
rect 3292 876 3300 884
rect 3180 836 3188 844
rect 3196 836 3204 844
rect 3260 836 3268 844
rect 3292 836 3300 844
rect 3228 796 3236 804
rect 3196 756 3204 764
rect 3180 716 3188 724
rect 3116 696 3124 704
rect 2812 656 2820 664
rect 2844 656 2852 664
rect 3052 636 3060 644
rect 3100 636 3108 644
rect 2700 616 2708 624
rect 2716 616 2724 624
rect 2828 616 2836 624
rect 2860 616 2868 624
rect 2684 556 2692 564
rect 2812 596 2820 604
rect 2876 596 2884 604
rect 2908 576 2916 584
rect 2764 556 2772 564
rect 2668 516 2676 524
rect 2684 516 2692 524
rect 2796 496 2804 504
rect 2844 496 2852 504
rect 2700 476 2708 484
rect 2428 456 2436 464
rect 2460 456 2468 464
rect 2636 456 2644 464
rect 2396 436 2404 444
rect 2700 436 2708 444
rect 2188 376 2196 384
rect 2332 376 2340 384
rect 2140 336 2148 344
rect 2268 336 2276 344
rect 2332 336 2340 344
rect 2620 336 2628 344
rect 2204 316 2212 324
rect 2140 296 2148 304
rect 2188 296 2196 304
rect 1964 276 1972 284
rect 1980 276 1988 284
rect 2108 276 2116 284
rect 2124 276 2132 284
rect 1980 236 1988 244
rect 1996 236 2004 244
rect 2028 236 2036 244
rect 2076 236 2084 244
rect 2092 236 2100 244
rect 1948 196 1956 204
rect 1868 136 1876 144
rect 1884 136 1892 144
rect 1820 36 1828 44
rect 2012 216 2020 224
rect 2092 196 2100 204
rect 2108 196 2116 204
rect 2028 176 2036 184
rect 2060 176 2068 184
rect 2508 316 2516 324
rect 2572 316 2580 324
rect 2604 316 2612 324
rect 2412 296 2420 304
rect 2524 296 2532 304
rect 2316 276 2324 284
rect 2204 256 2212 264
rect 2284 256 2292 264
rect 2236 196 2244 204
rect 2124 176 2132 184
rect 2220 176 2228 184
rect 2284 196 2292 204
rect 2428 276 2436 284
rect 2204 156 2212 164
rect 2044 136 2052 144
rect 2124 136 2132 144
rect 2172 136 2180 144
rect 1932 56 1940 64
rect 1980 56 1988 64
rect 2092 116 2100 124
rect 2396 256 2404 264
rect 2396 216 2404 224
rect 2476 276 2484 284
rect 2508 276 2516 284
rect 2444 216 2452 224
rect 2460 216 2468 224
rect 2476 196 2484 204
rect 2492 196 2500 204
rect 2428 176 2436 184
rect 2380 136 2388 144
rect 2172 96 2180 104
rect 2204 96 2212 104
rect 2412 96 2420 104
rect 2540 256 2548 264
rect 2604 256 2612 264
rect 2524 236 2532 244
rect 2572 236 2580 244
rect 2572 196 2580 204
rect 2940 556 2948 564
rect 3004 616 3012 624
rect 3052 576 3060 584
rect 3132 656 3140 664
rect 3148 636 3156 644
rect 3180 696 3188 704
rect 3452 1016 3460 1024
rect 3788 1156 3796 1164
rect 3900 1156 3908 1164
rect 3980 1156 3988 1164
rect 4060 1156 4068 1164
rect 3516 1096 3524 1104
rect 3532 1096 3540 1104
rect 3596 1096 3604 1104
rect 3772 1096 3780 1104
rect 3548 1076 3556 1084
rect 3612 1056 3620 1064
rect 3660 1056 3668 1064
rect 3676 1056 3684 1064
rect 3740 1056 3748 1064
rect 3756 1056 3764 1064
rect 3804 1056 3812 1064
rect 3516 1036 3524 1044
rect 3404 976 3412 984
rect 3468 976 3476 984
rect 3612 1016 3620 1024
rect 3628 1016 3636 1024
rect 3564 996 3572 1004
rect 3820 1036 3828 1044
rect 3484 956 3492 964
rect 3500 956 3508 964
rect 3532 956 3540 964
rect 3612 956 3620 964
rect 3660 956 3668 964
rect 3676 956 3684 964
rect 3436 936 3444 944
rect 3356 856 3364 864
rect 3372 796 3380 804
rect 3388 756 3396 764
rect 3292 716 3300 724
rect 3564 936 3572 944
rect 3500 836 3508 844
rect 3436 756 3444 764
rect 3212 636 3220 644
rect 3260 636 3268 644
rect 3132 616 3140 624
rect 3164 616 3172 624
rect 3228 616 3236 624
rect 3244 616 3252 624
rect 3148 596 3156 604
rect 3132 576 3140 584
rect 3020 556 3028 564
rect 2956 516 2964 524
rect 2972 496 2980 504
rect 3036 496 3044 504
rect 2924 476 2932 484
rect 2908 416 2916 424
rect 2924 416 2932 424
rect 2732 396 2740 404
rect 2828 396 2836 404
rect 2892 396 2900 404
rect 2652 356 2660 364
rect 2956 396 2964 404
rect 3036 396 3044 404
rect 3084 536 3092 544
rect 3084 516 3092 524
rect 3132 516 3140 524
rect 3116 496 3124 504
rect 3116 476 3124 484
rect 3084 436 3092 444
rect 3052 356 3060 364
rect 3068 356 3076 364
rect 2684 336 2692 344
rect 2668 316 2676 324
rect 2716 316 2724 324
rect 2812 316 2820 324
rect 2844 316 2852 324
rect 2940 316 2948 324
rect 3004 316 3012 324
rect 2684 276 2692 284
rect 2716 276 2724 284
rect 2732 276 2740 284
rect 2764 276 2772 284
rect 2796 256 2804 264
rect 2668 216 2676 224
rect 2732 216 2740 224
rect 2684 196 2692 204
rect 2652 156 2660 164
rect 2780 216 2788 224
rect 2844 276 2852 284
rect 2892 276 2900 284
rect 2828 256 2836 264
rect 2860 256 2868 264
rect 2892 256 2900 264
rect 2972 256 2980 264
rect 3004 256 3012 264
rect 3020 256 3028 264
rect 2764 196 2772 204
rect 2780 156 2788 164
rect 2892 216 2900 224
rect 2924 216 2932 224
rect 2956 216 2964 224
rect 2844 196 2852 204
rect 2876 196 2884 204
rect 2924 196 2932 204
rect 2524 116 2532 124
rect 2556 116 2564 124
rect 2572 116 2580 124
rect 2604 116 2612 124
rect 2684 116 2692 124
rect 2732 116 2740 124
rect 2796 116 2804 124
rect 2828 116 2836 124
rect 2428 76 2436 84
rect 2460 76 2468 84
rect 2540 76 2548 84
rect 1996 16 2004 24
rect 2012 16 2020 24
rect 2028 16 2036 24
rect 3004 216 3012 224
rect 3004 196 3012 204
rect 2972 176 2980 184
rect 3036 216 3044 224
rect 3196 576 3204 584
rect 3164 536 3172 544
rect 3260 556 3268 564
rect 3276 556 3284 564
rect 3308 536 3316 544
rect 3580 816 3588 824
rect 3532 796 3540 804
rect 3596 796 3604 804
rect 3564 776 3572 784
rect 3724 1016 3732 1024
rect 3836 1016 3844 1024
rect 3724 896 3732 904
rect 3756 956 3764 964
rect 3772 956 3780 964
rect 3804 956 3812 964
rect 4012 1096 4020 1104
rect 4380 1336 4388 1344
rect 4396 1336 4404 1344
rect 4956 1456 4964 1464
rect 4988 1456 4996 1464
rect 5020 1456 5028 1464
rect 5020 1376 5028 1384
rect 4972 1356 4980 1364
rect 4972 1336 4980 1344
rect 5004 1336 5012 1344
rect 4140 1316 4148 1324
rect 4172 1316 4180 1324
rect 4188 1316 4196 1324
rect 4124 1276 4132 1284
rect 4092 1176 4100 1184
rect 4108 1156 4116 1164
rect 3884 1056 3892 1064
rect 3932 1056 3940 1064
rect 3948 1056 3956 1064
rect 3868 1036 3876 1044
rect 3900 1036 3908 1044
rect 3884 1016 3892 1024
rect 3868 956 3876 964
rect 3756 896 3764 904
rect 3772 896 3780 904
rect 3804 896 3812 904
rect 3820 896 3828 904
rect 3852 896 3860 904
rect 4044 1016 4052 1024
rect 3916 976 3924 984
rect 3948 936 3956 944
rect 3964 936 3972 944
rect 4012 936 4020 944
rect 3900 916 3908 924
rect 3916 916 3924 924
rect 3932 916 3940 924
rect 3980 916 3988 924
rect 3996 916 4004 924
rect 3740 856 3748 864
rect 3948 896 3956 904
rect 3852 836 3860 844
rect 3660 776 3668 784
rect 3708 776 3716 784
rect 3596 736 3604 744
rect 3628 736 3636 744
rect 4012 816 4020 824
rect 4028 816 4036 824
rect 3788 796 3796 804
rect 3852 796 3860 804
rect 3996 776 4004 784
rect 3932 756 3940 764
rect 3948 756 3956 764
rect 4012 736 4020 744
rect 3836 716 3844 724
rect 3964 716 3972 724
rect 3980 716 3988 724
rect 3580 696 3588 704
rect 3628 696 3636 704
rect 3532 676 3540 684
rect 3452 656 3460 664
rect 3340 596 3348 604
rect 3468 616 3476 624
rect 3708 696 3716 704
rect 3692 676 3700 684
rect 3740 696 3748 704
rect 3740 676 3748 684
rect 3820 676 3828 684
rect 3516 616 3524 624
rect 3340 576 3348 584
rect 3436 576 3444 584
rect 3676 616 3684 624
rect 3708 616 3716 624
rect 3692 596 3700 604
rect 3580 556 3588 564
rect 3612 556 3620 564
rect 3276 516 3284 524
rect 3212 496 3220 504
rect 3132 456 3140 464
rect 3292 436 3300 444
rect 3148 416 3156 424
rect 3164 416 3172 424
rect 3100 296 3108 304
rect 3084 276 3092 284
rect 3244 396 3252 404
rect 3324 396 3332 404
rect 3180 376 3188 384
rect 3196 356 3204 364
rect 3308 376 3316 384
rect 3164 276 3172 284
rect 3212 276 3220 284
rect 3244 276 3252 284
rect 3068 236 3076 244
rect 3388 536 3396 544
rect 3404 536 3412 544
rect 3356 516 3364 524
rect 3644 536 3652 544
rect 3820 636 3828 644
rect 3852 636 3860 644
rect 3868 636 3876 644
rect 3756 616 3764 624
rect 3788 556 3796 564
rect 3820 556 3828 564
rect 3740 536 3748 544
rect 3756 536 3764 544
rect 3628 516 3636 524
rect 3660 516 3668 524
rect 3772 516 3780 524
rect 3372 496 3380 504
rect 3452 476 3460 484
rect 3548 476 3556 484
rect 3356 396 3364 404
rect 3372 396 3380 404
rect 3580 376 3588 384
rect 3612 376 3620 384
rect 3372 316 3380 324
rect 3452 316 3460 324
rect 3548 296 3556 304
rect 3612 296 3620 304
rect 3340 256 3348 264
rect 3468 256 3476 264
rect 3500 256 3508 264
rect 3420 216 3428 224
rect 3276 196 3284 204
rect 3292 196 3300 204
rect 3484 196 3492 204
rect 3148 176 3156 184
rect 3180 176 3188 184
rect 3356 176 3364 184
rect 3436 176 3444 184
rect 3596 176 3604 184
rect 3420 136 3428 144
rect 3564 136 3572 144
rect 3580 136 3588 144
rect 2956 116 2964 124
rect 3004 116 3012 124
rect 3020 116 3028 124
rect 3116 116 3124 124
rect 2972 56 2980 64
rect 2812 16 2820 24
rect 3052 76 3060 84
rect 3100 76 3108 84
rect 3692 476 3700 484
rect 3900 616 3908 624
rect 4236 1216 4244 1224
rect 4204 1196 4212 1204
rect 4204 1156 4212 1164
rect 4220 1156 4228 1164
rect 4540 1316 4548 1324
rect 4300 1296 4308 1304
rect 4316 1296 4324 1304
rect 4444 1296 4452 1304
rect 4572 1296 4580 1304
rect 4300 1276 4308 1284
rect 4316 1276 4324 1284
rect 4348 1276 4356 1284
rect 4460 1276 4468 1284
rect 4556 1276 4564 1284
rect 4348 1236 4356 1244
rect 4252 1176 4260 1184
rect 4220 1116 4228 1124
rect 4316 1116 4324 1124
rect 4204 1096 4212 1104
rect 4252 1096 4260 1104
rect 4156 1056 4164 1064
rect 4108 1016 4116 1024
rect 4124 1016 4132 1024
rect 4172 1016 4180 1024
rect 4140 976 4148 984
rect 4156 976 4164 984
rect 4108 956 4116 964
rect 4076 936 4084 944
rect 4204 996 4212 1004
rect 4284 996 4292 1004
rect 4300 996 4308 1004
rect 4524 1216 4532 1224
rect 4508 1176 4516 1184
rect 4540 1176 4548 1184
rect 4444 1156 4452 1164
rect 4652 1316 4660 1324
rect 4620 1296 4628 1304
rect 4700 1296 4708 1304
rect 4716 1296 4724 1304
rect 4764 1296 4772 1304
rect 4396 1136 4404 1144
rect 4460 1136 4468 1144
rect 4348 1116 4356 1124
rect 4364 1096 4372 1104
rect 4396 1096 4404 1104
rect 4444 1096 4452 1104
rect 4444 1076 4452 1084
rect 4588 1136 4596 1144
rect 4508 1096 4516 1104
rect 4444 1056 4452 1064
rect 4604 1076 4612 1084
rect 4540 1036 4548 1044
rect 4396 1016 4404 1024
rect 4508 1016 4516 1024
rect 4268 976 4276 984
rect 4332 976 4340 984
rect 4348 976 4356 984
rect 4588 1016 4596 1024
rect 4572 996 4580 1004
rect 4460 976 4468 984
rect 4860 1316 4868 1324
rect 4796 1296 4804 1304
rect 4876 1296 4884 1304
rect 4780 1276 4788 1284
rect 4812 1276 4820 1284
rect 4924 1276 4932 1284
rect 4956 1256 4964 1264
rect 4812 1236 4820 1244
rect 4860 1236 4868 1244
rect 4668 1196 4676 1204
rect 4732 1136 4740 1144
rect 4652 1116 4660 1124
rect 4796 1116 4804 1124
rect 4636 1076 4644 1084
rect 4684 1076 4692 1084
rect 4700 1076 4708 1084
rect 4764 1076 4772 1084
rect 4924 1116 4932 1124
rect 4828 1076 4836 1084
rect 4620 1016 4628 1024
rect 4716 996 4724 1004
rect 4668 976 4676 984
rect 4700 976 4708 984
rect 5068 1476 5076 1484
rect 5068 1436 5076 1444
rect 5084 1336 5092 1344
rect 5004 1236 5012 1244
rect 5004 1136 5012 1144
rect 4988 1096 4996 1104
rect 5020 1076 5028 1084
rect 4860 1056 4868 1064
rect 4924 1056 4932 1064
rect 4972 1056 4980 1064
rect 5036 1056 5044 1064
rect 4892 1036 4900 1044
rect 4764 996 4772 1004
rect 4732 976 4740 984
rect 4748 976 4756 984
rect 4780 976 4788 984
rect 4828 1016 4836 1024
rect 4876 1016 4884 1024
rect 4908 976 4916 984
rect 4156 936 4164 944
rect 4204 936 4212 944
rect 4236 936 4244 944
rect 4396 936 4404 944
rect 4492 936 4500 944
rect 4524 936 4532 944
rect 4604 936 4612 944
rect 4700 936 4708 944
rect 5068 1116 5076 1124
rect 4956 1016 4964 1024
rect 5052 1016 5060 1024
rect 5052 976 5060 984
rect 4956 956 4964 964
rect 5020 956 5028 964
rect 4076 916 4084 924
rect 4092 916 4100 924
rect 4060 856 4068 864
rect 4364 856 4372 864
rect 4300 836 4308 844
rect 4316 836 4324 844
rect 4044 796 4052 804
rect 4076 756 4084 764
rect 4092 756 4100 764
rect 4028 636 4036 644
rect 3996 616 4004 624
rect 4012 616 4020 624
rect 3964 596 3972 604
rect 3884 576 3892 584
rect 3932 576 3940 584
rect 3868 496 3876 504
rect 3884 496 3892 504
rect 3932 496 3940 504
rect 4028 596 4036 604
rect 4076 736 4084 744
rect 4060 716 4068 724
rect 4076 716 4084 724
rect 4156 716 4164 724
rect 4172 716 4180 724
rect 4076 636 4084 644
rect 4124 656 4132 664
rect 4108 636 4116 644
rect 4092 616 4100 624
rect 4044 576 4052 584
rect 4060 576 4068 584
rect 4076 556 4084 564
rect 4124 616 4132 624
rect 4140 616 4148 624
rect 4172 596 4180 604
rect 4156 556 4164 564
rect 4220 736 4228 744
rect 4284 736 4292 744
rect 4204 696 4212 704
rect 4252 696 4260 704
rect 4204 616 4212 624
rect 4300 636 4308 644
rect 4348 696 4356 704
rect 4604 916 4612 924
rect 4876 896 4884 904
rect 4908 896 4916 904
rect 5004 896 5012 904
rect 5020 896 5028 904
rect 5068 896 5076 904
rect 4604 876 4612 884
rect 4748 876 4756 884
rect 4764 876 4772 884
rect 5020 876 5028 884
rect 4444 836 4452 844
rect 4700 816 4708 824
rect 4428 776 4436 784
rect 4652 756 4660 764
rect 4396 736 4404 744
rect 4492 736 4500 744
rect 4636 736 4644 744
rect 4652 716 4660 724
rect 4380 696 4388 704
rect 4396 696 4404 704
rect 4492 696 4500 704
rect 4604 696 4612 704
rect 5052 816 5060 824
rect 4812 776 4820 784
rect 4892 756 4900 764
rect 4732 736 4740 744
rect 4796 736 4804 744
rect 4828 736 4836 744
rect 4876 736 4884 744
rect 4956 736 4964 744
rect 5036 736 5044 744
rect 4956 716 4964 724
rect 5148 1536 5156 1544
rect 5116 1516 5124 1524
rect 5132 1496 5140 1504
rect 5132 1476 5140 1484
rect 5100 1316 5108 1324
rect 5116 1316 5124 1324
rect 5100 1296 5108 1304
rect 5148 1456 5156 1464
rect 5148 1356 5156 1364
rect 5164 1296 5172 1304
rect 5132 1276 5140 1284
rect 5164 1276 5172 1284
rect 5100 1176 5108 1184
rect 5116 1156 5124 1164
rect 5116 1136 5124 1144
rect 5148 1096 5156 1104
rect 5132 976 5140 984
rect 5116 936 5124 944
rect 5148 956 5156 964
rect 5196 1336 5204 1344
rect 5196 1316 5204 1324
rect 5132 916 5140 924
rect 5132 756 5140 764
rect 5164 916 5172 924
rect 5196 1016 5204 1024
rect 5196 976 5204 984
rect 5196 896 5204 904
rect 5180 776 5188 784
rect 5148 736 5156 744
rect 4796 696 4804 704
rect 4908 696 4916 704
rect 5036 696 5044 704
rect 5084 696 5092 704
rect 4828 676 4836 684
rect 4924 676 4932 684
rect 4444 656 4452 664
rect 4524 656 4532 664
rect 4684 656 4692 664
rect 4716 656 4724 664
rect 4780 656 4788 664
rect 5004 656 5012 664
rect 4444 636 4452 644
rect 4204 596 4212 604
rect 4220 596 4228 604
rect 4252 596 4260 604
rect 4268 596 4276 604
rect 4316 596 4324 604
rect 4332 596 4340 604
rect 4492 596 4500 604
rect 4252 576 4260 584
rect 4316 576 4324 584
rect 4332 556 4340 564
rect 4524 556 4532 564
rect 4028 496 4036 504
rect 4044 496 4052 504
rect 4108 496 4116 504
rect 4156 496 4164 504
rect 3916 456 3924 464
rect 3836 436 3844 444
rect 3980 436 3988 444
rect 3852 376 3860 384
rect 3740 356 3748 364
rect 3644 336 3652 344
rect 3692 316 3700 324
rect 3660 296 3668 304
rect 3660 256 3668 264
rect 3772 336 3780 344
rect 3884 336 3892 344
rect 3676 216 3684 224
rect 3692 216 3700 224
rect 3804 316 3812 324
rect 3820 316 3828 324
rect 3836 316 3844 324
rect 3868 296 3876 304
rect 3964 316 3972 324
rect 3932 296 3940 304
rect 4060 396 4068 404
rect 4012 336 4020 344
rect 4076 316 4084 324
rect 4108 316 4116 324
rect 3852 236 3860 244
rect 3740 216 3748 224
rect 3772 216 3780 224
rect 3788 216 3796 224
rect 3804 216 3812 224
rect 3900 216 3908 224
rect 4188 436 4196 444
rect 4188 376 4196 384
rect 4236 536 4244 544
rect 4284 536 4292 544
rect 4364 536 4372 544
rect 4460 516 4468 524
rect 4428 496 4436 504
rect 4556 536 4564 544
rect 4604 596 4612 604
rect 4588 556 4596 564
rect 4972 616 4980 624
rect 4732 596 4740 604
rect 4796 596 4804 604
rect 4892 596 4900 604
rect 4924 596 4932 604
rect 4652 576 4660 584
rect 4716 576 4724 584
rect 4620 536 4628 544
rect 4652 536 4660 544
rect 4700 536 4708 544
rect 4540 496 4548 504
rect 4508 476 4516 484
rect 4476 456 4484 464
rect 4492 456 4500 464
rect 4252 436 4260 444
rect 4236 336 4244 344
rect 4460 416 4468 424
rect 4300 396 4308 404
rect 4396 396 4404 404
rect 4332 376 4340 384
rect 4316 336 4324 344
rect 4204 316 4212 324
rect 4428 336 4436 344
rect 4412 316 4420 324
rect 4332 296 4340 304
rect 4428 296 4436 304
rect 4156 276 4164 284
rect 4044 216 4052 224
rect 4012 196 4020 204
rect 4044 196 4052 204
rect 4092 196 4100 204
rect 4108 196 4116 204
rect 3964 176 3972 184
rect 4076 176 4084 184
rect 3740 156 3748 164
rect 3772 156 3780 164
rect 3868 156 3876 164
rect 4188 216 4196 224
rect 4140 196 4148 204
rect 4172 196 4180 204
rect 3756 136 3764 144
rect 3772 136 3780 144
rect 3788 136 3796 144
rect 3900 136 3908 144
rect 3292 116 3300 124
rect 3388 116 3396 124
rect 3564 116 3572 124
rect 3628 116 3636 124
rect 3900 116 3908 124
rect 4044 116 4052 124
rect 4076 116 4084 124
rect 4108 136 4116 144
rect 4172 136 4180 144
rect 3340 96 3348 104
rect 3532 96 3540 104
rect 3596 96 3604 104
rect 3644 96 3652 104
rect 3164 76 3172 84
rect 3196 76 3204 84
rect 3260 76 3268 84
rect 3148 56 3156 64
rect 3500 56 3508 64
rect 4220 196 4228 204
rect 4252 196 4260 204
rect 4364 276 4372 284
rect 4380 276 4388 284
rect 4412 276 4420 284
rect 4620 496 4628 504
rect 4588 476 4596 484
rect 4636 476 4644 484
rect 4620 436 4628 444
rect 4572 336 4580 344
rect 4604 336 4612 344
rect 4684 476 4692 484
rect 4716 476 4724 484
rect 4732 416 4740 424
rect 4828 576 4836 584
rect 4844 576 4852 584
rect 5036 596 5044 604
rect 5084 676 5092 684
rect 5148 656 5156 664
rect 5084 636 5092 644
rect 5068 616 5076 624
rect 5052 576 5060 584
rect 5116 596 5124 604
rect 5132 596 5140 604
rect 5212 616 5220 624
rect 4972 556 4980 564
rect 5052 556 5060 564
rect 5116 556 5124 564
rect 4812 536 4820 544
rect 4828 536 4836 544
rect 4876 536 4884 544
rect 4956 536 4964 544
rect 4924 516 4932 524
rect 5116 516 5124 524
rect 4764 396 4772 404
rect 4668 336 4676 344
rect 4556 316 4564 324
rect 4508 296 4516 304
rect 4620 296 4628 304
rect 4700 296 4708 304
rect 5084 496 5092 504
rect 4748 296 4756 304
rect 4796 296 4804 304
rect 4860 296 4868 304
rect 4524 276 4532 284
rect 4556 276 4564 284
rect 4652 276 4660 284
rect 4716 276 4724 284
rect 4780 276 4788 284
rect 4300 256 4308 264
rect 4348 256 4356 264
rect 4476 256 4484 264
rect 4604 256 4612 264
rect 4748 256 4756 264
rect 4460 236 4468 244
rect 4332 196 4340 204
rect 4412 196 4420 204
rect 4444 176 4452 184
rect 4476 156 4484 164
rect 4508 156 4516 164
rect 4828 276 4836 284
rect 4972 336 4980 344
rect 5020 336 5028 344
rect 5004 296 5012 304
rect 5020 276 5028 284
rect 4844 256 4852 264
rect 4876 256 4884 264
rect 4796 236 4804 244
rect 4972 236 4980 244
rect 4668 216 4676 224
rect 4780 216 4788 224
rect 4812 216 4820 224
rect 4668 196 4676 204
rect 4268 136 4276 144
rect 4284 136 4292 144
rect 4380 136 4388 144
rect 4396 136 4404 144
rect 4428 136 4436 144
rect 4860 196 4868 204
rect 4876 196 4884 204
rect 4764 156 4772 164
rect 4812 156 4820 164
rect 4844 156 4852 164
rect 4972 156 4980 164
rect 5004 156 5012 164
rect 5164 496 5172 504
rect 5164 416 5172 424
rect 5148 356 5156 364
rect 5100 336 5108 344
rect 5100 316 5108 324
rect 5132 296 5140 304
rect 5180 336 5188 344
rect 5052 276 5060 284
rect 5052 256 5060 264
rect 5180 176 5188 184
rect 5084 156 5092 164
rect 5132 156 5140 164
rect 5148 156 5156 164
rect 4684 136 4692 144
rect 4700 136 4708 144
rect 4812 136 4820 144
rect 4908 136 4916 144
rect 4940 136 4948 144
rect 5020 136 5028 144
rect 5068 136 5076 144
rect 4652 116 4660 124
rect 4732 116 4740 124
rect 4796 116 4804 124
rect 4892 116 4900 124
rect 5148 116 5156 124
rect 3948 96 3956 104
rect 4236 96 4244 104
rect 4476 96 4484 104
rect 4508 96 4516 104
rect 4556 96 4564 104
rect 4588 96 4596 104
rect 3772 76 3780 84
rect 4028 76 4036 84
rect 4060 76 4068 84
rect 4396 76 4404 84
<< metal3 >>
rect 2900 3617 3260 3623
rect 3380 3617 3388 3623
rect 4756 3617 4796 3623
rect 836 3597 1180 3603
rect 3652 3597 4028 3603
rect 4036 3597 4332 3603
rect 4340 3597 4652 3603
rect 4884 3597 4892 3603
rect 612 3577 1068 3583
rect 3668 3577 3676 3583
rect 3700 3577 3788 3583
rect 3796 3577 3884 3583
rect 3892 3577 4140 3583
rect 4148 3577 4508 3583
rect 708 3557 764 3563
rect 964 3557 972 3563
rect 1460 3557 1884 3563
rect 1924 3557 2060 3563
rect 2756 3557 3100 3563
rect 3108 3557 3308 3563
rect 3316 3557 4556 3563
rect 4564 3557 4796 3563
rect 4804 3557 4988 3563
rect 4996 3557 5052 3563
rect 324 3537 428 3543
rect 484 3537 492 3543
rect 564 3537 988 3543
rect 996 3537 1004 3543
rect 1012 3537 2380 3543
rect 2468 3537 2524 3543
rect 2900 3537 3356 3543
rect 3364 3537 4428 3543
rect 4436 3537 4748 3543
rect 340 3517 380 3523
rect 388 3517 1356 3523
rect 1389 3517 1404 3523
rect 1812 3517 1820 3523
rect 1956 3517 1964 3523
rect 2020 3517 2060 3523
rect 2116 3517 2156 3523
rect 2180 3517 2204 3523
rect 2228 3517 2332 3523
rect 2420 3517 2668 3523
rect 2676 3517 2684 3523
rect 2724 3517 2748 3523
rect 2845 3523 2851 3536
rect 2788 3517 2860 3523
rect 2884 3517 2908 3523
rect 2932 3517 3084 3523
rect 3092 3517 3404 3523
rect 3412 3517 3468 3523
rect 3476 3517 4380 3523
rect 4388 3517 4412 3523
rect 4452 3517 4460 3523
rect 4468 3517 4844 3523
rect 4852 3517 4956 3523
rect 4964 3517 4972 3523
rect 68 3497 108 3503
rect 116 3497 1148 3503
rect 1220 3497 1228 3503
rect 1268 3497 1308 3503
rect 1428 3497 1436 3503
rect 1444 3497 3068 3503
rect 3092 3497 3116 3503
rect 3124 3497 3276 3503
rect 3284 3497 3468 3503
rect 3492 3497 3564 3503
rect 3588 3497 4572 3503
rect 4612 3497 4716 3503
rect 4756 3497 4812 3503
rect 4836 3497 4844 3503
rect 4996 3497 5084 3503
rect 3069 3484 3075 3496
rect 228 3477 236 3483
rect 356 3477 380 3483
rect 420 3477 476 3483
rect 516 3477 652 3483
rect 676 3477 716 3483
rect 756 3477 1276 3483
rect 1348 3477 1388 3483
rect 1412 3477 1452 3483
rect 1492 3477 1724 3483
rect 1732 3477 1804 3483
rect 1844 3477 1852 3483
rect 1860 3477 2540 3483
rect 2660 3477 2764 3483
rect 2788 3477 3052 3483
rect 3108 3477 3404 3483
rect 3460 3477 3804 3483
rect 3812 3477 3820 3483
rect 3860 3477 3900 3483
rect 3924 3477 3932 3483
rect 4004 3477 4044 3483
rect 4084 3477 4300 3483
rect 4324 3477 4332 3483
rect 4388 3477 4396 3483
rect 4484 3477 4508 3483
rect 4516 3477 4556 3483
rect 4564 3477 4620 3483
rect 4660 3477 4860 3483
rect 4900 3477 5004 3483
rect 5044 3477 5052 3483
rect 2557 3464 2563 3476
rect 2573 3464 2579 3476
rect 148 3457 236 3463
rect 276 3457 716 3463
rect 804 3457 828 3463
rect 852 3457 860 3463
rect 932 3457 940 3463
rect 964 3457 972 3463
rect 980 3457 1180 3463
rect 1204 3457 1628 3463
rect 2036 3457 2044 3463
rect 2052 3457 2492 3463
rect 2708 3457 3148 3463
rect 3156 3457 3436 3463
rect 3460 3457 3500 3463
rect 3572 3457 3596 3463
rect 3620 3457 3628 3463
rect 3652 3457 3660 3463
rect 3716 3457 4236 3463
rect 4260 3457 4364 3463
rect 4372 3457 4460 3463
rect 4564 3457 4668 3463
rect 4676 3457 4684 3463
rect 4708 3457 4956 3463
rect 781 3444 787 3456
rect 2509 3444 2515 3456
rect 5165 3444 5171 3456
rect 132 3437 284 3443
rect 356 3437 364 3443
rect 468 3437 476 3443
rect 564 3437 572 3443
rect 644 3437 764 3443
rect 804 3437 812 3443
rect 1028 3437 1100 3443
rect 1172 3437 1244 3443
rect 1684 3437 1724 3443
rect 2228 3437 2236 3443
rect 2324 3437 2332 3443
rect 2372 3437 2380 3443
rect 2404 3437 2412 3443
rect 2484 3437 2492 3443
rect 2532 3437 2604 3443
rect 2612 3437 2732 3443
rect 2756 3437 3276 3443
rect 3284 3437 3308 3443
rect 3348 3437 3404 3443
rect 3412 3437 3548 3443
rect 3604 3437 4044 3443
rect 4068 3437 4156 3443
rect 4189 3437 4204 3443
rect 4276 3437 4396 3443
rect 4436 3437 4444 3443
rect 4468 3437 4492 3443
rect 4516 3437 4572 3443
rect 4580 3437 4604 3443
rect 4628 3437 4652 3443
rect 4676 3437 4684 3443
rect 4708 3437 4732 3443
rect 4836 3437 4892 3443
rect 4925 3424 4931 3436
rect 1108 3417 1228 3423
rect 1428 3417 1500 3423
rect 1508 3417 1644 3423
rect 1748 3417 1772 3423
rect 1780 3417 1980 3423
rect 1988 3417 2268 3423
rect 2324 3417 2764 3423
rect 2804 3417 2812 3423
rect 3044 3417 3052 3423
rect 3188 3417 3196 3423
rect 3236 3417 3372 3423
rect 3492 3417 3756 3423
rect 4180 3417 4444 3423
rect 4452 3417 4524 3423
rect 4532 3417 4780 3423
rect 628 3397 956 3403
rect 1156 3397 1164 3403
rect 1764 3397 1916 3403
rect 2276 3397 2316 3403
rect 2356 3397 2364 3403
rect 2516 3397 2620 3403
rect 2740 3397 2748 3403
rect 3028 3397 3100 3403
rect 3188 3397 3196 3403
rect 3220 3397 3228 3403
rect 3469 3397 3548 3403
rect 3133 3384 3139 3396
rect 20 3377 156 3383
rect 228 3377 348 3383
rect 548 3377 572 3383
rect 596 3377 636 3383
rect 740 3377 1324 3383
rect 1332 3377 1484 3383
rect 1508 3377 1516 3383
rect 1524 3377 3068 3383
rect 3156 3377 3260 3383
rect 3469 3383 3475 3397
rect 3572 3397 3708 3403
rect 4084 3397 4092 3403
rect 4164 3397 4172 3403
rect 4308 3397 4332 3403
rect 5108 3397 5116 3403
rect 3364 3377 3475 3383
rect 3492 3377 3731 3383
rect 20 3357 44 3363
rect 68 3357 108 3363
rect 212 3357 300 3363
rect 484 3357 540 3363
rect 548 3357 956 3363
rect 980 3357 1020 3363
rect 1060 3357 1100 3363
rect 1124 3357 1244 3363
rect 1300 3357 1308 3363
rect 1332 3357 1340 3363
rect 1396 3357 1468 3363
rect 1556 3357 1564 3363
rect 1581 3357 1612 3363
rect 100 3337 156 3343
rect 164 3337 284 3343
rect 292 3337 364 3343
rect 388 3337 396 3343
rect 484 3337 572 3343
rect 644 3337 700 3343
rect 724 3337 732 3343
rect 820 3337 828 3343
rect 852 3337 860 3343
rect 916 3337 1020 3343
rect 1037 3343 1043 3356
rect 1261 3344 1267 3356
rect 1037 3337 1052 3343
rect 1124 3337 1148 3343
rect 1172 3337 1212 3343
rect 1220 3337 1228 3343
rect 1581 3343 1587 3357
rect 1620 3357 1692 3363
rect 1732 3357 1740 3363
rect 1780 3357 2028 3363
rect 2164 3357 2380 3363
rect 2404 3357 2412 3363
rect 2484 3357 2508 3363
rect 2532 3357 2572 3363
rect 2612 3357 2620 3363
rect 2644 3357 2700 3363
rect 2724 3357 2844 3363
rect 2884 3357 2892 3363
rect 3060 3357 3084 3363
rect 3124 3357 3148 3363
rect 3172 3357 3180 3363
rect 3316 3357 3324 3363
rect 3396 3357 3484 3363
rect 3556 3357 3708 3363
rect 3725 3363 3731 3377
rect 3748 3377 4044 3383
rect 4052 3377 4268 3383
rect 4276 3377 4428 3383
rect 4468 3377 4476 3383
rect 4532 3377 4764 3383
rect 5108 3377 5116 3383
rect 4989 3364 4995 3376
rect 3725 3357 3756 3363
rect 3796 3357 3836 3363
rect 3860 3357 3948 3363
rect 3956 3357 3964 3363
rect 4013 3357 4028 3363
rect 4052 3357 4060 3363
rect 4180 3357 4380 3363
rect 4404 3357 4508 3363
rect 4708 3357 4748 3363
rect 4756 3357 4844 3363
rect 4884 3357 4940 3363
rect 5028 3357 5132 3363
rect 4093 3344 4099 3356
rect 1284 3337 1587 3343
rect 1604 3337 1788 3343
rect 1812 3337 1820 3343
rect 1860 3337 1868 3343
rect 1892 3337 2220 3343
rect 2244 3337 3036 3343
rect 3044 3337 3372 3343
rect 3460 3337 3852 3343
rect 3924 3337 3964 3343
rect 4004 3337 4076 3343
rect 4109 3337 4188 3343
rect 148 3317 1100 3323
rect 1108 3317 2748 3323
rect 2804 3317 2828 3323
rect 2868 3317 2876 3323
rect 2948 3317 3020 3323
rect 3124 3317 3132 3323
rect 3172 3317 3500 3323
rect 3508 3317 3532 3323
rect 3668 3317 3676 3323
rect 3764 3317 3900 3323
rect 4109 3323 4115 3337
rect 4212 3337 4284 3343
rect 4301 3337 4396 3343
rect 4036 3317 4115 3323
rect 4180 3317 4188 3323
rect 4301 3323 4307 3337
rect 4516 3337 4828 3343
rect 4868 3337 4972 3343
rect 4980 3337 5100 3343
rect 5124 3337 5164 3343
rect 4228 3317 4307 3323
rect 4324 3317 4332 3323
rect 4468 3317 4508 3323
rect 4692 3317 4732 3323
rect 4740 3317 4796 3323
rect 4916 3317 4924 3323
rect 5012 3317 5020 3323
rect 5028 3317 5068 3323
rect 2765 3304 2771 3316
rect 2925 3304 2931 3316
rect 116 3297 236 3303
rect 244 3297 252 3303
rect 356 3297 364 3303
rect 692 3297 876 3303
rect 900 3297 908 3303
rect 1076 3297 1116 3303
rect 1140 3297 1148 3303
rect 1156 3297 2556 3303
rect 2580 3297 2588 3303
rect 2628 3297 2636 3303
rect 2932 3297 3804 3303
rect 3828 3297 3852 3303
rect 3988 3297 3996 3303
rect 4052 3297 4060 3303
rect 4180 3297 4188 3303
rect 4260 3297 4316 3303
rect 4564 3297 4652 3303
rect 4660 3297 4972 3303
rect 5108 3297 5180 3303
rect 445 3284 451 3296
rect 493 3284 499 3296
rect 164 3277 284 3283
rect 516 3277 524 3283
rect 532 3277 956 3283
rect 964 3277 1180 3283
rect 1188 3277 1228 3283
rect 1460 3277 1596 3283
rect 1684 3277 1692 3283
rect 1732 3277 1740 3283
rect 2020 3277 2028 3283
rect 2180 3277 2188 3283
rect 2212 3277 2220 3283
rect 2276 3277 2364 3283
rect 2404 3277 2492 3283
rect 2532 3277 2540 3283
rect 2564 3277 3612 3283
rect 3620 3277 4268 3283
rect 4420 3277 4492 3283
rect 4500 3277 4636 3283
rect 4644 3277 4716 3283
rect 4980 3277 4988 3283
rect 4996 3277 5052 3283
rect 1837 3257 2044 3263
rect 1197 3244 1203 3256
rect 772 3237 780 3243
rect 1837 3243 1843 3257
rect 2084 3257 2124 3263
rect 2212 3257 2236 3263
rect 2292 3257 2300 3263
rect 3028 3257 3196 3263
rect 3252 3257 3260 3263
rect 3284 3257 3292 3263
rect 3396 3257 3436 3263
rect 4948 3257 5004 3263
rect 1604 3237 1843 3243
rect 1860 3237 1875 3243
rect 1940 3237 2732 3243
rect 2996 3237 3036 3243
rect 4612 3237 4620 3243
rect 4644 3237 4652 3243
rect 4660 3237 4668 3243
rect 4852 3237 4876 3243
rect 4964 3237 4972 3243
rect 5124 3237 5132 3243
rect 1901 3224 1907 3236
rect 4589 3224 4595 3236
rect 5037 3224 5043 3236
rect 196 3217 220 3223
rect 980 3217 988 3223
rect 1524 3217 1868 3223
rect 2964 3217 3132 3223
rect 3252 3217 3436 3223
rect 1348 3197 1932 3203
rect 1956 3197 2540 3203
rect 2548 3197 3036 3203
rect 3140 3197 3724 3203
rect 3844 3197 4524 3203
rect 1316 3177 1324 3183
rect 1364 3177 1372 3183
rect 1444 3177 2076 3183
rect 2196 3177 2220 3183
rect 2228 3177 2252 3183
rect 2276 3177 2828 3183
rect 3108 3177 3116 3183
rect 3780 3177 3836 3183
rect 3860 3177 4556 3183
rect 4836 3177 5036 3183
rect 5044 3177 5068 3183
rect 516 3157 524 3163
rect 708 3157 956 3163
rect 1028 3157 2316 3163
rect 2564 3157 2924 3163
rect 3005 3157 3020 3163
rect 212 3137 1084 3143
rect 1732 3137 2796 3143
rect 2804 3137 2812 3143
rect 3005 3143 3011 3157
rect 3524 3157 3692 3163
rect 3796 3157 3804 3163
rect 4308 3157 4396 3163
rect 4948 3157 4988 3163
rect 3037 3144 3043 3156
rect 2932 3137 3011 3143
rect 3060 3137 3068 3143
rect 3460 3137 3516 3143
rect 3540 3137 3932 3143
rect 4013 3137 4028 3143
rect 4116 3137 4316 3143
rect 4356 3137 4364 3143
rect 4692 3137 4700 3143
rect 4772 3137 4796 3143
rect 4820 3137 4892 3143
rect 1357 3124 1363 3136
rect 1405 3124 1411 3136
rect 4749 3124 4755 3136
rect 68 3117 172 3123
rect 260 3117 732 3123
rect 900 3117 1340 3123
rect 1508 3117 1660 3123
rect 1684 3117 1692 3123
rect 1796 3117 2108 3123
rect 2116 3117 2124 3123
rect 2132 3117 2220 3123
rect 2244 3117 2460 3123
rect 2468 3117 2476 3123
rect 2484 3117 3452 3123
rect 3524 3117 3532 3123
rect 3556 3117 3564 3123
rect 3636 3117 3644 3123
rect 4052 3117 4300 3123
rect 4436 3117 4444 3123
rect 4692 3117 4716 3123
rect 4772 3117 4844 3123
rect 4852 3117 4860 3123
rect 4900 3117 4908 3123
rect 4932 3117 5004 3123
rect 5012 3117 5164 3123
rect 189 3104 195 3116
rect 733 3104 739 3116
rect 4029 3104 4035 3116
rect 4557 3104 4563 3116
rect 20 3097 44 3103
rect 164 3097 172 3103
rect 196 3097 300 3103
rect 324 3097 364 3103
rect 404 3097 700 3103
rect 772 3097 780 3103
rect 804 3097 876 3103
rect 996 3097 1004 3103
rect 1076 3097 1100 3103
rect 1156 3097 1196 3103
rect 1284 3097 1292 3103
rect 1300 3097 1772 3103
rect 1796 3097 1852 3103
rect 1924 3097 1932 3103
rect 1972 3097 2012 3103
rect 2068 3097 2076 3103
rect 2180 3097 2188 3103
rect 2212 3097 2220 3103
rect 2260 3097 2332 3103
rect 2356 3097 2380 3103
rect 2420 3097 2620 3103
rect 2644 3097 3068 3103
rect 3140 3097 3356 3103
rect 3380 3097 3388 3103
rect 3412 3097 3932 3103
rect 3940 3097 3948 3103
rect 4068 3097 4076 3103
rect 4148 3097 4204 3103
rect 4404 3097 4444 3103
rect 4516 3097 4524 3103
rect 4596 3097 4604 3103
rect 4644 3097 4940 3103
rect 180 3077 204 3083
rect 228 3077 236 3083
rect 276 3077 316 3083
rect 356 3077 396 3083
rect 468 3077 588 3083
rect 612 3077 732 3083
rect 756 3077 780 3083
rect 820 3077 828 3083
rect 932 3077 940 3083
rect 948 3077 1020 3083
rect 1028 3077 1164 3083
rect 1188 3077 1196 3083
rect 1277 3077 1532 3083
rect 228 3057 828 3063
rect 836 3057 972 3063
rect 1277 3063 1283 3077
rect 1588 3077 2268 3083
rect 2308 3077 2371 3083
rect 1140 3057 1283 3063
rect 1316 3057 1628 3063
rect 1652 3057 2204 3063
rect 2228 3057 2348 3063
rect 2365 3063 2371 3077
rect 2388 3077 2652 3083
rect 2772 3077 2780 3083
rect 2804 3077 2844 3083
rect 2916 3077 2956 3083
rect 3028 3077 3292 3083
rect 3316 3077 3356 3083
rect 3396 3077 4124 3083
rect 4132 3077 4252 3083
rect 4356 3077 4604 3083
rect 4724 3077 4732 3083
rect 4740 3077 5020 3083
rect 2685 3064 2691 3076
rect 2973 3064 2979 3076
rect 2365 3057 2428 3063
rect 2484 3057 2668 3063
rect 2708 3057 2819 3063
rect 1117 3044 1123 3056
rect 2445 3044 2451 3056
rect 212 3037 556 3043
rect 612 3037 684 3043
rect 724 3037 796 3043
rect 820 3037 940 3043
rect 980 3037 1036 3043
rect 1076 3037 1084 3043
rect 1236 3037 1548 3043
rect 1556 3037 2156 3043
rect 2164 3037 2396 3043
rect 2468 3037 2492 3043
rect 2516 3037 2524 3043
rect 2548 3037 2588 3043
rect 2612 3037 2620 3043
rect 2660 3037 2796 3043
rect 2813 3043 2819 3057
rect 3076 3057 3084 3063
rect 3220 3057 3276 3063
rect 3380 3057 3388 3063
rect 3412 3057 3420 3063
rect 3460 3057 3468 3063
rect 3524 3057 3532 3063
rect 3549 3044 3555 3063
rect 3572 3057 3628 3063
rect 3700 3057 3811 3063
rect 3677 3044 3683 3056
rect 2813 3037 3084 3043
rect 3172 3037 3228 3043
rect 3300 3037 3436 3043
rect 3460 3037 3484 3043
rect 3805 3043 3811 3057
rect 3828 3057 3996 3063
rect 4068 3057 4476 3063
rect 4484 3057 4668 3063
rect 4708 3057 4796 3063
rect 4804 3057 4892 3063
rect 4900 3057 4940 3063
rect 4948 3057 4956 3063
rect 5060 3057 5084 3063
rect 4061 3044 4067 3056
rect 3805 3037 3868 3043
rect 4180 3037 4220 3043
rect 4308 3037 4332 3043
rect 4564 3037 4572 3043
rect 4653 3037 4668 3043
rect 4788 3037 4828 3043
rect 4884 3037 4988 3043
rect 4996 3037 5116 3043
rect 580 3017 652 3023
rect 676 3017 1196 3023
rect 1284 3017 1708 3023
rect 1860 3017 1964 3023
rect 1972 3017 2908 3023
rect 2932 3017 2988 3023
rect 3204 3017 3212 3023
rect 3444 3017 3596 3023
rect 4292 3017 4348 3023
rect 4660 3017 4716 3023
rect 84 2997 140 3003
rect 516 2997 892 3003
rect 948 2997 956 3003
rect 1012 2997 1036 3003
rect 1092 2997 1164 3003
rect 1476 2997 1964 3003
rect 1972 2997 2028 3003
rect 2100 2997 2108 3003
rect 2164 2997 2572 3003
rect 2580 2997 2636 3003
rect 2756 2997 2876 3003
rect 2900 2997 2908 3003
rect 2996 2997 3484 3003
rect 3492 2997 3523 3003
rect 292 2977 396 2983
rect 468 2977 524 2983
rect 564 2977 668 2983
rect 692 2977 764 2983
rect 788 2977 844 2983
rect 852 2977 1132 2983
rect 1156 2977 1228 2983
rect 1252 2977 1308 2983
rect 1316 2977 1324 2983
rect 1348 2977 1372 2983
rect 1412 2977 1420 2983
rect 1444 2977 1452 2983
rect 1476 2977 2364 2983
rect 2372 2977 3260 2983
rect 3460 2977 3468 2983
rect 3492 2977 3500 2983
rect 3517 2983 3523 2997
rect 3556 2997 3580 3003
rect 3620 2997 4044 3003
rect 4068 2997 4108 3003
rect 4132 2997 4268 3003
rect 4420 2997 4492 3003
rect 4900 2997 4908 3003
rect 3517 2977 3804 2983
rect 3908 2977 4940 2983
rect 5060 2977 5068 2983
rect 68 2957 172 2963
rect 324 2957 412 2963
rect 452 2957 460 2963
rect 484 2957 940 2963
rect 964 2957 972 2963
rect 996 2957 1356 2963
rect 1364 2957 2252 2963
rect 2260 2957 2476 2963
rect 2548 2957 2556 2963
rect 2628 2957 2652 2963
rect 2708 2957 2716 2963
rect 2836 2957 2844 2963
rect 2868 2957 3340 2963
rect 3348 2957 3564 2963
rect 3620 2957 3692 2963
rect 3796 2957 3900 2963
rect 3956 2957 4380 2963
rect 4388 2957 4732 2963
rect 4740 2957 4908 2963
rect 4948 2957 5052 2963
rect 5092 2957 5100 2963
rect 2477 2944 2483 2956
rect 52 2937 108 2943
rect 148 2937 252 2943
rect 260 2937 508 2943
rect 548 2937 556 2943
rect 660 2937 684 2943
rect 708 2937 716 2943
rect 724 2937 796 2943
rect 804 2937 1596 2943
rect 1668 2937 1916 2943
rect 1940 2937 1948 2943
rect 1972 2937 2028 2943
rect 2052 2937 2060 2943
rect 2148 2937 2444 2943
rect 2516 2937 2572 2943
rect 2596 2937 2620 2943
rect 2676 2937 3020 2943
rect 3044 2937 3052 2943
rect 3060 2937 3180 2943
rect 3188 2937 3292 2943
rect 3364 2937 3708 2943
rect 3716 2937 4028 2943
rect 4052 2937 4060 2943
rect 4100 2937 4204 2943
rect 4260 2937 4700 2943
rect 4724 2937 4732 2943
rect 4820 2937 4860 2943
rect 5101 2924 5107 2936
rect 148 2917 236 2923
rect 308 2917 316 2923
rect 356 2917 380 2923
rect 388 2917 524 2923
rect 548 2917 700 2923
rect 724 2917 764 2923
rect 788 2917 812 2923
rect 836 2917 844 2923
rect 852 2917 1836 2923
rect 1860 2917 1884 2923
rect 1908 2917 2076 2923
rect 2116 2917 2140 2923
rect 2196 2917 2204 2923
rect 2276 2917 2284 2923
rect 2292 2917 2764 2923
rect 2772 2917 3132 2923
rect 3156 2917 3180 2923
rect 3252 2917 3276 2923
rect 3316 2917 3468 2923
rect 3492 2917 3532 2923
rect 3556 2917 3596 2923
rect 3668 2917 3692 2923
rect 3860 2917 3875 2923
rect 109 2904 115 2916
rect 3629 2904 3635 2916
rect 3837 2904 3843 2916
rect 3869 2904 3875 2917
rect 3940 2917 3980 2923
rect 4004 2917 4012 2923
rect 4036 2917 4252 2923
rect 4260 2917 4268 2923
rect 4372 2917 4492 2923
rect 4516 2917 4524 2923
rect 4564 2917 4748 2923
rect 4756 2917 5020 2923
rect 5028 2917 5084 2923
rect 404 2897 412 2903
rect 436 2897 476 2903
rect 596 2897 604 2903
rect 660 2897 668 2903
rect 676 2897 780 2903
rect 788 2897 796 2903
rect 820 2897 860 2903
rect 884 2897 988 2903
rect 1076 2897 1084 2903
rect 1188 2897 1244 2903
rect 1268 2897 1404 2903
rect 1428 2897 1436 2903
rect 1460 2897 1468 2903
rect 1492 2897 1500 2903
rect 1508 2897 1580 2903
rect 1684 2897 1692 2903
rect 1700 2897 1708 2903
rect 1780 2897 1804 2903
rect 1828 2897 1836 2903
rect 1876 2897 1884 2903
rect 1924 2897 2316 2903
rect 2340 2897 2428 2903
rect 2452 2897 2940 2903
rect 3028 2897 3036 2903
rect 3108 2897 3116 2903
rect 3188 2897 3196 2903
rect 3236 2897 3308 2903
rect 3380 2897 3388 2903
rect 3412 2897 3420 2903
rect 3556 2897 3564 2903
rect 3748 2897 3756 2903
rect 3892 2897 3996 2903
rect 4052 2897 4124 2903
rect 4148 2897 4156 2903
rect 4436 2897 4460 2903
rect 4692 2897 4732 2903
rect 4756 2897 5004 2903
rect 5140 2897 5148 2903
rect 285 2884 291 2896
rect 340 2877 508 2883
rect 516 2877 908 2883
rect 964 2877 972 2883
rect 1252 2877 1292 2883
rect 1412 2877 1436 2883
rect 1636 2877 1772 2883
rect 1828 2877 1916 2883
rect 1988 2877 1996 2883
rect 2020 2877 2028 2883
rect 2068 2877 2220 2883
rect 2276 2877 2300 2883
rect 2372 2877 2380 2883
rect 2596 2877 2604 2883
rect 2644 2877 2668 2883
rect 2932 2877 2940 2883
rect 2996 2877 3004 2883
rect 3012 2877 3852 2883
rect 3860 2877 4012 2883
rect 4132 2877 4140 2883
rect 4452 2877 4476 2883
rect 4660 2877 4812 2883
rect 5124 2877 5132 2883
rect 1933 2864 1939 2876
rect 388 2857 412 2863
rect 788 2857 1004 2863
rect 1284 2857 1628 2863
rect 1716 2857 1724 2863
rect 1764 2857 1900 2863
rect 1956 2857 2108 2863
rect 2132 2857 2556 2863
rect 2580 2857 2588 2863
rect 2612 2857 2620 2863
rect 2676 2857 3036 2863
rect 3412 2857 3420 2863
rect 4180 2857 4812 2863
rect 4820 2857 4892 2863
rect 4900 2857 4956 2863
rect 5124 2857 5148 2863
rect 1188 2837 1580 2843
rect 1604 2837 1708 2843
rect 1716 2837 2172 2843
rect 2244 2837 2684 2843
rect 2836 2837 3644 2843
rect 3652 2837 3868 2843
rect 4148 2837 4172 2843
rect 461 2824 467 2836
rect 4317 2824 4323 2836
rect 5005 2824 5011 2836
rect 660 2817 1260 2823
rect 1332 2817 1388 2823
rect 1732 2817 1772 2823
rect 1796 2817 1804 2823
rect 1828 2817 1916 2823
rect 1988 2817 2268 2823
rect 2292 2817 2300 2823
rect 2660 2817 2716 2823
rect 2804 2817 2828 2823
rect 2964 2817 2972 2823
rect 3396 2817 3404 2823
rect 4244 2817 4300 2823
rect 5172 2817 5212 2823
rect 404 2797 476 2803
rect 692 2797 2508 2803
rect 2564 2797 2988 2803
rect 3092 2797 3356 2803
rect 3524 2797 3532 2803
rect 3892 2797 3900 2803
rect 4404 2797 4412 2803
rect 4436 2797 5164 2803
rect 580 2777 812 2783
rect 932 2777 1020 2783
rect 1252 2777 1436 2783
rect 1700 2777 1836 2783
rect 2068 2777 2092 2783
rect 2164 2777 2700 2783
rect 2756 2777 3276 2783
rect 3300 2777 3308 2783
rect 3492 2777 3516 2783
rect 3844 2777 3980 2783
rect 3988 2777 4620 2783
rect 340 2757 492 2763
rect 500 2757 2732 2763
rect 2740 2757 2892 2763
rect 2900 2757 3116 2763
rect 3172 2757 3180 2763
rect 3364 2757 3484 2763
rect 3492 2757 4012 2763
rect 4052 2757 4108 2763
rect 4164 2757 4172 2763
rect 4196 2757 4348 2763
rect 4404 2757 4412 2763
rect 4500 2757 4508 2763
rect 5156 2757 5164 2763
rect 4829 2744 4835 2756
rect 148 2737 188 2743
rect 196 2737 300 2743
rect 493 2737 508 2743
rect 644 2737 924 2743
rect 932 2737 1052 2743
rect 1204 2737 1788 2743
rect 1892 2737 1900 2743
rect 2004 2737 2012 2743
rect 2052 2737 2092 2743
rect 2148 2737 2156 2743
rect 2196 2737 2316 2743
rect 2436 2737 2492 2743
rect 2564 2737 2668 2743
rect 2708 2737 2780 2743
rect 2804 2737 2812 2743
rect 2836 2737 2924 2743
rect 2948 2737 2956 2743
rect 3028 2737 3052 2743
rect 3060 2737 3164 2743
rect 3428 2737 3660 2743
rect 3668 2737 3964 2743
rect 3972 2737 4124 2743
rect 4148 2737 4764 2743
rect 4900 2737 4908 2743
rect 5076 2737 5148 2743
rect 3197 2724 3203 2736
rect 52 2717 60 2723
rect 100 2717 108 2723
rect 244 2717 284 2723
rect 292 2717 636 2723
rect 708 2717 716 2723
rect 916 2717 924 2723
rect 996 2717 1004 2723
rect 1092 2717 1100 2723
rect 1284 2717 1292 2723
rect 1332 2717 1356 2723
rect 1460 2717 1516 2723
rect 1572 2717 1900 2723
rect 1908 2717 2252 2723
rect 2420 2717 2508 2723
rect 2612 2717 2620 2723
rect 2644 2717 3100 2723
rect 3220 2717 3228 2723
rect 3284 2717 3308 2723
rect 3364 2717 3388 2723
rect 3492 2717 3532 2723
rect 3556 2717 3564 2723
rect 3652 2717 3916 2723
rect 3924 2717 3932 2723
rect 4052 2717 4060 2723
rect 4100 2717 4140 2723
rect 4164 2717 4620 2723
rect 4628 2717 4828 2723
rect 4836 2717 4972 2723
rect 5092 2717 5100 2723
rect 20 2697 1148 2703
rect 1204 2697 1420 2703
rect 1508 2697 1516 2703
rect 1604 2697 1612 2703
rect 1620 2697 3004 2703
rect 3012 2697 3068 2703
rect 3108 2697 3676 2703
rect 3684 2697 3708 2703
rect 3764 2697 3852 2703
rect 3892 2697 3932 2703
rect 3940 2697 4540 2703
rect 4548 2697 4636 2703
rect 4676 2697 4684 2703
rect 4724 2697 4764 2703
rect 4788 2697 4844 2703
rect 4861 2697 4876 2703
rect 4884 2697 4908 2703
rect 116 2677 492 2683
rect 532 2677 540 2683
rect 564 2677 572 2683
rect 596 2677 700 2683
rect 804 2677 812 2683
rect 836 2677 940 2683
rect 948 2677 972 2683
rect 1012 2677 1020 2683
rect 1044 2677 1100 2683
rect 1124 2677 1132 2683
rect 1156 2677 1228 2683
rect 1236 2677 1244 2683
rect 1268 2677 1452 2683
rect 1460 2677 1500 2683
rect 1524 2677 1948 2683
rect 1956 2677 2380 2683
rect 2628 2677 2748 2683
rect 2964 2677 3148 2683
rect 3156 2677 4156 2683
rect 4164 2677 4220 2683
rect 4260 2677 4284 2683
rect 4324 2677 4332 2683
rect 4388 2677 4444 2683
rect 4468 2677 4492 2683
rect 4516 2677 4604 2683
rect 4644 2677 4940 2683
rect 4948 2677 4956 2683
rect 4980 2677 5052 2683
rect 5092 2677 5100 2683
rect 164 2657 172 2663
rect 244 2657 268 2663
rect 292 2657 300 2663
rect 324 2657 348 2663
rect 429 2657 444 2663
rect 196 2637 380 2643
rect 413 2637 419 2656
rect 429 2644 435 2657
rect 468 2657 652 2663
rect 804 2657 812 2663
rect 852 2657 860 2663
rect 884 2657 1132 2663
rect 1156 2657 1244 2663
rect 1316 2657 2652 2663
rect 2692 2657 2700 2663
rect 2708 2657 2860 2663
rect 2916 2657 2972 2663
rect 2980 2657 3068 2663
rect 3085 2657 3212 2663
rect 2893 2644 2899 2656
rect 484 2637 572 2643
rect 708 2637 748 2643
rect 996 2637 1356 2643
rect 1364 2637 1564 2643
rect 1652 2637 1708 2643
rect 1860 2637 2044 2643
rect 2068 2637 2268 2643
rect 2308 2637 2316 2643
rect 2500 2637 2524 2643
rect 2612 2637 2636 2643
rect 2676 2637 2700 2643
rect 2756 2637 2844 2643
rect 2916 2637 2988 2643
rect 3085 2643 3091 2657
rect 3252 2657 3260 2663
rect 3300 2657 3324 2663
rect 3396 2657 3452 2663
rect 3572 2657 3628 2663
rect 3668 2657 3740 2663
rect 3844 2657 4876 2663
rect 4884 2657 4972 2663
rect 4996 2657 5004 2663
rect 5060 2657 5068 2663
rect 3012 2637 3091 2643
rect 3140 2637 3564 2643
rect 3620 2637 3660 2643
rect 3684 2637 3724 2643
rect 3844 2637 3852 2643
rect 3860 2637 4092 2643
rect 4100 2637 4684 2643
rect 4900 2637 4924 2643
rect 5108 2637 5116 2643
rect 228 2617 995 2623
rect 68 2597 76 2603
rect 100 2597 124 2603
rect 132 2597 252 2603
rect 276 2597 284 2603
rect 340 2597 572 2603
rect 580 2597 620 2603
rect 989 2603 995 2617
rect 1012 2617 1036 2623
rect 1044 2617 1052 2623
rect 1332 2617 1340 2623
rect 1556 2617 1564 2623
rect 1956 2617 1964 2623
rect 2100 2617 2108 2623
rect 2164 2617 2172 2623
rect 2196 2617 2204 2623
rect 2276 2617 2300 2623
rect 2388 2617 2412 2623
rect 2436 2617 2444 2623
rect 2484 2617 3260 2623
rect 3364 2617 3436 2623
rect 3492 2617 3500 2623
rect 3588 2617 3596 2623
rect 3668 2617 3916 2623
rect 4036 2617 4044 2623
rect 4068 2617 4076 2623
rect 4148 2617 4204 2623
rect 4260 2617 4284 2623
rect 4468 2617 5020 2623
rect 5037 2617 5196 2623
rect 989 2597 1372 2603
rect 1380 2597 1708 2603
rect 1796 2597 2076 2603
rect 2100 2597 2188 2603
rect 2404 2597 2531 2603
rect 148 2577 236 2583
rect 468 2577 508 2583
rect 516 2577 540 2583
rect 692 2577 716 2583
rect 740 2577 764 2583
rect 836 2577 844 2583
rect 964 2577 1116 2583
rect 1140 2577 1260 2583
rect 1268 2577 1676 2583
rect 1732 2577 1980 2583
rect 2084 2577 2396 2583
rect 2420 2577 2460 2583
rect 2525 2583 2531 2597
rect 2564 2597 3148 2603
rect 3204 2597 3244 2603
rect 3268 2597 3692 2603
rect 4052 2597 4124 2603
rect 4148 2597 4172 2603
rect 4253 2597 4316 2603
rect 3869 2584 3875 2596
rect 4013 2584 4019 2596
rect 2525 2577 2732 2583
rect 2740 2577 2828 2583
rect 2964 2577 3532 2583
rect 3556 2577 3612 2583
rect 3716 2577 3740 2583
rect 4253 2583 4259 2597
rect 4452 2597 4492 2603
rect 5037 2603 5043 2617
rect 5012 2597 5043 2603
rect 5108 2597 5116 2603
rect 4084 2577 4259 2583
rect 4308 2577 4348 2583
rect 4372 2577 4380 2583
rect 4500 2577 4604 2583
rect 4740 2577 4972 2583
rect 5156 2577 5164 2583
rect 2029 2564 2035 2576
rect 116 2557 1356 2563
rect 1364 2557 1372 2563
rect 1380 2557 1724 2563
rect 1796 2557 1804 2563
rect 1828 2557 1836 2563
rect 1988 2557 1996 2563
rect 2052 2557 2060 2563
rect 2084 2557 2124 2563
rect 2164 2557 2179 2563
rect 2196 2557 2316 2563
rect 2340 2557 2380 2563
rect 2404 2557 2524 2563
rect 2708 2557 2748 2563
rect 2804 2557 2812 2563
rect 2884 2557 2908 2563
rect 2932 2557 2940 2563
rect 2980 2557 3004 2563
rect 3028 2557 3132 2563
rect 3156 2557 3212 2563
rect 3236 2557 3292 2563
rect 3316 2557 3452 2563
rect 3460 2557 3788 2563
rect 3924 2557 3932 2563
rect 3940 2557 4060 2563
rect 4084 2557 4108 2563
rect 4148 2557 4156 2563
rect 4260 2557 4604 2563
rect 4612 2557 4652 2563
rect 4804 2557 5084 2563
rect 5092 2557 5100 2563
rect 116 2537 796 2543
rect 932 2537 940 2543
rect 948 2537 1068 2543
rect 1172 2537 1196 2543
rect 1284 2537 1292 2543
rect 1332 2537 1340 2543
rect 1396 2537 1404 2543
rect 1444 2537 2316 2543
rect 2372 2537 2444 2543
rect 2500 2537 2524 2543
rect 2564 2537 2588 2543
rect 2644 2537 2668 2543
rect 2692 2537 2924 2543
rect 2932 2537 4108 2543
rect 4116 2537 4204 2543
rect 4260 2537 4924 2543
rect 4932 2537 5052 2543
rect 20 2517 108 2523
rect 324 2517 332 2523
rect 356 2517 540 2523
rect 548 2517 556 2523
rect 701 2517 716 2523
rect 756 2517 780 2523
rect 836 2517 1036 2523
rect 1060 2517 1212 2523
rect 1236 2517 1276 2523
rect 1300 2517 1308 2523
rect 1316 2517 1740 2523
rect 1892 2517 2908 2523
rect 2932 2517 3212 2523
rect 3220 2517 3372 2523
rect 3389 2517 3452 2523
rect 196 2497 204 2503
rect 212 2497 220 2503
rect 244 2497 428 2503
rect 452 2497 476 2503
rect 500 2497 508 2503
rect 516 2497 652 2503
rect 660 2497 924 2503
rect 980 2497 1020 2503
rect 1076 2497 1132 2503
rect 1156 2497 1388 2503
rect 1428 2497 1628 2503
rect 1732 2497 1740 2503
rect 1828 2497 1836 2503
rect 1908 2497 1916 2503
rect 2004 2497 2060 2503
rect 2132 2497 2188 2503
rect 2228 2497 2236 2503
rect 2276 2497 2291 2503
rect 2308 2497 2348 2503
rect 2356 2497 2364 2503
rect 2548 2497 2556 2503
rect 2676 2497 2684 2503
rect 2708 2497 2716 2503
rect 2756 2497 2764 2503
rect 2788 2497 2876 2503
rect 2884 2497 2924 2503
rect 2948 2497 2988 2503
rect 3044 2497 3052 2503
rect 3060 2497 3116 2503
rect 3124 2497 3180 2503
rect 3220 2497 3228 2503
rect 3252 2497 3260 2503
rect 3389 2503 3395 2517
rect 3460 2517 3484 2523
rect 3508 2517 3532 2523
rect 3572 2517 3612 2523
rect 3668 2517 3740 2523
rect 3860 2517 3916 2523
rect 3924 2517 3932 2523
rect 3956 2517 4060 2523
rect 4116 2517 4124 2523
rect 4164 2517 4172 2523
rect 4196 2517 4236 2523
rect 4340 2517 4444 2523
rect 4468 2517 4476 2523
rect 4500 2517 4508 2523
rect 4548 2517 4588 2523
rect 4685 2517 4716 2523
rect 3821 2504 3827 2516
rect 3332 2497 3395 2503
rect 3428 2497 3468 2503
rect 3540 2497 3564 2503
rect 3588 2497 3740 2503
rect 3748 2497 3756 2503
rect 3828 2497 3900 2503
rect 4004 2497 4012 2503
rect 4077 2503 4083 2516
rect 4077 2497 4092 2503
rect 4141 2503 4147 2516
rect 4285 2504 4291 2516
rect 4605 2504 4611 2516
rect 4132 2497 4147 2503
rect 4164 2497 4236 2503
rect 4484 2497 4508 2503
rect 2413 2484 2419 2496
rect 52 2477 140 2483
rect 148 2477 764 2483
rect 836 2477 860 2483
rect 948 2477 956 2483
rect 964 2477 1484 2483
rect 1508 2477 1516 2483
rect 1540 2477 1564 2483
rect 1636 2477 1644 2483
rect 1700 2477 1788 2483
rect 1844 2477 2204 2483
rect 2212 2477 2364 2483
rect 2548 2477 2668 2483
rect 2740 2477 2844 2483
rect 2964 2477 3004 2483
rect 3028 2477 3052 2483
rect 3076 2477 3084 2483
rect 3124 2477 3132 2483
rect 3156 2477 3660 2483
rect 3732 2477 3772 2483
rect 3812 2477 3868 2483
rect 4148 2477 4396 2483
rect 4468 2477 4556 2483
rect 4685 2483 4691 2517
rect 4772 2517 4780 2523
rect 4900 2517 4940 2523
rect 4964 2517 4988 2523
rect 4996 2517 5036 2523
rect 4708 2497 4748 2503
rect 4788 2497 4796 2503
rect 4884 2497 4908 2503
rect 4932 2497 4956 2503
rect 4980 2497 5132 2503
rect 5140 2497 5180 2503
rect 4685 2477 4700 2483
rect 4820 2477 4956 2483
rect 4964 2477 4972 2483
rect 5060 2477 5068 2483
rect 388 2457 1244 2463
rect 1252 2457 1404 2463
rect 1556 2457 1564 2463
rect 1588 2457 1836 2463
rect 1940 2457 2252 2463
rect 2260 2457 2428 2463
rect 2436 2457 3980 2463
rect 4100 2457 4716 2463
rect 628 2437 1660 2443
rect 1876 2437 1948 2443
rect 2020 2437 2028 2443
rect 2436 2437 2604 2443
rect 2676 2437 2780 2443
rect 2820 2437 2940 2443
rect 2980 2437 3020 2443
rect 3140 2437 3148 2443
rect 3204 2437 3292 2443
rect 3332 2437 3340 2443
rect 3364 2437 3372 2443
rect 3748 2437 4076 2443
rect 4516 2437 4828 2443
rect 564 2417 620 2423
rect 804 2417 972 2423
rect 1012 2417 1187 2423
rect 292 2397 540 2403
rect 628 2397 636 2403
rect 820 2397 1132 2403
rect 1181 2403 1187 2417
rect 1268 2417 1340 2423
rect 1524 2417 2396 2423
rect 2404 2417 2444 2423
rect 2676 2417 2739 2423
rect 1181 2397 1324 2403
rect 1444 2397 1660 2403
rect 1812 2397 1868 2403
rect 2052 2397 2332 2403
rect 2356 2397 2412 2403
rect 2452 2397 2540 2403
rect 2708 2397 2716 2403
rect 2733 2403 2739 2417
rect 2756 2417 2796 2423
rect 2852 2417 3244 2423
rect 3284 2417 3804 2423
rect 3876 2417 3996 2423
rect 4020 2417 4028 2423
rect 4084 2417 4268 2423
rect 4372 2417 4732 2423
rect 4756 2417 4860 2423
rect 2733 2397 2787 2403
rect 372 2377 460 2383
rect 548 2377 1436 2383
rect 1444 2377 2508 2383
rect 2612 2377 2764 2383
rect 2781 2383 2787 2397
rect 2804 2397 3020 2403
rect 3028 2397 3292 2403
rect 3620 2397 4252 2403
rect 2781 2377 3228 2383
rect 3252 2377 3436 2383
rect 3588 2377 4012 2383
rect 4068 2377 4076 2383
rect 4244 2377 4732 2383
rect 4740 2377 4812 2383
rect 308 2357 860 2363
rect 868 2357 1916 2363
rect 1924 2357 2044 2363
rect 2052 2357 2220 2363
rect 2244 2357 2300 2363
rect 2324 2357 2652 2363
rect 2708 2357 3052 2363
rect 3060 2357 3164 2363
rect 3172 2357 3612 2363
rect 3940 2357 4700 2363
rect 4948 2357 5036 2363
rect 516 2337 572 2343
rect 612 2337 620 2343
rect 772 2337 1020 2343
rect 1284 2337 1340 2343
rect 1364 2337 1404 2343
rect 1508 2337 1532 2343
rect 1556 2337 1580 2343
rect 1652 2337 1756 2343
rect 1796 2337 2412 2343
rect 2500 2337 2684 2343
rect 2708 2337 2748 2343
rect 2788 2337 2860 2343
rect 2996 2337 3100 2343
rect 3348 2337 3372 2343
rect 3380 2337 3388 2343
rect 3476 2337 3500 2343
rect 3524 2337 3580 2343
rect 3732 2337 3916 2343
rect 4004 2337 4140 2343
rect 4260 2337 4316 2343
rect 4436 2337 4732 2343
rect 4932 2337 5036 2343
rect 308 2317 348 2323
rect 468 2317 700 2323
rect 836 2317 844 2323
rect 852 2317 988 2323
rect 1044 2317 1100 2323
rect 1140 2317 1164 2323
rect 1236 2317 1331 2323
rect 13 2304 19 2316
rect 68 2297 412 2303
rect 436 2297 476 2303
rect 500 2297 508 2303
rect 580 2297 780 2303
rect 916 2297 1052 2303
rect 1108 2297 1212 2303
rect 1236 2297 1276 2303
rect 1300 2297 1308 2303
rect 1325 2303 1331 2317
rect 1348 2317 1580 2323
rect 1636 2317 1676 2323
rect 1844 2317 1852 2323
rect 1908 2317 1916 2323
rect 2068 2317 2316 2323
rect 2420 2317 2476 2323
rect 2484 2317 2956 2323
rect 2980 2317 3020 2323
rect 3364 2317 3580 2323
rect 3636 2317 3660 2323
rect 3700 2317 3740 2323
rect 3780 2317 3916 2323
rect 4100 2317 4108 2323
rect 4148 2317 4524 2323
rect 4644 2317 4652 2323
rect 4804 2317 4860 2323
rect 4900 2317 5180 2323
rect 1741 2304 1747 2316
rect 3037 2304 3043 2316
rect 3357 2304 3363 2316
rect 1325 2297 1404 2303
rect 1444 2297 1452 2303
rect 1476 2297 1516 2303
rect 1604 2297 1644 2303
rect 1876 2297 1916 2303
rect 2132 2297 2156 2303
rect 2180 2297 2220 2303
rect 2244 2297 2252 2303
rect 2452 2297 2460 2303
rect 2564 2297 2572 2303
rect 2596 2297 2780 2303
rect 2836 2297 2860 2303
rect 52 2277 364 2283
rect 372 2277 684 2283
rect 692 2277 796 2283
rect 804 2277 844 2283
rect 861 2277 867 2296
rect 916 2277 924 2283
rect 980 2277 988 2283
rect 1028 2277 1036 2283
rect 1060 2277 1244 2283
rect 1316 2277 1564 2283
rect 1588 2277 1820 2283
rect 1828 2277 1964 2283
rect 2004 2277 2012 2283
rect 2084 2277 2108 2283
rect 2132 2277 2236 2283
rect 2372 2277 2396 2283
rect 2452 2277 2492 2283
rect 2525 2277 2531 2296
rect 2797 2284 2803 2296
rect 2877 2284 2883 2303
rect 2948 2297 3020 2303
rect 3092 2297 3148 2303
rect 3220 2297 3228 2303
rect 3300 2297 3324 2303
rect 3412 2297 3548 2303
rect 3556 2297 4236 2303
rect 4244 2297 4252 2303
rect 4292 2297 4844 2303
rect 4852 2297 5004 2303
rect 5140 2297 5148 2303
rect 2580 2277 2588 2283
rect 2612 2277 2748 2283
rect 2756 2277 2764 2283
rect 2820 2277 2844 2283
rect 2916 2277 2940 2283
rect 3028 2277 3036 2283
rect 3092 2277 3132 2283
rect 3140 2277 3548 2283
rect 3588 2277 3596 2283
rect 3684 2277 3708 2283
rect 3844 2277 3884 2283
rect 3940 2277 4028 2283
rect 4036 2277 4156 2283
rect 4164 2277 4220 2283
rect 4244 2277 4268 2283
rect 4436 2277 4476 2283
rect 4548 2277 4556 2283
rect 4596 2277 4620 2283
rect 4644 2277 4652 2283
rect 4740 2277 4764 2283
rect 4836 2277 4892 2283
rect 4980 2277 4995 2283
rect 4989 2264 4995 2277
rect 5044 2277 5084 2283
rect 5149 2264 5155 2276
rect 36 2257 60 2263
rect 148 2257 172 2263
rect 196 2257 204 2263
rect 228 2257 300 2263
rect 340 2257 348 2263
rect 452 2257 460 2263
rect 477 2244 483 2263
rect 644 2257 652 2263
rect 852 2257 1580 2263
rect 1620 2257 1628 2263
rect 1732 2257 1804 2263
rect 1812 2257 1852 2263
rect 1876 2257 1884 2263
rect 1892 2257 3180 2263
rect 3220 2257 3260 2263
rect 3396 2257 3404 2263
rect 3325 2244 3331 2256
rect 3469 2244 3475 2263
rect 3796 2257 3804 2263
rect 3876 2257 3948 2263
rect 3972 2257 3980 2263
rect 4084 2257 4092 2263
rect 4196 2257 4268 2263
rect 4276 2257 4316 2263
rect 4340 2257 4652 2263
rect 4692 2257 4796 2263
rect 4868 2257 4924 2263
rect 3581 2244 3587 2256
rect 516 2237 540 2243
rect 612 2237 668 2243
rect 836 2237 1340 2243
rect 1348 2237 1420 2243
rect 1444 2237 1516 2243
rect 1572 2237 1628 2243
rect 1796 2237 1836 2243
rect 1860 2237 1900 2243
rect 1956 2237 2012 2243
rect 2052 2237 2300 2243
rect 2356 2237 2444 2243
rect 2484 2237 2572 2243
rect 2596 2237 3116 2243
rect 3268 2237 3308 2243
rect 3396 2237 3404 2243
rect 3492 2237 3564 2243
rect 3780 2237 3996 2243
rect 4084 2237 4140 2243
rect 4180 2237 4268 2243
rect 4372 2237 4764 2243
rect 4829 2237 4972 2243
rect 3661 2224 3667 2236
rect 388 2217 556 2223
rect 676 2217 956 2223
rect 1108 2217 1132 2223
rect 1172 2217 1708 2223
rect 1828 2217 1836 2223
rect 1860 2217 1884 2223
rect 1988 2217 2092 2223
rect 2180 2217 2204 2223
rect 2228 2217 2268 2223
rect 2388 2217 2396 2223
rect 2420 2217 2579 2223
rect 276 2197 284 2203
rect 644 2197 668 2203
rect 756 2197 940 2203
rect 980 2197 1228 2203
rect 1252 2197 1276 2203
rect 1524 2197 1532 2203
rect 1588 2197 1612 2203
rect 1636 2197 1756 2203
rect 1796 2197 1916 2203
rect 1988 2197 2076 2203
rect 2116 2197 2188 2203
rect 2244 2197 2252 2203
rect 2260 2197 2492 2203
rect 2573 2203 2579 2217
rect 2596 2217 2620 2223
rect 2676 2217 2700 2223
rect 2740 2217 2748 2223
rect 2804 2217 2844 2223
rect 2900 2217 2972 2223
rect 2996 2217 3004 2223
rect 3028 2217 3068 2223
rect 3316 2217 3324 2223
rect 3364 2217 3388 2223
rect 3396 2217 3564 2223
rect 3796 2217 3868 2223
rect 3924 2217 3932 2223
rect 3956 2217 4044 2223
rect 4205 2217 4380 2223
rect 4093 2204 4099 2216
rect 2573 2197 2828 2203
rect 2852 2197 2892 2203
rect 2948 2197 3420 2203
rect 3428 2197 3628 2203
rect 3636 2197 3788 2203
rect 3796 2197 3980 2203
rect 4205 2203 4211 2217
rect 4404 2217 4412 2223
rect 4484 2217 4508 2223
rect 4644 2217 4780 2223
rect 4829 2223 4835 2237
rect 5133 2243 5139 2256
rect 5133 2237 5148 2243
rect 4804 2217 4835 2223
rect 4884 2217 4956 2223
rect 4980 2217 5116 2223
rect 4132 2197 4211 2203
rect 4228 2197 4380 2203
rect 4420 2197 4444 2203
rect 4500 2197 4524 2203
rect 4596 2197 4636 2203
rect 4772 2197 4844 2203
rect 4884 2197 4892 2203
rect 5012 2197 5036 2203
rect 5060 2197 5267 2203
rect 244 2177 348 2183
rect 676 2177 684 2183
rect 724 2177 844 2183
rect 900 2177 1164 2183
rect 1172 2177 1740 2183
rect 1764 2177 1772 2183
rect 1780 2177 2508 2183
rect 2564 2177 2700 2183
rect 2756 2177 3148 2183
rect 3204 2177 3292 2183
rect 3364 2177 3404 2183
rect 3412 2177 4060 2183
rect 4068 2177 4332 2183
rect 4340 2177 4604 2183
rect 4724 2177 4780 2183
rect 4884 2177 5100 2183
rect 5261 2177 5267 2197
rect 61 2164 67 2176
rect 173 2157 179 2176
rect 3341 2164 3347 2176
rect 196 2157 220 2163
rect 260 2157 380 2163
rect 468 2157 604 2163
rect 628 2157 748 2163
rect 804 2157 844 2163
rect 948 2157 1116 2163
rect 1140 2157 1148 2163
rect 1220 2157 1260 2163
rect 1300 2157 1324 2163
rect 1348 2157 1356 2163
rect 1380 2157 1468 2163
rect 1524 2157 1564 2163
rect 1604 2157 1612 2163
rect 1636 2157 1644 2163
rect 1668 2157 1692 2163
rect 1716 2157 1724 2163
rect 1748 2157 1804 2163
rect 1812 2157 2572 2163
rect 2612 2157 2652 2163
rect 2676 2157 3340 2163
rect 3364 2157 3452 2163
rect 3460 2157 3516 2163
rect 3556 2157 3692 2163
rect 3716 2157 3740 2163
rect 3764 2157 3980 2163
rect 4020 2157 4028 2163
rect 4052 2157 4108 2163
rect 4148 2157 4204 2163
rect 4260 2157 4268 2163
rect 4308 2157 4316 2163
rect 4324 2157 4332 2163
rect 4356 2157 4604 2163
rect 4708 2157 4748 2163
rect 5060 2157 5100 2163
rect 5021 2144 5027 2156
rect -51 2137 12 2143
rect 52 2137 92 2143
rect 292 2137 316 2143
rect 324 2137 956 2143
rect 964 2137 1308 2143
rect 1316 2137 1996 2143
rect 2036 2137 2044 2143
rect 2068 2137 2140 2143
rect 2196 2137 2204 2143
rect 2221 2137 2460 2143
rect 100 2117 316 2123
rect 436 2117 444 2123
rect 500 2117 508 2123
rect 516 2117 796 2123
rect 948 2117 988 2123
rect 996 2117 1004 2123
rect 1044 2117 1052 2123
rect 1108 2117 1171 2123
rect 292 2097 300 2103
rect 308 2097 428 2103
rect 484 2097 572 2103
rect 596 2097 732 2103
rect 756 2097 764 2103
rect 1092 2097 1100 2103
rect 1165 2103 1171 2117
rect 1188 2117 1308 2123
rect 1316 2117 1868 2123
rect 1988 2117 2076 2123
rect 2084 2117 2156 2123
rect 2221 2123 2227 2137
rect 2500 2137 2844 2143
rect 2884 2137 3148 2143
rect 3188 2137 3196 2143
rect 3252 2137 3260 2143
rect 3268 2137 4284 2143
rect 4292 2137 4748 2143
rect 4756 2137 4796 2143
rect 4868 2137 4892 2143
rect 5060 2137 5116 2143
rect 2196 2117 2227 2123
rect 2276 2117 2284 2123
rect 2477 2117 2483 2136
rect 2861 2124 2867 2136
rect 4829 2124 4835 2136
rect 4941 2124 4947 2136
rect 2532 2117 2572 2123
rect 2660 2117 2668 2123
rect 2676 2117 2796 2123
rect 2836 2117 2844 2123
rect 2900 2117 2940 2123
rect 2980 2117 3004 2123
rect 3028 2117 3068 2123
rect 3124 2117 3132 2123
rect 3300 2117 3436 2123
rect 3460 2117 3468 2123
rect 3492 2117 3548 2123
rect 3604 2117 3660 2123
rect 3700 2117 3708 2123
rect 3732 2117 4204 2123
rect 4244 2117 4252 2123
rect 4356 2117 4412 2123
rect 4436 2117 4444 2123
rect 4468 2117 4476 2123
rect 4500 2117 4508 2123
rect 4548 2117 4556 2123
rect 4596 2117 4604 2123
rect 4644 2117 4652 2123
rect 4788 2117 4828 2123
rect 4948 2117 4988 2123
rect 5060 2117 5068 2123
rect 2381 2104 2387 2116
rect 3277 2104 3283 2116
rect 1165 2097 1340 2103
rect 1364 2097 1372 2103
rect 1492 2097 1500 2103
rect 1508 2097 2028 2103
rect 2036 2097 2236 2103
rect 2244 2097 2252 2103
rect 2420 2097 2492 2103
rect 2516 2097 2812 2103
rect 2820 2097 3244 2103
rect 3300 2097 3388 2103
rect 3476 2097 3500 2103
rect 3540 2097 3644 2103
rect 3668 2097 3692 2103
rect 3716 2097 3948 2103
rect 3956 2097 4076 2103
rect 4100 2097 4156 2103
rect 4180 2097 4188 2103
rect 4452 2097 4668 2103
rect 4676 2097 4700 2103
rect 5012 2097 5164 2103
rect 164 2077 460 2083
rect 468 2077 1596 2083
rect 1652 2077 1820 2083
rect 1844 2077 1852 2083
rect 1908 2077 1948 2083
rect 1956 2077 1980 2083
rect 2068 2077 2076 2083
rect 2100 2077 2332 2083
rect 2340 2077 2620 2083
rect 2644 2077 2668 2083
rect 2692 2077 2940 2083
rect 2980 2077 3740 2083
rect 3748 2077 4060 2083
rect 4068 2077 4396 2083
rect 4484 2077 4492 2083
rect 4564 2077 4684 2083
rect 4852 2077 4892 2083
rect 5012 2077 5116 2083
rect 388 2057 396 2063
rect 564 2057 604 2063
rect 660 2057 748 2063
rect 868 2057 1036 2063
rect 1044 2057 1484 2063
rect 1492 2057 1516 2063
rect 1613 2057 1628 2063
rect 1684 2057 1724 2063
rect 1748 2057 1788 2063
rect 1892 2057 1932 2063
rect 1972 2057 2012 2063
rect 2036 2057 2044 2063
rect 2068 2057 2092 2063
rect 2116 2057 2172 2063
rect 2452 2057 2732 2063
rect 2756 2057 2796 2063
rect 2836 2057 2844 2063
rect 2884 2057 2940 2063
rect 2964 2057 3820 2063
rect 3876 2057 3884 2063
rect 4004 2057 4092 2063
rect 4836 2057 5100 2063
rect 5124 2057 5148 2063
rect 1140 2037 1276 2043
rect 1284 2037 1420 2043
rect 1540 2037 1548 2043
rect 1700 2037 2124 2043
rect 2148 2037 2396 2043
rect 2420 2037 2460 2043
rect 2484 2037 3004 2043
rect 3012 2037 3340 2043
rect 3460 2037 3468 2043
rect 3636 2037 3644 2043
rect 3668 2037 3708 2043
rect 3732 2037 3772 2043
rect 4068 2037 4092 2043
rect 4452 2037 4780 2043
rect 3869 2024 3875 2036
rect 820 2017 828 2023
rect 1156 2017 1164 2023
rect 1204 2017 1244 2023
rect 1284 2017 1708 2023
rect 1716 2017 2060 2023
rect 2116 2017 2124 2023
rect 2148 2017 2172 2023
rect 2452 2017 2524 2023
rect 2564 2017 2604 2023
rect 2628 2017 2652 2023
rect 2724 2017 2892 2023
rect 2916 2017 2924 2023
rect 2948 2017 3036 2023
rect 3060 2017 3068 2023
rect 3140 2017 3148 2023
rect 3284 2017 3292 2023
rect 3444 2017 3468 2023
rect 3524 2017 3532 2023
rect 3604 2017 3740 2023
rect 3940 2017 4364 2023
rect 4516 2017 4556 2023
rect 4772 2017 5068 2023
rect 196 1997 412 2003
rect 420 1997 732 2003
rect 836 1997 844 2003
rect 852 1997 1020 2003
rect 1028 1997 1116 2003
rect 1124 1997 1276 2003
rect 1284 1997 1388 2003
rect 1396 1997 1900 2003
rect 1908 1997 2284 2003
rect 2292 1997 4044 2003
rect 4068 1997 4140 2003
rect 4980 1997 5084 2003
rect 804 1977 844 1983
rect 868 1977 908 1983
rect 916 1977 1756 1983
rect 1780 1977 1868 1983
rect 1924 1977 2876 1983
rect 2948 1977 3148 1983
rect 3332 1977 3404 1983
rect 3476 1977 3564 1983
rect 3588 1977 3612 1983
rect 3636 1977 3676 1983
rect 3924 1977 3980 1983
rect 4036 1977 4044 1983
rect 4420 1977 4444 1983
rect 4548 1977 4588 1983
rect 4772 1977 4876 1983
rect 5044 1977 5084 1983
rect 484 1957 492 1963
rect 916 1957 931 1963
rect 980 1957 1228 1963
rect 1268 1957 1356 1963
rect 1476 1957 1564 1963
rect 1572 1957 1852 1963
rect 1860 1957 2412 1963
rect 2484 1957 2556 1963
rect 2580 1957 2588 1963
rect 2612 1957 2652 1963
rect 2756 1957 2764 1963
rect 2820 1957 2876 1963
rect 2900 1957 3004 1963
rect 3060 1957 3132 1963
rect 3204 1957 3212 1963
rect 3252 1957 3724 1963
rect 3764 1957 3788 1963
rect 3924 1957 3932 1963
rect 4212 1957 4252 1963
rect 4301 1963 4307 1976
rect 4292 1957 4307 1963
rect 4356 1957 4428 1963
rect 4564 1957 4860 1963
rect 5108 1957 5132 1963
rect 5156 1957 5164 1963
rect 500 1937 732 1943
rect 740 1937 780 1943
rect 788 1937 1724 1943
rect 1732 1937 2188 1943
rect 2196 1937 2204 1943
rect 2228 1937 2268 1943
rect 2324 1937 3244 1943
rect 3252 1937 3404 1943
rect 3412 1937 3452 1943
rect 3476 1937 3836 1943
rect 3844 1937 4252 1943
rect 4260 1937 4300 1943
rect 4356 1937 4636 1943
rect 4660 1937 4748 1943
rect 148 1917 188 1923
rect 372 1917 396 1923
rect 564 1917 572 1923
rect 644 1917 668 1923
rect 692 1917 764 1923
rect 1060 1917 1164 1923
rect 1220 1917 1260 1923
rect 1341 1904 1347 1923
rect 1508 1917 1676 1923
rect 1684 1917 1692 1923
rect 1748 1917 1804 1923
rect 1860 1917 1868 1923
rect 1892 1917 1900 1923
rect 1940 1917 1948 1923
rect 2052 1917 2076 1923
rect 2093 1917 2588 1923
rect 1437 1904 1443 1916
rect 1821 1904 1827 1916
rect 100 1897 188 1903
rect 436 1897 531 1903
rect 381 1884 387 1896
rect 52 1877 348 1883
rect 397 1877 476 1883
rect 180 1857 188 1863
rect 308 1857 316 1863
rect 397 1863 403 1877
rect 525 1883 531 1897
rect 548 1897 588 1903
rect 788 1897 828 1903
rect 836 1897 860 1903
rect 900 1897 908 1903
rect 932 1897 988 1903
rect 996 1897 1036 1903
rect 1060 1897 1116 1903
rect 1364 1897 1404 1903
rect 1524 1897 1532 1903
rect 1556 1897 1564 1903
rect 1604 1897 1612 1903
rect 1636 1897 1724 1903
rect 1780 1897 1788 1903
rect 2093 1903 2099 1917
rect 2692 1917 2716 1923
rect 2740 1917 2940 1923
rect 2980 1917 3004 1923
rect 3044 1917 3180 1923
rect 3188 1917 3548 1923
rect 3556 1917 3772 1923
rect 3780 1917 3964 1923
rect 4004 1917 4012 1923
rect 4084 1917 4588 1923
rect 4596 1917 4604 1923
rect 4628 1917 4732 1923
rect 5108 1917 5267 1923
rect 2637 1904 2643 1916
rect 1860 1897 2099 1903
rect 2196 1897 2236 1903
rect 2308 1897 2508 1903
rect 2532 1897 2572 1903
rect 2708 1897 2716 1903
rect 2756 1897 2764 1903
rect 2868 1897 2876 1903
rect 2916 1897 2924 1903
rect 2948 1897 2956 1903
rect 2964 1897 3020 1903
rect 3060 1897 3164 1903
rect 3188 1897 3212 1903
rect 3300 1897 3468 1903
rect 3572 1897 3580 1903
rect 3604 1897 3628 1903
rect 3652 1897 3660 1903
rect 3668 1897 4220 1903
rect 4228 1897 4284 1903
rect 4308 1897 4316 1903
rect 4420 1897 4492 1903
rect 4868 1897 4892 1903
rect 4900 1897 4972 1903
rect 4980 1897 5116 1903
rect 525 1877 604 1883
rect 644 1877 684 1883
rect 804 1877 988 1883
rect 996 1877 1100 1883
rect 1108 1877 1788 1883
rect 1796 1877 2556 1883
rect 2564 1877 3500 1883
rect 3540 1877 3564 1883
rect 3604 1877 4540 1883
rect 4676 1877 4828 1883
rect 4868 1877 4876 1883
rect 5060 1877 5084 1883
rect 5124 1877 5148 1883
rect 372 1857 403 1863
rect 452 1857 460 1863
rect 708 1857 796 1863
rect 852 1857 876 1863
rect 916 1857 1052 1863
rect 1060 1857 1228 1863
rect 1252 1857 1324 1863
rect 1348 1857 2316 1863
rect 2340 1857 2364 1863
rect 2372 1857 3260 1863
rect 3268 1857 3484 1863
rect 3492 1857 3676 1863
rect 3732 1857 3747 1863
rect 269 1844 275 1856
rect 3741 1844 3747 1857
rect 3796 1857 3836 1863
rect 3876 1857 3884 1863
rect 3956 1857 4076 1863
rect 4100 1857 4108 1863
rect 4116 1857 4268 1863
rect 4372 1857 4444 1863
rect 4580 1857 4636 1863
rect 4644 1857 4652 1863
rect 4692 1857 4940 1863
rect 4996 1857 5052 1863
rect 4365 1844 4371 1856
rect 20 1837 60 1843
rect 340 1837 348 1843
rect 420 1837 1036 1843
rect 1060 1837 1100 1843
rect 1300 1837 1372 1843
rect 1412 1837 1516 1843
rect 1524 1837 1532 1843
rect 1604 1837 1612 1843
rect 1636 1837 1644 1843
rect 1652 1837 1820 1843
rect 1940 1837 2060 1843
rect 2125 1837 2140 1843
rect 1117 1824 1123 1836
rect 84 1817 956 1823
rect 1508 1817 1516 1823
rect 1540 1817 1564 1823
rect 1604 1817 1692 1823
rect 1764 1817 1772 1823
rect 1876 1817 1900 1823
rect 1972 1817 1980 1823
rect 2125 1823 2131 1837
rect 2340 1837 2348 1843
rect 2356 1837 3084 1843
rect 3236 1837 3260 1843
rect 3300 1837 3308 1843
rect 3348 1837 3372 1843
rect 3396 1837 3404 1843
rect 3476 1837 3500 1843
rect 3524 1837 3692 1843
rect 3876 1837 4348 1843
rect 4404 1837 4412 1843
rect 4484 1837 4572 1843
rect 4788 1837 4796 1843
rect 4852 1837 4860 1843
rect 4884 1837 4892 1843
rect 2020 1817 2131 1823
rect 2164 1817 2172 1823
rect 2196 1817 2444 1823
rect 2468 1817 2476 1823
rect 2516 1817 2540 1823
rect 2564 1817 2700 1823
rect 2772 1817 2860 1823
rect 2884 1817 2892 1823
rect 2916 1817 2947 1823
rect 1277 1804 1283 1816
rect 132 1797 172 1803
rect 180 1797 380 1803
rect 452 1797 460 1803
rect 772 1797 1036 1803
rect 1172 1797 1196 1803
rect 1524 1797 2092 1803
rect 2100 1797 2108 1803
rect 2132 1797 2556 1803
rect 2628 1797 2636 1803
rect 2724 1797 2748 1803
rect 2788 1797 2796 1803
rect 2836 1797 2892 1803
rect 2916 1797 2924 1803
rect 2941 1803 2947 1817
rect 2964 1817 2972 1823
rect 2996 1817 3004 1823
rect 3044 1817 3068 1823
rect 3076 1817 3100 1823
rect 3172 1817 3324 1823
rect 3364 1817 3596 1823
rect 3604 1817 3772 1823
rect 3780 1817 4412 1823
rect 4836 1817 4876 1823
rect 2941 1797 2956 1803
rect 2996 1797 3116 1803
rect 3156 1797 3196 1803
rect 3220 1797 3244 1803
rect 3348 1797 3356 1803
rect 3428 1797 3868 1803
rect 3956 1797 3964 1803
rect 4004 1797 4028 1803
rect 4045 1797 4172 1803
rect 1117 1784 1123 1796
rect 404 1777 476 1783
rect 516 1777 524 1783
rect 612 1777 652 1783
rect 740 1777 892 1783
rect 932 1777 1004 1783
rect 1124 1777 1308 1783
rect 1348 1777 1596 1783
rect 1636 1777 1644 1783
rect 1661 1777 1923 1783
rect 1325 1764 1331 1776
rect 148 1757 156 1763
rect 228 1757 604 1763
rect 612 1757 732 1763
rect 788 1757 844 1763
rect 932 1757 1228 1763
rect 1252 1757 1292 1763
rect 1508 1757 1516 1763
rect 1556 1757 1564 1763
rect 1661 1763 1667 1777
rect 1572 1757 1667 1763
rect 1684 1757 1692 1763
rect 1748 1757 1756 1763
rect 1828 1757 1884 1763
rect 1917 1763 1923 1777
rect 1940 1777 2380 1783
rect 2452 1777 2940 1783
rect 2948 1777 2956 1783
rect 2996 1777 3004 1783
rect 3108 1777 3500 1783
rect 3556 1777 3724 1783
rect 3748 1777 3756 1783
rect 3764 1777 3932 1783
rect 3972 1777 3980 1783
rect 4045 1783 4051 1797
rect 4196 1797 4220 1803
rect 4692 1797 4924 1803
rect 5076 1797 5084 1803
rect 4004 1777 4051 1783
rect 4084 1777 4364 1783
rect 4452 1777 4460 1783
rect 4500 1777 4588 1783
rect 4692 1777 4764 1783
rect 4804 1777 5100 1783
rect 5124 1777 5155 1783
rect 5149 1764 5155 1777
rect 1917 1757 1964 1763
rect 1988 1757 2012 1763
rect 2036 1757 2140 1763
rect 2180 1757 2236 1763
rect 2276 1757 2284 1763
rect 2324 1757 3452 1763
rect 3460 1757 3468 1763
rect 3492 1757 3500 1763
rect 3524 1757 3532 1763
rect 3620 1757 3628 1763
rect 3636 1757 3692 1763
rect 3821 1757 3884 1763
rect 212 1737 236 1743
rect 260 1737 332 1743
rect 372 1737 396 1743
rect 420 1737 444 1743
rect 500 1737 540 1743
rect 596 1737 796 1743
rect 804 1737 892 1743
rect 900 1737 1340 1743
rect 1389 1737 1395 1756
rect 1789 1744 1795 1756
rect 3725 1744 3731 1756
rect 3741 1744 3747 1756
rect 1508 1737 1708 1743
rect 1748 1737 1756 1743
rect 1876 1737 1916 1743
rect 1956 1737 2028 1743
rect 2132 1737 2188 1743
rect 2212 1737 2220 1743
rect 2244 1737 2588 1743
rect 2596 1737 3052 1743
rect 3076 1737 3180 1743
rect 3188 1737 3596 1743
rect 3636 1737 3660 1743
rect 3684 1737 3708 1743
rect 3764 1737 3788 1743
rect 3821 1743 3827 1757
rect 3924 1757 3948 1763
rect 4068 1757 4076 1763
rect 4084 1757 4124 1763
rect 4148 1757 4316 1763
rect 4340 1757 4876 1763
rect 4884 1757 4988 1763
rect 5028 1757 5116 1763
rect 3805 1737 3827 1743
rect 68 1717 108 1723
rect 260 1717 268 1723
rect 276 1717 492 1723
rect 676 1717 796 1723
rect 836 1717 844 1723
rect 1092 1717 1260 1723
rect 1300 1717 1340 1723
rect 1364 1717 1980 1723
rect 2020 1717 2524 1723
rect 2548 1717 2588 1723
rect 2660 1717 2684 1723
rect 2708 1717 2716 1723
rect 2788 1717 2803 1723
rect 292 1697 348 1703
rect 356 1697 412 1703
rect 484 1697 572 1703
rect 708 1697 828 1703
rect 852 1697 940 1703
rect 996 1697 1100 1703
rect 1220 1697 1228 1703
rect 1284 1697 1436 1703
rect 1460 1697 1788 1703
rect 1828 1697 1836 1703
rect 1924 1697 2252 1703
rect 2260 1697 2268 1703
rect 2292 1697 2364 1703
rect 2404 1697 2412 1703
rect 2452 1697 2476 1703
rect 2500 1697 2540 1703
rect 2580 1697 2588 1703
rect 2644 1697 2732 1703
rect 2749 1697 2755 1716
rect 2797 1704 2803 1717
rect 2900 1717 2908 1723
rect 3028 1717 3132 1723
rect 3172 1717 3260 1723
rect 3277 1717 3340 1723
rect 2877 1704 2883 1716
rect 2957 1704 2963 1716
rect 2900 1697 2908 1703
rect 3028 1697 3052 1703
rect 3076 1697 3212 1703
rect 3277 1703 3283 1717
rect 3364 1717 3692 1723
rect 3700 1717 3708 1723
rect 3805 1723 3811 1737
rect 3844 1737 3852 1743
rect 3876 1737 3916 1743
rect 4036 1737 4060 1743
rect 4084 1737 4092 1743
rect 4132 1737 4172 1743
rect 4228 1737 4460 1743
rect 4596 1737 4604 1743
rect 4644 1737 4652 1743
rect 4676 1737 4700 1743
rect 4788 1737 4908 1743
rect 4964 1737 4972 1743
rect 5012 1737 5020 1743
rect 5092 1737 5100 1743
rect 5133 1743 5139 1756
rect 5124 1737 5139 1743
rect 3748 1717 3811 1723
rect 3828 1717 3836 1723
rect 3844 1717 4124 1723
rect 4212 1717 4220 1723
rect 4276 1717 4316 1723
rect 4356 1717 4508 1723
rect 4660 1717 4684 1723
rect 4708 1717 5036 1723
rect 5044 1717 5068 1723
rect 5092 1717 5132 1723
rect 4125 1704 4131 1716
rect 3252 1697 3283 1703
rect 3300 1697 3308 1703
rect 3332 1697 3388 1703
rect 3444 1697 3452 1703
rect 3476 1697 3484 1703
rect 3508 1697 3644 1703
rect 3668 1697 3772 1703
rect 3860 1697 3916 1703
rect 3988 1697 4092 1703
rect 4164 1697 4220 1703
rect 4308 1697 4348 1703
rect 4356 1697 4364 1703
rect 4388 1697 4492 1703
rect 4548 1697 4796 1703
rect 4804 1697 5020 1703
rect 5092 1697 5164 1703
rect 116 1677 300 1683
rect 356 1677 364 1683
rect 532 1677 540 1683
rect 580 1677 636 1683
rect 644 1677 652 1683
rect 1284 1677 1292 1683
rect 1316 1677 1884 1683
rect 1892 1677 2140 1683
rect 2180 1677 2700 1683
rect 2708 1677 3084 1683
rect 3092 1677 3404 1683
rect 3412 1677 4204 1683
rect 4228 1677 4348 1683
rect 4388 1677 4412 1683
rect 4420 1677 4428 1683
rect 4804 1677 4844 1683
rect 4852 1677 5036 1683
rect 477 1664 483 1676
rect 612 1657 892 1663
rect 932 1657 1292 1663
rect 1524 1657 2156 1663
rect 2244 1657 2284 1663
rect 2308 1657 3020 1663
rect 3044 1657 3996 1663
rect 4100 1657 4396 1663
rect 4404 1657 4716 1663
rect 4724 1657 4796 1663
rect 4836 1657 4956 1663
rect 5012 1657 5052 1663
rect 660 1637 860 1643
rect 900 1637 956 1643
rect 1540 1637 1612 1643
rect 1716 1637 3004 1643
rect 3092 1637 3244 1643
rect 3268 1637 3708 1643
rect 3828 1637 4044 1643
rect 4196 1637 4204 1643
rect 4228 1637 4284 1643
rect 4372 1637 4524 1643
rect 4532 1637 4748 1643
rect 100 1617 124 1623
rect 276 1617 796 1623
rect 804 1617 2124 1623
rect 2148 1617 2236 1623
rect 2308 1617 2364 1623
rect 2388 1617 2924 1623
rect 2964 1617 2972 1623
rect 2996 1617 3068 1623
rect 3252 1617 3260 1623
rect 3652 1617 3772 1623
rect 3796 1617 3804 1623
rect 3876 1617 4892 1623
rect 1284 1597 1804 1603
rect 1892 1597 1916 1603
rect 1940 1597 1948 1603
rect 1956 1597 2044 1603
rect 2228 1597 2348 1603
rect 2356 1597 2739 1603
rect 228 1577 444 1583
rect 980 1577 1580 1583
rect 1604 1577 1788 1583
rect 1812 1577 1820 1583
rect 2004 1577 2188 1583
rect 2212 1577 2316 1583
rect 2340 1577 2412 1583
rect 2436 1577 2556 1583
rect 2612 1577 2668 1583
rect 2692 1577 2700 1583
rect 2733 1583 2739 1597
rect 2772 1597 2844 1603
rect 2868 1597 3084 1603
rect 3092 1597 3452 1603
rect 3540 1597 3692 1603
rect 3764 1597 3868 1603
rect 4052 1597 4060 1603
rect 4180 1597 4188 1603
rect 4196 1597 4204 1603
rect 4340 1597 4620 1603
rect 4820 1597 5068 1603
rect 2733 1577 2748 1583
rect 2772 1577 2860 1583
rect 2932 1577 2940 1583
rect 2996 1577 3004 1583
rect 3172 1577 3580 1583
rect 3588 1577 3596 1583
rect 3604 1577 4380 1583
rect 4740 1577 4764 1583
rect 4820 1577 4828 1583
rect 4852 1577 4892 1583
rect 228 1557 236 1563
rect 1204 1557 1244 1563
rect 1476 1557 1900 1563
rect 1908 1557 2092 1563
rect 2148 1557 2188 1563
rect 2244 1557 2428 1563
rect 2452 1557 2460 1563
rect 2484 1557 2508 1563
rect 2532 1557 3644 1563
rect 3652 1557 4460 1563
rect 4468 1557 4684 1563
rect 4708 1557 5020 1563
rect 5028 1557 5164 1563
rect 100 1537 284 1543
rect 292 1537 652 1543
rect 740 1537 924 1543
rect 932 1537 940 1543
rect 1060 1537 1180 1543
rect 1220 1537 1260 1543
rect 1300 1537 1404 1543
rect 1796 1537 1804 1543
rect 1812 1537 1852 1543
rect 1892 1537 1900 1543
rect 1924 1537 2188 1543
rect 2212 1537 2316 1543
rect 2324 1537 2652 1543
rect 2660 1537 2940 1543
rect 2964 1537 3100 1543
rect 3140 1537 3148 1543
rect 3220 1537 3228 1543
rect 3252 1537 3260 1543
rect 3284 1537 3292 1543
rect 3348 1537 3356 1543
rect 3380 1537 3500 1543
rect 3524 1537 3548 1543
rect 3636 1537 3660 1543
rect 3684 1537 3964 1543
rect 3972 1537 4268 1543
rect 4276 1537 4316 1543
rect 4404 1537 4412 1543
rect 4484 1537 4844 1543
rect 5092 1537 5148 1543
rect 84 1517 92 1523
rect 116 1517 124 1523
rect 196 1517 220 1523
rect 244 1517 252 1523
rect 340 1517 460 1523
rect 468 1517 556 1523
rect 596 1517 604 1523
rect 756 1517 780 1523
rect 884 1517 988 1523
rect 996 1517 1004 1523
rect 1028 1517 1116 1523
rect 1156 1517 1196 1523
rect 1252 1517 1468 1523
rect 1524 1517 1532 1523
rect 1716 1517 2172 1523
rect 2196 1517 2252 1523
rect 2308 1517 2332 1523
rect 2420 1517 2428 1523
rect 2452 1517 2572 1523
rect 2596 1517 2620 1523
rect 2628 1517 3244 1523
rect 3300 1517 3308 1523
rect 3348 1517 3404 1523
rect 3476 1517 3484 1523
rect 3572 1517 3932 1523
rect 4004 1517 4012 1523
rect 4036 1517 4060 1523
rect 4100 1517 4108 1523
rect 4132 1517 4268 1523
rect 4276 1517 4588 1523
rect 4596 1517 4940 1523
rect 5108 1517 5116 1523
rect 829 1504 835 1516
rect 1133 1504 1139 1516
rect 68 1497 204 1503
rect 244 1497 828 1503
rect 916 1497 924 1503
rect 948 1497 956 1503
rect 964 1497 1132 1503
rect 1236 1497 1372 1503
rect 1412 1497 1452 1503
rect 1460 1497 1548 1503
rect 1597 1497 1612 1503
rect 1668 1497 1740 1503
rect 1748 1497 1756 1503
rect 1780 1497 1788 1503
rect 1860 1497 1948 1503
rect 1972 1497 2044 1503
rect 2052 1497 2060 1503
rect 2068 1497 2140 1503
rect 2164 1497 2172 1503
rect 2196 1497 2444 1503
rect 2564 1497 2572 1503
rect 2596 1497 2652 1503
rect 2676 1497 2732 1503
rect 2756 1497 2780 1503
rect 2836 1497 2860 1503
rect 2884 1497 2908 1503
rect 2948 1497 3020 1503
rect 3060 1497 3580 1503
rect 3588 1497 3964 1503
rect 4004 1497 4140 1503
rect 4404 1497 4540 1503
rect 4564 1497 4604 1503
rect 4644 1497 4652 1503
rect 4692 1497 5068 1503
rect 5076 1497 5132 1503
rect -51 1477 12 1483
rect 212 1477 364 1483
rect 372 1477 620 1483
rect 756 1477 764 1483
rect 772 1477 876 1483
rect 948 1477 1564 1483
rect 1572 1477 1628 1483
rect 1652 1477 1660 1483
rect 1700 1477 1756 1483
rect 1796 1477 1804 1483
rect 1828 1477 1868 1483
rect 1876 1477 1900 1483
rect 1924 1477 1932 1483
rect 2004 1477 2012 1483
rect 2036 1477 2044 1483
rect 2100 1477 2236 1483
rect 2292 1477 2380 1483
rect 2420 1477 3532 1483
rect 3572 1477 3660 1483
rect 3844 1477 3868 1483
rect 3956 1477 4092 1483
rect 4116 1477 4156 1483
rect 4173 1477 4220 1483
rect 3805 1464 3811 1476
rect 164 1457 220 1463
rect 308 1457 316 1463
rect 356 1457 380 1463
rect 564 1457 860 1463
rect 884 1457 892 1463
rect 916 1457 972 1463
rect 1076 1457 1084 1463
rect 1092 1457 1260 1463
rect 1412 1457 1420 1463
rect 1604 1457 1612 1463
rect 1620 1457 2188 1463
rect 2244 1457 2268 1463
rect 2308 1457 2332 1463
rect 2372 1457 3628 1463
rect 3812 1457 3996 1463
rect 4052 1457 4076 1463
rect 4116 1457 4124 1463
rect 4173 1463 4179 1477
rect 4276 1477 4492 1483
rect 4500 1477 4556 1483
rect 4612 1477 4652 1483
rect 4836 1477 4924 1483
rect 4932 1477 4940 1483
rect 4996 1477 5059 1483
rect 4148 1457 4179 1463
rect 4212 1457 4220 1463
rect 4244 1457 4252 1463
rect 4276 1457 4284 1463
rect 4308 1457 4700 1463
rect 4724 1457 4748 1463
rect 4836 1457 4956 1463
rect 4973 1457 4988 1463
rect 5012 1457 5020 1463
rect 5053 1463 5059 1477
rect 5076 1477 5084 1483
rect 5140 1477 5148 1483
rect 5053 1457 5148 1463
rect 308 1437 316 1443
rect 548 1437 556 1443
rect 660 1437 684 1443
rect 948 1437 1132 1443
rect 1172 1437 2364 1443
rect 2484 1437 2524 1443
rect 2580 1437 2956 1443
rect 2964 1437 3260 1443
rect 3268 1437 3276 1443
rect 3300 1437 3308 1443
rect 3396 1437 3404 1443
rect 3476 1437 3516 1443
rect 3556 1437 4316 1443
rect 4324 1437 4412 1443
rect 4788 1437 4876 1443
rect 4980 1437 5068 1443
rect 3341 1424 3347 1436
rect 244 1417 364 1423
rect 420 1417 492 1423
rect 564 1417 572 1423
rect 1028 1417 1084 1423
rect 1092 1417 1148 1423
rect 1284 1417 1340 1423
rect 1364 1417 1388 1423
rect 1412 1417 2012 1423
rect 2020 1417 2108 1423
rect 2116 1417 2124 1423
rect 2148 1417 2220 1423
rect 2340 1417 2531 1423
rect 356 1397 364 1403
rect 388 1397 604 1403
rect 1188 1397 1244 1403
rect 1508 1397 1516 1403
rect 1556 1397 1596 1403
rect 1764 1397 1820 1403
rect 1860 1397 1932 1403
rect 2004 1397 2028 1403
rect 2148 1397 2156 1403
rect 2180 1397 2204 1403
rect 2260 1397 2284 1403
rect 2452 1397 2508 1403
rect 2525 1403 2531 1417
rect 2548 1417 2556 1423
rect 2580 1417 2588 1423
rect 2628 1417 2652 1423
rect 2676 1417 2700 1423
rect 2724 1417 2732 1423
rect 2756 1417 2796 1423
rect 2820 1417 2828 1423
rect 2868 1417 2876 1423
rect 2916 1417 3100 1423
rect 3156 1417 3164 1423
rect 3188 1417 3196 1423
rect 3588 1417 3644 1423
rect 3716 1417 3884 1423
rect 3956 1417 3980 1423
rect 4004 1417 4028 1423
rect 4052 1417 4060 1423
rect 4116 1417 4172 1423
rect 4276 1417 4380 1423
rect 2525 1397 3004 1403
rect 3076 1397 3164 1403
rect 3188 1397 3404 1403
rect 3469 1397 3596 1403
rect 1341 1384 1347 1396
rect 1645 1384 1651 1396
rect -51 1377 12 1383
rect 260 1377 380 1383
rect 452 1377 668 1383
rect 772 1377 1116 1383
rect 1124 1377 1324 1383
rect 1412 1377 1484 1383
rect 1556 1377 1564 1383
rect 1620 1377 1628 1383
rect 1700 1377 1708 1383
rect 1716 1377 2332 1383
rect 2388 1377 2572 1383
rect 2580 1377 2588 1383
rect 2660 1377 2924 1383
rect 2980 1377 2988 1383
rect 3028 1377 3068 1383
rect 3092 1377 3132 1383
rect 3204 1377 3260 1383
rect 3268 1377 3276 1383
rect 3300 1377 3340 1383
rect 3469 1383 3475 1397
rect 3620 1397 4460 1403
rect 4468 1397 4684 1403
rect 4836 1397 4876 1403
rect 3364 1377 3475 1383
rect 3492 1377 3660 1383
rect 3677 1377 3740 1383
rect 52 1357 76 1363
rect 109 1363 115 1376
rect 100 1357 115 1363
rect 164 1357 524 1363
rect 580 1357 588 1363
rect 596 1357 636 1363
rect 660 1357 668 1363
rect 788 1357 867 1363
rect 20 1337 76 1343
rect 148 1337 188 1343
rect 532 1337 668 1343
rect 708 1337 732 1343
rect 772 1337 812 1343
rect 861 1343 867 1357
rect 884 1357 972 1363
rect 1092 1357 1756 1363
rect 1764 1357 1852 1363
rect 1869 1357 1884 1363
rect 1924 1357 2044 1363
rect 2068 1357 2076 1363
rect 2100 1357 2115 1363
rect 2164 1357 2172 1363
rect 2244 1357 2252 1363
rect 2340 1357 2364 1363
rect 2420 1357 2652 1363
rect 2692 1357 2748 1363
rect 2884 1357 2908 1363
rect 2948 1357 3356 1363
rect 3380 1357 3500 1363
rect 3588 1357 3596 1363
rect 3677 1363 3683 1377
rect 3764 1377 3820 1383
rect 3908 1377 3955 1383
rect 3620 1357 3683 1363
rect 3716 1357 3724 1363
rect 3748 1357 3772 1363
rect 3844 1357 3852 1363
rect 3892 1357 3932 1363
rect 3949 1363 3955 1377
rect 3972 1377 4460 1383
rect 4468 1377 4732 1383
rect 4772 1377 5020 1383
rect 3949 1357 4028 1363
rect 4068 1357 4204 1363
rect 4276 1357 4284 1363
rect 4372 1357 4380 1363
rect 4404 1357 4412 1363
rect 4500 1357 4508 1363
rect 4580 1357 4604 1363
rect 4644 1357 4700 1363
rect 4724 1357 4828 1363
rect 4836 1357 4844 1363
rect 4868 1357 4972 1363
rect 2813 1344 2819 1356
rect 4045 1344 4051 1356
rect 5149 1344 5155 1356
rect 861 1337 892 1343
rect 948 1337 972 1343
rect 1028 1337 1036 1343
rect 1124 1337 1171 1343
rect 493 1324 499 1336
rect 132 1317 156 1323
rect 292 1317 332 1323
rect 516 1317 588 1323
rect 628 1317 652 1323
rect 676 1317 684 1323
rect 692 1317 844 1323
rect 868 1317 876 1323
rect 884 1317 1148 1323
rect 1165 1323 1171 1337
rect 1188 1337 1212 1343
rect 1220 1337 1244 1343
rect 1300 1337 1308 1343
rect 1332 1337 2300 1343
rect 2308 1337 2316 1343
rect 2340 1337 2380 1343
rect 2420 1337 2428 1343
rect 2532 1337 2588 1343
rect 2612 1337 2668 1343
rect 2692 1337 2732 1343
rect 2772 1337 2796 1343
rect 2852 1337 2892 1343
rect 2948 1337 2972 1343
rect 3012 1337 3052 1343
rect 3076 1337 3084 1343
rect 3108 1337 3228 1343
rect 3300 1337 3836 1343
rect 3892 1337 3955 1343
rect 1165 1317 1212 1323
rect 1220 1317 1468 1323
rect 1476 1317 1484 1323
rect 1508 1317 1724 1323
rect 1748 1317 1756 1323
rect 1837 1317 1852 1323
rect 1876 1317 1884 1323
rect 1908 1317 1916 1323
rect 1924 1317 2268 1323
rect 2276 1317 3660 1323
rect 3684 1317 3740 1323
rect 3780 1317 3788 1323
rect 3844 1317 3868 1323
rect 3892 1317 3900 1323
rect 3949 1323 3955 1337
rect 3972 1337 3996 1343
rect 4084 1337 4124 1343
rect 4148 1337 4380 1343
rect 4404 1337 4652 1343
rect 4660 1337 4972 1343
rect 4996 1337 5004 1343
rect 5092 1337 5100 1343
rect 4397 1324 4403 1336
rect 3949 1317 3980 1323
rect 4020 1317 4028 1323
rect 4052 1317 4124 1323
rect 4148 1317 4172 1323
rect 4196 1317 4332 1323
rect 4484 1317 4540 1323
rect 4644 1317 4652 1323
rect 4756 1317 4860 1323
rect 4445 1304 4451 1316
rect 4717 1304 4723 1316
rect 4765 1304 4771 1317
rect 5124 1317 5196 1323
rect 52 1297 60 1303
rect 276 1297 284 1303
rect 292 1297 1084 1303
rect 1124 1297 1212 1303
rect 1220 1297 1340 1303
rect 1428 1297 1484 1303
rect 1492 1297 1532 1303
rect 1812 1297 1884 1303
rect 1892 1297 1916 1303
rect 1940 1297 2076 1303
rect 2084 1297 2348 1303
rect 2436 1297 2444 1303
rect 2484 1297 2508 1303
rect 2532 1297 2604 1303
rect 2660 1297 2915 1303
rect 356 1277 764 1283
rect 772 1277 1420 1283
rect 1428 1277 1996 1283
rect 2004 1277 2636 1283
rect 2676 1277 2844 1283
rect 2909 1283 2915 1297
rect 2932 1297 2988 1303
rect 3012 1297 3036 1303
rect 3332 1297 3372 1303
rect 3444 1297 3548 1303
rect 3588 1297 3804 1303
rect 3844 1297 3948 1303
rect 3988 1297 4028 1303
rect 4052 1297 4300 1303
rect 4324 1297 4332 1303
rect 4580 1297 4588 1303
rect 4628 1297 4700 1303
rect 4804 1297 4876 1303
rect 5076 1297 5100 1303
rect 5156 1297 5164 1303
rect 2909 1277 3452 1283
rect 3508 1277 3939 1283
rect 340 1257 364 1263
rect 740 1257 780 1263
rect 1140 1257 1324 1263
rect 1332 1257 1580 1263
rect 1748 1257 1948 1263
rect 1972 1257 2028 1263
rect 2084 1257 2220 1263
rect 2324 1257 2860 1263
rect 2884 1257 3596 1263
rect 3933 1263 3939 1277
rect 4052 1277 4076 1283
rect 4084 1277 4124 1283
rect 4148 1277 4300 1283
rect 4324 1277 4348 1283
rect 4436 1277 4460 1283
rect 4564 1277 4780 1283
rect 4820 1277 4828 1283
rect 4884 1277 4924 1283
rect 5140 1277 5164 1283
rect 3933 1257 4060 1263
rect 4068 1257 4956 1263
rect 148 1237 476 1243
rect 484 1237 1324 1243
rect 1332 1237 1372 1243
rect 1588 1237 2348 1243
rect 2404 1237 2476 1243
rect 2532 1237 2748 1243
rect 2836 1237 2956 1243
rect 3044 1237 3100 1243
rect 3252 1237 3372 1243
rect 3524 1237 3628 1243
rect 3652 1237 3740 1243
rect 3748 1237 3868 1243
rect 3924 1237 4108 1243
rect 4116 1237 4348 1243
rect 2493 1224 2499 1236
rect 4525 1224 4531 1243
rect 4820 1237 4860 1243
rect 4996 1237 5004 1243
rect 388 1217 460 1223
rect 548 1217 684 1223
rect 724 1217 844 1223
rect 980 1217 1132 1223
rect 1348 1217 1500 1223
rect 1508 1217 1516 1223
rect 1524 1217 1948 1223
rect 2020 1217 2076 1223
rect 2228 1217 2284 1223
rect 2308 1217 2316 1223
rect 2404 1217 2412 1223
rect 2436 1217 2460 1223
rect 2644 1217 2652 1223
rect 2804 1217 3004 1223
rect 3028 1217 3116 1223
rect 3204 1217 3276 1223
rect 3316 1217 3340 1223
rect 3380 1217 3532 1223
rect 3796 1217 3820 1223
rect 4084 1217 4140 1223
rect 4244 1217 4252 1223
rect 3917 1204 3923 1216
rect 180 1197 204 1203
rect 420 1197 812 1203
rect 820 1197 860 1203
rect 868 1197 1436 1203
rect 1444 1197 2540 1203
rect 2548 1197 2604 1203
rect 2612 1197 2700 1203
rect 2708 1197 3324 1203
rect 3412 1197 3452 1203
rect 3636 1197 3676 1203
rect 3780 1197 3788 1203
rect 4212 1197 4668 1203
rect 708 1177 764 1183
rect 804 1177 812 1183
rect 852 1177 908 1183
rect 996 1177 1036 1183
rect 1060 1177 1740 1183
rect 1764 1177 1820 1183
rect 1844 1177 2531 1183
rect 36 1157 108 1163
rect 836 1157 1100 1163
rect 1460 1157 1484 1163
rect 1652 1157 1660 1163
rect 1876 1157 2140 1163
rect 2244 1157 2428 1163
rect 2436 1157 2508 1163
rect 2525 1163 2531 1177
rect 2548 1177 2556 1183
rect 2596 1177 2652 1183
rect 2676 1177 3020 1183
rect 3284 1177 4092 1183
rect 4148 1177 4252 1183
rect 4516 1177 4540 1183
rect 2525 1157 3004 1163
rect 3012 1157 3436 1163
rect 3444 1157 3532 1163
rect 3572 1157 3692 1163
rect 3716 1157 3740 1163
rect 3796 1157 3900 1163
rect 4004 1157 4060 1163
rect 4116 1157 4204 1163
rect 4228 1157 4284 1163
rect 5108 1157 5116 1163
rect 244 1137 636 1143
rect 644 1137 652 1143
rect 660 1137 1164 1143
rect 1188 1137 1260 1143
rect 1316 1137 1404 1143
rect 1421 1137 1427 1156
rect 1444 1137 1516 1143
rect 1540 1137 1564 1143
rect 1652 1137 1907 1143
rect 205 1123 211 1136
rect 205 1117 220 1123
rect 484 1117 492 1123
rect 516 1117 556 1123
rect 580 1117 588 1123
rect 772 1117 780 1123
rect 1124 1117 1132 1123
rect 1476 1117 1484 1123
rect 1572 1117 1580 1123
rect 1620 1117 1644 1123
rect 1652 1117 1692 1123
rect 1700 1117 1756 1123
rect 1764 1117 1884 1123
rect 1901 1123 1907 1137
rect 1972 1137 2124 1143
rect 2132 1137 2540 1143
rect 2564 1137 2924 1143
rect 3108 1137 3276 1143
rect 3316 1137 3324 1143
rect 3396 1137 3420 1143
rect 3444 1137 3628 1143
rect 3700 1137 4396 1143
rect 4404 1137 4460 1143
rect 4532 1137 4588 1143
rect 4612 1137 4732 1143
rect 5012 1137 5116 1143
rect 1901 1117 2076 1123
rect 2084 1117 2092 1123
rect 2100 1117 2108 1123
rect 2132 1117 2476 1123
rect 2564 1117 2572 1123
rect 2596 1117 2684 1123
rect 2820 1117 2860 1123
rect 2932 1117 3180 1123
rect 3220 1117 3228 1123
rect 3252 1117 4220 1123
rect 4228 1117 4300 1123
rect 4356 1117 4652 1123
rect 4660 1117 4668 1123
rect 4916 1117 4924 1123
rect 4932 1117 5068 1123
rect 1101 1104 1107 1116
rect 4317 1104 4323 1116
rect 116 1097 252 1103
rect 628 1097 716 1103
rect 900 1097 972 1103
rect 1108 1097 1612 1103
rect 1748 1097 2028 1103
rect 2036 1097 2044 1103
rect 2164 1097 2172 1103
rect 2196 1097 2220 1103
rect 2292 1097 2300 1103
rect 2388 1097 2396 1103
rect 2429 1097 2588 1103
rect 989 1084 995 1096
rect 20 1077 76 1083
rect 436 1077 524 1083
rect 628 1077 668 1083
rect 676 1077 844 1083
rect 1076 1077 1084 1083
rect 1140 1077 1148 1083
rect 1172 1077 1180 1083
rect 1204 1077 1212 1083
rect 1252 1077 1436 1083
rect 1460 1077 1500 1083
rect 2429 1083 2435 1097
rect 2628 1097 2636 1103
rect 2676 1097 2700 1103
rect 2724 1097 2732 1103
rect 2740 1097 2876 1103
rect 2884 1097 2892 1103
rect 3076 1097 3084 1103
rect 3101 1097 3164 1103
rect 1684 1077 2435 1083
rect 2468 1077 2924 1083
rect 2996 1077 3052 1083
rect 3101 1083 3107 1097
rect 3252 1097 3260 1103
rect 3284 1097 3516 1103
rect 3540 1097 3596 1103
rect 3668 1097 3772 1103
rect 3908 1097 4012 1103
rect 4020 1097 4204 1103
rect 4212 1097 4220 1103
rect 4260 1097 4268 1103
rect 4404 1097 4412 1103
rect 4452 1097 4467 1103
rect 3069 1077 3107 1083
rect 36 1057 44 1063
rect 68 1057 188 1063
rect 292 1057 380 1063
rect 516 1057 524 1063
rect 852 1057 908 1063
rect 1364 1057 1372 1063
rect 1396 1057 1724 1063
rect 1812 1057 1980 1063
rect 1988 1057 2252 1063
rect 2340 1057 2348 1063
rect 2372 1057 2380 1063
rect 2452 1057 2828 1063
rect 2868 1057 2956 1063
rect 3069 1063 3075 1077
rect 3124 1077 3148 1083
rect 3156 1077 3516 1083
rect 3556 1077 4444 1083
rect 4461 1083 4467 1097
rect 4516 1097 4940 1103
rect 4948 1097 4988 1103
rect 5076 1097 5148 1103
rect 4461 1077 4524 1083
rect 4612 1077 4636 1083
rect 4708 1077 4764 1083
rect 4836 1077 5020 1083
rect 4685 1064 4691 1076
rect 4829 1064 4835 1076
rect 3028 1057 3075 1063
rect 3092 1057 3100 1063
rect 3124 1057 3132 1063
rect 3204 1057 3500 1063
rect 3508 1057 3612 1063
rect 3636 1057 3660 1063
rect 3684 1057 3692 1063
rect 3732 1057 3740 1063
rect 3764 1057 3788 1063
rect 3924 1057 3932 1063
rect 3956 1057 4156 1063
rect 4452 1057 4684 1063
rect 4852 1057 4860 1063
rect 4932 1057 4972 1063
rect 5012 1057 5036 1063
rect 3885 1044 3891 1056
rect 52 1037 220 1043
rect 1028 1037 1228 1043
rect 1460 1037 2012 1043
rect 2084 1037 2108 1043
rect 2148 1037 2220 1043
rect 2244 1037 2332 1043
rect 2404 1037 2492 1043
rect 2516 1037 2524 1043
rect 2548 1037 2579 1043
rect 52 1017 60 1023
rect 740 1017 1116 1023
rect 1188 1017 1580 1023
rect 1684 1017 1916 1023
rect 1988 1017 1996 1023
rect 2036 1017 2108 1023
rect 2132 1017 2188 1023
rect 2212 1017 2332 1023
rect 2356 1017 2364 1023
rect 2388 1017 2524 1023
rect 2548 1017 2556 1023
rect 2573 1023 2579 1037
rect 2596 1037 2700 1043
rect 2724 1037 2876 1043
rect 2884 1037 3004 1043
rect 3060 1037 3196 1043
rect 3284 1037 3292 1043
rect 3364 1037 3372 1043
rect 3428 1037 3436 1043
rect 3524 1037 3820 1043
rect 3828 1037 3852 1043
rect 3908 1037 4236 1043
rect 4244 1037 4540 1043
rect 4548 1037 4716 1043
rect 4724 1037 4892 1043
rect 4900 1037 5004 1043
rect 5197 1024 5203 1036
rect 2573 1017 2780 1023
rect 2820 1017 2828 1023
rect 3012 1017 3308 1023
rect 3316 1017 3452 1023
rect 3492 1017 3612 1023
rect 3636 1017 3660 1023
rect 3716 1017 3724 1023
rect 3732 1017 3836 1023
rect 3860 1017 3884 1023
rect 4052 1017 4108 1023
rect 4132 1017 4172 1023
rect 4404 1017 4508 1023
rect 4596 1017 4620 1023
rect 4644 1017 4828 1023
rect 4884 1017 4956 1023
rect 1645 1004 1651 1016
rect 2797 1004 2803 1016
rect 36 997 60 1003
rect 132 997 156 1003
rect 196 997 252 1003
rect 660 997 860 1003
rect 1060 997 1132 1003
rect 1188 997 1244 1003
rect 1716 997 1827 1003
rect 1453 984 1459 996
rect 196 977 204 983
rect 212 977 460 983
rect 532 977 732 983
rect 756 977 764 983
rect 852 977 876 983
rect 1012 977 1116 983
rect 1156 977 1212 983
rect 1316 977 1404 983
rect 1476 977 1500 983
rect 1652 977 1660 983
rect 1684 977 1692 983
rect 1796 977 1804 983
rect 1821 983 1827 997
rect 1844 997 2460 1003
rect 2484 997 2508 1003
rect 2516 997 2764 1003
rect 2900 997 2908 1003
rect 2980 997 3100 1003
rect 3117 997 3155 1003
rect 1821 977 1852 983
rect 1892 977 2236 983
rect 2260 977 2460 983
rect 2532 977 2860 983
rect 3117 983 3123 997
rect 2932 977 3123 983
rect 3149 983 3155 997
rect 3188 997 3564 1003
rect 3636 997 4204 1003
rect 4260 997 4284 1003
rect 4580 997 4588 1003
rect 4724 997 4748 1003
rect 4772 997 5116 1003
rect 3149 977 3372 983
rect 3604 977 3916 983
rect 3940 977 4140 983
rect 4164 977 4268 983
rect 4356 977 4460 983
rect 4500 977 4668 983
rect 4708 977 4716 983
rect 4756 977 4780 983
rect 4900 977 4908 983
rect 5044 977 5052 983
rect 5140 977 5180 983
rect 5204 977 5267 983
rect 1869 964 1875 976
rect 3405 964 3411 976
rect 3469 964 3475 976
rect 260 957 268 963
rect 372 957 396 963
rect 452 957 476 963
rect 644 957 1740 963
rect 1748 957 1788 963
rect 1844 957 1852 963
rect 1892 957 1900 963
rect 1956 957 1964 963
rect 1988 957 2364 963
rect 2388 957 2396 963
rect 2596 957 2684 963
rect 2708 957 2732 963
rect 285 944 291 956
rect 621 944 627 956
rect 2429 944 2435 956
rect 2525 944 2531 956
rect 2797 944 2803 963
rect 2836 957 2908 963
rect 2932 957 3276 963
rect 3348 957 3372 963
rect 3508 957 3532 963
rect 3620 957 3628 963
rect 3652 957 3660 963
rect 3684 957 3756 963
rect 3780 957 3804 963
rect 3812 957 3868 963
rect 3876 957 3980 963
rect 4036 957 4108 963
rect 4148 957 4732 963
rect 4740 957 4956 963
rect 4964 957 4972 963
rect 5156 957 5164 963
rect 308 937 316 943
rect 468 937 540 943
rect 628 937 1196 943
rect 1476 937 1484 943
rect 1492 937 1980 943
rect 2004 937 2012 943
rect 2084 937 2092 943
rect 2116 937 2124 943
rect 2132 937 2412 943
rect 2452 937 2460 943
rect 2564 937 2572 943
rect 2724 937 2732 943
rect 2772 937 2780 943
rect 2813 937 2924 943
rect 13 924 19 936
rect 2653 924 2659 936
rect 2669 924 2675 936
rect 148 917 188 923
rect 196 917 444 923
rect 516 917 524 923
rect 548 917 572 923
rect 580 917 636 923
rect 804 917 1084 923
rect 1108 917 1292 923
rect 1300 917 1340 923
rect 1540 917 1628 923
rect 1684 917 1692 923
rect 1716 917 2156 923
rect 2180 917 2252 923
rect 2308 917 2316 923
rect 2420 917 2444 923
rect 2500 917 2636 923
rect 2813 923 2819 937
rect 2964 937 2972 943
rect 3108 937 3164 943
rect 3268 937 3372 943
rect 3444 937 3548 943
rect 3604 937 3948 943
rect 3972 937 4012 943
rect 4029 937 4076 943
rect 2756 917 2819 923
rect 2829 917 2844 923
rect 2900 917 3900 923
rect 3940 917 3980 923
rect 4029 923 4035 937
rect 4084 937 4156 943
rect 4196 937 4204 943
rect 4244 937 4396 943
rect 4404 937 4412 943
rect 4468 937 4492 943
rect 4500 937 4508 943
rect 4708 937 4876 943
rect 4932 937 5116 943
rect 4004 917 4035 923
rect 4068 917 4076 923
rect 4100 917 4604 923
rect 4612 917 5052 923
rect 5140 917 5164 923
rect 2285 904 2291 916
rect 116 897 124 903
rect 228 897 236 903
rect 244 897 940 903
rect 1060 897 1068 903
rect 1076 897 1340 903
rect 1492 897 1980 903
rect 2020 897 2092 903
rect 2180 897 2188 903
rect 2228 897 2236 903
rect 2260 897 2268 903
rect 2308 897 2764 903
rect 2788 897 2844 903
rect 2868 897 2988 903
rect 3012 897 3068 903
rect 3140 897 3148 903
rect 3220 897 3315 903
rect 3309 884 3315 897
rect 3348 897 3724 903
rect 3780 897 3788 903
rect 3828 897 3836 903
rect 3860 897 3948 903
rect 4036 897 4876 903
rect 4884 897 4892 903
rect 4916 897 5004 903
rect 5028 897 5068 903
rect 5188 897 5196 903
rect 340 877 348 883
rect 452 877 684 883
rect 772 877 828 883
rect 884 877 1164 883
rect 1245 877 1388 883
rect 180 857 300 863
rect 308 857 764 863
rect 1245 863 1251 877
rect 1572 877 1708 883
rect 1748 877 1804 883
rect 2004 877 2380 883
rect 2093 864 2099 877
rect 2388 877 2396 883
rect 2420 877 2860 883
rect 2996 877 3212 883
rect 3236 877 3292 883
rect 3316 877 4588 883
rect 4612 877 4748 883
rect 4772 877 4844 883
rect 1140 857 1251 863
rect 1380 857 1388 863
rect 1412 857 1644 863
rect 1652 857 1724 863
rect 1748 857 1756 863
rect 1940 857 1948 863
rect 2148 857 2796 863
rect 2820 857 3116 863
rect 3124 857 3260 863
rect 3364 857 3724 863
rect 3748 857 3820 863
rect 3837 857 3868 863
rect 388 837 1020 843
rect 1028 837 1084 843
rect 1156 837 1164 843
rect 1348 837 1548 843
rect 1556 837 1596 843
rect 1732 837 1804 843
rect 1812 837 1948 843
rect 1956 837 2988 843
rect 3172 837 3180 843
rect 3204 837 3260 843
rect 3300 837 3500 843
rect 3837 843 3843 857
rect 3892 857 4060 863
rect 4068 857 4364 863
rect 3508 837 3843 843
rect 3860 837 4188 843
rect 4324 837 4444 843
rect 4452 837 5148 843
rect 852 817 1356 823
rect 1716 817 1724 823
rect 2052 817 2108 823
rect 2164 817 2236 823
rect 2276 817 2652 823
rect 2788 817 2812 823
rect 2868 817 3004 823
rect 3044 817 3580 823
rect 3844 817 4012 823
rect 4036 817 4044 823
rect 164 797 172 803
rect 212 797 236 803
rect 308 797 316 803
rect 324 797 348 803
rect 1156 797 1644 803
rect 1780 797 1788 803
rect 2132 797 2140 803
rect 2180 797 2188 803
rect 2244 797 2252 803
rect 2340 797 2396 803
rect 2420 797 3212 803
rect 3236 797 3244 803
rect 3380 797 3388 803
rect 3540 797 3596 803
rect 3796 797 3852 803
rect 4045 784 4051 796
rect 436 777 451 783
rect 445 764 451 777
rect 1044 777 1180 783
rect 1364 777 1372 783
rect 1444 777 1580 783
rect 1588 777 1660 783
rect 1700 777 1964 783
rect 2004 777 2028 783
rect 2036 777 2060 783
rect 2068 777 2140 783
rect 2148 777 2332 783
rect 2340 777 3068 783
rect 3076 777 3564 783
rect 3668 777 3708 783
rect 3949 764 3955 783
rect 4260 777 4428 783
rect 4820 777 4940 783
rect 5165 777 5180 783
rect 3997 764 4003 776
rect 52 757 60 763
rect 68 757 252 763
rect 260 757 364 763
rect 852 757 1116 763
rect 1156 757 1324 763
rect 1332 757 1500 763
rect 1604 757 2156 763
rect 2228 757 2236 763
rect 2260 757 2636 763
rect 2676 757 3052 763
rect 3188 757 3196 763
rect 3380 757 3388 763
rect 3460 757 3900 763
rect 3924 757 3932 763
rect 4052 757 4076 763
rect 4100 757 4652 763
rect 4852 757 4892 763
rect 5140 757 5196 763
rect 276 737 284 743
rect 388 737 396 743
rect 404 737 460 743
rect 532 737 540 743
rect 820 737 988 743
rect 1012 737 1036 743
rect 1092 737 1324 743
rect 1396 737 1404 743
rect 1604 737 1644 743
rect 1860 737 2172 743
rect 2180 737 2188 743
rect 2228 737 2268 743
rect 2404 737 2428 743
rect 2484 737 2508 743
rect 2580 737 2588 743
rect 2756 737 3596 743
rect 3636 737 3644 743
rect 3652 737 4012 743
rect 4020 737 4028 743
rect 4084 737 4172 743
rect 4292 737 4396 743
rect 4628 737 4636 743
rect 4804 737 4828 743
rect 4884 737 4956 743
rect 5156 737 5164 743
rect 141 724 147 736
rect 189 724 195 736
rect 477 724 483 736
rect 2365 724 2371 736
rect 2653 724 2659 736
rect 5037 724 5043 736
rect 244 717 284 723
rect 292 717 476 723
rect 548 717 556 723
rect 612 717 828 723
rect 836 717 1484 723
rect 1508 717 1516 723
rect 1572 717 1580 723
rect 1620 717 1628 723
rect 1636 717 2012 723
rect 2036 717 2364 723
rect 2484 717 2540 723
rect 2724 717 2748 723
rect 2772 717 2780 723
rect 2788 717 3052 723
rect 3188 717 3292 723
rect 3396 717 3756 723
rect 3764 717 3836 723
rect 3844 717 3852 723
rect 3876 717 3964 723
rect 3988 717 4044 723
rect 4180 717 4316 723
rect 4324 717 4652 723
rect 4692 717 4956 723
rect 4964 717 4988 723
rect 20 697 796 703
rect 900 697 1004 703
rect 1044 697 1052 703
rect 1108 697 1148 703
rect 1188 697 1196 703
rect 1316 697 1324 703
rect 1348 697 1356 703
rect 1364 697 2716 703
rect 2772 697 2780 703
rect 2820 697 2972 703
rect 3124 697 3180 703
rect 3220 697 3580 703
rect 3588 697 3596 703
rect 3636 697 3708 703
rect 3716 697 3724 703
rect 3764 697 4204 703
rect 4260 697 4268 703
rect 4356 697 4380 703
rect 4404 697 4412 703
rect 4500 697 4508 703
rect 4628 697 4780 703
rect 4788 697 4796 703
rect 4916 697 5036 703
rect 4605 684 4611 696
rect 228 677 316 683
rect 340 677 403 683
rect 68 657 204 663
rect 340 657 380 663
rect 397 663 403 677
rect 420 677 492 683
rect 532 677 620 683
rect 644 677 652 683
rect 676 677 1452 683
rect 1588 677 1644 683
rect 1668 677 1772 683
rect 1780 677 2252 683
rect 2276 677 2332 683
rect 2340 677 2380 683
rect 2420 677 2428 683
rect 2468 677 2476 683
rect 2500 677 2524 683
rect 2580 677 2844 683
rect 2868 677 2876 683
rect 2916 677 2924 683
rect 2948 677 2956 683
rect 2980 677 3020 683
rect 3060 677 3516 683
rect 3540 677 3548 683
rect 3572 677 3692 683
rect 3700 677 3708 683
rect 3748 677 3820 683
rect 3828 677 4556 683
rect 4644 677 4828 683
rect 5092 677 5100 683
rect 4925 664 4931 676
rect 397 657 428 663
rect 516 657 684 663
rect 692 657 1052 663
rect 1092 657 1196 663
rect 1220 657 1692 663
rect 1732 657 1740 663
rect 1764 657 2812 663
rect 2820 657 2828 663
rect 2852 657 3036 663
rect 3140 657 3452 663
rect 3460 657 4124 663
rect 4132 657 4444 663
rect 4532 657 4540 663
rect 4692 657 4716 663
rect 4788 657 4796 663
rect 5044 657 5148 663
rect 3053 644 3059 656
rect 132 637 812 643
rect 820 637 1004 643
rect 1044 637 1228 643
rect 1236 637 1324 643
rect 1348 637 1596 643
rect 1668 637 1772 643
rect 1796 637 2044 643
rect 2052 637 2060 643
rect 2084 637 2108 643
rect 2164 637 2172 643
rect 2196 637 2220 643
rect 2276 637 2284 643
rect 2292 637 2908 643
rect 3108 637 3148 643
rect 3220 637 3228 643
rect 3268 637 3820 643
rect 3844 637 3852 643
rect 3876 637 4028 643
rect 4052 637 4076 643
rect 4148 637 4300 643
rect 4452 637 4828 643
rect 4836 637 5084 643
rect 180 617 204 623
rect 356 617 364 623
rect 708 617 844 623
rect 932 617 940 623
rect 964 617 972 623
rect 1092 617 1100 623
rect 1156 617 1164 623
rect 1204 617 1244 623
rect 1316 617 1324 623
rect 1348 617 1548 623
rect 1732 617 1756 623
rect 1764 617 1772 623
rect 1997 617 2140 623
rect 1005 604 1011 616
rect 452 597 460 603
rect 500 597 524 603
rect 548 597 556 603
rect 628 597 972 603
rect 1108 597 1116 603
rect 1140 597 1180 603
rect 1236 597 1244 603
rect 1300 597 1468 603
rect 1540 597 1548 603
rect 1997 603 2003 617
rect 2196 617 2220 623
rect 2244 617 2252 623
rect 2276 617 2300 623
rect 2388 617 2396 623
rect 2484 617 2492 623
rect 2516 617 2700 623
rect 2724 617 2732 623
rect 2756 617 2828 623
rect 2868 617 2988 623
rect 3012 617 3020 623
rect 3044 617 3091 623
rect 2365 604 2371 616
rect 1620 597 2003 603
rect 2100 597 2140 603
rect 2180 597 2332 603
rect 2388 597 2412 603
rect 2429 597 2476 603
rect 228 577 748 583
rect 788 577 812 583
rect 932 577 988 583
rect 1028 577 1932 583
rect 1956 577 1980 583
rect 2004 577 2012 583
rect 2020 577 2060 583
rect 2068 577 2252 583
rect 2429 583 2435 597
rect 2516 597 2540 603
rect 2580 597 2588 603
rect 2724 597 2812 603
rect 2868 597 2876 603
rect 2948 597 3068 603
rect 3085 603 3091 617
rect 3124 617 3132 623
rect 3140 617 3164 623
rect 3172 617 3228 623
rect 3332 617 3452 623
rect 3476 617 3484 623
rect 3508 617 3516 623
rect 3684 617 3692 623
rect 3716 617 3756 623
rect 3908 617 3916 623
rect 3956 617 3996 623
rect 4020 617 4044 623
rect 4100 617 4124 623
rect 4148 617 4156 623
rect 4212 617 4972 623
rect 5076 617 5212 623
rect 3245 604 3251 616
rect 4173 604 4179 616
rect 3085 597 3148 603
rect 3188 597 3235 603
rect 2276 577 2435 583
rect 2484 577 2908 583
rect 3060 577 3132 583
rect 3188 577 3196 583
rect 3229 583 3235 597
rect 3316 597 3340 603
rect 3444 597 3692 603
rect 3972 597 4012 603
rect 4036 597 4108 603
rect 4196 597 4204 603
rect 4276 597 4316 603
rect 4612 597 4732 603
rect 4804 597 4892 603
rect 5044 597 5116 603
rect 5133 584 5139 596
rect 3229 577 3324 583
rect 3348 577 3356 583
rect 3812 577 3884 583
rect 3940 577 4044 583
rect 4068 577 4076 583
rect 4132 577 4252 583
rect 4324 577 4348 583
rect 4644 577 4652 583
rect 4724 577 4828 583
rect 4852 577 5052 583
rect 52 557 156 563
rect 276 557 412 563
rect 516 557 572 563
rect 692 557 1036 563
rect 1076 557 1100 563
rect 1252 557 1676 563
rect 1700 557 1708 563
rect 1764 557 1788 563
rect 1812 557 1884 563
rect 1988 557 2028 563
rect 2068 557 2108 563
rect 2132 557 2140 563
rect 2148 557 2268 563
rect 2292 557 2300 563
rect 2340 557 2348 563
rect 2372 557 2412 563
rect 2436 557 2508 563
rect 2532 557 2556 563
rect 2580 557 2604 563
rect 2692 557 2764 563
rect 2772 557 2908 563
rect 2948 557 2988 563
rect 3012 557 3020 563
rect 3044 557 3260 563
rect 3284 557 3292 563
rect 3332 557 3580 563
rect 3620 557 3692 563
rect 3716 557 3788 563
rect 3828 557 4076 563
rect 4084 557 4092 563
rect 4116 557 4140 563
rect 4164 557 4188 563
rect 4212 557 4332 563
rect 4532 557 4547 563
rect 4580 557 4588 563
rect 4596 557 4972 563
rect 5060 557 5068 563
rect 100 537 108 543
rect 164 537 172 543
rect 196 537 236 543
rect 244 537 252 543
rect 372 537 860 543
rect 877 537 956 543
rect 877 524 883 537
rect 1092 537 1212 543
rect 1236 537 1276 543
rect 1412 537 1436 543
rect 1540 537 1548 543
rect 1604 537 1612 543
rect 1636 537 1644 543
rect 1668 537 1692 543
rect 1716 537 1740 543
rect 1748 537 1868 543
rect 1876 537 3020 543
rect 3076 537 3084 543
rect 3172 537 3308 543
rect 3325 537 3388 543
rect 1325 524 1331 536
rect 196 517 204 523
rect 340 517 396 523
rect 500 517 508 523
rect 564 517 764 523
rect 788 517 796 523
rect 836 517 844 523
rect 916 517 956 523
rect 996 517 1036 523
rect 1108 517 1116 523
rect 1236 517 1276 523
rect 1364 517 1372 523
rect 1444 517 1452 523
rect 1508 517 2460 523
rect 2500 517 2540 523
rect 2564 517 2668 523
rect 2692 517 2780 523
rect 2804 517 2956 523
rect 2996 517 3084 523
rect 3108 517 3132 523
rect 3268 517 3276 523
rect 3325 523 3331 537
rect 3412 537 3644 543
rect 3668 537 3740 543
rect 3764 537 3788 543
rect 3860 537 4236 543
rect 4372 537 4380 543
rect 4420 537 4556 543
rect 4612 537 4620 543
rect 4692 537 4700 543
rect 4804 537 4812 543
rect 4836 537 4876 543
rect 5117 543 5123 556
rect 5108 537 5123 543
rect 3645 524 3651 536
rect 4957 524 4963 536
rect 3300 517 3331 523
rect 3348 517 3356 523
rect 3364 517 3628 523
rect 3668 517 3772 523
rect 3892 517 4460 523
rect 4468 517 4924 523
rect 5124 517 5148 523
rect 2973 504 2979 516
rect 3213 504 3219 516
rect 68 497 268 503
rect 340 497 348 503
rect 596 497 652 503
rect 660 497 1020 503
rect 1412 497 1420 503
rect 1444 497 1628 503
rect 1636 497 1772 503
rect 1780 497 1900 503
rect 1908 497 2012 503
rect 2036 497 2060 503
rect 2100 497 2108 503
rect 2164 497 2796 503
rect 2804 497 2812 503
rect 2852 497 2860 503
rect 3044 497 3116 503
rect 3124 497 3132 503
rect 3236 497 3292 503
rect 3364 497 3372 503
rect 3460 497 3868 503
rect 3892 497 3932 503
rect 3956 497 4028 503
rect 4052 497 4092 503
rect 4116 497 4124 503
rect 4164 497 4428 503
rect 4500 497 4540 503
rect 4628 497 5084 503
rect 5108 497 5164 503
rect 324 477 636 483
rect 660 477 876 483
rect 948 477 956 483
rect 1396 477 1420 483
rect 1428 477 2524 483
rect 2532 477 2700 483
rect 2932 477 3036 483
rect 3124 477 3308 483
rect 3460 477 3484 483
rect 3540 477 3548 483
rect 3700 477 3708 483
rect 3732 477 4508 483
rect 4596 477 4636 483
rect 4692 477 4716 483
rect 893 457 899 476
rect 1012 457 1228 463
rect 1236 457 1244 463
rect 1668 457 1676 463
rect 1700 457 1820 463
rect 1828 457 2236 463
rect 2244 457 2300 463
rect 2324 457 2428 463
rect 2468 457 2492 463
rect 2685 457 3084 463
rect 580 437 1372 443
rect 1380 437 1868 443
rect 1988 437 1996 443
rect 2052 437 2060 443
rect 2068 437 2188 443
rect 2212 437 2268 443
rect 2276 437 2284 443
rect 2404 437 2412 443
rect 2685 443 2691 457
rect 3140 457 3916 463
rect 4020 457 4476 463
rect 4500 457 4812 463
rect 2468 437 2691 443
rect 2708 437 3084 443
rect 3300 437 3836 443
rect 3988 437 4188 443
rect 4260 437 4620 443
rect 20 417 28 423
rect 1108 417 1116 423
rect 1156 417 2908 423
rect 2932 417 3148 423
rect 3172 417 4460 423
rect 4740 417 4748 423
rect 1076 397 1212 403
rect 1220 397 1404 403
rect 1533 397 1644 403
rect 1533 383 1539 397
rect 2068 397 2716 403
rect 2740 397 2748 403
rect 2836 397 2860 403
rect 2900 397 2908 403
rect 2948 397 2956 403
rect 3044 397 3052 403
rect 3149 397 3244 403
rect 1661 384 1667 396
rect 2045 384 2051 396
rect 916 377 1539 383
rect 1556 377 1612 383
rect 1844 377 2028 383
rect 2196 377 2332 383
rect 3149 383 3155 397
rect 3332 397 3340 403
rect 3348 397 3356 403
rect 3364 397 3372 403
rect 4068 397 4300 403
rect 4404 397 4764 403
rect 2388 377 3155 383
rect 3172 377 3180 383
rect 3316 377 3580 383
rect 3620 377 3852 383
rect 4180 377 4188 383
rect 324 357 780 363
rect 788 357 828 363
rect 916 357 1116 363
rect 1220 357 1564 363
rect 1652 357 1996 363
rect 2020 357 2652 363
rect 2660 357 2892 363
rect 2900 357 3052 363
rect 3060 357 3068 363
rect 3124 357 3196 363
rect 3252 357 3740 363
rect 3844 357 5148 363
rect 548 337 604 343
rect 628 337 636 343
rect 676 337 700 343
rect 740 337 812 343
rect 820 337 1244 343
rect 1588 337 1596 343
rect 1620 337 1628 343
rect 1652 337 1660 343
rect 1684 337 1692 343
rect 1732 337 1740 343
rect 1796 337 1820 343
rect 1860 337 1868 343
rect 1892 337 1900 343
rect 1908 337 1932 343
rect 2068 337 2076 343
rect 2260 337 2268 343
rect 2276 337 2332 343
rect 2692 337 2796 343
rect 3044 337 3644 343
rect 3780 337 3820 343
rect 3860 337 3884 343
rect 4004 337 4012 343
rect 4244 337 4252 343
rect 4292 337 4316 343
rect 4324 337 4428 343
rect 4580 337 4604 343
rect 4644 337 4668 343
rect 4980 337 5020 343
rect 5108 337 5180 343
rect 1293 324 1299 336
rect 2621 324 2627 336
rect 2813 324 2819 336
rect 20 317 44 323
rect 276 317 284 323
rect 372 317 380 323
rect 468 317 796 323
rect 820 317 844 323
rect 868 317 908 323
rect 996 317 1036 323
rect 1076 317 1084 323
rect 1124 317 1148 323
rect 1204 317 1244 323
rect 1380 317 1916 323
rect 1924 317 2188 323
rect 2580 317 2604 323
rect 2644 317 2668 323
rect 2852 317 2924 323
rect 2948 317 3004 323
rect 3028 317 3372 323
rect 3380 317 3388 323
rect 3460 317 3468 323
rect 3508 317 3692 323
rect 3796 317 3804 323
rect 3844 317 3900 323
rect 3956 317 3964 323
rect 4116 317 4131 323
rect 4212 317 4412 323
rect 4724 317 5100 323
rect 2509 304 2515 316
rect 3821 304 3827 316
rect 4557 304 4563 316
rect 100 297 124 303
rect 148 297 172 303
rect 228 297 236 303
rect 292 297 332 303
rect 372 297 716 303
rect 724 297 1260 303
rect 1268 297 1324 303
rect 1332 297 2140 303
rect 2148 297 2156 303
rect 2173 297 2188 303
rect 2420 297 2428 303
rect 2612 297 3100 303
rect 3108 297 3548 303
rect 3668 297 3804 303
rect 3892 297 3932 303
rect 3988 297 4268 303
rect 4276 297 4332 303
rect 4436 297 4508 303
rect 4708 297 4748 303
rect 4772 297 4796 303
rect 4852 297 4860 303
rect 4996 297 5004 303
rect 2525 284 2531 296
rect 4621 284 4627 296
rect 52 277 124 283
rect 244 277 588 283
rect 317 264 323 277
rect 596 277 684 283
rect 701 277 1340 283
rect 196 257 268 263
rect 340 257 636 263
rect 413 244 419 257
rect 701 263 707 277
rect 1492 277 1900 283
rect 1956 277 1964 283
rect 1988 277 1996 283
rect 2052 277 2092 283
rect 2100 277 2108 283
rect 2132 277 2307 283
rect 644 257 707 263
rect 772 257 780 263
rect 852 257 2204 263
rect 2260 257 2284 263
rect 2301 263 2307 277
rect 2324 277 2380 283
rect 2404 277 2428 283
rect 2468 277 2476 283
rect 2516 277 2524 283
rect 2596 277 2684 283
rect 2708 277 2716 283
rect 2740 277 2764 283
rect 2804 277 2844 283
rect 2868 277 2883 283
rect 2301 257 2396 263
rect 2420 257 2540 263
rect 2612 257 2796 263
rect 2820 257 2828 263
rect 2852 257 2860 263
rect 2877 263 2883 277
rect 2900 277 2988 283
rect 2996 277 3068 283
rect 3092 277 3164 283
rect 3172 277 3180 283
rect 3204 277 3212 283
rect 3252 277 3260 283
rect 3284 277 4156 283
rect 4180 277 4364 283
rect 4388 277 4412 283
rect 4532 277 4556 283
rect 4644 277 4652 283
rect 4724 277 4771 283
rect 2877 257 2892 263
rect 2916 257 2972 263
rect 2980 257 3004 263
rect 3076 257 3212 263
rect 3220 257 3340 263
rect 3364 257 3468 263
rect 3492 257 3500 263
rect 3508 257 3660 263
rect 3684 257 4300 263
rect 4356 257 4476 263
rect 4612 257 4748 263
rect 4765 263 4771 277
rect 4788 277 4796 283
rect 4836 277 4876 283
rect 5028 277 5052 283
rect 5133 283 5139 296
rect 5124 277 5139 283
rect 4765 257 4844 263
rect 4884 257 4892 263
rect 5060 257 5084 263
rect 132 237 284 243
rect 516 237 796 243
rect 804 237 876 243
rect 900 237 988 243
rect 996 237 1068 243
rect 1076 237 1372 243
rect 1460 237 1651 243
rect 84 217 92 223
rect 404 217 556 223
rect 612 217 700 223
rect 724 217 828 223
rect 980 217 1244 223
rect 1268 217 1276 223
rect 1645 223 1651 237
rect 1668 237 1708 243
rect 1716 237 1836 243
rect 1876 237 1891 243
rect 1908 237 1964 243
rect 2004 237 2028 243
rect 2036 237 2044 243
rect 2061 237 2076 243
rect 2100 237 2508 243
rect 2532 237 2572 243
rect 2580 237 2972 243
rect 2980 237 3068 243
rect 3860 237 3916 243
rect 4468 237 4796 243
rect 4804 237 4972 243
rect 1981 224 1987 236
rect 1645 217 1692 223
rect 1764 217 1772 223
rect 1860 217 1868 223
rect 2004 217 2012 223
rect 2020 217 2028 223
rect 2468 217 2668 223
rect 2788 217 2860 223
rect 2948 217 2956 223
rect 3140 217 3420 223
rect 3444 217 3676 223
rect 3748 217 3772 223
rect 4004 217 4044 223
rect 4196 217 4668 223
rect 4772 217 4780 223
rect 4804 217 4812 223
rect 580 197 652 203
rect 932 197 956 203
rect 1572 197 1948 203
rect 1997 197 2092 203
rect 1133 184 1139 196
rect 308 177 332 183
rect 356 177 364 183
rect 580 177 604 183
rect 692 177 700 183
rect 756 177 972 183
rect 1156 177 1164 183
rect 1204 177 1244 183
rect 1268 177 1356 183
rect 1524 177 1612 183
rect 1636 177 1772 183
rect 1997 183 2003 197
rect 2244 197 2284 203
rect 2500 197 2508 203
rect 2692 197 2700 203
rect 2772 197 2844 203
rect 3012 197 3052 203
rect 3300 197 3468 203
rect 3492 197 4012 203
rect 4020 197 4044 203
rect 4148 197 4156 203
rect 4180 197 4188 203
rect 4212 197 4220 203
rect 4260 197 4300 203
rect 4324 197 4332 203
rect 4676 197 4844 203
rect 4884 197 5004 203
rect 1796 177 2003 183
rect 2020 177 2028 183
rect 2045 177 2060 183
rect 2109 183 2115 196
rect 4093 184 4099 196
rect 2100 177 2115 183
rect 2132 177 2220 183
rect 2228 177 2412 183
rect 2436 177 2972 183
rect 3140 177 3148 183
rect 3188 177 3196 183
rect 3364 177 3420 183
rect 3444 177 3452 183
rect 3540 177 3580 183
rect 3604 177 3948 183
rect 3988 177 4076 183
rect 4148 177 4428 183
rect 4436 177 4444 183
rect 4676 177 5180 183
rect 125 163 131 176
rect 445 164 451 176
rect 733 164 739 176
rect 3965 164 3971 176
rect 125 157 140 163
rect 276 157 428 163
rect 461 157 476 163
rect 564 157 716 163
rect 788 157 988 163
rect 1060 157 1068 163
rect 1092 157 1196 163
rect 1252 157 1340 163
rect 1428 157 1564 163
rect 1652 157 1692 163
rect 1812 157 2204 163
rect 2212 157 2620 163
rect 2756 157 2780 163
rect 2836 157 3740 163
rect 3748 157 3756 163
rect 3780 157 3868 163
rect 4068 157 4476 163
rect 4516 157 4524 163
rect 4772 157 4796 163
rect 4820 157 4835 163
rect 4852 157 4972 163
rect 4996 157 5004 163
rect 5092 157 5132 163
rect 5156 157 5171 163
rect 1757 144 1763 156
rect 5069 144 5075 156
rect 100 137 124 143
rect 196 137 300 143
rect 308 137 764 143
rect 772 137 860 143
rect 884 137 892 143
rect 916 137 924 143
rect 948 137 1020 143
rect 1044 137 1452 143
rect 1492 137 1548 143
rect 1604 137 1740 143
rect 1892 137 2012 143
rect 2036 137 2044 143
rect 2052 137 2124 143
rect 2180 137 2204 143
rect 2388 137 3404 143
rect 3412 137 3420 143
rect 3444 137 3532 143
rect 3556 137 3564 143
rect 3588 137 3603 143
rect 3620 137 3756 143
rect 3796 137 3900 143
rect 3956 137 4108 143
rect 4164 137 4172 143
rect 4196 137 4268 143
rect 4292 137 4380 143
rect 4404 137 4428 143
rect 4548 137 4684 143
rect 4708 137 4812 143
rect 4852 137 4908 143
rect 4948 137 5020 143
rect 3773 124 3779 136
rect 196 117 220 123
rect 292 117 300 123
rect 500 117 1180 123
rect 1716 117 2092 123
rect 2100 117 2524 123
rect 2580 117 2604 123
rect 2628 117 2684 123
rect 2708 117 2732 123
rect 2804 117 2812 123
rect 2836 117 2940 123
rect 2964 117 3004 123
rect 3028 117 3116 123
rect 3156 117 3292 123
rect 3380 117 3388 123
rect 3412 117 3564 123
rect 3572 117 3628 123
rect 3908 117 4028 123
rect 4052 117 4076 123
rect 4116 117 4652 123
rect 4660 117 4732 123
rect 4788 117 4796 123
rect 4900 117 4908 123
rect 5060 117 5148 123
rect 1181 104 1187 116
rect 228 97 268 103
rect 276 97 380 103
rect 525 97 540 103
rect 612 97 620 103
rect 628 97 636 103
rect 724 97 1084 103
rect 1092 97 1171 103
rect 669 84 675 96
rect 484 77 652 83
rect 788 77 812 83
rect 1165 83 1171 97
rect 1204 97 1452 103
rect 1572 97 1676 103
rect 1812 97 1900 103
rect 1908 97 2172 103
rect 2212 97 2220 103
rect 2420 97 3324 103
rect 3332 97 3340 103
rect 3540 97 3596 103
rect 3652 97 3660 103
rect 3956 97 3996 103
rect 4084 97 4236 103
rect 4484 97 4508 103
rect 4564 97 4588 103
rect 4061 84 4067 96
rect 1165 77 1260 83
rect 1748 77 2428 83
rect 2452 77 2460 83
rect 2468 77 2540 83
rect 2548 77 2908 83
rect 2948 77 3052 83
rect 3060 77 3068 83
rect 3092 77 3100 83
rect 3156 77 3164 83
rect 3268 77 3276 83
rect 3780 77 4028 83
rect 4404 77 5212 83
rect 925 57 931 76
rect 1652 57 1932 63
rect 1940 57 1980 63
rect 1988 57 2972 63
rect 2980 57 2988 63
rect 3156 57 3500 63
rect 1828 37 2428 43
rect 2813 24 2819 36
rect 1988 17 1996 23
rect 2020 17 2028 23
<< m4contact >>
rect 2300 3616 2308 3624
rect 2892 3616 2900 3624
rect 3372 3616 3380 3624
rect 4892 3596 4900 3604
rect 3676 3576 3684 3584
rect 956 3556 964 3564
rect 1884 3556 1892 3564
rect 3100 3556 3108 3564
rect 4556 3556 4564 3564
rect 4988 3556 4996 3564
rect 492 3536 500 3544
rect 988 3536 996 3544
rect 380 3516 388 3524
rect 1404 3516 1412 3524
rect 1820 3516 1828 3524
rect 1964 3516 1972 3524
rect 2060 3516 2068 3524
rect 2156 3516 2164 3524
rect 2204 3516 2212 3524
rect 2220 3516 2228 3524
rect 2684 3516 2692 3524
rect 2748 3516 2756 3524
rect 2860 3516 2868 3524
rect 2876 3516 2884 3524
rect 3084 3516 3092 3524
rect 4444 3516 4452 3524
rect 4972 3516 4980 3524
rect 108 3496 116 3504
rect 1228 3496 1236 3504
rect 1244 3496 1252 3504
rect 1420 3496 1428 3504
rect 3068 3496 3076 3504
rect 3116 3496 3124 3504
rect 3468 3496 3476 3504
rect 3580 3496 3588 3504
rect 4844 3496 4852 3504
rect 156 3476 164 3484
rect 220 3476 228 3484
rect 652 3476 660 3484
rect 1276 3476 1284 3484
rect 1804 3476 1812 3484
rect 1836 3476 1844 3484
rect 2540 3476 2548 3484
rect 2556 3476 2564 3484
rect 2572 3476 2580 3484
rect 2652 3476 2660 3484
rect 2780 3476 2788 3484
rect 3404 3476 3412 3484
rect 3452 3476 3460 3484
rect 3820 3476 3828 3484
rect 3852 3476 3860 3484
rect 3932 3476 3940 3484
rect 3948 3476 3956 3484
rect 3964 3476 3972 3484
rect 3980 3476 3988 3484
rect 4044 3476 4052 3484
rect 4076 3476 4084 3484
rect 4332 3476 4340 3484
rect 4380 3476 4388 3484
rect 4892 3476 4900 3484
rect 5052 3476 5060 3484
rect 5132 3476 5140 3484
rect 780 3456 788 3464
rect 796 3456 804 3464
rect 860 3456 868 3464
rect 940 3456 948 3464
rect 956 3456 964 3464
rect 1180 3456 1188 3464
rect 1708 3456 1716 3464
rect 2028 3456 2036 3464
rect 2492 3456 2500 3464
rect 2508 3456 2516 3464
rect 3148 3456 3156 3464
rect 3452 3456 3460 3464
rect 3500 3456 3508 3464
rect 3516 3456 3524 3464
rect 3532 3456 3540 3464
rect 3564 3456 3572 3464
rect 3628 3456 3636 3464
rect 3660 3456 3668 3464
rect 3708 3456 3716 3464
rect 4684 3456 4692 3464
rect 4700 3456 4708 3464
rect 5164 3456 5172 3464
rect 348 3436 356 3444
rect 476 3436 484 3444
rect 556 3436 564 3444
rect 796 3436 804 3444
rect 1916 3436 1924 3444
rect 2076 3436 2084 3444
rect 2236 3436 2244 3444
rect 2332 3436 2340 3444
rect 2380 3436 2388 3444
rect 2396 3436 2404 3444
rect 2492 3436 2500 3444
rect 2524 3436 2532 3444
rect 3308 3436 3316 3444
rect 3324 3436 3332 3444
rect 3548 3436 3556 3444
rect 3596 3436 3604 3444
rect 4060 3436 4068 3444
rect 4204 3436 4212 3444
rect 4268 3436 4276 3444
rect 4428 3436 4436 3444
rect 4460 3436 4468 3444
rect 4604 3436 4612 3444
rect 4620 3436 4628 3444
rect 4652 3436 4660 3444
rect 4668 3436 4676 3444
rect 4700 3436 4708 3444
rect 4924 3436 4932 3444
rect 4940 3436 4948 3444
rect 716 3416 724 3424
rect 1036 3416 1044 3424
rect 1084 3416 1092 3424
rect 1100 3416 1108 3424
rect 1740 3416 1748 3424
rect 2268 3416 2276 3424
rect 2300 3416 2308 3424
rect 2316 3416 2324 3424
rect 2764 3416 2772 3424
rect 2796 3416 2804 3424
rect 2972 3416 2980 3424
rect 3036 3416 3044 3424
rect 3180 3416 3188 3424
rect 3372 3416 3380 3424
rect 3484 3416 3492 3424
rect 3900 3416 3908 3424
rect 4092 3416 4100 3424
rect 1116 3396 1124 3404
rect 1164 3396 1172 3404
rect 1292 3396 1300 3404
rect 1756 3396 1764 3404
rect 2236 3396 2244 3404
rect 2364 3396 2372 3404
rect 2508 3396 2516 3404
rect 2748 3396 2756 3404
rect 2908 3396 2916 3404
rect 3004 3396 3012 3404
rect 3020 3396 3028 3404
rect 3196 3396 3204 3404
rect 3228 3396 3236 3404
rect 3244 3396 3252 3404
rect 3388 3396 3396 3404
rect 588 3376 596 3384
rect 1324 3376 1332 3384
rect 1500 3376 1508 3384
rect 3132 3376 3140 3384
rect 3564 3396 3572 3404
rect 3724 3396 3732 3404
rect 3804 3396 3812 3404
rect 4092 3396 4100 3404
rect 4108 3396 4116 3404
rect 4172 3396 4180 3404
rect 5100 3396 5108 3404
rect 956 3356 964 3364
rect 1020 3356 1028 3364
rect 1052 3356 1060 3364
rect 1100 3356 1108 3364
rect 1244 3356 1252 3364
rect 1260 3356 1268 3364
rect 1308 3356 1316 3364
rect 1340 3356 1348 3364
rect 1548 3356 1556 3364
rect 156 3336 164 3344
rect 364 3336 372 3344
rect 380 3336 388 3344
rect 476 3336 484 3344
rect 732 3336 740 3344
rect 764 3336 772 3344
rect 796 3336 804 3344
rect 828 3336 836 3344
rect 860 3336 868 3344
rect 908 3336 916 3344
rect 1052 3336 1060 3344
rect 1148 3336 1156 3344
rect 1212 3336 1220 3344
rect 1692 3356 1700 3364
rect 1724 3356 1732 3364
rect 2028 3356 2036 3364
rect 2124 3356 2132 3364
rect 2380 3356 2388 3364
rect 2412 3356 2420 3364
rect 2444 3356 2452 3364
rect 2508 3356 2516 3364
rect 2620 3356 2628 3364
rect 2636 3356 2644 3364
rect 2716 3356 2724 3364
rect 2892 3356 2900 3364
rect 3052 3356 3060 3364
rect 3116 3356 3124 3364
rect 3180 3356 3188 3364
rect 3324 3356 3332 3364
rect 3340 3356 3348 3364
rect 3500 3356 3508 3364
rect 4044 3376 4052 3384
rect 4428 3376 4436 3384
rect 4460 3376 4468 3384
rect 4524 3376 4532 3384
rect 5052 3376 5060 3384
rect 5116 3376 5124 3384
rect 3964 3356 3972 3364
rect 3996 3356 4004 3364
rect 4028 3356 4036 3364
rect 4060 3356 4068 3364
rect 4092 3356 4100 3364
rect 4172 3356 4180 3364
rect 4988 3356 4996 3364
rect 1788 3336 1796 3344
rect 1804 3336 1812 3344
rect 1852 3336 1860 3344
rect 1884 3336 1892 3344
rect 2236 3336 2244 3344
rect 3372 3336 3380 3344
rect 3404 3336 3412 3344
rect 3436 3336 3444 3344
rect 1100 3316 1108 3324
rect 2764 3316 2772 3324
rect 2860 3316 2868 3324
rect 2924 3316 2932 3324
rect 3020 3316 3028 3324
rect 3084 3316 3092 3324
rect 3116 3316 3124 3324
rect 3164 3316 3172 3324
rect 3564 3316 3572 3324
rect 3676 3316 3684 3324
rect 3740 3316 3748 3324
rect 4204 3336 4212 3344
rect 4188 3316 4196 3324
rect 4860 3336 4868 3344
rect 4972 3336 4980 3344
rect 5116 3336 5124 3344
rect 4332 3316 4340 3324
rect 4364 3316 4372 3324
rect 4908 3316 4916 3324
rect 5004 3316 5012 3324
rect 92 3296 100 3304
rect 252 3296 260 3304
rect 364 3296 372 3304
rect 396 3296 404 3304
rect 444 3296 452 3304
rect 492 3296 500 3304
rect 876 3296 884 3304
rect 892 3296 900 3304
rect 1116 3296 1124 3304
rect 1148 3296 1156 3304
rect 2556 3296 2564 3304
rect 2588 3296 2596 3304
rect 2636 3296 2644 3304
rect 3804 3296 3812 3304
rect 3996 3296 4004 3304
rect 4060 3296 4068 3304
rect 4172 3296 4180 3304
rect 5100 3296 5108 3304
rect 284 3276 292 3284
rect 508 3276 516 3284
rect 956 3276 964 3284
rect 1372 3276 1380 3284
rect 1452 3276 1460 3284
rect 1660 3276 1668 3284
rect 1676 3276 1684 3284
rect 1724 3276 1732 3284
rect 2012 3276 2020 3284
rect 2108 3276 2116 3284
rect 2172 3276 2180 3284
rect 2220 3276 2228 3284
rect 2364 3276 2372 3284
rect 2524 3276 2532 3284
rect 2556 3276 2564 3284
rect 4268 3276 4276 3284
rect 4716 3276 4724 3284
rect 844 3256 852 3264
rect 1196 3256 1204 3264
rect 1564 3256 1572 3264
rect 764 3236 772 3244
rect 2204 3256 2212 3264
rect 2236 3256 2244 3264
rect 2284 3256 2292 3264
rect 2988 3256 2996 3264
rect 3260 3256 3268 3264
rect 3292 3256 3300 3264
rect 3436 3256 3444 3264
rect 3484 3256 3492 3264
rect 4940 3256 4948 3264
rect 1852 3236 1860 3244
rect 1900 3236 1908 3244
rect 1932 3236 1940 3244
rect 3036 3236 3044 3244
rect 4588 3236 4596 3244
rect 4620 3236 4628 3244
rect 4636 3236 4644 3244
rect 4844 3236 4852 3244
rect 4972 3236 4980 3244
rect 5036 3236 5044 3244
rect 5116 3236 5124 3244
rect 332 3216 340 3224
rect 972 3216 980 3224
rect 1868 3216 1876 3224
rect 1980 3216 1988 3224
rect 2508 3216 2516 3224
rect 460 3196 468 3204
rect 1932 3196 1940 3204
rect 3116 3196 3124 3204
rect 3132 3196 3140 3204
rect 3772 3196 3780 3204
rect 4732 3196 4740 3204
rect 1308 3176 1316 3184
rect 1356 3176 1364 3184
rect 2188 3176 2196 3184
rect 2268 3176 2276 3184
rect 3100 3176 3108 3184
rect 3852 3176 3860 3184
rect 524 3156 532 3164
rect 1020 3156 1028 3164
rect 2556 3156 2564 3164
rect 204 3136 212 3144
rect 1308 3136 1316 3144
rect 1356 3136 1364 3144
rect 1404 3136 1412 3144
rect 1724 3136 1732 3144
rect 2812 3136 2820 3144
rect 3036 3156 3044 3164
rect 3788 3156 3796 3164
rect 3020 3136 3028 3144
rect 3052 3136 3060 3144
rect 3516 3136 3524 3144
rect 4028 3136 4036 3144
rect 4348 3136 4356 3144
rect 4684 3136 4692 3144
rect 4748 3136 4756 3144
rect 4764 3136 4772 3144
rect 4812 3136 4820 3144
rect 188 3116 196 3124
rect 252 3116 260 3124
rect 732 3116 740 3124
rect 892 3116 900 3124
rect 1340 3116 1348 3124
rect 1388 3116 1396 3124
rect 1484 3116 1492 3124
rect 1692 3116 1700 3124
rect 1788 3116 1796 3124
rect 2124 3116 2132 3124
rect 2220 3116 2228 3124
rect 2460 3116 2468 3124
rect 3516 3116 3524 3124
rect 3548 3116 3556 3124
rect 3580 3116 3588 3124
rect 3628 3116 3636 3124
rect 3740 3116 3748 3124
rect 4444 3116 4452 3124
rect 4764 3116 4772 3124
rect 4860 3116 4868 3124
rect 4892 3116 4900 3124
rect 5004 3116 5012 3124
rect 172 3096 180 3104
rect 316 3096 324 3104
rect 700 3096 708 3104
rect 764 3096 772 3104
rect 796 3096 804 3104
rect 908 3096 916 3104
rect 1004 3096 1012 3104
rect 1196 3096 1204 3104
rect 1276 3096 1284 3104
rect 1788 3096 1796 3104
rect 1932 3096 1940 3104
rect 2028 3096 2036 3104
rect 2076 3096 2084 3104
rect 2172 3096 2180 3104
rect 2204 3096 2212 3104
rect 2252 3096 2260 3104
rect 3132 3096 3140 3104
rect 3356 3096 3364 3104
rect 3372 3096 3380 3104
rect 3404 3096 3412 3104
rect 3948 3096 3956 3104
rect 4028 3096 4036 3104
rect 4060 3096 4068 3104
rect 4524 3096 4532 3104
rect 4556 3096 4564 3104
rect 4604 3096 4612 3104
rect 4636 3096 4644 3104
rect 204 3076 212 3084
rect 236 3076 244 3084
rect 748 3076 756 3084
rect 812 3076 820 3084
rect 924 3076 932 3084
rect 1180 3076 1188 3084
rect 1260 3076 1268 3084
rect 220 3056 228 3064
rect 972 3056 980 3064
rect 1116 3056 1124 3064
rect 1132 3056 1140 3064
rect 1532 3076 1540 3084
rect 2268 3076 2276 3084
rect 1308 3056 1316 3064
rect 1644 3056 1652 3064
rect 2204 3056 2212 3064
rect 2380 3076 2388 3084
rect 2652 3076 2660 3084
rect 2684 3076 2692 3084
rect 2716 3076 2724 3084
rect 2748 3076 2756 3084
rect 2780 3076 2788 3084
rect 3020 3076 3028 3084
rect 4716 3076 4724 3084
rect 2444 3056 2452 3064
rect 2476 3056 2484 3064
rect 2668 3056 2676 3064
rect 2700 3056 2708 3064
rect 684 3036 692 3044
rect 796 3036 804 3044
rect 940 3036 948 3044
rect 1036 3036 1044 3044
rect 1084 3036 1092 3044
rect 1228 3036 1236 3044
rect 2508 3036 2516 3044
rect 2604 3036 2612 3044
rect 2652 3036 2660 3044
rect 2796 3036 2804 3044
rect 2972 3056 2980 3064
rect 3084 3056 3092 3064
rect 3212 3056 3220 3064
rect 3340 3056 3348 3064
rect 3372 3056 3380 3064
rect 3404 3056 3412 3064
rect 3468 3056 3476 3064
rect 3532 3056 3540 3064
rect 3676 3056 3684 3064
rect 3292 3036 3300 3044
rect 3452 3036 3460 3044
rect 3548 3036 3556 3044
rect 3820 3056 3828 3064
rect 4060 3056 4068 3064
rect 4668 3056 4676 3064
rect 5052 3056 5060 3064
rect 3980 3036 3988 3044
rect 4172 3036 4180 3044
rect 4572 3036 4580 3044
rect 4604 3036 4612 3044
rect 4668 3036 4676 3044
rect 540 3016 548 3024
rect 1852 3016 1860 3024
rect 1964 3016 1972 3024
rect 2908 3016 2916 3024
rect 2924 3016 2932 3024
rect 3100 3016 3108 3024
rect 3196 3016 3204 3024
rect 3436 3016 3444 3024
rect 4172 3016 4180 3024
rect 4652 3016 4660 3024
rect 4716 3016 4724 3024
rect 4892 3016 4900 3024
rect 940 2996 948 3004
rect 2108 2996 2116 3004
rect 2140 2996 2148 3004
rect 2156 2996 2164 3004
rect 2876 2996 2884 3004
rect 2908 2996 2916 3004
rect 2956 2996 2964 3004
rect 460 2976 468 2984
rect 684 2976 692 2984
rect 780 2976 788 2984
rect 1132 2976 1140 2984
rect 1244 2976 1252 2984
rect 1308 2976 1316 2984
rect 1340 2976 1348 2984
rect 1404 2976 1412 2984
rect 1452 2976 1460 2984
rect 2364 2976 2372 2984
rect 3452 2976 3460 2984
rect 3484 2976 3492 2984
rect 3532 2996 3540 3004
rect 3580 2996 3588 3004
rect 3612 2996 3620 3004
rect 4572 2996 4580 3004
rect 4892 2996 4900 3004
rect 3900 2976 3908 2984
rect 5068 2976 5076 2984
rect 412 2956 420 2964
rect 460 2956 468 2964
rect 940 2956 948 2964
rect 972 2956 980 2964
rect 1356 2956 1364 2964
rect 2476 2956 2484 2964
rect 2524 2956 2532 2964
rect 2556 2956 2564 2964
rect 2668 2956 2676 2964
rect 2700 2956 2708 2964
rect 2764 2956 2772 2964
rect 2780 2956 2788 2964
rect 2828 2956 2836 2964
rect 2860 2956 2868 2964
rect 3564 2956 3572 2964
rect 3948 2956 3956 2964
rect 4732 2956 4740 2964
rect 4908 2956 4916 2964
rect 5084 2956 5092 2964
rect 508 2936 516 2944
rect 540 2936 548 2944
rect 716 2936 724 2944
rect 796 2936 804 2944
rect 1628 2936 1636 2944
rect 1660 2936 1668 2944
rect 1948 2936 1956 2944
rect 2044 2936 2052 2944
rect 2092 2936 2100 2944
rect 2140 2936 2148 2944
rect 2508 2936 2516 2944
rect 2588 2936 2596 2944
rect 3036 2936 3044 2944
rect 3180 2936 3188 2944
rect 3324 2936 3332 2944
rect 3356 2936 3364 2944
rect 4028 2936 4036 2944
rect 4044 2936 4052 2944
rect 4204 2936 4212 2944
rect 4220 2936 4228 2944
rect 4700 2936 4708 2944
rect 4732 2936 4740 2944
rect 4764 2936 4772 2944
rect 5100 2936 5108 2944
rect 140 2916 148 2924
rect 316 2916 324 2924
rect 380 2916 388 2924
rect 524 2916 532 2924
rect 540 2916 548 2924
rect 780 2916 788 2924
rect 844 2916 852 2924
rect 1836 2916 1844 2924
rect 1900 2916 1908 2924
rect 2140 2916 2148 2924
rect 2188 2916 2196 2924
rect 2268 2916 2276 2924
rect 2764 2916 2772 2924
rect 3132 2916 3140 2924
rect 3276 2916 3284 2924
rect 3308 2916 3316 2924
rect 3484 2916 3492 2924
rect 3548 2916 3556 2924
rect 3628 2916 3636 2924
rect 3692 2916 3700 2924
rect 3708 2916 3716 2924
rect 3836 2916 3844 2924
rect 3852 2916 3860 2924
rect 3980 2916 3988 2924
rect 3996 2916 4004 2924
rect 4268 2916 4276 2924
rect 4348 2916 4356 2924
rect 4364 2916 4372 2924
rect 4508 2916 4516 2924
rect 4748 2916 4756 2924
rect 108 2896 116 2904
rect 284 2896 292 2904
rect 412 2896 420 2904
rect 588 2896 596 2904
rect 652 2896 660 2904
rect 780 2896 788 2904
rect 1084 2896 1092 2904
rect 1132 2896 1140 2904
rect 1244 2896 1252 2904
rect 1404 2896 1412 2904
rect 1436 2896 1444 2904
rect 1452 2896 1460 2904
rect 1484 2896 1492 2904
rect 1580 2896 1588 2904
rect 1596 2896 1604 2904
rect 1644 2896 1652 2904
rect 1692 2896 1700 2904
rect 1708 2896 1716 2904
rect 1772 2896 1780 2904
rect 1820 2896 1828 2904
rect 1884 2896 1892 2904
rect 2316 2896 2324 2904
rect 2332 2896 2340 2904
rect 2428 2896 2436 2904
rect 2940 2896 2948 2904
rect 3020 2896 3028 2904
rect 3116 2896 3124 2904
rect 3148 2896 3156 2904
rect 3180 2896 3188 2904
rect 3308 2896 3316 2904
rect 3324 2896 3332 2904
rect 3388 2896 3396 2904
rect 3404 2896 3412 2904
rect 3564 2896 3572 2904
rect 3740 2896 3748 2904
rect 3996 2896 4004 2904
rect 4044 2896 4052 2904
rect 4140 2896 4148 2904
rect 4300 2896 4308 2904
rect 4460 2896 4468 2904
rect 5004 2896 5012 2904
rect 5148 2896 5156 2904
rect 332 2876 340 2884
rect 908 2876 916 2884
rect 972 2876 980 2884
rect 1340 2876 1348 2884
rect 1436 2876 1444 2884
rect 1532 2876 1540 2884
rect 1804 2876 1812 2884
rect 1980 2876 1988 2884
rect 2028 2876 2036 2884
rect 2220 2876 2228 2884
rect 2380 2876 2388 2884
rect 2428 2876 2436 2884
rect 2604 2876 2612 2884
rect 2924 2876 2932 2884
rect 2988 2876 2996 2884
rect 4012 2876 4020 2884
rect 4124 2876 4132 2884
rect 5116 2876 5124 2884
rect 412 2856 420 2864
rect 716 2856 724 2864
rect 1004 2856 1012 2864
rect 1628 2856 1636 2864
rect 1708 2856 1716 2864
rect 1900 2856 1908 2864
rect 1932 2856 1940 2864
rect 2108 2856 2116 2864
rect 2556 2856 2564 2864
rect 2588 2856 2596 2864
rect 2604 2856 2612 2864
rect 3036 2856 3044 2864
rect 3420 2856 3428 2864
rect 4892 2856 4900 2864
rect 4956 2856 4964 2864
rect 5148 2856 5156 2864
rect 460 2836 468 2844
rect 1580 2836 1588 2844
rect 2172 2836 2180 2844
rect 2236 2836 2244 2844
rect 2828 2836 2836 2844
rect 3868 2836 3876 2844
rect 4172 2836 4180 2844
rect 4316 2836 4324 2844
rect 5004 2836 5012 2844
rect 1612 2816 1620 2824
rect 1772 2816 1780 2824
rect 1804 2816 1812 2824
rect 1980 2816 1988 2824
rect 2284 2816 2292 2824
rect 2764 2816 2772 2824
rect 2796 2816 2804 2824
rect 2828 2816 2836 2824
rect 2972 2816 2980 2824
rect 3404 2816 3412 2824
rect 4300 2816 4308 2824
rect 4668 2816 4676 2824
rect 5212 2816 5220 2824
rect 476 2796 484 2804
rect 2508 2796 2516 2804
rect 2556 2796 2564 2804
rect 3036 2796 3044 2804
rect 3356 2796 3364 2804
rect 3532 2796 3540 2804
rect 3884 2796 3892 2804
rect 4412 2796 4420 2804
rect 4428 2796 4436 2804
rect 5180 2796 5188 2804
rect 812 2776 820 2784
rect 1020 2776 1028 2784
rect 1244 2776 1252 2784
rect 2092 2776 2100 2784
rect 2156 2776 2164 2784
rect 2700 2776 2708 2784
rect 2748 2776 2756 2784
rect 3308 2776 3316 2784
rect 3484 2776 3492 2784
rect 492 2756 500 2764
rect 2732 2756 2740 2764
rect 2892 2756 2900 2764
rect 3180 2756 3188 2764
rect 4156 2756 4164 2764
rect 4396 2756 4404 2764
rect 4492 2756 4500 2764
rect 4828 2756 4836 2764
rect 5164 2756 5172 2764
rect 188 2736 196 2744
rect 300 2736 308 2744
rect 508 2736 516 2744
rect 636 2736 644 2744
rect 924 2736 932 2744
rect 1196 2736 1204 2744
rect 1900 2736 1908 2744
rect 2012 2736 2020 2744
rect 2140 2736 2148 2744
rect 2188 2736 2196 2744
rect 2428 2736 2436 2744
rect 2556 2736 2564 2744
rect 2780 2736 2788 2744
rect 2796 2736 2804 2744
rect 2956 2736 2964 2744
rect 3020 2736 3028 2744
rect 3420 2736 3428 2744
rect 4140 2736 4148 2744
rect 4892 2736 4900 2744
rect 12 2716 20 2724
rect 44 2716 52 2724
rect 108 2716 116 2724
rect 284 2716 292 2724
rect 636 2716 644 2724
rect 700 2716 708 2724
rect 924 2716 932 2724
rect 1004 2716 1012 2724
rect 1084 2716 1092 2724
rect 1100 2716 1108 2724
rect 1292 2716 1300 2724
rect 1564 2716 1572 2724
rect 2252 2716 2260 2724
rect 2620 2716 2628 2724
rect 2636 2716 2644 2724
rect 3196 2716 3204 2724
rect 3228 2716 3236 2724
rect 3276 2716 3284 2724
rect 3436 2716 3444 2724
rect 3564 2716 3572 2724
rect 3644 2716 3652 2724
rect 3932 2716 3940 2724
rect 4044 2716 4052 2724
rect 4156 2716 4164 2724
rect 4620 2716 4628 2724
rect 4828 2716 4836 2724
rect 5084 2716 5092 2724
rect 1148 2696 1156 2704
rect 1196 2696 1204 2704
rect 1420 2696 1428 2704
rect 1516 2696 1524 2704
rect 1596 2696 1604 2704
rect 3004 2696 3012 2704
rect 3100 2696 3108 2704
rect 3676 2696 3684 2704
rect 3756 2696 3764 2704
rect 3852 2696 3860 2704
rect 3868 2696 3876 2704
rect 3932 2696 3940 2704
rect 4636 2696 4644 2704
rect 4684 2696 4692 2704
rect 4844 2696 4852 2704
rect 4876 2696 4884 2704
rect 492 2676 500 2684
rect 508 2676 516 2684
rect 540 2676 548 2684
rect 572 2676 580 2684
rect 588 2676 596 2684
rect 796 2676 804 2684
rect 828 2676 836 2684
rect 972 2676 980 2684
rect 1020 2676 1028 2684
rect 1132 2676 1140 2684
rect 1244 2676 1252 2684
rect 1452 2676 1460 2684
rect 1500 2676 1508 2684
rect 1516 2676 1524 2684
rect 2380 2676 2388 2684
rect 2748 2676 2756 2684
rect 2844 2676 2852 2684
rect 2940 2676 2948 2684
rect 2956 2676 2964 2684
rect 4220 2676 4228 2684
rect 4284 2676 4292 2684
rect 4300 2676 4308 2684
rect 4332 2676 4340 2684
rect 4364 2676 4372 2684
rect 4444 2676 4452 2684
rect 4460 2676 4468 2684
rect 4508 2676 4516 2684
rect 4940 2676 4948 2684
rect 5084 2676 5092 2684
rect 172 2656 180 2664
rect 204 2656 212 2664
rect 268 2656 276 2664
rect 284 2656 292 2664
rect 316 2656 324 2664
rect 412 2656 420 2664
rect 396 2636 404 2644
rect 460 2656 468 2664
rect 812 2656 820 2664
rect 860 2656 868 2664
rect 1244 2656 1252 2664
rect 2652 2656 2660 2664
rect 2700 2656 2708 2664
rect 2892 2656 2900 2664
rect 2972 2656 2980 2664
rect 3068 2656 3076 2664
rect 428 2636 436 2644
rect 748 2636 756 2644
rect 1708 2636 1716 2644
rect 1772 2636 1780 2644
rect 2044 2636 2052 2644
rect 2268 2636 2276 2644
rect 2300 2636 2308 2644
rect 2524 2636 2532 2644
rect 2844 2636 2852 2644
rect 2908 2636 2916 2644
rect 3260 2656 3268 2664
rect 3324 2656 3332 2664
rect 3452 2656 3460 2664
rect 3564 2656 3572 2664
rect 3660 2656 3668 2664
rect 3836 2656 3844 2664
rect 4972 2656 4980 2664
rect 4988 2656 4996 2664
rect 5052 2656 5060 2664
rect 3100 2636 3108 2644
rect 3852 2636 3860 2644
rect 4092 2636 4100 2644
rect 4892 2636 4900 2644
rect 4956 2636 4964 2644
rect 5116 2636 5124 2644
rect 60 2596 68 2604
rect 284 2596 292 2604
rect 748 2596 756 2604
rect 956 2596 964 2604
rect 1036 2616 1044 2624
rect 1052 2616 1060 2624
rect 1308 2616 1316 2624
rect 1340 2616 1348 2624
rect 1468 2616 1476 2624
rect 1564 2616 1572 2624
rect 1580 2616 1588 2624
rect 1628 2616 1636 2624
rect 1932 2616 1940 2624
rect 1964 2616 1972 2624
rect 1996 2616 2004 2624
rect 2092 2616 2100 2624
rect 2172 2616 2180 2624
rect 2188 2616 2196 2624
rect 2300 2616 2308 2624
rect 2412 2616 2420 2624
rect 2428 2616 2436 2624
rect 3356 2616 3364 2624
rect 3484 2616 3492 2624
rect 3580 2616 3588 2624
rect 3660 2616 3668 2624
rect 3916 2616 3924 2624
rect 3996 2616 4004 2624
rect 4028 2616 4036 2624
rect 4076 2616 4084 2624
rect 4140 2616 4148 2624
rect 4284 2616 4292 2624
rect 4428 2616 4436 2624
rect 4444 2616 4452 2624
rect 4460 2616 4468 2624
rect 1788 2596 1796 2604
rect 2188 2596 2196 2604
rect 2236 2596 2244 2604
rect 364 2576 372 2584
rect 540 2576 548 2584
rect 556 2576 564 2584
rect 764 2576 772 2584
rect 828 2576 836 2584
rect 1132 2576 1140 2584
rect 1676 2576 1684 2584
rect 1980 2576 1988 2584
rect 2076 2576 2084 2584
rect 2508 2576 2516 2584
rect 2540 2596 2548 2604
rect 2556 2596 2564 2604
rect 3148 2596 3156 2604
rect 3180 2596 3188 2604
rect 3196 2596 3204 2604
rect 4012 2596 4020 2604
rect 4028 2596 4036 2604
rect 4140 2596 4148 2604
rect 3532 2576 3540 2584
rect 3644 2576 3652 2584
rect 3708 2576 3716 2584
rect 3868 2576 3876 2584
rect 4444 2596 4452 2604
rect 4572 2596 4580 2604
rect 4892 2596 4900 2604
rect 5100 2596 5108 2604
rect 4380 2576 4388 2584
rect 4492 2576 4500 2584
rect 4972 2576 4980 2584
rect 5164 2576 5172 2584
rect 108 2556 116 2564
rect 1372 2556 1380 2564
rect 1724 2556 1732 2564
rect 1788 2556 1796 2564
rect 1836 2556 1844 2564
rect 1996 2556 2004 2564
rect 2028 2556 2036 2564
rect 2044 2556 2052 2564
rect 2156 2556 2164 2564
rect 2332 2556 2340 2564
rect 2524 2556 2532 2564
rect 2796 2556 2804 2564
rect 2924 2556 2932 2564
rect 3132 2556 3140 2564
rect 3212 2556 3220 2564
rect 3308 2556 3316 2564
rect 3452 2556 3460 2564
rect 3916 2556 3924 2564
rect 4140 2556 4148 2564
rect 4604 2556 4612 2564
rect 796 2536 804 2544
rect 828 2536 836 2544
rect 940 2536 948 2544
rect 1068 2536 1076 2544
rect 1292 2536 1300 2544
rect 1308 2536 1316 2544
rect 1340 2536 1348 2544
rect 1404 2536 1412 2544
rect 2316 2536 2324 2544
rect 2524 2536 2532 2544
rect 2588 2536 2596 2544
rect 2668 2536 2676 2544
rect 2684 2536 2692 2544
rect 2924 2536 2932 2544
rect 4108 2536 4116 2544
rect 4252 2536 4260 2544
rect 4924 2536 4932 2544
rect 108 2516 116 2524
rect 156 2516 164 2524
rect 332 2516 340 2524
rect 348 2516 356 2524
rect 556 2516 564 2524
rect 716 2516 724 2524
rect 1052 2516 1060 2524
rect 1292 2516 1300 2524
rect 1740 2516 1748 2524
rect 1884 2516 1892 2524
rect 2908 2516 2916 2524
rect 3212 2516 3220 2524
rect 3372 2516 3380 2524
rect 188 2496 196 2504
rect 220 2496 228 2504
rect 444 2496 452 2504
rect 492 2496 500 2504
rect 652 2496 660 2504
rect 924 2496 932 2504
rect 972 2496 980 2504
rect 1036 2496 1044 2504
rect 1148 2496 1156 2504
rect 1628 2496 1636 2504
rect 1708 2496 1716 2504
rect 1724 2496 1732 2504
rect 1836 2496 1844 2504
rect 1900 2496 1908 2504
rect 1980 2496 1988 2504
rect 2188 2496 2196 2504
rect 2236 2496 2244 2504
rect 2268 2496 2276 2504
rect 2364 2496 2372 2504
rect 2412 2496 2420 2504
rect 2556 2496 2564 2504
rect 2684 2496 2692 2504
rect 2700 2496 2708 2504
rect 2748 2496 2756 2504
rect 2876 2496 2884 2504
rect 2988 2496 2996 2504
rect 3036 2496 3044 2504
rect 3116 2496 3124 2504
rect 3180 2496 3188 2504
rect 3196 2496 3204 2504
rect 3228 2496 3236 2504
rect 3260 2496 3268 2504
rect 3548 2516 3556 2524
rect 3612 2516 3620 2524
rect 3628 2516 3636 2524
rect 3820 2516 3828 2524
rect 3852 2516 3860 2524
rect 3932 2516 3940 2524
rect 4076 2516 4084 2524
rect 4108 2516 4116 2524
rect 4140 2516 4148 2524
rect 4156 2516 4164 2524
rect 4284 2516 4292 2524
rect 4476 2516 4484 2524
rect 4508 2516 4516 2524
rect 4524 2516 4532 2524
rect 4540 2516 4548 2524
rect 4604 2516 4612 2524
rect 3404 2496 3412 2504
rect 3532 2496 3540 2504
rect 3740 2496 3748 2504
rect 3756 2496 3764 2504
rect 3900 2496 3908 2504
rect 3996 2496 4004 2504
rect 4156 2496 4164 2504
rect 44 2476 52 2484
rect 764 2476 772 2484
rect 828 2476 836 2484
rect 876 2476 884 2484
rect 940 2476 948 2484
rect 1484 2476 1492 2484
rect 1516 2476 1524 2484
rect 1564 2476 1572 2484
rect 1628 2476 1636 2484
rect 1836 2476 1844 2484
rect 2204 2476 2212 2484
rect 2668 2476 2676 2484
rect 2860 2476 2868 2484
rect 2876 2476 2884 2484
rect 3020 2476 3028 2484
rect 3068 2476 3076 2484
rect 3100 2476 3108 2484
rect 3116 2476 3124 2484
rect 3148 2476 3156 2484
rect 3660 2476 3668 2484
rect 3772 2476 3780 2484
rect 3884 2476 3892 2484
rect 4140 2476 4148 2484
rect 4460 2476 4468 2484
rect 4556 2476 4564 2484
rect 4780 2516 4788 2524
rect 4956 2516 4964 2524
rect 4988 2516 4996 2524
rect 4780 2496 4788 2504
rect 4876 2496 4884 2504
rect 4924 2496 4932 2504
rect 4972 2496 4980 2504
rect 4956 2476 4964 2484
rect 5052 2476 5060 2484
rect 1244 2456 1252 2464
rect 1564 2456 1572 2464
rect 1580 2456 1588 2464
rect 1932 2456 1940 2464
rect 2428 2456 2436 2464
rect 4092 2456 4100 2464
rect 1948 2436 1956 2444
rect 2028 2436 2036 2444
rect 2428 2436 2436 2444
rect 2780 2436 2788 2444
rect 3020 2436 3028 2444
rect 3132 2436 3140 2444
rect 3340 2436 3348 2444
rect 3356 2436 3364 2444
rect 3372 2436 3380 2444
rect 3740 2436 3748 2444
rect 972 2416 980 2424
rect 92 2396 100 2404
rect 540 2396 548 2404
rect 588 2396 596 2404
rect 620 2396 628 2404
rect 1132 2396 1140 2404
rect 1340 2416 1348 2424
rect 2604 2416 2612 2424
rect 2668 2416 2676 2424
rect 1436 2396 1444 2404
rect 1804 2396 1812 2404
rect 2044 2396 2052 2404
rect 2428 2396 2436 2404
rect 2700 2396 2708 2404
rect 2796 2416 2804 2424
rect 2844 2416 2852 2424
rect 4012 2416 4020 2424
rect 4332 2416 4340 2424
rect 4364 2416 4372 2424
rect 460 2376 468 2384
rect 540 2376 548 2384
rect 2604 2376 2612 2384
rect 2764 2376 2772 2384
rect 3612 2396 3620 2404
rect 3228 2376 3236 2384
rect 3580 2376 3588 2384
rect 4012 2376 4020 2384
rect 4076 2376 4084 2384
rect 4236 2376 4244 2384
rect 4732 2376 4740 2384
rect 300 2356 308 2364
rect 860 2356 868 2364
rect 1916 2356 1924 2364
rect 2220 2356 2228 2364
rect 2700 2356 2708 2364
rect 3052 2356 3060 2364
rect 3612 2356 3620 2364
rect 3932 2356 3940 2364
rect 508 2336 516 2344
rect 604 2336 612 2344
rect 1340 2336 1348 2344
rect 1404 2336 1412 2344
rect 1532 2336 1540 2344
rect 1580 2336 1588 2344
rect 1756 2336 1764 2344
rect 1788 2336 1796 2344
rect 2684 2336 2692 2344
rect 3340 2336 3348 2344
rect 3388 2336 3396 2344
rect 3468 2336 3476 2344
rect 3580 2336 3588 2344
rect 3916 2336 3924 2344
rect 828 2316 836 2324
rect 988 2316 996 2324
rect 1100 2316 1108 2324
rect 1132 2316 1140 2324
rect 12 2296 20 2304
rect 476 2296 484 2304
rect 492 2296 500 2304
rect 860 2296 868 2304
rect 1308 2296 1316 2304
rect 1580 2316 1588 2324
rect 1740 2316 1748 2324
rect 1852 2316 1860 2324
rect 1900 2316 1908 2324
rect 2476 2316 2484 2324
rect 3020 2316 3028 2324
rect 3356 2316 3364 2324
rect 3660 2316 3668 2324
rect 3772 2316 3780 2324
rect 4108 2316 4116 2324
rect 4124 2316 4132 2324
rect 4140 2316 4148 2324
rect 4636 2316 4644 2324
rect 4892 2316 4900 2324
rect 1436 2296 1444 2304
rect 1516 2296 1524 2304
rect 1532 2296 1540 2304
rect 1756 2296 1764 2304
rect 1868 2296 1876 2304
rect 2076 2296 2084 2304
rect 2124 2296 2132 2304
rect 2252 2296 2260 2304
rect 2460 2296 2468 2304
rect 2476 2296 2484 2304
rect 2524 2296 2532 2304
rect 2556 2296 2564 2304
rect 2796 2296 2804 2304
rect 2860 2296 2868 2304
rect 364 2276 372 2284
rect 844 2276 852 2284
rect 924 2276 932 2284
rect 972 2276 980 2284
rect 1036 2276 1044 2284
rect 1052 2276 1060 2284
rect 1564 2276 1572 2284
rect 1580 2276 1588 2284
rect 1820 2276 1828 2284
rect 2012 2276 2020 2284
rect 2108 2276 2116 2284
rect 2236 2276 2244 2284
rect 2396 2276 2404 2284
rect 2412 2276 2420 2284
rect 3036 2296 3044 2304
rect 3212 2296 3220 2304
rect 3292 2296 3300 2304
rect 3404 2296 3412 2304
rect 4252 2296 4260 2304
rect 4284 2296 4292 2304
rect 5004 2296 5012 2304
rect 5052 2296 5060 2304
rect 5148 2296 5156 2304
rect 2588 2276 2596 2284
rect 2748 2276 2756 2284
rect 2844 2276 2852 2284
rect 2876 2276 2884 2284
rect 2908 2276 2916 2284
rect 2988 2276 2996 2284
rect 3020 2276 3028 2284
rect 3084 2276 3092 2284
rect 3548 2276 3556 2284
rect 3596 2276 3604 2284
rect 3708 2276 3716 2284
rect 3740 2276 3748 2284
rect 3772 2276 3780 2284
rect 4236 2276 4244 2284
rect 4412 2276 4420 2284
rect 4428 2276 4436 2284
rect 4540 2276 4548 2284
rect 4652 2276 4660 2284
rect 4764 2276 4772 2284
rect 4972 2276 4980 2284
rect 5036 2276 5044 2284
rect 5148 2276 5156 2284
rect 172 2256 180 2264
rect 204 2256 212 2264
rect 220 2256 228 2264
rect 332 2256 340 2264
rect 460 2256 468 2264
rect 524 2256 532 2264
rect 540 2256 548 2264
rect 636 2256 644 2264
rect 668 2256 676 2264
rect 844 2256 852 2264
rect 1580 2256 1588 2264
rect 1628 2256 1636 2264
rect 1724 2256 1732 2264
rect 1852 2256 1860 2264
rect 1868 2256 1876 2264
rect 3180 2256 3188 2264
rect 3260 2256 3268 2264
rect 3324 2256 3332 2264
rect 3388 2256 3396 2264
rect 3580 2256 3588 2264
rect 3788 2256 3796 2264
rect 3868 2256 3876 2264
rect 3964 2256 3972 2264
rect 4092 2256 4100 2264
rect 4188 2256 4196 2264
rect 4316 2256 4324 2264
rect 4332 2256 4340 2264
rect 4860 2256 4868 2264
rect 332 2236 340 2244
rect 476 2236 484 2244
rect 540 2236 548 2244
rect 1788 2236 1796 2244
rect 1948 2236 1956 2244
rect 2028 2236 2036 2244
rect 2044 2236 2052 2244
rect 2300 2236 2308 2244
rect 2444 2236 2452 2244
rect 2476 2236 2484 2244
rect 2588 2236 2596 2244
rect 3308 2236 3316 2244
rect 3404 2236 3412 2244
rect 3468 2236 3476 2244
rect 3660 2236 3668 2244
rect 3996 2236 4004 2244
rect 4140 2236 4148 2244
rect 4268 2236 4276 2244
rect 1132 2216 1140 2224
rect 1708 2216 1716 2224
rect 1820 2216 1828 2224
rect 1852 2216 1860 2224
rect 1932 2216 1940 2224
rect 2172 2216 2180 2224
rect 2268 2216 2276 2224
rect 2284 2216 2292 2224
rect 2396 2216 2404 2224
rect 2412 2216 2420 2224
rect 284 2196 292 2204
rect 668 2196 676 2204
rect 1388 2196 1396 2204
rect 1516 2196 1524 2204
rect 1612 2196 1620 2204
rect 1916 2196 1924 2204
rect 1980 2196 1988 2204
rect 2188 2196 2196 2204
rect 2236 2196 2244 2204
rect 2556 2196 2564 2204
rect 2668 2216 2676 2224
rect 2748 2216 2756 2224
rect 2844 2216 2852 2224
rect 2988 2216 2996 2224
rect 3020 2216 3028 2224
rect 3324 2216 3332 2224
rect 3644 2216 3652 2224
rect 3772 2216 3780 2224
rect 3868 2216 3876 2224
rect 3916 2216 3924 2224
rect 3932 2216 3940 2224
rect 4092 2216 4100 2224
rect 4188 2216 4196 2224
rect 2908 2196 2916 2204
rect 2940 2196 2948 2204
rect 3628 2196 3636 2204
rect 3788 2196 3796 2204
rect 3980 2196 3988 2204
rect 4124 2196 4132 2204
rect 4396 2216 4404 2224
rect 4476 2216 4484 2224
rect 4508 2216 4516 2224
rect 4492 2196 4500 2204
rect 4636 2196 4644 2204
rect 4876 2196 4884 2204
rect 5036 2196 5044 2204
rect 172 2176 180 2184
rect 668 2176 676 2184
rect 700 2176 708 2184
rect 716 2176 724 2184
rect 1164 2176 1172 2184
rect 1740 2176 1748 2184
rect 1756 2176 1764 2184
rect 2556 2176 2564 2184
rect 2700 2176 2708 2184
rect 2748 2176 2756 2184
rect 3196 2176 3204 2184
rect 4604 2176 4612 2184
rect 4716 2176 4724 2184
rect 4876 2176 4884 2184
rect 60 2156 68 2164
rect 252 2156 260 2164
rect 604 2156 612 2164
rect 620 2156 628 2164
rect 748 2156 756 2164
rect 844 2156 852 2164
rect 1148 2156 1156 2164
rect 1260 2156 1268 2164
rect 1340 2156 1348 2164
rect 1372 2156 1380 2164
rect 1516 2156 1524 2164
rect 1612 2156 1620 2164
rect 1628 2156 1636 2164
rect 1724 2156 1732 2164
rect 1804 2156 1812 2164
rect 2572 2156 2580 2164
rect 2668 2156 2676 2164
rect 3340 2156 3348 2164
rect 3356 2156 3364 2164
rect 3692 2156 3700 2164
rect 3708 2156 3716 2164
rect 3980 2156 3988 2164
rect 4028 2156 4036 2164
rect 4124 2156 4132 2164
rect 4140 2156 4148 2164
rect 4236 2156 4244 2164
rect 4252 2156 4260 2164
rect 4300 2156 4308 2164
rect 4332 2156 4340 2164
rect 4348 2156 4356 2164
rect 5020 2156 5028 2164
rect 5052 2156 5060 2164
rect 284 2136 292 2144
rect 956 2136 964 2144
rect 1996 2136 2004 2144
rect 2044 2136 2052 2144
rect 2140 2136 2148 2144
rect 2188 2136 2196 2144
rect 316 2116 324 2124
rect 332 2116 340 2124
rect 364 2116 372 2124
rect 412 2116 420 2124
rect 428 2116 436 2124
rect 492 2116 500 2124
rect 796 2116 804 2124
rect 892 2116 900 2124
rect 988 2116 996 2124
rect 1036 2116 1044 2124
rect 300 2096 308 2104
rect 428 2096 436 2104
rect 572 2096 580 2104
rect 764 2096 772 2104
rect 1100 2096 1108 2104
rect 1180 2116 1188 2124
rect 1868 2116 1876 2124
rect 2076 2116 2084 2124
rect 2476 2136 2484 2144
rect 2844 2136 2852 2144
rect 2860 2136 2868 2144
rect 2876 2136 2884 2144
rect 3148 2136 3156 2144
rect 3180 2136 3188 2144
rect 3228 2136 3236 2144
rect 3260 2136 3268 2144
rect 4860 2136 4868 2144
rect 5116 2136 5124 2144
rect 2268 2116 2276 2124
rect 2572 2116 2580 2124
rect 2652 2116 2660 2124
rect 2796 2116 2804 2124
rect 2812 2116 2820 2124
rect 2844 2116 2852 2124
rect 2892 2116 2900 2124
rect 2940 2116 2948 2124
rect 2972 2116 2980 2124
rect 3100 2116 3108 2124
rect 3132 2116 3140 2124
rect 3148 2116 3156 2124
rect 3276 2116 3284 2124
rect 3452 2116 3460 2124
rect 3660 2116 3668 2124
rect 3692 2116 3700 2124
rect 3724 2116 3732 2124
rect 4252 2116 4260 2124
rect 4412 2116 4420 2124
rect 4444 2116 4452 2124
rect 4476 2116 4484 2124
rect 4492 2116 4500 2124
rect 4556 2116 4564 2124
rect 4604 2116 4612 2124
rect 4652 2116 4660 2124
rect 4780 2116 4788 2124
rect 4828 2116 4836 2124
rect 4940 2116 4948 2124
rect 5052 2116 5060 2124
rect 5116 2116 5124 2124
rect 1372 2096 1380 2104
rect 1484 2096 1492 2104
rect 2028 2096 2036 2104
rect 2236 2096 2244 2104
rect 2380 2096 2388 2104
rect 2412 2096 2420 2104
rect 2812 2096 2820 2104
rect 3292 2096 3300 2104
rect 3468 2096 3476 2104
rect 3644 2096 3652 2104
rect 3692 2096 3700 2104
rect 3708 2096 3716 2104
rect 3948 2096 3956 2104
rect 4092 2096 4100 2104
rect 4188 2096 4196 2104
rect 4444 2096 4452 2104
rect 4668 2096 4676 2104
rect 5004 2096 5012 2104
rect 156 2076 164 2084
rect 1596 2076 1604 2084
rect 1820 2076 1828 2084
rect 1852 2076 1860 2084
rect 2060 2076 2068 2084
rect 2092 2076 2100 2084
rect 2620 2076 2628 2084
rect 2684 2076 2692 2084
rect 2940 2076 2948 2084
rect 3740 2076 3748 2084
rect 4060 2076 4068 2084
rect 4396 2076 4404 2084
rect 4476 2076 4484 2084
rect 4556 2076 4564 2084
rect 396 2056 404 2064
rect 604 2056 612 2064
rect 1484 2056 1492 2064
rect 1564 2056 1572 2064
rect 1628 2056 1636 2064
rect 1724 2056 1732 2064
rect 1788 2056 1796 2064
rect 1884 2056 1892 2064
rect 1932 2056 1940 2064
rect 1964 2056 1972 2064
rect 2028 2056 2036 2064
rect 2092 2056 2100 2064
rect 2108 2056 2116 2064
rect 2444 2056 2452 2064
rect 2844 2056 2852 2064
rect 3820 2056 3828 2064
rect 3868 2056 3876 2064
rect 3980 2056 3988 2064
rect 5100 2056 5108 2064
rect 1132 2036 1140 2044
rect 1276 2036 1284 2044
rect 1532 2036 1540 2044
rect 1692 2036 1700 2044
rect 2124 2036 2132 2044
rect 2140 2036 2148 2044
rect 2476 2036 2484 2044
rect 3004 2036 3012 2044
rect 3452 2036 3460 2044
rect 3628 2036 3636 2044
rect 3772 2036 3780 2044
rect 3868 2036 3876 2044
rect 828 2016 836 2024
rect 1164 2016 1172 2024
rect 1244 2016 1252 2024
rect 1276 2016 1284 2024
rect 2060 2016 2068 2024
rect 2108 2016 2116 2024
rect 2300 2016 2308 2024
rect 2444 2016 2452 2024
rect 2668 2016 2676 2024
rect 2684 2016 2692 2024
rect 2892 2016 2900 2024
rect 2908 2016 2916 2024
rect 2940 2016 2948 2024
rect 3068 2016 3076 2024
rect 3148 2016 3156 2024
rect 3292 2016 3300 2024
rect 3308 2016 3316 2024
rect 3468 2016 3476 2024
rect 3516 2016 3524 2024
rect 3532 2016 3540 2024
rect 4364 2016 4372 2024
rect 4556 2016 4564 2024
rect 4764 2016 4772 2024
rect 188 1996 196 2004
rect 732 1996 740 2004
rect 828 1996 836 2004
rect 1116 1996 1124 2004
rect 1900 1996 1908 2004
rect 4044 1996 4052 2004
rect 4140 1996 4148 2004
rect 844 1976 852 1984
rect 860 1976 868 1984
rect 908 1976 916 1984
rect 1756 1976 1764 1984
rect 1916 1976 1924 1984
rect 2876 1976 2884 1984
rect 3404 1976 3412 1984
rect 3580 1976 3588 1984
rect 3916 1976 3924 1984
rect 4044 1976 4052 1984
rect 4300 1976 4308 1984
rect 4876 1976 4884 1984
rect 5036 1976 5044 1984
rect 476 1956 484 1964
rect 908 1956 916 1964
rect 1564 1956 1572 1964
rect 2412 1956 2420 1964
rect 2444 1956 2452 1964
rect 2572 1956 2580 1964
rect 2684 1956 2692 1964
rect 2748 1956 2756 1964
rect 2892 1956 2900 1964
rect 3196 1956 3204 1964
rect 3724 1956 3732 1964
rect 3756 1956 3764 1964
rect 3916 1956 3924 1964
rect 4076 1956 4084 1964
rect 4252 1956 4260 1964
rect 4428 1956 4436 1964
rect 4860 1956 4868 1964
rect 5164 1956 5172 1964
rect 780 1936 788 1944
rect 1724 1936 1732 1944
rect 2204 1936 2212 1944
rect 2268 1936 2276 1944
rect 3244 1936 3252 1944
rect 3404 1936 3412 1944
rect 3468 1936 3476 1944
rect 3836 1936 3844 1944
rect 4300 1936 4308 1944
rect 4348 1936 4356 1944
rect 572 1916 580 1924
rect 668 1916 676 1924
rect 764 1916 772 1924
rect 1164 1916 1172 1924
rect 1500 1916 1508 1924
rect 1692 1916 1700 1924
rect 1868 1916 1876 1924
rect 1900 1916 1908 1924
rect 1948 1916 1956 1924
rect 92 1896 100 1904
rect 380 1876 388 1884
rect 172 1856 180 1864
rect 268 1856 276 1864
rect 300 1856 308 1864
rect 476 1876 484 1884
rect 652 1896 660 1904
rect 908 1896 916 1904
rect 924 1896 932 1904
rect 1052 1896 1060 1904
rect 1340 1896 1348 1904
rect 1404 1896 1412 1904
rect 1436 1896 1444 1904
rect 1500 1896 1508 1904
rect 1516 1896 1524 1904
rect 1548 1896 1556 1904
rect 1612 1896 1620 1904
rect 1628 1896 1636 1904
rect 1788 1896 1796 1904
rect 1820 1896 1828 1904
rect 1852 1896 1860 1904
rect 2636 1916 2644 1924
rect 2732 1916 2740 1924
rect 2972 1916 2980 1924
rect 3036 1916 3044 1924
rect 3180 1916 3188 1924
rect 3772 1916 3780 1924
rect 3964 1916 3972 1924
rect 3996 1916 4004 1924
rect 4076 1916 4084 1924
rect 4588 1916 4596 1924
rect 4620 1916 4628 1924
rect 2108 1896 2116 1904
rect 2188 1896 2196 1904
rect 2572 1896 2580 1904
rect 2700 1896 2708 1904
rect 2748 1896 2756 1904
rect 2796 1896 2804 1904
rect 2876 1896 2884 1904
rect 2924 1896 2932 1904
rect 2940 1896 2948 1904
rect 3020 1896 3028 1904
rect 3052 1896 3060 1904
rect 3164 1896 3172 1904
rect 3212 1896 3220 1904
rect 3228 1896 3236 1904
rect 3292 1896 3300 1904
rect 3484 1896 3492 1904
rect 3564 1896 3572 1904
rect 3628 1896 3636 1904
rect 3660 1896 3668 1904
rect 4284 1896 4292 1904
rect 4316 1896 4324 1904
rect 4412 1896 4420 1904
rect 4860 1896 4868 1904
rect 4892 1896 4900 1904
rect 5116 1896 5124 1904
rect 796 1876 804 1884
rect 1100 1876 1108 1884
rect 1788 1876 1796 1884
rect 3500 1876 3508 1884
rect 3596 1876 3604 1884
rect 4876 1876 4884 1884
rect 5116 1876 5124 1884
rect 460 1856 468 1864
rect 844 1856 852 1864
rect 1052 1856 1060 1864
rect 1228 1856 1236 1864
rect 1340 1856 1348 1864
rect 2332 1856 2340 1864
rect 3260 1856 3268 1864
rect 3724 1856 3732 1864
rect 3836 1856 3844 1864
rect 3884 1856 3892 1864
rect 3948 1856 3956 1864
rect 4092 1856 4100 1864
rect 4268 1856 4276 1864
rect 4316 1856 4324 1864
rect 4364 1856 4372 1864
rect 4572 1856 4580 1864
rect 4636 1856 4644 1864
rect 4684 1856 4692 1864
rect 5052 1856 5060 1864
rect 348 1836 356 1844
rect 1036 1836 1044 1844
rect 1372 1836 1380 1844
rect 1516 1836 1524 1844
rect 1532 1836 1540 1844
rect 1548 1836 1556 1844
rect 1612 1836 1620 1844
rect 1628 1836 1636 1844
rect 1820 1836 1828 1844
rect 2060 1836 2068 1844
rect 956 1816 964 1824
rect 1116 1816 1124 1824
rect 1276 1816 1284 1824
rect 1372 1816 1380 1824
rect 1484 1816 1492 1824
rect 1500 1816 1508 1824
rect 1532 1816 1540 1824
rect 1596 1816 1604 1824
rect 1756 1816 1764 1824
rect 1900 1816 1908 1824
rect 1932 1816 1940 1824
rect 1980 1816 1988 1824
rect 1996 1816 2004 1824
rect 2140 1836 2148 1844
rect 2348 1836 2356 1844
rect 3084 1836 3092 1844
rect 3260 1836 3268 1844
rect 3308 1836 3316 1844
rect 3340 1836 3348 1844
rect 3388 1836 3396 1844
rect 3692 1836 3700 1844
rect 3868 1836 3876 1844
rect 4348 1836 4356 1844
rect 4412 1836 4420 1844
rect 4796 1836 4804 1844
rect 4860 1836 4868 1844
rect 4876 1836 4884 1844
rect 2140 1816 2148 1824
rect 2172 1816 2180 1824
rect 2188 1816 2196 1824
rect 2460 1816 2468 1824
rect 2508 1816 2516 1824
rect 2700 1816 2708 1824
rect 2732 1816 2740 1824
rect 2876 1816 2884 1824
rect 444 1796 452 1804
rect 748 1796 756 1804
rect 1036 1796 1044 1804
rect 1116 1796 1124 1804
rect 1164 1796 1172 1804
rect 1516 1796 1524 1804
rect 2108 1796 2116 1804
rect 2604 1796 2612 1804
rect 2620 1796 2628 1804
rect 2748 1796 2756 1804
rect 2796 1796 2804 1804
rect 2892 1796 2900 1804
rect 2908 1796 2916 1804
rect 2972 1816 2980 1824
rect 3004 1816 3012 1824
rect 3020 1816 3028 1824
rect 3068 1816 3076 1824
rect 3100 1816 3108 1824
rect 3324 1816 3332 1824
rect 2972 1796 2980 1804
rect 3116 1796 3124 1804
rect 3196 1796 3204 1804
rect 3244 1796 3252 1804
rect 3324 1796 3332 1804
rect 3340 1796 3348 1804
rect 3868 1796 3876 1804
rect 3964 1796 3972 1804
rect 3996 1796 4004 1804
rect 220 1776 228 1784
rect 476 1776 484 1784
rect 508 1776 516 1784
rect 924 1776 932 1784
rect 1644 1776 1652 1784
rect 156 1756 164 1764
rect 1324 1756 1332 1764
rect 1388 1756 1396 1764
rect 1516 1756 1524 1764
rect 1548 1756 1556 1764
rect 1676 1756 1684 1764
rect 1756 1756 1764 1764
rect 1820 1756 1828 1764
rect 1884 1756 1892 1764
rect 1932 1776 1940 1784
rect 2380 1776 2388 1784
rect 2396 1776 2404 1784
rect 2956 1776 2964 1784
rect 2988 1776 2996 1784
rect 3084 1776 3092 1784
rect 3724 1776 3732 1784
rect 3740 1776 3748 1784
rect 3980 1776 3988 1784
rect 3996 1776 4004 1784
rect 4188 1796 4196 1804
rect 4348 1796 4356 1804
rect 5084 1796 5092 1804
rect 4460 1776 4468 1784
rect 4764 1776 4772 1784
rect 2028 1756 2036 1764
rect 2268 1756 2276 1764
rect 2316 1756 2324 1764
rect 3468 1756 3476 1764
rect 3484 1756 3492 1764
rect 3516 1756 3524 1764
rect 3580 1756 3588 1764
rect 3612 1756 3620 1764
rect 3692 1756 3700 1764
rect 3724 1756 3732 1764
rect 3740 1756 3748 1764
rect 332 1736 340 1744
rect 540 1736 548 1744
rect 796 1736 804 1744
rect 1340 1736 1348 1744
rect 1708 1736 1716 1744
rect 1756 1736 1764 1744
rect 1788 1736 1796 1744
rect 2092 1736 2100 1744
rect 2108 1736 2116 1744
rect 2204 1736 2212 1744
rect 2236 1736 2244 1744
rect 3052 1736 3060 1744
rect 3068 1736 3076 1744
rect 3596 1736 3604 1744
rect 3628 1736 3636 1744
rect 3948 1756 3956 1764
rect 4060 1756 4068 1764
rect 4140 1756 4148 1764
rect 4332 1756 4340 1764
rect 4876 1756 4884 1764
rect 252 1716 260 1724
rect 492 1716 500 1724
rect 844 1716 852 1724
rect 1084 1716 1092 1724
rect 1980 1716 1988 1724
rect 1996 1716 2004 1724
rect 2012 1716 2020 1724
rect 2588 1716 2596 1724
rect 2652 1716 2660 1724
rect 2716 1716 2724 1724
rect 2748 1716 2756 1724
rect 476 1696 484 1704
rect 828 1696 836 1704
rect 844 1696 852 1704
rect 940 1696 948 1704
rect 1116 1696 1124 1704
rect 1164 1696 1172 1704
rect 1228 1696 1236 1704
rect 1276 1696 1284 1704
rect 1436 1696 1444 1704
rect 1788 1696 1796 1704
rect 1820 1696 1828 1704
rect 2252 1696 2260 1704
rect 2268 1696 2276 1704
rect 2380 1696 2388 1704
rect 2412 1696 2420 1704
rect 2444 1696 2452 1704
rect 2588 1696 2596 1704
rect 2732 1696 2740 1704
rect 2876 1716 2884 1724
rect 2892 1716 2900 1724
rect 3004 1716 3012 1724
rect 3132 1716 3140 1724
rect 2796 1696 2804 1704
rect 2908 1696 2916 1704
rect 2956 1696 2964 1704
rect 2988 1696 2996 1704
rect 3020 1696 3028 1704
rect 3068 1696 3076 1704
rect 3228 1696 3236 1704
rect 3244 1696 3252 1704
rect 3356 1716 3364 1724
rect 3708 1716 3716 1724
rect 3836 1736 3844 1744
rect 3916 1736 3924 1744
rect 3980 1736 3988 1744
rect 4092 1736 4100 1744
rect 4124 1736 4132 1744
rect 4220 1736 4228 1744
rect 4604 1736 4612 1744
rect 4652 1736 4660 1744
rect 4668 1736 4676 1744
rect 4908 1736 4916 1744
rect 4972 1736 4980 1744
rect 5004 1736 5012 1744
rect 5084 1736 5092 1744
rect 3820 1716 3828 1724
rect 4124 1716 4132 1724
rect 4220 1716 4228 1724
rect 4316 1716 4324 1724
rect 4348 1716 4356 1724
rect 4700 1716 4708 1724
rect 5084 1716 5092 1724
rect 3292 1696 3300 1704
rect 3388 1696 3396 1704
rect 3452 1696 3460 1704
rect 3468 1696 3476 1704
rect 3644 1696 3652 1704
rect 3660 1696 3668 1704
rect 4092 1696 4100 1704
rect 4348 1696 4356 1704
rect 4380 1696 4388 1704
rect 4492 1696 4500 1704
rect 4540 1696 4548 1704
rect 4796 1696 4804 1704
rect 108 1676 116 1684
rect 348 1676 356 1684
rect 524 1676 532 1684
rect 572 1676 580 1684
rect 652 1676 660 1684
rect 1276 1676 1284 1684
rect 1308 1676 1316 1684
rect 2140 1676 2148 1684
rect 2172 1676 2180 1684
rect 2700 1676 2708 1684
rect 3084 1676 3092 1684
rect 4204 1676 4212 1684
rect 4220 1676 4228 1684
rect 4380 1676 4388 1684
rect 4796 1676 4804 1684
rect 4844 1676 4852 1684
rect 5036 1676 5044 1684
rect 476 1656 484 1664
rect 892 1656 900 1664
rect 1292 1656 1300 1664
rect 1516 1656 1524 1664
rect 2300 1656 2308 1664
rect 3020 1656 3028 1664
rect 4092 1656 4100 1664
rect 4716 1656 4724 1664
rect 4828 1656 4836 1664
rect 5004 1656 5012 1664
rect 892 1636 900 1644
rect 1612 1636 1620 1644
rect 1644 1636 1652 1644
rect 1676 1636 1684 1644
rect 3004 1636 3012 1644
rect 3084 1636 3092 1644
rect 3244 1636 3252 1644
rect 3260 1636 3268 1644
rect 3708 1636 3716 1644
rect 4188 1636 4196 1644
rect 4220 1636 4228 1644
rect 4364 1636 4372 1644
rect 4524 1636 4532 1644
rect 268 1616 276 1624
rect 2236 1616 2244 1624
rect 2284 1616 2292 1624
rect 2364 1616 2372 1624
rect 2380 1616 2388 1624
rect 2956 1616 2964 1624
rect 3260 1616 3268 1624
rect 3388 1616 3396 1624
rect 3516 1616 3524 1624
rect 3644 1616 3652 1624
rect 3804 1616 3812 1624
rect 684 1596 692 1604
rect 1276 1596 1284 1604
rect 1804 1596 1812 1604
rect 1884 1596 1892 1604
rect 1916 1596 1924 1604
rect 220 1576 228 1584
rect 1788 1576 1796 1584
rect 1804 1576 1812 1584
rect 2188 1576 2196 1584
rect 2412 1576 2420 1584
rect 2684 1576 2692 1584
rect 2748 1596 2756 1604
rect 2764 1596 2772 1604
rect 3452 1596 3460 1604
rect 3484 1596 3492 1604
rect 4060 1596 4068 1604
rect 4140 1596 4148 1604
rect 4188 1596 4196 1604
rect 4764 1596 4772 1604
rect 4812 1596 4820 1604
rect 2748 1576 2756 1584
rect 2860 1576 2868 1584
rect 2940 1576 2948 1584
rect 3004 1576 3012 1584
rect 3148 1576 3156 1584
rect 3164 1576 3172 1584
rect 3580 1576 3588 1584
rect 4380 1576 4388 1584
rect 4828 1576 4836 1584
rect 4844 1576 4852 1584
rect 220 1556 228 1564
rect 1468 1556 1476 1564
rect 2092 1556 2100 1564
rect 2140 1556 2148 1564
rect 2236 1556 2244 1564
rect 2444 1556 2452 1564
rect 3644 1556 3652 1564
rect 4684 1556 4692 1564
rect 4700 1556 4708 1564
rect 5020 1556 5028 1564
rect 92 1536 100 1544
rect 652 1536 660 1544
rect 924 1536 932 1544
rect 1180 1536 1188 1544
rect 1260 1536 1268 1544
rect 1788 1536 1796 1544
rect 1852 1536 1860 1544
rect 1884 1536 1892 1544
rect 1916 1536 1924 1544
rect 2188 1536 2196 1544
rect 2204 1536 2212 1544
rect 2652 1536 2660 1544
rect 2940 1536 2948 1544
rect 2956 1536 2964 1544
rect 3132 1536 3140 1544
rect 3212 1536 3220 1544
rect 3244 1536 3252 1544
rect 3292 1536 3300 1544
rect 3340 1536 3348 1544
rect 3516 1536 3524 1544
rect 3628 1536 3636 1544
rect 4412 1536 4420 1544
rect 4476 1536 4484 1544
rect 4876 1536 4884 1544
rect 5084 1536 5092 1544
rect 76 1516 84 1524
rect 124 1516 132 1524
rect 220 1516 228 1524
rect 236 1516 244 1524
rect 460 1516 468 1524
rect 604 1516 612 1524
rect 748 1516 756 1524
rect 828 1516 836 1524
rect 988 1516 996 1524
rect 1132 1516 1140 1524
rect 1148 1516 1156 1524
rect 1468 1516 1476 1524
rect 1516 1516 1524 1524
rect 1708 1516 1716 1524
rect 2172 1516 2180 1524
rect 2300 1516 2308 1524
rect 2412 1516 2420 1524
rect 2588 1516 2596 1524
rect 3244 1516 3252 1524
rect 3292 1516 3300 1524
rect 3340 1516 3348 1524
rect 3484 1516 3492 1524
rect 3564 1516 3572 1524
rect 3996 1516 4004 1524
rect 4108 1516 4116 1524
rect 4124 1516 4132 1524
rect 4940 1516 4948 1524
rect 5036 1516 5044 1524
rect 5100 1516 5108 1524
rect 860 1496 868 1504
rect 924 1496 932 1504
rect 940 1496 948 1504
rect 1612 1496 1620 1504
rect 1756 1496 1764 1504
rect 1788 1496 1796 1504
rect 1948 1496 1956 1504
rect 2044 1496 2052 1504
rect 2172 1496 2180 1504
rect 2188 1496 2196 1504
rect 2444 1496 2452 1504
rect 2508 1496 2516 1504
rect 2572 1496 2580 1504
rect 2668 1496 2676 1504
rect 2748 1496 2756 1504
rect 2908 1496 2916 1504
rect 3052 1496 3060 1504
rect 3580 1496 3588 1504
rect 3996 1496 4004 1504
rect 4140 1496 4148 1504
rect 4188 1496 4196 1504
rect 4396 1496 4404 1504
rect 4652 1496 4660 1504
rect 4684 1496 4692 1504
rect 5068 1496 5076 1504
rect 364 1476 372 1484
rect 620 1476 628 1484
rect 748 1476 756 1484
rect 876 1476 884 1484
rect 1628 1476 1636 1484
rect 1644 1476 1652 1484
rect 1756 1476 1764 1484
rect 1788 1476 1796 1484
rect 1820 1476 1828 1484
rect 1932 1476 1940 1484
rect 1996 1476 2004 1484
rect 2028 1476 2036 1484
rect 2284 1476 2292 1484
rect 2412 1476 2420 1484
rect 3532 1476 3540 1484
rect 3660 1476 3668 1484
rect 3804 1476 3812 1484
rect 3868 1476 3876 1484
rect 3948 1476 3956 1484
rect 4108 1476 4116 1484
rect 316 1456 324 1464
rect 860 1456 868 1464
rect 892 1456 900 1464
rect 972 1456 980 1464
rect 1068 1456 1076 1464
rect 1260 1456 1268 1464
rect 1372 1456 1380 1464
rect 1420 1456 1428 1464
rect 1596 1456 1604 1464
rect 2188 1456 2196 1464
rect 2236 1456 2244 1464
rect 2300 1456 2308 1464
rect 2364 1456 2372 1464
rect 3996 1456 4004 1464
rect 4044 1456 4052 1464
rect 4124 1456 4132 1464
rect 4220 1476 4228 1484
rect 4268 1476 4276 1484
rect 4828 1476 4836 1484
rect 4924 1476 4932 1484
rect 4204 1456 4212 1464
rect 4252 1456 4260 1464
rect 4268 1456 4276 1464
rect 4300 1456 4308 1464
rect 4716 1456 4724 1464
rect 4988 1456 4996 1464
rect 5004 1456 5012 1464
rect 5084 1476 5092 1484
rect 5148 1476 5156 1484
rect 300 1436 308 1444
rect 556 1436 564 1444
rect 1132 1436 1140 1444
rect 1164 1436 1172 1444
rect 2364 1436 2372 1444
rect 2396 1436 2404 1444
rect 2572 1436 2580 1444
rect 3260 1436 3268 1444
rect 3292 1436 3300 1444
rect 3388 1436 3396 1444
rect 3452 1436 3460 1444
rect 3516 1436 3524 1444
rect 4316 1436 4324 1444
rect 4876 1436 4884 1444
rect 4972 1436 4980 1444
rect 236 1416 244 1424
rect 572 1416 580 1424
rect 1228 1416 1236 1424
rect 2108 1416 2116 1424
rect 2140 1416 2148 1424
rect 348 1396 356 1404
rect 1244 1396 1252 1404
rect 1340 1396 1348 1404
rect 1404 1396 1412 1404
rect 1516 1396 1524 1404
rect 1628 1396 1636 1404
rect 1676 1396 1684 1404
rect 1692 1396 1700 1404
rect 1836 1396 1844 1404
rect 1852 1396 1860 1404
rect 2028 1396 2036 1404
rect 2140 1396 2148 1404
rect 2172 1396 2180 1404
rect 2284 1396 2292 1404
rect 2412 1396 2420 1404
rect 2556 1416 2564 1424
rect 2572 1416 2580 1424
rect 2652 1416 2660 1424
rect 2668 1416 2676 1424
rect 2732 1416 2740 1424
rect 2796 1416 2804 1424
rect 2828 1416 2836 1424
rect 2876 1416 2884 1424
rect 2892 1416 2900 1424
rect 2908 1416 2916 1424
rect 3148 1416 3156 1424
rect 3180 1416 3188 1424
rect 3212 1416 3220 1424
rect 3340 1416 3348 1424
rect 4060 1416 4068 1424
rect 4108 1416 4116 1424
rect 4252 1416 4260 1424
rect 4268 1416 4276 1424
rect 4524 1416 4532 1424
rect 4668 1416 4676 1424
rect 4876 1416 4884 1424
rect 3068 1396 3076 1404
rect 380 1376 388 1384
rect 668 1376 676 1384
rect 1116 1376 1124 1384
rect 1324 1376 1332 1384
rect 1564 1376 1572 1384
rect 1580 1376 1588 1384
rect 1612 1376 1620 1384
rect 1644 1376 1652 1384
rect 1692 1376 1700 1384
rect 2332 1376 2340 1384
rect 2604 1376 2612 1384
rect 2988 1376 2996 1384
rect 3084 1376 3092 1384
rect 3196 1376 3204 1384
rect 3276 1376 3284 1384
rect 3340 1376 3348 1384
rect 4828 1396 4836 1404
rect 76 1356 84 1364
rect 156 1356 164 1364
rect 572 1356 580 1364
rect 588 1356 596 1364
rect 668 1356 676 1364
rect 428 1336 436 1344
rect 492 1336 500 1344
rect 524 1336 532 1344
rect 700 1336 708 1344
rect 1084 1356 1092 1364
rect 1756 1356 1764 1364
rect 1884 1356 1892 1364
rect 1900 1356 1908 1364
rect 2060 1356 2068 1364
rect 2092 1356 2100 1364
rect 2156 1356 2164 1364
rect 2236 1356 2244 1364
rect 2332 1356 2340 1364
rect 2412 1356 2420 1364
rect 2668 1356 2676 1364
rect 2748 1356 2756 1364
rect 2908 1356 2916 1364
rect 2940 1356 2948 1364
rect 3356 1356 3364 1364
rect 3372 1356 3380 1364
rect 3596 1356 3604 1364
rect 3612 1356 3620 1364
rect 3820 1376 3828 1384
rect 3708 1356 3716 1364
rect 3852 1356 3860 1364
rect 3884 1356 3892 1364
rect 3964 1376 3972 1384
rect 4460 1376 4468 1384
rect 4764 1376 4772 1384
rect 4284 1356 4292 1364
rect 4300 1356 4308 1364
rect 4380 1356 4388 1364
rect 4412 1356 4420 1364
rect 4444 1356 4452 1364
rect 4508 1356 4516 1364
rect 4572 1356 4580 1364
rect 4844 1356 4852 1364
rect 1036 1336 1044 1344
rect 92 1316 100 1324
rect 444 1316 452 1324
rect 588 1316 596 1324
rect 684 1316 692 1324
rect 860 1316 868 1324
rect 1148 1316 1156 1324
rect 1308 1336 1316 1344
rect 1324 1336 1332 1344
rect 2316 1336 2324 1344
rect 2396 1336 2404 1344
rect 2428 1336 2436 1344
rect 2492 1336 2500 1344
rect 2604 1336 2612 1344
rect 2732 1336 2740 1344
rect 2796 1336 2804 1344
rect 2812 1336 2820 1344
rect 2988 1336 2996 1344
rect 3004 1336 3012 1344
rect 3068 1336 3076 1344
rect 3100 1336 3108 1344
rect 1212 1316 1220 1324
rect 1484 1316 1492 1324
rect 1500 1316 1508 1324
rect 1740 1316 1748 1324
rect 1852 1316 1860 1324
rect 1868 1316 1876 1324
rect 1900 1316 1908 1324
rect 3660 1316 3668 1324
rect 3788 1316 3796 1324
rect 3836 1316 3844 1324
rect 3900 1316 3908 1324
rect 4044 1336 4052 1344
rect 4140 1336 4148 1344
rect 4652 1336 4660 1344
rect 4988 1336 4996 1344
rect 5100 1336 5108 1344
rect 5148 1336 5156 1344
rect 5196 1336 5204 1344
rect 3980 1316 3988 1324
rect 4012 1316 4020 1324
rect 4124 1316 4132 1324
rect 4332 1316 4340 1324
rect 4396 1316 4404 1324
rect 4444 1316 4452 1324
rect 4476 1316 4484 1324
rect 4636 1316 4644 1324
rect 4716 1316 4724 1324
rect 4748 1316 4756 1324
rect 5100 1316 5108 1324
rect 60 1296 68 1304
rect 268 1296 276 1304
rect 1084 1296 1092 1304
rect 1340 1296 1348 1304
rect 1388 1296 1396 1304
rect 1420 1296 1428 1304
rect 1884 1296 1892 1304
rect 1932 1296 1940 1304
rect 2348 1296 2356 1304
rect 2428 1296 2436 1304
rect 2508 1296 2516 1304
rect 2604 1296 2612 1304
rect 348 1276 356 1284
rect 764 1276 772 1284
rect 1996 1276 2004 1284
rect 2636 1276 2644 1284
rect 2668 1276 2676 1284
rect 2844 1276 2852 1284
rect 2924 1296 2932 1304
rect 3004 1296 3012 1304
rect 3212 1296 3220 1304
rect 3372 1296 3380 1304
rect 3388 1296 3396 1304
rect 3804 1296 3812 1304
rect 3836 1296 3844 1304
rect 4044 1296 4052 1304
rect 4332 1296 4340 1304
rect 4588 1296 4596 1304
rect 5068 1296 5076 1304
rect 5148 1296 5156 1304
rect 364 1256 372 1264
rect 524 1256 532 1264
rect 1068 1256 1076 1264
rect 1132 1256 1140 1264
rect 2028 1256 2036 1264
rect 2060 1256 2068 1264
rect 2316 1256 2324 1264
rect 2876 1256 2884 1264
rect 4140 1276 4148 1284
rect 4428 1276 4436 1284
rect 4828 1276 4836 1284
rect 4876 1276 4884 1284
rect 1324 1236 1332 1244
rect 1372 1236 1380 1244
rect 2396 1236 2404 1244
rect 2492 1236 2500 1244
rect 2748 1236 2756 1244
rect 3100 1236 3108 1244
rect 3628 1236 3636 1244
rect 3916 1236 3924 1244
rect 4108 1236 4116 1244
rect 4988 1236 4996 1244
rect 860 1216 868 1224
rect 1132 1216 1140 1224
rect 1948 1216 1956 1224
rect 1964 1216 1972 1224
rect 2140 1216 2148 1224
rect 2172 1216 2180 1224
rect 2300 1216 2308 1224
rect 2396 1216 2404 1224
rect 2428 1216 2436 1224
rect 2652 1216 2660 1224
rect 2748 1216 2756 1224
rect 2796 1216 2804 1224
rect 3004 1216 3012 1224
rect 3308 1216 3316 1224
rect 3340 1216 3348 1224
rect 3372 1216 3380 1224
rect 3708 1216 3716 1224
rect 3788 1216 3796 1224
rect 4140 1216 4148 1224
rect 4252 1216 4260 1224
rect 4524 1216 4532 1224
rect 812 1196 820 1204
rect 860 1196 868 1204
rect 2540 1196 2548 1204
rect 2604 1196 2612 1204
rect 3324 1196 3332 1204
rect 3452 1196 3460 1204
rect 3788 1196 3796 1204
rect 3836 1196 3844 1204
rect 3916 1196 3924 1204
rect 812 1176 820 1184
rect 1740 1176 1748 1184
rect 1820 1176 1828 1184
rect 1836 1176 1844 1184
rect 1260 1156 1268 1164
rect 1420 1156 1428 1164
rect 1484 1156 1492 1164
rect 1644 1156 1652 1164
rect 2140 1156 2148 1164
rect 2236 1156 2244 1164
rect 2428 1156 2436 1164
rect 2540 1176 2548 1184
rect 2652 1176 2660 1184
rect 3036 1176 3044 1184
rect 4140 1176 4148 1184
rect 5100 1176 5108 1184
rect 3436 1156 3444 1164
rect 3532 1156 3540 1164
rect 3564 1156 3572 1164
rect 3708 1156 3716 1164
rect 3980 1156 3988 1164
rect 3996 1156 4004 1164
rect 4284 1156 4292 1164
rect 4444 1156 4452 1164
rect 5100 1156 5108 1164
rect 636 1136 644 1144
rect 1164 1136 1172 1144
rect 1404 1136 1412 1144
rect 220 1116 228 1124
rect 460 1116 468 1124
rect 492 1116 500 1124
rect 588 1116 596 1124
rect 780 1116 788 1124
rect 1132 1116 1140 1124
rect 1164 1116 1172 1124
rect 1356 1116 1364 1124
rect 1468 1116 1476 1124
rect 1580 1116 1588 1124
rect 1644 1116 1652 1124
rect 1884 1116 1892 1124
rect 1916 1136 1924 1144
rect 1964 1136 1972 1144
rect 2540 1136 2548 1144
rect 3100 1136 3108 1144
rect 3308 1136 3316 1144
rect 3388 1136 3396 1144
rect 3628 1136 3636 1144
rect 3692 1136 3700 1144
rect 4524 1136 4532 1144
rect 4604 1136 4612 1144
rect 2076 1116 2084 1124
rect 2108 1116 2116 1124
rect 2476 1116 2484 1124
rect 2556 1116 2564 1124
rect 2812 1116 2820 1124
rect 3228 1116 3236 1124
rect 3244 1116 3252 1124
rect 4300 1116 4308 1124
rect 4668 1116 4676 1124
rect 4796 1116 4804 1124
rect 4908 1116 4916 1124
rect 252 1096 260 1104
rect 796 1096 804 1104
rect 988 1096 996 1104
rect 1100 1096 1108 1104
rect 2028 1096 2036 1104
rect 2044 1096 2052 1104
rect 2076 1096 2084 1104
rect 2156 1096 2164 1104
rect 2220 1096 2228 1104
rect 2236 1096 2244 1104
rect 2300 1096 2308 1104
rect 2348 1096 2356 1104
rect 2380 1096 2388 1104
rect 668 1076 676 1084
rect 844 1076 852 1084
rect 1084 1076 1092 1084
rect 1132 1076 1140 1084
rect 1164 1076 1172 1084
rect 1212 1076 1220 1084
rect 1500 1076 1508 1084
rect 2588 1096 2596 1104
rect 2636 1096 2644 1104
rect 2716 1096 2724 1104
rect 2892 1096 2900 1104
rect 3068 1096 3076 1104
rect 2924 1076 2932 1084
rect 3052 1076 3060 1084
rect 3244 1096 3252 1104
rect 3276 1096 3284 1104
rect 3660 1096 3668 1104
rect 3900 1096 3908 1104
rect 4220 1096 4228 1104
rect 4268 1096 4276 1104
rect 4316 1096 4324 1104
rect 4364 1096 4372 1104
rect 4412 1096 4420 1104
rect 44 1056 52 1064
rect 188 1056 196 1064
rect 524 1056 532 1064
rect 908 1056 916 1064
rect 1372 1056 1380 1064
rect 1804 1056 1812 1064
rect 2348 1056 2356 1064
rect 2380 1056 2388 1064
rect 2444 1056 2452 1064
rect 2956 1056 2964 1064
rect 3116 1076 3124 1084
rect 3516 1076 3524 1084
rect 3548 1076 3556 1084
rect 4940 1096 4948 1104
rect 5068 1096 5076 1104
rect 4524 1076 4532 1084
rect 3084 1056 3092 1064
rect 3100 1056 3108 1064
rect 3116 1056 3124 1064
rect 3180 1056 3188 1064
rect 3196 1056 3204 1064
rect 3500 1056 3508 1064
rect 3628 1056 3636 1064
rect 3692 1056 3700 1064
rect 3724 1056 3732 1064
rect 3788 1056 3796 1064
rect 3804 1056 3812 1064
rect 3916 1056 3924 1064
rect 4684 1056 4692 1064
rect 4828 1056 4836 1064
rect 4844 1056 4852 1064
rect 5004 1056 5012 1064
rect 220 1036 228 1044
rect 1020 1036 1028 1044
rect 1228 1036 1236 1044
rect 2012 1036 2020 1044
rect 2140 1036 2148 1044
rect 2220 1036 2228 1044
rect 2332 1036 2340 1044
rect 2396 1036 2404 1044
rect 2492 1036 2500 1044
rect 2524 1036 2532 1044
rect 44 1016 52 1024
rect 1148 1016 1156 1024
rect 1644 1016 1652 1024
rect 1676 1016 1684 1024
rect 1932 1016 1940 1024
rect 1980 1016 1988 1024
rect 2108 1016 2116 1024
rect 2364 1016 2372 1024
rect 2556 1016 2564 1024
rect 3004 1036 3012 1044
rect 3276 1036 3284 1044
rect 3324 1036 3332 1044
rect 3372 1036 3380 1044
rect 3436 1036 3444 1044
rect 3852 1036 3860 1044
rect 3868 1036 3876 1044
rect 3884 1036 3892 1044
rect 4236 1036 4244 1044
rect 4716 1036 4724 1044
rect 5004 1036 5012 1044
rect 5196 1036 5204 1044
rect 2796 1016 2804 1024
rect 2828 1016 2836 1024
rect 2876 1016 2884 1024
rect 3004 1016 3012 1024
rect 3484 1016 3492 1024
rect 3660 1016 3668 1024
rect 3708 1016 3716 1024
rect 3852 1016 3860 1024
rect 4636 1016 4644 1024
rect 5052 1016 5060 1024
rect 60 996 68 1004
rect 1244 996 1252 1004
rect 1308 996 1316 1004
rect 188 976 196 984
rect 460 976 468 984
rect 764 976 772 984
rect 876 976 884 984
rect 1148 976 1156 984
rect 1452 976 1460 984
rect 1468 976 1476 984
rect 1644 976 1652 984
rect 1676 976 1684 984
rect 1804 976 1812 984
rect 2508 996 2516 1004
rect 2764 996 2772 1004
rect 2908 996 2916 1004
rect 2972 996 2980 1004
rect 1884 976 1892 984
rect 2252 976 2260 984
rect 2524 976 2532 984
rect 2908 976 2916 984
rect 3180 996 3188 1004
rect 3628 996 3636 1004
rect 4252 996 4260 1004
rect 4300 996 4308 1004
rect 4588 996 4596 1004
rect 4748 996 4756 1004
rect 5116 996 5124 1004
rect 3596 976 3604 984
rect 3932 976 3940 984
rect 4332 976 4340 984
rect 4492 976 4500 984
rect 4716 976 4724 984
rect 4732 976 4740 984
rect 4892 976 4900 984
rect 5036 976 5044 984
rect 5180 976 5188 984
rect 140 956 148 964
rect 252 956 260 964
rect 636 956 644 964
rect 1788 956 1796 964
rect 1852 956 1860 964
rect 1868 956 1876 964
rect 1884 956 1892 964
rect 1948 956 1956 964
rect 1980 956 1988 964
rect 2380 956 2388 964
rect 2428 956 2436 964
rect 2524 956 2532 964
rect 2732 956 2740 964
rect 2828 956 2836 964
rect 2924 956 2932 964
rect 3276 956 3284 964
rect 3404 956 3412 964
rect 3468 956 3476 964
rect 3484 956 3492 964
rect 3628 956 3636 964
rect 3644 956 3652 964
rect 3980 956 3988 964
rect 4028 956 4036 964
rect 4140 956 4148 964
rect 4732 956 4740 964
rect 4972 956 4980 964
rect 5020 956 5028 964
rect 5164 956 5172 964
rect 12 936 20 944
rect 284 936 292 944
rect 300 936 308 944
rect 348 936 356 944
rect 460 936 468 944
rect 620 936 628 944
rect 1244 936 1252 944
rect 1276 936 1284 944
rect 1468 936 1476 944
rect 2012 936 2020 944
rect 2076 936 2084 944
rect 2108 936 2116 944
rect 2412 936 2420 944
rect 2460 936 2468 944
rect 2492 936 2500 944
rect 2556 936 2564 944
rect 2732 936 2740 944
rect 2780 936 2788 944
rect 2796 936 2804 944
rect 188 916 196 924
rect 444 916 452 924
rect 508 916 516 924
rect 540 916 548 924
rect 636 916 644 924
rect 716 916 724 924
rect 764 916 772 924
rect 1084 916 1092 924
rect 1100 916 1108 924
rect 1292 916 1300 924
rect 1628 916 1636 924
rect 1676 916 1684 924
rect 2156 916 2164 924
rect 2252 916 2260 924
rect 2284 916 2292 924
rect 2300 916 2308 924
rect 2412 916 2420 924
rect 2492 916 2500 924
rect 2636 916 2644 924
rect 2652 916 2660 924
rect 2668 916 2676 924
rect 2940 936 2948 944
rect 2956 936 2964 944
rect 3100 936 3108 944
rect 3372 936 3380 944
rect 3548 936 3556 944
rect 3564 936 3572 944
rect 3596 936 3604 944
rect 3948 936 3956 944
rect 2844 916 2852 924
rect 2892 916 2900 924
rect 3916 916 3924 924
rect 4188 936 4196 944
rect 4412 936 4420 944
rect 4460 936 4468 944
rect 4508 936 4516 944
rect 4524 936 4532 944
rect 4604 936 4612 944
rect 4876 936 4884 944
rect 4924 936 4932 944
rect 4060 916 4068 924
rect 5052 916 5060 924
rect 124 896 132 904
rect 220 896 228 904
rect 940 896 948 904
rect 956 896 964 904
rect 1052 896 1060 904
rect 1340 896 1348 904
rect 1468 896 1476 904
rect 2012 896 2020 904
rect 2172 896 2180 904
rect 2236 896 2244 904
rect 2252 896 2260 904
rect 2300 896 2308 904
rect 3148 896 3156 904
rect 3180 896 3188 904
rect 3756 896 3764 904
rect 3788 896 3796 904
rect 3804 896 3812 904
rect 3836 896 3844 904
rect 3948 896 3956 904
rect 4028 896 4036 904
rect 4892 896 4900 904
rect 5180 896 5188 904
rect 348 876 356 884
rect 444 876 452 884
rect 1164 876 1172 884
rect 1228 876 1236 884
rect 764 856 772 864
rect 1708 876 1716 884
rect 1740 876 1748 884
rect 1884 876 1892 884
rect 1932 876 1940 884
rect 2396 876 2404 884
rect 2412 876 2420 884
rect 2860 876 2868 884
rect 2892 876 2900 884
rect 2988 876 2996 884
rect 3212 876 3220 884
rect 3228 876 3236 884
rect 3308 876 3316 884
rect 4588 876 4596 884
rect 4844 876 4852 884
rect 5020 876 5028 884
rect 1388 856 1396 864
rect 1404 856 1412 864
rect 1740 856 1748 864
rect 1948 856 1956 864
rect 2140 856 2148 864
rect 2796 856 2804 864
rect 3260 856 3268 864
rect 3724 856 3732 864
rect 3820 856 3828 864
rect 1084 836 1092 844
rect 1148 836 1156 844
rect 1596 836 1604 844
rect 1708 836 1716 844
rect 2988 836 2996 844
rect 3164 836 3172 844
rect 3868 856 3876 864
rect 3884 856 3892 864
rect 4188 836 4196 844
rect 4300 836 4308 844
rect 5148 836 5156 844
rect 1356 816 1364 824
rect 1420 816 1428 824
rect 1724 816 1732 824
rect 2236 816 2244 824
rect 2652 816 2660 824
rect 2780 816 2788 824
rect 3004 816 3012 824
rect 3020 816 3028 824
rect 3036 816 3044 824
rect 3836 816 3844 824
rect 4044 816 4052 824
rect 4700 816 4708 824
rect 5052 816 5060 824
rect 172 796 180 804
rect 204 796 212 804
rect 236 796 244 804
rect 300 796 308 804
rect 1644 796 1652 804
rect 1740 796 1748 804
rect 1788 796 1796 804
rect 1916 796 1924 804
rect 2140 796 2148 804
rect 2172 796 2180 804
rect 2252 796 2260 804
rect 2332 796 2340 804
rect 3212 796 3220 804
rect 3244 796 3252 804
rect 3388 796 3396 804
rect 1356 776 1364 784
rect 1580 776 1588 784
rect 1964 776 1972 784
rect 4044 776 4052 784
rect 4252 776 4260 784
rect 4940 776 4948 784
rect 5180 776 5188 784
rect 364 756 372 764
rect 444 756 452 764
rect 844 756 852 764
rect 2236 756 2244 764
rect 2636 756 2644 764
rect 3180 756 3188 764
rect 3372 756 3380 764
rect 3436 756 3444 764
rect 3452 756 3460 764
rect 3900 756 3908 764
rect 3916 756 3924 764
rect 3948 756 3956 764
rect 3996 756 4004 764
rect 4044 756 4052 764
rect 4844 756 4852 764
rect 5196 756 5204 764
rect 284 736 292 744
rect 396 736 404 744
rect 460 736 468 744
rect 524 736 532 744
rect 764 736 772 744
rect 988 736 996 744
rect 1324 736 1332 744
rect 1404 736 1412 744
rect 1788 736 1796 744
rect 1852 736 1860 744
rect 2188 736 2196 744
rect 2220 736 2228 744
rect 2428 736 2436 744
rect 2556 736 2564 744
rect 2588 736 2596 744
rect 2748 736 2756 744
rect 3644 736 3652 744
rect 4028 736 4036 744
rect 4172 736 4180 744
rect 4220 736 4228 744
rect 4492 736 4500 744
rect 4620 736 4628 744
rect 4732 736 4740 744
rect 5164 736 5172 744
rect 140 716 148 724
rect 188 716 196 724
rect 476 716 484 724
rect 540 716 548 724
rect 828 716 836 724
rect 1500 716 1508 724
rect 1564 716 1572 724
rect 1612 716 1620 724
rect 2364 716 2372 724
rect 2412 716 2420 724
rect 2652 716 2660 724
rect 2748 716 2756 724
rect 2764 716 2772 724
rect 3052 716 3060 724
rect 3388 716 3396 724
rect 3756 716 3764 724
rect 3852 716 3860 724
rect 3868 716 3876 724
rect 4044 716 4052 724
rect 4060 716 4068 724
rect 4076 716 4084 724
rect 4156 716 4164 724
rect 4316 716 4324 724
rect 4684 716 4692 724
rect 4988 716 4996 724
rect 5036 716 5044 724
rect 796 696 804 704
rect 860 696 868 704
rect 1036 696 1044 704
rect 1084 696 1092 704
rect 1148 696 1156 704
rect 1196 696 1204 704
rect 1308 696 1316 704
rect 1340 696 1348 704
rect 2716 696 2724 704
rect 2780 696 2788 704
rect 2812 696 2820 704
rect 3212 696 3220 704
rect 3596 696 3604 704
rect 3724 696 3732 704
rect 3740 696 3748 704
rect 3756 696 3764 704
rect 4268 696 4276 704
rect 4412 696 4420 704
rect 4508 696 4516 704
rect 4620 696 4628 704
rect 4780 696 4788 704
rect 5084 696 5092 704
rect 316 676 324 684
rect 204 656 212 664
rect 492 676 500 684
rect 636 676 644 684
rect 668 676 676 684
rect 1644 676 1652 684
rect 1772 676 1780 684
rect 2380 676 2388 684
rect 2412 676 2420 684
rect 2476 676 2484 684
rect 2492 676 2500 684
rect 2572 676 2580 684
rect 2844 676 2852 684
rect 2860 676 2868 684
rect 2924 676 2932 684
rect 2940 676 2948 684
rect 2972 676 2980 684
rect 3516 676 3524 684
rect 3548 676 3556 684
rect 3564 676 3572 684
rect 3708 676 3716 684
rect 4556 676 4564 684
rect 4604 676 4612 684
rect 4636 676 4644 684
rect 5100 676 5108 684
rect 684 656 692 664
rect 1052 656 1060 664
rect 1084 656 1092 664
rect 1692 656 1700 664
rect 1724 656 1732 664
rect 1756 656 1764 664
rect 2828 656 2836 664
rect 3036 656 3044 664
rect 3052 656 3060 664
rect 4540 656 4548 664
rect 4796 656 4804 664
rect 4924 656 4932 664
rect 5004 656 5012 664
rect 5036 656 5044 664
rect 1004 636 1012 644
rect 1324 636 1332 644
rect 1340 636 1348 644
rect 1628 636 1636 644
rect 1660 636 1668 644
rect 1788 636 1796 644
rect 2060 636 2068 644
rect 2076 636 2084 644
rect 2172 636 2180 644
rect 2268 636 2276 644
rect 2908 636 2916 644
rect 3228 636 3236 644
rect 3836 636 3844 644
rect 4044 636 4052 644
rect 4108 636 4116 644
rect 4140 636 4148 644
rect 4828 636 4836 644
rect 172 616 180 624
rect 364 616 372 624
rect 844 616 852 624
rect 940 616 948 624
rect 956 616 964 624
rect 1084 616 1092 624
rect 1164 616 1172 624
rect 1196 616 1204 624
rect 1324 616 1332 624
rect 1548 616 1556 624
rect 1676 616 1684 624
rect 1772 616 1780 624
rect 1836 616 1844 624
rect 1916 616 1924 624
rect 1980 616 1988 624
rect 460 596 468 604
rect 556 596 564 604
rect 1004 596 1012 604
rect 1100 596 1108 604
rect 1244 596 1252 604
rect 1548 596 1556 604
rect 1612 596 1620 604
rect 2140 616 2148 624
rect 2220 616 2228 624
rect 2236 616 2244 624
rect 2268 616 2276 624
rect 2316 616 2324 624
rect 2380 616 2388 624
rect 2492 616 2500 624
rect 2732 616 2740 624
rect 2748 616 2756 624
rect 2988 616 2996 624
rect 3020 616 3028 624
rect 3036 616 3044 624
rect 2076 596 2084 604
rect 2140 596 2148 604
rect 2156 596 2164 604
rect 2172 596 2180 604
rect 2332 596 2340 604
rect 2364 596 2372 604
rect 2380 596 2388 604
rect 748 576 756 584
rect 764 576 772 584
rect 828 576 836 584
rect 1020 576 1028 584
rect 1932 576 1940 584
rect 1948 576 1956 584
rect 1996 576 2004 584
rect 2268 576 2276 584
rect 2476 596 2484 604
rect 2508 596 2516 604
rect 2588 596 2596 604
rect 2716 596 2724 604
rect 2860 596 2868 604
rect 2940 596 2948 604
rect 3068 596 3076 604
rect 3116 616 3124 624
rect 3324 616 3332 624
rect 3452 616 3460 624
rect 3484 616 3492 624
rect 3500 616 3508 624
rect 3692 616 3700 624
rect 3916 616 3924 624
rect 3948 616 3956 624
rect 4044 616 4052 624
rect 4156 616 4164 624
rect 4172 616 4180 624
rect 3180 596 3188 604
rect 2476 576 2484 584
rect 3180 576 3188 584
rect 3244 596 3252 604
rect 3308 596 3316 604
rect 3436 596 3444 604
rect 4012 596 4020 604
rect 4108 596 4116 604
rect 4188 596 4196 604
rect 4220 596 4228 604
rect 4252 596 4260 604
rect 4332 596 4340 604
rect 4492 596 4500 604
rect 4924 596 4932 604
rect 3324 576 3332 584
rect 3356 576 3364 584
rect 3436 576 3444 584
rect 3804 576 3812 584
rect 4076 576 4084 584
rect 4124 576 4132 584
rect 4348 576 4356 584
rect 4636 576 4644 584
rect 5052 576 5060 584
rect 5132 576 5140 584
rect 412 556 420 564
rect 684 556 692 564
rect 1036 556 1044 564
rect 1100 556 1108 564
rect 1244 556 1252 564
rect 1692 556 1700 564
rect 1724 556 1732 564
rect 1788 556 1796 564
rect 1932 556 1940 564
rect 1948 556 1956 564
rect 1964 556 1972 564
rect 1980 556 1988 564
rect 2044 556 2052 564
rect 2108 556 2116 564
rect 2124 556 2132 564
rect 2140 556 2148 564
rect 2268 556 2276 564
rect 2300 556 2308 564
rect 2348 556 2356 564
rect 2428 556 2436 564
rect 2556 556 2564 564
rect 2908 556 2916 564
rect 2988 556 2996 564
rect 3004 556 3012 564
rect 3036 556 3044 564
rect 3260 556 3268 564
rect 3292 556 3300 564
rect 3324 556 3332 564
rect 3580 556 3588 564
rect 3692 556 3700 564
rect 3708 556 3716 564
rect 4092 556 4100 564
rect 4108 556 4116 564
rect 4140 556 4148 564
rect 4188 556 4196 564
rect 4204 556 4212 564
rect 4524 556 4532 564
rect 4572 556 4580 564
rect 5068 556 5076 564
rect 108 536 116 544
rect 172 536 180 544
rect 252 536 260 544
rect 1084 536 1092 544
rect 1212 536 1220 544
rect 1228 536 1236 544
rect 1372 536 1380 544
rect 1404 536 1412 544
rect 1532 536 1540 544
rect 1580 536 1588 544
rect 1596 536 1604 544
rect 1644 536 1652 544
rect 1660 536 1668 544
rect 1740 536 1748 544
rect 3020 536 3028 544
rect 3068 536 3076 544
rect 188 516 196 524
rect 396 516 404 524
rect 508 516 516 524
rect 764 516 772 524
rect 780 516 788 524
rect 844 516 852 524
rect 892 516 900 524
rect 956 516 964 524
rect 1116 516 1124 524
rect 1276 516 1284 524
rect 1324 516 1332 524
rect 1356 516 1364 524
rect 1452 516 1460 524
rect 2460 516 2468 524
rect 2556 516 2564 524
rect 2780 516 2788 524
rect 2796 516 2804 524
rect 2956 516 2964 524
rect 2972 516 2980 524
rect 2988 516 2996 524
rect 3100 516 3108 524
rect 3212 516 3220 524
rect 3260 516 3268 524
rect 3292 516 3300 524
rect 3660 536 3668 544
rect 3788 536 3796 544
rect 3852 536 3860 544
rect 4284 536 4292 544
rect 4380 536 4388 544
rect 4412 536 4420 544
rect 4604 536 4612 544
rect 4652 536 4660 544
rect 4684 536 4692 544
rect 4796 536 4804 544
rect 5100 536 5108 544
rect 3340 516 3348 524
rect 3644 516 3652 524
rect 3884 516 3892 524
rect 4956 516 4964 524
rect 5148 516 5156 524
rect 268 496 276 504
rect 348 496 356 504
rect 588 496 596 504
rect 1404 496 1412 504
rect 1628 496 1636 504
rect 1772 496 1780 504
rect 2012 496 2020 504
rect 2060 496 2068 504
rect 2108 496 2116 504
rect 2124 496 2132 504
rect 2156 496 2164 504
rect 2812 496 2820 504
rect 2860 496 2868 504
rect 3132 496 3140 504
rect 3228 496 3236 504
rect 3292 496 3300 504
rect 3356 496 3364 504
rect 3452 496 3460 504
rect 3948 496 3956 504
rect 4092 496 4100 504
rect 4124 496 4132 504
rect 4492 496 4500 504
rect 5100 496 5108 504
rect 636 476 644 484
rect 876 476 884 484
rect 892 476 900 484
rect 940 476 948 484
rect 1420 476 1428 484
rect 2524 476 2532 484
rect 3036 476 3044 484
rect 3308 476 3316 484
rect 3484 476 3492 484
rect 3532 476 3540 484
rect 3708 476 3716 484
rect 3724 476 3732 484
rect 748 456 756 464
rect 1244 456 1252 464
rect 1644 456 1652 464
rect 1660 456 1668 464
rect 2316 456 2324 464
rect 2492 456 2500 464
rect 2636 456 2644 464
rect 572 436 580 444
rect 1868 436 1876 444
rect 1980 436 1988 444
rect 2060 436 2068 444
rect 2284 436 2292 444
rect 2412 436 2420 444
rect 2460 436 2468 444
rect 3084 456 3092 464
rect 4012 456 4020 464
rect 4812 456 4820 464
rect 12 416 20 424
rect 1100 416 1108 424
rect 1148 416 1156 424
rect 4748 416 4756 424
rect 5164 416 5172 424
rect 1212 396 1220 404
rect 908 376 916 384
rect 1660 396 1668 404
rect 2716 396 2724 404
rect 2748 396 2756 404
rect 2860 396 2868 404
rect 2908 396 2916 404
rect 2940 396 2948 404
rect 3052 396 3060 404
rect 1612 376 1620 384
rect 1836 376 1844 384
rect 2044 376 2052 384
rect 2380 376 2388 384
rect 3340 396 3348 404
rect 3164 376 3172 384
rect 4172 376 4180 384
rect 4332 376 4340 384
rect 1132 356 1140 364
rect 1564 356 1572 364
rect 1996 356 2004 364
rect 2012 356 2020 364
rect 2892 356 2900 364
rect 3116 356 3124 364
rect 3244 356 3252 364
rect 3836 356 3844 364
rect 620 336 628 344
rect 700 336 708 344
rect 812 336 820 344
rect 1244 336 1252 344
rect 1580 336 1588 344
rect 1628 336 1636 344
rect 1660 336 1668 344
rect 1692 336 1700 344
rect 1740 336 1748 344
rect 1820 336 1828 344
rect 1868 336 1876 344
rect 2060 336 2068 344
rect 2140 336 2148 344
rect 2252 336 2260 344
rect 2796 336 2804 344
rect 2812 336 2820 344
rect 3036 336 3044 344
rect 3820 336 3828 344
rect 3852 336 3860 344
rect 3996 336 4004 344
rect 4252 336 4260 344
rect 4284 336 4292 344
rect 4636 336 4644 344
rect 284 316 292 324
rect 364 316 372 324
rect 428 316 436 324
rect 796 316 804 324
rect 860 316 868 324
rect 940 316 948 324
rect 1084 316 1092 324
rect 1100 316 1108 324
rect 1116 316 1124 324
rect 1244 316 1252 324
rect 1292 316 1300 324
rect 1340 316 1348 324
rect 1372 316 1380 324
rect 2188 316 2196 324
rect 2204 316 2212 324
rect 2620 316 2628 324
rect 2636 316 2644 324
rect 2668 316 2676 324
rect 2716 316 2724 324
rect 2924 316 2932 324
rect 3020 316 3028 324
rect 3388 316 3396 324
rect 3468 316 3476 324
rect 3500 316 3508 324
rect 3788 316 3796 324
rect 3900 316 3908 324
rect 3948 316 3956 324
rect 4076 316 4084 324
rect 4108 316 4116 324
rect 4716 316 4724 324
rect 220 296 228 304
rect 716 296 724 304
rect 1260 296 1268 304
rect 2156 296 2164 304
rect 2188 296 2196 304
rect 2428 296 2436 304
rect 2508 296 2516 304
rect 2604 296 2612 304
rect 3548 296 3556 304
rect 3612 296 3620 304
rect 3804 296 3812 304
rect 3820 296 3828 304
rect 3868 296 3876 304
rect 3884 296 3892 304
rect 3980 296 3988 304
rect 4268 296 4276 304
rect 4556 296 4564 304
rect 4764 296 4772 304
rect 4844 296 4852 304
rect 4988 296 4996 304
rect 124 276 132 284
rect 684 276 692 284
rect 268 256 276 264
rect 332 256 340 264
rect 1356 276 1364 284
rect 1436 276 1444 284
rect 1468 276 1476 284
rect 1900 276 1908 284
rect 1948 276 1956 284
rect 1996 276 2004 284
rect 2044 276 2052 284
rect 2092 276 2100 284
rect 780 256 788 264
rect 2252 256 2260 264
rect 2380 276 2388 284
rect 2396 276 2404 284
rect 2460 276 2468 284
rect 2524 276 2532 284
rect 2588 276 2596 284
rect 2700 276 2708 284
rect 2796 276 2804 284
rect 2860 276 2868 284
rect 2412 256 2420 264
rect 2812 256 2820 264
rect 2844 256 2852 264
rect 2988 276 2996 284
rect 3068 276 3076 284
rect 3180 276 3188 284
rect 3196 276 3204 284
rect 3260 276 3268 284
rect 3276 276 3284 284
rect 4172 276 4180 284
rect 4620 276 4628 284
rect 4636 276 4644 284
rect 2908 256 2916 264
rect 3020 256 3028 264
rect 3068 256 3076 264
rect 3212 256 3220 264
rect 3356 256 3364 264
rect 3484 256 3492 264
rect 3676 256 3684 264
rect 4796 276 4804 284
rect 4876 276 4884 284
rect 5116 276 5124 284
rect 4892 256 4900 264
rect 5084 256 5092 264
rect 476 236 484 244
rect 876 236 884 244
rect 1068 236 1076 244
rect 1372 236 1380 244
rect 92 216 100 224
rect 828 216 836 224
rect 956 216 964 224
rect 972 216 980 224
rect 1260 216 1268 224
rect 1708 236 1716 244
rect 1868 236 1876 244
rect 1900 236 1908 244
rect 1964 236 1972 244
rect 2044 236 2052 244
rect 2076 236 2084 244
rect 2508 236 2516 244
rect 2972 236 2980 244
rect 3916 236 3924 244
rect 1724 216 1732 224
rect 1772 216 1780 224
rect 1804 216 1812 224
rect 1852 216 1860 224
rect 1980 216 1988 224
rect 1996 216 2004 224
rect 2028 216 2036 224
rect 2396 216 2404 224
rect 2444 216 2452 224
rect 2732 216 2740 224
rect 2860 216 2868 224
rect 2892 216 2900 224
rect 2924 216 2932 224
rect 2940 216 2948 224
rect 3004 216 3012 224
rect 3036 216 3044 224
rect 3132 216 3140 224
rect 3436 216 3444 224
rect 3692 216 3700 224
rect 3788 216 3796 224
rect 3804 216 3812 224
rect 3900 216 3908 224
rect 3996 216 4004 224
rect 4764 216 4772 224
rect 4796 216 4804 224
rect 924 196 932 204
rect 988 196 996 204
rect 1196 196 1204 204
rect 1564 196 1572 204
rect 348 176 356 184
rect 700 176 708 184
rect 748 176 756 184
rect 1132 176 1140 184
rect 1148 176 1156 184
rect 1628 176 1636 184
rect 2236 196 2244 204
rect 2476 196 2484 204
rect 2508 196 2516 204
rect 2572 196 2580 204
rect 2700 196 2708 204
rect 2876 196 2884 204
rect 2924 196 2932 204
rect 3052 196 3060 204
rect 3276 196 3284 204
rect 3468 196 3476 204
rect 4108 196 4116 204
rect 4156 196 4164 204
rect 4188 196 4196 204
rect 4204 196 4212 204
rect 4300 196 4308 204
rect 4316 196 4324 204
rect 4412 196 4420 204
rect 4844 196 4852 204
rect 4860 196 4868 204
rect 5004 196 5012 204
rect 2012 176 2020 184
rect 2060 176 2068 184
rect 2092 176 2100 184
rect 2412 176 2420 184
rect 3132 176 3140 184
rect 3196 176 3204 184
rect 3420 176 3428 184
rect 3452 176 3460 184
rect 3532 176 3540 184
rect 3580 176 3588 184
rect 3948 176 3956 184
rect 3980 176 3988 184
rect 4092 176 4100 184
rect 4140 176 4148 184
rect 4428 176 4436 184
rect 4668 176 4676 184
rect 140 156 148 164
rect 444 156 452 164
rect 476 156 484 164
rect 716 156 724 164
rect 732 156 740 164
rect 1052 156 1060 164
rect 1068 156 1076 164
rect 1196 156 1204 164
rect 1212 156 1220 164
rect 1228 156 1236 164
rect 1244 156 1252 164
rect 1804 156 1812 164
rect 2620 156 2628 164
rect 2652 156 2660 164
rect 2748 156 2756 164
rect 2828 156 2836 164
rect 3756 156 3764 164
rect 3964 156 3972 164
rect 4060 156 4068 164
rect 4524 156 4532 164
rect 4796 156 4804 164
rect 4812 156 4820 164
rect 4988 156 4996 164
rect 5068 156 5076 164
rect 5148 156 5156 164
rect 92 136 100 144
rect 300 136 308 144
rect 892 136 900 144
rect 908 136 916 144
rect 940 136 948 144
rect 1036 136 1044 144
rect 1484 136 1492 144
rect 1740 136 1748 144
rect 1756 136 1764 144
rect 1868 136 1876 144
rect 2012 136 2020 144
rect 2028 136 2036 144
rect 2204 136 2212 144
rect 3404 136 3412 144
rect 3436 136 3444 144
rect 3532 136 3540 144
rect 3548 136 3556 144
rect 3580 136 3588 144
rect 3612 136 3620 144
rect 3948 136 3956 144
rect 4156 136 4164 144
rect 4188 136 4196 144
rect 4540 136 4548 144
rect 4844 136 4852 144
rect 300 116 308 124
rect 492 116 500 124
rect 1660 116 1668 124
rect 2556 116 2564 124
rect 2604 116 2612 124
rect 2620 116 2628 124
rect 2684 116 2692 124
rect 2700 116 2708 124
rect 2812 116 2820 124
rect 2940 116 2948 124
rect 3148 116 3156 124
rect 3372 116 3380 124
rect 3404 116 3412 124
rect 3772 116 3780 124
rect 4028 116 4036 124
rect 4108 116 4116 124
rect 4780 116 4788 124
rect 4908 116 4916 124
rect 5052 116 5060 124
rect 268 96 276 104
rect 540 96 548 104
rect 604 96 612 104
rect 620 96 628 104
rect 668 96 676 104
rect 716 96 724 104
rect 924 76 932 84
rect 1180 96 1188 104
rect 1196 96 1204 104
rect 1676 96 1684 104
rect 1900 96 1908 104
rect 2220 96 2228 104
rect 3324 96 3332 104
rect 3660 96 3668 104
rect 3996 96 4004 104
rect 4060 96 4068 104
rect 4076 96 4084 104
rect 2444 76 2452 84
rect 2908 76 2916 84
rect 2940 76 2948 84
rect 3068 76 3076 84
rect 3084 76 3092 84
rect 3148 76 3156 84
rect 3196 76 3204 84
rect 3276 76 3284 84
rect 5212 76 5220 84
rect 1644 56 1652 64
rect 2988 56 2996 64
rect 2428 36 2436 44
rect 2812 36 2820 44
rect 1980 16 1988 24
rect 2012 16 2020 24
<< metal4 >>
rect 484 3537 492 3543
rect 93 3164 99 3296
rect 109 2904 115 3496
rect 157 3384 163 3476
rect 13 2304 19 2716
rect 45 2484 51 2716
rect 109 2704 115 2716
rect 61 2164 67 2596
rect 109 2524 115 2556
rect 93 1904 99 2396
rect 109 1684 115 2516
rect 77 1384 83 1516
rect 45 1024 51 1056
rect 61 1004 67 1296
rect 13 424 19 936
rect 77 724 83 1356
rect 93 1324 99 1536
rect 109 944 115 1676
rect 125 1364 131 1516
rect 141 964 147 2916
rect 157 2524 163 3336
rect 189 2744 195 3116
rect 205 3084 211 3136
rect 221 3064 227 3476
rect 253 3124 259 3296
rect 237 3064 243 3076
rect 205 2664 211 2676
rect 157 2084 163 2516
rect 221 2504 227 3056
rect 173 2164 179 2176
rect 189 2004 195 2496
rect 205 2184 211 2256
rect 173 1864 179 1896
rect 157 1744 163 1756
rect 221 1584 227 1776
rect 221 1524 227 1556
rect 237 1524 243 3056
rect 308 2917 316 2923
rect 285 2724 291 2896
rect 333 2884 339 3216
rect 285 2664 291 2696
rect 260 2657 268 2663
rect 285 2224 291 2596
rect 301 2364 307 2736
rect 276 2197 284 2203
rect 253 2164 259 2176
rect 237 1504 243 1516
rect 157 1364 163 1376
rect 212 1117 220 1123
rect 189 984 195 1056
rect 221 1024 227 1036
rect 109 544 115 936
rect 125 904 131 956
rect 141 724 147 956
rect 173 624 179 796
rect 189 724 195 916
rect 205 664 211 796
rect 125 284 131 576
rect 189 524 195 636
rect 221 304 227 896
rect 237 804 243 1416
rect 253 1104 259 1716
rect 269 1624 275 1856
rect 253 964 259 976
rect 253 324 259 536
rect 269 504 275 1296
rect 285 944 291 2136
rect 301 2104 307 2356
rect 317 2124 323 2656
rect 349 2524 355 3436
rect 381 3344 387 3516
rect 957 3484 963 3556
rect 381 2924 387 3336
rect 365 2584 371 2596
rect 333 2304 339 2516
rect 333 2144 339 2236
rect 317 1764 323 2116
rect 333 1744 339 2116
rect 349 1844 355 2436
rect 365 2124 371 2276
rect 308 1457 316 1463
rect 301 984 307 1436
rect 269 264 275 496
rect 285 324 291 736
rect 93 144 99 216
rect 132 157 140 163
rect 269 104 275 256
rect 301 144 307 796
rect 317 684 323 1456
rect 317 664 323 676
rect 333 264 339 1736
rect 349 1404 355 1676
rect 365 1484 371 2116
rect 381 1884 387 2676
rect 397 2644 403 3296
rect 413 2964 419 3456
rect 477 3444 483 3476
rect 557 3444 563 3456
rect 420 2897 428 2903
rect 413 2724 419 2856
rect 413 2644 419 2656
rect 429 2644 435 2656
rect 445 2544 451 3296
rect 461 3164 467 3196
rect 461 2984 467 3156
rect 461 2964 467 2976
rect 461 2704 467 2836
rect 477 2804 483 3336
rect 493 3284 499 3296
rect 461 2384 467 2656
rect 461 2264 467 2336
rect 477 2304 483 2796
rect 493 2764 499 3276
rect 509 2944 515 3276
rect 525 3104 531 3156
rect 541 2944 547 3016
rect 500 2737 508 2743
rect 493 2504 499 2676
rect 509 2664 515 2676
rect 509 2304 515 2336
rect 493 2284 499 2296
rect 525 2264 531 2916
rect 653 2904 659 3476
rect 797 3464 803 3476
rect 852 3457 860 3463
rect 701 3104 707 3116
rect 685 2984 691 3036
rect 596 2897 604 2903
rect 637 2724 643 2736
rect 589 2684 595 2696
rect 541 2644 547 2676
rect 541 2564 547 2576
rect 557 2544 563 2576
rect 541 2384 547 2396
rect 541 2264 547 2376
rect 477 2244 483 2263
rect 429 2124 435 2136
rect 381 1564 387 1876
rect 349 944 355 1276
rect 365 1264 371 1436
rect 349 884 355 916
rect 349 504 355 876
rect 365 624 371 756
rect 397 744 403 2056
rect 413 1124 419 2116
rect 429 1344 435 2096
rect 477 1964 483 2136
rect 477 1884 483 1956
rect 445 1324 451 1796
rect 461 1784 467 1856
rect 477 1704 483 1776
rect 493 1724 499 2116
rect 509 1764 515 1776
rect 541 1744 547 2236
rect 477 1664 483 1683
rect 372 317 380 323
rect 397 284 403 516
rect 413 364 419 556
rect 429 324 435 936
rect 445 924 451 1316
rect 461 1124 467 1516
rect 461 984 467 1116
rect 445 884 451 916
rect 445 764 451 776
rect 461 744 467 936
rect 477 724 483 1476
rect 493 1344 499 1376
rect 525 1344 531 1676
rect 493 984 499 1116
rect 525 1064 531 1256
rect 541 924 547 1736
rect 557 1464 563 2516
rect 573 2324 579 2676
rect 573 2104 579 2296
rect 573 1924 579 2096
rect 573 1684 579 1916
rect 557 1404 563 1436
rect 573 1424 579 1596
rect 589 1364 595 2396
rect 621 2164 627 2396
rect 637 2264 643 2716
rect 605 2124 611 2156
rect 605 1544 611 2056
rect 605 1524 611 1536
rect 516 917 524 923
rect 525 724 531 736
rect 548 717 556 723
rect 452 597 460 603
rect 429 304 435 316
rect 477 244 483 276
rect 349 164 355 176
rect 468 157 476 163
rect 445 144 451 156
rect 285 123 291 136
rect 493 124 499 676
rect 548 597 556 603
rect 573 444 579 1356
rect 589 504 595 1116
rect 285 117 300 123
rect 605 104 611 1516
rect 621 944 627 1476
rect 637 1144 643 2256
rect 653 1904 659 2496
rect 669 2244 675 2256
rect 669 2204 675 2216
rect 669 2124 675 2176
rect 653 1544 659 1676
rect 685 1604 691 2976
rect 717 2944 723 3416
rect 733 3344 739 3376
rect 765 3324 771 3336
rect 733 3124 739 3276
rect 765 3224 771 3236
rect 717 2864 723 2876
rect 701 2724 707 2756
rect 708 2517 716 2523
rect 733 2304 739 3116
rect 756 3077 764 3083
rect 781 2984 787 3456
rect 797 3344 803 3436
rect 941 3364 947 3456
rect 957 3364 963 3456
rect 829 3304 835 3336
rect 797 3044 803 3096
rect 797 2963 803 2996
rect 781 2957 803 2963
rect 781 2924 787 2957
rect 749 2664 755 2696
rect 749 2624 755 2636
rect 701 2184 707 2236
rect 749 2184 755 2596
rect 653 1104 659 1536
rect 669 1384 675 1416
rect 669 1344 675 1356
rect 701 1324 707 1336
rect 637 924 643 956
rect 669 684 675 1076
rect 644 677 652 683
rect 621 284 627 336
rect 669 104 675 676
rect 685 664 691 1316
rect 685 284 691 556
rect 701 224 707 336
rect 717 304 723 916
rect 733 244 739 1996
rect 749 1964 755 2156
rect 765 2104 771 2476
rect 765 1924 771 2096
rect 781 1944 787 2896
rect 797 2684 803 2936
rect 813 2864 819 3076
rect 829 2684 835 3296
rect 845 2924 851 3256
rect 797 2544 803 2676
rect 797 2124 803 2536
rect 749 1524 755 1796
rect 749 584 755 1476
rect 765 1284 771 1916
rect 765 984 771 1236
rect 781 1124 787 1936
rect 797 1884 803 2116
rect 765 924 771 936
rect 765 744 771 756
rect 781 744 787 1116
rect 797 1104 803 1736
rect 813 1204 819 2656
rect 829 2564 835 2576
rect 829 2524 835 2536
rect 829 2044 835 2316
rect 845 2284 851 2916
rect 861 2684 867 3336
rect 893 3304 899 3316
rect 861 2364 867 2656
rect 877 2564 883 3296
rect 893 3144 899 3296
rect 877 2484 883 2556
rect 861 2284 867 2296
rect 845 2064 851 2156
rect 836 2017 844 2023
rect 829 1704 835 1996
rect 845 1724 851 1796
rect 829 1524 835 1696
rect 797 704 803 1096
rect 765 564 771 576
rect 749 543 755 556
rect 781 543 787 596
rect 749 537 787 543
rect 749 324 755 456
rect 765 264 771 516
rect 797 324 803 696
rect 813 344 819 1176
rect 829 724 835 1516
rect 845 1084 851 1696
rect 861 1504 867 1976
rect 861 1484 867 1496
rect 877 1484 883 2436
rect 893 2124 899 3116
rect 909 3104 915 3336
rect 909 2884 915 3096
rect 909 1984 915 2876
rect 925 2744 931 3076
rect 941 3044 947 3136
rect 925 2504 931 2716
rect 941 2544 947 2956
rect 957 2604 963 3276
rect 973 3224 979 3496
rect 973 3064 979 3216
rect 973 2944 979 2956
rect 973 2884 979 2916
rect 973 2664 979 2676
rect 925 2364 931 2496
rect 916 1957 924 1963
rect 909 1884 915 1896
rect 893 1644 899 1656
rect 893 1464 899 1636
rect 925 1544 931 1756
rect 941 1704 947 2476
rect 957 2144 963 2596
rect 973 2504 979 2636
rect 989 2324 995 3536
rect 1396 3517 1404 3523
rect 1821 3504 1827 3516
rect 1037 3424 1043 3456
rect 1085 3424 1091 3436
rect 1005 3377 1043 3383
rect 1005 3364 1011 3377
rect 1037 3363 1043 3377
rect 1101 3364 1107 3416
rect 1037 3357 1052 3363
rect 1117 3344 1123 3396
rect 1044 3337 1052 3343
rect 1005 3084 1011 3096
rect 1005 2864 1011 3016
rect 1021 2784 1027 3156
rect 1037 3044 1043 3096
rect 973 2284 979 2296
rect 957 1824 963 1856
rect 861 1324 867 1456
rect 861 1224 867 1296
rect 845 624 851 756
rect 861 704 867 1196
rect 909 1044 915 1056
rect 772 257 780 263
rect 701 164 707 176
rect 733 164 739 236
rect 829 224 835 576
rect 717 144 723 156
rect 845 144 851 516
rect 877 484 883 976
rect 893 524 899 556
rect 893 464 899 476
rect 909 344 915 376
rect 877 244 883 316
rect 925 204 931 1496
rect 941 904 947 1496
rect 973 1464 979 1976
rect 989 1964 995 2116
rect 989 1484 995 1516
rect 989 1464 995 1476
rect 1005 1284 1011 2716
rect 1021 1904 1027 2676
rect 1037 2624 1043 2916
rect 1076 2897 1084 2903
rect 1101 2724 1107 3316
rect 1117 3064 1123 3296
rect 1133 3064 1139 3096
rect 1053 2524 1059 2616
rect 1037 2284 1043 2496
rect 1053 2244 1059 2276
rect 1037 1844 1043 2116
rect 1053 1904 1059 1916
rect 1037 1344 1043 1556
rect 989 1084 995 1096
rect 957 904 963 936
rect 989 744 995 1056
rect 941 604 947 616
rect 941 484 947 556
rect 957 524 963 616
rect 941 324 947 336
rect 909 144 915 156
rect 884 137 892 143
rect 941 124 947 136
rect 957 124 963 216
rect 989 204 995 736
rect 1005 604 1011 616
rect 1021 584 1027 1036
rect 1037 704 1043 1336
rect 1053 904 1059 1856
rect 1069 1464 1075 2536
rect 1085 1724 1091 2716
rect 1101 2284 1107 2316
rect 1101 1924 1107 2096
rect 1117 2004 1123 3056
rect 1133 2904 1139 2916
rect 1149 2704 1155 3296
rect 1133 2684 1139 2696
rect 1133 2444 1139 2576
rect 1149 2504 1155 2696
rect 1133 2384 1139 2396
rect 1133 2324 1139 2336
rect 1133 2104 1139 2216
rect 1149 2164 1155 2496
rect 1165 2184 1171 3396
rect 1181 3084 1187 3456
rect 1197 3264 1203 3336
rect 1085 1364 1091 1716
rect 1085 1304 1091 1356
rect 1069 1264 1075 1276
rect 1037 564 1043 696
rect 1037 144 1043 556
rect 1053 164 1059 656
rect 1069 244 1075 1256
rect 1085 1084 1091 1296
rect 1101 1104 1107 1876
rect 1117 1824 1123 1836
rect 1117 1784 1123 1796
rect 1117 1704 1123 1716
rect 1133 1524 1139 2036
rect 1149 1524 1155 2156
rect 1181 2124 1187 3076
rect 1197 2724 1203 2736
rect 1165 2004 1171 2016
rect 1165 1744 1171 1796
rect 1085 924 1091 1076
rect 1101 924 1107 1096
rect 1085 704 1091 836
rect 1085 644 1091 656
rect 1092 617 1100 623
rect 1085 544 1091 556
rect 1117 524 1123 1376
rect 1133 1303 1139 1436
rect 1149 1324 1155 1516
rect 1165 1464 1171 1696
rect 1181 1544 1187 2116
rect 1133 1297 1155 1303
rect 1149 1264 1155 1297
rect 1133 1124 1139 1216
rect 1133 1064 1139 1076
rect 1101 344 1107 416
rect 1133 364 1139 1036
rect 1149 1024 1155 1236
rect 1165 1144 1171 1436
rect 1165 1124 1171 1136
rect 1165 1064 1171 1076
rect 1149 944 1155 976
rect 1165 884 1171 936
rect 1156 837 1164 843
rect 1165 624 1171 796
rect 1149 424 1155 576
rect 1101 324 1107 336
rect 1085 303 1091 316
rect 1117 303 1123 316
rect 1085 297 1123 303
rect 1133 184 1139 196
rect 1156 177 1164 183
rect 1069 144 1075 156
rect 717 104 723 116
rect 532 97 540 103
rect 621 84 627 96
rect 957 84 963 116
rect 1181 104 1187 1536
rect 1197 704 1203 2696
rect 1213 2244 1219 3336
rect 1229 3044 1235 3496
rect 1245 3484 1251 3496
rect 1213 1324 1219 2236
rect 1229 1864 1235 3036
rect 1245 2984 1251 3356
rect 1261 3344 1267 3356
rect 1277 3104 1283 3476
rect 1293 3264 1299 3396
rect 1309 3164 1315 3176
rect 1309 3124 1315 3136
rect 1245 2884 1251 2896
rect 1245 2684 1251 2776
rect 1245 2024 1251 2456
rect 1261 2184 1267 3076
rect 1261 2124 1267 2156
rect 1277 2044 1283 3096
rect 1309 3044 1315 3056
rect 1309 2624 1315 2976
rect 1293 2544 1299 2596
rect 1309 2544 1315 2556
rect 1268 2017 1276 2023
rect 1229 1424 1235 1576
rect 1261 1544 1267 1816
rect 1277 1804 1283 1816
rect 1277 1704 1283 1716
rect 1293 1704 1299 2516
rect 1309 2304 1315 2516
rect 1309 1924 1315 2016
rect 1325 1764 1331 3376
rect 1341 3124 1347 3356
rect 1357 3164 1363 3176
rect 1357 3124 1363 3136
rect 1341 2944 1347 2976
rect 1341 2884 1347 2916
rect 1341 2604 1347 2616
rect 1341 2424 1347 2456
rect 1341 2204 1347 2336
rect 1341 2104 1347 2156
rect 1341 1904 1347 1923
rect 1277 1664 1283 1676
rect 1293 1664 1299 1696
rect 1213 1084 1219 1156
rect 1213 904 1219 1076
rect 1229 1044 1235 1416
rect 1245 1004 1251 1316
rect 1261 1164 1267 1456
rect 1229 884 1235 896
rect 1245 604 1251 936
rect 1213 544 1219 576
rect 1197 184 1203 196
rect 1213 164 1219 396
rect 1229 264 1235 536
rect 1245 464 1251 556
rect 1245 264 1251 316
rect 1261 304 1267 1156
rect 1277 944 1283 1596
rect 1309 1504 1315 1676
rect 1309 1344 1315 1496
rect 1325 1384 1331 1756
rect 1341 1744 1347 1856
rect 1341 1384 1347 1396
rect 1325 1344 1331 1376
rect 1277 524 1283 876
rect 1293 324 1299 916
rect 1309 884 1315 996
rect 1325 744 1331 1236
rect 1357 1124 1363 2956
rect 1373 2724 1379 3276
rect 1405 3124 1411 3136
rect 1389 2584 1395 3116
rect 1405 2904 1411 2976
rect 1405 2564 1411 2896
rect 1421 2704 1427 3496
rect 1453 3284 1459 3336
rect 1485 3044 1491 3116
rect 1453 2944 1459 2976
rect 1437 2904 1443 2916
rect 1444 2877 1452 2883
rect 1373 2164 1379 2556
rect 1389 2484 1395 2556
rect 1405 2344 1411 2536
rect 1437 2404 1443 2576
rect 1421 2304 1427 2316
rect 1389 2204 1395 2216
rect 1380 2097 1388 2103
rect 1373 1844 1379 1896
rect 1389 1864 1395 1916
rect 1405 1864 1411 1896
rect 1373 1804 1379 1816
rect 1389 1744 1395 1756
rect 1421 1464 1427 2296
rect 1437 2284 1443 2296
rect 1437 1904 1443 1936
rect 1373 1244 1379 1456
rect 1373 1064 1379 1196
rect 1341 704 1347 896
rect 1389 884 1395 1296
rect 1405 1144 1411 1396
rect 1421 1224 1427 1296
rect 1421 1144 1427 1156
rect 1357 784 1363 816
rect 1316 697 1324 703
rect 1316 617 1324 623
rect 1325 524 1331 536
rect 1341 324 1347 636
rect 1373 424 1379 536
rect 1389 404 1395 856
rect 1405 684 1411 736
rect 1405 544 1411 576
rect 1405 384 1411 496
rect 1421 484 1427 816
rect 1357 264 1363 276
rect 1229 164 1235 256
rect 1373 244 1379 316
rect 1437 284 1443 1696
rect 1453 984 1459 2676
rect 1469 2544 1475 2616
rect 1469 2104 1475 2536
rect 1485 2503 1491 2896
rect 1501 2684 1507 3376
rect 1533 3044 1539 3076
rect 1485 2497 1507 2503
rect 1485 2104 1491 2476
rect 1485 1824 1491 2056
rect 1501 1924 1507 2497
rect 1517 2484 1523 2496
rect 1533 2444 1539 2876
rect 1533 2304 1539 2316
rect 1517 2284 1523 2296
rect 1524 2197 1532 2203
rect 1517 2164 1523 2176
rect 1517 1904 1523 1956
rect 1501 1864 1507 1896
rect 1533 1844 1539 2036
rect 1549 1904 1555 3356
rect 1565 2724 1571 3256
rect 1645 3064 1651 3376
rect 1677 3284 1683 3336
rect 1629 2944 1635 3056
rect 1661 2944 1667 3276
rect 1693 3144 1699 3356
rect 1684 3117 1692 3123
rect 1597 2904 1603 2916
rect 1581 2824 1587 2836
rect 1565 2584 1571 2616
rect 1581 2584 1587 2616
rect 1565 2484 1571 2556
rect 1581 2464 1587 2476
rect 1565 2444 1571 2456
rect 1581 2344 1587 2436
rect 1565 2184 1571 2276
rect 1581 2264 1587 2276
rect 1565 2064 1571 2136
rect 1549 1844 1555 1856
rect 1517 1804 1523 1836
rect 1517 1664 1523 1756
rect 1469 1524 1475 1556
rect 1517 1524 1523 1656
rect 1469 1124 1475 1516
rect 1501 1324 1507 1356
rect 1485 1204 1491 1316
rect 1469 964 1475 976
rect 1469 924 1475 936
rect 1469 884 1475 896
rect 1453 504 1459 516
rect 1469 264 1475 276
rect 1268 217 1283 223
rect 1245 164 1251 216
rect 1197 104 1203 156
rect 1357 124 1363 176
rect 1485 144 1491 1156
rect 1501 1024 1507 1076
rect 1508 717 1516 723
rect 1533 684 1539 1816
rect 1549 1764 1555 1816
rect 1533 544 1539 676
rect 1549 624 1555 1676
rect 1565 1384 1571 1956
rect 1581 1504 1587 2256
rect 1597 2084 1603 2696
rect 1613 2204 1619 2816
rect 1629 2624 1635 2756
rect 1629 2464 1635 2476
rect 1629 2204 1635 2256
rect 1613 2104 1619 2156
rect 1620 2057 1628 2063
rect 1629 1944 1635 2016
rect 1613 1904 1619 1936
rect 1645 1844 1651 2896
rect 1661 2044 1667 2936
rect 1709 2904 1715 3456
rect 1725 3364 1731 3376
rect 1725 3144 1731 3276
rect 1677 2464 1683 2576
rect 1693 2044 1699 2896
rect 1709 2864 1715 2876
rect 1709 2504 1715 2576
rect 1725 2564 1731 3136
rect 1741 2524 1747 3416
rect 1725 2264 1731 2496
rect 1757 2344 1763 3396
rect 1805 3344 1811 3476
rect 1789 3124 1795 3336
rect 1773 3044 1779 3096
rect 1773 2904 1779 2936
rect 1789 2823 1795 3096
rect 1821 2904 1827 2936
rect 1837 2924 1843 3476
rect 1885 3344 1891 3556
rect 1917 3444 1923 3496
rect 1860 3337 1868 3343
rect 1860 3237 1868 3243
rect 1869 3044 1875 3076
rect 1805 2864 1811 2876
rect 1780 2817 1795 2823
rect 1805 2704 1811 2816
rect 1709 2204 1715 2216
rect 1741 2184 1747 2316
rect 1757 2264 1763 2296
rect 1716 2157 1724 2163
rect 1604 1837 1612 1843
rect 1597 1804 1603 1816
rect 1613 1644 1619 1656
rect 1604 1497 1612 1503
rect 1629 1484 1635 1836
rect 1645 1644 1651 1736
rect 1645 1584 1651 1636
rect 1645 1484 1651 1556
rect 1581 1364 1587 1376
rect 1581 964 1587 1116
rect 1597 844 1603 1456
rect 1613 1384 1619 1396
rect 1629 1324 1635 1396
rect 1645 1384 1651 1396
rect 1565 704 1571 716
rect 1533 524 1539 536
rect 1549 164 1555 596
rect 1581 544 1587 776
rect 1613 724 1619 1196
rect 1645 1144 1651 1156
rect 1645 1043 1651 1116
rect 1629 1037 1651 1043
rect 1629 924 1635 1037
rect 1645 1004 1651 1016
rect 1645 804 1651 976
rect 1645 684 1651 796
rect 1661 644 1667 2016
rect 1693 1904 1699 1916
rect 1677 1524 1683 1636
rect 1677 1404 1683 1476
rect 1693 1404 1699 1896
rect 1709 1744 1715 2116
rect 1725 2024 1731 2056
rect 1709 1624 1715 1736
rect 1677 1064 1683 1396
rect 1677 1024 1683 1036
rect 1677 964 1683 976
rect 1677 864 1683 916
rect 1613 384 1619 596
rect 1629 504 1635 636
rect 1677 624 1683 676
rect 1693 664 1699 1376
rect 1709 1124 1715 1516
rect 1709 884 1715 1116
rect 1645 544 1651 596
rect 1661 544 1667 556
rect 1565 204 1571 356
rect 1581 344 1587 376
rect 1629 264 1635 336
rect 1629 164 1635 176
rect 925 64 931 76
rect 1645 64 1651 456
rect 1661 384 1667 396
rect 1661 284 1667 336
rect 1661 124 1667 156
rect 1677 124 1683 616
rect 1693 564 1699 576
rect 1693 284 1699 336
rect 1709 244 1715 836
rect 1725 824 1731 1936
rect 1741 1924 1747 2176
rect 1757 1984 1763 2176
rect 1741 1324 1747 1856
rect 1757 1824 1763 1936
rect 1757 1504 1763 1596
rect 1741 1144 1747 1176
rect 1741 884 1747 916
rect 1741 844 1747 856
rect 1725 644 1731 656
rect 1725 544 1731 556
rect 1741 544 1747 796
rect 1757 664 1763 1356
rect 1773 684 1779 2636
rect 1789 2564 1795 2576
rect 1805 2404 1811 2416
rect 1789 2264 1795 2336
rect 1789 2064 1795 2236
rect 1805 2223 1811 2376
rect 1821 2284 1827 2896
rect 1837 2584 1843 2656
rect 1853 2644 1859 3016
rect 1837 2564 1843 2576
rect 1837 2504 1843 2536
rect 1805 2217 1820 2223
rect 1789 1904 1795 1936
rect 1789 1744 1795 1876
rect 1789 1704 1795 1716
rect 1805 1604 1811 2156
rect 1821 1884 1827 1896
rect 1821 1864 1827 1876
rect 1821 1764 1827 1836
rect 1789 1564 1795 1576
rect 1789 1504 1795 1516
rect 1789 964 1795 1476
rect 1805 1284 1811 1576
rect 1821 1484 1827 1696
rect 1837 1404 1843 2476
rect 1853 2324 1859 2636
rect 1869 2304 1875 2996
rect 1885 2904 1891 3336
rect 1901 3004 1907 3236
rect 1901 2904 1907 2916
rect 1885 2524 1891 2896
rect 1901 2704 1907 2736
rect 1869 2124 1875 2256
rect 1853 1904 1859 2076
rect 1885 2064 1891 2516
rect 1917 2364 1923 3436
rect 1933 3204 1939 3236
rect 1933 3004 1939 3096
rect 1965 3024 1971 3516
rect 2061 3504 2067 3516
rect 2029 3364 2035 3456
rect 1933 2864 1939 2876
rect 1933 2464 1939 2616
rect 1949 2564 1955 2936
rect 1981 2884 1987 3216
rect 2013 2944 2019 3276
rect 2029 3104 2035 3156
rect 1965 2624 1971 2796
rect 1981 2584 1987 2816
rect 2004 2737 2012 2743
rect 1997 2624 2003 2676
rect 1981 2504 1987 2536
rect 1901 2004 1907 2316
rect 1933 2224 1939 2356
rect 1949 2244 1955 2436
rect 1917 2204 1923 2216
rect 1885 1917 1900 1923
rect 1853 1544 1859 1896
rect 1869 1824 1875 1916
rect 1885 1804 1891 1917
rect 1885 1604 1891 1696
rect 1885 1464 1891 1536
rect 1837 1384 1843 1396
rect 1901 1384 1907 1816
rect 1917 1624 1923 1976
rect 1933 1824 1939 2056
rect 1949 1964 1955 2236
rect 1965 2064 1971 2476
rect 1981 2164 1987 2196
rect 1997 2164 2003 2556
rect 2013 2284 2019 2716
rect 2029 2684 2035 2876
rect 2045 2664 2051 2936
rect 2045 2564 2051 2596
rect 2029 2544 2035 2556
rect 2029 2403 2035 2436
rect 2029 2397 2044 2403
rect 1997 2144 2003 2156
rect 1917 1544 1923 1596
rect 1933 1484 1939 1776
rect 1949 1504 1955 1916
rect 1933 1444 1939 1476
rect 1901 1364 1907 1376
rect 1876 1357 1884 1363
rect 1885 1344 1891 1356
rect 1869 1324 1875 1336
rect 1965 1324 1971 1896
rect 1997 1824 2003 1876
rect 1981 1744 1987 1816
rect 1997 1744 2003 1776
rect 2013 1724 2019 2276
rect 2029 2104 2035 2236
rect 2045 2204 2051 2236
rect 2045 2144 2051 2176
rect 2029 2024 2035 2056
rect 2045 2003 2051 2136
rect 2061 2103 2067 3496
rect 2077 3444 2083 3456
rect 2109 3284 2115 3356
rect 2125 3344 2131 3356
rect 2173 3284 2179 3356
rect 2109 3104 2115 3276
rect 2189 3184 2195 3336
rect 2205 3264 2211 3516
rect 2228 3437 2236 3443
rect 2301 3424 2307 3616
rect 2509 3444 2515 3456
rect 2525 3444 2531 3536
rect 2740 3517 2748 3523
rect 2852 3517 2860 3523
rect 2653 3484 2659 3496
rect 2685 3484 2691 3516
rect 2829 3503 2835 3516
rect 2877 3503 2883 3516
rect 2765 3497 2819 3503
rect 2829 3497 2883 3503
rect 2541 3444 2547 3476
rect 2372 3437 2380 3443
rect 2237 3364 2243 3396
rect 2221 3337 2236 3343
rect 2221 3284 2227 3337
rect 2077 2824 2083 3096
rect 2100 2997 2108 3003
rect 2093 2904 2099 2936
rect 2109 2864 2115 2876
rect 2084 2777 2092 2783
rect 2093 2624 2099 2636
rect 2077 2464 2083 2576
rect 2077 2124 2083 2296
rect 2061 2097 2083 2103
rect 2029 1997 2051 2003
rect 2029 1764 2035 1997
rect 1844 1317 1852 1323
rect 1885 1284 1891 1296
rect 1805 1064 1811 1076
rect 1789 804 1795 916
rect 1789 744 1795 756
rect 1805 684 1811 976
rect 1741 304 1747 336
rect 1725 224 1731 296
rect 1757 144 1763 656
rect 1789 644 1795 656
rect 1773 504 1779 616
rect 1821 344 1827 1176
rect 1837 904 1843 1176
rect 1853 964 1859 1036
rect 1869 964 1875 1156
rect 1885 984 1891 1116
rect 1885 944 1891 956
rect 1837 644 1843 896
rect 1885 884 1891 896
rect 1837 624 1843 636
rect 1805 224 1811 296
rect 1853 224 1859 736
rect 1869 344 1875 376
rect 1901 284 1907 1316
rect 1917 1124 1923 1136
rect 1933 1024 1939 1296
rect 1965 1224 1971 1236
rect 1981 1204 1987 1716
rect 1997 1704 2003 1716
rect 1997 1364 2003 1476
rect 1949 984 1955 1196
rect 1949 964 1955 976
rect 1917 804 1923 816
rect 1917 764 1923 796
rect 1933 784 1939 876
rect 1949 804 1955 856
rect 1917 624 1923 636
rect 1949 584 1955 796
rect 1965 784 1971 1136
rect 1981 964 1987 1016
rect 1981 684 1987 956
rect 1981 624 1987 656
rect 1997 584 2003 1276
rect 2013 1044 2019 1716
rect 2045 1504 2051 1956
rect 2061 1904 2067 2016
rect 2061 1483 2067 1836
rect 2045 1477 2067 1483
rect 2029 1404 2035 1456
rect 2029 1264 2035 1356
rect 2045 1264 2051 1477
rect 2061 1264 2067 1356
rect 2045 1104 2051 1256
rect 2013 904 2019 936
rect 1933 484 1939 556
rect 1949 544 1955 556
rect 1949 264 1955 276
rect 1965 244 1971 556
rect 1981 504 1987 556
rect 2013 504 2019 896
rect 1981 444 1987 456
rect 1997 364 2003 376
rect 2013 364 2019 396
rect 1997 264 2003 276
rect 1876 237 1884 243
rect 1677 104 1683 116
rect 1741 44 1747 136
rect 1805 104 1811 156
rect 1869 104 1875 136
rect 1901 104 1907 236
rect 1981 224 1987 236
rect 1997 24 2003 216
rect 2013 184 2019 356
rect 2029 224 2035 1096
rect 2045 964 2051 1036
rect 2061 644 2067 1156
rect 2077 1124 2083 2097
rect 2093 2084 2099 2616
rect 2125 2384 2131 3116
rect 2141 2944 2147 2996
rect 2141 2924 2147 2936
rect 2173 2844 2179 3096
rect 2205 3084 2211 3096
rect 2221 3084 2227 3116
rect 2189 2864 2195 2916
rect 2125 2304 2131 2316
rect 2109 2064 2115 2276
rect 2141 2184 2147 2736
rect 2157 2664 2163 2776
rect 2173 2624 2179 2656
rect 2189 2564 2195 2596
rect 2164 2557 2172 2563
rect 2205 2484 2211 3056
rect 2221 2864 2227 2876
rect 2237 2844 2243 3256
rect 2269 3184 2275 3416
rect 2333 3384 2339 3436
rect 2365 3344 2371 3396
rect 2253 2724 2259 3096
rect 2269 2924 2275 3076
rect 2237 2544 2243 2596
rect 2141 2144 2147 2176
rect 2093 1904 2099 2056
rect 2109 2004 2115 2016
rect 2093 1744 2099 1896
rect 2109 1884 2115 1896
rect 2109 1804 2115 1816
rect 2093 1564 2099 1736
rect 2109 1424 2115 1736
rect 2100 1357 2108 1363
rect 2077 1084 2083 1096
rect 2077 644 2083 656
rect 2045 564 2051 636
rect 2077 564 2083 596
rect 2045 384 2051 496
rect 2061 444 2067 496
rect 2077 344 2083 556
rect 2061 304 2067 336
rect 2093 284 2099 1316
rect 2109 1024 2115 1096
rect 2109 564 2115 936
rect 2125 564 2131 2036
rect 2141 1844 2147 1996
rect 2141 1784 2147 1816
rect 2141 1664 2147 1676
rect 2141 1564 2147 1616
rect 2141 1324 2147 1396
rect 2157 1364 2163 2376
rect 2173 1984 2179 2216
rect 2189 2124 2195 2136
rect 2205 2084 2211 2316
rect 2173 1883 2179 1936
rect 2189 1904 2195 1996
rect 2205 1944 2211 2076
rect 2173 1877 2195 1883
rect 2189 1824 2195 1877
rect 2173 1684 2179 1816
rect 2173 1524 2179 1676
rect 2189 1584 2195 1616
rect 2205 1604 2211 1736
rect 2189 1504 2195 1536
rect 2173 1464 2179 1496
rect 2173 1364 2179 1396
rect 2157 1304 2163 1356
rect 2141 1224 2147 1256
rect 2173 1224 2179 1256
rect 2141 1044 2147 1156
rect 2157 924 2163 1096
rect 2173 1084 2179 1216
rect 2141 864 2147 916
rect 2173 904 2179 956
rect 2173 804 2179 816
rect 2141 784 2147 796
rect 2141 624 2147 636
rect 2157 604 2163 796
rect 2189 764 2195 1416
rect 2173 644 2179 736
rect 2141 583 2147 596
rect 2173 583 2179 596
rect 2141 577 2179 583
rect 2125 464 2131 496
rect 2141 344 2147 556
rect 2189 504 2195 736
rect 2157 304 2163 496
rect 2205 324 2211 1536
rect 2221 1104 2227 2356
rect 2237 2284 2243 2496
rect 2253 2304 2259 2716
rect 2269 2644 2275 2916
rect 2285 2824 2291 3256
rect 2365 2984 2371 3276
rect 2381 3084 2387 3356
rect 2301 2917 2339 2923
rect 2301 2904 2307 2917
rect 2333 2904 2339 2917
rect 2308 2637 2316 2643
rect 2301 2504 2307 2616
rect 2333 2564 2339 2596
rect 2276 2497 2284 2503
rect 2237 2204 2243 2276
rect 2237 1744 2243 2096
rect 2253 1704 2259 2296
rect 2269 2224 2275 2376
rect 2269 2124 2275 2196
rect 2285 2004 2291 2216
rect 2301 2204 2307 2236
rect 2269 1944 2275 1976
rect 2269 1764 2275 1776
rect 2237 1564 2243 1616
rect 2237 1444 2243 1456
rect 2237 1164 2243 1356
rect 2237 1104 2243 1136
rect 2221 764 2227 1036
rect 2253 984 2259 1676
rect 2253 924 2259 976
rect 2237 904 2243 916
rect 2237 804 2243 816
rect 2221 624 2227 736
rect 2237 664 2243 756
rect 2180 297 2188 303
rect 2045 244 2051 276
rect 2068 237 2076 243
rect 2052 177 2060 183
rect 2100 177 2108 183
rect 2013 144 2019 176
rect 2029 124 2035 136
rect 2205 124 2211 136
rect 2221 104 2227 496
rect 2237 484 2243 616
rect 2237 204 2243 456
rect 2253 344 2259 796
rect 2269 644 2275 1696
rect 2285 1624 2291 1756
rect 2301 1664 2307 2016
rect 2317 1784 2323 2536
rect 2365 2504 2371 2976
rect 2381 2884 2387 2936
rect 2301 1644 2307 1656
rect 2285 1484 2291 1516
rect 2301 1404 2307 1456
rect 2285 1184 2291 1396
rect 2317 1344 2323 1756
rect 2333 1384 2339 1856
rect 2349 1304 2355 1836
rect 2365 1684 2371 2496
rect 2381 2104 2387 2656
rect 2397 2324 2403 3436
rect 2413 3224 2419 3356
rect 2445 3344 2451 3356
rect 2429 2904 2435 2936
rect 2429 2824 2435 2876
rect 2429 2724 2435 2736
rect 2413 2604 2419 2616
rect 2413 2284 2419 2496
rect 2445 2444 2451 3056
rect 2397 2144 2403 2216
rect 2381 1804 2387 2096
rect 2413 2044 2419 2096
rect 2413 1964 2419 1976
rect 2397 1784 2403 1956
rect 2413 1704 2419 1956
rect 2381 1644 2387 1696
rect 2365 1524 2371 1616
rect 2365 1444 2371 1456
rect 2317 1204 2323 1256
rect 2349 1104 2355 1136
rect 2292 1097 2300 1103
rect 2317 964 2323 1036
rect 2301 924 2307 956
rect 2269 584 2275 596
rect 2285 564 2291 916
rect 2301 564 2307 896
rect 2333 804 2339 1036
rect 2317 604 2323 616
rect 2269 543 2275 556
rect 2301 544 2307 556
rect 2269 537 2291 543
rect 2285 523 2291 537
rect 2317 523 2323 556
rect 2285 517 2323 523
rect 2333 484 2339 596
rect 2349 564 2355 1056
rect 2365 1024 2371 1436
rect 2381 1104 2387 1616
rect 2397 1604 2403 1636
rect 2413 1584 2419 1596
rect 2413 1524 2419 1536
rect 2413 1444 2419 1476
rect 2397 1384 2403 1436
rect 2413 1364 2419 1396
rect 2397 1324 2403 1336
rect 2381 1044 2387 1056
rect 2397 1044 2403 1176
rect 2381 944 2387 956
rect 2397 903 2403 956
rect 2413 944 2419 1356
rect 2429 1344 2435 2396
rect 2461 2304 2467 3116
rect 2477 3044 2483 3056
rect 2477 2324 2483 2956
rect 2445 2064 2451 2236
rect 2445 2024 2451 2036
rect 2445 1944 2451 1956
rect 2461 1884 2467 2296
rect 2477 2284 2483 2296
rect 2477 2204 2483 2236
rect 2477 2124 2483 2136
rect 2445 1704 2451 1836
rect 2461 1824 2467 1836
rect 2445 1504 2451 1516
rect 2429 1284 2435 1296
rect 2429 1204 2435 1216
rect 2429 1164 2435 1176
rect 2445 1064 2451 1356
rect 2429 937 2435 956
rect 2420 917 2428 923
rect 2397 897 2419 903
rect 2413 884 2419 897
rect 2365 684 2371 716
rect 2381 664 2387 676
rect 2381 624 2387 656
rect 2365 604 2371 616
rect 2285 444 2291 456
rect 2381 424 2387 596
rect 2253 284 2259 336
rect 2397 284 2403 876
rect 2413 724 2419 736
rect 2429 663 2435 676
rect 2413 657 2435 663
rect 2413 604 2419 657
rect 2429 564 2435 596
rect 2413 264 2419 436
rect 2397 224 2403 256
rect 2013 24 2019 96
rect 2429 44 2435 296
rect 2445 224 2451 1056
rect 2461 944 2467 1676
rect 2477 1124 2483 2036
rect 2493 1364 2499 3436
rect 2509 3384 2515 3396
rect 2516 3357 2531 3363
rect 2525 3284 2531 3357
rect 2557 3304 2563 3476
rect 2557 3284 2563 3296
rect 2509 3044 2515 3216
rect 2541 3044 2547 3156
rect 2525 2964 2531 3016
rect 2557 2964 2563 3156
rect 2509 2584 2515 2796
rect 2541 2623 2547 2936
rect 2557 2804 2563 2856
rect 2557 2704 2563 2736
rect 2525 2617 2547 2623
rect 2525 2564 2531 2617
rect 2516 2537 2524 2543
rect 2525 2284 2531 2296
rect 2509 1824 2515 1956
rect 2509 1504 2515 1556
rect 2493 1264 2499 1336
rect 2493 1217 2499 1236
rect 2461 544 2467 936
rect 2477 684 2483 1116
rect 2493 1044 2499 1196
rect 2509 1004 2515 1296
rect 2525 1044 2531 2196
rect 2541 1204 2547 2596
rect 2557 2564 2563 2596
rect 2557 2484 2563 2496
rect 2557 2264 2563 2296
rect 2573 2223 2579 3476
rect 2765 3424 2771 3497
rect 2740 3397 2748 3403
rect 2589 3304 2595 3376
rect 2612 3357 2620 3363
rect 2637 3304 2643 3356
rect 2717 3144 2723 3356
rect 2765 3324 2771 3356
rect 2669 3097 2707 3103
rect 2653 3044 2659 3076
rect 2669 3064 2675 3097
rect 2589 2944 2595 2996
rect 2605 2884 2611 3036
rect 2669 2964 2675 3036
rect 2589 2724 2595 2856
rect 2589 2304 2595 2536
rect 2605 2424 2611 2856
rect 2621 2724 2627 2736
rect 2589 2264 2595 2276
rect 2573 2217 2595 2223
rect 2557 2204 2563 2216
rect 2557 1424 2563 2176
rect 2573 2144 2579 2156
rect 2573 2044 2579 2116
rect 2589 2024 2595 2217
rect 2573 1944 2579 1956
rect 2573 1884 2579 1896
rect 2573 1504 2579 1856
rect 2589 1743 2595 1896
rect 2605 1804 2611 2376
rect 2621 2084 2627 2696
rect 2621 1804 2627 2076
rect 2637 1924 2643 2716
rect 2669 2664 2675 2956
rect 2653 2124 2659 2656
rect 2685 2544 2691 3076
rect 2701 3064 2707 3097
rect 2717 3084 2723 3136
rect 2781 3084 2787 3476
rect 2813 3424 2819 3497
rect 2893 3483 2899 3616
rect 2877 3477 2899 3483
rect 2701 2924 2707 2956
rect 2701 2744 2707 2776
rect 2701 2644 2707 2656
rect 2685 2504 2691 2516
rect 2701 2504 2707 2556
rect 2669 2464 2675 2476
rect 2669 2344 2675 2416
rect 2701 2404 2707 2416
rect 2669 2224 2675 2276
rect 2589 1737 2611 1743
rect 2589 1644 2595 1696
rect 2573 1444 2579 1456
rect 2573 1364 2579 1416
rect 2541 1144 2547 1176
rect 2525 964 2531 976
rect 2493 944 2499 956
rect 2493 804 2499 916
rect 2493 684 2499 736
rect 2484 617 2492 623
rect 2509 604 2515 936
rect 2461 524 2467 536
rect 2461 404 2467 436
rect 2461 264 2467 276
rect 2477 204 2483 496
rect 2493 464 2499 576
rect 2445 84 2451 116
rect 2493 24 2499 396
rect 2509 304 2515 596
rect 2525 484 2531 956
rect 2541 304 2547 1136
rect 2557 1104 2563 1116
rect 2557 1024 2563 1076
rect 2557 924 2563 936
rect 2557 744 2563 796
rect 2573 684 2579 1296
rect 2589 1104 2595 1516
rect 2605 1384 2611 1737
rect 2589 1004 2595 1076
rect 2589 744 2595 756
rect 2580 597 2588 603
rect 2557 564 2563 576
rect 2557 504 2563 516
rect 2605 304 2611 1196
rect 2621 324 2627 1736
rect 2637 1284 2643 1916
rect 2653 1724 2659 2116
rect 2669 2024 2675 2156
rect 2685 2084 2691 2256
rect 2701 2184 2707 2356
rect 2685 2024 2691 2036
rect 2653 1544 2659 1716
rect 2669 1504 2675 2016
rect 2685 1964 2691 1996
rect 2685 1584 2691 1916
rect 2701 1904 2707 1936
rect 2717 1784 2723 3076
rect 2749 3024 2755 3076
rect 2781 3064 2787 3076
rect 2797 3044 2803 3056
rect 2765 2944 2771 2956
rect 2765 2824 2771 2916
rect 2781 2884 2787 2956
rect 2797 2824 2803 3036
rect 2733 1924 2739 2756
rect 2749 2724 2755 2776
rect 2749 2564 2755 2676
rect 2765 2384 2771 2816
rect 2781 2444 2787 2736
rect 2797 2664 2803 2736
rect 2797 2544 2803 2556
rect 2797 2424 2803 2476
rect 2749 2284 2755 2296
rect 2749 2224 2755 2236
rect 2749 2104 2755 2176
rect 2749 2004 2755 2036
rect 2765 1964 2771 2216
rect 2749 1924 2755 1956
rect 2733 1824 2739 1916
rect 2749 1804 2755 1856
rect 2717 1724 2723 1756
rect 2669 1424 2675 1456
rect 2669 1344 2675 1356
rect 2644 1217 2652 1223
rect 2637 1064 2643 1096
rect 2637 924 2643 996
rect 2653 964 2659 1176
rect 2669 924 2675 1276
rect 2653 824 2659 916
rect 2637 624 2643 756
rect 2653 724 2659 736
rect 2637 404 2643 456
rect 2525 284 2531 296
rect 2509 244 2515 256
rect 2509 144 2515 196
rect 2573 164 2579 196
rect 2605 124 2611 296
rect 2653 264 2659 476
rect 2669 324 2675 916
rect 2653 164 2659 256
rect 2621 124 2627 156
rect 2685 124 2691 1576
rect 2701 284 2707 1676
rect 2717 1124 2723 1716
rect 2749 1704 2755 1716
rect 2733 1424 2739 1696
rect 2749 1604 2755 1656
rect 2765 1644 2771 1896
rect 2749 1504 2755 1536
rect 2749 1364 2755 1416
rect 2733 1304 2739 1336
rect 2717 704 2723 1096
rect 2733 1004 2739 1156
rect 2749 1064 2755 1216
rect 2765 1144 2771 1596
rect 2733 924 2739 936
rect 2749 884 2755 1056
rect 2717 604 2723 676
rect 2733 624 2739 756
rect 2749 744 2755 776
rect 2765 724 2771 996
rect 2781 944 2787 2276
rect 2797 2124 2803 2296
rect 2813 2284 2819 3136
rect 2829 2944 2835 2956
rect 2813 2124 2819 2236
rect 2797 1904 2803 2036
rect 2797 1844 2803 1896
rect 2797 1764 2803 1796
rect 2797 1704 2803 1716
rect 2797 1424 2803 1596
rect 2813 1344 2819 2096
rect 2829 1484 2835 2816
rect 2845 2684 2851 3076
rect 2861 2964 2867 3316
rect 2877 3004 2883 3477
rect 2877 2844 2883 2916
rect 2845 2424 2851 2636
rect 2877 2504 2883 2836
rect 2893 2764 2899 3356
rect 2909 3024 2915 3396
rect 2973 3384 2979 3416
rect 2925 3304 2931 3316
rect 2989 3264 2995 3296
rect 2957 2944 2963 2996
rect 2973 2964 2979 3056
rect 2925 2864 2931 2876
rect 2941 2684 2947 2896
rect 2989 2884 2995 3116
rect 2964 2817 2972 2823
rect 2861 2484 2867 2496
rect 2877 2464 2883 2476
rect 2893 2424 2899 2656
rect 2909 2624 2915 2636
rect 2877 2324 2883 2416
rect 2852 2297 2860 2303
rect 2877 2284 2883 2296
rect 2909 2284 2915 2516
rect 2845 2264 2851 2276
rect 2845 2224 2851 2236
rect 2845 2157 2899 2163
rect 2845 2144 2851 2157
rect 2845 2104 2851 2116
rect 2845 1964 2851 2056
rect 2813 1124 2819 1336
rect 2829 1304 2835 1416
rect 2845 1284 2851 1896
rect 2861 1824 2867 2136
rect 2877 2124 2883 2136
rect 2893 2124 2899 2157
rect 2909 2124 2915 2196
rect 2925 2164 2931 2536
rect 2941 2204 2947 2676
rect 2957 2364 2963 2676
rect 2909 2024 2915 2096
rect 2877 1964 2883 1976
rect 2893 1964 2899 2016
rect 2877 1864 2883 1896
rect 2877 1764 2883 1816
rect 2909 1804 2915 2016
rect 2925 1904 2931 2156
rect 2941 2124 2947 2156
rect 2941 2024 2947 2076
rect 2893 1784 2899 1796
rect 2861 1704 2867 1756
rect 2900 1717 2908 1723
rect 2877 1684 2883 1716
rect 2909 1644 2915 1696
rect 2861 1584 2867 1636
rect 2909 1424 2915 1496
rect 2868 1417 2876 1423
rect 2893 1364 2899 1416
rect 2925 1304 2931 1896
rect 2941 1884 2947 1896
rect 2941 1584 2947 1836
rect 2957 1784 2963 2356
rect 2973 2124 2979 2656
rect 2989 2504 2995 2876
rect 3005 2704 3011 3396
rect 3021 3144 3027 3316
rect 3037 3244 3043 3416
rect 3037 3144 3043 3156
rect 3021 3084 3027 3136
rect 3021 2904 3027 2936
rect 3037 2864 3043 2936
rect 2989 2284 2995 2456
rect 2989 1884 2995 2216
rect 3005 2044 3011 2696
rect 3037 2664 3043 2796
rect 3021 2484 3027 2516
rect 3021 2444 3027 2456
rect 3037 2304 3043 2496
rect 3053 2364 3059 3136
rect 3069 2664 3075 3496
rect 3085 3324 3091 3516
rect 3101 3184 3107 3556
rect 3117 3504 3123 3516
rect 3133 3424 3139 3516
rect 3117 3364 3123 3396
rect 3133 3384 3139 3403
rect 3124 3317 3132 3323
rect 3069 2484 3075 2596
rect 3085 2284 3091 3056
rect 3101 2744 3107 3016
rect 3117 2924 3123 3196
rect 3133 2924 3139 3096
rect 3149 2904 3155 3456
rect 3213 3424 3219 3516
rect 3325 3444 3331 3516
rect 3188 3417 3203 3423
rect 3188 3397 3196 3403
rect 3229 3384 3235 3396
rect 3101 2684 3107 2696
rect 3101 2524 3107 2636
rect 3117 2504 3123 2896
rect 3133 2564 3139 2716
rect 3133 2484 3139 2556
rect 3149 2484 3155 2596
rect 3021 2264 3027 2276
rect 3021 1884 3027 1896
rect 2973 1824 2979 1856
rect 3005 1824 3011 1876
rect 3021 1824 3027 1836
rect 2957 1704 2963 1716
rect 2957 1624 2963 1676
rect 2941 1364 2947 1536
rect 2957 1464 2963 1536
rect 2973 1464 2979 1796
rect 2989 1764 2995 1776
rect 3005 1724 3011 1756
rect 2989 1664 2995 1696
rect 3021 1664 3027 1676
rect 3005 1644 3011 1656
rect 3005 1524 3011 1576
rect 2989 1384 2995 1516
rect 2797 1004 2803 1016
rect 2797 944 2803 956
rect 2781 824 2787 836
rect 2797 824 2803 856
rect 2749 684 2755 716
rect 2781 684 2787 696
rect 2797 664 2803 736
rect 2813 704 2819 1116
rect 2829 1024 2835 1136
rect 2877 1024 2883 1096
rect 2829 944 2835 956
rect 2836 917 2844 923
rect 2861 884 2867 956
rect 2749 624 2755 636
rect 2781 504 2787 516
rect 2813 504 2819 516
rect 2717 244 2723 316
rect 2733 224 2739 236
rect 2701 124 2707 196
rect 2749 164 2755 396
rect 2797 284 2803 336
rect 2813 324 2819 336
rect 2813 244 2819 256
rect 2813 124 2819 176
rect 2829 164 2835 656
rect 2845 264 2851 676
rect 2861 604 2867 656
rect 2861 324 2867 396
rect 2861 224 2867 236
rect 2877 204 2883 936
rect 2893 924 2899 1096
rect 2909 1004 2915 1256
rect 2925 1084 2931 1296
rect 2893 884 2899 896
rect 2893 464 2899 876
rect 2909 684 2915 976
rect 2925 964 2931 1076
rect 2941 944 2947 1356
rect 2989 1344 2995 1356
rect 3005 1344 3011 1396
rect 2957 1064 2963 1136
rect 3005 1124 3011 1216
rect 2973 1004 2979 1116
rect 3005 1044 3011 1076
rect 2941 684 2947 876
rect 2909 644 2915 676
rect 2909 564 2915 576
rect 2925 404 2931 676
rect 2941 604 2947 616
rect 2957 524 2963 896
rect 2973 684 2979 996
rect 2989 844 2995 876
rect 3005 824 3011 836
rect 3021 824 3027 1656
rect 3037 1184 3043 1916
rect 3053 1744 3059 1896
rect 3069 1824 3075 2016
rect 3085 1844 3091 2276
rect 3101 2124 3107 2476
rect 3117 2404 3123 2476
rect 3133 2444 3139 2456
rect 3133 2124 3139 2156
rect 3149 2144 3155 2156
rect 3149 2084 3155 2116
rect 3053 1504 3059 1736
rect 3069 1483 3075 1696
rect 3085 1684 3091 1776
rect 3053 1477 3075 1483
rect 3053 1084 3059 1477
rect 3069 1344 3075 1396
rect 3069 1044 3075 1096
rect 3085 1064 3091 1376
rect 3101 1344 3107 1816
rect 3117 1804 3123 1856
rect 3133 1724 3139 1736
rect 3149 1724 3155 2016
rect 3165 1904 3171 3316
rect 3181 3244 3187 3356
rect 3181 2944 3187 3236
rect 3197 2964 3203 3016
rect 3181 2904 3187 2916
rect 3181 2744 3187 2756
rect 3197 2684 3203 2716
rect 3181 2564 3187 2596
rect 3197 2504 3203 2596
rect 3213 2564 3219 3056
rect 3229 2724 3235 2736
rect 3213 2304 3219 2516
rect 3229 2504 3235 2516
rect 3181 2144 3187 2256
rect 3197 2184 3203 2196
rect 3181 1924 3187 2136
rect 3197 1944 3203 1956
rect 3213 1904 3219 2296
rect 3229 2204 3235 2376
rect 3229 1923 3235 2136
rect 3245 1944 3251 3396
rect 3293 3264 3299 3296
rect 3261 2984 3267 3256
rect 3277 2924 3283 2936
rect 3277 2724 3283 2756
rect 3261 2644 3267 2656
rect 3261 2504 3267 2536
rect 3261 2264 3267 2456
rect 3293 2304 3299 3036
rect 3309 2924 3315 3436
rect 3373 3424 3379 3616
rect 3677 3544 3683 3576
rect 3469 3484 3475 3496
rect 3405 3444 3411 3476
rect 3517 3464 3523 3516
rect 3533 3464 3539 3536
rect 3389 3404 3395 3436
rect 3453 3424 3459 3456
rect 3501 3443 3507 3456
rect 3549 3444 3555 3516
rect 3565 3464 3571 3496
rect 3501 3437 3523 3443
rect 3517 3424 3523 3437
rect 3492 3417 3500 3423
rect 3325 3364 3331 3376
rect 3341 3344 3347 3356
rect 3341 3044 3347 3056
rect 3357 2944 3363 3096
rect 3373 3084 3379 3096
rect 3325 2924 3331 2936
rect 3309 2884 3315 2896
rect 3309 2564 3315 2776
rect 3325 2704 3331 2896
rect 3357 2624 3363 2796
rect 3309 2464 3315 2516
rect 3325 2444 3331 2516
rect 3341 2444 3347 2536
rect 3357 2444 3363 2536
rect 3373 2524 3379 3056
rect 3389 2904 3395 3396
rect 3565 3384 3571 3396
rect 3405 3104 3411 3336
rect 3437 3304 3443 3336
rect 3485 3264 3491 3276
rect 3405 3044 3411 3056
rect 3437 3024 3443 3256
rect 3453 3044 3459 3056
rect 3453 2984 3459 3016
rect 3412 2897 3420 2903
rect 3277 2264 3283 2296
rect 3325 2244 3331 2256
rect 3229 1917 3251 1923
rect 3229 1884 3235 1896
rect 3245 1804 3251 1917
rect 3261 1864 3267 2136
rect 3277 2104 3283 2116
rect 3293 2084 3299 2096
rect 3309 2024 3315 2236
rect 3284 2017 3292 2023
rect 3309 1964 3315 2016
rect 3293 1864 3299 1896
rect 3325 1844 3331 2216
rect 3341 2164 3347 2336
rect 3357 2184 3363 2316
rect 3341 1844 3347 1936
rect 3101 1244 3107 1256
rect 3101 1144 3107 1176
rect 3117 1084 3123 1636
rect 3149 1564 3155 1576
rect 3149 1424 3155 1436
rect 3101 944 3107 1056
rect 2973 524 2979 676
rect 3021 624 3027 796
rect 3037 624 3043 656
rect 2989 524 2995 556
rect 2941 404 2947 476
rect 2893 224 2899 356
rect 2909 264 2915 396
rect 2925 284 2931 316
rect 2925 224 2931 236
rect 2941 224 2947 236
rect 2877 184 2883 196
rect 2893 163 2899 176
rect 2925 164 2931 196
rect 2957 164 2963 516
rect 2973 244 2979 516
rect 3005 324 3011 556
rect 3021 324 3027 536
rect 3037 484 3043 556
rect 3037 344 3043 476
rect 3053 464 3059 656
rect 3069 604 3075 816
rect 3069 504 3075 536
rect 2868 157 2899 163
rect 2557 84 2563 116
rect 2813 44 2819 96
rect 2941 84 2947 116
rect 2989 64 2995 276
rect 3005 224 3011 276
rect 3021 264 3027 316
rect 3037 304 3043 336
rect 3037 224 3043 296
rect 3053 204 3059 396
rect 3069 284 3075 496
rect 3085 464 3091 796
rect 3117 624 3123 1056
rect 3140 897 3148 903
rect 3165 844 3171 1576
rect 3181 1424 3187 1436
rect 3197 1384 3203 1796
rect 3229 1704 3235 1736
rect 3245 1644 3251 1696
rect 3261 1644 3267 1836
rect 3245 1544 3251 1576
rect 3220 1537 3228 1543
rect 3261 1524 3267 1616
rect 3293 1544 3299 1696
rect 3213 1424 3219 1456
rect 3181 1064 3187 1076
rect 3181 904 3187 916
rect 3181 764 3187 776
rect 3181 604 3187 616
rect 3181 564 3187 576
rect 3101 484 3107 516
rect 3133 484 3139 496
rect 3085 304 3091 396
rect 3165 324 3171 376
rect 3069 84 3075 256
rect 3085 84 3091 296
rect 3181 284 3187 316
rect 3197 284 3203 1056
rect 3213 884 3219 1296
rect 3245 1124 3251 1516
rect 3293 1484 3299 1516
rect 3309 1464 3315 1836
rect 3325 1824 3331 1836
rect 3325 1484 3331 1796
rect 3229 1084 3235 1116
rect 3245 1104 3251 1116
rect 3229 864 3235 876
rect 3261 864 3267 1436
rect 3277 1104 3283 1376
rect 3277 1044 3283 1076
rect 3236 797 3244 803
rect 3213 704 3219 796
rect 3213 524 3219 696
rect 3245 604 3251 616
rect 3213 264 3219 516
rect 3229 504 3235 596
rect 3261 564 3267 776
rect 3261 484 3267 516
rect 3133 224 3139 236
rect 3229 224 3235 356
rect 3245 284 3251 356
rect 3277 284 3283 956
rect 3293 784 3299 1436
rect 3309 1224 3315 1456
rect 3325 1204 3331 1476
rect 3341 1424 3347 1436
rect 3341 1344 3347 1376
rect 3357 1364 3363 1716
rect 3373 1644 3379 2436
rect 3389 2344 3395 2896
rect 3421 2864 3427 2876
rect 3405 2564 3411 2816
rect 3405 2304 3411 2496
rect 3389 1984 3395 2256
rect 3405 2224 3411 2236
rect 3389 1844 3395 1876
rect 3389 1704 3395 1756
rect 3389 1604 3395 1616
rect 3389 1444 3395 1556
rect 3373 1323 3379 1356
rect 3357 1317 3379 1323
rect 3357 1304 3363 1317
rect 3309 1144 3315 1156
rect 3325 1044 3331 1156
rect 3293 524 3299 556
rect 3293 484 3299 496
rect 3309 484 3315 596
rect 3325 584 3331 616
rect 3133 104 3139 176
rect 3197 144 3203 176
rect 3149 124 3155 136
rect 3277 84 3283 196
rect 3325 104 3331 556
rect 3341 524 3347 1216
rect 3373 1204 3379 1216
rect 3389 1204 3395 1296
rect 3357 584 3363 1076
rect 3373 1024 3379 1036
rect 3389 804 3395 1136
rect 3405 964 3411 1936
rect 3373 664 3379 756
rect 3364 497 3372 503
rect 3092 77 3100 83
rect 3156 77 3164 83
rect 3197 64 3203 76
rect 3341 44 3347 396
rect 3373 284 3379 496
rect 3389 324 3395 716
rect 3357 264 3363 276
rect 3405 144 3411 956
rect 3421 584 3427 2736
rect 3437 1164 3443 2716
rect 3453 2624 3459 2656
rect 3453 2124 3459 2556
rect 3469 2404 3475 3056
rect 3485 2984 3491 3256
rect 3485 2924 3491 2936
rect 3485 2724 3491 2776
rect 3469 2324 3475 2336
rect 3485 2324 3491 2616
rect 3469 2244 3475 2256
rect 3453 2084 3459 2116
rect 3469 2104 3475 2176
rect 3460 2037 3468 2043
rect 3453 1704 3459 1816
rect 3469 1764 3475 1936
rect 3485 1904 3491 2276
rect 3501 1884 3507 3356
rect 3524 3137 3555 3143
rect 3549 3124 3555 3137
rect 3517 2064 3523 3116
rect 3533 3064 3539 3076
rect 3549 3044 3555 3063
rect 3533 2984 3539 2996
rect 3565 2964 3571 3316
rect 3581 3124 3587 3496
rect 3629 3464 3635 3496
rect 3645 3464 3651 3536
rect 3853 3484 3859 3516
rect 3997 3497 4099 3503
rect 3965 3484 3971 3496
rect 3997 3483 4003 3497
rect 3988 3477 4003 3483
rect 3652 3457 3660 3463
rect 3597 3444 3603 3456
rect 3581 3104 3587 3116
rect 3533 2584 3539 2796
rect 3549 2563 3555 2916
rect 3565 2904 3571 2936
rect 3533 2557 3555 2563
rect 3533 2504 3539 2557
rect 3533 2024 3539 2336
rect 3549 2284 3555 2516
rect 3517 1944 3523 2016
rect 3453 1444 3459 1596
rect 3453 1204 3459 1396
rect 3437 1044 3443 1056
rect 3469 964 3475 1696
rect 3485 1544 3491 1596
rect 3501 1064 3507 1876
rect 3517 1624 3523 1756
rect 3517 1544 3523 1596
rect 3517 1444 3523 1516
rect 3533 1484 3539 1996
rect 3517 1064 3523 1076
rect 3485 944 3491 956
rect 3437 624 3443 756
rect 3453 744 3459 756
rect 3453 604 3459 616
rect 3437 244 3443 576
rect 3421 223 3427 236
rect 3421 217 3436 223
rect 3453 184 3459 496
rect 3469 344 3475 656
rect 3517 644 3523 676
rect 3508 617 3516 623
rect 3485 484 3491 616
rect 3533 484 3539 1156
rect 3549 1084 3555 2276
rect 3565 1904 3571 2656
rect 3581 2624 3587 2996
rect 3581 2384 3587 2616
rect 3597 2284 3603 3436
rect 3677 3324 3683 3376
rect 3629 3084 3635 3116
rect 3677 3024 3683 3056
rect 3629 2924 3635 2936
rect 3709 2924 3715 3456
rect 3613 2524 3619 2596
rect 3645 2584 3651 2716
rect 3613 2364 3619 2396
rect 3581 2104 3587 2256
rect 3581 1924 3587 1976
rect 3572 1897 3580 1903
rect 3565 1524 3571 1896
rect 3597 1884 3603 2276
rect 3581 1764 3587 1876
rect 3597 1744 3603 1876
rect 3613 1764 3619 2356
rect 3629 2204 3635 2516
rect 3661 2484 3667 2616
rect 3645 2224 3651 2256
rect 3661 2224 3667 2236
rect 3629 2044 3635 2176
rect 3645 2104 3651 2176
rect 3661 1904 3667 2116
rect 3629 1744 3635 1776
rect 3581 1584 3587 1736
rect 3661 1704 3667 1896
rect 3645 1684 3651 1696
rect 3645 1604 3651 1616
rect 3629 1524 3635 1536
rect 3565 1144 3571 1156
rect 3565 944 3571 996
rect 3549 884 3555 936
rect 3469 324 3475 336
rect 3549 304 3555 676
rect 3581 564 3587 1496
rect 3597 1244 3603 1356
rect 3613 1344 3619 1356
rect 3597 984 3603 1236
rect 3613 1057 3628 1063
rect 3613 964 3619 1057
rect 3629 1004 3635 1036
rect 3645 964 3651 1556
rect 3661 1484 3667 1696
rect 3661 1324 3667 1476
rect 3661 1104 3667 1316
rect 3661 1024 3667 1096
rect 3597 704 3603 936
rect 3645 904 3651 956
rect 3645 524 3651 736
rect 3613 284 3619 296
rect 3677 264 3683 2696
rect 3709 2584 3715 2596
rect 3700 2277 3708 2283
rect 3693 2124 3699 2156
rect 3725 2124 3731 3396
rect 3741 3324 3747 3396
rect 3805 3384 3811 3396
rect 3741 3124 3747 3256
rect 3773 3104 3779 3196
rect 3789 3144 3795 3156
rect 3741 2504 3747 2896
rect 3757 2644 3763 2696
rect 3741 2424 3747 2436
rect 3693 2004 3699 2096
rect 3693 1844 3699 1896
rect 3693 1144 3699 1756
rect 3709 1724 3715 2096
rect 3725 1964 3731 2116
rect 3741 2084 3747 2276
rect 3757 2164 3763 2496
rect 3773 2324 3779 2336
rect 3773 2224 3779 2276
rect 3789 2224 3795 2256
rect 3757 1964 3763 2116
rect 3732 1857 3747 1863
rect 3741 1784 3747 1796
rect 3725 1764 3731 1776
rect 3725 1724 3731 1756
rect 3709 1364 3715 1636
rect 3709 1224 3715 1316
rect 3693 1064 3699 1136
rect 3709 1124 3715 1156
rect 3725 1104 3731 1716
rect 3741 1204 3747 1756
rect 3725 1064 3731 1096
rect 3693 624 3699 1036
rect 3709 984 3715 1016
rect 3725 964 3731 1056
rect 3709 684 3715 936
rect 3741 724 3747 1196
rect 3757 904 3763 1956
rect 3757 724 3763 896
rect 3741 704 3747 716
rect 3693 584 3699 616
rect 3693 544 3699 556
rect 3709 484 3715 556
rect 3492 257 3500 263
rect 3421 143 3427 176
rect 3421 137 3436 143
rect 3469 124 3475 196
rect 3533 144 3539 176
rect 3581 164 3587 176
rect 3549 144 3555 156
rect 3588 137 3596 143
rect 3620 137 3628 143
rect 3380 117 3388 123
rect 3405 24 3411 116
rect 3661 104 3667 216
rect 3693 164 3699 216
rect 3757 164 3763 696
rect 3773 124 3779 1916
rect 3789 1324 3795 2196
rect 3805 1724 3811 3296
rect 3821 3064 3827 3476
rect 3933 3444 3939 3476
rect 3949 3464 3955 3476
rect 3901 3424 3907 3436
rect 4045 3384 4051 3476
rect 4061 3444 4067 3476
rect 4061 3364 4067 3376
rect 4020 3357 4028 3363
rect 3860 2917 3868 2923
rect 3837 2664 3843 2916
rect 3869 2704 3875 2836
rect 3853 2683 3859 2696
rect 3853 2677 3875 2683
rect 3821 2304 3827 2516
rect 3821 2224 3827 2256
rect 3821 2124 3827 2176
rect 3821 1724 3827 2056
rect 3837 1944 3843 2656
rect 3869 2644 3875 2677
rect 3860 2597 3875 2603
rect 3869 2584 3875 2597
rect 3885 2524 3891 2796
rect 3853 2404 3859 2516
rect 3901 2504 3907 2976
rect 3949 2964 3955 3096
rect 3933 2724 3939 2956
rect 3917 2604 3923 2616
rect 3885 2484 3891 2496
rect 3805 1604 3811 1616
rect 3789 1304 3795 1316
rect 3805 1304 3811 1476
rect 3821 1264 3827 1376
rect 3853 1364 3859 2396
rect 3869 2184 3875 2216
rect 3869 2064 3875 2076
rect 3869 1844 3875 2036
rect 3885 1884 3891 2476
rect 3917 2344 3923 2556
rect 3933 2524 3939 2696
rect 3869 1484 3875 1796
rect 3885 1744 3891 1856
rect 3853 1344 3859 1356
rect 3837 1324 3843 1336
rect 3901 1324 3907 2296
rect 3917 2224 3923 2336
rect 3933 2144 3939 2216
rect 3917 1984 3923 2016
rect 3917 1744 3923 1956
rect 3805 1243 3811 1256
rect 3837 1243 3843 1296
rect 3805 1237 3843 1243
rect 3789 1164 3795 1196
rect 3789 1064 3795 1156
rect 3837 1144 3843 1196
rect 3805 1064 3811 1136
rect 3853 1044 3859 1196
rect 3901 1104 3907 1316
rect 3917 1244 3923 1736
rect 3917 1204 3923 1216
rect 3901 1084 3907 1096
rect 3917 1064 3923 1096
rect 3805 904 3811 976
rect 3789 884 3795 896
rect 3821 883 3827 1036
rect 3853 1004 3859 1016
rect 3837 904 3843 976
rect 3805 877 3827 883
rect 3805 584 3811 877
rect 3869 864 3875 1036
rect 3885 884 3891 1036
rect 3933 984 3939 2136
rect 3949 2104 3955 2956
rect 3965 2264 3971 3356
rect 3997 3304 4003 3356
rect 4052 3297 4060 3303
rect 4020 3137 4028 3143
rect 3981 2924 3987 3036
rect 3965 1924 3971 2256
rect 3981 2204 3987 2916
rect 3997 2904 4003 2916
rect 3997 2624 4003 2896
rect 4013 2884 4019 3016
rect 4029 2944 4035 3096
rect 4045 2924 4051 2936
rect 4045 2724 4051 2896
rect 4029 2624 4035 2636
rect 3997 2584 4003 2616
rect 4013 2584 4019 2596
rect 3997 2244 4003 2496
rect 3981 2144 3987 2156
rect 3949 1864 3955 1916
rect 3965 1804 3971 1856
rect 3981 1824 3987 2056
rect 3997 2004 4003 2236
rect 3997 1804 4003 1816
rect 3949 1764 3955 1796
rect 3972 1777 3980 1783
rect 3997 1744 4003 1776
rect 3981 1564 3987 1736
rect 3997 1524 4003 1536
rect 3917 924 3923 976
rect 3949 944 3955 1476
rect 3997 1464 4003 1496
rect 3949 884 3955 896
rect 3821 843 3827 856
rect 3821 837 3843 843
rect 3837 824 3843 837
rect 3789 504 3795 536
rect 3821 344 3827 776
rect 3949 764 3955 776
rect 3924 757 3932 763
rect 3869 724 3875 756
rect 3837 684 3843 696
rect 3837 644 3843 676
rect 3853 544 3859 716
rect 3901 704 3907 756
rect 3949 624 3955 696
rect 3901 617 3916 623
rect 3965 564 3971 1376
rect 4013 1324 4019 2376
rect 4029 2164 4035 2596
rect 3981 1224 3987 1316
rect 3981 1124 3987 1156
rect 3981 964 3987 976
rect 3997 744 4003 756
rect 3981 704 3987 736
rect 3997 724 4003 736
rect 4013 724 4019 1316
rect 4029 964 4035 2156
rect 4045 2004 4051 2716
rect 4061 2084 4067 3056
rect 4077 2624 4083 3476
rect 4093 3444 4099 3497
rect 4317 3484 4323 3496
rect 4324 3477 4332 3483
rect 4381 3464 4387 3476
rect 4196 3437 4204 3443
rect 4093 3424 4099 3436
rect 4164 3397 4172 3403
rect 4093 3384 4099 3396
rect 4093 2644 4099 3356
rect 4109 2544 4115 3396
rect 4173 3304 4179 3356
rect 4189 3324 4195 3336
rect 4141 2904 4147 2936
rect 4077 2504 4083 2516
rect 4093 2464 4099 2516
rect 4109 2464 4115 2516
rect 4077 2384 4083 2396
rect 4045 1764 4051 1976
rect 4077 1964 4083 2356
rect 4093 2264 4099 2456
rect 4125 2364 4131 2876
rect 4173 2844 4179 3016
rect 4141 2684 4147 2736
rect 4141 2624 4147 2636
rect 4157 2564 4163 2716
rect 4148 2557 4156 2563
rect 4141 2504 4147 2516
rect 4157 2324 4163 2496
rect 4093 2197 4099 2216
rect 4093 2104 4099 2116
rect 4109 1984 4115 2316
rect 4125 2304 4131 2316
rect 4125 2204 4131 2256
rect 4141 2244 4147 2316
rect 4125 2164 4131 2176
rect 4141 2004 4147 2156
rect 4157 2124 4163 2316
rect 4061 1764 4067 1956
rect 4077 1944 4083 1956
rect 4077 1884 4083 1916
rect 4061 1604 4067 1736
rect 4052 1457 4060 1463
rect 4045 1344 4051 1356
rect 4029 744 4035 896
rect 4045 824 4051 1296
rect 4061 924 4067 1416
rect 4045 784 4051 796
rect 4061 724 4067 896
rect 4077 724 4083 1876
rect 4093 1744 4099 1856
rect 4093 1684 4099 1696
rect 4045 704 4051 716
rect 4029 643 4035 696
rect 4029 637 4044 643
rect 4013 604 4019 616
rect 3837 364 3843 376
rect 3789 264 3795 316
rect 3805 304 3811 316
rect 3821 284 3827 296
rect 3853 244 3859 336
rect 3901 324 3907 516
rect 3949 324 3955 336
rect 3869 264 3875 296
rect 3885 284 3891 296
rect 3901 224 3907 236
rect 3789 144 3795 216
rect 3805 204 3811 216
rect 3949 144 3955 176
rect 3965 164 3971 556
rect 4029 504 4035 596
rect 4045 564 4051 616
rect 4013 464 4019 476
rect 3997 344 4003 356
rect 3981 124 3987 176
rect 3997 104 4003 216
rect 4061 164 4067 716
rect 4077 704 4083 716
rect 4077 584 4083 596
rect 4093 564 4099 1656
rect 4109 1524 4115 1836
rect 4125 1744 4131 1776
rect 4141 1744 4147 1756
rect 4125 1524 4131 1716
rect 4141 1524 4147 1596
rect 4109 1464 4115 1476
rect 4109 1404 4115 1416
rect 4125 1364 4131 1456
rect 4141 1344 4147 1496
rect 4132 1317 4147 1323
rect 4141 1304 4147 1317
rect 4109 824 4115 1236
rect 4109 644 4115 816
rect 4125 584 4131 1296
rect 4141 1224 4147 1276
rect 4141 1044 4147 1176
rect 4141 704 4147 756
rect 4157 724 4163 2116
rect 4173 744 4179 2676
rect 4189 2264 4195 3316
rect 4205 2944 4211 3336
rect 4269 3284 4275 3436
rect 4429 3384 4435 3436
rect 4365 3324 4371 3336
rect 4189 2224 4195 2236
rect 4189 1804 4195 2096
rect 4205 1684 4211 2936
rect 4221 2684 4227 2936
rect 4269 2924 4275 3276
rect 4333 2944 4339 3316
rect 4349 3144 4355 3156
rect 4445 3124 4451 3516
rect 4461 3424 4467 3436
rect 4525 3344 4531 3376
rect 4557 3104 4563 3556
rect 4829 3497 4844 3503
rect 4653 3477 4723 3483
rect 4589 3457 4627 3463
rect 4589 3444 4595 3457
rect 4621 3444 4627 3457
rect 4653 3444 4659 3477
rect 4717 3464 4723 3477
rect 4829 3464 4835 3497
rect 4893 3484 4899 3596
rect 4349 2924 4355 2956
rect 4221 1744 4227 2676
rect 4237 2384 4243 2836
rect 4301 2824 4307 2896
rect 4285 2684 4291 2716
rect 4301 2664 4307 2676
rect 4317 2643 4323 2836
rect 4333 2664 4339 2676
rect 4285 2637 4323 2643
rect 4285 2624 4291 2637
rect 4253 2304 4259 2536
rect 4237 2284 4243 2296
rect 4269 2244 4275 2516
rect 4285 2304 4291 2516
rect 4349 2444 4355 2916
rect 4365 2744 4371 2916
rect 4461 2904 4467 2976
rect 4509 2924 4515 2956
rect 4365 2684 4371 2716
rect 4397 2664 4403 2756
rect 4372 2577 4380 2583
rect 4413 2564 4419 2796
rect 4429 2624 4435 2796
rect 4500 2757 4515 2763
rect 4509 2744 4515 2757
rect 4525 2724 4531 3096
rect 4564 3037 4572 3043
rect 4573 2984 4579 2996
rect 4468 2677 4476 2683
rect 4445 2664 4451 2676
rect 4509 2664 4515 2676
rect 4445 2624 4451 2636
rect 4253 2164 4259 2176
rect 4221 1684 4227 1716
rect 4189 1504 4195 1536
rect 4205 1464 4211 1676
rect 4221 1624 4227 1636
rect 4189 944 4195 1456
rect 4189 924 4195 936
rect 4189 844 4195 876
rect 4141 644 4147 676
rect 4157 664 4163 716
rect 4148 617 4156 623
rect 4173 604 4179 616
rect 4189 604 4195 836
rect 4109 543 4115 556
rect 4093 537 4115 543
rect 4093 504 4099 537
rect 4125 504 4131 576
rect 4205 564 4211 1456
rect 4221 1224 4227 1476
rect 4221 1084 4227 1096
rect 4237 1044 4243 2156
rect 4253 1944 4259 1956
rect 4253 1464 4259 1876
rect 4269 1864 4275 2236
rect 4285 1904 4291 2296
rect 4333 2264 4339 2416
rect 4301 1964 4307 1976
rect 4269 1524 4275 1856
rect 4269 1484 4275 1496
rect 4269 1444 4275 1456
rect 4253 1224 4259 1416
rect 4269 1184 4275 1416
rect 4285 1384 4291 1856
rect 4301 1464 4307 1936
rect 4317 1904 4323 2256
rect 4317 1884 4323 1896
rect 4317 1844 4323 1856
rect 4333 1764 4339 2156
rect 4349 2144 4355 2156
rect 4365 2024 4371 2416
rect 4413 2124 4419 2276
rect 4445 2143 4451 2596
rect 4429 2137 4451 2143
rect 4349 1844 4355 1936
rect 4365 1864 4371 1896
rect 4317 1684 4323 1716
rect 4333 1464 4339 1756
rect 4349 1743 4355 1796
rect 4349 1737 4371 1743
rect 4365 1724 4371 1737
rect 4381 1704 4387 2056
rect 4285 1364 4291 1376
rect 4301 1364 4307 1456
rect 4260 1097 4268 1103
rect 4285 1064 4291 1156
rect 4317 1104 4323 1436
rect 4333 1324 4339 1396
rect 4333 1244 4339 1296
rect 4253 1004 4259 1036
rect 4301 844 4307 996
rect 4221 744 4227 796
rect 4221 604 4227 616
rect 4253 604 4259 776
rect 4317 724 4323 1096
rect 4333 904 4339 976
rect 4189 544 4195 556
rect 4077 324 4083 416
rect 4173 384 4179 396
rect 4244 337 4252 343
rect 4116 317 4124 323
rect 4269 304 4275 696
rect 4285 344 4291 536
rect 4333 384 4339 596
rect 4349 584 4355 1696
rect 4365 1204 4371 1636
rect 4381 1584 4387 1596
rect 4381 1364 4387 1576
rect 4397 1504 4403 2076
rect 4413 1904 4419 2116
rect 4429 1964 4435 2137
rect 4413 1564 4419 1836
rect 4461 1784 4467 2476
rect 4477 2224 4483 2516
rect 4493 2504 4499 2576
rect 4541 2524 4547 2556
rect 4509 2504 4515 2516
rect 4493 2204 4499 2476
rect 4477 2144 4483 2196
rect 4477 2124 4483 2136
rect 4477 2044 4483 2076
rect 4493 2004 4499 2116
rect 4509 2104 4515 2216
rect 4493 1883 4499 1996
rect 4477 1877 4499 1883
rect 4397 1324 4403 1496
rect 4413 1464 4419 1536
rect 4461 1384 4467 1776
rect 4477 1544 4483 1877
rect 4445 1364 4451 1376
rect 4413 1324 4419 1356
rect 4477 1324 4483 1356
rect 4445 1284 4451 1316
rect 4429 1264 4435 1276
rect 4365 1104 4371 1196
rect 4413 1104 4419 1116
rect 4381 544 4387 956
rect 4413 924 4419 936
rect 4413 704 4419 716
rect 4413 544 4419 696
rect 4445 664 4451 1156
rect 4493 984 4499 1696
rect 4525 1644 4531 2516
rect 4557 2484 4563 2936
rect 4573 2604 4579 2636
rect 4548 2277 4556 2283
rect 4548 2117 4556 2123
rect 4557 2084 4563 2116
rect 4509 1364 4515 1416
rect 4525 1364 4531 1416
rect 4493 964 4499 976
rect 4509 944 4515 1316
rect 4525 1224 4531 1236
rect 4525 1084 4531 1136
rect 4525 924 4531 936
rect 4493 684 4499 736
rect 4509 704 4515 736
rect 4541 664 4547 1696
rect 4557 1384 4563 2016
rect 4573 1864 4579 2596
rect 4589 1924 4595 3236
rect 4605 3084 4611 3096
rect 4605 2564 4611 3036
rect 4621 2724 4627 3236
rect 4637 2704 4643 3096
rect 4669 3064 4675 3436
rect 4685 3144 4691 3456
rect 4829 3444 4835 3456
rect 4941 3444 4947 3456
rect 4685 3084 4691 3136
rect 4660 3037 4668 3043
rect 4701 2944 4707 3436
rect 4717 3084 4723 3276
rect 4605 2184 4611 2516
rect 4637 2204 4643 2316
rect 4653 2284 4659 2796
rect 4644 2117 4652 2123
rect 4605 2104 4611 2116
rect 4669 2104 4675 2816
rect 4685 2704 4691 2716
rect 4669 2084 4675 2096
rect 4685 1864 4691 2696
rect 4605 1744 4611 1796
rect 4637 1604 4643 1856
rect 4653 1744 4659 1776
rect 4685 1564 4691 1856
rect 4701 1724 4707 2936
rect 4717 2184 4723 3016
rect 4733 2964 4739 3196
rect 4749 3124 4755 3136
rect 4765 2944 4771 3116
rect 4717 1664 4723 2176
rect 4701 1564 4707 1596
rect 4573 1364 4579 1396
rect 4653 1384 4659 1496
rect 4589 1304 4595 1376
rect 4637 1324 4643 1376
rect 4557 684 4563 1096
rect 4541 644 4547 656
rect 4493 504 4499 596
rect 4532 557 4540 563
rect 4205 204 4211 216
rect 4301 204 4307 216
rect 4413 204 4419 216
rect 4324 197 4332 203
rect 4093 184 4099 196
rect 4045 137 4083 143
rect 4045 123 4051 137
rect 4036 117 4051 123
rect 4061 104 4067 116
rect 4077 104 4083 137
rect 4109 124 4115 196
rect 4157 163 4163 196
rect 4189 183 4195 196
rect 4429 184 4435 476
rect 4557 304 4563 676
rect 4573 564 4579 1076
rect 4589 884 4595 996
rect 4605 684 4611 936
rect 4628 737 4636 743
rect 4605 524 4611 536
rect 4621 284 4627 696
rect 4637 504 4643 576
rect 4653 544 4659 1336
rect 4669 1304 4675 1416
rect 4644 277 4652 283
rect 4669 184 4675 1116
rect 4685 1064 4691 1496
rect 4685 724 4691 1056
rect 4701 824 4707 1556
rect 4717 1044 4723 1316
rect 4733 1024 4739 2376
rect 4749 1324 4755 2916
rect 4772 2517 4780 2523
rect 4765 2264 4771 2276
rect 4781 2244 4787 2496
rect 4765 1784 4771 2016
rect 4765 1604 4771 1756
rect 4765 1384 4771 1596
rect 4756 1317 4764 1323
rect 4749 1004 4755 1056
rect 4733 984 4739 996
rect 4685 544 4691 556
rect 4717 324 4723 976
rect 4733 744 4739 956
rect 4749 424 4755 836
rect 4765 304 4771 1016
rect 4781 704 4787 2116
rect 4797 1844 4803 2696
rect 4813 2024 4819 3136
rect 4829 2737 4835 2756
rect 4829 2124 4835 2716
rect 4845 2704 4851 3236
rect 4861 3124 4867 3336
rect 4893 3024 4899 3116
rect 4893 2864 4899 2996
rect 4868 2697 4876 2703
rect 4797 1704 4803 1816
rect 4797 1124 4803 1676
rect 4829 1664 4835 1696
rect 4845 1684 4851 2696
rect 4893 2684 4899 2736
rect 4877 2204 4883 2336
rect 4893 2324 4899 2596
rect 4877 1984 4883 2176
rect 4909 1964 4915 2956
rect 4925 2544 4931 3436
rect 4941 3264 4947 3436
rect 4973 3344 4979 3516
rect 4989 3364 4995 3556
rect 5044 3477 5052 3483
rect 5053 3364 5059 3376
rect 4861 1904 4867 1956
rect 4877 1844 4883 1876
rect 4861 1824 4867 1836
rect 4797 1104 4803 1116
rect 4797 624 4803 656
rect 4813 464 4819 1596
rect 4845 1544 4851 1576
rect 4829 1384 4835 1396
rect 4845 1364 4851 1516
rect 4829 1264 4835 1276
rect 4845 1064 4851 1076
rect 4829 644 4835 1056
rect 4845 764 4851 876
rect 4788 277 4796 283
rect 4845 224 4851 296
rect 4772 217 4780 223
rect 4189 177 4211 183
rect 4157 157 4195 163
rect 4189 144 4195 157
rect 4157 124 4163 136
rect 4205 124 4211 177
rect 4525 164 4531 176
rect 4541 124 4547 136
rect 4781 124 4787 176
rect 4797 164 4803 216
rect 4861 204 4867 1796
rect 4877 1544 4883 1756
rect 4877 1324 4883 1416
rect 4893 1043 4899 1896
rect 4909 1124 4915 1736
rect 4925 1484 4931 2496
rect 4941 2124 4947 2676
rect 4957 2644 4963 2856
rect 4973 2664 4979 3236
rect 5005 3124 5011 3316
rect 5101 3304 5107 3396
rect 5117 3364 5123 3376
rect 5005 2844 5011 2896
rect 4957 2524 4963 2536
rect 4973 2504 4979 2576
rect 4989 2524 4995 2656
rect 4957 2484 4963 2496
rect 5005 2304 5011 2836
rect 4980 2277 4988 2283
rect 4941 1524 4947 2116
rect 4893 1037 4915 1043
rect 4877 544 4883 936
rect 4877 284 4883 536
rect 4893 264 4899 896
rect 4820 157 4828 163
rect 4845 144 4851 196
rect 4909 124 4915 1037
rect 4925 944 4931 1456
rect 4941 1104 4947 1516
rect 4925 664 4931 936
rect 4941 784 4947 956
rect 4925 584 4931 596
rect 4957 524 4963 1956
rect 4973 1744 4979 2116
rect 5005 2104 5011 2296
rect 5037 2284 5043 3236
rect 5053 2784 5059 3056
rect 5053 2644 5059 2656
rect 5053 2484 5059 2496
rect 5005 1724 5011 1736
rect 5021 1564 5027 2156
rect 5037 1984 5043 2196
rect 5053 2164 5059 2296
rect 5053 1864 5059 2116
rect 5037 1524 5043 1676
rect 5069 1504 5075 2976
rect 5085 2744 5091 2956
rect 5085 2704 5091 2716
rect 5101 2663 5107 2936
rect 5117 2884 5123 3236
rect 5117 2664 5123 2736
rect 5085 2657 5107 2663
rect 5085 1804 5091 2657
rect 5101 2064 5107 2596
rect 5117 2144 5123 2636
rect 5101 2004 5107 2036
rect 5085 1744 5091 1776
rect 5085 1504 5091 1536
rect 5101 1524 5107 1976
rect 5117 1904 5123 2116
rect 4980 1457 4988 1463
rect 5005 1444 5011 1456
rect 4973 964 4979 1436
rect 4996 1337 5004 1343
rect 4989 1064 4995 1236
rect 5005 1064 5011 1336
rect 5069 1104 5075 1116
rect 4989 304 4995 716
rect 5005 664 5011 1036
rect 5037 984 5043 996
rect 5021 884 5027 956
rect 5053 924 5059 1016
rect 5053 824 5059 916
rect 5085 844 5091 1476
rect 5101 1344 5107 1496
rect 5101 1184 5107 1316
rect 5101 964 5107 1156
rect 5117 1004 5123 1876
rect 5037 724 5043 776
rect 5005 204 5011 636
rect 4989 144 4995 156
rect 5053 124 5059 576
rect 5085 503 5091 696
rect 5101 684 5107 696
rect 5133 644 5139 3476
rect 5165 3444 5171 3456
rect 5149 2884 5155 2896
rect 5149 2304 5155 2856
rect 5165 2584 5171 2756
rect 5149 1484 5155 2276
rect 5149 1344 5155 1356
rect 5149 844 5155 1296
rect 5165 964 5171 1956
rect 5181 984 5187 2796
rect 5197 1064 5203 1336
rect 5133 584 5139 596
rect 5108 537 5116 543
rect 5149 524 5155 816
rect 5172 777 5180 783
rect 5197 764 5203 1036
rect 5085 497 5100 503
rect 5165 424 5171 736
rect 5124 277 5132 283
rect 5076 257 5084 263
rect 5069 164 5075 176
rect 5156 157 5164 163
rect 5213 84 5219 2816
rect 1988 17 1996 23
<< m5contact >>
rect 476 3536 484 3544
rect 92 3156 100 3164
rect 156 3376 164 3384
rect 108 2696 116 2704
rect 76 1376 84 1384
rect 124 1356 132 1364
rect 172 3096 180 3104
rect 284 3276 292 3284
rect 316 3096 324 3104
rect 236 3056 244 3064
rect 204 2676 212 2684
rect 172 2656 180 2664
rect 172 2256 180 2264
rect 172 2156 180 2164
rect 220 2256 228 2264
rect 204 2176 212 2184
rect 172 1896 180 1904
rect 156 1736 164 1744
rect 300 2916 308 2924
rect 284 2696 292 2704
rect 252 2656 260 2664
rect 284 2216 292 2224
rect 268 2196 276 2204
rect 252 2176 260 2184
rect 236 1496 244 1504
rect 156 1376 164 1384
rect 204 1116 212 1124
rect 220 1016 228 1024
rect 124 956 132 964
rect 108 936 116 944
rect 76 716 84 724
rect 188 636 196 644
rect 124 576 132 584
rect 172 536 180 544
rect 252 976 260 984
rect 972 3496 980 3504
rect 476 3476 484 3484
rect 796 3476 804 3484
rect 956 3476 964 3484
rect 412 3456 420 3464
rect 364 3336 372 3344
rect 364 3296 372 3304
rect 380 2676 388 2684
rect 364 2596 372 2604
rect 348 2436 356 2444
rect 332 2296 340 2304
rect 332 2256 340 2264
rect 332 2136 340 2144
rect 300 1856 308 1864
rect 316 1756 324 1764
rect 300 1456 308 1464
rect 300 976 308 984
rect 300 936 308 944
rect 284 736 292 744
rect 252 316 260 324
rect 124 156 132 164
rect 316 656 324 664
rect 556 3456 564 3464
rect 588 3376 596 3384
rect 428 2896 436 2904
rect 412 2716 420 2724
rect 428 2656 436 2664
rect 412 2636 420 2644
rect 460 3156 468 3164
rect 492 3276 500 3284
rect 460 2696 468 2704
rect 444 2536 452 2544
rect 444 2496 452 2504
rect 460 2336 468 2344
rect 524 3096 532 3104
rect 540 2916 548 2924
rect 492 2736 500 2744
rect 508 2656 516 2664
rect 508 2296 516 2304
rect 492 2276 500 2284
rect 844 3456 852 3464
rect 700 3116 708 3124
rect 604 2896 612 2904
rect 588 2696 596 2704
rect 540 2636 548 2644
rect 540 2556 548 2564
rect 556 2536 564 2544
rect 476 2236 484 2244
rect 428 2136 436 2144
rect 476 2136 484 2144
rect 380 1556 388 1564
rect 364 1436 372 1444
rect 380 1376 388 1384
rect 348 916 356 924
rect 460 1776 468 1784
rect 508 1756 516 1764
rect 476 1656 484 1664
rect 412 1116 420 1124
rect 428 936 436 944
rect 380 316 388 324
rect 412 356 420 364
rect 476 1476 484 1484
rect 444 776 452 784
rect 492 1376 500 1384
rect 492 976 500 984
rect 572 2316 580 2324
rect 572 2296 580 2304
rect 572 1596 580 1604
rect 556 1456 564 1464
rect 556 1396 564 1404
rect 604 2336 612 2344
rect 604 2116 612 2124
rect 604 1536 612 1544
rect 524 916 532 924
rect 524 716 532 724
rect 556 716 564 724
rect 444 596 452 604
rect 428 296 436 304
rect 396 276 404 284
rect 476 276 484 284
rect 348 156 356 164
rect 460 156 468 164
rect 284 136 292 144
rect 444 136 452 144
rect 540 596 548 604
rect 508 516 516 524
rect 588 1316 596 1324
rect 668 2236 676 2244
rect 668 2216 676 2224
rect 668 2116 676 2124
rect 668 1916 676 1924
rect 732 3376 740 3384
rect 764 3316 772 3324
rect 732 3276 740 3284
rect 764 3216 772 3224
rect 716 2876 724 2884
rect 700 2756 708 2764
rect 700 2516 708 2524
rect 764 3096 772 3104
rect 764 3076 772 3084
rect 940 3356 948 3364
rect 828 3296 836 3304
rect 796 2996 804 3004
rect 748 2696 756 2704
rect 748 2656 756 2664
rect 748 2616 756 2624
rect 732 2296 740 2304
rect 700 2236 708 2244
rect 764 2576 772 2584
rect 716 2176 724 2184
rect 748 2176 756 2184
rect 668 1416 676 1424
rect 668 1336 676 1344
rect 700 1316 708 1324
rect 652 1096 660 1104
rect 652 676 660 684
rect 636 476 644 484
rect 620 276 628 284
rect 748 1956 756 1964
rect 812 2856 820 2864
rect 812 2776 820 2784
rect 764 1236 772 1244
rect 764 936 772 944
rect 764 856 772 864
rect 764 756 772 764
rect 828 2556 836 2564
rect 828 2516 836 2524
rect 828 2476 836 2484
rect 892 3316 900 3324
rect 860 2676 868 2684
rect 892 3136 900 3144
rect 876 2556 884 2564
rect 876 2436 884 2444
rect 860 2276 868 2284
rect 844 2256 852 2264
rect 844 2056 852 2064
rect 828 2036 836 2044
rect 844 2016 852 2024
rect 844 1976 852 1984
rect 844 1856 852 1864
rect 844 1796 852 1804
rect 812 1176 820 1184
rect 780 736 788 744
rect 780 596 788 604
rect 748 556 756 564
rect 764 556 772 564
rect 780 516 788 524
rect 748 316 756 324
rect 940 3136 948 3144
rect 940 2996 948 3004
rect 940 2956 948 2964
rect 972 2936 980 2944
rect 972 2916 980 2924
rect 972 2656 980 2664
rect 972 2636 980 2644
rect 924 2356 932 2364
rect 924 2276 932 2284
rect 924 1956 932 1964
rect 924 1896 932 1904
rect 908 1876 916 1884
rect 924 1776 932 1784
rect 924 1756 932 1764
rect 860 1476 868 1484
rect 972 2416 980 2424
rect 1388 3516 1396 3524
rect 1820 3496 1828 3504
rect 1036 3456 1044 3464
rect 1084 3436 1092 3444
rect 1004 3356 1012 3364
rect 1020 3356 1028 3364
rect 1036 3336 1044 3344
rect 1116 3336 1124 3344
rect 1148 3336 1156 3344
rect 1004 3076 1012 3084
rect 1004 3016 1012 3024
rect 1036 3096 1044 3104
rect 1084 3036 1092 3044
rect 1036 2916 1044 2924
rect 972 2296 980 2304
rect 972 1976 980 1984
rect 956 1856 964 1864
rect 860 1296 868 1304
rect 908 1036 916 1044
rect 764 256 772 264
rect 732 236 740 244
rect 700 216 708 224
rect 748 176 756 184
rect 700 156 708 164
rect 892 556 900 564
rect 892 456 900 464
rect 908 336 916 344
rect 860 316 868 324
rect 876 316 884 324
rect 988 1956 996 1964
rect 988 1476 996 1484
rect 988 1456 996 1464
rect 1068 2896 1076 2904
rect 1132 3096 1140 3104
rect 1052 2236 1060 2244
rect 1020 1896 1028 1904
rect 1052 1916 1060 1924
rect 1036 1796 1044 1804
rect 1036 1556 1044 1564
rect 1004 1276 1012 1284
rect 988 1076 996 1084
rect 988 1056 996 1064
rect 956 936 964 944
rect 940 596 948 604
rect 940 556 948 564
rect 940 336 948 344
rect 972 216 980 224
rect 908 156 916 164
rect 716 136 724 144
rect 844 136 852 144
rect 876 136 884 144
rect 1004 636 1012 644
rect 1004 616 1012 624
rect 1100 2276 1108 2284
rect 1132 2976 1140 2984
rect 1132 2916 1140 2924
rect 1132 2696 1140 2704
rect 1132 2436 1140 2444
rect 1132 2376 1140 2384
rect 1132 2336 1140 2344
rect 1196 3336 1204 3344
rect 1196 3096 1204 3104
rect 1132 2096 1140 2104
rect 1100 1916 1108 1924
rect 1068 1276 1076 1284
rect 1052 656 1060 664
rect 1116 1836 1124 1844
rect 1116 1776 1124 1784
rect 1116 1716 1124 1724
rect 1196 2716 1204 2724
rect 1164 1996 1172 2004
rect 1164 1916 1172 1924
rect 1164 1736 1172 1744
rect 1084 636 1092 644
rect 1100 616 1108 624
rect 1100 596 1108 604
rect 1084 556 1092 564
rect 1100 556 1108 564
rect 1164 1456 1172 1464
rect 1132 1256 1140 1264
rect 1148 1256 1156 1264
rect 1148 1236 1156 1244
rect 1132 1216 1140 1224
rect 1132 1056 1140 1064
rect 1132 1036 1140 1044
rect 1164 1056 1172 1064
rect 1148 936 1156 944
rect 1164 936 1172 944
rect 1164 836 1172 844
rect 1164 796 1172 804
rect 1148 696 1156 704
rect 1148 576 1156 584
rect 1100 336 1108 344
rect 1132 196 1140 204
rect 1164 176 1172 184
rect 1068 136 1076 144
rect 716 116 724 124
rect 940 116 948 124
rect 956 116 964 124
rect 524 96 532 104
rect 1244 3476 1252 3484
rect 1212 2236 1220 2244
rect 1260 3336 1268 3344
rect 1308 3356 1316 3364
rect 1292 3256 1300 3264
rect 1308 3156 1316 3164
rect 1308 3116 1316 3124
rect 1244 2876 1252 2884
rect 1244 2656 1252 2664
rect 1260 2176 1268 2184
rect 1260 2116 1268 2124
rect 1308 3036 1316 3044
rect 1292 2716 1300 2724
rect 1292 2596 1300 2604
rect 1308 2556 1316 2564
rect 1308 2516 1316 2524
rect 1260 2016 1268 2024
rect 1260 1816 1268 1824
rect 1228 1696 1236 1704
rect 1228 1576 1236 1584
rect 1276 1796 1284 1804
rect 1276 1716 1284 1724
rect 1308 2016 1316 2024
rect 1308 1916 1316 1924
rect 1340 3356 1348 3364
rect 1356 3156 1364 3164
rect 1356 3116 1364 3124
rect 1340 2936 1348 2944
rect 1340 2916 1348 2924
rect 1340 2596 1348 2604
rect 1340 2536 1348 2544
rect 1340 2456 1348 2464
rect 1340 2196 1348 2204
rect 1340 2096 1348 2104
rect 1340 1896 1348 1904
rect 1292 1696 1300 1704
rect 1276 1656 1284 1664
rect 1212 1156 1220 1164
rect 1244 1396 1252 1404
rect 1244 1316 1252 1324
rect 1212 896 1220 904
rect 1228 896 1236 904
rect 1196 616 1204 624
rect 1212 576 1220 584
rect 1196 176 1204 184
rect 1244 336 1252 344
rect 1308 1496 1316 1504
rect 1340 1376 1348 1384
rect 1340 1296 1348 1304
rect 1276 876 1284 884
rect 1308 876 1316 884
rect 1404 3116 1412 3124
rect 1372 2716 1380 2724
rect 1388 2576 1396 2584
rect 1644 3376 1652 3384
rect 1452 3336 1460 3344
rect 1484 3036 1492 3044
rect 1452 2936 1460 2944
rect 1436 2916 1444 2924
rect 1452 2896 1460 2904
rect 1452 2876 1460 2884
rect 1436 2576 1444 2584
rect 1388 2556 1396 2564
rect 1404 2556 1412 2564
rect 1388 2476 1396 2484
rect 1420 2316 1428 2324
rect 1420 2296 1428 2304
rect 1388 2216 1396 2224
rect 1388 2096 1396 2104
rect 1388 1916 1396 1924
rect 1372 1896 1380 1904
rect 1388 1856 1396 1864
rect 1404 1856 1412 1864
rect 1372 1796 1380 1804
rect 1388 1736 1396 1744
rect 1436 2276 1444 2284
rect 1436 1936 1444 1944
rect 1372 1196 1380 1204
rect 1420 1216 1428 1224
rect 1420 1136 1428 1144
rect 1388 876 1396 884
rect 1404 856 1412 864
rect 1356 816 1364 824
rect 1324 696 1332 704
rect 1324 636 1332 644
rect 1308 616 1316 624
rect 1324 536 1332 544
rect 1356 516 1364 524
rect 1372 416 1380 424
rect 1404 676 1412 684
rect 1404 576 1412 584
rect 1388 396 1396 404
rect 1404 376 1412 384
rect 1228 256 1236 264
rect 1244 256 1252 264
rect 1356 256 1364 264
rect 1468 2536 1476 2544
rect 1532 3036 1540 3044
rect 1516 2696 1524 2704
rect 1516 2676 1524 2684
rect 1468 2096 1476 2104
rect 1516 2496 1524 2504
rect 1532 2436 1540 2444
rect 1532 2336 1540 2344
rect 1532 2316 1540 2324
rect 1516 2276 1524 2284
rect 1532 2196 1540 2204
rect 1516 2176 1524 2184
rect 1516 1956 1524 1964
rect 1500 1856 1508 1864
rect 1676 3336 1684 3344
rect 1628 3056 1636 3064
rect 1692 3136 1700 3144
rect 1676 3116 1684 3124
rect 1596 2916 1604 2924
rect 1580 2896 1588 2904
rect 1628 2856 1636 2864
rect 1580 2816 1588 2824
rect 1564 2576 1572 2584
rect 1580 2576 1588 2584
rect 1564 2556 1572 2564
rect 1580 2476 1588 2484
rect 1564 2436 1572 2444
rect 1580 2436 1588 2444
rect 1580 2316 1588 2324
rect 1564 2176 1572 2184
rect 1564 2136 1572 2144
rect 1548 1856 1556 1864
rect 1500 1816 1508 1824
rect 1548 1816 1556 1824
rect 1516 1396 1524 1404
rect 1500 1356 1508 1364
rect 1484 1196 1492 1204
rect 1468 956 1476 964
rect 1468 916 1476 924
rect 1468 876 1476 884
rect 1452 496 1460 504
rect 1468 256 1476 264
rect 1244 216 1252 224
rect 1260 216 1268 224
rect 1356 176 1364 184
rect 1500 1016 1508 1024
rect 1516 716 1524 724
rect 1548 1676 1556 1684
rect 1532 676 1540 684
rect 1628 2756 1636 2764
rect 1628 2496 1636 2504
rect 1628 2456 1636 2464
rect 1628 2196 1636 2204
rect 1628 2156 1636 2164
rect 1612 2096 1620 2104
rect 1612 2056 1620 2064
rect 1628 2016 1636 2024
rect 1612 1936 1620 1944
rect 1628 1936 1636 1944
rect 1628 1896 1636 1904
rect 1724 3376 1732 3384
rect 1676 2456 1684 2464
rect 1708 2876 1716 2884
rect 1708 2636 1716 2644
rect 1708 2576 1716 2584
rect 1772 3096 1780 3104
rect 1772 3036 1780 3044
rect 1772 2936 1780 2944
rect 1820 2936 1828 2944
rect 2060 3516 2068 3524
rect 2156 3516 2164 3524
rect 2220 3516 2228 3524
rect 1916 3496 1924 3504
rect 1868 3336 1876 3344
rect 1868 3236 1876 3244
rect 1868 3216 1876 3224
rect 1868 3076 1876 3084
rect 1868 3036 1876 3044
rect 1804 2856 1812 2864
rect 1804 2696 1812 2704
rect 1708 2196 1716 2204
rect 1756 2256 1764 2264
rect 1708 2156 1716 2164
rect 1708 2116 1716 2124
rect 1660 2036 1668 2044
rect 1660 2016 1668 2024
rect 1596 1836 1604 1844
rect 1644 1836 1652 1844
rect 1596 1796 1604 1804
rect 1612 1656 1620 1664
rect 1580 1496 1588 1504
rect 1596 1496 1604 1504
rect 1644 1776 1652 1784
rect 1644 1736 1652 1744
rect 1644 1576 1652 1584
rect 1644 1556 1652 1564
rect 1580 1356 1588 1364
rect 1580 956 1588 964
rect 1612 1396 1620 1404
rect 1644 1396 1652 1404
rect 1628 1316 1636 1324
rect 1612 1196 1620 1204
rect 1564 696 1572 704
rect 1532 516 1540 524
rect 1644 1136 1652 1144
rect 1644 996 1652 1004
rect 1692 1896 1700 1904
rect 1676 1756 1684 1764
rect 1676 1516 1684 1524
rect 1676 1476 1684 1484
rect 1724 2016 1732 2024
rect 1708 1616 1716 1624
rect 1676 1056 1684 1064
rect 1676 1036 1684 1044
rect 1676 956 1684 964
rect 1676 856 1684 864
rect 1676 676 1684 684
rect 1596 536 1604 544
rect 1708 1116 1716 1124
rect 1644 596 1652 604
rect 1660 556 1668 564
rect 1660 456 1668 464
rect 1580 376 1588 384
rect 1628 256 1636 264
rect 1548 156 1556 164
rect 1628 156 1636 164
rect 1356 116 1364 124
rect 620 76 628 84
rect 956 76 964 84
rect 1660 376 1668 384
rect 1660 276 1668 284
rect 1660 156 1668 164
rect 1692 576 1700 584
rect 1692 276 1700 284
rect 1756 1936 1764 1944
rect 1740 1916 1748 1924
rect 1740 1856 1748 1864
rect 1756 1756 1764 1764
rect 1756 1736 1764 1744
rect 1756 1596 1764 1604
rect 1756 1476 1764 1484
rect 1740 1136 1748 1144
rect 1740 916 1748 924
rect 1740 836 1748 844
rect 1724 636 1732 644
rect 1788 2596 1796 2604
rect 1788 2576 1796 2584
rect 1804 2416 1812 2424
rect 1804 2376 1812 2384
rect 1788 2256 1796 2264
rect 1836 2656 1844 2664
rect 1868 2996 1876 3004
rect 1852 2636 1860 2644
rect 1836 2576 1844 2584
rect 1836 2536 1844 2544
rect 1788 1936 1796 1944
rect 1788 1716 1796 1724
rect 1820 2076 1828 2084
rect 1820 1876 1828 1884
rect 1820 1856 1828 1864
rect 1788 1556 1796 1564
rect 1788 1536 1796 1544
rect 1788 1516 1796 1524
rect 1900 2996 1908 3004
rect 1900 2896 1908 2904
rect 1900 2856 1908 2864
rect 1900 2696 1908 2704
rect 1852 2256 1860 2264
rect 1852 2216 1860 2224
rect 1900 2496 1908 2504
rect 2060 3496 2068 3504
rect 1932 2996 1940 3004
rect 1932 2876 1940 2884
rect 2028 3156 2036 3164
rect 2012 2936 2020 2944
rect 1964 2796 1972 2804
rect 1996 2736 2004 2744
rect 2012 2716 2020 2724
rect 1996 2676 2004 2684
rect 1948 2556 1956 2564
rect 1980 2536 1988 2544
rect 1964 2476 1972 2484
rect 1932 2356 1940 2364
rect 1916 2216 1924 2224
rect 1868 1816 1876 1824
rect 1884 1796 1892 1804
rect 1884 1756 1892 1764
rect 1884 1696 1892 1704
rect 1884 1456 1892 1464
rect 1852 1396 1860 1404
rect 2028 2676 2036 2684
rect 2044 2656 2052 2664
rect 2044 2636 2052 2644
rect 2044 2596 2052 2604
rect 2028 2536 2036 2544
rect 1980 2156 1988 2164
rect 1996 2156 2004 2164
rect 1948 1956 1956 1964
rect 1916 1616 1924 1624
rect 1964 1896 1972 1904
rect 1932 1436 1940 1444
rect 1836 1376 1844 1384
rect 1900 1376 1908 1384
rect 1868 1356 1876 1364
rect 1868 1336 1876 1344
rect 1884 1336 1892 1344
rect 1996 1876 2004 1884
rect 1996 1776 2004 1784
rect 1980 1736 1988 1744
rect 1996 1736 2004 1744
rect 2044 2196 2052 2204
rect 2044 2176 2052 2184
rect 2028 2016 2036 2024
rect 2076 3456 2084 3464
rect 2108 3356 2116 3364
rect 2172 3356 2180 3364
rect 2124 3336 2132 3344
rect 2188 3336 2196 3344
rect 2220 3436 2228 3444
rect 2524 3536 2532 3544
rect 2492 3456 2500 3464
rect 2732 3516 2740 3524
rect 2828 3516 2836 3524
rect 2844 3516 2852 3524
rect 2652 3496 2660 3504
rect 2684 3476 2692 3484
rect 2364 3436 2372 3444
rect 2508 3436 2516 3444
rect 2540 3436 2548 3444
rect 2316 3416 2324 3424
rect 2236 3356 2244 3364
rect 2108 3096 2116 3104
rect 2092 2996 2100 3004
rect 2092 2896 2100 2904
rect 2108 2876 2116 2884
rect 2076 2816 2084 2824
rect 2076 2776 2084 2784
rect 2092 2636 2100 2644
rect 2076 2456 2084 2464
rect 2060 2076 2068 2084
rect 2060 2016 2068 2024
rect 2044 1956 2052 1964
rect 1836 1316 1844 1324
rect 1964 1316 1972 1324
rect 1804 1276 1812 1284
rect 1884 1276 1892 1284
rect 1804 1076 1812 1084
rect 1788 916 1796 924
rect 1788 756 1796 764
rect 1804 676 1812 684
rect 1788 656 1796 664
rect 1724 536 1732 544
rect 1724 296 1732 304
rect 1740 296 1748 304
rect 1788 556 1796 564
rect 1868 1156 1876 1164
rect 1852 1036 1860 1044
rect 1884 936 1892 944
rect 1836 896 1844 904
rect 1884 896 1892 904
rect 1836 636 1844 644
rect 1836 376 1844 384
rect 1804 296 1812 304
rect 1868 436 1876 444
rect 1868 376 1876 384
rect 1916 1116 1924 1124
rect 1964 1236 1972 1244
rect 1948 1216 1956 1224
rect 1996 1696 2004 1704
rect 1996 1356 2004 1364
rect 1948 1196 1956 1204
rect 1980 1196 1988 1204
rect 1948 976 1956 984
rect 1916 816 1924 824
rect 1948 796 1956 804
rect 1932 776 1940 784
rect 1916 756 1924 764
rect 1916 636 1924 644
rect 1980 676 1988 684
rect 1980 656 1988 664
rect 2060 1896 2068 1904
rect 2028 1476 2036 1484
rect 2028 1456 2036 1464
rect 2028 1356 2036 1364
rect 2044 1256 2052 1264
rect 2060 1156 2068 1164
rect 1932 576 1940 584
rect 1948 536 1956 544
rect 1932 476 1940 484
rect 1948 256 1956 264
rect 1980 496 1988 504
rect 1980 456 1988 464
rect 2012 396 2020 404
rect 1996 376 2004 384
rect 1996 256 2004 264
rect 1884 236 1892 244
rect 1980 236 1988 244
rect 1772 216 1780 224
rect 1676 116 1684 124
rect 924 56 932 64
rect 1804 96 1812 104
rect 1868 96 1876 104
rect 1740 36 1748 44
rect 2044 1036 2052 1044
rect 2044 956 2052 964
rect 2156 2996 2164 3004
rect 2204 3076 2212 3084
rect 2220 3076 2228 3084
rect 2188 2856 2196 2864
rect 2124 2376 2132 2384
rect 2124 2316 2132 2324
rect 2188 2736 2196 2744
rect 2156 2656 2164 2664
rect 2172 2656 2180 2664
rect 2188 2616 2196 2624
rect 2172 2556 2180 2564
rect 2188 2556 2196 2564
rect 2188 2496 2196 2504
rect 2220 2856 2228 2864
rect 2332 3376 2340 3384
rect 2364 3336 2372 3344
rect 2236 2536 2244 2544
rect 2156 2376 2164 2384
rect 2140 2176 2148 2184
rect 2140 2036 2148 2044
rect 2108 1996 2116 2004
rect 2092 1896 2100 1904
rect 2108 1876 2116 1884
rect 2108 1816 2116 1824
rect 2108 1356 2116 1364
rect 2092 1316 2100 1324
rect 2076 1076 2084 1084
rect 2076 936 2084 944
rect 2076 656 2084 664
rect 2044 636 2052 644
rect 2076 556 2084 564
rect 2044 496 2052 504
rect 2076 336 2084 344
rect 2060 296 2068 304
rect 2108 1116 2116 1124
rect 2108 1096 2116 1104
rect 2140 1996 2148 2004
rect 2140 1776 2148 1784
rect 2140 1656 2148 1664
rect 2140 1616 2148 1624
rect 2140 1416 2148 1424
rect 2204 2316 2212 2324
rect 2188 2196 2196 2204
rect 2188 2116 2196 2124
rect 2204 2076 2212 2084
rect 2188 1996 2196 2004
rect 2172 1976 2180 1984
rect 2172 1936 2180 1944
rect 2188 1616 2196 1624
rect 2204 1596 2212 1604
rect 2172 1456 2180 1464
rect 2188 1456 2196 1464
rect 2188 1416 2196 1424
rect 2172 1356 2180 1364
rect 2140 1316 2148 1324
rect 2156 1296 2164 1304
rect 2140 1256 2148 1264
rect 2172 1256 2180 1264
rect 2172 1076 2180 1084
rect 2172 956 2180 964
rect 2140 916 2148 924
rect 2172 816 2180 824
rect 2156 796 2164 804
rect 2140 776 2148 784
rect 2140 636 2148 644
rect 2188 756 2196 764
rect 2172 736 2180 744
rect 2108 496 2116 504
rect 2124 456 2132 464
rect 2188 496 2196 504
rect 2300 2896 2308 2904
rect 2316 2896 2324 2904
rect 2316 2636 2324 2644
rect 2332 2596 2340 2604
rect 2284 2496 2292 2504
rect 2300 2496 2308 2504
rect 2268 2376 2276 2384
rect 2268 2196 2276 2204
rect 2300 2196 2308 2204
rect 2284 1996 2292 2004
rect 2268 1976 2276 1984
rect 2268 1776 2276 1784
rect 2284 1756 2292 1764
rect 2252 1676 2260 1684
rect 2236 1436 2244 1444
rect 2236 1136 2244 1144
rect 2236 916 2244 924
rect 2252 896 2260 904
rect 2236 796 2244 804
rect 2220 756 2228 764
rect 2236 656 2244 664
rect 2220 496 2228 504
rect 2188 316 2196 324
rect 2172 296 2180 304
rect 2060 236 2068 244
rect 2044 176 2052 184
rect 2108 176 2116 184
rect 2028 116 2036 124
rect 2204 116 2212 124
rect 2236 476 2244 484
rect 2236 456 2244 464
rect 2380 2936 2388 2944
rect 2380 2676 2388 2684
rect 2380 2656 2388 2664
rect 2316 1776 2324 1784
rect 2300 1636 2308 1644
rect 2284 1516 2292 1524
rect 2300 1516 2308 1524
rect 2300 1396 2308 1404
rect 2348 1836 2356 1844
rect 2332 1356 2340 1364
rect 2444 3336 2452 3344
rect 2412 3216 2420 3224
rect 2428 2936 2436 2944
rect 2428 2816 2436 2824
rect 2428 2716 2436 2724
rect 2428 2616 2436 2624
rect 2412 2596 2420 2604
rect 2396 2316 2404 2324
rect 2428 2456 2436 2464
rect 2428 2436 2436 2444
rect 2444 2436 2452 2444
rect 2396 2276 2404 2284
rect 2412 2216 2420 2224
rect 2396 2136 2404 2144
rect 2412 2036 2420 2044
rect 2412 1976 2420 1984
rect 2396 1956 2404 1964
rect 2380 1796 2388 1804
rect 2380 1776 2388 1784
rect 2364 1676 2372 1684
rect 2380 1636 2388 1644
rect 2396 1636 2404 1644
rect 2364 1516 2372 1524
rect 2300 1216 2308 1224
rect 2316 1196 2324 1204
rect 2284 1176 2292 1184
rect 2348 1136 2356 1144
rect 2284 1096 2292 1104
rect 2316 1036 2324 1044
rect 2300 956 2308 964
rect 2316 956 2324 964
rect 2268 616 2276 624
rect 2268 596 2276 604
rect 2316 596 2324 604
rect 2284 556 2292 564
rect 2316 556 2324 564
rect 2300 536 2308 544
rect 2396 1596 2404 1604
rect 2412 1596 2420 1604
rect 2412 1536 2420 1544
rect 2412 1436 2420 1444
rect 2396 1376 2404 1384
rect 2396 1316 2404 1324
rect 2396 1236 2404 1244
rect 2396 1216 2404 1224
rect 2396 1176 2404 1184
rect 2380 1036 2388 1044
rect 2396 956 2404 964
rect 2380 936 2388 944
rect 2476 3036 2484 3044
rect 2444 2036 2452 2044
rect 2444 1936 2452 1944
rect 2476 2276 2484 2284
rect 2476 2196 2484 2204
rect 2476 2116 2484 2124
rect 2460 1876 2468 1884
rect 2444 1836 2452 1844
rect 2460 1836 2468 1844
rect 2460 1676 2468 1684
rect 2444 1556 2452 1564
rect 2444 1516 2452 1524
rect 2444 1356 2452 1364
rect 2428 1276 2436 1284
rect 2428 1196 2436 1204
rect 2428 1176 2436 1184
rect 2444 1056 2452 1064
rect 2428 956 2436 964
rect 2428 916 2436 924
rect 2364 676 2372 684
rect 2380 656 2388 664
rect 2364 616 2372 624
rect 2332 476 2340 484
rect 2284 456 2292 464
rect 2316 456 2324 464
rect 2380 416 2388 424
rect 2380 376 2388 384
rect 2412 736 2420 744
rect 2428 736 2436 744
rect 2412 676 2420 684
rect 2428 676 2436 684
rect 2412 596 2420 604
rect 2428 596 2436 604
rect 2252 276 2260 284
rect 2380 276 2388 284
rect 2252 256 2260 264
rect 2396 256 2404 264
rect 2412 176 2420 184
rect 2012 96 2020 104
rect 2508 3376 2516 3384
rect 2540 3156 2548 3164
rect 2540 3036 2548 3044
rect 2524 3016 2532 3024
rect 2508 2936 2516 2944
rect 2540 2936 2548 2944
rect 2524 2636 2532 2644
rect 2556 2696 2564 2704
rect 2508 2536 2516 2544
rect 2524 2276 2532 2284
rect 2524 2196 2532 2204
rect 2508 1956 2516 1964
rect 2508 1556 2516 1564
rect 2492 1356 2500 1364
rect 2492 1256 2500 1264
rect 2492 1236 2500 1244
rect 2492 1196 2500 1204
rect 2556 2556 2564 2564
rect 2556 2476 2564 2484
rect 2556 2256 2564 2264
rect 2556 2216 2564 2224
rect 2732 3396 2740 3404
rect 2588 3376 2596 3384
rect 2604 3356 2612 3364
rect 2764 3356 2772 3364
rect 2716 3136 2724 3144
rect 2668 3036 2676 3044
rect 2588 2996 2596 3004
rect 2588 2716 2596 2724
rect 2620 2736 2628 2744
rect 2620 2696 2628 2704
rect 2588 2296 2596 2304
rect 2588 2256 2596 2264
rect 2588 2236 2596 2244
rect 2572 2136 2580 2144
rect 2572 2036 2580 2044
rect 2588 2016 2596 2024
rect 2572 1936 2580 1944
rect 2588 1896 2596 1904
rect 2572 1876 2580 1884
rect 2572 1856 2580 1864
rect 2668 2656 2676 2664
rect 2796 3416 2804 3424
rect 2812 3416 2820 3424
rect 2700 2916 2708 2924
rect 2700 2736 2708 2744
rect 2700 2636 2708 2644
rect 2700 2556 2708 2564
rect 2668 2536 2676 2544
rect 2684 2516 2692 2524
rect 2668 2456 2676 2464
rect 2700 2416 2708 2424
rect 2668 2336 2676 2344
rect 2684 2336 2692 2344
rect 2668 2276 2676 2284
rect 2684 2256 2692 2264
rect 2588 1716 2596 1724
rect 2588 1636 2596 1644
rect 2572 1456 2580 1464
rect 2572 1356 2580 1364
rect 2572 1296 2580 1304
rect 2492 956 2500 964
rect 2508 936 2516 944
rect 2492 796 2500 804
rect 2492 736 2500 744
rect 2476 616 2484 624
rect 2476 596 2484 604
rect 2476 576 2484 584
rect 2492 576 2500 584
rect 2460 536 2468 544
rect 2476 496 2484 504
rect 2460 396 2468 404
rect 2460 256 2468 264
rect 2492 396 2500 404
rect 2444 116 2452 124
rect 2556 1096 2564 1104
rect 2556 1076 2564 1084
rect 2556 916 2564 924
rect 2556 796 2564 804
rect 2620 1736 2628 1744
rect 2604 1336 2612 1344
rect 2604 1296 2612 1304
rect 2588 1076 2596 1084
rect 2588 996 2596 1004
rect 2588 756 2596 764
rect 2572 596 2580 604
rect 2556 576 2564 584
rect 2556 496 2564 504
rect 2684 2036 2692 2044
rect 2684 1996 2692 2004
rect 2700 1936 2708 1944
rect 2684 1916 2692 1924
rect 2700 1816 2708 1824
rect 2780 3056 2788 3064
rect 2796 3056 2804 3064
rect 2748 3016 2756 3024
rect 2764 2936 2772 2944
rect 2780 2876 2788 2884
rect 2748 2716 2756 2724
rect 2748 2556 2756 2564
rect 2748 2496 2756 2504
rect 2796 2656 2804 2664
rect 2796 2536 2804 2544
rect 2796 2476 2804 2484
rect 2748 2296 2756 2304
rect 2780 2276 2788 2284
rect 2748 2236 2756 2244
rect 2764 2216 2772 2224
rect 2748 2096 2756 2104
rect 2748 2036 2756 2044
rect 2748 1996 2756 2004
rect 2764 1956 2772 1964
rect 2748 1916 2756 1924
rect 2748 1896 2756 1904
rect 2764 1896 2772 1904
rect 2748 1856 2756 1864
rect 2716 1776 2724 1784
rect 2716 1756 2724 1764
rect 2668 1456 2676 1464
rect 2652 1416 2660 1424
rect 2668 1336 2676 1344
rect 2636 1216 2644 1224
rect 2636 1056 2644 1064
rect 2636 996 2644 1004
rect 2652 956 2660 964
rect 2652 736 2660 744
rect 2636 616 2644 624
rect 2652 476 2660 484
rect 2636 396 2644 404
rect 2636 316 2644 324
rect 2524 296 2532 304
rect 2540 296 2548 304
rect 2588 276 2596 284
rect 2508 256 2516 264
rect 2572 156 2580 164
rect 2508 136 2516 144
rect 2652 256 2660 264
rect 2748 1696 2756 1704
rect 2748 1656 2756 1664
rect 2764 1636 2772 1644
rect 2748 1576 2756 1584
rect 2748 1536 2756 1544
rect 2748 1416 2756 1424
rect 2732 1296 2740 1304
rect 2748 1236 2756 1244
rect 2732 1156 2740 1164
rect 2716 1116 2724 1124
rect 2764 1136 2772 1144
rect 2748 1056 2756 1064
rect 2732 996 2740 1004
rect 2732 956 2740 964
rect 2732 916 2740 924
rect 2748 876 2756 884
rect 2748 776 2756 784
rect 2732 756 2740 764
rect 2716 676 2724 684
rect 2844 3076 2852 3084
rect 2828 2936 2836 2944
rect 2828 2836 2836 2844
rect 2812 2276 2820 2284
rect 2812 2236 2820 2244
rect 2796 2036 2804 2044
rect 2796 1836 2804 1844
rect 2796 1756 2804 1764
rect 2796 1716 2804 1724
rect 2796 1596 2804 1604
rect 2860 2956 2868 2964
rect 2876 2916 2884 2924
rect 2876 2836 2884 2844
rect 3020 3396 3028 3404
rect 2972 3376 2980 3384
rect 2924 3296 2932 3304
rect 2988 3296 2996 3304
rect 2988 3116 2996 3124
rect 2924 3016 2932 3024
rect 2908 2996 2916 3004
rect 2972 2956 2980 2964
rect 2956 2936 2964 2944
rect 2924 2856 2932 2864
rect 2956 2816 2964 2824
rect 2956 2736 2964 2744
rect 2860 2496 2868 2504
rect 2876 2456 2884 2464
rect 2908 2616 2916 2624
rect 2924 2556 2932 2564
rect 2876 2416 2884 2424
rect 2892 2416 2900 2424
rect 2876 2316 2884 2324
rect 2844 2296 2852 2304
rect 2876 2296 2884 2304
rect 2844 2256 2852 2264
rect 2844 2236 2852 2244
rect 2844 2096 2852 2104
rect 2844 1956 2852 1964
rect 2844 1896 2852 1904
rect 2828 1476 2836 1484
rect 2796 1336 2804 1344
rect 2796 1216 2804 1224
rect 2828 1296 2836 1304
rect 2956 2356 2964 2364
rect 2940 2196 2948 2204
rect 2924 2156 2932 2164
rect 2940 2156 2948 2164
rect 2876 2116 2884 2124
rect 2908 2116 2916 2124
rect 2908 2096 2916 2104
rect 2876 1956 2884 1964
rect 2876 1856 2884 1864
rect 2860 1816 2868 1824
rect 2892 1776 2900 1784
rect 2860 1756 2868 1764
rect 2876 1756 2884 1764
rect 2908 1716 2916 1724
rect 2860 1696 2868 1704
rect 2876 1676 2884 1684
rect 2860 1636 2868 1644
rect 2908 1636 2916 1644
rect 2860 1416 2868 1424
rect 2892 1356 2900 1364
rect 2908 1356 2916 1364
rect 2940 1876 2948 1884
rect 2940 1836 2948 1844
rect 3052 3356 3060 3364
rect 3036 3136 3044 3144
rect 3020 2936 3028 2944
rect 3020 2736 3028 2744
rect 2988 2456 2996 2464
rect 2972 1916 2980 1924
rect 3036 2656 3044 2664
rect 3020 2516 3028 2524
rect 3020 2456 3028 2464
rect 3020 2316 3028 2324
rect 3116 3516 3124 3524
rect 3132 3516 3140 3524
rect 3212 3516 3220 3524
rect 3324 3516 3332 3524
rect 3132 3416 3140 3424
rect 3116 3396 3124 3404
rect 3132 3376 3140 3384
rect 3132 3316 3140 3324
rect 3132 3196 3140 3204
rect 3068 2596 3076 2604
rect 3116 2916 3124 2924
rect 3180 3416 3188 3424
rect 3212 3416 3220 3424
rect 3180 3396 3188 3404
rect 3228 3376 3236 3384
rect 3116 2896 3124 2904
rect 3100 2736 3108 2744
rect 3100 2676 3108 2684
rect 3100 2516 3108 2524
rect 3132 2716 3140 2724
rect 3132 2476 3140 2484
rect 3020 2256 3028 2264
rect 3020 2216 3028 2224
rect 2988 1876 2996 1884
rect 3004 1876 3012 1884
rect 3020 1876 3028 1884
rect 2972 1856 2980 1864
rect 3020 1836 3028 1844
rect 2956 1716 2964 1724
rect 2956 1676 2964 1684
rect 2988 1756 2996 1764
rect 3004 1756 3012 1764
rect 3020 1696 3028 1704
rect 3020 1676 3028 1684
rect 2988 1656 2996 1664
rect 3004 1656 3012 1664
rect 2988 1516 2996 1524
rect 3004 1516 3012 1524
rect 2956 1456 2964 1464
rect 2972 1456 2980 1464
rect 3004 1396 3012 1404
rect 2988 1356 2996 1364
rect 2876 1256 2884 1264
rect 2908 1256 2916 1264
rect 2828 1136 2836 1144
rect 2796 996 2804 1004
rect 2796 956 2804 964
rect 2780 836 2788 844
rect 2796 816 2804 824
rect 2796 736 2804 744
rect 2748 676 2756 684
rect 2780 676 2788 684
rect 2876 1096 2884 1104
rect 2860 956 2868 964
rect 2828 936 2836 944
rect 2828 916 2836 924
rect 2876 936 2884 944
rect 2860 676 2868 684
rect 2796 656 2804 664
rect 2748 636 2756 644
rect 2796 516 2804 524
rect 2812 516 2820 524
rect 2780 496 2788 504
rect 2716 396 2724 404
rect 2716 236 2724 244
rect 2732 236 2740 244
rect 2812 316 2820 324
rect 2812 236 2820 244
rect 2812 176 2820 184
rect 2860 656 2868 664
rect 2860 496 2868 504
rect 2860 316 2868 324
rect 2860 276 2868 284
rect 2860 236 2868 244
rect 2908 996 2916 1004
rect 2892 896 2900 904
rect 3004 1296 3012 1304
rect 2956 1136 2964 1144
rect 2972 1116 2980 1124
rect 3004 1116 3012 1124
rect 3004 1076 3012 1084
rect 3004 1016 3012 1024
rect 2956 936 2964 944
rect 2956 896 2964 904
rect 2940 876 2948 884
rect 2908 676 2916 684
rect 2908 576 2916 584
rect 2892 456 2900 464
rect 2940 616 2948 624
rect 3004 836 3012 844
rect 3132 2456 3140 2464
rect 3116 2396 3124 2404
rect 3132 2156 3140 2164
rect 3148 2156 3156 2164
rect 3148 2076 3156 2084
rect 3116 1856 3124 1864
rect 3068 1736 3076 1744
rect 3084 1636 3092 1644
rect 3132 1736 3140 1744
rect 3180 3236 3188 3244
rect 3196 2956 3204 2964
rect 3180 2916 3188 2924
rect 3180 2736 3188 2744
rect 3196 2676 3204 2684
rect 3180 2556 3188 2564
rect 3228 2736 3236 2744
rect 3228 2516 3236 2524
rect 3180 2496 3188 2504
rect 3196 2196 3204 2204
rect 3196 1936 3204 1944
rect 3228 2196 3236 2204
rect 3292 3296 3300 3304
rect 3260 2976 3268 2984
rect 3276 2936 3284 2944
rect 3276 2756 3284 2764
rect 3260 2636 3268 2644
rect 3260 2536 3268 2544
rect 3260 2456 3268 2464
rect 3532 3536 3540 3544
rect 3644 3536 3652 3544
rect 3676 3536 3684 3544
rect 3516 3516 3524 3524
rect 3452 3476 3460 3484
rect 3468 3476 3476 3484
rect 3548 3516 3556 3524
rect 3388 3436 3396 3444
rect 3404 3436 3412 3444
rect 3564 3496 3572 3504
rect 3628 3496 3636 3504
rect 3452 3416 3460 3424
rect 3500 3416 3508 3424
rect 3516 3416 3524 3424
rect 3324 3376 3332 3384
rect 3340 3336 3348 3344
rect 3372 3336 3380 3344
rect 3340 3036 3348 3044
rect 3372 3076 3380 3084
rect 3324 2916 3332 2924
rect 3324 2896 3332 2904
rect 3308 2876 3316 2884
rect 3324 2696 3332 2704
rect 3324 2656 3332 2664
rect 3340 2536 3348 2544
rect 3356 2536 3364 2544
rect 3308 2516 3316 2524
rect 3324 2516 3332 2524
rect 3308 2456 3316 2464
rect 3564 3376 3572 3384
rect 3436 3296 3444 3304
rect 3484 3276 3492 3284
rect 3404 3036 3412 3044
rect 3452 3056 3460 3064
rect 3452 3016 3460 3024
rect 3420 2896 3428 2904
rect 3324 2436 3332 2444
rect 3276 2296 3284 2304
rect 3292 2296 3300 2304
rect 3276 2256 3284 2264
rect 3324 2236 3332 2244
rect 3228 1876 3236 1884
rect 3276 2096 3284 2104
rect 3292 2076 3300 2084
rect 3276 2016 3284 2024
rect 3308 1956 3316 1964
rect 3292 1856 3300 1864
rect 3356 2176 3364 2184
rect 3356 2156 3364 2164
rect 3340 1936 3348 1944
rect 3324 1836 3332 1844
rect 3148 1716 3156 1724
rect 3116 1636 3124 1644
rect 3100 1256 3108 1264
rect 3100 1176 3108 1184
rect 3148 1556 3156 1564
rect 3132 1536 3140 1544
rect 3148 1436 3156 1444
rect 3116 1056 3124 1064
rect 3068 1036 3076 1044
rect 3036 816 3044 824
rect 3068 816 3076 824
rect 3020 796 3028 804
rect 3052 716 3060 724
rect 2988 616 2996 624
rect 2940 476 2948 484
rect 2924 396 2932 404
rect 2924 276 2932 284
rect 2924 236 2932 244
rect 2940 236 2948 244
rect 2876 176 2884 184
rect 2892 176 2900 184
rect 2860 156 2868 164
rect 3084 796 3092 804
rect 3068 496 3076 504
rect 3052 456 3060 464
rect 3004 316 3012 324
rect 3004 276 3012 284
rect 2924 156 2932 164
rect 2956 156 2964 164
rect 2620 116 2628 124
rect 2812 96 2820 104
rect 2556 76 2564 84
rect 2908 76 2916 84
rect 3036 296 3044 304
rect 3132 896 3140 904
rect 3180 1436 3188 1444
rect 3228 1736 3236 1744
rect 3244 1576 3252 1584
rect 3228 1536 3236 1544
rect 3260 1516 3268 1524
rect 3212 1456 3220 1464
rect 3180 1076 3188 1084
rect 3180 996 3188 1004
rect 3180 916 3188 924
rect 3180 776 3188 784
rect 3180 616 3188 624
rect 3180 556 3188 564
rect 3100 476 3108 484
rect 3132 476 3140 484
rect 3084 396 3092 404
rect 3116 356 3124 364
rect 3164 316 3172 324
rect 3180 316 3188 324
rect 3084 296 3092 304
rect 3292 1476 3300 1484
rect 3340 1796 3348 1804
rect 3340 1536 3348 1544
rect 3340 1516 3348 1524
rect 3324 1476 3332 1484
rect 3308 1456 3316 1464
rect 3228 1076 3236 1084
rect 3276 1076 3284 1084
rect 3228 856 3236 864
rect 3228 796 3236 804
rect 3260 776 3268 784
rect 3228 636 3236 644
rect 3244 616 3252 624
rect 3228 596 3236 604
rect 3260 476 3268 484
rect 3228 356 3236 364
rect 3132 236 3140 244
rect 3340 1436 3348 1444
rect 3420 2876 3428 2884
rect 3404 2556 3412 2564
rect 3404 2216 3412 2224
rect 3388 1976 3396 1984
rect 3404 1976 3412 1984
rect 3388 1876 3396 1884
rect 3388 1756 3396 1764
rect 3372 1636 3380 1644
rect 3388 1596 3396 1604
rect 3388 1556 3396 1564
rect 3340 1336 3348 1344
rect 3356 1296 3364 1304
rect 3372 1296 3380 1304
rect 3308 1156 3316 1164
rect 3324 1156 3332 1164
rect 3308 876 3316 884
rect 3292 776 3300 784
rect 3292 476 3300 484
rect 3244 276 3252 284
rect 3260 276 3268 284
rect 3228 216 3236 224
rect 3132 176 3140 184
rect 3148 136 3156 144
rect 3196 136 3204 144
rect 3132 96 3140 104
rect 3372 1196 3380 1204
rect 3388 1196 3396 1204
rect 3356 1076 3364 1084
rect 3372 1016 3380 1024
rect 3372 936 3380 944
rect 3372 656 3380 664
rect 3372 496 3380 504
rect 3100 76 3108 84
rect 3164 76 3172 84
rect 3196 56 3204 64
rect 3356 276 3364 284
rect 3372 276 3380 284
rect 3452 2616 3460 2624
rect 3484 2936 3492 2944
rect 3484 2716 3492 2724
rect 3468 2396 3476 2404
rect 3468 2316 3476 2324
rect 3484 2316 3492 2324
rect 3484 2276 3492 2284
rect 3468 2256 3476 2264
rect 3468 2176 3476 2184
rect 3452 2076 3460 2084
rect 3468 2036 3476 2044
rect 3468 2016 3476 2024
rect 3452 1816 3460 1824
rect 3532 3076 3540 3084
rect 3548 3036 3556 3044
rect 3532 2976 3540 2984
rect 3852 3516 3860 3524
rect 3964 3496 3972 3504
rect 4060 3476 4068 3484
rect 3596 3456 3604 3464
rect 3644 3456 3652 3464
rect 3580 3096 3588 3104
rect 3564 2936 3572 2944
rect 3564 2716 3572 2724
rect 3532 2336 3540 2344
rect 3516 2056 3524 2064
rect 3532 1996 3540 2004
rect 3516 1936 3524 1944
rect 3484 1756 3492 1764
rect 3452 1396 3460 1404
rect 3436 1056 3444 1064
rect 3484 1536 3492 1544
rect 3484 1516 3492 1524
rect 3516 1756 3524 1764
rect 3516 1596 3524 1604
rect 3516 1516 3524 1524
rect 3516 1056 3524 1064
rect 3484 1016 3492 1024
rect 3484 936 3492 944
rect 3452 736 3460 744
rect 3468 656 3476 664
rect 3436 616 3444 624
rect 3436 596 3444 604
rect 3452 596 3460 604
rect 3420 576 3428 584
rect 3420 236 3428 244
rect 3436 236 3444 244
rect 3516 636 3524 644
rect 3516 616 3524 624
rect 3580 2336 3588 2344
rect 3676 3376 3684 3384
rect 3628 3076 3636 3084
rect 3676 3016 3684 3024
rect 3612 2996 3620 3004
rect 3628 2936 3636 2944
rect 3740 3396 3748 3404
rect 3692 2916 3700 2924
rect 3612 2596 3620 2604
rect 3660 2656 3668 2664
rect 3580 2096 3588 2104
rect 3580 1916 3588 1924
rect 3580 1896 3588 1904
rect 3580 1876 3588 1884
rect 3660 2316 3668 2324
rect 3644 2256 3652 2264
rect 3660 2216 3668 2224
rect 3628 2176 3636 2184
rect 3644 2176 3652 2184
rect 3628 1896 3636 1904
rect 3628 1776 3636 1784
rect 3580 1736 3588 1744
rect 3644 1676 3652 1684
rect 3644 1596 3652 1604
rect 3628 1516 3636 1524
rect 3564 1136 3572 1144
rect 3564 996 3572 1004
rect 3548 876 3556 884
rect 3564 676 3572 684
rect 3468 336 3476 344
rect 3500 316 3508 324
rect 3612 1336 3620 1344
rect 3596 1236 3604 1244
rect 3628 1236 3636 1244
rect 3628 1136 3636 1144
rect 3628 1036 3636 1044
rect 3612 956 3620 964
rect 3628 956 3636 964
rect 3644 896 3652 904
rect 3660 536 3668 544
rect 3612 276 3620 284
rect 3708 2596 3716 2604
rect 3692 2276 3700 2284
rect 3708 2156 3716 2164
rect 3804 3376 3812 3384
rect 3740 3256 3748 3264
rect 3788 3136 3796 3144
rect 3772 3096 3780 3104
rect 3756 2636 3764 2644
rect 3740 2416 3748 2424
rect 3692 1996 3700 2004
rect 3692 1896 3700 1904
rect 3772 2476 3780 2484
rect 3772 2336 3780 2344
rect 3788 2216 3796 2224
rect 3756 2156 3764 2164
rect 3756 2116 3764 2124
rect 3772 2036 3780 2044
rect 3724 1856 3732 1864
rect 3740 1796 3748 1804
rect 3724 1776 3732 1784
rect 3724 1716 3732 1724
rect 3708 1316 3716 1324
rect 3708 1116 3716 1124
rect 3740 1196 3748 1204
rect 3724 1096 3732 1104
rect 3692 1036 3700 1044
rect 3708 976 3716 984
rect 3724 956 3732 964
rect 3708 936 3716 944
rect 3724 856 3732 864
rect 3740 716 3748 724
rect 3724 696 3732 704
rect 3692 576 3700 584
rect 3692 536 3700 544
rect 3724 476 3732 484
rect 3500 256 3508 264
rect 3660 216 3668 224
rect 3548 156 3556 164
rect 3580 156 3588 164
rect 3596 136 3604 144
rect 3628 136 3636 144
rect 3388 116 3396 124
rect 3468 116 3476 124
rect 3340 36 3348 44
rect 3692 156 3700 164
rect 3948 3456 3956 3464
rect 3900 3436 3908 3444
rect 3932 3436 3940 3444
rect 4060 3376 4068 3384
rect 4012 3356 4020 3364
rect 3852 3176 3860 3184
rect 3868 2916 3876 2924
rect 3820 2296 3828 2304
rect 3820 2256 3828 2264
rect 3820 2216 3828 2224
rect 3820 2176 3828 2184
rect 3820 2116 3828 2124
rect 3852 2636 3860 2644
rect 3868 2636 3876 2644
rect 3852 2596 3860 2604
rect 3884 2516 3892 2524
rect 3932 2956 3940 2964
rect 3916 2596 3924 2604
rect 3884 2496 3892 2504
rect 3852 2396 3860 2404
rect 3836 1856 3844 1864
rect 3836 1736 3844 1744
rect 3804 1716 3812 1724
rect 3804 1596 3812 1604
rect 3788 1296 3796 1304
rect 3868 2256 3876 2264
rect 3868 2176 3876 2184
rect 3868 2076 3876 2084
rect 3932 2356 3940 2364
rect 3900 2296 3908 2304
rect 3884 1876 3892 1884
rect 3884 1736 3892 1744
rect 3884 1356 3892 1364
rect 3836 1336 3844 1344
rect 3852 1336 3860 1344
rect 3932 2136 3940 2144
rect 3916 2016 3924 2024
rect 3804 1256 3812 1264
rect 3820 1256 3828 1264
rect 3788 1216 3796 1224
rect 3852 1196 3860 1204
rect 3788 1156 3796 1164
rect 3804 1136 3812 1144
rect 3836 1136 3844 1144
rect 3916 1216 3924 1224
rect 3916 1096 3924 1104
rect 3900 1076 3908 1084
rect 3820 1036 3828 1044
rect 3804 976 3812 984
rect 3788 876 3796 884
rect 3852 996 3860 1004
rect 3836 976 3844 984
rect 4044 3296 4052 3304
rect 4012 3136 4020 3144
rect 4060 3096 4068 3104
rect 3980 3036 3988 3044
rect 4012 3016 4020 3024
rect 4044 2916 4052 2924
rect 4028 2636 4036 2644
rect 3996 2576 4004 2584
rect 4012 2576 4020 2584
rect 4012 2416 4020 2424
rect 3980 2136 3988 2144
rect 3948 1916 3956 1924
rect 3964 1856 3972 1864
rect 3996 1996 4004 2004
rect 3996 1916 4004 1924
rect 3980 1816 3988 1824
rect 3996 1816 4004 1824
rect 3948 1796 3956 1804
rect 3964 1776 3972 1784
rect 3996 1736 4004 1744
rect 3980 1556 3988 1564
rect 3996 1536 4004 1544
rect 3916 976 3924 984
rect 3884 876 3892 884
rect 3948 876 3956 884
rect 3884 856 3892 864
rect 3820 776 3828 784
rect 3948 776 3956 784
rect 3788 496 3796 504
rect 3868 756 3876 764
rect 3932 756 3940 764
rect 3836 696 3844 704
rect 3836 676 3844 684
rect 3900 696 3908 704
rect 3948 696 3956 704
rect 3916 616 3924 624
rect 3980 1216 3988 1224
rect 3996 1156 4004 1164
rect 3980 1116 3988 1124
rect 3980 976 3988 984
rect 3980 736 3988 744
rect 3996 736 4004 744
rect 4316 3496 4324 3504
rect 4316 3476 4324 3484
rect 4380 3456 4388 3464
rect 4092 3436 4100 3444
rect 4188 3436 4196 3444
rect 4156 3396 4164 3404
rect 4092 3376 4100 3384
rect 4188 3336 4196 3344
rect 4172 3036 4180 3044
rect 4140 2936 4148 2944
rect 4092 2516 4100 2524
rect 4076 2496 4084 2504
rect 4108 2456 4116 2464
rect 4076 2396 4084 2404
rect 4076 2356 4084 2364
rect 4156 2756 4164 2764
rect 4140 2676 4148 2684
rect 4140 2636 4148 2644
rect 4140 2596 4148 2604
rect 4172 2676 4180 2684
rect 4156 2556 4164 2564
rect 4156 2516 4164 2524
rect 4140 2496 4148 2504
rect 4140 2476 4148 2484
rect 4124 2356 4132 2364
rect 4156 2316 4164 2324
rect 4092 2216 4100 2224
rect 4092 2116 4100 2124
rect 4124 2296 4132 2304
rect 4124 2256 4132 2264
rect 4124 2176 4132 2184
rect 4156 2116 4164 2124
rect 4108 1976 4116 1984
rect 4060 1956 4068 1964
rect 4076 1936 4084 1944
rect 4076 1876 4084 1884
rect 4044 1756 4052 1764
rect 4060 1736 4068 1744
rect 4060 1456 4068 1464
rect 4044 1356 4052 1364
rect 4060 896 4068 904
rect 4044 796 4052 804
rect 4044 756 4052 764
rect 4108 1836 4116 1844
rect 4092 1676 4100 1684
rect 3996 716 4004 724
rect 4012 716 4020 724
rect 3980 696 3988 704
rect 4028 696 4036 704
rect 4044 696 4052 704
rect 4012 616 4020 624
rect 4028 596 4036 604
rect 3964 556 3972 564
rect 3884 516 3892 524
rect 3900 516 3908 524
rect 3836 376 3844 384
rect 3804 316 3812 324
rect 3820 276 3828 284
rect 3788 256 3796 264
rect 3948 496 3956 504
rect 3948 336 3956 344
rect 3884 276 3892 284
rect 3868 256 3876 264
rect 3852 236 3860 244
rect 3900 236 3908 244
rect 3916 236 3924 244
rect 3804 196 3812 204
rect 4044 556 4052 564
rect 4028 496 4036 504
rect 4012 476 4020 484
rect 3996 356 4004 364
rect 3980 296 3988 304
rect 3788 136 3796 144
rect 3980 116 3988 124
rect 4076 696 4084 704
rect 4076 596 4084 604
rect 4124 1776 4132 1784
rect 4140 1736 4148 1744
rect 4140 1516 4148 1524
rect 4108 1456 4116 1464
rect 4108 1396 4116 1404
rect 4124 1356 4132 1364
rect 4124 1296 4132 1304
rect 4140 1296 4148 1304
rect 4108 816 4116 824
rect 4108 596 4116 604
rect 4140 1036 4148 1044
rect 4140 956 4148 964
rect 4140 756 4148 764
rect 4364 3336 4372 3344
rect 4188 2236 4196 2244
rect 4348 3156 4356 3164
rect 4460 3416 4468 3424
rect 4460 3376 4468 3384
rect 4524 3336 4532 3344
rect 4700 3456 4708 3464
rect 4716 3456 4724 3464
rect 4828 3456 4836 3464
rect 4940 3456 4948 3464
rect 4588 3436 4596 3444
rect 4604 3436 4612 3444
rect 4636 3236 4644 3244
rect 4460 2976 4468 2984
rect 4348 2956 4356 2964
rect 4332 2936 4340 2944
rect 4236 2836 4244 2844
rect 4284 2716 4292 2724
rect 4300 2656 4308 2664
rect 4332 2656 4340 2664
rect 4268 2516 4276 2524
rect 4236 2296 4244 2304
rect 4508 2956 4516 2964
rect 4364 2736 4372 2744
rect 4364 2716 4372 2724
rect 4396 2656 4404 2664
rect 4364 2576 4372 2584
rect 4508 2736 4516 2744
rect 4556 3036 4564 3044
rect 4572 2976 4580 2984
rect 4556 2936 4564 2944
rect 4524 2716 4532 2724
rect 4476 2676 4484 2684
rect 4444 2656 4452 2664
rect 4508 2656 4516 2664
rect 4444 2636 4452 2644
rect 4460 2616 4468 2624
rect 4412 2556 4420 2564
rect 4348 2436 4356 2444
rect 4252 2176 4260 2184
rect 4188 1636 4196 1644
rect 4188 1596 4196 1604
rect 4188 1536 4196 1544
rect 4220 1616 4228 1624
rect 4188 1456 4196 1464
rect 4188 916 4196 924
rect 4188 876 4196 884
rect 4140 696 4148 704
rect 4140 676 4148 684
rect 4156 656 4164 664
rect 4140 616 4148 624
rect 4172 596 4180 604
rect 4220 1216 4228 1224
rect 4220 1076 4228 1084
rect 4252 2116 4260 2124
rect 4252 1936 4260 1944
rect 4252 1876 4260 1884
rect 4332 2256 4340 2264
rect 4300 2156 4308 2164
rect 4300 1956 4308 1964
rect 4284 1856 4292 1864
rect 4268 1516 4276 1524
rect 4268 1496 4276 1504
rect 4268 1436 4276 1444
rect 4316 1876 4324 1884
rect 4316 1836 4324 1844
rect 4348 2136 4356 2144
rect 4428 2276 4436 2284
rect 4396 2216 4404 2224
rect 4380 2056 4388 2064
rect 4364 1896 4372 1904
rect 4316 1676 4324 1684
rect 4348 1716 4356 1724
rect 4364 1716 4372 1724
rect 4332 1456 4340 1464
rect 4284 1376 4292 1384
rect 4268 1176 4276 1184
rect 4252 1096 4260 1104
rect 4300 1116 4308 1124
rect 4332 1396 4340 1404
rect 4332 1236 4340 1244
rect 4284 1056 4292 1064
rect 4252 1036 4260 1044
rect 4220 796 4228 804
rect 4220 616 4228 624
rect 4332 896 4340 904
rect 4140 556 4148 564
rect 4188 536 4196 544
rect 4076 416 4084 424
rect 4172 396 4180 404
rect 4236 336 4244 344
rect 4124 316 4132 324
rect 4380 1676 4388 1684
rect 4380 1596 4388 1604
rect 4444 2116 4452 2124
rect 4444 2096 4452 2104
rect 4540 2556 4548 2564
rect 4492 2496 4500 2504
rect 4508 2496 4516 2504
rect 4492 2476 4500 2484
rect 4476 2196 4484 2204
rect 4476 2136 4484 2144
rect 4476 2036 4484 2044
rect 4508 2096 4516 2104
rect 4492 1996 4500 2004
rect 4412 1556 4420 1564
rect 4412 1456 4420 1464
rect 4444 1376 4452 1384
rect 4476 1356 4484 1364
rect 4412 1316 4420 1324
rect 4444 1276 4452 1284
rect 4428 1256 4436 1264
rect 4364 1196 4372 1204
rect 4412 1116 4420 1124
rect 4380 956 4388 964
rect 4412 916 4420 924
rect 4412 716 4420 724
rect 4572 2636 4580 2644
rect 4556 2276 4564 2284
rect 4540 2116 4548 2124
rect 4508 1416 4516 1424
rect 4524 1356 4532 1364
rect 4508 1316 4516 1324
rect 4492 956 4500 964
rect 4524 1236 4532 1244
rect 4460 936 4468 944
rect 4524 916 4532 924
rect 4508 736 4516 744
rect 4492 676 4500 684
rect 4604 3076 4612 3084
rect 4828 3436 4836 3444
rect 4684 3076 4692 3084
rect 4652 3036 4660 3044
rect 4652 3016 4660 3024
rect 4652 2796 4660 2804
rect 4636 2116 4644 2124
rect 4684 2716 4692 2724
rect 4604 2096 4612 2104
rect 4668 2076 4676 2084
rect 4620 1916 4628 1924
rect 4604 1796 4612 1804
rect 4652 1776 4660 1784
rect 4668 1736 4676 1744
rect 4636 1596 4644 1604
rect 4764 3136 4772 3144
rect 4748 3116 4756 3124
rect 4732 2936 4740 2944
rect 4700 1596 4708 1604
rect 4572 1396 4580 1404
rect 4556 1376 4564 1384
rect 4588 1376 4596 1384
rect 4636 1376 4644 1384
rect 4652 1376 4660 1384
rect 4604 1136 4612 1144
rect 4556 1096 4564 1104
rect 4572 1076 4580 1084
rect 4444 656 4452 664
rect 4540 636 4548 644
rect 4540 556 4548 564
rect 4428 476 4436 484
rect 4172 276 4180 284
rect 4204 216 4212 224
rect 4300 216 4308 224
rect 4412 216 4420 224
rect 4092 196 4100 204
rect 4332 196 4340 204
rect 4060 116 4068 124
rect 4140 176 4148 184
rect 4636 1016 4644 1024
rect 4636 736 4644 744
rect 4604 516 4612 524
rect 4636 676 4644 684
rect 4668 1296 4676 1304
rect 4636 496 4644 504
rect 4636 336 4644 344
rect 4652 276 4660 284
rect 4716 1456 4724 1464
rect 4796 2696 4804 2704
rect 4764 2516 4772 2524
rect 4764 2256 4772 2264
rect 4780 2236 4788 2244
rect 4764 1756 4772 1764
rect 4764 1316 4772 1324
rect 4748 1056 4756 1064
rect 4732 1016 4740 1024
rect 4764 1016 4772 1024
rect 4732 996 4740 1004
rect 4684 556 4692 564
rect 4748 836 4756 844
rect 4828 2756 4836 2764
rect 4908 3316 4916 3324
rect 4860 2696 4868 2704
rect 4812 2016 4820 2024
rect 4796 1816 4804 1824
rect 4828 1696 4836 1704
rect 4892 2676 4900 2684
rect 4892 2636 4900 2644
rect 4876 2496 4884 2504
rect 4876 2336 4884 2344
rect 4860 2256 4868 2264
rect 4860 2136 4868 2144
rect 5036 3476 5044 3484
rect 5052 3356 5060 3364
rect 4908 1956 4916 1964
rect 4860 1816 4868 1824
rect 4860 1796 4868 1804
rect 4796 1096 4804 1104
rect 4796 616 4804 624
rect 4796 536 4804 544
rect 4828 1576 4836 1584
rect 4844 1536 4852 1544
rect 4844 1516 4852 1524
rect 4828 1476 4836 1484
rect 4828 1376 4836 1384
rect 4828 1256 4836 1264
rect 4844 1076 4852 1084
rect 4780 276 4788 284
rect 4780 216 4788 224
rect 4844 216 4852 224
rect 4524 176 4532 184
rect 4780 176 4788 184
rect 4876 1436 4884 1444
rect 4876 1316 4884 1324
rect 4876 1276 4884 1284
rect 5116 3356 5124 3364
rect 5116 3336 5124 3344
rect 4956 2536 4964 2544
rect 4956 2496 4964 2504
rect 4988 2276 4996 2284
rect 4972 2116 4980 2124
rect 4956 1956 4964 1964
rect 4924 1456 4932 1464
rect 4892 976 4900 984
rect 4876 536 4884 544
rect 4828 156 4836 164
rect 4940 956 4948 964
rect 4924 576 4932 584
rect 5052 2776 5060 2784
rect 5052 2636 5060 2644
rect 5052 2496 5060 2504
rect 5004 1716 5012 1724
rect 5004 1656 5012 1664
rect 5084 2736 5092 2744
rect 5084 2696 5092 2704
rect 5084 2676 5092 2684
rect 5116 2736 5124 2744
rect 5116 2656 5124 2664
rect 5100 2036 5108 2044
rect 5100 1996 5108 2004
rect 5100 1976 5108 1984
rect 5084 1776 5092 1784
rect 5084 1716 5092 1724
rect 5084 1496 5092 1504
rect 5100 1496 5108 1504
rect 4972 1456 4980 1464
rect 5004 1436 5012 1444
rect 5004 1336 5012 1344
rect 5068 1296 5076 1304
rect 5068 1116 5076 1124
rect 4988 1056 4996 1064
rect 5036 996 5044 1004
rect 5100 956 5108 964
rect 5084 836 5092 844
rect 5036 776 5044 784
rect 5100 696 5108 704
rect 5036 656 5044 664
rect 5004 636 5012 644
rect 4988 136 4996 144
rect 5068 556 5076 564
rect 5164 3436 5172 3444
rect 5148 2876 5156 2884
rect 5148 1356 5156 1364
rect 5196 1056 5204 1064
rect 5180 896 5188 904
rect 5148 816 5156 824
rect 5132 636 5140 644
rect 5132 596 5140 604
rect 5116 536 5124 544
rect 5164 776 5172 784
rect 5132 276 5140 284
rect 5068 256 5076 264
rect 5068 176 5076 184
rect 5164 156 5172 164
rect 4156 116 4164 124
rect 4204 116 4212 124
rect 4540 116 4548 124
rect 1996 16 2004 24
rect 2492 16 2500 24
rect 3404 16 3412 24
<< metal5 >>
rect 484 3537 2524 3543
rect 3540 3537 3644 3543
rect 3669 3537 3676 3543
rect 1396 3517 2060 3523
rect 2164 3517 2220 3523
rect 2740 3517 2828 3523
rect 2852 3517 3116 3523
rect 3140 3517 3212 3523
rect 3332 3517 3515 3523
rect 3556 3517 3852 3523
rect 980 3497 1811 3503
rect 484 3477 796 3483
rect 964 3477 1244 3483
rect 1805 3483 1811 3497
rect 1828 3497 1916 3503
rect 2068 3497 2652 3503
rect 2669 3497 3564 3503
rect 2669 3483 2675 3497
rect 3572 3497 3611 3503
rect 3636 3497 3964 3503
rect 3972 3497 4316 3503
rect 1805 3477 2675 3483
rect 2692 3477 3452 3483
rect 3476 3477 4060 3483
rect 4324 3477 5036 3483
rect 420 3457 556 3463
rect 852 3457 1036 3463
rect 2084 3457 2475 3463
rect 2500 3457 3596 3463
rect 3652 3457 3948 3463
rect 3956 3457 4380 3463
rect 4388 3457 4700 3463
rect 4724 3457 4811 3463
rect 4836 3457 4940 3463
rect 1092 3437 1267 3443
rect 1261 3423 1267 3437
rect 2228 3437 2235 3443
rect 2372 3437 2395 3443
rect 2516 3437 2523 3443
rect 2548 3437 3388 3443
rect 3412 3437 3900 3443
rect 3940 3437 4092 3443
rect 4100 3437 4188 3443
rect 4453 3437 4588 3443
rect 4612 3437 4828 3443
rect 4869 3437 5164 3443
rect 1261 3417 2316 3423
rect 2725 3417 2796 3423
rect 2820 3417 3132 3423
rect 3188 3417 3195 3423
rect 3220 3417 3452 3423
rect 3493 3417 3500 3423
rect 3524 3417 4460 3423
rect 2740 3397 3020 3403
rect 3045 3397 3116 3403
rect 3188 3397 3347 3403
rect 3133 3384 3139 3395
rect 164 3377 588 3383
rect 740 3377 1644 3383
rect 2340 3377 2508 3383
rect 2596 3377 2787 3383
rect 948 3357 1004 3363
rect 1028 3357 1308 3363
rect 1348 3357 2108 3363
rect 2180 3357 2236 3363
rect 2612 3357 2764 3363
rect 2781 3363 2787 3377
rect 2980 3377 3091 3383
rect 2781 3357 3035 3363
rect 3060 3357 3067 3363
rect 3085 3363 3091 3377
rect 3341 3383 3347 3397
rect 3397 3397 3707 3403
rect 3748 3397 4156 3403
rect 3341 3377 3564 3383
rect 3589 3377 3659 3383
rect 3684 3377 3804 3383
rect 3829 3377 4060 3383
rect 4100 3377 4460 3383
rect 3085 3357 4012 3363
rect 4037 3357 5052 3363
rect 372 3337 1036 3343
rect 1156 3337 1196 3343
rect 1268 3337 1452 3343
rect 1684 3337 1851 3343
rect 1876 3337 1883 3343
rect 2132 3337 2188 3343
rect 2372 3337 2444 3343
rect 2509 3337 3340 3343
rect 772 3317 827 3323
rect 2509 3323 2515 3337
rect 3380 3337 4188 3343
rect 4372 3337 4524 3343
rect 4933 3337 5116 3343
rect 900 3317 2515 3323
rect 2533 3317 3132 3323
rect 4901 3317 4908 3323
rect 372 3297 828 3303
rect 836 3297 2924 3303
rect 2996 3297 3131 3303
rect 3300 3297 3419 3303
rect 3444 3297 4044 3303
rect 4052 3297 4251 3303
rect 292 3277 492 3283
rect 740 3277 3484 3283
rect 1300 3257 3067 3263
rect 3077 3257 3740 3263
rect 1861 3237 1868 3243
rect 3188 3237 4636 3243
rect 765 3224 771 3235
rect 1876 3217 2412 3223
rect 1605 3197 3132 3203
rect 2693 3177 3852 3183
rect 100 3157 460 3163
rect 1364 3157 1371 3163
rect 1389 3157 2028 3163
rect 1389 3143 1395 3157
rect 2548 3157 4348 3163
rect 948 3137 1395 3143
rect 1765 3137 2716 3143
rect 3044 3137 3788 3143
rect 4020 3137 4764 3143
rect 708 3117 1308 3123
rect 1364 3117 1404 3123
rect 1669 3117 1676 3123
rect 1684 3117 2988 3123
rect 3077 3117 4748 3123
rect 4756 3117 4763 3123
rect 180 3097 316 3103
rect 532 3097 764 3103
rect 1044 3097 1132 3103
rect 1204 3097 1755 3103
rect 1780 3097 1891 3103
rect 772 3077 1004 3083
rect 1012 3077 1868 3083
rect 1885 3083 1891 3097
rect 2116 3097 3580 3103
rect 3780 3097 4060 3103
rect 1885 3077 2204 3083
rect 2228 3077 2844 3083
rect 2852 3077 3372 3083
rect 3540 3077 3628 3083
rect 4612 3077 4684 3083
rect 244 3057 1628 3063
rect 1636 3057 2780 3063
rect 2804 3057 3452 3063
rect 1092 3037 1308 3043
rect 1445 3037 1484 3043
rect 1540 3037 1772 3043
rect 1876 3037 2476 3043
rect 2501 3037 2540 3043
rect 2676 3037 3067 3043
rect 3549 3044 3555 3055
rect 3348 3037 3404 3043
rect 3988 3037 4172 3043
rect 4564 3037 4652 3043
rect 1012 3017 2524 3023
rect 2756 3017 2924 3023
rect 3460 3017 3676 3023
rect 4020 3017 4652 3023
rect 804 2997 940 3003
rect 1876 2997 1900 3003
rect 1940 2997 2075 3003
rect 2100 2997 2156 3003
rect 2181 2997 2588 3003
rect 2916 2997 3612 3003
rect 1140 2977 3131 2983
rect 3268 2977 3532 2983
rect 4468 2977 4572 2983
rect 948 2957 2860 2963
rect 2980 2957 3196 2963
rect 3940 2957 4348 2963
rect 4356 2957 4508 2963
rect 980 2937 1340 2943
rect 1460 2937 1772 2943
rect 1828 2937 2012 2943
rect 2388 2937 2411 2943
rect 2436 2937 2508 2943
rect 2548 2937 2723 2943
rect 308 2917 540 2923
rect 980 2917 1036 2923
rect 1140 2917 1267 2923
rect 413 2897 428 2903
rect 436 2897 604 2903
rect 1076 2897 1179 2903
rect 1261 2903 1267 2917
rect 1348 2917 1371 2923
rect 1444 2917 1596 2923
rect 1733 2917 2203 2923
rect 2213 2917 2459 2923
rect 2501 2917 2700 2923
rect 2717 2923 2723 2937
rect 2772 2937 2828 2943
rect 2964 2937 3020 2943
rect 3284 2937 3484 2943
rect 3572 2937 3628 2943
rect 4045 2937 4140 2943
rect 2717 2917 2876 2923
rect 4045 2924 4051 2937
rect 4340 2937 4556 2943
rect 4564 2937 4732 2943
rect 3109 2917 3116 2923
rect 3188 2917 3323 2923
rect 3700 2917 3868 2923
rect 1261 2897 1452 2903
rect 1588 2897 1900 2903
rect 2100 2897 2300 2903
rect 2324 2897 3116 2903
rect 3332 2897 3420 2903
rect 724 2877 1051 2883
rect 1245 2884 1251 2895
rect 1445 2877 1452 2883
rect 1716 2877 1723 2883
rect 1925 2877 1932 2883
rect 2116 2877 2780 2883
rect 3316 2877 3420 2883
rect 3428 2877 3451 2883
rect 5149 2884 5155 2895
rect 805 2857 812 2863
rect 1636 2857 1804 2863
rect 1908 2857 2188 2863
rect 2228 2857 2924 2863
rect 1893 2837 2828 2843
rect 2884 2837 4236 2843
rect 1588 2817 2043 2823
rect 2436 2817 2956 2823
rect 1972 2797 2235 2803
rect 2245 2797 4652 2803
rect 820 2777 2076 2783
rect 2373 2777 5052 2783
rect 708 2757 763 2763
rect 1636 2757 3276 2763
rect 3301 2757 4156 2763
rect 485 2737 492 2743
rect 2004 2737 2188 2743
rect 2628 2737 2683 2743
rect 2708 2737 2939 2743
rect 2964 2737 3020 2743
rect 3108 2737 3171 2743
rect 420 2717 1196 2723
rect 1300 2717 1372 2723
rect 1380 2717 2012 2723
rect 2053 2717 2428 2723
rect 2596 2717 2748 2723
rect 3165 2723 3171 2737
rect 3188 2737 3228 2743
rect 4509 2744 4515 2755
rect 4829 2745 4835 2756
rect 4325 2737 4364 2743
rect 5092 2737 5116 2743
rect 3165 2717 3484 2723
rect 3525 2717 3564 2723
rect 4292 2717 4364 2723
rect 4532 2717 4684 2723
rect 116 2697 284 2703
rect 468 2697 588 2703
rect 756 2697 1132 2703
rect 1509 2697 1516 2703
rect 1812 2697 1900 2703
rect 5085 2704 5091 2715
rect 2277 2697 2556 2703
rect 2628 2697 3324 2703
rect 3332 2697 4796 2703
rect 4804 2697 4860 2703
rect 212 2677 380 2683
rect 388 2677 860 2683
rect 868 2677 1516 2683
rect 1541 2677 1996 2683
rect 2036 2677 2235 2683
rect 2388 2677 3100 2683
rect 3204 2677 4140 2683
rect 4180 2677 4476 2683
rect 4900 2677 5084 2683
rect 180 2657 252 2663
rect 436 2657 475 2663
rect 516 2657 748 2663
rect 965 2657 972 2663
rect 1252 2657 1836 2663
rect 1861 2657 2044 2663
rect 2052 2657 2156 2663
rect 2180 2657 2380 2663
rect 2388 2657 2668 2663
rect 2804 2657 3036 2663
rect 3332 2657 3660 2663
rect 3668 2657 4300 2663
rect 4340 2657 4396 2663
rect 4452 2657 4508 2663
rect 420 2637 540 2643
rect 980 2637 1467 2643
rect 1509 2637 1531 2643
rect 1716 2637 1852 2643
rect 2052 2637 2092 2643
rect 2309 2637 2316 2643
rect 2532 2637 2700 2643
rect 3268 2637 3756 2643
rect 3845 2637 3852 2643
rect 3876 2637 3995 2643
rect 4036 2637 4140 2643
rect 4148 2637 4155 2643
rect 5053 2644 5059 2655
rect 4197 2637 4444 2643
rect 4580 2637 4892 2643
rect 756 2617 2188 2623
rect 2436 2617 2459 2623
rect 2501 2617 2908 2623
rect 3460 2617 4460 2623
rect 372 2597 819 2603
rect 772 2577 795 2583
rect 813 2583 819 2597
rect 1300 2597 1340 2603
rect 1357 2597 1788 2603
rect 1357 2583 1363 2597
rect 2052 2597 2332 2603
rect 2420 2597 3068 2603
rect 3620 2597 3708 2603
rect 3860 2597 3867 2603
rect 3924 2597 4140 2603
rect 813 2577 1363 2583
rect 1396 2577 1436 2583
rect 1588 2577 1708 2583
rect 1765 2577 1788 2583
rect 1844 2577 3996 2583
rect 4020 2577 4364 2583
rect 548 2557 828 2563
rect 884 2557 923 2563
rect 1316 2557 1388 2563
rect 1412 2557 1435 2563
rect 1477 2557 1564 2563
rect 1956 2557 2172 2563
rect 2196 2557 2556 2563
rect 2597 2557 2700 2563
rect 2757 2557 2924 2563
rect 3077 2557 3180 2563
rect 3412 2557 4156 2563
rect 4420 2557 4540 2563
rect 453 2537 556 2543
rect 564 2537 891 2543
rect 1348 2537 1468 2543
rect 1844 2537 1980 2543
rect 2021 2537 2028 2543
rect 2244 2537 2508 2543
rect 2676 2537 2796 2543
rect 2853 2537 3251 2543
rect 708 2517 795 2523
rect 836 2517 1308 2523
rect 1325 2517 2491 2523
rect 1325 2503 1331 2517
rect 2509 2517 2587 2523
rect 452 2497 1331 2503
rect 1373 2497 1516 2503
rect 1373 2483 1379 2497
rect 1636 2497 1900 2503
rect 2196 2497 2284 2503
rect 2509 2503 2515 2517
rect 2692 2517 3020 2523
rect 3108 2517 3228 2523
rect 3245 2523 3251 2537
rect 3268 2537 3340 2543
rect 3364 2537 4956 2543
rect 3245 2517 3308 2523
rect 3332 2517 3884 2523
rect 3892 2517 4092 2523
rect 4164 2517 4187 2523
rect 4261 2517 4268 2523
rect 4276 2517 4764 2523
rect 2308 2497 2515 2503
rect 2661 2497 2748 2503
rect 2868 2497 2875 2503
rect 2885 2497 2971 2503
rect 3013 2497 3131 2503
rect 3188 2497 3884 2503
rect 3909 2497 4076 2503
rect 4148 2497 4492 2503
rect 4516 2497 4876 2503
rect 4964 2497 5052 2503
rect 836 2477 1379 2483
rect 1396 2477 1580 2483
rect 2557 2484 2563 2495
rect 1972 2477 2547 2483
rect 413 2457 1275 2463
rect 413 2443 419 2457
rect 1629 2464 1635 2475
rect 1348 2457 1619 2463
rect 356 2437 419 2443
rect 884 2437 1132 2443
rect 1588 2437 1595 2443
rect 1613 2443 1619 2457
rect 1684 2457 2076 2463
rect 2436 2457 2459 2463
rect 2541 2463 2547 2477
rect 2653 2477 2779 2483
rect 2653 2463 2659 2477
rect 2804 2477 2883 2483
rect 2541 2457 2659 2463
rect 2676 2457 2843 2463
rect 2877 2464 2883 2477
rect 2917 2477 3132 2483
rect 3140 2477 3739 2483
rect 3780 2477 4140 2483
rect 4500 2477 4507 2483
rect 2981 2457 2988 2463
rect 3013 2457 3020 2463
rect 3268 2457 3291 2463
rect 3316 2457 4108 2463
rect 1613 2437 2428 2443
rect 2452 2437 2811 2443
rect 2821 2437 3324 2443
rect 4293 2437 4348 2443
rect 980 2417 1804 2423
rect 1893 2417 1915 2423
rect 1925 2417 2700 2423
rect 2789 2417 2876 2423
rect 2900 2417 3740 2423
rect 4020 2417 4027 2423
rect 1285 2397 3116 2403
rect 3476 2397 3852 2403
rect 4069 2397 4076 2403
rect 1140 2377 1804 2383
rect 2132 2377 2156 2383
rect 2276 2377 3091 2383
rect 932 2357 1932 2363
rect 1940 2357 2956 2363
rect 3085 2363 3091 2377
rect 3109 2377 4091 2383
rect 4101 2377 4699 2383
rect 3085 2357 3932 2363
rect 4084 2357 4124 2363
rect 468 2337 604 2343
rect 1125 2337 1132 2343
rect 1540 2337 2668 2343
rect 2692 2337 3532 2343
rect 3588 2337 3772 2343
rect 4005 2337 4876 2343
rect 580 2317 1420 2323
rect 1509 2317 1532 2323
rect 1588 2317 2124 2323
rect 2212 2317 2396 2323
rect 2413 2317 2779 2323
rect 340 2297 508 2303
rect 580 2297 732 2303
rect 749 2297 972 2303
rect 749 2283 755 2297
rect 2413 2303 2419 2317
rect 2884 2317 3003 2323
rect 3028 2317 3468 2323
rect 3668 2317 4156 2323
rect 1428 2297 2419 2303
rect 2437 2297 2588 2303
rect 2756 2297 2844 2303
rect 2884 2297 3276 2303
rect 3300 2297 3820 2303
rect 3828 2297 3900 2303
rect 4132 2297 4236 2303
rect 500 2277 755 2283
rect 868 2277 924 2283
rect 1108 2277 1436 2283
rect 1524 2277 2003 2283
rect 180 2257 220 2263
rect 340 2257 347 2263
rect 837 2257 844 2263
rect 869 2257 1723 2263
rect 1860 2257 1979 2263
rect 1997 2263 2003 2277
rect 2404 2277 2476 2283
rect 2532 2277 2668 2283
rect 2788 2277 2812 2283
rect 2820 2277 3484 2283
rect 3492 2277 3692 2283
rect 3709 2277 4428 2283
rect 1997 2257 2556 2263
rect 2596 2257 2684 2263
rect 2852 2257 3020 2263
rect 3284 2257 3468 2263
rect 3709 2263 3715 2277
rect 4564 2277 4988 2283
rect 3652 2257 3715 2263
rect 3781 2257 3820 2263
rect 3876 2257 3883 2263
rect 3973 2257 4124 2263
rect 4189 2257 4332 2263
rect 477 2244 483 2255
rect 708 2237 1052 2243
rect 1220 2237 2588 2243
rect 4189 2244 4195 2257
rect 4772 2257 4860 2263
rect 2629 2237 2691 2243
rect 676 2217 859 2223
rect 1396 2217 1819 2223
rect 1860 2217 1883 2223
rect 1924 2217 2412 2223
rect 2564 2217 2651 2223
rect 2685 2223 2691 2237
rect 2756 2237 2812 2243
rect 2852 2237 3324 2243
rect 3405 2237 4179 2243
rect 2685 2217 2764 2223
rect 3405 2224 3411 2237
rect 2853 2217 3020 2223
rect 3668 2217 3771 2223
rect 3796 2217 3803 2223
rect 3828 2217 3963 2223
rect 4173 2223 4179 2237
rect 4788 2237 4795 2243
rect 4173 2217 4396 2223
rect 4093 2205 4099 2216
rect 276 2197 1299 2203
rect 212 2177 252 2183
rect 293 2177 716 2183
rect 741 2177 748 2183
rect 1268 2177 1275 2183
rect 1293 2183 1299 2197
rect 1348 2197 1467 2203
rect 1540 2197 1628 2203
rect 1716 2197 2044 2203
rect 2196 2197 2268 2203
rect 2308 2197 2476 2203
rect 2532 2197 2940 2203
rect 2981 2197 3196 2203
rect 3236 2197 3995 2203
rect 4109 2197 4476 2203
rect 1293 2177 1516 2183
rect 1573 2177 2044 2183
rect 2148 2177 3356 2183
rect 3476 2177 3628 2183
rect 3652 2177 3820 2183
rect 4109 2183 4115 2197
rect 5117 2203 5123 2656
rect 5101 2197 5123 2203
rect 3876 2177 4115 2183
rect 4165 2177 4252 2183
rect 180 2157 1587 2163
rect 340 2137 428 2143
rect 484 2137 1564 2143
rect 1581 2143 1587 2157
rect 1605 2157 1628 2163
rect 1701 2157 1708 2163
rect 1829 2157 1980 2163
rect 2004 2157 2924 2163
rect 2948 2157 2971 2163
rect 3156 2157 3356 2163
rect 3461 2157 3708 2163
rect 3764 2157 4300 2163
rect 1581 2137 2395 2143
rect 2580 2137 3932 2143
rect 3988 2137 4348 2143
rect 4484 2137 4860 2143
rect 612 2117 668 2123
rect 1268 2117 1708 2123
rect 1716 2117 2188 2123
rect 2484 2117 2491 2123
rect 2501 2117 2876 2123
rect 2916 2117 3756 2123
rect 3828 2117 4092 2123
rect 4164 2117 4252 2123
rect 4452 2117 4540 2123
rect 4644 2117 4923 2123
rect 4933 2117 4972 2123
rect 1140 2097 1340 2103
rect 1381 2097 1388 2103
rect 1476 2097 1595 2103
rect 1620 2097 2748 2103
rect 2916 2097 3276 2103
rect 3749 2097 4444 2103
rect 4516 2097 4604 2103
rect 837 2077 1723 2083
rect 3293 2084 3299 2095
rect 1828 2077 2060 2083
rect 2212 2077 3148 2083
rect 3621 2077 3868 2083
rect 4676 2077 4923 2083
rect 852 2057 1612 2063
rect 1645 2057 2683 2063
rect 1645 2043 1651 2057
rect 2693 2057 3516 2063
rect 3524 2057 4380 2063
rect 836 2037 1651 2043
rect 837 2017 844 2023
rect 1268 2017 1275 2023
rect 1316 2017 1628 2023
rect 1645 2023 1651 2037
rect 1668 2037 1691 2043
rect 1733 2037 2140 2043
rect 2181 2037 2412 2043
rect 2437 2037 2444 2043
rect 2580 2037 2587 2043
rect 2629 2037 2684 2043
rect 2725 2037 2748 2043
rect 2804 2037 2811 2043
rect 2853 2037 2939 2043
rect 5101 2044 5107 2197
rect 3013 2037 3468 2043
rect 3780 2037 4476 2043
rect 1645 2017 1660 2023
rect 1732 2017 2028 2023
rect 2068 2017 2588 2023
rect 2596 2017 3276 2023
rect 3284 2017 3291 2023
rect 3476 2017 3916 2023
rect 3941 2017 4812 2023
rect 1172 1997 1499 2003
rect 2085 1997 2108 2003
rect 2148 1997 2171 2003
rect 2196 1997 2284 2003
rect 2301 1997 2651 2003
rect 773 1977 844 1983
rect 980 1977 1851 1983
rect 2301 1983 2307 1997
rect 2692 1997 2715 2003
rect 2756 1997 2843 2003
rect 3540 1997 3692 2003
rect 4004 1997 4492 2003
rect 5108 1997 5123 2003
rect 2276 1977 2307 1983
rect 2420 1977 3388 1983
rect 3412 1977 4108 1983
rect 4116 1977 5100 1983
rect 756 1957 859 1963
rect 869 1957 924 1963
rect 996 1957 1516 1963
rect 1605 1957 1659 1963
rect 1956 1957 2044 1963
rect 2245 1957 2396 1963
rect 2404 1957 2508 1963
rect 2772 1957 2844 1963
rect 2884 1957 2939 1963
rect 3077 1957 3195 1963
rect 3316 1957 4060 1963
rect 4916 1957 4956 1963
rect 5117 1963 5123 1997
rect 5101 1957 5123 1963
rect 453 1937 1436 1943
rect 1477 1937 1612 1943
rect 1636 1937 1756 1943
rect 1796 1937 2172 1943
rect 2213 1937 2444 1943
rect 2580 1937 2700 1943
rect 2725 1937 2995 1943
rect 676 1917 1052 1923
rect 1108 1917 1115 1923
rect 1172 1917 1308 1923
rect 1396 1917 1659 1923
rect 1748 1917 2523 1923
rect 2533 1917 2684 1923
rect 2756 1917 2972 1923
rect 2989 1923 2995 1937
rect 3204 1937 3340 1943
rect 3524 1937 4076 1943
rect 4301 1943 4307 1956
rect 4260 1937 4307 1943
rect 2989 1917 3580 1923
rect 3717 1917 3948 1923
rect 4004 1917 4620 1923
rect 1341 1904 1347 1915
rect 180 1897 924 1903
rect 1380 1897 1628 1903
rect 1700 1897 1964 1903
rect 2068 1897 2075 1903
rect 2100 1897 2588 1903
rect 2596 1897 2748 1903
rect 2772 1897 2811 1903
rect 2852 1897 3580 1903
rect 3621 1897 3628 1903
rect 3700 1897 4364 1903
rect 916 1877 1820 1883
rect 1861 1877 1996 1883
rect 2116 1877 2460 1883
rect 2533 1877 2555 1883
rect 2580 1877 2940 1883
rect 2981 1877 2988 1883
rect 3028 1877 3228 1883
rect 3396 1877 3515 1883
rect 3588 1877 3884 1883
rect 3892 1877 4076 1883
rect 4260 1877 4316 1883
rect 308 1857 844 1863
rect 964 1857 1388 1863
rect 1412 1857 1500 1863
rect 1556 1857 1595 1863
rect 1605 1857 1740 1863
rect 1828 1857 2572 1863
rect 2661 1857 2748 1863
rect 2765 1857 2811 1863
rect 1124 1837 1555 1843
rect 1189 1817 1260 1823
rect 1549 1824 1555 1837
rect 1604 1837 1644 1843
rect 1652 1837 2348 1843
rect 2373 1837 2444 1843
rect 2461 1825 2467 1836
rect 2765 1843 2771 1857
rect 2884 1857 2963 1863
rect 2565 1837 2771 1843
rect 2804 1837 2940 1843
rect 2957 1843 2963 1857
rect 2980 1857 3099 1863
rect 3124 1857 3292 1863
rect 3309 1857 3707 1863
rect 2957 1837 3020 1843
rect 3309 1843 3315 1857
rect 3732 1857 3739 1863
rect 3844 1857 3867 1863
rect 3972 1857 4275 1863
rect 3045 1837 3315 1843
rect 3332 1837 4108 1843
rect 4269 1843 4275 1857
rect 4269 1837 4316 1843
rect 1317 1817 1500 1823
rect 1765 1817 1851 1823
rect 1876 1817 1883 1823
rect 2116 1817 2331 1823
rect 2373 1817 2427 1823
rect 2708 1817 2860 1823
rect 2868 1817 3452 1823
rect 3460 1817 3980 1823
rect 4004 1817 4187 1823
rect 805 1797 844 1803
rect 1044 1797 1276 1803
rect 1380 1797 1596 1803
rect 1669 1797 1884 1803
rect 2181 1797 2380 1803
rect 2469 1797 2587 1803
rect 2701 1797 3340 1803
rect 468 1777 924 1783
rect 1061 1777 1116 1783
rect 1652 1777 1996 1783
rect 2148 1777 2235 1783
rect 2276 1777 2299 1783
rect 2388 1777 2491 1783
rect 324 1757 508 1763
rect 1445 1757 1676 1763
rect 1764 1757 1819 1763
rect 1892 1757 2267 1763
rect 2277 1757 2284 1763
rect 2317 1763 2323 1776
rect 2701 1783 2707 1797
rect 3357 1797 3740 1803
rect 2597 1777 2707 1783
rect 3357 1783 3363 1797
rect 3956 1797 4604 1803
rect 4773 1797 4860 1803
rect 2900 1777 3363 1783
rect 3373 1777 3628 1783
rect 2317 1757 2716 1763
rect 2804 1757 2860 1763
rect 2884 1757 2988 1763
rect 3373 1763 3379 1777
rect 3732 1777 3835 1783
rect 3972 1777 4124 1783
rect 4149 1777 4652 1783
rect 3012 1757 3379 1763
rect 3396 1757 3484 1763
rect 3524 1757 4044 1763
rect 4052 1757 4764 1763
rect 5101 1763 5107 1957
rect 5093 1757 5107 1763
rect 164 1737 1164 1743
rect 1285 1737 1388 1743
rect 1652 1737 1756 1743
rect 1957 1737 1980 1743
rect 2004 1737 2555 1743
rect 2628 1737 3068 1743
rect 3140 1737 3228 1743
rect 3621 1737 3836 1743
rect 3892 1737 3996 1743
rect 4068 1737 4140 1743
rect 4676 1737 4699 1743
rect 4869 1737 5091 1743
rect 1124 1717 1276 1723
rect 1796 1717 2491 1723
rect 2565 1717 2588 1723
rect 2596 1717 2796 1723
rect 5085 1724 5091 1737
rect 2853 1717 2908 1723
rect 2964 1717 3139 1723
rect 1236 1697 1243 1703
rect 1300 1697 1884 1703
rect 2004 1697 2139 1703
rect 2349 1697 2748 1703
rect 1556 1677 2011 1683
rect 2349 1683 2355 1697
rect 2868 1697 3020 1703
rect 3133 1703 3139 1717
rect 3156 1717 3724 1723
rect 3812 1717 4348 1723
rect 4372 1717 5004 1723
rect 3133 1697 4828 1703
rect 2260 1677 2355 1683
rect 2372 1677 2460 1683
rect 2501 1677 2876 1683
rect 2949 1677 2956 1683
rect 3028 1677 3547 1683
rect 3652 1677 4059 1683
rect 4100 1677 4155 1683
rect 4229 1677 4316 1683
rect 4324 1677 4380 1683
rect 477 1664 483 1675
rect 1277 1664 1283 1675
rect 1620 1657 2107 1663
rect 2148 1657 2651 1663
rect 2756 1657 2779 1663
rect 2821 1657 2988 1663
rect 3012 1657 4059 1663
rect 4173 1657 5004 1663
rect 1541 1637 1755 1643
rect 1765 1637 2300 1643
rect 2373 1637 2380 1643
rect 2404 1637 2491 1643
rect 2596 1637 2619 1643
rect 2772 1637 2860 1643
rect 2916 1637 3084 1643
rect 3124 1637 3372 1643
rect 4173 1643 4179 1657
rect 3429 1637 4179 1643
rect 4196 1637 4251 1643
rect 1716 1617 1723 1623
rect 1741 1617 1916 1623
rect 1741 1603 1747 1617
rect 2196 1617 2227 1623
rect 580 1597 1747 1603
rect 1764 1597 2204 1603
rect 2221 1603 2227 1617
rect 2245 1617 4220 1623
rect 2221 1597 2396 1603
rect 2420 1597 2779 1603
rect 2804 1597 3388 1603
rect 3461 1597 3515 1603
rect 3621 1597 3644 1603
rect 3812 1597 3931 1603
rect 4005 1597 4188 1603
rect 4388 1597 4636 1603
rect 4644 1597 4700 1603
rect 965 1577 1228 1583
rect 1652 1577 2579 1583
rect 388 1557 1036 1563
rect 1637 1557 1644 1563
rect 1796 1557 2363 1563
rect 2373 1557 2444 1563
rect 2477 1557 2508 1563
rect 612 1537 1788 1543
rect 1989 1537 2412 1543
rect 2477 1543 2483 1557
rect 2573 1563 2579 1577
rect 2756 1577 3244 1583
rect 3373 1577 3419 1583
rect 2573 1557 3148 1563
rect 3373 1563 3379 1577
rect 3453 1577 4828 1583
rect 3237 1557 3379 1563
rect 3453 1563 3459 1577
rect 3396 1557 3459 1563
rect 3988 1557 4019 1563
rect 2437 1537 2483 1543
rect 2501 1537 2587 1543
rect 2629 1537 2748 1543
rect 2789 1537 3091 1543
rect 1669 1517 1676 1523
rect 2021 1517 2284 1523
rect 2308 1517 2331 1523
rect 2372 1517 2427 1523
rect 2452 1517 2587 1523
rect 2789 1517 2988 1523
rect 3085 1523 3091 1537
rect 3109 1537 3132 1543
rect 3236 1537 3340 1543
rect 3492 1537 3996 1543
rect 4013 1543 4019 1557
rect 4420 1557 4435 1563
rect 4013 1537 4188 1543
rect 4429 1543 4435 1557
rect 4429 1537 4844 1543
rect 3085 1517 3227 1523
rect 3268 1517 3340 1523
rect 3461 1517 3484 1523
rect 3524 1517 3628 1523
rect 3653 1517 4091 1523
rect 4133 1517 4140 1523
rect 4276 1517 4844 1523
rect 5093 1517 5107 1523
rect 5101 1504 5107 1517
rect 244 1497 1308 1503
rect 1588 1497 1596 1503
rect 1604 1497 4268 1503
rect 484 1477 860 1483
rect 996 1477 1676 1483
rect 1764 1477 2011 1483
rect 2036 1477 2043 1483
rect 2117 1477 2811 1483
rect 2836 1477 3292 1483
rect 3332 1477 4828 1483
rect 308 1457 556 1463
rect 564 1457 988 1463
rect 1157 1457 1164 1463
rect 1221 1457 1884 1463
rect 2036 1457 2172 1463
rect 2196 1457 2572 1463
rect 2676 1457 2956 1463
rect 2980 1457 3212 1463
rect 3316 1457 4060 1463
rect 4101 1457 4108 1463
rect 4196 1457 4332 1463
rect 4420 1457 4716 1463
rect 4965 1457 4972 1463
rect 357 1437 364 1443
rect 1797 1437 1932 1443
rect 2053 1437 2236 1443
rect 2277 1437 2412 1443
rect 2437 1437 3148 1443
rect 3173 1437 3180 1443
rect 3348 1437 4268 1443
rect 4884 1437 5004 1443
rect 676 1417 2140 1423
rect 2196 1417 2652 1423
rect 2756 1417 2779 1423
rect 2868 1417 3643 1423
rect 3685 1417 4508 1423
rect 564 1397 1211 1403
rect 1252 1397 1516 1403
rect 1524 1397 1612 1403
rect 1652 1397 1852 1403
rect 2149 1397 2235 1403
rect 2308 1397 3004 1403
rect 3460 1397 4108 1403
rect 4340 1397 4572 1403
rect 84 1377 156 1383
rect 388 1377 492 1383
rect 1348 1377 1836 1383
rect 1908 1377 2396 1383
rect 2404 1377 4284 1383
rect 4452 1377 4556 1383
rect 4596 1377 4636 1383
rect 4660 1377 4828 1383
rect 132 1357 1500 1363
rect 1588 1357 1868 1363
rect 1925 1357 1947 1363
rect 2004 1357 2028 1363
rect 2116 1357 2172 1363
rect 2340 1357 2363 1363
rect 2452 1357 2492 1363
rect 2580 1357 2619 1363
rect 2629 1357 2892 1363
rect 2916 1357 2988 1363
rect 3013 1357 3195 1363
rect 3301 1357 3884 1363
rect 4052 1357 4059 1363
rect 4132 1357 4476 1363
rect 4532 1357 5148 1363
rect 676 1337 1868 1343
rect 1892 1337 2555 1343
rect 2565 1337 2604 1343
rect 2676 1337 2779 1343
rect 2804 1337 3067 1343
rect 3348 1337 3612 1343
rect 3781 1337 3836 1343
rect 3860 1337 5004 1343
rect 596 1317 700 1323
rect 1252 1317 1628 1323
rect 1844 1317 1964 1323
rect 1972 1317 2092 1323
rect 2100 1317 2140 1323
rect 2148 1317 2396 1323
rect 2437 1317 3675 1323
rect 3716 1317 4412 1323
rect 4420 1317 4443 1323
rect 4516 1317 4764 1323
rect 4869 1317 4876 1323
rect 1348 1297 2139 1303
rect 2164 1297 2572 1303
rect 2597 1297 2604 1303
rect 2740 1297 2828 1303
rect 2853 1297 3004 1303
rect 3012 1297 3035 1303
rect 3077 1297 3356 1303
rect 3380 1297 3771 1303
rect 3796 1297 4124 1303
rect 4148 1297 4443 1303
rect 4677 1297 5068 1303
rect 749 1277 763 1283
rect 749 1243 755 1277
rect 1012 1277 1068 1283
rect 1076 1277 1804 1283
rect 1892 1277 2428 1283
rect 2477 1277 4444 1283
rect 773 1257 1132 1263
rect 1156 1257 2011 1263
rect 2052 1257 2140 1263
rect 2477 1263 2483 1277
rect 4805 1277 4876 1283
rect 2245 1257 2483 1263
rect 2500 1257 2523 1263
rect 2533 1257 2587 1263
rect 2605 1257 2876 1263
rect 749 1237 764 1243
rect 1972 1237 2396 1243
rect 2413 1237 2427 1243
rect 1140 1217 1420 1223
rect 1956 1217 2300 1223
rect 2413 1223 2419 1237
rect 2493 1225 2499 1236
rect 2605 1243 2611 1257
rect 2949 1257 3003 1263
rect 3108 1257 3804 1263
rect 3828 1257 4428 1263
rect 4453 1257 4828 1263
rect 2565 1237 2611 1243
rect 2756 1237 3596 1243
rect 3636 1237 4332 1243
rect 4532 1237 4539 1243
rect 2404 1217 2419 1223
rect 2629 1217 2636 1223
rect 2789 1217 2796 1223
rect 2821 1217 3611 1223
rect 3781 1217 3788 1223
rect 3877 1217 3916 1223
rect 3988 1217 4220 1223
rect 1492 1197 1612 1203
rect 1956 1197 1980 1203
rect 2429 1204 2435 1215
rect 2021 1197 2316 1203
rect 2500 1197 3372 1203
rect 3396 1197 3740 1203
rect 3860 1197 4364 1203
rect 820 1177 1339 1183
rect 1669 1177 2235 1183
rect 2292 1177 2396 1183
rect 2436 1177 3100 1183
rect 3301 1177 4268 1183
rect 1125 1157 1212 1163
rect 1876 1157 2060 1163
rect 2068 1157 2715 1163
rect 2740 1157 3308 1163
rect 3332 1157 3788 1163
rect 3796 1157 3996 1163
rect 4197 1157 4667 1163
rect 1061 1137 1420 1143
rect 1652 1137 1659 1143
rect 1748 1137 2171 1143
rect 2244 1137 2348 1143
rect 2356 1137 2427 1143
rect 2629 1137 2764 1143
rect 2836 1137 2939 1143
rect 2964 1137 3564 1143
rect 3636 1137 3804 1143
rect 3844 1137 4604 1143
rect 212 1117 412 1123
rect 420 1117 1708 1123
rect 1924 1117 2067 1123
rect 660 1097 1187 1103
rect 996 1077 1147 1083
rect 1181 1083 1187 1097
rect 1205 1097 1723 1103
rect 1733 1097 2043 1103
rect 2061 1103 2067 1117
rect 2116 1117 2491 1123
rect 2724 1117 2972 1123
rect 3012 1117 3291 1123
rect 3716 1117 3980 1123
rect 3988 1117 3995 1123
rect 4308 1117 4412 1123
rect 4901 1117 5068 1123
rect 2061 1097 2108 1103
rect 2181 1097 2267 1103
rect 2292 1097 2523 1103
rect 2564 1097 2876 1103
rect 2884 1097 3724 1103
rect 3924 1097 4219 1103
rect 4260 1097 4556 1103
rect 4564 1097 4796 1103
rect 1181 1077 1804 1083
rect 2053 1077 2076 1083
rect 2180 1077 2556 1083
rect 2596 1077 2939 1083
rect 3012 1077 3180 1083
rect 3236 1077 3276 1083
rect 3364 1077 3900 1083
rect 4228 1077 4572 1083
rect 4805 1077 4844 1083
rect 996 1057 1019 1063
rect 1029 1057 1132 1063
rect 1149 1057 1164 1063
rect 916 1037 1051 1043
rect 1149 1043 1155 1057
rect 1172 1057 1563 1063
rect 1684 1057 2444 1063
rect 2533 1057 2636 1063
rect 2756 1057 3116 1063
rect 3444 1057 3451 1063
rect 3524 1057 3699 1063
rect 1140 1037 1155 1043
rect 1165 1037 1676 1043
rect 1165 1023 1171 1037
rect 1860 1037 2011 1043
rect 3693 1044 3699 1057
rect 4165 1057 4284 1063
rect 4756 1057 4988 1063
rect 5189 1057 5196 1063
rect 2052 1037 2316 1043
rect 2388 1037 3068 1043
rect 3076 1037 3628 1043
rect 3813 1037 3820 1043
rect 4148 1037 4155 1043
rect 228 1017 1171 1023
rect 1508 1017 3004 1023
rect 3380 1017 3484 1023
rect 3653 1017 4636 1023
rect 4740 1017 4764 1023
rect 1637 997 1644 1003
rect 2021 997 2588 1003
rect 2644 997 2732 1003
rect 2789 997 2796 1003
rect 2949 997 3180 1003
rect 3572 997 3852 1003
rect 3973 997 4732 1003
rect 5044 997 5051 1003
rect 260 977 300 983
rect 500 977 1699 983
rect 132 957 1468 963
rect 1588 957 1676 963
rect 1693 963 1699 977
rect 1956 977 3708 983
rect 3812 977 3819 983
rect 3844 977 3916 983
rect 3988 977 4892 983
rect 1693 957 2044 963
rect 2180 957 2300 963
rect 2324 957 2396 963
rect 2501 957 2652 963
rect 2429 945 2435 956
rect 2693 957 2732 963
rect 2804 957 2811 963
rect 2868 957 3612 963
rect 3636 957 3643 963
rect 3732 957 4140 963
rect 4388 957 4492 963
rect 4948 957 5100 963
rect 116 937 300 943
rect 436 937 443 943
rect 453 937 764 943
rect 964 937 1148 943
rect 1172 937 1811 943
rect 356 917 524 923
rect 532 917 1468 923
rect 1637 917 1740 923
rect 1805 923 1811 937
rect 2085 937 2380 943
rect 2469 937 2508 943
rect 2725 937 2828 943
rect 2884 937 2956 943
rect 3380 937 3484 943
rect 3716 937 4460 943
rect 1805 917 2140 923
rect 2244 917 2428 923
rect 2436 917 2556 923
rect 2564 917 2732 923
rect 2836 917 3180 923
rect 3188 917 4188 923
rect 4420 917 4524 923
rect 1220 897 1228 903
rect 1236 897 1836 903
rect 1892 897 2075 903
rect 2260 897 2267 903
rect 2277 897 2892 903
rect 2964 897 2971 903
rect 3140 897 3515 903
rect 3652 897 4060 903
rect 4340 897 5180 903
rect 1284 877 1308 883
rect 1396 877 1468 883
rect 1476 877 2748 883
rect 2948 877 3308 883
rect 3556 877 3788 883
rect 3892 877 3931 883
rect 3956 877 3963 883
rect 4196 877 4955 883
rect 772 857 1404 863
rect 1684 857 3228 863
rect 3732 857 3884 863
rect 1172 837 1740 843
rect 2085 837 2715 843
rect 3012 837 4748 843
rect 4756 837 5084 843
rect 2781 825 2787 836
rect 1364 817 1659 823
rect 2117 817 2172 823
rect 2245 817 2619 823
rect 2804 817 3036 823
rect 3076 817 4108 823
rect 1172 797 1948 803
rect 1956 797 2156 803
rect 2244 797 2492 803
rect 2564 797 3011 803
rect 452 777 1915 783
rect 1940 777 2107 783
rect 2148 777 2748 783
rect 3005 783 3011 797
rect 3028 797 3035 803
rect 3092 797 3228 803
rect 4052 797 4059 803
rect 4077 797 4220 803
rect 3005 777 3180 783
rect 3268 777 3292 783
rect 3781 777 3820 783
rect 4077 783 4083 797
rect 3956 777 4083 783
rect 4101 777 5036 783
rect 5172 777 5179 783
rect 1924 757 2188 763
rect 2228 757 2555 763
rect 1789 745 1795 756
rect 2597 757 2732 763
rect 2789 757 3868 763
rect 3940 757 4044 763
rect 4133 757 4140 763
rect 292 737 780 743
rect 1925 737 2172 743
rect 2213 737 2412 743
rect 2436 737 2492 743
rect 2660 737 2747 743
rect 2804 737 3452 743
rect 3589 737 3980 743
rect 4004 737 4508 743
rect 4644 737 4795 743
rect 84 717 524 723
rect 564 717 571 723
rect 1524 717 2931 723
rect 1156 697 1324 703
rect 1572 697 2907 703
rect 2925 703 2931 717
rect 3060 717 3740 723
rect 3781 717 3996 723
rect 4020 717 4412 723
rect 2925 697 3587 703
rect 660 677 667 683
rect 1412 677 1532 683
rect 1684 677 1804 683
rect 1812 677 1980 683
rect 2021 677 2331 683
rect 2372 677 2412 683
rect 2436 677 2716 683
rect 2788 677 2860 683
rect 2916 677 3564 683
rect 3581 683 3587 697
rect 3732 697 3836 703
rect 3908 697 3948 703
rect 3988 697 4028 703
rect 4052 697 4076 703
rect 4148 697 5100 703
rect 3581 677 3771 683
rect 3844 677 4140 683
rect 4500 677 4636 683
rect 293 657 316 663
rect 1060 657 1788 663
rect 1821 657 1980 663
rect 196 637 371 643
rect 365 623 371 637
rect 1012 637 1084 643
rect 1332 637 1724 643
rect 1821 643 1827 657
rect 1988 657 2076 663
rect 2244 657 2380 663
rect 2533 657 2796 663
rect 2868 657 2875 663
rect 3213 657 3355 663
rect 1732 637 1827 643
rect 1844 637 1916 643
rect 1924 637 2044 643
rect 2148 637 2748 643
rect 3213 643 3219 657
rect 3380 657 3451 663
rect 3476 657 4156 663
rect 4452 657 5036 663
rect 2885 637 3219 643
rect 3236 637 3483 643
rect 3524 637 4540 643
rect 5012 637 5132 643
rect 365 617 1004 623
rect 1108 617 1196 623
rect 1316 617 2268 623
rect 2372 617 2476 623
rect 2644 617 2940 623
rect 2996 617 3180 623
rect 3252 617 3259 623
rect 3365 617 3419 623
rect 3444 617 3516 623
rect 3909 617 3916 623
rect 4020 617 4140 623
rect 4157 617 4220 623
rect 452 597 540 603
rect 788 597 795 603
rect 948 597 1100 603
rect 1652 597 2268 603
rect 2309 597 2316 603
rect 2341 597 2412 603
rect 2484 597 2572 603
rect 2597 597 3228 603
rect 3429 597 3436 603
rect 3460 597 4028 603
rect 4084 597 4091 603
rect 4157 603 4163 617
rect 4517 617 4796 623
rect 4116 597 4163 603
rect 4180 597 4187 603
rect 4709 597 5132 603
rect 132 577 1148 583
rect 1220 577 1404 583
rect 1940 577 2476 583
rect 2500 577 2523 583
rect 1693 565 1699 576
rect 2564 577 2843 583
rect 2916 577 3420 583
rect 3700 577 4924 583
rect 581 557 748 563
rect 772 557 892 563
rect 948 557 1084 563
rect 1108 557 1660 563
rect 1765 557 1788 563
rect 1829 557 2011 563
rect 2084 557 2284 563
rect 2324 557 3180 563
rect 3188 557 3964 563
rect 4052 557 4123 563
rect 4148 557 4507 563
rect 4548 557 4684 563
rect 5076 557 5083 563
rect 180 537 1324 543
rect 1604 537 1724 543
rect 1956 537 2300 543
rect 2468 537 3660 543
rect 3700 537 4188 543
rect 4196 537 4796 543
rect 4884 537 5116 543
rect 516 517 780 523
rect 805 517 1356 523
rect 1540 517 2796 523
rect 2820 517 3884 523
rect 3908 517 4604 523
rect 1460 497 1980 503
rect 2116 497 2188 503
rect 2196 497 2220 503
rect 2228 497 2476 503
rect 2484 497 2556 503
rect 2788 497 2860 503
rect 3076 497 3372 503
rect 3461 497 3779 503
rect 644 477 1932 483
rect 2340 477 2587 483
rect 2948 477 3100 483
rect 3300 477 3724 483
rect 3773 483 3779 497
rect 3796 497 3948 503
rect 4036 497 4636 503
rect 3773 477 4012 483
rect 4037 477 4428 483
rect 900 457 1660 463
rect 1988 457 2124 463
rect 2244 457 2267 463
rect 2292 457 2316 463
rect 2341 457 2875 463
rect 2900 457 3052 463
rect 3060 457 4059 463
rect 1876 437 2811 443
rect 1380 417 2380 423
rect 2388 417 4076 423
rect 1396 397 2012 403
rect 2245 397 2460 403
rect 2629 397 2636 403
rect 2724 397 2907 403
rect 2932 397 3084 403
rect 3109 397 4172 403
rect 1412 377 1563 383
rect 1588 377 1660 383
rect 1685 377 1836 383
rect 1861 377 1868 383
rect 2004 377 2380 383
rect 2405 377 3836 383
rect 420 357 3116 363
rect 3236 357 3996 363
rect 741 337 908 343
rect 948 337 955 343
rect 1061 337 1100 343
rect 1252 337 2076 343
rect 2084 337 3468 343
rect 3493 337 3948 343
rect 4244 337 4636 343
rect 260 317 380 323
rect 756 317 860 323
rect 884 317 2171 323
rect 2196 317 2636 323
rect 2661 317 2812 323
rect 2868 317 2971 323
rect 3012 317 3164 323
rect 3188 317 3500 323
rect 3812 317 4124 323
rect 436 297 1724 303
rect 1748 297 1804 303
rect 2068 297 2172 303
rect 2532 297 2540 303
rect 2548 297 3036 303
rect 3092 297 3980 303
rect 404 277 476 283
rect 628 277 1660 283
rect 1700 277 2252 283
rect 2388 277 2588 283
rect 2629 277 2860 283
rect 2932 277 2939 283
rect 3045 277 3244 283
rect 3268 277 3356 283
rect 3380 277 3612 283
rect 3828 277 3884 283
rect 4069 277 4172 283
rect 4660 277 4780 283
rect 4837 277 5132 283
rect 772 257 1228 263
rect 1252 257 1356 263
rect 1381 257 1468 263
rect 1636 257 1787 263
rect 1956 257 1979 263
rect 2004 257 2252 263
rect 2404 257 2460 263
rect 2516 257 2635 263
rect 2660 257 3500 263
rect 3796 257 3851 263
rect 3876 257 4315 263
rect 4869 257 5068 263
rect 740 237 1884 243
rect 1892 237 1980 243
rect 2021 237 2060 243
rect 2181 237 2716 243
rect 2740 237 2812 243
rect 2868 237 2924 243
rect 2948 237 3132 243
rect 3173 237 3420 243
rect 3444 237 3852 243
rect 3877 237 3900 243
rect 3924 237 3931 243
rect 708 217 972 223
rect 1268 217 1275 223
rect 1780 217 3228 223
rect 3668 217 4204 223
rect 4308 217 4412 223
rect 4788 217 4844 223
rect 1140 197 3804 203
rect 4100 197 4332 203
rect 301 177 748 183
rect 301 163 307 177
rect 1172 177 1196 183
rect 1364 177 2044 183
rect 2116 177 2395 183
rect 2420 177 2812 183
rect 2820 177 2876 183
rect 2900 177 3115 183
rect 3140 177 4140 183
rect 4165 177 4524 183
rect 4788 177 5068 183
rect 132 157 307 163
rect 356 157 460 163
rect 708 157 908 163
rect 1556 157 1628 163
rect 1668 157 2572 163
rect 2597 157 2860 163
rect 2885 157 2924 163
rect 2932 157 2939 163
rect 2964 157 3548 163
rect 3588 157 3683 163
rect 452 137 699 143
rect 285 125 291 136
rect 724 137 844 143
rect 852 137 876 143
rect 1076 137 2508 143
rect 2516 137 3148 143
rect 3204 137 3596 143
rect 3621 137 3628 143
rect 3677 143 3683 157
rect 3700 157 4828 163
rect 5125 157 5164 163
rect 3677 137 3771 143
rect 3796 137 4988 143
rect 293 117 716 123
rect 741 117 940 123
rect 964 117 1356 123
rect 1684 117 2028 123
rect 2212 117 2444 123
rect 2628 117 3388 123
rect 3476 117 3980 123
rect 4068 117 4156 123
rect 4212 117 4540 123
rect 532 97 1804 103
rect 1876 97 2012 103
rect 2821 97 3132 103
rect 628 77 956 83
rect 2564 77 2875 83
rect 2916 77 3100 83
rect 3141 77 3164 83
rect 932 57 3196 63
rect 1748 37 3340 43
rect 2004 17 2492 23
rect 2500 17 3404 23
<< m6contact >>
rect 3659 3535 3669 3545
rect 3515 3524 3525 3525
rect 3515 3516 3516 3524
rect 3516 3516 3524 3524
rect 3524 3516 3525 3524
rect 3515 3515 3525 3516
rect 3611 3495 3621 3505
rect 2475 3455 2485 3465
rect 4811 3455 4821 3465
rect 2235 3435 2245 3445
rect 2395 3435 2405 3445
rect 2523 3435 2533 3445
rect 4443 3435 4453 3445
rect 4859 3435 4869 3445
rect 2715 3415 2725 3425
rect 3195 3415 3205 3425
rect 3483 3415 3493 3425
rect 3035 3395 3045 3405
rect 3131 3395 3141 3405
rect 1723 3384 1733 3385
rect 3227 3384 3237 3385
rect 1723 3376 1724 3384
rect 1724 3376 1732 3384
rect 1732 3376 1733 3384
rect 1723 3375 1733 3376
rect 3035 3355 3045 3365
rect 3067 3355 3077 3365
rect 3227 3376 3228 3384
rect 3228 3376 3236 3384
rect 3236 3376 3237 3384
rect 3227 3375 3237 3376
rect 3323 3384 3333 3385
rect 3323 3376 3324 3384
rect 3324 3376 3332 3384
rect 3332 3376 3333 3384
rect 3387 3395 3397 3405
rect 3707 3395 3717 3405
rect 3323 3375 3333 3376
rect 3579 3375 3589 3385
rect 3659 3375 3669 3385
rect 3819 3375 3829 3385
rect 4027 3355 4037 3365
rect 5115 3364 5125 3365
rect 5115 3356 5116 3364
rect 5116 3356 5124 3364
rect 5124 3356 5125 3364
rect 5115 3355 5125 3356
rect 1115 3344 1125 3345
rect 1115 3336 1116 3344
rect 1116 3336 1124 3344
rect 1124 3336 1125 3344
rect 1115 3335 1125 3336
rect 1851 3335 1861 3345
rect 1883 3335 1893 3345
rect 827 3315 837 3325
rect 4923 3335 4933 3345
rect 2523 3315 2533 3325
rect 4891 3315 4901 3325
rect 3131 3295 3141 3305
rect 3419 3295 3429 3305
rect 4251 3295 4261 3305
rect 3067 3255 3077 3265
rect 763 3235 773 3245
rect 1851 3235 1861 3245
rect 1595 3195 1605 3205
rect 2683 3175 2693 3185
rect 1307 3164 1317 3165
rect 1307 3156 1308 3164
rect 1308 3156 1316 3164
rect 1316 3156 1317 3164
rect 1307 3155 1317 3156
rect 1371 3155 1381 3165
rect 891 3144 901 3145
rect 891 3136 892 3144
rect 892 3136 900 3144
rect 900 3136 901 3144
rect 1691 3144 1701 3145
rect 1691 3136 1692 3144
rect 1692 3136 1700 3144
rect 1700 3136 1701 3144
rect 891 3135 901 3136
rect 1691 3135 1701 3136
rect 1755 3135 1765 3145
rect 1659 3115 1669 3125
rect 3067 3115 3077 3125
rect 4763 3115 4773 3125
rect 1755 3095 1765 3105
rect 3547 3055 3557 3065
rect 1435 3035 1445 3045
rect 2491 3035 2501 3045
rect 3067 3035 3077 3045
rect 2075 2995 2085 3005
rect 2171 2995 2181 3005
rect 3131 2975 3141 2985
rect 2411 2935 2421 2945
rect 1179 2895 1189 2905
rect 1243 2895 1253 2905
rect 1371 2915 1381 2925
rect 1723 2915 1733 2925
rect 2203 2915 2213 2925
rect 2459 2915 2469 2925
rect 2491 2915 2501 2925
rect 3099 2915 3109 2925
rect 3323 2924 3333 2925
rect 3323 2916 3324 2924
rect 3324 2916 3332 2924
rect 3332 2916 3333 2924
rect 3323 2915 3333 2916
rect 5147 2895 5157 2905
rect 1051 2875 1061 2885
rect 1435 2875 1445 2885
rect 1723 2875 1733 2885
rect 1915 2875 1925 2885
rect 3451 2875 3461 2885
rect 795 2855 805 2865
rect 1883 2835 1893 2845
rect 2043 2815 2053 2825
rect 2075 2824 2085 2825
rect 2075 2816 2076 2824
rect 2076 2816 2084 2824
rect 2084 2816 2085 2824
rect 2075 2815 2085 2816
rect 2235 2795 2245 2805
rect 2363 2775 2373 2785
rect 763 2755 773 2765
rect 3291 2755 3301 2765
rect 4507 2755 4517 2765
rect 475 2735 485 2745
rect 2683 2735 2693 2745
rect 2939 2735 2949 2745
rect 2043 2715 2053 2725
rect 3131 2724 3141 2725
rect 3131 2716 3132 2724
rect 3132 2716 3140 2724
rect 3140 2716 3141 2724
rect 4315 2735 4325 2745
rect 4827 2735 4837 2745
rect 3131 2715 3141 2716
rect 3515 2715 3525 2725
rect 5083 2715 5093 2725
rect 1499 2695 1509 2705
rect 2267 2695 2277 2705
rect 1531 2675 1541 2685
rect 2235 2675 2245 2685
rect 475 2655 485 2665
rect 955 2655 965 2665
rect 1851 2655 1861 2665
rect 5051 2655 5061 2665
rect 1467 2635 1477 2645
rect 1499 2635 1509 2645
rect 1531 2635 1541 2645
rect 2299 2635 2309 2645
rect 3835 2635 3845 2645
rect 3995 2635 4005 2645
rect 4155 2635 4165 2645
rect 4187 2635 4197 2645
rect 2459 2615 2469 2625
rect 2491 2615 2501 2625
rect 795 2575 805 2585
rect 3867 2595 3877 2605
rect 1563 2584 1573 2585
rect 1563 2576 1564 2584
rect 1564 2576 1572 2584
rect 1572 2576 1573 2584
rect 1563 2575 1573 2576
rect 1755 2575 1765 2585
rect 923 2555 933 2565
rect 1435 2555 1445 2565
rect 1467 2555 1477 2565
rect 2587 2555 2597 2565
rect 2747 2564 2757 2565
rect 2747 2556 2748 2564
rect 2748 2556 2756 2564
rect 2756 2556 2757 2564
rect 2747 2555 2757 2556
rect 3067 2555 3077 2565
rect 443 2544 453 2545
rect 443 2536 444 2544
rect 444 2536 452 2544
rect 452 2536 453 2544
rect 443 2535 453 2536
rect 891 2535 901 2545
rect 2011 2535 2021 2545
rect 2843 2535 2853 2545
rect 795 2515 805 2525
rect 2491 2515 2501 2525
rect 2587 2515 2597 2525
rect 4187 2515 4197 2525
rect 4251 2515 4261 2525
rect 2555 2495 2565 2505
rect 2651 2495 2661 2505
rect 2875 2495 2885 2505
rect 2971 2495 2981 2505
rect 3003 2495 3013 2505
rect 3131 2495 3141 2505
rect 3899 2495 3909 2505
rect 1627 2475 1637 2485
rect 1275 2455 1285 2465
rect 1531 2444 1541 2445
rect 1531 2436 1532 2444
rect 1532 2436 1540 2444
rect 1540 2436 1541 2444
rect 1531 2435 1541 2436
rect 1563 2444 1573 2445
rect 1563 2436 1564 2444
rect 1564 2436 1572 2444
rect 1572 2436 1573 2444
rect 1563 2435 1573 2436
rect 1595 2435 1605 2445
rect 2459 2455 2469 2465
rect 2779 2475 2789 2485
rect 2843 2455 2853 2465
rect 2907 2475 2917 2485
rect 3739 2475 3749 2485
rect 4507 2475 4517 2485
rect 2971 2455 2981 2465
rect 3003 2455 3013 2465
rect 3131 2464 3141 2465
rect 3131 2456 3132 2464
rect 3132 2456 3140 2464
rect 3140 2456 3141 2464
rect 3131 2455 3141 2456
rect 3291 2455 3301 2465
rect 2811 2435 2821 2445
rect 4283 2435 4293 2445
rect 1883 2415 1893 2425
rect 1915 2415 1925 2425
rect 2779 2415 2789 2425
rect 4027 2415 4037 2425
rect 1275 2395 1285 2405
rect 4059 2395 4069 2405
rect 3099 2375 3109 2385
rect 4091 2375 4101 2385
rect 4699 2375 4709 2385
rect 1115 2335 1125 2345
rect 3995 2335 4005 2345
rect 1499 2315 1509 2325
rect 2779 2315 2789 2325
rect 3003 2315 3013 2325
rect 3483 2324 3493 2325
rect 3483 2316 3484 2324
rect 3484 2316 3492 2324
rect 3492 2316 3493 2324
rect 3483 2315 3493 2316
rect 2427 2295 2437 2305
rect 347 2255 357 2265
rect 475 2255 485 2265
rect 827 2255 837 2265
rect 859 2255 869 2265
rect 1723 2255 1733 2265
rect 1755 2264 1765 2265
rect 1755 2256 1756 2264
rect 1756 2256 1764 2264
rect 1764 2256 1765 2264
rect 1755 2255 1765 2256
rect 1787 2264 1797 2265
rect 1787 2256 1788 2264
rect 1788 2256 1796 2264
rect 1796 2256 1797 2264
rect 1787 2255 1797 2256
rect 1979 2255 1989 2265
rect 3771 2255 3781 2265
rect 3883 2255 3893 2265
rect 3963 2255 3973 2265
rect 667 2244 677 2245
rect 667 2236 668 2244
rect 668 2236 676 2244
rect 676 2236 677 2244
rect 667 2235 677 2236
rect 2619 2235 2629 2245
rect 283 2224 293 2225
rect 283 2216 284 2224
rect 284 2216 292 2224
rect 292 2216 293 2224
rect 283 2215 293 2216
rect 859 2215 869 2225
rect 1819 2215 1829 2225
rect 1883 2215 1893 2225
rect 2651 2215 2661 2225
rect 2843 2215 2853 2225
rect 3771 2215 3781 2225
rect 3803 2215 3813 2225
rect 3963 2215 3973 2225
rect 4795 2235 4805 2245
rect 283 2175 293 2185
rect 731 2175 741 2185
rect 1275 2175 1285 2185
rect 1467 2195 1477 2205
rect 2971 2195 2981 2205
rect 3995 2195 4005 2205
rect 4091 2195 4101 2205
rect 1563 2184 1573 2185
rect 1563 2176 1564 2184
rect 1564 2176 1572 2184
rect 1572 2176 1573 2184
rect 4123 2184 4133 2185
rect 4123 2176 4124 2184
rect 4124 2176 4132 2184
rect 4132 2176 4133 2184
rect 1563 2175 1573 2176
rect 4123 2175 4133 2176
rect 4155 2175 4165 2185
rect 1595 2155 1605 2165
rect 1691 2155 1701 2165
rect 1819 2155 1829 2165
rect 2971 2155 2981 2165
rect 3131 2164 3141 2165
rect 3131 2156 3132 2164
rect 3132 2156 3140 2164
rect 3140 2156 3141 2164
rect 3131 2155 3141 2156
rect 3451 2155 3461 2165
rect 2395 2144 2405 2145
rect 2395 2136 2396 2144
rect 2396 2136 2404 2144
rect 2404 2136 2405 2144
rect 2395 2135 2405 2136
rect 2491 2115 2501 2125
rect 4923 2115 4933 2125
rect 1371 2095 1381 2105
rect 1595 2095 1605 2105
rect 2843 2104 2853 2105
rect 2843 2096 2844 2104
rect 2844 2096 2852 2104
rect 2852 2096 2853 2104
rect 2843 2095 2853 2096
rect 3291 2095 3301 2105
rect 3579 2104 3589 2105
rect 3579 2096 3580 2104
rect 3580 2096 3588 2104
rect 3588 2096 3589 2104
rect 3579 2095 3589 2096
rect 3739 2095 3749 2105
rect 827 2075 837 2085
rect 1723 2075 1733 2085
rect 3451 2084 3461 2085
rect 3451 2076 3452 2084
rect 3452 2076 3460 2084
rect 3460 2076 3461 2084
rect 3451 2075 3461 2076
rect 3611 2075 3621 2085
rect 4923 2075 4933 2085
rect 2683 2055 2693 2065
rect 827 2015 837 2025
rect 1275 2015 1285 2025
rect 1691 2035 1701 2045
rect 1723 2035 1733 2045
rect 2171 2035 2181 2045
rect 2427 2035 2437 2045
rect 2587 2035 2597 2045
rect 2619 2035 2629 2045
rect 2715 2035 2725 2045
rect 2811 2035 2821 2045
rect 2843 2035 2853 2045
rect 2939 2035 2949 2045
rect 3003 2035 3013 2045
rect 3291 2015 3301 2025
rect 3931 2015 3941 2025
rect 1499 1995 1509 2005
rect 2075 1995 2085 2005
rect 2171 1995 2181 2005
rect 763 1975 773 1985
rect 1851 1975 1861 1985
rect 2171 1984 2181 1985
rect 2171 1976 2172 1984
rect 2172 1976 2180 1984
rect 2180 1976 2181 1984
rect 2651 1995 2661 2005
rect 2715 1995 2725 2005
rect 2843 1995 2853 2005
rect 2171 1975 2181 1976
rect 859 1955 869 1965
rect 1595 1955 1605 1965
rect 1659 1955 1669 1965
rect 2235 1955 2245 1965
rect 2939 1955 2949 1965
rect 3067 1955 3077 1965
rect 3195 1955 3205 1965
rect 443 1935 453 1945
rect 1467 1935 1477 1945
rect 2203 1935 2213 1945
rect 2715 1935 2725 1945
rect 1115 1915 1125 1925
rect 1339 1915 1349 1925
rect 1659 1915 1669 1925
rect 2523 1915 2533 1925
rect 3707 1915 3717 1925
rect 1019 1904 1029 1905
rect 1019 1896 1020 1904
rect 1020 1896 1028 1904
rect 1028 1896 1029 1904
rect 1019 1895 1029 1896
rect 2075 1895 2085 1905
rect 2811 1895 2821 1905
rect 3611 1895 3621 1905
rect 1851 1875 1861 1885
rect 2523 1875 2533 1885
rect 2555 1875 2565 1885
rect 2971 1875 2981 1885
rect 3003 1884 3013 1885
rect 3003 1876 3004 1884
rect 3004 1876 3012 1884
rect 3012 1876 3013 1884
rect 3003 1875 3013 1876
rect 3515 1875 3525 1885
rect 1595 1855 1605 1865
rect 2651 1855 2661 1865
rect 1179 1815 1189 1825
rect 1307 1815 1317 1825
rect 2363 1835 2373 1845
rect 2555 1835 2565 1845
rect 2811 1855 2821 1865
rect 3099 1855 3109 1865
rect 3035 1835 3045 1845
rect 3707 1855 3717 1865
rect 3739 1855 3749 1865
rect 3867 1855 3877 1865
rect 4283 1864 4293 1865
rect 4283 1856 4284 1864
rect 4284 1856 4292 1864
rect 4292 1856 4293 1864
rect 4283 1855 4293 1856
rect 1755 1815 1765 1825
rect 1851 1815 1861 1825
rect 1883 1815 1893 1825
rect 2331 1815 2341 1825
rect 2363 1815 2373 1825
rect 2427 1815 2437 1825
rect 2459 1815 2469 1825
rect 4187 1815 4197 1825
rect 4795 1824 4805 1825
rect 4795 1816 4796 1824
rect 4796 1816 4804 1824
rect 4804 1816 4805 1824
rect 4795 1815 4805 1816
rect 4859 1824 4869 1825
rect 4859 1816 4860 1824
rect 4860 1816 4868 1824
rect 4868 1816 4869 1824
rect 4859 1815 4869 1816
rect 795 1795 805 1805
rect 1659 1795 1669 1805
rect 2171 1795 2181 1805
rect 2459 1795 2469 1805
rect 2587 1795 2597 1805
rect 1051 1775 1061 1785
rect 2235 1775 2245 1785
rect 2299 1775 2309 1785
rect 923 1764 933 1765
rect 923 1756 924 1764
rect 924 1756 932 1764
rect 932 1756 933 1764
rect 923 1755 933 1756
rect 1435 1755 1445 1765
rect 1819 1755 1829 1765
rect 2267 1755 2277 1765
rect 2491 1775 2501 1785
rect 2587 1775 2597 1785
rect 2715 1784 2725 1785
rect 2715 1776 2716 1784
rect 2716 1776 2724 1784
rect 2724 1776 2725 1784
rect 4763 1795 4773 1805
rect 2715 1775 2725 1776
rect 3835 1775 3845 1785
rect 4139 1775 4149 1785
rect 5083 1784 5093 1785
rect 5083 1776 5084 1784
rect 5084 1776 5092 1784
rect 5092 1776 5093 1784
rect 5083 1775 5093 1776
rect 5083 1755 5093 1765
rect 1275 1735 1285 1745
rect 1947 1735 1957 1745
rect 2555 1735 2565 1745
rect 3579 1744 3589 1745
rect 3579 1736 3580 1744
rect 3580 1736 3588 1744
rect 3588 1736 3589 1744
rect 3579 1735 3589 1736
rect 3611 1735 3621 1745
rect 4699 1735 4709 1745
rect 4859 1735 4869 1745
rect 2491 1715 2501 1725
rect 2555 1715 2565 1725
rect 2843 1715 2853 1725
rect 1243 1695 1253 1705
rect 2139 1695 2149 1705
rect 475 1675 485 1685
rect 1275 1675 1285 1685
rect 2011 1675 2021 1685
rect 2491 1675 2501 1685
rect 2939 1675 2949 1685
rect 3547 1675 3557 1685
rect 4059 1675 4069 1685
rect 4155 1675 4165 1685
rect 4219 1675 4229 1685
rect 2107 1655 2117 1665
rect 2651 1655 2661 1665
rect 2779 1655 2789 1665
rect 2811 1655 2821 1665
rect 4059 1655 4069 1665
rect 1531 1635 1541 1645
rect 1755 1635 1765 1645
rect 2363 1635 2373 1645
rect 2491 1635 2501 1645
rect 2619 1635 2629 1645
rect 3419 1635 3429 1645
rect 4251 1635 4261 1645
rect 1723 1615 1733 1625
rect 2139 1624 2149 1625
rect 2139 1616 2140 1624
rect 2140 1616 2148 1624
rect 2148 1616 2149 1624
rect 2139 1615 2149 1616
rect 2235 1615 2245 1625
rect 2779 1595 2789 1605
rect 3451 1595 3461 1605
rect 3515 1604 3525 1605
rect 3515 1596 3516 1604
rect 3516 1596 3524 1604
rect 3524 1596 3525 1604
rect 3515 1595 3525 1596
rect 3611 1595 3621 1605
rect 3931 1595 3941 1605
rect 3995 1595 4005 1605
rect 955 1575 965 1585
rect 1627 1555 1637 1565
rect 2363 1555 2373 1565
rect 1979 1535 1989 1545
rect 2427 1535 2437 1545
rect 3227 1555 3237 1565
rect 3419 1575 3429 1585
rect 2491 1535 2501 1545
rect 2587 1535 2597 1545
rect 2619 1535 2629 1545
rect 2779 1535 2789 1545
rect 1659 1515 1669 1525
rect 1787 1524 1797 1525
rect 1787 1516 1788 1524
rect 1788 1516 1796 1524
rect 1796 1516 1797 1524
rect 1787 1515 1797 1516
rect 2011 1515 2021 1525
rect 2331 1515 2341 1525
rect 2427 1515 2437 1525
rect 2587 1515 2597 1525
rect 2779 1515 2789 1525
rect 3003 1524 3013 1525
rect 3003 1516 3004 1524
rect 3004 1516 3012 1524
rect 3012 1516 3013 1524
rect 3099 1535 3109 1545
rect 3003 1515 3013 1516
rect 3227 1515 3237 1525
rect 3451 1515 3461 1525
rect 3643 1515 3653 1525
rect 4091 1515 4101 1525
rect 4123 1515 4133 1525
rect 5083 1515 5093 1525
rect 5083 1504 5093 1505
rect 5083 1496 5084 1504
rect 5084 1496 5092 1504
rect 5092 1496 5093 1504
rect 5083 1495 5093 1496
rect 2011 1475 2021 1485
rect 2043 1475 2053 1485
rect 2107 1475 2117 1485
rect 2811 1475 2821 1485
rect 1147 1455 1157 1465
rect 1211 1455 1221 1465
rect 4091 1455 4101 1465
rect 4923 1464 4933 1465
rect 4923 1456 4924 1464
rect 4924 1456 4932 1464
rect 4932 1456 4933 1464
rect 4923 1455 4933 1456
rect 4955 1455 4965 1465
rect 347 1435 357 1445
rect 1787 1435 1797 1445
rect 2043 1435 2053 1445
rect 2267 1435 2277 1445
rect 2427 1435 2437 1445
rect 3163 1435 3173 1445
rect 2779 1415 2789 1425
rect 3643 1415 3653 1425
rect 3675 1415 3685 1425
rect 1211 1395 1221 1405
rect 2139 1395 2149 1405
rect 2235 1395 2245 1405
rect 1915 1355 1925 1365
rect 1947 1355 1957 1365
rect 2363 1355 2373 1365
rect 2619 1355 2629 1365
rect 3003 1355 3013 1365
rect 3195 1355 3205 1365
rect 3291 1355 3301 1365
rect 4059 1355 4069 1365
rect 2555 1335 2565 1345
rect 2779 1335 2789 1345
rect 3067 1335 3077 1345
rect 3771 1335 3781 1345
rect 2427 1315 2437 1325
rect 3675 1315 3685 1325
rect 4443 1315 4453 1325
rect 4859 1315 4869 1325
rect 859 1304 869 1305
rect 859 1296 860 1304
rect 860 1296 868 1304
rect 868 1296 869 1304
rect 859 1295 869 1296
rect 2139 1295 2149 1305
rect 2587 1295 2597 1305
rect 2843 1295 2853 1305
rect 3035 1295 3045 1305
rect 3067 1295 3077 1305
rect 3771 1295 3781 1305
rect 4443 1295 4453 1305
rect 4667 1304 4677 1305
rect 4667 1296 4668 1304
rect 4668 1296 4676 1304
rect 4676 1296 4677 1304
rect 4667 1295 4677 1296
rect 763 1275 773 1285
rect 763 1255 773 1265
rect 2011 1255 2021 1265
rect 2171 1264 2181 1265
rect 2171 1256 2172 1264
rect 2172 1256 2180 1264
rect 2180 1256 2181 1264
rect 2171 1255 2181 1256
rect 2235 1255 2245 1265
rect 4795 1275 4805 1285
rect 2523 1255 2533 1265
rect 2587 1255 2597 1265
rect 2907 1264 2917 1265
rect 1147 1244 1157 1245
rect 1147 1236 1148 1244
rect 1148 1236 1156 1244
rect 1156 1236 1157 1244
rect 1147 1235 1157 1236
rect 2427 1235 2437 1245
rect 2555 1235 2565 1245
rect 2907 1256 2908 1264
rect 2908 1256 2916 1264
rect 2916 1256 2917 1264
rect 2907 1255 2917 1256
rect 2939 1255 2949 1265
rect 3003 1255 3013 1265
rect 4443 1255 4453 1265
rect 4539 1235 4549 1245
rect 2427 1215 2437 1225
rect 2491 1215 2501 1225
rect 2619 1215 2629 1225
rect 2779 1215 2789 1225
rect 2811 1215 2821 1225
rect 3611 1215 3621 1225
rect 3771 1215 3781 1225
rect 3867 1215 3877 1225
rect 1371 1204 1381 1205
rect 1371 1196 1372 1204
rect 1372 1196 1380 1204
rect 1380 1196 1381 1204
rect 1371 1195 1381 1196
rect 2011 1195 2021 1205
rect 1339 1175 1349 1185
rect 1659 1175 1669 1185
rect 2235 1175 2245 1185
rect 3291 1175 3301 1185
rect 1115 1155 1125 1165
rect 2715 1155 2725 1165
rect 4187 1155 4197 1165
rect 4667 1155 4677 1165
rect 1051 1135 1061 1145
rect 1659 1135 1669 1145
rect 2171 1135 2181 1145
rect 2427 1135 2437 1145
rect 2619 1135 2629 1145
rect 2939 1135 2949 1145
rect 1147 1075 1157 1085
rect 1195 1095 1205 1105
rect 1723 1095 1733 1105
rect 2043 1095 2053 1105
rect 2491 1115 2501 1125
rect 3291 1115 3301 1125
rect 3995 1115 4005 1125
rect 4891 1115 4901 1125
rect 2171 1095 2181 1105
rect 2267 1095 2277 1105
rect 2523 1095 2533 1105
rect 4219 1095 4229 1105
rect 2043 1075 2053 1085
rect 2939 1075 2949 1085
rect 4795 1075 4805 1085
rect 1019 1055 1029 1065
rect 1051 1035 1061 1045
rect 1563 1055 1573 1065
rect 2523 1055 2533 1065
rect 3451 1055 3461 1065
rect 2011 1035 2021 1045
rect 4155 1055 4165 1065
rect 5179 1055 5189 1065
rect 3803 1035 3813 1045
rect 4155 1035 4165 1045
rect 4251 1044 4261 1045
rect 4251 1036 4252 1044
rect 4252 1036 4260 1044
rect 4260 1036 4261 1044
rect 4251 1035 4261 1036
rect 3643 1015 3653 1025
rect 1627 995 1637 1005
rect 2011 995 2021 1005
rect 2779 995 2789 1005
rect 2907 1004 2917 1005
rect 2907 996 2908 1004
rect 2908 996 2916 1004
rect 2916 996 2917 1004
rect 2907 995 2917 996
rect 2939 995 2949 1005
rect 3963 995 3973 1005
rect 5051 995 5061 1005
rect 3819 975 3829 985
rect 2491 964 2501 965
rect 2491 956 2492 964
rect 2492 956 2500 964
rect 2500 956 2501 964
rect 2491 955 2501 956
rect 2683 955 2693 965
rect 2811 955 2821 965
rect 3643 955 3653 965
rect 443 935 453 945
rect 1883 944 1893 945
rect 1627 915 1637 925
rect 1787 924 1797 925
rect 1787 916 1788 924
rect 1788 916 1796 924
rect 1796 916 1797 924
rect 1883 936 1884 944
rect 1884 936 1892 944
rect 1892 936 1893 944
rect 1883 935 1893 936
rect 2075 944 2085 945
rect 2075 936 2076 944
rect 2076 936 2084 944
rect 2084 936 2085 944
rect 2075 935 2085 936
rect 2427 935 2437 945
rect 2459 935 2469 945
rect 2715 935 2725 945
rect 1787 915 1797 916
rect 2075 895 2085 905
rect 2267 895 2277 905
rect 2971 895 2981 905
rect 3515 895 3525 905
rect 3931 875 3941 885
rect 3963 875 3973 885
rect 4955 875 4965 885
rect 2075 835 2085 845
rect 2715 835 2725 845
rect 1659 815 1669 825
rect 1915 824 1925 825
rect 1915 816 1916 824
rect 1916 816 1924 824
rect 1924 816 1925 824
rect 1915 815 1925 816
rect 2107 815 2117 825
rect 2235 815 2245 825
rect 2619 815 2629 825
rect 2779 815 2789 825
rect 5147 824 5157 825
rect 5147 816 5148 824
rect 5148 816 5156 824
rect 5156 816 5157 824
rect 5147 815 5157 816
rect 1915 775 1925 785
rect 2107 775 2117 785
rect 3035 795 3045 805
rect 4059 795 4069 805
rect 3771 775 3781 785
rect 4091 775 4101 785
rect 5179 775 5189 785
rect 763 764 773 765
rect 763 756 764 764
rect 764 756 772 764
rect 772 756 773 764
rect 763 755 773 756
rect 2555 755 2565 765
rect 2587 764 2597 765
rect 2587 756 2588 764
rect 2588 756 2596 764
rect 2596 756 2597 764
rect 2587 755 2597 756
rect 2779 755 2789 765
rect 4123 755 4133 765
rect 1787 735 1797 745
rect 1915 735 1925 745
rect 2203 735 2213 745
rect 2747 735 2757 745
rect 3579 735 3589 745
rect 4795 735 4805 745
rect 571 715 581 725
rect 2907 695 2917 705
rect 3771 715 3781 725
rect 667 675 677 685
rect 2011 675 2021 685
rect 2331 675 2341 685
rect 2747 684 2757 685
rect 2747 676 2748 684
rect 2748 676 2756 684
rect 2756 676 2757 684
rect 2747 675 2757 676
rect 3771 675 3781 685
rect 283 655 293 665
rect 2523 655 2533 665
rect 2875 655 2885 665
rect 2875 635 2885 645
rect 3355 655 3365 665
rect 3451 655 3461 665
rect 3483 635 3493 645
rect 3259 615 3269 625
rect 3355 615 3365 625
rect 3419 615 3429 625
rect 3899 615 3909 625
rect 795 595 805 605
rect 2299 595 2309 605
rect 2331 595 2341 605
rect 2427 604 2437 605
rect 2427 596 2428 604
rect 2428 596 2436 604
rect 2436 596 2437 604
rect 2427 595 2437 596
rect 2587 595 2597 605
rect 3419 595 3429 605
rect 4091 595 4101 605
rect 4507 615 4517 625
rect 4187 595 4197 605
rect 4699 595 4709 605
rect 2523 575 2533 585
rect 2843 575 2853 585
rect 571 555 581 565
rect 1691 555 1701 565
rect 1755 555 1765 565
rect 1819 555 1829 565
rect 2011 555 2021 565
rect 4123 555 4133 565
rect 4507 555 4517 565
rect 5083 555 5093 565
rect 795 515 805 525
rect 2043 504 2053 505
rect 2043 496 2044 504
rect 2044 496 2052 504
rect 2052 496 2053 504
rect 2043 495 2053 496
rect 3451 495 3461 505
rect 2235 484 2245 485
rect 2235 476 2236 484
rect 2236 476 2244 484
rect 2244 476 2245 484
rect 2235 475 2245 476
rect 2587 475 2597 485
rect 2651 484 2661 485
rect 3131 484 3141 485
rect 2651 476 2652 484
rect 2652 476 2660 484
rect 2660 476 2661 484
rect 3131 476 3132 484
rect 3132 476 3140 484
rect 3140 476 3141 484
rect 2651 475 2661 476
rect 3131 475 3141 476
rect 3259 484 3269 485
rect 3259 476 3260 484
rect 3260 476 3268 484
rect 3268 476 3269 484
rect 3259 475 3269 476
rect 4027 475 4037 485
rect 2267 455 2277 465
rect 2331 455 2341 465
rect 2875 455 2885 465
rect 4059 455 4069 465
rect 2811 435 2821 445
rect 2235 395 2245 405
rect 2491 404 2501 405
rect 2491 396 2492 404
rect 2492 396 2500 404
rect 2500 396 2501 404
rect 2491 395 2501 396
rect 2619 395 2629 405
rect 2907 395 2917 405
rect 3099 395 3109 405
rect 1563 375 1573 385
rect 1675 375 1685 385
rect 1851 375 1861 385
rect 2395 375 2405 385
rect 731 335 741 345
rect 955 335 965 345
rect 1051 335 1061 345
rect 3483 335 3493 345
rect 2171 315 2181 325
rect 2651 315 2661 325
rect 2971 315 2981 325
rect 2619 275 2629 285
rect 2939 275 2949 285
rect 3003 284 3013 285
rect 3003 276 3004 284
rect 3004 276 3012 284
rect 3012 276 3013 284
rect 3003 275 3013 276
rect 3035 275 3045 285
rect 4059 275 4069 285
rect 4827 275 4837 285
rect 1371 255 1381 265
rect 1787 255 1797 265
rect 1979 255 1989 265
rect 2635 255 2645 265
rect 3851 255 3861 265
rect 4315 255 4325 265
rect 4859 255 4869 265
rect 2011 235 2021 245
rect 2171 235 2181 245
rect 3163 235 3173 245
rect 3867 235 3877 245
rect 3931 235 3941 245
rect 1243 224 1253 225
rect 1243 216 1244 224
rect 1244 216 1252 224
rect 1252 216 1253 224
rect 1243 215 1253 216
rect 1275 215 1285 225
rect 2395 175 2405 185
rect 3115 175 3125 185
rect 4155 175 4165 185
rect 2587 155 2597 165
rect 2875 155 2885 165
rect 2939 155 2949 165
rect 699 135 709 145
rect 3611 135 3621 145
rect 5115 155 5125 165
rect 3771 135 3781 145
rect 283 115 293 125
rect 731 115 741 125
rect 2811 104 2821 105
rect 2811 96 2812 104
rect 2812 96 2820 104
rect 2820 96 2821 104
rect 2811 95 2821 96
rect 2875 75 2885 85
rect 3131 75 3141 85
<< metal6 >>
rect 3515 3535 3659 3545
rect 3515 3525 3525 3535
rect 2485 3455 3205 3465
rect 763 2765 773 3235
rect 475 2665 485 2735
rect 795 2585 805 2855
rect 283 2185 293 2215
rect 347 1445 357 2255
rect 443 1945 453 2535
rect 443 945 453 1935
rect 475 1685 485 2255
rect 283 125 293 655
rect 571 565 581 715
rect 667 685 677 2235
rect 731 345 741 2175
rect 763 1285 773 1975
rect 795 1805 805 2515
rect 827 2265 837 3315
rect 891 2545 901 3135
rect 859 2225 869 2255
rect 827 2025 837 2075
rect 859 1305 869 1955
rect 923 1765 933 2555
rect 955 1585 965 2655
rect 763 765 773 1255
rect 1019 1065 1029 1895
rect 1051 1785 1061 2875
rect 1115 2345 1125 3335
rect 1115 1165 1125 1915
rect 1179 1825 1189 2895
rect 1243 1705 1253 2895
rect 1275 2405 1285 2455
rect 1275 2025 1285 2175
rect 1307 1825 1317 3155
rect 1371 2925 1381 3155
rect 1435 2885 1445 3035
rect 1499 2645 1509 2695
rect 1531 2645 1541 2675
rect 1467 2565 1477 2635
rect 1147 1245 1157 1455
rect 1211 1405 1221 1455
rect 1051 1045 1061 1135
rect 1147 1095 1195 1105
rect 1147 1085 1157 1095
rect 795 525 805 595
rect 955 305 965 335
rect 1051 305 1061 335
rect 955 295 1061 305
rect 1243 225 1253 1695
rect 1275 1685 1285 1735
rect 1339 1185 1349 1915
rect 1371 1205 1381 2095
rect 1435 1765 1445 2555
rect 1563 2445 1573 2575
rect 1595 2445 1605 3195
rect 1467 1945 1477 2195
rect 1499 2005 1509 2315
rect 1531 1645 1541 2435
rect 1563 1065 1573 2175
rect 1595 2105 1605 2155
rect 1595 1865 1605 1955
rect 1627 1565 1637 2475
rect 1659 1965 1669 3115
rect 1691 2165 1701 3135
rect 1723 3065 1733 3375
rect 1851 3245 1861 3335
rect 1755 3105 1765 3135
rect 1723 3055 1765 3065
rect 1723 2885 1733 2915
rect 1755 2585 1765 3055
rect 1883 2845 1893 3335
rect 2075 2985 2085 2995
rect 2171 2985 2181 2995
rect 2075 2975 2181 2985
rect 1723 2295 1797 2305
rect 1723 2265 1733 2295
rect 1787 2265 1797 2295
rect 1723 2045 1733 2075
rect 1659 1805 1669 1915
rect 1659 1185 1669 1515
rect 1627 925 1637 995
rect 1659 825 1669 1135
rect 1691 565 1701 2035
rect 1755 1825 1765 2255
rect 1819 2165 1829 2215
rect 1851 1985 1861 2655
rect 1915 2425 1925 2875
rect 2043 2725 2053 2815
rect 1883 2225 1893 2415
rect 1851 1865 1861 1875
rect 1787 1855 1861 1865
rect 1723 1105 1733 1615
rect 1755 565 1765 1635
rect 1787 1525 1797 1855
rect 1787 925 1797 1435
rect 1573 375 1675 385
rect 1787 265 1797 735
rect 1819 565 1829 1755
rect 1851 385 1861 1815
rect 1883 945 1893 1815
rect 1947 1365 1957 1735
rect 1979 1545 1989 2255
rect 2011 1685 2021 2535
rect 2075 2005 2085 2815
rect 2171 2005 2181 2035
rect 2011 1485 2021 1515
rect 2043 1445 2053 1475
rect 1915 825 1925 1355
rect 2011 1205 2021 1255
rect 2043 1085 2053 1095
rect 2011 1005 2021 1035
rect 1915 745 1925 775
rect 2011 565 2021 675
rect 2043 505 2053 1075
rect 2075 945 2085 1895
rect 2171 1825 2181 1975
rect 2203 1945 2213 2915
rect 2235 2805 2245 3435
rect 2395 3105 2405 3435
rect 2523 3325 2533 3435
rect 3195 3425 3205 3455
rect 2395 3095 2501 3105
rect 2491 3045 2501 3095
rect 2421 2935 2501 2945
rect 2491 2925 2501 2935
rect 2235 1965 2245 2675
rect 2171 1815 2213 1825
rect 2107 1485 2117 1655
rect 2139 1625 2149 1695
rect 2139 1305 2149 1395
rect 2171 1265 2181 1795
rect 2171 1105 2181 1135
rect 2075 845 2085 895
rect 2107 785 2117 815
rect 2203 745 2213 1815
rect 2235 1625 2245 1775
rect 2267 1765 2277 2695
rect 2299 1785 2309 2635
rect 2363 1845 2373 2775
rect 2459 2625 2469 2915
rect 2491 2525 2501 2615
rect 2331 1525 2341 1815
rect 2363 1645 2373 1815
rect 2235 1265 2245 1395
rect 2235 825 2245 1175
rect 2267 1105 2277 1435
rect 2363 1365 2373 1555
rect 2235 405 2245 475
rect 2267 465 2277 895
rect 2331 605 2341 675
rect 2299 465 2309 595
rect 2299 455 2331 465
rect 2395 385 2405 2135
rect 2427 2045 2437 2295
rect 2459 1825 2469 2455
rect 2427 1545 2437 1815
rect 2427 1445 2437 1515
rect 2427 1245 2437 1315
rect 2427 1145 2437 1215
rect 2459 945 2469 1795
rect 2491 1785 2501 2115
rect 2523 1925 2533 3315
rect 3323 3455 3493 3465
rect 2683 2745 2693 3175
rect 2587 2525 2597 2555
rect 2555 1885 2565 2495
rect 2619 2045 2629 2235
rect 2651 2225 2661 2495
rect 2491 1685 2501 1715
rect 2491 1545 2501 1635
rect 2523 1265 2533 1875
rect 2555 1745 2565 1835
rect 2587 1805 2597 2035
rect 2651 1865 2661 1995
rect 2555 1345 2565 1715
rect 2587 1545 2597 1775
rect 2619 1545 2629 1635
rect 2587 1305 2597 1515
rect 2491 1125 2501 1215
rect 2523 1065 2533 1095
rect 2427 605 2437 935
rect 2491 405 2501 955
rect 2555 765 2565 1235
rect 2587 765 2597 1255
rect 2619 1225 2629 1355
rect 2619 825 2629 1135
rect 2523 585 2533 655
rect 2587 485 2597 595
rect 2651 485 2661 1655
rect 2683 965 2693 2055
rect 2715 2045 2725 3415
rect 3035 3365 3045 3395
rect 3067 3265 3077 3355
rect 3131 3305 3141 3395
rect 3323 3385 3333 3455
rect 3483 3425 3493 3455
rect 3227 3345 3237 3375
rect 3387 3345 3397 3395
rect 3227 3335 3397 3345
rect 3419 3375 3579 3385
rect 3419 3305 3429 3375
rect 3067 3045 3077 3115
rect 3131 2985 3141 3295
rect 2715 1945 2725 1995
rect 2715 1165 2725 1775
rect 2715 845 2725 935
rect 2747 745 2757 2555
rect 2779 2425 2789 2475
rect 2843 2465 2853 2535
rect 2779 1665 2789 2315
rect 2811 2045 2821 2435
rect 2843 2105 2853 2215
rect 2843 2025 2853 2035
rect 2811 2015 2853 2025
rect 2811 1905 2821 2015
rect 2811 1665 2821 1855
rect 2843 1725 2853 1995
rect 2779 1545 2789 1595
rect 2779 1425 2789 1515
rect 2779 1225 2789 1335
rect 2811 1225 2821 1475
rect 2779 825 2789 995
rect 2779 705 2789 755
rect 2747 695 2789 705
rect 2747 685 2757 695
rect 2811 445 2821 955
rect 2843 585 2853 1295
rect 2875 665 2885 2495
rect 2907 1265 2917 2475
rect 2939 2045 2949 2735
rect 2971 2465 2981 2495
rect 3003 2465 3013 2495
rect 2971 2165 2981 2195
rect 3003 2045 3013 2315
rect 3067 1965 3077 2555
rect 3099 2385 3109 2915
rect 3131 2725 3141 2975
rect 3131 2465 3141 2495
rect 3291 2465 3301 2755
rect 3131 2145 3141 2155
rect 3131 2135 3301 2145
rect 3291 2105 3301 2135
rect 2939 1685 2949 1955
rect 2939 1145 2949 1255
rect 2939 1005 2949 1075
rect 2907 705 2917 995
rect 2971 905 2981 1875
rect 3003 1865 3013 1875
rect 3003 1855 3045 1865
rect 3035 1845 3045 1855
rect 3099 1545 3109 1855
rect 3003 1465 3013 1515
rect 3003 1455 3173 1465
rect 3163 1445 3173 1455
rect 3195 1365 3205 1955
rect 3227 1525 3237 1555
rect 3291 1365 3301 2015
rect 3323 1505 3333 2915
rect 3451 2165 3461 2875
rect 3419 1585 3429 1635
rect 3451 1605 3461 2075
rect 3451 1505 3461 1515
rect 3323 1495 3461 1505
rect 3003 1265 3013 1355
rect 3067 1305 3077 1335
rect 3035 805 3045 1295
rect 3291 1125 3301 1175
rect 3483 1105 3493 2315
rect 3515 1885 3525 2715
rect 3547 1685 3557 3055
rect 3579 1745 3589 2095
rect 3611 2085 3621 3495
rect 4821 3455 4869 3465
rect 4859 3445 4869 3455
rect 3707 3385 3717 3395
rect 3669 3375 3685 3385
rect 3707 3375 3819 3385
rect 3675 3345 3685 3375
rect 4027 3345 4037 3355
rect 3675 3335 4037 3345
rect 3995 2655 4197 2665
rect 3995 2645 4005 2655
rect 4187 2645 4197 2655
rect 3739 2105 3749 2475
rect 3771 2225 3781 2255
rect 3611 1745 3621 1895
rect 3707 1865 3717 1915
rect 3739 1865 3749 2095
rect 3451 1095 3493 1105
rect 3451 1065 3461 1095
rect 3515 905 3525 1595
rect 3611 1225 3621 1595
rect 3643 1425 3653 1515
rect 3675 1325 3685 1415
rect 3771 1305 3781 1335
rect 3643 965 3653 1015
rect 3771 785 3781 1215
rect 3803 1045 3813 2215
rect 3835 1785 3845 2635
rect 3867 2505 3877 2595
rect 3867 2495 3899 2505
rect 3867 2255 3883 2265
rect 3867 1865 3877 2255
rect 3963 2225 3973 2255
rect 3995 2205 4005 2335
rect 3931 1605 3941 2015
rect 3867 985 3877 1215
rect 3995 1125 4005 1595
rect 3829 975 3877 985
rect 3963 885 3973 995
rect 3579 705 3589 735
rect 3451 695 3589 705
rect 3451 665 3461 695
rect 3771 685 3781 715
rect 3483 655 3909 665
rect 2875 465 2885 635
rect 3355 625 3365 655
rect 3483 645 3493 655
rect 3899 625 3909 655
rect 3429 615 3461 625
rect 3259 585 3269 615
rect 3419 585 3429 595
rect 3259 575 3429 585
rect 3451 505 3461 615
rect 3131 495 3269 505
rect 3131 485 3141 495
rect 3259 485 3269 495
rect 1275 255 1371 265
rect 1989 255 2021 265
rect 1275 225 1285 255
rect 2011 245 2021 255
rect 2171 245 2181 315
rect 2619 285 2629 395
rect 2651 265 2661 315
rect 2645 255 2661 265
rect 2405 175 2597 185
rect 2587 165 2597 175
rect 709 135 741 145
rect 731 125 741 135
rect 2811 105 2821 435
rect 2907 385 2917 395
rect 3099 385 3109 395
rect 2907 375 3109 385
rect 3387 335 3483 345
rect 2939 225 2949 275
rect 2971 265 2981 315
rect 3387 305 3397 335
rect 3003 295 3397 305
rect 3003 285 3013 295
rect 3035 265 3045 275
rect 2971 255 3045 265
rect 3861 255 3877 265
rect 3867 245 3877 255
rect 3931 245 3941 875
rect 4027 485 4037 2415
rect 4059 2185 4069 2395
rect 4091 2205 4101 2375
rect 4155 2185 4165 2635
rect 4251 2525 4261 3295
rect 4059 2175 4123 2185
rect 4187 1825 4197 2515
rect 4283 1865 4293 2435
rect 4059 1775 4139 1785
rect 4059 1685 4069 1775
rect 4059 1365 4069 1655
rect 4091 1465 4101 1515
rect 4059 465 4069 795
rect 4091 605 4101 775
rect 4123 765 4133 1515
rect 4155 1065 4165 1675
rect 4155 745 4165 1035
rect 4123 735 4165 745
rect 4123 565 4133 735
rect 4187 605 4197 1155
rect 4219 1105 4229 1675
rect 4251 1045 4261 1635
rect 4059 285 4069 455
rect 4315 265 4325 2735
rect 4443 1325 4453 3435
rect 4507 2485 4517 2755
rect 4699 1745 4709 2375
rect 4763 1805 4773 3115
rect 4795 1825 4805 2235
rect 4443 1265 4453 1295
rect 4507 565 4517 615
rect 4539 585 4549 1235
rect 4667 1165 4677 1295
rect 4795 1085 4805 1275
rect 4795 745 4805 1075
rect 4699 585 4709 595
rect 4539 575 4709 585
rect 4827 285 4837 2735
rect 4859 1745 4869 1815
rect 4859 265 4869 1315
rect 4891 1125 4901 3315
rect 4923 2125 4933 3335
rect 4923 1465 4933 2075
rect 4955 885 4965 1455
rect 5051 1005 5061 2655
rect 5083 1785 5093 2715
rect 5083 1525 5093 1755
rect 5083 565 5093 1495
rect 3163 225 3173 235
rect 2939 215 3173 225
rect 3125 175 3333 185
rect 2875 85 2885 155
rect 2939 145 2949 155
rect 3323 145 3333 175
rect 4123 175 4155 185
rect 4123 145 4133 175
rect 5115 165 5125 3355
rect 5147 825 5157 2895
rect 5179 785 5189 1055
rect 2939 135 3109 145
rect 3323 135 3611 145
rect 3781 135 4133 145
rect 3099 105 3109 135
rect 3099 95 3141 105
rect 3131 85 3141 95
use NAND2X1  NAND2X1_302
timestamp 1598350056
transform 1 0 5096 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_21
timestamp 1598350056
transform -1 0 5096 0 1 3410
box -16 -6 64 210
use INVX1  INVX1_140
timestamp 1598350056
transform -1 0 5176 0 1 3410
box -18 -6 52 210
use FILL  FILL_18_2
timestamp 1598350056
transform 1 0 5192 0 1 3410
box -16 -6 32 210
use FILL  FILL_18_1
timestamp 1598350056
transform 1 0 5176 0 1 3410
box -16 -6 32 210
use NAND2X1  NAND2X1_408
timestamp 1598350056
transform 1 0 5000 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_30
timestamp 1598350056
transform -1 0 5000 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_36
timestamp 1598350056
transform -1 0 4952 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_17
timestamp 1598350056
transform 1 0 4856 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_21
timestamp 1598350056
transform -1 0 4856 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_30
timestamp 1598350056
transform -1 0 4808 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_31
timestamp 1598350056
transform -1 0 4760 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_51
timestamp 1598350056
transform 1 0 4664 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_1
timestamp 1598350056
transform -1 0 4664 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_22
timestamp 1598350056
transform 1 0 4568 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_11
timestamp 1598350056
transform 1 0 4424 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_51
timestamp 1598350056
transform 1 0 4376 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_50
timestamp 1598350056
transform 1 0 4520 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_408
timestamp 1598350056
transform -1 0 4520 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_50
timestamp 1598350056
transform -1 0 4376 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_22
timestamp 1598350056
transform 1 0 4280 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_18
timestamp 1598350056
transform -1 0 4280 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_1
timestamp 1598350056
transform -1 0 4232 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_17
timestamp 1598350056
transform 1 0 4136 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_36
timestamp 1598350056
transform -1 0 4136 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_12
timestamp 1598350056
transform -1 0 4088 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_429
timestamp 1598350056
transform -1 0 4040 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_31
timestamp 1598350056
transform -1 0 3992 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_3
timestamp 1598350056
transform -1 0 3944 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_581
timestamp 1598350056
transform -1 0 3896 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_582
timestamp 1598350056
transform 1 0 3800 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_762
timestamp 1598350056
transform -1 0 3800 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_59
timestamp 1598350056
transform -1 0 3752 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_25
timestamp 1598350056
transform -1 0 3704 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_587
timestamp 1598350056
transform -1 0 3656 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_588
timestamp 1598350056
transform -1 0 3608 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_40
timestamp 1598350056
transform -1 0 3560 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_26
timestamp 1598350056
transform 1 0 3464 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_70
timestamp 1598350056
transform 1 0 3416 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_64
timestamp 1598350056
transform 1 0 3368 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_2
timestamp 1598350056
transform -1 0 3368 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_157
timestamp 1598350056
transform -1 0 3320 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_47
timestamp 1598350056
transform -1 0 3272 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_769
timestamp 1598350056
transform -1 0 3224 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_467
timestamp 1598350056
transform 1 0 3080 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_44
timestamp 1598350056
transform -1 0 3032 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_764
timestamp 1598350056
transform 1 0 3128 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_163
timestamp 1598350056
transform 1 0 3032 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_452
timestamp 1598350056
transform 1 0 2936 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_328
timestamp 1598350056
transform 1 0 2888 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_386
timestamp 1598350056
transform -1 0 2888 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_387
timestamp 1598350056
transform 1 0 2792 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_425
timestamp 1598350056
transform 1 0 2744 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_427
timestamp 1598350056
transform -1 0 2712 0 1 3410
box -16 -6 64 210
use INVX1  INVX1_192
timestamp 1598350056
transform 1 0 2712 0 1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_450
timestamp 1598350056
transform -1 0 2664 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_426
timestamp 1598350056
transform 1 0 2568 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_163
timestamp 1598350056
transform -1 0 2568 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_160
timestamp 1598350056
transform -1 0 2520 0 1 3410
box -16 -6 64 210
use INVX1  INVX1_115
timestamp 1598350056
transform -1 0 2328 0 1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_162
timestamp 1598350056
transform 1 0 2424 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_161
timestamp 1598350056
transform 1 0 2376 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_466
timestamp 1598350056
transform -1 0 2376 0 1 3410
box -16 -6 64 210
use INVX1  INVX1_103
timestamp 1598350056
transform 1 0 2216 0 1 3410
box -18 -6 52 210
use INVX1  INVX1_189
timestamp 1598350056
transform -1 0 2168 0 1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_221
timestamp 1598350056
transform -1 0 2296 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_223
timestamp 1598350056
transform 1 0 2168 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_422
timestamp 1598350056
transform -1 0 2056 0 1 3410
box -16 -6 64 210
use INVX1  INVX1_295
timestamp 1598350056
transform -1 0 2088 0 1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_453
timestamp 1598350056
transform -1 0 2136 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_448
timestamp 1598350056
transform -1 0 2008 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_421
timestamp 1598350056
transform 1 0 1912 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_766
timestamp 1598350056
transform -1 0 1864 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_771
timestamp 1598350056
transform 1 0 1864 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_770
timestamp 1598350056
transform -1 0 1816 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_375
timestamp 1598350056
transform -1 0 1768 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_459
timestamp 1598350056
transform -1 0 1672 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_376
timestamp 1598350056
transform 1 0 1672 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_378
timestamp 1598350056
transform -1 0 1624 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_259
timestamp 1598350056
transform -1 0 1544 0 1 3410
box -16 -6 64 210
use INVX1  INVX1_32
timestamp 1598350056
transform -1 0 1576 0 1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_258
timestamp 1598350056
transform -1 0 1496 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_145
timestamp 1598350056
transform 1 0 1400 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_628
timestamp 1598350056
transform 1 0 1352 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_148
timestamp 1598350056
transform -1 0 1352 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_149
timestamp 1598350056
transform 1 0 1256 0 1 3410
box -16 -6 64 210
use INVX1  INVX1_193
timestamp 1598350056
transform -1 0 1208 0 1 3410
box -18 -6 52 210
use INVX1  INVX1_75
timestamp 1598350056
transform 1 0 1144 0 1 3410
box -18 -6 52 210
use INVX1  INVX1_174
timestamp 1598350056
transform -1 0 1096 0 1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_146
timestamp 1598350056
transform -1 0 1256 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_546
timestamp 1598350056
transform 1 0 1096 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_526
timestamp 1598350056
transform 1 0 968 0 1 3410
box -16 -6 64 210
use INVX1  INVX1_86
timestamp 1598350056
transform 1 0 936 0 1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_705
timestamp 1598350056
transform 1 0 1016 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_706
timestamp 1598350056
transform -1 0 936 0 1 3410
box -16 -6 64 210
use INVX1  INVX1_76
timestamp 1598350056
transform -1 0 792 0 1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_713
timestamp 1598350056
transform -1 0 888 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_463
timestamp 1598350056
transform 1 0 792 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_379
timestamp 1598350056
transform 1 0 712 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_380
timestamp 1598350056
transform -1 0 712 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_409
timestamp 1598350056
transform 1 0 568 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_460
timestamp 1598350056
transform 1 0 616 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_682
timestamp 1598350056
transform 1 0 520 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_694
timestamp 1598350056
transform -1 0 520 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_725
timestamp 1598350056
transform -1 0 472 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_707
timestamp 1598350056
transform 1 0 376 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_695
timestamp 1598350056
transform -1 0 376 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_696
timestamp 1598350056
transform -1 0 280 0 1 3410
box -16 -6 64 210
use INVX1  INVX1_287
timestamp 1598350056
transform -1 0 232 0 1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_712
timestamp 1598350056
transform 1 0 280 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_782
timestamp 1598350056
transform -1 0 200 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_744
timestamp 1598350056
transform -1 0 104 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_708
timestamp 1598350056
transform 1 0 104 0 1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_780
timestamp 1598350056
transform -1 0 56 0 1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_303
timestamp 1598350056
transform 1 0 5144 0 -1 3410
box -16 -6 64 210
use INVX1  INVX1_173
timestamp 1598350056
transform -1 0 5144 0 -1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_2
timestamp 1598350056
transform -1 0 5112 0 -1 3410
box -16 -6 64 210
use FILL  FILL_17_1
timestamp 1598350056
transform -1 0 5208 0 -1 3410
box -16 -6 32 210
use NAND2X1  NAND2X1_737
timestamp 1598350056
transform -1 0 4936 0 -1 3410
box -16 -6 64 210
use INVX1  INVX1_296
timestamp 1598350056
transform -1 0 5064 0 -1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_11
timestamp 1598350056
transform 1 0 4984 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_157
timestamp 1598350056
transform 1 0 4936 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_44
timestamp 1598350056
transform 1 0 4840 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_25
timestamp 1598350056
transform 1 0 4792 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_587
timestamp 1598350056
transform 1 0 4744 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_47
timestamp 1598350056
transform 1 0 4696 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_40
timestamp 1598350056
transform -1 0 4696 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_12
timestamp 1598350056
transform -1 0 4648 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_3
timestamp 1598350056
transform 1 0 4552 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_581
timestamp 1598350056
transform -1 0 4552 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_762
timestamp 1598350056
transform -1 0 4504 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_429
timestamp 1598350056
transform 1 0 4408 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_582
timestamp 1598350056
transform -1 0 4408 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_95
timestamp 1598350056
transform 1 0 4264 0 -1 3410
box -16 -6 64 210
use INVX1  INVX1_244
timestamp 1598350056
transform -1 0 4264 0 -1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_588
timestamp 1598350056
transform -1 0 4360 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_430
timestamp 1598350056
transform -1 0 4232 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_635
timestamp 1598350056
transform 1 0 4136 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_428
timestamp 1598350056
transform 1 0 4088 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_763
timestamp 1598350056
transform -1 0 4088 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_451
timestamp 1598350056
transform 1 0 3992 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_430
timestamp 1598350056
transform 1 0 3944 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_451
timestamp 1598350056
transform -1 0 3944 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_452
timestamp 1598350056
transform -1 0 3896 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_583
timestamp 1598350056
transform -1 0 3848 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_639
timestamp 1598350056
transform -1 0 3752 0 -1 3410
box -16 -6 64 210
use INVX1  INVX1_262
timestamp 1598350056
transform 1 0 3672 0 -1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_635
timestamp 1598350056
transform -1 0 3800 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_584
timestamp 1598350056
transform 1 0 3576 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_651
timestamp 1598350056
transform 1 0 3496 0 -1 3410
box -16 -6 64 210
use INVX1  INVX1_243
timestamp 1598350056
transform -1 0 3576 0 -1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_636
timestamp 1598350056
transform 1 0 3624 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_428
timestamp 1598350056
transform 1 0 3448 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_638
timestamp 1598350056
transform 1 0 3352 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_48
timestamp 1598350056
transform 1 0 3400 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_763
timestamp 1598350056
transform -1 0 3352 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_663
timestamp 1598350056
transform 1 0 3208 0 -1 3410
box -16 -6 64 210
use INVX1  INVX1_268
timestamp 1598350056
transform -1 0 3208 0 -1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_769
timestamp 1598350056
transform 1 0 3256 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_764
timestamp 1598350056
transform -1 0 3176 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_209
timestamp 1598350056
transform 1 0 3080 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_161
timestamp 1598350056
transform -1 0 3080 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_162
timestamp 1598350056
transform 1 0 2984 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_160
timestamp 1598350056
transform 1 0 2936 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_155
timestamp 1598350056
transform 1 0 2888 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_154
timestamp 1598350056
transform 1 0 2840 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_156
timestamp 1598350056
transform -1 0 2840 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_158
timestamp 1598350056
transform -1 0 2792 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_213
timestamp 1598350056
transform -1 0 2744 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_220
timestamp 1598350056
transform -1 0 2664 0 -1 3410
box -16 -6 64 210
use INVX1  INVX1_114
timestamp 1598350056
transform 1 0 2664 0 -1 3410
box -18 -6 52 210
use INVX1  INVX1_199
timestamp 1598350056
transform -1 0 2520 0 -1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_210
timestamp 1598350056
transform 1 0 2568 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_467
timestamp 1598350056
transform -1 0 2568 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_470
timestamp 1598350056
transform -1 0 2488 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_480
timestamp 1598350056
transform 1 0 2264 0 -1 3410
box -16 -6 64 210
use INVX1  INVX1_204
timestamp 1598350056
transform -1 0 2344 0 -1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_477
timestamp 1598350056
transform 1 0 2392 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_478
timestamp 1598350056
transform 1 0 2344 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_449
timestamp 1598350056
transform -1 0 2216 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_424
timestamp 1598350056
transform 1 0 2216 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_589
timestamp 1598350056
transform -1 0 2168 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_592
timestamp 1598350056
transform -1 0 2120 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_76
timestamp 1598350056
transform -1 0 1992 0 -1 3410
box -16 -6 64 210
use INVX1  INVX1_245
timestamp 1598350056
transform -1 0 2072 0 -1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_74
timestamp 1598350056
transform -1 0 2040 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_260
timestamp 1598350056
transform 1 0 1784 0 -1 3410
box -16 -6 64 210
use INVX1  INVX1_55
timestamp 1598350056
transform -1 0 1944 0 -1 3410
box -18 -6 52 210
use INVX1  INVX1_298
timestamp 1598350056
transform 1 0 1880 0 -1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_261
timestamp 1598350056
transform 1 0 1832 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_765
timestamp 1598350056
transform -1 0 1784 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_345
timestamp 1598350056
transform 1 0 1656 0 -1 3410
box -16 -6 64 210
use INVX1  INVX1_153
timestamp 1598350056
transform 1 0 1704 0 -1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_377
timestamp 1598350056
transform 1 0 1608 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_630
timestamp 1598350056
transform 1 0 1464 0 -1 3410
box -16 -6 64 210
use INVX1  INVX1_259
timestamp 1598350056
transform -1 0 1464 0 -1 3410
box -18 -6 52 210
use INVX1  INVX1_121
timestamp 1598350056
transform -1 0 1432 0 -1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_684
timestamp 1598350056
transform 1 0 1560 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_257
timestamp 1598350056
transform 1 0 1512 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_686
timestamp 1598350056
transform -1 0 1320 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_693
timestamp 1598350056
transform -1 0 1272 0 -1 3410
box -16 -6 64 210
use INVX1  INVX1_257
timestamp 1598350056
transform 1 0 1368 0 -1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_683
timestamp 1598350056
transform 1 0 1320 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_484
timestamp 1598350056
transform -1 0 1224 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_525
timestamp 1598350056
transform -1 0 1176 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_486
timestamp 1598350056
transform 1 0 1080 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_485
timestamp 1598350056
transform 1 0 1032 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_144
timestamp 1598350056
transform -1 0 1032 0 -1 3410
box -16 -6 64 210
use INVX1  INVX1_275
timestamp 1598350056
transform -1 0 984 0 -1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_147
timestamp 1598350056
transform -1 0 952 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_692
timestamp 1598350056
transform 1 0 856 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_142
timestamp 1598350056
transform 1 0 808 0 -1 3410
box -16 -6 64 210
use INVX1  INVX1_198
timestamp 1598350056
transform -1 0 808 0 -1 3410
box -18 -6 52 210
use NOR2X1  NOR2X1_746
timestamp 1598350056
transform 1 0 728 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_781
timestamp 1598350056
transform -1 0 680 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_745
timestamp 1598350056
transform -1 0 728 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_687
timestamp 1598350056
transform -1 0 632 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_685
timestamp 1598350056
transform -1 0 584 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_681
timestamp 1598350056
transform -1 0 536 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_511
timestamp 1598350056
transform -1 0 488 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_732
timestamp 1598350056
transform -1 0 440 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_747
timestamp 1598350056
transform -1 0 392 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_700
timestamp 1598350056
transform -1 0 344 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_701
timestamp 1598350056
transform -1 0 296 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_710
timestamp 1598350056
transform -1 0 248 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_743
timestamp 1598350056
transform -1 0 200 0 -1 3410
box -16 -6 64 210
use NAND2X1  NAND2X1_697
timestamp 1598350056
transform -1 0 152 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_779
timestamp 1598350056
transform 1 0 56 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_783
timestamp 1598350056
transform 1 0 8 0 -1 3410
box -16 -6 64 210
use NOR2X1  NOR2X1_386
timestamp 1598350056
transform 1 0 5128 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_571
timestamp 1598350056
transform 1 0 5080 0 1 3010
box -16 -6 64 210
use FILL  FILL_16_2
timestamp 1598350056
transform 1 0 5192 0 1 3010
box -16 -6 32 210
use FILL  FILL_16_1
timestamp 1598350056
transform 1 0 5176 0 1 3010
box -16 -6 32 210
use NOR2X1  NOR2X1_59
timestamp 1598350056
transform -1 0 5080 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_18
timestamp 1598350056
transform 1 0 4984 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_70
timestamp 1598350056
transform 1 0 4936 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_328
timestamp 1598350056
transform 1 0 4888 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_425
timestamp 1598350056
transform -1 0 4888 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_694
timestamp 1598350056
transform -1 0 4840 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_426
timestamp 1598350056
transform -1 0 4792 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_450
timestamp 1598350056
transform -1 0 4696 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_95
timestamp 1598350056
transform 1 0 4696 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_427
timestamp 1598350056
transform 1 0 4600 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_752
timestamp 1598350056
transform -1 0 4600 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_752
timestamp 1598350056
transform -1 0 4440 0 1 3010
box -16 -6 64 210
use INVX1  INVX1_191
timestamp 1598350056
transform -1 0 4552 0 1 3010
box -18 -6 52 210
use INVX1  INVX1_187
timestamp 1598350056
transform -1 0 4472 0 1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_418
timestamp 1598350056
transform 1 0 4472 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_636
timestamp 1598350056
transform 1 0 4264 0 1 3010
box -16 -6 64 210
use INVX1  INVX1_261
timestamp 1598350056
transform -1 0 4344 0 1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_454
timestamp 1598350056
transform 1 0 4344 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_583
timestamp 1598350056
transform 1 0 4216 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_638
timestamp 1598350056
transform 1 0 4168 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_651
timestamp 1598350056
transform 1 0 4120 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_639
timestamp 1598350056
transform -1 0 4120 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_584
timestamp 1598350056
transform -1 0 4072 0 1 3010
box -16 -6 64 210
use INVX1  INVX1_77
timestamp 1598350056
transform 1 0 3992 0 1 3010
box -18 -6 52 210
use INVX1  INVX1_288
timestamp 1598350056
transform -1 0 3944 0 1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_747
timestamp 1598350056
transform -1 0 3992 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_782
timestamp 1598350056
transform 1 0 3864 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_797
timestamp 1598350056
transform 1 0 3736 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_654
timestamp 1598350056
transform -1 0 3736 0 1 3010
box -16 -6 64 210
use INVX1  INVX1_302
timestamp 1598350056
transform -1 0 3864 0 1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_158
timestamp 1598350056
transform -1 0 3832 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_637
timestamp 1598350056
transform -1 0 3640 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_745
timestamp 1598350056
transform 1 0 3496 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_781
timestamp 1598350056
transform -1 0 3688 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_585
timestamp 1598350056
transform 1 0 3544 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_586
timestamp 1598350056
transform -1 0 3496 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_229
timestamp 1598350056
transform -1 0 3448 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_230
timestamp 1598350056
transform -1 0 3400 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_231
timestamp 1598350056
transform -1 0 3352 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_196
timestamp 1598350056
transform 1 0 3208 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_199
timestamp 1598350056
transform -1 0 3208 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_45
timestamp 1598350056
transform 1 0 3256 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_53
timestamp 1598350056
transform -1 0 3128 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_210
timestamp 1598350056
transform -1 0 3032 0 1 3010
box -16 -6 64 210
use INVX1  INVX1_107
timestamp 1598350056
transform -1 0 3160 0 1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_75
timestamp 1598350056
transform -1 0 3080 0 1 3010
box -16 -6 64 210
use INVX1  INVX1_105
timestamp 1598350056
transform -1 0 2984 0 1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_207
timestamp 1598350056
transform 1 0 2904 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_200
timestamp 1598350056
transform 1 0 2856 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_194
timestamp 1598350056
transform 1 0 2808 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_16
timestamp 1598350056
transform 1 0 2760 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_39
timestamp 1598350056
transform 1 0 2680 0 1 3010
box -16 -6 64 210
use INVX1  INVX1_113
timestamp 1598350056
transform -1 0 2760 0 1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_300
timestamp 1598350056
transform -1 0 2680 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_831
timestamp 1598350056
transform -1 0 2632 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_301
timestamp 1598350056
transform 1 0 2536 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_841
timestamp 1598350056
transform -1 0 2536 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_433
timestamp 1598350056
transform 1 0 2440 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_435
timestamp 1598350056
transform -1 0 2344 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_273
timestamp 1598350056
transform -1 0 2440 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_432
timestamp 1598350056
transform -1 0 2392 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_832
timestamp 1598350056
transform 1 0 2248 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_605
timestamp 1598350056
transform 1 0 2152 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_604
timestamp 1598350056
transform 1 0 2200 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_603
timestamp 1598350056
transform -1 0 2152 0 1 3010
box -16 -6 64 210
use INVX1  INVX1_139
timestamp 1598350056
transform -1 0 2104 0 1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_737
timestamp 1598350056
transform -1 0 2072 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_741
timestamp 1598350056
transform -1 0 2024 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_733
timestamp 1598350056
transform -1 0 1976 0 1 3010
box -16 -6 64 210
use INVX1  INVX1_281
timestamp 1598350056
transform -1 0 1928 0 1 3010
box -18 -6 52 210
use INVX1  INVX1_283
timestamp 1598350056
transform 1 0 1768 0 1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_723
timestamp 1598350056
transform 1 0 1848 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_722
timestamp 1598350056
transform -1 0 1848 0 1 3010
box -16 -6 64 210
use INVX1  INVX1_249
timestamp 1598350056
transform 1 0 1688 0 1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_718
timestamp 1598350056
transform -1 0 1768 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_626
timestamp 1598350056
transform 1 0 1640 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_593
timestamp 1598350056
transform 1 0 1592 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_629
timestamp 1598350056
transform 1 0 1496 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_627
timestamp 1598350056
transform 1 0 1544 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_632
timestamp 1598350056
transform -1 0 1496 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_303
timestamp 1598350056
transform 1 0 1400 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_299
timestamp 1598350056
transform -1 0 1304 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_555
timestamp 1598350056
transform -1 0 1400 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_213
timestamp 1598350056
transform -1 0 1352 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_298
timestamp 1598350056
transform -1 0 1208 0 1 3010
box -16 -6 64 210
use INVX1  INVX1_85
timestamp 1598350056
transform -1 0 1112 0 1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_302
timestamp 1598350056
transform -1 0 1256 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_590
timestamp 1598350056
transform 1 0 1112 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_591
timestamp 1598350056
transform 1 0 1032 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_56
timestamp 1598350056
transform 1 0 984 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_252
timestamp 1598350056
transform -1 0 952 0 1 3010
box -16 -6 64 210
use INVX1  INVX1_311
timestamp 1598350056
transform -1 0 984 0 1 3010
box -18 -6 52 210
use NAND2X1  NAND2X1_304
timestamp 1598350056
transform -1 0 776 0 1 3010
box -16 -6 64 210
use INVX1  INVX1_83
timestamp 1598350056
transform 1 0 824 0 1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_306
timestamp 1598350056
transform 1 0 856 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_742
timestamp 1598350056
transform -1 0 824 0 1 3010
box -16 -6 64 210
use INVX1  INVX1_142
timestamp 1598350056
transform -1 0 728 0 1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_308
timestamp 1598350056
transform 1 0 648 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_727
timestamp 1598350056
transform 1 0 600 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_307
timestamp 1598350056
transform 1 0 552 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_740
timestamp 1598350056
transform -1 0 552 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_738
timestamp 1598350056
transform -1 0 504 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_731
timestamp 1598350056
transform -1 0 456 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_209
timestamp 1598350056
transform -1 0 408 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_305
timestamp 1598350056
transform -1 0 232 0 1 3010
box -16 -6 64 210
use INVX1  INVX1_277
timestamp 1598350056
transform -1 0 312 0 1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_726
timestamp 1598350056
transform 1 0 312 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_711
timestamp 1598350056
transform 1 0 232 0 1 3010
box -16 -6 64 210
use INVX1  INVX1_301
timestamp 1598350056
transform 1 0 56 0 1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_149
timestamp 1598350056
transform 1 0 136 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_797
timestamp 1598350056
transform 1 0 88 0 1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_796
timestamp 1598350056
transform -1 0 56 0 1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_460
timestamp 1598350056
transform -1 0 5192 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_732
timestamp 1598350056
transform 1 0 5096 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_505
timestamp 1598350056
transform 1 0 5048 0 -1 3010
box -16 -6 64 210
use FILL  FILL_15_1
timestamp 1598350056
transform -1 0 5208 0 -1 3010
box -16 -6 32 210
use NOR2X1  NOR2X1_26
timestamp 1598350056
transform -1 0 5048 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_64
timestamp 1598350056
transform 1 0 4952 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_695
timestamp 1598350056
transform 1 0 4904 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_707
timestamp 1598350056
transform 1 0 4856 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_712
timestamp 1598350056
transform -1 0 4856 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_53
timestamp 1598350056
transform -1 0 4808 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_696
timestamp 1598350056
transform 1 0 4712 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_708
timestamp 1598350056
transform -1 0 4664 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_227
timestamp 1598350056
transform -1 0 4616 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_224
timestamp 1598350056
transform 1 0 4664 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_446
timestamp 1598350056
transform -1 0 4488 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_509
timestamp 1598350056
transform -1 0 4440 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_289
timestamp 1598350056
transform 1 0 4488 0 -1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_226
timestamp 1598350056
transform 1 0 4520 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_211
timestamp 1598350056
transform -1 0 4344 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_146
timestamp 1598350056
transform -1 0 4216 0 -1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_417
timestamp 1598350056
transform 1 0 4344 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_447
timestamp 1598350056
transform 1 0 4264 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_330
timestamp 1598350056
transform 1 0 4216 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_420
timestamp 1598350056
transform 1 0 4088 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_356
timestamp 1598350056
transform -1 0 4088 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_329
timestamp 1598350056
transform -1 0 4184 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_355
timestamp 1598350056
transform -1 0 4040 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_155
timestamp 1598350056
transform -1 0 3944 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_331
timestamp 1598350056
transform 1 0 3944 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_594
timestamp 1598350056
transform -1 0 3896 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_156
timestamp 1598350056
transform 1 0 3752 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_154
timestamp 1598350056
transform 1 0 3704 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_653
timestamp 1598350056
transform 1 0 3656 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_697
timestamp 1598350056
transform 1 0 3800 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_661
timestamp 1598350056
transform -1 0 3656 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_662
timestamp 1598350056
transform -1 0 3608 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_43
timestamp 1598350056
transform 1 0 3512 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_746
timestamp 1598350056
transform 1 0 3432 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_423
timestamp 1598350056
transform 1 0 3336 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_117
timestamp 1598350056
transform -1 0 3512 0 -1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_13
timestamp 1598350056
transform 1 0 3384 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_195
timestamp 1598350056
transform -1 0 3288 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_193
timestamp 1598350056
transform 1 0 3192 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_341
timestamp 1598350056
transform 1 0 3144 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_41
timestamp 1598350056
transform 1 0 3288 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_228
timestamp 1598350056
transform -1 0 3096 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_758
timestamp 1598350056
transform -1 0 3048 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_7
timestamp 1598350056
transform -1 0 3144 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_159
timestamp 1598350056
transform -1 0 2904 0 -1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_759
timestamp 1598350056
transform 1 0 2952 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_659
timestamp 1598350056
transform -1 0 2952 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_365
timestamp 1598350056
transform 1 0 2824 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_716
timestamp 1598350056
transform -1 0 2680 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_364
timestamp 1598350056
transform -1 0 2824 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_367
timestamp 1598350056
transform 1 0 2728 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_222
timestamp 1598350056
transform -1 0 2728 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_212
timestamp 1598350056
transform 1 0 2584 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_469
timestamp 1598350056
transform 1 0 2536 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_214
timestamp 1598350056
transform 1 0 2488 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_142
timestamp 1598350056
transform -1 0 2488 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_206
timestamp 1598350056
transform 1 0 2392 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_219
timestamp 1598350056
transform 1 0 2344 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_215
timestamp 1598350056
transform -1 0 2344 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_52
timestamp 1598350056
transform 1 0 2168 0 -1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_423
timestamp 1598350056
transform 1 0 2248 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_202
timestamp 1598350056
transform -1 0 2248 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_69
timestamp 1598350056
transform 1 0 2120 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_68
timestamp 1598350056
transform 1 0 2072 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_658
timestamp 1598350056
transform 1 0 2024 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_736
timestamp 1598350056
transform 1 0 1976 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_735
timestamp 1598350056
transform -1 0 1976 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_664
timestamp 1598350056
transform 1 0 1832 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_719
timestamp 1598350056
transform -1 0 1832 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_665
timestamp 1598350056
transform 1 0 1880 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_67
timestamp 1598350056
transform 1 0 1736 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_147
timestamp 1598350056
transform -1 0 1736 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_144
timestamp 1598350056
transform -1 0 1688 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_66
timestamp 1598350056
transform 1 0 1592 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_625
timestamp 1598350056
transform -1 0 1592 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_136
timestamp 1598350056
transform -1 0 1544 0 -1 3010
box -18 -6 52 210
use INVX1  INVX1_96
timestamp 1598350056
transform 1 0 1432 0 -1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_57
timestamp 1598350056
transform 1 0 1464 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_631
timestamp 1598350056
transform -1 0 1432 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_556
timestamp 1598350056
transform 1 0 1336 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_562
timestamp 1598350056
transform 1 0 1288 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_357
timestamp 1598350056
transform 1 0 1240 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_44
timestamp 1598350056
transform -1 0 1144 0 -1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_353
timestamp 1598350056
transform 1 0 1192 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_208
timestamp 1598350056
transform 1 0 1144 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_198
timestamp 1598350056
transform 1 0 1064 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_50
timestamp 1598350056
transform 1 0 984 0 -1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_197
timestamp 1598350056
transform 1 0 1016 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_254
timestamp 1598350056
transform 1 0 936 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_483
timestamp 1598350056
transform 1 0 888 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_253
timestamp 1598350056
transform -1 0 840 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_709
timestamp 1598350056
transform -1 0 760 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_186
timestamp 1598350056
transform 1 0 760 0 -1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_698
timestamp 1598350056
transform 1 0 840 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_677
timestamp 1598350056
transform -1 0 712 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_851
timestamp 1598350056
transform -1 0 664 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_840
timestamp 1598350056
transform 1 0 568 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_482
timestamp 1598350056
transform 1 0 472 0 -1 3010
box -16 -6 64 210
use INVX1  INVX1_213
timestamp 1598350056
transform 1 0 440 0 -1 3010
box -18 -6 52 210
use NOR2X1  NOR2X1_834
timestamp 1598350056
transform -1 0 568 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_833
timestamp 1598350056
transform 1 0 392 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_152
timestamp 1598350056
transform 1 0 344 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_495
timestamp 1598350056
transform 1 0 248 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_407
timestamp 1598350056
transform -1 0 344 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_777
timestamp 1598350056
transform 1 0 200 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_146
timestamp 1598350056
transform -1 0 152 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_784
timestamp 1598350056
transform 1 0 152 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_148
timestamp 1598350056
transform -1 0 104 0 -1 3010
box -16 -6 64 210
use NOR2X1  NOR2X1_803
timestamp 1598350056
transform -1 0 56 0 -1 3010
box -16 -6 64 210
use NAND2X1  NAND2X1_507
timestamp 1598350056
transform 1 0 5112 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_857
timestamp 1598350056
transform 1 0 5064 0 1 2610
box -16 -6 64 210
use INVX1  INVX1_209
timestamp 1598350056
transform 1 0 5160 0 1 2610
box -18 -6 52 210
use FILL  FILL_14_1
timestamp 1598350056
transform 1 0 5192 0 1 2610
box -16 -6 32 210
use NAND2X1  NAND2X1_448
timestamp 1598350056
transform -1 0 5064 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_422
timestamp 1598350056
transform -1 0 5016 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_421
timestamp 1598350056
transform -1 0 4968 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_596
timestamp 1598350056
transform 1 0 4776 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_504
timestamp 1598350056
transform 1 0 4872 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_597
timestamp 1598350056
transform 1 0 4824 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_56
timestamp 1598350056
transform 1 0 4728 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_317
timestamp 1598350056
transform 1 0 4584 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_304
timestamp 1598350056
transform 1 0 4680 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_314
timestamp 1598350056
transform 1 0 4632 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_313
timestamp 1598350056
transform -1 0 4584 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_704
timestamp 1598350056
transform -1 0 4536 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_340
timestamp 1598350056
transform -1 0 4488 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_508
timestamp 1598350056
transform -1 0 4440 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_319
timestamp 1598350056
transform -1 0 4392 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_798
timestamp 1598350056
transform -1 0 4344 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_510
timestamp 1598350056
transform 1 0 4248 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_506
timestamp 1598350056
transform -1 0 4248 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_586
timestamp 1598350056
transform -1 0 4168 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_239
timestamp 1598350056
transform 1 0 4024 0 1 2610
box -16 -6 64 210
use INVX1  INVX1_144
timestamp 1598350056
transform 1 0 4168 0 1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_637
timestamp 1598350056
transform -1 0 4120 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_589
timestamp 1598350056
transform 1 0 3928 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_814
timestamp 1598350056
transform 1 0 3880 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_592
timestamp 1598350056
transform 1 0 3976 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_431
timestamp 1598350056
transform 1 0 3832 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_434
timestamp 1598350056
transform 1 0 3784 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_436
timestamp 1598350056
transform -1 0 3784 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_432
timestamp 1598350056
transform -1 0 3704 0 1 2610
box -16 -6 64 210
use INVX1  INVX1_180
timestamp 1598350056
transform 1 0 3704 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_63
timestamp 1598350056
transform 1 0 3624 0 1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_435
timestamp 1598350056
transform 1 0 3576 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_832
timestamp 1598350056
transform -1 0 3576 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_470
timestamp 1598350056
transform 1 0 3480 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_453
timestamp 1598350056
transform -1 0 3400 0 1 2610
box -16 -6 64 210
use INVX1  INVX1_190
timestamp 1598350056
transform -1 0 3432 0 1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_449
timestamp 1598350056
transform 1 0 3432 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_466
timestamp 1598350056
transform -1 0 3352 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_468
timestamp 1598350056
transform -1 0 3304 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_350
timestamp 1598350056
transform -1 0 3256 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_197
timestamp 1598350056
transform 1 0 3160 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_433
timestamp 1598350056
transform -1 0 3160 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_424
timestamp 1598350056
transform 1 0 3064 0 1 2610
box -16 -6 64 210
use INVX1  INVX1_157
timestamp 1598350056
transform -1 0 3016 0 1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_358
timestamp 1598350056
transform -1 0 3064 0 1 2610
box -16 -6 64 210
use INVX1  INVX1_109
timestamp 1598350056
transform -1 0 2984 0 1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_52
timestamp 1598350056
transform 1 0 2904 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_657
timestamp 1598350056
transform -1 0 2904 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_131
timestamp 1598350056
transform 1 0 2808 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_130
timestamp 1598350056
transform 1 0 2760 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_140
timestamp 1598350056
transform 1 0 2712 0 1 2610
box -16 -6 64 210
use INVX1  INVX1_81
timestamp 1598350056
transform -1 0 2664 0 1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_141
timestamp 1598350056
transform 1 0 2664 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_274
timestamp 1598350056
transform -1 0 2632 0 1 2610
box -16 -6 64 210
use INVX1  INVX1_130
timestamp 1598350056
transform -1 0 2536 0 1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_275
timestamp 1598350056
transform -1 0 2584 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_217
timestamp 1598350056
transform -1 0 2504 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_271
timestamp 1598350056
transform -1 0 2376 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_479
timestamp 1598350056
transform -1 0 2328 0 1 2610
box -16 -6 64 210
use INVX1  INVX1_73
timestamp 1598350056
transform 1 0 2424 0 1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_276
timestamp 1598350056
transform -1 0 2424 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_476
timestamp 1598350056
transform 1 0 2200 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_121
timestamp 1598350056
transform 1 0 2152 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_120
timestamp 1598350056
transform 1 0 2104 0 1 2610
box -16 -6 64 210
use INVX1  INVX1_202
timestamp 1598350056
transform -1 0 2280 0 1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_368
timestamp 1598350056
transform -1 0 2040 0 1 2610
box -16 -6 64 210
use INVX1  INVX1_271
timestamp 1598350056
transform -1 0 2104 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_6
timestamp 1598350056
transform -1 0 2072 0 1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_270
timestamp 1598350056
transform -1 0 1992 0 1 2610
box -16 -6 64 210
use INVX1  INVX1_88
timestamp 1598350056
transform -1 0 1944 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_10
timestamp 1598350056
transform -1 0 1864 0 1 2610
box -18 -6 52 210
use INVX1  INVX1_42
timestamp 1598350056
transform -1 0 1784 0 1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_666
timestamp 1598350056
transform 1 0 1864 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_151
timestamp 1598350056
transform -1 0 1832 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_597
timestamp 1598350056
transform -1 0 1704 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_717
timestamp 1598350056
transform -1 0 1752 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_596
timestamp 1598350056
transform -1 0 1656 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_645
timestamp 1598350056
transform 1 0 1560 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_471
timestamp 1598350056
transform -1 0 1560 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_457
timestamp 1598350056
transform 1 0 1464 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_464
timestamp 1598350056
transform 1 0 1416 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_602
timestamp 1598350056
transform 1 0 1320 0 1 2610
box -16 -6 64 210
use INVX1  INVX1_78
timestamp 1598350056
transform -1 0 1272 0 1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_458
timestamp 1598350056
transform 1 0 1368 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_601
timestamp 1598350056
transform -1 0 1320 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_178
timestamp 1598350056
transform 1 0 1048 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_352
timestamp 1598350056
transform 1 0 1192 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_680
timestamp 1598350056
transform 1 0 1144 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_182
timestamp 1598350056
transform 1 0 1096 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_179
timestamp 1598350056
transform 1 0 952 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_177
timestamp 1598350056
transform -1 0 952 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_181
timestamp 1598350056
transform 1 0 1000 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_176
timestamp 1598350056
transform 1 0 808 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_512
timestamp 1598350056
transform -1 0 808 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_513
timestamp 1598350056
transform 1 0 712 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_180
timestamp 1598350056
transform -1 0 904 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_472
timestamp 1598350056
transform 1 0 664 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_679
timestamp 1598350056
transform -1 0 616 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_676
timestamp 1598350056
transform 1 0 616 0 1 2610
box -16 -6 64 210
use INVX1  INVX1_274
timestamp 1598350056
transform -1 0 520 0 1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_739
timestamp 1598350056
transform 1 0 520 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_728
timestamp 1598350056
transform 1 0 440 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_730
timestamp 1598350056
transform 1 0 392 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_496
timestamp 1598350056
transform 1 0 200 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_729
timestamp 1598350056
transform 1 0 344 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_828
timestamp 1598350056
transform -1 0 344 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_499
timestamp 1598350056
transform 1 0 248 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_145
timestamp 1598350056
transform 1 0 8 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_313
timestamp 1598350056
transform 1 0 104 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_829
timestamp 1598350056
transform 1 0 56 0 1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_778
timestamp 1598350056
transform 1 0 152 0 1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_828
timestamp 1598350056
transform -1 0 5144 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_409
timestamp 1598350056
transform 1 0 5144 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_599
timestamp 1598350056
transform -1 0 5096 0 -1 2610
box -16 -6 64 210
use FILL  FILL_13_1
timestamp 1598350056
transform -1 0 5208 0 -1 2610
box -16 -6 32 210
use NAND2X1  NAND2X1_809
timestamp 1598350056
transform 1 0 4904 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_387
timestamp 1598350056
transform 1 0 5000 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_761
timestamp 1598350056
transform -1 0 5000 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_801
timestamp 1598350056
transform -1 0 4904 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_644
timestamp 1598350056
transform -1 0 4856 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_598
timestamp 1598350056
transform 1 0 4760 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_407
timestamp 1598350056
transform -1 0 4760 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_676
timestamp 1598350056
transform 1 0 4664 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_679
timestamp 1598350056
transform 1 0 4616 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_503
timestamp 1598350056
transform 1 0 4568 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_502
timestamp 1598350056
transform 1 0 4520 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_802
timestamp 1598350056
transform 1 0 4472 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_799
timestamp 1598350056
transform -1 0 4472 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_593
timestamp 1598350056
transform -1 0 4424 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_354
timestamp 1598350056
transform 1 0 4296 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_419
timestamp 1598350056
transform 1 0 4200 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_246
timestamp 1598350056
transform 1 0 4344 0 -1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_677
timestamp 1598350056
transform 1 0 4248 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_678
timestamp 1598350056
transform 1 0 4152 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_175
timestamp 1598350056
transform -1 0 4120 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_585
timestamp 1598350056
transform -1 0 4072 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_272
timestamp 1598350056
transform 1 0 4120 0 -1 2610
box -18 -6 52 210
use NAND2X1  NAND2X1_186
timestamp 1598350056
transform 1 0 3976 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_174
timestamp 1598350056
transform 1 0 3832 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_173
timestamp 1598350056
transform -1 0 3976 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_815
timestamp 1598350056
transform -1 0 3928 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_333
timestamp 1598350056
transform -1 0 3784 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_652
timestamp 1598350056
transform 1 0 3688 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_171
timestamp 1598350056
transform 1 0 3784 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_61
timestamp 1598350056
transform -1 0 3544 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_289
timestamp 1598350056
transform 1 0 3640 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_58
timestamp 1598350056
transform -1 0 3640 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_60
timestamp 1598350056
transform 1 0 3544 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_201
timestamp 1598350056
transform -1 0 3464 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_147
timestamp 1598350056
transform -1 0 3496 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_128
timestamp 1598350056
transform -1 0 3368 0 -1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_268
timestamp 1598350056
transform 1 0 3368 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_339
timestamp 1598350056
transform -1 0 3336 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_151
timestamp 1598350056
transform -1 0 3288 0 -1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_351
timestamp 1598350056
transform -1 0 3256 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_338
timestamp 1598350056
transform 1 0 3160 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_702
timestamp 1598350056
transform -1 0 3160 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_715
timestamp 1598350056
transform -1 0 3016 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_269
timestamp 1598350056
transform 1 0 3064 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_127
timestamp 1598350056
transform 1 0 3016 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_272
timestamp 1598350056
transform -1 0 2968 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_362
timestamp 1598350056
transform -1 0 2920 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_361
timestamp 1598350056
transform 1 0 2824 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_128
timestamp 1598350056
transform 1 0 2632 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_125
timestamp 1598350056
transform 1 0 2776 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_473
timestamp 1598350056
transform 1 0 2728 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_366
timestamp 1598350056
transform 1 0 2680 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_440
timestamp 1598350056
transform -1 0 2504 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_290
timestamp 1598350056
transform -1 0 2632 0 -1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_218
timestamp 1598350056
transform -1 0 2600 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_678
timestamp 1598350056
transform 1 0 2504 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_124
timestamp 1598350056
transform -1 0 2456 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_756
timestamp 1598350056
transform -1 0 2408 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_122
timestamp 1598350056
transform 1 0 2312 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_757
timestamp 1598350056
transform 1 0 2264 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_791
timestamp 1598350056
transform -1 0 2168 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_437
timestamp 1598350056
transform -1 0 2264 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_755
timestamp 1598350056
transform 1 0 2168 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_792
timestamp 1598350056
transform -1 0 2120 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_192
timestamp 1598350056
transform -1 0 1976 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_363
timestamp 1598350056
transform 1 0 2024 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_359
timestamp 1598350056
transform -1 0 2024 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_191
timestamp 1598350056
transform 1 0 1880 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_187
timestamp 1598350056
transform 1 0 1832 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_348
timestamp 1598350056
transform 1 0 1784 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_454
timestamp 1598350056
transform 1 0 1608 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_263
timestamp 1598350056
transform 1 0 1704 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_188
timestamp 1598350056
transform 1 0 1576 0 -1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_648
timestamp 1598350056
transform 1 0 1736 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_644
timestamp 1598350056
transform 1 0 1656 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_372
timestamp 1598350056
transform -1 0 1448 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_182
timestamp 1598350056
transform 1 0 1496 0 -1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_465
timestamp 1598350056
transform 1 0 1528 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_446
timestamp 1598350056
transform -1 0 1496 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_418
timestamp 1598350056
transform 1 0 1352 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_787
timestamp 1598350056
transform 1 0 1304 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_600
timestamp 1598350056
transform 1 0 1256 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_190
timestamp 1598350056
transform -1 0 1208 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_97
timestamp 1598350056
transform 1 0 1128 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_99
timestamp 1598350056
transform 1 0 1048 0 -1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_344
timestamp 1598350056
transform -1 0 1256 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_540
timestamp 1598350056
transform -1 0 1128 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_183
timestamp 1598350056
transform 1 0 920 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_247
timestamp 1598350056
transform -1 0 1000 0 -1 2610
box -18 -6 52 210
use INVX1  INVX1_179
timestamp 1598350056
transform -1 0 920 0 -1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_456
timestamp 1598350056
transform 1 0 1000 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_439
timestamp 1598350056
transform 1 0 840 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_842
timestamp 1598350056
transform 1 0 792 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_850
timestamp 1598350056
transform -1 0 792 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_599
timestamp 1598350056
transform -1 0 648 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_830
timestamp 1598350056
transform -1 0 744 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_858
timestamp 1598350056
transform 1 0 648 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_598
timestamp 1598350056
transform -1 0 600 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_438
timestamp 1598350056
transform -1 0 552 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_279
timestamp 1598350056
transform -1 0 504 0 -1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_544
timestamp 1598350056
transform -1 0 472 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_724
timestamp 1598350056
transform -1 0 424 0 -1 2610
box -16 -6 64 210
use INVX1  INVX1_307
timestamp 1598350056
transform -1 0 376 0 -1 2610
box -18 -6 52 210
use NOR2X1  NOR2X1_714
timestamp 1598350056
transform 1 0 296 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_704
timestamp 1598350056
transform -1 0 296 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_374
timestamp 1598350056
transform -1 0 248 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_314
timestamp 1598350056
transform 1 0 8 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_322
timestamp 1598350056
transform 1 0 152 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_373
timestamp 1598350056
transform 1 0 104 0 -1 2610
box -16 -6 64 210
use NOR2X1  NOR2X1_317
timestamp 1598350056
transform 1 0 56 0 -1 2610
box -16 -6 64 210
use NAND2X1  NAND2X1_741
timestamp 1598350056
transform 1 0 5144 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_742
timestamp 1598350056
transform 1 0 5096 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_771
timestamp 1598350056
transform -1 0 5096 0 1 2210
box -16 -6 64 210
use FILL  FILL_12_1
timestamp 1598350056
transform 1 0 5192 0 1 2210
box -16 -6 32 210
use NAND2X1  NAND2X1_810
timestamp 1598350056
transform 1 0 5000 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_730
timestamp 1598350056
transform -1 0 5000 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_389
timestamp 1598350056
transform 1 0 4904 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_800
timestamp 1598350056
transform -1 0 4776 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_231
timestamp 1598350056
transform 1 0 4776 0 1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_578
timestamp 1598350056
transform -1 0 4904 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_385
timestamp 1598350056
transform 1 0 4808 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_739
timestamp 1598350056
transform 1 0 4648 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_568
timestamp 1598350056
transform 1 0 4600 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_728
timestamp 1598350056
transform -1 0 4600 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_161
timestamp 1598350056
transform -1 0 4728 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_648
timestamp 1598350056
transform -1 0 4520 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_273
timestamp 1598350056
transform 1 0 4520 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_264
timestamp 1598350056
transform 1 0 4440 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_291
timestamp 1598350056
transform 1 0 4408 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_276
timestamp 1598350056
transform -1 0 4408 0 1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_687
timestamp 1598350056
transform 1 0 4328 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_685
timestamp 1598350056
transform 1 0 4280 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_834
timestamp 1598350056
transform -1 0 4232 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_682
timestamp 1598350056
transform -1 0 4280 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_214
timestamp 1598350056
transform -1 0 4040 0 1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_511
timestamp 1598350056
transform -1 0 4184 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_681
timestamp 1598350056
transform 1 0 4088 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_574
timestamp 1598350056
transform 1 0 4040 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_779
timestamp 1598350056
transform 1 0 3928 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_516
timestamp 1598350056
transform 1 0 3880 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_21
timestamp 1598350056
transform 1 0 3976 0 1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_513
timestamp 1598350056
transform 1 0 3832 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_846
timestamp 1598350056
transform -1 0 3832 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_683
timestamp 1598350056
transform 1 0 3688 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_816
timestamp 1598350056
transform -1 0 3784 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_684
timestamp 1598350056
transform 1 0 3592 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_324
timestamp 1598350056
transform -1 0 3544 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_686
timestamp 1598350056
transform 1 0 3640 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_320
timestamp 1598350056
transform -1 0 3592 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_760
timestamp 1598350056
transform 1 0 3368 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_249
timestamp 1598350056
transform 1 0 3320 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_215
timestamp 1598350056
transform 1 0 3464 0 1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_65
timestamp 1598350056
transform 1 0 3416 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_112
timestamp 1598350056
transform -1 0 3320 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_332
timestamp 1598350056
transform -1 0 3224 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_111
timestamp 1598350056
transform -1 0 3272 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_138
timestamp 1598350056
transform -1 0 3096 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_9
timestamp 1598350056
transform -1 0 3128 0 1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_135
timestamp 1598350056
transform -1 0 3176 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_136
timestamp 1598350056
transform 1 0 3000 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_514
timestamp 1598350056
transform 1 0 2904 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_515
timestamp 1598350056
transform 1 0 2856 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_321
timestamp 1598350056
transform 1 0 2952 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_106
timestamp 1598350056
transform -1 0 2856 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_115
timestamp 1598350056
transform 1 0 2760 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_133
timestamp 1598350056
transform 1 0 2728 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_79
timestamp 1598350056
transform -1 0 2728 0 1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_139
timestamp 1598350056
transform -1 0 2696 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_554
timestamp 1598350056
transform 1 0 2600 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_67
timestamp 1598350056
transform -1 0 2600 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_313
timestamp 1598350056
transform -1 0 2568 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_177
timestamp 1598350056
transform 1 0 2504 0 1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_674
timestamp 1598350056
transform -1 0 2504 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_675
timestamp 1598350056
transform -1 0 2408 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_155
timestamp 1598350056
transform -1 0 2360 0 1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_760
timestamp 1598350056
transform -1 0 2456 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_137
timestamp 1598350056
transform 1 0 2280 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_646
timestamp 1598350056
transform -1 0 2184 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_607
timestamp 1598350056
transform -1 0 2280 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_390
timestamp 1598350056
transform -1 0 2232 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_132
timestamp 1598350056
transform 1 0 2040 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_608
timestamp 1598350056
transform -1 0 2008 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_29
timestamp 1598350056
transform -1 0 2040 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_101
timestamp 1598350056
transform 1 0 1928 0 1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_609
timestamp 1598350056
transform 1 0 2088 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_491
timestamp 1598350056
transform 1 0 1880 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_329
timestamp 1598350056
transform -1 0 1880 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_493
timestamp 1598350056
transform 1 0 1784 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_492
timestamp 1598350056
transform -1 0 1784 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_206
timestamp 1598350056
transform -1 0 1688 0 1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_205
timestamp 1598350056
transform -1 0 1736 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_203
timestamp 1598350056
transform -1 0 1656 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_266
timestamp 1598350056
transform 1 0 1528 0 1 2210
box -18 -6 52 210
use INVX1  INVX1_227
timestamp 1598350056
transform -1 0 1480 0 1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_455
timestamp 1598350056
transform 1 0 1560 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_577
timestamp 1598350056
transform -1 0 1528 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_563
timestamp 1598350056
transform -1 0 1448 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_753
timestamp 1598350056
transform -1 0 1304 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_570
timestamp 1598350056
transform -1 0 1400 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_388
timestamp 1598350056
transform 1 0 1304 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_553
timestamp 1598350056
transform -1 0 1256 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_550
timestamp 1598350056
transform -1 0 1208 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_565
timestamp 1598350056
transform -1 0 1160 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_549
timestamp 1598350056
transform -1 0 1112 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_220
timestamp 1598350056
transform 1 0 888 0 1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_569
timestamp 1598350056
transform -1 0 1064 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_794
timestamp 1598350056
transform 1 0 968 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_788
timestamp 1598350056
transform -1 0 968 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_167
timestamp 1598350056
transform 1 0 792 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_531
timestamp 1598350056
transform 1 0 840 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_564
timestamp 1598350056
transform -1 0 792 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_312
timestamp 1598350056
transform 1 0 648 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_292
timestamp 1598350056
transform -1 0 648 0 1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_551
timestamp 1598350056
transform -1 0 744 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_703
timestamp 1598350056
transform -1 0 616 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_761
timestamp 1598350056
transform 1 0 520 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_804
timestamp 1598350056
transform 1 0 472 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_800
timestamp 1598350056
transform -1 0 472 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_801
timestamp 1598350056
transform -1 0 424 0 1 2210
box -16 -6 64 210
use INVX1  INVX1_196
timestamp 1598350056
transform 1 0 344 0 1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_805
timestamp 1598350056
transform -1 0 344 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_324
timestamp 1598350056
transform 1 0 248 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_326
timestamp 1598350056
transform 1 0 200 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_325
timestamp 1598350056
transform -1 0 200 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_807
timestamp 1598350056
transform 1 0 104 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_811
timestamp 1598350056
transform 1 0 56 0 1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_808
timestamp 1598350056
transform -1 0 56 0 1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_379
timestamp 1598350056
transform 1 0 5128 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_770
timestamp 1598350056
transform 1 0 5080 0 -1 2210
box -16 -6 64 210
use FILL  FILL_11_2
timestamp 1598350056
transform -1 0 5208 0 -1 2210
box -16 -6 32 210
use FILL  FILL_11_1
timestamp 1598350056
transform -1 0 5192 0 -1 2210
box -16 -6 32 210
use NAND2X1  NAND2X1_812
timestamp 1598350056
transform 1 0 5032 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_537
timestamp 1598350056
transform -1 0 4936 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_766
timestamp 1598350056
transform -1 0 5032 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_829
timestamp 1598350056
transform -1 0 4984 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_729
timestamp 1598350056
transform 1 0 4840 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_536
timestamp 1598350056
transform 1 0 4792 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_533
timestamp 1598350056
transform 1 0 4744 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_532
timestamp 1598350056
transform -1 0 4744 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_854
timestamp 1598350056
transform 1 0 4648 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_566
timestamp 1598350056
transform 1 0 4600 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_567
timestamp 1598350056
transform 1 0 4552 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_539
timestamp 1598350056
transform 1 0 4456 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_535
timestamp 1598350056
transform -1 0 4456 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_221
timestamp 1598350056
transform 1 0 4376 0 -1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_753
timestamp 1598350056
transform -1 0 4552 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_590
timestamp 1598350056
transform -1 0 4328 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_534
timestamp 1598350056
transform -1 0 4248 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_119
timestamp 1598350056
transform 1 0 4248 0 -1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_591
timestamp 1598350056
transform -1 0 4376 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_326
timestamp 1598350056
transform 1 0 4152 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_236
timestamp 1598350056
transform 1 0 4120 0 -1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_152
timestamp 1598350056
transform -1 0 4120 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_667
timestamp 1598350056
transform 1 0 4024 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_680
timestamp 1598350056
transform -1 0 4024 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_151
timestamp 1598350056
transform 1 0 3928 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_306
timestamp 1598350056
transform -1 0 3928 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_141
timestamp 1598350056
transform 1 0 3848 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_643
timestamp 1598350056
transform -1 0 3800 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_538
timestamp 1598350056
transform -1 0 3752 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_649
timestamp 1598350056
transform 1 0 3656 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_512
timestamp 1598350056
transform -1 0 3848 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_655
timestamp 1598350056
transform -1 0 3656 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_327
timestamp 1598350056
transform 1 0 3512 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_595
timestamp 1598350056
transform 1 0 3560 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_660
timestamp 1598350056
transform -1 0 3512 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_49
timestamp 1598350056
transform 1 0 3336 0 -1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_441
timestamp 1598350056
transform 1 0 3416 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_250
timestamp 1598350056
transform -1 0 3416 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_211
timestamp 1598350056
transform 1 0 3288 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_315
timestamp 1598350056
transform -1 0 3192 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_172
timestamp 1598350056
transform 1 0 3240 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_318
timestamp 1598350056
transform -1 0 3240 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_343
timestamp 1598350056
transform -1 0 3112 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_843
timestamp 1598350056
transform 1 0 3016 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_118
timestamp 1598350056
transform -1 0 3144 0 -1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_251
timestamp 1598350056
transform 1 0 2968 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_330
timestamp 1598350056
transform -1 0 2968 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_105
timestamp 1598350056
transform 1 0 2872 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_331
timestamp 1598350056
transform -1 0 2872 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_145
timestamp 1598350056
transform -1 0 2824 0 -1 2210
box -18 -6 52 210
use NAND2X1  NAND2X1_349
timestamp 1598350056
transform 1 0 2744 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_545
timestamp 1598350056
transform -1 0 2664 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_208
timestamp 1598350056
transform 1 0 2712 0 -1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_524
timestamp 1598350056
transform -1 0 2712 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_45
timestamp 1598350056
transform -1 0 2520 0 -1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_116
timestamp 1598350056
transform 1 0 2568 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_216
timestamp 1598350056
transform -1 0 2568 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_117
timestamp 1598350056
transform 1 0 2440 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_123
timestamp 1598350056
transform -1 0 2440 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_606
timestamp 1598350056
transform 1 0 2344 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_294
timestamp 1598350056
transform -1 0 2344 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_310
timestamp 1598350056
transform 1 0 2200 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_94
timestamp 1598350056
transform 1 0 2168 0 -1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_295
timestamp 1598350056
transform -1 0 2296 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_335
timestamp 1598350056
transform -1 0 2168 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_189
timestamp 1598350056
transform -1 0 1992 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_28
timestamp 1598350056
transform -1 0 2072 0 -1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_481
timestamp 1598350056
transform -1 0 2120 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_188
timestamp 1598350056
transform -1 0 2040 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_498
timestamp 1598350056
transform -1 0 1944 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_309
timestamp 1598350056
transform 1 0 1800 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_501
timestamp 1598350056
transform 1 0 1848 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_355
timestamp 1598350056
transform -1 0 1800 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_369
timestamp 1598350056
transform -1 0 1752 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_370
timestamp 1598350056
transform -1 0 1704 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_543
timestamp 1598350056
transform -1 0 1656 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_72
timestamp 1598350056
transform -1 0 1560 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_166
timestamp 1598350056
transform 1 0 1464 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_445
timestamp 1598350056
transform -1 0 1608 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_169
timestamp 1598350056
transform 1 0 1416 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_530
timestamp 1598350056
transform -1 0 1320 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_170
timestamp 1598350056
transform -1 0 1416 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_548
timestamp 1598350056
transform 1 0 1320 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_337
timestamp 1598350056
transform 1 0 1224 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_371
timestamp 1598350056
transform -1 0 1224 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_165
timestamp 1598350056
transform -1 0 1144 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_223
timestamp 1598350056
transform -1 0 1176 0 -1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_168
timestamp 1598350056
transform -1 0 1096 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_184
timestamp 1598350056
transform -1 0 1048 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_533
timestamp 1598350056
transform -1 0 952 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_336
timestamp 1598350056
transform 1 0 952 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_532
timestamp 1598350056
transform -1 0 904 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_500
timestamp 1598350056
transform -1 0 856 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_552
timestamp 1598350056
transform -1 0 808 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_614
timestamp 1598350056
transform 1 0 712 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_754
timestamp 1598350056
transform 1 0 616 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_790
timestamp 1598350056
transform 1 0 664 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_542
timestamp 1598350056
transform -1 0 616 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_417
timestamp 1598350056
transform 1 0 520 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_237
timestamp 1598350056
transform -1 0 520 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_323
timestamp 1598350056
transform -1 0 424 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_793
timestamp 1598350056
transform -1 0 472 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_321
timestamp 1598350056
transform 1 0 328 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_320
timestamp 1598350056
transform -1 0 328 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_356
timestamp 1598350056
transform -1 0 280 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_354
timestamp 1598350056
transform 1 0 184 0 -1 2210
box -16 -6 64 210
use INVX1  INVX1_269
timestamp 1598350056
transform -1 0 184 0 -1 2210
box -18 -6 52 210
use NOR2X1  NOR2X1_806
timestamp 1598350056
transform -1 0 152 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_855
timestamp 1598350056
transform 1 0 56 0 -1 2210
box -16 -6 64 210
use NOR2X1  NOR2X1_812
timestamp 1598350056
transform -1 0 56 0 -1 2210
box -16 -6 64 210
use NAND2X1  NAND2X1_723
timestamp 1598350056
transform -1 0 5192 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_864
timestamp 1598350056
transform 1 0 5096 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_300
timestamp 1598350056
transform 1 0 5064 0 1 1810
box -18 -6 52 210
use FILL  FILL_10_1
timestamp 1598350056
transform 1 0 5192 0 1 1810
box -16 -6 32 210
use NAND2X1  NAND2X1_855
timestamp 1598350056
transform 1 0 4888 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_297
timestamp 1598350056
transform 1 0 4984 0 1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_774
timestamp 1598350056
transform -1 0 5064 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_765
timestamp 1598350056
transform 1 0 4936 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_856
timestamp 1598350056
transform 1 0 4840 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_738
timestamp 1598350056
transform 1 0 4792 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_740
timestamp 1598350056
transform -1 0 4792 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_307
timestamp 1598350056
transform 1 0 4696 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_308
timestamp 1598350056
transform 1 0 4648 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_250
timestamp 1598350056
transform 1 0 4568 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_11
timestamp 1598350056
transform 1 0 4536 0 1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_305
timestamp 1598350056
transform -1 0 4648 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_718
timestamp 1598350056
transform 1 0 4488 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_788
timestamp 1598350056
transform -1 0 4440 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_248
timestamp 1598350056
transform 1 0 4360 0 1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_645
timestamp 1598350056
transform -1 0 4488 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_714
timestamp 1598350056
transform 1 0 4312 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_668
timestamp 1598350056
transform 1 0 4216 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_669
timestamp 1598350056
transform 1 0 4264 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_720
timestamp 1598350056
transform 1 0 4168 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_575
timestamp 1598350056
transform 1 0 4120 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_405
timestamp 1598350056
transform -1 0 4120 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_840
timestamp 1598350056
transform 1 0 4024 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_851
timestamp 1598350056
transform -1 0 4024 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_777
timestamp 1598350056
transform 1 0 3928 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_803
timestamp 1598350056
transform 1 0 3880 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_796
timestamp 1598350056
transform 1 0 3832 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_783
timestamp 1598350056
transform 1 0 3784 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_780
timestamp 1598350056
transform 1 0 3688 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_744
timestamp 1598350056
transform 1 0 3736 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_336
timestamp 1598350056
transform -1 0 3640 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_600
timestamp 1598350056
transform 1 0 3544 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_311
timestamp 1598350056
transform -1 0 3688 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_602
timestamp 1598350056
transform 1 0 3496 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_601
timestamp 1598350056
transform -1 0 3496 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_312
timestamp 1598350056
transform 1 0 3416 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_33
timestamp 1598350056
transform 1 0 3336 0 1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_841
timestamp 1598350056
transform -1 0 3416 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_300
timestamp 1598350056
transform 1 0 3240 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_110
timestamp 1598350056
transform 1 0 3288 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_831
timestamp 1598350056
transform -1 0 3240 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_109
timestamp 1598350056
transform 1 0 3144 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_759
timestamp 1598350056
transform 1 0 3096 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_286
timestamp 1598350056
transform 1 0 3000 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_758
timestamp 1598350056
transform -1 0 3096 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_573
timestamp 1598350056
transform 1 0 2952 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_273
timestamp 1598350056
transform 1 0 2904 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_288
timestamp 1598350056
transform 1 0 2856 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_806
timestamp 1598350056
transform -1 0 2856 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_337
timestamp 1598350056
transform 1 0 2680 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_107
timestamp 1598350056
transform -1 0 2680 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_131
timestamp 1598350056
transform 1 0 2728 0 1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_743
timestamp 1598350056
transform -1 0 2808 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_283
timestamp 1598350056
transform 1 0 2552 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_270
timestamp 1598350056
transform 1 0 2600 0 1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_113
timestamp 1598350056
transform -1 0 2552 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_114
timestamp 1598350056
transform -1 0 2504 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_830
timestamp 1598350056
transform 1 0 2408 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_103
timestamp 1598350056
transform -1 0 2328 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_66
timestamp 1598350056
transform -1 0 2408 0 1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_108
timestamp 1598350056
transform -1 0 2376 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_134
timestamp 1598350056
transform 1 0 2152 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_150
timestamp 1598350056
transform -1 0 2232 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_285
timestamp 1598350056
transform -1 0 2152 0 1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_768
timestamp 1598350056
transform 1 0 2232 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_647
timestamp 1598350056
transform -1 0 2088 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_656
timestamp 1598350056
transform 1 0 1992 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_699
timestamp 1598350056
transform -1 0 1992 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_54
timestamp 1598350056
transform -1 0 2120 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_774
timestamp 1598350056
transform -1 0 1912 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_14
timestamp 1598350056
transform -1 0 1944 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_111
timestamp 1598350056
transform -1 0 1864 0 1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_309
timestamp 1598350056
transform 1 0 1784 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_335
timestamp 1598350056
transform -1 0 1736 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_225
timestamp 1598350056
transform -1 0 1640 0 1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_274
timestamp 1598350056
transform -1 0 1784 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_310
timestamp 1598350056
transform 1 0 1640 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_406
timestamp 1598350056
transform -1 0 1528 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_58
timestamp 1598350056
transform -1 0 1560 0 1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_534
timestamp 1598350056
transform -1 0 1608 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_405
timestamp 1598350056
transform -1 0 1480 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_536
timestamp 1598350056
transform -1 0 1432 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_272
timestamp 1598350056
transform 1 0 1304 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_149
timestamp 1598350056
transform -1 0 1384 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_222
timestamp 1598350056
transform -1 0 1256 0 1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_541
timestamp 1598350056
transform -1 0 1304 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_256
timestamp 1598350056
transform 1 0 1176 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_650
timestamp 1598350056
transform -1 0 1176 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_799
timestamp 1598350056
transform -1 0 1128 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_311
timestamp 1598350056
transform 1 0 984 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_24
timestamp 1598350056
transform 1 0 904 0 1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_567
timestamp 1598350056
transform -1 0 1080 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_535
timestamp 1598350056
transform -1 0 984 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_497
timestamp 1598350056
transform 1 0 824 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_615
timestamp 1598350056
transform -1 0 792 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_18
timestamp 1598350056
transform -1 0 904 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_69
timestamp 1598350056
transform 1 0 792 0 1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_118
timestamp 1598350056
transform 1 0 648 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_280
timestamp 1598350056
transform -1 0 600 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_633
timestamp 1598350056
transform -1 0 744 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_640
timestamp 1598350056
transform 1 0 600 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_279
timestamp 1598350056
transform 1 0 456 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_164
timestamp 1598350056
transform 1 0 376 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_305
timestamp 1598350056
transform -1 0 456 0 1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_284
timestamp 1598350056
transform -1 0 552 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_809
timestamp 1598350056
transform 1 0 328 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_802
timestamp 1598350056
transform -1 0 328 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_798
timestamp 1598350056
transform -1 0 280 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_319
timestamp 1598350056
transform -1 0 232 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_299
timestamp 1598350056
transform -1 0 88 0 1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_854
timestamp 1598350056
transform -1 0 184 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_856
timestamp 1598350056
transform 1 0 88 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_810
timestamp 1598350056
transform -1 0 56 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_863
timestamp 1598350056
transform 1 0 5128 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_689
timestamp 1598350056
transform -1 0 5128 0 -1 1810
box -16 -6 64 210
use FILL  FILL_9_2
timestamp 1598350056
transform -1 0 5208 0 -1 1810
box -16 -6 32 210
use FILL  FILL_9_1
timestamp 1598350056
transform -1 0 5192 0 -1 1810
box -16 -6 32 210
use NAND2X1  NAND2X1_724
timestamp 1598350056
transform 1 0 5032 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_688
timestamp 1598350056
transform 1 0 4984 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_353
timestamp 1598350056
transform -1 0 4984 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_727
timestamp 1598350056
transform -1 0 4936 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_731
timestamp 1598350056
transform 1 0 4840 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_691
timestamp 1598350056
transform 1 0 4792 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_264
timestamp 1598350056
transform -1 0 4792 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_726
timestamp 1598350056
transform 1 0 4696 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_811
timestamp 1598350056
transform 1 0 4648 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_808
timestamp 1598350056
transform 1 0 4600 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_605
timestamp 1598350056
transform -1 0 4600 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_603
timestamp 1598350056
transform -1 0 4552 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_604
timestamp 1598350056
transform 1 0 4456 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_322
timestamp 1598350056
transform -1 0 4456 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_406
timestamp 1598350056
transform 1 0 4360 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_721
timestamp 1598350056
transform 1 0 4312 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_734
timestamp 1598350056
transform -1 0 4312 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_325
timestamp 1598350056
transform -1 0 4264 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_784
timestamp 1598350056
transform 1 0 4168 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_323
timestamp 1598350056
transform 1 0 4120 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_527
timestamp 1598350056
transform 1 0 4072 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_654
timestamp 1598350056
transform -1 0 4072 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_547
timestamp 1598350056
transform -1 0 4024 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_703
timestamp 1598350056
transform -1 0 3976 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_542
timestamp 1598350056
transform 1 0 3880 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_312
timestamp 1598350056
transform 1 0 3832 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_661
timestamp 1598350056
transform -1 0 3832 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_245
timestamp 1598350056
transform 1 0 3736 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_280
timestamp 1598350056
transform -1 0 3736 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_284
timestamp 1598350056
transform 1 0 3640 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_285
timestamp 1598350056
transform -1 0 3544 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_279
timestamp 1598350056
transform -1 0 3640 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_281
timestamp 1598350056
transform 1 0 3544 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_594
timestamp 1598350056
transform 1 0 3400 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_282
timestamp 1598350056
transform 1 0 3448 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_653
timestamp 1598350056
transform 1 0 3352 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_807
timestamp 1598350056
transform 1 0 3304 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_805
timestamp 1598350056
transform 1 0 3256 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_316
timestamp 1598350056
transform 1 0 3176 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_162
timestamp 1598350056
transform 1 0 3224 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_308
timestamp 1598350056
transform 1 0 3144 0 -1 1810
box -18 -6 52 210
use NAND2X1  NAND2X1_352
timestamp 1598350056
transform -1 0 3096 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_287
timestamp 1598350056
transform -1 0 3048 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_792
timestamp 1598350056
transform 1 0 3096 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_357
timestamp 1598350056
transform -1 0 3000 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_53
timestamp 1598350056
transform -1 0 2952 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_95
timestamp 1598350056
transform -1 0 2872 0 -1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_389
timestamp 1598350056
transform -1 0 2920 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_246
timestamp 1598350056
transform -1 0 2840 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_342
timestamp 1598350056
transform 1 0 2744 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_153
timestamp 1598350056
transform 1 0 2696 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_248
timestamp 1598350056
transform 1 0 2648 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_247
timestamp 1598350056
transform 1 0 2600 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_187
timestamp 1598350056
transform -1 0 2600 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_15
timestamp 1598350056
transform 1 0 2504 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_150
timestamp 1598350056
transform 1 0 2456 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_674
timestamp 1598350056
transform -1 0 2456 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_475
timestamp 1598350056
transform 1 0 2264 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_675
timestamp 1598350056
transform -1 0 2408 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_773
timestamp 1598350056
transform -1 0 2360 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_294
timestamp 1598350056
transform 1 0 2184 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_171
timestamp 1598350056
transform 1 0 2152 0 -1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_772
timestamp 1598350056
transform -1 0 2264 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_186
timestamp 1598350056
transform -1 0 2152 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_78
timestamp 1598350056
transform 1 0 2008 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_767
timestamp 1598350056
transform 1 0 2056 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_652
timestamp 1598350056
transform 1 0 1960 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_204
timestamp 1598350056
transform -1 0 1880 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_385
timestamp 1598350056
transform 1 0 1784 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_1
timestamp 1598350056
transform 1 0 1880 0 -1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_79
timestamp 1598350056
transform -1 0 1960 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_568
timestamp 1598350056
transform -1 0 1784 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_566
timestamp 1598350056
transform 1 0 1688 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_212
timestamp 1598350056
transform 1 0 1640 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_211
timestamp 1598350056
transform 1 0 1592 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_71
timestamp 1598350056
transform -1 0 1512 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_116
timestamp 1598350056
transform -1 0 1544 0 -1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_220
timestamp 1598350056
transform -1 0 1592 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_537
timestamp 1598350056
transform 1 0 1416 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_173
timestamp 1598350056
transform -1 0 1416 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_255
timestamp 1598350056
transform 1 0 1224 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_699
timestamp 1598350056
transform 1 0 1320 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_175
timestamp 1598350056
transform 1 0 1272 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_853
timestamp 1598350056
transform 1 0 1176 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_748
timestamp 1598350056
transform 1 0 1128 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_539
timestamp 1598350056
transform 1 0 1080 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_789
timestamp 1598350056
transform 1 0 984 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_278
timestamp 1598350056
transform -1 0 984 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_277
timestamp 1598350056
transform -1 0 936 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_538
timestamp 1598350056
transform 1 0 1032 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_171
timestamp 1598350056
transform -1 0 888 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_436
timestamp 1598350056
transform -1 0 840 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_174
timestamp 1598350056
transform 1 0 744 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_172
timestamp 1598350056
transform -1 0 744 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_431
timestamp 1598350056
transform 1 0 600 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_434
timestamp 1598350056
transform 1 0 648 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_287
timestamp 1598350056
transform 1 0 552 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_690
timestamp 1598350056
transform -1 0 504 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_691
timestamp 1598350056
transform 1 0 504 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_634
timestamp 1598350056
transform -1 0 456 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_288
timestamp 1598350056
transform -1 0 408 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_290
timestamp 1598350056
transform -1 0 312 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_821
timestamp 1598350056
transform -1 0 264 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_160
timestamp 1598350056
transform -1 0 216 0 -1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_334
timestamp 1598350056
transform 1 0 312 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_134
timestamp 1598350056
transform -1 0 184 0 -1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_857
timestamp 1598350056
transform -1 0 152 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_863
timestamp 1598350056
transform -1 0 104 0 -1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_864
timestamp 1598350056
transform -1 0 56 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_853
timestamp 1598350056
transform 1 0 5080 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_700
timestamp 1598350056
transform -1 0 5176 0 1 1410
box -16 -6 64 210
use FILL  FILL_8_2
timestamp 1598350056
transform 1 0 5192 0 1 1410
box -16 -6 32 210
use FILL  FILL_8_1
timestamp 1598350056
transform 1 0 5176 0 1 1410
box -16 -6 32 210
use NAND2X1  NAND2X1_710
timestamp 1598350056
transform 1 0 4984 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_794
timestamp 1598350056
transform -1 0 4936 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_701
timestamp 1598350056
transform -1 0 5080 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_690
timestamp 1598350056
transform -1 0 4984 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_188
timestamp 1598350056
transform -1 0 4888 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_711
timestamp 1598350056
transform 1 0 4744 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_189
timestamp 1598350056
transform -1 0 4840 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_520
timestamp 1598350056
transform 1 0 4648 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_168
timestamp 1598350056
transform -1 0 4648 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_519
timestamp 1598350056
transform 1 0 4696 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_518
timestamp 1598350056
transform 1 0 4552 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_185
timestamp 1598350056
transform 1 0 4456 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_278
timestamp 1598350056
transform 1 0 4376 0 1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_165
timestamp 1598350056
transform 1 0 4504 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_166
timestamp 1598350056
transform 1 0 4408 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_169
timestamp 1598350056
transform -1 0 4376 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_170
timestamp 1598350056
transform -1 0 4328 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_57
timestamp 1598350056
transform -1 0 4232 0 1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_167
timestamp 1598350056
transform 1 0 4232 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_858
timestamp 1598350056
transform 1 0 4152 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_775
timestamp 1598350056
transform -1 0 4152 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_265
timestamp 1598350056
transform -1 0 4056 0 1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_46
timestamp 1598350056
transform 1 0 4056 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_650
timestamp 1598350056
transform 1 0 3976 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_442
timestamp 1598350056
transform -1 0 3976 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_444
timestamp 1598350056
transform -1 0 3896 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_183
timestamp 1598350056
transform -1 0 3928 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_443
timestamp 1598350056
transform 1 0 3800 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_286
timestamp 1598350056
transform 1 0 3768 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_185
timestamp 1598350056
transform -1 0 3768 0 1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_469
timestamp 1598350056
transform 1 0 3688 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_388
timestamp 1598350056
transform -1 0 3688 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_41
timestamp 1598350056
transform -1 0 3640 0 1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_176
timestamp 1598350056
transform -1 0 3608 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_265
timestamp 1598350056
transform 1 0 3512 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_641
timestamp 1598350056
transform 1 0 3464 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_390
timestamp 1598350056
transform -1 0 3464 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_102
timestamp 1598350056
transform -1 0 3416 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_126
timestamp 1598350056
transform -1 0 3384 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_93
timestamp 1598350056
transform -1 0 3352 0 1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_474
timestamp 1598350056
transform -1 0 3192 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_181
timestamp 1598350056
transform -1 0 3272 0 1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_129
timestamp 1598350056
transform 1 0 3272 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_267
timestamp 1598350056
transform 1 0 3192 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_842
timestamp 1598350056
transform -1 0 3144 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_100
timestamp 1598350056
transform -1 0 3096 0 1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_190
timestamp 1598350056
transform -1 0 3064 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_266
timestamp 1598350056
transform 1 0 2968 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_850
timestamp 1598350056
transform -1 0 2888 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_98
timestamp 1598350056
transform 1 0 2888 0 1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_153
timestamp 1598350056
transform -1 0 2968 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_191
timestamp 1598350056
transform -1 0 2840 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_698
timestamp 1598350056
transform -1 0 2744 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_124
timestamp 1598350056
transform 1 0 2664 0 1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_192
timestamp 1598350056
transform -1 0 2792 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_709
timestamp 1598350056
transform 1 0 2616 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_183
timestamp 1598350056
transform 1 0 2568 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_263
timestamp 1598350056
transform 1 0 2520 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_561
timestamp 1598350056
transform -1 0 2520 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_117
timestamp 1598350056
transform -1 0 2376 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_610
timestamp 1598350056
transform 1 0 2280 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_558
timestamp 1598350056
transform -1 0 2472 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_225
timestamp 1598350056
transform 1 0 2376 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_346
timestamp 1598350056
transform 1 0 2232 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_87
timestamp 1598350056
transform -1 0 2136 0 1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_440
timestamp 1598350056
transform -1 0 2232 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_468
timestamp 1598350056
transform -1 0 2184 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_266
timestamp 1598350056
transform 1 0 1960 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_292
timestamp 1598350056
transform -1 0 2104 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_612
timestamp 1598350056
transform 1 0 2008 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_786
timestamp 1598350056
transform 1 0 1864 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_488
timestamp 1598350056
transform -1 0 1864 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_275
timestamp 1598350056
transform -1 0 1816 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_262
timestamp 1598350056
transform 1 0 1912 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_487
timestamp 1598350056
transform 1 0 1672 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_489
timestamp 1598350056
transform -1 0 1768 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_557
timestamp 1598350056
transform 1 0 1624 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_73
timestamp 1598350056
transform -1 0 1624 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_221
timestamp 1598350056
transform 1 0 1448 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_47
timestamp 1598350056
transform 1 0 1544 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_104
timestamp 1598350056
transform 1 0 1416 0 1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_734
timestamp 1598350056
transform 1 0 1496 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_150
timestamp 1598350056
transform 1 0 1368 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_63
timestamp 1598350056
transform -1 0 1336 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_8
timestamp 1598350056
transform -1 0 1368 0 1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_751
timestamp 1598350056
transform -1 0 1288 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_52
timestamp 1598350056
transform -1 0 1240 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_13
timestamp 1598350056
transform 1 0 1096 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_230
timestamp 1598350056
transform -1 0 1096 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_641
timestamp 1598350056
transform -1 0 1192 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_229
timestamp 1598350056
transform 1 0 952 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_314
timestamp 1598350056
transform 1 0 920 0 1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_231
timestamp 1598350056
transform -1 0 1048 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_843
timestamp 1598350056
transform 1 0 872 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_108
timestamp 1598350056
transform -1 0 872 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_623
timestamp 1598350056
transform -1 0 824 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_442
timestamp 1598350056
transform -1 0 776 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_289
timestamp 1598350056
transform 1 0 552 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_184
timestamp 1598350056
transform -1 0 728 0 1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_444
timestamp 1598350056
transform 1 0 648 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_333
timestamp 1598350056
transform 1 0 600 0 1 1410
box -16 -6 64 210
use INVX1  INVX1_303
timestamp 1598350056
transform -1 0 552 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_143
timestamp 1598350056
transform -1 0 472 0 1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_795
timestamp 1598350056
transform -1 0 520 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_776
timestamp 1598350056
transform 1 0 392 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_238
timestamp 1598350056
transform 1 0 296 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_281
timestamp 1598350056
transform 1 0 248 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_822
timestamp 1598350056
transform 1 0 200 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_241
timestamp 1598350056
transform 1 0 344 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_362
timestamp 1598350056
transform -1 0 152 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_365
timestamp 1598350056
transform 1 0 56 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_835
timestamp 1598350056
transform 1 0 152 0 1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_866
timestamp 1598350056
transform -1 0 56 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_560
timestamp 1598350056
transform 1 0 5160 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_722
timestamp 1598350056
transform -1 0 5160 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_559
timestamp 1598350056
transform 1 0 5064 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_787
timestamp 1598350056
transform -1 0 4968 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_517
timestamp 1598350056
transform 1 0 5016 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_498
timestamp 1598350056
transform 1 0 4968 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_804
timestamp 1598350056
transform -1 0 4920 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_795
timestamp 1598350056
transform 1 0 4776 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_692
timestamp 1598350056
transform 1 0 4824 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_164
timestamp 1598350056
transform 1 0 4728 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_776
timestamp 1598350056
transform 1 0 4632 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_833
timestamp 1598350056
transform 1 0 4584 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_785
timestamp 1598350056
transform 1 0 4536 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_495
timestamp 1598350056
transform 1 0 4680 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_790
timestamp 1598350056
transform 1 0 4456 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_233
timestamp 1598350056
transform 1 0 4504 0 -1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_716
timestamp 1598350056
transform 1 0 4408 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_91
timestamp 1598350056
transform 1 0 4360 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_865
timestamp 1598350056
transform 1 0 4312 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_862
timestamp 1598350056
transform 1 0 4216 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_488
timestamp 1598350056
transform 1 0 4264 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_552
timestamp 1598350056
transform -1 0 4216 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_543
timestamp 1598350056
transform 1 0 4088 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_370
timestamp 1598350056
transform 1 0 4040 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_200
timestamp 1598350056
transform 1 0 4136 0 -1 1410
box -18 -6 52 210
use NAND2X1  NAND2X1_640
timestamp 1598350056
transform 1 0 3880 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_304
timestamp 1598350056
transform 1 0 3960 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_71
timestamp 1598350056
transform 1 0 3928 0 -1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_369
timestamp 1598350056
transform 1 0 3992 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_438
timestamp 1598350056
transform 1 0 3832 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_439
timestamp 1598350056
transform -1 0 3784 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_177
timestamp 1598350056
transform -1 0 3832 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_301
timestamp 1598350056
transform -1 0 3736 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_180
timestamp 1598350056
transform 1 0 3640 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_793
timestamp 1598350056
transform 1 0 3592 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_860
timestamp 1598350056
transform -1 0 3592 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_861
timestamp 1598350056
transform 1 0 3496 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_182
timestamp 1598350056
transform -1 0 3496 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_392
timestamp 1598350056
transform -1 0 3448 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_277
timestamp 1598350056
transform 1 0 3352 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_633
timestamp 1598350056
transform 1 0 3304 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_70
timestamp 1598350056
transform -1 0 3208 0 -1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_118
timestamp 1598350056
transform 1 0 3256 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_278
timestamp 1598350056
transform -1 0 3256 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_404
timestamp 1598350056
transform 1 0 3128 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_168
timestamp 1598350056
transform 1 0 3096 0 -1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_123
timestamp 1598350056
transform -1 0 3096 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_786
timestamp 1598350056
transform 1 0 3000 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_396
timestamp 1598350056
transform 1 0 2952 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_395
timestamp 1598350056
transform 1 0 2808 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_401
timestamp 1598350056
transform -1 0 2952 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_402
timestamp 1598350056
transform -1 0 2904 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_164
timestamp 1598350056
transform 1 0 2776 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_256
timestamp 1598350056
transform 1 0 2744 0 -1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_10
timestamp 1598350056
transform 1 0 2696 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_9
timestamp 1598350056
transform 1 0 2648 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_494
timestamp 1598350056
transform -1 0 2504 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_397
timestamp 1598350056
transform -1 0 2648 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_82
timestamp 1598350056
transform 1 0 2552 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_315
timestamp 1598350056
transform -1 0 2552 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_572
timestamp 1598350056
transform 1 0 2408 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_262
timestamp 1598350056
transform 1 0 2312 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_71
timestamp 1598350056
transform 1 0 2360 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_83
timestamp 1598350056
transform -1 0 2312 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_318
timestamp 1598350056
transform -1 0 2264 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_316
timestamp 1598350056
transform -1 0 2216 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_80
timestamp 1598350056
transform 1 0 2120 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_84
timestamp 1598350056
transform 1 0 2024 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_437
timestamp 1598350056
transform 1 0 1976 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_267
timestamp 1598350056
transform 1 0 1928 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_81
timestamp 1598350056
transform -1 0 2120 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_361
timestamp 1598350056
transform -1 0 1800 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_129
timestamp 1598350056
transform -1 0 1832 0 -1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_283
timestamp 1598350056
transform 1 0 1880 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_159
timestamp 1598350056
transform -1 0 1880 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_447
timestamp 1598350056
transform 1 0 1656 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_62
timestamp 1598350056
transform 1 0 1576 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_125
timestamp 1598350056
transform 1 0 1624 0 -1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_420
timestamp 1598350056
transform 1 0 1704 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_265
timestamp 1598350056
transform -1 0 1528 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_327
timestamp 1598350056
transform 1 0 1528 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_264
timestamp 1598350056
transform 1 0 1432 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_750
timestamp 1598350056
transform 1 0 1336 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_7
timestamp 1598350056
transform -1 0 1304 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_92
timestamp 1598350056
transform -1 0 1336 0 -1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_749
timestamp 1598350056
transform 1 0 1384 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_106
timestamp 1598350056
transform 1 0 1176 0 -1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_228
timestamp 1598350056
transform -1 0 1256 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_193
timestamp 1598350056
transform 1 0 1128 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_341
timestamp 1598350056
transform 1 0 1080 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_616
timestamp 1598350056
transform 1 0 1032 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_621
timestamp 1598350056
transform 1 0 984 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_622
timestamp 1598350056
transform 1 0 936 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_624
timestamp 1598350056
transform 1 0 888 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_617
timestamp 1598350056
transform 1 0 840 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_65
timestamp 1598350056
transform -1 0 840 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_31
timestamp 1598350056
transform -1 0 808 0 -1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_827
timestamp 1598350056
transform -1 0 776 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_689
timestamp 1598350056
transform -1 0 728 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_132
timestamp 1598350056
transform -1 0 632 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_148
timestamp 1598350056
transform -1 0 600 0 -1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_688
timestamp 1598350056
transform 1 0 632 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_364
timestamp 1598350056
transform -1 0 568 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_412
timestamp 1598350056
transform -1 0 488 0 -1 1410
box -16 -6 64 210
use INVX1  INVX1_310
timestamp 1598350056
transform -1 0 520 0 -1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_785
timestamp 1598350056
transform -1 0 440 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_282
timestamp 1598350056
transform 1 0 248 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_286
timestamp 1598350056
transform 1 0 344 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_285
timestamp 1598350056
transform 1 0 296 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_838
timestamp 1598350056
transform 1 0 200 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_367
timestamp 1598350056
transform -1 0 56 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_366
timestamp 1598350056
transform -1 0 104 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_852
timestamp 1598350056
transform 1 0 152 0 -1 1410
box -16 -6 64 210
use NOR2X1  NOR2X1_839
timestamp 1598350056
transform 1 0 104 0 -1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_866
timestamp 1598350056
transform 1 0 5160 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_733
timestamp 1598350056
transform 1 0 5128 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_835
timestamp 1598350056
transform 1 0 5080 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_839
timestamp 1598350056
transform -1 0 5112 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_238
timestamp 1598350056
transform 1 0 5176 0 1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_380
timestamp 1598350056
transform -1 0 5160 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_852
timestamp 1598350056
transform 1 0 5016 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_836
timestamp 1598350056
transform 1 0 4968 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_821
timestamp 1598350056
transform 1 0 5032 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_822
timestamp 1598350056
transform -1 0 5032 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_525
timestamp 1598350056
transform -1 0 4984 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_484
timestamp 1598350056
transform 1 0 4888 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_823
timestamp 1598350056
transform -1 0 4968 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_486
timestamp 1598350056
transform -1 0 4888 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_706
timestamp 1598350056
transform -1 0 4792 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_546
timestamp 1598350056
transform -1 0 4872 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_705
timestamp 1598350056
transform -1 0 4824 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_717
timestamp 1598350056
transform 1 0 4728 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_485
timestamp 1598350056
transform -1 0 4840 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_824
timestamp 1598350056
transform -1 0 4920 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_713
timestamp 1598350056
transform -1 0 4744 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_483
timestamp 1598350056
transform -1 0 4648 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_254
timestamp 1598350056
transform -1 0 4600 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_501
timestamp 1598350056
transform -1 0 4728 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_499
timestamp 1598350056
transform -1 0 4600 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_91
timestamp 1598350056
transform -1 0 4680 0 -1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_252
timestamp 1598350056
transform -1 0 4696 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_526
timestamp 1598350056
transform -1 0 4648 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_614
timestamp 1598350056
transform 1 0 4360 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_500
timestamp 1598350056
transform 1 0 4504 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_844
timestamp 1598350056
transform 1 0 4408 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_754
timestamp 1598350056
transform 1 0 4504 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_253
timestamp 1598350056
transform 1 0 4456 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_482
timestamp 1598350056
transform -1 0 4456 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_496
timestamp 1598350056
transform 1 0 4456 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_615
timestamp 1598350056
transform -1 0 4408 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_620
timestamp 1598350056
transform 1 0 4264 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_623
timestamp 1598350056
transform 1 0 4312 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_778
timestamp 1598350056
transform 1 0 4264 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_613
timestamp 1598350056
transform -1 0 4360 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_528
timestamp 1598350056
transform -1 0 4264 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_497
timestamp 1598350056
transform 1 0 4216 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_242
timestamp 1598350056
transform -1 0 4168 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_241
timestamp 1598350056
transform 1 0 4072 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_489
timestamp 1598350056
transform 1 0 4024 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_244
timestamp 1598350056
transform -1 0 4056 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_17
timestamp 1598350056
transform 1 0 4136 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_37
timestamp 1598350056
transform 1 0 4104 0 -1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_238
timestamp 1598350056
transform 1 0 4168 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_617
timestamp 1598350056
transform 1 0 4168 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_371
timestamp 1598350056
transform -1 0 4104 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_374
timestamp 1598350056
transform 1 0 3928 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_478
timestamp 1598350056
transform -1 0 3928 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_458
timestamp 1598350056
transform 1 0 3912 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_487
timestamp 1598350056
transform 1 0 3976 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_693
timestamp 1598350056
transform -1 0 3880 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_372
timestamp 1598350056
transform -1 0 4008 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_291
timestamp 1598350056
transform 1 0 3864 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_634
timestamp 1598350056
transform 1 0 3816 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_334
timestamp 1598350056
transform 1 0 3672 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_373
timestamp 1598350056
transform -1 0 3832 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_237
timestamp 1598350056
transform 1 0 3736 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_134
timestamp 1598350056
transform 1 0 3688 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_234
timestamp 1598350056
transform -1 0 3816 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_233
timestamp 1598350056
transform 1 0 3720 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_544
timestamp 1598350056
transform -1 0 3688 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_97
timestamp 1598350056
transform -1 0 3608 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_550
timestamp 1598350056
transform -1 0 3624 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_464
timestamp 1598350056
transform 1 0 3528 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_19
timestamp 1598350056
transform 1 0 3608 0 1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_89
timestamp 1598350056
transform 1 0 3512 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_290
timestamp 1598350056
transform 1 0 3624 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_457
timestamp 1598350056
transform 1 0 3464 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_477
timestamp 1598350056
transform 1 0 3416 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_564
timestamp 1598350056
transform 1 0 3368 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_551
timestamp 1598350056
transform -1 0 3368 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_471
timestamp 1598350056
transform -1 0 3528 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_772
timestamp 1598350056
transform 1 0 3352 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_35
timestamp 1598350056
transform 1 0 3400 0 -1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_103
timestamp 1598350056
transform -1 0 3480 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_445
timestamp 1598350056
transform -1 0 3320 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_455
timestamp 1598350056
transform 1 0 3176 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_768
timestamp 1598350056
transform 1 0 3304 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_465
timestamp 1598350056
transform 1 0 3224 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_456
timestamp 1598350056
transform 1 0 3176 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_170
timestamp 1598350056
transform 1 0 3144 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_23
timestamp 1598350056
transform 1 0 3272 0 -1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_368
timestamp 1598350056
transform 1 0 3224 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_74
timestamp 1598350056
transform -1 0 3048 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_400
timestamp 1598350056
transform -1 0 3128 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_165
timestamp 1598350056
transform -1 0 3080 0 -1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_92
timestamp 1598350056
transform -1 0 3144 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_184
timestamp 1598350056
transform 1 0 3048 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_393
timestamp 1598350056
transform 1 0 3128 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_403
timestamp 1598350056
transform -1 0 3048 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_270
timestamp 1598350056
transform -1 0 2920 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_75
timestamp 1598350056
transform 1 0 2824 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_80
timestamp 1598350056
transform 1 0 2952 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_56
timestamp 1598350056
transform -1 0 2952 0 1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_76
timestamp 1598350056
transform 1 0 2952 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_394
timestamp 1598350056
transform 1 0 2904 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_236
timestamp 1598350056
transform 1 0 2856 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_38
timestamp 1598350056
transform 1 0 2808 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_198
timestamp 1598350056
transform 1 0 2776 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_181
timestamp 1598350056
transform 1 0 2632 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_399
timestamp 1598350056
transform 1 0 2712 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_179
timestamp 1598350056
transform -1 0 2776 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_271
timestamp 1598350056
transform -1 0 2728 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_398
timestamp 1598350056
transform -1 0 2808 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_756
timestamp 1598350056
transform -1 0 2712 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_791
timestamp 1598350056
transform 1 0 2616 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_540
timestamp 1598350056
transform 1 0 2584 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_269
timestamp 1598350056
transform -1 0 2584 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_268
timestamp 1598350056
transform 1 0 2456 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_757
timestamp 1598350056
transform 1 0 2568 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_127
timestamp 1598350056
transform 1 0 2504 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_72
timestamp 1598350056
transform 1 0 2536 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_25
timestamp 1598350056
transform 1 0 2456 0 -1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_49
timestamp 1598350056
transform -1 0 2536 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_203
timestamp 1598350056
transform 1 0 2408 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_384
timestamp 1598350056
transform 1 0 2312 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_119
timestamp 1598350056
transform -1 0 2424 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_55
timestamp 1598350056
transform -1 0 2376 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_34
timestamp 1598350056
transform -1 0 2456 0 -1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_72
timestamp 1598350056
transform 1 0 2360 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_178
timestamp 1598350056
transform -1 0 2312 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_296
timestamp 1598350056
transform -1 0 2328 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_297
timestamp 1598350056
transform -1 0 2232 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_90
timestamp 1598350056
transform -1 0 2184 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_43
timestamp 1598350056
transform 1 0 2184 0 1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_383
timestamp 1598350056
transform -1 0 2264 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_119
timestamp 1598350056
transform 1 0 2136 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_55
timestamp 1598350056
transform 1 0 2232 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_57
timestamp 1598350056
transform 1 0 2088 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_347
timestamp 1598350056
transform -1 0 2056 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_236
timestamp 1598350056
transform -1 0 2008 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_92
timestamp 1598350056
transform -1 0 2136 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_102
timestamp 1598350056
transform 1 0 1992 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_137
timestamp 1598350056
transform -1 0 2088 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_13
timestamp 1598350056
transform -1 0 1992 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_46
timestamp 1598350056
transform 1 0 1928 0 -1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_606
timestamp 1598350056
transform -1 0 2088 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_360
timestamp 1598350056
transform -1 0 1960 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_276
timestamp 1598350056
transform -1 0 1848 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_611
timestamp 1598350056
transform -1 0 1800 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_773
timestamp 1598350056
transform -1 0 1928 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_99
timestamp 1598350056
transform -1 0 1848 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_101
timestamp 1598350056
transform -1 0 1800 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_251
timestamp 1598350056
transform 1 0 1880 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_306
timestamp 1598350056
transform 1 0 1848 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_27
timestamp 1598350056
transform -1 0 1880 0 -1 1010
box -18 -6 52 210
use NAND2X1  NAND2X1_93
timestamp 1598350056
transform 1 0 1608 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_9
timestamp 1598350056
transform -1 0 1752 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_224
timestamp 1598350056
transform 1 0 1576 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_60
timestamp 1598350056
transform 1 0 1624 0 -1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_77
timestamp 1598350056
transform 1 0 1704 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_6
timestamp 1598350056
transform -1 0 1704 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_39
timestamp 1598350056
transform 1 0 1656 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_98
timestamp 1598350056
transform 1 0 1576 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_194
timestamp 1598350056
transform 1 0 1528 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_113
timestamp 1598350056
transform -1 0 1448 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_96
timestamp 1598350056
transform 1 0 1528 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_94
timestamp 1598350056
transform 1 0 1480 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_30
timestamp 1598350056
transform -1 0 1528 0 1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_16
timestamp 1598350056
transform 1 0 1448 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_133
timestamp 1598350056
transform 1 0 1432 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_292
timestamp 1598350056
transform -1 0 1352 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_669
timestamp 1598350056
transform -1 0 1304 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_529
timestamp 1598350056
transform -1 0 1384 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_107
timestamp 1598350056
transform -1 0 1400 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_618
timestamp 1598350056
transform -1 0 1432 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_721
timestamp 1598350056
transform 1 0 1288 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_720
timestamp 1598350056
transform -1 0 1288 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_200
timestamp 1598350056
transform 1 0 1208 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_667
timestamp 1598350056
transform -1 0 1160 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_518
timestamp 1598350056
transform 1 0 1192 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_490
timestamp 1598350056
transform 1 0 1144 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_218
timestamp 1598350056
transform 1 0 1112 0 -1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_185
timestamp 1598350056
transform -1 0 1208 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_668
timestamp 1598350056
transform 1 0 1064 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_619
timestamp 1598350056
transform -1 0 1112 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_517
timestamp 1598350056
transform 1 0 936 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_642
timestamp 1598350056
transform 1 0 1016 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_254
timestamp 1598350056
transform -1 0 1064 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_22
timestamp 1598350056
transform -1 0 936 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_51
timestamp 1598350056
transform 1 0 888 0 -1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_68
timestamp 1598350056
transform -1 0 1032 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_559
timestamp 1598350056
transform -1 0 1016 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_520
timestamp 1598350056
transform 1 0 920 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_69
timestamp 1598350056
transform 1 0 856 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_114
timestamp 1598350056
transform 1 0 808 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_524
timestamp 1598350056
transform -1 0 808 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_519
timestamp 1598350056
transform 1 0 760 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_226
timestamp 1598350056
transform 1 0 856 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_158
timestamp 1598350056
transform -1 0 760 0 -1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_545
timestamp 1598350056
transform -1 0 760 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_350
timestamp 1598350056
transform -1 0 856 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_613
timestamp 1598350056
transform 1 0 616 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_441
timestamp 1598350056
transform -1 0 616 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_528
timestamp 1598350056
transform -1 0 728 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_527
timestamp 1598350056
transform -1 0 632 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_110
timestamp 1598350056
transform -1 0 584 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_620
timestamp 1598350056
transform 1 0 664 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_547
timestamp 1598350056
transform -1 0 680 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_338
timestamp 1598350056
transform -1 0 520 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_91
timestamp 1598350056
transform -1 0 472 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_413
timestamp 1598350056
transform -1 0 424 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_358
timestamp 1598350056
transform -1 0 536 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_351
timestamp 1598350056
transform 1 0 440 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_443
timestamp 1598350056
transform -1 0 568 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_775
timestamp 1598350056
transform 1 0 392 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_826
timestamp 1598350056
transform -1 0 248 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_109
timestamp 1598350056
transform -1 0 392 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_15
timestamp 1598350056
transform 1 0 296 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_291
timestamp 1598350056
transform -1 0 296 0 -1 1010
box -16 -6 64 210
use INVX1  INVX1_176
timestamp 1598350056
transform -1 0 376 0 1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_462
timestamp 1598350056
transform 1 0 296 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_461
timestamp 1598350056
transform -1 0 296 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_410
timestamp 1598350056
transform 1 0 200 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_363
timestamp 1598350056
transform 1 0 8 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_245
timestamp 1598350056
transform 1 0 104 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_823
timestamp 1598350056
transform 1 0 56 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_411
timestamp 1598350056
transform 1 0 152 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_825
timestamp 1598350056
transform -1 0 152 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_824
timestamp 1598350056
transform -1 0 104 0 -1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_837
timestamp 1598350056
transform -1 0 200 0 1 1010
box -16 -6 64 210
use NOR2X1  NOR2X1_836
timestamp 1598350056
transform -1 0 56 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_579
timestamp 1598350056
transform 1 0 5096 0 1 610
box -16 -6 64 210
use INVX1  INVX1_282
timestamp 1598350056
transform 1 0 5144 0 1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_491
timestamp 1598350056
transform -1 0 5096 0 1 610
box -16 -6 64 210
use FILL  FILL_4_2
timestamp 1598350056
transform 1 0 5192 0 1 610
box -16 -6 32 210
use FILL  FILL_4_1
timestamp 1598350056
transform 1 0 5176 0 1 610
box -16 -6 32 210
use NAND2X1  NAND2X1_838
timestamp 1598350056
transform 1 0 5000 0 1 610
box -16 -6 64 210
use INVX1  INVX1_309
timestamp 1598350056
transform 1 0 4968 0 1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_492
timestamp 1598350056
transform 1 0 4920 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_493
timestamp 1598350056
transform -1 0 4920 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_558
timestamp 1598350056
transform -1 0 4872 0 1 610
box -16 -6 64 210
use INVX1  INVX1_284
timestamp 1598350056
transform 1 0 4792 0 1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_494
timestamp 1598350056
transform 1 0 4744 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_383
timestamp 1598350056
transform 1 0 4696 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_556
timestamp 1598350056
transform 1 0 4600 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_631
timestamp 1598350056
transform -1 0 4600 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_384
timestamp 1598350056
transform -1 0 4696 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_561
timestamp 1598350056
transform 1 0 4456 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_557
timestamp 1598350056
transform 1 0 4360 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_625
timestamp 1598350056
transform -1 0 4552 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_522
timestamp 1598350056
transform -1 0 4456 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_523
timestamp 1598350056
transform 1 0 4312 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_849
timestamp 1598350056
transform -1 0 4264 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_490
timestamp 1598350056
transform -1 0 4312 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_827
timestamp 1598350056
transform 1 0 4168 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_670
timestamp 1598350056
transform 1 0 4120 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_88
timestamp 1598350056
transform -1 0 4120 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_232
timestamp 1598350056
transform 1 0 4024 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_66
timestamp 1598350056
transform 1 0 3976 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_845
timestamp 1598350056
transform 1 0 3928 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_100
timestamp 1598350056
transform 1 0 3880 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_86
timestamp 1598350056
transform -1 0 3880 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_240
timestamp 1598350056
transform -1 0 3784 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_412
timestamp 1598350056
transform -1 0 3832 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_85
timestamp 1598350056
transform -1 0 3736 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_243
timestamp 1598350056
transform 1 0 3640 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_54
timestamp 1598350056
transform 1 0 3544 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_565
timestamp 1598350056
transform 1 0 3496 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_235
timestamp 1598350056
transform -1 0 3640 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_569
timestamp 1598350056
transform 1 0 3400 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_391
timestamp 1598350056
transform 1 0 3352 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_530
timestamp 1598350056
transform 1 0 3448 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_137
timestamp 1598350056
transform 1 0 3304 0 1 610
box -16 -6 64 210
use INVX1  INVX1_59
timestamp 1598350056
transform -1 0 3256 0 1 610
box -18 -6 52 210
use INVX1  INVX1_61
timestamp 1598350056
transform -1 0 3224 0 1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_132
timestamp 1598350056
transform 1 0 3256 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_90
timestamp 1598350056
transform 1 0 3144 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_81
timestamp 1598350056
transform 1 0 2968 0 1 610
box -16 -6 64 210
use INVX1  INVX1_39
timestamp 1598350056
transform 1 0 3064 0 1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_102
timestamp 1598350056
transform 1 0 3096 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_293
timestamp 1598350056
transform -1 0 3064 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_344
timestamp 1598350056
transform -1 0 2968 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_208
timestamp 1598350056
transform -1 0 2872 0 1 610
box -16 -6 64 210
use INVX1  INVX1_89
timestamp 1598350056
transform -1 0 2824 0 1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_256
timestamp 1598350056
transform 1 0 2872 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_541
timestamp 1598350056
transform -1 0 2696 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_255
timestamp 1598350056
transform 1 0 2744 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_813
timestamp 1598350056
transform 1 0 2696 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_553
timestamp 1598350056
transform 1 0 2600 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_122
timestamp 1598350056
transform 1 0 2472 0 1 610
box -16 -6 64 210
use INVX1  INVX1_12
timestamp 1598350056
transform 1 0 2568 0 1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_101
timestamp 1598350056
transform -1 0 2568 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_666
timestamp 1598350056
transform 1 0 2328 0 1 610
box -16 -6 64 210
use INVX1  INVX1_123
timestamp 1598350056
transform 1 0 2296 0 1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_121
timestamp 1598350056
transform 1 0 2424 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_392
timestamp 1598350056
transform 1 0 2376 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_607
timestamp 1598350056
transform -1 0 2184 0 1 610
box -16 -6 64 210
use INVX1  INVX1_16
timestamp 1598350056
transform -1 0 2296 0 1 610
box -18 -6 52 210
use INVX1  INVX1_293
timestamp 1598350056
transform -1 0 2216 0 1 610
box -18 -6 52 210
use INVX1  INVX1_48
timestamp 1598350056
transform 1 0 2104 0 1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_99
timestamp 1598350056
transform -1 0 2264 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_77
timestamp 1598350056
transform -1 0 2104 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_120
timestamp 1598350056
transform -1 0 2056 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_62
timestamp 1598350056
transform -1 0 2008 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_748
timestamp 1598350056
transform -1 0 1960 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_73
timestamp 1598350056
transform 1 0 1816 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_789
timestamp 1598350056
transform 1 0 1864 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_63
timestamp 1598350056
transform -1 0 1816 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_133
timestamp 1598350056
transform -1 0 1736 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_159
timestamp 1598350056
transform -1 0 1688 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_10
timestamp 1598350056
transform -1 0 1640 0 1 610
box -16 -6 64 210
use INVX1  INVX1_7
timestamp 1598350056
transform -1 0 1768 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_670
timestamp 1598350056
transform 1 0 1448 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_126
timestamp 1598350056
transform 1 0 1544 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_673
timestamp 1598350056
transform -1 0 1544 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_67
timestamp 1598350056
transform 1 0 1400 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_263
timestamp 1598350056
transform 1 0 1272 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_813
timestamp 1598350056
transform 1 0 1224 0 1 610
box -16 -6 64 210
use INVX1  INVX1_26
timestamp 1598350056
transform -1 0 1352 0 1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_419
timestamp 1598350056
transform -1 0 1400 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_85
timestamp 1598350056
transform 1 0 1048 0 1 610
box -16 -6 64 210
use INVX1  INVX1_62
timestamp 1598350056
transform 1 0 1144 0 1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_239
timestamp 1598350056
transform -1 0 1224 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_845
timestamp 1598350056
transform 1 0 1096 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_235
timestamp 1598350056
transform -1 0 1048 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_202
timestamp 1598350056
transform -1 0 1000 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_100
timestamp 1598350056
transform -1 0 952 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_86
timestamp 1598350056
transform 1 0 856 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_506
timestamp 1598350056
transform 1 0 808 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_65
timestamp 1598350056
transform 1 0 760 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_862
timestamp 1598350056
transform 1 0 712 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_522
timestamp 1598350056
transform 1 0 568 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_849
timestamp 1598350056
transform -1 0 712 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_844
timestamp 1598350056
transform 1 0 616 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_60
timestamp 1598350056
transform -1 0 520 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_111
timestamp 1598350056
transform -1 0 424 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_865
timestamp 1598350056
transform 1 0 520 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_97
timestamp 1598350056
transform -1 0 472 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_89
timestamp 1598350056
transform 1 0 280 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_135
timestamp 1598350056
transform 1 0 232 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_45
timestamp 1598350056
transform -1 0 232 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_112
timestamp 1598350056
transform 1 0 328 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_234
timestamp 1598350056
transform 1 0 8 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_246
timestamp 1598350056
transform -1 0 184 0 1 610
box -16 -6 64 210
use INVX1  INVX1_120
timestamp 1598350056
transform -1 0 136 0 1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_242
timestamp 1598350056
transform 1 0 56 0 1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_735
timestamp 1598350056
transform -1 0 5128 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_576
timestamp 1598350056
transform 1 0 5128 0 -1 610
box -16 -6 64 210
use FILL  FILL_3_2
timestamp 1598350056
transform -1 0 5208 0 -1 610
box -16 -6 32 210
use FILL  FILL_3_1
timestamp 1598350056
transform -1 0 5192 0 -1 610
box -16 -6 32 210
use INVX1  INVX1_229
timestamp 1598350056
transform -1 0 5080 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_241
timestamp 1598350056
transform -1 0 5048 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_258
timestamp 1598350056
transform -1 0 4920 0 -1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_396
timestamp 1598350056
transform -1 0 5016 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_628
timestamp 1598350056
transform 1 0 4920 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_237
timestamp 1598350056
transform -1 0 4888 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_260
timestamp 1598350056
transform -1 0 4760 0 -1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_32
timestamp 1598350056
transform -1 0 4856 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_630
timestamp 1598350056
transform 1 0 4760 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_576
timestamp 1598350056
transform 1 0 4680 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_632
timestamp 1598350056
transform 1 0 4600 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_234
timestamp 1598350056
transform 1 0 4648 0 -1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_24
timestamp 1598350056
transform -1 0 4600 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_571
timestamp 1598350056
transform 1 0 4504 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_627
timestamp 1598350056
transform -1 0 4472 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_280
timestamp 1598350056
transform 1 0 4472 0 -1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_629
timestamp 1598350056
transform -1 0 4424 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_626
timestamp 1598350056
transform 1 0 4328 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_172
timestamp 1598350056
transform -1 0 4328 0 -1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_521
timestamp 1598350056
transform 1 0 4248 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_413
timestamp 1598350056
transform 1 0 4200 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_87
timestamp 1598350056
transform -1 0 4168 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_837
timestamp 1598350056
transform 1 0 4024 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_217
timestamp 1598350056
transform 1 0 4168 0 -1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_826
timestamp 1598350056
transform 1 0 4072 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_859
timestamp 1598350056
transform 1 0 3976 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_673
timestamp 1598350056
transform -1 0 3976 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_848
timestamp 1598350056
transform 1 0 3880 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_672
timestamp 1598350056
transform 1 0 3832 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_98
timestamp 1598350056
transform -1 0 3736 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_96
timestamp 1598350056
transform -1 0 3832 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_825
timestamp 1598350056
transform -1 0 3784 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_531
timestamp 1598350056
transform -1 0 3592 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_219
timestamp 1598350056
transform -1 0 3544 0 -1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_93
timestamp 1598350056
transform -1 0 3688 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_94
timestamp 1598350056
transform 1 0 3592 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_549
timestamp 1598350056
transform -1 0 3512 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_548
timestamp 1598350056
transform 1 0 3416 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_529
timestamp 1598350056
transform -1 0 3416 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_23
timestamp 1598350056
transform -1 0 3368 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_671
timestamp 1598350056
transform -1 0 3320 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_29
timestamp 1598350056
transform -1 0 3272 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_143
timestamp 1598350056
transform 1 0 3176 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_104
timestamp 1598350056
transform 1 0 3128 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_37
timestamp 1598350056
transform 1 0 3080 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_8
timestamp 1598350056
transform -1 0 3080 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_84
timestamp 1598350056
transform -1 0 3032 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_49
timestamp 1598350056
transform 1 0 2888 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_232
timestamp 1598350056
transform 1 0 2808 0 -1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_42
timestamp 1598350056
transform 1 0 2936 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_572
timestamp 1598350056
transform -1 0 2888 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_131
timestamp 1598350056
transform 1 0 2712 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_129
timestamp 1598350056
transform -1 0 2712 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_130
timestamp 1598350056
transform 1 0 2760 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_124
timestamp 1598350056
transform -1 0 2664 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_205
timestamp 1598350056
transform -1 0 2616 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_112
timestamp 1598350056
transform 1 0 2536 0 -1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_204
timestamp 1598350056
transform -1 0 2536 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_719
timestamp 1598350056
transform -1 0 2488 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_79
timestamp 1598350056
transform 1 0 2392 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_665
timestamp 1598350056
transform 1 0 2296 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_391
timestamp 1598350056
transform 1 0 2344 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_767
timestamp 1598350056
transform -1 0 2248 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_755
timestamp 1598350056
transform 1 0 2152 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_78
timestamp 1598350056
transform 1 0 2248 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_646
timestamp 1598350056
transform 1 0 2104 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_42
timestamp 1598350056
transform 1 0 2056 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_609
timestamp 1598350056
transform 1 0 1960 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_664
timestamp 1598350056
transform 1 0 2008 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_749
timestamp 1598350056
transform 1 0 1864 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_751
timestamp 1598350056
transform 1 0 1816 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_608
timestamp 1598350056
transform 1 0 1912 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_750
timestamp 1598350056
transform -1 0 1816 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_415
timestamp 1598350056
transform -1 0 1768 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_215
timestamp 1598350056
transform 1 0 1640 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_2
timestamp 1598350056
transform -1 0 1720 0 -1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_414
timestamp 1598350056
transform 1 0 1592 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_296
timestamp 1598350056
transform 1 0 1544 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_138
timestamp 1598350056
transform -1 0 1496 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_230
timestamp 1598350056
transform 1 0 1432 0 -1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_297
timestamp 1598350056
transform -1 0 1544 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_861
timestamp 1598350056
transform 1 0 1384 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_860
timestamp 1598350056
transform -1 0 1384 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_360
timestamp 1598350056
transform 1 0 1288 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_347
timestamp 1598350056
transform 1 0 1240 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_295
timestamp 1598350056
transform 1 0 1144 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_38
timestamp 1598350056
transform -1 0 1144 0 -1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_346
timestamp 1598350056
transform 1 0 1192 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_416
timestamp 1598350056
transform 1 0 1064 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_88
timestamp 1598350056
transform -1 0 1016 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_206
timestamp 1598350056
transform 1 0 872 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_87
timestamp 1598350056
transform 1 0 1016 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_560
timestamp 1598350056
transform 1 0 920 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_110
timestamp 1598350056
transform 1 0 744 0 -1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_340
timestamp 1598350056
transform 1 0 824 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_201
timestamp 1598350056
transform -1 0 824 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_521
timestamp 1598350056
transform -1 0 696 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_58
timestamp 1598350056
transform 1 0 552 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_859
timestamp 1598350056
transform 1 0 696 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_523
timestamp 1598350056
transform 1 0 600 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_152
timestamp 1598350056
transform -1 0 552 0 -1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_61
timestamp 1598350056
transform 1 0 472 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_339
timestamp 1598350056
transform 1 0 424 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_332
timestamp 1598350056
transform -1 0 424 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_233
timestamp 1598350056
transform -1 0 376 0 -1 610
box -16 -6 64 210
use INVX1  INVX1_64
timestamp 1598350056
transform -1 0 232 0 -1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_715
timestamp 1598350056
transform 1 0 280 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_702
timestamp 1598350056
transform -1 0 280 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_232
timestamp 1598350056
transform -1 0 104 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_243
timestamp 1598350056
transform 1 0 152 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_244
timestamp 1598350056
transform -1 0 152 0 -1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_240
timestamp 1598350056
transform 1 0 8 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_736
timestamp 1598350056
transform 1 0 5144 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_725
timestamp 1598350056
transform -1 0 5144 0 1 210
box -16 -6 64 210
use INVX1  INVX1_240
timestamp 1598350056
transform 1 0 5064 0 1 210
box -18 -6 52 210
use FILL  FILL_2_1
timestamp 1598350056
transform 1 0 5192 0 1 210
box -16 -6 32 210
use NAND2X1  NAND2X1_401
timestamp 1598350056
transform -1 0 5064 0 1 210
box -16 -6 64 210
use INVX1  INVX1_5
timestamp 1598350056
transform 1 0 4936 0 1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_395
timestamp 1598350056
transform 1 0 4968 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_27
timestamp 1598350056
transform 1 0 4888 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_34
timestamp 1598350056
transform -1 0 4888 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_35
timestamp 1598350056
transform -1 0 4760 0 1 210
box -16 -6 64 210
use INVX1  INVX1_207
timestamp 1598350056
transform -1 0 4840 0 1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_411
timestamp 1598350056
transform 1 0 4760 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_461
timestamp 1598350056
transform -1 0 4712 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_410
timestamp 1598350056
transform 1 0 4616 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_33
timestamp 1598350056
transform 1 0 4568 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_621
timestamp 1598350056
transform 1 0 4376 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_399
timestamp 1598350056
transform 1 0 4520 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_20
timestamp 1598350056
transform 1 0 4472 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_616
timestamp 1598350056
transform -1 0 4472 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_624
timestamp 1598350056
transform 1 0 4248 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_658
timestamp 1598350056
transform 1 0 4200 0 1 210
box -16 -6 64 210
use INVX1  INVX1_15
timestamp 1598350056
transform 1 0 4296 0 1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_19
timestamp 1598350056
transform -1 0 4376 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_619
timestamp 1598350056
transform -1 0 4168 0 1 210
box -16 -6 64 210
use INVX1  INVX1_255
timestamp 1598350056
transform -1 0 4200 0 1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_474
timestamp 1598350056
transform -1 0 4120 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_475
timestamp 1598350056
transform 1 0 4024 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_570
timestamp 1598350056
transform 1 0 3928 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_577
timestamp 1598350056
transform 1 0 3880 0 1 210
box -16 -6 64 210
use INVX1  INVX1_178
timestamp 1598350056
transform -1 0 3880 0 1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_642
timestamp 1598350056
transform 1 0 3976 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_562
timestamp 1598350056
transform 1 0 3800 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_578
timestamp 1598350056
transform 1 0 3752 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_397
timestamp 1598350056
transform 1 0 3656 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_662
timestamp 1598350056
transform -1 0 3752 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_618
timestamp 1598350056
transform 1 0 3608 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_515
timestamp 1598350056
transform 1 0 3560 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_514
timestamp 1598350056
transform 1 0 3512 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_136
timestamp 1598350056
transform -1 0 3512 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_139
timestamp 1598350056
transform -1 0 3464 0 1 210
box -16 -6 64 210
use INVX1  INVX1_80
timestamp 1598350056
transform 1 0 3384 0 1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_4
timestamp 1598350056
transform 1 0 3336 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_83
timestamp 1598350056
transform -1 0 3208 0 1 210
box -16 -6 64 210
use INVX1  INVX1_216
timestamp 1598350056
transform -1 0 3336 0 1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_516
timestamp 1598350056
transform -1 0 3304 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_138
timestamp 1598350056
transform -1 0 3256 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_82
timestamp 1598350056
transform 1 0 3016 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_563
timestamp 1598350056
transform 1 0 2968 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_382
timestamp 1598350056
transform -1 0 3160 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_28
timestamp 1598350056
transform 1 0 3064 0 1 210
box -16 -6 64 210
use INVX1  INVX1_316
timestamp 1598350056
transform 1 0 2936 0 1 210
box -18 -6 52 210
use INVX1  INVX1_228
timestamp 1598350056
transform 1 0 2904 0 1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_381
timestamp 1598350056
transform 1 0 2856 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_817
timestamp 1598350056
transform -1 0 2856 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_125
timestamp 1598350056
transform -1 0 2712 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_381
timestamp 1598350056
transform -1 0 2664 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_847
timestamp 1598350056
transform 1 0 2760 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_554
timestamp 1598350056
transform -1 0 2760 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_817
timestamp 1598350056
transform 1 0 2568 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_382
timestamp 1598350056
transform 1 0 2520 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_656
timestamp 1598350056
transform 1 0 2472 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_819
timestamp 1598350056
transform -1 0 2376 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_820
timestamp 1598350056
transform 1 0 2280 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_660
timestamp 1598350056
transform -1 0 2472 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_647
timestamp 1598350056
transform -1 0 2424 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_818
timestamp 1598350056
transform 1 0 2104 0 1 210
box -16 -6 64 210
use INVX1  INVX1_40
timestamp 1598350056
transform -1 0 2280 0 1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_819
timestamp 1598350056
transform -1 0 2248 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_820
timestamp 1598350056
transform -1 0 2200 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_847
timestamp 1598350056
transform -1 0 2104 0 1 210
box -16 -6 64 210
use INVX1  INVX1_4
timestamp 1598350056
transform 1 0 2024 0 1 210
box -18 -6 52 210
use INVX1  INVX1_315
timestamp 1598350056
transform -1 0 1976 0 1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_818
timestamp 1598350056
transform 1 0 1976 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_104
timestamp 1598350056
transform 1 0 1896 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_143
timestamp 1598350056
transform 1 0 1848 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_473
timestamp 1598350056
transform 1 0 1752 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_655
timestamp 1598350056
transform 1 0 1800 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_216
timestamp 1598350056
transform 1 0 1608 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_649
timestamp 1598350056
transform 1 0 1704 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_54
timestamp 1598350056
transform 1 0 1656 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_219
timestamp 1598350056
transform 1 0 1560 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_214
timestamp 1598350056
transform 1 0 1512 0 1 210
box -16 -6 64 210
use INVX1  INVX1_20
timestamp 1598350056
transform 1 0 1480 0 1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_643
timestamp 1598350056
transform -1 0 1480 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_29
timestamp 1598350056
transform -1 0 1432 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_27
timestamp 1598350056
transform -1 0 1336 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_207
timestamp 1598350056
transform 1 0 1240 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_294
timestamp 1598350056
transform -1 0 1384 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_481
timestamp 1598350056
transform -1 0 1240 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_816
timestamp 1598350056
transform 1 0 1096 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_848
timestamp 1598350056
transform -1 0 1192 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_846
timestamp 1598350056
transform -1 0 1096 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_815
timestamp 1598350056
transform 1 0 1000 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_251
timestamp 1598350056
transform -1 0 952 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_814
timestamp 1598350056
transform 1 0 952 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_106
timestamp 1598350056
transform 1 0 776 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_43
timestamp 1598350056
transform -1 0 776 0 1 210
box -16 -6 64 210
use INVX1  INVX1_36
timestamp 1598350056
transform -1 0 856 0 1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_105
timestamp 1598350056
transform -1 0 904 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_116
timestamp 1598350056
transform -1 0 648 0 1 210
box -16 -6 64 210
use INVX1  INVX1_108
timestamp 1598350056
transform 1 0 648 0 1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_195
timestamp 1598350056
transform -1 0 728 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_199
timestamp 1598350056
transform 1 0 552 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_48
timestamp 1598350056
transform 1 0 424 0 1 210
box -16 -6 64 210
use INVX1  INVX1_68
timestamp 1598350056
transform 1 0 520 0 1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_115
timestamp 1598350056
transform 1 0 472 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_196
timestamp 1598350056
transform -1 0 424 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_248
timestamp 1598350056
transform -1 0 328 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_257
timestamp 1598350056
transform 1 0 232 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_247
timestamp 1598350056
transform 1 0 328 0 1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_260
timestamp 1598350056
transform 1 0 184 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_348
timestamp 1598350056
transform -1 0 56 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_261
timestamp 1598350056
transform -1 0 184 0 1 210
box -16 -6 64 210
use INVX1  INVX1_154
timestamp 1598350056
transform -1 0 88 0 1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_342
timestamp 1598350056
transform -1 0 136 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_580
timestamp 1598350056
transform -1 0 5144 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_242
timestamp 1598350056
transform 1 0 5064 0 -1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_298
timestamp 1598350056
transform -1 0 5192 0 -1 210
box -16 -6 64 210
use FILL  FILL_1_1
timestamp 1598350056
transform -1 0 5208 0 -1 210
box -16 -6 32 210
use NAND2X1  NAND2X1_402
timestamp 1598350056
transform -1 0 4984 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_239
timestamp 1598350056
transform 1 0 4984 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_167
timestamp 1598350056
transform -1 0 4936 0 -1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_580
timestamp 1598350056
transform -1 0 5064 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_163
timestamp 1598350056
transform 1 0 4824 0 -1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_299
timestamp 1598350056
transform 1 0 4856 0 -1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_579
timestamp 1598350056
transform 1 0 4776 0 -1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_573
timestamp 1598350056
transform -1 0 4776 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_403
timestamp 1598350056
transform 1 0 4552 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_169
timestamp 1598350056
transform 1 0 4600 0 -1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_575
timestamp 1598350056
transform 1 0 4680 0 -1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_404
timestamp 1598350056
transform 1 0 4632 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_398
timestamp 1598350056
transform 1 0 4472 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_463
timestamp 1598350056
transform 1 0 4360 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_166
timestamp 1598350056
transform 1 0 4520 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_135
timestamp 1598350056
transform 1 0 4440 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_197
timestamp 1598350056
transform -1 0 4440 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_622
timestamp 1598350056
transform -1 0 4328 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_194
timestamp 1598350056
transform 1 0 4328 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_195
timestamp 1598350056
transform 1 0 4200 0 -1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_472
timestamp 1598350056
transform -1 0 4280 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_462
timestamp 1598350056
transform 1 0 4152 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_253
timestamp 1598350056
transform 1 0 4120 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_175
timestamp 1598350056
transform 1 0 4040 0 -1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_459
timestamp 1598350056
transform -1 0 4120 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_376
timestamp 1598350056
transform 1 0 3992 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_84
timestamp 1598350056
transform 1 0 3960 0 -1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_479
timestamp 1598350056
transform 1 0 3912 0 -1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_476
timestamp 1598350056
transform 1 0 3864 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_203
timestamp 1598350056
transform -1 0 3864 0 -1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_480
timestamp 1598350056
transform 1 0 3784 0 -1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_375
timestamp 1598350056
transform 1 0 3736 0 -1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_663
timestamp 1598350056
transform -1 0 3736 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_659
timestamp 1598350056
transform 1 0 3608 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_378
timestamp 1598350056
transform 1 0 3560 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_377
timestamp 1598350056
transform 1 0 3512 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_267
timestamp 1598350056
transform 1 0 3656 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_416
timestamp 1598350056
transform 1 0 3464 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_394
timestamp 1598350056
transform -1 0 3432 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_90
timestamp 1598350056
transform 1 0 3432 0 -1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_400
timestamp 1598350056
transform -1 0 3384 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_393
timestamp 1598350056
transform 1 0 3288 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_574
timestamp 1598350056
transform 1 0 3208 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_657
timestamp 1598350056
transform 1 0 3160 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_235
timestamp 1598350056
transform 1 0 3256 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_414
timestamp 1598350056
transform 1 0 3064 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_28
timestamp 1598350056
transform 1 0 3016 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_14
timestamp 1598350056
transform -1 0 3016 0 -1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_415
timestamp 1598350056
transform 1 0 3112 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_141
timestamp 1598350056
transform -1 0 2968 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_5
timestamp 1598350056
transform -1 0 2920 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_293
timestamp 1598350056
transform -1 0 2840 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_82
timestamp 1598350056
transform 1 0 2840 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_127
timestamp 1598350056
transform 1 0 2648 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_74
timestamp 1598350056
transform -1 0 2648 0 -1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_140
timestamp 1598350056
transform -1 0 2792 0 -1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_128
timestamp 1598350056
transform 1 0 2696 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_217
timestamp 1598350056
transform -1 0 2616 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_4
timestamp 1598350056
transform -1 0 2568 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_38
timestamp 1598350056
transform -1 0 2520 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_23
timestamp 1598350056
transform -1 0 2472 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_612
timestamp 1598350056
transform -1 0 2376 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_252
timestamp 1598350056
transform 1 0 2296 0 -1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_610
timestamp 1598350056
transform 1 0 2376 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_126
timestamp 1598350056
transform 1 0 2168 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_6
timestamp 1598350056
transform -1 0 2168 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_3
timestamp 1598350056
transform 1 0 2216 0 -1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_611
timestamp 1598350056
transform 1 0 2248 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_225
timestamp 1598350056
transform -1 0 2088 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_201
timestamp 1598350056
transform 1 0 2088 0 -1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_14
timestamp 1598350056
transform -1 0 2040 0 -1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_5
timestamp 1598350056
transform -1 0 1992 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_8
timestamp 1598350056
transform 1 0 1896 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_37
timestamp 1598350056
transform 1 0 1848 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_671
timestamp 1598350056
transform -1 0 1848 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_672
timestamp 1598350056
transform 1 0 1752 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_46
timestamp 1598350056
transform 1 0 1704 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_218
timestamp 1598350056
transform -1 0 1704 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_222
timestamp 1598350056
transform -1 0 1656 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_19
timestamp 1598350056
transform -1 0 1608 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_223
timestamp 1598350056
transform -1 0 1560 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_595
timestamp 1598350056
transform -1 0 1512 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_20
timestamp 1598350056
transform -1 0 1464 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_24
timestamp 1598350056
transform 1 0 1224 0 -1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_33
timestamp 1598350056
transform 1 0 1368 0 -1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_35
timestamp 1598350056
transform 1 0 1320 0 -1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_34
timestamp 1598350056
transform 1 0 1272 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_32
timestamp 1598350056
transform -1 0 1224 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_555
timestamp 1598350056
transform 1 0 1096 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_205
timestamp 1598350056
transform -1 0 1176 0 -1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_249
timestamp 1598350056
transform 1 0 1048 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_250
timestamp 1598350056
transform 1 0 1000 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_510
timestamp 1598350056
transform 1 0 904 0 -1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_343
timestamp 1598350056
transform 1 0 952 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_503
timestamp 1598350056
transform 1 0 776 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_212
timestamp 1598350056
transform 1 0 872 0 -1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_509
timestamp 1598350056
transform 1 0 824 0 -1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_502
timestamp 1598350056
transform 1 0 728 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_508
timestamp 1598350056
transform -1 0 728 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_41
timestamp 1598350056
transform 1 0 632 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_226
timestamp 1598350056
transform 1 0 584 0 -1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_227
timestamp 1598350056
transform -1 0 584 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_224
timestamp 1598350056
transform 1 0 488 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_504
timestamp 1598350056
transform -1 0 424 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_210
timestamp 1598350056
transform 1 0 456 0 -1 210
box -18 -6 52 210
use INVX1  INVX1_122
timestamp 1598350056
transform 1 0 424 0 -1 210
box -18 -6 52 210
use NAND2X1  NAND2X1_505
timestamp 1598350056
transform -1 0 328 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_258
timestamp 1598350056
transform 1 0 184 0 -1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_507
timestamp 1598350056
transform 1 0 328 0 -1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_259
timestamp 1598350056
transform 1 0 232 0 -1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_359
timestamp 1598350056
transform 1 0 8 0 -1 210
box -16 -6 64 210
use INVX1  INVX1_156
timestamp 1598350056
transform -1 0 88 0 -1 210
box -18 -6 52 210
use NOR2X1  NOR2X1_345
timestamp 1598350056
transform 1 0 136 0 -1 210
box -16 -6 64 210
use NOR2X1  NOR2X1_349
timestamp 1598350056
transform -1 0 136 0 -1 210
box -16 -6 64 210
<< labels >>
rlabel metal2 s 2608 -40 2608 -40 8 INPUT_0
port 0 nsew
rlabel metal2 s 3136 -40 3136 -40 8 D_INPUT_0
port 1 nsew
rlabel metal2 s 3056 -40 3056 -40 8 INPUT_1
port 2 nsew
rlabel metal2 s 2528 -40 2528 -40 8 D_INPUT_1
port 3 nsew
rlabel metal2 s 2032 -40 2032 -40 8 INPUT_2
port 4 nsew
rlabel metal2 s 3008 -40 3008 -40 8 D_INPUT_2
port 5 nsew
rlabel metal2 s 1888 -40 1888 -40 8 INPUT_3
port 6 nsew
rlabel metal2 s 2976 -40 2976 -40 8 D_INPUT_3
port 7 nsew
rlabel metal2 s 4992 3680 4992 3680 6 INPUT_4
port 8 nsew
rlabel metal2 s 4800 3680 4800 3680 6 D_INPUT_4
port 9 nsew
rlabel metal2 s 4960 3680 4960 3680 6 INPUT_5
port 10 nsew
rlabel metal2 s 5056 3680 5056 3680 6 D_INPUT_5
port 11 nsew
rlabel metal2 s 4512 3680 4512 3680 6 INPUT_6
port 12 nsew
rlabel metal2 s 4880 3680 4880 3680 6 D_INPUT_6
port 13 nsew
rlabel metal2 s 4176 3680 4176 3680 6 INPUT_7
port 14 nsew
rlabel metal2 s 4336 3680 4336 3680 6 D_INPUT_7
port 15 nsew
rlabel metal2 s 2192 3680 2192 3680 6 D_GATE_222
port 16 nsew
rlabel metal2 s 3264 3680 3264 3680 6 D_GATE_366
port 17 nsew
rlabel metal2 s 3808 -40 3808 -40 8 D_GATE_479
port 18 nsew
rlabel metal2 s 5008 -40 5008 -40 8 D_GATE_579
port 19 nsew
rlabel metal2 s 3728 -40 3728 -40 8 D_GATE_662
port 20 nsew
rlabel metal2 s 816 3680 816 3680 6 D_GATE_741
port 21 nsew
rlabel metal3 s -48 2140 -48 2140 4 D_GATE_811
port 22 nsew
rlabel metal3 s -48 1480 -48 1480 4 D_GATE_865
port 23 nsew
rlabel metal2 s 1552 -40 1552 -40 8 GATE_222
port 24 nsew
rlabel metal3 s -48 1380 -48 1380 4 GATE_366
port 25 nsew
rlabel metal2 s 2304 3680 2304 3680 6 GATE_479
port 26 nsew
rlabel metal2 s 5088 -40 5088 -40 8 GATE_579
port 27 nsew
rlabel metal2 s 3392 3680 3392 3680 6 GATE_662
port 28 nsew
rlabel metal3 s -48 560 -48 560 4 gate
port 32 nsew
rlabel metal3 s -48 580 -48 580 4 type:
port 33 nsew
rlabel metal3 s -48 1680 -48 1680 4 NAND;
port 34 nsew
rlabel metal3 s -48 2180 -48 2180 4 name:
port 35 nsew
rlabel metal3 s -48 60 -48 60 4 GATE_0_I0
port 36 nsew
rlabel metal3 s 5264 980 5264 980 6 GATE_865
port 31 nsew
rlabel metal3 s 5264 2180 5264 2180 6 GATE_811
port 30 nsew
rlabel metal3 s 5264 1920 5264 1920 6 GATE_741
port 29 nsew
rlabel space -408 -43 5626 3740 1 vdd
rlabel space -408 -43 5626 3740 1 gnd
<< end >>
