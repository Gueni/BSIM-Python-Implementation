magic
tech scmos
magscale 1 2
timestamp 1602346068
<< checkpaint >>
rect 40000 8000 45032 11464
rect 40800 800 45032 8000
rect 29244 145 45032 800
rect 29600 0 45032 145
rect 29204 -59 45032 0
rect 29600 -102 45032 -59
<< error_s >>
rect 32096 11277 32104 11285
rect 32160 11277 32168 11285
rect 34416 11277 34424 11285
rect 34368 11237 34376 11245
rect 38096 11237 38104 11245
rect 34688 11217 34696 11225
rect 35408 11217 35416 11225
rect 35696 11217 35704 11225
rect 39408 11217 39416 11225
rect 31200 11197 31208 11205
rect 36224 11197 36232 11205
rect 29936 11177 29944 11185
rect 29984 11177 29992 11185
rect 30432 11177 30440 11185
rect 30480 11177 30488 11185
rect 30912 11177 30920 11185
rect 31408 11177 31416 11185
rect 31632 11177 31640 11185
rect 31840 11177 31848 11185
rect 32752 11177 32760 11185
rect 33008 11177 33016 11185
rect 33744 11177 33752 11185
rect 34016 11177 34024 11185
rect 35104 11177 35112 11185
rect 36912 11177 36920 11185
rect 37024 11177 37032 11185
rect 38384 11177 38392 11185
rect 38464 11177 38472 11185
rect 38624 11177 38632 11185
rect 39088 11177 39096 11185
rect 39264 11177 39272 11185
rect 39360 11177 39368 11185
rect 39520 11177 39528 11185
rect 30320 11157 30328 11165
rect 31568 11157 31576 11165
rect 33952 11157 33960 11165
rect 34768 11157 34776 11165
rect 36064 11157 36072 11165
rect 36240 11157 36248 11165
rect 36636 11164 36638 11165
rect 36636 11157 36638 11158
rect 37984 11157 37992 11165
rect 38096 11157 38104 11165
rect 39456 11157 39464 11165
rect 29408 11137 29416 11145
rect 29488 11137 29496 11145
rect 30512 11137 30520 11145
rect 31040 11137 31048 11145
rect 31200 11137 31208 11145
rect 32000 11137 32008 11145
rect 32640 11137 32648 11145
rect 32864 11137 32872 11145
rect 33840 11137 33848 11145
rect 34384 11137 34392 11145
rect 34560 11137 34568 11145
rect 34784 11137 34792 11145
rect 35408 11137 35416 11145
rect 35584 11137 35592 11145
rect 35760 11137 35768 11145
rect 29504 11117 29512 11125
rect 29616 11117 29624 11125
rect 30176 11117 30184 11125
rect 30256 11117 30264 11125
rect 30512 11117 30520 11125
rect 30720 11117 30728 11125
rect 31008 11117 31016 11125
rect 31056 11117 31064 11125
rect 31920 11117 31928 11125
rect 32080 11117 32088 11125
rect 32304 11117 32312 11125
rect 32384 11117 32392 11125
rect 33248 11117 33256 11125
rect 33584 11117 33592 11125
rect 33648 11117 33656 11125
rect 33824 11117 33832 11125
rect 33888 11117 33896 11125
rect 33984 11117 33992 11125
rect 34144 11117 34152 11125
rect 34608 11117 34616 11125
rect 35232 11117 35240 11125
rect 35296 11117 35304 11125
rect 36064 11117 36072 11125
rect 37552 11117 37560 11125
rect 38320 11117 38328 11125
rect 38560 11117 38568 11125
rect 38704 11117 38712 11125
rect 32072 11105 32073 11110
rect 34112 11097 34120 11105
rect 35248 11097 35256 11105
rect 36672 11097 36680 11105
rect 36992 11097 37000 11105
rect 38880 11097 38888 11105
rect 38896 11097 38904 11105
rect 38976 11097 38984 11105
rect 39728 11097 39736 11105
rect 31440 11077 31448 11085
rect 38016 11077 38024 11085
rect 38336 11077 38344 11085
rect 39536 11077 39544 11085
rect 29380 11067 29392 11075
rect 29412 11067 29424 11075
rect 29428 11067 29432 11075
rect 29448 11067 29464 11075
rect 29480 11067 29512 11075
rect 29528 11067 29552 11075
rect 29568 11067 29572 11075
rect 29576 11067 29588 11075
rect 29604 11067 29628 11075
rect 29644 11067 29660 11075
rect 29676 11067 29688 11075
rect 29700 11067 29704 11075
rect 29708 11067 29712 11075
rect 29724 11067 29736 11075
rect 29748 11067 29752 11075
rect 29756 11067 29760 11075
rect 29772 11067 29784 11075
rect 29896 11067 29908 11075
rect 29920 11067 29924 11075
rect 29928 11067 29932 11075
rect 29944 11067 29956 11075
rect 30108 11067 30112 11075
rect 30116 11067 30120 11075
rect 30140 11067 30144 11075
rect 30148 11067 30152 11075
rect 30164 11067 30176 11075
rect 30184 11067 30200 11075
rect 30216 11067 30220 11075
rect 30224 11067 30228 11075
rect 30240 11067 30252 11075
rect 30260 11067 30276 11075
rect 30292 11067 30296 11075
rect 30300 11067 30304 11075
rect 30316 11067 30328 11075
rect 30336 11067 30352 11075
rect 30368 11067 30372 11075
rect 30376 11067 30380 11075
rect 30392 11067 30400 11075
rect 30412 11067 30428 11075
rect 30444 11067 30460 11075
rect 30468 11067 30480 11075
rect 30492 11067 30496 11075
rect 30500 11067 30504 11075
rect 30516 11067 30528 11075
rect 30540 11067 30544 11075
rect 30548 11067 30552 11075
rect 30568 11067 30600 11075
rect 30616 11067 30632 11075
rect 30648 11067 30664 11075
rect 30680 11067 30696 11075
rect 30712 11067 30744 11075
rect 30760 11067 30772 11075
rect 30792 11067 30804 11075
rect 30816 11067 30820 11075
rect 30824 11067 30828 11075
rect 30916 11067 30928 11075
rect 30984 11067 30988 11075
rect 30992 11067 30996 11075
rect 31016 11067 31020 11075
rect 31024 11067 31028 11075
rect 31040 11067 31052 11075
rect 31068 11067 31084 11075
rect 31100 11067 31132 11075
rect 31140 11067 31156 11075
rect 31172 11067 31184 11075
rect 31188 11067 31200 11075
rect 31204 11067 31216 11075
rect 31264 11067 31276 11075
rect 31280 11067 31292 11075
rect 31296 11067 31308 11075
rect 31356 11067 31368 11075
rect 31372 11067 31384 11075
rect 31388 11067 31400 11075
rect 31420 11067 31432 11075
rect 31448 11067 31472 11075
rect 31480 11067 31496 11075
rect 31512 11067 31560 11075
rect 31576 11067 31588 11075
rect 31604 11067 31652 11075
rect 31668 11067 31684 11075
rect 31696 11067 31744 11075
rect 31760 11067 31776 11075
rect 31792 11067 31796 11075
rect 31800 11067 31812 11075
rect 31824 11067 31828 11075
rect 31832 11067 31836 11075
rect 31856 11067 31860 11075
rect 31864 11067 31868 11075
rect 31932 11067 31936 11075
rect 31940 11067 31944 11075
rect 31964 11067 31968 11075
rect 31972 11067 31976 11075
rect 31988 11067 32000 11075
rect 32004 11067 32008 11075
rect 32028 11067 32032 11075
rect 32036 11067 32048 11075
rect 32060 11067 32064 11075
rect 32068 11067 32072 11075
rect 32092 11067 32096 11075
rect 32100 11067 32112 11075
rect 32124 11067 32128 11075
rect 32132 11067 32136 11075
rect 32184 11067 32188 11075
rect 32192 11067 32204 11075
rect 32216 11067 32220 11075
rect 32224 11067 32228 11075
rect 32240 11067 32252 11075
rect 32256 11067 32268 11075
rect 32280 11067 32284 11075
rect 32288 11067 32292 11075
rect 32312 11067 32316 11075
rect 32320 11067 32332 11075
rect 32344 11067 32348 11075
rect 32352 11067 32356 11075
rect 32376 11067 32380 11075
rect 32384 11067 32388 11075
rect 32452 11067 32456 11075
rect 32460 11067 32472 11075
rect 32484 11067 32488 11075
rect 32492 11067 32496 11075
rect 32508 11067 32520 11075
rect 32524 11067 32528 11075
rect 32548 11067 32552 11075
rect 32556 11067 32560 11075
rect 32576 11067 32592 11075
rect 32600 11067 32632 11075
rect 32640 11067 32652 11075
rect 32668 11067 32684 11075
rect 32692 11067 32724 11075
rect 32732 11067 32748 11075
rect 32764 11067 32776 11075
rect 32784 11067 32816 11075
rect 32824 11067 32840 11075
rect 32856 11067 32868 11075
rect 32880 11067 32884 11075
rect 32888 11067 32900 11075
rect 33036 11067 33040 11075
rect 33044 11067 33056 11075
rect 33060 11067 33064 11075
rect 33076 11067 33088 11075
rect 33328 11067 33340 11075
rect 33352 11067 33356 11075
rect 33360 11067 33372 11075
rect 33376 11067 33380 11075
rect 33392 11067 33404 11075
rect 33424 11067 33436 11075
rect 33440 11067 33444 11075
rect 33456 11067 33468 11075
rect 33488 11067 33500 11075
rect 33504 11067 33516 11075
rect 33520 11067 33532 11075
rect 33552 11067 33564 11075
rect 33580 11067 33600 11075
rect 33612 11067 33628 11075
rect 33644 11067 33648 11075
rect 33652 11067 33656 11075
rect 33668 11067 33680 11075
rect 33684 11067 33696 11075
rect 33708 11067 33712 11075
rect 33716 11067 33720 11075
rect 33848 11067 33852 11075
rect 33856 11067 33860 11075
rect 33872 11067 33884 11075
rect 33888 11067 33900 11075
rect 33912 11067 33916 11075
rect 33920 11067 33924 11075
rect 33940 11067 33988 11075
rect 34000 11067 34016 11075
rect 34032 11067 34080 11075
rect 34096 11067 34108 11075
rect 34128 11067 34140 11075
rect 34152 11067 34156 11075
rect 34160 11067 34172 11075
rect 34244 11067 34248 11075
rect 34252 11067 34264 11075
rect 34460 11067 34464 11075
rect 34468 11067 34480 11075
rect 34500 11067 34512 11075
rect 34516 11067 34520 11075
rect 34532 11067 34544 11075
rect 34564 11067 34576 11075
rect 34592 11067 34640 11075
rect 34656 11067 34672 11075
rect 34680 11067 34692 11075
rect 34696 11067 34708 11075
rect 34720 11067 34724 11075
rect 34728 11067 34732 11075
rect 34748 11067 34752 11075
rect 34756 11067 34760 11075
rect 34772 11067 34784 11075
rect 34788 11067 34800 11075
rect 34812 11067 34816 11075
rect 34820 11067 34824 11075
rect 34840 11067 34856 11075
rect 34864 11067 34876 11075
rect 34880 11067 34892 11075
rect 34904 11067 34908 11075
rect 34912 11067 34916 11075
rect 34936 11067 34940 11075
rect 34944 11067 34948 11075
rect 35044 11067 35048 11075
rect 35052 11067 35056 11075
rect 35068 11067 35080 11075
rect 35084 11067 35096 11075
rect 35108 11067 35112 11075
rect 35116 11067 35120 11075
rect 35136 11067 35152 11075
rect 35160 11067 35172 11075
rect 35176 11067 35188 11075
rect 35200 11067 35204 11075
rect 35208 11067 35212 11075
rect 35228 11067 35244 11075
rect 35252 11067 35276 11075
rect 35292 11067 35308 11075
rect 35324 11067 35348 11075
rect 35356 11067 35372 11075
rect 35388 11067 35436 11075
rect 35448 11067 35464 11075
rect 35480 11067 35528 11075
rect 35544 11067 35560 11075
rect 35572 11067 35620 11075
rect 35636 11067 35652 11075
rect 35664 11067 35712 11075
rect 35728 11067 35752 11075
rect 35760 11067 35776 11075
rect 35792 11067 35808 11075
rect 35824 11067 35828 11075
rect 35832 11067 35844 11075
rect 35848 11067 35860 11075
rect 35864 11067 35868 11075
rect 35888 11067 35892 11075
rect 35896 11067 35900 11075
rect 35964 11067 35968 11075
rect 35972 11067 35976 11075
rect 35996 11067 36000 11075
rect 36004 11067 36016 11075
rect 36020 11067 36032 11075
rect 36036 11067 36040 11075
rect 36060 11067 36064 11075
rect 36068 11067 36072 11075
rect 36184 11067 36188 11075
rect 36192 11067 36196 11075
rect 36216 11067 36220 11075
rect 36224 11067 36228 11075
rect 36240 11067 36252 11075
rect 36256 11067 36268 11075
rect 36280 11067 36284 11075
rect 36288 11067 36292 11075
rect 36304 11067 36316 11075
rect 36320 11067 36332 11075
rect 36344 11067 36348 11075
rect 36352 11067 36356 11075
rect 36376 11067 36380 11075
rect 36384 11067 36396 11075
rect 36408 11067 36412 11075
rect 36416 11067 36420 11075
rect 36500 11067 36504 11075
rect 36508 11067 36512 11075
rect 36532 11067 36536 11075
rect 36540 11067 36544 11075
rect 36640 11067 36644 11075
rect 36648 11067 36652 11075
rect 36664 11067 36676 11075
rect 36680 11067 36684 11075
rect 36704 11067 36708 11075
rect 36712 11067 36724 11075
rect 36732 11067 36748 11075
rect 36756 11067 36780 11075
rect 36800 11067 36808 11075
rect 36828 11067 36840 11075
rect 36852 11067 36856 11075
rect 36860 11067 36872 11075
rect 36876 11067 36880 11075
rect 36944 11067 36948 11075
rect 36952 11067 36964 11075
rect 36968 11067 36972 11075
rect 37012 11067 37024 11075
rect 37036 11067 37040 11075
rect 37044 11067 37056 11075
rect 37060 11067 37064 11075
rect 37076 11067 37088 11075
rect 37128 11067 37132 11075
rect 37136 11067 37148 11075
rect 37152 11067 37156 11075
rect 37168 11067 37180 11075
rect 37192 11067 37196 11075
rect 37200 11067 37212 11075
rect 37228 11067 37252 11075
rect 37260 11067 37276 11075
rect 37292 11067 37308 11075
rect 37324 11067 37328 11075
rect 37332 11067 37344 11075
rect 37348 11067 37360 11075
rect 37364 11067 37368 11075
rect 37388 11067 37392 11075
rect 37396 11067 37400 11075
rect 37412 11067 37424 11075
rect 37428 11067 37432 11075
rect 37448 11067 37464 11075
rect 37480 11067 37528 11075
rect 37544 11067 37592 11075
rect 37608 11067 37612 11075
rect 37616 11067 37620 11075
rect 37640 11067 37644 11075
rect 37648 11067 37660 11075
rect 37672 11067 37676 11075
rect 37680 11067 37684 11075
rect 37704 11067 37708 11075
rect 37712 11067 37724 11075
rect 37728 11067 37740 11075
rect 37744 11067 37748 11075
rect 37768 11067 37772 11075
rect 37776 11067 37780 11075
rect 37796 11067 37812 11075
rect 37820 11067 37844 11075
rect 37860 11067 37872 11075
rect 37876 11067 37880 11075
rect 37892 11067 37904 11075
rect 37912 11067 37936 11075
rect 37952 11067 37964 11075
rect 37968 11067 37972 11075
rect 37984 11067 37996 11075
rect 38008 11067 38012 11075
rect 38016 11067 38028 11075
rect 38032 11067 38036 11075
rect 38048 11067 38060 11075
rect 38140 11067 38152 11075
rect 38164 11067 38168 11075
rect 38172 11067 38184 11075
rect 38188 11067 38192 11075
rect 38204 11067 38216 11075
rect 38228 11067 38232 11075
rect 38236 11067 38248 11075
rect 38264 11067 38288 11075
rect 38296 11067 38312 11075
rect 38328 11067 38344 11075
rect 38360 11067 38364 11075
rect 38368 11067 38380 11075
rect 38384 11067 38396 11075
rect 38400 11067 38404 11075
rect 38424 11067 38428 11075
rect 38432 11067 38436 11075
rect 38456 11067 38460 11075
rect 38464 11067 38468 11075
rect 38488 11067 38492 11075
rect 38496 11067 38500 11075
rect 38520 11067 38524 11075
rect 38528 11067 38540 11075
rect 38544 11067 38556 11075
rect 38560 11067 38564 11075
rect 38660 11067 38664 11075
rect 38668 11067 38672 11075
rect 38752 11067 38756 11075
rect 38760 11067 38764 11075
rect 38844 11067 38848 11075
rect 38852 11067 38856 11075
rect 38876 11067 38880 11075
rect 38884 11067 38888 11075
rect 38900 11067 38912 11075
rect 38916 11067 38920 11075
rect 38940 11067 38944 11075
rect 38948 11067 38960 11075
rect 38968 11067 38984 11075
rect 38992 11067 39004 11075
rect 39008 11067 39012 11075
rect 39028 11067 39052 11075
rect 39060 11067 39076 11075
rect 39084 11067 39108 11075
rect 39120 11067 39144 11075
rect 39152 11067 39168 11075
rect 39176 11067 39200 11075
rect 39216 11067 39220 11075
rect 39224 11067 39236 11075
rect 39240 11067 39252 11075
rect 39256 11067 39260 11075
rect 39280 11067 39284 11075
rect 39288 11067 39292 11075
rect 39388 11067 39392 11075
rect 39396 11067 39408 11075
rect 39412 11067 39424 11075
rect 39428 11067 39432 11075
rect 39452 11067 39456 11075
rect 39460 11067 39472 11075
rect 39476 11067 39488 11075
rect 39492 11067 39496 11075
rect 39516 11067 39520 11075
rect 39524 11067 39528 11075
rect 39540 11067 39552 11075
rect 39556 11067 39560 11075
rect 39580 11067 39584 11075
rect 39588 11067 39592 11075
rect 39604 11067 39616 11075
rect 39620 11067 39632 11075
rect 39644 11067 39648 11075
rect 39652 11067 39656 11075
rect 39676 11067 39680 11075
rect 39684 11067 39696 11075
rect 39708 11067 39712 11075
rect 39716 11067 39720 11075
rect 39800 11067 39804 11075
rect 39808 11067 39812 11075
rect 39892 11067 39896 11075
rect 39900 11067 39904 11075
rect 39924 11067 39928 11075
rect 39932 11067 39936 11075
rect 39948 11067 39960 11075
rect 39964 11067 39968 11075
rect 39988 11067 39992 11075
rect 39996 11067 40000 11075
rect 38784 11057 38792 11065
rect 39136 11057 39144 11065
rect 29408 11037 29416 11045
rect 29920 11037 29928 11045
rect 30048 11037 30056 11045
rect 30384 11037 30392 11045
rect 30672 11037 30680 11045
rect 30816 11037 30824 11045
rect 30960 11037 30968 11045
rect 31184 11037 31192 11045
rect 31520 11037 31528 11045
rect 31536 11037 31544 11045
rect 31696 11037 31704 11045
rect 31904 11037 31912 11045
rect 32288 11037 32296 11045
rect 32848 11037 32856 11045
rect 33232 11037 33240 11045
rect 33568 11037 33576 11045
rect 34144 11037 34152 11045
rect 34416 11037 34424 11045
rect 34528 11037 34536 11045
rect 34672 11037 34680 11045
rect 35584 11037 35592 11045
rect 35680 11037 35688 11045
rect 36256 11037 36264 11045
rect 36320 11037 36328 11045
rect 36736 11037 36744 11045
rect 36944 11037 36952 11045
rect 36960 11037 36968 11045
rect 37328 11037 37336 11045
rect 37504 11037 37512 11045
rect 37792 11037 37800 11045
rect 38080 11037 38088 11045
rect 38480 11037 38488 11045
rect 39360 11037 39368 11045
rect 39520 11037 39528 11045
rect 39664 11037 39672 11045
rect 39984 11037 39992 11045
rect 29424 11017 29432 11025
rect 29600 11017 29608 11025
rect 29728 11017 29736 11025
rect 30624 11017 30632 11025
rect 31168 11017 31176 11025
rect 32240 11017 32248 11025
rect 32272 11017 32280 11025
rect 32320 11017 32328 11025
rect 33440 11017 33448 11025
rect 33856 11017 33864 11025
rect 34720 11017 34728 11025
rect 29616 10997 29624 11005
rect 30464 10997 30472 11005
rect 30640 10997 30648 11005
rect 30864 10997 30872 11005
rect 31616 10997 31624 11005
rect 34320 10997 34328 11005
rect 34816 10997 34824 11005
rect 35184 10997 35192 11005
rect 35328 10997 35336 11005
rect 37104 10997 37112 11005
rect 37248 10997 37256 11005
rect 37984 10997 37992 11005
rect 38432 10997 38440 11005
rect 38608 10997 38616 11005
rect 38880 10997 38888 11005
rect 39232 10997 39240 11005
rect 35600 10977 35608 10985
rect 29568 10957 29576 10965
rect 29648 10957 29656 10965
rect 29760 10957 29768 10965
rect 29824 10957 29832 10965
rect 29904 10957 29912 10965
rect 30128 10957 30136 10965
rect 30784 10957 30792 10965
rect 30928 10957 30936 10965
rect 31008 10957 31016 10965
rect 32272 10957 32280 10965
rect 32480 10957 32488 10965
rect 32736 10957 32744 10965
rect 32816 10957 32824 10965
rect 32928 10957 32936 10965
rect 33072 10957 33080 10965
rect 33344 10957 33352 10965
rect 33536 10957 33544 10965
rect 33648 10957 33656 10965
rect 34288 10957 34296 10965
rect 35168 10957 35176 10965
rect 35200 10957 35208 10965
rect 35632 10957 35640 10965
rect 36816 10957 36824 10965
rect 36992 10957 37000 10965
rect 38032 10957 38040 10965
rect 38144 10957 38152 10965
rect 38592 10957 38600 10965
rect 38768 10957 38776 10965
rect 39840 10957 39848 10965
rect 32944 10937 32952 10945
rect 39152 10937 39160 10945
rect 31088 10917 31096 10925
rect 34288 10917 34296 10925
rect 34560 10877 34568 10885
rect 29380 10867 29392 10875
rect 29412 10867 29424 10875
rect 29428 10867 29432 10875
rect 29448 10867 29464 10875
rect 29480 10867 29512 10875
rect 29528 10867 29540 10875
rect 29544 10867 29548 10875
rect 29568 10867 29572 10875
rect 29576 10867 29588 10875
rect 29604 10867 29616 10875
rect 29620 10867 29624 10875
rect 29644 10867 29648 10875
rect 29652 10867 29664 10875
rect 29680 10867 29704 10875
rect 29720 10867 29724 10875
rect 29728 10867 29740 10875
rect 29744 10867 29748 10875
rect 29796 10867 29800 10875
rect 29804 10867 29816 10875
rect 29820 10867 29832 10875
rect 29888 10867 29892 10875
rect 29896 10867 29908 10875
rect 29920 10867 29924 10875
rect 29928 10867 29932 10875
rect 30184 10867 30188 10875
rect 30192 10867 30196 10875
rect 30344 10867 30356 10875
rect 30368 10867 30372 10875
rect 30376 10867 30388 10875
rect 30392 10867 30396 10875
rect 30412 10867 30428 10875
rect 30444 10867 30448 10875
rect 30452 10867 30464 10875
rect 30468 10867 30472 10875
rect 30492 10867 30496 10875
rect 30500 10867 30512 10875
rect 30516 10867 30528 10875
rect 30576 10867 30588 10875
rect 30592 10867 30604 10875
rect 30624 10867 30636 10875
rect 30648 10867 30652 10875
rect 30656 10867 30668 10875
rect 30688 10867 30700 10875
rect 30720 10867 30732 10875
rect 30736 10867 30740 10875
rect 30756 10867 30772 10875
rect 30788 10867 30828 10875
rect 30844 10867 30848 10875
rect 30852 10867 30856 10875
rect 30868 10867 30880 10875
rect 30892 10867 30896 10875
rect 30900 10867 30904 10875
rect 30984 10867 30988 10875
rect 30992 10867 30996 10875
rect 31016 10867 31020 10875
rect 31024 10867 31028 10875
rect 31040 10867 31052 10875
rect 31060 10867 31076 10875
rect 31092 10867 31124 10875
rect 31140 10867 31156 10875
rect 31168 10867 31200 10875
rect 31208 10867 31224 10875
rect 31240 10867 31244 10875
rect 31248 10867 31252 10875
rect 31272 10867 31276 10875
rect 31280 10867 31292 10875
rect 31304 10867 31308 10875
rect 31312 10867 31316 10875
rect 31572 10867 31576 10875
rect 31580 10867 31584 10875
rect 31604 10867 31608 10875
rect 31612 10867 31616 10875
rect 31696 10867 31700 10875
rect 31704 10867 31708 10875
rect 31720 10867 31732 10875
rect 31736 10867 31740 10875
rect 31760 10867 31764 10875
rect 31768 10867 31772 10875
rect 31792 10867 31796 10875
rect 31800 10867 31812 10875
rect 31824 10867 31828 10875
rect 31832 10867 31836 10875
rect 31856 10867 31860 10875
rect 31864 10867 31868 10875
rect 31880 10867 31892 10875
rect 31896 10867 31900 10875
rect 31920 10867 31924 10875
rect 31928 10867 31932 10875
rect 31952 10867 31956 10875
rect 31960 10867 31972 10875
rect 31984 10867 31988 10875
rect 31992 10867 31996 10875
rect 32124 10867 32128 10875
rect 32132 10867 32136 10875
rect 32392 10867 32396 10875
rect 32400 10867 32404 10875
rect 32416 10867 32428 10875
rect 32432 10867 32436 10875
rect 32452 10867 32468 10875
rect 32484 10867 32500 10875
rect 32508 10867 32540 10875
rect 32548 10867 32564 10875
rect 32580 10867 32592 10875
rect 32604 10867 32608 10875
rect 32612 10867 32624 10875
rect 32760 10867 32764 10875
rect 32768 10867 32780 10875
rect 32784 10867 32788 10875
rect 32800 10867 32812 10875
rect 32824 10867 32828 10875
rect 32832 10867 32844 10875
rect 32860 10867 32884 10875
rect 32892 10867 32908 10875
rect 32924 10867 32928 10875
rect 32932 10867 32936 10875
rect 32956 10867 32960 10875
rect 32964 10867 32976 10875
rect 32980 10867 32992 10875
rect 32996 10867 33000 10875
rect 33020 10867 33024 10875
rect 33028 10867 33040 10875
rect 33044 10867 33056 10875
rect 33060 10867 33064 10875
rect 33084 10867 33088 10875
rect 33092 10867 33096 10875
rect 33112 10867 33116 10875
rect 33120 10867 33132 10875
rect 33136 10867 33148 10875
rect 33152 10867 33156 10875
rect 33176 10867 33180 10875
rect 33184 10867 33188 10875
rect 33204 10867 33220 10875
rect 33228 10867 33252 10875
rect 33268 10867 33292 10875
rect 33300 10867 33312 10875
rect 33320 10867 33344 10875
rect 33360 10867 33384 10875
rect 33392 10867 33404 10875
rect 33416 10867 33420 10875
rect 33424 10867 33436 10875
rect 33440 10867 33444 10875
rect 33456 10867 33468 10875
rect 33580 10867 33592 10875
rect 33596 10867 33600 10875
rect 33612 10867 33624 10875
rect 33640 10867 33656 10875
rect 33664 10867 33696 10875
rect 33704 10867 33720 10875
rect 33736 10867 33740 10875
rect 33744 10867 33748 10875
rect 33768 10867 33772 10875
rect 33776 10867 33788 10875
rect 33800 10867 33804 10875
rect 33808 10867 33812 10875
rect 33824 10867 33836 10875
rect 33840 10867 33844 10875
rect 33940 10867 33944 10875
rect 33948 10867 33952 10875
rect 33964 10867 33976 10875
rect 33980 10867 33992 10875
rect 34000 10867 34016 10875
rect 34032 10867 34080 10875
rect 34096 10867 34108 10875
rect 34112 10867 34116 10875
rect 34128 10867 34140 10875
rect 34152 10867 34156 10875
rect 34160 10867 34172 10875
rect 34276 10867 34280 10875
rect 34284 10867 34296 10875
rect 34316 10867 34328 10875
rect 34332 10867 34344 10875
rect 34348 10867 34360 10875
rect 34380 10867 34392 10875
rect 34400 10867 34432 10875
rect 34440 10867 34456 10875
rect 34464 10867 34476 10875
rect 34480 10867 34484 10875
rect 34504 10867 34508 10875
rect 34512 10867 34524 10875
rect 34532 10867 34548 10875
rect 34556 10867 34580 10875
rect 34596 10867 34600 10875
rect 34604 10867 34616 10875
rect 34620 10867 34632 10875
rect 34636 10867 34640 10875
rect 34660 10867 34664 10875
rect 34668 10867 34672 10875
rect 34736 10867 34740 10875
rect 34744 10867 34756 10875
rect 34768 10867 34772 10875
rect 34776 10867 34780 10875
rect 34792 10867 34804 10875
rect 34808 10867 34812 10875
rect 34832 10867 34836 10875
rect 34840 10867 34844 10875
rect 34860 10867 34876 10875
rect 34884 10867 34916 10875
rect 34924 10867 34940 10875
rect 34956 10867 34968 10875
rect 34972 10867 34984 10875
rect 34996 10867 35000 10875
rect 35004 10867 35008 10875
rect 35020 10867 35032 10875
rect 35036 10867 35040 10875
rect 35136 10867 35140 10875
rect 35144 10867 35148 10875
rect 35160 10867 35172 10875
rect 35176 10867 35188 10875
rect 35200 10867 35204 10875
rect 35208 10867 35212 10875
rect 35228 10867 35276 10875
rect 35292 10867 35308 10875
rect 35324 10867 35328 10875
rect 35332 10867 35344 10875
rect 35356 10867 35360 10875
rect 35364 10867 35368 10875
rect 35388 10867 35392 10875
rect 35396 10867 35400 10875
rect 35412 10867 35424 10875
rect 35428 10867 35432 10875
rect 35448 10867 35464 10875
rect 35480 10867 35528 10875
rect 35544 10867 35560 10875
rect 35576 10867 35588 10875
rect 35600 10867 35604 10875
rect 35608 10867 35620 10875
rect 35640 10867 35652 10875
rect 35656 10867 35660 10875
rect 36084 10867 36096 10875
rect 36100 10867 36112 10875
rect 36116 10867 36128 10875
rect 36148 10867 36160 10875
rect 36172 10867 36176 10875
rect 36180 10867 36192 10875
rect 36212 10867 36224 10875
rect 36244 10867 36256 10875
rect 36260 10867 36264 10875
rect 36276 10867 36288 10875
rect 36308 10867 36320 10875
rect 36324 10867 36336 10875
rect 36340 10867 36352 10875
rect 36424 10867 36428 10875
rect 36432 10867 36444 10875
rect 36556 10867 36568 10875
rect 36572 10867 36584 10875
rect 36588 10867 36600 10875
rect 36620 10867 36632 10875
rect 36648 10867 36672 10875
rect 36680 10867 36696 10875
rect 36712 10867 36728 10875
rect 36736 10867 36748 10875
rect 36752 10867 36764 10875
rect 36776 10867 36780 10875
rect 36784 10867 36788 10875
rect 36884 10867 36888 10875
rect 36892 10867 36904 10875
rect 36916 10867 36920 10875
rect 36924 10867 36928 10875
rect 36940 10867 36952 10875
rect 36956 10867 36968 10875
rect 36976 10867 36992 10875
rect 37008 10867 37056 10875
rect 37072 10867 37076 10875
rect 37080 10867 37084 10875
rect 37100 10867 37148 10875
rect 37164 10867 37168 10875
rect 37172 10867 37176 10875
rect 37188 10867 37200 10875
rect 37204 10867 37216 10875
rect 37228 10867 37232 10875
rect 37236 10867 37240 10875
rect 37260 10867 37264 10875
rect 37268 10867 37272 10875
rect 37292 10867 37296 10875
rect 37300 10867 37304 10875
rect 37324 10867 37328 10875
rect 37332 10867 37336 10875
rect 37348 10867 37360 10875
rect 37364 10867 37376 10875
rect 37388 10867 37392 10875
rect 37396 10867 37400 10875
rect 37448 10867 37452 10875
rect 37456 10867 37468 10875
rect 37480 10867 37484 10875
rect 37488 10867 37492 10875
rect 37504 10867 37516 10875
rect 37520 10867 37532 10875
rect 37544 10867 37548 10875
rect 37552 10867 37556 10875
rect 37568 10867 37580 10875
rect 37584 10867 37588 10875
rect 37684 10867 37688 10875
rect 37692 10867 37696 10875
rect 37708 10867 37720 10875
rect 37724 10867 37736 10875
rect 37748 10867 37752 10875
rect 37756 10867 37760 10875
rect 37780 10867 37784 10875
rect 37788 10867 37792 10875
rect 37856 10867 37860 10875
rect 37864 10867 37876 10875
rect 37888 10867 37892 10875
rect 37896 10867 37900 10875
rect 37948 10867 37952 10875
rect 37956 10867 37968 10875
rect 37988 10867 38000 10875
rect 38004 10867 38008 10875
rect 38020 10867 38032 10875
rect 38052 10867 38064 10875
rect 38080 10867 38120 10875
rect 38136 10867 38148 10875
rect 38152 10867 38156 10875
rect 38176 10867 38180 10875
rect 38184 10867 38196 10875
rect 38204 10867 38220 10875
rect 38228 10867 38244 10875
rect 38260 10867 38272 10875
rect 38284 10867 38288 10875
rect 38292 10867 38304 10875
rect 38324 10867 38336 10875
rect 38392 10867 38396 10875
rect 38400 10867 38404 10875
rect 38424 10867 38428 10875
rect 38432 10867 38436 10875
rect 38448 10867 38460 10875
rect 38476 10867 38492 10875
rect 38508 10867 38540 10875
rect 38548 10867 38560 10875
rect 38576 10867 38592 10875
rect 38600 10867 38632 10875
rect 38640 10867 38656 10875
rect 38668 10867 38684 10875
rect 38692 10867 38724 10875
rect 38732 10867 38748 10875
rect 38764 10867 38768 10875
rect 38772 10867 38776 10875
rect 38796 10867 38800 10875
rect 38804 10867 38816 10875
rect 38828 10867 38832 10875
rect 38836 10867 38840 10875
rect 38968 10867 38972 10875
rect 38976 10867 38980 10875
rect 38992 10867 39004 10875
rect 39008 10867 39020 10875
rect 39028 10867 39044 10875
rect 39060 10867 39064 10875
rect 39068 10867 39072 10875
rect 39084 10867 39096 10875
rect 39100 10867 39112 10875
rect 39120 10867 39136 10875
rect 39152 10867 39156 10875
rect 39160 10867 39164 10875
rect 39176 10867 39188 10875
rect 39192 10867 39200 10875
rect 39216 10867 39220 10875
rect 39224 10867 39228 10875
rect 39240 10867 39252 10875
rect 39256 10867 39268 10875
rect 39280 10867 39284 10875
rect 39288 10867 39292 10875
rect 39312 10867 39316 10875
rect 39320 10867 39324 10875
rect 39420 10867 39424 10875
rect 39428 10867 39432 10875
rect 39444 10867 39456 10875
rect 39460 10867 39472 10875
rect 39484 10867 39488 10875
rect 39492 10867 39496 10875
rect 39516 10867 39520 10875
rect 39524 10867 39528 10875
rect 39548 10867 39552 10875
rect 39556 10867 39560 10875
rect 39580 10867 39584 10875
rect 39588 10867 39592 10875
rect 39604 10867 39616 10875
rect 39620 10867 39632 10875
rect 39644 10867 39648 10875
rect 39652 10867 39656 10875
rect 39676 10867 39680 10875
rect 39684 10867 39696 10875
rect 39708 10867 39712 10875
rect 39716 10867 39720 10875
rect 39816 10867 39820 10875
rect 39824 10867 39836 10875
rect 39848 10867 39852 10875
rect 39856 10867 39860 10875
rect 39872 10867 39884 10875
rect 39888 10867 39892 10875
rect 39912 10867 39916 10875
rect 39920 10867 39924 10875
rect 39944 10867 39948 10875
rect 39952 10867 39956 10875
rect 39976 10867 39980 10875
rect 39984 10867 39996 10875
rect 36176 10837 36184 10845
rect 32304 10817 32312 10825
rect 37520 10817 37528 10825
rect 39264 10817 39272 10825
rect 29968 10797 29976 10805
rect 33296 10797 33304 10805
rect 38512 10797 38520 10805
rect 29392 10777 29400 10785
rect 29872 10777 29880 10785
rect 29952 10777 29960 10785
rect 30288 10777 30296 10785
rect 30560 10777 30568 10785
rect 32128 10777 32136 10785
rect 32160 10777 32168 10785
rect 32832 10777 32840 10785
rect 33168 10777 33176 10785
rect 33456 10777 33464 10785
rect 34496 10777 34504 10785
rect 35632 10777 35640 10785
rect 37120 10777 37128 10785
rect 37632 10777 37640 10785
rect 37680 10777 37688 10785
rect 38176 10777 38184 10785
rect 38560 10777 38568 10785
rect 39168 10777 39176 10785
rect 31264 10757 31272 10765
rect 35104 10757 35112 10765
rect 35392 10757 35400 10765
rect 35888 10757 35896 10765
rect 39520 10757 39528 10765
rect 39632 10757 39640 10765
rect 39648 10757 39656 10765
rect 29968 10737 29976 10745
rect 30064 10737 30072 10745
rect 30304 10737 30312 10745
rect 30576 10737 30584 10745
rect 32656 10737 32664 10745
rect 33888 10737 33896 10745
rect 34464 10737 34472 10745
rect 35264 10737 35272 10745
rect 36640 10737 36648 10745
rect 37120 10737 37128 10745
rect 37440 10737 37448 10745
rect 37952 10737 37960 10745
rect 30016 10717 30024 10725
rect 30352 10717 30360 10725
rect 30720 10717 30728 10725
rect 30800 10717 30808 10725
rect 30912 10717 30920 10725
rect 30992 10717 31000 10725
rect 31392 10717 31400 10725
rect 31472 10717 31480 10725
rect 32352 10717 32360 10725
rect 32480 10717 32488 10725
rect 32736 10717 32744 10725
rect 32912 10717 32920 10725
rect 33392 10717 33400 10725
rect 33552 10717 33560 10725
rect 33680 10717 33688 10725
rect 34048 10717 34056 10725
rect 35376 10717 35384 10725
rect 36624 10717 36632 10725
rect 37008 10717 37016 10725
rect 37328 10717 37336 10725
rect 38368 10717 38376 10725
rect 39616 10717 39624 10725
rect 31736 10705 31737 10710
rect 29712 10697 29720 10705
rect 32576 10697 32584 10705
rect 33840 10697 33848 10705
rect 35008 10697 35016 10705
rect 35088 10697 35096 10705
rect 35696 10697 35704 10705
rect 39984 10697 39992 10705
rect 35472 10677 35480 10685
rect 37680 10677 37688 10685
rect 37808 10677 37816 10685
rect 38544 10677 38552 10685
rect 29380 10667 29392 10675
rect 29412 10667 29424 10675
rect 29428 10667 29432 10675
rect 29448 10667 29464 10675
rect 29480 10667 29512 10675
rect 29528 10667 29540 10675
rect 29560 10667 29572 10675
rect 29584 10667 29588 10675
rect 29592 10667 29596 10675
rect 29708 10667 29712 10675
rect 29716 10667 29728 10675
rect 29732 10667 29736 10675
rect 29752 10667 29768 10675
rect 29784 10667 29788 10675
rect 29792 10667 29804 10675
rect 29808 10667 29820 10675
rect 29824 10667 29828 10675
rect 29844 10667 29860 10675
rect 29876 10667 29892 10675
rect 29900 10667 29924 10675
rect 29940 10667 29952 10675
rect 29956 10667 29960 10675
rect 29972 10667 29984 10675
rect 29992 10667 30008 10675
rect 30024 10667 30072 10675
rect 30088 10667 30100 10675
rect 30116 10667 30164 10675
rect 30180 10667 30196 10675
rect 30212 10667 30216 10675
rect 30220 10667 30232 10675
rect 30244 10667 30248 10675
rect 30252 10667 30256 10675
rect 30540 10667 30544 10675
rect 30548 10667 30552 10675
rect 30572 10667 30576 10675
rect 30580 10667 30584 10675
rect 30596 10667 30608 10675
rect 30620 10667 30624 10675
rect 30628 10667 30640 10675
rect 30644 10667 30648 10675
rect 30752 10667 30764 10675
rect 30784 10667 30796 10675
rect 30800 10667 30812 10675
rect 30816 10667 30828 10675
rect 30844 10667 30860 10675
rect 30868 10667 30884 10675
rect 30892 10667 30908 10675
rect 30916 10667 30928 10675
rect 30948 10667 30960 10675
rect 30972 10667 30976 10675
rect 30980 10667 30984 10675
rect 31064 10667 31068 10675
rect 31072 10667 31076 10675
rect 31096 10667 31100 10675
rect 31104 10667 31116 10675
rect 31120 10667 31124 10675
rect 31144 10667 31148 10675
rect 31152 10667 31156 10675
rect 31172 10667 31176 10675
rect 31180 10667 31192 10675
rect 31196 10667 31200 10675
rect 31220 10667 31224 10675
rect 31228 10667 31232 10675
rect 31248 10667 31264 10675
rect 31272 10667 31296 10675
rect 31312 10667 31336 10675
rect 31344 10667 31356 10675
rect 31368 10667 31372 10675
rect 31376 10667 31388 10675
rect 31408 10667 31420 10675
rect 31492 10667 31496 10675
rect 31500 10667 31512 10675
rect 31532 10667 31544 10675
rect 31548 10667 31560 10675
rect 31564 10667 31576 10675
rect 31596 10667 31608 10675
rect 31624 10667 31636 10675
rect 31640 10667 31652 10675
rect 31656 10667 31668 10675
rect 31688 10667 31700 10675
rect 31704 10667 31708 10675
rect 31720 10667 31732 10675
rect 31748 10667 31764 10675
rect 31780 10667 31828 10675
rect 31844 10667 31860 10675
rect 31876 10667 31880 10675
rect 31884 10667 31896 10675
rect 31908 10667 31912 10675
rect 31916 10667 31920 10675
rect 31940 10667 31944 10675
rect 31948 10667 31960 10675
rect 31964 10667 31976 10675
rect 31980 10667 31984 10675
rect 32000 10667 32016 10675
rect 32032 10667 32036 10675
rect 32040 10667 32052 10675
rect 32056 10667 32068 10675
rect 32072 10667 32076 10675
rect 32124 10667 32128 10675
rect 32132 10667 32144 10675
rect 32148 10667 32160 10675
rect 32164 10667 32168 10675
rect 32188 10667 32192 10675
rect 32196 10667 32200 10675
rect 32264 10667 32268 10675
rect 32272 10667 32276 10675
rect 32296 10667 32300 10675
rect 32304 10667 32316 10675
rect 32320 10667 32332 10675
rect 32336 10667 32340 10675
rect 32360 10667 32364 10675
rect 32368 10667 32380 10675
rect 32388 10667 32404 10675
rect 32412 10667 32436 10675
rect 32452 10667 32464 10675
rect 32484 10667 32496 10675
rect 32508 10667 32512 10675
rect 32516 10667 32528 10675
rect 32532 10667 32536 10675
rect 32548 10667 32560 10675
rect 32640 10667 32652 10675
rect 32672 10667 32684 10675
rect 32688 10667 32700 10675
rect 32704 10667 32716 10675
rect 32732 10667 32748 10675
rect 32756 10667 32788 10675
rect 32800 10667 32812 10675
rect 32820 10667 32844 10675
rect 32860 10667 32864 10675
rect 32868 10667 32880 10675
rect 32892 10667 32896 10675
rect 32900 10667 32904 10675
rect 33032 10667 33036 10675
rect 33040 10667 33052 10675
rect 33056 10667 33068 10675
rect 33072 10667 33076 10675
rect 33096 10667 33100 10675
rect 33104 10667 33108 10675
rect 33124 10667 33128 10675
rect 33132 10667 33144 10675
rect 33148 10667 33160 10675
rect 33164 10667 33168 10675
rect 33188 10667 33192 10675
rect 33196 10667 33200 10675
rect 33296 10667 33300 10675
rect 33304 10667 33316 10675
rect 33320 10667 33332 10675
rect 33336 10667 33340 10675
rect 33360 10667 33364 10675
rect 33368 10667 33380 10675
rect 33388 10667 33404 10675
rect 33412 10667 33436 10675
rect 33452 10667 33456 10675
rect 33460 10667 33472 10675
rect 33480 10667 33496 10675
rect 33504 10667 33528 10675
rect 33544 10667 33548 10675
rect 33552 10667 33564 10675
rect 33576 10667 33580 10675
rect 33584 10667 33588 10675
rect 33608 10667 33612 10675
rect 33616 10667 33620 10675
rect 33716 10667 33720 10675
rect 33724 10667 33728 10675
rect 33740 10667 33752 10675
rect 33756 10667 33760 10675
rect 33780 10667 33784 10675
rect 33788 10667 33792 10675
rect 33808 10667 33856 10675
rect 33872 10667 33888 10675
rect 33904 10667 33916 10675
rect 33928 10667 33932 10675
rect 33936 10667 33948 10675
rect 33968 10667 33980 10675
rect 33984 10667 33996 10675
rect 34000 10667 34012 10675
rect 34156 10667 34168 10675
rect 34172 10667 34176 10675
rect 34188 10667 34200 10675
rect 34220 10667 34232 10675
rect 34236 10667 34240 10675
rect 34252 10667 34264 10675
rect 34272 10667 34296 10675
rect 34312 10667 34360 10675
rect 34376 10667 34392 10675
rect 34400 10667 34412 10675
rect 34416 10667 34428 10675
rect 34440 10667 34444 10675
rect 34448 10667 34452 10675
rect 34464 10667 34476 10675
rect 34480 10667 34484 10675
rect 34532 10667 34536 10675
rect 34540 10667 34544 10675
rect 34556 10667 34568 10675
rect 34572 10667 34576 10675
rect 34596 10667 34600 10675
rect 34604 10667 34608 10675
rect 34620 10667 34632 10675
rect 34636 10667 34640 10675
rect 34660 10667 34664 10675
rect 34668 10667 34680 10675
rect 34684 10667 34696 10675
rect 34700 10667 34704 10675
rect 34724 10667 34728 10675
rect 34732 10667 34736 10675
rect 34832 10667 34836 10675
rect 34840 10667 34844 10675
rect 34856 10667 34868 10675
rect 34872 10667 34876 10675
rect 34892 10667 34916 10675
rect 34924 10667 34940 10675
rect 34948 10667 34980 10675
rect 34996 10667 35012 10675
rect 35020 10667 35032 10675
rect 35036 10667 35048 10675
rect 35060 10667 35064 10675
rect 35068 10667 35072 10675
rect 35092 10667 35096 10675
rect 35100 10667 35104 10675
rect 35168 10667 35172 10675
rect 35176 10667 35188 10675
rect 35200 10667 35204 10675
rect 35208 10667 35212 10675
rect 35224 10667 35236 10675
rect 35240 10667 35252 10675
rect 35264 10667 35268 10675
rect 35272 10667 35276 10675
rect 35292 10667 35308 10675
rect 35316 10667 35328 10675
rect 35332 10667 35344 10675
rect 35356 10667 35360 10675
rect 35364 10667 35368 10675
rect 35384 10667 35400 10675
rect 35408 10667 35432 10675
rect 35448 10667 35460 10675
rect 35480 10667 35492 10675
rect 35496 10667 35508 10675
rect 35512 10667 35524 10675
rect 35544 10667 35556 10675
rect 35660 10667 35664 10675
rect 35668 10667 35680 10675
rect 35684 10667 35688 10675
rect 35700 10667 35712 10675
rect 35728 10667 35744 10675
rect 35760 10667 35784 10675
rect 35792 10667 35808 10675
rect 35816 10667 35828 10675
rect 35832 10667 35836 10675
rect 35856 10667 35860 10675
rect 35864 10667 35876 10675
rect 35880 10667 35892 10675
rect 35896 10667 35900 10675
rect 36028 10667 36032 10675
rect 36036 10667 36040 10675
rect 36052 10667 36064 10675
rect 36068 10667 36072 10675
rect 36088 10667 36112 10675
rect 36120 10667 36136 10675
rect 36144 10667 36176 10675
rect 36184 10667 36196 10675
rect 36216 10667 36228 10675
rect 36240 10667 36244 10675
rect 36248 10667 36260 10675
rect 36280 10667 36292 10675
rect 36304 10667 36308 10675
rect 36312 10667 36324 10675
rect 36328 10667 36332 10675
rect 36344 10667 36356 10675
rect 36364 10667 36388 10675
rect 36404 10667 36416 10675
rect 36420 10667 36424 10675
rect 36436 10667 36448 10675
rect 36456 10667 36480 10675
rect 36496 10667 36520 10675
rect 36528 10667 36540 10675
rect 36552 10667 36556 10675
rect 36560 10667 36572 10675
rect 36576 10667 36580 10675
rect 36592 10667 36604 10675
rect 36684 10667 36696 10675
rect 36716 10667 36728 10675
rect 36732 10667 36744 10675
rect 36748 10667 36760 10675
rect 36780 10667 36792 10675
rect 36808 10667 36832 10675
rect 36840 10667 36856 10675
rect 36872 10667 36876 10675
rect 36880 10667 36884 10675
rect 36896 10667 36908 10675
rect 36912 10667 36924 10675
rect 36936 10667 36940 10675
rect 36944 10667 36948 10675
rect 36960 10667 36972 10675
rect 36976 10667 36980 10675
rect 37000 10667 37004 10675
rect 37008 10667 37012 10675
rect 37024 10667 37036 10675
rect 37040 10667 37044 10675
rect 37060 10667 37084 10675
rect 37092 10667 37108 10675
rect 37116 10667 37128 10675
rect 37132 10667 37136 10675
rect 37152 10667 37176 10675
rect 37184 10667 37200 10675
rect 37208 10667 37232 10675
rect 37248 10667 37252 10675
rect 37256 10667 37268 10675
rect 37280 10667 37284 10675
rect 37288 10667 37292 10675
rect 37668 10667 37672 10675
rect 37676 10667 37680 10675
rect 37888 10667 37892 10675
rect 37896 10667 37900 10675
rect 37964 10667 37968 10675
rect 37972 10667 37976 10675
rect 37988 10667 38000 10675
rect 38020 10667 38032 10675
rect 38048 10667 38072 10675
rect 38080 10667 38096 10675
rect 38104 10667 38120 10675
rect 38136 10667 38148 10675
rect 38152 10667 38164 10675
rect 38184 10667 38196 10675
rect 38212 10667 38236 10675
rect 38252 10667 38268 10675
rect 38284 10667 38308 10675
rect 38324 10667 38336 10675
rect 38356 10667 38368 10675
rect 38372 10667 38384 10675
rect 38400 10667 38412 10675
rect 38432 10667 38444 10675
rect 38448 10667 38460 10675
rect 38468 10667 38484 10675
rect 38500 10667 38516 10675
rect 38524 10667 38536 10675
rect 38544 10667 38568 10675
rect 38584 10667 38596 10675
rect 38600 10667 38604 10675
rect 38616 10667 38628 10675
rect 38640 10667 38644 10675
rect 38648 10667 38660 10675
rect 38676 10667 38700 10675
rect 38708 10667 38720 10675
rect 38732 10667 38736 10675
rect 38740 10667 38752 10675
rect 38772 10667 38784 10675
rect 38896 10667 38908 10675
rect 38912 10667 38916 10675
rect 38928 10667 38940 10675
rect 38960 10667 38972 10675
rect 38976 10667 38980 10675
rect 38992 10667 39004 10675
rect 39016 10667 39020 10675
rect 39024 10667 39036 10675
rect 39052 10667 39064 10675
rect 39068 10667 39072 10675
rect 39084 10667 39096 10675
rect 39108 10667 39112 10675
rect 39116 10667 39128 10675
rect 39304 10667 39316 10675
rect 39320 10667 39324 10675
rect 39428 10667 39440 10675
rect 39444 10667 39448 10675
rect 39552 10667 39564 10675
rect 39568 10667 39572 10675
rect 39584 10667 39596 10675
rect 39608 10667 39612 10675
rect 39616 10667 39628 10675
rect 39644 10667 39668 10675
rect 39676 10667 39692 10675
rect 39708 10667 39712 10675
rect 39716 10667 39720 10675
rect 39740 10667 39744 10675
rect 39748 10667 39760 10675
rect 39764 10667 39776 10675
rect 39780 10667 39784 10675
rect 39804 10667 39808 10675
rect 39812 10667 39816 10675
rect 39912 10667 39916 10675
rect 39920 10667 39924 10675
rect 39936 10667 39948 10675
rect 39952 10667 39956 10675
rect 39976 10667 39980 10675
rect 39984 10667 39996 10675
rect 34256 10657 34264 10665
rect 29888 10637 29896 10645
rect 33984 10637 33992 10645
rect 35664 10637 35672 10645
rect 35872 10637 35880 10645
rect 36240 10637 36248 10645
rect 37056 10637 37064 10645
rect 37648 10637 37656 10645
rect 37776 10637 37784 10645
rect 39840 10637 39848 10645
rect 29904 10617 29912 10625
rect 30208 10617 30216 10625
rect 30288 10617 30296 10625
rect 36304 10617 36312 10625
rect 36352 10617 36360 10625
rect 37568 10617 37576 10625
rect 38208 10617 38216 10625
rect 38256 10617 38264 10625
rect 38272 10617 38280 10625
rect 38368 10617 38376 10625
rect 38912 10617 38920 10625
rect 39104 10617 39112 10625
rect 39232 10617 39240 10625
rect 29728 10597 29736 10605
rect 30240 10597 30248 10605
rect 30784 10597 30792 10605
rect 30880 10597 30888 10605
rect 31296 10597 31304 10605
rect 32528 10597 32536 10605
rect 32800 10597 32808 10605
rect 35248 10597 35256 10605
rect 35488 10597 35496 10605
rect 35616 10597 35624 10605
rect 35856 10597 35864 10605
rect 35984 10597 35992 10605
rect 36480 10597 36488 10605
rect 37712 10597 37720 10605
rect 37792 10597 37800 10605
rect 39488 10597 39496 10605
rect 39728 10597 39736 10605
rect 29584 10577 29592 10585
rect 29872 10577 29880 10585
rect 30848 10577 30856 10585
rect 31504 10577 31512 10585
rect 32976 10577 32984 10585
rect 34416 10577 34424 10585
rect 38220 10584 38222 10585
rect 38220 10577 38222 10578
rect 39408 10577 39416 10585
rect 30928 10557 30936 10565
rect 32544 10557 32552 10565
rect 32656 10557 32664 10565
rect 33504 10557 33512 10565
rect 33680 10557 33688 10565
rect 34288 10557 34296 10565
rect 34704 10557 34712 10565
rect 34784 10557 34792 10565
rect 35344 10557 35352 10565
rect 35536 10557 35544 10565
rect 35632 10557 35640 10565
rect 35744 10557 35752 10565
rect 36000 10557 36008 10565
rect 36496 10557 36504 10565
rect 37376 10557 37384 10565
rect 37936 10557 37944 10565
rect 38000 10557 38008 10565
rect 38096 10557 38104 10565
rect 38768 10557 38776 10565
rect 38992 10557 39000 10565
rect 39424 10557 39432 10565
rect 30496 10517 30504 10525
rect 31216 10517 31224 10525
rect 29644 10467 29648 10475
rect 29652 10467 29664 10475
rect 29684 10467 29696 10475
rect 29700 10467 29712 10475
rect 29716 10467 29728 10475
rect 29744 10467 29760 10475
rect 29776 10467 29788 10475
rect 29792 10467 29804 10475
rect 29808 10467 29820 10475
rect 29840 10467 29852 10475
rect 29872 10467 29884 10475
rect 29904 10467 29916 10475
rect 29936 10467 29948 10475
rect 29952 10467 29964 10475
rect 29968 10467 29980 10475
rect 29996 10467 30008 10475
rect 30028 10467 30040 10475
rect 30044 10467 30056 10475
rect 30060 10467 30072 10475
rect 30248 10467 30260 10475
rect 30280 10467 30292 10475
rect 30296 10467 30308 10475
rect 30312 10467 30324 10475
rect 30344 10467 30356 10475
rect 30368 10467 30372 10475
rect 30376 10467 30388 10475
rect 30408 10467 30420 10475
rect 30660 10467 30672 10475
rect 30684 10467 30688 10475
rect 30692 10467 30704 10475
rect 30708 10467 30712 10475
rect 30752 10467 30764 10475
rect 30776 10467 30780 10475
rect 30784 10467 30796 10475
rect 30800 10467 30804 10475
rect 30816 10467 30828 10475
rect 30836 10467 30852 10475
rect 30868 10467 30884 10475
rect 30892 10467 30908 10475
rect 30924 10467 30928 10475
rect 30932 10467 30936 10475
rect 30956 10467 30960 10475
rect 30964 10467 30976 10475
rect 30980 10467 30984 10475
rect 31000 10467 31004 10475
rect 31008 10467 31012 10475
rect 31032 10467 31036 10475
rect 31040 10467 31052 10475
rect 31056 10467 31060 10475
rect 31172 10467 31176 10475
rect 31180 10467 31184 10475
rect 31200 10467 31208 10475
rect 31220 10467 31224 10475
rect 31228 10467 31240 10475
rect 31256 10467 31280 10475
rect 31288 10467 31304 10475
rect 31320 10467 31336 10475
rect 31352 10467 31356 10475
rect 31360 10467 31372 10475
rect 31376 10467 31388 10475
rect 31392 10467 31396 10475
rect 31412 10467 31428 10475
rect 31444 10467 31448 10475
rect 31452 10467 31464 10475
rect 31468 10467 31480 10475
rect 31484 10467 31488 10475
rect 31536 10467 31540 10475
rect 31544 10467 31556 10475
rect 31560 10467 31572 10475
rect 31576 10467 31580 10475
rect 31600 10467 31604 10475
rect 31608 10467 31612 10475
rect 31740 10467 31744 10475
rect 31748 10467 31752 10475
rect 31772 10467 31776 10475
rect 31780 10467 31784 10475
rect 31796 10467 31808 10475
rect 31812 10467 31816 10475
rect 31836 10467 31840 10475
rect 31844 10467 31848 10475
rect 31864 10467 31912 10475
rect 31928 10467 31976 10475
rect 32000 10467 32016 10475
rect 32024 10467 32036 10475
rect 32048 10467 32052 10475
rect 32056 10467 32068 10475
rect 32212 10467 32224 10475
rect 32228 10467 32240 10475
rect 32244 10467 32256 10475
rect 32272 10467 32288 10475
rect 32304 10467 32328 10475
rect 32336 10467 32352 10475
rect 32368 10467 32384 10475
rect 32392 10467 32404 10475
rect 32408 10467 32420 10475
rect 32432 10467 32436 10475
rect 32440 10467 32444 10475
rect 32572 10467 32576 10475
rect 32580 10467 32584 10475
rect 32596 10467 32608 10475
rect 32612 10467 32624 10475
rect 32632 10467 32648 10475
rect 32664 10467 32712 10475
rect 32728 10467 32740 10475
rect 32744 10467 32748 10475
rect 32760 10467 32772 10475
rect 32784 10467 32788 10475
rect 32792 10467 32804 10475
rect 32808 10467 32812 10475
rect 32824 10467 32836 10475
rect 32852 10467 32864 10475
rect 32876 10467 32880 10475
rect 32884 10467 32896 10475
rect 32900 10467 32904 10475
rect 32968 10467 32972 10475
rect 32976 10467 32988 10475
rect 32992 10467 32996 10475
rect 33008 10467 33020 10475
rect 33060 10467 33064 10475
rect 33068 10467 33080 10475
rect 33084 10467 33088 10475
rect 33100 10467 33112 10475
rect 33192 10467 33204 10475
rect 33224 10467 33236 10475
rect 33240 10467 33244 10475
rect 33256 10467 33268 10475
rect 33288 10467 33300 10475
rect 33308 10467 33340 10475
rect 33348 10467 33364 10475
rect 33372 10467 33396 10475
rect 33412 10467 33428 10475
rect 33444 10467 33456 10475
rect 33468 10467 33472 10475
rect 33476 10467 33488 10475
rect 33492 10467 33496 10475
rect 33508 10467 33520 10475
rect 33536 10467 33548 10475
rect 33560 10467 33564 10475
rect 33568 10467 33580 10475
rect 33584 10467 33588 10475
rect 33600 10467 33612 10475
rect 33724 10467 33736 10475
rect 33740 10467 33752 10475
rect 33756 10467 33768 10475
rect 33788 10467 33800 10475
rect 33808 10467 33840 10475
rect 33848 10467 33864 10475
rect 33880 10467 33896 10475
rect 33912 10467 33916 10475
rect 33920 10467 33932 10475
rect 33944 10467 33948 10475
rect 33952 10467 33956 10475
rect 33968 10467 33980 10475
rect 33984 10467 33996 10475
rect 34008 10467 34012 10475
rect 34016 10467 34020 10475
rect 34148 10467 34152 10475
rect 34156 10467 34160 10475
rect 34172 10467 34184 10475
rect 34188 10467 34200 10475
rect 34212 10467 34216 10475
rect 34220 10467 34224 10475
rect 34236 10467 34248 10475
rect 34252 10467 34264 10475
rect 34272 10467 34288 10475
rect 34304 10467 34320 10475
rect 34328 10467 34352 10475
rect 34368 10467 34384 10475
rect 34400 10467 34412 10475
rect 34416 10467 34428 10475
rect 34432 10467 34444 10475
rect 34460 10467 34476 10475
rect 34492 10467 34504 10475
rect 34508 10467 34520 10475
rect 34524 10467 34536 10475
rect 34556 10467 34568 10475
rect 34572 10467 34576 10475
rect 34588 10467 34600 10475
rect 34620 10467 34632 10475
rect 34636 10467 34640 10475
rect 34652 10467 34664 10475
rect 34676 10467 34680 10475
rect 34684 10467 34696 10475
rect 34716 10467 34728 10475
rect 34840 10467 34852 10475
rect 34856 10467 34860 10475
rect 34892 10467 34896 10475
rect 34900 10467 34912 10475
rect 34932 10467 34944 10475
rect 34948 10467 34952 10475
rect 34964 10467 34976 10475
rect 34996 10467 35008 10475
rect 35024 10467 35072 10475
rect 35088 10467 35100 10475
rect 35116 10467 35164 10475
rect 35176 10467 35192 10475
rect 35208 10467 35256 10475
rect 35272 10467 35284 10475
rect 35300 10467 35348 10475
rect 35364 10467 35376 10475
rect 35392 10467 35440 10475
rect 35452 10467 35468 10475
rect 35484 10467 35532 10475
rect 35548 10467 35564 10475
rect 35580 10467 35584 10475
rect 35588 10467 35600 10475
rect 35612 10467 35616 10475
rect 35620 10467 35624 10475
rect 35644 10467 35648 10475
rect 35652 10467 35656 10475
rect 35720 10467 35724 10475
rect 35728 10467 35740 10475
rect 35752 10467 35756 10475
rect 35760 10467 35764 10475
rect 35776 10467 35788 10475
rect 35792 10467 35796 10475
rect 35812 10467 35816 10475
rect 35820 10467 35832 10475
rect 35844 10467 35848 10475
rect 35852 10467 35856 10475
rect 35868 10467 35880 10475
rect 35884 10467 35888 10475
rect 35904 10467 35920 10475
rect 35936 10467 35952 10475
rect 35960 10467 35992 10475
rect 36000 10467 36016 10475
rect 36028 10467 36044 10475
rect 36052 10467 36084 10475
rect 36092 10467 36104 10475
rect 36120 10467 36136 10475
rect 36144 10467 36176 10475
rect 36184 10467 36196 10475
rect 36216 10467 36228 10475
rect 36240 10467 36244 10475
rect 36248 10467 36260 10475
rect 36280 10467 36292 10475
rect 36304 10467 36308 10475
rect 36312 10467 36324 10475
rect 36328 10467 36332 10475
rect 36344 10467 36356 10475
rect 36368 10467 36372 10475
rect 36376 10467 36388 10475
rect 36392 10467 36396 10475
rect 36460 10467 36464 10475
rect 36468 10467 36480 10475
rect 36484 10467 36488 10475
rect 36500 10467 36512 10475
rect 36624 10467 36636 10475
rect 36640 10467 36652 10475
rect 36656 10467 36668 10475
rect 36684 10467 36700 10475
rect 36708 10467 36740 10475
rect 36748 10467 36764 10475
rect 36772 10467 36796 10475
rect 36812 10467 36816 10475
rect 36820 10467 36832 10475
rect 36836 10467 36848 10475
rect 36852 10467 36856 10475
rect 36968 10467 36972 10475
rect 36976 10467 36980 10475
rect 36992 10467 37004 10475
rect 37008 10467 37012 10475
rect 37032 10467 37036 10475
rect 37040 10467 37044 10475
rect 37060 10467 37108 10475
rect 37124 10467 37128 10475
rect 37132 10467 37136 10475
rect 37156 10467 37160 10475
rect 37164 10467 37176 10475
rect 37188 10467 37192 10475
rect 37196 10467 37200 10475
rect 37220 10467 37224 10475
rect 37228 10467 37232 10475
rect 37296 10467 37300 10475
rect 37304 10467 37308 10475
rect 37328 10467 37332 10475
rect 37336 10467 37340 10475
rect 37352 10467 37364 10475
rect 37384 10467 37396 10475
rect 37404 10467 37436 10475
rect 37452 10467 37476 10475
rect 37484 10467 37500 10475
rect 37516 10467 37540 10475
rect 37548 10467 37564 10475
rect 37572 10467 37588 10475
rect 37600 10467 37608 10475
rect 37612 10467 37616 10475
rect 37632 10467 37656 10475
rect 37672 10467 37684 10475
rect 37688 10467 37692 10475
rect 37712 10467 37716 10475
rect 37720 10467 37732 10475
rect 37736 10467 37748 10475
rect 37752 10467 37756 10475
rect 37776 10467 37780 10475
rect 37784 10467 37796 10475
rect 37800 10467 37804 10475
rect 37816 10467 37828 10475
rect 37840 10467 37844 10475
rect 37848 10467 37852 10475
rect 37872 10467 37876 10475
rect 37880 10467 37884 10475
rect 37964 10467 37968 10475
rect 37972 10467 37984 10475
rect 37988 10467 37992 10475
rect 38040 10467 38044 10475
rect 38048 10467 38060 10475
rect 38064 10467 38076 10475
rect 38080 10467 38084 10475
rect 38132 10467 38136 10475
rect 38140 10467 38152 10475
rect 38156 10467 38168 10475
rect 38188 10467 38200 10475
rect 38212 10467 38216 10475
rect 38220 10467 38232 10475
rect 38252 10467 38264 10475
rect 38320 10467 38324 10475
rect 38328 10467 38332 10475
rect 38352 10467 38356 10475
rect 38360 10467 38364 10475
rect 38376 10467 38388 10475
rect 38404 10467 38420 10475
rect 38436 10467 38484 10475
rect 38500 10467 38516 10475
rect 38528 10467 38576 10475
rect 38592 10467 38596 10475
rect 38600 10467 38604 10475
rect 38624 10467 38628 10475
rect 38632 10467 38644 10475
rect 38656 10467 38660 10475
rect 38664 10467 38668 10475
rect 38688 10467 38692 10475
rect 38696 10467 38700 10475
rect 38780 10467 38784 10475
rect 38788 10467 38792 10475
rect 38888 10467 38892 10475
rect 38896 10467 38900 10475
rect 38912 10467 38924 10475
rect 38928 10467 38932 10475
rect 38952 10467 38956 10475
rect 38960 10467 38972 10475
rect 38976 10467 38988 10475
rect 38992 10467 38996 10475
rect 39044 10467 39048 10475
rect 39052 10467 39064 10475
rect 39068 10467 39080 10475
rect 39084 10467 39088 10475
rect 39184 10467 39188 10475
rect 39192 10467 39196 10475
rect 39216 10467 39220 10475
rect 39224 10467 39236 10475
rect 39240 10467 39252 10475
rect 39256 10467 39260 10475
rect 39276 10467 39292 10475
rect 39308 10467 39312 10475
rect 39316 10467 39328 10475
rect 39332 10467 39344 10475
rect 39348 10467 39352 10475
rect 39372 10467 39376 10475
rect 39380 10467 39392 10475
rect 39396 10467 39408 10475
rect 39412 10467 39416 10475
rect 39436 10467 39440 10475
rect 39444 10467 39448 10475
rect 39544 10467 39548 10475
rect 39552 10467 39564 10475
rect 39568 10467 39580 10475
rect 39584 10467 39588 10475
rect 39636 10467 39640 10475
rect 39644 10467 39656 10475
rect 39660 10467 39672 10475
rect 39676 10467 39680 10475
rect 39696 10467 39712 10475
rect 39728 10467 39744 10475
rect 39752 10467 39776 10475
rect 39792 10467 39816 10475
rect 39824 10467 39836 10475
rect 39844 10467 39868 10475
rect 39884 10467 39908 10475
rect 39916 10467 39928 10475
rect 39940 10467 39944 10475
rect 39948 10467 39960 10475
rect 39980 10467 39992 10475
rect 31680 10457 31688 10465
rect 32784 10437 32792 10445
rect 35344 10437 35352 10445
rect 36768 10437 36776 10445
rect 32752 10417 32760 10425
rect 38528 10397 38536 10405
rect 30016 10377 30024 10385
rect 30736 10377 30744 10385
rect 38784 10377 38792 10385
rect 39136 10377 39144 10385
rect 39200 10377 39208 10385
rect 39296 10377 39304 10385
rect 31152 10357 31160 10365
rect 32704 10357 32712 10365
rect 33888 10357 33896 10365
rect 34688 10357 34696 10365
rect 37152 10357 37160 10365
rect 30352 10337 30360 10345
rect 30752 10337 30760 10345
rect 36992 10337 37000 10345
rect 37104 10337 37112 10345
rect 37680 10337 37688 10345
rect 37840 10337 37848 10345
rect 37872 10337 37880 10345
rect 38352 10337 38360 10345
rect 38432 10337 38440 10345
rect 38736 10337 38744 10345
rect 38864 10337 38872 10345
rect 39216 10337 39224 10345
rect 29696 10317 29704 10325
rect 29904 10317 29912 10325
rect 30496 10317 30504 10325
rect 30672 10317 30680 10325
rect 31888 10317 31896 10325
rect 32704 10317 32712 10325
rect 32816 10317 32824 10325
rect 33376 10317 33384 10325
rect 33440 10317 33448 10325
rect 33856 10317 33864 10325
rect 34304 10317 34312 10325
rect 34368 10317 34376 10325
rect 34928 10317 34936 10325
rect 35936 10317 35944 10325
rect 36720 10317 36728 10325
rect 37488 10317 37496 10325
rect 29600 10297 29608 10305
rect 31328 10297 31336 10305
rect 31744 10297 31752 10305
rect 33152 10297 33160 10305
rect 33200 10297 33208 10305
rect 33216 10297 33224 10305
rect 34128 10297 34136 10305
rect 34192 10297 34200 10305
rect 37776 10297 37784 10305
rect 38912 10297 38920 10305
rect 39056 10297 39064 10305
rect 30880 10277 30888 10285
rect 33136 10277 33144 10285
rect 37936 10277 37944 10285
rect 39712 10277 39720 10285
rect 39728 10277 39736 10285
rect 29508 10267 29520 10275
rect 29540 10267 29552 10275
rect 29556 10267 29568 10275
rect 29588 10267 29600 10275
rect 29604 10267 29616 10275
rect 29620 10267 29632 10275
rect 29648 10267 29660 10275
rect 29680 10267 29692 10275
rect 29696 10267 29708 10275
rect 29712 10267 29724 10275
rect 29772 10267 29784 10275
rect 29788 10267 29800 10275
rect 29804 10267 29816 10275
rect 29836 10267 29848 10275
rect 29852 10267 29856 10275
rect 29868 10267 29880 10275
rect 29900 10267 29912 10275
rect 29916 10267 29920 10275
rect 29932 10267 29944 10275
rect 29952 10267 29976 10275
rect 29992 10267 30004 10275
rect 30008 10267 30012 10275
rect 30024 10267 30036 10275
rect 30044 10267 30068 10275
rect 30084 10267 30108 10275
rect 30116 10267 30132 10275
rect 30148 10267 30164 10275
rect 30180 10267 30184 10275
rect 30188 10267 30200 10275
rect 30204 10267 30216 10275
rect 30220 10267 30224 10275
rect 30240 10267 30244 10275
rect 30248 10267 30252 10275
rect 30272 10267 30276 10275
rect 30280 10267 30292 10275
rect 30296 10267 30308 10275
rect 30312 10267 30316 10275
rect 30336 10267 30340 10275
rect 30344 10267 30348 10275
rect 30412 10267 30416 10275
rect 30420 10267 30424 10275
rect 30444 10267 30448 10275
rect 30452 10267 30464 10275
rect 30468 10267 30480 10275
rect 30484 10267 30488 10275
rect 30508 10267 30512 10275
rect 30516 10267 30520 10275
rect 30536 10267 30552 10275
rect 30560 10267 30584 10275
rect 30600 10267 30624 10275
rect 30632 10267 30644 10275
rect 30656 10267 30660 10275
rect 30664 10267 30668 10275
rect 30680 10267 30692 10275
rect 30696 10267 30700 10275
rect 30716 10267 30720 10275
rect 30724 10267 30736 10275
rect 30756 10267 30768 10275
rect 30772 10267 30776 10275
rect 30864 10267 30876 10275
rect 30880 10267 30884 10275
rect 30904 10267 30908 10275
rect 30912 10267 30916 10275
rect 30928 10267 30940 10275
rect 30944 10267 30948 10275
rect 30968 10267 30972 10275
rect 30976 10267 30988 10275
rect 30992 10267 30996 10275
rect 31060 10267 31064 10275
rect 31068 10267 31080 10275
rect 31084 10267 31088 10275
rect 31100 10267 31112 10275
rect 31132 10267 31144 10275
rect 31160 10267 31184 10275
rect 31216 10267 31240 10275
rect 31256 10267 31260 10275
rect 31264 10267 31276 10275
rect 31288 10267 31292 10275
rect 31296 10267 31300 10275
rect 31412 10267 31416 10275
rect 31420 10267 31424 10275
rect 31520 10267 31524 10275
rect 31528 10267 31532 10275
rect 31612 10267 31616 10275
rect 31620 10267 31624 10275
rect 31636 10267 31648 10275
rect 31652 10267 31656 10275
rect 31672 10267 31688 10275
rect 31704 10267 31752 10275
rect 31768 10267 31784 10275
rect 31800 10267 31812 10275
rect 31824 10267 31828 10275
rect 31832 10267 31844 10275
rect 31988 10267 32000 10275
rect 32004 10267 32016 10275
rect 32020 10267 32032 10275
rect 32052 10267 32064 10275
rect 32080 10267 32104 10275
rect 32112 10267 32128 10275
rect 32144 10267 32160 10275
rect 32168 10267 32180 10275
rect 32184 10267 32196 10275
rect 32208 10267 32212 10275
rect 32216 10267 32220 10275
rect 32232 10267 32244 10275
rect 32248 10267 32252 10275
rect 32348 10267 32352 10275
rect 32356 10267 32360 10275
rect 32372 10267 32384 10275
rect 32388 10267 32400 10275
rect 32408 10267 32424 10275
rect 32440 10267 32488 10275
rect 32504 10267 32520 10275
rect 32536 10267 32548 10275
rect 32560 10267 32564 10275
rect 32568 10267 32580 10275
rect 32600 10267 32612 10275
rect 32616 10267 32620 10275
rect 32976 10267 32988 10275
rect 32992 10267 32996 10275
rect 33008 10267 33020 10275
rect 33040 10267 33052 10275
rect 33060 10267 33092 10275
rect 33100 10267 33116 10275
rect 33124 10267 33156 10275
rect 33164 10267 33180 10275
rect 33192 10267 33208 10275
rect 33216 10267 33248 10275
rect 33256 10267 33272 10275
rect 33288 10267 33300 10275
rect 33308 10267 33340 10275
rect 33348 10267 33364 10275
rect 33380 10267 33392 10275
rect 33404 10267 33408 10275
rect 33412 10267 33424 10275
rect 33444 10267 33456 10275
rect 33536 10267 33548 10275
rect 33660 10267 33672 10275
rect 33676 10267 33680 10275
rect 33692 10267 33704 10275
rect 33724 10267 33736 10275
rect 33744 10267 33776 10275
rect 33784 10267 33800 10275
rect 33808 10267 33832 10275
rect 33848 10267 33852 10275
rect 33856 10267 33868 10275
rect 33880 10267 33884 10275
rect 33888 10267 33892 10275
rect 33912 10267 33916 10275
rect 33920 10267 33924 10275
rect 34020 10267 34024 10275
rect 34028 10267 34032 10275
rect 34044 10267 34056 10275
rect 34060 10267 34064 10275
rect 34084 10267 34088 10275
rect 34092 10267 34096 10275
rect 34112 10267 34160 10275
rect 34176 10267 34200 10275
rect 34208 10267 34220 10275
rect 34232 10267 34236 10275
rect 34240 10267 34252 10275
rect 34256 10267 34260 10275
rect 34400 10267 34408 10275
rect 34412 10267 34424 10275
rect 34428 10267 34440 10275
rect 34616 10267 34628 10275
rect 34640 10267 34644 10275
rect 34648 10267 34660 10275
rect 34664 10267 34668 10275
rect 34680 10267 34692 10275
rect 34712 10267 34724 10275
rect 34740 10267 34764 10275
rect 34772 10267 34788 10275
rect 34796 10267 34808 10275
rect 34812 10267 34816 10275
rect 34836 10267 34840 10275
rect 34844 10267 34856 10275
rect 34864 10267 34880 10275
rect 34888 10267 34912 10275
rect 34928 10267 34932 10275
rect 34936 10267 34948 10275
rect 34960 10267 34964 10275
rect 34968 10267 34972 10275
rect 34992 10267 34996 10275
rect 35000 10267 35012 10275
rect 35024 10267 35028 10275
rect 35032 10267 35036 10275
rect 35048 10267 35060 10275
rect 35064 10267 35076 10275
rect 35084 10267 35100 10275
rect 35116 10267 35132 10275
rect 35140 10267 35164 10275
rect 35180 10267 35192 10275
rect 35212 10267 35224 10275
rect 35228 10267 35240 10275
rect 35244 10267 35256 10275
rect 35552 10267 35564 10275
rect 35568 10267 35572 10275
rect 35584 10267 35596 10275
rect 35616 10267 35628 10275
rect 35644 10267 35692 10275
rect 35708 10267 35724 10275
rect 35732 10267 35744 10275
rect 35748 10267 35760 10275
rect 35772 10267 35776 10275
rect 35780 10267 35784 10275
rect 35800 10267 35816 10275
rect 35824 10267 35836 10275
rect 35840 10267 35852 10275
rect 35864 10267 35868 10275
rect 35872 10267 35876 10275
rect 35896 10267 35900 10275
rect 35904 10267 35908 10275
rect 35928 10267 35932 10275
rect 35936 10267 35940 10275
rect 35960 10267 35964 10275
rect 35968 10267 35972 10275
rect 35984 10267 35996 10275
rect 36000 10267 36012 10275
rect 36020 10267 36036 10275
rect 36052 10267 36100 10275
rect 36112 10267 36128 10275
rect 36144 10267 36192 10275
rect 36208 10267 36224 10275
rect 36240 10267 36244 10275
rect 36248 10267 36260 10275
rect 36272 10267 36276 10275
rect 36280 10267 36284 10275
rect 36304 10267 36308 10275
rect 36312 10267 36316 10275
rect 36412 10267 36416 10275
rect 36420 10267 36424 10275
rect 36436 10267 36448 10275
rect 36452 10267 36456 10275
rect 36504 10267 36508 10275
rect 36512 10267 36516 10275
rect 36528 10267 36540 10275
rect 36544 10267 36548 10275
rect 36568 10267 36572 10275
rect 36576 10267 36580 10275
rect 36596 10267 36612 10275
rect 36620 10267 36652 10275
rect 36660 10267 36676 10275
rect 36692 10267 36704 10275
rect 36708 10267 36720 10275
rect 36724 10267 36736 10275
rect 36756 10267 36768 10275
rect 36772 10267 36776 10275
rect 36788 10267 36800 10275
rect 36820 10267 36832 10275
rect 36836 10267 36840 10275
rect 36852 10267 36864 10275
rect 36876 10267 36880 10275
rect 36884 10267 36896 10275
rect 36900 10267 36904 10275
rect 36968 10267 36972 10275
rect 36976 10267 36988 10275
rect 36992 10267 36996 10275
rect 37008 10267 37020 10275
rect 37060 10267 37064 10275
rect 37068 10267 37080 10275
rect 37084 10267 37088 10275
rect 37100 10267 37112 10275
rect 37192 10267 37204 10275
rect 37224 10267 37236 10275
rect 37240 10267 37252 10275
rect 37256 10267 37268 10275
rect 37284 10267 37300 10275
rect 37316 10267 37340 10275
rect 37348 10267 37364 10275
rect 37380 10267 37384 10275
rect 37388 10267 37392 10275
rect 37404 10267 37416 10275
rect 37420 10267 37432 10275
rect 37444 10267 37448 10275
rect 37452 10267 37456 10275
rect 37468 10267 37480 10275
rect 37484 10267 37488 10275
rect 37632 10267 37636 10275
rect 37640 10267 37644 10275
rect 37664 10267 37668 10275
rect 37672 10267 37684 10275
rect 37688 10267 37700 10275
rect 37876 10267 37888 10275
rect 37908 10267 37920 10275
rect 37924 10267 37928 10275
rect 37940 10267 37952 10275
rect 37964 10267 37968 10275
rect 37972 10267 37984 10275
rect 38000 10267 38012 10275
rect 38016 10267 38020 10275
rect 38032 10267 38044 10275
rect 38056 10267 38060 10275
rect 38064 10267 38076 10275
rect 38092 10267 38104 10275
rect 38108 10267 38112 10275
rect 38124 10267 38136 10275
rect 38148 10267 38152 10275
rect 38156 10267 38168 10275
rect 38188 10267 38200 10275
rect 38212 10267 38216 10275
rect 38220 10267 38232 10275
rect 38252 10267 38264 10275
rect 38268 10267 38272 10275
rect 38304 10267 38308 10275
rect 38312 10267 38324 10275
rect 38344 10267 38356 10275
rect 38360 10267 38364 10275
rect 38376 10267 38388 10275
rect 38408 10267 38420 10275
rect 38424 10267 38428 10275
rect 38440 10267 38452 10275
rect 38464 10267 38468 10275
rect 38472 10267 38484 10275
rect 38500 10267 38524 10275
rect 38532 10267 38544 10275
rect 38552 10267 38576 10275
rect 38592 10267 38616 10275
rect 38624 10267 38640 10275
rect 38656 10267 38672 10275
rect 38688 10267 38692 10275
rect 38696 10267 38708 10275
rect 38712 10267 38724 10275
rect 38728 10267 38732 10275
rect 38752 10267 38756 10275
rect 38760 10267 38772 10275
rect 38780 10267 38796 10275
rect 38804 10267 38828 10275
rect 38844 10267 38848 10275
rect 38852 10267 38864 10275
rect 38876 10267 38880 10275
rect 38884 10267 38888 10275
rect 38908 10267 38912 10275
rect 38916 10267 38920 10275
rect 38940 10267 38944 10275
rect 38948 10267 38952 10275
rect 38964 10267 38976 10275
rect 38980 10267 38984 10275
rect 39000 10267 39024 10275
rect 39032 10267 39048 10275
rect 39056 10267 39088 10275
rect 39096 10267 39108 10275
rect 39124 10267 39140 10275
rect 39148 10267 39180 10275
rect 39188 10267 39200 10275
rect 39220 10267 39232 10275
rect 39240 10267 39272 10275
rect 39280 10267 39292 10275
rect 39312 10267 39324 10275
rect 39328 10267 39340 10275
rect 39344 10267 39356 10275
rect 39376 10267 39388 10275
rect 39396 10267 39428 10275
rect 39436 10267 39452 10275
rect 39468 10267 39472 10275
rect 39476 10267 39480 10275
rect 39500 10267 39504 10275
rect 39508 10267 39520 10275
rect 39532 10267 39536 10275
rect 39540 10267 39544 10275
rect 39556 10267 39568 10275
rect 39572 10267 39576 10275
rect 39592 10267 39596 10275
rect 39600 10267 39612 10275
rect 39624 10267 39628 10275
rect 39632 10267 39636 10275
rect 39648 10267 39660 10275
rect 39664 10267 39668 10275
rect 39732 10267 39736 10275
rect 39740 10267 39744 10275
rect 39764 10267 39768 10275
rect 39772 10267 39776 10275
rect 39788 10267 39800 10275
rect 39804 10267 39816 10275
rect 39828 10267 39832 10275
rect 39836 10267 39840 10275
rect 39856 10267 39860 10275
rect 39864 10267 39868 10275
rect 39880 10267 39892 10275
rect 39896 10267 39908 10275
rect 39920 10267 39924 10275
rect 39928 10267 39932 10275
rect 39948 10267 39964 10275
rect 39972 10267 39996 10275
rect 30704 10257 30712 10265
rect 32256 10257 32264 10265
rect 29408 10237 29416 10245
rect 29808 10237 29816 10245
rect 31408 10237 31416 10245
rect 33120 10237 33128 10245
rect 35648 10237 35656 10245
rect 35936 10237 35944 10245
rect 29856 10217 29864 10225
rect 35024 10217 35032 10225
rect 35072 10217 35080 10225
rect 35184 10217 35192 10225
rect 36672 10217 36680 10225
rect 36832 10217 36840 10225
rect 37600 10217 37608 10225
rect 37792 10217 37800 10225
rect 37840 10217 37848 10225
rect 29376 10197 29384 10205
rect 29712 10197 29720 10205
rect 30080 10197 30088 10205
rect 31472 10197 31480 10205
rect 31696 10197 31704 10205
rect 31872 10197 31880 10205
rect 31936 10197 31944 10205
rect 32576 10197 32584 10205
rect 32880 10197 32888 10205
rect 32976 10197 32984 10205
rect 33136 10197 33144 10205
rect 33424 10197 33432 10205
rect 34240 10197 34248 10205
rect 34272 10197 34280 10205
rect 34336 10197 34344 10205
rect 34464 10197 34472 10205
rect 34528 10197 34536 10205
rect 34832 10197 34840 10205
rect 35168 10197 35176 10205
rect 35488 10197 35496 10205
rect 35584 10197 35592 10205
rect 35776 10197 35784 10205
rect 36176 10197 36184 10205
rect 36976 10197 36984 10205
rect 37248 10197 37256 10205
rect 37936 10197 37944 10205
rect 38848 10197 38856 10205
rect 39904 10197 39912 10205
rect 30896 10177 30904 10185
rect 30928 10177 30936 10185
rect 38000 10177 38008 10185
rect 29968 10157 29976 10165
rect 30320 10157 30328 10165
rect 30512 10157 30520 10165
rect 31216 10157 31224 10165
rect 31584 10157 31592 10165
rect 31760 10157 31768 10165
rect 32480 10157 32488 10165
rect 32496 10157 32504 10165
rect 32864 10157 32872 10165
rect 33344 10157 33352 10165
rect 33520 10157 33528 10165
rect 33616 10157 33624 10165
rect 33696 10157 33704 10165
rect 33984 10157 33992 10165
rect 34352 10157 34360 10165
rect 36288 10157 36296 10165
rect 36384 10157 36392 10165
rect 36480 10157 36488 10165
rect 36656 10157 36664 10165
rect 37200 10157 37208 10165
rect 37296 10157 37304 10165
rect 38640 10157 38648 10165
rect 39472 10157 39480 10165
rect 39648 10157 39656 10165
rect 30656 10117 30664 10125
rect 30800 10117 30808 10125
rect 33440 10117 33448 10125
rect 36960 10117 36968 10125
rect 37088 10117 37096 10125
rect 33152 10097 33160 10105
rect 34960 10097 34968 10105
rect 29500 10067 29504 10075
rect 29508 10067 29512 10075
rect 29608 10067 29612 10075
rect 29616 10067 29628 10075
rect 29772 10067 29784 10075
rect 29788 10067 29792 10075
rect 29804 10067 29816 10075
rect 29836 10067 29848 10075
rect 29852 10067 29856 10075
rect 29868 10067 29880 10075
rect 29892 10067 29896 10075
rect 29900 10067 29912 10075
rect 29916 10067 29920 10075
rect 29960 10067 29972 10075
rect 29984 10067 29988 10075
rect 29992 10067 30004 10075
rect 30008 10067 30012 10075
rect 30024 10067 30036 10075
rect 30052 10067 30064 10075
rect 30076 10067 30080 10075
rect 30084 10067 30096 10075
rect 30100 10067 30104 10075
rect 30168 10067 30172 10075
rect 30176 10067 30188 10075
rect 30192 10067 30196 10075
rect 30208 10067 30220 10075
rect 30236 10067 30252 10075
rect 30268 10067 30292 10075
rect 30300 10067 30316 10075
rect 30324 10067 30348 10075
rect 30364 10067 30368 10075
rect 30372 10067 30384 10075
rect 30416 10067 30428 10075
rect 30432 10067 30436 10075
rect 30456 10067 30460 10075
rect 30464 10067 30476 10075
rect 30484 10067 30500 10075
rect 30508 10067 30532 10075
rect 30548 10067 30552 10075
rect 30556 10067 30568 10075
rect 30576 10067 30592 10075
rect 30600 10067 30624 10075
rect 30640 10067 30644 10075
rect 30648 10067 30660 10075
rect 30680 10067 30692 10075
rect 30780 10067 30784 10075
rect 30788 10067 30792 10075
rect 30856 10067 30860 10075
rect 30864 10067 30868 10075
rect 30880 10067 30892 10075
rect 30912 10067 30924 10075
rect 30928 10067 30932 10075
rect 30944 10067 30956 10075
rect 30976 10067 30988 10075
rect 30992 10067 31004 10075
rect 31008 10067 31012 10075
rect 31032 10067 31036 10075
rect 31040 10067 31044 10075
rect 31060 10067 31064 10075
rect 31068 10067 31080 10075
rect 31084 10067 31088 10075
rect 31100 10067 31112 10075
rect 31124 10067 31128 10075
rect 31132 10067 31136 10075
rect 31152 10067 31168 10075
rect 31176 10067 31200 10075
rect 31216 10067 31232 10075
rect 31248 10067 31260 10075
rect 31264 10067 31276 10075
rect 31284 10067 31300 10075
rect 31316 10067 31320 10075
rect 31324 10067 31328 10075
rect 31340 10067 31352 10075
rect 31360 10067 31384 10075
rect 31400 10067 31424 10075
rect 31432 10067 31444 10075
rect 31456 10067 31460 10075
rect 31464 10067 31476 10075
rect 31492 10067 31516 10075
rect 31524 10067 31536 10075
rect 31548 10067 31552 10075
rect 31556 10067 31568 10075
rect 31584 10067 31608 10075
rect 31616 10067 31628 10075
rect 31640 10067 31644 10075
rect 31648 10067 31660 10075
rect 31664 10067 31668 10075
rect 31804 10067 31816 10075
rect 31820 10067 31832 10075
rect 31836 10067 31848 10075
rect 31864 10067 31880 10075
rect 31896 10067 31908 10075
rect 31912 10067 31924 10075
rect 31928 10067 31940 10075
rect 31960 10067 31972 10075
rect 31988 10067 32012 10075
rect 32020 10067 32036 10075
rect 32052 10067 32068 10075
rect 32076 10067 32088 10075
rect 32092 10067 32104 10075
rect 32112 10067 32128 10075
rect 32144 10067 32160 10075
rect 32168 10067 32180 10075
rect 32184 10067 32196 10075
rect 32208 10067 32212 10075
rect 32216 10067 32220 10075
rect 32236 10067 32252 10075
rect 32260 10067 32272 10075
rect 32276 10067 32288 10075
rect 32300 10067 32304 10075
rect 32308 10067 32312 10075
rect 32328 10067 32344 10075
rect 32352 10067 32364 10075
rect 32368 10067 32380 10075
rect 32392 10067 32396 10075
rect 32400 10067 32404 10075
rect 32420 10067 32424 10075
rect 32428 10067 32432 10075
rect 32444 10067 32456 10075
rect 32460 10067 32472 10075
rect 32484 10067 32488 10075
rect 32492 10067 32496 10075
rect 32512 10067 32528 10075
rect 32536 10067 32548 10075
rect 32552 10067 32564 10075
rect 32576 10067 32580 10075
rect 32584 10067 32588 10075
rect 32604 10067 32620 10075
rect 32628 10067 32640 10075
rect 32644 10067 32656 10075
rect 32668 10067 32672 10075
rect 32676 10067 32680 10075
rect 32696 10067 32712 10075
rect 32720 10067 32744 10075
rect 32760 10067 32776 10075
rect 32792 10067 32804 10075
rect 32808 10067 32820 10075
rect 32824 10067 32836 10075
rect 32852 10067 32868 10075
rect 32876 10067 32908 10075
rect 32916 10067 32932 10075
rect 32948 10067 32964 10075
rect 32980 10067 32996 10075
rect 33012 10067 33028 10075
rect 33036 10067 33068 10075
rect 33076 10067 33092 10075
rect 33108 10067 33120 10075
rect 33124 10067 33136 10075
rect 33140 10067 33152 10075
rect 33172 10067 33184 10075
rect 33200 10067 33212 10075
rect 33216 10067 33228 10075
rect 33232 10067 33236 10075
rect 33256 10067 33260 10075
rect 33264 10067 33276 10075
rect 33284 10067 33300 10075
rect 33308 10067 33320 10075
rect 33324 10067 33328 10075
rect 33348 10067 33352 10075
rect 33356 10067 33368 10075
rect 33376 10067 33392 10075
rect 33400 10067 33424 10075
rect 33440 10067 33444 10075
rect 33448 10067 33460 10075
rect 33468 10067 33484 10075
rect 33492 10067 33516 10075
rect 33532 10067 33548 10075
rect 33564 10067 33576 10075
rect 33588 10067 33592 10075
rect 33596 10067 33608 10075
rect 33612 10067 33616 10075
rect 33628 10067 33640 10075
rect 33844 10067 33856 10075
rect 33860 10067 33864 10075
rect 33876 10067 33888 10075
rect 33908 10067 33920 10075
rect 33928 10067 33960 10075
rect 33968 10067 33984 10075
rect 33992 10067 34016 10075
rect 34032 10067 34036 10075
rect 34040 10067 34052 10075
rect 34064 10067 34068 10075
rect 34072 10067 34076 10075
rect 34096 10067 34100 10075
rect 34104 10067 34108 10075
rect 34204 10067 34208 10075
rect 34212 10067 34224 10075
rect 34228 10067 34240 10075
rect 34244 10067 34248 10075
rect 34264 10067 34288 10075
rect 34296 10067 34312 10075
rect 34320 10067 34344 10075
rect 34360 10067 34376 10075
rect 34392 10067 34400 10075
rect 34416 10067 34420 10075
rect 34424 10067 34436 10075
rect 34440 10067 34444 10075
rect 34456 10067 34468 10075
rect 34488 10067 34500 10075
rect 34504 10067 34508 10075
rect 34520 10067 34532 10075
rect 34552 10067 34564 10075
rect 34572 10067 34604 10075
rect 34612 10067 34624 10075
rect 34644 10067 34656 10075
rect 34668 10067 34672 10075
rect 34676 10067 34688 10075
rect 34708 10067 34720 10075
rect 34800 10067 34812 10075
rect 34832 10067 34844 10075
rect 34848 10067 34852 10075
rect 34864 10067 34876 10075
rect 34896 10067 34908 10075
rect 34916 10067 34948 10075
rect 34956 10067 34972 10075
rect 34988 10067 35000 10075
rect 35004 10067 35016 10075
rect 35020 10067 35032 10075
rect 35052 10067 35064 10075
rect 35068 10067 35072 10075
rect 35176 10067 35188 10075
rect 35192 10067 35196 10075
rect 35208 10067 35220 10075
rect 35228 10067 35252 10075
rect 35268 10067 35316 10075
rect 35332 10067 35348 10075
rect 35360 10067 35408 10075
rect 35424 10067 35440 10075
rect 35452 10067 35500 10075
rect 35516 10067 35540 10075
rect 35548 10067 35560 10075
rect 35572 10067 35576 10075
rect 35580 10067 35592 10075
rect 35612 10067 35624 10075
rect 35736 10067 35748 10075
rect 35752 10067 35764 10075
rect 35768 10067 35780 10075
rect 35800 10067 35812 10075
rect 35828 10067 35840 10075
rect 35844 10067 35856 10075
rect 35860 10067 35872 10075
rect 36008 10067 36012 10075
rect 36016 10067 36028 10075
rect 36032 10067 36036 10075
rect 36048 10067 36060 10075
rect 36072 10067 36076 10075
rect 36080 10067 36092 10075
rect 36236 10067 36248 10075
rect 36252 10067 36256 10075
rect 36328 10067 36340 10075
rect 36344 10067 36348 10075
rect 36360 10067 36372 10075
rect 36392 10067 36404 10075
rect 36420 10067 36468 10075
rect 36484 10067 36500 10075
rect 36508 10067 36520 10075
rect 36524 10067 36536 10075
rect 36548 10067 36552 10075
rect 36556 10067 36560 10075
rect 36576 10067 36592 10075
rect 36600 10067 36612 10075
rect 36616 10067 36628 10075
rect 36640 10067 36644 10075
rect 36648 10067 36652 10075
rect 36672 10067 36676 10075
rect 36680 10067 36684 10075
rect 36796 10067 36800 10075
rect 36804 10067 36808 10075
rect 36828 10067 36832 10075
rect 36836 10067 36840 10075
rect 36852 10067 36864 10075
rect 36868 10067 36880 10075
rect 36892 10067 36896 10075
rect 36900 10067 36904 10075
rect 36920 10067 36924 10075
rect 36928 10067 36932 10075
rect 36944 10067 36956 10075
rect 36960 10067 36972 10075
rect 36984 10067 36988 10075
rect 36992 10067 36996 10075
rect 37008 10067 37020 10075
rect 37024 10067 37028 10075
rect 37124 10067 37128 10075
rect 37132 10067 37144 10075
rect 37148 10067 37160 10075
rect 37164 10067 37168 10075
rect 37184 10067 37208 10075
rect 37216 10067 37232 10075
rect 37240 10067 37272 10075
rect 37280 10067 37292 10075
rect 37312 10067 37324 10075
rect 37336 10067 37340 10075
rect 37344 10067 37356 10075
rect 37720 10067 37732 10075
rect 37744 10067 37748 10075
rect 37752 10067 37764 10075
rect 37768 10067 37772 10075
rect 37784 10067 37796 10075
rect 37808 10067 37812 10075
rect 37816 10067 37828 10075
rect 37832 10067 37836 10075
rect 37848 10067 37860 10075
rect 37876 10067 37888 10075
rect 37900 10067 37904 10075
rect 37908 10067 37920 10075
rect 37924 10067 37928 10075
rect 37992 10067 37996 10075
rect 38000 10067 38012 10075
rect 38016 10067 38020 10075
rect 38032 10067 38044 10075
rect 38056 10067 38060 10075
rect 38064 10067 38076 10075
rect 38092 10067 38116 10075
rect 38124 10067 38140 10075
rect 38156 10067 38172 10075
rect 38188 10067 38204 10075
rect 38212 10067 38236 10075
rect 38252 10067 38300 10075
rect 38316 10067 38320 10075
rect 38324 10067 38328 10075
rect 38340 10067 38352 10075
rect 38356 10067 38368 10075
rect 38376 10067 38392 10075
rect 38408 10067 38456 10075
rect 38472 10067 38484 10075
rect 38500 10067 38548 10075
rect 38560 10067 38576 10075
rect 38592 10067 38640 10075
rect 38656 10067 38672 10075
rect 38684 10067 38732 10075
rect 38748 10067 38760 10075
rect 38764 10067 38768 10075
rect 38780 10067 38792 10075
rect 38804 10067 38808 10075
rect 38812 10067 38824 10075
rect 38840 10067 38888 10075
rect 38904 10067 38920 10075
rect 38936 10067 38952 10075
rect 38968 10067 38984 10075
rect 39000 10067 39048 10075
rect 39064 10067 39076 10075
rect 39080 10067 39084 10075
rect 39096 10067 39108 10075
rect 39116 10067 39140 10075
rect 39156 10067 39200 10075
rect 39220 10067 39236 10075
rect 39252 10067 39256 10075
rect 39260 10067 39272 10075
rect 39284 10067 39288 10075
rect 39292 10067 39296 10075
rect 39316 10067 39320 10075
rect 39324 10067 39336 10075
rect 39340 10067 39352 10075
rect 39356 10067 39360 10075
rect 39376 10067 39392 10075
rect 39408 10067 39412 10075
rect 39416 10067 39428 10075
rect 39432 10067 39444 10075
rect 39448 10067 39452 10075
rect 39500 10067 39504 10075
rect 39508 10067 39520 10075
rect 39524 10067 39536 10075
rect 39540 10067 39544 10075
rect 39564 10067 39568 10075
rect 39572 10067 39576 10075
rect 39672 10067 39676 10075
rect 39680 10067 39692 10075
rect 39696 10067 39708 10075
rect 39712 10067 39716 10075
rect 39732 10067 39756 10075
rect 39764 10067 39780 10075
rect 39788 10067 39812 10075
rect 39828 10067 39844 10075
rect 39860 10067 39872 10075
rect 39884 10067 39888 10075
rect 39892 10067 39904 10075
rect 39908 10067 39912 10075
rect 39924 10067 39936 10075
rect 39952 10067 39964 10075
rect 39976 10067 39980 10075
rect 39984 10067 39996 10075
rect 33984 10057 33992 10065
rect 35312 10057 35320 10065
rect 29584 10037 29592 10045
rect 31616 10037 31624 10045
rect 37088 10037 37096 10045
rect 30976 10017 30984 10025
rect 31344 10017 31352 10025
rect 34512 10017 34520 10025
rect 34656 10017 34664 10025
rect 34672 10017 34680 10025
rect 34704 10017 34712 10025
rect 31072 9997 31080 10005
rect 32080 9997 32088 10005
rect 39344 9997 39352 10005
rect 29536 9977 29544 9985
rect 29808 9977 29816 9985
rect 30448 9977 30456 9985
rect 31600 9977 31608 9985
rect 31632 9977 31640 9985
rect 31856 9977 31864 9985
rect 32128 9977 32136 9985
rect 32304 9977 32312 9985
rect 32736 9977 32744 9985
rect 34224 9977 34232 9985
rect 34272 9977 34280 9985
rect 34544 9977 34552 9985
rect 36544 9977 36552 9985
rect 36816 9977 36824 9985
rect 37248 9977 37256 9985
rect 37952 9977 37960 9985
rect 38496 9977 38504 9985
rect 38656 9977 38664 9985
rect 38784 9977 38792 9985
rect 39472 9977 39480 9985
rect 33808 9957 33816 9965
rect 33856 9957 33864 9965
rect 37648 9957 37656 9965
rect 37968 9957 37976 9965
rect 29968 9937 29976 9945
rect 30528 9937 30536 9945
rect 31296 9937 31304 9945
rect 31328 9937 31336 9945
rect 31392 9937 31400 9945
rect 31520 9937 31528 9945
rect 32192 9937 32200 9945
rect 32464 9937 32472 9945
rect 34528 9937 34536 9945
rect 29824 9917 29832 9925
rect 30640 9917 30648 9925
rect 31968 9917 31976 9925
rect 32032 9917 32040 9925
rect 33248 9917 33256 9925
rect 33344 9917 33352 9925
rect 36720 9917 36728 9925
rect 37152 9917 37160 9925
rect 37488 9917 37496 9925
rect 37600 9917 37608 9925
rect 37664 9917 37672 9925
rect 38256 9917 38264 9925
rect 39008 9917 39016 9925
rect 29680 9897 29688 9905
rect 30752 9897 30760 9905
rect 30944 9897 30952 9905
rect 32816 9897 32824 9905
rect 33568 9897 33576 9905
rect 33840 9897 33848 9905
rect 34064 9897 34072 9905
rect 34576 9897 34584 9905
rect 34928 9897 34936 9905
rect 35520 9897 35528 9905
rect 35600 9897 35608 9905
rect 34352 9877 34360 9885
rect 29452 9867 29456 9875
rect 29460 9867 29464 9875
rect 29476 9867 29488 9875
rect 29496 9867 29512 9875
rect 29528 9867 29532 9875
rect 29536 9867 29540 9875
rect 29552 9867 29564 9875
rect 29572 9867 29596 9875
rect 29612 9867 29624 9875
rect 29628 9867 29632 9875
rect 29652 9867 29656 9875
rect 29660 9867 29672 9875
rect 29680 9867 29696 9875
rect 29704 9867 29720 9875
rect 29728 9867 29752 9875
rect 29768 9867 29784 9875
rect 29800 9867 29816 9875
rect 29832 9867 29856 9875
rect 29872 9867 29896 9875
rect 29904 9867 29916 9875
rect 29924 9867 29948 9875
rect 29964 9867 29976 9875
rect 29980 9867 29984 9875
rect 29996 9867 30008 9875
rect 30020 9867 30024 9875
rect 30028 9867 30040 9875
rect 30056 9867 30080 9875
rect 30088 9867 30100 9875
rect 30108 9867 30132 9875
rect 30148 9867 30196 9875
rect 30212 9867 30228 9875
rect 30244 9867 30260 9875
rect 30276 9867 30292 9875
rect 30308 9867 30356 9875
rect 30372 9867 30388 9875
rect 30400 9867 30408 9875
rect 30412 9867 30424 9875
rect 30432 9867 30448 9875
rect 30464 9867 30480 9875
rect 30488 9867 30500 9875
rect 30504 9867 30516 9875
rect 30524 9867 30540 9875
rect 30556 9867 30572 9875
rect 30580 9867 30592 9875
rect 30596 9867 30608 9875
rect 30616 9867 30632 9875
rect 30648 9867 30664 9875
rect 30672 9867 30696 9875
rect 30712 9867 30728 9875
rect 30736 9867 30768 9875
rect 30776 9867 30792 9875
rect 30808 9867 30812 9875
rect 30816 9867 30820 9875
rect 30840 9867 30844 9875
rect 30848 9867 30860 9875
rect 30880 9867 30892 9875
rect 30896 9867 30900 9875
rect 30912 9867 30924 9875
rect 30940 9867 30956 9875
rect 30972 9867 31012 9875
rect 31028 9867 31040 9875
rect 31056 9867 31088 9875
rect 31104 9867 31128 9875
rect 31144 9867 31160 9875
rect 31176 9867 31192 9875
rect 31208 9867 31232 9875
rect 31248 9867 31260 9875
rect 31264 9867 31268 9875
rect 31284 9867 31308 9875
rect 31324 9867 31336 9875
rect 31340 9867 31344 9875
rect 31360 9867 31384 9875
rect 31400 9867 31412 9875
rect 31416 9867 31420 9875
rect 31432 9867 31444 9875
rect 31456 9867 31460 9875
rect 31464 9867 31468 9875
rect 31484 9867 31500 9875
rect 31508 9867 31520 9875
rect 31524 9867 31536 9875
rect 31584 9867 31596 9875
rect 31600 9867 31612 9875
rect 31616 9867 31628 9875
rect 31648 9867 31660 9875
rect 31664 9867 31668 9875
rect 31680 9867 31692 9875
rect 31712 9867 31724 9875
rect 31744 9867 31756 9875
rect 31768 9867 31772 9875
rect 31776 9867 31788 9875
rect 31808 9867 31820 9875
rect 31824 9867 31836 9875
rect 31840 9867 31852 9875
rect 31900 9867 31912 9875
rect 31916 9867 31928 9875
rect 31932 9867 31944 9875
rect 32212 9867 32224 9875
rect 32304 9867 32316 9875
rect 32428 9867 32440 9875
rect 32444 9867 32448 9875
rect 32460 9867 32472 9875
rect 32492 9867 32504 9875
rect 32512 9867 32544 9875
rect 32552 9867 32564 9875
rect 32584 9867 32596 9875
rect 32604 9867 32636 9875
rect 32644 9867 32660 9875
rect 32676 9867 32692 9875
rect 32708 9867 32712 9875
rect 32716 9867 32728 9875
rect 32740 9867 32744 9875
rect 32748 9867 32752 9875
rect 32764 9867 32776 9875
rect 32780 9867 32784 9875
rect 32928 9867 32932 9875
rect 32936 9867 32940 9875
rect 32960 9867 32964 9875
rect 32968 9867 32972 9875
rect 32984 9867 32996 9875
rect 33000 9867 33004 9875
rect 33024 9867 33028 9875
rect 33032 9867 33044 9875
rect 33048 9867 33060 9875
rect 33064 9867 33068 9875
rect 33088 9867 33092 9875
rect 33096 9867 33100 9875
rect 33116 9867 33120 9875
rect 33124 9867 33136 9875
rect 33140 9867 33152 9875
rect 33156 9867 33160 9875
rect 33180 9867 33184 9875
rect 33188 9867 33192 9875
rect 33304 9867 33308 9875
rect 33312 9867 33324 9875
rect 33344 9867 33356 9875
rect 33360 9867 33372 9875
rect 33376 9867 33388 9875
rect 33408 9867 33420 9875
rect 33436 9867 33460 9875
rect 33468 9867 33484 9875
rect 33500 9867 33516 9875
rect 33524 9867 33548 9875
rect 33564 9867 33580 9875
rect 33588 9867 33620 9875
rect 33628 9867 33644 9875
rect 33660 9867 33672 9875
rect 33676 9867 33688 9875
rect 33692 9867 33704 9875
rect 33752 9867 33764 9875
rect 33768 9867 33780 9875
rect 33784 9867 33796 9875
rect 33908 9867 33920 9875
rect 33932 9867 33936 9875
rect 33940 9867 33952 9875
rect 33956 9867 33960 9875
rect 33972 9867 33984 9875
rect 33996 9867 34000 9875
rect 34004 9867 34016 9875
rect 34032 9867 34056 9875
rect 34064 9867 34080 9875
rect 34096 9867 34112 9875
rect 34128 9867 34132 9875
rect 34136 9867 34148 9875
rect 34152 9867 34164 9875
rect 34168 9867 34172 9875
rect 34268 9867 34272 9875
rect 34276 9867 34288 9875
rect 34300 9867 34304 9875
rect 34308 9867 34312 9875
rect 34324 9867 34336 9875
rect 34340 9867 34344 9875
rect 34364 9867 34368 9875
rect 34372 9867 34376 9875
rect 34416 9867 34448 9875
rect 34456 9867 34468 9875
rect 34488 9867 34500 9875
rect 34504 9867 34516 9875
rect 34520 9867 34532 9875
rect 34580 9867 34592 9875
rect 34596 9867 34608 9875
rect 34612 9867 34624 9875
rect 34644 9867 34656 9875
rect 34760 9867 34764 9875
rect 34768 9867 34780 9875
rect 34784 9867 34788 9875
rect 34800 9867 34812 9875
rect 34828 9867 34844 9875
rect 34860 9867 34884 9875
rect 34892 9867 34908 9875
rect 34916 9867 34928 9875
rect 34932 9867 34936 9875
rect 34956 9867 34960 9875
rect 34964 9867 34976 9875
rect 34984 9867 35000 9875
rect 35008 9867 35020 9875
rect 35024 9867 35028 9875
rect 35048 9867 35052 9875
rect 35056 9867 35068 9875
rect 35076 9867 35092 9875
rect 35100 9867 35112 9875
rect 35116 9867 35120 9875
rect 35140 9867 35144 9875
rect 35148 9867 35160 9875
rect 35168 9867 35184 9875
rect 35200 9867 35216 9875
rect 35232 9867 35244 9875
rect 35264 9867 35276 9875
rect 35288 9867 35292 9875
rect 35296 9867 35308 9875
rect 35312 9867 35316 9875
rect 35328 9867 35340 9875
rect 35452 9867 35464 9875
rect 35468 9867 35480 9875
rect 35484 9867 35496 9875
rect 35640 9867 35652 9875
rect 35656 9867 35660 9875
rect 35672 9867 35684 9875
rect 35692 9867 35716 9875
rect 35732 9867 35780 9875
rect 35796 9867 35812 9875
rect 35828 9867 35840 9875
rect 35852 9867 35856 9875
rect 35860 9867 35872 9875
rect 35944 9867 35948 9875
rect 35952 9867 35964 9875
rect 35984 9867 35996 9875
rect 36000 9867 36004 9875
rect 36076 9867 36088 9875
rect 36092 9867 36096 9875
rect 36108 9867 36120 9875
rect 36140 9867 36152 9875
rect 36156 9867 36160 9875
rect 36172 9867 36184 9875
rect 36192 9867 36216 9875
rect 36232 9867 36256 9875
rect 36264 9867 36276 9875
rect 36288 9867 36292 9875
rect 36296 9867 36308 9875
rect 36324 9867 36348 9875
rect 36356 9867 36372 9875
rect 36388 9867 36412 9875
rect 36420 9867 36436 9875
rect 36444 9867 36476 9875
rect 36484 9867 36500 9875
rect 36508 9867 36540 9875
rect 36548 9867 36564 9875
rect 36580 9867 36592 9875
rect 36600 9867 36632 9875
rect 36640 9867 36656 9875
rect 36672 9867 36676 9875
rect 36680 9867 36684 9875
rect 36704 9867 36708 9875
rect 36712 9867 36724 9875
rect 36736 9867 36740 9875
rect 36744 9867 36748 9875
rect 36760 9867 36772 9875
rect 36776 9867 36780 9875
rect 36796 9867 36800 9875
rect 36804 9867 36816 9875
rect 36828 9867 36832 9875
rect 36836 9867 36840 9875
rect 36852 9867 36864 9875
rect 36868 9867 36872 9875
rect 36892 9867 36896 9875
rect 36900 9867 36904 9875
rect 36920 9867 36936 9875
rect 36944 9867 36976 9875
rect 36984 9867 37000 9875
rect 37008 9867 37020 9875
rect 37024 9867 37028 9875
rect 37048 9867 37052 9875
rect 37056 9867 37068 9875
rect 37072 9867 37084 9875
rect 37088 9867 37092 9875
rect 37112 9867 37116 9875
rect 37120 9867 37124 9875
rect 37136 9867 37148 9875
rect 37152 9867 37156 9875
rect 37176 9867 37180 9875
rect 37184 9867 37188 9875
rect 37200 9867 37212 9875
rect 37216 9867 37228 9875
rect 37240 9867 37244 9875
rect 37248 9867 37252 9875
rect 37380 9867 37384 9875
rect 37388 9867 37392 9875
rect 37404 9867 37416 9875
rect 37420 9867 37432 9875
rect 37444 9867 37448 9875
rect 37452 9867 37456 9875
rect 37472 9867 37488 9875
rect 37496 9867 37508 9875
rect 37512 9867 37524 9875
rect 37532 9867 37548 9875
rect 37564 9867 37612 9875
rect 37628 9867 37640 9875
rect 37660 9867 37672 9875
rect 37684 9867 37688 9875
rect 37692 9867 37704 9875
rect 37848 9867 37860 9875
rect 37864 9867 37868 9875
rect 37940 9867 37952 9875
rect 37972 9867 37984 9875
rect 37988 9867 37992 9875
rect 38004 9867 38016 9875
rect 38028 9867 38032 9875
rect 38036 9867 38048 9875
rect 38052 9867 38056 9875
rect 38068 9867 38080 9875
rect 38092 9867 38096 9875
rect 38100 9867 38112 9875
rect 38132 9867 38144 9875
rect 38216 9867 38220 9875
rect 38224 9867 38236 9875
rect 38256 9867 38268 9875
rect 38272 9867 38284 9875
rect 38288 9867 38300 9875
rect 38316 9867 38332 9875
rect 38340 9867 38372 9875
rect 38380 9867 38392 9875
rect 38412 9867 38424 9875
rect 38436 9867 38440 9875
rect 38444 9867 38456 9875
rect 38692 9867 38704 9875
rect 38708 9867 38712 9875
rect 38724 9867 38736 9875
rect 38752 9867 38768 9875
rect 38776 9867 38808 9875
rect 38816 9867 38832 9875
rect 38840 9867 38872 9875
rect 38880 9867 38896 9875
rect 38912 9867 38928 9875
rect 38944 9867 38960 9875
rect 38976 9867 38992 9875
rect 39000 9867 39032 9875
rect 39040 9867 39052 9875
rect 39068 9867 39084 9875
rect 39092 9867 39124 9875
rect 39132 9867 39144 9875
rect 39164 9867 39176 9875
rect 39180 9867 39192 9875
rect 39196 9867 39208 9875
rect 39228 9867 39240 9875
rect 39344 9867 39348 9875
rect 39352 9867 39364 9875
rect 39368 9867 39372 9875
rect 39412 9867 39424 9875
rect 39436 9867 39440 9875
rect 39444 9867 39456 9875
rect 39460 9867 39464 9875
rect 39476 9867 39488 9875
rect 39504 9867 39516 9875
rect 39528 9867 39532 9875
rect 39536 9867 39548 9875
rect 39552 9867 39556 9875
rect 39568 9867 39580 9875
rect 39596 9867 39612 9875
rect 39628 9867 39652 9875
rect 39660 9867 39676 9875
rect 39684 9867 39696 9875
rect 39700 9867 39704 9875
rect 39724 9867 39728 9875
rect 39732 9867 39744 9875
rect 39748 9867 39760 9875
rect 39764 9867 39768 9875
rect 39788 9867 39792 9875
rect 39796 9867 39808 9875
rect 39820 9867 39824 9875
rect 39828 9867 39832 9875
rect 39852 9867 39856 9875
rect 39860 9867 39864 9875
rect 39928 9867 39932 9875
rect 39936 9867 39940 9875
rect 31456 9857 31464 9865
rect 33584 9857 33592 9865
rect 34688 9857 34696 9865
rect 34976 9857 34984 9865
rect 39664 9857 39672 9865
rect 29744 9837 29752 9845
rect 29904 9837 29912 9845
rect 30400 9837 30408 9845
rect 30480 9837 30488 9845
rect 30992 9837 31000 9845
rect 31008 9837 31016 9845
rect 31072 9837 31080 9845
rect 31520 9837 31528 9845
rect 31808 9837 31816 9845
rect 32048 9837 32056 9845
rect 32224 9837 32232 9845
rect 32272 9837 32280 9845
rect 32832 9837 32840 9845
rect 33664 9837 33672 9845
rect 33680 9837 33688 9845
rect 33776 9837 33784 9845
rect 34160 9837 34168 9845
rect 34512 9837 34520 9845
rect 34880 9837 34888 9845
rect 36160 9837 36168 9845
rect 37488 9837 37496 9845
rect 38672 9837 38680 9845
rect 39104 9837 39112 9845
rect 29344 9817 29352 9825
rect 29536 9817 29544 9825
rect 30112 9817 30120 9825
rect 31216 9817 31224 9825
rect 31296 9817 31304 9825
rect 31648 9817 31656 9825
rect 32080 9817 32088 9825
rect 34224 9817 34232 9825
rect 36480 9817 36488 9825
rect 37472 9817 37480 9825
rect 38480 9817 38488 9825
rect 38608 9817 38616 9825
rect 38800 9817 38808 9825
rect 39360 9817 39368 9825
rect 39728 9817 39736 9825
rect 39776 9817 39784 9825
rect 39888 9817 39896 9825
rect 39920 9817 39928 9825
rect 39952 9817 39960 9825
rect 29536 9797 29544 9805
rect 29744 9797 29752 9805
rect 30224 9797 30232 9805
rect 31056 9797 31064 9805
rect 32608 9797 32616 9805
rect 33600 9797 33608 9805
rect 33840 9797 33848 9805
rect 33968 9797 33976 9805
rect 34304 9797 34312 9805
rect 34672 9797 34680 9805
rect 35040 9797 35048 9805
rect 36272 9797 36280 9805
rect 36640 9797 36648 9805
rect 36864 9797 36872 9805
rect 37040 9797 37048 9805
rect 37328 9797 37336 9805
rect 37568 9797 37576 9805
rect 39536 9797 39544 9805
rect 39712 9797 39720 9805
rect 30112 9777 30120 9785
rect 30224 9777 30232 9785
rect 30560 9777 30568 9785
rect 30720 9777 30728 9785
rect 30816 9777 30824 9785
rect 31152 9777 31160 9785
rect 31584 9777 31592 9785
rect 36880 9777 36888 9785
rect 37056 9777 37064 9785
rect 29632 9757 29640 9765
rect 30640 9757 30648 9765
rect 31040 9757 31048 9765
rect 31472 9757 31480 9765
rect 31824 9757 31832 9765
rect 31968 9757 31976 9765
rect 32944 9757 32952 9765
rect 33920 9757 33928 9765
rect 34368 9757 34376 9765
rect 34560 9757 34568 9765
rect 35968 9757 35976 9765
rect 37024 9757 37032 9765
rect 37280 9757 37288 9765
rect 39696 9757 39704 9765
rect 37664 9737 37672 9745
rect 30544 9717 30552 9725
rect 32864 9717 32872 9725
rect 38128 9717 38136 9725
rect 38240 9717 38248 9725
rect 29404 9667 29408 9675
rect 29412 9667 29416 9675
rect 29428 9667 29440 9675
rect 29496 9667 29500 9675
rect 29504 9667 29508 9675
rect 29528 9667 29532 9675
rect 29536 9667 29540 9675
rect 29552 9667 29564 9675
rect 29572 9667 29588 9675
rect 29604 9667 29620 9675
rect 29628 9667 29640 9675
rect 29652 9667 29656 9675
rect 29660 9667 29664 9675
rect 29680 9667 29696 9675
rect 29704 9667 29716 9675
rect 29728 9667 29732 9675
rect 29736 9667 29740 9675
rect 29760 9667 29764 9675
rect 29768 9667 29780 9675
rect 29792 9667 29796 9675
rect 29800 9667 29804 9675
rect 29824 9667 29828 9675
rect 29832 9667 29836 9675
rect 29900 9667 29904 9675
rect 29908 9667 29920 9675
rect 29924 9667 29936 9675
rect 29940 9667 29944 9675
rect 29960 9667 29976 9675
rect 29992 9667 29996 9675
rect 30000 9667 30012 9675
rect 30016 9667 30028 9675
rect 30032 9667 30036 9675
rect 30056 9667 30060 9675
rect 30064 9667 30076 9675
rect 30084 9667 30100 9675
rect 30108 9667 30132 9675
rect 30148 9667 30164 9675
rect 30172 9667 30196 9675
rect 30212 9667 30236 9675
rect 30244 9667 30260 9675
rect 30276 9667 30280 9675
rect 30284 9667 30288 9675
rect 30308 9667 30312 9675
rect 30316 9667 30328 9675
rect 30332 9667 30344 9675
rect 30348 9667 30352 9675
rect 30432 9667 30436 9675
rect 30440 9667 30444 9675
rect 30524 9667 30528 9675
rect 30532 9667 30536 9675
rect 30616 9667 30620 9675
rect 30624 9667 30628 9675
rect 30648 9667 30652 9675
rect 30656 9667 30660 9675
rect 30756 9667 30760 9675
rect 30764 9667 30768 9675
rect 30780 9667 30792 9675
rect 30796 9667 30800 9675
rect 30820 9667 30824 9675
rect 30828 9667 30832 9675
rect 30844 9667 30856 9675
rect 30860 9667 30864 9675
rect 30884 9667 30888 9675
rect 30892 9667 30904 9675
rect 30916 9667 30920 9675
rect 30924 9667 30928 9675
rect 31024 9667 31028 9675
rect 31032 9667 31036 9675
rect 31140 9667 31152 9675
rect 31172 9667 31184 9675
rect 31188 9667 31192 9675
rect 31204 9667 31216 9675
rect 31224 9667 31240 9675
rect 31256 9667 31260 9675
rect 31264 9667 31268 9675
rect 31280 9667 31292 9675
rect 31296 9667 31308 9675
rect 31396 9667 31400 9675
rect 31404 9667 31408 9675
rect 31428 9667 31432 9675
rect 31436 9667 31448 9675
rect 31452 9667 31464 9675
rect 31484 9667 31496 9675
rect 31504 9667 31536 9675
rect 31552 9667 31564 9675
rect 31580 9667 31628 9675
rect 31644 9667 31648 9675
rect 31652 9667 31656 9675
rect 31676 9667 31680 9675
rect 31684 9667 31696 9675
rect 31708 9667 31712 9675
rect 31716 9667 31720 9675
rect 31740 9667 31744 9675
rect 31748 9667 31752 9675
rect 31816 9667 31820 9675
rect 31824 9667 31836 9675
rect 31848 9667 31852 9675
rect 31856 9667 31860 9675
rect 31908 9667 31912 9675
rect 31916 9667 31928 9675
rect 31940 9667 31944 9675
rect 31948 9667 31952 9675
rect 32000 9667 32004 9675
rect 32008 9667 32020 9675
rect 32032 9667 32036 9675
rect 32040 9667 32044 9675
rect 32056 9667 32068 9675
rect 32072 9667 32084 9675
rect 32092 9667 32108 9675
rect 32124 9667 32128 9675
rect 32132 9667 32136 9675
rect 32148 9667 32160 9675
rect 32164 9667 32176 9675
rect 32188 9667 32192 9675
rect 32196 9667 32200 9675
rect 32296 9667 32300 9675
rect 32304 9667 32316 9675
rect 32328 9667 32332 9675
rect 32336 9667 32340 9675
rect 32352 9667 32364 9675
rect 32368 9667 32372 9675
rect 32548 9667 32552 9675
rect 32556 9667 32568 9675
rect 32580 9667 32584 9675
rect 32588 9667 32592 9675
rect 32720 9667 32724 9675
rect 32728 9667 32732 9675
rect 32744 9667 32756 9675
rect 32760 9667 32772 9675
rect 32780 9667 32796 9675
rect 32812 9667 32860 9675
rect 32876 9667 32900 9675
rect 32908 9667 32920 9675
rect 32928 9667 32952 9675
rect 32968 9667 32992 9675
rect 33000 9667 33016 9675
rect 33032 9667 33056 9675
rect 33064 9667 33080 9675
rect 33088 9667 33112 9675
rect 33128 9667 33132 9675
rect 33136 9667 33148 9675
rect 33156 9667 33172 9675
rect 33180 9667 33204 9675
rect 33220 9667 33236 9675
rect 33244 9667 33268 9675
rect 33284 9667 33296 9675
rect 33300 9667 33304 9675
rect 33316 9667 33328 9675
rect 33340 9667 33344 9675
rect 33348 9667 33360 9675
rect 33364 9667 33368 9675
rect 33380 9667 33392 9675
rect 33404 9667 33408 9675
rect 33412 9667 33424 9675
rect 33444 9667 33456 9675
rect 33528 9667 33532 9675
rect 33536 9667 33548 9675
rect 33568 9667 33580 9675
rect 33584 9667 33596 9675
rect 33600 9667 33612 9675
rect 33632 9667 33644 9675
rect 33724 9667 33736 9675
rect 33748 9667 33752 9675
rect 33756 9667 33768 9675
rect 33772 9667 33776 9675
rect 33788 9667 33800 9675
rect 33808 9667 33832 9675
rect 33848 9667 33896 9675
rect 33912 9667 33916 9675
rect 33920 9667 33924 9675
rect 33936 9667 33948 9675
rect 33952 9667 33964 9675
rect 33976 9667 33980 9675
rect 33984 9667 33988 9675
rect 34000 9667 34012 9675
rect 34016 9667 34020 9675
rect 34116 9667 34120 9675
rect 34124 9667 34128 9675
rect 34140 9667 34152 9675
rect 34156 9667 34168 9675
rect 34176 9667 34192 9675
rect 34208 9667 34224 9675
rect 34232 9667 34256 9675
rect 34272 9667 34284 9675
rect 34304 9667 34316 9675
rect 34320 9667 34332 9675
rect 34336 9667 34348 9675
rect 34368 9667 34380 9675
rect 34384 9667 34388 9675
rect 34452 9667 34456 9675
rect 34460 9667 34472 9675
rect 34492 9667 34504 9675
rect 34508 9667 34512 9675
rect 34524 9667 34536 9675
rect 34552 9667 34568 9675
rect 34584 9667 34632 9675
rect 34648 9667 34660 9675
rect 34676 9667 34716 9675
rect 34732 9667 34748 9675
rect 34764 9667 34776 9675
rect 34788 9667 34792 9675
rect 34796 9667 34808 9675
rect 34912 9667 34916 9675
rect 34920 9667 34924 9675
rect 34944 9667 34948 9675
rect 34952 9667 34956 9675
rect 34968 9667 34980 9675
rect 34984 9667 34996 9675
rect 35004 9667 35020 9675
rect 35036 9667 35040 9675
rect 35044 9667 35048 9675
rect 35060 9667 35072 9675
rect 35076 9667 35088 9675
rect 35104 9667 35120 9675
rect 35136 9667 35160 9675
rect 35168 9667 35184 9675
rect 35200 9667 35216 9675
rect 35224 9667 35240 9675
rect 35256 9667 35260 9675
rect 35264 9667 35268 9675
rect 35288 9667 35292 9675
rect 35296 9667 35308 9675
rect 35312 9667 35316 9675
rect 35328 9667 35340 9675
rect 35396 9667 35400 9675
rect 35404 9667 35408 9675
rect 35428 9667 35432 9675
rect 35436 9667 35440 9675
rect 35452 9667 35464 9675
rect 35468 9667 35480 9675
rect 35492 9667 35496 9675
rect 35500 9667 35504 9675
rect 35632 9667 35636 9675
rect 35640 9667 35644 9675
rect 35692 9667 35696 9675
rect 35700 9667 35712 9675
rect 35724 9667 35728 9675
rect 35732 9667 35736 9675
rect 35748 9667 35760 9675
rect 35764 9667 35768 9675
rect 35788 9667 35792 9675
rect 35796 9667 35800 9675
rect 35820 9667 35824 9675
rect 35828 9667 35832 9675
rect 35852 9667 35856 9675
rect 35860 9667 35872 9675
rect 35884 9667 35888 9675
rect 35892 9667 35896 9675
rect 35944 9667 35948 9675
rect 35952 9667 35964 9675
rect 35976 9667 35980 9675
rect 35984 9667 35988 9675
rect 36068 9667 36072 9675
rect 36076 9667 36080 9675
rect 36192 9667 36196 9675
rect 36200 9667 36204 9675
rect 36224 9667 36228 9675
rect 36232 9667 36244 9675
rect 36248 9667 36252 9675
rect 36264 9667 36276 9675
rect 36288 9667 36292 9675
rect 36296 9667 36308 9675
rect 36324 9667 36348 9675
rect 36356 9667 36368 9675
rect 36380 9667 36384 9675
rect 36388 9667 36400 9675
rect 36404 9667 36408 9675
rect 36420 9667 36432 9675
rect 36452 9667 36464 9675
rect 36468 9667 36472 9675
rect 36484 9667 36496 9675
rect 36516 9667 36528 9675
rect 36532 9667 36544 9675
rect 36548 9667 36560 9675
rect 36580 9667 36592 9675
rect 36600 9667 36632 9675
rect 36640 9667 36652 9675
rect 36668 9667 36684 9675
rect 36692 9667 36724 9675
rect 36732 9667 36748 9675
rect 36764 9667 36776 9675
rect 36784 9667 36816 9675
rect 36824 9667 36840 9675
rect 36848 9667 36872 9675
rect 36888 9667 36900 9675
rect 36920 9667 36932 9675
rect 36944 9667 36948 9675
rect 36952 9667 36964 9675
rect 36968 9667 36972 9675
rect 37012 9667 37024 9675
rect 37036 9667 37040 9675
rect 37044 9667 37056 9675
rect 37060 9667 37064 9675
rect 37076 9667 37088 9675
rect 37264 9667 37276 9675
rect 37288 9667 37292 9675
rect 37296 9667 37308 9675
rect 37312 9667 37316 9675
rect 37328 9667 37340 9675
rect 37352 9667 37356 9675
rect 37360 9667 37364 9675
rect 37380 9667 37396 9675
rect 37404 9667 37428 9675
rect 37444 9667 37460 9675
rect 37476 9667 37488 9675
rect 37492 9667 37504 9675
rect 37508 9667 37520 9675
rect 37624 9667 37628 9675
rect 37632 9667 37636 9675
rect 37656 9667 37660 9675
rect 37664 9667 37668 9675
rect 37680 9667 37692 9675
rect 37696 9667 37708 9675
rect 37716 9667 37732 9675
rect 37748 9667 37780 9675
rect 37788 9667 37804 9675
rect 37820 9667 37832 9675
rect 37840 9667 37856 9675
rect 37864 9667 37888 9675
rect 37904 9667 37920 9675
rect 37936 9667 37952 9675
rect 37968 9667 37992 9675
rect 38008 9667 38020 9675
rect 38024 9667 38028 9675
rect 38040 9667 38052 9675
rect 38064 9667 38068 9675
rect 38072 9667 38084 9675
rect 38088 9667 38092 9675
rect 38104 9667 38116 9675
rect 38128 9667 38132 9675
rect 38136 9667 38140 9675
rect 38156 9667 38188 9675
rect 38196 9667 38212 9675
rect 38224 9667 38240 9675
rect 38248 9667 38264 9675
rect 38272 9667 38284 9675
rect 38288 9667 38292 9675
rect 38308 9667 38332 9675
rect 38348 9667 38372 9675
rect 38380 9667 38392 9675
rect 38404 9667 38408 9675
rect 38412 9667 38416 9675
rect 38504 9667 38516 9675
rect 38528 9667 38532 9675
rect 38536 9667 38548 9675
rect 38552 9667 38556 9675
rect 38844 9667 38848 9675
rect 38852 9667 38864 9675
rect 38884 9667 38896 9675
rect 38900 9667 38904 9675
rect 38916 9667 38928 9675
rect 38948 9667 38960 9675
rect 38976 9667 39024 9675
rect 39040 9667 39052 9675
rect 39068 9667 39116 9675
rect 39132 9667 39144 9675
rect 39164 9667 39176 9675
rect 39188 9667 39192 9675
rect 39196 9667 39208 9675
rect 39228 9667 39240 9675
rect 39244 9667 39248 9675
rect 39280 9667 39284 9675
rect 39288 9667 39300 9675
rect 39320 9667 39332 9675
rect 39336 9667 39340 9675
rect 39496 9667 39500 9675
rect 39504 9667 39508 9675
rect 39528 9667 39532 9675
rect 39536 9667 39540 9675
rect 39552 9667 39564 9675
rect 39568 9667 39580 9675
rect 39588 9667 39604 9675
rect 39620 9667 39636 9675
rect 39644 9667 39668 9675
rect 39684 9667 39696 9675
rect 39716 9667 39728 9675
rect 39732 9667 39744 9675
rect 39748 9667 39760 9675
rect 39780 9667 39792 9675
rect 39796 9667 39808 9675
rect 39812 9667 39824 9675
rect 39844 9667 39856 9675
rect 39936 9667 39948 9675
rect 39960 9667 39964 9675
rect 39968 9667 39980 9675
rect 39984 9667 39988 9675
rect 29712 9637 29720 9645
rect 33168 9637 33176 9645
rect 33184 9637 33192 9645
rect 33328 9637 33336 9645
rect 29552 9617 29560 9625
rect 29808 9617 29816 9625
rect 31920 9617 31928 9625
rect 32880 9617 32888 9625
rect 36192 9617 36200 9625
rect 36464 9617 36472 9625
rect 38112 9617 38120 9625
rect 38480 9617 38488 9625
rect 34992 9597 35000 9605
rect 39264 9597 39272 9605
rect 29664 9577 29672 9585
rect 29952 9577 29960 9585
rect 30992 9577 31000 9585
rect 31056 9577 31064 9585
rect 31648 9577 31656 9585
rect 31728 9577 31736 9585
rect 34672 9577 34680 9585
rect 35328 9577 35336 9585
rect 35600 9577 35608 9585
rect 36272 9577 36280 9585
rect 36720 9577 36728 9585
rect 36960 9577 36968 9585
rect 37648 9577 37656 9585
rect 37664 9577 37672 9585
rect 37840 9577 37848 9585
rect 38192 9577 38200 9585
rect 39024 9577 39032 9585
rect 39424 9577 39432 9585
rect 39872 9577 39880 9585
rect 35552 9557 35560 9565
rect 30480 9537 30488 9545
rect 30576 9537 30584 9545
rect 31344 9537 31352 9545
rect 31664 9537 31672 9545
rect 31936 9537 31944 9545
rect 31952 9537 31960 9545
rect 32128 9537 32136 9545
rect 33424 9537 33432 9545
rect 35296 9537 35304 9545
rect 36128 9537 36136 9545
rect 36240 9537 36248 9545
rect 36272 9537 36280 9545
rect 37184 9537 37192 9545
rect 37920 9537 37928 9545
rect 38048 9537 38056 9545
rect 38176 9537 38184 9545
rect 38464 9537 38472 9545
rect 30224 9517 30232 9525
rect 30752 9517 30760 9525
rect 30864 9517 30872 9525
rect 30912 9517 30920 9525
rect 33056 9517 33064 9525
rect 33760 9517 33768 9525
rect 34224 9517 34232 9525
rect 34304 9517 34312 9525
rect 34528 9517 34536 9525
rect 34560 9517 34568 9525
rect 34720 9517 34728 9525
rect 35360 9517 35368 9525
rect 30784 9497 30792 9505
rect 31184 9497 31192 9505
rect 31568 9497 31576 9505
rect 32512 9497 32520 9505
rect 36144 9497 36152 9505
rect 37328 9497 37336 9505
rect 37344 9497 37352 9505
rect 37360 9497 37368 9505
rect 37440 9497 37448 9505
rect 38480 9497 38488 9505
rect 38768 9497 38776 9505
rect 39136 9497 39144 9505
rect 39776 9497 39784 9505
rect 39856 9497 39864 9505
rect 33392 9477 33400 9485
rect 29404 9467 29408 9475
rect 29412 9467 29416 9475
rect 29428 9467 29440 9475
rect 29496 9467 29500 9475
rect 29504 9467 29508 9475
rect 29528 9467 29532 9475
rect 29536 9467 29540 9475
rect 29552 9467 29564 9475
rect 29576 9467 29580 9475
rect 29584 9467 29588 9475
rect 29604 9467 29620 9475
rect 29628 9467 29640 9475
rect 29652 9467 29656 9475
rect 29660 9467 29664 9475
rect 29684 9467 29688 9475
rect 29692 9467 29696 9475
rect 29980 9467 29984 9475
rect 29988 9467 29992 9475
rect 30004 9467 30016 9475
rect 30020 9467 30032 9475
rect 30052 9467 30064 9475
rect 30068 9467 30080 9475
rect 30084 9467 30096 9475
rect 30116 9467 30128 9475
rect 30140 9467 30144 9475
rect 30148 9467 30160 9475
rect 30364 9467 30376 9475
rect 30400 9467 30408 9475
rect 30412 9467 30416 9475
rect 30428 9467 30440 9475
rect 30456 9467 30472 9475
rect 30480 9467 30512 9475
rect 30520 9467 30536 9475
rect 30548 9467 30564 9475
rect 30572 9467 30604 9475
rect 30612 9467 30628 9475
rect 30644 9467 30660 9475
rect 30676 9467 30680 9475
rect 30684 9467 30696 9475
rect 30708 9467 30712 9475
rect 30716 9467 30720 9475
rect 30732 9467 30744 9475
rect 30748 9467 30752 9475
rect 30768 9467 30772 9475
rect 30776 9467 30788 9475
rect 30800 9467 30804 9475
rect 30808 9467 30812 9475
rect 30824 9467 30836 9475
rect 30840 9467 30852 9475
rect 30864 9467 30868 9475
rect 30872 9467 30876 9475
rect 30892 9467 30908 9475
rect 30916 9467 30940 9475
rect 30956 9467 30972 9475
rect 30988 9467 31012 9475
rect 31020 9467 31036 9475
rect 31052 9467 31056 9475
rect 31060 9467 31064 9475
rect 31076 9467 31088 9475
rect 31092 9467 31104 9475
rect 31116 9467 31120 9475
rect 31124 9467 31128 9475
rect 31176 9467 31180 9475
rect 31184 9467 31196 9475
rect 31208 9467 31212 9475
rect 31216 9467 31220 9475
rect 31300 9467 31304 9475
rect 31308 9467 31312 9475
rect 31324 9467 31336 9475
rect 31340 9467 31344 9475
rect 31360 9467 31376 9475
rect 31392 9467 31408 9475
rect 31416 9467 31448 9475
rect 31456 9467 31472 9475
rect 31480 9467 31512 9475
rect 31520 9467 31536 9475
rect 31552 9467 31564 9475
rect 31572 9467 31604 9475
rect 31612 9467 31628 9475
rect 31636 9467 31648 9475
rect 31652 9467 31656 9475
rect 31676 9467 31680 9475
rect 31684 9467 31696 9475
rect 31708 9467 31712 9475
rect 31716 9467 31720 9475
rect 31740 9467 31744 9475
rect 31748 9467 31752 9475
rect 31816 9467 31820 9475
rect 31824 9467 31828 9475
rect 31848 9467 31852 9475
rect 31856 9467 31860 9475
rect 31872 9467 31884 9475
rect 31888 9467 31892 9475
rect 31908 9467 31924 9475
rect 31940 9467 31988 9475
rect 32004 9467 32016 9475
rect 32020 9467 32024 9475
rect 32036 9467 32048 9475
rect 32056 9467 32080 9475
rect 32096 9467 32108 9475
rect 32112 9467 32116 9475
rect 32128 9467 32140 9475
rect 32152 9467 32156 9475
rect 32160 9467 32172 9475
rect 32188 9467 32212 9475
rect 32220 9467 32236 9475
rect 32252 9467 32256 9475
rect 32260 9467 32264 9475
rect 32284 9467 32288 9475
rect 32292 9467 32304 9475
rect 32308 9467 32320 9475
rect 32324 9467 32328 9475
rect 32348 9467 32352 9475
rect 32356 9467 32368 9475
rect 32376 9467 32392 9475
rect 32400 9467 32424 9475
rect 32440 9467 32444 9475
rect 32448 9467 32460 9475
rect 32472 9467 32476 9475
rect 32480 9467 32484 9475
rect 32504 9467 32508 9475
rect 32512 9467 32524 9475
rect 32536 9467 32540 9475
rect 32544 9467 32548 9475
rect 32560 9467 32572 9475
rect 32576 9467 32580 9475
rect 32596 9467 32600 9475
rect 32604 9467 32616 9475
rect 32628 9467 32632 9475
rect 32636 9467 32640 9475
rect 32652 9467 32664 9475
rect 32668 9467 32672 9475
rect 32692 9467 32696 9475
rect 32700 9467 32704 9475
rect 32720 9467 32736 9475
rect 32744 9467 32776 9475
rect 32784 9467 32796 9475
rect 32816 9467 32828 9475
rect 32832 9467 32844 9475
rect 32848 9467 32860 9475
rect 32880 9467 32892 9475
rect 32908 9467 32920 9475
rect 32924 9467 32936 9475
rect 32940 9467 32952 9475
rect 32972 9467 32984 9475
rect 33000 9467 33024 9475
rect 33032 9467 33048 9475
rect 33064 9467 33068 9475
rect 33072 9467 33076 9475
rect 33088 9467 33100 9475
rect 33104 9467 33116 9475
rect 33128 9467 33132 9475
rect 33136 9467 33140 9475
rect 33156 9467 33172 9475
rect 33180 9467 33204 9475
rect 33220 9467 33236 9475
rect 33244 9467 33276 9475
rect 33284 9467 33296 9475
rect 33316 9467 33328 9475
rect 33332 9467 33344 9475
rect 33348 9467 33360 9475
rect 33380 9467 33392 9475
rect 33400 9467 33432 9475
rect 33440 9467 33456 9475
rect 33472 9467 33484 9475
rect 33496 9467 33500 9475
rect 33504 9467 33516 9475
rect 33660 9467 33672 9475
rect 33676 9467 33680 9475
rect 33692 9467 33704 9475
rect 33720 9467 33736 9475
rect 33744 9467 33776 9475
rect 33784 9467 33800 9475
rect 33808 9467 33820 9475
rect 33824 9467 33828 9475
rect 33848 9467 33852 9475
rect 33856 9467 33868 9475
rect 33872 9467 33884 9475
rect 33888 9467 33892 9475
rect 33912 9467 33916 9475
rect 33920 9467 33932 9475
rect 33936 9467 33948 9475
rect 33952 9467 33956 9475
rect 33976 9467 33980 9475
rect 33984 9467 33988 9475
rect 34052 9467 34056 9475
rect 34060 9467 34064 9475
rect 34084 9467 34088 9475
rect 34092 9467 34096 9475
rect 34108 9467 34120 9475
rect 34124 9467 34128 9475
rect 34144 9467 34168 9475
rect 34176 9467 34192 9475
rect 34200 9467 34224 9475
rect 34240 9467 34252 9475
rect 34272 9467 34284 9475
rect 34296 9467 34300 9475
rect 34304 9467 34316 9475
rect 34320 9467 34324 9475
rect 34452 9467 34456 9475
rect 34460 9467 34472 9475
rect 34476 9467 34480 9475
rect 34492 9467 34504 9475
rect 34520 9467 34536 9475
rect 34552 9467 34576 9475
rect 34592 9467 34604 9475
rect 34608 9467 34612 9475
rect 34624 9467 34636 9475
rect 34644 9467 34660 9475
rect 34676 9467 34692 9475
rect 34700 9467 34712 9475
rect 34724 9467 34728 9475
rect 34732 9467 34736 9475
rect 34756 9467 34760 9475
rect 34764 9467 34768 9475
rect 34848 9467 34852 9475
rect 34856 9467 34860 9475
rect 34872 9467 34884 9475
rect 34904 9467 34916 9475
rect 34932 9467 34956 9475
rect 34972 9467 34984 9475
rect 34988 9467 34992 9475
rect 35004 9467 35016 9475
rect 35024 9467 35040 9475
rect 35056 9467 35060 9475
rect 35064 9467 35068 9475
rect 35080 9467 35092 9475
rect 35104 9467 35108 9475
rect 35112 9467 35116 9475
rect 35136 9467 35140 9475
rect 35144 9467 35148 9475
rect 35244 9467 35248 9475
rect 35252 9467 35256 9475
rect 35276 9467 35280 9475
rect 35284 9467 35288 9475
rect 35300 9467 35312 9475
rect 35324 9467 35328 9475
rect 35332 9467 35336 9475
rect 35352 9467 35356 9475
rect 35360 9467 35364 9475
rect 35376 9467 35388 9475
rect 35396 9467 35420 9475
rect 35436 9467 35448 9475
rect 35452 9467 35456 9475
rect 35468 9467 35480 9475
rect 35492 9467 35496 9475
rect 35500 9467 35512 9475
rect 35532 9467 35544 9475
rect 35748 9467 35760 9475
rect 35764 9467 35768 9475
rect 35780 9467 35792 9475
rect 35808 9467 35824 9475
rect 35840 9467 35888 9475
rect 35904 9467 35916 9475
rect 35936 9467 35948 9475
rect 35960 9467 35964 9475
rect 35968 9467 35980 9475
rect 36084 9467 36088 9475
rect 36092 9467 36104 9475
rect 36124 9467 36136 9475
rect 36140 9467 36144 9475
rect 36240 9467 36244 9475
rect 36248 9467 36252 9475
rect 36264 9467 36276 9475
rect 36280 9467 36292 9475
rect 36304 9467 36308 9475
rect 36312 9467 36316 9475
rect 36332 9467 36348 9475
rect 36356 9467 36368 9475
rect 36372 9467 36384 9475
rect 36396 9467 36400 9475
rect 36404 9467 36408 9475
rect 36424 9467 36440 9475
rect 36448 9467 36472 9475
rect 36488 9467 36504 9475
rect 36520 9467 36532 9475
rect 36536 9467 36548 9475
rect 36552 9467 36564 9475
rect 36584 9467 36596 9475
rect 36600 9467 36604 9475
rect 36616 9467 36628 9475
rect 36644 9467 36660 9475
rect 36676 9467 36724 9475
rect 36740 9467 36756 9475
rect 36768 9467 36816 9475
rect 36832 9467 36856 9475
rect 36864 9467 36880 9475
rect 36896 9467 36900 9475
rect 36904 9467 36908 9475
rect 36928 9467 36932 9475
rect 36936 9467 36948 9475
rect 36952 9467 36964 9475
rect 36968 9467 36972 9475
rect 37020 9467 37024 9475
rect 37028 9467 37040 9475
rect 37044 9467 37056 9475
rect 37060 9467 37064 9475
rect 37084 9467 37088 9475
rect 37092 9467 37096 9475
rect 37112 9467 37116 9475
rect 37120 9467 37132 9475
rect 37136 9467 37148 9475
rect 37152 9467 37156 9475
rect 37176 9467 37180 9475
rect 37184 9467 37188 9475
rect 37204 9467 37220 9475
rect 37228 9467 37252 9475
rect 37268 9467 37292 9475
rect 37300 9467 37316 9475
rect 37332 9467 37356 9475
rect 37372 9467 37396 9475
rect 37404 9467 37420 9475
rect 37436 9467 37440 9475
rect 37444 9467 37448 9475
rect 37468 9467 37472 9475
rect 37476 9467 37488 9475
rect 37492 9467 37496 9475
rect 37616 9467 37628 9475
rect 37632 9467 37636 9475
rect 37652 9467 37668 9475
rect 37684 9467 37724 9475
rect 37740 9467 37744 9475
rect 37748 9467 37752 9475
rect 37764 9467 37776 9475
rect 37788 9467 37792 9475
rect 37796 9467 37800 9475
rect 37816 9467 37820 9475
rect 37824 9467 37828 9475
rect 37840 9467 37852 9475
rect 37864 9467 37868 9475
rect 37872 9467 37876 9475
rect 37896 9467 37900 9475
rect 37904 9467 37908 9475
rect 37964 9467 37976 9475
rect 37988 9467 37992 9475
rect 37996 9467 38000 9475
rect 38224 9467 38228 9475
rect 38232 9467 38236 9475
rect 38248 9467 38260 9475
rect 38276 9467 38292 9475
rect 38308 9467 38340 9475
rect 38356 9467 38372 9475
rect 38380 9467 38392 9475
rect 38404 9467 38408 9475
rect 38412 9467 38416 9475
rect 38504 9467 38516 9475
rect 38528 9467 38532 9475
rect 38536 9467 38540 9475
rect 38660 9467 38672 9475
rect 38676 9467 38680 9475
rect 38696 9467 38712 9475
rect 38728 9467 38768 9475
rect 38784 9467 38800 9475
rect 38808 9467 38820 9475
rect 38824 9467 38836 9475
rect 38844 9467 38860 9475
rect 38876 9467 38892 9475
rect 38900 9467 38912 9475
rect 38916 9467 38928 9475
rect 38940 9467 38944 9475
rect 38948 9467 38952 9475
rect 38968 9467 38984 9475
rect 38992 9467 39016 9475
rect 39032 9467 39048 9475
rect 39064 9467 39076 9475
rect 39080 9467 39092 9475
rect 39096 9467 39108 9475
rect 39124 9467 39140 9475
rect 39156 9467 39180 9475
rect 39188 9467 39200 9475
rect 39220 9467 39224 9475
rect 39228 9467 39232 9475
rect 39244 9467 39256 9475
rect 39260 9467 39272 9475
rect 39280 9467 39296 9475
rect 39312 9467 39316 9475
rect 39320 9467 39324 9475
rect 39336 9467 39348 9475
rect 39352 9467 39364 9475
rect 39376 9467 39380 9475
rect 39384 9467 39388 9475
rect 39404 9467 39444 9475
rect 39460 9467 39476 9475
rect 39484 9467 39500 9475
rect 39516 9467 39520 9475
rect 39524 9467 39528 9475
rect 39548 9467 39552 9475
rect 39556 9467 39568 9475
rect 39572 9467 39576 9475
rect 39656 9467 39660 9475
rect 39664 9467 39668 9475
rect 39688 9467 39692 9475
rect 39696 9467 39700 9475
rect 39712 9467 39724 9475
rect 39728 9467 39740 9475
rect 39748 9467 39764 9475
rect 39780 9467 39828 9475
rect 39844 9467 39856 9475
rect 39876 9467 39888 9475
rect 39900 9467 39904 9475
rect 39908 9467 39920 9475
rect 39992 9467 39996 9475
rect 34512 9457 34520 9465
rect 30640 9437 30648 9445
rect 33328 9437 33336 9445
rect 34944 9437 34952 9445
rect 35424 9437 35432 9445
rect 36448 9437 36456 9445
rect 37136 9437 37144 9445
rect 38032 9437 38040 9445
rect 38096 9437 38104 9445
rect 38480 9437 38488 9445
rect 38656 9437 38664 9445
rect 38800 9437 38808 9445
rect 39152 9437 39160 9445
rect 39280 9437 39288 9445
rect 39632 9437 39640 9445
rect 39808 9437 39816 9445
rect 29360 9417 29368 9425
rect 29376 9417 29384 9425
rect 29680 9417 29688 9425
rect 30080 9417 30088 9425
rect 30400 9417 30408 9425
rect 30608 9417 30616 9425
rect 30624 9417 30632 9425
rect 30832 9417 30840 9425
rect 31088 9417 31096 9425
rect 31632 9417 31640 9425
rect 31872 9417 31880 9425
rect 31968 9417 31976 9425
rect 32000 9417 32008 9425
rect 32464 9417 32472 9425
rect 32704 9417 32712 9425
rect 32768 9417 32776 9425
rect 35232 9417 35240 9425
rect 35280 9417 35288 9425
rect 35952 9417 35960 9425
rect 36000 9417 36008 9425
rect 37344 9417 37352 9425
rect 37744 9417 37752 9425
rect 39264 9417 39272 9425
rect 39376 9417 39384 9425
rect 39424 9417 39432 9425
rect 39984 9417 39992 9425
rect 29408 9397 29416 9405
rect 31248 9397 31256 9405
rect 32096 9397 32104 9405
rect 32272 9397 32280 9405
rect 33168 9397 33176 9405
rect 33696 9397 33704 9405
rect 33936 9397 33944 9405
rect 34176 9397 34184 9405
rect 36192 9397 36200 9405
rect 36448 9397 36456 9405
rect 37456 9397 37464 9405
rect 37696 9397 37704 9405
rect 37760 9397 37768 9405
rect 37840 9397 37848 9405
rect 37856 9397 37864 9405
rect 38128 9397 38136 9405
rect 38288 9397 38296 9405
rect 39024 9397 39032 9405
rect 39472 9397 39480 9405
rect 39616 9397 39624 9405
rect 30848 9377 30856 9385
rect 31392 9377 31400 9385
rect 31712 9377 31720 9385
rect 32640 9377 32648 9385
rect 32688 9377 32696 9385
rect 33184 9377 33192 9385
rect 35936 9377 35944 9385
rect 37040 9377 37048 9385
rect 38560 9377 38568 9385
rect 39008 9377 39016 9385
rect 29808 9357 29816 9365
rect 31200 9357 31208 9365
rect 31264 9357 31272 9365
rect 32960 9357 32968 9365
rect 33824 9357 33832 9365
rect 34256 9357 34264 9365
rect 36736 9357 36744 9365
rect 37088 9357 37096 9365
rect 37168 9357 37176 9365
rect 37440 9357 37448 9365
rect 38128 9357 38136 9365
rect 38256 9357 38264 9365
rect 38592 9357 38600 9365
rect 38624 9357 38632 9365
rect 38864 9357 38872 9365
rect 39136 9357 39144 9365
rect 39936 9357 39944 9365
rect 30864 9337 30872 9345
rect 32880 9337 32888 9345
rect 34576 9337 34584 9345
rect 32720 9297 32728 9305
rect 29452 9267 29456 9275
rect 29460 9267 29472 9275
rect 29476 9267 29480 9275
rect 29496 9267 29500 9275
rect 29504 9267 29508 9275
rect 29528 9267 29532 9275
rect 29536 9267 29548 9275
rect 29552 9267 29556 9275
rect 29576 9267 29580 9275
rect 29584 9267 29596 9275
rect 29604 9267 29620 9275
rect 29628 9267 29640 9275
rect 29660 9267 29672 9275
rect 29684 9267 29688 9275
rect 29692 9267 29704 9275
rect 29724 9267 29736 9275
rect 29908 9267 29920 9275
rect 29940 9267 29952 9275
rect 29956 9267 29960 9275
rect 29972 9267 29984 9275
rect 30004 9267 30016 9275
rect 30020 9267 30032 9275
rect 30036 9267 30040 9275
rect 30060 9267 30064 9275
rect 30068 9267 30080 9275
rect 30092 9267 30096 9275
rect 30100 9267 30104 9275
rect 30124 9267 30128 9275
rect 30132 9267 30144 9275
rect 30156 9267 30160 9275
rect 30164 9267 30168 9275
rect 30216 9267 30220 9275
rect 30224 9267 30236 9275
rect 30248 9267 30252 9275
rect 30256 9267 30260 9275
rect 30372 9267 30376 9275
rect 30380 9267 30384 9275
rect 30404 9267 30408 9275
rect 30412 9267 30416 9275
rect 30428 9267 30440 9275
rect 30444 9267 30448 9275
rect 30468 9267 30472 9275
rect 30476 9267 30488 9275
rect 30492 9267 30504 9275
rect 30508 9267 30512 9275
rect 30532 9267 30536 9275
rect 30540 9267 30544 9275
rect 30688 9267 30692 9275
rect 30696 9267 30700 9275
rect 30720 9267 30724 9275
rect 30728 9267 30740 9275
rect 30744 9267 30756 9275
rect 30760 9267 30764 9275
rect 30892 9267 30896 9275
rect 30900 9267 30912 9275
rect 30916 9267 30928 9275
rect 30932 9267 30936 9275
rect 30956 9267 30960 9275
rect 30964 9267 30976 9275
rect 30988 9267 30992 9275
rect 30996 9267 31000 9275
rect 31020 9267 31024 9275
rect 31028 9267 31032 9275
rect 31176 9267 31180 9275
rect 31184 9267 31188 9275
rect 31208 9267 31212 9275
rect 31216 9267 31228 9275
rect 31232 9267 31244 9275
rect 31248 9267 31252 9275
rect 31272 9267 31276 9275
rect 31280 9267 31292 9275
rect 31300 9267 31316 9275
rect 31324 9267 31336 9275
rect 31340 9267 31344 9275
rect 31360 9267 31384 9275
rect 31392 9267 31408 9275
rect 31416 9267 31440 9275
rect 31456 9267 31460 9275
rect 31464 9267 31476 9275
rect 31480 9267 31492 9275
rect 31496 9267 31500 9275
rect 31548 9267 31552 9275
rect 31556 9267 31568 9275
rect 31572 9267 31584 9275
rect 31588 9267 31592 9275
rect 31848 9267 31852 9275
rect 31856 9267 31860 9275
rect 31880 9267 31884 9275
rect 31888 9267 31892 9275
rect 31904 9267 31916 9275
rect 31920 9267 31924 9275
rect 31940 9267 31964 9275
rect 31972 9267 31988 9275
rect 32000 9267 32028 9275
rect 32036 9267 32052 9275
rect 32064 9267 32080 9275
rect 32088 9267 32120 9275
rect 32128 9267 32144 9275
rect 32152 9267 32176 9275
rect 32192 9267 32196 9275
rect 32200 9267 32212 9275
rect 32220 9267 32236 9275
rect 32244 9267 32256 9275
rect 32260 9267 32264 9275
rect 32284 9267 32288 9275
rect 32292 9267 32304 9275
rect 32312 9267 32328 9275
rect 32336 9267 32368 9275
rect 32376 9267 32392 9275
rect 32408 9267 32424 9275
rect 32440 9267 32444 9275
rect 32448 9267 32460 9275
rect 32472 9267 32476 9275
rect 32480 9267 32484 9275
rect 32496 9267 32508 9275
rect 32512 9267 32524 9275
rect 32532 9267 32548 9275
rect 32564 9267 32580 9275
rect 32588 9267 32600 9275
rect 32604 9267 32616 9275
rect 32628 9267 32632 9275
rect 32636 9267 32640 9275
rect 32652 9267 32664 9275
rect 32668 9267 32672 9275
rect 32688 9267 32704 9275
rect 32720 9267 32736 9275
rect 32744 9267 32776 9275
rect 32784 9267 32800 9275
rect 32816 9267 32828 9275
rect 32832 9267 32844 9275
rect 32848 9267 32860 9275
rect 32880 9267 32892 9275
rect 32908 9267 32920 9275
rect 32924 9267 32936 9275
rect 32940 9267 32952 9275
rect 32972 9267 32984 9275
rect 33000 9267 33024 9275
rect 33032 9267 33048 9275
rect 33064 9267 33068 9275
rect 33072 9267 33076 9275
rect 33088 9267 33100 9275
rect 33104 9267 33116 9275
rect 33128 9267 33132 9275
rect 33136 9267 33140 9275
rect 33160 9267 33164 9275
rect 33168 9267 33172 9275
rect 33192 9267 33196 9275
rect 33200 9267 33204 9275
rect 33224 9267 33228 9275
rect 33232 9267 33236 9275
rect 33248 9267 33260 9275
rect 33264 9267 33276 9275
rect 33288 9267 33292 9275
rect 33296 9267 33300 9275
rect 33316 9267 33364 9275
rect 33380 9267 33396 9275
rect 33412 9267 33416 9275
rect 33420 9267 33432 9275
rect 33444 9267 33448 9275
rect 33452 9267 33456 9275
rect 33476 9267 33480 9275
rect 33484 9267 33488 9275
rect 33500 9267 33512 9275
rect 33516 9267 33520 9275
rect 33540 9267 33544 9275
rect 33548 9267 33552 9275
rect 33564 9267 33576 9275
rect 33580 9267 33592 9275
rect 33604 9267 33608 9275
rect 33612 9267 33616 9275
rect 33632 9267 33648 9275
rect 33656 9267 33668 9275
rect 33672 9267 33684 9275
rect 33696 9267 33700 9275
rect 33704 9267 33708 9275
rect 33788 9267 33792 9275
rect 33796 9267 33800 9275
rect 33992 9267 33996 9275
rect 34000 9267 34004 9275
rect 34016 9267 34028 9275
rect 34032 9267 34044 9275
rect 34052 9267 34068 9275
rect 34084 9267 34088 9275
rect 34092 9267 34096 9275
rect 34108 9267 34120 9275
rect 34124 9267 34136 9275
rect 34144 9267 34160 9275
rect 34176 9267 34180 9275
rect 34184 9267 34188 9275
rect 34200 9267 34212 9275
rect 34216 9267 34228 9275
rect 34236 9267 34252 9275
rect 34268 9267 34284 9275
rect 34292 9267 34316 9275
rect 34332 9267 34344 9275
rect 34364 9267 34376 9275
rect 34380 9267 34392 9275
rect 34396 9267 34408 9275
rect 34428 9267 34440 9275
rect 34444 9267 34448 9275
rect 34572 9267 34576 9275
rect 34580 9267 34584 9275
rect 34772 9267 34776 9275
rect 34780 9267 34784 9275
rect 34856 9267 34868 9275
rect 34872 9267 34876 9275
rect 34924 9267 34928 9275
rect 34932 9267 34936 9275
rect 34948 9267 34960 9275
rect 34976 9267 34992 9275
rect 35008 9267 35032 9275
rect 35048 9267 35060 9275
rect 35064 9267 35068 9275
rect 35080 9267 35092 9275
rect 35104 9267 35108 9275
rect 35112 9267 35116 9275
rect 35128 9267 35140 9275
rect 35432 9267 35436 9275
rect 35440 9267 35444 9275
rect 35464 9267 35468 9275
rect 35472 9267 35476 9275
rect 35488 9267 35500 9275
rect 35504 9267 35516 9275
rect 35528 9267 35532 9275
rect 35536 9267 35540 9275
rect 35556 9267 35588 9275
rect 35596 9267 35608 9275
rect 35628 9267 35640 9275
rect 35648 9267 35664 9275
rect 35672 9267 35696 9275
rect 35712 9267 35728 9275
rect 35744 9267 35756 9275
rect 35768 9267 35772 9275
rect 35776 9267 35788 9275
rect 35792 9267 35796 9275
rect 35900 9267 35912 9275
rect 35932 9267 35944 9275
rect 35948 9267 35952 9275
rect 35964 9267 35976 9275
rect 36000 9267 36008 9275
rect 36016 9267 36048 9275
rect 36056 9267 36072 9275
rect 36080 9267 36092 9275
rect 36096 9267 36100 9275
rect 36120 9267 36124 9275
rect 36128 9267 36140 9275
rect 36148 9267 36164 9275
rect 36172 9267 36196 9275
rect 36212 9267 36216 9275
rect 36220 9267 36232 9275
rect 36240 9267 36256 9275
rect 36264 9267 36288 9275
rect 36304 9267 36308 9275
rect 36312 9267 36324 9275
rect 36332 9267 36348 9275
rect 36356 9267 36380 9275
rect 36396 9267 36412 9275
rect 36428 9267 36440 9275
rect 36452 9267 36456 9275
rect 36460 9267 36472 9275
rect 36476 9267 36480 9275
rect 36492 9267 36504 9275
rect 36520 9267 36532 9275
rect 36544 9267 36548 9275
rect 36552 9267 36564 9275
rect 36568 9267 36572 9275
rect 36584 9267 36596 9275
rect 36616 9267 36628 9275
rect 36632 9267 36636 9275
rect 36648 9267 36660 9275
rect 36680 9267 36692 9275
rect 36704 9267 36708 9275
rect 36712 9267 36724 9275
rect 36744 9267 36756 9275
rect 36836 9267 36848 9275
rect 36868 9267 36880 9275
rect 36884 9267 36888 9275
rect 36900 9267 36912 9275
rect 36932 9267 36944 9275
rect 36948 9267 36960 9275
rect 36972 9267 36976 9275
rect 36980 9267 36984 9275
rect 37000 9267 37016 9275
rect 37024 9267 37036 9275
rect 37048 9267 37052 9275
rect 37056 9267 37068 9275
rect 37088 9267 37100 9275
rect 37188 9267 37192 9275
rect 37196 9267 37200 9275
rect 37424 9267 37428 9275
rect 37432 9267 37436 9275
rect 37456 9267 37460 9275
rect 37464 9267 37468 9275
rect 37480 9267 37492 9275
rect 37500 9267 37524 9275
rect 37540 9267 37564 9275
rect 37580 9267 37584 9275
rect 37588 9267 37600 9275
rect 37608 9267 37624 9275
rect 37632 9267 37648 9275
rect 37660 9267 37676 9275
rect 37684 9267 37716 9275
rect 37732 9267 37744 9275
rect 37764 9267 37776 9275
rect 37788 9267 37792 9275
rect 37796 9267 37800 9275
rect 37920 9267 37932 9275
rect 37936 9267 37940 9275
rect 37956 9267 37972 9275
rect 37988 9267 38004 9275
rect 38012 9267 38044 9275
rect 38052 9267 38068 9275
rect 38076 9267 38088 9275
rect 38092 9267 38096 9275
rect 38116 9267 38120 9275
rect 38124 9267 38136 9275
rect 38140 9267 38152 9275
rect 38172 9267 38184 9275
rect 38188 9267 38192 9275
rect 38360 9267 38372 9275
rect 38376 9267 38388 9275
rect 38392 9267 38396 9275
rect 38412 9267 38428 9275
rect 38444 9267 38460 9275
rect 38468 9267 38492 9275
rect 38508 9267 38540 9275
rect 38548 9267 38560 9275
rect 38580 9267 38592 9275
rect 38596 9267 38608 9275
rect 38612 9267 38616 9275
rect 38636 9267 38640 9275
rect 38644 9267 38648 9275
rect 38664 9267 38668 9275
rect 38672 9267 38684 9275
rect 38688 9267 38692 9275
rect 38732 9267 38744 9275
rect 38756 9267 38760 9275
rect 38764 9267 38768 9275
rect 38780 9267 38792 9275
rect 38796 9267 38800 9275
rect 38816 9267 38820 9275
rect 38824 9267 38836 9275
rect 38848 9267 38852 9275
rect 38856 9267 38860 9275
rect 38872 9267 38884 9275
rect 38888 9267 38892 9275
rect 39100 9267 39104 9275
rect 39108 9267 39112 9275
rect 39208 9267 39212 9275
rect 39216 9267 39220 9275
rect 39240 9267 39244 9275
rect 39248 9267 39252 9275
rect 39264 9267 39276 9275
rect 39280 9267 39292 9275
rect 39308 9267 39324 9275
rect 39340 9267 39364 9275
rect 39372 9267 39388 9275
rect 39404 9267 39444 9275
rect 39460 9267 39464 9275
rect 39468 9267 39472 9275
rect 39484 9267 39496 9275
rect 39504 9267 39520 9275
rect 39536 9267 39540 9275
rect 39544 9267 39548 9275
rect 39560 9267 39572 9275
rect 39580 9267 39596 9275
rect 39612 9267 39616 9275
rect 39620 9267 39624 9275
rect 39636 9267 39648 9275
rect 39656 9267 39680 9275
rect 39696 9267 39744 9275
rect 39760 9267 39764 9275
rect 39768 9267 39772 9275
rect 39788 9267 39836 9275
rect 39848 9267 39864 9275
rect 39880 9267 39928 9275
rect 39940 9267 39956 9275
rect 39972 9267 40000 9275
rect 30192 9237 30200 9245
rect 31456 9237 31464 9245
rect 31232 9217 31240 9225
rect 34448 9217 34456 9225
rect 36752 9217 36760 9225
rect 39584 9217 39592 9225
rect 30256 9197 30264 9205
rect 29504 9177 29512 9185
rect 29712 9177 29720 9185
rect 30640 9177 30648 9185
rect 31120 9177 31128 9185
rect 31344 9177 31352 9185
rect 32272 9177 32280 9185
rect 33760 9177 33768 9185
rect 34592 9177 34600 9185
rect 34848 9177 34856 9185
rect 35904 9177 35912 9185
rect 36848 9177 36856 9185
rect 38800 9177 38808 9185
rect 39760 9177 39768 9185
rect 39952 9177 39960 9185
rect 33008 9157 33016 9165
rect 34944 9157 34952 9165
rect 34992 9157 35000 9165
rect 29520 9137 29528 9145
rect 29792 9137 29800 9145
rect 29936 9137 29944 9145
rect 30720 9137 30728 9145
rect 31344 9137 31352 9145
rect 31392 9137 31400 9145
rect 31888 9137 31896 9145
rect 32240 9137 32248 9145
rect 32400 9137 32408 9145
rect 33744 9137 33752 9145
rect 35968 9137 35976 9145
rect 36112 9137 36120 9145
rect 36864 9137 36872 9145
rect 38768 9137 38776 9145
rect 38880 9137 38888 9145
rect 39104 9137 39112 9145
rect 39328 9137 39336 9145
rect 39488 9137 39496 9145
rect 39568 9137 39576 9145
rect 39888 9137 39896 9145
rect 29568 9117 29576 9125
rect 30128 9117 30136 9125
rect 30448 9117 30456 9125
rect 30848 9117 30856 9125
rect 30976 9117 30984 9125
rect 32112 9117 32120 9125
rect 32976 9117 32984 9125
rect 33008 9117 33016 9125
rect 33632 9117 33640 9125
rect 36384 9117 36392 9125
rect 37744 9117 37752 9125
rect 37920 9117 37928 9125
rect 39392 9117 39400 9125
rect 39408 9117 39416 9125
rect 30112 9097 30120 9105
rect 30496 9097 30504 9105
rect 31792 9097 31800 9105
rect 32672 9097 32680 9105
rect 33520 9097 33528 9105
rect 34144 9097 34152 9105
rect 34336 9097 34344 9105
rect 34720 9097 34728 9105
rect 35024 9097 35032 9105
rect 35072 9097 35080 9105
rect 35120 9097 35128 9105
rect 38224 9097 38232 9105
rect 39216 9097 39224 9105
rect 39408 9097 39416 9105
rect 39904 9097 39912 9105
rect 34064 9077 34072 9085
rect 29484 9067 29488 9075
rect 29492 9067 29504 9075
rect 29624 9067 29628 9075
rect 29632 9067 29636 9075
rect 29656 9067 29660 9075
rect 29664 9067 29668 9075
rect 29680 9067 29692 9075
rect 29696 9067 29700 9075
rect 29720 9067 29724 9075
rect 29728 9067 29740 9075
rect 29748 9067 29764 9075
rect 29772 9067 29796 9075
rect 29812 9067 29828 9075
rect 29844 9067 29856 9075
rect 29868 9067 29872 9075
rect 29876 9067 29888 9075
rect 29892 9067 29896 9075
rect 30000 9067 30012 9075
rect 30024 9067 30028 9075
rect 30032 9067 30044 9075
rect 30048 9067 30052 9075
rect 30064 9067 30076 9075
rect 30092 9067 30108 9075
rect 30124 9067 30148 9075
rect 30156 9067 30172 9075
rect 30180 9067 30204 9075
rect 30216 9067 30240 9075
rect 30248 9067 30264 9075
rect 30272 9067 30296 9075
rect 30312 9067 30328 9075
rect 30336 9067 30360 9075
rect 30376 9067 30388 9075
rect 30392 9067 30396 9075
rect 30408 9067 30420 9075
rect 30432 9067 30436 9075
rect 30440 9067 30452 9075
rect 30468 9067 30516 9075
rect 30532 9067 30548 9075
rect 30564 9067 30568 9075
rect 30572 9067 30584 9075
rect 30596 9067 30600 9075
rect 30604 9067 30608 9075
rect 30688 9067 30692 9075
rect 30696 9067 30700 9075
rect 30720 9067 30724 9075
rect 30728 9067 30732 9075
rect 30796 9067 30800 9075
rect 30804 9067 30808 9075
rect 30828 9067 30832 9075
rect 30836 9067 30840 9075
rect 30852 9067 30864 9075
rect 30868 9067 30872 9075
rect 30888 9067 30912 9075
rect 30920 9067 30936 9075
rect 30944 9067 30976 9075
rect 30984 9067 31000 9075
rect 31016 9067 31028 9075
rect 31036 9067 31068 9075
rect 31076 9067 31092 9075
rect 31108 9067 31120 9075
rect 31132 9067 31136 9075
rect 31140 9067 31152 9075
rect 31172 9067 31184 9075
rect 31328 9067 31340 9075
rect 31360 9067 31372 9075
rect 31376 9067 31388 9075
rect 31392 9067 31404 9075
rect 31424 9067 31436 9075
rect 31444 9067 31476 9075
rect 31484 9067 31500 9075
rect 31516 9067 31520 9075
rect 31524 9067 31528 9075
rect 31548 9067 31552 9075
rect 31556 9067 31568 9075
rect 31580 9067 31584 9075
rect 31588 9067 31592 9075
rect 31672 9067 31676 9075
rect 31680 9067 31684 9075
rect 31696 9067 31708 9075
rect 31712 9067 31716 9075
rect 31736 9067 31740 9075
rect 31744 9067 31748 9075
rect 31764 9067 31780 9075
rect 31788 9067 31820 9075
rect 31828 9067 31844 9075
rect 31860 9067 31864 9075
rect 31868 9067 31872 9075
rect 31892 9067 31896 9075
rect 31900 9067 31912 9075
rect 31924 9067 31928 9075
rect 31932 9067 31936 9075
rect 31984 9067 31988 9075
rect 31992 9067 32000 9075
rect 32016 9067 32020 9075
rect 32024 9067 32028 9075
rect 32040 9067 32052 9075
rect 32056 9067 32060 9075
rect 32108 9067 32112 9075
rect 32116 9067 32120 9075
rect 32132 9067 32144 9075
rect 32148 9067 32160 9075
rect 32172 9067 32176 9075
rect 32180 9067 32184 9075
rect 32200 9067 32216 9075
rect 32224 9067 32236 9075
rect 32240 9067 32252 9075
rect 32264 9067 32268 9075
rect 32272 9067 32276 9075
rect 32292 9067 32308 9075
rect 32316 9067 32328 9075
rect 32332 9067 32344 9075
rect 32356 9067 32360 9075
rect 32364 9067 32368 9075
rect 32380 9067 32392 9075
rect 32396 9067 32400 9075
rect 32420 9067 32424 9075
rect 32428 9067 32432 9075
rect 32452 9067 32456 9075
rect 32460 9067 32464 9075
rect 32484 9067 32488 9075
rect 32492 9067 32504 9075
rect 32516 9067 32520 9075
rect 32524 9067 32528 9075
rect 32608 9067 32612 9075
rect 32616 9067 32620 9075
rect 32632 9067 32644 9075
rect 32648 9067 32660 9075
rect 32672 9067 32676 9075
rect 32680 9067 32684 9075
rect 32812 9067 32816 9075
rect 32820 9067 32824 9075
rect 32904 9067 32908 9075
rect 32912 9067 32916 9075
rect 33044 9067 33048 9075
rect 33052 9067 33056 9075
rect 33068 9067 33080 9075
rect 33084 9067 33096 9075
rect 33104 9067 33120 9075
rect 33136 9067 33152 9075
rect 33160 9067 33184 9075
rect 33200 9067 33212 9075
rect 33232 9067 33244 9075
rect 33248 9067 33260 9075
rect 33264 9067 33276 9075
rect 33296 9067 33308 9075
rect 33324 9067 33336 9075
rect 33340 9067 33352 9075
rect 33356 9067 33368 9075
rect 33388 9067 33400 9075
rect 33412 9067 33416 9075
rect 33420 9067 33432 9075
rect 33452 9067 33464 9075
rect 33476 9067 33480 9075
rect 33484 9067 33496 9075
rect 33500 9067 33504 9075
rect 33796 9067 33808 9075
rect 33812 9067 33824 9075
rect 33828 9067 33840 9075
rect 33860 9067 33872 9075
rect 33876 9067 33888 9075
rect 33892 9067 33904 9075
rect 34016 9067 34028 9075
rect 34040 9067 34044 9075
rect 34048 9067 34060 9075
rect 34064 9067 34068 9075
rect 34108 9067 34120 9075
rect 34132 9067 34136 9075
rect 34140 9067 34152 9075
rect 34156 9067 34160 9075
rect 34296 9067 34308 9075
rect 34312 9067 34316 9075
rect 34328 9067 34340 9075
rect 34356 9067 34372 9075
rect 34380 9067 34412 9075
rect 34420 9067 34436 9075
rect 34444 9067 34468 9075
rect 34484 9067 34488 9075
rect 34492 9067 34504 9075
rect 34512 9067 34528 9075
rect 34536 9067 34560 9075
rect 34576 9067 34588 9075
rect 34608 9067 34620 9075
rect 34632 9067 34636 9075
rect 34640 9067 34652 9075
rect 34656 9067 34660 9075
rect 34672 9067 34684 9075
rect 34888 9067 34900 9075
rect 34904 9067 34908 9075
rect 34920 9067 34932 9075
rect 34952 9067 34964 9075
rect 34976 9067 34980 9075
rect 34984 9067 34996 9075
rect 35016 9067 35028 9075
rect 35040 9067 35044 9075
rect 35048 9067 35060 9075
rect 35064 9067 35068 9075
rect 35204 9067 35216 9075
rect 35220 9067 35232 9075
rect 35236 9067 35240 9075
rect 35260 9067 35264 9075
rect 35268 9067 35280 9075
rect 35288 9067 35304 9075
rect 35312 9067 35336 9075
rect 35352 9067 35356 9075
rect 35360 9067 35372 9075
rect 35392 9067 35404 9075
rect 35424 9067 35436 9075
rect 35456 9067 35468 9075
rect 35472 9067 35476 9075
rect 35492 9067 35516 9075
rect 35524 9067 35540 9075
rect 35548 9067 35564 9075
rect 35572 9067 35584 9075
rect 35600 9067 35616 9075
rect 35624 9067 35656 9075
rect 35672 9067 35696 9075
rect 35712 9067 35724 9075
rect 35744 9067 35756 9075
rect 35768 9067 35772 9075
rect 35776 9067 35780 9075
rect 35860 9067 35864 9075
rect 35868 9067 35880 9075
rect 36024 9067 36036 9075
rect 36040 9067 36044 9075
rect 36056 9067 36068 9075
rect 36084 9067 36100 9075
rect 36116 9067 36164 9075
rect 36180 9067 36196 9075
rect 36208 9067 36256 9075
rect 36272 9067 36288 9075
rect 36304 9067 36308 9075
rect 36312 9067 36324 9075
rect 36336 9067 36340 9075
rect 36344 9067 36348 9075
rect 36368 9067 36372 9075
rect 36376 9067 36380 9075
rect 36392 9067 36404 9075
rect 36408 9067 36412 9075
rect 36432 9067 36436 9075
rect 36440 9067 36444 9075
rect 36456 9067 36468 9075
rect 36472 9067 36484 9075
rect 36492 9067 36508 9075
rect 36524 9067 36528 9075
rect 36532 9067 36536 9075
rect 36548 9067 36560 9075
rect 36564 9067 36576 9075
rect 36588 9067 36592 9075
rect 36596 9067 36600 9075
rect 36616 9067 36664 9075
rect 36680 9067 36696 9075
rect 36712 9067 36724 9075
rect 36736 9067 36740 9075
rect 36744 9067 36756 9075
rect 36828 9067 36832 9075
rect 36836 9067 36848 9075
rect 36868 9067 36880 9075
rect 36884 9067 36888 9075
rect 36952 9067 36956 9075
rect 36960 9067 36964 9075
rect 36984 9067 36988 9075
rect 36992 9067 36996 9075
rect 37188 9067 37192 9075
rect 37196 9067 37200 9075
rect 37320 9067 37332 9075
rect 37336 9067 37348 9075
rect 37352 9067 37364 9075
rect 37384 9067 37396 9075
rect 37412 9067 37436 9075
rect 37444 9067 37460 9075
rect 37476 9067 37492 9075
rect 37500 9067 37512 9075
rect 37516 9067 37528 9075
rect 37540 9067 37544 9075
rect 37548 9067 37552 9075
rect 37568 9067 37584 9075
rect 37592 9067 37604 9075
rect 37608 9067 37620 9075
rect 37632 9067 37636 9075
rect 37640 9067 37644 9075
rect 37660 9067 37676 9075
rect 37684 9067 37696 9075
rect 37700 9067 37712 9075
rect 37732 9067 37744 9075
rect 37832 9067 37836 9075
rect 37840 9067 37852 9075
rect 37856 9067 37860 9075
rect 37880 9067 37884 9075
rect 37888 9067 37900 9075
rect 37916 9067 37940 9075
rect 37948 9067 37964 9075
rect 37980 9067 37996 9075
rect 38012 9067 38016 9075
rect 38020 9067 38032 9075
rect 38036 9067 38048 9075
rect 38052 9067 38056 9075
rect 38072 9067 38088 9075
rect 38104 9067 38120 9075
rect 38128 9067 38152 9075
rect 38168 9067 38192 9075
rect 38200 9067 38212 9075
rect 38224 9067 38228 9075
rect 38232 9067 38244 9075
rect 38248 9067 38252 9075
rect 38264 9067 38276 9075
rect 38288 9067 38292 9075
rect 38296 9067 38308 9075
rect 38324 9067 38348 9075
rect 38356 9067 38368 9075
rect 38380 9067 38384 9075
rect 38388 9067 38400 9075
rect 38640 9067 38652 9075
rect 38656 9067 38660 9075
rect 38732 9067 38744 9075
rect 38764 9067 38776 9075
rect 38780 9067 38784 9075
rect 38796 9067 38808 9075
rect 38816 9067 38840 9075
rect 38856 9067 38904 9075
rect 38920 9067 38932 9075
rect 38952 9067 38964 9075
rect 38976 9067 38980 9075
rect 38984 9067 38996 9075
rect 39108 9067 39120 9075
rect 39124 9067 39128 9075
rect 39232 9067 39244 9075
rect 39248 9067 39252 9075
rect 39264 9067 39276 9075
rect 39288 9067 39292 9075
rect 39296 9067 39300 9075
rect 39316 9067 39332 9075
rect 39340 9067 39364 9075
rect 39380 9067 39396 9075
rect 39412 9067 39436 9075
rect 39452 9067 39464 9075
rect 39484 9067 39496 9075
rect 39500 9067 39512 9075
rect 39516 9067 39520 9075
rect 39536 9067 39540 9075
rect 39544 9067 39548 9075
rect 39568 9067 39572 9075
rect 39576 9067 39588 9075
rect 39592 9067 39596 9075
rect 39636 9067 39648 9075
rect 39660 9067 39664 9075
rect 39668 9067 39680 9075
rect 39684 9067 39688 9075
rect 39700 9067 39712 9075
rect 39724 9067 39728 9075
rect 39732 9067 39744 9075
rect 39748 9067 39752 9075
rect 39764 9067 39776 9075
rect 39856 9067 39868 9075
rect 39888 9067 39900 9075
rect 39904 9067 39916 9075
rect 39920 9067 39932 9075
rect 39948 9067 39964 9075
rect 39972 9067 40000 9075
rect 33136 9057 33144 9065
rect 37072 9057 37080 9065
rect 37168 9057 37176 9065
rect 29904 9037 29912 9045
rect 30464 9037 30472 9045
rect 31328 9037 31336 9045
rect 32224 9037 32232 9045
rect 32736 9037 32744 9045
rect 33360 9037 33368 9045
rect 33872 9037 33880 9045
rect 34080 9037 34088 9045
rect 34224 9037 34232 9045
rect 35456 9037 35464 9045
rect 35936 9037 35944 9045
rect 38880 9037 38888 9045
rect 31920 9017 31928 9025
rect 32336 9017 32344 9025
rect 32464 9017 32472 9025
rect 32880 9017 32888 9025
rect 33696 9017 33704 9025
rect 35984 9017 35992 9025
rect 36064 9017 36072 9025
rect 29664 8997 29672 9005
rect 30128 8997 30136 9005
rect 30496 8997 30504 9005
rect 30656 8997 30664 9005
rect 31232 8997 31240 9005
rect 31616 8997 31624 9005
rect 31712 8997 31720 9005
rect 32224 8997 32232 9005
rect 32992 8997 33000 9005
rect 33264 8997 33272 9005
rect 33728 8997 33736 9005
rect 36848 8997 36856 9005
rect 36928 8997 36936 9005
rect 37776 8997 37784 9005
rect 37952 8997 37960 9005
rect 38144 8997 38152 9005
rect 38272 8997 38280 9005
rect 38576 8997 38584 9005
rect 38976 8997 38984 9005
rect 39168 8997 39176 9005
rect 39472 8997 39480 9005
rect 39840 8997 39848 9005
rect 31888 8977 31896 8985
rect 36048 8977 36056 8985
rect 36912 8977 36920 8985
rect 37088 8977 37096 8985
rect 37408 8977 37416 8985
rect 37744 8977 37752 8985
rect 39392 8977 39400 8985
rect 39424 8977 39432 8985
rect 30176 8957 30184 8965
rect 30816 8957 30824 8965
rect 31520 8957 31528 8965
rect 31648 8957 31656 8965
rect 32256 8957 32264 8965
rect 33536 8957 33544 8965
rect 34032 8957 34040 8965
rect 34720 8957 34728 8965
rect 35088 8957 35096 8965
rect 35584 8957 35592 8965
rect 35728 8957 35736 8965
rect 36512 8957 36520 8965
rect 36656 8957 36664 8965
rect 36784 8957 36792 8965
rect 36864 8957 36872 8965
rect 36976 8957 36984 8965
rect 37856 8957 37864 8965
rect 38048 8957 38056 8965
rect 39648 8957 39656 8965
rect 35680 8917 35688 8925
rect 38128 8917 38136 8925
rect 39904 8897 39912 8905
rect 29592 8867 29596 8875
rect 29600 8867 29604 8875
rect 29624 8867 29628 8875
rect 29632 8867 29636 8875
rect 29648 8867 29660 8875
rect 29676 8867 29692 8875
rect 29708 8867 29740 8875
rect 29748 8867 29764 8875
rect 29780 8867 29796 8875
rect 29812 8867 29828 8875
rect 29844 8867 29860 8875
rect 29868 8867 29884 8875
rect 29892 8867 29924 8875
rect 29940 8867 29952 8875
rect 29956 8867 29960 8875
rect 29972 8867 29984 8875
rect 29992 8867 30008 8875
rect 30024 8867 30056 8875
rect 30064 8867 30080 8875
rect 30096 8867 30100 8875
rect 30104 8867 30108 8875
rect 30128 8867 30132 8875
rect 30136 8867 30148 8875
rect 30160 8867 30164 8875
rect 30168 8867 30172 8875
rect 30184 8867 30196 8875
rect 30460 8867 30464 8875
rect 30468 8867 30480 8875
rect 30484 8867 30488 8875
rect 30552 8867 30556 8875
rect 30560 8867 30564 8875
rect 30612 8867 30616 8875
rect 30620 8867 30632 8875
rect 30744 8867 30756 8875
rect 30760 8867 30764 8875
rect 30796 8867 30800 8875
rect 30804 8867 30816 8875
rect 30836 8867 30848 8875
rect 30852 8867 30856 8875
rect 30888 8867 30892 8875
rect 30896 8867 30908 8875
rect 30928 8867 30940 8875
rect 30944 8867 30956 8875
rect 30960 8867 30972 8875
rect 31020 8867 31032 8875
rect 31036 8867 31048 8875
rect 31052 8867 31064 8875
rect 31112 8867 31124 8875
rect 31128 8867 31140 8875
rect 31144 8867 31156 8875
rect 31204 8867 31216 8875
rect 31220 8867 31232 8875
rect 31236 8867 31248 8875
rect 31268 8867 31280 8875
rect 31608 8867 31612 8875
rect 31616 8867 31628 8875
rect 31632 8867 31636 8875
rect 31648 8867 31660 8875
rect 31676 8867 31688 8875
rect 31700 8867 31704 8875
rect 31708 8867 31720 8875
rect 31724 8867 31728 8875
rect 31744 8867 31760 8875
rect 31776 8867 31780 8875
rect 31784 8867 31796 8875
rect 31800 8867 31812 8875
rect 31832 8867 31844 8875
rect 31860 8867 31884 8875
rect 31892 8867 31908 8875
rect 31924 8867 31928 8875
rect 31932 8867 31936 8875
rect 31948 8867 31960 8875
rect 31964 8867 31976 8875
rect 31984 8867 32000 8875
rect 32016 8867 32032 8875
rect 32040 8867 32064 8875
rect 32080 8867 32096 8875
rect 32112 8867 32124 8875
rect 32128 8867 32140 8875
rect 32144 8867 32156 8875
rect 32176 8867 32188 8875
rect 32192 8867 32196 8875
rect 32228 8867 32232 8875
rect 32236 8867 32248 8875
rect 32268 8867 32280 8875
rect 32284 8867 32288 8875
rect 32544 8867 32548 8875
rect 32552 8867 32564 8875
rect 32584 8867 32596 8875
rect 32600 8867 32604 8875
rect 32636 8867 32640 8875
rect 32644 8867 32656 8875
rect 32676 8867 32688 8875
rect 32692 8867 32696 8875
rect 32708 8867 32720 8875
rect 32740 8867 32752 8875
rect 32768 8867 32816 8875
rect 32828 8867 32844 8875
rect 32860 8867 32908 8875
rect 32924 8867 32936 8875
rect 32940 8867 32944 8875
rect 32956 8867 32968 8875
rect 32976 8867 33000 8875
rect 33016 8867 33040 8875
rect 33048 8867 33060 8875
rect 33068 8867 33092 8875
rect 33108 8867 33120 8875
rect 33124 8867 33128 8875
rect 33140 8867 33152 8875
rect 33164 8867 33168 8875
rect 33172 8867 33184 8875
rect 33188 8867 33192 8875
rect 33232 8867 33244 8875
rect 33256 8867 33260 8875
rect 33264 8867 33276 8875
rect 33280 8867 33284 8875
rect 33296 8867 33308 8875
rect 33508 8867 33512 8875
rect 33516 8867 33528 8875
rect 33548 8867 33560 8875
rect 33564 8867 33568 8875
rect 33916 8867 33920 8875
rect 33924 8867 33936 8875
rect 34008 8867 34012 8875
rect 34016 8867 34028 8875
rect 34048 8867 34060 8875
rect 34064 8867 34068 8875
rect 34100 8867 34104 8875
rect 34108 8867 34120 8875
rect 34140 8867 34152 8875
rect 34156 8867 34160 8875
rect 34172 8867 34184 8875
rect 34204 8867 34216 8875
rect 34220 8867 34224 8875
rect 34236 8867 34248 8875
rect 34260 8867 34264 8875
rect 34268 8867 34280 8875
rect 34296 8867 34344 8875
rect 34356 8867 34372 8875
rect 34388 8867 34436 8875
rect 34452 8867 34464 8875
rect 34480 8867 34528 8875
rect 34544 8867 34560 8875
rect 34576 8867 34592 8875
rect 34608 8867 34624 8875
rect 34640 8867 34688 8875
rect 34704 8867 34716 8875
rect 34720 8867 34724 8875
rect 34736 8867 34748 8875
rect 34760 8867 34764 8875
rect 34768 8867 34780 8875
rect 34796 8867 34820 8875
rect 34828 8867 34840 8875
rect 34852 8867 34856 8875
rect 34860 8867 34872 8875
rect 34892 8867 34904 8875
rect 34924 8867 34936 8875
rect 34956 8867 34968 8875
rect 34972 8867 34976 8875
rect 34988 8867 35000 8875
rect 35012 8867 35016 8875
rect 35020 8867 35024 8875
rect 35072 8867 35076 8875
rect 35080 8867 35092 8875
rect 35104 8867 35108 8875
rect 35112 8867 35116 8875
rect 35204 8867 35216 8875
rect 35220 8867 35224 8875
rect 35236 8867 35248 8875
rect 35268 8867 35280 8875
rect 35296 8867 35336 8875
rect 35352 8867 35376 8875
rect 35392 8867 35404 8875
rect 35424 8867 35436 8875
rect 35448 8867 35452 8875
rect 35456 8867 35460 8875
rect 35500 8867 35512 8875
rect 35524 8867 35528 8875
rect 35532 8867 35544 8875
rect 35548 8867 35552 8875
rect 35568 8867 35584 8875
rect 35600 8867 35616 8875
rect 35624 8867 35648 8875
rect 35664 8867 35704 8875
rect 35716 8867 35732 8875
rect 35748 8867 35780 8875
rect 35788 8867 35800 8875
rect 35816 8867 35832 8875
rect 35840 8867 35856 8875
rect 35864 8867 35876 8875
rect 35880 8867 35884 8875
rect 35904 8867 35908 8875
rect 35912 8867 35924 8875
rect 35936 8867 35940 8875
rect 35944 8867 35948 8875
rect 35968 8867 35972 8875
rect 35976 8867 35988 8875
rect 36000 8867 36004 8875
rect 36008 8867 36012 8875
rect 36024 8867 36036 8875
rect 36040 8867 36044 8875
rect 36060 8867 36076 8875
rect 36092 8867 36108 8875
rect 36116 8867 36148 8875
rect 36156 8867 36172 8875
rect 36180 8867 36204 8875
rect 36216 8867 36240 8875
rect 36248 8867 36264 8875
rect 36272 8867 36296 8875
rect 36312 8867 36324 8875
rect 36344 8867 36356 8875
rect 36368 8867 36372 8875
rect 36376 8867 36380 8875
rect 36392 8867 36404 8875
rect 36408 8867 36420 8875
rect 36432 8867 36436 8875
rect 36440 8867 36444 8875
rect 36456 8867 36468 8875
rect 36472 8867 36476 8875
rect 36492 8867 36496 8875
rect 36500 8867 36512 8875
rect 36524 8867 36528 8875
rect 36532 8867 36536 8875
rect 36548 8867 36560 8875
rect 36564 8867 36568 8875
rect 36616 8867 36620 8875
rect 36624 8867 36628 8875
rect 36708 8867 36712 8875
rect 36716 8867 36720 8875
rect 36732 8867 36744 8875
rect 36748 8867 36760 8875
rect 36768 8867 36784 8875
rect 36800 8867 36816 8875
rect 36824 8867 36836 8875
rect 36840 8867 36852 8875
rect 36864 8867 36868 8875
rect 36872 8867 36876 8875
rect 36892 8867 36908 8875
rect 36916 8867 36928 8875
rect 36932 8867 36944 8875
rect 36952 8867 36968 8875
rect 36984 8867 37032 8875
rect 37048 8867 37064 8875
rect 37080 8867 37084 8875
rect 37088 8867 37100 8875
rect 37112 8867 37116 8875
rect 37120 8867 37124 8875
rect 37144 8867 37148 8875
rect 37152 8867 37156 8875
rect 37168 8867 37180 8875
rect 37184 8867 37188 8875
rect 37204 8867 37220 8875
rect 37236 8867 37276 8875
rect 37292 8867 37308 8875
rect 37316 8867 37328 8875
rect 37332 8867 37344 8875
rect 37352 8867 37368 8875
rect 37384 8867 37400 8875
rect 37408 8867 37420 8875
rect 37424 8867 37436 8875
rect 37448 8867 37452 8875
rect 37456 8867 37460 8875
rect 37472 8867 37484 8875
rect 37488 8867 37492 8875
rect 37540 8867 37544 8875
rect 37548 8867 37552 8875
rect 37564 8867 37576 8875
rect 37580 8867 37584 8875
rect 37680 8867 37684 8875
rect 37688 8867 37692 8875
rect 37704 8867 37716 8875
rect 37728 8867 37732 8875
rect 37736 8867 37748 8875
rect 37764 8867 37788 8875
rect 37804 8867 37820 8875
rect 37836 8867 37848 8875
rect 37860 8867 37864 8875
rect 37868 8867 37872 8875
rect 37884 8867 37896 8875
rect 37900 8867 37904 8875
rect 37920 8867 37924 8875
rect 37928 8867 37940 8875
rect 37952 8867 37956 8875
rect 37960 8867 37964 8875
rect 37976 8867 37988 8875
rect 37992 8867 37996 8875
rect 38012 8867 38016 8875
rect 38020 8867 38032 8875
rect 38044 8867 38048 8875
rect 38052 8867 38056 8875
rect 38068 8867 38080 8875
rect 38084 8867 38088 8875
rect 38104 8867 38120 8875
rect 38136 8867 38152 8875
rect 38160 8867 38192 8875
rect 38200 8867 38212 8875
rect 38232 8867 38244 8875
rect 38248 8867 38260 8875
rect 38264 8867 38276 8875
rect 38296 8867 38308 8875
rect 38316 8867 38348 8875
rect 38356 8867 38368 8875
rect 38388 8867 38400 8875
rect 38412 8867 38416 8875
rect 38420 8867 38432 8875
rect 38568 8867 38572 8875
rect 38576 8867 38588 8875
rect 38592 8867 38596 8875
rect 38608 8867 38620 8875
rect 38636 8867 38648 8875
rect 38660 8867 38664 8875
rect 38668 8867 38680 8875
rect 38684 8867 38688 8875
rect 38700 8867 38712 8875
rect 38728 8867 38744 8875
rect 38760 8867 38784 8875
rect 38792 8867 38808 8875
rect 38816 8867 38828 8875
rect 38832 8867 38836 8875
rect 38856 8867 38860 8875
rect 38864 8867 38876 8875
rect 38880 8867 38892 8875
rect 38896 8867 38900 8875
rect 38916 8867 38940 8875
rect 38948 8867 38964 8875
rect 38972 8867 38996 8875
rect 39012 8867 39024 8875
rect 39044 8867 39056 8875
rect 39068 8867 39072 8875
rect 39076 8867 39088 8875
rect 39092 8867 39096 8875
rect 39108 8867 39120 8875
rect 39136 8867 39148 8875
rect 39160 8867 39164 8875
rect 39168 8867 39180 8875
rect 39184 8867 39188 8875
rect 39200 8867 39212 8875
rect 39228 8867 39240 8875
rect 39252 8867 39256 8875
rect 39260 8867 39272 8875
rect 39276 8867 39280 8875
rect 39292 8867 39304 8875
rect 39320 8867 39332 8875
rect 39344 8867 39348 8875
rect 39352 8867 39364 8875
rect 39368 8867 39372 8875
rect 39384 8867 39396 8875
rect 39416 8867 39428 8875
rect 39432 8867 39436 8875
rect 39448 8867 39460 8875
rect 39476 8867 39492 8875
rect 39500 8867 39532 8875
rect 39540 8867 39552 8875
rect 39572 8867 39584 8875
rect 39592 8867 39624 8875
rect 39632 8867 39644 8875
rect 39664 8867 39676 8875
rect 39688 8867 39692 8875
rect 39696 8867 39708 8875
rect 39728 8867 39740 8875
rect 39752 8867 39756 8875
rect 39760 8867 39772 8875
rect 39776 8867 39780 8875
rect 39792 8867 39804 8875
rect 39820 8867 39836 8875
rect 39852 8867 39876 8875
rect 39884 8867 39900 8875
rect 39908 8867 39932 8875
rect 39948 8867 39964 8875
rect 39972 8867 39996 8875
rect 36160 8857 36168 8865
rect 36960 8857 36968 8865
rect 31888 8837 31896 8845
rect 29920 8817 29928 8825
rect 32192 8817 32200 8825
rect 33600 8817 33608 8825
rect 36928 8817 36936 8825
rect 38736 8817 38744 8825
rect 38864 8817 38872 8825
rect 39280 8817 39288 8825
rect 30384 8797 30392 8805
rect 32112 8797 32120 8805
rect 35088 8797 35096 8805
rect 35760 8797 35768 8805
rect 29904 8777 29912 8785
rect 29952 8777 29960 8785
rect 30832 8777 30840 8785
rect 31104 8777 31112 8785
rect 31264 8777 31272 8785
rect 31680 8777 31688 8785
rect 31856 8777 31864 8785
rect 32512 8777 32520 8785
rect 33536 8777 33544 8785
rect 33648 8777 33656 8785
rect 34048 8777 34056 8785
rect 34416 8777 34424 8785
rect 35488 8777 35496 8785
rect 35728 8777 35736 8785
rect 36656 8777 36664 8785
rect 38208 8777 38216 8785
rect 38368 8777 38376 8785
rect 38464 8777 38472 8785
rect 38528 8777 38536 8785
rect 39552 8777 39560 8785
rect 30864 8757 30872 8765
rect 31360 8757 31368 8765
rect 29552 8737 29560 8745
rect 29632 8737 29640 8745
rect 29712 8737 29720 8745
rect 29968 8737 29976 8745
rect 29984 8737 29992 8745
rect 30400 8737 30408 8745
rect 30816 8737 30824 8745
rect 31408 8737 31416 8745
rect 31712 8737 31720 8745
rect 36096 8737 36104 8745
rect 37552 8737 37560 8745
rect 37952 8737 37960 8745
rect 38048 8737 38056 8745
rect 38256 8737 38264 8745
rect 38608 8737 38616 8745
rect 39504 8737 39512 8745
rect 39856 8737 39864 8745
rect 29488 8717 29496 8725
rect 29568 8717 29576 8725
rect 30064 8717 30072 8725
rect 30624 8717 30632 8725
rect 31408 8717 31416 8725
rect 31456 8717 31464 8725
rect 34320 8717 34328 8725
rect 34816 8717 34824 8725
rect 35760 8717 35768 8725
rect 35936 8717 35944 8725
rect 36000 8717 36008 8725
rect 36080 8717 36088 8725
rect 36128 8717 36136 8725
rect 36976 8717 36984 8725
rect 37744 8717 37752 8725
rect 38320 8717 38328 8725
rect 39744 8717 39752 8725
rect 39952 8717 39960 8725
rect 29472 8697 29480 8705
rect 29760 8697 29768 8705
rect 30432 8697 30440 8705
rect 30960 8697 30968 8705
rect 31136 8697 31144 8705
rect 31872 8697 31880 8705
rect 32016 8697 32024 8705
rect 32192 8697 32200 8705
rect 32336 8697 32344 8705
rect 32592 8697 32600 8705
rect 32784 8697 32792 8705
rect 33184 8697 33192 8705
rect 33568 8697 33576 8705
rect 33664 8697 33672 8705
rect 33808 8697 33816 8705
rect 33888 8697 33896 8705
rect 33968 8697 33976 8705
rect 34416 8697 34424 8705
rect 36544 8697 36552 8705
rect 36880 8697 36888 8705
rect 37488 8697 37496 8705
rect 38768 8697 38776 8705
rect 39088 8697 39096 8705
rect 39712 8697 39720 8705
rect 29440 8677 29448 8685
rect 29808 8677 29816 8685
rect 33008 8677 33016 8685
rect 33408 8677 33416 8685
rect 33424 8677 33432 8685
rect 35264 8677 35272 8685
rect 35376 8677 35384 8685
rect 37600 8677 37608 8685
rect 29420 8667 29424 8675
rect 29428 8667 29432 8675
rect 29444 8667 29456 8675
rect 29472 8667 29488 8675
rect 29496 8667 29512 8675
rect 29520 8667 29532 8675
rect 29548 8667 29564 8675
rect 29572 8667 29588 8675
rect 29600 8667 29608 8675
rect 29628 8667 29640 8675
rect 29648 8667 29664 8675
rect 29672 8667 29684 8675
rect 29704 8667 29716 8675
rect 29724 8667 29740 8675
rect 29748 8667 29764 8675
rect 29780 8667 29796 8675
rect 29812 8667 29816 8675
rect 29820 8667 29832 8675
rect 29852 8667 29864 8675
rect 29868 8667 29872 8675
rect 29944 8667 29956 8675
rect 30076 8667 30080 8675
rect 30084 8667 30088 8675
rect 30108 8667 30112 8675
rect 30116 8667 30120 8675
rect 30132 8667 30144 8675
rect 30160 8667 30176 8675
rect 30184 8667 30200 8675
rect 30208 8667 30232 8675
rect 30248 8667 30264 8675
rect 30272 8667 30288 8675
rect 30304 8667 30320 8675
rect 30328 8667 30340 8675
rect 30352 8667 30356 8675
rect 30360 8667 30364 8675
rect 30492 8667 30496 8675
rect 30500 8667 30512 8675
rect 30532 8667 30544 8675
rect 30548 8667 30560 8675
rect 30568 8667 30584 8675
rect 30600 8667 30616 8675
rect 30624 8667 30640 8675
rect 30656 8667 30660 8675
rect 30664 8667 30668 8675
rect 30688 8667 30692 8675
rect 30696 8667 30708 8675
rect 30712 8667 30724 8675
rect 30728 8667 30732 8675
rect 30752 8667 30756 8675
rect 30760 8667 30764 8675
rect 30860 8667 30864 8675
rect 30868 8667 30880 8675
rect 30884 8667 30896 8675
rect 30900 8667 30904 8675
rect 30924 8667 30928 8675
rect 30932 8667 30936 8675
rect 30984 8667 30988 8675
rect 30992 8667 30996 8675
rect 31016 8667 31020 8675
rect 31024 8667 31028 8675
rect 31040 8667 31052 8675
rect 31056 8667 31060 8675
rect 31076 8667 31092 8675
rect 31108 8667 31156 8675
rect 31172 8667 31184 8675
rect 31188 8667 31192 8675
rect 31204 8667 31216 8675
rect 31228 8667 31232 8675
rect 31236 8667 31248 8675
rect 31264 8667 31288 8675
rect 31296 8667 31308 8675
rect 31320 8667 31324 8675
rect 31328 8667 31340 8675
rect 31360 8667 31372 8675
rect 31392 8667 31404 8675
rect 31424 8667 31436 8675
rect 31440 8667 31444 8675
rect 31456 8667 31468 8675
rect 31476 8667 31500 8675
rect 31516 8667 31548 8675
rect 31556 8667 31572 8675
rect 31588 8667 31600 8675
rect 31608 8667 31624 8675
rect 31632 8667 31664 8675
rect 31680 8667 31684 8675
rect 31688 8667 31692 8675
rect 31712 8667 31716 8675
rect 31720 8667 31732 8675
rect 31836 8667 31840 8675
rect 31844 8667 31848 8675
rect 31912 8667 31916 8675
rect 31920 8667 31924 8675
rect 31944 8667 31948 8675
rect 31952 8667 31964 8675
rect 31968 8667 31980 8675
rect 31984 8667 31988 8675
rect 32008 8667 32012 8675
rect 32016 8667 32020 8675
rect 32148 8667 32152 8675
rect 32156 8667 32160 8675
rect 32180 8667 32184 8675
rect 32188 8667 32200 8675
rect 32204 8667 32216 8675
rect 32220 8667 32224 8675
rect 32272 8667 32276 8675
rect 32280 8667 32292 8675
rect 32296 8667 32308 8675
rect 32312 8667 32316 8675
rect 32336 8667 32340 8675
rect 32344 8667 32348 8675
rect 32360 8667 32372 8675
rect 32376 8667 32380 8675
rect 32400 8667 32404 8675
rect 32408 8667 32412 8675
rect 32432 8667 32436 8675
rect 32440 8667 32452 8675
rect 32464 8667 32468 8675
rect 32472 8667 32476 8675
rect 32496 8667 32500 8675
rect 32504 8667 32516 8675
rect 32520 8667 32532 8675
rect 32536 8667 32540 8675
rect 32636 8667 32640 8675
rect 32644 8667 32648 8675
rect 32744 8667 32748 8675
rect 32752 8667 32756 8675
rect 32820 8667 32824 8675
rect 32828 8667 32832 8675
rect 32852 8667 32856 8675
rect 32860 8667 32864 8675
rect 32876 8667 32888 8675
rect 32892 8667 32896 8675
rect 32916 8667 32920 8675
rect 32924 8667 32936 8675
rect 32940 8667 32952 8675
rect 32956 8667 32960 8675
rect 32976 8667 32980 8675
rect 32984 8667 32988 8675
rect 33008 8667 33012 8675
rect 33016 8667 33028 8675
rect 33032 8667 33044 8675
rect 33048 8667 33052 8675
rect 33068 8667 33084 8675
rect 33100 8667 33104 8675
rect 33108 8667 33120 8675
rect 33124 8667 33136 8675
rect 33140 8667 33144 8675
rect 33164 8667 33168 8675
rect 33172 8667 33184 8675
rect 33188 8667 33200 8675
rect 33204 8667 33208 8675
rect 33224 8667 33240 8675
rect 33256 8667 33272 8675
rect 33280 8667 33304 8675
rect 33320 8667 33368 8675
rect 33384 8667 33388 8675
rect 33392 8667 33396 8675
rect 33416 8667 33420 8675
rect 33424 8667 33436 8675
rect 33448 8667 33452 8675
rect 33456 8667 33460 8675
rect 33572 8667 33576 8675
rect 33580 8667 33584 8675
rect 33632 8667 33636 8675
rect 33640 8667 33644 8675
rect 33664 8667 33668 8675
rect 33672 8667 33676 8675
rect 33688 8667 33700 8675
rect 33704 8667 33708 8675
rect 33728 8667 33732 8675
rect 33736 8667 33740 8675
rect 33752 8667 33764 8675
rect 33768 8667 33780 8675
rect 33792 8667 33796 8675
rect 33800 8667 33804 8675
rect 33932 8667 33936 8675
rect 33940 8667 33944 8675
rect 34236 8667 34248 8675
rect 34252 8667 34264 8675
rect 34268 8667 34280 8675
rect 34300 8667 34312 8675
rect 34324 8667 34328 8675
rect 34332 8667 34344 8675
rect 34456 8667 34468 8675
rect 34548 8667 34560 8675
rect 34580 8667 34592 8675
rect 34596 8667 34600 8675
rect 34612 8667 34624 8675
rect 34640 8667 34656 8675
rect 34664 8667 34696 8675
rect 34712 8667 34716 8675
rect 34720 8667 34724 8675
rect 34736 8667 34748 8675
rect 34752 8667 34764 8675
rect 34776 8667 34780 8675
rect 34784 8667 34788 8675
rect 34804 8667 34820 8675
rect 34828 8667 34840 8675
rect 34844 8667 34856 8675
rect 34868 8667 34872 8675
rect 34876 8667 34880 8675
rect 34896 8667 34912 8675
rect 34920 8667 34936 8675
rect 34952 8667 34968 8675
rect 34984 8667 35000 8675
rect 35008 8667 35024 8675
rect 35040 8667 35044 8675
rect 35048 8667 35052 8675
rect 35064 8667 35076 8675
rect 35084 8667 35108 8675
rect 35124 8667 35136 8675
rect 35140 8667 35144 8675
rect 35160 8667 35184 8675
rect 35200 8667 35224 8675
rect 35240 8667 35256 8675
rect 35272 8667 35284 8675
rect 35296 8667 35300 8675
rect 35304 8667 35316 8675
rect 35320 8667 35324 8675
rect 35344 8667 35348 8675
rect 35352 8667 35356 8675
rect 35388 8667 35392 8675
rect 35396 8667 35408 8675
rect 35428 8667 35440 8675
rect 35444 8667 35448 8675
rect 35464 8667 35468 8675
rect 35472 8667 35484 8675
rect 35496 8667 35500 8675
rect 35504 8667 35508 8675
rect 35520 8667 35532 8675
rect 35536 8667 35540 8675
rect 35636 8667 35640 8675
rect 35644 8667 35648 8675
rect 35660 8667 35672 8675
rect 35676 8667 35688 8675
rect 35700 8667 35704 8675
rect 35708 8667 35712 8675
rect 35808 8667 35812 8675
rect 35816 8667 35828 8675
rect 35840 8667 35844 8675
rect 35848 8667 35852 8675
rect 35864 8667 35876 8675
rect 35880 8667 35884 8675
rect 35948 8667 35952 8675
rect 35956 8667 35960 8675
rect 35980 8667 35984 8675
rect 35988 8667 35992 8675
rect 36004 8667 36016 8675
rect 36020 8667 36032 8675
rect 36044 8667 36048 8675
rect 36052 8667 36056 8675
rect 36072 8667 36076 8675
rect 36080 8667 36084 8675
rect 36096 8667 36108 8675
rect 36112 8667 36124 8675
rect 36136 8667 36140 8675
rect 36144 8667 36148 8675
rect 36160 8667 36172 8675
rect 36176 8667 36188 8675
rect 36200 8667 36204 8675
rect 36208 8667 36212 8675
rect 36308 8667 36312 8675
rect 36316 8667 36328 8675
rect 36340 8667 36344 8675
rect 36348 8667 36352 8675
rect 36364 8667 36376 8675
rect 36388 8667 36392 8675
rect 36396 8667 36408 8675
rect 36412 8667 36416 8675
rect 36428 8667 36440 8675
rect 36452 8667 36456 8675
rect 36460 8667 36472 8675
rect 36488 8667 36512 8675
rect 36520 8667 36536 8675
rect 36552 8667 36568 8675
rect 36584 8667 36588 8675
rect 36592 8667 36604 8675
rect 36608 8667 36620 8675
rect 36624 8667 36628 8675
rect 36740 8667 36744 8675
rect 36748 8667 36760 8675
rect 36764 8667 36776 8675
rect 36780 8667 36784 8675
rect 36804 8667 36808 8675
rect 36812 8667 36816 8675
rect 36912 8667 36916 8675
rect 36920 8667 36932 8675
rect 36936 8667 36948 8675
rect 36952 8667 36956 8675
rect 37068 8667 37072 8675
rect 37076 8667 37080 8675
rect 37176 8667 37180 8675
rect 37184 8667 37188 8675
rect 37200 8667 37212 8675
rect 37216 8667 37220 8675
rect 37240 8667 37244 8675
rect 37248 8667 37260 8675
rect 37272 8667 37276 8675
rect 37280 8667 37284 8675
rect 37304 8667 37308 8675
rect 37312 8667 37324 8675
rect 37336 8667 37340 8675
rect 37344 8667 37348 8675
rect 37396 8667 37400 8675
rect 37404 8667 37416 8675
rect 37428 8667 37432 8675
rect 37436 8667 37440 8675
rect 37452 8667 37464 8675
rect 37468 8667 37480 8675
rect 37492 8667 37496 8675
rect 37500 8667 37504 8675
rect 37520 8667 37536 8675
rect 37544 8667 37556 8675
rect 37560 8667 37572 8675
rect 37584 8667 37588 8675
rect 37592 8667 37596 8675
rect 37612 8667 37628 8675
rect 37636 8667 37660 8675
rect 37676 8667 37692 8675
rect 37708 8667 37720 8675
rect 37724 8667 37736 8675
rect 37740 8667 37752 8675
rect 37772 8667 37784 8675
rect 37928 8667 37940 8675
rect 37960 8667 37972 8675
rect 37976 8667 37988 8675
rect 37992 8667 38004 8675
rect 38020 8667 38036 8675
rect 38044 8667 38076 8675
rect 38084 8667 38100 8675
rect 38116 8667 38120 8675
rect 38124 8667 38128 8675
rect 38148 8667 38152 8675
rect 38156 8667 38168 8675
rect 38180 8667 38184 8675
rect 38188 8667 38192 8675
rect 38352 8667 38356 8675
rect 38360 8667 38364 8675
rect 38384 8667 38388 8675
rect 38392 8667 38396 8675
rect 38408 8667 38420 8675
rect 38424 8667 38436 8675
rect 38444 8667 38460 8675
rect 38476 8667 38480 8675
rect 38484 8667 38488 8675
rect 38500 8667 38512 8675
rect 38516 8667 38528 8675
rect 38540 8667 38544 8675
rect 38548 8667 38552 8675
rect 38568 8667 38584 8675
rect 38592 8667 38616 8675
rect 38632 8667 38644 8675
rect 38664 8667 38676 8675
rect 38680 8667 38692 8675
rect 38696 8667 38708 8675
rect 38820 8667 38832 8675
rect 38852 8667 38864 8675
rect 38868 8667 38872 8675
rect 38884 8667 38896 8675
rect 38908 8667 38912 8675
rect 38916 8667 38928 8675
rect 38932 8667 38936 8675
rect 39072 8667 39084 8675
rect 39088 8667 39100 8675
rect 39104 8667 39116 8675
rect 39132 8667 39144 8675
rect 39164 8667 39176 8675
rect 39180 8667 39192 8675
rect 39196 8667 39208 8675
rect 39256 8667 39268 8675
rect 39272 8667 39284 8675
rect 39288 8667 39300 8675
rect 39476 8667 39488 8675
rect 39500 8667 39504 8675
rect 39508 8667 39520 8675
rect 39524 8667 39528 8675
rect 39540 8667 39552 8675
rect 39564 8667 39568 8675
rect 39572 8667 39584 8675
rect 39600 8667 39648 8675
rect 39664 8667 39676 8675
rect 39696 8667 39708 8675
rect 39720 8667 39724 8675
rect 39728 8667 39740 8675
rect 39812 8667 39816 8675
rect 39820 8667 39832 8675
rect 39852 8667 39864 8675
rect 39868 8667 39872 8675
rect 39976 8667 39988 8675
rect 39992 8667 39996 8675
rect 30480 8657 30488 8665
rect 33920 8657 33928 8665
rect 33952 8657 33960 8665
rect 31296 8637 31304 8645
rect 31424 8637 31432 8645
rect 31728 8637 31736 8645
rect 32368 8637 32376 8645
rect 34272 8637 34280 8645
rect 34528 8637 34536 8645
rect 35008 8637 35016 8645
rect 35024 8637 35032 8645
rect 36240 8637 36248 8645
rect 36512 8637 36520 8645
rect 36656 8637 36664 8645
rect 38096 8637 38104 8645
rect 39088 8637 39096 8645
rect 39312 8637 39320 8645
rect 31904 8617 31912 8625
rect 32592 8617 32600 8625
rect 36400 8617 36408 8625
rect 36496 8617 36504 8625
rect 29376 8597 29384 8605
rect 29920 8597 29928 8605
rect 31200 8597 31208 8605
rect 33360 8597 33368 8605
rect 33424 8597 33432 8605
rect 33936 8597 33944 8605
rect 34016 8597 34024 8605
rect 34352 8597 34360 8605
rect 34672 8597 34680 8605
rect 34720 8597 34728 8605
rect 35312 8597 35320 8605
rect 35584 8597 35592 8605
rect 35696 8597 35704 8605
rect 36016 8597 36024 8605
rect 37040 8597 37048 8605
rect 37744 8597 37752 8605
rect 37888 8597 37896 8605
rect 38112 8597 38120 8605
rect 38368 8597 38376 8605
rect 39168 8597 39176 8605
rect 39696 8597 39704 8605
rect 30208 8577 30216 8585
rect 30304 8577 30312 8585
rect 31600 8577 31608 8585
rect 33264 8577 33272 8585
rect 33376 8577 33384 8585
rect 34288 8577 34296 8585
rect 34336 8577 34344 8585
rect 35008 8577 35016 8585
rect 36096 8577 36104 8585
rect 36240 8577 36248 8585
rect 36816 8577 36824 8585
rect 37856 8577 37864 8585
rect 38128 8577 38136 8585
rect 29392 8557 29400 8565
rect 29840 8557 29848 8565
rect 29936 8557 29944 8565
rect 32112 8557 32120 8565
rect 32240 8557 32248 8565
rect 32720 8557 32728 8565
rect 33392 8557 33400 8565
rect 34992 8557 35000 8565
rect 35104 8557 35112 8565
rect 35744 8557 35752 8565
rect 35984 8557 35992 8565
rect 39040 8557 39048 8565
rect 39840 8557 39848 8565
rect 30768 8537 30776 8545
rect 36976 8537 36984 8545
rect 37072 8517 37080 8525
rect 37088 8517 37096 8525
rect 29396 8467 29408 8475
rect 29464 8467 29468 8475
rect 29472 8467 29476 8475
rect 29540 8467 29544 8475
rect 29548 8467 29560 8475
rect 29648 8467 29652 8475
rect 29656 8467 29660 8475
rect 29724 8467 29728 8475
rect 29732 8467 29744 8475
rect 29748 8467 29752 8475
rect 29772 8467 29776 8475
rect 29780 8467 29792 8475
rect 29800 8467 29816 8475
rect 29824 8467 29840 8475
rect 29856 8467 29868 8475
rect 29876 8467 29908 8475
rect 29916 8467 29932 8475
rect 29940 8467 29964 8475
rect 29980 8467 29984 8475
rect 29988 8467 30000 8475
rect 30012 8467 30016 8475
rect 30020 8467 30024 8475
rect 30044 8467 30048 8475
rect 30052 8467 30064 8475
rect 30136 8467 30140 8475
rect 30144 8467 30148 8475
rect 30228 8467 30232 8475
rect 30236 8467 30240 8475
rect 30260 8467 30264 8475
rect 30268 8467 30280 8475
rect 30284 8467 30288 8475
rect 30300 8467 30312 8475
rect 30328 8467 30340 8475
rect 30352 8467 30356 8475
rect 30360 8467 30364 8475
rect 30412 8467 30416 8475
rect 30420 8467 30432 8475
rect 30444 8467 30448 8475
rect 30452 8467 30456 8475
rect 30468 8467 30480 8475
rect 30484 8467 30496 8475
rect 30504 8467 30520 8475
rect 30536 8467 30584 8475
rect 30600 8467 30612 8475
rect 30632 8467 30644 8475
rect 30656 8467 30660 8475
rect 30664 8467 30676 8475
rect 30860 8467 30864 8475
rect 30868 8467 30880 8475
rect 30884 8467 30896 8475
rect 30916 8467 30928 8475
rect 30932 8467 30936 8475
rect 31072 8467 31084 8475
rect 31088 8467 31092 8475
rect 31112 8467 31116 8475
rect 31120 8467 31132 8475
rect 31144 8467 31148 8475
rect 31152 8467 31156 8475
rect 31176 8467 31180 8475
rect 31184 8467 31196 8475
rect 31208 8467 31212 8475
rect 31216 8467 31220 8475
rect 31232 8467 31244 8475
rect 31284 8467 31288 8475
rect 31292 8467 31304 8475
rect 31308 8467 31312 8475
rect 31332 8467 31336 8475
rect 31340 8467 31344 8475
rect 31364 8467 31368 8475
rect 31372 8467 31376 8475
rect 31396 8467 31400 8475
rect 31404 8467 31408 8475
rect 31428 8467 31432 8475
rect 31436 8467 31448 8475
rect 31452 8467 31464 8475
rect 31468 8467 31472 8475
rect 31488 8467 31492 8475
rect 31496 8467 31500 8475
rect 31520 8467 31524 8475
rect 31528 8467 31540 8475
rect 31544 8467 31548 8475
rect 31564 8467 31580 8475
rect 31596 8467 31600 8475
rect 31604 8467 31616 8475
rect 31620 8467 31624 8475
rect 31640 8467 31664 8475
rect 31680 8467 31704 8475
rect 31720 8467 31732 8475
rect 31752 8467 31764 8475
rect 31776 8467 31780 8475
rect 31784 8467 31788 8475
rect 31800 8467 31812 8475
rect 31816 8467 31820 8475
rect 31836 8467 31840 8475
rect 31844 8467 31856 8475
rect 31868 8467 31872 8475
rect 31876 8467 31880 8475
rect 31892 8467 31904 8475
rect 31908 8467 31920 8475
rect 31932 8467 31936 8475
rect 31940 8467 31944 8475
rect 31956 8467 31968 8475
rect 31972 8467 31976 8475
rect 31996 8467 32000 8475
rect 32004 8467 32008 8475
rect 32024 8467 32040 8475
rect 32048 8467 32080 8475
rect 32088 8467 32104 8475
rect 32112 8467 32124 8475
rect 32128 8467 32132 8475
rect 32148 8467 32172 8475
rect 32188 8467 32200 8475
rect 32204 8467 32208 8475
rect 32220 8467 32232 8475
rect 32244 8467 32248 8475
rect 32252 8467 32256 8475
rect 32272 8467 32276 8475
rect 32280 8467 32284 8475
rect 32296 8467 32308 8475
rect 32312 8467 32324 8475
rect 32336 8467 32340 8475
rect 32344 8467 32348 8475
rect 32360 8467 32372 8475
rect 32376 8467 32388 8475
rect 32400 8467 32404 8475
rect 32408 8467 32412 8475
rect 32432 8467 32436 8475
rect 32440 8467 32444 8475
rect 32464 8467 32468 8475
rect 32472 8467 32476 8475
rect 32496 8467 32500 8475
rect 32504 8467 32508 8475
rect 32520 8467 32532 8475
rect 32536 8467 32548 8475
rect 32560 8467 32564 8475
rect 32568 8467 32572 8475
rect 32652 8467 32656 8475
rect 32660 8467 32664 8475
rect 32676 8467 32688 8475
rect 32692 8467 32696 8475
rect 32716 8467 32720 8475
rect 32724 8467 32728 8475
rect 32744 8467 32760 8475
rect 32768 8467 32800 8475
rect 32808 8467 32824 8475
rect 32840 8467 32864 8475
rect 32872 8467 32888 8475
rect 32904 8467 32908 8475
rect 32912 8467 32916 8475
rect 32928 8467 32940 8475
rect 32944 8467 32956 8475
rect 32964 8467 32980 8475
rect 32996 8467 33044 8475
rect 33060 8467 33084 8475
rect 33092 8467 33104 8475
rect 33116 8467 33120 8475
rect 33124 8467 33136 8475
rect 33152 8467 33200 8475
rect 33216 8467 33232 8475
rect 33248 8467 33264 8475
rect 33280 8467 33296 8475
rect 33312 8467 33360 8475
rect 33376 8467 33388 8475
rect 33392 8467 33396 8475
rect 33408 8467 33420 8475
rect 33428 8467 33452 8475
rect 33468 8467 33480 8475
rect 33484 8467 33488 8475
rect 33504 8467 33528 8475
rect 33536 8467 33552 8475
rect 33560 8467 33576 8475
rect 33588 8467 33600 8475
rect 33612 8467 33644 8475
rect 33660 8467 33676 8475
rect 33692 8467 33704 8475
rect 33716 8467 33720 8475
rect 33724 8467 33728 8475
rect 33748 8467 33752 8475
rect 33756 8467 33760 8475
rect 34072 8467 34076 8475
rect 34080 8467 34084 8475
rect 34096 8467 34108 8475
rect 34112 8467 34124 8475
rect 34136 8467 34140 8475
rect 34144 8467 34148 8475
rect 34228 8467 34232 8475
rect 34236 8467 34240 8475
rect 34252 8467 34264 8475
rect 34268 8467 34272 8475
rect 34368 8467 34372 8475
rect 34376 8467 34380 8475
rect 34392 8467 34404 8475
rect 34408 8467 34420 8475
rect 34432 8467 34436 8475
rect 34440 8467 34444 8475
rect 34460 8467 34476 8475
rect 34484 8467 34496 8475
rect 34500 8467 34512 8475
rect 34520 8467 34536 8475
rect 34552 8467 34556 8475
rect 34560 8467 34564 8475
rect 34576 8467 34588 8475
rect 34592 8467 34604 8475
rect 34616 8467 34620 8475
rect 34624 8467 34628 8475
rect 34644 8467 34648 8475
rect 34652 8467 34656 8475
rect 34668 8467 34680 8475
rect 34684 8467 34696 8475
rect 34716 8467 34728 8475
rect 34740 8467 34744 8475
rect 34748 8467 34760 8475
rect 34780 8467 34792 8475
rect 34904 8467 34916 8475
rect 34920 8467 34924 8475
rect 34944 8467 34948 8475
rect 34952 8467 34956 8475
rect 34976 8467 34980 8475
rect 34984 8467 34996 8475
rect 35016 8467 35028 8475
rect 35048 8467 35060 8475
rect 35064 8467 35068 8475
rect 35084 8467 35100 8475
rect 35116 8467 35148 8475
rect 35164 8467 35176 8475
rect 35180 8467 35184 8475
rect 35204 8467 35208 8475
rect 35212 8467 35224 8475
rect 35228 8467 35232 8475
rect 35252 8467 35256 8475
rect 35260 8467 35264 8475
rect 35280 8467 35284 8475
rect 35288 8467 35300 8475
rect 35304 8467 35316 8475
rect 35336 8467 35348 8475
rect 35452 8467 35456 8475
rect 35460 8467 35472 8475
rect 35476 8467 35480 8475
rect 35492 8467 35504 8475
rect 35544 8467 35548 8475
rect 35552 8467 35556 8475
rect 35568 8467 35580 8475
rect 35584 8467 35596 8475
rect 35608 8467 35612 8475
rect 35616 8467 35620 8475
rect 35636 8467 35640 8475
rect 35644 8467 35648 8475
rect 35660 8467 35672 8475
rect 35676 8467 35688 8475
rect 35896 8467 35908 8475
rect 35912 8467 35924 8475
rect 35928 8467 35940 8475
rect 35956 8467 35968 8475
rect 35988 8467 36000 8475
rect 36004 8467 36016 8475
rect 36020 8467 36024 8475
rect 36044 8467 36048 8475
rect 36052 8467 36056 8475
rect 36072 8467 36088 8475
rect 36096 8467 36120 8475
rect 36136 8467 36184 8475
rect 36200 8467 36216 8475
rect 36232 8467 36248 8475
rect 36264 8467 36280 8475
rect 36296 8467 36344 8475
rect 36360 8467 36364 8475
rect 36368 8467 36372 8475
rect 36384 8467 36396 8475
rect 36400 8467 36412 8475
rect 36432 8467 36444 8475
rect 36448 8467 36452 8475
rect 36464 8467 36476 8475
rect 36496 8467 36508 8475
rect 36528 8467 36540 8475
rect 36552 8467 36556 8475
rect 36560 8467 36572 8475
rect 36592 8467 36604 8475
rect 36608 8467 36612 8475
rect 36740 8467 36744 8475
rect 36748 8467 36752 8475
rect 36764 8467 36776 8475
rect 36780 8467 36792 8475
rect 36804 8467 36808 8475
rect 36812 8467 36816 8475
rect 36836 8467 36840 8475
rect 36844 8467 36848 8475
rect 36960 8467 36964 8475
rect 36968 8467 36972 8475
rect 36992 8467 36996 8475
rect 37000 8467 37004 8475
rect 37016 8467 37028 8475
rect 37032 8467 37044 8475
rect 37056 8467 37060 8475
rect 37064 8467 37068 8475
rect 37084 8467 37088 8475
rect 37092 8467 37096 8475
rect 37108 8467 37120 8475
rect 37124 8467 37136 8475
rect 37148 8467 37152 8475
rect 37156 8467 37160 8475
rect 37176 8467 37224 8475
rect 37240 8467 37244 8475
rect 37248 8467 37252 8475
rect 37272 8467 37276 8475
rect 37280 8467 37292 8475
rect 37304 8467 37308 8475
rect 37312 8467 37316 8475
rect 37396 8467 37400 8475
rect 37404 8467 37408 8475
rect 37428 8467 37432 8475
rect 37436 8467 37440 8475
rect 37520 8467 37524 8475
rect 37528 8467 37540 8475
rect 37544 8467 37556 8475
rect 37560 8467 37564 8475
rect 37584 8467 37588 8475
rect 37592 8467 37596 8475
rect 37612 8467 37628 8475
rect 37636 8467 37660 8475
rect 37676 8467 37700 8475
rect 37708 8467 37720 8475
rect 37732 8467 37736 8475
rect 37740 8467 37752 8475
rect 37768 8467 37792 8475
rect 37800 8467 37812 8475
rect 37820 8467 37844 8475
rect 37860 8467 37884 8475
rect 37892 8467 37908 8475
rect 37924 8467 37948 8475
rect 37956 8467 37972 8475
rect 37980 8467 38004 8475
rect 38020 8467 38036 8475
rect 38044 8467 38068 8475
rect 38084 8467 38108 8475
rect 38116 8467 38132 8475
rect 38148 8467 38164 8475
rect 38180 8467 38184 8475
rect 38188 8467 38200 8475
rect 38204 8467 38216 8475
rect 38220 8467 38224 8475
rect 38244 8467 38248 8475
rect 38252 8467 38264 8475
rect 38268 8467 38280 8475
rect 38284 8467 38288 8475
rect 38384 8467 38388 8475
rect 38392 8467 38396 8475
rect 38416 8467 38420 8475
rect 38424 8467 38436 8475
rect 38440 8467 38452 8475
rect 38456 8467 38460 8475
rect 38508 8467 38512 8475
rect 38516 8467 38528 8475
rect 38532 8467 38544 8475
rect 38548 8467 38552 8475
rect 38572 8467 38576 8475
rect 38580 8467 38584 8475
rect 38600 8467 38616 8475
rect 38624 8467 38648 8475
rect 38664 8467 38688 8475
rect 38696 8467 38708 8475
rect 38720 8467 38724 8475
rect 38728 8467 38740 8475
rect 38744 8467 38748 8475
rect 38760 8467 38772 8475
rect 38792 8467 38804 8475
rect 38824 8467 38836 8475
rect 38856 8467 38868 8475
rect 38880 8467 38884 8475
rect 38888 8467 38900 8475
rect 38904 8467 38908 8475
rect 38920 8467 38932 8475
rect 38940 8467 38964 8475
rect 38980 8467 38992 8475
rect 38996 8467 39000 8475
rect 39012 8467 39024 8475
rect 39036 8467 39040 8475
rect 39044 8467 39056 8475
rect 39072 8467 39084 8475
rect 39088 8467 39092 8475
rect 39104 8467 39116 8475
rect 39124 8467 39148 8475
rect 39164 8467 39176 8475
rect 39180 8467 39184 8475
rect 39200 8467 39208 8475
rect 39220 8467 39224 8475
rect 39228 8467 39240 8475
rect 39256 8467 39280 8475
rect 39288 8467 39304 8475
rect 39320 8467 39336 8475
rect 39352 8467 39368 8475
rect 39376 8467 39400 8475
rect 39416 8467 39428 8475
rect 39432 8467 39436 8475
rect 39448 8467 39460 8475
rect 39472 8467 39476 8475
rect 39480 8467 39492 8475
rect 39496 8467 39500 8475
rect 39628 8467 39632 8475
rect 39636 8467 39648 8475
rect 39652 8467 39656 8475
rect 39760 8467 39772 8475
rect 39792 8467 39804 8475
rect 39808 8467 39812 8475
rect 39824 8467 39836 8475
rect 39856 8467 39868 8475
rect 39876 8467 39908 8475
rect 39916 8467 39932 8475
rect 39940 8467 39964 8475
rect 39980 8467 39984 8475
rect 39988 8467 40000 8475
rect 31472 8457 31480 8465
rect 32336 8437 32344 8445
rect 37392 8437 37400 8445
rect 30864 8417 30872 8425
rect 31856 8417 31864 8425
rect 29680 8377 29688 8385
rect 29872 8377 29880 8385
rect 30656 8377 30664 8385
rect 30704 8377 30712 8385
rect 30832 8377 30840 8385
rect 32128 8377 32136 8385
rect 32208 8377 32216 8385
rect 32528 8377 32536 8385
rect 32912 8377 32920 8385
rect 33120 8377 33128 8385
rect 34384 8377 34392 8385
rect 34432 8377 34440 8385
rect 34512 8377 34520 8385
rect 35008 8377 35016 8385
rect 35488 8377 35496 8385
rect 35648 8377 35656 8385
rect 37248 8377 37256 8385
rect 38256 8377 38264 8385
rect 38304 8377 38312 8385
rect 38560 8377 38568 8385
rect 38944 8377 38952 8385
rect 39184 8377 39192 8385
rect 39456 8377 39464 8385
rect 29712 8357 29720 8365
rect 30048 8357 30056 8365
rect 31040 8357 31048 8365
rect 34720 8357 34728 8365
rect 35056 8357 35064 8365
rect 35328 8357 35336 8365
rect 35472 8357 35480 8365
rect 35520 8357 35528 8365
rect 35840 8357 35848 8365
rect 38800 8357 38808 8365
rect 29696 8337 29704 8345
rect 31520 8337 31528 8345
rect 32224 8337 32232 8345
rect 32608 8337 32616 8345
rect 33088 8337 33096 8345
rect 34048 8337 34056 8345
rect 35824 8337 35832 8345
rect 36560 8337 36568 8345
rect 36768 8337 36776 8345
rect 37264 8337 37272 8345
rect 38080 8337 38088 8345
rect 38464 8337 38472 8345
rect 38544 8337 38552 8345
rect 39008 8337 39016 8345
rect 39200 8337 39208 8345
rect 39632 8337 39640 8345
rect 29856 8317 29864 8325
rect 37984 8317 37992 8325
rect 38832 8317 38840 8325
rect 39264 8317 39272 8325
rect 39328 8317 39336 8325
rect 39664 8317 39672 8325
rect 39760 8317 39768 8325
rect 32472 8311 32480 8313
rect 32466 8305 32480 8311
rect 30192 8297 30200 8305
rect 30368 8297 30376 8305
rect 30656 8297 30664 8305
rect 31616 8297 31624 8305
rect 31936 8297 31944 8305
rect 32064 8297 32072 8305
rect 32464 8297 32472 8305
rect 35120 8297 35128 8305
rect 35184 8297 35192 8305
rect 35616 8297 35624 8305
rect 36304 8297 36312 8305
rect 36640 8297 36648 8305
rect 37184 8297 37192 8305
rect 37600 8297 37608 8305
rect 38032 8297 38040 8305
rect 38688 8297 38696 8305
rect 38784 8297 38792 8305
rect 39120 8297 39128 8305
rect 39376 8297 39384 8305
rect 36208 8277 36216 8285
rect 39440 8277 39448 8285
rect 29396 8267 29408 8275
rect 29428 8267 29440 8275
rect 29444 8267 29448 8275
rect 29460 8267 29472 8275
rect 29488 8267 29504 8275
rect 29512 8267 29544 8275
rect 29552 8267 29568 8275
rect 29584 8267 29588 8275
rect 29592 8267 29596 8275
rect 29616 8267 29620 8275
rect 29624 8267 29636 8275
rect 29648 8267 29652 8275
rect 29656 8267 29660 8275
rect 29852 8267 29856 8275
rect 29860 8267 29864 8275
rect 29960 8267 29964 8275
rect 29968 8267 29972 8275
rect 29992 8267 29996 8275
rect 30000 8267 30004 8275
rect 30016 8267 30028 8275
rect 30032 8267 30036 8275
rect 30052 8267 30068 8275
rect 30084 8267 30132 8275
rect 30148 8267 30152 8275
rect 30156 8267 30160 8275
rect 30180 8267 30184 8275
rect 30188 8267 30200 8275
rect 30212 8267 30216 8275
rect 30220 8267 30224 8275
rect 30304 8267 30308 8275
rect 30312 8267 30316 8275
rect 30412 8267 30416 8275
rect 30420 8267 30432 8275
rect 30444 8267 30448 8275
rect 30452 8267 30456 8275
rect 30468 8267 30480 8275
rect 30484 8267 30488 8275
rect 30504 8267 30520 8275
rect 30536 8267 30552 8275
rect 30560 8267 30592 8275
rect 30600 8267 30612 8275
rect 30628 8267 30644 8275
rect 30652 8267 30684 8275
rect 30700 8267 30704 8275
rect 30708 8267 30712 8275
rect 30732 8267 30736 8275
rect 30740 8267 30752 8275
rect 30772 8267 30784 8275
rect 30796 8267 30800 8275
rect 30804 8267 30816 8275
rect 30820 8267 30824 8275
rect 30840 8267 30856 8275
rect 30872 8267 30876 8275
rect 30880 8267 30892 8275
rect 30896 8267 30900 8275
rect 30916 8267 30940 8275
rect 30948 8267 30964 8275
rect 30972 8267 30988 8275
rect 30996 8267 31020 8275
rect 31036 8267 31040 8275
rect 31044 8267 31056 8275
rect 31072 8267 31096 8275
rect 31112 8267 31116 8275
rect 31120 8267 31132 8275
rect 31152 8267 31164 8275
rect 31284 8267 31288 8275
rect 31292 8267 31296 8275
rect 31400 8267 31412 8275
rect 31432 8267 31444 8275
rect 31448 8267 31460 8275
rect 31472 8267 31476 8275
rect 31480 8267 31484 8275
rect 31572 8267 31584 8275
rect 31596 8267 31600 8275
rect 31604 8267 31608 8275
rect 31620 8267 31632 8275
rect 31640 8267 31656 8275
rect 31672 8267 31688 8275
rect 31696 8267 31708 8275
rect 31716 8267 31732 8275
rect 31748 8267 31764 8275
rect 31772 8267 31784 8275
rect 31796 8267 31800 8275
rect 31804 8267 31808 8275
rect 31824 8267 31840 8275
rect 31848 8267 31872 8275
rect 31888 8267 31904 8275
rect 31912 8267 31944 8275
rect 31960 8267 31976 8275
rect 31984 8267 32000 8275
rect 32024 8267 32036 8275
rect 32056 8267 32068 8275
rect 32072 8267 32084 8275
rect 32088 8267 32092 8275
rect 32108 8267 32124 8275
rect 32140 8267 32156 8275
rect 32164 8267 32180 8275
rect 32196 8267 32200 8275
rect 32204 8267 32208 8275
rect 32220 8267 32232 8275
rect 32240 8267 32256 8275
rect 32272 8267 32276 8275
rect 32280 8267 32284 8275
rect 32296 8267 32308 8275
rect 32312 8267 32324 8275
rect 32336 8267 32340 8275
rect 32344 8267 32348 8275
rect 32364 8267 32412 8275
rect 32428 8267 32444 8275
rect 32460 8267 32472 8275
rect 32484 8267 32488 8275
rect 32492 8267 32504 8275
rect 32524 8267 32536 8275
rect 32540 8267 32544 8275
rect 32576 8267 32580 8275
rect 32584 8267 32596 8275
rect 32616 8267 32628 8275
rect 32632 8267 32636 8275
rect 32740 8267 32752 8275
rect 32756 8267 32760 8275
rect 32772 8267 32784 8275
rect 32800 8267 32816 8275
rect 32832 8267 32880 8275
rect 32896 8267 32908 8275
rect 32928 8267 32940 8275
rect 32952 8267 32956 8275
rect 32960 8267 32972 8275
rect 32992 8267 33004 8275
rect 33008 8267 33020 8275
rect 33024 8267 33036 8275
rect 33056 8267 33068 8275
rect 33076 8267 33108 8275
rect 33116 8267 33132 8275
rect 33148 8267 33160 8275
rect 33168 8267 33200 8275
rect 33208 8267 33224 8275
rect 33240 8267 33256 8275
rect 33272 8267 33288 8275
rect 33304 8267 33320 8275
rect 33328 8267 33360 8275
rect 33368 8267 33384 8275
rect 33392 8267 33416 8275
rect 33428 8267 33452 8275
rect 33468 8267 33492 8275
rect 33508 8267 33520 8275
rect 33540 8267 33552 8275
rect 33564 8267 33568 8275
rect 33572 8267 33576 8275
rect 33616 8267 33628 8275
rect 33640 8267 33644 8275
rect 33648 8267 33652 8275
rect 33664 8267 33676 8275
rect 33772 8267 33784 8275
rect 33788 8267 33792 8275
rect 33808 8267 33824 8275
rect 33840 8267 33888 8275
rect 33904 8267 33920 8275
rect 33932 8267 33980 8275
rect 33996 8267 34000 8275
rect 34004 8267 34008 8275
rect 34028 8267 34032 8275
rect 34036 8267 34048 8275
rect 34060 8267 34064 8275
rect 34068 8267 34072 8275
rect 34152 8267 34156 8275
rect 34160 8267 34164 8275
rect 34184 8267 34188 8275
rect 34192 8267 34196 8275
rect 34276 8267 34280 8275
rect 34284 8267 34288 8275
rect 34300 8267 34312 8275
rect 34316 8267 34320 8275
rect 34340 8267 34344 8275
rect 34348 8267 34352 8275
rect 34368 8267 34416 8275
rect 34432 8267 34448 8275
rect 34464 8267 34476 8275
rect 34488 8267 34492 8275
rect 34496 8267 34508 8275
rect 34652 8267 34664 8275
rect 34668 8267 34672 8275
rect 34808 8267 34820 8275
rect 34832 8267 34836 8275
rect 34840 8267 34852 8275
rect 34856 8267 34860 8275
rect 34872 8267 34884 8275
rect 34900 8267 34916 8275
rect 34932 8267 34956 8275
rect 34964 8267 34980 8275
rect 34988 8267 35004 8275
rect 35012 8267 35036 8275
rect 35052 8267 35064 8275
rect 35084 8267 35096 8275
rect 35108 8267 35112 8275
rect 35116 8267 35128 8275
rect 35132 8267 35136 8275
rect 35216 8267 35220 8275
rect 35224 8267 35236 8275
rect 35256 8267 35268 8275
rect 35272 8267 35276 8275
rect 35332 8267 35344 8275
rect 35348 8267 35352 8275
rect 35368 8267 35384 8275
rect 35400 8267 35416 8275
rect 35424 8267 35440 8275
rect 35448 8267 35472 8275
rect 35488 8267 35492 8275
rect 35496 8267 35508 8275
rect 35524 8267 35536 8275
rect 35540 8267 35544 8275
rect 35564 8267 35568 8275
rect 35572 8267 35584 8275
rect 35588 8267 35592 8275
rect 35604 8267 35616 8275
rect 35624 8267 35640 8275
rect 35656 8267 35672 8275
rect 35680 8267 35696 8275
rect 35712 8267 35716 8275
rect 35720 8267 35724 8275
rect 35744 8267 35748 8275
rect 35752 8267 35764 8275
rect 35768 8267 35780 8275
rect 35796 8267 35812 8275
rect 35828 8267 35852 8275
rect 35868 8267 35880 8275
rect 35900 8267 35912 8275
rect 35916 8267 35928 8275
rect 35932 8267 35936 8275
rect 35952 8267 35968 8275
rect 35984 8267 35988 8275
rect 35992 8267 36004 8275
rect 36008 8267 36012 8275
rect 36032 8267 36036 8275
rect 36040 8267 36044 8275
rect 36132 8267 36144 8275
rect 36148 8267 36160 8275
rect 36164 8267 36176 8275
rect 36196 8267 36208 8275
rect 36224 8267 36248 8275
rect 36256 8267 36272 8275
rect 36288 8267 36336 8275
rect 36348 8267 36364 8275
rect 36380 8267 36412 8275
rect 36428 8267 36444 8275
rect 36460 8267 36464 8275
rect 36468 8267 36480 8275
rect 36568 8267 36572 8275
rect 36576 8267 36580 8275
rect 36600 8267 36604 8275
rect 36608 8267 36612 8275
rect 36676 8267 36680 8275
rect 36684 8267 36688 8275
rect 36700 8267 36712 8275
rect 36728 8267 36744 8275
rect 36760 8267 36792 8275
rect 36800 8267 36816 8275
rect 36832 8267 36844 8275
rect 36852 8267 36884 8275
rect 36892 8267 36908 8275
rect 36916 8267 36932 8275
rect 36948 8267 36972 8275
rect 36980 8267 36996 8275
rect 37012 8267 37028 8275
rect 37036 8267 37048 8275
rect 37052 8267 37064 8275
rect 37072 8267 37088 8275
rect 37104 8267 37120 8275
rect 37128 8267 37152 8275
rect 37168 8267 37184 8275
rect 37192 8267 37224 8275
rect 37232 8267 37244 8275
rect 37260 8267 37276 8275
rect 37284 8267 37316 8275
rect 37324 8267 37336 8275
rect 37356 8267 37368 8275
rect 37376 8267 37408 8275
rect 37416 8267 37432 8275
rect 37448 8267 37460 8275
rect 37468 8267 37500 8275
rect 37508 8267 37524 8275
rect 37532 8267 37556 8275
rect 37572 8267 37576 8275
rect 37580 8267 37592 8275
rect 37604 8267 37608 8275
rect 37612 8267 37616 8275
rect 37636 8267 37640 8275
rect 37644 8267 37656 8275
rect 37668 8267 37672 8275
rect 37676 8267 37680 8275
rect 37692 8267 37704 8275
rect 37708 8267 37712 8275
rect 37732 8267 37736 8275
rect 37740 8267 37744 8275
rect 37760 8267 37776 8275
rect 37784 8267 37816 8275
rect 37824 8267 37836 8275
rect 37856 8267 37868 8275
rect 37876 8267 37908 8275
rect 37916 8267 37932 8275
rect 37940 8267 37964 8275
rect 37980 8267 37984 8275
rect 37988 8267 38000 8275
rect 38012 8267 38016 8275
rect 38020 8267 38024 8275
rect 38152 8267 38156 8275
rect 38160 8267 38164 8275
rect 38292 8267 38296 8275
rect 38300 8267 38304 8275
rect 38324 8267 38328 8275
rect 38332 8267 38344 8275
rect 38348 8267 38360 8275
rect 38364 8267 38368 8275
rect 38384 8267 38400 8275
rect 38416 8267 38432 8275
rect 38440 8267 38452 8275
rect 38456 8267 38460 8275
rect 38480 8267 38484 8275
rect 38488 8267 38500 8275
rect 38508 8267 38524 8275
rect 38532 8267 38556 8275
rect 38572 8267 38588 8275
rect 38604 8267 38616 8275
rect 38628 8267 38632 8275
rect 38636 8267 38648 8275
rect 38652 8267 38656 8275
rect 38668 8267 38680 8275
rect 38720 8267 38724 8275
rect 38728 8267 38740 8275
rect 38744 8267 38748 8275
rect 38760 8267 38772 8275
rect 38792 8267 38804 8275
rect 38820 8267 38844 8275
rect 38852 8267 38868 8275
rect 38876 8267 38900 8275
rect 38916 8267 38932 8275
rect 38940 8267 38964 8275
rect 38980 8267 38992 8275
rect 38996 8267 39000 8275
rect 39012 8267 39024 8275
rect 39036 8267 39040 8275
rect 39044 8267 39056 8275
rect 39060 8267 39064 8275
rect 39128 8267 39132 8275
rect 39136 8267 39148 8275
rect 39152 8267 39156 8275
rect 39200 8267 39208 8275
rect 39220 8267 39224 8275
rect 39228 8267 39240 8275
rect 39244 8267 39248 8275
rect 39260 8267 39272 8275
rect 39292 8267 39304 8275
rect 39320 8267 39344 8275
rect 39352 8267 39368 8275
rect 39376 8267 39400 8275
rect 39416 8267 39428 8275
rect 39448 8267 39460 8275
rect 39472 8267 39476 8275
rect 39480 8267 39492 8275
rect 39496 8267 39500 8275
rect 39696 8267 39708 8275
rect 39720 8267 39724 8275
rect 39728 8267 39740 8275
rect 39744 8267 39748 8275
rect 39760 8267 39772 8275
rect 39788 8267 39804 8275
rect 39820 8267 39844 8275
rect 39852 8267 39868 8275
rect 39876 8267 39900 8275
rect 39916 8267 39920 8275
rect 39924 8267 39936 8275
rect 39940 8267 39952 8275
rect 39956 8267 39960 8275
rect 39980 8267 39984 8275
rect 39988 8267 39992 8275
rect 35200 8257 35208 8265
rect 35280 8257 35288 8265
rect 37520 8257 37528 8265
rect 37888 8257 37896 8265
rect 30735 8238 30742 8243
rect 31536 8237 31544 8245
rect 34448 8237 34456 8245
rect 34720 8237 34728 8245
rect 34848 8237 34856 8245
rect 29920 8217 29928 8225
rect 30384 8217 30392 8225
rect 30576 8217 30584 8225
rect 30896 8217 30904 8225
rect 31376 8217 31384 8225
rect 31984 8217 31992 8225
rect 32096 8217 32104 8225
rect 33360 8217 33368 8225
rect 33424 8217 33432 8225
rect 33568 8217 33576 8225
rect 33696 8217 33704 8225
rect 33792 8217 33800 8225
rect 34272 8217 34280 8225
rect 35840 8217 35848 8225
rect 36128 8217 36136 8225
rect 36912 8217 36920 8225
rect 38288 8217 38296 8225
rect 38384 8217 38392 8225
rect 30976 8197 30984 8205
rect 31056 8197 31064 8205
rect 31200 8197 31208 8205
rect 31248 8197 31256 8205
rect 32064 8197 32072 8205
rect 32496 8197 32504 8205
rect 32688 8197 32696 8205
rect 33136 8197 33144 8205
rect 33472 8197 33480 8205
rect 33648 8197 33656 8205
rect 34144 8197 34152 8205
rect 35472 8197 35480 8205
rect 35552 8197 35560 8205
rect 35920 8197 35928 8205
rect 37296 8197 37304 8205
rect 37504 8197 37512 8205
rect 37920 8197 37928 8205
rect 38912 8197 38920 8205
rect 39072 8197 39080 8205
rect 39584 8197 39592 8205
rect 39920 8197 39928 8205
rect 29600 8177 29608 8185
rect 32224 8177 32232 8185
rect 33136 8177 33144 8185
rect 33168 8177 33176 8185
rect 33664 8177 33672 8185
rect 35088 8177 35096 8185
rect 35472 8177 35480 8185
rect 35504 8177 35512 8185
rect 37696 8177 37704 8185
rect 38880 8177 38888 8185
rect 30656 8157 30664 8165
rect 30992 8157 31000 8165
rect 31360 8157 31368 8165
rect 31408 8157 31416 8165
rect 31728 8157 31736 8165
rect 32704 8157 32712 8165
rect 33632 8157 33640 8165
rect 34000 8157 34008 8165
rect 34912 8157 34920 8165
rect 36096 8157 36104 8165
rect 38048 8157 38056 8165
rect 38128 8157 38136 8165
rect 39360 8157 39368 8165
rect 39968 8157 39976 8165
rect 30176 8137 30184 8145
rect 29396 8067 29408 8075
rect 29428 8067 29440 8075
rect 29444 8067 29448 8075
rect 29460 8067 29472 8075
rect 29492 8067 29504 8075
rect 29516 8067 29520 8075
rect 29524 8067 29536 8075
rect 29556 8067 29568 8075
rect 29588 8067 29600 8075
rect 29604 8067 29608 8075
rect 29620 8067 29632 8075
rect 29652 8067 29664 8075
rect 29668 8067 29680 8075
rect 29684 8067 29696 8075
rect 29712 8067 29728 8075
rect 29744 8067 29768 8075
rect 29776 8067 29792 8075
rect 29808 8067 29824 8075
rect 29832 8067 29856 8075
rect 29872 8067 29884 8075
rect 29904 8067 29916 8075
rect 29920 8067 29932 8075
rect 29936 8067 29948 8075
rect 30060 8067 30072 8075
rect 30092 8067 30104 8075
rect 30108 8067 30112 8075
rect 30124 8067 30136 8075
rect 30148 8067 30152 8075
rect 30156 8067 30168 8075
rect 30312 8067 30324 8075
rect 30344 8067 30356 8075
rect 30360 8067 30364 8075
rect 30376 8067 30388 8075
rect 30400 8067 30404 8075
rect 30408 8067 30420 8075
rect 30424 8067 30428 8075
rect 30440 8067 30452 8075
rect 30472 8067 30484 8075
rect 30504 8067 30516 8075
rect 30536 8067 30548 8075
rect 30560 8067 30564 8075
rect 30568 8067 30580 8075
rect 30584 8067 30588 8075
rect 30600 8067 30612 8075
rect 30628 8067 30644 8075
rect 30660 8067 30684 8075
rect 30700 8067 30724 8075
rect 30732 8067 30748 8075
rect 30764 8067 30788 8075
rect 30804 8067 30816 8075
rect 30820 8067 30824 8075
rect 30840 8067 30864 8075
rect 30880 8067 30912 8075
rect 30928 8067 30932 8075
rect 30936 8067 30940 8075
rect 30960 8067 30964 8075
rect 30968 8067 30980 8075
rect 31000 8067 31012 8075
rect 31100 8067 31104 8075
rect 31108 8067 31112 8075
rect 31124 8067 31136 8075
rect 31156 8067 31168 8075
rect 31184 8067 31200 8075
rect 31224 8067 31256 8075
rect 31272 8067 31288 8075
rect 31300 8067 31332 8075
rect 31348 8067 31364 8075
rect 31372 8067 31384 8075
rect 31392 8067 31408 8075
rect 31424 8067 31440 8075
rect 31448 8067 31464 8075
rect 31480 8067 31496 8075
rect 31512 8067 31528 8075
rect 31536 8067 31552 8075
rect 31568 8067 31600 8075
rect 31616 8067 31620 8075
rect 31624 8067 31628 8075
rect 31640 8067 31652 8075
rect 31664 8067 31668 8075
rect 31672 8067 31676 8075
rect 31692 8067 31708 8075
rect 31716 8067 31728 8075
rect 31740 8067 31744 8075
rect 31748 8067 31752 8075
rect 31768 8067 31800 8075
rect 31816 8067 31832 8075
rect 31848 8067 31864 8075
rect 31880 8067 31896 8075
rect 31912 8067 31944 8075
rect 31960 8067 31976 8075
rect 31984 8067 31996 8075
rect 32000 8067 32012 8075
rect 32028 8067 32044 8075
rect 32060 8067 32072 8075
rect 32076 8067 32088 8075
rect 32100 8067 32104 8075
rect 32108 8067 32112 8075
rect 32340 8067 32352 8075
rect 32356 8067 32360 8075
rect 32464 8067 32476 8075
rect 32480 8067 32484 8075
rect 32496 8067 32508 8075
rect 32520 8067 32524 8075
rect 32528 8067 32540 8075
rect 32556 8067 32580 8075
rect 32588 8067 32604 8075
rect 32620 8067 32636 8075
rect 32652 8067 32656 8075
rect 32660 8067 32672 8075
rect 32676 8067 32688 8075
rect 32692 8067 32696 8075
rect 32716 8067 32720 8075
rect 32724 8067 32728 8075
rect 32792 8067 32796 8075
rect 32800 8067 32804 8075
rect 33076 8067 33080 8075
rect 33084 8067 33088 8075
rect 33100 8067 33112 8075
rect 33116 8067 33120 8075
rect 33140 8067 33144 8075
rect 33148 8067 33152 8075
rect 33168 8067 33184 8075
rect 33192 8067 33224 8075
rect 33232 8067 33248 8075
rect 33264 8067 33280 8075
rect 33296 8067 33312 8075
rect 33328 8067 33344 8075
rect 33352 8067 33384 8075
rect 33392 8067 33408 8075
rect 33420 8067 33436 8075
rect 33444 8067 33460 8075
rect 33468 8067 33492 8075
rect 33508 8067 33524 8075
rect 33540 8067 33552 8075
rect 33564 8067 33568 8075
rect 33572 8067 33584 8075
rect 33588 8067 33592 8075
rect 33608 8067 33624 8075
rect 33640 8067 33656 8075
rect 33664 8067 33680 8075
rect 33696 8067 33728 8075
rect 33736 8067 33752 8075
rect 33768 8067 33792 8075
rect 33800 8067 33816 8075
rect 33832 8067 33848 8075
rect 33856 8067 33868 8075
rect 33872 8067 33884 8075
rect 33896 8067 33900 8075
rect 33904 8067 33908 8075
rect 33924 8067 33972 8075
rect 33988 8067 34000 8075
rect 34016 8067 34064 8075
rect 34080 8067 34092 8075
rect 34108 8067 34156 8075
rect 34172 8067 34188 8075
rect 34200 8067 34248 8075
rect 34264 8067 34280 8075
rect 34296 8067 34300 8075
rect 34304 8067 34316 8075
rect 34328 8067 34332 8075
rect 34336 8067 34340 8075
rect 34360 8067 34364 8075
rect 34368 8067 34372 8075
rect 34468 8067 34472 8075
rect 34476 8067 34480 8075
rect 34492 8067 34504 8075
rect 34508 8067 34512 8075
rect 34528 8067 34552 8075
rect 34560 8067 34576 8075
rect 34584 8067 34616 8075
rect 34624 8067 34640 8075
rect 34656 8067 34672 8075
rect 34688 8067 34692 8075
rect 34696 8067 34708 8075
rect 34720 8067 34724 8075
rect 34728 8067 34732 8075
rect 34744 8067 34756 8075
rect 34760 8067 34772 8075
rect 34780 8067 34796 8075
rect 34812 8067 34816 8075
rect 34820 8067 34824 8075
rect 34836 8067 34848 8075
rect 34856 8067 34880 8075
rect 34896 8067 34908 8075
rect 34912 8067 34916 8075
rect 34936 8067 34940 8075
rect 34944 8067 34956 8075
rect 34964 8067 34980 8075
rect 34988 8067 35004 8075
rect 35012 8067 35044 8075
rect 35052 8067 35064 8075
rect 35084 8067 35096 8075
rect 35104 8067 35136 8075
rect 35152 8067 35156 8075
rect 35160 8067 35164 8075
rect 35180 8067 35212 8075
rect 35228 8067 35232 8075
rect 35236 8067 35240 8075
rect 35256 8067 35288 8075
rect 35304 8067 35320 8075
rect 35328 8067 35340 8075
rect 35344 8067 35356 8075
rect 35404 8067 35416 8075
rect 35420 8067 35432 8075
rect 35452 8067 35464 8075
rect 35480 8067 35492 8075
rect 35496 8067 35508 8075
rect 35788 8067 35792 8075
rect 35796 8067 35800 8075
rect 35820 8067 35824 8075
rect 35828 8067 35840 8075
rect 35844 8067 35848 8075
rect 35864 8067 35888 8075
rect 35896 8067 35912 8075
rect 35920 8067 35936 8075
rect 35952 8067 35968 8075
rect 35984 8067 35988 8075
rect 35992 8067 36000 8075
rect 36024 8067 36036 8075
rect 36040 8067 36044 8075
rect 36124 8067 36128 8075
rect 36132 8067 36136 8075
rect 36216 8067 36220 8075
rect 36224 8067 36228 8075
rect 36240 8067 36252 8075
rect 36256 8067 36268 8075
rect 36280 8067 36284 8075
rect 36288 8067 36292 8075
rect 36304 8067 36316 8075
rect 36320 8067 36324 8075
rect 36340 8067 36356 8075
rect 36372 8067 36388 8075
rect 36396 8067 36412 8075
rect 36420 8067 36444 8075
rect 36460 8067 36464 8075
rect 36468 8067 36480 8075
rect 36484 8067 36488 8075
rect 36552 8067 36556 8075
rect 36560 8067 36564 8075
rect 36652 8067 36664 8075
rect 36668 8067 36672 8075
rect 36720 8067 36724 8075
rect 36728 8067 36732 8075
rect 36920 8067 36924 8075
rect 36928 8067 36932 8075
rect 36944 8067 36956 8075
rect 36960 8067 36972 8075
rect 36984 8067 36988 8075
rect 36992 8067 36996 8075
rect 37012 8067 37028 8075
rect 37036 8067 37048 8075
rect 37052 8067 37064 8075
rect 37076 8067 37080 8075
rect 37084 8067 37088 8075
rect 37100 8067 37112 8075
rect 37116 8067 37120 8075
rect 37140 8067 37144 8075
rect 37148 8067 37152 8075
rect 37164 8067 37176 8075
rect 37180 8067 37184 8075
rect 37204 8067 37208 8075
rect 37212 8067 37224 8075
rect 37232 8067 37248 8075
rect 37256 8067 37268 8075
rect 37272 8067 37276 8075
rect 37296 8067 37300 8075
rect 37304 8067 37316 8075
rect 37328 8067 37332 8075
rect 37336 8067 37340 8075
rect 37360 8067 37364 8075
rect 37368 8067 37372 8075
rect 37468 8067 37472 8075
rect 37476 8067 37488 8075
rect 37492 8067 37504 8075
rect 37508 8067 37512 8075
rect 37560 8067 37564 8075
rect 37568 8067 37580 8075
rect 37584 8067 37596 8075
rect 37600 8067 37604 8075
rect 37624 8067 37628 8075
rect 37632 8067 37644 8075
rect 37648 8067 37660 8075
rect 37664 8067 37668 8075
rect 37688 8067 37692 8075
rect 37696 8067 37700 8075
rect 37720 8067 37724 8075
rect 37728 8067 37732 8075
rect 37752 8067 37756 8075
rect 37760 8067 37764 8075
rect 37784 8067 37788 8075
rect 37792 8067 37804 8075
rect 37808 8067 37820 8075
rect 37824 8067 37828 8075
rect 37848 8067 37852 8075
rect 37856 8067 37860 8075
rect 37876 8067 37892 8075
rect 37900 8067 37924 8075
rect 37940 8067 37964 8075
rect 37972 8067 37984 8075
rect 37996 8067 38000 8075
rect 38004 8067 38016 8075
rect 38032 8067 38044 8075
rect 38048 8067 38052 8075
rect 38064 8067 38076 8075
rect 38088 8067 38092 8075
rect 38096 8067 38108 8075
rect 38128 8067 38140 8075
rect 38404 8067 38408 8075
rect 38412 8067 38424 8075
rect 38728 8067 38740 8075
rect 38744 8067 38748 8075
rect 38760 8067 38772 8075
rect 38784 8067 38788 8075
rect 38792 8067 38804 8075
rect 38820 8067 38832 8075
rect 38836 8067 38840 8075
rect 38852 8067 38864 8075
rect 38876 8067 38880 8075
rect 38884 8067 38896 8075
rect 39136 8067 39148 8075
rect 39152 8067 39156 8075
rect 39168 8067 39180 8075
rect 39188 8067 39212 8075
rect 39228 8067 39252 8075
rect 39260 8067 39272 8075
rect 39284 8067 39288 8075
rect 39292 8067 39304 8075
rect 39320 8067 39344 8075
rect 39352 8067 39364 8075
rect 39376 8067 39380 8075
rect 39384 8067 39396 8075
rect 39416 8067 39428 8075
rect 39628 8067 39632 8075
rect 39636 8067 39648 8075
rect 39652 8067 39656 8075
rect 39668 8067 39680 8075
rect 39688 8067 39712 8075
rect 39728 8067 39752 8075
rect 39760 8067 39776 8075
rect 39792 8067 39796 8075
rect 39800 8067 39804 8075
rect 39824 8067 39828 8075
rect 39832 8067 39844 8075
rect 39848 8067 39860 8075
rect 39864 8067 39868 8075
rect 39888 8067 39892 8075
rect 39896 8067 39900 8075
rect 39948 8067 39952 8075
rect 39956 8067 39960 8075
rect 39980 8067 39984 8075
rect 39988 8067 39992 8075
rect 30512 8057 30520 8065
rect 33312 8057 33320 8065
rect 36480 8037 36488 8045
rect 31984 8017 31992 8025
rect 32208 8017 32216 8025
rect 35072 8017 35080 8025
rect 36112 8017 36120 8025
rect 36864 8017 36872 8025
rect 37104 8017 37112 8025
rect 38784 8017 38792 8025
rect 31728 7997 31736 8005
rect 34688 7997 34696 8005
rect 34752 7997 34760 8005
rect 37792 7997 37800 8005
rect 30208 7977 30216 7985
rect 31264 7977 31272 7985
rect 32304 7977 32312 7985
rect 32832 7977 32840 7985
rect 33488 7977 33496 7985
rect 33648 7977 33656 7985
rect 34064 7977 34072 7985
rect 35488 7977 35496 7985
rect 38064 7977 38072 7985
rect 38832 7977 38840 7985
rect 39408 7977 39416 7985
rect 40128 7977 40136 7985
rect 40752 7977 40760 7985
rect 29680 7957 29688 7965
rect 29840 7957 29848 7965
rect 30320 7957 30328 7965
rect 30480 7957 30488 7965
rect 33008 7957 33016 7965
rect 33040 7957 33048 7965
rect 39968 7957 39976 7965
rect 29424 7937 29432 7945
rect 30992 7937 31000 7945
rect 31248 7937 31256 7945
rect 31312 7937 31320 7945
rect 32464 7937 32472 7945
rect 32624 7937 32632 7945
rect 33808 7937 33816 7945
rect 35344 7937 35352 7945
rect 35616 7937 35624 7945
rect 35952 7937 35960 7945
rect 36176 7937 36184 7945
rect 36592 7937 36600 7945
rect 36688 7937 36696 7945
rect 36960 7937 36968 7945
rect 37040 7937 37048 7945
rect 37184 7937 37192 7945
rect 37552 7937 37560 7945
rect 38560 7937 38568 7945
rect 38848 7937 38856 7945
rect 38944 7937 38952 7945
rect 39200 7937 39208 7945
rect 39296 7937 39304 7945
rect 39520 7937 39528 7945
rect 40416 7937 40424 7945
rect 40512 7937 40520 7945
rect 40736 7937 40744 7945
rect 29520 7917 29528 7925
rect 29584 7917 29592 7925
rect 29840 7917 29848 7925
rect 29904 7917 29912 7925
rect 30624 7917 30632 7925
rect 30704 7917 30712 7925
rect 31296 7917 31304 7925
rect 31584 7917 31592 7925
rect 32768 7917 32776 7925
rect 33952 7917 33960 7925
rect 34512 7917 34520 7925
rect 39504 7917 39512 7925
rect 39904 7917 39912 7925
rect 33600 7897 33608 7905
rect 33680 7897 33688 7905
rect 37120 7897 37128 7905
rect 39632 7897 39640 7905
rect 33408 7877 33416 7885
rect 33712 7877 33720 7885
rect 34400 7877 34408 7885
rect 36336 7877 36344 7885
rect 36352 7877 36360 7885
rect 36368 7877 36376 7885
rect 37680 7877 37688 7885
rect 39856 7877 39864 7885
rect 29396 7867 29408 7875
rect 29428 7867 29440 7875
rect 29444 7867 29448 7875
rect 29460 7867 29472 7875
rect 29492 7867 29504 7875
rect 29516 7867 29520 7875
rect 29524 7867 29536 7875
rect 29648 7867 29660 7875
rect 29672 7867 29676 7875
rect 29680 7867 29692 7875
rect 29696 7867 29700 7875
rect 29740 7867 29752 7875
rect 29764 7867 29768 7875
rect 29772 7867 29784 7875
rect 29788 7867 29792 7875
rect 29804 7867 29816 7875
rect 29832 7867 29848 7875
rect 29864 7867 29888 7875
rect 29896 7867 29912 7875
rect 29920 7867 29932 7875
rect 29936 7867 29940 7875
rect 29960 7867 29964 7875
rect 29968 7867 29980 7875
rect 29984 7867 29996 7875
rect 30000 7867 30004 7875
rect 30100 7867 30104 7875
rect 30108 7867 30112 7875
rect 30132 7867 30136 7875
rect 30140 7867 30152 7875
rect 30156 7867 30168 7875
rect 30172 7867 30176 7875
rect 30320 7867 30324 7875
rect 30328 7867 30332 7875
rect 30352 7867 30356 7875
rect 30360 7867 30364 7875
rect 30376 7867 30388 7875
rect 30392 7867 30400 7875
rect 30412 7867 30428 7875
rect 30444 7867 30460 7875
rect 30468 7867 30492 7875
rect 30508 7867 30520 7875
rect 30540 7867 30552 7875
rect 30556 7867 30568 7875
rect 30572 7867 30584 7875
rect 30604 7867 30616 7875
rect 30696 7867 30708 7875
rect 30720 7867 30724 7875
rect 30728 7867 30740 7875
rect 30744 7867 30748 7875
rect 30760 7867 30772 7875
rect 30780 7867 30796 7875
rect 30812 7867 30816 7875
rect 30820 7867 30824 7875
rect 30836 7867 30848 7875
rect 30852 7867 30864 7875
rect 30884 7867 30896 7875
rect 30904 7867 30920 7875
rect 30928 7867 30952 7875
rect 30968 7867 30980 7875
rect 31000 7867 31012 7875
rect 31024 7867 31028 7875
rect 31032 7867 31044 7875
rect 31048 7867 31052 7875
rect 31156 7867 31168 7875
rect 31188 7867 31200 7875
rect 31204 7867 31208 7875
rect 31224 7867 31248 7875
rect 31264 7867 31288 7875
rect 31300 7867 31324 7875
rect 31340 7867 31364 7875
rect 31376 7867 31400 7875
rect 31416 7867 31440 7875
rect 31456 7867 31468 7875
rect 31488 7867 31500 7875
rect 31512 7867 31516 7875
rect 31520 7867 31524 7875
rect 31712 7867 31716 7875
rect 31720 7867 31724 7875
rect 31736 7867 31748 7875
rect 31768 7867 31780 7875
rect 31784 7867 31788 7875
rect 31808 7867 31812 7875
rect 31816 7867 31820 7875
rect 31840 7867 31844 7875
rect 31848 7867 31860 7875
rect 31880 7867 31892 7875
rect 31904 7867 31908 7875
rect 31912 7867 31916 7875
rect 31980 7867 31984 7875
rect 31988 7867 31992 7875
rect 32056 7867 32060 7875
rect 32064 7867 32068 7875
rect 32080 7867 32092 7875
rect 32096 7867 32108 7875
rect 32124 7867 32140 7875
rect 32156 7867 32168 7875
rect 32172 7867 32184 7875
rect 32188 7867 32192 7875
rect 32212 7867 32216 7875
rect 32220 7867 32224 7875
rect 32240 7867 32256 7875
rect 32264 7867 32288 7875
rect 32304 7867 32328 7875
rect 32344 7867 32348 7875
rect 32352 7867 32364 7875
rect 32372 7867 32388 7875
rect 32396 7867 32412 7875
rect 32428 7867 32432 7875
rect 32436 7867 32440 7875
rect 32460 7867 32464 7875
rect 32468 7867 32480 7875
rect 32492 7867 32496 7875
rect 32500 7867 32504 7875
rect 32516 7867 32528 7875
rect 32532 7867 32536 7875
rect 32556 7867 32560 7875
rect 32564 7867 32568 7875
rect 32588 7867 32592 7875
rect 32596 7867 32600 7875
rect 32620 7867 32624 7875
rect 32628 7867 32640 7875
rect 32652 7867 32656 7875
rect 32660 7867 32664 7875
rect 32676 7867 32688 7875
rect 32692 7867 32704 7875
rect 32716 7867 32720 7875
rect 32724 7867 32728 7875
rect 32808 7867 32812 7875
rect 32816 7867 32820 7875
rect 32916 7867 32920 7875
rect 32924 7867 32928 7875
rect 32948 7867 32952 7875
rect 32956 7867 32960 7875
rect 32972 7867 32984 7875
rect 32988 7867 32992 7875
rect 33008 7867 33024 7875
rect 33040 7867 33088 7875
rect 33104 7867 33120 7875
rect 33136 7867 33148 7875
rect 33160 7867 33164 7875
rect 33168 7867 33180 7875
rect 33292 7867 33304 7875
rect 33324 7867 33336 7875
rect 33340 7867 33344 7875
rect 33356 7867 33368 7875
rect 33376 7867 33400 7875
rect 33416 7867 33428 7875
rect 33432 7867 33436 7875
rect 33448 7867 33460 7875
rect 33468 7867 33492 7875
rect 33508 7867 33532 7875
rect 33540 7867 33552 7875
rect 33560 7867 33584 7875
rect 33600 7867 33624 7875
rect 33632 7867 33648 7875
rect 33664 7867 33668 7875
rect 33672 7867 33676 7875
rect 33696 7867 33700 7875
rect 33704 7867 33716 7875
rect 33720 7867 33732 7875
rect 33736 7867 33740 7875
rect 33836 7867 33840 7875
rect 33844 7867 33848 7875
rect 33928 7867 33932 7875
rect 33936 7867 33948 7875
rect 33960 7867 33964 7875
rect 33968 7867 33972 7875
rect 33984 7867 33996 7875
rect 34000 7867 34004 7875
rect 34052 7867 34056 7875
rect 34060 7867 34064 7875
rect 34076 7867 34088 7875
rect 34092 7867 34096 7875
rect 34176 7867 34180 7875
rect 34184 7867 34188 7875
rect 34284 7867 34288 7875
rect 34292 7867 34296 7875
rect 34376 7867 34380 7875
rect 34384 7867 34388 7875
rect 34400 7867 34412 7875
rect 34416 7867 34420 7875
rect 34440 7867 34444 7875
rect 34448 7867 34452 7875
rect 34468 7867 34516 7875
rect 34532 7867 34544 7875
rect 34548 7867 34552 7875
rect 34564 7867 34576 7875
rect 34588 7867 34592 7875
rect 34596 7867 34608 7875
rect 34628 7867 34640 7875
rect 34660 7867 34672 7875
rect 34692 7867 34704 7875
rect 34708 7867 34712 7875
rect 34724 7867 34736 7875
rect 34748 7867 34752 7875
rect 34756 7867 34768 7875
rect 34784 7867 34796 7875
rect 34800 7867 34804 7875
rect 34816 7867 34828 7875
rect 34840 7867 34844 7875
rect 34848 7867 34852 7875
rect 34964 7867 34968 7875
rect 34972 7867 34976 7875
rect 34988 7867 35000 7875
rect 35020 7867 35032 7875
rect 35036 7867 35040 7875
rect 35052 7867 35064 7875
rect 35084 7867 35096 7875
rect 35104 7867 35120 7875
rect 35128 7867 35140 7875
rect 35160 7867 35172 7875
rect 35180 7867 35196 7875
rect 35204 7867 35220 7875
rect 35236 7867 35248 7875
rect 35256 7867 35272 7875
rect 35280 7867 35296 7875
rect 35312 7867 35336 7875
rect 35344 7867 35360 7875
rect 35376 7867 35392 7875
rect 35400 7867 35412 7875
rect 35416 7867 35428 7875
rect 35444 7867 35460 7875
rect 35476 7867 35488 7875
rect 35492 7867 35504 7875
rect 35524 7867 35536 7875
rect 35548 7867 35552 7875
rect 35556 7867 35560 7875
rect 35580 7867 35584 7875
rect 35588 7867 35592 7875
rect 35612 7867 35616 7875
rect 35620 7867 35624 7875
rect 35636 7867 35648 7875
rect 35664 7867 35680 7875
rect 35688 7867 35704 7875
rect 35712 7867 35728 7875
rect 35744 7867 35748 7875
rect 35752 7867 35756 7875
rect 35776 7867 35780 7875
rect 35784 7867 35796 7875
rect 35884 7867 35888 7875
rect 35892 7867 35904 7875
rect 35924 7867 35936 7875
rect 35940 7867 35944 7875
rect 35960 7867 35976 7875
rect 36016 7867 36032 7875
rect 36040 7867 36072 7875
rect 36088 7867 36112 7875
rect 36120 7867 36132 7875
rect 36140 7867 36156 7875
rect 36172 7867 36176 7875
rect 36180 7867 36184 7875
rect 36196 7867 36208 7875
rect 36212 7867 36224 7875
rect 36488 7867 36492 7875
rect 36496 7867 36508 7875
rect 36528 7867 36540 7875
rect 36544 7867 36548 7875
rect 36620 7867 36632 7875
rect 36636 7867 36640 7875
rect 36672 7867 36676 7875
rect 36680 7867 36692 7875
rect 36712 7867 36724 7875
rect 36728 7867 36732 7875
rect 36764 7867 36768 7875
rect 36772 7867 36784 7875
rect 36804 7867 36816 7875
rect 36820 7867 36824 7875
rect 36856 7867 36860 7875
rect 36864 7867 36876 7875
rect 36896 7867 36908 7875
rect 36912 7867 36916 7875
rect 37020 7867 37032 7875
rect 37036 7867 37040 7875
rect 37052 7867 37064 7875
rect 37076 7867 37080 7875
rect 37084 7867 37096 7875
rect 37100 7867 37104 7875
rect 37116 7867 37128 7875
rect 37140 7867 37144 7875
rect 37148 7867 37160 7875
rect 37164 7867 37168 7875
rect 37180 7867 37192 7875
rect 37204 7867 37208 7875
rect 37212 7867 37224 7875
rect 37240 7867 37264 7875
rect 37272 7867 37284 7875
rect 37296 7867 37300 7875
rect 37304 7867 37316 7875
rect 37336 7867 37348 7875
rect 37360 7867 37364 7875
rect 37368 7867 37380 7875
rect 37400 7867 37412 7875
rect 37416 7867 37420 7875
rect 37432 7867 37444 7875
rect 37464 7867 37476 7875
rect 37480 7867 37484 7875
rect 37496 7867 37508 7875
rect 37516 7867 37540 7875
rect 37556 7867 37568 7875
rect 37572 7867 37576 7875
rect 37588 7867 37600 7875
rect 37612 7867 37616 7875
rect 37620 7867 37632 7875
rect 37636 7867 37640 7875
rect 37652 7867 37664 7875
rect 37744 7867 37756 7875
rect 37776 7867 37788 7875
rect 37792 7867 37804 7875
rect 37808 7867 37820 7875
rect 37836 7867 37852 7875
rect 37868 7867 37892 7875
rect 37900 7867 37916 7875
rect 37932 7867 37936 7875
rect 37940 7867 37944 7875
rect 37956 7867 37968 7875
rect 37972 7867 37984 7875
rect 37996 7867 38000 7875
rect 38004 7867 38008 7875
rect 38024 7867 38028 7875
rect 38032 7867 38036 7875
rect 38048 7867 38060 7875
rect 38064 7867 38076 7875
rect 38088 7867 38092 7875
rect 38096 7867 38100 7875
rect 38228 7867 38232 7875
rect 38236 7867 38240 7875
rect 38252 7867 38264 7875
rect 38268 7867 38272 7875
rect 38288 7867 38304 7875
rect 38320 7867 38336 7875
rect 38344 7867 38376 7875
rect 38384 7867 38396 7875
rect 38412 7867 38428 7875
rect 38436 7867 38468 7875
rect 38476 7867 38488 7875
rect 38508 7867 38520 7875
rect 38532 7867 38536 7875
rect 38540 7867 38552 7875
rect 38664 7867 38676 7875
rect 38696 7867 38708 7875
rect 38712 7867 38716 7875
rect 38728 7867 38740 7875
rect 38756 7867 38772 7875
rect 38780 7867 38812 7875
rect 38820 7867 38832 7875
rect 38848 7867 38864 7875
rect 38872 7867 38904 7875
rect 38912 7867 38924 7875
rect 38944 7867 38956 7875
rect 38964 7867 38996 7875
rect 39004 7867 39020 7875
rect 39028 7867 39040 7875
rect 39044 7867 39048 7875
rect 39068 7867 39072 7875
rect 39076 7867 39088 7875
rect 39100 7867 39104 7875
rect 39108 7867 39112 7875
rect 39208 7867 39212 7875
rect 39216 7867 39220 7875
rect 39240 7867 39244 7875
rect 39248 7867 39252 7875
rect 39332 7867 39336 7875
rect 39340 7867 39344 7875
rect 39424 7867 39428 7875
rect 39432 7867 39436 7875
rect 39516 7867 39520 7875
rect 39524 7867 39528 7875
rect 39540 7867 39552 7875
rect 39556 7867 39560 7875
rect 39580 7867 39584 7875
rect 39588 7867 39592 7875
rect 39612 7867 39616 7875
rect 39620 7867 39632 7875
rect 39644 7867 39648 7875
rect 39652 7867 39656 7875
rect 39676 7867 39680 7875
rect 39684 7867 39696 7875
rect 39700 7867 39712 7875
rect 39716 7867 39720 7875
rect 39740 7867 39744 7875
rect 39748 7867 39752 7875
rect 39768 7867 39784 7875
rect 39792 7867 39816 7875
rect 39832 7867 39844 7875
rect 39848 7867 39852 7875
rect 39864 7867 39876 7875
rect 39888 7867 39892 7875
rect 39896 7867 39908 7875
rect 39912 7867 39916 7875
rect 39928 7867 39940 7875
rect 39956 7867 39968 7875
rect 39980 7867 39984 7875
rect 39988 7867 40000 7875
rect 40004 7867 40008 7875
rect 40020 7867 40032 7875
rect 40044 7867 40048 7875
rect 40052 7867 40064 7875
rect 40068 7867 40072 7875
rect 40084 7867 40096 7875
rect 40112 7867 40128 7875
rect 40144 7867 40168 7875
rect 40176 7867 40192 7875
rect 40200 7867 40212 7875
rect 40216 7867 40220 7875
rect 40236 7867 40260 7875
rect 40268 7867 40284 7875
rect 40292 7867 40316 7875
rect 40332 7867 40336 7875
rect 40340 7867 40352 7875
rect 40364 7867 40368 7875
rect 40372 7867 40376 7875
rect 40472 7867 40476 7875
rect 40480 7867 40484 7875
rect 40504 7867 40508 7875
rect 40512 7867 40516 7875
rect 40596 7867 40600 7875
rect 40604 7867 40608 7875
rect 40620 7867 40632 7875
rect 40636 7867 40640 7875
rect 40656 7867 40672 7875
rect 40688 7867 40736 7875
rect 40752 7867 40776 7875
rect 40784 7867 40796 7875
rect 32208 7857 32216 7865
rect 32256 7857 32264 7865
rect 32272 7857 32280 7865
rect 32816 7857 32824 7865
rect 37024 7857 37032 7865
rect 29792 7837 29800 7845
rect 30288 7837 30296 7845
rect 30368 7837 30376 7845
rect 30624 7837 30632 7845
rect 30656 7837 30664 7845
rect 30864 7837 30872 7845
rect 30912 7837 30920 7845
rect 30992 7837 31000 7845
rect 31200 7837 31208 7845
rect 31664 7837 31672 7845
rect 32704 7837 32712 7845
rect 34399 7838 34406 7843
rect 35360 7837 35368 7845
rect 36400 7837 36408 7845
rect 36816 7837 36824 7845
rect 37264 7837 37272 7845
rect 37472 7837 37480 7845
rect 37920 7837 37928 7845
rect 37952 7837 37960 7845
rect 38000 7837 38008 7845
rect 38256 7837 38264 7845
rect 38624 7837 38632 7845
rect 38800 7837 38808 7845
rect 39008 7837 39016 7845
rect 40112 7837 40120 7845
rect 40224 7837 40232 7845
rect 40352 7837 40360 7845
rect 40384 7837 40392 7845
rect 40768 7837 40776 7845
rect 29488 7817 29496 7825
rect 29600 7817 29608 7825
rect 34448 7817 34456 7825
rect 34512 7817 34520 7825
rect 34784 7817 34792 7825
rect 35936 7817 35944 7825
rect 36720 7817 36728 7825
rect 36992 7817 37000 7825
rect 37120 7817 37128 7825
rect 37296 7817 37304 7825
rect 38704 7817 38712 7825
rect 29776 7797 29784 7805
rect 30048 7797 30056 7805
rect 33040 7797 33048 7805
rect 33056 7797 33064 7805
rect 33136 7797 33144 7805
rect 33968 7797 33976 7805
rect 34224 7797 34232 7805
rect 36096 7797 36104 7805
rect 36144 7797 36152 7805
rect 36272 7797 36280 7805
rect 36640 7797 36648 7805
rect 37776 7797 37784 7805
rect 38416 7797 38424 7805
rect 38688 7797 38696 7805
rect 38912 7797 38920 7805
rect 39152 7797 39160 7805
rect 39360 7797 39368 7805
rect 39600 7797 39608 7805
rect 39888 7797 39896 7805
rect 40352 7797 40360 7805
rect 40784 7797 40792 7805
rect 29440 7777 29448 7785
rect 34224 7777 34232 7785
rect 34368 7777 34376 7785
rect 36016 7777 36024 7785
rect 37232 7777 37240 7785
rect 38176 7777 38184 7785
rect 39616 7777 39624 7785
rect 40624 7777 40632 7785
rect 30032 7757 30040 7765
rect 30112 7757 30120 7765
rect 30336 7757 30344 7765
rect 32848 7757 32856 7765
rect 33392 7757 33400 7765
rect 34016 7757 34024 7765
rect 37568 7757 37576 7765
rect 38496 7757 38504 7765
rect 38576 7757 38584 7765
rect 38768 7757 38776 7765
rect 38864 7757 38872 7765
rect 39040 7757 39048 7765
rect 39392 7757 39400 7765
rect 40256 7757 40264 7765
rect 36000 7737 36008 7745
rect 38032 7737 38040 7745
rect 39136 7737 39144 7745
rect 30864 7717 30872 7725
rect 31072 7717 31080 7725
rect 31168 7717 31176 7725
rect 31184 7717 31192 7725
rect 38496 7717 38504 7725
rect 30592 7697 30600 7705
rect 30800 7697 30808 7705
rect 31296 7677 31304 7685
rect 32880 7677 32888 7685
rect 29548 7667 29552 7675
rect 29556 7667 29560 7675
rect 29580 7667 29584 7675
rect 29588 7667 29592 7675
rect 29604 7667 29616 7675
rect 29620 7667 29632 7675
rect 29648 7667 29664 7675
rect 29672 7667 29704 7675
rect 29712 7667 29728 7675
rect 29736 7667 29748 7675
rect 29752 7667 29756 7675
rect 29772 7667 29796 7675
rect 29804 7667 29820 7675
rect 29828 7667 29840 7675
rect 29844 7667 29848 7675
rect 29868 7667 29872 7675
rect 29876 7667 29888 7675
rect 29900 7667 29904 7675
rect 29908 7667 29912 7675
rect 30008 7667 30012 7675
rect 30016 7667 30020 7675
rect 30040 7667 30044 7675
rect 30048 7667 30052 7675
rect 30100 7667 30104 7675
rect 30108 7667 30112 7675
rect 30132 7667 30136 7675
rect 30140 7667 30152 7675
rect 30156 7667 30168 7675
rect 30172 7667 30176 7675
rect 30196 7667 30200 7675
rect 30204 7667 30208 7675
rect 30220 7667 30232 7675
rect 30236 7667 30240 7675
rect 30260 7667 30264 7675
rect 30268 7667 30272 7675
rect 30284 7667 30296 7675
rect 30300 7667 30312 7675
rect 30320 7667 30336 7675
rect 30352 7667 30368 7675
rect 30376 7667 30388 7675
rect 30392 7667 30400 7675
rect 30412 7667 30428 7675
rect 30444 7667 30448 7675
rect 30452 7667 30456 7675
rect 30468 7667 30480 7675
rect 30484 7667 30496 7675
rect 30504 7667 30520 7675
rect 30536 7667 30540 7675
rect 30544 7667 30548 7675
rect 30560 7667 30572 7675
rect 30576 7667 30588 7675
rect 30600 7667 30604 7675
rect 30608 7667 30612 7675
rect 30628 7667 30632 7675
rect 30636 7667 30640 7675
rect 30652 7667 30664 7675
rect 30668 7667 30680 7675
rect 30688 7667 30704 7675
rect 30720 7667 30736 7675
rect 30744 7667 30756 7675
rect 30760 7667 30772 7675
rect 30780 7667 30796 7675
rect 30812 7667 30860 7675
rect 30876 7667 30880 7675
rect 30884 7667 30888 7675
rect 30904 7667 30952 7675
rect 30968 7667 30980 7675
rect 30984 7667 30988 7675
rect 31000 7667 31012 7675
rect 31024 7667 31028 7675
rect 31032 7667 31044 7675
rect 31148 7667 31152 7675
rect 31156 7667 31168 7675
rect 31224 7667 31228 7675
rect 31232 7667 31244 7675
rect 31256 7667 31260 7675
rect 31264 7667 31268 7675
rect 31280 7667 31292 7675
rect 31308 7667 31320 7675
rect 31332 7667 31336 7675
rect 31340 7667 31352 7675
rect 31356 7667 31360 7675
rect 31376 7667 31392 7675
rect 31408 7667 31412 7675
rect 31416 7667 31428 7675
rect 31432 7667 31444 7675
rect 31460 7667 31476 7675
rect 31492 7667 31516 7675
rect 31532 7667 31544 7675
rect 31564 7667 31576 7675
rect 31580 7667 31592 7675
rect 31596 7667 31600 7675
rect 31808 7667 31812 7675
rect 31816 7667 31820 7675
rect 31840 7667 31844 7675
rect 31848 7667 31860 7675
rect 31864 7667 31868 7675
rect 31884 7667 31908 7675
rect 31924 7667 31936 7675
rect 31940 7667 31944 7675
rect 31964 7667 31968 7675
rect 31972 7667 31984 7675
rect 32000 7667 32012 7675
rect 32016 7667 32020 7675
rect 32032 7667 32044 7675
rect 32052 7667 32068 7675
rect 32084 7667 32116 7675
rect 32124 7667 32140 7675
rect 32152 7667 32168 7675
rect 32176 7667 32192 7675
rect 32200 7667 32224 7675
rect 32240 7667 32256 7675
rect 32264 7667 32288 7675
rect 32304 7667 32336 7675
rect 32344 7667 32360 7675
rect 32372 7667 32388 7675
rect 32396 7667 32412 7675
rect 32420 7667 32432 7675
rect 32452 7667 32464 7675
rect 32468 7667 32480 7675
rect 32484 7667 32496 7675
rect 32516 7667 32528 7675
rect 32532 7667 32536 7675
rect 32548 7667 32560 7675
rect 32576 7667 32592 7675
rect 32608 7667 32640 7675
rect 32648 7667 32664 7675
rect 32680 7667 32692 7675
rect 32696 7667 32708 7675
rect 32712 7667 32724 7675
rect 32740 7667 32756 7675
rect 32772 7667 32796 7675
rect 32804 7667 32820 7675
rect 32836 7667 32840 7675
rect 32844 7667 32848 7675
rect 32860 7667 32872 7675
rect 32876 7667 32888 7675
rect 32900 7667 32904 7675
rect 32908 7667 32912 7675
rect 32928 7667 32932 7675
rect 32936 7667 32940 7675
rect 32952 7667 32964 7675
rect 32968 7667 32980 7675
rect 32992 7667 32996 7675
rect 33000 7667 33004 7675
rect 33020 7667 33024 7675
rect 33028 7667 33032 7675
rect 33044 7667 33056 7675
rect 33060 7667 33072 7675
rect 33084 7667 33088 7675
rect 33092 7667 33096 7675
rect 33112 7667 33128 7675
rect 33136 7667 33148 7675
rect 33152 7667 33164 7675
rect 33176 7667 33180 7675
rect 33184 7667 33188 7675
rect 33284 7667 33288 7675
rect 33292 7667 33304 7675
rect 33316 7667 33320 7675
rect 33324 7667 33328 7675
rect 33340 7667 33352 7675
rect 33356 7667 33368 7675
rect 33376 7667 33392 7675
rect 33408 7667 33412 7675
rect 33416 7667 33420 7675
rect 33432 7667 33444 7675
rect 33448 7667 33460 7675
rect 33468 7667 33484 7675
rect 33500 7667 33516 7675
rect 33524 7667 33536 7675
rect 33540 7667 33552 7675
rect 33560 7667 33576 7675
rect 33616 7667 33628 7675
rect 33632 7667 33644 7675
rect 33652 7667 33668 7675
rect 33684 7667 33700 7675
rect 33708 7667 33732 7675
rect 33748 7667 33760 7675
rect 33780 7667 33792 7675
rect 33796 7667 33808 7675
rect 33812 7667 33824 7675
rect 33936 7667 33948 7675
rect 33968 7667 33980 7675
rect 33984 7667 33988 7675
rect 34000 7667 34012 7675
rect 34024 7667 34028 7675
rect 34032 7667 34044 7675
rect 34060 7667 34072 7675
rect 34076 7667 34080 7675
rect 34092 7667 34104 7675
rect 34116 7667 34120 7675
rect 34124 7667 34136 7675
rect 34140 7667 34144 7675
rect 34156 7667 34168 7675
rect 34184 7667 34200 7675
rect 34216 7667 34240 7675
rect 34248 7667 34264 7675
rect 34272 7667 34296 7675
rect 34312 7667 34316 7675
rect 34320 7667 34332 7675
rect 34336 7667 34348 7675
rect 34352 7667 34356 7675
rect 34372 7667 34388 7675
rect 34404 7667 34420 7675
rect 34428 7667 34452 7675
rect 34468 7667 34492 7675
rect 34500 7667 34512 7675
rect 34524 7667 34528 7675
rect 34532 7667 34544 7675
rect 34548 7667 34552 7675
rect 34564 7667 34576 7675
rect 34784 7667 34796 7675
rect 34800 7667 34804 7675
rect 34816 7667 34828 7675
rect 34840 7667 34844 7675
rect 34848 7667 34860 7675
rect 34948 7667 34952 7675
rect 34956 7667 34968 7675
rect 34988 7667 35000 7675
rect 35004 7667 35008 7675
rect 35028 7667 35032 7675
rect 35036 7667 35040 7675
rect 35056 7667 35072 7675
rect 35080 7667 35096 7675
rect 35104 7667 35120 7675
rect 35128 7667 35140 7675
rect 35160 7667 35172 7675
rect 35184 7667 35188 7675
rect 35192 7667 35196 7675
rect 35216 7667 35220 7675
rect 35224 7667 35228 7675
rect 35388 7667 35392 7675
rect 35396 7667 35408 7675
rect 35412 7667 35424 7675
rect 35428 7667 35432 7675
rect 35480 7667 35484 7675
rect 35488 7667 35500 7675
rect 35504 7667 35508 7675
rect 35528 7667 35532 7675
rect 35536 7667 35540 7675
rect 35560 7667 35564 7675
rect 35568 7667 35572 7675
rect 35592 7667 35596 7675
rect 35600 7667 35604 7675
rect 35624 7667 35628 7675
rect 35632 7667 35644 7675
rect 35648 7667 35652 7675
rect 35668 7667 35672 7675
rect 35676 7667 35680 7675
rect 35700 7667 35704 7675
rect 35708 7667 35720 7675
rect 35724 7667 35728 7675
rect 35884 7667 35888 7675
rect 35892 7667 35896 7675
rect 35960 7667 35964 7675
rect 35968 7667 35980 7675
rect 36000 7667 36012 7675
rect 36016 7667 36020 7675
rect 36092 7667 36104 7675
rect 36160 7667 36164 7675
rect 36168 7667 36172 7675
rect 36192 7667 36196 7675
rect 36200 7667 36204 7675
rect 36216 7667 36228 7675
rect 36244 7667 36260 7675
rect 36276 7667 36324 7675
rect 36340 7667 36352 7675
rect 36372 7667 36384 7675
rect 36396 7667 36400 7675
rect 36404 7667 36416 7675
rect 36436 7667 36448 7675
rect 36452 7667 36464 7675
rect 36468 7667 36480 7675
rect 36496 7667 36508 7675
rect 36528 7667 36540 7675
rect 36544 7667 36556 7675
rect 36560 7667 36572 7675
rect 36592 7667 36604 7675
rect 36620 7667 36644 7675
rect 36652 7667 36668 7675
rect 36684 7667 36688 7675
rect 36692 7667 36696 7675
rect 36708 7667 36720 7675
rect 36724 7667 36736 7675
rect 36748 7667 36752 7675
rect 36756 7667 36760 7675
rect 36856 7667 36860 7675
rect 36864 7667 36868 7675
rect 36888 7667 36892 7675
rect 36896 7667 36900 7675
rect 36912 7667 36924 7675
rect 36928 7667 36940 7675
rect 36952 7667 36956 7675
rect 36960 7667 36964 7675
rect 36984 7667 36988 7675
rect 36992 7667 36996 7675
rect 37060 7667 37064 7675
rect 37068 7667 37080 7675
rect 37092 7667 37096 7675
rect 37100 7667 37104 7675
rect 37116 7667 37128 7675
rect 37132 7667 37144 7675
rect 37156 7667 37160 7675
rect 37164 7667 37168 7675
rect 37188 7667 37192 7675
rect 37196 7667 37208 7675
rect 37220 7667 37224 7675
rect 37228 7667 37232 7675
rect 37252 7667 37256 7675
rect 37260 7667 37264 7675
rect 37552 7667 37556 7675
rect 37560 7667 37572 7675
rect 37584 7667 37588 7675
rect 37592 7667 37596 7675
rect 37608 7667 37620 7675
rect 37624 7667 37628 7675
rect 37648 7667 37652 7675
rect 37656 7667 37660 7675
rect 37676 7667 37692 7675
rect 37700 7667 37732 7675
rect 37740 7667 37752 7675
rect 37772 7667 37784 7675
rect 37788 7667 37800 7675
rect 37804 7667 37816 7675
rect 37864 7667 37876 7675
rect 37880 7667 37892 7675
rect 37896 7667 37908 7675
rect 37956 7667 37968 7675
rect 37972 7667 37984 7675
rect 37988 7667 38000 7675
rect 38016 7667 38028 7675
rect 38048 7667 38060 7675
rect 38064 7667 38076 7675
rect 38080 7667 38092 7675
rect 38228 7667 38232 7675
rect 38236 7667 38248 7675
rect 38252 7667 38256 7675
rect 38268 7667 38280 7675
rect 38296 7667 38308 7675
rect 38320 7667 38324 7675
rect 38328 7667 38340 7675
rect 38344 7667 38348 7675
rect 38388 7667 38400 7675
rect 38412 7667 38416 7675
rect 38420 7667 38432 7675
rect 38436 7667 38440 7675
rect 38480 7667 38492 7675
rect 38504 7667 38508 7675
rect 38512 7667 38516 7675
rect 38528 7667 38540 7675
rect 38544 7667 38556 7675
rect 38572 7667 38588 7675
rect 38604 7667 38628 7675
rect 38636 7667 38652 7675
rect 38668 7667 38672 7675
rect 38676 7667 38680 7675
rect 38692 7667 38704 7675
rect 38712 7667 38736 7675
rect 38752 7667 38764 7675
rect 38768 7667 38772 7675
rect 38792 7667 38796 7675
rect 38800 7667 38812 7675
rect 38820 7667 38836 7675
rect 38844 7667 38856 7675
rect 38876 7667 38888 7675
rect 38900 7667 38904 7675
rect 38908 7667 38920 7675
rect 38940 7667 38952 7675
rect 39024 7667 39028 7675
rect 39032 7667 39036 7675
rect 39116 7667 39120 7675
rect 39124 7667 39128 7675
rect 39192 7667 39196 7675
rect 39200 7667 39204 7675
rect 39316 7667 39320 7675
rect 39324 7667 39328 7675
rect 39424 7667 39428 7675
rect 39432 7667 39436 7675
rect 39448 7667 39460 7675
rect 39464 7667 39468 7675
rect 39488 7667 39492 7675
rect 39496 7667 39508 7675
rect 39516 7667 39532 7675
rect 39540 7667 39572 7675
rect 39580 7667 39596 7675
rect 39612 7667 39636 7675
rect 39644 7667 39660 7675
rect 39676 7667 39724 7675
rect 39740 7667 39764 7675
rect 39772 7667 39784 7675
rect 39796 7667 39800 7675
rect 39804 7667 39816 7675
rect 40044 7667 40048 7675
rect 40052 7667 40064 7675
rect 40084 7667 40096 7675
rect 40100 7667 40104 7675
rect 40116 7667 40128 7675
rect 40144 7667 40160 7675
rect 40176 7667 40224 7675
rect 40236 7667 40252 7675
rect 40268 7667 40316 7675
rect 40332 7667 40336 7675
rect 40340 7667 40344 7675
rect 40364 7667 40368 7675
rect 40372 7667 40384 7675
rect 40396 7667 40400 7675
rect 40404 7667 40408 7675
rect 40504 7667 40508 7675
rect 40512 7667 40516 7675
rect 40756 7667 40760 7675
rect 40764 7667 40776 7675
rect 40788 7667 40792 7675
rect 40796 7667 40800 7675
rect 31104 7657 31112 7665
rect 35760 7657 35768 7665
rect 36112 7657 36120 7665
rect 37856 7657 37864 7665
rect 38416 7657 38424 7665
rect 29408 7637 29416 7645
rect 32272 7637 32280 7645
rect 37568 7637 37576 7645
rect 32464 7617 32472 7625
rect 37344 7617 37352 7625
rect 39136 7617 39144 7625
rect 39696 7617 39704 7625
rect 32896 7597 32904 7605
rect 38832 7597 38840 7605
rect 38912 7597 38920 7605
rect 30448 7577 30456 7585
rect 31824 7577 31832 7585
rect 32080 7577 32088 7585
rect 33424 7577 33432 7585
rect 33440 7577 33448 7585
rect 33488 7577 33496 7585
rect 34608 7577 34616 7585
rect 34960 7577 34968 7585
rect 35360 7577 35368 7585
rect 35696 7577 35704 7585
rect 37024 7577 37032 7585
rect 37824 7577 37832 7585
rect 38368 7577 38376 7585
rect 38464 7577 38472 7585
rect 38560 7577 38568 7585
rect 38784 7577 38792 7585
rect 39904 7577 39912 7585
rect 31552 7557 31560 7565
rect 32544 7557 32552 7565
rect 36064 7557 36072 7565
rect 36112 7557 36120 7565
rect 36208 7557 36216 7565
rect 36224 7557 36232 7565
rect 37408 7557 37416 7565
rect 38288 7557 38296 7565
rect 38656 7557 38664 7565
rect 39104 7557 39112 7565
rect 30000 7537 30008 7545
rect 31472 7537 31480 7545
rect 31680 7537 31688 7545
rect 32672 7537 32680 7545
rect 34544 7537 34552 7545
rect 35584 7537 35592 7545
rect 35840 7537 35848 7545
rect 39056 7537 39064 7545
rect 39264 7537 39272 7545
rect 40176 7537 40184 7545
rect 40544 7537 40552 7545
rect 29712 7517 29720 7525
rect 30272 7517 30280 7525
rect 30784 7517 30792 7525
rect 30976 7517 30984 7525
rect 32208 7517 32216 7525
rect 32224 7517 32232 7525
rect 33712 7517 33720 7525
rect 33776 7517 33784 7525
rect 36608 7517 36616 7525
rect 36688 7517 36696 7525
rect 37040 7517 37048 7525
rect 37120 7517 37128 7525
rect 37280 7517 37288 7525
rect 37488 7517 37496 7525
rect 37680 7517 37688 7525
rect 29728 7497 29736 7505
rect 30832 7497 30840 7505
rect 31040 7497 31048 7505
rect 31648 7497 31656 7505
rect 32432 7497 32440 7505
rect 33312 7497 33320 7505
rect 33376 7497 33384 7505
rect 33904 7497 33912 7505
rect 35184 7497 35192 7505
rect 35552 7497 35560 7505
rect 36208 7497 36216 7505
rect 37968 7497 37976 7505
rect 39616 7497 39624 7505
rect 39680 7497 39688 7505
rect 40656 7497 40664 7505
rect 32032 7477 32040 7485
rect 34304 7477 34312 7485
rect 29396 7467 29408 7475
rect 29420 7467 29424 7475
rect 29428 7467 29432 7475
rect 29444 7467 29456 7475
rect 29460 7467 29472 7475
rect 29484 7467 29488 7475
rect 29492 7467 29496 7475
rect 29508 7467 29520 7475
rect 29524 7467 29528 7475
rect 29548 7467 29552 7475
rect 29556 7467 29560 7475
rect 29572 7467 29584 7475
rect 29588 7467 29592 7475
rect 29608 7467 29632 7475
rect 29648 7467 29696 7475
rect 29712 7467 29716 7475
rect 29720 7467 29724 7475
rect 29736 7467 29748 7475
rect 29752 7467 29764 7475
rect 29772 7467 29788 7475
rect 29804 7467 29820 7475
rect 29828 7467 29840 7475
rect 29844 7467 29856 7475
rect 29868 7467 29872 7475
rect 29876 7467 29880 7475
rect 29900 7467 29904 7475
rect 29908 7467 29912 7475
rect 30008 7467 30012 7475
rect 30016 7467 30020 7475
rect 30032 7467 30044 7475
rect 30048 7467 30052 7475
rect 30068 7467 30072 7475
rect 30076 7467 30088 7475
rect 30100 7467 30104 7475
rect 30108 7467 30112 7475
rect 30124 7467 30136 7475
rect 30140 7467 30152 7475
rect 30164 7467 30168 7475
rect 30172 7467 30176 7475
rect 30188 7467 30200 7475
rect 30204 7467 30208 7475
rect 30228 7467 30232 7475
rect 30236 7467 30240 7475
rect 30260 7467 30264 7475
rect 30268 7467 30272 7475
rect 30292 7467 30296 7475
rect 30300 7467 30312 7475
rect 30324 7467 30328 7475
rect 30332 7467 30336 7475
rect 30348 7467 30360 7475
rect 30364 7467 30368 7475
rect 30432 7467 30436 7475
rect 30440 7467 30444 7475
rect 30464 7467 30468 7475
rect 30472 7467 30476 7475
rect 30524 7467 30528 7475
rect 30532 7467 30536 7475
rect 30556 7467 30560 7475
rect 30564 7467 30568 7475
rect 30580 7467 30592 7475
rect 30596 7467 30600 7475
rect 30616 7467 30632 7475
rect 30648 7467 30696 7475
rect 30712 7467 30736 7475
rect 30744 7467 30756 7475
rect 30764 7467 30788 7475
rect 30804 7467 30852 7475
rect 30868 7467 30880 7475
rect 30896 7467 30944 7475
rect 30960 7467 30976 7475
rect 30984 7467 30996 7475
rect 31000 7467 31012 7475
rect 31024 7467 31028 7475
rect 31032 7467 31036 7475
rect 31180 7467 31184 7475
rect 31188 7467 31192 7475
rect 31212 7467 31216 7475
rect 31220 7467 31224 7475
rect 31236 7467 31248 7475
rect 31252 7467 31264 7475
rect 31276 7467 31280 7475
rect 31284 7467 31288 7475
rect 31304 7467 31308 7475
rect 31312 7467 31316 7475
rect 31328 7467 31340 7475
rect 31344 7467 31356 7475
rect 31368 7467 31372 7475
rect 31376 7467 31380 7475
rect 31396 7467 31412 7475
rect 31420 7467 31432 7475
rect 31436 7467 31448 7475
rect 31460 7467 31464 7475
rect 31468 7467 31472 7475
rect 31568 7467 31572 7475
rect 31576 7467 31588 7475
rect 31600 7467 31604 7475
rect 31608 7467 31612 7475
rect 31624 7467 31636 7475
rect 31640 7467 31644 7475
rect 31664 7467 31668 7475
rect 31672 7467 31676 7475
rect 31692 7467 31708 7475
rect 31716 7467 31732 7475
rect 31740 7467 31756 7475
rect 31772 7467 31796 7475
rect 31812 7467 31824 7475
rect 31844 7467 31856 7475
rect 31860 7467 31872 7475
rect 31888 7467 31900 7475
rect 31920 7467 31932 7475
rect 31936 7467 31948 7475
rect 31952 7467 31956 7475
rect 31976 7467 31980 7475
rect 31984 7467 31988 7475
rect 32052 7467 32056 7475
rect 32060 7467 32064 7475
rect 32084 7467 32088 7475
rect 32092 7467 32104 7475
rect 32108 7467 32120 7475
rect 32124 7467 32128 7475
rect 32144 7467 32148 7475
rect 32152 7467 32156 7475
rect 32176 7467 32180 7475
rect 32184 7467 32196 7475
rect 32200 7467 32212 7475
rect 32216 7467 32220 7475
rect 32240 7467 32244 7475
rect 32248 7467 32252 7475
rect 32364 7467 32368 7475
rect 32372 7467 32376 7475
rect 32396 7467 32400 7475
rect 32404 7467 32408 7475
rect 32420 7467 32432 7475
rect 32444 7467 32448 7475
rect 32452 7467 32464 7475
rect 32468 7467 32472 7475
rect 32568 7467 32572 7475
rect 32576 7467 32588 7475
rect 32608 7467 32620 7475
rect 32624 7467 32628 7475
rect 32648 7467 32652 7475
rect 32656 7467 32660 7475
rect 32676 7467 32692 7475
rect 32700 7467 32732 7475
rect 32748 7467 32760 7475
rect 32780 7467 32792 7475
rect 32804 7467 32808 7475
rect 32812 7467 32816 7475
rect 32912 7467 32916 7475
rect 32920 7467 32924 7475
rect 33004 7467 33008 7475
rect 33012 7467 33016 7475
rect 33112 7467 33116 7475
rect 33120 7467 33124 7475
rect 33136 7467 33148 7475
rect 33152 7467 33156 7475
rect 33176 7467 33180 7475
rect 33184 7467 33188 7475
rect 33208 7467 33212 7475
rect 33216 7467 33228 7475
rect 33240 7467 33244 7475
rect 33248 7467 33252 7475
rect 33272 7467 33276 7475
rect 33280 7467 33292 7475
rect 33296 7467 33308 7475
rect 33312 7467 33316 7475
rect 33396 7467 33400 7475
rect 33404 7467 33408 7475
rect 33428 7467 33432 7475
rect 33436 7467 33440 7475
rect 33504 7467 33508 7475
rect 33512 7467 33516 7475
rect 33612 7467 33616 7475
rect 33620 7467 33624 7475
rect 33848 7467 33852 7475
rect 33856 7467 33868 7475
rect 33880 7467 33884 7475
rect 33888 7467 33892 7475
rect 33904 7467 33916 7475
rect 33920 7467 33924 7475
rect 33940 7467 33956 7475
rect 33972 7467 33988 7475
rect 33996 7467 34028 7475
rect 34036 7467 34052 7475
rect 34060 7467 34072 7475
rect 34076 7467 34080 7475
rect 34100 7467 34104 7475
rect 34108 7467 34120 7475
rect 34128 7467 34144 7475
rect 34152 7467 34176 7475
rect 34192 7467 34208 7475
rect 34224 7467 34236 7475
rect 34248 7467 34252 7475
rect 34256 7467 34268 7475
rect 34272 7467 34276 7475
rect 34288 7467 34300 7475
rect 34380 7467 34392 7475
rect 34472 7467 34484 7475
rect 34596 7467 34608 7475
rect 34612 7467 34616 7475
rect 34628 7467 34640 7475
rect 34660 7467 34672 7475
rect 34676 7467 34688 7475
rect 34692 7467 34704 7475
rect 34816 7467 34828 7475
rect 34840 7467 34844 7475
rect 34848 7467 34860 7475
rect 34864 7467 34868 7475
rect 34956 7467 34968 7475
rect 35064 7467 35076 7475
rect 35080 7467 35084 7475
rect 35104 7467 35108 7475
rect 35112 7467 35116 7475
rect 35128 7467 35140 7475
rect 35152 7467 35156 7475
rect 35160 7467 35164 7475
rect 35252 7467 35264 7475
rect 35276 7467 35280 7475
rect 35284 7467 35288 7475
rect 35300 7467 35312 7475
rect 35320 7467 35344 7475
rect 35360 7467 35384 7475
rect 35392 7467 35404 7475
rect 35416 7467 35420 7475
rect 35424 7467 35436 7475
rect 35452 7467 35476 7475
rect 35484 7467 35496 7475
rect 35508 7467 35512 7475
rect 35516 7467 35520 7475
rect 35540 7467 35544 7475
rect 35548 7467 35552 7475
rect 35572 7467 35576 7475
rect 35580 7467 35584 7475
rect 35604 7467 35608 7475
rect 35612 7467 35616 7475
rect 35628 7467 35640 7475
rect 35644 7467 35656 7475
rect 35712 7467 35716 7475
rect 35720 7467 35732 7475
rect 35752 7467 35764 7475
rect 35768 7467 35780 7475
rect 35788 7467 35804 7475
rect 35820 7467 35824 7475
rect 35828 7467 35832 7475
rect 35844 7467 35856 7475
rect 35860 7467 35872 7475
rect 35884 7467 35888 7475
rect 35892 7467 35896 7475
rect 36024 7467 36028 7475
rect 36032 7467 36036 7475
rect 36084 7467 36088 7475
rect 36092 7467 36104 7475
rect 36116 7467 36120 7475
rect 36124 7467 36128 7475
rect 36336 7467 36340 7475
rect 36344 7467 36356 7475
rect 36368 7467 36372 7475
rect 36376 7467 36380 7475
rect 36476 7467 36480 7475
rect 36484 7467 36488 7475
rect 36600 7467 36604 7475
rect 36608 7467 36612 7475
rect 36624 7467 36636 7475
rect 36640 7467 36644 7475
rect 36660 7467 36676 7475
rect 36692 7467 36740 7475
rect 36756 7467 36800 7475
rect 36820 7467 36836 7475
rect 36844 7467 36868 7475
rect 36884 7467 36896 7475
rect 36916 7467 36928 7475
rect 36932 7467 36944 7475
rect 36948 7467 36960 7475
rect 37008 7467 37020 7475
rect 37024 7467 37036 7475
rect 37040 7467 37052 7475
rect 37068 7467 37080 7475
rect 37100 7467 37112 7475
rect 37116 7467 37128 7475
rect 37132 7467 37144 7475
rect 37164 7467 37176 7475
rect 37280 7467 37284 7475
rect 37288 7467 37300 7475
rect 37304 7467 37308 7475
rect 37320 7467 37332 7475
rect 37344 7467 37348 7475
rect 37352 7467 37364 7475
rect 37380 7467 37404 7475
rect 37412 7467 37428 7475
rect 37444 7467 37460 7475
rect 37476 7467 37480 7475
rect 37484 7467 37496 7475
rect 37500 7467 37512 7475
rect 37516 7467 37520 7475
rect 37648 7467 37652 7475
rect 37656 7467 37660 7475
rect 37672 7467 37684 7475
rect 37688 7467 37692 7475
rect 37712 7467 37716 7475
rect 37720 7467 37732 7475
rect 37736 7467 37748 7475
rect 37752 7467 37756 7475
rect 37772 7467 37796 7475
rect 37804 7467 37820 7475
rect 37828 7467 37852 7475
rect 37868 7467 37872 7475
rect 37876 7467 37888 7475
rect 37900 7467 37904 7475
rect 37908 7467 37912 7475
rect 37932 7467 37936 7475
rect 37940 7467 37944 7475
rect 38008 7467 38012 7475
rect 38016 7467 38020 7475
rect 38040 7467 38044 7475
rect 38048 7467 38052 7475
rect 38116 7467 38120 7475
rect 38124 7467 38128 7475
rect 38148 7467 38152 7475
rect 38156 7467 38160 7475
rect 38172 7467 38184 7475
rect 38188 7467 38192 7475
rect 38212 7467 38216 7475
rect 38220 7467 38232 7475
rect 38236 7467 38248 7475
rect 38252 7467 38256 7475
rect 38276 7467 38280 7475
rect 38284 7467 38288 7475
rect 38352 7467 38356 7475
rect 38360 7467 38364 7475
rect 38384 7467 38388 7475
rect 38392 7467 38404 7475
rect 38408 7467 38420 7475
rect 38424 7467 38428 7475
rect 38444 7467 38460 7475
rect 38476 7467 38480 7475
rect 38484 7467 38496 7475
rect 38500 7467 38512 7475
rect 38532 7467 38544 7475
rect 38548 7467 38552 7475
rect 38572 7467 38576 7475
rect 38580 7467 38584 7475
rect 38604 7467 38608 7475
rect 38612 7467 38616 7475
rect 38636 7467 38640 7475
rect 38644 7467 38656 7475
rect 38712 7467 38716 7475
rect 38720 7467 38732 7475
rect 38752 7467 38764 7475
rect 38768 7467 38772 7475
rect 38828 7467 38840 7475
rect 38844 7467 38848 7475
rect 38912 7467 38916 7475
rect 38920 7467 38924 7475
rect 38944 7467 38948 7475
rect 38952 7467 38956 7475
rect 38968 7467 38980 7475
rect 38984 7467 38996 7475
rect 39016 7467 39028 7475
rect 39044 7467 39056 7475
rect 39060 7467 39072 7475
rect 39076 7467 39088 7475
rect 39104 7467 39120 7475
rect 39136 7467 39148 7475
rect 39152 7467 39164 7475
rect 39168 7467 39180 7475
rect 39324 7467 39336 7475
rect 39340 7467 39344 7475
rect 39608 7467 39620 7475
rect 39624 7467 39636 7475
rect 39640 7467 39652 7475
rect 39672 7467 39684 7475
rect 39692 7467 39724 7475
rect 39732 7467 39748 7475
rect 39756 7467 39788 7475
rect 39796 7467 39812 7475
rect 39828 7467 39844 7475
rect 39860 7467 39876 7475
rect 39892 7467 39908 7475
rect 39916 7467 39948 7475
rect 39956 7467 39968 7475
rect 39988 7467 40000 7475
rect 40004 7467 40016 7475
rect 40020 7467 40032 7475
rect 40048 7467 40060 7475
rect 40080 7467 40092 7475
rect 40096 7467 40108 7475
rect 40112 7467 40124 7475
rect 40236 7467 40248 7475
rect 40260 7467 40264 7475
rect 40268 7467 40280 7475
rect 40284 7467 40288 7475
rect 40300 7467 40312 7475
rect 40320 7467 40344 7475
rect 40360 7467 40384 7475
rect 40392 7467 40408 7475
rect 40424 7467 40428 7475
rect 40432 7467 40436 7475
rect 40456 7467 40460 7475
rect 40464 7467 40476 7475
rect 40480 7467 40492 7475
rect 40496 7467 40500 7475
rect 40548 7467 40552 7475
rect 40556 7467 40568 7475
rect 40572 7467 40584 7475
rect 40588 7467 40592 7475
rect 40608 7467 40624 7475
rect 40640 7467 40656 7475
rect 40664 7467 40688 7475
rect 40704 7467 40716 7475
rect 40720 7467 40724 7475
rect 40736 7467 40748 7475
rect 40756 7467 40780 7475
rect 29680 7457 29688 7465
rect 30592 7457 30600 7465
rect 35712 7457 35720 7465
rect 40016 7457 40024 7465
rect 40032 7457 40040 7465
rect 29680 7437 29688 7445
rect 29824 7437 29832 7445
rect 30752 7437 30760 7445
rect 31775 7438 31782 7443
rect 32880 7437 32888 7445
rect 33024 7437 33032 7445
rect 33440 7437 33448 7445
rect 33536 7437 33544 7445
rect 33760 7437 33768 7445
rect 34064 7437 34072 7445
rect 34512 7437 34520 7445
rect 34640 7437 34648 7445
rect 35088 7437 35096 7445
rect 35680 7437 35688 7445
rect 36112 7437 36120 7445
rect 36848 7437 36856 7445
rect 36928 7437 36936 7445
rect 37024 7437 37032 7445
rect 37744 7437 37752 7445
rect 38000 7437 38008 7445
rect 38256 7437 38264 7445
rect 39664 7437 39672 7445
rect 39776 7437 39784 7445
rect 39904 7437 39912 7445
rect 39920 7437 39928 7445
rect 40032 7437 40040 7445
rect 40336 7437 40344 7445
rect 29488 7417 29496 7425
rect 30176 7417 30184 7425
rect 30256 7417 30264 7425
rect 30336 7417 30344 7425
rect 31856 7417 31864 7425
rect 32528 7417 32536 7425
rect 32576 7417 32584 7425
rect 33232 7417 33240 7425
rect 33280 7417 33288 7425
rect 38192 7417 38200 7425
rect 38528 7417 38536 7425
rect 38576 7417 38584 7425
rect 38784 7417 38792 7425
rect 38896 7417 38904 7425
rect 39264 7417 39272 7425
rect 39360 7417 39368 7425
rect 39408 7417 39416 7425
rect 39552 7417 39560 7425
rect 29648 7397 29656 7405
rect 29776 7397 29784 7405
rect 30832 7397 30840 7405
rect 31072 7397 31080 7405
rect 33360 7397 33368 7405
rect 33376 7397 33384 7405
rect 33488 7397 33496 7405
rect 33712 7397 33720 7405
rect 34080 7397 34088 7405
rect 35280 7397 35288 7405
rect 35744 7397 35752 7405
rect 35920 7397 35928 7405
rect 36016 7397 36024 7405
rect 36176 7397 36184 7405
rect 36416 7397 36424 7405
rect 36704 7397 36712 7405
rect 36800 7397 36808 7405
rect 36912 7397 36920 7405
rect 37008 7397 37016 7405
rect 32016 7377 32024 7385
rect 32320 7377 32328 7385
rect 32368 7377 32376 7385
rect 32832 7377 32840 7385
rect 33408 7377 33416 7385
rect 37904 7377 37912 7385
rect 37968 7377 37976 7385
rect 38096 7377 38104 7385
rect 39040 7377 39048 7385
rect 39072 7377 39080 7385
rect 29408 7357 29416 7365
rect 30944 7357 30952 7365
rect 31584 7357 31592 7365
rect 32224 7357 32232 7365
rect 33520 7357 33528 7365
rect 34736 7357 34744 7365
rect 35184 7357 35192 7365
rect 35200 7357 35208 7365
rect 35808 7357 35816 7365
rect 36144 7357 36152 7365
rect 36512 7357 36520 7365
rect 37616 7357 37624 7365
rect 38032 7357 38040 7365
rect 38144 7357 38152 7365
rect 38672 7357 38680 7365
rect 38688 7357 38696 7365
rect 38928 7357 38936 7365
rect 39312 7357 39320 7365
rect 39568 7357 39576 7365
rect 36480 7337 36488 7345
rect 37104 7337 37112 7345
rect 40496 7337 40504 7345
rect 32928 7317 32936 7325
rect 33024 7317 33032 7325
rect 33056 7317 33064 7325
rect 34992 7317 35000 7325
rect 36064 7317 36072 7325
rect 36400 7317 36408 7325
rect 39856 7277 39864 7285
rect 21008 7260 21016 7268
rect 23488 7260 23496 7268
rect 23712 7260 23720 7268
rect 23904 7260 23912 7268
rect 24320 7260 24328 7268
rect 25776 7260 25784 7268
rect 27520 7260 27528 7268
rect 28048 7260 28056 7268
rect 29488 7267 29500 7275
rect 29512 7267 29516 7275
rect 29520 7267 29532 7275
rect 29536 7267 29540 7275
rect 29552 7267 29564 7275
rect 29572 7267 29596 7275
rect 29612 7267 29624 7275
rect 29628 7267 29632 7275
rect 29644 7267 29656 7275
rect 29668 7267 29672 7275
rect 29676 7267 29688 7275
rect 29704 7267 29716 7275
rect 29720 7267 29724 7275
rect 29736 7267 29748 7275
rect 29760 7267 29764 7275
rect 29768 7267 29780 7275
rect 29796 7267 29820 7275
rect 29828 7267 29840 7275
rect 29852 7267 29856 7275
rect 29860 7267 29872 7275
rect 29892 7267 29904 7275
rect 30016 7267 30028 7275
rect 30032 7267 30044 7275
rect 30048 7267 30060 7275
rect 30076 7267 30088 7275
rect 30108 7267 30120 7275
rect 30124 7267 30136 7275
rect 30140 7267 30152 7275
rect 30488 7267 30500 7275
rect 30504 7267 30508 7275
rect 30520 7267 30532 7275
rect 30544 7267 30548 7275
rect 30552 7267 30564 7275
rect 30584 7267 30596 7275
rect 30608 7267 30612 7275
rect 30616 7267 30628 7275
rect 30648 7267 30660 7275
rect 30664 7267 30676 7275
rect 30680 7267 30692 7275
rect 30764 7267 30768 7275
rect 30772 7267 30784 7275
rect 30804 7267 30816 7275
rect 30820 7267 30832 7275
rect 30836 7267 30848 7275
rect 30868 7267 30880 7275
rect 30896 7267 30908 7275
rect 30912 7267 30924 7275
rect 30928 7267 30940 7275
rect 30960 7267 30972 7275
rect 30988 7267 31012 7275
rect 31020 7267 31036 7275
rect 31052 7267 31056 7275
rect 31060 7267 31064 7275
rect 31076 7267 31088 7275
rect 31092 7267 31104 7275
rect 31116 7267 31120 7275
rect 31124 7267 31128 7275
rect 31140 7267 31152 7275
rect 31156 7267 31160 7275
rect 31176 7267 31192 7275
rect 31208 7267 31224 7275
rect 31232 7267 31264 7275
rect 31272 7267 31284 7275
rect 31300 7267 31316 7275
rect 31324 7267 31356 7275
rect 31364 7267 31380 7275
rect 31388 7267 31412 7275
rect 31424 7267 31448 7275
rect 31456 7267 31472 7275
rect 31480 7267 31492 7275
rect 31496 7267 31500 7275
rect 31516 7267 31540 7275
rect 31548 7267 31564 7275
rect 31572 7267 31584 7275
rect 31588 7267 31592 7275
rect 31612 7267 31616 7275
rect 31620 7267 31632 7275
rect 31640 7267 31656 7275
rect 31664 7267 31688 7275
rect 31704 7267 31708 7275
rect 31712 7267 31724 7275
rect 31744 7267 31756 7275
rect 31776 7267 31788 7275
rect 31808 7267 31820 7275
rect 31824 7267 31828 7275
rect 31840 7267 31852 7275
rect 31860 7267 31876 7275
rect 31892 7267 31896 7275
rect 31900 7267 31904 7275
rect 31916 7267 31928 7275
rect 31932 7267 31944 7275
rect 31952 7267 31968 7275
rect 31984 7267 32000 7275
rect 32008 7267 32024 7275
rect 32040 7267 32064 7275
rect 32080 7267 32128 7275
rect 32140 7267 32156 7275
rect 32172 7267 32220 7275
rect 32236 7267 32252 7275
rect 32264 7267 32312 7275
rect 32328 7267 32340 7275
rect 32360 7267 32372 7275
rect 32384 7267 32388 7275
rect 32392 7267 32404 7275
rect 32424 7267 32436 7275
rect 32440 7267 32452 7275
rect 32456 7267 32468 7275
rect 32484 7267 32500 7275
rect 32516 7267 32540 7275
rect 32556 7267 32572 7275
rect 32580 7267 32596 7275
rect 32604 7267 32628 7275
rect 32644 7267 32660 7275
rect 32668 7267 32684 7275
rect 32700 7267 32716 7275
rect 32724 7267 32740 7275
rect 32756 7267 32760 7275
rect 32764 7267 32768 7275
rect 32788 7267 32792 7275
rect 32796 7267 32808 7275
rect 32812 7267 32816 7275
rect 32912 7267 32916 7275
rect 32920 7267 32924 7275
rect 32944 7267 32948 7275
rect 32952 7267 32964 7275
rect 32968 7267 32980 7275
rect 32984 7267 32988 7275
rect 33004 7267 33028 7275
rect 33044 7267 33084 7275
rect 33100 7267 33116 7275
rect 33132 7267 33136 7275
rect 33140 7267 33152 7275
rect 33172 7267 33184 7275
rect 33204 7267 33216 7275
rect 33220 7267 33224 7275
rect 33236 7267 33248 7275
rect 33268 7267 33280 7275
rect 33284 7267 33296 7275
rect 33300 7267 33304 7275
rect 33320 7267 33336 7275
rect 33352 7267 33368 7275
rect 33376 7267 33400 7275
rect 33416 7267 33440 7275
rect 33456 7267 33460 7275
rect 33464 7267 33476 7275
rect 33484 7267 33500 7275
rect 33508 7267 33520 7275
rect 33524 7267 33528 7275
rect 33548 7267 33552 7275
rect 33556 7267 33568 7275
rect 33580 7267 33584 7275
rect 33588 7267 33592 7275
rect 33612 7267 33616 7275
rect 33620 7267 33624 7275
rect 33736 7267 33740 7275
rect 33744 7267 33748 7275
rect 33760 7267 33772 7275
rect 33776 7267 33780 7275
rect 33800 7267 33804 7275
rect 33808 7267 33820 7275
rect 33832 7267 33836 7275
rect 33840 7267 33844 7275
rect 33940 7267 33944 7275
rect 33948 7267 33952 7275
rect 34048 7267 34052 7275
rect 34056 7267 34068 7275
rect 34080 7267 34084 7275
rect 34088 7267 34092 7275
rect 34104 7267 34116 7275
rect 34120 7267 34124 7275
rect 34140 7267 34144 7275
rect 34148 7267 34160 7275
rect 34172 7267 34176 7275
rect 34180 7267 34184 7275
rect 34196 7267 34208 7275
rect 34212 7267 34216 7275
rect 34312 7267 34316 7275
rect 34320 7267 34324 7275
rect 34336 7267 34348 7275
rect 34352 7267 34356 7275
rect 34376 7267 34380 7275
rect 34384 7267 34388 7275
rect 34404 7267 34452 7275
rect 34468 7267 34480 7275
rect 34496 7267 34544 7275
rect 34560 7267 34576 7275
rect 34592 7267 34608 7275
rect 34624 7267 34640 7275
rect 34656 7267 34704 7275
rect 34716 7267 34732 7275
rect 34748 7267 34796 7275
rect 34812 7267 34824 7275
rect 34828 7267 34832 7275
rect 34844 7267 34856 7275
rect 34868 7267 34872 7275
rect 34876 7267 34888 7275
rect 34904 7267 34944 7275
rect 34960 7267 34972 7275
rect 34988 7267 35020 7275
rect 35028 7267 35044 7275
rect 35060 7267 35076 7275
rect 35092 7267 35096 7275
rect 35100 7267 35112 7275
rect 35124 7267 35128 7275
rect 35132 7267 35136 7275
rect 35148 7267 35160 7275
rect 35176 7267 35192 7275
rect 35208 7267 35232 7275
rect 35248 7267 35260 7275
rect 35264 7267 35268 7275
rect 35280 7267 35292 7275
rect 35300 7267 35316 7275
rect 35332 7267 35336 7275
rect 35340 7267 35344 7275
rect 35356 7267 35368 7275
rect 35372 7267 35384 7275
rect 35396 7267 35400 7275
rect 35404 7267 35408 7275
rect 35424 7267 35440 7275
rect 35448 7267 35460 7275
rect 35464 7267 35476 7275
rect 35488 7267 35492 7275
rect 35496 7267 35500 7275
rect 35512 7267 35524 7275
rect 35528 7267 35532 7275
rect 35552 7267 35556 7275
rect 35560 7267 35564 7275
rect 35580 7267 35596 7275
rect 35604 7267 35636 7275
rect 35644 7267 35660 7275
rect 35676 7267 35700 7275
rect 35716 7267 35728 7275
rect 35748 7267 35760 7275
rect 35764 7267 35776 7275
rect 35780 7267 35784 7275
rect 35800 7267 35804 7275
rect 35808 7267 35812 7275
rect 35832 7267 35836 7275
rect 35840 7267 35852 7275
rect 35856 7267 35868 7275
rect 35872 7267 35876 7275
rect 35896 7267 35900 7275
rect 35904 7267 35908 7275
rect 35928 7267 35932 7275
rect 35936 7267 35940 7275
rect 35960 7267 35964 7275
rect 35968 7267 35972 7275
rect 35992 7267 35996 7275
rect 36000 7267 36012 7275
rect 36016 7267 36028 7275
rect 36032 7267 36036 7275
rect 36084 7267 36088 7275
rect 36092 7267 36104 7275
rect 36108 7267 36120 7275
rect 36124 7267 36128 7275
rect 36384 7267 36388 7275
rect 36392 7267 36396 7275
rect 36416 7267 36420 7275
rect 36424 7267 36436 7275
rect 36440 7267 36452 7275
rect 36456 7267 36460 7275
rect 36476 7267 36480 7275
rect 36484 7267 36488 7275
rect 36508 7267 36512 7275
rect 36516 7267 36528 7275
rect 36532 7267 36544 7275
rect 36548 7267 36552 7275
rect 36572 7267 36576 7275
rect 36580 7267 36584 7275
rect 36600 7267 36616 7275
rect 36624 7267 36648 7275
rect 36664 7267 36676 7275
rect 36680 7267 36684 7275
rect 36696 7267 36708 7275
rect 36720 7267 36724 7275
rect 36728 7267 36740 7275
rect 36744 7267 36748 7275
rect 36760 7267 36772 7275
rect 36784 7267 36788 7275
rect 36792 7267 36800 7275
rect 36824 7267 36836 7275
rect 36848 7267 36852 7275
rect 36856 7267 36868 7275
rect 36940 7267 36944 7275
rect 36948 7267 36960 7275
rect 37072 7267 37084 7275
rect 37104 7267 37116 7275
rect 37120 7267 37124 7275
rect 37136 7267 37148 7275
rect 37160 7267 37164 7275
rect 37168 7267 37180 7275
rect 37196 7267 37208 7275
rect 37212 7267 37216 7275
rect 37228 7267 37240 7275
rect 37252 7267 37256 7275
rect 37260 7267 37272 7275
rect 37288 7267 37300 7275
rect 37304 7267 37308 7275
rect 37320 7267 37332 7275
rect 37344 7267 37348 7275
rect 37352 7267 37364 7275
rect 37380 7267 37392 7275
rect 37396 7267 37400 7275
rect 37412 7267 37424 7275
rect 37436 7267 37440 7275
rect 37444 7267 37456 7275
rect 37472 7267 37496 7275
rect 37504 7267 37516 7275
rect 37524 7267 37548 7275
rect 37564 7267 37588 7275
rect 37600 7267 37612 7275
rect 37628 7267 37644 7275
rect 37660 7267 37664 7275
rect 37668 7267 37680 7275
rect 37684 7267 37696 7275
rect 37700 7267 37704 7275
rect 37724 7267 37728 7275
rect 37732 7267 37744 7275
rect 37748 7267 37760 7275
rect 37764 7267 37768 7275
rect 38040 7267 38044 7275
rect 38048 7267 38052 7275
rect 38116 7267 38120 7275
rect 38124 7267 38128 7275
rect 38224 7267 38228 7275
rect 38232 7267 38244 7275
rect 38248 7267 38260 7275
rect 38264 7267 38268 7275
rect 38288 7267 38292 7275
rect 38296 7267 38300 7275
rect 38312 7267 38324 7275
rect 38328 7267 38332 7275
rect 38352 7267 38356 7275
rect 38360 7267 38364 7275
rect 38384 7267 38388 7275
rect 38392 7267 38400 7275
rect 38416 7267 38420 7275
rect 38424 7267 38428 7275
rect 38448 7267 38452 7275
rect 38456 7267 38460 7275
rect 38508 7267 38512 7275
rect 38516 7267 38520 7275
rect 38540 7267 38544 7275
rect 38548 7267 38552 7275
rect 38564 7267 38576 7275
rect 38580 7267 38584 7275
rect 38604 7267 38608 7275
rect 38612 7267 38616 7275
rect 38628 7267 38640 7275
rect 38644 7267 38656 7275
rect 38776 7267 38780 7275
rect 38784 7267 38796 7275
rect 38800 7267 38812 7275
rect 38832 7267 38844 7275
rect 38860 7267 38884 7275
rect 38892 7267 38908 7275
rect 38924 7267 38928 7275
rect 38932 7267 38936 7275
rect 38948 7267 38960 7275
rect 38964 7267 38976 7275
rect 38984 7267 39000 7275
rect 39016 7267 39032 7275
rect 39040 7267 39052 7275
rect 39056 7267 39068 7275
rect 39076 7267 39092 7275
rect 39108 7267 39112 7275
rect 39116 7267 39120 7275
rect 39132 7267 39144 7275
rect 39148 7267 39160 7275
rect 39168 7267 39184 7275
rect 39200 7267 39248 7275
rect 39264 7267 39312 7275
rect 39328 7267 39344 7275
rect 39352 7267 39364 7275
rect 39368 7267 39380 7275
rect 39392 7267 39396 7275
rect 39400 7267 39404 7275
rect 39424 7267 39428 7275
rect 39432 7267 39436 7275
rect 39456 7267 39460 7275
rect 39464 7267 39468 7275
rect 39488 7267 39492 7275
rect 39496 7267 39500 7275
rect 39512 7267 39524 7275
rect 39528 7267 39540 7275
rect 39548 7267 39564 7275
rect 39580 7267 39596 7275
rect 39604 7267 39616 7275
rect 39620 7267 39632 7275
rect 39640 7267 39656 7275
rect 39672 7267 39688 7275
rect 39696 7267 39708 7275
rect 39712 7267 39724 7275
rect 39736 7267 39740 7275
rect 39744 7267 39748 7275
rect 39760 7267 39772 7275
rect 39776 7267 39788 7275
rect 39796 7267 39812 7275
rect 39828 7267 39844 7275
rect 39852 7267 39876 7275
rect 39892 7267 39908 7275
rect 39916 7267 39948 7275
rect 39956 7267 39972 7275
rect 39988 7267 40000 7275
rect 40004 7267 40016 7275
rect 40020 7267 40032 7275
rect 40048 7267 40060 7275
rect 40080 7267 40092 7275
rect 40096 7267 40108 7275
rect 40112 7267 40124 7275
rect 40144 7267 40156 7275
rect 40260 7267 40264 7275
rect 40268 7267 40280 7275
rect 40284 7267 40288 7275
rect 40300 7267 40312 7275
rect 40324 7267 40328 7275
rect 40332 7267 40344 7275
rect 40360 7267 40384 7275
rect 40392 7267 40408 7275
rect 40424 7267 40440 7275
rect 40456 7267 40472 7275
rect 40480 7267 40504 7275
rect 40520 7267 40544 7275
rect 40552 7267 40564 7275
rect 40576 7267 40580 7275
rect 40584 7267 40596 7275
rect 40600 7267 40604 7275
rect 40644 7267 40656 7275
rect 40668 7267 40672 7275
rect 40676 7267 40688 7275
rect 40692 7267 40696 7275
rect 40736 7267 40748 7275
rect 40760 7267 40764 7275
rect 40768 7267 40780 7275
rect 40784 7267 40788 7275
rect 33472 7257 33480 7265
rect 32656 7237 32664 7245
rect 40656 7237 40664 7245
rect 31392 7217 31400 7225
rect 31664 7217 31672 7225
rect 33488 7217 33496 7225
rect 35520 7217 35528 7225
rect 36560 7217 36568 7225
rect 39136 7217 39144 7225
rect 40608 7197 40616 7205
rect 21136 7180 21144 7188
rect 24672 7180 24680 7188
rect 29504 7177 29512 7185
rect 30096 7177 30104 7185
rect 30512 7177 30520 7185
rect 31872 7177 31880 7185
rect 32224 7177 32232 7185
rect 32448 7177 32456 7185
rect 33456 7177 33464 7185
rect 34784 7177 34792 7185
rect 36224 7177 36232 7185
rect 39664 7177 39672 7185
rect 19056 7161 19066 7166
rect 19264 7160 19272 7168
rect 19872 7160 19880 7168
rect 20688 7160 20696 7168
rect 21568 7160 21576 7168
rect 22608 7160 22616 7168
rect 23712 7160 23720 7168
rect 23904 7160 23912 7168
rect 24320 7160 24328 7168
rect 25796 7161 25799 7166
rect 26416 7160 26424 7168
rect 27856 7160 27864 7168
rect 29712 7157 29720 7165
rect 40192 7157 40200 7165
rect 40288 7157 40296 7165
rect 18864 7140 18872 7148
rect 19456 7140 19464 7148
rect 28240 7140 28248 7148
rect 30112 7137 30120 7145
rect 31312 7137 31320 7145
rect 31456 7137 31464 7145
rect 31904 7137 31912 7145
rect 32368 7137 32376 7145
rect 32752 7137 32760 7145
rect 34080 7137 34088 7145
rect 34176 7137 34184 7145
rect 34560 7137 34568 7145
rect 34592 7137 34600 7145
rect 34752 7137 34760 7145
rect 35648 7137 35656 7145
rect 35696 7137 35704 7145
rect 36032 7137 36040 7145
rect 36160 7137 36168 7145
rect 36208 7137 36216 7145
rect 37232 7137 37240 7145
rect 38080 7137 38088 7145
rect 39680 7137 39688 7145
rect 40112 7137 40120 7145
rect 40304 7137 40312 7145
rect 40432 7137 40440 7145
rect 19248 7120 19256 7128
rect 20064 7120 20072 7128
rect 20480 7120 20488 7128
rect 21296 7120 21304 7128
rect 21920 7120 21928 7128
rect 22592 7120 22600 7128
rect 22992 7120 23000 7128
rect 23520 7120 23528 7128
rect 23904 7120 23912 7128
rect 24144 7120 24152 7128
rect 24752 7120 24760 7128
rect 24960 7120 24968 7128
rect 27440 7120 27448 7128
rect 27520 7120 27528 7128
rect 28064 7120 28072 7128
rect 29856 7117 29864 7125
rect 30336 7117 30344 7125
rect 30624 7117 30632 7125
rect 30800 7117 30808 7125
rect 31008 7117 31016 7125
rect 32528 7117 32536 7125
rect 32592 7117 32600 7125
rect 33584 7117 33592 7125
rect 33632 7117 33640 7125
rect 33872 7117 33880 7125
rect 35760 7117 35768 7125
rect 36864 7117 36872 7125
rect 37648 7117 37656 7125
rect 37744 7117 37752 7125
rect 37840 7117 37848 7125
rect 37984 7117 37992 7125
rect 38000 7117 38008 7125
rect 38496 7117 38504 7125
rect 38672 7117 38680 7125
rect 18624 7100 18632 7108
rect 19696 7100 19704 7108
rect 21728 7100 21736 7108
rect 23728 7100 23736 7108
rect 24064 7100 24072 7108
rect 25136 7100 25144 7108
rect 25376 7100 25384 7108
rect 25584 7100 25592 7108
rect 26128 7100 26136 7108
rect 26144 7100 26152 7108
rect 35688 7105 35689 7110
rect 30128 7097 30136 7105
rect 32864 7097 32872 7105
rect 33920 7097 33928 7105
rect 34656 7097 34664 7105
rect 36800 7097 36808 7105
rect 37088 7097 37096 7105
rect 38720 7097 38728 7105
rect 39040 7097 39048 7105
rect 39472 7097 39480 7105
rect 39600 7097 39608 7105
rect 19488 7080 19496 7088
rect 20720 7080 20728 7088
rect 21120 7080 21128 7088
rect 21744 7080 21752 7088
rect 22176 7080 22184 7088
rect 22816 7080 22824 7088
rect 26592 7080 26600 7088
rect 23248 7060 23256 7068
rect 25968 7060 25976 7068
rect 29396 7067 29408 7075
rect 29420 7067 29424 7075
rect 29428 7067 29440 7075
rect 29444 7067 29448 7075
rect 29460 7067 29472 7075
rect 29488 7067 29504 7075
rect 29520 7067 29544 7075
rect 29552 7067 29568 7075
rect 29576 7067 29588 7075
rect 29592 7067 29596 7075
rect 29616 7067 29620 7075
rect 29624 7067 29636 7075
rect 29640 7067 29652 7075
rect 29656 7067 29660 7075
rect 29680 7067 29684 7075
rect 29688 7067 29692 7075
rect 29708 7067 29712 7075
rect 29716 7067 29728 7075
rect 29732 7067 29744 7075
rect 29748 7067 29752 7075
rect 29772 7067 29776 7075
rect 29780 7067 29784 7075
rect 29832 7067 29836 7075
rect 29840 7067 29844 7075
rect 29864 7067 29868 7075
rect 29872 7067 29876 7075
rect 29888 7067 29900 7075
rect 29904 7067 29908 7075
rect 29928 7067 29932 7075
rect 29936 7067 29940 7075
rect 29960 7067 29964 7075
rect 29968 7067 29980 7075
rect 29992 7067 29996 7075
rect 30000 7067 30004 7075
rect 30024 7067 30028 7075
rect 30032 7067 30044 7075
rect 30048 7067 30060 7075
rect 30064 7067 30068 7075
rect 30116 7067 30120 7075
rect 30124 7067 30136 7075
rect 30140 7067 30152 7075
rect 30156 7067 30160 7075
rect 30208 7067 30212 7075
rect 30216 7067 30228 7075
rect 30232 7067 30244 7075
rect 30248 7067 30252 7075
rect 30272 7067 30276 7075
rect 30280 7067 30284 7075
rect 30300 7067 30316 7075
rect 30324 7067 30348 7075
rect 30364 7067 30376 7075
rect 30380 7067 30384 7075
rect 30400 7067 30408 7075
rect 30420 7067 30424 7075
rect 30428 7067 30440 7075
rect 30804 7067 30816 7075
rect 30828 7067 30832 7075
rect 30836 7067 30848 7075
rect 30852 7067 30856 7075
rect 30868 7067 30880 7075
rect 30920 7067 30924 7075
rect 30928 7067 30940 7075
rect 30944 7067 30948 7075
rect 30960 7067 30972 7075
rect 30992 7067 31004 7075
rect 31020 7067 31044 7075
rect 31052 7067 31068 7075
rect 31076 7067 31100 7075
rect 31116 7067 31132 7075
rect 31140 7067 31164 7075
rect 31180 7067 31192 7075
rect 31196 7067 31200 7075
rect 31212 7067 31224 7075
rect 31232 7067 31256 7075
rect 31272 7067 31284 7075
rect 31288 7067 31292 7075
rect 31304 7067 31316 7075
rect 31324 7067 31348 7075
rect 31364 7067 31412 7075
rect 31428 7067 31440 7075
rect 31460 7067 31472 7075
rect 31484 7067 31488 7075
rect 31492 7067 31504 7075
rect 31648 7067 31660 7075
rect 31664 7067 31668 7075
rect 31740 7067 31752 7075
rect 31772 7067 31784 7075
rect 31788 7067 31792 7075
rect 31804 7067 31816 7075
rect 31828 7067 31832 7075
rect 31836 7067 31848 7075
rect 31852 7067 31856 7075
rect 31960 7067 31972 7075
rect 31992 7067 32004 7075
rect 32008 7067 32020 7075
rect 32032 7067 32036 7075
rect 32040 7067 32044 7075
rect 32056 7067 32068 7075
rect 32080 7067 32084 7075
rect 32088 7067 32100 7075
rect 32104 7067 32108 7075
rect 32120 7067 32132 7075
rect 32148 7067 32160 7075
rect 32172 7067 32176 7075
rect 32180 7067 32192 7075
rect 32196 7067 32200 7075
rect 32212 7067 32224 7075
rect 32236 7067 32240 7075
rect 32244 7067 32256 7075
rect 32272 7067 32296 7075
rect 32304 7067 32320 7075
rect 32336 7067 32340 7075
rect 32344 7067 32348 7075
rect 32368 7067 32372 7075
rect 32376 7067 32388 7075
rect 32392 7067 32404 7075
rect 32408 7067 32412 7075
rect 32432 7067 32436 7075
rect 32440 7067 32452 7075
rect 32460 7067 32476 7075
rect 32484 7067 32508 7075
rect 32524 7067 32540 7075
rect 32556 7067 32568 7075
rect 32580 7067 32584 7075
rect 32588 7067 32600 7075
rect 32604 7067 32608 7075
rect 32620 7067 32632 7075
rect 32696 7067 32708 7075
rect 32728 7067 32740 7075
rect 32744 7067 32748 7075
rect 32764 7067 32780 7075
rect 32800 7067 32828 7075
rect 32844 7067 32856 7075
rect 32876 7067 32888 7075
rect 32900 7067 32904 7075
rect 32908 7067 32912 7075
rect 33000 7067 33012 7075
rect 33024 7067 33028 7075
rect 33032 7067 33036 7075
rect 33048 7067 33060 7075
rect 33068 7067 33084 7075
rect 33100 7067 33116 7075
rect 33124 7067 33136 7075
rect 33148 7067 33152 7075
rect 33156 7067 33160 7075
rect 33172 7067 33184 7075
rect 33200 7067 33216 7075
rect 33232 7067 33256 7075
rect 33272 7067 33284 7075
rect 33288 7067 33292 7075
rect 33312 7067 33316 7075
rect 33320 7067 33332 7075
rect 33468 7067 33472 7075
rect 33476 7067 33480 7075
rect 33592 7067 33596 7075
rect 33600 7067 33604 7075
rect 33616 7067 33628 7075
rect 33632 7067 33636 7075
rect 33652 7067 33676 7075
rect 33684 7067 33700 7075
rect 33708 7067 33732 7075
rect 33744 7067 33768 7075
rect 33776 7067 33792 7075
rect 33800 7067 33824 7075
rect 33840 7067 33852 7075
rect 33872 7067 33884 7075
rect 33896 7067 33900 7075
rect 33904 7067 33916 7075
rect 33920 7067 33924 7075
rect 33936 7067 33948 7075
rect 33956 7067 33980 7075
rect 33996 7067 34020 7075
rect 34028 7067 34040 7075
rect 34048 7067 34072 7075
rect 34088 7067 34112 7075
rect 34120 7067 34136 7075
rect 34152 7067 34156 7075
rect 34160 7067 34164 7075
rect 34184 7067 34188 7075
rect 34192 7067 34204 7075
rect 34208 7067 34220 7075
rect 34224 7067 34228 7075
rect 34244 7067 34268 7075
rect 34276 7067 34292 7075
rect 34300 7067 34324 7075
rect 34340 7067 34356 7075
rect 34372 7067 34384 7075
rect 34396 7067 34400 7075
rect 34404 7067 34416 7075
rect 34420 7067 34424 7075
rect 34488 7067 34492 7075
rect 34496 7067 34508 7075
rect 34512 7067 34516 7075
rect 34528 7067 34540 7075
rect 34552 7067 34556 7075
rect 34560 7067 34572 7075
rect 34592 7067 34604 7075
rect 34616 7067 34620 7075
rect 34624 7067 34636 7075
rect 34708 7067 34712 7075
rect 34716 7067 34728 7075
rect 34748 7067 34760 7075
rect 34764 7067 34776 7075
rect 34780 7067 34792 7075
rect 34812 7067 34824 7075
rect 34828 7067 34832 7075
rect 34904 7067 34916 7075
rect 34920 7067 34924 7075
rect 34936 7067 34948 7075
rect 34964 7067 34980 7075
rect 34996 7067 35044 7075
rect 35060 7067 35076 7075
rect 35084 7067 35096 7075
rect 35100 7067 35112 7075
rect 35124 7067 35128 7075
rect 35132 7067 35136 7075
rect 35152 7067 35168 7075
rect 35176 7067 35200 7075
rect 35216 7067 35232 7075
rect 35240 7067 35272 7075
rect 35280 7067 35292 7075
rect 35308 7067 35324 7075
rect 35332 7067 35364 7075
rect 35372 7067 35388 7075
rect 35404 7067 35420 7075
rect 35436 7067 35440 7075
rect 35444 7067 35456 7075
rect 35468 7067 35472 7075
rect 35476 7067 35480 7075
rect 35492 7067 35504 7075
rect 35508 7067 35520 7075
rect 35528 7067 35544 7075
rect 35560 7067 35576 7075
rect 35584 7067 35596 7075
rect 35600 7067 35612 7075
rect 35624 7067 35628 7075
rect 35632 7067 35636 7075
rect 35648 7067 35660 7075
rect 35664 7067 35668 7075
rect 35688 7067 35692 7075
rect 35696 7067 35700 7075
rect 35712 7067 35724 7075
rect 35728 7067 35732 7075
rect 35748 7067 35772 7075
rect 35780 7067 35796 7075
rect 35804 7067 35816 7075
rect 35820 7067 35824 7075
rect 35844 7067 35848 7075
rect 35852 7067 35864 7075
rect 35868 7067 35880 7075
rect 35884 7067 35888 7075
rect 35908 7067 35912 7075
rect 35916 7067 35920 7075
rect 35936 7067 35952 7075
rect 35960 7067 35984 7075
rect 36000 7067 36012 7075
rect 36016 7067 36020 7075
rect 36032 7067 36044 7075
rect 36056 7067 36060 7075
rect 36064 7067 36076 7075
rect 36092 7067 36104 7075
rect 36108 7067 36112 7075
rect 36124 7067 36136 7075
rect 36148 7067 36152 7075
rect 36156 7067 36168 7075
rect 36188 7067 36200 7075
rect 36312 7067 36324 7075
rect 36328 7067 36332 7075
rect 36344 7067 36356 7075
rect 36376 7067 36388 7075
rect 36404 7067 36452 7075
rect 36464 7067 36480 7075
rect 36496 7067 36544 7075
rect 36560 7067 36576 7075
rect 36592 7067 36596 7075
rect 36600 7067 36612 7075
rect 36624 7067 36628 7075
rect 36632 7067 36636 7075
rect 36656 7067 36660 7075
rect 36664 7067 36668 7075
rect 36764 7067 36768 7075
rect 36772 7067 36776 7075
rect 36788 7067 36800 7075
rect 36804 7067 36808 7075
rect 36824 7067 36840 7075
rect 36856 7067 36872 7075
rect 36880 7067 36912 7075
rect 36920 7067 36932 7075
rect 36948 7067 36964 7075
rect 36972 7067 37004 7075
rect 37012 7067 37028 7075
rect 37036 7067 37060 7075
rect 37076 7067 37088 7075
rect 37108 7067 37120 7075
rect 37132 7067 37136 7075
rect 37140 7067 37152 7075
rect 37156 7067 37160 7075
rect 37200 7067 37212 7075
rect 37224 7067 37228 7075
rect 37232 7067 37244 7075
rect 37248 7067 37252 7075
rect 37292 7067 37304 7075
rect 37316 7067 37320 7075
rect 37324 7067 37336 7075
rect 37340 7067 37344 7075
rect 37356 7067 37368 7075
rect 37384 7067 37400 7075
rect 37416 7067 37440 7075
rect 37448 7067 37464 7075
rect 37472 7067 37496 7075
rect 37512 7067 37516 7075
rect 37520 7067 37532 7075
rect 37536 7067 37548 7075
rect 37552 7067 37556 7075
rect 37576 7067 37580 7075
rect 37584 7067 37588 7075
rect 37600 7067 37612 7075
rect 37616 7067 37620 7075
rect 37636 7067 37652 7075
rect 37668 7067 37716 7075
rect 37732 7067 37744 7075
rect 37748 7067 37752 7075
rect 37764 7067 37776 7075
rect 37788 7067 37792 7075
rect 37796 7067 37808 7075
rect 37812 7067 37816 7075
rect 37828 7067 37840 7075
rect 37920 7067 37932 7075
rect 37952 7067 37964 7075
rect 37968 7067 37980 7075
rect 37984 7067 37996 7075
rect 38012 7067 38028 7075
rect 38044 7067 38056 7075
rect 38060 7067 38072 7075
rect 38076 7067 38088 7075
rect 38108 7067 38120 7075
rect 38136 7067 38148 7075
rect 38152 7067 38164 7075
rect 38168 7067 38180 7075
rect 38200 7067 38212 7075
rect 38452 7067 38464 7075
rect 38468 7067 38480 7075
rect 38484 7067 38496 7075
rect 38512 7067 38524 7075
rect 38544 7067 38556 7075
rect 38560 7067 38572 7075
rect 38576 7067 38588 7075
rect 38608 7067 38620 7075
rect 38624 7067 38636 7075
rect 38640 7067 38652 7075
rect 38672 7067 38684 7075
rect 38700 7067 38724 7075
rect 38732 7067 38748 7075
rect 38764 7067 38768 7075
rect 38772 7067 38776 7075
rect 38788 7067 38800 7075
rect 38804 7067 38816 7075
rect 38828 7067 38832 7075
rect 38836 7067 38840 7075
rect 38860 7067 38864 7075
rect 38868 7067 38880 7075
rect 38892 7067 38896 7075
rect 38900 7067 38904 7075
rect 38924 7067 38928 7075
rect 38932 7067 38936 7075
rect 38948 7067 38960 7075
rect 38964 7067 38968 7075
rect 38984 7067 39000 7075
rect 39016 7067 39064 7075
rect 39076 7067 39092 7075
rect 39108 7067 39156 7075
rect 39168 7067 39184 7075
rect 39200 7067 39248 7075
rect 39264 7067 39268 7075
rect 39272 7067 39276 7075
rect 39288 7067 39300 7075
rect 39304 7067 39316 7075
rect 39328 7067 39332 7075
rect 39336 7067 39340 7075
rect 39436 7067 39440 7075
rect 39444 7067 39448 7075
rect 39468 7067 39472 7075
rect 39476 7067 39480 7075
rect 39492 7067 39504 7075
rect 39508 7067 39520 7075
rect 39532 7067 39536 7075
rect 39540 7067 39544 7075
rect 39640 7067 39644 7075
rect 39648 7067 39660 7075
rect 39672 7067 39676 7075
rect 39680 7067 39684 7075
rect 39780 7067 39784 7075
rect 39788 7067 39792 7075
rect 39904 7067 39908 7075
rect 39912 7067 39924 7075
rect 39928 7067 39940 7075
rect 39944 7067 39948 7075
rect 39968 7067 39972 7075
rect 39976 7067 39980 7075
rect 40044 7067 40048 7075
rect 40052 7067 40056 7075
rect 40076 7067 40080 7075
rect 40084 7067 40096 7075
rect 40100 7067 40112 7075
rect 40116 7067 40120 7075
rect 40140 7067 40144 7075
rect 40148 7067 40152 7075
rect 40168 7067 40172 7075
rect 40176 7067 40188 7075
rect 40192 7067 40204 7075
rect 40208 7067 40212 7075
rect 40232 7067 40236 7075
rect 40240 7067 40244 7075
rect 40260 7067 40276 7075
rect 40284 7067 40308 7075
rect 40324 7067 40348 7075
rect 40356 7067 40368 7075
rect 40380 7067 40384 7075
rect 40388 7067 40400 7075
rect 40404 7067 40408 7075
rect 40420 7067 40432 7075
rect 40452 7067 40464 7075
rect 40480 7067 40504 7075
rect 40512 7067 40528 7075
rect 40536 7067 40560 7075
rect 40576 7067 40580 7075
rect 40584 7067 40596 7075
rect 40600 7067 40612 7075
rect 40616 7067 40620 7075
rect 40636 7067 40652 7075
rect 40668 7067 40684 7075
rect 40692 7067 40716 7075
rect 40732 7067 40744 7075
rect 40748 7067 40752 7075
rect 40764 7067 40776 7075
rect 40788 7067 40792 7075
rect 40796 7067 40800 7075
rect 18536 7056 18538 7060
rect 18948 7056 18950 7060
rect 19574 7056 19576 7060
rect 19772 7056 19774 7060
rect 19986 7056 19988 7060
rect 18542 7052 18544 7056
rect 18954 7052 18956 7056
rect 19580 7052 19582 7056
rect 19778 7052 19780 7056
rect 19992 7052 19994 7056
rect 20152 7050 20160 7058
rect 20302 7050 20308 7058
rect 20906 7050 20920 7058
rect 21174 7050 21182 7058
rect 21326 7050 21332 7058
rect 21334 7050 21348 7058
rect 21388 7050 21402 7058
rect 21800 7050 21808 7058
rect 21952 7050 21958 7058
rect 21960 7050 21966 7058
rect 22228 7050 22236 7058
rect 22316 7050 22322 7058
rect 22324 7050 22330 7058
rect 22594 7050 22600 7058
rect 22602 7050 22608 7058
rect 22656 7050 22664 7058
rect 22744 7050 22750 7058
rect 22752 7050 22758 7058
rect 23022 7050 23028 7058
rect 23030 7050 23036 7058
rect 23322 7050 23328 7058
rect 23330 7050 23336 7058
rect 23480 7050 23486 7058
rect 23750 7050 23756 7058
rect 23758 7050 23764 7058
rect 23948 7050 23954 7058
rect 23956 7050 23962 7058
rect 24106 7050 24112 7058
rect 24154 7050 24168 7058
rect 24304 7050 24310 7058
rect 24360 7050 24366 7058
rect 24368 7050 24374 7058
rect 24986 7050 24992 7058
rect 24994 7050 25000 7058
rect 25248 7050 25254 7058
rect 25256 7050 25262 7058
rect 25342 7050 25348 7058
rect 25398 7050 25404 7058
rect 25406 7050 25412 7058
rect 25556 7050 25562 7058
rect 25612 7050 25618 7058
rect 25620 7050 25626 7058
rect 25770 7050 25776 7058
rect 26016 7050 26024 7058
rect 26104 7050 26110 7058
rect 26112 7050 26118 7058
rect 26452 7050 26458 7058
rect 26460 7050 26466 7058
rect 27156 7050 27162 7058
rect 27564 7050 27574 7058
rect 27778 7050 27788 7058
rect 27876 7050 27880 7058
rect 27884 7050 27888 7058
rect 28082 7050 28094 7058
rect 28172 7050 28180 7058
rect 28386 7050 28394 7058
rect 33728 7057 33736 7065
rect 34032 7057 34040 7065
rect 38048 7057 38056 7065
rect 20992 7040 21000 7048
rect 26448 7040 26456 7048
rect 29984 7037 29992 7045
rect 31312 7037 31320 7045
rect 31792 7037 31800 7045
rect 33952 7037 33960 7045
rect 34144 7037 34152 7045
rect 34560 7037 34568 7045
rect 35568 7037 35576 7045
rect 36768 7037 36776 7045
rect 38800 7037 38808 7045
rect 18880 7020 18888 7028
rect 19488 7020 19496 7028
rect 19728 7020 19736 7028
rect 20752 7020 20760 7028
rect 21184 7020 21192 7028
rect 22032 7020 22040 7028
rect 25808 7020 25816 7028
rect 27408 7020 27416 7028
rect 27600 7020 27608 7028
rect 27728 7020 27736 7028
rect 28000 7020 28008 7028
rect 29376 7017 29384 7025
rect 29648 7017 29656 7025
rect 30752 7017 30760 7025
rect 34240 7017 34248 7025
rect 35024 7017 35032 7025
rect 35072 7017 35080 7025
rect 35280 7017 35288 7025
rect 35824 7017 35832 7025
rect 35872 7017 35880 7025
rect 36400 7017 36408 7025
rect 39136 7017 39144 7025
rect 39600 7017 39608 7025
rect 40400 7017 40408 7025
rect 21840 7000 21848 7008
rect 22416 7000 22424 7008
rect 22432 7000 22440 7008
rect 23072 7000 23080 7008
rect 24768 7000 24776 7008
rect 25168 7000 25176 7008
rect 28560 7000 28568 7008
rect 29808 6997 29816 7005
rect 29952 6997 29960 7005
rect 30608 6997 30616 7005
rect 31456 6997 31464 7005
rect 33376 6997 33384 7005
rect 33536 6997 33544 7005
rect 33696 6997 33704 7005
rect 33776 6997 33784 7005
rect 33968 6997 33976 7005
rect 35104 6997 35112 7005
rect 35408 6997 35416 7005
rect 35792 6997 35800 7005
rect 36352 6997 36360 7005
rect 37680 6997 37688 7005
rect 37952 6997 37960 7005
rect 38544 6997 38552 7005
rect 39376 6997 39384 7005
rect 39728 6997 39736 7005
rect 39872 6997 39880 7005
rect 19680 6980 19688 6988
rect 21520 6980 21528 6988
rect 23536 6980 23544 6988
rect 23696 6980 23704 6988
rect 24288 6980 24296 6988
rect 24368 6980 24376 6988
rect 24400 6980 24408 6988
rect 25120 6980 25128 6988
rect 25456 6980 25464 6988
rect 25648 6980 25656 6988
rect 26080 6980 26088 6988
rect 26896 6980 26904 6988
rect 27136 6980 27144 6988
rect 27296 6980 27304 6988
rect 28208 6980 28216 6988
rect 29488 6977 29496 6985
rect 31632 6977 31640 6985
rect 31936 6977 31944 6985
rect 20496 6960 20504 6968
rect 20720 6960 20728 6968
rect 30080 6957 30088 6965
rect 32864 6957 32872 6965
rect 33008 6957 33016 6965
rect 33088 6957 33096 6965
rect 33760 6957 33768 6965
rect 34000 6957 34008 6965
rect 34448 6957 34456 6965
rect 35552 6957 35560 6965
rect 35776 6957 35784 6965
rect 36480 6957 36488 6965
rect 36848 6957 36856 6965
rect 36944 6957 36952 6965
rect 37232 6957 37240 6965
rect 37936 6957 37944 6965
rect 38656 6957 38664 6965
rect 19072 6948 19076 6953
rect 23970 6948 23974 6953
rect 27899 6948 27908 6953
rect 18720 6940 18728 6948
rect 21152 6940 21160 6948
rect 21568 6940 21576 6948
rect 22208 6940 22216 6948
rect 22688 6940 22696 6948
rect 23040 6940 23048 6948
rect 23344 6940 23352 6948
rect 23712 6940 23720 6948
rect 23952 6940 23960 6948
rect 24608 6940 24616 6948
rect 24944 6940 24952 6948
rect 25216 6940 25224 6948
rect 26912 6940 26920 6948
rect 27472 6940 27480 6948
rect 27696 6940 27704 6948
rect 36960 6937 36968 6945
rect 22880 6920 22888 6928
rect 37312 6917 37320 6925
rect 37712 6917 37720 6925
rect 37728 6917 37736 6925
rect 37520 6897 37528 6905
rect 32976 6877 32984 6885
rect 29524 6867 29536 6875
rect 29556 6867 29568 6875
rect 29572 6867 29584 6875
rect 29596 6867 29600 6875
rect 29604 6867 29608 6875
rect 29628 6867 29632 6875
rect 29636 6867 29648 6875
rect 29660 6867 29664 6875
rect 29668 6867 29672 6875
rect 29692 6867 29696 6875
rect 29700 6867 29704 6875
rect 29832 6867 29836 6875
rect 29840 6867 29844 6875
rect 29864 6867 29868 6875
rect 29872 6867 29876 6875
rect 29888 6867 29900 6875
rect 29904 6867 29908 6875
rect 29928 6867 29932 6875
rect 29936 6867 29948 6875
rect 29960 6867 29964 6875
rect 29968 6867 29972 6875
rect 29992 6867 29996 6875
rect 30000 6867 30004 6875
rect 30024 6867 30028 6875
rect 30032 6867 30036 6875
rect 30048 6867 30060 6875
rect 30064 6867 30068 6875
rect 30088 6867 30092 6875
rect 30096 6867 30108 6875
rect 30116 6867 30132 6875
rect 30140 6867 30152 6875
rect 30156 6867 30160 6875
rect 30180 6867 30184 6875
rect 30188 6867 30200 6875
rect 30208 6867 30224 6875
rect 30232 6867 30244 6875
rect 30248 6867 30252 6875
rect 30272 6867 30276 6875
rect 30280 6867 30292 6875
rect 30300 6867 30316 6875
rect 30324 6867 30348 6875
rect 30360 6867 30384 6875
rect 30416 6867 30440 6875
rect 30452 6867 30476 6875
rect 30484 6867 30500 6875
rect 30508 6867 30540 6875
rect 30548 6867 30564 6875
rect 30580 6867 30596 6875
rect 30612 6867 30616 6875
rect 30620 6867 30632 6875
rect 30644 6867 30648 6875
rect 30652 6867 30656 6875
rect 30668 6867 30680 6875
rect 30684 6867 30688 6875
rect 30704 6867 30720 6875
rect 30736 6867 30752 6875
rect 30760 6867 30792 6875
rect 30800 6867 30812 6875
rect 30832 6867 30844 6875
rect 30848 6867 30860 6875
rect 30864 6867 30876 6875
rect 30896 6867 30908 6875
rect 30912 6867 30916 6875
rect 31020 6867 31032 6875
rect 31036 6867 31040 6875
rect 31052 6867 31064 6875
rect 31076 6867 31080 6875
rect 31084 6867 31096 6875
rect 31116 6867 31128 6875
rect 31148 6867 31160 6875
rect 31180 6867 31192 6875
rect 31196 6867 31200 6875
rect 31212 6867 31224 6875
rect 31232 6867 31256 6875
rect 31272 6867 31320 6875
rect 31332 6867 31348 6875
rect 31364 6867 31412 6875
rect 31428 6867 31440 6875
rect 31460 6867 31472 6875
rect 31484 6867 31488 6875
rect 31492 6867 31504 6875
rect 31648 6867 31660 6875
rect 31664 6867 31668 6875
rect 31700 6867 31704 6875
rect 31708 6867 31720 6875
rect 31832 6867 31844 6875
rect 31848 6867 31860 6875
rect 31864 6867 31876 6875
rect 31892 6867 31908 6875
rect 31924 6867 31948 6875
rect 31956 6867 31972 6875
rect 31988 6867 32000 6875
rect 32012 6867 32036 6875
rect 32052 6867 32068 6875
rect 32076 6867 32108 6875
rect 32116 6867 32132 6875
rect 32144 6867 32160 6875
rect 32168 6867 32200 6875
rect 32208 6867 32224 6875
rect 32232 6867 32256 6875
rect 32272 6867 32276 6875
rect 32280 6867 32292 6875
rect 32304 6867 32308 6875
rect 32312 6867 32316 6875
rect 32336 6867 32340 6875
rect 32344 6867 32348 6875
rect 32368 6867 32372 6875
rect 32376 6867 32380 6875
rect 32392 6867 32404 6875
rect 32408 6867 32412 6875
rect 32432 6867 32436 6875
rect 32440 6867 32452 6875
rect 32460 6867 32476 6875
rect 32484 6867 32508 6875
rect 32524 6867 32528 6875
rect 32532 6867 32544 6875
rect 32552 6867 32568 6875
rect 32576 6867 32608 6875
rect 32616 6867 32632 6875
rect 32648 6867 32660 6875
rect 32672 6867 32676 6875
rect 32680 6867 32684 6875
rect 32764 6867 32768 6875
rect 32772 6867 32784 6875
rect 32804 6867 32816 6875
rect 32820 6867 32824 6875
rect 32840 6867 32844 6875
rect 32848 6867 32860 6875
rect 32872 6867 32876 6875
rect 32880 6867 32884 6875
rect 32896 6867 32908 6875
rect 32924 6867 32940 6875
rect 32956 6867 32980 6875
rect 32996 6867 33008 6875
rect 33012 6867 33016 6875
rect 33028 6867 33040 6875
rect 33052 6867 33056 6875
rect 33060 6867 33064 6875
rect 33192 6867 33196 6875
rect 33200 6867 33204 6875
rect 33224 6867 33228 6875
rect 33232 6867 33244 6875
rect 33248 6867 33260 6875
rect 33276 6867 33292 6875
rect 33300 6867 33316 6875
rect 33324 6867 33340 6875
rect 33356 6867 33360 6875
rect 33364 6867 33368 6875
rect 33388 6867 33392 6875
rect 33396 6867 33408 6875
rect 33428 6867 33440 6875
rect 33444 6867 33456 6875
rect 33504 6867 33516 6875
rect 33520 6867 33532 6875
rect 33544 6867 33548 6875
rect 33552 6867 33556 6875
rect 33576 6867 33580 6875
rect 33584 6867 33588 6875
rect 33652 6867 33656 6875
rect 33660 6867 33672 6875
rect 33684 6867 33688 6875
rect 33692 6867 33696 6875
rect 33708 6867 33720 6875
rect 33724 6867 33736 6875
rect 33744 6867 33760 6875
rect 33776 6867 33792 6875
rect 33800 6867 33824 6875
rect 33840 6867 33852 6875
rect 33872 6867 33884 6875
rect 33888 6867 33900 6875
rect 33912 6867 33916 6875
rect 33920 6867 33924 6875
rect 33940 6867 33980 6875
rect 33996 6867 34012 6875
rect 34024 6867 34056 6875
rect 34064 6867 34080 6875
rect 34096 6867 34112 6875
rect 34128 6867 34144 6875
rect 34160 6867 34176 6875
rect 34184 6867 34216 6875
rect 34224 6867 34236 6875
rect 34252 6867 34268 6875
rect 34276 6867 34308 6875
rect 34316 6867 34328 6875
rect 34348 6867 34360 6875
rect 34368 6867 34400 6875
rect 34408 6867 34424 6875
rect 34436 6867 34452 6875
rect 34460 6867 34492 6875
rect 34500 6867 34516 6875
rect 34532 6867 34544 6875
rect 34548 6867 34560 6875
rect 34564 6867 34576 6875
rect 34596 6867 34608 6875
rect 34612 6867 34624 6875
rect 34628 6867 34640 6875
rect 34656 6867 34672 6875
rect 34688 6867 34712 6875
rect 34720 6867 34736 6875
rect 34752 6867 34800 6875
rect 34816 6867 34828 6875
rect 34844 6867 34892 6875
rect 34908 6867 34924 6875
rect 34940 6867 34952 6875
rect 34964 6867 34968 6875
rect 34972 6867 34984 6875
rect 35088 6867 35092 6875
rect 35096 6867 35108 6875
rect 35128 6867 35140 6875
rect 35144 6867 35148 6875
rect 35284 6867 35296 6875
rect 35308 6867 35312 6875
rect 35316 6867 35328 6875
rect 35332 6867 35336 6875
rect 35348 6867 35360 6875
rect 35536 6867 35548 6875
rect 35560 6867 35564 6875
rect 35568 6867 35580 6875
rect 35584 6867 35588 6875
rect 35600 6867 35612 6875
rect 35632 6867 35644 6875
rect 35648 6867 35652 6875
rect 35664 6867 35676 6875
rect 35696 6867 35708 6875
rect 35712 6867 35724 6875
rect 35728 6867 35740 6875
rect 35756 6867 35768 6875
rect 35788 6867 35800 6875
rect 35804 6867 35816 6875
rect 35820 6867 35832 6875
rect 35852 6867 35864 6875
rect 35868 6867 35872 6875
rect 35884 6867 35896 6875
rect 35916 6867 35928 6875
rect 35944 6867 35992 6875
rect 36008 6867 36012 6875
rect 36016 6867 36020 6875
rect 36036 6867 36084 6875
rect 36100 6867 36104 6875
rect 36108 6867 36112 6875
rect 36128 6867 36176 6875
rect 36192 6867 36208 6875
rect 36224 6867 36228 6875
rect 36232 6867 36244 6875
rect 36256 6867 36260 6875
rect 36264 6867 36268 6875
rect 36288 6867 36292 6875
rect 36296 6867 36300 6875
rect 36396 6867 36400 6875
rect 36404 6867 36408 6875
rect 36420 6867 36432 6875
rect 36436 6867 36440 6875
rect 36456 6867 36472 6875
rect 36488 6867 36504 6875
rect 36512 6867 36544 6875
rect 36552 6867 36568 6875
rect 36584 6867 36596 6875
rect 36600 6867 36612 6875
rect 36616 6867 36628 6875
rect 36648 6867 36660 6875
rect 36764 6867 36768 6875
rect 36772 6867 36784 6875
rect 36788 6867 36792 6875
rect 36832 6867 36844 6875
rect 36856 6867 36860 6875
rect 36864 6867 36876 6875
rect 36880 6867 36884 6875
rect 36896 6867 36908 6875
rect 36916 6867 36940 6875
rect 36956 6867 37004 6875
rect 37020 6867 37032 6875
rect 37036 6867 37040 6875
rect 37052 6867 37064 6875
rect 37072 6867 37096 6875
rect 37112 6867 37160 6875
rect 37176 6867 37180 6875
rect 37184 6867 37188 6875
rect 37200 6867 37212 6875
rect 37216 6867 37228 6875
rect 37236 6867 37252 6875
rect 37268 6867 37272 6875
rect 37276 6867 37280 6875
rect 37292 6867 37304 6875
rect 37308 6867 37320 6875
rect 37328 6867 37344 6875
rect 37360 6867 37376 6875
rect 37384 6867 37408 6875
rect 37424 6867 37440 6875
rect 37456 6867 37480 6875
rect 37488 6867 37504 6875
rect 37520 6867 37568 6875
rect 37584 6867 37632 6875
rect 37648 6867 37652 6875
rect 37656 6867 37660 6875
rect 37676 6867 37724 6875
rect 37740 6867 37744 6875
rect 37748 6867 37752 6875
rect 37768 6867 37816 6875
rect 37832 6867 37848 6875
rect 37856 6867 37868 6875
rect 37872 6867 37884 6875
rect 37892 6867 37908 6875
rect 37924 6867 37928 6875
rect 37932 6867 37936 6875
rect 37948 6867 37960 6875
rect 37964 6867 37976 6875
rect 37984 6867 38000 6875
rect 38016 6867 38020 6875
rect 38024 6867 38028 6875
rect 38040 6867 38052 6875
rect 38056 6867 38068 6875
rect 38080 6867 38084 6875
rect 38088 6867 38092 6875
rect 38108 6867 38124 6875
rect 38132 6867 38144 6875
rect 38148 6867 38160 6875
rect 38172 6867 38176 6875
rect 38180 6867 38184 6875
rect 38200 6867 38216 6875
rect 38224 6867 38248 6875
rect 38264 6867 38276 6875
rect 38296 6867 38308 6875
rect 38312 6867 38324 6875
rect 38328 6867 38340 6875
rect 38360 6867 38372 6875
rect 38376 6867 38380 6875
rect 38452 6867 38464 6875
rect 38468 6867 38472 6875
rect 38504 6867 38508 6875
rect 38512 6867 38524 6875
rect 38544 6867 38556 6875
rect 38560 6867 38564 6875
rect 38700 6867 38712 6875
rect 38716 6867 38720 6875
rect 38732 6867 38744 6875
rect 38752 6867 38776 6875
rect 38792 6867 38804 6875
rect 38808 6867 38812 6875
rect 38824 6867 38836 6875
rect 38848 6867 38852 6875
rect 38856 6867 38868 6875
rect 38872 6867 38876 6875
rect 38980 6867 38992 6875
rect 39012 6867 39024 6875
rect 39028 6867 39040 6875
rect 39044 6867 39056 6875
rect 39072 6867 39084 6875
rect 39104 6867 39116 6875
rect 39120 6867 39132 6875
rect 39136 6867 39148 6875
rect 39260 6867 39272 6875
rect 39292 6867 39304 6875
rect 39308 6867 39312 6875
rect 39324 6867 39336 6875
rect 39344 6867 39368 6875
rect 39384 6867 39408 6875
rect 39416 6867 39428 6875
rect 39436 6867 39460 6875
rect 39476 6867 39524 6875
rect 39540 6867 39556 6875
rect 39572 6867 39584 6875
rect 39596 6867 39600 6875
rect 39604 6867 39616 6875
rect 39636 6867 39648 6875
rect 39652 6867 39656 6875
rect 39668 6867 39680 6875
rect 39696 6867 39712 6875
rect 39728 6867 39776 6875
rect 39788 6867 39804 6875
rect 39820 6867 39868 6875
rect 39884 6867 39896 6875
rect 39912 6867 39960 6875
rect 39976 6867 39992 6875
rect 40008 6867 40020 6875
rect 40032 6867 40036 6875
rect 40040 6867 40052 6875
rect 40164 6867 40176 6875
rect 40180 6867 40192 6875
rect 40196 6867 40208 6875
rect 40228 6867 40240 6875
rect 40260 6867 40272 6875
rect 40292 6867 40304 6875
rect 40324 6867 40336 6875
rect 40340 6867 40352 6875
rect 40356 6867 40368 6875
rect 40480 6867 40492 6875
rect 40496 6867 40500 6875
rect 40664 6867 40676 6875
rect 40696 6867 40708 6875
rect 40712 6867 40716 6875
rect 40728 6867 40740 6875
rect 40748 6867 40772 6875
rect 40788 6867 40800 6875
rect 20234 6850 20236 6858
rect 20242 6850 20244 6858
rect 21514 6850 21518 6858
rect 21522 6850 21526 6858
rect 21720 6850 21732 6858
rect 22262 6850 22268 6858
rect 22270 6850 22276 6858
rect 22338 6850 22344 6858
rect 22346 6850 22352 6858
rect 22690 6850 22696 6858
rect 22698 6850 22704 6858
rect 22766 6850 22772 6858
rect 22774 6850 22780 6858
rect 23012 6850 23016 6858
rect 23020 6850 23024 6858
rect 23088 6850 23092 6858
rect 23096 6850 23100 6858
rect 23332 6850 23338 6858
rect 23340 6850 23346 6858
rect 23408 6850 23414 6858
rect 23416 6850 23422 6858
rect 23654 6850 23658 6858
rect 23662 6850 23666 6858
rect 23730 6850 23734 6858
rect 23738 6850 23742 6858
rect 23952 6850 23964 6858
rect 24158 6850 24162 6858
rect 24166 6850 24170 6858
rect 24372 6850 24376 6858
rect 24380 6850 24384 6858
rect 24586 6850 24590 6858
rect 24594 6850 24598 6858
rect 24998 6850 25002 6858
rect 25006 6850 25010 6858
rect 26052 6850 26056 6858
rect 26060 6850 26064 6858
rect 26258 6850 26270 6858
rect 26464 6850 26468 6858
rect 26472 6850 26476 6858
rect 26678 6850 26682 6858
rect 26686 6850 26690 6858
rect 27418 6850 27430 6858
rect 27434 6850 27438 6858
rect 27502 6850 27506 6858
rect 27510 6850 27514 6858
rect 27632 6850 27644 6858
rect 27708 6850 27720 6858
rect 28060 6850 28072 6858
rect 28136 6850 28148 6858
rect 34208 6857 34216 6865
rect 35024 6857 35032 6865
rect 20336 6840 20344 6848
rect 29712 6837 29720 6845
rect 32560 6837 32568 6845
rect 36912 6837 36920 6845
rect 26352 6820 26360 6828
rect 37680 6817 37688 6825
rect 37952 6817 37960 6825
rect 40032 6817 40040 6825
rect 28000 6800 28008 6808
rect 29392 6797 29400 6805
rect 35232 6797 35240 6805
rect 35632 6797 35640 6805
rect 37680 6797 37688 6805
rect 22736 6780 22744 6788
rect 25536 6780 25544 6788
rect 26416 6780 26424 6788
rect 27248 6780 27256 6788
rect 29536 6777 29544 6785
rect 30416 6777 30424 6785
rect 31536 6777 31544 6785
rect 31776 6777 31784 6785
rect 32928 6777 32936 6785
rect 33904 6777 33912 6785
rect 33984 6777 33992 6785
rect 37728 6777 37736 6785
rect 37856 6777 37864 6785
rect 38000 6777 38008 6785
rect 38032 6777 38040 6785
rect 38128 6777 38136 6785
rect 38448 6777 38456 6785
rect 38544 6777 38552 6785
rect 38816 6777 38824 6785
rect 38896 6777 38904 6785
rect 39008 6777 39016 6785
rect 39088 6777 39096 6785
rect 39664 6777 39672 6785
rect 39968 6777 39976 6785
rect 40400 6777 40408 6785
rect 40768 6777 40776 6785
rect 19072 6761 19082 6766
rect 19280 6760 19288 6768
rect 20096 6760 20104 6768
rect 20304 6760 20312 6768
rect 21150 6761 21160 6766
rect 21710 6761 21720 6766
rect 22113 6761 22114 6766
rect 22464 6760 22472 6768
rect 22752 6760 22760 6768
rect 23040 6760 23048 6768
rect 23648 6760 23656 6768
rect 23680 6760 23688 6768
rect 24112 6760 24120 6768
rect 24944 6760 24952 6768
rect 26208 6760 26216 6768
rect 27408 6761 27418 6766
rect 27442 6761 27452 6766
rect 18720 6740 18728 6748
rect 19888 6740 19896 6748
rect 20480 6740 20488 6748
rect 21888 6740 21896 6748
rect 22320 6740 22328 6748
rect 24896 6740 24904 6748
rect 25712 6740 25720 6748
rect 26000 6740 26008 6748
rect 30544 6737 30552 6745
rect 32208 6737 32216 6745
rect 33376 6737 33384 6745
rect 37936 6737 37944 6745
rect 38016 6737 38024 6745
rect 38656 6737 38664 6745
rect 39920 6737 39928 6745
rect 40688 6737 40696 6745
rect 18640 6720 18648 6728
rect 18736 6720 18744 6728
rect 19456 6720 19464 6728
rect 19680 6720 19688 6728
rect 22096 6720 22104 6728
rect 23488 6720 23496 6728
rect 23904 6720 23912 6728
rect 24096 6720 24104 6728
rect 24128 6720 24136 6728
rect 24960 6720 24968 6728
rect 26976 6720 26984 6728
rect 27808 6720 27816 6728
rect 28096 6720 28104 6728
rect 29792 6717 29800 6725
rect 29872 6717 29880 6725
rect 30192 6717 30200 6725
rect 31280 6717 31288 6725
rect 32256 6717 32264 6725
rect 32528 6717 32536 6725
rect 32592 6717 32600 6725
rect 33120 6717 33128 6725
rect 33616 6717 33624 6725
rect 33808 6717 33816 6725
rect 34096 6717 34104 6725
rect 34240 6717 34248 6725
rect 34736 6717 34744 6725
rect 34944 6717 34952 6725
rect 36032 6717 36040 6725
rect 36192 6717 36200 6725
rect 36352 6717 36360 6725
rect 36464 6717 36472 6725
rect 36720 6717 36728 6725
rect 37152 6717 37160 6725
rect 38112 6717 38120 6725
rect 18480 6700 18488 6708
rect 23216 6700 23224 6708
rect 24720 6700 24728 6708
rect 26576 6700 26584 6708
rect 26608 6700 26616 6708
rect 26624 6700 26632 6708
rect 32528 6697 32536 6705
rect 32656 6697 32664 6705
rect 33040 6697 33048 6705
rect 33056 6697 33064 6705
rect 33952 6697 33960 6705
rect 34064 6697 34072 6705
rect 34688 6697 34696 6705
rect 34752 6697 34760 6705
rect 35056 6697 35064 6705
rect 35200 6697 35208 6705
rect 36688 6697 36696 6705
rect 36864 6697 36872 6705
rect 37312 6697 37320 6705
rect 38928 6697 38936 6705
rect 39408 6697 39416 6705
rect 39712 6697 39720 6705
rect 40000 6697 40008 6705
rect 40304 6697 40312 6705
rect 19504 6680 19512 6688
rect 21344 6680 21352 6688
rect 22576 6680 22584 6688
rect 24272 6680 24280 6688
rect 25104 6680 25112 6688
rect 25568 6680 25576 6688
rect 25584 6680 25592 6688
rect 34736 6677 34744 6685
rect 39760 6677 39768 6685
rect 26784 6660 26792 6668
rect 29380 6667 29392 6675
rect 29412 6667 29424 6675
rect 29428 6667 29432 6675
rect 29448 6667 29464 6675
rect 29480 6667 29512 6675
rect 29528 6667 29532 6675
rect 29536 6667 29540 6675
rect 29556 6667 29588 6675
rect 29604 6667 29616 6675
rect 29636 6667 29648 6675
rect 29660 6667 29664 6675
rect 29668 6667 29672 6675
rect 29692 6667 29696 6675
rect 29700 6667 29704 6675
rect 29800 6667 29804 6675
rect 29808 6667 29812 6675
rect 29824 6667 29836 6675
rect 29840 6667 29844 6675
rect 29860 6667 29876 6675
rect 29892 6667 29908 6675
rect 29916 6667 29948 6675
rect 29956 6667 29968 6675
rect 29988 6667 30000 6675
rect 30012 6667 30016 6675
rect 30020 6667 30032 6675
rect 30052 6667 30064 6675
rect 30076 6667 30080 6675
rect 30084 6667 30096 6675
rect 30100 6667 30104 6675
rect 30144 6667 30156 6675
rect 30168 6667 30172 6675
rect 30176 6667 30188 6675
rect 30192 6667 30196 6675
rect 30208 6667 30220 6675
rect 30228 6667 30252 6675
rect 30268 6667 30292 6675
rect 30300 6667 30312 6675
rect 30324 6667 30328 6675
rect 30332 6667 30344 6675
rect 30360 6667 30400 6675
rect 30424 6667 30440 6675
rect 30456 6667 30460 6675
rect 30464 6667 30476 6675
rect 30488 6667 30492 6675
rect 30496 6667 30500 6675
rect 30520 6667 30524 6675
rect 30528 6667 30540 6675
rect 30544 6667 30556 6675
rect 30560 6667 30564 6675
rect 30584 6667 30588 6675
rect 30592 6667 30596 6675
rect 30612 6667 30616 6675
rect 30620 6667 30632 6675
rect 30636 6667 30648 6675
rect 30652 6667 30656 6675
rect 30676 6667 30680 6675
rect 30684 6667 30688 6675
rect 30704 6667 30720 6675
rect 30728 6667 30752 6675
rect 30768 6667 30780 6675
rect 30784 6667 30788 6675
rect 30800 6667 30812 6675
rect 30824 6667 30828 6675
rect 30832 6667 30844 6675
rect 30848 6667 30852 6675
rect 30864 6667 30876 6675
rect 30988 6667 31000 6675
rect 31004 6667 31008 6675
rect 31020 6667 31032 6675
rect 31048 6667 31064 6675
rect 31072 6667 31104 6675
rect 31112 6667 31128 6675
rect 31144 6667 31160 6675
rect 31176 6667 31180 6675
rect 31184 6667 31196 6675
rect 31208 6667 31212 6675
rect 31216 6667 31220 6675
rect 31332 6667 31336 6675
rect 31340 6667 31344 6675
rect 31424 6667 31428 6675
rect 31432 6667 31436 6675
rect 31456 6667 31460 6675
rect 31464 6667 31468 6675
rect 31480 6667 31492 6675
rect 31496 6667 31500 6675
rect 31516 6667 31540 6675
rect 31548 6667 31564 6675
rect 31572 6667 31596 6675
rect 31612 6667 31628 6675
rect 31644 6667 31656 6675
rect 31668 6667 31672 6675
rect 31676 6667 31688 6675
rect 31692 6667 31696 6675
rect 31736 6667 31748 6675
rect 31760 6667 31764 6675
rect 31768 6667 31780 6675
rect 31784 6667 31788 6675
rect 31800 6667 31812 6675
rect 31892 6667 31904 6675
rect 31924 6667 31936 6675
rect 31940 6667 31952 6675
rect 31956 6667 31968 6675
rect 31988 6667 32000 6675
rect 32260 6667 32264 6675
rect 32268 6667 32280 6675
rect 32284 6667 32288 6675
rect 32300 6667 32312 6675
rect 32424 6667 32436 6675
rect 32440 6667 32452 6675
rect 32456 6667 32468 6675
rect 32488 6667 32500 6675
rect 32504 6667 32508 6675
rect 32540 6667 32544 6675
rect 32548 6667 32560 6675
rect 32580 6667 32592 6675
rect 32596 6667 32608 6675
rect 32612 6667 32624 6675
rect 32644 6667 32656 6675
rect 32672 6667 32696 6675
rect 32704 6667 32720 6675
rect 32736 6667 32740 6675
rect 32744 6667 32748 6675
rect 32760 6667 32772 6675
rect 32776 6667 32788 6675
rect 32800 6667 32804 6675
rect 32808 6667 32812 6675
rect 32828 6667 32844 6675
rect 32852 6667 32864 6675
rect 32868 6667 32880 6675
rect 32892 6667 32896 6675
rect 32900 6667 32904 6675
rect 32924 6667 32928 6675
rect 32932 6667 32936 6675
rect 33000 6667 33004 6675
rect 33008 6667 33020 6675
rect 33032 6667 33036 6675
rect 33040 6667 33044 6675
rect 33056 6667 33068 6675
rect 33072 6667 33084 6675
rect 33096 6667 33100 6675
rect 33104 6667 33108 6675
rect 33124 6667 33140 6675
rect 33148 6667 33172 6675
rect 33188 6667 33200 6675
rect 33220 6667 33232 6675
rect 33236 6667 33248 6675
rect 33252 6667 33256 6675
rect 33276 6667 33280 6675
rect 33284 6667 33288 6675
rect 33336 6667 33340 6675
rect 33344 6667 33348 6675
rect 33368 6667 33372 6675
rect 33376 6667 33380 6675
rect 33392 6667 33404 6675
rect 33420 6667 33436 6675
rect 33444 6667 33460 6675
rect 33468 6667 33484 6675
rect 33500 6667 33512 6675
rect 33520 6667 33536 6675
rect 33544 6667 33560 6675
rect 33576 6667 33592 6675
rect 33608 6667 33612 6675
rect 33616 6667 33628 6675
rect 33648 6667 33660 6675
rect 33664 6667 33676 6675
rect 33680 6667 33692 6675
rect 33712 6667 33724 6675
rect 33728 6667 33732 6675
rect 33804 6667 33816 6675
rect 33836 6667 33848 6675
rect 33852 6667 33856 6675
rect 33868 6667 33880 6675
rect 33892 6667 33896 6675
rect 33900 6667 33904 6675
rect 33920 6667 33936 6675
rect 33944 6667 33956 6675
rect 33960 6667 33972 6675
rect 33992 6667 34004 6675
rect 34008 6667 34012 6675
rect 34028 6667 34032 6675
rect 34036 6667 34048 6675
rect 34068 6667 34080 6675
rect 34084 6667 34088 6675
rect 34100 6667 34112 6675
rect 34132 6667 34144 6675
rect 34164 6667 34176 6675
rect 34188 6667 34192 6675
rect 34196 6667 34208 6675
rect 34280 6667 34284 6675
rect 34288 6667 34300 6675
rect 34412 6667 34424 6675
rect 34428 6667 34432 6675
rect 34536 6667 34548 6675
rect 34552 6667 34556 6675
rect 34568 6667 34580 6675
rect 34592 6667 34596 6675
rect 34600 6667 34612 6675
rect 34616 6667 34620 6675
rect 34632 6667 34644 6675
rect 34944 6667 34956 6675
rect 34960 6667 34964 6675
rect 34976 6667 34988 6675
rect 34996 6667 35020 6675
rect 35036 6667 35084 6675
rect 35096 6667 35112 6675
rect 35128 6667 35176 6675
rect 35192 6667 35200 6675
rect 35224 6667 35236 6675
rect 35248 6667 35252 6675
rect 35256 6667 35268 6675
rect 35380 6667 35392 6675
rect 35396 6667 35400 6675
rect 35472 6667 35484 6675
rect 35504 6667 35516 6675
rect 35520 6667 35524 6675
rect 35536 6667 35548 6675
rect 35560 6667 35564 6675
rect 35568 6667 35580 6675
rect 35584 6667 35588 6675
rect 35600 6667 35612 6675
rect 35628 6667 35644 6675
rect 35660 6667 35684 6675
rect 35692 6667 35708 6675
rect 35716 6667 35728 6675
rect 35732 6667 35736 6675
rect 35752 6667 35776 6675
rect 35784 6667 35800 6675
rect 35808 6667 35840 6675
rect 35848 6667 35864 6675
rect 35880 6667 35884 6675
rect 35888 6667 35892 6675
rect 35912 6667 35916 6675
rect 35920 6667 35932 6675
rect 35944 6667 35948 6675
rect 35952 6667 35956 6675
rect 36036 6667 36040 6675
rect 36044 6667 36048 6675
rect 36060 6667 36072 6675
rect 36076 6667 36080 6675
rect 36128 6667 36132 6675
rect 36136 6667 36140 6675
rect 36152 6667 36164 6675
rect 36168 6667 36172 6675
rect 36332 6667 36336 6675
rect 36340 6667 36344 6675
rect 36356 6667 36368 6675
rect 36372 6667 36384 6675
rect 36396 6667 36400 6675
rect 36404 6667 36408 6675
rect 36424 6667 36440 6675
rect 36448 6667 36472 6675
rect 36488 6667 36500 6675
rect 36520 6667 36532 6675
rect 36536 6667 36548 6675
rect 36552 6667 36564 6675
rect 36584 6667 36596 6675
rect 36600 6667 36604 6675
rect 36708 6667 36720 6675
rect 36724 6667 36728 6675
rect 36740 6667 36752 6675
rect 36764 6667 36768 6675
rect 36772 6667 36784 6675
rect 36920 6667 36924 6675
rect 36928 6667 36940 6675
rect 36960 6667 36972 6675
rect 36976 6667 36988 6675
rect 36992 6667 37004 6675
rect 37244 6667 37256 6675
rect 37268 6667 37272 6675
rect 37276 6667 37288 6675
rect 37292 6667 37296 6675
rect 37336 6667 37348 6675
rect 37360 6667 37364 6675
rect 37368 6667 37380 6675
rect 37384 6667 37388 6675
rect 37524 6667 37536 6675
rect 37540 6667 37552 6675
rect 37556 6667 37568 6675
rect 37588 6667 37600 6675
rect 37604 6667 37616 6675
rect 37620 6667 37632 6675
rect 37652 6667 37664 6675
rect 37768 6667 37772 6675
rect 37776 6667 37788 6675
rect 37792 6667 37796 6675
rect 37808 6667 37820 6675
rect 37840 6667 37852 6675
rect 37856 6667 37860 6675
rect 37872 6667 37884 6675
rect 37900 6667 37916 6675
rect 37924 6667 37956 6675
rect 37964 6667 37976 6675
rect 37992 6667 38008 6675
rect 38016 6667 38048 6675
rect 38056 6667 38072 6675
rect 38088 6667 38100 6675
rect 38108 6667 38140 6675
rect 38148 6667 38164 6675
rect 38180 6667 38196 6675
rect 38212 6667 38216 6675
rect 38220 6667 38232 6675
rect 38244 6667 38248 6675
rect 38252 6667 38256 6675
rect 38304 6667 38308 6675
rect 38312 6667 38324 6675
rect 38336 6667 38340 6675
rect 38344 6667 38348 6675
rect 38360 6667 38372 6675
rect 38376 6667 38380 6675
rect 38428 6667 38432 6675
rect 38436 6667 38440 6675
rect 38452 6667 38464 6675
rect 38468 6667 38472 6675
rect 38568 6667 38572 6675
rect 38576 6667 38580 6675
rect 38592 6667 38604 6675
rect 38608 6667 38620 6675
rect 38632 6667 38636 6675
rect 38640 6667 38644 6675
rect 38664 6667 38668 6675
rect 38672 6667 38684 6675
rect 38696 6667 38700 6675
rect 38704 6667 38708 6675
rect 38788 6667 38792 6675
rect 38796 6667 38800 6675
rect 38820 6667 38824 6675
rect 38828 6667 38832 6675
rect 38844 6667 38856 6675
rect 38860 6667 38864 6675
rect 38880 6667 38896 6675
rect 38912 6667 38960 6675
rect 38976 6667 38988 6675
rect 38992 6667 38996 6675
rect 39008 6667 39020 6675
rect 39032 6667 39036 6675
rect 39040 6667 39052 6675
rect 39056 6667 39060 6675
rect 39124 6667 39128 6675
rect 39132 6667 39144 6675
rect 39148 6667 39152 6675
rect 39164 6667 39176 6675
rect 39188 6667 39192 6675
rect 39196 6667 39208 6675
rect 39224 6667 39248 6675
rect 39256 6667 39272 6675
rect 39288 6667 39312 6675
rect 39320 6667 39336 6675
rect 39344 6667 39368 6675
rect 39384 6667 39388 6675
rect 39392 6667 39404 6675
rect 39412 6667 39428 6675
rect 39436 6667 39460 6675
rect 39476 6667 39492 6675
rect 39500 6667 39524 6675
rect 39540 6667 39564 6675
rect 39572 6667 39584 6675
rect 39596 6667 39600 6675
rect 39604 6667 39616 6675
rect 39632 6667 39656 6675
rect 39664 6667 39680 6675
rect 39696 6667 39712 6675
rect 39728 6667 39732 6675
rect 39736 6667 39748 6675
rect 39752 6667 39764 6675
rect 39768 6667 39772 6675
rect 39788 6667 39804 6675
rect 39820 6667 39836 6675
rect 39844 6667 39868 6675
rect 39884 6667 39896 6675
rect 39900 6667 39904 6675
rect 39916 6667 39928 6675
rect 39936 6667 39960 6675
rect 39976 6667 40000 6675
rect 40008 6667 40020 6675
rect 40028 6667 40052 6675
rect 40068 6667 40080 6675
rect 40084 6667 40088 6675
rect 40100 6667 40112 6675
rect 40124 6667 40128 6675
rect 40132 6667 40144 6675
rect 40160 6667 40208 6675
rect 40224 6667 40240 6675
rect 40256 6667 40260 6675
rect 40264 6667 40276 6675
rect 40288 6667 40292 6675
rect 40296 6667 40300 6675
rect 40320 6667 40324 6675
rect 40328 6667 40340 6675
rect 40344 6667 40356 6675
rect 40360 6667 40364 6675
rect 40380 6667 40404 6675
rect 40412 6667 40428 6675
rect 40436 6667 40460 6675
rect 40476 6667 40492 6675
rect 40508 6667 40520 6675
rect 40532 6667 40536 6675
rect 40540 6667 40552 6675
rect 40556 6667 40560 6675
rect 40664 6667 40676 6675
rect 40696 6667 40708 6675
rect 40712 6667 40716 6675
rect 40728 6667 40740 6675
rect 40756 6667 40772 6675
rect 40780 6667 40800 6675
rect 20002 6656 20004 6660
rect 20008 6652 20010 6656
rect 20708 6650 20722 6658
rect 21120 6650 21134 6658
rect 21372 6650 21380 6658
rect 21524 6650 21530 6658
rect 21532 6650 21538 6658
rect 22720 6650 22734 6658
rect 23362 6650 23376 6658
rect 23718 6650 23724 6658
rect 23726 6650 23732 6658
rect 23876 6650 23882 6658
rect 23924 6650 23938 6658
rect 24138 6650 24152 6658
rect 25198 6650 25202 6658
rect 25288 6650 25296 6658
rect 25620 6656 25622 6660
rect 26316 6656 26318 6660
rect 25626 6652 25628 6656
rect 26322 6652 26324 6656
rect 26450 6650 26454 6658
rect 26540 6650 26548 6658
rect 26664 6650 26668 6658
rect 26754 6650 26762 6658
rect 28398 6652 28400 6660
rect 28648 6648 28652 6660
rect 29568 6637 29576 6645
rect 30000 6637 30008 6645
rect 32192 6637 32200 6645
rect 32416 6637 32424 6645
rect 32512 6637 32520 6645
rect 33936 6637 33944 6645
rect 34144 6637 34152 6645
rect 34192 6637 34200 6645
rect 34496 6637 34504 6645
rect 35248 6637 35256 6645
rect 35520 6637 35528 6645
rect 37536 6637 37544 6645
rect 37839 6638 37846 6643
rect 20976 6620 20984 6628
rect 24096 6620 24104 6628
rect 24928 6620 24936 6628
rect 26416 6620 26424 6628
rect 28432 6620 28440 6628
rect 29712 6617 29720 6625
rect 30400 6617 30408 6625
rect 30464 6617 30472 6625
rect 31648 6617 31656 6625
rect 32096 6617 32104 6625
rect 34928 6617 34936 6625
rect 35008 6617 35016 6625
rect 35056 6617 35064 6625
rect 35920 6617 35928 6625
rect 36816 6617 36824 6625
rect 38016 6617 38024 6625
rect 38080 6617 38088 6625
rect 38176 6617 38184 6625
rect 21360 6600 21368 6608
rect 22176 6600 22184 6608
rect 23488 6600 23496 6608
rect 29408 6597 29416 6605
rect 29504 6597 29512 6605
rect 29744 6597 29752 6605
rect 31072 6597 31080 6605
rect 31392 6597 31400 6605
rect 31664 6597 31672 6605
rect 32016 6597 32024 6605
rect 32768 6597 32776 6605
rect 33248 6597 33256 6605
rect 33296 6597 33304 6605
rect 33344 6597 33352 6605
rect 33472 6597 33480 6605
rect 33920 6597 33928 6605
rect 34320 6597 34328 6605
rect 34480 6597 34488 6605
rect 34528 6597 34536 6605
rect 35744 6597 35752 6605
rect 36656 6597 36664 6605
rect 36768 6597 36776 6605
rect 37664 6597 37672 6605
rect 37888 6597 37896 6605
rect 38288 6597 38296 6605
rect 38688 6597 38696 6605
rect 38848 6597 38856 6605
rect 39072 6597 39080 6605
rect 39440 6597 39448 6605
rect 39488 6597 39496 6605
rect 39792 6597 39800 6605
rect 39968 6597 39976 6605
rect 18528 6580 18536 6588
rect 19360 6580 19368 6588
rect 20320 6580 20328 6588
rect 20736 6580 20744 6588
rect 20832 6580 20840 6588
rect 21776 6580 21784 6588
rect 22848 6580 22856 6588
rect 23136 6580 23144 6588
rect 23568 6580 23576 6588
rect 26560 6580 26568 6588
rect 26880 6580 26888 6588
rect 27024 6580 27032 6588
rect 27888 6580 27896 6588
rect 28096 6580 28104 6588
rect 28288 6580 28296 6588
rect 30320 6577 30328 6585
rect 30464 6577 30472 6585
rect 34160 6577 34168 6585
rect 34512 6577 34520 6585
rect 37680 6577 37688 6585
rect 19952 6560 19960 6568
rect 24320 6560 24328 6568
rect 29392 6557 29400 6565
rect 29472 6557 29480 6565
rect 29968 6557 29976 6565
rect 31744 6557 31752 6565
rect 32752 6557 32760 6565
rect 33200 6557 33208 6565
rect 33376 6557 33384 6565
rect 33440 6557 33448 6565
rect 33568 6557 33576 6565
rect 33616 6557 33624 6565
rect 34304 6557 34312 6565
rect 34848 6557 34856 6565
rect 35216 6557 35224 6565
rect 36672 6557 36680 6565
rect 36944 6557 36952 6565
rect 38320 6557 38328 6565
rect 39680 6557 39688 6565
rect 40208 6557 40216 6565
rect 40704 6557 40712 6565
rect 19072 6548 19076 6553
rect 19540 6548 19544 6553
rect 18864 6540 18872 6548
rect 19792 6540 19800 6548
rect 19952 6540 19960 6548
rect 20816 6540 20824 6548
rect 21152 6540 21160 6548
rect 21360 6540 21368 6548
rect 21776 6540 21784 6548
rect 23552 6540 23560 6548
rect 23744 6540 23752 6548
rect 23936 6540 23944 6548
rect 25520 6540 25528 6548
rect 26016 6540 26024 6548
rect 26576 6540 26584 6548
rect 26864 6540 26872 6548
rect 28080 6540 28088 6548
rect 39072 6537 39080 6545
rect 40512 6537 40520 6545
rect 24784 6520 24792 6528
rect 27888 6520 27896 6528
rect 31696 6517 31704 6525
rect 33696 6517 33704 6525
rect 35792 6517 35800 6525
rect 24512 6500 24520 6508
rect 27824 6500 27832 6508
rect 36272 6497 36280 6505
rect 33760 6477 33768 6485
rect 34784 6477 34792 6485
rect 36336 6477 36344 6485
rect 36576 6477 36584 6485
rect 29372 6467 29376 6475
rect 29380 6467 29384 6475
rect 29404 6467 29408 6475
rect 29412 6467 29416 6475
rect 29428 6467 29440 6475
rect 29456 6467 29472 6475
rect 29488 6467 29520 6475
rect 29528 6467 29544 6475
rect 29560 6467 29572 6475
rect 29576 6467 29588 6475
rect 29592 6467 29596 6475
rect 29716 6467 29728 6475
rect 29732 6467 29744 6475
rect 29748 6467 29760 6475
rect 29780 6467 29792 6475
rect 29808 6467 29832 6475
rect 29840 6467 29856 6475
rect 29872 6467 29876 6475
rect 29880 6467 29884 6475
rect 29896 6467 29908 6475
rect 29912 6467 29924 6475
rect 29936 6467 29940 6475
rect 29944 6467 29948 6475
rect 30028 6467 30032 6475
rect 30036 6467 30040 6475
rect 30052 6467 30064 6475
rect 30068 6467 30080 6475
rect 30092 6467 30096 6475
rect 30100 6467 30104 6475
rect 30248 6467 30252 6475
rect 30256 6467 30260 6475
rect 30280 6467 30284 6475
rect 30288 6467 30292 6475
rect 30372 6467 30376 6475
rect 30380 6467 30392 6475
rect 30396 6467 30408 6475
rect 30412 6467 30416 6475
rect 30436 6467 30440 6475
rect 30444 6467 30448 6475
rect 30464 6467 30480 6475
rect 30488 6467 30512 6475
rect 30528 6467 30576 6475
rect 30592 6467 30608 6475
rect 30624 6467 30628 6475
rect 30632 6467 30644 6475
rect 30656 6467 30660 6475
rect 30664 6467 30668 6475
rect 30688 6467 30692 6475
rect 30696 6467 30700 6475
rect 30764 6467 30768 6475
rect 30772 6467 30784 6475
rect 30796 6467 30800 6475
rect 30804 6467 30808 6475
rect 30820 6467 30832 6475
rect 30836 6467 30840 6475
rect 30888 6467 30892 6475
rect 30896 6467 30900 6475
rect 30912 6467 30924 6475
rect 30928 6467 30932 6475
rect 30980 6467 30984 6475
rect 30988 6467 30992 6475
rect 31040 6467 31044 6475
rect 31048 6467 31060 6475
rect 31072 6467 31076 6475
rect 31080 6467 31084 6475
rect 31096 6467 31108 6475
rect 31112 6467 31116 6475
rect 31136 6467 31140 6475
rect 31144 6467 31148 6475
rect 31164 6467 31180 6475
rect 31188 6467 31220 6475
rect 31228 6467 31240 6475
rect 31256 6467 31272 6475
rect 31280 6467 31312 6475
rect 31320 6467 31336 6475
rect 31352 6467 31364 6475
rect 31372 6467 31404 6475
rect 31412 6467 31428 6475
rect 31444 6467 31448 6475
rect 31452 6467 31456 6475
rect 31476 6467 31480 6475
rect 31484 6467 31496 6475
rect 31508 6467 31512 6475
rect 31516 6467 31520 6475
rect 31532 6467 31544 6475
rect 31548 6467 31552 6475
rect 31728 6467 31732 6475
rect 31736 6467 31748 6475
rect 31760 6467 31764 6475
rect 31768 6467 31772 6475
rect 31784 6467 31796 6475
rect 31800 6467 31804 6475
rect 32012 6467 32016 6475
rect 32020 6467 32024 6475
rect 32036 6467 32048 6475
rect 32052 6467 32056 6475
rect 32136 6467 32140 6475
rect 32144 6467 32148 6475
rect 32168 6467 32172 6475
rect 32176 6467 32180 6475
rect 32192 6467 32204 6475
rect 32208 6467 32212 6475
rect 32232 6467 32236 6475
rect 32240 6467 32252 6475
rect 32256 6467 32268 6475
rect 32272 6467 32276 6475
rect 32296 6467 32300 6475
rect 32304 6467 32316 6475
rect 32324 6467 32340 6475
rect 32348 6467 32360 6475
rect 32364 6467 32368 6475
rect 32388 6467 32392 6475
rect 32396 6467 32408 6475
rect 32416 6467 32432 6475
rect 32440 6467 32464 6475
rect 32480 6467 32484 6475
rect 32488 6467 32500 6475
rect 32504 6467 32516 6475
rect 32520 6467 32524 6475
rect 32540 6467 32544 6475
rect 32548 6467 32552 6475
rect 32572 6467 32576 6475
rect 32580 6467 32592 6475
rect 32596 6467 32608 6475
rect 32612 6467 32616 6475
rect 32636 6467 32640 6475
rect 32644 6467 32648 6475
rect 32664 6467 32668 6475
rect 32672 6467 32684 6475
rect 32688 6467 32700 6475
rect 32704 6467 32708 6475
rect 32724 6467 32728 6475
rect 32732 6467 32736 6475
rect 32756 6467 32760 6475
rect 32764 6467 32776 6475
rect 32780 6467 32792 6475
rect 32796 6467 32800 6475
rect 32848 6467 32852 6475
rect 32856 6467 32868 6475
rect 32872 6467 32876 6475
rect 32888 6467 32900 6475
rect 32920 6467 32932 6475
rect 32948 6467 32972 6475
rect 32980 6467 32996 6475
rect 33004 6467 33016 6475
rect 33036 6467 33048 6475
rect 33052 6467 33064 6475
rect 33076 6467 33080 6475
rect 33084 6467 33088 6475
rect 33104 6467 33120 6475
rect 33128 6467 33140 6475
rect 33152 6467 33156 6475
rect 33160 6467 33172 6475
rect 33300 6467 33312 6475
rect 33316 6467 33328 6475
rect 33336 6467 33352 6475
rect 33368 6467 33384 6475
rect 33392 6467 33404 6475
rect 33412 6467 33436 6475
rect 33452 6467 33476 6475
rect 33492 6467 33496 6475
rect 33500 6467 33512 6475
rect 33520 6467 33536 6475
rect 33544 6467 33560 6475
rect 33576 6467 33592 6475
rect 33608 6467 33612 6475
rect 33616 6467 33628 6475
rect 33648 6467 33660 6475
rect 33664 6467 33676 6475
rect 33680 6467 33692 6475
rect 33708 6467 33724 6475
rect 33740 6467 33752 6475
rect 33756 6467 33768 6475
rect 33772 6467 33784 6475
rect 33832 6467 33844 6475
rect 33848 6467 33860 6475
rect 33864 6467 33876 6475
rect 33896 6467 33908 6475
rect 34028 6467 34032 6475
rect 34036 6467 34040 6475
rect 34168 6467 34172 6475
rect 34176 6467 34180 6475
rect 34192 6467 34204 6475
rect 34208 6467 34212 6475
rect 34232 6467 34236 6475
rect 34240 6467 34252 6475
rect 34256 6467 34268 6475
rect 34272 6467 34276 6475
rect 34404 6467 34408 6475
rect 34412 6467 34424 6475
rect 34428 6467 34440 6475
rect 34444 6467 34448 6475
rect 34468 6467 34472 6475
rect 34476 6467 34488 6475
rect 34500 6467 34504 6475
rect 34508 6467 34512 6475
rect 34532 6467 34536 6475
rect 34540 6467 34544 6475
rect 34608 6467 34612 6475
rect 34616 6467 34620 6475
rect 34640 6467 34644 6475
rect 34648 6467 34652 6475
rect 34700 6467 34704 6475
rect 34708 6467 34712 6475
rect 34732 6467 34736 6475
rect 34740 6467 34752 6475
rect 34756 6467 34768 6475
rect 34788 6467 34800 6475
rect 34804 6467 34808 6475
rect 34840 6467 34844 6475
rect 34848 6467 34860 6475
rect 34880 6467 34892 6475
rect 34896 6467 34900 6475
rect 34912 6467 34924 6475
rect 34944 6467 34956 6475
rect 34972 6467 35020 6475
rect 35036 6467 35040 6475
rect 35044 6467 35048 6475
rect 35060 6467 35072 6475
rect 35076 6467 35088 6475
rect 35096 6467 35112 6475
rect 35128 6467 35144 6475
rect 35152 6467 35176 6475
rect 35192 6467 35200 6475
rect 35224 6467 35236 6475
rect 35240 6467 35252 6475
rect 35256 6467 35268 6475
rect 35284 6467 35296 6475
rect 35316 6467 35328 6475
rect 35332 6467 35344 6475
rect 35348 6467 35360 6475
rect 35380 6467 35392 6475
rect 35472 6467 35484 6475
rect 35496 6467 35500 6475
rect 35504 6467 35516 6475
rect 35520 6467 35524 6475
rect 35536 6467 35548 6475
rect 35720 6467 35732 6475
rect 35744 6467 35748 6475
rect 35752 6467 35764 6475
rect 35768 6467 35772 6475
rect 35784 6467 35796 6475
rect 35808 6467 35812 6475
rect 35816 6467 35828 6475
rect 35832 6467 35836 6475
rect 35848 6467 35860 6475
rect 35876 6467 35892 6475
rect 35908 6467 35932 6475
rect 35940 6467 35956 6475
rect 35964 6467 35976 6475
rect 35980 6467 35984 6475
rect 36004 6467 36008 6475
rect 36012 6467 36024 6475
rect 36028 6467 36040 6475
rect 36044 6467 36048 6475
rect 36068 6467 36072 6475
rect 36076 6467 36080 6475
rect 36176 6467 36180 6475
rect 36184 6467 36188 6475
rect 36200 6467 36212 6475
rect 36216 6467 36220 6475
rect 36240 6467 36244 6475
rect 36248 6467 36252 6475
rect 36264 6467 36276 6475
rect 36280 6467 36284 6475
rect 36304 6467 36308 6475
rect 36312 6467 36324 6475
rect 36332 6467 36348 6475
rect 36356 6467 36368 6475
rect 36372 6467 36376 6475
rect 36396 6467 36400 6475
rect 36404 6467 36416 6475
rect 36424 6467 36440 6475
rect 36448 6467 36472 6475
rect 36488 6467 36500 6475
rect 36520 6467 36532 6475
rect 36544 6467 36548 6475
rect 36552 6467 36564 6475
rect 36568 6467 36572 6475
rect 36584 6467 36596 6475
rect 36676 6467 36688 6475
rect 36928 6467 36940 6475
rect 36960 6467 36972 6475
rect 36976 6467 36980 6475
rect 36992 6467 37004 6475
rect 37024 6467 37036 6475
rect 37040 6467 37052 6475
rect 37056 6467 37068 6475
rect 37300 6467 37304 6475
rect 37308 6467 37320 6475
rect 37392 6467 37396 6475
rect 37400 6467 37412 6475
rect 37648 6467 37660 6475
rect 37664 6467 37668 6475
rect 37680 6467 37692 6475
rect 37712 6467 37724 6475
rect 37740 6467 37788 6475
rect 37804 6467 37808 6475
rect 37812 6467 37816 6475
rect 37836 6467 37840 6475
rect 37844 6467 37856 6475
rect 37868 6467 37872 6475
rect 37876 6467 37880 6475
rect 37900 6467 37904 6475
rect 37908 6467 37912 6475
rect 37960 6467 37964 6475
rect 37968 6467 37972 6475
rect 37992 6467 37996 6475
rect 38000 6467 38012 6475
rect 38016 6467 38028 6475
rect 38032 6467 38036 6475
rect 38056 6467 38060 6475
rect 38064 6467 38076 6475
rect 38084 6467 38100 6475
rect 38108 6467 38120 6475
rect 38124 6467 38128 6475
rect 38148 6467 38152 6475
rect 38156 6467 38168 6475
rect 38180 6467 38184 6475
rect 38188 6467 38192 6475
rect 38212 6467 38216 6475
rect 38220 6467 38224 6475
rect 38304 6467 38308 6475
rect 38312 6467 38316 6475
rect 38380 6467 38384 6475
rect 38388 6467 38392 6475
rect 38412 6467 38416 6475
rect 38420 6467 38424 6475
rect 38472 6467 38476 6475
rect 38480 6467 38484 6475
rect 38504 6467 38508 6475
rect 38512 6467 38516 6475
rect 38528 6467 38540 6475
rect 38544 6467 38548 6475
rect 38568 6467 38572 6475
rect 38576 6467 38580 6475
rect 38596 6467 38644 6475
rect 38660 6467 38684 6475
rect 38692 6467 38704 6475
rect 38712 6467 38736 6475
rect 38752 6467 38776 6475
rect 38784 6467 38796 6475
rect 38808 6467 38812 6475
rect 38816 6467 38828 6475
rect 38848 6467 38860 6475
rect 38872 6467 38876 6475
rect 38880 6467 38892 6475
rect 38912 6467 38924 6475
rect 38928 6467 38932 6475
rect 39036 6467 39048 6475
rect 39052 6467 39064 6475
rect 39068 6467 39080 6475
rect 39100 6467 39112 6475
rect 39128 6467 39140 6475
rect 39144 6467 39156 6475
rect 39160 6467 39172 6475
rect 39188 6467 39200 6475
rect 39220 6467 39232 6475
rect 39236 6467 39248 6475
rect 39252 6467 39264 6475
rect 39284 6467 39296 6475
rect 39304 6467 39336 6475
rect 39344 6467 39360 6475
rect 39376 6467 39388 6475
rect 39396 6467 39428 6475
rect 39436 6467 39452 6475
rect 39468 6467 39492 6475
rect 39500 6467 39516 6475
rect 39532 6467 39536 6475
rect 39540 6467 39544 6475
rect 39556 6467 39568 6475
rect 39572 6467 39584 6475
rect 39596 6467 39600 6475
rect 39604 6467 39608 6475
rect 39624 6467 39628 6475
rect 39632 6467 39636 6475
rect 39648 6467 39660 6475
rect 39664 6467 39676 6475
rect 39688 6467 39692 6475
rect 39696 6467 39700 6475
rect 39716 6467 39720 6475
rect 39724 6467 39728 6475
rect 39740 6467 39752 6475
rect 39756 6467 39768 6475
rect 39780 6467 39784 6475
rect 39788 6467 39792 6475
rect 39888 6467 39892 6475
rect 39896 6467 39908 6475
rect 39920 6467 39924 6475
rect 39928 6467 39932 6475
rect 40028 6467 40032 6475
rect 40036 6467 40040 6475
rect 40060 6467 40064 6475
rect 40068 6467 40072 6475
rect 40084 6467 40096 6475
rect 40100 6467 40112 6475
rect 40124 6467 40128 6475
rect 40132 6467 40136 6475
rect 40152 6467 40200 6475
rect 40216 6467 40232 6475
rect 40248 6467 40260 6475
rect 40272 6467 40276 6475
rect 40280 6467 40292 6475
rect 40312 6467 40324 6475
rect 40328 6467 40340 6475
rect 40344 6467 40356 6475
rect 40376 6467 40388 6475
rect 40396 6467 40428 6475
rect 40436 6467 40452 6475
rect 40468 6467 40492 6475
rect 40500 6467 40516 6475
rect 40532 6467 40580 6475
rect 40596 6467 40612 6475
rect 40620 6467 40632 6475
rect 40636 6467 40648 6475
rect 40660 6467 40664 6475
rect 40668 6467 40672 6475
rect 18472 6448 18476 6460
rect 18570 6450 18572 6458
rect 18578 6450 18580 6458
rect 24656 6450 24666 6458
rect 25258 6450 25260 6458
rect 25266 6450 25268 6458
rect 25464 6450 25474 6458
rect 25678 6450 25688 6458
rect 26518 6450 26528 6458
rect 28128 6450 28132 6458
rect 28136 6450 28140 6458
rect 28334 6450 28346 6458
rect 38000 6457 38008 6465
rect 38992 6457 39000 6465
rect 30544 6437 30552 6445
rect 35808 6437 35816 6445
rect 20960 6420 20968 6428
rect 30336 6417 30344 6425
rect 31456 6417 31464 6425
rect 32432 6417 32440 6425
rect 33952 6417 33960 6425
rect 34752 6417 34760 6425
rect 35008 6417 35016 6425
rect 39776 6417 39784 6425
rect 40400 6417 40408 6425
rect 21536 6400 21544 6408
rect 39488 6397 39496 6405
rect 22512 6380 22520 6388
rect 27264 6380 27272 6388
rect 30272 6377 30280 6385
rect 31200 6377 31208 6385
rect 32032 6377 32040 6385
rect 33072 6377 33080 6385
rect 33520 6377 33528 6385
rect 34064 6377 34072 6385
rect 34512 6377 34520 6385
rect 36096 6377 36104 6385
rect 36672 6377 36680 6385
rect 37344 6377 37352 6385
rect 37360 6377 37368 6385
rect 37440 6377 37448 6385
rect 37696 6377 37704 6385
rect 37808 6377 37816 6385
rect 37888 6377 37896 6385
rect 38128 6377 38136 6385
rect 38800 6377 38808 6385
rect 39200 6377 39208 6385
rect 40576 6377 40584 6385
rect 18640 6360 18648 6368
rect 18704 6360 18712 6368
rect 19120 6360 19128 6368
rect 19552 6360 19560 6368
rect 20352 6360 20360 6368
rect 21120 6360 21128 6368
rect 22416 6360 22424 6368
rect 22688 6360 22696 6368
rect 23056 6360 23064 6368
rect 23120 6360 23128 6368
rect 23472 6360 23480 6368
rect 23486 6361 23496 6366
rect 24528 6360 24536 6368
rect 25844 6361 25847 6366
rect 26400 6360 26408 6368
rect 26832 6360 26840 6368
rect 31872 6357 31880 6365
rect 33200 6357 33208 6365
rect 34080 6357 34088 6365
rect 34304 6357 34312 6365
rect 36236 6364 36238 6365
rect 36236 6357 36238 6358
rect 40464 6357 40472 6365
rect 27648 6340 27656 6348
rect 29984 6337 29992 6345
rect 30304 6337 30312 6345
rect 31072 6337 31080 6345
rect 31280 6337 31288 6345
rect 31632 6337 31640 6345
rect 31680 6337 31688 6345
rect 32016 6337 32024 6345
rect 32128 6337 32136 6345
rect 32176 6337 32184 6345
rect 32416 6337 32424 6345
rect 32752 6337 32760 6345
rect 32912 6337 32920 6345
rect 33216 6337 33224 6345
rect 34912 6337 34920 6345
rect 35136 6337 35144 6345
rect 35504 6337 35512 6345
rect 35872 6337 35880 6345
rect 36384 6337 36392 6345
rect 36704 6337 36712 6345
rect 36976 6337 36984 6345
rect 37376 6337 37384 6345
rect 37680 6337 37688 6345
rect 39344 6337 39352 6345
rect 19728 6320 19736 6328
rect 19760 6320 19768 6328
rect 19904 6320 19912 6328
rect 21104 6320 21112 6328
rect 21200 6320 21208 6328
rect 23504 6320 23512 6328
rect 23984 6320 23992 6328
rect 24224 6320 24232 6328
rect 24368 6320 24376 6328
rect 25200 6320 25208 6328
rect 25296 6320 25304 6328
rect 25856 6320 25864 6328
rect 26032 6320 26040 6328
rect 26064 6320 26072 6328
rect 26480 6320 26488 6328
rect 27952 6320 27960 6328
rect 29424 6317 29432 6325
rect 29488 6317 29496 6325
rect 29792 6317 29800 6325
rect 29808 6317 29816 6325
rect 29872 6317 29880 6325
rect 30160 6317 30168 6325
rect 32960 6317 32968 6325
rect 33216 6317 33224 6325
rect 33648 6317 33656 6325
rect 35200 6317 35208 6325
rect 35376 6317 35384 6325
rect 35488 6317 35496 6325
rect 36048 6317 36056 6325
rect 36176 6317 36184 6325
rect 36848 6317 36856 6325
rect 36992 6317 37000 6325
rect 21376 6300 21384 6308
rect 21632 6300 21640 6308
rect 22880 6300 22888 6308
rect 24784 6300 24792 6308
rect 28384 6300 28392 6308
rect 30144 6297 30152 6305
rect 30656 6297 30664 6305
rect 31184 6297 31192 6305
rect 31936 6297 31944 6305
rect 36464 6297 36472 6305
rect 37248 6297 37256 6305
rect 37952 6297 37960 6305
rect 18912 6280 18920 6288
rect 22896 6280 22904 6288
rect 23296 6280 23304 6288
rect 23920 6280 23928 6288
rect 30784 6277 30792 6285
rect 33904 6277 33912 6285
rect 35584 6277 35592 6285
rect 38288 6277 38296 6285
rect 38336 6277 38344 6285
rect 18880 6260 18888 6268
rect 19504 6260 19512 6268
rect 20944 6260 20952 6268
rect 26672 6260 26680 6268
rect 27472 6260 27480 6268
rect 29396 6267 29408 6275
rect 29428 6267 29440 6275
rect 29444 6267 29448 6275
rect 29460 6267 29472 6275
rect 29488 6267 29504 6275
rect 29512 6267 29544 6275
rect 29552 6267 29568 6275
rect 29576 6267 29588 6275
rect 29592 6267 29596 6275
rect 29616 6267 29620 6275
rect 29624 6267 29636 6275
rect 29648 6267 29652 6275
rect 29656 6267 29660 6275
rect 29788 6267 29792 6275
rect 29796 6267 29800 6275
rect 29812 6267 29824 6275
rect 29828 6267 29832 6275
rect 29852 6267 29856 6275
rect 29860 6267 29864 6275
rect 29880 6267 29928 6275
rect 29944 6267 29956 6275
rect 29960 6267 29964 6275
rect 29976 6267 29988 6275
rect 30000 6267 30004 6275
rect 30008 6267 30020 6275
rect 30036 6267 30048 6275
rect 30052 6267 30056 6275
rect 30068 6267 30080 6275
rect 30092 6267 30096 6275
rect 30100 6267 30112 6275
rect 30132 6267 30144 6275
rect 30156 6267 30160 6275
rect 30164 6267 30176 6275
rect 30248 6267 30252 6275
rect 30256 6267 30268 6275
rect 30380 6267 30392 6275
rect 30396 6267 30400 6275
rect 30412 6267 30424 6275
rect 30444 6267 30456 6275
rect 30472 6267 30520 6275
rect 30536 6267 30548 6275
rect 30552 6267 30556 6275
rect 30568 6267 30580 6275
rect 30592 6267 30596 6275
rect 30600 6267 30612 6275
rect 30632 6267 30644 6275
rect 30756 6267 30768 6275
rect 30772 6267 30784 6275
rect 30788 6267 30800 6275
rect 30820 6267 30832 6275
rect 30836 6267 30840 6275
rect 30944 6267 30956 6275
rect 30960 6267 30964 6275
rect 30976 6267 30988 6275
rect 30996 6267 31020 6275
rect 31036 6267 31048 6275
rect 31052 6267 31056 6275
rect 31068 6267 31080 6275
rect 31092 6267 31096 6275
rect 31100 6267 31112 6275
rect 31248 6267 31252 6275
rect 31256 6267 31268 6275
rect 31288 6267 31300 6275
rect 31304 6267 31308 6275
rect 31380 6267 31392 6275
rect 31396 6267 31408 6275
rect 31412 6267 31424 6275
rect 31440 6267 31456 6275
rect 31472 6267 31484 6275
rect 31488 6267 31500 6275
rect 31504 6267 31516 6275
rect 31536 6267 31548 6275
rect 31564 6267 31588 6275
rect 31596 6267 31612 6275
rect 31628 6267 31644 6275
rect 31652 6267 31676 6275
rect 31692 6267 31708 6275
rect 31716 6267 31748 6275
rect 31756 6267 31768 6275
rect 31788 6267 31800 6275
rect 31808 6267 31840 6275
rect 31848 6267 31864 6275
rect 31872 6267 31896 6275
rect 31912 6267 31924 6275
rect 31944 6267 31956 6275
rect 31968 6267 31972 6275
rect 31976 6267 31988 6275
rect 31992 6267 31996 6275
rect 32060 6267 32064 6275
rect 32068 6267 32080 6275
rect 32084 6267 32088 6275
rect 32100 6267 32112 6275
rect 32224 6267 32236 6275
rect 32240 6267 32252 6275
rect 32256 6267 32268 6275
rect 32288 6267 32300 6275
rect 32308 6267 32340 6275
rect 32348 6267 32360 6275
rect 32380 6267 32392 6275
rect 32396 6267 32408 6275
rect 32412 6267 32424 6275
rect 32444 6267 32456 6275
rect 32536 6267 32548 6275
rect 32560 6267 32564 6275
rect 32568 6267 32580 6275
rect 32584 6267 32588 6275
rect 32600 6267 32612 6275
rect 32624 6267 32628 6275
rect 32632 6267 32644 6275
rect 32660 6267 32684 6275
rect 32692 6267 32708 6275
rect 32724 6267 32728 6275
rect 32732 6267 32736 6275
rect 32756 6267 32760 6275
rect 32764 6267 32776 6275
rect 32780 6267 32792 6275
rect 32840 6267 32852 6275
rect 32856 6267 32868 6275
rect 32888 6267 32900 6275
rect 32916 6267 32940 6275
rect 32956 6267 32968 6275
rect 32988 6267 33000 6275
rect 33004 6267 33016 6275
rect 33036 6267 33048 6275
rect 33052 6267 33056 6275
rect 33228 6267 33232 6275
rect 33236 6267 33240 6275
rect 33252 6267 33264 6275
rect 33268 6267 33280 6275
rect 33300 6267 33312 6275
rect 33320 6267 33352 6275
rect 33360 6267 33376 6275
rect 33392 6267 33404 6275
rect 33416 6267 33420 6275
rect 33424 6267 33436 6275
rect 33456 6267 33468 6275
rect 33612 6267 33624 6275
rect 33644 6267 33656 6275
rect 33660 6267 33672 6275
rect 33676 6267 33688 6275
rect 33800 6267 33812 6275
rect 33816 6267 33820 6275
rect 33892 6267 33904 6275
rect 33908 6267 33912 6275
rect 33924 6267 33936 6275
rect 33956 6267 33968 6275
rect 33984 6267 34032 6275
rect 34048 6267 34060 6275
rect 34080 6267 34092 6275
rect 34104 6267 34108 6275
rect 34112 6267 34124 6275
rect 34144 6267 34156 6275
rect 34160 6267 34164 6275
rect 34260 6267 34264 6275
rect 34268 6267 34280 6275
rect 34300 6267 34312 6275
rect 34316 6267 34320 6275
rect 34332 6267 34344 6275
rect 34360 6267 34376 6275
rect 34400 6267 34440 6275
rect 34456 6267 34472 6275
rect 34480 6267 34492 6275
rect 34496 6267 34508 6275
rect 34520 6267 34524 6275
rect 34528 6267 34532 6275
rect 34548 6267 34564 6275
rect 34572 6267 34596 6275
rect 34612 6267 34624 6275
rect 34644 6267 34656 6275
rect 34660 6267 34672 6275
rect 34676 6267 34688 6275
rect 34840 6267 34844 6275
rect 34848 6267 34852 6275
rect 34872 6267 34876 6275
rect 34880 6267 34892 6275
rect 34896 6267 34908 6275
rect 34912 6267 34916 6275
rect 34936 6267 34940 6275
rect 34944 6267 34948 6275
rect 34964 6267 34968 6275
rect 34972 6267 34984 6275
rect 34988 6267 35000 6275
rect 35004 6267 35008 6275
rect 35024 6267 35040 6275
rect 35056 6267 35060 6275
rect 35064 6267 35076 6275
rect 35080 6267 35092 6275
rect 35096 6267 35100 6275
rect 35120 6267 35124 6275
rect 35128 6267 35140 6275
rect 35152 6267 35156 6275
rect 35160 6267 35164 6275
rect 35184 6267 35188 6275
rect 35192 6267 35196 6275
rect 35276 6267 35280 6275
rect 35284 6267 35288 6275
rect 35384 6267 35388 6275
rect 35392 6267 35396 6275
rect 35408 6267 35420 6275
rect 35424 6267 35428 6275
rect 35444 6267 35460 6275
rect 35476 6267 35524 6275
rect 35540 6267 35556 6275
rect 35572 6267 35576 6275
rect 35580 6267 35592 6275
rect 35604 6267 35608 6275
rect 35612 6267 35616 6275
rect 35792 6267 35796 6275
rect 35800 6267 35812 6275
rect 35816 6267 35828 6275
rect 35832 6267 35836 6275
rect 35856 6267 35860 6275
rect 35864 6267 35868 6275
rect 35884 6267 35900 6275
rect 35908 6267 35932 6275
rect 35948 6267 35960 6275
rect 35964 6267 35968 6275
rect 35980 6267 35992 6275
rect 36004 6267 36008 6275
rect 36012 6267 36024 6275
rect 36028 6267 36032 6275
rect 36044 6267 36056 6275
rect 36068 6267 36072 6275
rect 36076 6267 36088 6275
rect 36092 6267 36096 6275
rect 36200 6267 36212 6275
rect 36232 6267 36244 6275
rect 36248 6267 36252 6275
rect 36264 6267 36276 6275
rect 36292 6267 36308 6275
rect 36316 6267 36348 6275
rect 36356 6267 36368 6275
rect 36388 6267 36400 6275
rect 36408 6267 36440 6275
rect 36448 6267 36464 6275
rect 36480 6267 36484 6275
rect 36488 6267 36492 6275
rect 36512 6267 36516 6275
rect 36520 6267 36532 6275
rect 36544 6267 36548 6275
rect 36552 6267 36556 6275
rect 36568 6267 36580 6275
rect 36584 6267 36596 6275
rect 36608 6267 36612 6275
rect 36616 6267 36620 6275
rect 36668 6267 36672 6275
rect 36676 6267 36688 6275
rect 36700 6267 36704 6275
rect 36708 6267 36712 6275
rect 36724 6267 36736 6275
rect 36740 6267 36744 6275
rect 36840 6267 36844 6275
rect 36848 6267 36852 6275
rect 36864 6267 36876 6275
rect 36880 6267 36892 6275
rect 36904 6267 36908 6275
rect 36912 6267 36916 6275
rect 36932 6267 36948 6275
rect 36956 6267 36980 6275
rect 36996 6267 37008 6275
rect 37028 6267 37040 6275
rect 37044 6267 37056 6275
rect 37060 6267 37072 6275
rect 37088 6267 37104 6275
rect 37120 6267 37132 6275
rect 37136 6267 37148 6275
rect 37152 6267 37164 6275
rect 37184 6267 37196 6275
rect 37208 6267 37212 6275
rect 37216 6267 37228 6275
rect 37340 6267 37352 6275
rect 37432 6267 37444 6275
rect 37464 6267 37476 6275
rect 37480 6267 37484 6275
rect 37496 6267 37508 6275
rect 37524 6267 37540 6275
rect 37548 6267 37580 6275
rect 37588 6267 37600 6275
rect 37612 6267 37636 6275
rect 37652 6267 37656 6275
rect 37660 6267 37672 6275
rect 37684 6267 37688 6275
rect 37692 6267 37696 6275
rect 37716 6267 37720 6275
rect 37724 6267 37728 6275
rect 37792 6267 37796 6275
rect 37800 6267 37804 6275
rect 37824 6267 37828 6275
rect 37832 6267 37836 6275
rect 37848 6267 37860 6275
rect 37864 6267 37868 6275
rect 37888 6267 37892 6275
rect 37896 6267 37900 6275
rect 37916 6267 37964 6275
rect 37980 6267 37984 6275
rect 37988 6267 37992 6275
rect 38004 6267 38016 6275
rect 38020 6267 38032 6275
rect 38044 6267 38048 6275
rect 38052 6267 38056 6275
rect 38068 6267 38080 6275
rect 38084 6267 38088 6275
rect 38104 6267 38108 6275
rect 38112 6267 38124 6275
rect 38136 6267 38140 6275
rect 38144 6267 38148 6275
rect 38228 6267 38232 6275
rect 38236 6267 38240 6275
rect 38252 6267 38264 6275
rect 38268 6267 38272 6275
rect 38292 6267 38296 6275
rect 38300 6267 38304 6275
rect 38320 6267 38336 6275
rect 38344 6267 38376 6275
rect 38384 6267 38396 6275
rect 38416 6267 38428 6275
rect 38432 6267 38444 6275
rect 38448 6267 38460 6275
rect 38604 6267 38616 6275
rect 38620 6267 38624 6275
rect 38636 6267 38648 6275
rect 38660 6267 38664 6275
rect 38668 6267 38680 6275
rect 38696 6267 38744 6275
rect 38760 6267 38776 6275
rect 38792 6267 38796 6275
rect 38800 6267 38812 6275
rect 38824 6267 38828 6275
rect 38832 6267 38836 6275
rect 38856 6267 38860 6275
rect 38864 6267 38876 6275
rect 38880 6267 38892 6275
rect 38896 6267 38900 6275
rect 38920 6267 38924 6275
rect 38928 6267 38932 6275
rect 38980 6267 38984 6275
rect 38988 6267 38992 6275
rect 39012 6267 39016 6275
rect 39020 6267 39024 6275
rect 39120 6267 39124 6275
rect 39128 6267 39132 6275
rect 39144 6267 39156 6275
rect 39160 6267 39164 6275
rect 39180 6267 39200 6275
rect 39212 6267 39228 6275
rect 39236 6267 39260 6275
rect 39276 6267 39292 6275
rect 39308 6267 39320 6275
rect 39332 6267 39336 6275
rect 39340 6267 39352 6275
rect 39356 6267 39360 6275
rect 39372 6267 39384 6275
rect 39424 6267 39428 6275
rect 39432 6267 39444 6275
rect 39448 6267 39452 6275
rect 39464 6267 39476 6275
rect 39484 6267 39508 6275
rect 39524 6267 39536 6275
rect 39540 6267 39544 6275
rect 39556 6267 39568 6275
rect 39580 6267 39584 6275
rect 39588 6267 39600 6275
rect 39704 6267 39708 6275
rect 39712 6267 39724 6275
rect 39744 6267 39756 6275
rect 39760 6267 39764 6275
rect 39776 6267 39788 6275
rect 39804 6267 39820 6275
rect 39836 6267 39884 6275
rect 39900 6267 39904 6275
rect 39908 6267 39912 6275
rect 39924 6267 39936 6275
rect 39940 6267 39952 6275
rect 39964 6267 39968 6275
rect 39972 6267 39976 6275
rect 40016 6267 40040 6275
rect 40056 6267 40068 6275
rect 40088 6267 40100 6275
rect 40104 6267 40116 6275
rect 40120 6267 40132 6275
rect 40152 6267 40164 6275
rect 40168 6267 40172 6275
rect 40184 6267 40196 6275
rect 40216 6267 40228 6275
rect 40248 6267 40260 6275
rect 40272 6267 40276 6275
rect 40280 6267 40292 6275
rect 40528 6267 40540 6275
rect 40544 6267 40556 6275
rect 40560 6267 40572 6275
rect 40592 6267 40604 6275
rect 40620 6267 40632 6275
rect 40636 6267 40648 6275
rect 40652 6267 40664 6275
rect 18536 6256 18538 6260
rect 18542 6252 18544 6256
rect 18740 6250 18744 6258
rect 18830 6250 18838 6258
rect 18964 6256 18966 6260
rect 18970 6252 18972 6256
rect 19366 6250 19370 6258
rect 19456 6250 19464 6258
rect 19778 6250 19782 6258
rect 19868 6250 19876 6258
rect 20682 6256 20684 6260
rect 20688 6252 20690 6256
rect 20816 6250 20820 6258
rect 20906 6250 20914 6258
rect 21442 6252 21444 6260
rect 21870 6252 21872 6260
rect 22458 6250 22466 6258
rect 22608 6250 22614 6258
rect 22672 6250 22680 6258
rect 22822 6250 22828 6258
rect 23742 6250 23756 6258
rect 23892 6250 23898 6258
rect 23948 6250 23954 6258
rect 23956 6250 23962 6258
rect 24218 6250 24232 6258
rect 24418 6256 24422 6258
rect 24488 6250 24494 6258
rect 24496 6250 24502 6258
rect 24542 6250 24548 6258
rect 24550 6250 24556 6258
rect 24636 6250 24642 6258
rect 24738 6250 24740 6258
rect 24900 6250 24906 6258
rect 24908 6250 24914 6258
rect 24954 6250 24960 6258
rect 24962 6250 24968 6258
rect 25028 6256 25032 6258
rect 25098 6250 25104 6258
rect 25106 6250 25112 6258
rect 25152 6250 25158 6258
rect 25160 6250 25166 6258
rect 25872 6250 25878 6258
rect 25966 6250 25978 6258
rect 26188 6250 26190 6258
rect 26350 6250 26356 6258
rect 26358 6250 26364 6258
rect 26404 6250 26410 6258
rect 26412 6250 26418 6258
rect 26498 6250 26504 6258
rect 26592 6250 26604 6258
rect 26690 6250 26698 6258
rect 27028 6250 27030 6258
rect 27124 6250 27130 6258
rect 27338 6250 27344 6258
rect 27618 6250 27624 6258
rect 27626 6250 27632 6258
rect 27672 6250 27678 6258
rect 27680 6250 27686 6258
rect 27746 6256 27750 6258
rect 28058 6250 28070 6258
rect 28392 6250 28398 6258
rect 30528 6257 30536 6265
rect 34704 6257 34712 6265
rect 35168 6257 35176 6265
rect 35328 6257 35336 6265
rect 36048 6257 36056 6265
rect 38992 6257 39000 6265
rect 19136 6240 19144 6248
rect 20736 6240 20744 6248
rect 22224 6240 22232 6248
rect 29376 6237 29384 6245
rect 29792 6237 29800 6245
rect 30016 6237 30024 6245
rect 30480 6237 30488 6245
rect 30576 6237 30584 6245
rect 30768 6237 30776 6245
rect 31424 6237 31432 6245
rect 32128 6237 32136 6245
rect 32224 6237 32232 6245
rect 32496 6237 32504 6245
rect 33424 6237 33432 6245
rect 34112 6237 34120 6245
rect 40224 6237 40232 6245
rect 40464 6237 40472 6245
rect 19920 6220 19928 6228
rect 23024 6220 23032 6228
rect 23408 6220 23416 6228
rect 31184 6217 31192 6225
rect 32400 6217 32408 6225
rect 32624 6217 32632 6225
rect 32704 6217 32712 6225
rect 33664 6217 33672 6225
rect 33952 6217 33960 6225
rect 34064 6217 34072 6225
rect 39584 6217 39592 6225
rect 39696 6217 39704 6225
rect 39872 6217 39880 6225
rect 18640 6200 18648 6208
rect 18928 6200 18936 6208
rect 20768 6200 20776 6208
rect 22192 6200 22200 6208
rect 28416 6200 28424 6208
rect 29616 6197 29624 6205
rect 29824 6197 29832 6205
rect 30096 6197 30104 6205
rect 30304 6197 30312 6205
rect 30320 6197 30328 6205
rect 30608 6197 30616 6205
rect 30720 6197 30728 6205
rect 30752 6197 30760 6205
rect 31200 6197 31208 6205
rect 31952 6197 31960 6205
rect 32256 6197 32264 6205
rect 33264 6197 33272 6205
rect 33744 6197 33752 6205
rect 34432 6197 34440 6205
rect 34896 6197 34904 6205
rect 35424 6197 35432 6205
rect 35488 6197 35496 6205
rect 35840 6197 35848 6205
rect 36144 6197 36152 6205
rect 36512 6197 36520 6205
rect 37024 6197 37032 6205
rect 37440 6197 37448 6205
rect 37664 6197 37672 6205
rect 37872 6197 37880 6205
rect 37952 6197 37960 6205
rect 38192 6197 38200 6205
rect 38336 6197 38344 6205
rect 38352 6197 38360 6205
rect 38560 6197 38568 6205
rect 38784 6197 38792 6205
rect 39024 6197 39032 6205
rect 40016 6197 40024 6205
rect 40144 6197 40152 6205
rect 40464 6197 40472 6205
rect 40496 6197 40504 6205
rect 40560 6197 40568 6205
rect 19072 6180 19080 6188
rect 19280 6180 19288 6188
rect 19760 6180 19768 6188
rect 20112 6180 20120 6188
rect 21168 6180 21176 6188
rect 21328 6180 21336 6188
rect 21824 6180 21832 6188
rect 22208 6180 22216 6188
rect 22784 6180 22792 6188
rect 22880 6180 22888 6188
rect 23248 6180 23256 6188
rect 24288 6180 24296 6188
rect 24720 6180 24728 6188
rect 25344 6180 25352 6188
rect 25568 6180 25576 6188
rect 26240 6180 26248 6188
rect 26928 6180 26936 6188
rect 27184 6180 27192 6188
rect 28160 6180 28168 6188
rect 28480 6180 28488 6188
rect 31568 6177 31576 6185
rect 33424 6177 33432 6185
rect 38576 6177 38584 6185
rect 39616 6177 39624 6185
rect 29440 6157 29448 6165
rect 29840 6157 29848 6165
rect 30000 6157 30008 6165
rect 30304 6157 30312 6165
rect 31776 6157 31784 6165
rect 32192 6157 32200 6165
rect 32272 6157 32280 6165
rect 32880 6157 32888 6165
rect 33856 6157 33864 6165
rect 34672 6157 34680 6165
rect 35344 6157 35352 6165
rect 35856 6157 35864 6165
rect 36208 6157 36216 6165
rect 36768 6157 36776 6165
rect 37088 6157 37096 6165
rect 37328 6157 37336 6165
rect 37984 6157 37992 6165
rect 40080 6157 40088 6165
rect 40544 6157 40552 6165
rect 19088 6148 19092 6153
rect 19500 6148 19504 6153
rect 21346 6148 21350 6153
rect 26148 6148 26152 6153
rect 19296 6140 19304 6148
rect 19696 6140 19704 6148
rect 20192 6140 20200 6148
rect 20528 6140 20536 6148
rect 20576 6140 20584 6148
rect 22592 6140 22600 6148
rect 23520 6140 23528 6148
rect 24496 6140 24504 6148
rect 25744 6140 25752 6148
rect 26944 6140 26952 6148
rect 26992 6140 27000 6148
rect 31328 6137 31336 6145
rect 36480 6137 36488 6145
rect 36704 6137 36712 6145
rect 36784 6137 36792 6145
rect 20192 6120 20200 6128
rect 22176 6120 22184 6128
rect 27808 6120 27816 6128
rect 35584 6117 35592 6125
rect 35744 6117 35752 6125
rect 36880 6117 36888 6125
rect 38080 6117 38088 6125
rect 38096 6117 38104 6125
rect 21760 6100 21768 6108
rect 25120 6100 25128 6108
rect 31312 6097 31320 6105
rect 25904 6080 25912 6088
rect 27808 6080 27816 6088
rect 27824 6080 27832 6088
rect 36224 6077 36232 6085
rect 37856 6077 37864 6085
rect 18496 6060 18504 6068
rect 20736 6060 20744 6068
rect 27168 6060 27176 6068
rect 29396 6067 29408 6075
rect 29428 6067 29440 6075
rect 29444 6067 29448 6075
rect 29460 6067 29472 6075
rect 29488 6067 29504 6075
rect 29512 6067 29544 6075
rect 29552 6067 29568 6075
rect 29576 6067 29588 6075
rect 29592 6067 29596 6075
rect 29616 6067 29620 6075
rect 29624 6067 29636 6075
rect 29640 6067 29652 6075
rect 29656 6067 29660 6075
rect 29708 6067 29712 6075
rect 29716 6067 29728 6075
rect 29732 6067 29744 6075
rect 29748 6067 29752 6075
rect 29768 6067 29784 6075
rect 29800 6067 29804 6075
rect 29808 6067 29820 6075
rect 29824 6067 29836 6075
rect 29840 6067 29844 6075
rect 29860 6067 29876 6075
rect 29892 6067 29896 6075
rect 29900 6067 29912 6075
rect 29916 6067 29928 6075
rect 29932 6067 29936 6075
rect 29984 6067 29988 6075
rect 29992 6067 30004 6075
rect 30008 6067 30020 6075
rect 30024 6067 30028 6075
rect 30188 6067 30192 6075
rect 30196 6067 30200 6075
rect 30288 6067 30300 6075
rect 30312 6067 30316 6075
rect 30320 6067 30332 6075
rect 30336 6067 30340 6075
rect 30444 6067 30456 6075
rect 30476 6067 30488 6075
rect 30492 6067 30504 6075
rect 30508 6067 30520 6075
rect 30592 6067 30596 6075
rect 30600 6067 30612 6075
rect 30632 6067 30644 6075
rect 30648 6067 30652 6075
rect 30684 6067 30688 6075
rect 30692 6067 30704 6075
rect 30724 6067 30736 6075
rect 30740 6067 30744 6075
rect 30776 6067 30780 6075
rect 30784 6067 30796 6075
rect 30816 6067 30828 6075
rect 30832 6067 30844 6075
rect 30848 6067 30860 6075
rect 30876 6067 30892 6075
rect 30908 6067 30932 6075
rect 30940 6067 30956 6075
rect 30972 6067 30988 6075
rect 30996 6067 31020 6075
rect 31036 6067 31048 6075
rect 31068 6067 31080 6075
rect 31084 6067 31096 6075
rect 31100 6067 31112 6075
rect 31128 6067 31140 6075
rect 31160 6067 31172 6075
rect 31176 6067 31188 6075
rect 31192 6067 31200 6075
rect 31224 6067 31236 6075
rect 31244 6067 31276 6075
rect 31284 6067 31300 6075
rect 31316 6067 31328 6075
rect 31340 6067 31344 6075
rect 31348 6067 31360 6075
rect 31380 6067 31392 6075
rect 31404 6067 31408 6075
rect 31412 6067 31424 6075
rect 31428 6067 31432 6075
rect 31444 6067 31456 6075
rect 31472 6067 31484 6075
rect 31496 6067 31500 6075
rect 31504 6067 31516 6075
rect 31520 6067 31524 6075
rect 31536 6067 31548 6075
rect 31564 6067 31580 6075
rect 31596 6067 31620 6075
rect 31628 6067 31644 6075
rect 31652 6067 31664 6075
rect 31668 6067 31672 6075
rect 31692 6067 31696 6075
rect 31700 6067 31712 6075
rect 31716 6067 31728 6075
rect 31732 6067 31736 6075
rect 31752 6067 31756 6075
rect 31760 6067 31764 6075
rect 31784 6067 31788 6075
rect 31792 6067 31804 6075
rect 31808 6067 31820 6075
rect 31824 6067 31828 6075
rect 31848 6067 31852 6075
rect 31856 6067 31860 6075
rect 31908 6067 31912 6075
rect 31916 6067 31920 6075
rect 31940 6067 31944 6075
rect 31948 6067 31952 6075
rect 32000 6067 32004 6075
rect 32008 6067 32012 6075
rect 32124 6067 32128 6075
rect 32132 6067 32144 6075
rect 32148 6067 32160 6075
rect 32164 6067 32168 6075
rect 32188 6067 32192 6075
rect 32196 6067 32200 6075
rect 32216 6067 32232 6075
rect 32240 6067 32264 6075
rect 32280 6067 32304 6075
rect 32312 6067 32324 6075
rect 32336 6067 32340 6075
rect 32344 6067 32356 6075
rect 32376 6067 32388 6075
rect 32400 6067 32404 6075
rect 32408 6067 32420 6075
rect 32440 6067 32452 6075
rect 32456 6067 32460 6075
rect 32472 6067 32484 6075
rect 32500 6067 32516 6075
rect 32532 6067 32580 6075
rect 32596 6067 32612 6075
rect 32620 6067 32644 6075
rect 32660 6067 32676 6075
rect 32692 6067 32716 6075
rect 32724 6067 32740 6075
rect 32756 6067 32760 6075
rect 32764 6067 32768 6075
rect 32780 6067 32792 6075
rect 32804 6067 32808 6075
rect 32812 6067 32824 6075
rect 32840 6067 32872 6075
rect 32888 6067 32904 6075
rect 32912 6067 32924 6075
rect 32936 6067 32940 6075
rect 32944 6067 32948 6075
rect 33060 6067 33064 6075
rect 33068 6067 33072 6075
rect 33084 6067 33096 6075
rect 33104 6067 33120 6075
rect 33136 6067 33152 6075
rect 33160 6067 33184 6075
rect 33200 6067 33216 6075
rect 33232 6067 33244 6075
rect 33248 6067 33260 6075
rect 33264 6067 33276 6075
rect 33292 6067 33308 6075
rect 33324 6067 33336 6075
rect 33340 6067 33352 6075
rect 33356 6067 33368 6075
rect 33384 6067 33400 6075
rect 33416 6067 33440 6075
rect 33448 6067 33464 6075
rect 33480 6067 33484 6075
rect 33488 6067 33492 6075
rect 33504 6067 33516 6075
rect 33520 6067 33532 6075
rect 33544 6067 33548 6075
rect 33552 6067 33556 6075
rect 33604 6067 33608 6075
rect 33612 6067 33624 6075
rect 33636 6067 33640 6075
rect 33644 6067 33648 6075
rect 33660 6067 33672 6075
rect 33676 6067 33688 6075
rect 33700 6067 33704 6075
rect 33708 6067 33712 6075
rect 33724 6067 33736 6075
rect 33740 6067 33744 6075
rect 33792 6067 33796 6075
rect 33800 6067 33804 6075
rect 33816 6067 33828 6075
rect 33832 6067 33836 6075
rect 33856 6067 33860 6075
rect 33864 6067 33868 6075
rect 33884 6067 33900 6075
rect 33908 6067 33940 6075
rect 33948 6067 33964 6075
rect 33980 6067 33992 6075
rect 34000 6067 34032 6075
rect 34040 6067 34056 6075
rect 34072 6067 34076 6075
rect 34080 6067 34084 6075
rect 34104 6067 34108 6075
rect 34112 6067 34124 6075
rect 34136 6067 34140 6075
rect 34144 6067 34148 6075
rect 34160 6067 34172 6075
rect 34176 6067 34180 6075
rect 34200 6067 34204 6075
rect 34208 6067 34212 6075
rect 34224 6067 34236 6075
rect 34240 6067 34244 6075
rect 34260 6067 34284 6075
rect 34292 6067 34308 6075
rect 34316 6067 34328 6075
rect 34332 6067 34336 6075
rect 34352 6067 34376 6075
rect 34384 6067 34400 6075
rect 34408 6067 34420 6075
rect 34424 6067 34428 6075
rect 34448 6067 34452 6075
rect 34456 6067 34468 6075
rect 34476 6067 34492 6075
rect 34500 6067 34512 6075
rect 34516 6067 34520 6075
rect 34540 6067 34544 6075
rect 34548 6067 34560 6075
rect 34572 6067 34576 6075
rect 34580 6067 34584 6075
rect 34680 6067 34684 6075
rect 34688 6067 34692 6075
rect 34712 6067 34716 6075
rect 34720 6067 34732 6075
rect 34736 6067 34748 6075
rect 34752 6067 34756 6075
rect 34776 6067 34780 6075
rect 34784 6067 34788 6075
rect 34804 6067 34820 6075
rect 34828 6067 34852 6075
rect 34868 6067 34880 6075
rect 34884 6067 34888 6075
rect 34900 6067 34912 6075
rect 34924 6067 34928 6075
rect 34932 6067 34944 6075
rect 34960 6067 34972 6075
rect 34976 6067 34980 6075
rect 34992 6067 35004 6075
rect 35016 6067 35020 6075
rect 35024 6067 35036 6075
rect 35052 6067 35064 6075
rect 35068 6067 35072 6075
rect 35084 6067 35096 6075
rect 35108 6067 35112 6075
rect 35116 6067 35128 6075
rect 35132 6067 35136 6075
rect 35148 6067 35160 6075
rect 35200 6067 35204 6075
rect 35208 6067 35220 6075
rect 35224 6067 35228 6075
rect 35292 6067 35296 6075
rect 35300 6067 35312 6075
rect 35316 6067 35320 6075
rect 35384 6067 35388 6075
rect 35392 6067 35404 6075
rect 35408 6067 35412 6075
rect 35424 6067 35436 6075
rect 35452 6067 35468 6075
rect 35484 6067 35508 6075
rect 35516 6067 35532 6075
rect 35540 6067 35564 6075
rect 35580 6067 35596 6075
rect 35612 6067 35624 6075
rect 35636 6067 35640 6075
rect 35644 6067 35656 6075
rect 35660 6067 35664 6075
rect 35676 6067 35688 6075
rect 35792 6067 35796 6075
rect 35800 6067 35812 6075
rect 35816 6067 35820 6075
rect 35884 6067 35888 6075
rect 35892 6067 35904 6075
rect 35908 6067 35912 6075
rect 35952 6067 35964 6075
rect 35976 6067 35980 6075
rect 35984 6067 35996 6075
rect 36000 6067 36004 6075
rect 36200 6067 36212 6075
rect 36416 6067 36428 6075
rect 36432 6067 36436 6075
rect 36448 6067 36460 6075
rect 36476 6067 36492 6075
rect 36500 6067 36532 6075
rect 36540 6067 36552 6075
rect 36572 6067 36584 6075
rect 36588 6067 36600 6075
rect 36604 6067 36616 6075
rect 36632 6067 36648 6075
rect 36656 6067 36688 6075
rect 36696 6067 36712 6075
rect 36728 6067 36744 6075
rect 36760 6067 36764 6075
rect 36768 6067 36780 6075
rect 36792 6067 36796 6075
rect 36800 6067 36804 6075
rect 36816 6067 36828 6075
rect 36832 6067 36836 6075
rect 36932 6067 36936 6075
rect 36940 6067 36944 6075
rect 36956 6067 36968 6075
rect 36972 6067 36984 6075
rect 36992 6067 37008 6075
rect 37024 6067 37040 6075
rect 37048 6067 37060 6075
rect 37064 6067 37076 6075
rect 37088 6067 37092 6075
rect 37096 6067 37100 6075
rect 37116 6067 37132 6075
rect 37140 6067 37164 6075
rect 37180 6067 37196 6075
rect 37204 6067 37236 6075
rect 37244 6067 37256 6075
rect 37276 6067 37288 6075
rect 37292 6067 37304 6075
rect 37308 6067 37320 6075
rect 37340 6067 37352 6075
rect 37356 6067 37360 6075
rect 37392 6067 37396 6075
rect 37400 6067 37412 6075
rect 37432 6067 37444 6075
rect 37448 6067 37452 6075
rect 37464 6067 37476 6075
rect 37492 6067 37508 6075
rect 37524 6067 37572 6075
rect 37588 6067 37592 6075
rect 37596 6067 37600 6075
rect 37612 6067 37624 6075
rect 37628 6067 37640 6075
rect 37652 6067 37656 6075
rect 37660 6067 37664 6075
rect 37684 6067 37688 6075
rect 37692 6067 37696 6075
rect 37792 6067 37796 6075
rect 37800 6067 37804 6075
rect 37816 6067 37828 6075
rect 37832 6067 37836 6075
rect 37852 6067 37868 6075
rect 37884 6067 37900 6075
rect 37908 6067 37940 6075
rect 37948 6067 37964 6075
rect 37976 6067 37992 6075
rect 38000 6067 38032 6075
rect 38040 6067 38052 6075
rect 38072 6067 38084 6075
rect 38092 6067 38124 6075
rect 38132 6067 38148 6075
rect 38160 6067 38176 6075
rect 38184 6067 38216 6075
rect 38224 6067 38236 6075
rect 38256 6067 38268 6075
rect 38280 6067 38284 6075
rect 38288 6067 38300 6075
rect 38320 6067 38332 6075
rect 38352 6067 38364 6075
rect 38368 6067 38372 6075
rect 38384 6067 38396 6075
rect 38416 6067 38428 6075
rect 38432 6067 38444 6075
rect 38448 6067 38460 6075
rect 38480 6067 38492 6075
rect 38496 6067 38508 6075
rect 38512 6067 38524 6075
rect 38544 6067 38556 6075
rect 38576 6067 38588 6075
rect 38608 6067 38620 6075
rect 38640 6067 38652 6075
rect 38656 6067 38668 6075
rect 38672 6067 38684 6075
rect 38828 6067 38840 6075
rect 38844 6067 38848 6075
rect 38860 6067 38872 6075
rect 38884 6067 38888 6075
rect 38892 6067 38904 6075
rect 38908 6067 38912 6075
rect 38924 6067 38936 6075
rect 38948 6067 38952 6075
rect 38956 6067 38968 6075
rect 39176 6067 39188 6075
rect 39200 6067 39204 6075
rect 39208 6067 39220 6075
rect 39224 6067 39228 6075
rect 39240 6067 39252 6075
rect 39268 6067 39284 6075
rect 39300 6067 39324 6075
rect 39332 6067 39348 6075
rect 39356 6067 39380 6075
rect 39396 6067 39400 6075
rect 39404 6067 39416 6075
rect 39424 6067 39440 6075
rect 39448 6067 39472 6075
rect 39488 6067 39500 6075
rect 39520 6067 39532 6075
rect 39544 6067 39548 6075
rect 39552 6067 39564 6075
rect 39568 6067 39572 6075
rect 39584 6067 39596 6075
rect 39612 6067 39628 6075
rect 39644 6067 39668 6075
rect 39676 6067 39692 6075
rect 39700 6067 39712 6075
rect 39716 6067 39720 6075
rect 39740 6067 39744 6075
rect 39748 6067 39760 6075
rect 39772 6067 39776 6075
rect 39780 6067 39784 6075
rect 39804 6067 39808 6075
rect 39812 6067 39824 6075
rect 39836 6067 39840 6075
rect 39844 6067 39848 6075
rect 39860 6067 39872 6075
rect 39876 6067 39880 6075
rect 39976 6067 39980 6075
rect 39984 6067 39988 6075
rect 40052 6067 40056 6075
rect 40060 6067 40064 6075
rect 40084 6067 40088 6075
rect 40092 6067 40096 6075
rect 40108 6067 40120 6075
rect 40124 6067 40128 6075
rect 40148 6067 40152 6075
rect 40156 6067 40168 6075
rect 40180 6067 40184 6075
rect 40188 6067 40192 6075
rect 40212 6067 40216 6075
rect 40220 6067 40224 6075
rect 40244 6067 40248 6075
rect 40252 6067 40256 6075
rect 40268 6067 40280 6075
rect 40284 6067 40288 6075
rect 40304 6067 40328 6075
rect 40336 6067 40352 6075
rect 40360 6067 40372 6075
rect 40376 6067 40380 6075
rect 40396 6067 40420 6075
rect 40428 6067 40444 6075
rect 40452 6067 40476 6075
rect 40492 6067 40496 6075
rect 40500 6067 40512 6075
rect 40520 6067 40536 6075
rect 40544 6067 40556 6075
rect 40560 6067 40564 6075
rect 40584 6067 40588 6075
rect 40592 6067 40604 6075
rect 40612 6067 40628 6075
rect 40636 6067 40660 6075
rect 40676 6067 40692 6075
rect 40708 6067 40724 6075
rect 40740 6067 40764 6075
rect 40772 6067 40788 6075
rect 20242 6050 20252 6058
rect 21050 6050 21060 6058
rect 22928 6050 22938 6058
rect 23142 6050 23152 6058
rect 23356 6050 23366 6058
rect 23570 6050 23580 6058
rect 26660 6050 26662 6058
rect 26668 6050 26670 6058
rect 26874 6050 26876 6058
rect 26882 6050 26884 6058
rect 36016 6037 36024 6045
rect 39824 6037 39832 6045
rect 34832 6017 34840 6025
rect 35280 6017 35288 6025
rect 35296 6017 35304 6025
rect 40368 6017 40376 6025
rect 19456 6000 19464 6008
rect 19936 6000 19944 6008
rect 26400 6000 26408 6008
rect 32704 5997 32712 6005
rect 34752 5997 34760 6005
rect 37648 5997 37656 6005
rect 38128 5997 38136 6005
rect 40560 5997 40568 6005
rect 26784 5980 26792 5988
rect 30224 5977 30232 5985
rect 30608 5977 30616 5985
rect 30896 5977 30904 5985
rect 31664 5977 31672 5985
rect 31920 5977 31928 5985
rect 32064 5977 32072 5985
rect 33392 5977 33400 5985
rect 34608 5977 34616 5985
rect 35456 5977 35464 5985
rect 35648 5977 35656 5985
rect 35664 5977 35672 5985
rect 35936 5977 35944 5985
rect 36304 5977 36312 5985
rect 36736 5977 36744 5985
rect 37360 5977 37368 5985
rect 37408 5977 37416 5985
rect 37664 5977 37672 5985
rect 37872 5977 37880 5985
rect 39184 5977 39192 5985
rect 39344 5977 39352 5985
rect 18496 5960 18504 5968
rect 18849 5961 18850 5966
rect 19888 5960 19896 5968
rect 20752 5960 20760 5968
rect 21104 5960 21112 5968
rect 22368 5961 22378 5966
rect 22994 5961 23004 5966
rect 23200 5960 23208 5968
rect 24304 5960 24312 5968
rect 24528 5960 24536 5968
rect 24736 5960 24744 5968
rect 24912 5960 24920 5968
rect 25088 5960 25096 5968
rect 25504 5960 25512 5968
rect 26560 5960 26568 5968
rect 26816 5960 26824 5968
rect 27456 5960 27464 5968
rect 27809 5961 27812 5966
rect 28448 5960 28456 5968
rect 30048 5957 30056 5965
rect 30096 5957 30104 5965
rect 31344 5957 31352 5965
rect 31856 5957 31864 5965
rect 32176 5957 32184 5965
rect 32416 5957 32424 5965
rect 33152 5957 33160 5965
rect 33184 5957 33192 5965
rect 21936 5940 21944 5948
rect 22176 5940 22184 5948
rect 23696 5940 23704 5948
rect 27776 5940 27784 5948
rect 30640 5937 30648 5945
rect 31104 5937 31112 5945
rect 31328 5937 31336 5945
rect 31600 5937 31608 5945
rect 32048 5937 32056 5945
rect 32960 5937 32968 5945
rect 32992 5937 33000 5945
rect 33056 5937 33064 5945
rect 34896 5937 34904 5945
rect 35552 5937 35560 5945
rect 36224 5937 36232 5945
rect 37424 5937 37432 5945
rect 37616 5937 37624 5945
rect 37920 5937 37928 5945
rect 39328 5937 39336 5945
rect 39888 5937 39896 5945
rect 40064 5937 40072 5945
rect 40224 5937 40232 5945
rect 40240 5937 40248 5945
rect 40432 5937 40440 5945
rect 18512 5920 18520 5928
rect 19680 5920 19688 5928
rect 19872 5920 19880 5928
rect 21072 5920 21080 5928
rect 21312 5920 21320 5928
rect 22976 5920 22984 5928
rect 23616 5920 23624 5928
rect 23904 5920 23912 5928
rect 24224 5920 24232 5928
rect 24304 5920 24312 5928
rect 24528 5920 24536 5928
rect 25488 5920 25496 5928
rect 25904 5920 25912 5928
rect 25936 5920 25944 5928
rect 26096 5920 26104 5928
rect 26320 5920 26328 5928
rect 26608 5920 26616 5928
rect 26832 5920 26840 5928
rect 27248 5920 27256 5928
rect 27632 5920 27640 5928
rect 28016 5920 28024 5928
rect 28448 5920 28456 5928
rect 29728 5917 29736 5925
rect 30256 5917 30264 5925
rect 31712 5917 31720 5925
rect 32624 5917 32632 5925
rect 32816 5917 32824 5925
rect 36704 5917 36712 5925
rect 37120 5917 37128 5925
rect 37984 5917 37992 5925
rect 38192 5917 38200 5925
rect 38864 5917 38872 5925
rect 40176 5917 40184 5925
rect 40368 5917 40376 5925
rect 40672 5917 40680 5925
rect 19520 5900 19528 5908
rect 20928 5900 20936 5908
rect 21168 5900 21176 5908
rect 21536 5900 21544 5908
rect 23184 5900 23192 5908
rect 25088 5900 25096 5908
rect 26576 5900 26584 5908
rect 29456 5897 29464 5905
rect 30400 5897 30408 5905
rect 30992 5897 31000 5905
rect 31520 5897 31528 5905
rect 34000 5897 34008 5905
rect 34224 5897 34232 5905
rect 34464 5897 34472 5905
rect 34640 5897 34648 5905
rect 34656 5897 34664 5905
rect 34800 5897 34808 5905
rect 35008 5897 35016 5905
rect 35312 5897 35320 5905
rect 35536 5897 35544 5905
rect 36064 5897 36072 5905
rect 38704 5897 38712 5905
rect 19088 5880 19096 5888
rect 19296 5880 19304 5888
rect 20928 5880 20936 5888
rect 21968 5880 21976 5888
rect 23472 5880 23480 5888
rect 23872 5880 23880 5888
rect 25552 5880 25560 5888
rect 27024 5880 27032 5888
rect 27632 5880 27640 5888
rect 37552 5877 37560 5885
rect 37664 5877 37672 5885
rect 40304 5877 40312 5885
rect 19712 5860 19720 5868
rect 24080 5860 24088 5868
rect 28288 5860 28296 5868
rect 29428 5867 29440 5875
rect 29444 5867 29448 5875
rect 29460 5867 29472 5875
rect 29488 5867 29504 5875
rect 29512 5867 29544 5875
rect 29552 5867 29568 5875
rect 29576 5867 29600 5875
rect 29616 5867 29620 5875
rect 29624 5867 29636 5875
rect 29640 5867 29652 5875
rect 29656 5867 29660 5875
rect 29680 5867 29684 5875
rect 29688 5867 29692 5875
rect 29708 5867 29724 5875
rect 29732 5867 29756 5875
rect 29772 5867 29784 5875
rect 29788 5867 29792 5875
rect 29804 5867 29816 5875
rect 29828 5867 29832 5875
rect 29836 5867 29848 5875
rect 29852 5867 29856 5875
rect 29984 5867 29988 5875
rect 29992 5867 30004 5875
rect 30008 5867 30012 5875
rect 30024 5867 30036 5875
rect 30212 5867 30224 5875
rect 30236 5867 30240 5875
rect 30244 5867 30256 5875
rect 30260 5867 30264 5875
rect 30344 5867 30348 5875
rect 30352 5867 30356 5875
rect 30376 5867 30380 5875
rect 30384 5867 30388 5875
rect 30436 5867 30440 5875
rect 30444 5867 30448 5875
rect 30468 5867 30472 5875
rect 30476 5867 30480 5875
rect 30492 5867 30504 5875
rect 30508 5867 30512 5875
rect 30532 5867 30536 5875
rect 30540 5867 30544 5875
rect 30556 5867 30568 5875
rect 30572 5867 30584 5875
rect 30592 5867 30608 5875
rect 30624 5867 30640 5875
rect 30648 5867 30660 5875
rect 30664 5867 30676 5875
rect 30684 5867 30700 5875
rect 30716 5867 30732 5875
rect 30740 5867 30764 5875
rect 30780 5867 30792 5875
rect 30812 5867 30824 5875
rect 30828 5867 30840 5875
rect 30844 5867 30856 5875
rect 30928 5867 30932 5875
rect 30936 5867 30948 5875
rect 30968 5867 30980 5875
rect 30984 5867 30988 5875
rect 31000 5867 31012 5875
rect 31032 5867 31044 5875
rect 31048 5867 31052 5875
rect 31064 5867 31076 5875
rect 31084 5867 31108 5875
rect 31124 5867 31136 5875
rect 31140 5867 31144 5875
rect 31156 5867 31168 5875
rect 31176 5867 31200 5875
rect 31216 5867 31240 5875
rect 31248 5867 31260 5875
rect 31272 5867 31276 5875
rect 31280 5867 31292 5875
rect 31312 5867 31324 5875
rect 31344 5867 31356 5875
rect 31376 5867 31388 5875
rect 31392 5867 31396 5875
rect 31408 5867 31420 5875
rect 31432 5867 31436 5875
rect 31440 5867 31452 5875
rect 31556 5867 31560 5875
rect 31564 5867 31576 5875
rect 31596 5867 31608 5875
rect 31612 5867 31624 5875
rect 31628 5867 31640 5875
rect 31656 5867 31672 5875
rect 31688 5867 31712 5875
rect 31720 5867 31736 5875
rect 31752 5867 31756 5875
rect 31760 5867 31764 5875
rect 31776 5867 31788 5875
rect 31792 5867 31804 5875
rect 31812 5867 31828 5875
rect 31844 5867 31860 5875
rect 31868 5867 31880 5875
rect 31884 5867 31896 5875
rect 31908 5867 31912 5875
rect 31916 5867 31920 5875
rect 31936 5867 31952 5875
rect 31960 5867 31972 5875
rect 31976 5867 31988 5875
rect 32000 5867 32004 5875
rect 32008 5867 32012 5875
rect 32028 5867 32032 5875
rect 32036 5867 32040 5875
rect 32052 5867 32064 5875
rect 32068 5867 32080 5875
rect 32092 5867 32096 5875
rect 32100 5867 32104 5875
rect 32120 5867 32168 5875
rect 32184 5867 32200 5875
rect 32216 5867 32228 5875
rect 32240 5867 32244 5875
rect 32248 5867 32260 5875
rect 32280 5867 32292 5875
rect 32296 5867 32300 5875
rect 32404 5867 32416 5875
rect 32420 5867 32424 5875
rect 32436 5867 32448 5875
rect 32460 5867 32464 5875
rect 32468 5867 32480 5875
rect 32496 5867 32508 5875
rect 32512 5867 32516 5875
rect 32532 5867 32556 5875
rect 32564 5867 32580 5875
rect 32588 5867 32604 5875
rect 32620 5867 32636 5875
rect 32652 5867 32656 5875
rect 32660 5867 32672 5875
rect 32744 5867 32748 5875
rect 32752 5867 32756 5875
rect 32868 5867 32872 5875
rect 32876 5867 32880 5875
rect 32892 5867 32904 5875
rect 32916 5867 32920 5875
rect 32924 5867 32928 5875
rect 32944 5867 32960 5875
rect 32968 5867 32992 5875
rect 33008 5867 33020 5875
rect 33040 5867 33052 5875
rect 33056 5867 33068 5875
rect 33080 5867 33084 5875
rect 33088 5867 33092 5875
rect 33104 5867 33116 5875
rect 33292 5867 33304 5875
rect 33316 5867 33320 5875
rect 33324 5867 33336 5875
rect 33340 5867 33344 5875
rect 33356 5867 33368 5875
rect 33376 5867 33400 5875
rect 33416 5867 33440 5875
rect 33448 5867 33464 5875
rect 33480 5867 33484 5875
rect 33488 5867 33492 5875
rect 33512 5867 33516 5875
rect 33520 5867 33532 5875
rect 33536 5867 33548 5875
rect 33552 5867 33556 5875
rect 33668 5867 33672 5875
rect 33676 5867 33688 5875
rect 33692 5867 33704 5875
rect 33708 5867 33712 5875
rect 33732 5867 33736 5875
rect 33740 5867 33744 5875
rect 33760 5867 33764 5875
rect 33768 5867 33780 5875
rect 33784 5867 33796 5875
rect 33800 5867 33804 5875
rect 33824 5867 33828 5875
rect 33832 5867 33836 5875
rect 33852 5867 33868 5875
rect 33876 5867 33900 5875
rect 33916 5867 33964 5875
rect 33980 5867 33996 5875
rect 34012 5867 34016 5875
rect 34020 5867 34032 5875
rect 34044 5867 34048 5875
rect 34052 5867 34056 5875
rect 34168 5867 34172 5875
rect 34176 5867 34180 5875
rect 34192 5867 34204 5875
rect 34208 5867 34212 5875
rect 34232 5867 34236 5875
rect 34240 5867 34244 5875
rect 34256 5867 34268 5875
rect 34272 5867 34284 5875
rect 34296 5867 34300 5875
rect 34304 5867 34308 5875
rect 34404 5867 34408 5875
rect 34412 5867 34424 5875
rect 34436 5867 34440 5875
rect 34444 5867 34448 5875
rect 34460 5867 34472 5875
rect 34476 5867 34488 5875
rect 34496 5867 34512 5875
rect 34528 5867 34544 5875
rect 34552 5867 34576 5875
rect 34592 5867 34604 5875
rect 34624 5867 34636 5875
rect 34640 5867 34652 5875
rect 34656 5867 34668 5875
rect 34684 5867 34696 5875
rect 34716 5867 34728 5875
rect 34732 5867 34744 5875
rect 34748 5867 34760 5875
rect 34780 5867 34792 5875
rect 34796 5867 34800 5875
rect 34872 5867 34884 5875
rect 34904 5867 34916 5875
rect 34920 5867 34924 5875
rect 34936 5867 34948 5875
rect 34956 5867 34980 5875
rect 34996 5867 35020 5875
rect 35028 5867 35040 5875
rect 35048 5867 35072 5875
rect 35088 5867 35136 5875
rect 35152 5867 35168 5875
rect 35184 5867 35188 5875
rect 35192 5867 35200 5875
rect 35216 5867 35220 5875
rect 35224 5867 35228 5875
rect 35324 5867 35328 5875
rect 35332 5867 35336 5875
rect 35432 5867 35436 5875
rect 35440 5867 35444 5875
rect 35456 5867 35468 5875
rect 35472 5867 35476 5875
rect 35496 5867 35500 5875
rect 35504 5867 35508 5875
rect 35524 5867 35572 5875
rect 35588 5867 35604 5875
rect 35620 5867 35624 5875
rect 35628 5867 35640 5875
rect 35652 5867 35656 5875
rect 35660 5867 35664 5875
rect 35684 5867 35688 5875
rect 35692 5867 35696 5875
rect 35824 5867 35828 5875
rect 35832 5867 35836 5875
rect 35856 5867 35860 5875
rect 35864 5867 35876 5875
rect 35880 5867 35892 5875
rect 35896 5867 35900 5875
rect 35916 5867 35932 5875
rect 35948 5867 35964 5875
rect 35972 5867 35996 5875
rect 36012 5867 36024 5875
rect 36028 5867 36032 5875
rect 36044 5867 36056 5875
rect 36068 5867 36072 5875
rect 36076 5867 36088 5875
rect 36092 5867 36096 5875
rect 36136 5867 36148 5875
rect 36160 5867 36164 5875
rect 36168 5867 36180 5875
rect 36184 5867 36188 5875
rect 36200 5867 36212 5875
rect 36228 5867 36240 5875
rect 36252 5867 36256 5875
rect 36260 5867 36272 5875
rect 36276 5867 36280 5875
rect 36320 5867 36332 5875
rect 36344 5867 36348 5875
rect 36352 5867 36364 5875
rect 36368 5867 36372 5875
rect 36384 5867 36396 5875
rect 36412 5867 36428 5875
rect 36444 5867 36468 5875
rect 36476 5867 36492 5875
rect 36500 5867 36524 5875
rect 36536 5867 36560 5875
rect 36568 5867 36584 5875
rect 36592 5867 36616 5875
rect 36632 5867 36636 5875
rect 36640 5867 36652 5875
rect 36656 5867 36668 5875
rect 36672 5867 36676 5875
rect 36804 5867 36808 5875
rect 36812 5867 36824 5875
rect 36828 5867 36840 5875
rect 36844 5867 36848 5875
rect 36868 5867 36872 5875
rect 36876 5867 36880 5875
rect 36896 5867 36912 5875
rect 36920 5867 36944 5875
rect 36960 5867 36984 5875
rect 36992 5867 37004 5875
rect 37016 5867 37020 5875
rect 37024 5867 37036 5875
rect 37052 5867 37076 5875
rect 37084 5867 37096 5875
rect 37108 5867 37112 5875
rect 37116 5867 37128 5875
rect 37148 5867 37160 5875
rect 37180 5867 37192 5875
rect 37212 5867 37224 5875
rect 37228 5867 37232 5875
rect 37244 5867 37256 5875
rect 37268 5867 37272 5875
rect 37276 5867 37288 5875
rect 37292 5867 37296 5875
rect 37308 5867 37320 5875
rect 37492 5867 37504 5875
rect 37524 5867 37536 5875
rect 37540 5867 37544 5875
rect 37556 5867 37568 5875
rect 37584 5867 37600 5875
rect 37608 5867 37640 5875
rect 37648 5867 37664 5875
rect 37680 5867 37692 5875
rect 37700 5867 37732 5875
rect 37740 5867 37756 5875
rect 37772 5867 37788 5875
rect 37804 5867 37808 5875
rect 37812 5867 37824 5875
rect 37836 5867 37840 5875
rect 37844 5867 37848 5875
rect 37976 5867 37980 5875
rect 37984 5867 37988 5875
rect 38000 5867 38012 5875
rect 38016 5867 38020 5875
rect 38036 5867 38052 5875
rect 38068 5867 38116 5875
rect 38132 5867 38136 5875
rect 38140 5867 38144 5875
rect 38160 5867 38208 5875
rect 38224 5867 38236 5875
rect 38252 5867 38300 5875
rect 38316 5867 38340 5875
rect 38348 5867 38364 5875
rect 38380 5867 38400 5875
rect 38412 5867 38428 5875
rect 38436 5867 38468 5875
rect 38476 5867 38492 5875
rect 38500 5867 38524 5875
rect 38540 5867 38544 5875
rect 38548 5867 38560 5875
rect 38572 5867 38576 5875
rect 38580 5867 38584 5875
rect 38696 5867 38700 5875
rect 38704 5867 38708 5875
rect 38804 5867 38808 5875
rect 38812 5867 38816 5875
rect 38864 5867 38868 5875
rect 38872 5867 38876 5875
rect 38896 5867 38900 5875
rect 38904 5867 38916 5875
rect 38920 5867 38932 5875
rect 38936 5867 38940 5875
rect 38960 5867 38964 5875
rect 38968 5867 38972 5875
rect 38988 5867 39004 5875
rect 39012 5867 39036 5875
rect 39052 5867 39076 5875
rect 39084 5867 39100 5875
rect 39116 5867 39140 5875
rect 39148 5867 39164 5875
rect 39172 5867 39184 5875
rect 39188 5867 39192 5875
rect 39212 5867 39216 5875
rect 39220 5867 39232 5875
rect 39236 5867 39248 5875
rect 39252 5867 39256 5875
rect 39272 5867 39276 5875
rect 39280 5867 39284 5875
rect 39304 5867 39308 5875
rect 39312 5867 39324 5875
rect 39328 5867 39340 5875
rect 39344 5867 39348 5875
rect 39368 5867 39372 5875
rect 39376 5867 39380 5875
rect 39396 5867 39400 5875
rect 39404 5867 39416 5875
rect 39420 5867 39432 5875
rect 39436 5867 39440 5875
rect 39460 5867 39464 5875
rect 39468 5867 39472 5875
rect 39492 5867 39496 5875
rect 39500 5867 39504 5875
rect 39524 5867 39528 5875
rect 39532 5867 39536 5875
rect 39556 5867 39560 5875
rect 39564 5867 39576 5875
rect 39580 5867 39592 5875
rect 39596 5867 39600 5875
rect 39648 5867 39652 5875
rect 39656 5867 39668 5875
rect 39672 5867 39684 5875
rect 39688 5867 39692 5875
rect 39708 5867 39712 5875
rect 39716 5867 39720 5875
rect 39740 5867 39744 5875
rect 39748 5867 39760 5875
rect 39764 5867 39776 5875
rect 39780 5867 39784 5875
rect 39804 5867 39808 5875
rect 39812 5867 39824 5875
rect 39832 5867 39848 5875
rect 39856 5867 39880 5875
rect 39896 5867 39900 5875
rect 39904 5867 39916 5875
rect 39924 5867 39940 5875
rect 39948 5867 39972 5875
rect 39988 5867 39992 5875
rect 39996 5867 40008 5875
rect 40016 5867 40032 5875
rect 40040 5867 40064 5875
rect 40080 5867 40096 5875
rect 40112 5867 40128 5875
rect 40144 5867 40168 5875
rect 40176 5867 40192 5875
rect 40200 5867 40224 5875
rect 40240 5867 40252 5875
rect 40272 5867 40284 5875
rect 40296 5867 40300 5875
rect 40304 5867 40316 5875
rect 40320 5867 40324 5875
rect 40336 5867 40348 5875
rect 40364 5867 40376 5875
rect 40388 5867 40392 5875
rect 40396 5867 40408 5875
rect 40412 5867 40416 5875
rect 40428 5867 40440 5875
rect 40460 5867 40472 5875
rect 40488 5867 40512 5875
rect 40520 5867 40536 5875
rect 40544 5867 40556 5875
rect 40560 5867 40564 5875
rect 40584 5867 40588 5875
rect 40592 5867 40604 5875
rect 40612 5867 40628 5875
rect 40636 5867 40660 5875
rect 40676 5867 40692 5875
rect 40708 5867 40720 5875
rect 40732 5867 40736 5875
rect 40740 5867 40752 5875
rect 40756 5867 40760 5875
rect 40772 5867 40784 5875
rect 18526 5850 18530 5858
rect 18616 5850 18624 5858
rect 19564 5852 19566 5860
rect 19762 5850 19766 5858
rect 19852 5850 19860 5858
rect 20046 5852 20048 5860
rect 20174 5850 20178 5858
rect 20264 5850 20272 5858
rect 20458 5852 20460 5860
rect 20656 5852 20658 5860
rect 20998 5852 21000 5860
rect 22860 5850 22864 5858
rect 22950 5850 22958 5858
rect 23074 5850 23078 5858
rect 23164 5850 23172 5858
rect 23304 5852 23306 5860
rect 24112 5850 24116 5858
rect 24202 5850 24210 5858
rect 24502 5850 24510 5858
rect 24652 5850 24658 5858
rect 24716 5850 24724 5858
rect 24866 5850 24872 5858
rect 25144 5850 25158 5858
rect 25578 5850 25582 5858
rect 25668 5850 25676 5858
rect 26364 5850 26372 5858
rect 26514 5850 26520 5858
rect 26578 5850 26586 5858
rect 26728 5850 26734 5858
rect 26792 5850 26800 5858
rect 26942 5850 26948 5858
rect 27220 5850 27228 5858
rect 27370 5850 27376 5858
rect 27434 5850 27442 5858
rect 27584 5850 27590 5858
rect 31936 5857 31944 5865
rect 21936 5840 21944 5848
rect 28432 5840 28440 5848
rect 29440 5837 29448 5845
rect 29728 5837 29736 5845
rect 30720 5837 30728 5845
rect 30896 5837 30904 5845
rect 31760 5837 31768 5845
rect 33488 5837 33496 5845
rect 34192 5837 34200 5845
rect 38016 5837 38024 5845
rect 38112 5837 38120 5845
rect 38288 5837 38296 5845
rect 38384 5837 38392 5845
rect 39056 5837 39064 5845
rect 39232 5837 39240 5845
rect 20928 5820 20936 5828
rect 22592 5820 22600 5828
rect 24432 5820 24440 5828
rect 27152 5820 27160 5828
rect 27408 5820 27416 5828
rect 29968 5817 29976 5825
rect 30064 5817 30072 5825
rect 30224 5817 30232 5825
rect 31040 5817 31048 5825
rect 31376 5817 31384 5825
rect 33200 5817 33208 5825
rect 33424 5817 33432 5825
rect 33456 5817 33464 5825
rect 33872 5817 33880 5825
rect 36096 5817 36104 5825
rect 36672 5817 36680 5825
rect 40224 5817 40232 5825
rect 40256 5817 40264 5825
rect 21136 5800 21144 5808
rect 23216 5800 23224 5808
rect 24080 5800 24088 5808
rect 26768 5800 26776 5808
rect 27008 5800 27016 5808
rect 27200 5800 27208 5808
rect 30000 5797 30008 5805
rect 30464 5797 30472 5805
rect 30496 5797 30504 5805
rect 30736 5797 30744 5805
rect 32256 5797 32264 5805
rect 32432 5797 32440 5805
rect 32720 5797 32728 5805
rect 32800 5797 32808 5805
rect 33072 5797 33080 5805
rect 33616 5797 33624 5805
rect 35472 5797 35480 5805
rect 35936 5797 35944 5805
rect 36096 5797 36104 5805
rect 36368 5797 36376 5805
rect 36576 5797 36584 5805
rect 36752 5797 36760 5805
rect 37024 5797 37032 5805
rect 37280 5797 37288 5805
rect 37568 5797 37576 5805
rect 38896 5797 38904 5805
rect 39088 5797 39096 5805
rect 39472 5797 39480 5805
rect 39520 5797 39528 5805
rect 39760 5797 39768 5805
rect 39872 5797 39880 5805
rect 40096 5797 40104 5805
rect 40752 5797 40760 5805
rect 18736 5780 18744 5788
rect 19440 5780 19448 5788
rect 19936 5780 19944 5788
rect 21296 5780 21304 5788
rect 21568 5780 21576 5788
rect 21776 5780 21784 5788
rect 22192 5780 22200 5788
rect 22416 5780 22424 5788
rect 22464 5780 22472 5788
rect 22736 5780 22744 5788
rect 23424 5780 23432 5788
rect 25360 5780 25368 5788
rect 25952 5780 25960 5788
rect 26144 5780 26152 5788
rect 26560 5780 26568 5788
rect 26688 5780 26696 5788
rect 27344 5780 27352 5788
rect 28480 5780 28488 5788
rect 31696 5777 31704 5785
rect 33456 5777 33464 5785
rect 35488 5777 35496 5785
rect 20016 5760 20024 5768
rect 21984 5760 21992 5768
rect 25760 5760 25768 5768
rect 30016 5757 30024 5765
rect 30352 5757 30360 5765
rect 30944 5757 30952 5765
rect 31200 5757 31208 5765
rect 31904 5757 31912 5765
rect 32448 5757 32456 5765
rect 32576 5757 32584 5765
rect 32832 5757 32840 5765
rect 32896 5757 32904 5765
rect 33024 5757 33032 5765
rect 33632 5757 33640 5765
rect 34704 5757 34712 5765
rect 35072 5757 35080 5765
rect 35312 5757 35320 5765
rect 36864 5757 36872 5765
rect 36960 5757 36968 5765
rect 37040 5757 37048 5765
rect 37424 5757 37432 5765
rect 37712 5757 37720 5765
rect 38496 5757 38504 5765
rect 38768 5757 38776 5765
rect 38880 5757 38888 5765
rect 39296 5757 39304 5765
rect 39888 5757 39896 5765
rect 19468 5748 19472 5753
rect 20530 5748 20534 5753
rect 21766 5748 21770 5753
rect 26699 5748 26710 5753
rect 19728 5740 19736 5748
rect 19920 5740 19928 5748
rect 21088 5740 21096 5748
rect 21296 5740 21304 5748
rect 23456 5740 23464 5748
rect 23808 5740 23816 5748
rect 24848 5740 24856 5748
rect 25744 5740 25752 5748
rect 27632 5740 27640 5748
rect 28064 5740 28072 5748
rect 31680 5737 31688 5745
rect 32240 5737 32248 5745
rect 32544 5737 32552 5745
rect 33872 5737 33880 5745
rect 36912 5737 36920 5745
rect 18496 5720 18504 5728
rect 28224 5720 28232 5728
rect 38336 5717 38344 5725
rect 21968 5700 21976 5708
rect 27648 5700 27656 5708
rect 27856 5700 27864 5708
rect 32000 5697 32008 5705
rect 38464 5697 38472 5705
rect 36656 5677 36664 5685
rect 37408 5677 37416 5685
rect 38848 5677 38856 5685
rect 20912 5660 20920 5668
rect 23616 5660 23624 5668
rect 23648 5660 23656 5668
rect 29420 5667 29424 5675
rect 29428 5667 29440 5675
rect 29444 5667 29448 5675
rect 29460 5667 29472 5675
rect 29480 5667 29504 5675
rect 29520 5667 29532 5675
rect 29536 5667 29540 5675
rect 29552 5667 29564 5675
rect 29576 5667 29580 5675
rect 29584 5667 29596 5675
rect 29612 5667 29636 5675
rect 29644 5667 29656 5675
rect 29668 5667 29672 5675
rect 29676 5667 29688 5675
rect 29792 5667 29796 5675
rect 29800 5667 29812 5675
rect 29832 5667 29844 5675
rect 29848 5667 29860 5675
rect 29864 5667 29876 5675
rect 29896 5667 29908 5675
rect 29916 5667 29948 5675
rect 29956 5667 29972 5675
rect 29980 5667 30004 5675
rect 30020 5667 30024 5675
rect 30028 5667 30040 5675
rect 30048 5667 30064 5675
rect 30072 5667 30096 5675
rect 30112 5667 30116 5675
rect 30120 5667 30132 5675
rect 30144 5667 30148 5675
rect 30152 5667 30156 5675
rect 30176 5667 30180 5675
rect 30184 5667 30196 5675
rect 30208 5667 30212 5675
rect 30216 5667 30220 5675
rect 30232 5667 30244 5675
rect 30248 5667 30252 5675
rect 30268 5667 30272 5675
rect 30276 5667 30288 5675
rect 30300 5667 30304 5675
rect 30308 5667 30312 5675
rect 30324 5667 30336 5675
rect 30340 5667 30344 5675
rect 30364 5667 30368 5675
rect 30372 5667 30376 5675
rect 30416 5667 30448 5675
rect 30456 5667 30472 5675
rect 30488 5667 30512 5675
rect 30520 5667 30536 5675
rect 30552 5667 30556 5675
rect 30560 5667 30564 5675
rect 30576 5667 30588 5675
rect 30592 5667 30604 5675
rect 30616 5667 30620 5675
rect 30624 5667 30628 5675
rect 30644 5667 30660 5675
rect 30668 5667 30692 5675
rect 30708 5667 30724 5675
rect 30740 5667 30764 5675
rect 30772 5667 30788 5675
rect 30804 5667 30820 5675
rect 30828 5667 30840 5675
rect 30844 5667 30856 5675
rect 30868 5667 30872 5675
rect 30876 5667 30880 5675
rect 30892 5667 30904 5675
rect 30908 5667 30912 5675
rect 30928 5667 30932 5675
rect 30936 5667 30948 5675
rect 30960 5667 30964 5675
rect 30968 5667 30972 5675
rect 31084 5667 31088 5675
rect 31092 5667 31104 5675
rect 31116 5667 31120 5675
rect 31124 5667 31128 5675
rect 31176 5667 31180 5675
rect 31184 5667 31196 5675
rect 31208 5667 31212 5675
rect 31216 5667 31220 5675
rect 31232 5667 31244 5675
rect 31248 5667 31260 5675
rect 31272 5667 31276 5675
rect 31280 5667 31284 5675
rect 31304 5667 31308 5675
rect 31312 5667 31316 5675
rect 31380 5667 31384 5675
rect 31388 5667 31400 5675
rect 31412 5667 31416 5675
rect 31420 5667 31424 5675
rect 31436 5667 31448 5675
rect 31452 5667 31456 5675
rect 31472 5667 31488 5675
rect 31504 5667 31520 5675
rect 31528 5667 31560 5675
rect 31568 5667 31584 5675
rect 31600 5667 31612 5675
rect 31616 5667 31628 5675
rect 31632 5667 31644 5675
rect 31664 5667 31676 5675
rect 31688 5667 31692 5675
rect 31696 5667 31708 5675
rect 31728 5667 31740 5675
rect 31812 5667 31816 5675
rect 31820 5667 31824 5675
rect 31912 5667 31924 5675
rect 31928 5667 31932 5675
rect 32028 5667 32032 5675
rect 32036 5667 32040 5675
rect 32052 5667 32064 5675
rect 32068 5667 32080 5675
rect 32100 5667 32112 5675
rect 32120 5667 32136 5675
rect 32144 5667 32168 5675
rect 32184 5667 32188 5675
rect 32192 5667 32204 5675
rect 32220 5667 32268 5675
rect 32284 5667 32300 5675
rect 32312 5667 32360 5675
rect 32376 5667 32392 5675
rect 32404 5667 32452 5675
rect 32468 5667 32484 5675
rect 32492 5667 32504 5675
rect 32508 5667 32520 5675
rect 32648 5667 32660 5675
rect 32664 5667 32676 5675
rect 32692 5667 32708 5675
rect 32724 5667 32748 5675
rect 32764 5667 32776 5675
rect 32800 5667 32808 5675
rect 32812 5667 32824 5675
rect 32840 5667 32856 5675
rect 32872 5667 32884 5675
rect 32888 5667 32900 5675
rect 32920 5667 32932 5675
rect 32936 5667 32940 5675
rect 32988 5667 32992 5675
rect 32996 5667 33000 5675
rect 33040 5667 33052 5675
rect 33064 5667 33068 5675
rect 33072 5667 33084 5675
rect 33088 5667 33092 5675
rect 33104 5667 33116 5675
rect 33316 5667 33320 5675
rect 33324 5667 33336 5675
rect 33340 5667 33344 5675
rect 33356 5667 33368 5675
rect 33380 5667 33384 5675
rect 33388 5667 33400 5675
rect 33420 5667 33432 5675
rect 33452 5667 33464 5675
rect 33484 5667 33496 5675
rect 33500 5667 33504 5675
rect 33516 5667 33528 5675
rect 33540 5667 33544 5675
rect 33548 5667 33560 5675
rect 33580 5667 33592 5675
rect 33604 5667 33608 5675
rect 33612 5667 33624 5675
rect 33644 5667 33656 5675
rect 33660 5667 33664 5675
rect 33696 5667 33700 5675
rect 33704 5667 33716 5675
rect 33736 5667 33748 5675
rect 33752 5667 33756 5675
rect 33788 5667 33792 5675
rect 33796 5667 33808 5675
rect 33828 5667 33840 5675
rect 33844 5667 33848 5675
rect 33960 5667 33964 5675
rect 33968 5667 33972 5675
rect 33984 5667 33996 5675
rect 34000 5667 34004 5675
rect 34020 5667 34036 5675
rect 34052 5667 34068 5675
rect 34076 5667 34108 5675
rect 34116 5667 34132 5675
rect 34148 5667 34160 5675
rect 34168 5667 34200 5675
rect 34208 5667 34224 5675
rect 34240 5667 34252 5675
rect 34256 5667 34268 5675
rect 34272 5667 34284 5675
rect 34304 5667 34316 5675
rect 34336 5667 34348 5675
rect 34368 5667 34380 5675
rect 34400 5667 34412 5675
rect 34416 5667 34428 5675
rect 34432 5667 34444 5675
rect 34464 5667 34476 5675
rect 34480 5667 34484 5675
rect 34676 5667 34680 5675
rect 34684 5667 34688 5675
rect 34708 5667 34712 5675
rect 34716 5667 34728 5675
rect 34732 5667 34736 5675
rect 34748 5667 34760 5675
rect 34780 5667 34792 5675
rect 34796 5667 34800 5675
rect 34812 5667 34824 5675
rect 34844 5667 34856 5675
rect 34868 5667 34872 5675
rect 34876 5667 34888 5675
rect 34908 5667 34920 5675
rect 35000 5667 35012 5675
rect 35116 5667 35120 5675
rect 35124 5667 35136 5675
rect 35140 5667 35144 5675
rect 35156 5667 35168 5675
rect 35188 5667 35200 5675
rect 35216 5667 35240 5675
rect 35248 5667 35264 5675
rect 35272 5667 35296 5675
rect 35312 5667 35316 5675
rect 35320 5667 35332 5675
rect 35340 5667 35356 5675
rect 35364 5667 35396 5675
rect 35404 5667 35420 5675
rect 35436 5667 35448 5675
rect 35456 5667 35488 5675
rect 35496 5667 35512 5675
rect 35528 5667 35540 5675
rect 35552 5667 35556 5675
rect 35560 5667 35572 5675
rect 35592 5667 35604 5675
rect 35624 5667 35636 5675
rect 35640 5667 35644 5675
rect 35656 5667 35668 5675
rect 35684 5667 35700 5675
rect 35708 5667 35740 5675
rect 35748 5667 35764 5675
rect 35780 5667 35796 5675
rect 35812 5667 35828 5675
rect 35844 5667 35860 5675
rect 35868 5667 35900 5675
rect 35908 5667 35924 5675
rect 35940 5667 35964 5675
rect 35972 5667 35988 5675
rect 36004 5667 36008 5675
rect 36012 5667 36016 5675
rect 36028 5667 36040 5675
rect 36044 5667 36056 5675
rect 36068 5667 36072 5675
rect 36076 5667 36080 5675
rect 36128 5667 36132 5675
rect 36136 5667 36148 5675
rect 36160 5667 36164 5675
rect 36168 5667 36172 5675
rect 36220 5667 36224 5675
rect 36228 5667 36240 5675
rect 36252 5667 36256 5675
rect 36260 5667 36264 5675
rect 36276 5667 36288 5675
rect 36292 5667 36296 5675
rect 36312 5667 36328 5675
rect 36344 5667 36360 5675
rect 36368 5667 36400 5675
rect 36408 5667 36420 5675
rect 36440 5667 36452 5675
rect 36456 5667 36468 5675
rect 36472 5667 36484 5675
rect 36504 5667 36516 5675
rect 36620 5667 36624 5675
rect 36628 5667 36640 5675
rect 36644 5667 36648 5675
rect 36660 5667 36672 5675
rect 36680 5667 36704 5675
rect 36720 5667 36744 5675
rect 36752 5667 36764 5675
rect 36776 5667 36780 5675
rect 36784 5667 36796 5675
rect 36812 5667 36836 5675
rect 36844 5667 36856 5675
rect 36868 5667 36872 5675
rect 36876 5667 36888 5675
rect 36904 5667 36928 5675
rect 36936 5667 36952 5675
rect 36968 5667 36984 5675
rect 37000 5667 37004 5675
rect 37008 5667 37020 5675
rect 37024 5667 37036 5675
rect 37040 5667 37044 5675
rect 37064 5667 37068 5675
rect 37072 5667 37076 5675
rect 37332 5667 37336 5675
rect 37340 5667 37352 5675
rect 37356 5667 37368 5675
rect 37372 5667 37376 5675
rect 37392 5667 37408 5675
rect 37424 5667 37428 5675
rect 37432 5667 37444 5675
rect 37448 5667 37460 5675
rect 37464 5667 37468 5675
rect 37488 5667 37492 5675
rect 37496 5667 37500 5675
rect 37520 5667 37524 5675
rect 37528 5667 37532 5675
rect 37552 5667 37556 5675
rect 37560 5667 37564 5675
rect 37584 5667 37588 5675
rect 37592 5667 37604 5675
rect 37608 5667 37620 5675
rect 37624 5667 37628 5675
rect 37648 5667 37652 5675
rect 37656 5667 37668 5675
rect 37676 5667 37692 5675
rect 37700 5667 37724 5675
rect 37740 5667 37756 5675
rect 37772 5667 37788 5675
rect 37804 5667 37828 5675
rect 37836 5667 37852 5675
rect 37860 5667 37884 5675
rect 37900 5667 37904 5675
rect 37908 5667 37920 5675
rect 37924 5667 37936 5675
rect 37940 5667 37944 5675
rect 38040 5667 38044 5675
rect 38048 5667 38052 5675
rect 38072 5667 38076 5675
rect 38080 5667 38092 5675
rect 38096 5667 38108 5675
rect 38112 5667 38116 5675
rect 38164 5667 38168 5675
rect 38172 5667 38184 5675
rect 38188 5667 38200 5675
rect 38204 5667 38208 5675
rect 38228 5667 38232 5675
rect 38236 5667 38240 5675
rect 38256 5667 38260 5675
rect 38264 5667 38276 5675
rect 38280 5667 38292 5675
rect 38296 5667 38300 5675
rect 38320 5667 38324 5675
rect 38328 5667 38340 5675
rect 38348 5667 38364 5675
rect 38372 5667 38400 5675
rect 38412 5667 38428 5675
rect 38444 5667 38456 5675
rect 38460 5667 38472 5675
rect 38476 5667 38488 5675
rect 38508 5667 38520 5675
rect 38528 5667 38560 5675
rect 38568 5667 38584 5675
rect 38596 5667 38612 5675
rect 38620 5667 38652 5675
rect 38660 5667 38676 5675
rect 38684 5667 38708 5675
rect 38724 5667 38728 5675
rect 38732 5667 38744 5675
rect 38748 5667 38760 5675
rect 38764 5667 38768 5675
rect 38788 5667 38792 5675
rect 38796 5667 38800 5675
rect 38816 5667 38820 5675
rect 38824 5667 38836 5675
rect 38840 5667 38852 5675
rect 38856 5667 38860 5675
rect 38988 5667 38992 5675
rect 38996 5667 39000 5675
rect 39012 5667 39024 5675
rect 39028 5667 39032 5675
rect 39052 5667 39056 5675
rect 39060 5667 39072 5675
rect 39084 5667 39088 5675
rect 39092 5667 39096 5675
rect 39272 5667 39276 5675
rect 39280 5667 39292 5675
rect 39304 5667 39308 5675
rect 39312 5667 39316 5675
rect 39396 5667 39400 5675
rect 39404 5667 39408 5675
rect 39648 5667 39652 5675
rect 39656 5667 39660 5675
rect 39672 5667 39684 5675
rect 39688 5667 39692 5675
rect 39708 5667 39712 5675
rect 39716 5667 39728 5675
rect 39740 5667 39744 5675
rect 39748 5667 39752 5675
rect 39764 5667 39776 5675
rect 39780 5667 39784 5675
rect 39832 5667 39836 5675
rect 39840 5667 39844 5675
rect 39856 5667 39868 5675
rect 39872 5667 39876 5675
rect 39924 5667 39928 5675
rect 39932 5667 39936 5675
rect 39948 5667 39960 5675
rect 39964 5667 39968 5675
rect 40016 5667 40020 5675
rect 40024 5667 40028 5675
rect 40188 5667 40192 5675
rect 40196 5667 40208 5675
rect 40220 5667 40224 5675
rect 40228 5667 40232 5675
rect 40280 5667 40284 5675
rect 40288 5667 40300 5675
rect 40312 5667 40316 5675
rect 40320 5667 40324 5675
rect 40336 5667 40348 5675
rect 40352 5667 40356 5675
rect 40404 5667 40408 5675
rect 40412 5667 40416 5675
rect 40428 5667 40440 5675
rect 40444 5667 40448 5675
rect 40468 5667 40472 5675
rect 40476 5667 40480 5675
rect 40492 5667 40504 5675
rect 40508 5667 40512 5675
rect 40528 5667 40552 5675
rect 40560 5667 40576 5675
rect 40584 5667 40608 5675
rect 40624 5667 40628 5675
rect 40632 5667 40644 5675
rect 40656 5667 40660 5675
rect 40664 5667 40668 5675
rect 40688 5667 40692 5675
rect 40696 5667 40700 5675
rect 40780 5667 40784 5675
rect 40788 5667 40792 5675
rect 26112 5658 26116 5660
rect 21110 5650 21122 5658
rect 21546 5650 21550 5658
rect 21554 5650 21558 5658
rect 21622 5650 21626 5658
rect 21630 5650 21634 5658
rect 21752 5650 21764 5658
rect 21828 5650 21840 5658
rect 21942 5650 21948 5658
rect 21950 5650 21956 5658
rect 22476 5650 22482 5658
rect 22484 5650 22490 5658
rect 22690 5650 22696 5658
rect 22698 5650 22704 5658
rect 22798 5650 22804 5658
rect 22806 5650 22812 5658
rect 23432 5650 23446 5658
rect 24058 5650 24072 5658
rect 24256 5650 24270 5658
rect 24576 5650 24590 5658
rect 24790 5650 24800 5658
rect 26112 5650 26126 5658
rect 26188 5650 26202 5658
rect 26646 5650 26660 5658
rect 26722 5650 26736 5658
rect 27288 5650 27302 5658
rect 27364 5650 27378 5658
rect 27502 5650 27516 5658
rect 27578 5650 27592 5658
rect 27610 5650 27624 5658
rect 27686 5650 27700 5658
rect 28038 5650 28052 5658
rect 28114 5650 28128 5658
rect 28458 5650 28464 5658
rect 28466 5650 28472 5658
rect 28534 5650 28540 5658
rect 28542 5650 28548 5658
rect 26112 5648 26116 5650
rect 38528 5637 38536 5645
rect 32816 5617 32824 5625
rect 34560 5617 34568 5625
rect 36192 5617 36200 5625
rect 38304 5617 38312 5625
rect 39168 5617 39176 5625
rect 20736 5600 20744 5608
rect 25056 5600 25064 5608
rect 35328 5597 35336 5605
rect 35424 5597 35432 5605
rect 21888 5580 21896 5588
rect 29584 5577 29592 5585
rect 29888 5577 29896 5585
rect 30800 5577 30808 5585
rect 30880 5577 30888 5585
rect 31088 5577 31096 5585
rect 31152 5577 31160 5585
rect 31488 5577 31496 5585
rect 31728 5577 31736 5585
rect 31792 5577 31800 5585
rect 31872 5577 31880 5585
rect 32368 5577 32376 5585
rect 33488 5577 33496 5585
rect 34480 5577 34488 5585
rect 34896 5577 34904 5585
rect 35264 5577 35272 5585
rect 35728 5577 35736 5585
rect 37376 5577 37384 5585
rect 38064 5577 38072 5585
rect 38784 5577 38792 5585
rect 39552 5577 39560 5585
rect 39760 5577 39768 5585
rect 39936 5577 39944 5585
rect 40048 5577 40056 5585
rect 40368 5577 40376 5585
rect 40432 5577 40440 5585
rect 18720 5560 18728 5568
rect 18928 5560 18936 5568
rect 19136 5560 19144 5568
rect 19296 5560 19304 5568
rect 19472 5560 19480 5568
rect 19680 5560 19688 5568
rect 19888 5560 19896 5568
rect 21392 5560 21400 5568
rect 22464 5561 22474 5566
rect 22672 5560 22680 5568
rect 23104 5560 23112 5568
rect 24000 5560 24008 5568
rect 24784 5560 24792 5568
rect 24848 5560 24856 5568
rect 26128 5560 26136 5568
rect 26704 5560 26712 5568
rect 27344 5560 27352 5568
rect 27568 5561 27578 5566
rect 28416 5560 28424 5568
rect 30320 5557 30328 5565
rect 30368 5557 30376 5565
rect 33392 5557 33400 5565
rect 33424 5557 33432 5565
rect 36912 5557 36920 5565
rect 37104 5557 37112 5565
rect 38640 5557 38648 5565
rect 24528 5540 24536 5548
rect 24864 5540 24872 5548
rect 29584 5537 29592 5545
rect 30512 5537 30520 5545
rect 30576 5537 30584 5545
rect 30768 5537 30776 5545
rect 31552 5537 31560 5545
rect 31776 5537 31784 5545
rect 32352 5537 32360 5545
rect 32944 5537 32952 5545
rect 33728 5537 33736 5545
rect 33824 5537 33832 5545
rect 34192 5537 34200 5545
rect 35808 5537 35816 5545
rect 36032 5537 36040 5545
rect 36768 5537 36776 5545
rect 37120 5537 37128 5545
rect 37360 5537 37368 5545
rect 38544 5537 38552 5545
rect 38768 5537 38776 5545
rect 39296 5537 39304 5545
rect 39328 5537 39336 5545
rect 39360 5537 39368 5545
rect 40512 5537 40520 5545
rect 18736 5520 18744 5528
rect 19456 5520 19464 5528
rect 19872 5520 19880 5528
rect 20400 5520 20408 5528
rect 21376 5520 21384 5528
rect 21584 5520 21592 5528
rect 22656 5520 22664 5528
rect 22752 5520 22760 5528
rect 23408 5520 23416 5528
rect 25280 5520 25288 5528
rect 27328 5520 27336 5528
rect 27552 5520 27560 5528
rect 27648 5520 27656 5528
rect 27968 5520 27976 5528
rect 28496 5520 28504 5528
rect 30176 5517 30184 5525
rect 30368 5517 30376 5525
rect 30432 5517 30440 5525
rect 31184 5517 31192 5525
rect 33152 5517 33160 5525
rect 36320 5517 36328 5525
rect 36384 5517 36392 5525
rect 23184 5500 23192 5508
rect 23616 5500 23624 5508
rect 23808 5500 23816 5508
rect 26688 5500 26696 5508
rect 27184 5500 27192 5508
rect 31952 5497 31960 5505
rect 32016 5497 32024 5505
rect 33152 5497 33160 5505
rect 33744 5497 33752 5505
rect 33840 5497 33848 5505
rect 34000 5497 34008 5505
rect 34976 5497 34984 5505
rect 35472 5497 35480 5505
rect 35520 5497 35528 5505
rect 35536 5497 35544 5505
rect 35664 5497 35672 5505
rect 36560 5497 36568 5505
rect 37760 5497 37768 5505
rect 37936 5497 37944 5505
rect 38480 5497 38488 5505
rect 38736 5497 38744 5505
rect 39024 5497 39032 5505
rect 39392 5497 39400 5505
rect 40144 5497 40152 5505
rect 40272 5497 40280 5505
rect 40704 5497 40712 5505
rect 19920 5480 19928 5488
rect 24592 5480 24600 5488
rect 25008 5480 25016 5488
rect 28640 5480 28648 5488
rect 29680 5477 29688 5485
rect 32928 5477 32936 5485
rect 23344 5460 23352 5468
rect 23552 5460 23560 5468
rect 23760 5460 23768 5468
rect 25424 5460 25432 5468
rect 26096 5460 26104 5468
rect 26512 5460 26520 5468
rect 29524 5467 29536 5475
rect 29556 5467 29568 5475
rect 29572 5467 29584 5475
rect 29588 5467 29600 5475
rect 29620 5467 29632 5475
rect 29648 5467 29672 5475
rect 29680 5467 29696 5475
rect 29712 5467 29716 5475
rect 29720 5467 29724 5475
rect 29736 5467 29748 5475
rect 29752 5467 29764 5475
rect 29772 5467 29788 5475
rect 29804 5467 29808 5475
rect 29812 5467 29816 5475
rect 29828 5467 29840 5475
rect 29844 5467 29856 5475
rect 29864 5467 29880 5475
rect 29896 5467 29912 5475
rect 29920 5467 29932 5475
rect 29936 5467 29948 5475
rect 29956 5467 29972 5475
rect 29988 5467 30004 5475
rect 30012 5467 30024 5475
rect 30028 5467 30040 5475
rect 30052 5467 30056 5475
rect 30060 5467 30064 5475
rect 30084 5467 30088 5475
rect 30092 5467 30096 5475
rect 30256 5467 30260 5475
rect 30264 5467 30268 5475
rect 30280 5467 30292 5475
rect 30296 5467 30300 5475
rect 30320 5467 30324 5475
rect 30328 5467 30340 5475
rect 30352 5467 30356 5475
rect 30360 5467 30364 5475
rect 30460 5467 30464 5475
rect 30468 5467 30472 5475
rect 30492 5467 30496 5475
rect 30500 5467 30512 5475
rect 30516 5467 30528 5475
rect 30532 5467 30536 5475
rect 30552 5467 30556 5475
rect 30560 5467 30564 5475
rect 30584 5467 30588 5475
rect 30592 5467 30604 5475
rect 30608 5467 30620 5475
rect 30624 5467 30628 5475
rect 30648 5467 30652 5475
rect 30656 5467 30660 5475
rect 30672 5467 30684 5475
rect 30688 5467 30692 5475
rect 30708 5467 30724 5475
rect 30740 5467 30788 5475
rect 30804 5467 30816 5475
rect 30832 5467 30880 5475
rect 30896 5467 30908 5475
rect 30924 5467 30972 5475
rect 30988 5467 30992 5475
rect 30996 5467 31000 5475
rect 31012 5467 31024 5475
rect 31028 5467 31040 5475
rect 31052 5467 31056 5475
rect 31060 5467 31064 5475
rect 31080 5467 31128 5475
rect 31144 5467 31148 5475
rect 31152 5467 31156 5475
rect 31176 5467 31180 5475
rect 31184 5467 31196 5475
rect 31208 5467 31212 5475
rect 31216 5467 31220 5475
rect 31240 5467 31244 5475
rect 31248 5467 31260 5475
rect 31264 5467 31276 5475
rect 31280 5467 31284 5475
rect 31304 5467 31308 5475
rect 31312 5467 31316 5475
rect 31380 5467 31384 5475
rect 31388 5467 31392 5475
rect 31412 5467 31416 5475
rect 31420 5467 31424 5475
rect 31436 5467 31448 5475
rect 31452 5467 31456 5475
rect 31472 5467 31496 5475
rect 31504 5467 31520 5475
rect 31528 5467 31560 5475
rect 31568 5467 31584 5475
rect 31600 5467 31612 5475
rect 31624 5467 31628 5475
rect 31632 5467 31644 5475
rect 31664 5467 31676 5475
rect 31688 5467 31692 5475
rect 31696 5467 31708 5475
rect 31712 5467 31716 5475
rect 31728 5467 31740 5475
rect 31756 5467 31768 5475
rect 31780 5467 31784 5475
rect 31788 5467 31792 5475
rect 31804 5467 31816 5475
rect 31820 5467 31824 5475
rect 31912 5467 31924 5475
rect 31928 5467 31932 5475
rect 31952 5467 31956 5475
rect 31960 5467 31972 5475
rect 31984 5467 31988 5475
rect 31992 5467 31996 5475
rect 32016 5467 32020 5475
rect 32024 5467 32036 5475
rect 32124 5467 32128 5475
rect 32132 5467 32136 5475
rect 32156 5467 32160 5475
rect 32164 5467 32168 5475
rect 32312 5467 32316 5475
rect 32320 5467 32332 5475
rect 32336 5467 32340 5475
rect 32404 5467 32408 5475
rect 32412 5467 32424 5475
rect 32428 5467 32432 5475
rect 32444 5467 32456 5475
rect 32476 5467 32488 5475
rect 32492 5467 32496 5475
rect 32508 5467 32520 5475
rect 32540 5467 32552 5475
rect 32556 5467 32568 5475
rect 32572 5467 32584 5475
rect 32696 5467 32708 5475
rect 32728 5467 32740 5475
rect 32744 5467 32748 5475
rect 32764 5467 32780 5475
rect 32800 5467 32828 5475
rect 32840 5467 32856 5475
rect 32872 5467 32904 5475
rect 32912 5467 32928 5475
rect 32936 5467 32952 5475
rect 32960 5467 32976 5475
rect 32992 5467 33004 5475
rect 33016 5467 33020 5475
rect 33024 5467 33028 5475
rect 33132 5467 33144 5475
rect 33164 5467 33176 5475
rect 33180 5467 33184 5475
rect 33196 5467 33208 5475
rect 33224 5467 33240 5475
rect 33248 5467 33280 5475
rect 33288 5467 33304 5475
rect 33316 5467 33332 5475
rect 33340 5467 33372 5475
rect 33380 5467 33396 5475
rect 33412 5467 33416 5475
rect 33420 5467 33424 5475
rect 33444 5467 33448 5475
rect 33452 5467 33464 5475
rect 33476 5467 33480 5475
rect 33484 5467 33488 5475
rect 33584 5467 33588 5475
rect 33592 5467 33596 5475
rect 33616 5467 33620 5475
rect 33624 5467 33628 5475
rect 33640 5467 33652 5475
rect 33656 5467 33668 5475
rect 33680 5467 33684 5475
rect 33688 5467 33692 5475
rect 33788 5467 33792 5475
rect 33796 5467 33800 5475
rect 33968 5467 33980 5475
rect 33984 5467 33988 5475
rect 34020 5467 34024 5475
rect 34028 5467 34040 5475
rect 34060 5467 34072 5475
rect 34076 5467 34080 5475
rect 34152 5467 34164 5475
rect 34168 5467 34172 5475
rect 34184 5467 34196 5475
rect 34216 5467 34228 5475
rect 34244 5467 34292 5475
rect 34308 5467 34324 5475
rect 34340 5467 34352 5475
rect 34364 5467 34368 5475
rect 34372 5467 34384 5475
rect 34404 5467 34416 5475
rect 34420 5467 34424 5475
rect 34436 5467 34448 5475
rect 34468 5467 34480 5475
rect 34496 5467 34544 5475
rect 34560 5467 34592 5475
rect 34608 5467 34620 5475
rect 34640 5467 34652 5475
rect 34664 5467 34668 5475
rect 34672 5467 34676 5475
rect 34788 5467 34792 5475
rect 34796 5467 34800 5475
rect 34812 5467 34824 5475
rect 34840 5467 34856 5475
rect 34864 5467 34896 5475
rect 34912 5467 34924 5475
rect 34940 5467 34980 5475
rect 34992 5467 35008 5475
rect 35024 5467 35072 5475
rect 35088 5467 35092 5475
rect 35096 5467 35100 5475
rect 35116 5467 35164 5475
rect 35180 5467 35196 5475
rect 35212 5467 35224 5475
rect 35236 5467 35240 5475
rect 35244 5467 35256 5475
rect 35276 5467 35288 5475
rect 35292 5467 35296 5475
rect 35464 5467 35476 5475
rect 35480 5467 35484 5475
rect 35496 5467 35508 5475
rect 35520 5467 35524 5475
rect 35528 5467 35540 5475
rect 35560 5467 35572 5475
rect 35584 5467 35588 5475
rect 35592 5467 35604 5475
rect 35676 5467 35680 5475
rect 35684 5467 35696 5475
rect 35808 5467 35820 5475
rect 35840 5467 35852 5475
rect 35856 5467 35860 5475
rect 35872 5467 35884 5475
rect 35892 5467 35916 5475
rect 35932 5467 35980 5475
rect 36000 5467 36008 5475
rect 36024 5467 36072 5475
rect 36088 5467 36100 5475
rect 36120 5467 36132 5475
rect 36144 5467 36148 5475
rect 36152 5467 36164 5475
rect 36340 5467 36352 5475
rect 36356 5467 36360 5475
rect 36372 5467 36384 5475
rect 36392 5467 36416 5475
rect 36432 5467 36480 5475
rect 36496 5467 36520 5475
rect 36528 5467 36544 5475
rect 36560 5467 36564 5475
rect 36568 5467 36572 5475
rect 36592 5467 36596 5475
rect 36600 5467 36612 5475
rect 36616 5467 36628 5475
rect 36632 5467 36636 5475
rect 36748 5467 36752 5475
rect 36756 5467 36760 5475
rect 36824 5467 36828 5475
rect 36832 5467 36836 5475
rect 36916 5467 36920 5475
rect 36924 5467 36928 5475
rect 36948 5467 36952 5475
rect 36956 5467 36960 5475
rect 36972 5467 36984 5475
rect 36988 5467 36992 5475
rect 37008 5467 37032 5475
rect 37040 5467 37056 5475
rect 37064 5467 37088 5475
rect 37104 5467 37120 5475
rect 37136 5467 37148 5475
rect 37160 5467 37164 5475
rect 37168 5467 37180 5475
rect 37184 5467 37188 5475
rect 37292 5467 37304 5475
rect 37324 5467 37336 5475
rect 37340 5467 37352 5475
rect 37356 5467 37368 5475
rect 37384 5467 37400 5475
rect 37416 5467 37428 5475
rect 37432 5467 37444 5475
rect 37448 5467 37460 5475
rect 37480 5467 37492 5475
rect 37496 5467 37500 5475
rect 37512 5467 37524 5475
rect 37540 5467 37556 5475
rect 37572 5467 37620 5475
rect 37636 5467 37640 5475
rect 37644 5467 37648 5475
rect 37660 5467 37672 5475
rect 37676 5467 37688 5475
rect 37700 5467 37704 5475
rect 37708 5467 37712 5475
rect 37732 5467 37736 5475
rect 37740 5467 37744 5475
rect 37808 5467 37812 5475
rect 37816 5467 37828 5475
rect 37840 5467 37844 5475
rect 37848 5467 37852 5475
rect 37864 5467 37876 5475
rect 37880 5467 37884 5475
rect 37932 5467 37936 5475
rect 37940 5467 37944 5475
rect 37992 5467 37996 5475
rect 38000 5467 38012 5475
rect 38024 5467 38028 5475
rect 38032 5467 38036 5475
rect 38164 5467 38168 5475
rect 38172 5467 38176 5475
rect 38188 5467 38200 5475
rect 38204 5467 38216 5475
rect 38228 5467 38232 5475
rect 38236 5467 38240 5475
rect 38256 5467 38272 5475
rect 38280 5467 38304 5475
rect 38320 5467 38336 5475
rect 38352 5467 38364 5475
rect 38368 5467 38380 5475
rect 38384 5467 38396 5475
rect 38416 5467 38428 5475
rect 38444 5467 38456 5475
rect 38460 5467 38472 5475
rect 38476 5467 38488 5475
rect 38508 5467 38520 5475
rect 38532 5467 38536 5475
rect 38540 5467 38552 5475
rect 38572 5467 38584 5475
rect 38664 5467 38676 5475
rect 38688 5467 38692 5475
rect 38696 5467 38708 5475
rect 38712 5467 38716 5475
rect 38728 5467 38740 5475
rect 38752 5467 38756 5475
rect 38760 5467 38772 5475
rect 38788 5467 38812 5475
rect 38820 5467 38832 5475
rect 38844 5467 38848 5475
rect 38852 5467 38864 5475
rect 38884 5467 38896 5475
rect 38908 5467 38912 5475
rect 38916 5467 38928 5475
rect 38948 5467 38960 5475
rect 38964 5467 38968 5475
rect 38980 5467 38992 5475
rect 39008 5467 39024 5475
rect 39040 5467 39088 5475
rect 39100 5467 39116 5475
rect 39132 5467 39180 5475
rect 39200 5467 39212 5475
rect 39220 5467 39244 5475
rect 39260 5467 39276 5475
rect 39284 5467 39316 5475
rect 39324 5467 39336 5475
rect 39356 5467 39368 5475
rect 39376 5467 39408 5475
rect 39416 5467 39428 5475
rect 39448 5467 39460 5475
rect 39464 5467 39476 5475
rect 39480 5467 39492 5475
rect 39512 5467 39524 5475
rect 39540 5467 39564 5475
rect 39572 5467 39588 5475
rect 39604 5467 39652 5475
rect 39668 5467 39672 5475
rect 39676 5467 39680 5475
rect 39696 5467 39744 5475
rect 39760 5467 39776 5475
rect 39792 5467 39804 5475
rect 39816 5467 39820 5475
rect 39824 5467 39836 5475
rect 39856 5467 39868 5475
rect 39872 5467 39876 5475
rect 39908 5467 39912 5475
rect 39916 5467 39928 5475
rect 39948 5467 39960 5475
rect 39964 5467 39968 5475
rect 40040 5467 40052 5475
rect 40072 5467 40084 5475
rect 40088 5467 40092 5475
rect 40104 5467 40116 5475
rect 40128 5467 40132 5475
rect 40136 5467 40148 5475
rect 40152 5467 40156 5475
rect 40168 5467 40180 5475
rect 40196 5467 40208 5475
rect 40220 5467 40224 5475
rect 40228 5467 40240 5475
rect 40244 5467 40248 5475
rect 40260 5467 40272 5475
rect 40288 5467 40300 5475
rect 40312 5467 40316 5475
rect 40320 5467 40332 5475
rect 40336 5467 40340 5475
rect 40352 5467 40364 5475
rect 40384 5467 40396 5475
rect 40412 5467 40436 5475
rect 40444 5467 40460 5475
rect 40468 5467 40500 5475
rect 40508 5467 40524 5475
rect 40540 5467 40544 5475
rect 40548 5467 40552 5475
rect 40572 5467 40576 5475
rect 40580 5467 40592 5475
rect 40604 5467 40608 5475
rect 40612 5467 40616 5475
rect 40628 5467 40640 5475
rect 40644 5467 40648 5475
rect 40664 5467 40680 5475
rect 40696 5467 40712 5475
rect 40720 5467 40752 5475
rect 40760 5467 40772 5475
rect 40788 5467 40800 5475
rect 19992 5452 19994 5460
rect 20152 5450 20160 5458
rect 20302 5450 20308 5458
rect 20366 5450 20374 5458
rect 20516 5450 20522 5458
rect 20762 5450 20770 5458
rect 20914 5450 20920 5458
rect 20922 5450 20928 5458
rect 20976 5450 20984 5458
rect 21128 5450 21134 5458
rect 21136 5450 21150 5458
rect 21190 5450 21204 5458
rect 21272 5456 21276 5458
rect 21342 5450 21348 5458
rect 21350 5450 21356 5458
rect 21396 5450 21402 5458
rect 21404 5450 21410 5458
rect 21572 5450 21574 5458
rect 21786 5450 21788 5458
rect 22012 5450 22014 5458
rect 22210 5450 22214 5458
rect 22218 5450 22222 5458
rect 22420 5450 22422 5458
rect 23148 5450 23162 5458
rect 23362 5450 23376 5458
rect 23576 5450 23590 5458
rect 23790 5450 23804 5458
rect 24186 5450 24194 5458
rect 24524 5450 24536 5458
rect 24952 5452 24954 5460
rect 25470 5450 25484 5458
rect 25684 5450 25698 5458
rect 25898 5450 25912 5458
rect 26112 5450 26126 5458
rect 26578 5450 26582 5458
rect 26722 5450 26730 5458
rect 27006 5450 27010 5458
rect 27150 5450 27158 5458
rect 27396 5448 27400 5460
rect 27610 5448 27614 5460
rect 27824 5448 27828 5460
rect 28038 5448 28042 5460
rect 28252 5448 28256 5460
rect 28466 5448 28470 5460
rect 30976 5457 30984 5465
rect 31152 5457 31160 5465
rect 31328 5457 31336 5465
rect 31840 5457 31848 5465
rect 35232 5457 35240 5465
rect 35392 5457 35400 5465
rect 37664 5457 37672 5465
rect 38352 5457 38360 5465
rect 38464 5457 38472 5465
rect 23184 5440 23192 5448
rect 29936 5437 29944 5445
rect 30240 5437 30248 5445
rect 30432 5437 30440 5445
rect 30768 5437 30776 5445
rect 30848 5437 30856 5445
rect 31008 5437 31016 5445
rect 31536 5437 31544 5445
rect 31664 5437 31672 5445
rect 32096 5437 32104 5445
rect 32176 5437 32184 5445
rect 32272 5437 32280 5445
rect 32656 5437 32664 5445
rect 33072 5437 33080 5445
rect 33280 5437 33288 5445
rect 33312 5437 33320 5445
rect 33360 5437 33368 5445
rect 33552 5437 33560 5445
rect 33760 5437 33768 5445
rect 34560 5437 34568 5445
rect 34880 5437 34888 5445
rect 35456 5437 35464 5445
rect 35664 5437 35672 5445
rect 36464 5437 36472 5445
rect 36768 5437 36776 5445
rect 37504 5437 37512 5445
rect 38512 5437 38520 5445
rect 38576 5437 38584 5445
rect 38608 5437 38616 5445
rect 38879 5438 38886 5443
rect 39056 5437 39064 5445
rect 39184 5437 39192 5445
rect 39376 5437 39384 5445
rect 39472 5437 39480 5445
rect 19504 5420 19512 5428
rect 19920 5420 19928 5428
rect 20912 5420 20920 5428
rect 24240 5420 24248 5428
rect 29488 5417 29496 5425
rect 29840 5417 29848 5425
rect 30016 5417 30024 5425
rect 30192 5417 30200 5425
rect 30224 5417 30232 5425
rect 30240 5417 30248 5425
rect 30288 5417 30296 5425
rect 30512 5417 30520 5425
rect 30848 5417 30856 5425
rect 31120 5417 31128 5425
rect 31360 5417 31368 5425
rect 31504 5417 31512 5425
rect 31616 5417 31624 5425
rect 32032 5417 32040 5425
rect 33728 5417 33736 5425
rect 34016 5417 34024 5425
rect 34112 5417 34120 5425
rect 34960 5417 34968 5425
rect 35584 5417 35592 5425
rect 37152 5417 37160 5425
rect 39552 5417 39560 5425
rect 39648 5417 39656 5425
rect 39872 5417 39880 5425
rect 40128 5417 40136 5425
rect 40480 5417 40488 5425
rect 20896 5400 20904 5408
rect 21008 5400 21016 5408
rect 21104 5400 21112 5408
rect 23552 5400 23560 5408
rect 24672 5400 24680 5408
rect 25232 5400 25240 5408
rect 25264 5400 25272 5408
rect 26288 5400 26296 5408
rect 26368 5400 26376 5408
rect 30000 5397 30008 5405
rect 30496 5397 30504 5405
rect 30592 5397 30600 5405
rect 30928 5397 30936 5405
rect 31872 5397 31880 5405
rect 32720 5397 32728 5405
rect 33280 5397 33288 5405
rect 33504 5397 33512 5405
rect 34416 5397 34424 5405
rect 34864 5397 34872 5405
rect 35648 5397 35656 5405
rect 36672 5397 36680 5405
rect 37088 5397 37096 5405
rect 37344 5397 37352 5405
rect 37568 5397 37576 5405
rect 37664 5397 37672 5405
rect 37888 5397 37896 5405
rect 38144 5397 38152 5405
rect 38736 5397 38744 5405
rect 38896 5397 38904 5405
rect 40704 5397 40712 5405
rect 18528 5380 18536 5388
rect 19856 5380 19864 5388
rect 20064 5380 20072 5388
rect 20480 5380 20488 5388
rect 21984 5380 21992 5388
rect 22192 5380 22200 5388
rect 22368 5380 22376 5388
rect 22800 5380 22808 5388
rect 22960 5380 22968 5388
rect 23120 5380 23128 5388
rect 24080 5380 24088 5388
rect 24480 5380 24488 5388
rect 25872 5380 25880 5388
rect 26512 5380 26520 5388
rect 28064 5380 28072 5388
rect 28096 5380 28104 5388
rect 28208 5380 28216 5388
rect 29664 5377 29672 5385
rect 31232 5377 31240 5385
rect 32448 5377 32456 5385
rect 34352 5377 34360 5385
rect 36080 5377 36088 5385
rect 36112 5377 36120 5385
rect 38848 5377 38856 5385
rect 39792 5377 39800 5385
rect 39920 5377 39928 5385
rect 40272 5377 40280 5385
rect 40304 5377 40312 5385
rect 27008 5360 27016 5368
rect 30384 5357 30392 5365
rect 30672 5357 30680 5365
rect 32368 5357 32376 5365
rect 32784 5357 32792 5365
rect 32864 5357 32872 5365
rect 34752 5357 34760 5365
rect 35104 5357 35112 5365
rect 35920 5357 35928 5365
rect 37104 5357 37112 5365
rect 39936 5357 39944 5365
rect 40512 5357 40520 5365
rect 19072 5348 19076 5353
rect 19682 5348 19686 5353
rect 24068 5348 24077 5353
rect 25451 5348 25458 5353
rect 18864 5340 18872 5348
rect 20288 5340 20296 5348
rect 20496 5340 20504 5348
rect 21104 5340 21112 5348
rect 21920 5340 21928 5348
rect 23344 5340 23352 5348
rect 23776 5340 23784 5348
rect 25040 5340 25048 5348
rect 25888 5340 25896 5348
rect 26528 5340 26536 5348
rect 27024 5340 27032 5348
rect 27648 5340 27656 5348
rect 28080 5340 28088 5348
rect 28304 5340 28312 5348
rect 31408 5337 31416 5345
rect 39104 5337 39112 5345
rect 39232 5337 39240 5345
rect 39728 5337 39736 5345
rect 40400 5337 40408 5345
rect 22976 5320 22984 5328
rect 26096 5320 26104 5328
rect 30736 5317 30744 5325
rect 33920 5317 33928 5325
rect 37920 5317 37928 5325
rect 37936 5317 37944 5325
rect 20720 5300 20728 5308
rect 22736 5300 22744 5308
rect 27888 5300 27896 5308
rect 33776 5297 33784 5305
rect 31184 5277 31192 5285
rect 18912 5260 18920 5268
rect 19088 5260 19096 5268
rect 21744 5260 21752 5268
rect 25296 5260 25304 5268
rect 25696 5260 25704 5268
rect 29420 5267 29424 5275
rect 29428 5267 29440 5275
rect 29444 5267 29448 5275
rect 29460 5267 29472 5275
rect 29488 5267 29504 5275
rect 29520 5267 29544 5275
rect 29552 5267 29568 5275
rect 29576 5267 29600 5275
rect 29616 5267 29620 5275
rect 29624 5267 29636 5275
rect 29648 5267 29652 5275
rect 29656 5267 29660 5275
rect 29680 5267 29684 5275
rect 29688 5267 29692 5275
rect 29712 5267 29716 5275
rect 29720 5267 29724 5275
rect 29736 5267 29748 5275
rect 29752 5267 29756 5275
rect 29772 5267 29796 5275
rect 29804 5267 29820 5275
rect 29828 5267 29840 5275
rect 29844 5267 29848 5275
rect 29864 5267 29888 5275
rect 29896 5267 29912 5275
rect 29920 5267 29932 5275
rect 29936 5267 29940 5275
rect 29956 5267 29980 5275
rect 29988 5267 30004 5275
rect 30012 5267 30024 5275
rect 30028 5267 30032 5275
rect 30052 5267 30056 5275
rect 30060 5267 30072 5275
rect 30084 5267 30088 5275
rect 30092 5267 30096 5275
rect 30192 5267 30196 5275
rect 30200 5267 30204 5275
rect 30224 5267 30228 5275
rect 30232 5267 30236 5275
rect 30248 5267 30260 5275
rect 30264 5267 30268 5275
rect 30284 5267 30300 5275
rect 30316 5267 30364 5275
rect 30380 5267 30384 5275
rect 30388 5267 30392 5275
rect 30408 5267 30456 5275
rect 30468 5267 30484 5275
rect 30500 5267 30548 5275
rect 30564 5267 30568 5275
rect 30572 5267 30576 5275
rect 30592 5267 30640 5275
rect 30656 5267 30680 5275
rect 30688 5267 30704 5275
rect 30720 5267 30724 5275
rect 30728 5267 30732 5275
rect 30752 5267 30756 5275
rect 30760 5267 30772 5275
rect 30776 5267 30788 5275
rect 30792 5267 30796 5275
rect 30812 5267 30816 5275
rect 30820 5267 30824 5275
rect 30844 5267 30848 5275
rect 30852 5267 30864 5275
rect 30868 5267 30880 5275
rect 30884 5267 30888 5275
rect 30936 5267 30940 5275
rect 30944 5267 30956 5275
rect 30960 5267 30972 5275
rect 30976 5267 30980 5275
rect 31000 5267 31004 5275
rect 31008 5267 31020 5275
rect 31024 5267 31036 5275
rect 31040 5267 31044 5275
rect 31064 5267 31068 5275
rect 31072 5267 31076 5275
rect 31284 5267 31288 5275
rect 31292 5267 31296 5275
rect 31316 5267 31320 5275
rect 31324 5267 31336 5275
rect 31340 5267 31352 5275
rect 31356 5267 31360 5275
rect 31380 5267 31384 5275
rect 31388 5267 31392 5275
rect 31404 5267 31416 5275
rect 31436 5267 31448 5275
rect 31452 5267 31456 5275
rect 31468 5267 31480 5275
rect 31492 5267 31496 5275
rect 31500 5267 31512 5275
rect 31516 5267 31520 5275
rect 31532 5267 31544 5275
rect 31556 5267 31560 5275
rect 31564 5267 31576 5275
rect 31592 5267 31616 5275
rect 31624 5267 31640 5275
rect 31656 5267 31672 5275
rect 31688 5267 31704 5275
rect 31712 5267 31736 5275
rect 31752 5267 31764 5275
rect 31768 5267 31772 5275
rect 31784 5267 31796 5275
rect 31804 5267 31828 5275
rect 31844 5267 31868 5275
rect 31876 5267 31892 5275
rect 31908 5267 31912 5275
rect 31916 5267 31920 5275
rect 31940 5267 31944 5275
rect 31948 5267 31960 5275
rect 31964 5267 31976 5275
rect 31980 5267 31984 5275
rect 32004 5267 32008 5275
rect 32012 5267 32016 5275
rect 32028 5267 32040 5275
rect 32056 5267 32072 5275
rect 32088 5267 32120 5275
rect 32128 5267 32140 5275
rect 32160 5267 32172 5275
rect 32184 5267 32188 5275
rect 32192 5267 32196 5275
rect 32216 5267 32220 5275
rect 32224 5267 32228 5275
rect 32248 5267 32252 5275
rect 32256 5267 32260 5275
rect 32272 5267 32284 5275
rect 32288 5267 32292 5275
rect 32308 5267 32332 5275
rect 32348 5267 32360 5275
rect 32364 5267 32368 5275
rect 32380 5267 32392 5275
rect 32404 5267 32408 5275
rect 32412 5267 32424 5275
rect 32444 5267 32456 5275
rect 32476 5267 32488 5275
rect 32508 5267 32520 5275
rect 32524 5267 32528 5275
rect 32540 5267 32552 5275
rect 32560 5267 32584 5275
rect 32600 5267 32612 5275
rect 32616 5267 32620 5275
rect 32632 5267 32644 5275
rect 32656 5267 32660 5275
rect 32664 5267 32676 5275
rect 32764 5267 32768 5275
rect 32772 5267 32784 5275
rect 32796 5267 32800 5275
rect 32804 5267 32808 5275
rect 32820 5267 32832 5275
rect 32848 5267 32860 5275
rect 32872 5267 32876 5275
rect 32880 5267 32892 5275
rect 32896 5267 32900 5275
rect 32912 5267 32924 5275
rect 32944 5267 32956 5275
rect 32960 5267 32964 5275
rect 32984 5267 32988 5275
rect 32992 5267 32996 5275
rect 33016 5267 33020 5275
rect 33024 5267 33036 5275
rect 33048 5267 33052 5275
rect 33056 5267 33060 5275
rect 33080 5267 33084 5275
rect 33088 5267 33092 5275
rect 33124 5267 33128 5275
rect 33132 5267 33144 5275
rect 33164 5267 33176 5275
rect 33180 5267 33184 5275
rect 33196 5267 33208 5275
rect 33224 5267 33240 5275
rect 33256 5267 33304 5275
rect 33320 5267 33324 5275
rect 33328 5267 33332 5275
rect 33344 5267 33356 5275
rect 33360 5267 33372 5275
rect 33384 5267 33388 5275
rect 33392 5267 33396 5275
rect 33492 5267 33496 5275
rect 33500 5267 33512 5275
rect 33524 5267 33528 5275
rect 33532 5267 33536 5275
rect 33548 5267 33560 5275
rect 33564 5267 33568 5275
rect 33584 5267 33588 5275
rect 33592 5267 33600 5275
rect 33616 5267 33620 5275
rect 33624 5267 33628 5275
rect 33756 5267 33760 5275
rect 33764 5267 33776 5275
rect 33780 5267 33792 5275
rect 33796 5267 33800 5275
rect 33992 5267 33996 5275
rect 34000 5267 34012 5275
rect 34016 5267 34028 5275
rect 34032 5267 34036 5275
rect 34056 5267 34060 5275
rect 34064 5267 34076 5275
rect 34084 5267 34100 5275
rect 34108 5267 34132 5275
rect 34148 5267 34164 5275
rect 34180 5267 34196 5275
rect 34212 5267 34236 5275
rect 34244 5267 34260 5275
rect 34268 5267 34300 5275
rect 34308 5267 34324 5275
rect 34336 5267 34352 5275
rect 34360 5267 34392 5275
rect 34400 5267 34416 5275
rect 34432 5267 34436 5275
rect 34440 5267 34444 5275
rect 34464 5267 34468 5275
rect 34472 5267 34484 5275
rect 34496 5267 34500 5275
rect 34504 5267 34508 5275
rect 34680 5267 34684 5275
rect 34688 5267 34692 5275
rect 34712 5267 34716 5275
rect 34720 5267 34724 5275
rect 34796 5267 34808 5275
rect 34812 5267 34816 5275
rect 34832 5267 34836 5275
rect 34840 5267 34852 5275
rect 34864 5267 34868 5275
rect 34872 5267 34876 5275
rect 34888 5267 34900 5275
rect 34916 5267 34928 5275
rect 34940 5267 34944 5275
rect 34948 5267 34960 5275
rect 34964 5267 34968 5275
rect 34984 5267 35008 5275
rect 35016 5267 35032 5275
rect 35040 5267 35052 5275
rect 35056 5267 35060 5275
rect 35076 5267 35100 5275
rect 35108 5267 35124 5275
rect 35132 5267 35156 5275
rect 35172 5267 35188 5275
rect 35204 5267 35220 5275
rect 35236 5267 35260 5275
rect 35268 5267 35284 5275
rect 35292 5267 35304 5275
rect 35308 5267 35312 5275
rect 35332 5267 35336 5275
rect 35340 5267 35352 5275
rect 35356 5267 35368 5275
rect 35372 5267 35376 5275
rect 35396 5267 35400 5275
rect 35404 5267 35416 5275
rect 35428 5267 35432 5275
rect 35436 5267 35440 5275
rect 35460 5267 35464 5275
rect 35468 5267 35472 5275
rect 35492 5267 35496 5275
rect 35500 5267 35504 5275
rect 35516 5267 35528 5275
rect 35532 5267 35536 5275
rect 35556 5267 35560 5275
rect 35564 5267 35576 5275
rect 35580 5267 35592 5275
rect 35596 5267 35600 5275
rect 35616 5267 35640 5275
rect 35648 5267 35664 5275
rect 35672 5267 35704 5275
rect 35712 5267 35724 5275
rect 35744 5267 35756 5275
rect 35764 5267 35796 5275
rect 35804 5267 35816 5275
rect 35832 5267 35848 5275
rect 35856 5267 35888 5275
rect 35896 5267 35908 5275
rect 35928 5267 35940 5275
rect 35948 5267 35980 5275
rect 35988 5267 36000 5275
rect 36016 5267 36032 5275
rect 36040 5267 36072 5275
rect 36080 5267 36096 5275
rect 36112 5267 36136 5275
rect 36144 5267 36160 5275
rect 36176 5267 36224 5275
rect 36240 5267 36288 5275
rect 36304 5267 36308 5275
rect 36312 5267 36316 5275
rect 36332 5267 36380 5275
rect 36396 5267 36408 5275
rect 36424 5267 36472 5275
rect 36488 5267 36504 5275
rect 36512 5267 36536 5275
rect 36552 5267 36564 5275
rect 36584 5267 36596 5275
rect 36600 5267 36612 5275
rect 36616 5267 36628 5275
rect 36772 5267 36784 5275
rect 36788 5267 36800 5275
rect 36804 5267 36816 5275
rect 36832 5267 36848 5275
rect 36864 5267 36888 5275
rect 36896 5267 36912 5275
rect 36928 5267 36932 5275
rect 36936 5267 36940 5275
rect 36952 5267 36964 5275
rect 36968 5267 36980 5275
rect 36988 5267 37004 5275
rect 37020 5267 37024 5275
rect 37028 5267 37032 5275
rect 37044 5267 37056 5275
rect 37060 5267 37072 5275
rect 37084 5267 37088 5275
rect 37092 5267 37096 5275
rect 37116 5267 37120 5275
rect 37124 5267 37128 5275
rect 37192 5267 37196 5275
rect 37200 5267 37212 5275
rect 37224 5267 37228 5275
rect 37232 5267 37236 5275
rect 37284 5267 37288 5275
rect 37292 5267 37304 5275
rect 37316 5267 37320 5275
rect 37324 5267 37328 5275
rect 37376 5267 37380 5275
rect 37384 5267 37396 5275
rect 37408 5267 37412 5275
rect 37416 5267 37420 5275
rect 37432 5267 37444 5275
rect 37448 5267 37460 5275
rect 37472 5267 37476 5275
rect 37480 5267 37484 5275
rect 37496 5267 37508 5275
rect 37512 5267 37524 5275
rect 37532 5267 37548 5275
rect 37564 5267 37612 5275
rect 37628 5267 37640 5275
rect 37644 5267 37648 5275
rect 37660 5267 37672 5275
rect 37684 5267 37688 5275
rect 37692 5267 37704 5275
rect 37724 5267 37736 5275
rect 37808 5267 37812 5275
rect 37816 5267 37828 5275
rect 37940 5267 37952 5275
rect 37956 5267 37960 5275
rect 37972 5267 37984 5275
rect 38000 5267 38016 5275
rect 38032 5267 38080 5275
rect 38096 5267 38112 5275
rect 38120 5267 38144 5275
rect 38160 5267 38172 5275
rect 38192 5267 38204 5275
rect 38208 5267 38220 5275
rect 38224 5267 38236 5275
rect 38256 5267 38268 5275
rect 38348 5267 38360 5275
rect 38372 5267 38376 5275
rect 38380 5267 38392 5275
rect 38396 5267 38400 5275
rect 38412 5267 38424 5275
rect 38600 5267 38612 5275
rect 38624 5267 38628 5275
rect 38632 5267 38644 5275
rect 38648 5267 38652 5275
rect 38788 5267 38800 5275
rect 38804 5267 38816 5275
rect 38820 5267 38832 5275
rect 39008 5267 39020 5275
rect 39040 5267 39052 5275
rect 39056 5267 39068 5275
rect 39072 5267 39084 5275
rect 39100 5267 39116 5275
rect 39124 5267 39156 5275
rect 39164 5267 39180 5275
rect 39200 5267 39208 5275
rect 39220 5267 39224 5275
rect 39228 5267 39240 5275
rect 39260 5267 39272 5275
rect 39292 5267 39304 5275
rect 39308 5267 39312 5275
rect 39324 5267 39336 5275
rect 39356 5267 39368 5275
rect 39376 5267 39408 5275
rect 39416 5267 39428 5275
rect 39448 5267 39460 5275
rect 39464 5267 39476 5275
rect 39480 5267 39492 5275
rect 39512 5267 39524 5275
rect 39540 5267 39564 5275
rect 39572 5267 39588 5275
rect 39604 5267 39652 5275
rect 39668 5267 39672 5275
rect 39676 5267 39680 5275
rect 39692 5267 39704 5275
rect 39708 5267 39720 5275
rect 39732 5267 39736 5275
rect 39740 5267 39744 5275
rect 39760 5267 39776 5275
rect 39784 5267 39808 5275
rect 39824 5267 39840 5275
rect 39856 5267 39868 5275
rect 39872 5267 39884 5275
rect 39888 5267 39900 5275
rect 39916 5267 39932 5275
rect 39948 5267 39972 5275
rect 39980 5267 39996 5275
rect 40012 5267 40028 5275
rect 40036 5267 40060 5275
rect 40076 5267 40092 5275
rect 40100 5267 40132 5275
rect 40140 5267 40156 5275
rect 40164 5267 40188 5275
rect 40200 5267 40224 5275
rect 40232 5267 40248 5275
rect 40256 5267 40280 5275
rect 40292 5267 40316 5275
rect 40324 5267 40340 5275
rect 40348 5267 40372 5275
rect 40388 5267 40404 5275
rect 40412 5267 40436 5275
rect 40452 5267 40464 5275
rect 40468 5267 40472 5275
rect 40484 5267 40496 5275
rect 40508 5267 40512 5275
rect 40516 5267 40528 5275
rect 40724 5267 40728 5275
rect 40732 5267 40744 5275
rect 20020 5250 20022 5258
rect 20028 5250 20030 5258
rect 20226 5250 20236 5258
rect 20440 5250 20450 5258
rect 21218 5250 21230 5258
rect 21416 5250 21428 5258
rect 21850 5250 21856 5258
rect 21858 5250 21864 5258
rect 21926 5250 21932 5258
rect 21934 5250 21940 5258
rect 22476 5250 22482 5258
rect 22484 5250 22490 5258
rect 22552 5250 22558 5258
rect 22560 5250 22566 5258
rect 22774 5250 22786 5258
rect 22850 5250 22862 5258
rect 23820 5250 23826 5258
rect 23828 5250 23834 5258
rect 24034 5250 24040 5258
rect 24042 5250 24048 5258
rect 24248 5250 24254 5258
rect 24256 5250 24262 5258
rect 24462 5250 24468 5258
rect 24470 5250 24476 5258
rect 26150 5250 26164 5258
rect 26470 5250 26484 5258
rect 26792 5250 26806 5258
rect 27006 5250 27020 5258
rect 27632 5250 27646 5258
rect 30752 5237 30760 5245
rect 31200 5237 31208 5245
rect 31216 5237 31224 5245
rect 31344 5237 31352 5245
rect 36192 5237 36200 5245
rect 36592 5237 36600 5245
rect 36768 5237 36776 5245
rect 31456 5217 31464 5225
rect 32848 5217 32856 5225
rect 34544 5217 34552 5225
rect 34640 5217 34648 5225
rect 34768 5217 34776 5225
rect 35312 5217 35320 5225
rect 35664 5217 35672 5225
rect 35952 5217 35960 5225
rect 36752 5217 36760 5225
rect 37312 5217 37320 5225
rect 23296 5200 23304 5208
rect 25696 5200 25704 5208
rect 28208 5200 28216 5208
rect 32320 5197 32328 5205
rect 38368 5197 38376 5205
rect 39696 5197 39704 5205
rect 19952 5180 19960 5188
rect 29568 5177 29576 5185
rect 30208 5177 30216 5185
rect 30304 5177 30312 5185
rect 31920 5177 31928 5185
rect 32816 5177 32824 5185
rect 33472 5177 33480 5185
rect 33648 5177 33656 5185
rect 34624 5177 34632 5185
rect 35056 5177 35064 5185
rect 35728 5177 35736 5185
rect 35840 5177 35848 5185
rect 36064 5177 36072 5185
rect 36512 5177 36520 5185
rect 37856 5177 37864 5185
rect 18656 5160 18664 5168
rect 18848 5160 18856 5168
rect 18892 5161 18902 5166
rect 19744 5160 19752 5168
rect 20592 5160 20600 5168
rect 20800 5160 20808 5168
rect 20816 5160 20824 5168
rect 21024 5160 21032 5168
rect 21184 5160 21192 5168
rect 21230 5161 21240 5166
rect 21440 5160 21448 5168
rect 21824 5160 21832 5168
rect 22048 5160 22056 5168
rect 22080 5160 22088 5168
rect 22432 5161 22442 5166
rect 23840 5160 23848 5168
rect 24144 5160 24152 5168
rect 24400 5160 24408 5168
rect 24624 5160 24632 5168
rect 25840 5160 25848 5168
rect 26096 5160 26104 5168
rect 26736 5160 26744 5168
rect 26960 5160 26968 5168
rect 28160 5160 28168 5168
rect 30704 5157 30712 5165
rect 31648 5157 31656 5165
rect 31696 5157 31704 5165
rect 32032 5157 32040 5165
rect 32704 5157 32712 5165
rect 38512 5157 38520 5165
rect 39920 5157 39928 5165
rect 39952 5157 39960 5165
rect 23008 5140 23016 5148
rect 25920 5140 25928 5148
rect 26256 5140 26264 5148
rect 29712 5137 29720 5145
rect 29952 5137 29960 5145
rect 30544 5137 30552 5145
rect 30688 5137 30696 5145
rect 30880 5137 30888 5145
rect 31328 5137 31336 5145
rect 32928 5137 32936 5145
rect 35072 5137 35080 5145
rect 35712 5137 35720 5145
rect 36640 5137 36648 5145
rect 37824 5137 37832 5145
rect 38000 5137 38008 5145
rect 38096 5137 38104 5145
rect 38192 5137 38200 5145
rect 38992 5137 39000 5145
rect 39136 5137 39144 5145
rect 39456 5137 39464 5145
rect 39712 5137 39720 5145
rect 40336 5137 40344 5145
rect 40608 5137 40616 5145
rect 18640 5120 18648 5128
rect 19536 5120 19544 5128
rect 19760 5120 19768 5128
rect 20400 5120 20408 5128
rect 20608 5120 20616 5128
rect 21888 5120 21896 5128
rect 22096 5120 22104 5128
rect 23056 5120 23064 5128
rect 23136 5120 23144 5128
rect 23984 5120 23992 5128
rect 24416 5120 24424 5128
rect 24848 5120 24856 5128
rect 25248 5120 25256 5128
rect 26112 5120 26120 5128
rect 26176 5120 26184 5128
rect 26752 5120 26760 5128
rect 27520 5120 27528 5128
rect 28352 5120 28360 5128
rect 29376 5117 29384 5125
rect 31248 5117 31256 5125
rect 31424 5117 31432 5125
rect 31440 5117 31448 5125
rect 31504 5117 31512 5125
rect 31600 5117 31608 5125
rect 32224 5117 32232 5125
rect 32544 5117 32552 5125
rect 32912 5117 32920 5125
rect 35136 5117 35144 5125
rect 35456 5117 35464 5125
rect 36176 5117 36184 5125
rect 36704 5117 36712 5125
rect 36912 5117 36920 5125
rect 39072 5117 39080 5125
rect 39472 5117 39480 5125
rect 39760 5117 39768 5125
rect 40368 5117 40376 5125
rect 18912 5100 18920 5108
rect 19120 5100 19128 5108
rect 21616 5100 21624 5108
rect 23120 5100 23128 5108
rect 25824 5100 25832 5108
rect 26624 5100 26632 5108
rect 26896 5100 26904 5108
rect 27536 5100 27544 5108
rect 31056 5097 31064 5105
rect 31088 5097 31096 5105
rect 34128 5097 34136 5105
rect 34912 5097 34920 5105
rect 35232 5097 35240 5105
rect 20784 5080 20792 5088
rect 24560 5080 24568 5088
rect 33456 5077 33464 5085
rect 33584 5077 33592 5085
rect 33888 5077 33896 5085
rect 33904 5077 33912 5085
rect 33952 5077 33960 5085
rect 34224 5077 34232 5085
rect 34832 5077 34840 5085
rect 35264 5077 35272 5085
rect 37440 5077 37448 5085
rect 38032 5077 38040 5085
rect 38144 5077 38152 5085
rect 38160 5077 38168 5085
rect 19056 5060 19064 5068
rect 19280 5060 19288 5068
rect 19472 5060 19480 5068
rect 27984 5060 27992 5068
rect 29428 5067 29440 5075
rect 29444 5067 29448 5075
rect 29460 5067 29472 5075
rect 29488 5067 29504 5075
rect 29512 5067 29544 5075
rect 29552 5067 29564 5075
rect 29584 5067 29596 5075
rect 29604 5067 29636 5075
rect 29644 5067 29660 5075
rect 29676 5067 29688 5075
rect 29700 5067 29704 5075
rect 29708 5067 29720 5075
rect 29740 5067 29752 5075
rect 29832 5067 29844 5075
rect 29856 5067 29860 5075
rect 29864 5067 29876 5075
rect 29880 5067 29884 5075
rect 29896 5067 29908 5075
rect 29924 5067 29940 5075
rect 29956 5067 29980 5075
rect 29988 5067 30004 5075
rect 30012 5067 30024 5075
rect 30028 5067 30032 5075
rect 30052 5067 30056 5075
rect 30060 5067 30072 5075
rect 30080 5067 30096 5075
rect 30104 5067 30116 5075
rect 30120 5067 30124 5075
rect 30144 5067 30148 5075
rect 30152 5067 30164 5075
rect 30176 5067 30180 5075
rect 30184 5067 30188 5075
rect 30284 5067 30288 5075
rect 30292 5067 30296 5075
rect 30316 5067 30320 5075
rect 30324 5067 30336 5075
rect 30340 5067 30352 5075
rect 30356 5067 30360 5075
rect 30380 5067 30384 5075
rect 30388 5067 30392 5075
rect 30408 5067 30424 5075
rect 30432 5067 30456 5075
rect 30472 5067 30484 5075
rect 30488 5067 30492 5075
rect 30504 5067 30516 5075
rect 30528 5067 30532 5075
rect 30536 5067 30548 5075
rect 30564 5067 30588 5075
rect 30596 5067 30608 5075
rect 30620 5067 30624 5075
rect 30628 5067 30640 5075
rect 30656 5067 30680 5075
rect 30688 5067 30704 5075
rect 30720 5067 30736 5075
rect 30752 5067 30756 5075
rect 30760 5067 30772 5075
rect 30776 5067 30788 5075
rect 30792 5067 30796 5075
rect 30812 5067 30828 5075
rect 30844 5067 30848 5075
rect 30852 5067 30864 5075
rect 30868 5067 30880 5075
rect 30884 5067 30888 5075
rect 30908 5067 30912 5075
rect 30916 5067 30920 5075
rect 30936 5067 30952 5075
rect 30960 5067 30984 5075
rect 31000 5067 31048 5075
rect 31064 5067 31080 5075
rect 31096 5067 31100 5075
rect 31104 5067 31116 5075
rect 31128 5067 31132 5075
rect 31136 5067 31140 5075
rect 31284 5067 31288 5075
rect 31292 5067 31296 5075
rect 31316 5067 31320 5075
rect 31324 5067 31328 5075
rect 31340 5067 31352 5075
rect 31356 5067 31360 5075
rect 31380 5067 31384 5075
rect 31388 5067 31392 5075
rect 31404 5067 31416 5075
rect 31428 5067 31432 5075
rect 31436 5067 31448 5075
rect 31452 5067 31456 5075
rect 31560 5067 31572 5075
rect 31652 5067 31664 5075
rect 31684 5067 31696 5075
rect 31700 5067 31704 5075
rect 31716 5067 31728 5075
rect 31748 5067 31760 5075
rect 31768 5067 31800 5075
rect 31808 5067 31820 5075
rect 31840 5067 31852 5075
rect 31860 5067 31892 5075
rect 31900 5067 31912 5075
rect 31932 5067 31944 5075
rect 31948 5067 31960 5075
rect 31964 5067 31976 5075
rect 32000 5067 32008 5075
rect 32024 5067 32048 5075
rect 32056 5067 32072 5075
rect 32088 5067 32136 5075
rect 32152 5067 32156 5075
rect 32160 5067 32164 5075
rect 32184 5067 32188 5075
rect 32192 5067 32204 5075
rect 32216 5067 32220 5075
rect 32224 5067 32228 5075
rect 32308 5067 32312 5075
rect 32316 5067 32320 5075
rect 32340 5067 32344 5075
rect 32348 5067 32352 5075
rect 32416 5067 32420 5075
rect 32424 5067 32428 5075
rect 32448 5067 32452 5075
rect 32456 5067 32460 5075
rect 32472 5067 32484 5075
rect 32488 5067 32492 5075
rect 32512 5067 32516 5075
rect 32520 5067 32532 5075
rect 32540 5067 32556 5075
rect 32564 5067 32576 5075
rect 32580 5067 32584 5075
rect 32604 5067 32608 5075
rect 32612 5067 32624 5075
rect 32632 5067 32648 5075
rect 32656 5067 32680 5075
rect 32696 5067 32712 5075
rect 32728 5067 32740 5075
rect 32752 5067 32756 5075
rect 32760 5067 32772 5075
rect 32776 5067 32780 5075
rect 32792 5067 32800 5075
rect 32844 5067 32848 5075
rect 32852 5067 32864 5075
rect 32868 5067 32872 5075
rect 33008 5067 33020 5075
rect 33024 5067 33036 5075
rect 33040 5067 33052 5075
rect 33072 5067 33084 5075
rect 33100 5067 33112 5075
rect 33116 5067 33128 5075
rect 33132 5067 33144 5075
rect 33164 5067 33176 5075
rect 33192 5067 33216 5075
rect 33224 5067 33240 5075
rect 33256 5067 33272 5075
rect 33280 5067 33292 5075
rect 33296 5067 33308 5075
rect 33320 5067 33324 5075
rect 33328 5067 33332 5075
rect 33344 5067 33356 5075
rect 33360 5067 33364 5075
rect 33460 5067 33464 5075
rect 33468 5067 33472 5075
rect 33484 5067 33496 5075
rect 33500 5067 33512 5075
rect 33524 5067 33528 5075
rect 33532 5067 33536 5075
rect 33552 5067 33568 5075
rect 33576 5067 33588 5075
rect 33592 5067 33600 5075
rect 33616 5067 33620 5075
rect 33624 5067 33628 5075
rect 33756 5067 33760 5075
rect 33764 5067 33768 5075
rect 33780 5067 33792 5075
rect 33796 5067 33800 5075
rect 33896 5067 33900 5075
rect 33904 5067 33908 5075
rect 33920 5067 33932 5075
rect 33936 5067 33940 5075
rect 33960 5067 33964 5075
rect 33968 5067 33972 5075
rect 33988 5067 34036 5075
rect 34052 5067 34076 5075
rect 34084 5067 34096 5075
rect 34108 5067 34112 5075
rect 34116 5067 34128 5075
rect 34148 5067 34160 5075
rect 34172 5067 34176 5075
rect 34180 5067 34192 5075
rect 34212 5067 34224 5075
rect 34228 5067 34240 5075
rect 34244 5067 34256 5075
rect 34276 5067 34288 5075
rect 34292 5067 34296 5075
rect 34308 5067 34320 5075
rect 34336 5067 34352 5075
rect 34368 5067 34416 5075
rect 34432 5067 34436 5075
rect 34440 5067 34444 5075
rect 34456 5067 34468 5075
rect 34472 5067 34484 5075
rect 34496 5067 34500 5075
rect 34504 5067 34508 5075
rect 34604 5067 34608 5075
rect 34612 5067 34624 5075
rect 34636 5067 34640 5075
rect 34644 5067 34648 5075
rect 34660 5067 34672 5075
rect 34676 5067 34688 5075
rect 34700 5067 34704 5075
rect 34708 5067 34712 5075
rect 34728 5067 34744 5075
rect 34752 5067 34776 5075
rect 34792 5067 34808 5075
rect 34824 5067 34836 5075
rect 34840 5067 34852 5075
rect 34856 5067 34868 5075
rect 34888 5067 34900 5075
rect 34904 5067 34908 5075
rect 34980 5067 34992 5075
rect 34996 5067 35008 5075
rect 35012 5067 35024 5075
rect 35072 5067 35084 5075
rect 35088 5067 35100 5075
rect 35104 5067 35116 5075
rect 35136 5067 35148 5075
rect 35164 5067 35188 5075
rect 35200 5067 35212 5075
rect 35228 5067 35244 5075
rect 35252 5067 35264 5075
rect 35268 5067 35280 5075
rect 35288 5067 35304 5075
rect 35320 5067 35336 5075
rect 35344 5067 35356 5075
rect 35360 5067 35372 5075
rect 35384 5067 35388 5075
rect 35392 5067 35396 5075
rect 35408 5067 35420 5075
rect 35424 5067 35428 5075
rect 35764 5067 35768 5075
rect 35772 5067 35776 5075
rect 35788 5067 35800 5075
rect 35804 5067 35816 5075
rect 35824 5067 35840 5075
rect 35856 5067 35872 5075
rect 35880 5067 35904 5075
rect 35920 5067 35936 5075
rect 35952 5067 35964 5075
rect 35968 5067 35980 5075
rect 35984 5067 35996 5075
rect 36012 5067 36024 5075
rect 36044 5067 36056 5075
rect 36060 5067 36072 5075
rect 36076 5067 36088 5075
rect 36108 5067 36120 5075
rect 36128 5067 36160 5075
rect 36168 5067 36184 5075
rect 36192 5067 36216 5075
rect 36232 5067 36248 5075
rect 36256 5067 36280 5075
rect 36296 5067 36308 5075
rect 36312 5067 36316 5075
rect 36328 5067 36340 5075
rect 36352 5067 36356 5075
rect 36360 5067 36372 5075
rect 36388 5067 36412 5075
rect 36420 5067 36432 5075
rect 36440 5067 36464 5075
rect 36480 5067 36504 5075
rect 36512 5067 36528 5075
rect 36544 5067 36548 5075
rect 36552 5067 36556 5075
rect 36576 5067 36580 5075
rect 36584 5067 36596 5075
rect 36600 5067 36612 5075
rect 36616 5067 36620 5075
rect 36640 5067 36644 5075
rect 36648 5067 36652 5075
rect 36812 5067 36816 5075
rect 36820 5067 36824 5075
rect 36836 5067 36848 5075
rect 36852 5067 36856 5075
rect 36872 5067 36888 5075
rect 36904 5067 36920 5075
rect 36928 5067 36960 5075
rect 36968 5067 36984 5075
rect 36996 5067 37012 5075
rect 37020 5067 37052 5075
rect 37060 5067 37076 5075
rect 37092 5067 37104 5075
rect 37116 5067 37120 5075
rect 37124 5067 37136 5075
rect 37156 5067 37168 5075
rect 37180 5067 37184 5075
rect 37188 5067 37200 5075
rect 37204 5067 37208 5075
rect 37248 5067 37260 5075
rect 37272 5067 37276 5075
rect 37280 5067 37292 5075
rect 37296 5067 37300 5075
rect 37312 5067 37324 5075
rect 37340 5067 37352 5075
rect 37364 5067 37368 5075
rect 37372 5067 37384 5075
rect 37388 5067 37392 5075
rect 37404 5067 37416 5075
rect 37648 5067 37652 5075
rect 37656 5067 37668 5075
rect 37688 5067 37700 5075
rect 37704 5067 37708 5075
rect 37720 5067 37732 5075
rect 37748 5067 37764 5075
rect 37780 5067 37828 5075
rect 37844 5067 37856 5075
rect 37872 5067 37920 5075
rect 37936 5067 37952 5075
rect 37968 5067 37972 5075
rect 37976 5067 37988 5075
rect 38000 5067 38004 5075
rect 38008 5067 38012 5075
rect 38032 5067 38036 5075
rect 38040 5067 38052 5075
rect 38056 5067 38068 5075
rect 38072 5067 38076 5075
rect 38156 5067 38160 5075
rect 38164 5067 38168 5075
rect 38280 5067 38284 5075
rect 38288 5067 38292 5075
rect 38304 5067 38316 5075
rect 38320 5067 38324 5075
rect 38340 5067 38356 5075
rect 38372 5067 38420 5075
rect 38436 5067 38440 5075
rect 38444 5067 38448 5075
rect 38468 5067 38472 5075
rect 38476 5067 38488 5075
rect 38500 5067 38504 5075
rect 38508 5067 38512 5075
rect 38592 5067 38596 5075
rect 38600 5067 38604 5075
rect 38732 5067 38736 5075
rect 38740 5067 38744 5075
rect 38756 5067 38768 5075
rect 38772 5067 38776 5075
rect 38796 5067 38800 5075
rect 38804 5067 38816 5075
rect 38824 5067 38840 5075
rect 38848 5067 38860 5075
rect 38864 5067 38868 5075
rect 38888 5067 38892 5075
rect 38896 5067 38908 5075
rect 38916 5067 38932 5075
rect 38940 5067 38964 5075
rect 38980 5067 38992 5075
rect 39012 5067 39024 5075
rect 39036 5067 39040 5075
rect 39044 5067 39056 5075
rect 39060 5067 39064 5075
rect 39292 5067 39304 5075
rect 39308 5067 39312 5075
rect 39324 5067 39336 5075
rect 39356 5067 39368 5075
rect 39372 5067 39384 5075
rect 39388 5067 39400 5075
rect 39448 5067 39460 5075
rect 39464 5067 39476 5075
rect 39480 5067 39492 5075
rect 39512 5067 39524 5075
rect 39540 5067 39564 5075
rect 39572 5067 39588 5075
rect 39604 5067 39620 5075
rect 39628 5067 39640 5075
rect 39644 5067 39656 5075
rect 39668 5067 39672 5075
rect 39676 5067 39680 5075
rect 39760 5067 39764 5075
rect 39768 5067 39772 5075
rect 39784 5067 39796 5075
rect 39800 5067 39804 5075
rect 39852 5067 39856 5075
rect 39860 5067 39864 5075
rect 39876 5067 39888 5075
rect 39892 5067 39896 5075
rect 39916 5067 39920 5075
rect 39924 5067 39928 5075
rect 39948 5067 39952 5075
rect 39956 5067 39960 5075
rect 39980 5067 39984 5075
rect 39988 5067 40000 5075
rect 40012 5067 40016 5075
rect 40020 5067 40024 5075
rect 40036 5067 40048 5075
rect 40052 5067 40056 5075
rect 40200 5067 40204 5075
rect 40208 5067 40212 5075
rect 40232 5067 40236 5075
rect 40240 5067 40252 5075
rect 40256 5067 40268 5075
rect 40272 5067 40276 5075
rect 40292 5067 40308 5075
rect 40324 5067 40340 5075
rect 40348 5067 40372 5075
rect 40388 5067 40436 5075
rect 40452 5067 40464 5075
rect 40468 5067 40472 5075
rect 40484 5067 40496 5075
rect 40504 5067 40528 5075
rect 40544 5067 40556 5075
rect 40560 5067 40564 5075
rect 40576 5067 40588 5075
rect 40600 5067 40604 5075
rect 40608 5067 40620 5075
rect 40624 5067 40628 5075
rect 40640 5067 40652 5075
rect 40732 5067 40744 5075
rect 40764 5067 40776 5075
rect 40780 5067 40792 5075
rect 40796 5067 40800 5075
rect 18938 5050 18942 5058
rect 19028 5050 19036 5058
rect 19136 5050 19140 5058
rect 19226 5050 19234 5058
rect 19724 5050 19732 5058
rect 19874 5050 19880 5058
rect 19938 5050 19946 5058
rect 20088 5050 20094 5058
rect 20152 5050 20160 5058
rect 20302 5050 20308 5058
rect 20366 5050 20380 5058
rect 21008 5050 21022 5058
rect 21222 5050 21236 5058
rect 21420 5050 21428 5058
rect 21570 5050 21576 5058
rect 22474 5050 22482 5058
rect 22624 5050 22630 5058
rect 22710 5050 22714 5058
rect 22800 5050 22808 5058
rect 23224 5052 23226 5060
rect 24080 5052 24082 5060
rect 24294 5052 24296 5060
rect 24508 5052 24510 5060
rect 24722 5052 24724 5060
rect 25048 5050 25052 5058
rect 25138 5050 25146 5058
rect 25348 5052 25350 5060
rect 25562 5052 25564 5060
rect 25776 5052 25778 5060
rect 26722 5050 26730 5058
rect 26872 5050 26878 5058
rect 28332 5050 28346 5058
rect 28418 5050 28432 5058
rect 22224 5040 22232 5048
rect 22832 5040 22840 5048
rect 28160 5040 28168 5048
rect 31024 5037 31032 5045
rect 31600 5037 31608 5045
rect 32064 5037 32072 5045
rect 37152 5037 37160 5045
rect 40464 5037 40472 5045
rect 19488 5020 19496 5028
rect 21376 5020 21384 5028
rect 21776 5020 21784 5028
rect 23504 5020 23512 5028
rect 24736 5020 24744 5028
rect 26176 5020 26184 5028
rect 27344 5020 27352 5028
rect 27744 5020 27752 5028
rect 29488 5017 29496 5025
rect 29872 5017 29880 5025
rect 30768 5017 30776 5025
rect 30880 5017 30888 5025
rect 31376 5017 31384 5025
rect 31536 5017 31544 5025
rect 33696 5017 33704 5025
rect 33744 5017 33752 5025
rect 35296 5017 35304 5025
rect 35504 5017 35512 5025
rect 35536 5017 35544 5025
rect 35600 5017 35608 5025
rect 35648 5017 35656 5025
rect 35824 5017 35832 5025
rect 35984 5017 35992 5025
rect 36000 5017 36008 5025
rect 36144 5017 36152 5025
rect 38304 5017 38312 5025
rect 40016 5017 40024 5025
rect 40176 5017 40184 5025
rect 40576 5017 40584 5025
rect 20512 5000 20520 5008
rect 20544 5000 20552 5008
rect 22176 5000 22184 5008
rect 22432 5000 22440 5008
rect 25168 5000 25176 5008
rect 26288 5000 26296 5008
rect 27344 5000 27352 5008
rect 29616 4997 29624 5005
rect 29712 4997 29720 5005
rect 29792 4997 29800 5005
rect 30592 4997 30600 5005
rect 31328 4997 31336 5005
rect 31584 4997 31592 5005
rect 31712 4997 31720 5005
rect 32768 4997 32776 5005
rect 33312 4997 33320 5005
rect 34560 4997 34568 5005
rect 35008 4997 35016 5005
rect 35104 4997 35112 5005
rect 35200 4997 35208 5005
rect 35376 4997 35384 5005
rect 35504 4997 35512 5005
rect 36384 4997 36392 5005
rect 36944 4997 36952 5005
rect 37280 4997 37288 5005
rect 37376 4997 37384 5005
rect 37904 4997 37912 5005
rect 38048 4997 38056 5005
rect 38288 4997 38296 5005
rect 38464 4997 38472 5005
rect 38992 4997 39000 5005
rect 39136 4997 39144 5005
rect 39232 4997 39240 5005
rect 39568 4997 39576 5005
rect 18720 4980 18728 4988
rect 19056 4980 19064 4988
rect 20272 4980 20280 4988
rect 21536 4980 21544 4988
rect 21616 4980 21624 4988
rect 22160 4980 22168 4988
rect 22592 4980 22600 4988
rect 23872 4980 23880 4988
rect 24160 4980 24168 4988
rect 24192 4980 24200 4988
rect 24208 4980 24216 4988
rect 24608 4980 24616 4988
rect 24816 4980 24824 4988
rect 25632 4980 25640 4988
rect 25664 4980 25672 4988
rect 25888 4980 25896 4988
rect 26848 4980 26856 4988
rect 28112 4980 28120 4988
rect 28288 4980 28296 4988
rect 28400 4980 28408 4988
rect 34176 4977 34184 4985
rect 34240 4977 34248 4985
rect 34544 4977 34552 4985
rect 34752 4977 34760 4985
rect 36192 4977 36200 4985
rect 36240 4977 36248 4985
rect 39392 4977 39400 4985
rect 39648 4977 39656 4985
rect 40096 4977 40104 4985
rect 40304 4977 40312 4985
rect 27488 4960 27496 4968
rect 27504 4960 27512 4968
rect 27696 4960 27704 4968
rect 29632 4957 29640 4965
rect 30048 4957 30056 4965
rect 30528 4957 30536 4965
rect 30608 4957 30616 4965
rect 31168 4957 31176 4965
rect 31824 4957 31832 4965
rect 32048 4957 32056 4965
rect 32160 4957 32168 4965
rect 32784 4957 32792 4965
rect 32960 4957 32968 4965
rect 33952 4957 33960 4965
rect 34048 4957 34056 4965
rect 35040 4957 35048 4965
rect 35408 4957 35416 4965
rect 35456 4957 35464 4965
rect 36464 4957 36472 4965
rect 36624 4957 36632 4965
rect 37664 4957 37672 4965
rect 37840 4957 37848 4965
rect 37920 4957 37928 4965
rect 38448 4957 38456 4965
rect 38800 4957 38808 4965
rect 39408 4957 39416 4965
rect 39696 4957 39704 4965
rect 39712 4957 39720 4965
rect 22400 4948 22404 4953
rect 18656 4940 18664 4948
rect 20336 4940 20344 4948
rect 20896 4940 20904 4948
rect 20912 4940 20920 4948
rect 23456 4940 23464 4948
rect 23888 4940 23896 4948
rect 24176 4940 24184 4948
rect 24576 4940 24584 4948
rect 24592 4940 24600 4948
rect 24800 4940 24808 4948
rect 25856 4940 25864 4948
rect 27904 4940 27912 4948
rect 33856 4937 33864 4945
rect 18704 4920 18712 4928
rect 19456 4920 19464 4928
rect 20512 4920 20520 4928
rect 20800 4920 20808 4928
rect 27136 4920 27144 4928
rect 40320 4917 40328 4925
rect 18688 4900 18696 4908
rect 25232 4900 25240 4908
rect 25440 4900 25448 4908
rect 25456 4900 25464 4908
rect 38880 4897 38888 4905
rect 29548 4867 29552 4875
rect 29556 4867 29560 4875
rect 29580 4867 29584 4875
rect 29588 4867 29600 4875
rect 29604 4867 29616 4875
rect 29620 4867 29624 4875
rect 29672 4867 29676 4875
rect 29680 4867 29692 4875
rect 29696 4867 29708 4875
rect 29712 4867 29716 4875
rect 29736 4867 29740 4875
rect 29744 4867 29748 4875
rect 29764 4867 29768 4875
rect 29772 4867 29784 4875
rect 29788 4867 29800 4875
rect 29804 4867 29808 4875
rect 29904 4867 29908 4875
rect 29912 4867 29916 4875
rect 29936 4867 29940 4875
rect 29944 4867 29948 4875
rect 29960 4867 29972 4875
rect 29976 4867 29980 4875
rect 30000 4867 30004 4875
rect 30008 4867 30020 4875
rect 30028 4867 30044 4875
rect 30052 4867 30076 4875
rect 30092 4867 30096 4875
rect 30100 4867 30112 4875
rect 30120 4867 30136 4875
rect 30144 4867 30168 4875
rect 30184 4867 30200 4875
rect 30208 4867 30232 4875
rect 30248 4867 30296 4875
rect 30312 4867 30336 4875
rect 30344 4867 30360 4875
rect 30376 4867 30392 4875
rect 30408 4867 30424 4875
rect 30432 4867 30456 4875
rect 30472 4867 30520 4875
rect 30536 4867 30552 4875
rect 30568 4867 30572 4875
rect 30576 4867 30588 4875
rect 30600 4867 30604 4875
rect 30608 4867 30612 4875
rect 30632 4867 30636 4875
rect 30640 4867 30644 4875
rect 30740 4867 30744 4875
rect 30748 4867 30752 4875
rect 30764 4867 30776 4875
rect 30780 4867 30784 4875
rect 30832 4867 30836 4875
rect 30840 4867 30844 4875
rect 30856 4867 30868 4875
rect 30872 4867 30884 4875
rect 30896 4867 30900 4875
rect 30904 4867 30908 4875
rect 30928 4867 30932 4875
rect 30936 4867 30940 4875
rect 31036 4867 31040 4875
rect 31044 4867 31048 4875
rect 31060 4867 31072 4875
rect 31076 4867 31080 4875
rect 31128 4867 31132 4875
rect 31136 4867 31140 4875
rect 31348 4867 31352 4875
rect 31356 4867 31360 4875
rect 31380 4867 31384 4875
rect 31388 4867 31392 4875
rect 31404 4867 31416 4875
rect 31420 4867 31432 4875
rect 31440 4867 31456 4875
rect 31472 4867 31476 4875
rect 31480 4867 31484 4875
rect 31496 4867 31508 4875
rect 31512 4867 31524 4875
rect 31536 4867 31540 4875
rect 31544 4867 31548 4875
rect 31564 4867 31568 4875
rect 31572 4867 31576 4875
rect 31588 4867 31600 4875
rect 31604 4867 31616 4875
rect 31628 4867 31632 4875
rect 31636 4867 31640 4875
rect 31656 4867 31660 4875
rect 31664 4867 31668 4875
rect 31680 4867 31692 4875
rect 31696 4867 31708 4875
rect 31720 4867 31724 4875
rect 31728 4867 31732 4875
rect 31748 4867 31764 4875
rect 31772 4867 31784 4875
rect 31788 4867 31800 4875
rect 31808 4867 31824 4875
rect 31840 4867 31856 4875
rect 31864 4867 31876 4875
rect 31880 4867 31892 4875
rect 31904 4867 31908 4875
rect 31912 4867 31916 4875
rect 31928 4867 31940 4875
rect 31944 4867 31956 4875
rect 31968 4867 31972 4875
rect 31976 4867 31980 4875
rect 32000 4867 32004 4875
rect 32008 4867 32012 4875
rect 32124 4867 32128 4875
rect 32132 4867 32136 4875
rect 32232 4867 32236 4875
rect 32240 4867 32244 4875
rect 32340 4867 32344 4875
rect 32348 4867 32352 4875
rect 32400 4867 32404 4875
rect 32408 4867 32412 4875
rect 32540 4867 32544 4875
rect 32548 4867 32552 4875
rect 32564 4867 32576 4875
rect 32580 4867 32584 4875
rect 32604 4867 32608 4875
rect 32612 4867 32616 4875
rect 32632 4867 32648 4875
rect 32656 4867 32688 4875
rect 32696 4867 32712 4875
rect 32728 4867 32740 4875
rect 32748 4867 32780 4875
rect 32788 4867 32800 4875
rect 32820 4867 32832 4875
rect 32844 4867 32848 4875
rect 32852 4867 32864 4875
rect 32976 4867 32988 4875
rect 33804 4867 33808 4875
rect 33812 4867 33824 4875
rect 33828 4867 33832 4875
rect 33844 4867 33856 4875
rect 33896 4867 33900 4875
rect 33904 4867 33916 4875
rect 33920 4867 33924 4875
rect 33936 4867 33948 4875
rect 33968 4867 33980 4875
rect 33996 4867 34020 4875
rect 34028 4867 34044 4875
rect 34052 4867 34076 4875
rect 34092 4867 34096 4875
rect 34100 4867 34112 4875
rect 34124 4867 34128 4875
rect 34132 4867 34136 4875
rect 34156 4867 34160 4875
rect 34164 4867 34176 4875
rect 34188 4867 34192 4875
rect 34196 4867 34200 4875
rect 34212 4867 34224 4875
rect 34228 4867 34240 4875
rect 34252 4867 34256 4875
rect 34260 4867 34264 4875
rect 34284 4867 34288 4875
rect 34292 4867 34296 4875
rect 34316 4867 34320 4875
rect 34324 4867 34328 4875
rect 34348 4867 34352 4875
rect 34356 4867 34360 4875
rect 34372 4867 34384 4875
rect 34388 4867 34400 4875
rect 34408 4867 34424 4875
rect 34440 4867 34488 4875
rect 34504 4867 34516 4875
rect 34536 4867 34548 4875
rect 34560 4867 34564 4875
rect 34568 4867 34580 4875
rect 34788 4867 34800 4875
rect 34804 4867 34808 4875
rect 34820 4867 34832 4875
rect 34844 4867 34848 4875
rect 34852 4867 34864 4875
rect 34884 4867 34896 4875
rect 34908 4867 34912 4875
rect 34916 4867 34928 4875
rect 34948 4867 34960 4875
rect 34964 4867 34968 4875
rect 35072 4867 35084 4875
rect 35088 4867 35092 4875
rect 35256 4867 35268 4875
rect 35272 4867 35276 4875
rect 35348 4867 35360 4875
rect 35364 4867 35368 4875
rect 35440 4867 35452 4875
rect 35456 4867 35460 4875
rect 35524 4867 35528 4875
rect 35532 4867 35544 4875
rect 35564 4867 35576 4875
rect 35580 4867 35592 4875
rect 35596 4867 35608 4875
rect 35624 4867 35640 4875
rect 35648 4867 35680 4875
rect 35688 4867 35704 4875
rect 35720 4867 35724 4875
rect 35728 4867 35732 4875
rect 35752 4867 35756 4875
rect 35760 4867 35772 4875
rect 35784 4867 35788 4875
rect 35792 4867 35796 4875
rect 35808 4867 35820 4875
rect 35824 4867 35828 4875
rect 35924 4867 35928 4875
rect 35932 4867 35936 4875
rect 35948 4867 35960 4875
rect 35964 4867 35976 4875
rect 35984 4867 36000 4875
rect 36016 4867 36020 4875
rect 36024 4867 36028 4875
rect 36040 4867 36052 4875
rect 36056 4867 36068 4875
rect 36080 4867 36084 4875
rect 36088 4867 36092 4875
rect 36104 4867 36116 4875
rect 36120 4867 36124 4875
rect 36140 4867 36144 4875
rect 36148 4867 36160 4875
rect 36172 4867 36176 4875
rect 36180 4867 36184 4875
rect 36196 4867 36208 4875
rect 36212 4867 36216 4875
rect 36232 4867 36248 4875
rect 36264 4867 36280 4875
rect 36288 4867 36320 4875
rect 36328 4867 36340 4875
rect 36360 4867 36372 4875
rect 36380 4867 36412 4875
rect 36420 4867 36432 4875
rect 36448 4867 36464 4875
rect 36472 4867 36504 4875
rect 36512 4867 36528 4875
rect 36540 4867 36556 4875
rect 36564 4867 36596 4875
rect 36604 4867 36620 4875
rect 36636 4867 36648 4875
rect 36656 4867 36688 4875
rect 36696 4867 36708 4875
rect 36728 4867 36740 4875
rect 36744 4867 36756 4875
rect 36760 4867 36772 4875
rect 36820 4867 36832 4875
rect 36836 4867 36848 4875
rect 36852 4867 36864 4875
rect 36880 4867 36896 4875
rect 36912 4867 36924 4875
rect 36928 4867 36940 4875
rect 36944 4867 36956 4875
rect 37004 4867 37016 4875
rect 37020 4867 37032 4875
rect 37036 4867 37048 4875
rect 37068 4867 37080 4875
rect 37096 4867 37108 4875
rect 37112 4867 37124 4875
rect 37128 4867 37140 4875
rect 37212 4867 37216 4875
rect 37220 4867 37232 4875
rect 37252 4867 37264 4875
rect 37268 4867 37272 4875
rect 37344 4867 37356 4875
rect 37360 4867 37364 4875
rect 37376 4867 37388 4875
rect 37408 4867 37420 4875
rect 37436 4867 37484 4875
rect 37500 4867 37516 4875
rect 37532 4867 37548 4875
rect 37564 4867 37580 4875
rect 37600 4867 37644 4875
rect 37660 4867 37664 4875
rect 37668 4867 37672 4875
rect 37692 4867 37696 4875
rect 37700 4867 37712 4875
rect 37724 4867 37728 4875
rect 37732 4867 37736 4875
rect 37864 4867 37868 4875
rect 37872 4867 37876 4875
rect 37888 4867 37900 4875
rect 37904 4867 37908 4875
rect 37956 4867 37960 4875
rect 37964 4867 37968 4875
rect 37980 4867 37992 4875
rect 37996 4867 38000 4875
rect 38020 4867 38024 4875
rect 38028 4867 38032 4875
rect 38044 4867 38056 4875
rect 38060 4867 38064 4875
rect 38080 4867 38104 4875
rect 38112 4867 38128 4875
rect 38136 4867 38168 4875
rect 38176 4867 38188 4875
rect 38204 4867 38220 4875
rect 38228 4867 38260 4875
rect 38268 4867 38284 4875
rect 38300 4867 38304 4875
rect 38308 4867 38312 4875
rect 38332 4867 38336 4875
rect 38340 4867 38352 4875
rect 38364 4867 38368 4875
rect 38372 4867 38376 4875
rect 38388 4867 38400 4875
rect 38404 4867 38408 4875
rect 38424 4867 38428 4875
rect 38432 4867 38444 4875
rect 38456 4867 38460 4875
rect 38464 4867 38468 4875
rect 38480 4867 38492 4875
rect 38496 4867 38500 4875
rect 38516 4867 38520 4875
rect 38524 4867 38536 4875
rect 38548 4867 38552 4875
rect 38556 4867 38560 4875
rect 38572 4867 38584 4875
rect 38588 4867 38600 4875
rect 38608 4867 38624 4875
rect 38640 4867 38656 4875
rect 38664 4867 38676 4875
rect 38680 4867 38692 4875
rect 38704 4867 38708 4875
rect 38712 4867 38716 4875
rect 38732 4867 38736 4875
rect 38740 4867 38744 4875
rect 38756 4867 38768 4875
rect 38772 4867 38784 4875
rect 38796 4867 38800 4875
rect 38804 4867 38808 4875
rect 38824 4867 38840 4875
rect 38848 4867 38860 4875
rect 38864 4867 38876 4875
rect 38888 4867 38892 4875
rect 38896 4867 38900 4875
rect 38916 4867 38932 4875
rect 38940 4867 38964 4875
rect 38980 4867 38992 4875
rect 39012 4867 39024 4875
rect 39028 4867 39040 4875
rect 39044 4867 39056 4875
rect 39128 4867 39132 4875
rect 39136 4867 39148 4875
rect 39168 4867 39180 4875
rect 39184 4867 39188 4875
rect 39292 4867 39304 4875
rect 39308 4867 39312 4875
rect 39324 4867 39336 4875
rect 39348 4867 39352 4875
rect 39356 4867 39368 4875
rect 39372 4867 39376 4875
rect 39440 4867 39444 4875
rect 39448 4867 39460 4875
rect 39464 4867 39468 4875
rect 39532 4867 39536 4875
rect 39540 4867 39552 4875
rect 39556 4867 39560 4875
rect 39624 4867 39628 4875
rect 39632 4867 39644 4875
rect 39648 4867 39652 4875
rect 39692 4867 39704 4875
rect 39716 4867 39720 4875
rect 39724 4867 39736 4875
rect 39740 4867 39744 4875
rect 39808 4867 39812 4875
rect 39816 4867 39828 4875
rect 39832 4867 39836 4875
rect 39848 4867 39860 4875
rect 39872 4867 39876 4875
rect 39880 4867 39892 4875
rect 40068 4867 40080 4875
rect 40084 4867 40088 4875
rect 40100 4867 40112 4875
rect 40124 4867 40128 4875
rect 40132 4867 40144 4875
rect 40164 4867 40176 4875
rect 40196 4867 40208 4875
rect 40228 4867 40240 4875
rect 40244 4867 40248 4875
rect 40260 4867 40272 4875
rect 40284 4867 40288 4875
rect 40292 4867 40304 4875
rect 40324 4867 40336 4875
rect 40348 4867 40352 4875
rect 40356 4867 40368 4875
rect 40472 4867 40476 4875
rect 40480 4867 40492 4875
rect 40604 4867 40616 4875
rect 40620 4867 40632 4875
rect 40636 4867 40648 4875
rect 40668 4867 40680 4875
rect 40696 4867 40720 4875
rect 40728 4867 40744 4875
rect 40760 4867 40776 4875
rect 40784 4867 40796 4875
rect 18472 4848 18474 4860
rect 21668 4850 21670 4858
rect 21676 4850 21678 4858
rect 23622 4850 23626 4858
rect 23630 4850 23634 4858
rect 23944 4850 23948 4858
rect 23952 4850 23956 4858
rect 24158 4850 24162 4858
rect 24166 4850 24170 4858
rect 21360 4840 21368 4848
rect 29440 4837 29448 4845
rect 31216 4837 31224 4845
rect 35728 4817 35736 4825
rect 35888 4817 35896 4825
rect 36016 4817 36024 4825
rect 36256 4817 36264 4825
rect 36720 4817 36728 4825
rect 39872 4817 39880 4825
rect 40080 4817 40088 4825
rect 19472 4800 19480 4808
rect 26672 4800 26680 4808
rect 39104 4797 39112 4805
rect 39280 4797 39288 4805
rect 21200 4780 21208 4788
rect 27520 4780 27528 4788
rect 29536 4777 29544 4785
rect 29840 4777 29848 4785
rect 29920 4777 29928 4785
rect 30096 4777 30104 4785
rect 30144 4777 30152 4785
rect 30496 4777 30504 4785
rect 30912 4777 30920 4785
rect 31104 4777 31112 4785
rect 32720 4777 32728 4785
rect 33056 4777 33064 4785
rect 33248 4777 33256 4785
rect 33424 4777 33432 4785
rect 33840 4777 33848 4785
rect 34528 4777 34536 4785
rect 34848 4777 34856 4785
rect 37056 4777 37064 4785
rect 38304 4777 38312 4785
rect 39072 4777 39080 4785
rect 39152 4777 39160 4785
rect 39168 4777 39176 4785
rect 39920 4777 39928 4785
rect 39936 4777 39944 4785
rect 40496 4777 40504 4785
rect 40752 4777 40760 4785
rect 18640 4760 18648 4768
rect 20112 4760 20120 4768
rect 22208 4760 22216 4768
rect 22432 4760 22440 4768
rect 23408 4760 23416 4768
rect 23680 4760 23688 4768
rect 25824 4760 25832 4768
rect 26256 4760 26264 4768
rect 26880 4760 26888 4768
rect 27728 4760 27736 4768
rect 31824 4757 31832 4765
rect 32432 4757 32440 4765
rect 33936 4757 33944 4765
rect 34624 4757 34632 4765
rect 37376 4757 37384 4765
rect 19888 4740 19896 4748
rect 27072 4740 27080 4748
rect 29664 4737 29672 4745
rect 29984 4737 29992 4745
rect 31072 4737 31080 4745
rect 31520 4737 31528 4745
rect 31840 4737 31848 4745
rect 32192 4737 32200 4745
rect 32288 4737 32296 4745
rect 33824 4737 33832 4745
rect 34544 4737 34552 4745
rect 35536 4737 35544 4745
rect 35552 4737 35560 4745
rect 35568 4737 35576 4745
rect 36576 4737 36584 4745
rect 36816 4737 36824 4745
rect 37552 4737 37560 4745
rect 38368 4737 38376 4745
rect 38448 4737 38456 4745
rect 39600 4737 39608 4745
rect 40736 4737 40744 4745
rect 18832 4720 18840 4728
rect 19520 4720 19528 4728
rect 20112 4720 20120 4728
rect 23056 4720 23064 4728
rect 23408 4720 23416 4728
rect 23600 4720 23608 4728
rect 24128 4720 24136 4728
rect 24768 4720 24776 4728
rect 25616 4720 25624 4728
rect 26480 4720 26488 4728
rect 27104 4720 27112 4728
rect 27312 4720 27320 4728
rect 27552 4720 27560 4728
rect 27568 4720 27576 4728
rect 27712 4720 27720 4728
rect 27744 4720 27752 4728
rect 30784 4717 30792 4725
rect 30864 4717 30872 4725
rect 31200 4717 31208 4725
rect 31232 4717 31240 4725
rect 32064 4717 32072 4725
rect 33760 4717 33768 4725
rect 34576 4717 34584 4725
rect 34848 4717 34856 4725
rect 36544 4717 36552 4725
rect 37696 4717 37704 4725
rect 37776 4717 37784 4725
rect 38144 4717 38152 4725
rect 39264 4717 39272 4725
rect 39312 4717 39320 4725
rect 39856 4717 39864 4725
rect 40000 4717 40008 4725
rect 40016 4717 40024 4725
rect 20176 4700 20184 4708
rect 20320 4700 20328 4708
rect 21728 4700 21736 4708
rect 21936 4700 21944 4708
rect 22624 4700 22632 4708
rect 23744 4700 23752 4708
rect 24288 4700 24296 4708
rect 25120 4700 25128 4708
rect 31200 4697 31208 4705
rect 32864 4697 32872 4705
rect 35776 4697 35784 4705
rect 35872 4697 35880 4705
rect 36000 4697 36008 4705
rect 36960 4697 36968 4705
rect 39760 4697 39768 4705
rect 21376 4680 21384 4688
rect 23232 4680 23240 4688
rect 25552 4680 25560 4688
rect 19968 4660 19976 4668
rect 24064 4660 24072 4668
rect 26400 4660 26408 4668
rect 27888 4660 27896 4668
rect 29548 4667 29552 4675
rect 29556 4667 29560 4675
rect 29580 4667 29584 4675
rect 29588 4667 29600 4675
rect 29604 4667 29616 4675
rect 29620 4667 29624 4675
rect 29640 4667 29644 4675
rect 29648 4667 29652 4675
rect 29672 4667 29676 4675
rect 29680 4667 29692 4675
rect 29696 4667 29708 4675
rect 29712 4667 29716 4675
rect 29736 4667 29740 4675
rect 29744 4667 29748 4675
rect 29812 4667 29816 4675
rect 29820 4667 29824 4675
rect 29844 4667 29848 4675
rect 29852 4667 29856 4675
rect 29868 4667 29880 4675
rect 29884 4667 29888 4675
rect 29904 4667 29928 4675
rect 29936 4667 29952 4675
rect 29960 4667 29984 4675
rect 30000 4667 30016 4675
rect 30032 4667 30044 4675
rect 30056 4667 30060 4675
rect 30064 4667 30076 4675
rect 30080 4667 30084 4675
rect 30096 4667 30108 4675
rect 30124 4667 30136 4675
rect 30148 4667 30152 4675
rect 30156 4667 30168 4675
rect 30172 4667 30176 4675
rect 30188 4667 30200 4675
rect 30212 4667 30216 4675
rect 30220 4667 30232 4675
rect 30236 4667 30240 4675
rect 30252 4667 30264 4675
rect 30276 4667 30280 4675
rect 30284 4667 30296 4675
rect 30312 4667 30336 4675
rect 30344 4667 30360 4675
rect 30376 4667 30392 4675
rect 30408 4667 30424 4675
rect 30432 4667 30456 4675
rect 30472 4667 30520 4675
rect 30536 4667 30540 4675
rect 30544 4667 30548 4675
rect 30568 4667 30572 4675
rect 30576 4667 30588 4675
rect 30600 4667 30604 4675
rect 30608 4667 30612 4675
rect 30708 4667 30712 4675
rect 30716 4667 30728 4675
rect 30740 4667 30744 4675
rect 30748 4667 30752 4675
rect 30764 4667 30776 4675
rect 30780 4667 30784 4675
rect 30800 4667 30804 4675
rect 30808 4667 30820 4675
rect 30832 4667 30836 4675
rect 30840 4667 30844 4675
rect 30856 4667 30868 4675
rect 30872 4667 30884 4675
rect 30892 4667 30908 4675
rect 30924 4667 30940 4675
rect 30948 4667 30960 4675
rect 30964 4667 30976 4675
rect 30988 4667 30992 4675
rect 30996 4667 31000 4675
rect 31012 4667 31024 4675
rect 31028 4667 31032 4675
rect 31128 4667 31132 4675
rect 31136 4667 31140 4675
rect 31152 4667 31164 4675
rect 31168 4667 31180 4675
rect 31192 4667 31196 4675
rect 31200 4667 31204 4675
rect 31348 4667 31352 4675
rect 31356 4667 31360 4675
rect 31440 4667 31444 4675
rect 31448 4667 31452 4675
rect 31564 4667 31568 4675
rect 31572 4667 31576 4675
rect 31588 4667 31600 4675
rect 31604 4667 31608 4675
rect 31628 4667 31632 4675
rect 31636 4667 31640 4675
rect 31656 4667 31704 4675
rect 31720 4667 31744 4675
rect 31752 4667 31764 4675
rect 31776 4667 31780 4675
rect 31784 4667 31796 4675
rect 32036 4667 32048 4675
rect 32052 4667 32056 4675
rect 32068 4667 32080 4675
rect 32088 4667 32112 4675
rect 32128 4667 32140 4675
rect 32144 4667 32148 4675
rect 32160 4667 32172 4675
rect 32184 4667 32188 4675
rect 32192 4667 32204 4675
rect 32208 4667 32212 4675
rect 32224 4667 32236 4675
rect 32348 4667 32360 4675
rect 32364 4667 32376 4675
rect 32380 4667 32392 4675
rect 32408 4667 32424 4675
rect 32432 4667 32464 4675
rect 32472 4667 32488 4675
rect 32496 4667 32528 4675
rect 32536 4667 32552 4675
rect 32568 4667 32580 4675
rect 32592 4667 32596 4675
rect 32600 4667 32612 4675
rect 32724 4667 32736 4675
rect 32816 4667 32828 4675
rect 32848 4667 32860 4675
rect 32864 4667 32868 4675
rect 32880 4667 32892 4675
rect 32912 4667 32924 4675
rect 32928 4667 32940 4675
rect 32944 4667 32956 4675
rect 32972 4667 32984 4675
rect 33004 4667 33016 4675
rect 33020 4667 33032 4675
rect 33036 4667 33048 4675
rect 33068 4667 33080 4675
rect 33184 4667 33188 4675
rect 33192 4667 33204 4675
rect 33208 4667 33212 4675
rect 33276 4667 33280 4675
rect 33284 4667 33296 4675
rect 33300 4667 33304 4675
rect 33316 4667 33328 4675
rect 33348 4667 33360 4675
rect 33376 4667 33400 4675
rect 33408 4667 33424 4675
rect 33432 4667 33456 4675
rect 33468 4667 33492 4675
rect 33500 4667 33516 4675
rect 33524 4667 33548 4675
rect 33564 4667 33568 4675
rect 33572 4667 33584 4675
rect 33596 4667 33600 4675
rect 33604 4667 33608 4675
rect 33628 4667 33632 4675
rect 33636 4667 33640 4675
rect 33660 4667 33664 4675
rect 33668 4667 33672 4675
rect 33684 4667 33696 4675
rect 33700 4667 33704 4675
rect 33720 4667 33744 4675
rect 33752 4667 33768 4675
rect 33776 4667 33808 4675
rect 33816 4667 33828 4675
rect 33848 4667 33860 4675
rect 33868 4667 33900 4675
rect 33908 4667 33924 4675
rect 33940 4667 33952 4675
rect 33964 4667 33968 4675
rect 33972 4667 33984 4675
rect 34004 4667 34016 4675
rect 34128 4667 34140 4675
rect 34144 4667 34148 4675
rect 34160 4667 34172 4675
rect 34192 4667 34204 4675
rect 34212 4667 34244 4675
rect 34252 4667 34268 4675
rect 34284 4667 34288 4675
rect 34292 4667 34296 4675
rect 34316 4667 34320 4675
rect 34324 4667 34336 4675
rect 34348 4667 34352 4675
rect 34356 4667 34360 4675
rect 34372 4667 34384 4675
rect 34388 4667 34392 4675
rect 34408 4667 34412 4675
rect 34416 4667 34428 4675
rect 34440 4667 34444 4675
rect 34448 4667 34452 4675
rect 34464 4667 34476 4675
rect 34480 4667 34492 4675
rect 34500 4667 34516 4675
rect 34532 4667 34548 4675
rect 34556 4667 34568 4675
rect 34572 4667 34584 4675
rect 34592 4667 34608 4675
rect 34624 4667 34640 4675
rect 34648 4667 34660 4675
rect 34664 4667 34676 4675
rect 34688 4667 34692 4675
rect 34696 4667 34700 4675
rect 34712 4667 34724 4675
rect 34728 4667 34732 4675
rect 34752 4667 34756 4675
rect 34760 4667 34764 4675
rect 34780 4667 34796 4675
rect 34804 4667 34836 4675
rect 34844 4667 34860 4675
rect 34876 4667 34880 4675
rect 34884 4667 34888 4675
rect 34908 4667 34912 4675
rect 34916 4667 34928 4675
rect 34940 4667 34944 4675
rect 34948 4667 34952 4675
rect 34964 4667 34976 4675
rect 34980 4667 34992 4675
rect 35004 4667 35008 4675
rect 35012 4667 35016 4675
rect 35028 4667 35040 4675
rect 35044 4667 35056 4675
rect 35068 4667 35072 4675
rect 35076 4667 35080 4675
rect 35096 4667 35112 4675
rect 35120 4667 35144 4675
rect 35160 4667 35172 4675
rect 35192 4667 35204 4675
rect 35208 4667 35220 4675
rect 35224 4667 35236 4675
rect 35252 4667 35268 4675
rect 35284 4667 35296 4675
rect 35300 4667 35312 4675
rect 35316 4667 35328 4675
rect 35348 4667 35360 4675
rect 35464 4667 35468 4675
rect 35472 4667 35484 4675
rect 35488 4667 35492 4675
rect 35504 4667 35516 4675
rect 35524 4667 35548 4675
rect 35564 4667 35612 4675
rect 35628 4667 35632 4675
rect 35636 4667 35640 4675
rect 35660 4667 35664 4675
rect 35668 4667 35680 4675
rect 35692 4667 35696 4675
rect 35700 4667 35704 4675
rect 35832 4667 35836 4675
rect 35840 4667 35844 4675
rect 35856 4667 35868 4675
rect 35872 4667 35884 4675
rect 35896 4667 35900 4675
rect 35904 4667 35908 4675
rect 35924 4667 35940 4675
rect 35948 4667 35972 4675
rect 35988 4667 36000 4675
rect 36020 4667 36032 4675
rect 36036 4667 36048 4675
rect 36052 4667 36064 4675
rect 36084 4667 36096 4675
rect 36100 4667 36112 4675
rect 36116 4667 36128 4675
rect 36240 4667 36252 4675
rect 36264 4667 36268 4675
rect 36272 4667 36284 4675
rect 36288 4667 36292 4675
rect 36304 4667 36316 4675
rect 36332 4667 36348 4675
rect 36364 4667 36388 4675
rect 36396 4667 36412 4675
rect 36420 4667 36432 4675
rect 36436 4667 36440 4675
rect 36456 4667 36480 4675
rect 36488 4667 36504 4675
rect 36512 4667 36536 4675
rect 36552 4667 36556 4675
rect 36560 4667 36572 4675
rect 36576 4667 36588 4675
rect 36592 4667 36596 4675
rect 36616 4667 36620 4675
rect 36624 4667 36628 4675
rect 36692 4667 36696 4675
rect 36700 4667 36704 4675
rect 36724 4667 36728 4675
rect 36732 4667 36744 4675
rect 36748 4667 36760 4675
rect 36764 4667 36768 4675
rect 36784 4667 36800 4675
rect 36816 4667 36820 4675
rect 36824 4667 36836 4675
rect 36840 4667 36852 4675
rect 36856 4667 36860 4675
rect 36880 4667 36884 4675
rect 36888 4667 36892 4675
rect 36908 4667 36924 4675
rect 36932 4667 36956 4675
rect 36972 4667 36984 4675
rect 36988 4667 36992 4675
rect 37004 4667 37016 4675
rect 37028 4667 37032 4675
rect 37036 4667 37048 4675
rect 37052 4667 37056 4675
rect 37068 4667 37080 4675
rect 37160 4667 37172 4675
rect 37192 4667 37204 4675
rect 37208 4667 37220 4675
rect 37224 4667 37236 4675
rect 37256 4667 37268 4675
rect 37276 4667 37308 4675
rect 37316 4667 37332 4675
rect 37348 4667 37360 4675
rect 37372 4667 37376 4675
rect 37380 4667 37392 4675
rect 37412 4667 37424 4675
rect 37436 4667 37440 4675
rect 37444 4667 37456 4675
rect 37460 4667 37464 4675
rect 37476 4667 37488 4675
rect 37600 4667 37612 4675
rect 37616 4667 37628 4675
rect 37632 4667 37644 4675
rect 37664 4667 37676 4675
rect 37692 4667 37716 4675
rect 37724 4667 37740 4675
rect 37756 4667 37760 4675
rect 37764 4667 37768 4675
rect 37780 4667 37792 4675
rect 37796 4667 37808 4675
rect 37820 4667 37824 4675
rect 37828 4667 37832 4675
rect 37844 4667 37856 4675
rect 37860 4667 37864 4675
rect 37912 4667 37916 4675
rect 37920 4667 37924 4675
rect 37936 4667 37948 4675
rect 37952 4667 37956 4675
rect 38020 4667 38024 4675
rect 38028 4667 38032 4675
rect 38052 4667 38056 4675
rect 38060 4667 38064 4675
rect 38076 4667 38088 4675
rect 38092 4667 38104 4675
rect 38116 4667 38120 4675
rect 38124 4667 38128 4675
rect 38148 4667 38152 4675
rect 38156 4667 38168 4675
rect 38180 4667 38184 4675
rect 38188 4667 38192 4675
rect 38272 4667 38276 4675
rect 38280 4667 38284 4675
rect 38396 4667 38400 4675
rect 38404 4667 38408 4675
rect 38504 4667 38508 4675
rect 38512 4667 38516 4675
rect 38528 4667 38540 4675
rect 38544 4667 38548 4675
rect 38568 4667 38572 4675
rect 38576 4667 38588 4675
rect 38592 4667 38604 4675
rect 38608 4667 38612 4675
rect 38632 4667 38636 4675
rect 38640 4667 38644 4675
rect 38660 4667 38676 4675
rect 38684 4667 38708 4675
rect 38724 4667 38736 4675
rect 38740 4667 38744 4675
rect 38756 4667 38768 4675
rect 38780 4667 38784 4675
rect 38788 4667 38800 4675
rect 38816 4667 38840 4675
rect 38848 4667 38860 4675
rect 38872 4667 38876 4675
rect 38880 4667 38892 4675
rect 38908 4667 38932 4675
rect 38940 4667 38956 4675
rect 38972 4667 38976 4675
rect 38980 4667 38984 4675
rect 39004 4667 39008 4675
rect 39012 4667 39024 4675
rect 39028 4667 39040 4675
rect 39044 4667 39048 4675
rect 39068 4667 39072 4675
rect 39076 4667 39088 4675
rect 39092 4667 39104 4675
rect 39108 4667 39112 4675
rect 39128 4667 39144 4675
rect 39160 4667 39164 4675
rect 39168 4667 39180 4675
rect 39184 4667 39196 4675
rect 39200 4667 39204 4675
rect 39224 4667 39228 4675
rect 39232 4667 39236 4675
rect 39380 4667 39384 4675
rect 39388 4667 39392 4675
rect 39412 4667 39416 4675
rect 39420 4667 39424 4675
rect 39436 4667 39448 4675
rect 39452 4667 39456 4675
rect 39472 4667 39496 4675
rect 39504 4667 39520 4675
rect 39528 4667 39552 4675
rect 39568 4667 39580 4675
rect 39600 4667 39612 4675
rect 39624 4667 39628 4675
rect 39632 4667 39644 4675
rect 39648 4667 39652 4675
rect 39716 4667 39720 4675
rect 39724 4667 39736 4675
rect 39740 4667 39744 4675
rect 39784 4667 39796 4675
rect 39808 4667 39812 4675
rect 39816 4667 39828 4675
rect 39832 4667 39836 4675
rect 39848 4667 39860 4675
rect 39872 4667 39876 4675
rect 39880 4667 39892 4675
rect 39908 4667 39920 4675
rect 39924 4667 39928 4675
rect 39940 4667 39952 4675
rect 39964 4667 39968 4675
rect 39972 4667 39984 4675
rect 40000 4667 40024 4675
rect 40032 4667 40048 4675
rect 40064 4667 40080 4675
rect 40096 4667 40100 4675
rect 40104 4667 40116 4675
rect 40120 4667 40132 4675
rect 40136 4667 40140 4675
rect 40160 4667 40164 4675
rect 40168 4667 40172 4675
rect 40268 4667 40272 4675
rect 40276 4667 40288 4675
rect 40292 4667 40304 4675
rect 40308 4667 40312 4675
rect 40332 4667 40336 4675
rect 40340 4667 40352 4675
rect 40364 4667 40368 4675
rect 40372 4667 40376 4675
rect 40472 4667 40476 4675
rect 40480 4667 40484 4675
rect 40504 4667 40508 4675
rect 40512 4667 40516 4675
rect 40596 4667 40600 4675
rect 40604 4667 40608 4675
rect 40688 4667 40692 4675
rect 40696 4667 40700 4675
rect 40712 4667 40724 4675
rect 40728 4667 40732 4675
rect 40752 4667 40756 4675
rect 40760 4667 40764 4675
rect 40780 4667 40800 4675
rect 18740 4652 18742 4660
rect 18938 4652 18940 4660
rect 20634 4652 20636 4660
rect 21634 4656 21636 4660
rect 21640 4652 21642 4656
rect 22464 4650 22468 4658
rect 22554 4650 22562 4658
rect 22886 4656 22888 4660
rect 23100 4656 23102 4660
rect 23314 4656 23316 4660
rect 22892 4652 22894 4656
rect 23106 4652 23108 4656
rect 23320 4652 23322 4656
rect 23480 4650 23488 4658
rect 23630 4650 23636 4658
rect 24336 4650 24344 4658
rect 24486 4650 24492 4658
rect 24550 4650 24558 4658
rect 24700 4650 24706 4658
rect 24786 4650 24790 4658
rect 24876 4650 24884 4658
rect 25080 4656 25082 4660
rect 25224 4656 25226 4660
rect 25086 4652 25088 4656
rect 25230 4652 25232 4656
rect 25428 4650 25432 4658
rect 25518 4650 25526 4658
rect 25722 4656 25724 4660
rect 25936 4656 25938 4660
rect 25728 4652 25730 4656
rect 25942 4652 25944 4656
rect 26070 4650 26074 4658
rect 26160 4650 26168 4658
rect 26284 4650 26288 4658
rect 26374 4650 26382 4658
rect 26578 4656 26580 4660
rect 27418 4656 27420 4660
rect 27632 4656 27634 4660
rect 26584 4652 26586 4656
rect 27424 4652 27426 4656
rect 27638 4652 27640 4656
rect 27766 4650 27770 4658
rect 27856 4650 27864 4658
rect 28060 4656 28062 4660
rect 28274 4656 28276 4660
rect 28488 4656 28490 4660
rect 33568 4657 33576 4665
rect 38032 4657 38040 4665
rect 39712 4657 39720 4665
rect 28066 4652 28068 4656
rect 28280 4652 28282 4656
rect 28494 4652 28496 4656
rect 20112 4640 20120 4648
rect 23680 4640 23688 4648
rect 25120 4640 25128 4648
rect 25760 4640 25768 4648
rect 28112 4640 28120 4648
rect 30064 4637 30072 4645
rect 30784 4637 30792 4645
rect 30960 4637 30968 4645
rect 19472 4620 19480 4628
rect 19680 4620 19688 4628
rect 20352 4620 20360 4628
rect 21568 4620 21576 4628
rect 22608 4620 22616 4628
rect 23248 4620 23256 4628
rect 23904 4620 23912 4628
rect 24128 4620 24136 4628
rect 25136 4620 25144 4628
rect 26224 4620 26232 4628
rect 28656 4620 28664 4628
rect 29600 4617 29608 4625
rect 29744 4617 29752 4625
rect 29872 4617 29880 4625
rect 30336 4617 30344 4625
rect 30448 4617 30456 4625
rect 31056 4617 31064 4625
rect 31120 4617 31128 4625
rect 31424 4617 31432 4625
rect 31552 4617 31560 4625
rect 33024 4617 33032 4625
rect 34240 4617 34248 4625
rect 35008 4617 35016 4625
rect 35168 4617 35176 4625
rect 35536 4617 35544 4625
rect 35680 4617 35688 4625
rect 35824 4617 35832 4625
rect 35872 4617 35880 4625
rect 35984 4617 35992 4625
rect 36112 4617 36120 4625
rect 36192 4617 36200 4625
rect 36400 4617 36408 4625
rect 38464 4617 38472 4625
rect 38640 4617 38648 4625
rect 39040 4617 39048 4625
rect 39344 4617 39352 4625
rect 39392 4617 39400 4625
rect 20928 4600 20936 4608
rect 20944 4600 20952 4608
rect 22176 4600 22184 4608
rect 23008 4600 23016 4608
rect 27264 4600 27272 4608
rect 28176 4600 28184 4608
rect 29600 4597 29608 4605
rect 29744 4597 29752 4605
rect 29968 4597 29976 4605
rect 30832 4597 30840 4605
rect 30928 4597 30936 4605
rect 31680 4597 31688 4605
rect 32304 4597 32312 4605
rect 33088 4597 33096 4605
rect 33136 4597 33144 4605
rect 33584 4597 33592 4605
rect 33856 4597 33864 4605
rect 34928 4597 34936 4605
rect 35664 4597 35672 4605
rect 35968 4597 35976 4605
rect 40192 4597 40200 4605
rect 40688 4597 40696 4605
rect 40768 4597 40776 4605
rect 18512 4580 18520 4588
rect 18816 4580 18824 4588
rect 19728 4580 19736 4588
rect 19856 4580 19864 4588
rect 20176 4580 20184 4588
rect 20736 4580 20744 4588
rect 21728 4580 21736 4588
rect 22032 4580 22040 4588
rect 22160 4580 22168 4588
rect 22768 4580 22776 4588
rect 22992 4580 23000 4588
rect 23200 4580 23208 4588
rect 25632 4580 25640 4588
rect 26192 4580 26200 4588
rect 27328 4580 27336 4588
rect 27360 4580 27368 4588
rect 27488 4580 27496 4588
rect 27968 4580 27976 4588
rect 28192 4580 28200 4588
rect 28528 4580 28536 4588
rect 30000 4577 30008 4585
rect 30400 4577 30408 4585
rect 31088 4577 31096 4585
rect 31760 4577 31768 4585
rect 34416 4577 34424 4585
rect 36576 4577 36584 4585
rect 36864 4577 36872 4585
rect 37104 4577 37112 4585
rect 39264 4577 39272 4585
rect 39408 4577 39416 4585
rect 40336 4577 40344 4585
rect 40544 4577 40552 4585
rect 40688 4577 40696 4585
rect 25328 4560 25336 4568
rect 25536 4560 25544 4568
rect 27296 4560 27304 4568
rect 29568 4557 29576 4565
rect 30544 4557 30552 4565
rect 30640 4557 30648 4565
rect 31232 4557 31240 4565
rect 32000 4557 32008 4565
rect 32112 4557 32120 4565
rect 32528 4557 32536 4565
rect 34480 4557 34488 4565
rect 34880 4557 34888 4565
rect 36768 4557 36776 4565
rect 37312 4557 37320 4565
rect 39216 4557 39224 4565
rect 39872 4557 39880 4565
rect 39968 4557 39976 4565
rect 40144 4557 40152 4565
rect 19040 4548 19044 4553
rect 19666 4548 19670 4553
rect 23010 4548 23014 4553
rect 18496 4540 18504 4548
rect 18832 4540 18840 4548
rect 18864 4540 18872 4548
rect 19088 4540 19096 4548
rect 20160 4540 20168 4548
rect 21200 4540 21208 4548
rect 23216 4540 23224 4548
rect 23504 4540 23512 4548
rect 24352 4540 24360 4548
rect 24960 4540 24968 4548
rect 24976 4540 24984 4548
rect 25616 4540 25624 4548
rect 25792 4540 25800 4548
rect 26480 4540 26488 4548
rect 27312 4540 27320 4548
rect 27712 4540 27720 4548
rect 27888 4540 27896 4548
rect 28384 4540 28392 4548
rect 30272 4537 30280 4545
rect 35936 4537 35944 4545
rect 37296 4537 37304 4545
rect 22592 4520 22600 4528
rect 24720 4520 24728 4528
rect 26416 4520 26424 4528
rect 37600 4517 37608 4525
rect 37744 4517 37752 4525
rect 23872 4500 23880 4508
rect 24912 4500 24920 4508
rect 25552 4500 25560 4508
rect 18640 4460 18648 4468
rect 30060 4467 30072 4475
rect 30076 4467 30088 4475
rect 30092 4467 30104 4475
rect 30120 4467 30132 4475
rect 30152 4467 30164 4475
rect 30168 4467 30180 4475
rect 30184 4467 30196 4475
rect 30212 4467 30228 4475
rect 30236 4467 30268 4475
rect 30276 4467 30292 4475
rect 30304 4467 30320 4475
rect 30328 4467 30360 4475
rect 30368 4467 30384 4475
rect 30400 4467 30404 4475
rect 30408 4467 30412 4475
rect 30432 4467 30436 4475
rect 30440 4467 30452 4475
rect 30472 4467 30484 4475
rect 30488 4467 30492 4475
rect 30504 4467 30516 4475
rect 30532 4467 30548 4475
rect 30564 4467 30604 4475
rect 30616 4467 30632 4475
rect 30648 4467 30696 4475
rect 30712 4467 30724 4475
rect 30740 4467 30788 4475
rect 30804 4467 30816 4475
rect 30836 4467 30848 4475
rect 30860 4467 30864 4475
rect 30868 4467 30880 4475
rect 30992 4467 31004 4475
rect 31008 4467 31020 4475
rect 31024 4467 31036 4475
rect 31056 4467 31068 4475
rect 31084 4467 31108 4475
rect 31116 4467 31132 4475
rect 31148 4467 31152 4475
rect 31156 4467 31160 4475
rect 31172 4467 31184 4475
rect 31188 4467 31200 4475
rect 31208 4467 31224 4475
rect 31240 4467 31244 4475
rect 31248 4467 31252 4475
rect 31264 4467 31276 4475
rect 31280 4467 31292 4475
rect 31304 4467 31308 4475
rect 31312 4467 31316 4475
rect 31328 4467 31340 4475
rect 31344 4467 31348 4475
rect 31364 4467 31368 4475
rect 31372 4467 31384 4475
rect 31396 4467 31400 4475
rect 31404 4467 31408 4475
rect 31420 4467 31432 4475
rect 31436 4467 31440 4475
rect 31456 4467 31460 4475
rect 31464 4467 31476 4475
rect 31488 4467 31492 4475
rect 31496 4467 31500 4475
rect 31512 4467 31524 4475
rect 31528 4467 31532 4475
rect 31788 4467 31792 4475
rect 31796 4467 31800 4475
rect 31812 4467 31824 4475
rect 31828 4467 31832 4475
rect 31852 4467 31856 4475
rect 31860 4467 31864 4475
rect 31876 4467 31888 4475
rect 31892 4467 31904 4475
rect 31916 4467 31920 4475
rect 31924 4467 31928 4475
rect 31940 4467 31952 4475
rect 31956 4467 31968 4475
rect 31980 4467 31984 4475
rect 31988 4467 31992 4475
rect 32012 4467 32016 4475
rect 32020 4467 32024 4475
rect 32088 4467 32092 4475
rect 32096 4467 32108 4475
rect 32120 4467 32124 4475
rect 32128 4467 32132 4475
rect 32228 4467 32232 4475
rect 32236 4467 32240 4475
rect 32260 4467 32264 4475
rect 32268 4467 32272 4475
rect 32284 4467 32296 4475
rect 32300 4467 32304 4475
rect 32320 4467 32336 4475
rect 32352 4467 32400 4475
rect 32416 4467 32428 4475
rect 32432 4467 32436 4475
rect 32448 4467 32460 4475
rect 32472 4467 32476 4475
rect 32480 4467 32492 4475
rect 32496 4467 32500 4475
rect 32564 4467 32568 4475
rect 32572 4467 32584 4475
rect 32588 4467 32592 4475
rect 32632 4467 32644 4475
rect 32656 4467 32660 4475
rect 32664 4467 32676 4475
rect 32680 4467 32684 4475
rect 32724 4467 32736 4475
rect 32748 4467 32752 4475
rect 32756 4467 32768 4475
rect 32772 4467 32776 4475
rect 32788 4467 32800 4475
rect 32816 4467 32828 4475
rect 32840 4467 32844 4475
rect 32848 4467 32860 4475
rect 32864 4467 32868 4475
rect 32880 4467 32892 4475
rect 32912 4467 32924 4475
rect 32928 4467 32932 4475
rect 32944 4467 32956 4475
rect 32972 4467 32988 4475
rect 32996 4467 33028 4475
rect 33036 4467 33052 4475
rect 33068 4467 33080 4475
rect 33092 4467 33096 4475
rect 33100 4467 33112 4475
rect 33132 4467 33144 4475
rect 33164 4467 33176 4475
rect 33180 4467 33184 4475
rect 33196 4467 33208 4475
rect 33224 4467 33240 4475
rect 33248 4467 33280 4475
rect 33288 4467 33304 4475
rect 33320 4467 33332 4475
rect 33344 4467 33348 4475
rect 33352 4467 33364 4475
rect 33384 4467 33396 4475
rect 33408 4467 33412 4475
rect 33416 4467 33428 4475
rect 33432 4467 33436 4475
rect 33476 4467 33488 4475
rect 33500 4467 33504 4475
rect 33508 4467 33520 4475
rect 33524 4467 33528 4475
rect 33540 4467 33552 4475
rect 33728 4467 33740 4475
rect 33752 4467 33756 4475
rect 33760 4467 33772 4475
rect 33776 4467 33780 4475
rect 33820 4467 33832 4475
rect 33844 4467 33848 4475
rect 33852 4467 33864 4475
rect 33868 4467 33872 4475
rect 33936 4467 33940 4475
rect 33944 4467 33956 4475
rect 33960 4467 33964 4475
rect 34028 4467 34032 4475
rect 34036 4467 34048 4475
rect 34052 4467 34056 4475
rect 34068 4467 34080 4475
rect 34092 4467 34096 4475
rect 34100 4467 34112 4475
rect 34128 4467 34152 4475
rect 34160 4467 34172 4475
rect 34184 4467 34188 4475
rect 34192 4467 34204 4475
rect 34220 4467 34244 4475
rect 34252 4467 34268 4475
rect 34284 4467 34288 4475
rect 34292 4467 34296 4475
rect 34316 4467 34320 4475
rect 34324 4467 34336 4475
rect 34340 4467 34352 4475
rect 34356 4467 34360 4475
rect 34376 4467 34392 4475
rect 34408 4467 34412 4475
rect 34416 4467 34428 4475
rect 34432 4467 34444 4475
rect 34448 4467 34452 4475
rect 34472 4467 34476 4475
rect 34480 4467 34492 4475
rect 34504 4467 34508 4475
rect 34512 4467 34516 4475
rect 34536 4467 34540 4475
rect 34544 4467 34548 4475
rect 34644 4467 34648 4475
rect 34652 4467 34664 4475
rect 34668 4467 34680 4475
rect 34684 4467 34688 4475
rect 34708 4467 34712 4475
rect 34716 4467 34728 4475
rect 34740 4467 34744 4475
rect 34748 4467 34752 4475
rect 34864 4467 34868 4475
rect 34872 4467 34876 4475
rect 34940 4467 34944 4475
rect 34948 4467 34952 4475
rect 34972 4467 34976 4475
rect 34980 4467 34992 4475
rect 34996 4467 35008 4475
rect 35012 4467 35016 4475
rect 35036 4467 35040 4475
rect 35044 4467 35056 4475
rect 35064 4467 35080 4475
rect 35088 4467 35112 4475
rect 35128 4467 35140 4475
rect 35160 4467 35172 4475
rect 35184 4467 35188 4475
rect 35192 4467 35204 4475
rect 35208 4467 35212 4475
rect 35224 4467 35236 4475
rect 35252 4467 35268 4475
rect 35284 4467 35308 4475
rect 35316 4467 35332 4475
rect 35340 4467 35364 4475
rect 35380 4467 35396 4475
rect 35412 4467 35424 4475
rect 35436 4467 35440 4475
rect 35444 4467 35456 4475
rect 35460 4467 35464 4475
rect 35476 4467 35488 4475
rect 35500 4467 35504 4475
rect 35508 4467 35520 4475
rect 35524 4467 35528 4475
rect 35816 4467 35820 4475
rect 35824 4467 35836 4475
rect 35840 4467 35844 4475
rect 35856 4467 35868 4475
rect 35876 4467 35900 4475
rect 35916 4467 35940 4475
rect 35948 4467 35964 4475
rect 35980 4467 35996 4475
rect 36012 4467 36016 4475
rect 36020 4467 36032 4475
rect 36036 4467 36048 4475
rect 36052 4467 36056 4475
rect 36076 4467 36080 4475
rect 36084 4467 36096 4475
rect 36100 4467 36112 4475
rect 36116 4467 36120 4475
rect 36140 4467 36144 4475
rect 36148 4467 36152 4475
rect 36248 4467 36252 4475
rect 36256 4467 36268 4475
rect 36272 4467 36284 4475
rect 36288 4467 36292 4475
rect 36312 4467 36316 4475
rect 36320 4467 36324 4475
rect 36340 4467 36356 4475
rect 36364 4467 36388 4475
rect 36404 4467 36428 4475
rect 36436 4467 36452 4475
rect 36468 4467 36472 4475
rect 36476 4467 36480 4475
rect 36500 4467 36504 4475
rect 36508 4467 36520 4475
rect 36524 4467 36536 4475
rect 36540 4467 36544 4475
rect 36560 4467 36584 4475
rect 36592 4467 36608 4475
rect 36616 4467 36640 4475
rect 36656 4467 36668 4475
rect 36688 4467 36700 4475
rect 36712 4467 36716 4475
rect 36720 4467 36732 4475
rect 36736 4467 36740 4475
rect 36752 4467 36764 4475
rect 36776 4467 36780 4475
rect 36784 4467 36796 4475
rect 36812 4467 36836 4475
rect 36844 4467 36860 4475
rect 36876 4467 36892 4475
rect 36908 4467 36924 4475
rect 36932 4467 36956 4475
rect 36972 4467 36984 4475
rect 36988 4467 36992 4475
rect 37004 4467 37016 4475
rect 37028 4467 37032 4475
rect 37036 4467 37048 4475
rect 37052 4467 37056 4475
rect 37068 4467 37080 4475
rect 37092 4467 37096 4475
rect 37100 4467 37112 4475
rect 37132 4467 37144 4475
rect 37164 4467 37176 4475
rect 37196 4467 37208 4475
rect 37212 4467 37216 4475
rect 37228 4467 37240 4475
rect 37252 4467 37256 4475
rect 37260 4467 37272 4475
rect 37276 4467 37280 4475
rect 37292 4467 37304 4475
rect 37316 4467 37320 4475
rect 37324 4467 37336 4475
rect 37352 4467 37364 4475
rect 37368 4467 37372 4475
rect 37384 4467 37396 4475
rect 37408 4467 37412 4475
rect 37416 4467 37428 4475
rect 37432 4467 37436 4475
rect 37500 4467 37504 4475
rect 37508 4467 37520 4475
rect 37524 4467 37528 4475
rect 37540 4467 37552 4475
rect 37572 4467 37584 4475
rect 37600 4467 37624 4475
rect 37632 4467 37648 4475
rect 37656 4467 37680 4475
rect 37692 4467 37716 4475
rect 37724 4467 37740 4475
rect 37748 4467 37760 4475
rect 37764 4467 37768 4475
rect 37784 4467 37808 4475
rect 37816 4467 37832 4475
rect 37840 4467 37864 4475
rect 37880 4467 37884 4475
rect 37888 4467 37900 4475
rect 37912 4467 37916 4475
rect 37920 4467 37924 4475
rect 37944 4467 37948 4475
rect 37952 4467 37956 4475
rect 38020 4467 38024 4475
rect 38028 4467 38032 4475
rect 38160 4467 38164 4475
rect 38168 4467 38172 4475
rect 38184 4467 38196 4475
rect 38200 4467 38204 4475
rect 38220 4467 38244 4475
rect 38252 4467 38268 4475
rect 38276 4467 38288 4475
rect 38292 4467 38296 4475
rect 38312 4467 38336 4475
rect 38344 4467 38360 4475
rect 38368 4467 38392 4475
rect 38408 4467 38412 4475
rect 38416 4467 38428 4475
rect 38432 4467 38444 4475
rect 38448 4467 38452 4475
rect 38472 4467 38476 4475
rect 38480 4467 38484 4475
rect 38500 4467 38516 4475
rect 38524 4467 38548 4475
rect 38564 4467 38588 4475
rect 38596 4467 38612 4475
rect 38628 4467 38644 4475
rect 38660 4467 38676 4475
rect 38684 4467 38708 4475
rect 38724 4467 38748 4475
rect 38756 4467 38768 4475
rect 38780 4467 38784 4475
rect 38788 4467 38800 4475
rect 38816 4467 38840 4475
rect 38848 4467 38860 4475
rect 38872 4467 38876 4475
rect 38880 4467 38892 4475
rect 38908 4467 38920 4475
rect 38924 4467 38928 4475
rect 38940 4467 38952 4475
rect 38960 4467 38984 4475
rect 39000 4467 39012 4475
rect 39016 4467 39020 4475
rect 39032 4467 39044 4475
rect 39056 4467 39060 4475
rect 39064 4467 39076 4475
rect 39080 4467 39084 4475
rect 39096 4467 39108 4475
rect 39128 4467 39140 4475
rect 39156 4467 39180 4475
rect 39188 4467 39200 4475
rect 39212 4467 39236 4475
rect 39252 4467 39256 4475
rect 39260 4467 39272 4475
rect 39276 4467 39288 4475
rect 39292 4467 39296 4475
rect 39316 4467 39320 4475
rect 39324 4467 39336 4475
rect 39344 4467 39360 4475
rect 39368 4467 39392 4475
rect 39408 4467 39424 4475
rect 39440 4467 39452 4475
rect 39464 4467 39468 4475
rect 39472 4467 39484 4475
rect 39488 4467 39492 4475
rect 39716 4467 39720 4475
rect 39724 4467 39736 4475
rect 39740 4467 39744 4475
rect 39756 4467 39768 4475
rect 39776 4467 39800 4475
rect 39816 4467 39864 4475
rect 39880 4467 39892 4475
rect 39908 4467 39956 4475
rect 39972 4467 39988 4475
rect 40000 4467 40008 4475
rect 40012 4467 40024 4475
rect 40036 4467 40040 4475
rect 40044 4467 40048 4475
rect 40060 4467 40072 4475
rect 40076 4467 40080 4475
rect 40176 4467 40180 4475
rect 40184 4467 40188 4475
rect 40200 4467 40212 4475
rect 40216 4467 40220 4475
rect 40240 4467 40244 4475
rect 40248 4467 40252 4475
rect 40268 4467 40316 4475
rect 40332 4467 40356 4475
rect 40364 4467 40380 4475
rect 40396 4467 40420 4475
rect 40428 4467 40444 4475
rect 40452 4467 40476 4475
rect 40492 4467 40496 4475
rect 40500 4467 40512 4475
rect 40520 4467 40536 4475
rect 40544 4467 40556 4475
rect 40560 4467 40564 4475
rect 40584 4467 40588 4475
rect 40592 4467 40604 4475
rect 40612 4467 40628 4475
rect 40636 4467 40648 4475
rect 40652 4467 40656 4475
rect 40676 4467 40680 4475
rect 40684 4467 40696 4475
rect 40708 4467 40712 4475
rect 40716 4467 40720 4475
rect 40740 4467 40744 4475
rect 40748 4467 40752 4475
rect 24410 4450 24420 4458
rect 24624 4450 24634 4458
rect 25900 4450 25902 4458
rect 25908 4450 25910 4458
rect 33280 4457 33288 4465
rect 40480 4457 40488 4465
rect 18672 4440 18680 4448
rect 19296 4440 19304 4448
rect 29760 4437 29768 4445
rect 31504 4437 31512 4445
rect 32816 4437 32824 4445
rect 37424 4437 37432 4445
rect 30128 4417 30136 4425
rect 30592 4417 30600 4425
rect 31264 4417 31272 4425
rect 31872 4417 31880 4425
rect 32288 4417 32296 4425
rect 33408 4417 33416 4425
rect 33936 4417 33944 4425
rect 35488 4417 35496 4425
rect 20336 4400 20344 4408
rect 31792 4397 31800 4405
rect 33808 4397 33816 4405
rect 36288 4397 36296 4405
rect 38640 4397 38648 4405
rect 39616 4397 39624 4405
rect 25760 4380 25768 4388
rect 26688 4380 26696 4388
rect 27744 4380 27752 4388
rect 29568 4377 29576 4385
rect 30704 4377 30712 4385
rect 30960 4377 30968 4385
rect 32656 4377 32664 4385
rect 33536 4377 33544 4385
rect 33984 4377 33992 4385
rect 34672 4377 34680 4385
rect 34768 4377 34776 4385
rect 34960 4377 34968 4385
rect 36256 4377 36264 4385
rect 37664 4377 37672 4385
rect 39888 4377 39896 4385
rect 40688 4377 40696 4385
rect 18832 4360 18840 4368
rect 19104 4360 19112 4368
rect 19456 4360 19464 4368
rect 19520 4360 19528 4368
rect 20544 4360 20552 4368
rect 21100 4361 21110 4366
rect 21296 4360 21304 4368
rect 21312 4360 21320 4368
rect 21360 4360 21368 4368
rect 23040 4360 23048 4368
rect 23392 4360 23400 4368
rect 24116 4361 24119 4366
rect 24465 4361 24468 4366
rect 24960 4360 24968 4368
rect 25596 4361 25606 4366
rect 26672 4360 26680 4368
rect 27104 4360 27112 4368
rect 27472 4360 27480 4368
rect 27744 4360 27752 4368
rect 31056 4357 31064 4365
rect 34496 4357 34504 4365
rect 38464 4357 38472 4365
rect 21760 4340 21768 4348
rect 23696 4340 23704 4348
rect 27280 4340 27288 4348
rect 29680 4337 29688 4345
rect 30688 4337 30696 4345
rect 31264 4337 31272 4345
rect 31392 4337 31400 4345
rect 31488 4337 31496 4345
rect 32000 4337 32008 4345
rect 32960 4337 32968 4345
rect 33472 4337 33480 4345
rect 33504 4337 33512 4345
rect 33520 4337 33528 4345
rect 33760 4337 33768 4345
rect 33824 4337 33832 4345
rect 33920 4337 33928 4345
rect 34336 4337 34344 4345
rect 34352 4337 34360 4345
rect 34560 4337 34568 4345
rect 34672 4337 34680 4345
rect 35648 4337 35656 4345
rect 36176 4337 36184 4345
rect 36192 4337 36200 4345
rect 36592 4337 36600 4345
rect 36832 4337 36840 4345
rect 37392 4337 37400 4345
rect 37584 4337 37592 4345
rect 37600 4337 37608 4345
rect 37824 4337 37832 4345
rect 38352 4337 38360 4345
rect 39040 4337 39048 4345
rect 39296 4337 39304 4345
rect 39712 4337 39720 4345
rect 18624 4320 18632 4328
rect 19120 4320 19128 4328
rect 19696 4320 19704 4328
rect 19728 4320 19736 4328
rect 20352 4320 20360 4328
rect 21584 4320 21592 4328
rect 22000 4320 22008 4328
rect 22432 4320 22440 4328
rect 22576 4320 22584 4328
rect 22624 4320 22632 4328
rect 23056 4320 23064 4328
rect 23392 4320 23400 4328
rect 24128 4320 24136 4328
rect 24288 4320 24296 4328
rect 24976 4320 24984 4328
rect 25952 4320 25960 4328
rect 26480 4320 26488 4328
rect 26688 4320 26696 4328
rect 28160 4320 28168 4328
rect 28192 4320 28200 4328
rect 28528 4320 28536 4328
rect 29440 4317 29448 4325
rect 29616 4317 29624 4325
rect 35216 4317 35224 4325
rect 35344 4317 35352 4325
rect 36048 4317 36056 4325
rect 36528 4317 36536 4325
rect 36816 4317 36824 4325
rect 37776 4317 37784 4325
rect 38160 4317 38168 4325
rect 39648 4317 39656 4325
rect 19328 4300 19336 4308
rect 20128 4300 20136 4308
rect 20880 4300 20888 4308
rect 21280 4300 21288 4308
rect 22816 4300 22824 4308
rect 23488 4300 23496 4308
rect 23920 4300 23928 4308
rect 24528 4300 24536 4308
rect 24688 4300 24696 4308
rect 24880 4300 24888 4308
rect 25200 4300 25208 4308
rect 26240 4300 26248 4308
rect 27280 4300 27288 4308
rect 30520 4305 30521 4310
rect 31824 4297 31832 4305
rect 32576 4297 32584 4305
rect 33200 4297 33208 4305
rect 33328 4297 33336 4305
rect 33392 4297 33400 4305
rect 33840 4297 33848 4305
rect 34000 4297 34008 4305
rect 34016 4297 34024 4305
rect 37936 4297 37944 4305
rect 37952 4297 37960 4305
rect 38272 4297 38280 4305
rect 38800 4297 38808 4305
rect 39344 4297 39352 4305
rect 39440 4297 39448 4305
rect 40496 4297 40504 4305
rect 40576 4297 40584 4305
rect 18464 4280 18472 4288
rect 23840 4280 23848 4288
rect 24736 4280 24744 4288
rect 25728 4280 25736 4288
rect 27392 4280 27400 4288
rect 29904 4277 29912 4285
rect 30224 4277 30232 4285
rect 31792 4277 31800 4285
rect 32368 4277 32376 4285
rect 37264 4277 37272 4285
rect 37392 4277 37400 4285
rect 39616 4277 39624 4285
rect 40048 4277 40056 4285
rect 40208 4277 40216 4285
rect 40224 4277 40232 4285
rect 40272 4277 40280 4285
rect 19488 4260 19496 4268
rect 24288 4260 24296 4268
rect 26832 4260 26840 4268
rect 27056 4260 27064 4268
rect 28336 4260 28344 4268
rect 28384 4260 28392 4268
rect 29428 4267 29440 4275
rect 29444 4267 29448 4275
rect 29460 4267 29472 4275
rect 29488 4267 29504 4275
rect 29512 4267 29544 4275
rect 29552 4267 29564 4275
rect 29584 4267 29596 4275
rect 29600 4267 29612 4275
rect 29616 4267 29628 4275
rect 29644 4267 29656 4275
rect 29676 4267 29688 4275
rect 29692 4267 29704 4275
rect 29708 4267 29720 4275
rect 29740 4267 29752 4275
rect 29760 4267 29792 4275
rect 29800 4267 29816 4275
rect 29824 4267 29836 4275
rect 29840 4267 29844 4275
rect 29864 4267 29868 4275
rect 29872 4267 29884 4275
rect 29896 4267 29900 4275
rect 29904 4267 29908 4275
rect 30052 4267 30056 4275
rect 30060 4267 30064 4275
rect 30076 4267 30088 4275
rect 30092 4267 30096 4275
rect 30112 4267 30136 4275
rect 30144 4267 30160 4275
rect 30168 4267 30200 4275
rect 30216 4267 30220 4275
rect 30224 4267 30228 4275
rect 30248 4267 30252 4275
rect 30256 4267 30268 4275
rect 30280 4267 30284 4275
rect 30288 4267 30292 4275
rect 30356 4267 30360 4275
rect 30364 4267 30376 4275
rect 30432 4267 30436 4275
rect 30440 4267 30452 4275
rect 30472 4267 30484 4275
rect 30488 4267 30492 4275
rect 30508 4267 30524 4275
rect 30540 4267 30556 4275
rect 30564 4267 30580 4275
rect 30588 4267 30600 4275
rect 30616 4267 30632 4275
rect 30640 4267 30672 4275
rect 30680 4267 30696 4275
rect 30712 4267 30724 4275
rect 30732 4267 30764 4275
rect 30772 4267 30788 4275
rect 30796 4267 30820 4275
rect 30836 4267 30852 4275
rect 30868 4267 30880 4275
rect 30892 4267 30896 4275
rect 30900 4267 30912 4275
rect 30916 4267 30920 4275
rect 30984 4267 30988 4275
rect 30992 4267 31004 4275
rect 31008 4267 31012 4275
rect 31024 4267 31036 4275
rect 31056 4267 31068 4275
rect 31084 4267 31108 4275
rect 31116 4267 31132 4275
rect 31140 4267 31152 4275
rect 31156 4267 31160 4275
rect 31180 4267 31184 4275
rect 31188 4267 31200 4275
rect 31204 4267 31216 4275
rect 31220 4267 31224 4275
rect 31272 4267 31276 4275
rect 31280 4267 31292 4275
rect 31296 4267 31308 4275
rect 31312 4267 31316 4275
rect 31336 4267 31340 4275
rect 31344 4267 31348 4275
rect 31444 4267 31448 4275
rect 31452 4267 31464 4275
rect 31468 4267 31480 4275
rect 31484 4267 31488 4275
rect 31508 4267 31512 4275
rect 31516 4267 31520 4275
rect 31536 4267 31540 4275
rect 31544 4267 31556 4275
rect 31560 4267 31572 4275
rect 31576 4267 31580 4275
rect 31788 4267 31792 4275
rect 31796 4267 31808 4275
rect 31812 4267 31824 4275
rect 31828 4267 31832 4275
rect 32136 4267 32140 4275
rect 32144 4267 32148 4275
rect 32168 4267 32172 4275
rect 32176 4267 32188 4275
rect 32192 4267 32204 4275
rect 32208 4267 32212 4275
rect 32228 4267 32244 4275
rect 32260 4267 32264 4275
rect 32268 4267 32280 4275
rect 32284 4267 32296 4275
rect 32300 4267 32304 4275
rect 32320 4267 32336 4275
rect 32352 4267 32356 4275
rect 32360 4267 32372 4275
rect 32376 4267 32388 4275
rect 32392 4267 32396 4275
rect 32412 4267 32428 4275
rect 32444 4267 32460 4275
rect 32468 4267 32492 4275
rect 32508 4267 32520 4275
rect 32524 4267 32528 4275
rect 32540 4267 32552 4275
rect 32564 4267 32568 4275
rect 32572 4267 32584 4275
rect 32688 4267 32692 4275
rect 32696 4267 32708 4275
rect 32912 4267 32924 4275
rect 32944 4267 32956 4275
rect 32960 4267 32964 4275
rect 32976 4267 32988 4275
rect 33000 4267 33004 4275
rect 33008 4267 33020 4275
rect 33036 4267 33060 4275
rect 33068 4267 33080 4275
rect 33092 4267 33096 4275
rect 33100 4267 33112 4275
rect 33116 4267 33120 4275
rect 33132 4267 33144 4275
rect 33164 4267 33176 4275
rect 33192 4267 33216 4275
rect 33224 4267 33240 4275
rect 33248 4267 33280 4275
rect 33288 4267 33304 4275
rect 33320 4267 33332 4275
rect 33336 4267 33348 4275
rect 33352 4267 33364 4275
rect 33384 4267 33396 4275
rect 33404 4267 33436 4275
rect 33444 4267 33456 4275
rect 33476 4267 33488 4275
rect 33496 4267 33528 4275
rect 33536 4267 33552 4275
rect 33568 4267 33580 4275
rect 33592 4267 33596 4275
rect 33600 4267 33612 4275
rect 33632 4267 33644 4275
rect 33664 4267 33676 4275
rect 33680 4267 33684 4275
rect 33696 4267 33708 4275
rect 33728 4267 33740 4275
rect 33744 4267 33756 4275
rect 33760 4267 33772 4275
rect 33876 4267 33880 4275
rect 33884 4267 33896 4275
rect 33916 4267 33928 4275
rect 33932 4267 33944 4275
rect 33948 4267 33960 4275
rect 33976 4267 33992 4275
rect 34008 4267 34020 4275
rect 34024 4267 34036 4275
rect 34040 4267 34052 4275
rect 34072 4267 34084 4275
rect 34088 4267 34092 4275
rect 34164 4267 34176 4275
rect 34180 4267 34184 4275
rect 34288 4267 34300 4275
rect 34304 4267 34308 4275
rect 34320 4267 34332 4275
rect 34344 4267 34348 4275
rect 34352 4267 34364 4275
rect 34380 4267 34392 4275
rect 34396 4267 34400 4275
rect 34412 4267 34424 4275
rect 34432 4267 34456 4275
rect 34472 4267 34496 4275
rect 34504 4267 34520 4275
rect 34536 4267 34552 4275
rect 34568 4267 34584 4275
rect 34592 4267 34616 4275
rect 34632 4267 34680 4275
rect 34696 4267 34700 4275
rect 34704 4267 34708 4275
rect 34720 4267 34732 4275
rect 34736 4267 34748 4275
rect 34756 4267 34772 4275
rect 34788 4267 34804 4275
rect 34812 4267 34824 4275
rect 34828 4267 34840 4275
rect 34852 4267 34856 4275
rect 34860 4267 34864 4275
rect 34880 4267 34896 4275
rect 34904 4267 34928 4275
rect 34944 4267 34956 4275
rect 34976 4267 34988 4275
rect 34992 4267 35004 4275
rect 35008 4267 35020 4275
rect 35036 4267 35052 4275
rect 35068 4267 35080 4275
rect 35084 4267 35096 4275
rect 35100 4267 35112 4275
rect 35128 4267 35140 4275
rect 35160 4267 35172 4275
rect 35176 4267 35188 4275
rect 35192 4267 35200 4275
rect 35224 4267 35236 4275
rect 35252 4267 35276 4275
rect 35284 4267 35300 4275
rect 35316 4267 35332 4275
rect 35340 4267 35364 4275
rect 35380 4267 35396 4275
rect 35412 4267 35424 4275
rect 35428 4267 35440 4275
rect 35444 4267 35456 4275
rect 35476 4267 35488 4275
rect 35492 4267 35504 4275
rect 35508 4267 35520 4275
rect 35536 4267 35548 4275
rect 35568 4267 35580 4275
rect 35584 4267 35596 4275
rect 35600 4267 35612 4275
rect 35632 4267 35644 4275
rect 35660 4267 35684 4275
rect 35692 4267 35708 4275
rect 35724 4267 35728 4275
rect 35732 4267 35736 4275
rect 35748 4267 35760 4275
rect 35764 4267 35776 4275
rect 35788 4267 35792 4275
rect 35796 4267 35800 4275
rect 35816 4267 35832 4275
rect 35840 4267 35864 4275
rect 35880 4267 35892 4275
rect 35912 4267 35924 4275
rect 35928 4267 35940 4275
rect 35944 4267 35956 4275
rect 35976 4267 35988 4275
rect 36004 4267 36016 4275
rect 36020 4267 36032 4275
rect 36036 4267 36048 4275
rect 36068 4267 36080 4275
rect 36092 4267 36096 4275
rect 36100 4267 36112 4275
rect 36132 4267 36144 4275
rect 36256 4267 36268 4275
rect 36272 4267 36276 4275
rect 36288 4267 36300 4275
rect 36320 4267 36332 4275
rect 36340 4267 36372 4275
rect 36380 4267 36396 4275
rect 36404 4267 36428 4275
rect 36444 4267 36460 4275
rect 36468 4267 36492 4275
rect 36508 4267 36556 4275
rect 36572 4267 36576 4275
rect 36580 4267 36584 4275
rect 36596 4267 36608 4275
rect 36612 4267 36624 4275
rect 36636 4267 36640 4275
rect 36644 4267 36648 4275
rect 36664 4267 36668 4275
rect 36672 4267 36676 4275
rect 36688 4267 36700 4275
rect 36704 4267 36716 4275
rect 36728 4267 36732 4275
rect 36736 4267 36740 4275
rect 36756 4267 36800 4275
rect 36820 4267 36832 4275
rect 36852 4267 36864 4275
rect 36876 4267 36880 4275
rect 36884 4267 36896 4275
rect 36916 4267 36928 4275
rect 36932 4267 36936 4275
rect 36968 4267 36972 4275
rect 36976 4267 36988 4275
rect 37008 4267 37020 4275
rect 37024 4267 37028 4275
rect 37132 4267 37144 4275
rect 37148 4267 37152 4275
rect 37164 4267 37176 4275
rect 37196 4267 37208 4275
rect 37224 4267 37272 4275
rect 37288 4267 37304 4275
rect 37312 4267 37336 4275
rect 37352 4267 37364 4275
rect 37384 4267 37396 4275
rect 37400 4267 37412 4275
rect 37416 4267 37428 4275
rect 37444 4267 37456 4275
rect 37476 4267 37488 4275
rect 37492 4267 37504 4275
rect 37508 4267 37520 4275
rect 37540 4267 37552 4275
rect 37568 4267 37592 4275
rect 37600 4267 37616 4275
rect 37632 4267 37636 4275
rect 37640 4267 37644 4275
rect 37656 4267 37668 4275
rect 37672 4267 37684 4275
rect 37692 4267 37708 4275
rect 37724 4267 37740 4275
rect 37748 4267 37760 4275
rect 37764 4267 37776 4275
rect 37784 4267 37800 4275
rect 37816 4267 37832 4275
rect 37840 4267 37852 4275
rect 37856 4267 37868 4275
rect 37880 4267 37884 4275
rect 37888 4267 37892 4275
rect 37912 4267 37916 4275
rect 37920 4267 37932 4275
rect 37944 4267 37948 4275
rect 37952 4267 37956 4275
rect 37976 4267 37980 4275
rect 37984 4267 37988 4275
rect 38000 4267 38012 4275
rect 38016 4267 38020 4275
rect 38036 4267 38052 4275
rect 38068 4267 38116 4275
rect 38132 4267 38136 4275
rect 38140 4267 38144 4275
rect 38160 4267 38208 4275
rect 38224 4267 38236 4275
rect 38240 4267 38244 4275
rect 38256 4267 38268 4275
rect 38280 4267 38284 4275
rect 38288 4267 38300 4275
rect 38316 4267 38328 4275
rect 38332 4267 38336 4275
rect 38348 4267 38360 4275
rect 38368 4267 38392 4275
rect 38408 4267 38456 4275
rect 38472 4267 38488 4275
rect 38504 4267 38516 4275
rect 38528 4267 38532 4275
rect 38536 4267 38548 4275
rect 38568 4267 38580 4275
rect 38584 4267 38588 4275
rect 38600 4267 38612 4275
rect 38628 4267 38644 4275
rect 38660 4267 38708 4275
rect 38724 4267 38740 4275
rect 38752 4267 38800 4275
rect 38816 4267 38832 4275
rect 38848 4267 38860 4275
rect 38872 4267 38876 4275
rect 38880 4267 38892 4275
rect 39160 4267 39172 4275
rect 39176 4267 39180 4275
rect 39192 4267 39200 4275
rect 39212 4267 39236 4275
rect 39252 4267 39300 4275
rect 39316 4267 39320 4275
rect 39324 4267 39328 4275
rect 39344 4267 39392 4275
rect 39408 4267 39424 4275
rect 39436 4267 39484 4275
rect 39500 4267 39512 4275
rect 39528 4267 39576 4275
rect 39592 4267 39608 4275
rect 39624 4267 39640 4275
rect 39656 4267 39672 4275
rect 39688 4267 39736 4275
rect 39752 4267 39768 4275
rect 39776 4267 39800 4275
rect 39816 4267 39832 4275
rect 39840 4267 39872 4275
rect 39880 4267 39892 4275
rect 39908 4267 39924 4275
rect 39932 4267 39964 4275
rect 39972 4267 39988 4275
rect 40000 4267 40008 4275
rect 40012 4267 40016 4275
rect 40036 4267 40040 4275
rect 40044 4267 40056 4275
rect 40060 4267 40072 4275
rect 40076 4267 40080 4275
rect 40100 4267 40104 4275
rect 40108 4267 40112 4275
rect 40176 4267 40180 4275
rect 40184 4267 40188 4275
rect 40208 4267 40212 4275
rect 40216 4267 40220 4275
rect 40232 4267 40244 4275
rect 40248 4267 40252 4275
rect 40272 4267 40276 4275
rect 40280 4267 40292 4275
rect 40304 4267 40308 4275
rect 40312 4267 40316 4275
rect 40336 4267 40340 4275
rect 40344 4267 40356 4275
rect 40368 4267 40372 4275
rect 40376 4267 40380 4275
rect 40392 4267 40404 4275
rect 40408 4267 40420 4275
rect 40432 4267 40436 4275
rect 40440 4267 40444 4275
rect 40456 4267 40468 4275
rect 40472 4267 40476 4275
rect 40492 4267 40496 4275
rect 40500 4267 40512 4275
rect 40524 4267 40528 4275
rect 40532 4267 40536 4275
rect 40632 4267 40636 4275
rect 40640 4267 40644 4275
rect 40664 4267 40668 4275
rect 40672 4267 40684 4275
rect 40688 4267 40700 4275
rect 40704 4267 40708 4275
rect 40756 4267 40760 4275
rect 40764 4267 40776 4275
rect 40780 4267 40792 4275
rect 40796 4267 40800 4275
rect 19816 4252 19818 4260
rect 20768 4250 20772 4258
rect 20858 4250 20866 4258
rect 20982 4252 20984 4260
rect 21164 4250 21168 4258
rect 21254 4250 21262 4258
rect 21340 4250 21348 4258
rect 21490 4250 21496 4258
rect 21554 4250 21562 4258
rect 21704 4250 21710 4258
rect 22304 4252 22306 4260
rect 22518 4252 22520 4260
rect 23272 4250 23276 4258
rect 23362 4250 23370 4258
rect 23448 4250 23456 4258
rect 23598 4250 23604 4258
rect 24090 4250 24104 4258
rect 24946 4250 24960 4258
rect 25160 4250 25174 4258
rect 25930 4250 25944 4258
rect 26016 4250 26030 4258
rect 26444 4250 26458 4258
rect 26658 4250 26672 4258
rect 27086 4250 27100 4258
rect 27728 4250 27742 4258
rect 27942 4250 27956 4258
rect 28156 4250 28170 4258
rect 35840 4257 35848 4265
rect 39200 4257 39208 4265
rect 21920 4240 21928 4248
rect 27424 4240 27432 4248
rect 27472 4240 27480 4248
rect 30032 4237 30040 4245
rect 30224 4237 30232 4245
rect 30320 4237 30328 4245
rect 31568 4237 31576 4245
rect 31776 4237 31784 4245
rect 32416 4237 32424 4245
rect 32592 4237 32600 4245
rect 32624 4237 32632 4245
rect 32672 4237 32680 4245
rect 33216 4237 33224 4245
rect 33600 4237 33608 4245
rect 34208 4237 34216 4245
rect 34624 4237 34632 4245
rect 35408 4237 35416 4245
rect 35472 4237 35480 4245
rect 35872 4237 35880 4245
rect 36032 4237 36040 4245
rect 36064 4237 36072 4245
rect 36400 4237 36408 4245
rect 37072 4237 37080 4245
rect 38224 4237 38232 4245
rect 19040 4220 19048 4228
rect 20112 4220 20120 4228
rect 20496 4220 20504 4228
rect 21312 4220 21320 4228
rect 24224 4220 24232 4228
rect 24432 4220 24440 4228
rect 24448 4220 24456 4228
rect 26144 4220 26152 4228
rect 28656 4220 28664 4228
rect 30736 4217 30744 4225
rect 30784 4217 30792 4225
rect 31184 4217 31192 4225
rect 36096 4217 36104 4225
rect 36416 4217 36424 4225
rect 36592 4217 36600 4225
rect 38096 4217 38104 4225
rect 38368 4217 38376 4225
rect 38544 4217 38552 4225
rect 38608 4217 38616 4225
rect 38816 4217 38824 4225
rect 39040 4217 39048 4225
rect 39840 4217 39848 4225
rect 39952 4217 39960 4225
rect 20720 4200 20728 4208
rect 25808 4200 25816 4208
rect 29856 4197 29864 4205
rect 29952 4197 29960 4205
rect 30960 4197 30968 4205
rect 31472 4197 31480 4205
rect 32752 4197 32760 4205
rect 33136 4197 33144 4205
rect 33616 4197 33624 4205
rect 33648 4197 33656 4205
rect 33792 4197 33800 4205
rect 34144 4197 34152 4205
rect 34224 4197 34232 4205
rect 34720 4197 34728 4205
rect 35104 4197 35112 4205
rect 35200 4197 35208 4205
rect 35600 4197 35608 4205
rect 36288 4197 36296 4205
rect 36800 4197 36808 4205
rect 37072 4197 37080 4205
rect 37328 4197 37336 4205
rect 37488 4197 37496 4205
rect 38400 4197 38408 4205
rect 39280 4197 39288 4205
rect 39376 4197 39384 4205
rect 39568 4197 39576 4205
rect 40064 4197 40072 4205
rect 40304 4197 40312 4205
rect 18624 4180 18632 4188
rect 18704 4180 18712 4188
rect 18896 4180 18904 4188
rect 19216 4180 19224 4188
rect 19712 4180 19720 4188
rect 19920 4180 19928 4188
rect 21136 4180 21144 4188
rect 21456 4180 21464 4188
rect 21664 4180 21672 4188
rect 22192 4180 22200 4188
rect 23152 4180 23160 4188
rect 23248 4180 23256 4188
rect 23760 4180 23768 4188
rect 24928 4180 24936 4188
rect 25472 4180 25480 4188
rect 25744 4180 25752 4188
rect 26000 4180 26008 4188
rect 26432 4180 26440 4188
rect 26640 4180 26648 4188
rect 27392 4180 27400 4188
rect 27616 4180 27624 4188
rect 28144 4180 28152 4188
rect 30256 4177 30264 4185
rect 30816 4177 30824 4185
rect 32448 4177 32456 4185
rect 33456 4177 33464 4185
rect 33568 4177 33576 4185
rect 33600 4177 33608 4185
rect 34912 4177 34920 4185
rect 35856 4177 35864 4185
rect 36096 4177 36104 4185
rect 37856 4177 37864 4185
rect 21072 4160 21080 4168
rect 27024 4160 27032 4168
rect 27216 4160 27224 4168
rect 29392 4157 29400 4165
rect 29504 4157 29512 4165
rect 29728 4157 29736 4165
rect 30384 4157 30392 4165
rect 30608 4157 30616 4165
rect 30832 4157 30840 4165
rect 31600 4157 31608 4165
rect 32288 4157 32296 4165
rect 34160 4157 34168 4165
rect 34240 4157 34248 4165
rect 34336 4157 34344 4165
rect 34784 4157 34792 4165
rect 35136 4157 35144 4165
rect 36720 4157 36728 4165
rect 36832 4157 36840 4165
rect 38384 4157 38392 4165
rect 38528 4157 38536 4165
rect 38928 4157 38936 4165
rect 39120 4157 39128 4165
rect 39232 4157 39240 4165
rect 39328 4157 39336 4165
rect 39488 4157 39496 4165
rect 40080 4157 40088 4165
rect 40592 4157 40600 4165
rect 20688 4148 20692 4153
rect 21694 4148 21698 4153
rect 22962 4148 22966 4153
rect 25712 4148 25716 4153
rect 28134 4148 28141 4153
rect 18880 4140 18888 4148
rect 19280 4140 19288 4148
rect 20272 4140 20280 4148
rect 22160 4140 22168 4148
rect 22176 4140 22184 4148
rect 22400 4140 22408 4148
rect 23232 4140 23240 4148
rect 23408 4140 23416 4148
rect 23584 4140 23592 4148
rect 24000 4140 24008 4148
rect 24496 4140 24504 4148
rect 25984 4140 25992 4148
rect 26416 4140 26424 4148
rect 27056 4140 27064 4148
rect 27264 4140 27272 4148
rect 28336 4140 28344 4148
rect 37280 4137 37288 4145
rect 40288 4117 40296 4125
rect 18672 4100 18680 4108
rect 19888 4100 19896 4108
rect 26208 4100 26216 4108
rect 26352 4100 26360 4108
rect 33664 4097 33672 4105
rect 39344 4097 39352 4105
rect 39376 4097 39384 4105
rect 40544 4097 40552 4105
rect 19904 4080 19912 4088
rect 26576 4080 26584 4088
rect 29808 4077 29816 4085
rect 23200 4060 23208 4068
rect 29420 4067 29424 4075
rect 29428 4067 29440 4075
rect 29444 4067 29448 4075
rect 29488 4067 29500 4075
rect 29512 4067 29516 4075
rect 29520 4067 29532 4075
rect 29536 4067 29540 4075
rect 29644 4067 29656 4075
rect 29736 4067 29748 4075
rect 29828 4067 29840 4075
rect 29852 4067 29856 4075
rect 29860 4067 29872 4075
rect 29876 4067 29880 4075
rect 29892 4067 29904 4075
rect 29920 4067 29936 4075
rect 29952 4067 29976 4075
rect 29984 4067 30000 4075
rect 30008 4067 30032 4075
rect 30048 4067 30060 4075
rect 30080 4067 30092 4075
rect 30104 4067 30108 4075
rect 30112 4067 30124 4075
rect 30128 4067 30132 4075
rect 30144 4067 30156 4075
rect 30168 4067 30172 4075
rect 30176 4067 30188 4075
rect 30192 4067 30196 4075
rect 30292 4067 30296 4075
rect 30300 4067 30304 4075
rect 30324 4067 30328 4075
rect 30332 4067 30344 4075
rect 30348 4067 30352 4075
rect 30392 4067 30400 4075
rect 30416 4067 30420 4075
rect 30424 4067 30428 4075
rect 30476 4067 30480 4075
rect 30484 4067 30496 4075
rect 30584 4067 30588 4075
rect 30592 4067 30596 4075
rect 30616 4067 30620 4075
rect 30624 4067 30628 4075
rect 30640 4067 30652 4075
rect 30656 4067 30660 4075
rect 30680 4067 30684 4075
rect 30688 4067 30700 4075
rect 30708 4067 30724 4075
rect 30732 4067 30744 4075
rect 30748 4067 30752 4075
rect 30772 4067 30776 4075
rect 30780 4067 30792 4075
rect 30796 4067 30808 4075
rect 30812 4067 30816 4075
rect 30864 4067 30868 4075
rect 30872 4067 30884 4075
rect 30888 4067 30892 4075
rect 30904 4067 30916 4075
rect 30932 4067 30944 4075
rect 30956 4067 30960 4075
rect 30964 4067 30976 4075
rect 30980 4067 30984 4075
rect 30996 4067 31008 4075
rect 31028 4067 31040 4075
rect 31060 4067 31072 4075
rect 31092 4067 31104 4075
rect 31116 4067 31120 4075
rect 31124 4067 31136 4075
rect 31140 4067 31144 4075
rect 31156 4067 31168 4075
rect 31248 4067 31260 4075
rect 31532 4067 31544 4075
rect 31548 4067 31552 4075
rect 31564 4067 31576 4075
rect 31584 4067 31608 4075
rect 31624 4067 31648 4075
rect 31656 4067 31668 4075
rect 31680 4067 31684 4075
rect 31688 4067 31700 4075
rect 31720 4067 31732 4075
rect 31744 4067 31748 4075
rect 31752 4067 31764 4075
rect 31836 4067 31840 4075
rect 31844 4067 31856 4075
rect 31876 4067 31888 4075
rect 31892 4067 31896 4075
rect 32008 4067 32012 4075
rect 32016 4067 32020 4075
rect 32040 4067 32044 4075
rect 32048 4067 32052 4075
rect 32064 4067 32076 4075
rect 32080 4067 32084 4075
rect 32100 4067 32124 4075
rect 32132 4067 32148 4075
rect 32156 4067 32188 4075
rect 32196 4067 32208 4075
rect 32228 4067 32240 4075
rect 32248 4067 32280 4075
rect 32288 4067 32300 4075
rect 32320 4067 32332 4075
rect 32340 4067 32372 4075
rect 32380 4067 32392 4075
rect 32412 4067 32424 4075
rect 32436 4067 32440 4075
rect 32444 4067 32456 4075
rect 32600 4067 32612 4075
rect 32616 4067 32620 4075
rect 32632 4067 32644 4075
rect 32664 4067 32676 4075
rect 32684 4067 32716 4075
rect 32724 4067 32736 4075
rect 32752 4067 32768 4075
rect 32776 4067 32800 4075
rect 32816 4067 32828 4075
rect 32844 4067 32860 4075
rect 32868 4067 32900 4075
rect 32908 4067 32920 4075
rect 32940 4067 32952 4075
rect 32960 4067 32992 4075
rect 33000 4067 33016 4075
rect 33032 4067 33044 4075
rect 33056 4067 33060 4075
rect 33064 4067 33076 4075
rect 33096 4067 33108 4075
rect 33120 4067 33124 4075
rect 33128 4067 33140 4075
rect 33144 4067 33148 4075
rect 33160 4067 33172 4075
rect 33188 4067 33200 4075
rect 33212 4067 33216 4075
rect 33220 4067 33232 4075
rect 33236 4067 33240 4075
rect 33252 4067 33264 4075
rect 33276 4067 33280 4075
rect 33284 4067 33296 4075
rect 33312 4067 33360 4075
rect 33376 4067 33400 4075
rect 33408 4067 33420 4075
rect 33432 4067 33436 4075
rect 33440 4067 33452 4075
rect 33456 4067 33460 4075
rect 33472 4067 33484 4075
rect 33500 4067 33512 4075
rect 33524 4067 33528 4075
rect 33532 4067 33544 4075
rect 33548 4067 33552 4075
rect 33564 4067 33576 4075
rect 33600 4067 33608 4075
rect 33624 4067 33648 4075
rect 33656 4067 33672 4075
rect 33680 4067 33704 4075
rect 33720 4067 33736 4075
rect 33744 4067 33768 4075
rect 33784 4067 33832 4075
rect 33848 4067 33896 4075
rect 33912 4067 33928 4075
rect 33936 4067 33960 4075
rect 33976 4067 33992 4075
rect 34008 4067 34020 4075
rect 34024 4067 34036 4075
rect 34040 4067 34052 4075
rect 34072 4067 34084 4075
rect 34088 4067 34092 4075
rect 34164 4067 34176 4075
rect 34180 4067 34184 4075
rect 34288 4067 34300 4075
rect 34304 4067 34308 4075
rect 34320 4067 34332 4075
rect 34344 4067 34348 4075
rect 34352 4067 34364 4075
rect 34380 4067 34392 4075
rect 34396 4067 34400 4075
rect 34412 4067 34424 4075
rect 34432 4067 34456 4075
rect 34472 4067 34496 4075
rect 34504 4067 34516 4075
rect 34528 4067 34532 4075
rect 34536 4067 34548 4075
rect 34652 4067 34656 4075
rect 34660 4067 34672 4075
rect 34784 4067 34796 4075
rect 34800 4067 34804 4075
rect 34836 4067 34840 4075
rect 34844 4067 34856 4075
rect 34876 4067 34888 4075
rect 34892 4067 34896 4075
rect 34908 4067 34920 4075
rect 34940 4067 34952 4075
rect 34956 4067 34960 4075
rect 34972 4067 34984 4075
rect 34996 4067 35000 4075
rect 35004 4067 35016 4075
rect 35032 4067 35044 4075
rect 35048 4067 35052 4075
rect 35064 4067 35076 4075
rect 35088 4067 35092 4075
rect 35096 4067 35108 4075
rect 35252 4067 35264 4075
rect 35268 4067 35272 4075
rect 35284 4067 35296 4075
rect 35316 4067 35328 4075
rect 35348 4067 35360 4075
rect 35372 4067 35376 4075
rect 35380 4067 35392 4075
rect 35412 4067 35424 4075
rect 35428 4067 35432 4075
rect 35444 4067 35456 4075
rect 35476 4067 35488 4075
rect 35492 4067 35496 4075
rect 35508 4067 35520 4075
rect 35528 4067 35552 4075
rect 35568 4067 35580 4075
rect 35584 4067 35588 4075
rect 35600 4067 35612 4075
rect 35624 4067 35628 4075
rect 35632 4067 35644 4075
rect 35660 4067 35708 4075
rect 35720 4067 35736 4075
rect 35752 4067 35800 4075
rect 35816 4067 35832 4075
rect 35848 4067 35864 4075
rect 35880 4067 35896 4075
rect 35912 4067 35960 4075
rect 35976 4067 35992 4075
rect 36000 4067 36012 4075
rect 36016 4067 36028 4075
rect 36040 4067 36044 4075
rect 36048 4067 36052 4075
rect 36072 4067 36076 4075
rect 36080 4067 36084 4075
rect 36104 4067 36108 4075
rect 36112 4067 36116 4075
rect 36136 4067 36140 4075
rect 36144 4067 36148 4075
rect 36160 4067 36172 4075
rect 36176 4067 36188 4075
rect 36196 4067 36212 4075
rect 36228 4067 36244 4075
rect 36252 4067 36276 4075
rect 36292 4067 36304 4075
rect 36324 4067 36336 4075
rect 36340 4067 36352 4075
rect 36356 4067 36368 4075
rect 36388 4067 36400 4075
rect 36404 4067 36416 4075
rect 36420 4067 36432 4075
rect 36452 4067 36464 4075
rect 36468 4067 36472 4075
rect 36484 4067 36496 4075
rect 36516 4067 36528 4075
rect 36532 4067 36536 4075
rect 36548 4067 36560 4075
rect 36572 4067 36576 4075
rect 36580 4067 36592 4075
rect 36596 4067 36600 4075
rect 36612 4067 36624 4075
rect 36636 4067 36640 4075
rect 36644 4067 36656 4075
rect 36672 4067 36720 4075
rect 36736 4067 36752 4075
rect 36764 4067 36812 4075
rect 36824 4067 36840 4075
rect 36856 4067 36904 4075
rect 36920 4067 36936 4075
rect 36948 4067 36996 4075
rect 37012 4067 37028 4075
rect 37044 4067 37048 4075
rect 37052 4067 37064 4075
rect 37076 4067 37080 4075
rect 37084 4067 37088 4075
rect 37108 4067 37112 4075
rect 37116 4067 37120 4075
rect 37200 4067 37204 4075
rect 37208 4067 37212 4075
rect 37436 4067 37440 4075
rect 37444 4067 37456 4075
rect 37468 4067 37472 4075
rect 37476 4067 37480 4075
rect 37492 4067 37504 4075
rect 37508 4067 37512 4075
rect 37532 4067 37536 4075
rect 37540 4067 37544 4075
rect 37560 4067 37576 4075
rect 37584 4067 37616 4075
rect 37624 4067 37636 4075
rect 37656 4067 37668 4075
rect 37672 4067 37684 4075
rect 37688 4067 37700 4075
rect 37720 4067 37732 4075
rect 37736 4067 37740 4075
rect 38088 4067 38092 4075
rect 38096 4067 38108 4075
rect 38180 4067 38184 4075
rect 38188 4067 38200 4075
rect 38220 4067 38232 4075
rect 38236 4067 38248 4075
rect 38252 4067 38264 4075
rect 38284 4067 38296 4075
rect 38312 4067 38324 4075
rect 38328 4067 38340 4075
rect 38344 4067 38356 4075
rect 38588 4067 38592 4075
rect 38596 4067 38608 4075
rect 38752 4067 38764 4075
rect 38768 4067 38772 4075
rect 38784 4067 38796 4075
rect 38808 4067 38812 4075
rect 38816 4067 38828 4075
rect 38972 4067 38984 4075
rect 38988 4067 38992 4075
rect 39024 4067 39028 4075
rect 39032 4067 39044 4075
rect 39064 4067 39076 4075
rect 39080 4067 39092 4075
rect 39096 4067 39108 4075
rect 39128 4067 39140 4075
rect 39156 4067 39168 4075
rect 39172 4067 39184 4075
rect 39188 4067 39200 4075
rect 39312 4067 39324 4075
rect 39336 4067 39340 4075
rect 39344 4067 39356 4075
rect 39360 4067 39364 4075
rect 39376 4067 39388 4075
rect 39400 4067 39404 4075
rect 39408 4067 39420 4075
rect 39436 4067 39448 4075
rect 39452 4067 39456 4075
rect 39468 4067 39480 4075
rect 39492 4067 39496 4075
rect 39500 4067 39512 4075
rect 39528 4067 39576 4075
rect 39592 4067 39608 4075
rect 39624 4067 39640 4075
rect 39656 4067 39672 4075
rect 39688 4067 39736 4075
rect 39752 4067 39768 4075
rect 39784 4067 39800 4075
rect 39816 4067 39832 4075
rect 39848 4067 39896 4075
rect 39912 4067 39916 4075
rect 39920 4067 39924 4075
rect 39940 4067 39988 4075
rect 40004 4067 40008 4075
rect 40012 4067 40016 4075
rect 40028 4067 40040 4075
rect 40044 4067 40056 4075
rect 40068 4067 40072 4075
rect 40076 4067 40080 4075
rect 40100 4067 40104 4075
rect 40108 4067 40112 4075
rect 40176 4067 40180 4075
rect 40184 4067 40196 4075
rect 40208 4067 40212 4075
rect 40216 4067 40220 4075
rect 40476 4067 40480 4075
rect 40484 4067 40488 4075
rect 40712 4067 40716 4075
rect 40720 4067 40724 4075
rect 40744 4067 40748 4075
rect 40752 4067 40764 4075
rect 40768 4067 40780 4075
rect 40784 4067 40788 4075
rect 19958 4050 19962 4058
rect 19966 4050 19970 4058
rect 20278 4050 20282 4058
rect 20286 4050 20290 4058
rect 20690 4050 20694 4058
rect 20698 4050 20702 4058
rect 20790 4050 20800 4058
rect 21110 4050 21122 4058
rect 21186 4050 21198 4058
rect 21406 4050 21412 4058
rect 21414 4050 21420 4058
rect 21620 4050 21626 4058
rect 21628 4050 21634 4058
rect 22132 4050 22144 4058
rect 22454 4050 22466 4058
rect 22766 4050 22770 4058
rect 22774 4050 22778 4058
rect 24002 4050 24006 4058
rect 24010 4050 24014 4058
rect 24110 4050 24114 4058
rect 24118 4050 24122 4058
rect 24324 4050 24328 4058
rect 24332 4050 24336 4058
rect 24752 4050 24756 4058
rect 24760 4050 24764 4058
rect 24966 4050 24970 4058
rect 24974 4050 24978 4058
rect 25180 4050 25184 4058
rect 25188 4050 25192 4058
rect 26036 4050 26040 4058
rect 26044 4050 26048 4058
rect 26250 4050 26254 4058
rect 26258 4050 26262 4058
rect 26678 4050 26682 4058
rect 26686 4050 26690 4058
rect 33440 4057 33448 4065
rect 36448 4057 36456 4065
rect 33872 4037 33880 4045
rect 37456 4037 37464 4045
rect 39504 4037 39512 4045
rect 12490 4019 12498 4027
rect 13594 4019 13602 4027
rect 31680 4017 31688 4025
rect 40624 4017 40632 4025
rect 12170 3999 12178 4007
rect 13786 3999 13794 4007
rect 20080 4000 20088 4008
rect 26448 4000 26456 4008
rect 27680 4000 27688 4008
rect 31136 3997 31144 4005
rect 31152 3997 31160 4005
rect 40320 3997 40328 4005
rect 15370 3979 15378 3987
rect 15626 3979 15634 3987
rect 15946 3979 15954 3987
rect 16138 3979 16146 3987
rect 16330 3979 16338 3987
rect 17050 3979 17058 3987
rect 24096 3980 24104 3988
rect 27264 3980 27272 3988
rect 29472 3977 29480 3985
rect 29744 3977 29752 3985
rect 30160 3977 30168 3985
rect 30400 3977 30408 3985
rect 31152 3977 31160 3985
rect 31280 3977 31288 3985
rect 31728 3977 31736 3985
rect 32112 3977 32120 3985
rect 32768 3977 32776 3985
rect 33584 3977 33592 3985
rect 34848 3977 34856 3985
rect 36912 3977 36920 3985
rect 40496 3977 40504 3985
rect 40528 3977 40536 3985
rect 12250 3959 12258 3967
rect 13018 3959 13026 3967
rect 13418 3959 13426 3967
rect 13466 3959 13474 3967
rect 13562 3959 13570 3967
rect 13834 3959 13842 3967
rect 13898 3959 13906 3967
rect 14410 3959 14418 3967
rect 14538 3959 14546 3967
rect 15114 3959 15122 3967
rect 15162 3959 15170 3967
rect 16026 3959 16034 3967
rect 16170 3959 16178 3967
rect 16618 3959 16626 3967
rect 16666 3959 16674 3967
rect 16906 3959 16914 3967
rect 16986 3959 16994 3967
rect 17178 3959 17186 3967
rect 17274 3959 17282 3967
rect 19072 3961 19082 3966
rect 19714 3961 19724 3966
rect 19920 3960 19928 3968
rect 20336 3960 20344 3968
rect 21392 3960 21400 3968
rect 22480 3960 22488 3968
rect 22862 3961 22872 3966
rect 23216 3960 23224 3968
rect 23424 3960 23432 3968
rect 23840 3960 23848 3968
rect 24064 3960 24072 3968
rect 25840 3960 25848 3968
rect 26624 3960 26632 3968
rect 28384 3960 28392 3968
rect 31344 3957 31352 3965
rect 31520 3957 31528 3965
rect 33376 3957 33384 3965
rect 35184 3957 35192 3965
rect 35456 3957 35464 3965
rect 35856 3957 35864 3965
rect 39248 3957 39256 3965
rect 39632 3957 39640 3965
rect 39968 3957 39976 3965
rect 40208 3957 40216 3965
rect 13210 3939 13218 3947
rect 13882 3939 13890 3947
rect 14346 3939 14354 3947
rect 14362 3939 14370 3947
rect 14986 3939 14994 3947
rect 15130 3939 15138 3947
rect 15242 3939 15250 3947
rect 15322 3939 15330 3947
rect 15434 3939 15442 3947
rect 15530 3939 15538 3947
rect 16474 3939 16482 3947
rect 18832 3940 18840 3948
rect 20528 3940 20536 3948
rect 22192 3940 22200 3948
rect 25392 3940 25400 3948
rect 31072 3937 31080 3945
rect 31488 3937 31496 3945
rect 31856 3937 31864 3945
rect 32144 3937 32152 3945
rect 32224 3937 32232 3945
rect 32320 3937 32328 3945
rect 32608 3937 32616 3945
rect 32912 3937 32920 3945
rect 33072 3937 33080 3945
rect 34976 3937 34984 3945
rect 35760 3937 35768 3945
rect 36688 3937 36696 3945
rect 36896 3937 36904 3945
rect 37296 3937 37304 3945
rect 38128 3937 38136 3945
rect 38256 3937 38264 3945
rect 38272 3937 38280 3945
rect 12122 3919 12130 3927
rect 12282 3919 12290 3927
rect 12682 3919 12690 3927
rect 12730 3919 12738 3927
rect 12970 3919 12978 3927
rect 13050 3919 13058 3927
rect 13322 3919 13330 3927
rect 13898 3919 13906 3927
rect 14074 3919 14082 3927
rect 14090 3919 14098 3927
rect 14170 3919 14178 3927
rect 14394 3919 14402 3927
rect 14938 3919 14946 3927
rect 17114 3919 17122 3927
rect 17306 3919 17314 3927
rect 17370 3919 17378 3927
rect 18624 3920 18632 3928
rect 18864 3920 18872 3928
rect 19056 3920 19064 3928
rect 19296 3920 19304 3928
rect 19472 3920 19480 3928
rect 19984 3920 19992 3928
rect 20832 3920 20840 3928
rect 21376 3920 21384 3928
rect 23200 3920 23208 3928
rect 23408 3920 23416 3928
rect 25200 3920 25208 3928
rect 25424 3920 25432 3928
rect 25856 3920 25864 3928
rect 26384 3920 26392 3928
rect 27664 3920 27672 3928
rect 28400 3920 28408 3928
rect 29888 3917 29896 3925
rect 30016 3917 30024 3925
rect 30112 3917 30120 3925
rect 30576 3917 30584 3925
rect 30992 3917 31000 3925
rect 37264 3917 37272 3925
rect 37536 3917 37544 3925
rect 37584 3917 37592 3925
rect 37824 3917 37832 3925
rect 37936 3917 37944 3925
rect 38640 3917 38648 3925
rect 38784 3917 38792 3925
rect 39792 3917 39800 3925
rect 40464 3917 40472 3925
rect 40704 3917 40712 3925
rect 14426 3899 14434 3907
rect 14554 3899 14562 3907
rect 14730 3899 14738 3907
rect 14778 3899 14786 3907
rect 15002 3899 15010 3907
rect 22000 3900 22008 3908
rect 22400 3900 22408 3908
rect 23056 3900 23064 3908
rect 26064 3900 26072 3908
rect 27952 3900 27960 3908
rect 28288 3900 28296 3908
rect 29824 3897 29832 3905
rect 30160 3897 30168 3905
rect 31648 3897 31656 3905
rect 31664 3897 31672 3905
rect 32160 3897 32168 3905
rect 32432 3897 32440 3905
rect 32800 3897 32808 3905
rect 33392 3897 33400 3905
rect 33408 3897 33416 3905
rect 33840 3897 33848 3905
rect 34064 3897 34072 3905
rect 35168 3897 35176 3905
rect 35888 3897 35896 3905
rect 38576 3897 38584 3905
rect 39984 3897 39992 3905
rect 40080 3897 40088 3905
rect 12234 3879 12242 3887
rect 12394 3879 12402 3887
rect 12682 3879 12690 3887
rect 14234 3879 14242 3887
rect 16458 3879 16466 3887
rect 18656 3880 18664 3888
rect 19520 3880 19528 3888
rect 22016 3880 22024 3888
rect 22656 3880 22664 3888
rect 23232 3880 23240 3888
rect 23904 3880 23912 3888
rect 24928 3880 24936 3888
rect 26848 3880 26856 3888
rect 27088 3880 27096 3888
rect 28544 3880 28552 3888
rect 31696 3877 31704 3885
rect 32784 3877 32792 3885
rect 34320 3877 34328 3885
rect 34624 3877 34632 3885
rect 34912 3877 34920 3885
rect 39888 3877 39896 3885
rect 15770 3859 15778 3867
rect 15882 3859 15890 3867
rect 16106 3859 16114 3867
rect 20176 3860 20184 3868
rect 23040 3860 23048 3868
rect 24512 3860 24520 3868
rect 25168 3860 25176 3868
rect 27072 3860 27080 3868
rect 27904 3860 27912 3868
rect 29460 3867 29472 3875
rect 29492 3867 29504 3875
rect 29508 3867 29520 3875
rect 29524 3867 29536 3875
rect 29552 3867 29568 3875
rect 29584 3867 29596 3875
rect 29600 3867 29612 3875
rect 29616 3867 29628 3875
rect 29648 3867 29660 3875
rect 29668 3867 29700 3875
rect 29708 3867 29724 3875
rect 29740 3867 29744 3875
rect 29748 3867 29752 3875
rect 29772 3867 29776 3875
rect 29780 3867 29792 3875
rect 29804 3867 29808 3875
rect 29812 3867 29816 3875
rect 29828 3867 29840 3875
rect 29844 3867 29856 3875
rect 29864 3867 29880 3875
rect 29896 3867 29912 3875
rect 29920 3867 29944 3875
rect 29960 3867 29976 3875
rect 29992 3867 30016 3875
rect 30024 3867 30040 3875
rect 30056 3867 30060 3875
rect 30064 3867 30068 3875
rect 30080 3867 30092 3875
rect 30096 3867 30108 3875
rect 30120 3867 30124 3875
rect 30128 3867 30132 3875
rect 30144 3867 30156 3875
rect 30160 3867 30172 3875
rect 30184 3867 30188 3875
rect 30192 3867 30196 3875
rect 30292 3867 30296 3875
rect 30300 3867 30304 3875
rect 30324 3867 30328 3875
rect 30332 3867 30336 3875
rect 30348 3867 30360 3875
rect 30364 3867 30376 3875
rect 30384 3867 30400 3875
rect 30416 3867 30420 3875
rect 30424 3867 30428 3875
rect 30440 3867 30452 3875
rect 30456 3867 30468 3875
rect 30476 3867 30492 3875
rect 30508 3867 30524 3875
rect 30532 3867 30544 3875
rect 30548 3867 30560 3875
rect 30572 3867 30576 3875
rect 30580 3867 30584 3875
rect 30604 3867 30608 3875
rect 30612 3867 30616 3875
rect 30712 3867 30716 3875
rect 30720 3867 30724 3875
rect 30804 3867 30808 3875
rect 30812 3867 30816 3875
rect 30864 3867 30868 3875
rect 30872 3867 30884 3875
rect 30904 3867 30916 3875
rect 30920 3867 30924 3875
rect 31240 3867 31244 3875
rect 31248 3867 31260 3875
rect 31280 3867 31292 3875
rect 31296 3867 31300 3875
rect 31532 3867 31544 3875
rect 31564 3867 31576 3875
rect 31580 3867 31592 3875
rect 31596 3867 31608 3875
rect 31628 3867 31640 3875
rect 31656 3867 31668 3875
rect 31672 3867 31684 3875
rect 31688 3867 31700 3875
rect 31720 3867 31732 3875
rect 31744 3867 31748 3875
rect 31752 3867 31764 3875
rect 31908 3867 31920 3875
rect 31924 3867 31928 3875
rect 31948 3867 31952 3875
rect 31956 3867 31960 3875
rect 31972 3867 31984 3875
rect 31988 3867 32000 3875
rect 32008 3867 32024 3875
rect 32040 3867 32044 3875
rect 32048 3867 32052 3875
rect 32064 3867 32076 3875
rect 32080 3867 32092 3875
rect 32100 3867 32116 3875
rect 32132 3867 32148 3875
rect 32156 3867 32180 3875
rect 32196 3867 32208 3875
rect 32228 3867 32240 3875
rect 32244 3867 32256 3875
rect 32260 3867 32272 3875
rect 32344 3867 32348 3875
rect 32352 3867 32364 3875
rect 32600 3867 32612 3875
rect 32616 3867 32620 3875
rect 32632 3867 32644 3875
rect 32656 3867 32660 3875
rect 32664 3867 32676 3875
rect 32692 3867 32716 3875
rect 32724 3867 32740 3875
rect 32756 3867 32760 3875
rect 32764 3867 32768 3875
rect 32788 3867 32792 3875
rect 32796 3867 32808 3875
rect 32812 3867 32824 3875
rect 32828 3867 32832 3875
rect 32848 3867 32852 3875
rect 32856 3867 32860 3875
rect 32880 3867 32884 3875
rect 32888 3867 32900 3875
rect 32904 3867 32916 3875
rect 32920 3867 32924 3875
rect 32944 3867 32948 3875
rect 32952 3867 32956 3875
rect 32972 3867 32976 3875
rect 32980 3867 32992 3875
rect 32996 3867 33008 3875
rect 33012 3867 33016 3875
rect 33032 3867 33048 3875
rect 33064 3867 33080 3875
rect 33088 3867 33112 3875
rect 33128 3867 33152 3875
rect 33160 3867 33176 3875
rect 33192 3867 33196 3875
rect 33200 3867 33204 3875
rect 33224 3867 33228 3875
rect 33232 3867 33244 3875
rect 33248 3867 33260 3875
rect 33264 3867 33268 3875
rect 33288 3867 33292 3875
rect 33296 3867 33300 3875
rect 33348 3867 33352 3875
rect 33356 3867 33360 3875
rect 33380 3867 33384 3875
rect 33388 3867 33400 3875
rect 33404 3867 33416 3875
rect 33420 3867 33424 3875
rect 33440 3867 33464 3875
rect 33472 3867 33488 3875
rect 33496 3867 33508 3875
rect 33512 3867 33516 3875
rect 33536 3867 33540 3875
rect 33544 3867 33556 3875
rect 33560 3867 33572 3875
rect 33576 3867 33580 3875
rect 33600 3867 33604 3875
rect 33608 3867 33612 3875
rect 33628 3867 33632 3875
rect 33636 3867 33648 3875
rect 33652 3867 33664 3875
rect 33668 3867 33672 3875
rect 33692 3867 33696 3875
rect 33700 3867 33704 3875
rect 33720 3867 33736 3875
rect 33744 3867 33768 3875
rect 33784 3867 33796 3875
rect 33800 3867 33804 3875
rect 33816 3867 33828 3875
rect 33840 3867 33844 3875
rect 33848 3867 33860 3875
rect 33864 3867 33868 3875
rect 33880 3867 33892 3875
rect 34004 3867 34016 3875
rect 34020 3867 34032 3875
rect 34036 3867 34048 3875
rect 34068 3867 34080 3875
rect 34092 3867 34096 3875
rect 34100 3867 34112 3875
rect 34132 3867 34144 3875
rect 34288 3867 34300 3875
rect 34320 3867 34332 3875
rect 34336 3867 34348 3875
rect 34352 3867 34364 3875
rect 34500 3867 34504 3875
rect 34508 3867 34520 3875
rect 34524 3867 34528 3875
rect 34540 3867 34552 3875
rect 34560 3867 34584 3875
rect 34600 3867 34624 3875
rect 34632 3867 34644 3875
rect 34652 3867 34676 3875
rect 34692 3867 34716 3875
rect 34724 3867 34736 3875
rect 34748 3867 34752 3875
rect 34756 3867 34768 3875
rect 34784 3867 34808 3875
rect 34816 3867 34828 3875
rect 34836 3867 34860 3875
rect 34876 3867 34900 3875
rect 34908 3867 34920 3875
rect 34932 3867 34936 3875
rect 34940 3867 34952 3875
rect 34956 3867 34960 3875
rect 34972 3867 34984 3875
rect 35024 3867 35028 3875
rect 35032 3867 35044 3875
rect 35048 3867 35052 3875
rect 35188 3867 35200 3875
rect 35204 3867 35216 3875
rect 35220 3867 35232 3875
rect 35248 3867 35264 3875
rect 35280 3867 35304 3875
rect 35312 3867 35328 3875
rect 35344 3867 35348 3875
rect 35352 3867 35356 3875
rect 35368 3867 35380 3875
rect 35384 3867 35396 3875
rect 35408 3867 35412 3875
rect 35416 3867 35420 3875
rect 35440 3867 35444 3875
rect 35448 3867 35452 3875
rect 35548 3867 35552 3875
rect 35556 3867 35560 3875
rect 35640 3867 35644 3875
rect 35648 3867 35652 3875
rect 35664 3867 35676 3875
rect 35680 3867 35692 3875
rect 35704 3867 35708 3875
rect 35712 3867 35716 3875
rect 35732 3867 35736 3875
rect 35740 3867 35744 3875
rect 35756 3867 35768 3875
rect 35772 3867 35784 3875
rect 35796 3867 35800 3875
rect 35804 3867 35808 3875
rect 35828 3867 35832 3875
rect 35836 3867 35840 3875
rect 35860 3867 35864 3875
rect 35868 3867 35872 3875
rect 35892 3867 35896 3875
rect 35900 3867 35904 3875
rect 35916 3867 35928 3875
rect 35932 3867 35944 3875
rect 35956 3867 35960 3875
rect 35964 3867 35968 3875
rect 35984 3867 36032 3875
rect 36048 3867 36064 3875
rect 36072 3867 36096 3875
rect 36112 3867 36128 3875
rect 36136 3867 36168 3875
rect 36176 3867 36192 3875
rect 36208 3867 36212 3875
rect 36216 3867 36220 3875
rect 36240 3867 36244 3875
rect 36248 3867 36260 3875
rect 36272 3867 36276 3875
rect 36280 3867 36284 3875
rect 36332 3867 36336 3875
rect 36340 3867 36352 3875
rect 36364 3867 36368 3875
rect 36372 3867 36376 3875
rect 36388 3867 36400 3875
rect 36404 3867 36416 3875
rect 36428 3867 36432 3875
rect 36436 3867 36440 3875
rect 36456 3867 36472 3875
rect 36480 3867 36504 3875
rect 36520 3867 36532 3875
rect 36552 3867 36564 3875
rect 36568 3867 36580 3875
rect 36584 3867 36596 3875
rect 36700 3867 36704 3875
rect 36708 3867 36720 3875
rect 36740 3867 36752 3875
rect 36756 3867 36760 3875
rect 36792 3867 36796 3875
rect 36800 3867 36812 3875
rect 36956 3867 36968 3875
rect 36972 3867 36976 3875
rect 36988 3867 37000 3875
rect 37012 3867 37016 3875
rect 37020 3867 37032 3875
rect 37052 3867 37064 3875
rect 37076 3867 37080 3875
rect 37084 3867 37096 3875
rect 37116 3867 37128 3875
rect 37132 3867 37144 3875
rect 37148 3867 37160 3875
rect 37180 3867 37192 3875
rect 37208 3867 37220 3875
rect 37224 3867 37236 3875
rect 37240 3867 37252 3875
rect 37364 3867 37376 3875
rect 37388 3867 37392 3875
rect 37396 3867 37408 3875
rect 37412 3867 37416 3875
rect 37428 3867 37440 3875
rect 37452 3867 37456 3875
rect 37460 3867 37472 3875
rect 37476 3867 37480 3875
rect 37492 3867 37504 3875
rect 37524 3867 37536 3875
rect 37552 3867 37576 3875
rect 37584 3867 37600 3875
rect 37608 3867 37620 3875
rect 37624 3867 37628 3875
rect 37648 3867 37652 3875
rect 37656 3867 37668 3875
rect 37672 3867 37684 3875
rect 37688 3867 37692 3875
rect 37788 3867 37792 3875
rect 37796 3867 37808 3875
rect 37820 3867 37824 3875
rect 37828 3867 37832 3875
rect 37912 3867 37916 3875
rect 37920 3867 37924 3875
rect 37936 3867 37948 3875
rect 37952 3867 37956 3875
rect 37976 3867 37980 3875
rect 37984 3867 37988 3875
rect 38000 3867 38012 3875
rect 38016 3867 38020 3875
rect 38040 3867 38044 3875
rect 38048 3867 38060 3875
rect 38068 3867 38084 3875
rect 38092 3867 38104 3875
rect 38108 3867 38112 3875
rect 38132 3867 38136 3875
rect 38140 3867 38152 3875
rect 38156 3867 38168 3875
rect 38172 3867 38176 3875
rect 38288 3867 38292 3875
rect 38296 3867 38300 3875
rect 38540 3867 38544 3875
rect 38548 3867 38560 3875
rect 38564 3867 38576 3875
rect 38580 3867 38584 3875
rect 38600 3867 38604 3875
rect 38608 3867 38612 3875
rect 38632 3867 38636 3875
rect 38640 3867 38652 3875
rect 38656 3867 38668 3875
rect 38672 3867 38676 3875
rect 38696 3867 38700 3875
rect 38704 3867 38708 3875
rect 38724 3867 38740 3875
rect 38748 3867 38772 3875
rect 38788 3867 38800 3875
rect 38804 3867 38808 3875
rect 38820 3867 38832 3875
rect 38840 3867 38864 3875
rect 38880 3867 38904 3875
rect 38912 3867 38924 3875
rect 38936 3867 38940 3875
rect 38944 3867 38956 3875
rect 38972 3867 38996 3875
rect 39004 3867 39020 3875
rect 39036 3867 39040 3875
rect 39044 3867 39048 3875
rect 39068 3867 39072 3875
rect 39076 3867 39088 3875
rect 39092 3867 39104 3875
rect 39108 3867 39112 3875
rect 39132 3867 39136 3875
rect 39140 3867 39144 3875
rect 39192 3867 39196 3875
rect 39200 3867 39204 3875
rect 39224 3867 39228 3875
rect 39232 3867 39236 3875
rect 39248 3867 39260 3875
rect 39264 3867 39268 3875
rect 39288 3867 39292 3875
rect 39296 3867 39300 3875
rect 39312 3867 39324 3875
rect 39328 3867 39340 3875
rect 39352 3867 39356 3875
rect 39360 3867 39364 3875
rect 39384 3867 39388 3875
rect 39392 3867 39404 3875
rect 39416 3867 39420 3875
rect 39424 3867 39428 3875
rect 39604 3867 39608 3875
rect 39612 3867 39616 3875
rect 39628 3867 39640 3875
rect 39644 3867 39648 3875
rect 39668 3867 39672 3875
rect 39676 3867 39680 3875
rect 39696 3867 39744 3875
rect 39760 3867 39772 3875
rect 39792 3867 39804 3875
rect 39816 3867 39820 3875
rect 39824 3867 39836 3875
rect 39856 3867 39868 3875
rect 39872 3867 39884 3875
rect 39888 3867 39900 3875
rect 39948 3867 39960 3875
rect 39964 3867 39976 3875
rect 39980 3867 39992 3875
rect 40136 3867 40148 3875
rect 40152 3867 40156 3875
rect 40168 3867 40180 3875
rect 40192 3867 40196 3875
rect 40200 3867 40212 3875
rect 40228 3867 40240 3875
rect 40244 3867 40248 3875
rect 40260 3867 40272 3875
rect 40280 3867 40304 3875
rect 40320 3867 40344 3875
rect 40352 3867 40368 3875
rect 40384 3867 40388 3875
rect 40392 3867 40396 3875
rect 40416 3867 40420 3875
rect 40424 3867 40436 3875
rect 40440 3867 40452 3875
rect 40456 3867 40460 3875
rect 40476 3867 40480 3875
rect 40484 3867 40488 3875
rect 40508 3867 40512 3875
rect 40516 3867 40528 3875
rect 40532 3867 40544 3875
rect 40548 3867 40552 3875
rect 40572 3867 40576 3875
rect 40580 3867 40584 3875
rect 40680 3867 40684 3875
rect 40688 3867 40692 3875
rect 40704 3867 40716 3875
rect 40720 3867 40724 3875
rect 40740 3867 40764 3875
rect 40772 3867 40788 3875
rect 18536 3856 18538 3860
rect 18750 3856 18752 3860
rect 18964 3856 18966 3860
rect 19178 3856 19180 3860
rect 19392 3856 19394 3860
rect 18542 3852 18544 3856
rect 18756 3852 18758 3856
rect 18970 3852 18972 3856
rect 19184 3852 19186 3856
rect 19398 3852 19400 3856
rect 20008 3850 20012 3858
rect 20098 3850 20106 3858
rect 20232 3856 20234 3860
rect 20446 3856 20448 3860
rect 20238 3852 20240 3856
rect 20452 3852 20454 3856
rect 20848 3850 20852 3858
rect 20938 3850 20946 3858
rect 21072 3856 21074 3860
rect 21078 3852 21080 3856
rect 22206 3850 22220 3858
rect 22420 3850 22434 3858
rect 22688 3850 22696 3858
rect 22832 3850 22846 3858
rect 23180 3850 23194 3858
rect 23386 3850 23392 3858
rect 23394 3850 23400 3858
rect 23600 3856 23604 3858
rect 23672 3850 23686 3858
rect 23726 3850 23740 3858
rect 23814 3856 23818 3858
rect 24020 3850 24034 3858
rect 24162 3850 24168 3858
rect 24170 3850 24176 3858
rect 24320 3850 24326 3858
rect 24566 3850 24574 3858
rect 24718 3850 24724 3858
rect 24726 3850 24732 3858
rect 24804 3850 24810 3858
rect 24812 3850 24818 3858
rect 24962 3850 24968 3858
rect 25224 3850 25238 3858
rect 26492 3850 26500 3858
rect 26642 3850 26648 3858
rect 28418 3850 28432 3858
rect 34512 3857 34520 3865
rect 35472 3857 35480 3865
rect 36592 3857 36600 3865
rect 40096 3857 40104 3865
rect 12762 3839 12770 3847
rect 12938 3839 12946 3847
rect 13450 3839 13458 3847
rect 13642 3839 13650 3847
rect 14602 3839 14610 3847
rect 14938 3839 14946 3847
rect 16090 3839 16098 3847
rect 26912 3840 26920 3848
rect 29984 3837 29992 3845
rect 31136 3837 31144 3845
rect 31472 3837 31480 3845
rect 32752 3837 32760 3845
rect 33248 3837 33256 3845
rect 33312 3837 33320 3845
rect 36128 3837 36136 3845
rect 36656 3837 36664 3845
rect 36784 3837 36792 3845
rect 37200 3837 37208 3845
rect 37504 3837 37512 3845
rect 37552 3837 37560 3845
rect 37664 3837 37672 3845
rect 38544 3837 38552 3845
rect 38976 3837 38984 3845
rect 39696 3837 39704 3845
rect 39872 3837 39880 3845
rect 40192 3837 40200 3845
rect 40256 3837 40264 3845
rect 40688 3837 40696 3845
rect 13706 3819 13714 3827
rect 13770 3819 13778 3827
rect 16858 3819 16866 3827
rect 17322 3819 17330 3827
rect 18464 3820 18472 3828
rect 21024 3820 21032 3828
rect 22512 3820 22520 3828
rect 22816 3820 22824 3828
rect 23552 3820 23560 3828
rect 24576 3820 24584 3828
rect 25648 3820 25656 3828
rect 26384 3820 26392 3828
rect 26400 3820 26408 3828
rect 27520 3820 27528 3828
rect 29600 3817 29608 3825
rect 37232 3817 37240 3825
rect 37744 3817 37752 3825
rect 37952 3817 37960 3825
rect 39712 3817 39720 3825
rect 40080 3817 40088 3825
rect 40224 3817 40232 3825
rect 40400 3817 40408 3825
rect 40592 3817 40600 3825
rect 12874 3799 12882 3807
rect 14554 3799 14562 3807
rect 14682 3799 14690 3807
rect 14746 3799 14754 3807
rect 14858 3799 14866 3807
rect 14890 3799 14898 3807
rect 15018 3799 15026 3807
rect 15338 3799 15346 3807
rect 15370 3799 15378 3807
rect 15562 3799 15570 3807
rect 15722 3799 15730 3807
rect 16282 3799 16290 3807
rect 16426 3799 16434 3807
rect 16714 3799 16722 3807
rect 17434 3799 17442 3807
rect 17498 3799 17506 3807
rect 18864 3800 18872 3808
rect 20352 3800 20360 3808
rect 21232 3800 21240 3808
rect 29904 3797 29912 3805
rect 31216 3797 31224 3805
rect 31600 3797 31608 3805
rect 32160 3797 32168 3805
rect 32304 3797 32312 3805
rect 32368 3797 32376 3805
rect 32416 3797 32424 3805
rect 33536 3797 33544 3805
rect 33584 3797 33592 3805
rect 33824 3797 33832 3805
rect 33920 3797 33928 3805
rect 33936 3797 33944 3805
rect 34096 3797 34104 3805
rect 34256 3797 34264 3805
rect 34576 3797 34584 3805
rect 34848 3797 34856 3805
rect 35408 3797 35416 3805
rect 35936 3797 35944 3805
rect 36016 3797 36024 3805
rect 36560 3797 36568 3805
rect 36640 3797 36648 3805
rect 36912 3797 36920 3805
rect 37856 3797 37864 3805
rect 38496 3797 38504 3805
rect 39792 3797 39800 3805
rect 40048 3797 40056 3805
rect 40624 3797 40632 3805
rect 12458 3779 12466 3787
rect 12474 3779 12482 3787
rect 13322 3779 13330 3787
rect 13658 3779 13666 3787
rect 13834 3779 13842 3787
rect 14890 3779 14898 3787
rect 15850 3779 15858 3787
rect 16234 3779 16242 3787
rect 16298 3779 16306 3787
rect 16314 3779 16322 3787
rect 16938 3779 16946 3787
rect 19488 3780 19496 3788
rect 20336 3780 20344 3788
rect 21168 3780 21176 3788
rect 21584 3780 21592 3788
rect 21680 3780 21688 3788
rect 22016 3780 22024 3788
rect 23072 3780 23080 3788
rect 24208 3780 24216 3788
rect 24528 3780 24536 3788
rect 25744 3780 25752 3788
rect 25888 3780 25896 3788
rect 26208 3780 26216 3788
rect 26448 3780 26456 3788
rect 26912 3780 26920 3788
rect 27584 3780 27592 3788
rect 27920 3780 27928 3788
rect 27952 3780 27960 3788
rect 28240 3780 28248 3788
rect 29600 3777 29608 3785
rect 29744 3777 29752 3785
rect 30832 3777 30840 3785
rect 31072 3777 31080 3785
rect 31408 3777 31416 3785
rect 31744 3777 31752 3785
rect 31920 3777 31928 3785
rect 31936 3777 31944 3785
rect 32544 3777 32552 3785
rect 32736 3777 32744 3785
rect 32768 3777 32776 3785
rect 33008 3777 33016 3785
rect 33056 3777 33064 3785
rect 36928 3777 36936 3785
rect 39168 3777 39176 3785
rect 14602 3759 14610 3767
rect 16794 3759 16802 3767
rect 16906 3759 16914 3767
rect 17146 3759 17154 3767
rect 26048 3760 26056 3768
rect 28384 3760 28392 3768
rect 30768 3757 30776 3765
rect 32048 3757 32056 3765
rect 32432 3757 32440 3765
rect 33168 3757 33176 3765
rect 33360 3757 33368 3765
rect 33456 3757 33464 3765
rect 33600 3757 33608 3765
rect 33872 3757 33880 3765
rect 34240 3757 34248 3765
rect 34560 3757 34568 3765
rect 34752 3757 34760 3765
rect 34800 3757 34808 3765
rect 34864 3757 34872 3765
rect 35520 3757 35528 3765
rect 35616 3757 35624 3765
rect 35952 3757 35960 3765
rect 36048 3757 36056 3765
rect 36432 3757 36440 3765
rect 36720 3757 36728 3765
rect 37168 3757 37176 3765
rect 37872 3757 37880 3765
rect 39216 3757 39224 3765
rect 39568 3757 39576 3765
rect 40096 3757 40104 3765
rect 40304 3757 40312 3765
rect 40480 3757 40488 3765
rect 40656 3757 40664 3765
rect 19088 3748 19092 3753
rect 24184 3748 24188 3753
rect 27588 3748 27597 3753
rect 12378 3739 12386 3747
rect 12634 3739 12642 3747
rect 13130 3739 13138 3747
rect 13370 3739 13378 3747
rect 14186 3739 14194 3747
rect 14522 3739 14530 3747
rect 15050 3739 15058 3747
rect 15498 3739 15506 3747
rect 15578 3739 15586 3747
rect 15658 3739 15666 3747
rect 15706 3739 15714 3747
rect 15754 3739 15762 3747
rect 15994 3739 16002 3747
rect 16106 3739 16114 3747
rect 16202 3739 16210 3747
rect 16346 3739 16354 3747
rect 16362 3739 16370 3747
rect 16618 3739 16626 3747
rect 16666 3739 16674 3747
rect 16778 3739 16786 3747
rect 17210 3739 17218 3747
rect 17290 3739 17298 3747
rect 17370 3739 17378 3747
rect 17418 3739 17426 3747
rect 17498 3739 17506 3747
rect 18864 3740 18872 3748
rect 19504 3740 19512 3748
rect 20128 3740 20136 3748
rect 20352 3740 20360 3748
rect 23152 3740 23160 3748
rect 24768 3740 24776 3748
rect 25168 3740 25176 3748
rect 25792 3740 25800 3748
rect 26512 3740 26520 3748
rect 26704 3740 26712 3748
rect 28224 3740 28232 3748
rect 14410 3719 14418 3727
rect 15306 3719 15314 3727
rect 17050 3719 17058 3727
rect 18848 3720 18856 3728
rect 19712 3720 19720 3728
rect 25872 3720 25880 3728
rect 27936 3720 27944 3728
rect 37712 3717 37720 3725
rect 38624 3717 38632 3725
rect 13306 3699 13314 3707
rect 14170 3699 14178 3707
rect 23504 3700 23512 3708
rect 28016 3700 28024 3708
rect 34752 3697 34760 3705
rect 14010 3679 14018 3687
rect 15194 3679 15202 3687
rect 24352 3680 24360 3688
rect 26496 3680 26504 3688
rect 29556 3667 29568 3675
rect 29808 3667 29820 3675
rect 29832 3667 29836 3675
rect 29840 3667 29852 3675
rect 29856 3667 29860 3675
rect 29964 3667 29976 3675
rect 29996 3667 30008 3675
rect 30012 3667 30016 3675
rect 30028 3667 30040 3675
rect 30056 3667 30072 3675
rect 30080 3667 30112 3675
rect 30120 3667 30136 3675
rect 30144 3667 30168 3675
rect 30184 3667 30200 3675
rect 30208 3667 30232 3675
rect 30248 3667 30272 3675
rect 30280 3667 30296 3675
rect 30312 3667 30316 3675
rect 30320 3667 30324 3675
rect 30344 3667 30348 3675
rect 30352 3667 30364 3675
rect 30368 3667 30380 3675
rect 30384 3667 30388 3675
rect 30404 3667 30420 3675
rect 30436 3667 30440 3675
rect 30444 3667 30456 3675
rect 30460 3667 30472 3675
rect 30476 3667 30480 3675
rect 30528 3667 30532 3675
rect 30536 3667 30548 3675
rect 30552 3667 30564 3675
rect 30568 3667 30572 3675
rect 30620 3667 30624 3675
rect 30628 3667 30640 3675
rect 30644 3667 30656 3675
rect 30660 3667 30664 3675
rect 30684 3667 30688 3675
rect 30692 3667 30696 3675
rect 30712 3667 30716 3675
rect 30720 3667 30732 3675
rect 30736 3667 30748 3675
rect 30752 3667 30756 3675
rect 30804 3667 30808 3675
rect 30812 3667 30824 3675
rect 30828 3667 30840 3675
rect 30844 3667 30848 3675
rect 30864 3667 30880 3675
rect 30896 3667 30900 3675
rect 30904 3667 30916 3675
rect 30920 3667 30932 3675
rect 30936 3667 30940 3675
rect 30960 3667 30964 3675
rect 30968 3667 30972 3675
rect 31068 3667 31072 3675
rect 31076 3667 31080 3675
rect 31092 3667 31104 3675
rect 31108 3667 31112 3675
rect 31132 3667 31136 3675
rect 31140 3667 31152 3675
rect 31156 3667 31168 3675
rect 31172 3667 31176 3675
rect 31192 3667 31196 3675
rect 31200 3667 31204 3675
rect 31224 3667 31228 3675
rect 31232 3667 31244 3675
rect 31248 3667 31260 3675
rect 31264 3667 31268 3675
rect 31284 3667 31300 3675
rect 31316 3667 31320 3675
rect 31324 3667 31336 3675
rect 31340 3667 31352 3675
rect 31356 3667 31360 3675
rect 31376 3667 31392 3675
rect 31408 3667 31424 3675
rect 31432 3667 31456 3675
rect 31472 3667 31496 3675
rect 31504 3667 31516 3675
rect 31524 3667 31548 3675
rect 31564 3667 31588 3675
rect 31596 3667 31608 3675
rect 31620 3667 31624 3675
rect 31628 3667 31640 3675
rect 31656 3667 31668 3675
rect 31672 3667 31676 3675
rect 31688 3667 31700 3675
rect 31712 3667 31716 3675
rect 31720 3667 31732 3675
rect 31876 3667 31888 3675
rect 31892 3667 31896 3675
rect 31908 3667 31920 3675
rect 31936 3667 31952 3675
rect 31968 3667 32016 3675
rect 32028 3667 32044 3675
rect 32060 3667 32108 3675
rect 32124 3667 32128 3675
rect 32132 3667 32136 3675
rect 32156 3667 32160 3675
rect 32164 3667 32176 3675
rect 32188 3667 32192 3675
rect 32196 3667 32200 3675
rect 32296 3667 32300 3675
rect 32304 3667 32316 3675
rect 32328 3667 32332 3675
rect 32336 3667 32340 3675
rect 32388 3667 32392 3675
rect 32396 3667 32408 3675
rect 32420 3667 32424 3675
rect 32428 3667 32432 3675
rect 32444 3667 32456 3675
rect 32460 3667 32464 3675
rect 32512 3667 32516 3675
rect 32520 3667 32524 3675
rect 32536 3667 32548 3675
rect 32552 3667 32556 3675
rect 32572 3667 32588 3675
rect 32604 3667 32620 3675
rect 32628 3667 32660 3675
rect 32668 3667 32680 3675
rect 32700 3667 32712 3675
rect 32724 3667 32728 3675
rect 32732 3667 32744 3675
rect 32764 3667 32776 3675
rect 32788 3667 32792 3675
rect 32796 3667 32808 3675
rect 32812 3667 32816 3675
rect 32828 3667 32840 3675
rect 32848 3667 32872 3675
rect 32888 3667 32912 3675
rect 32920 3667 32936 3675
rect 32952 3667 32968 3675
rect 32984 3667 32988 3675
rect 32992 3667 33004 3675
rect 33008 3667 33020 3675
rect 33024 3667 33028 3675
rect 33332 3667 33336 3675
rect 33340 3667 33344 3675
rect 33440 3667 33444 3675
rect 33448 3667 33452 3675
rect 33628 3667 33632 3675
rect 33636 3667 33648 3675
rect 33652 3667 33664 3675
rect 33668 3667 33672 3675
rect 33692 3667 33696 3675
rect 33700 3667 33712 3675
rect 33720 3667 33736 3675
rect 33744 3667 33776 3675
rect 33784 3667 33796 3675
rect 33816 3667 33828 3675
rect 33840 3667 33844 3675
rect 33848 3667 33860 3675
rect 33880 3667 33892 3675
rect 33996 3667 34000 3675
rect 34004 3667 34016 3675
rect 34020 3667 34024 3675
rect 34036 3667 34048 3675
rect 34068 3667 34080 3675
rect 34100 3667 34112 3675
rect 34132 3667 34144 3675
rect 34156 3667 34160 3675
rect 34164 3667 34176 3675
rect 34180 3667 34184 3675
rect 34196 3667 34208 3675
rect 34288 3667 34300 3675
rect 34312 3667 34316 3675
rect 34320 3667 34332 3675
rect 34336 3667 34340 3675
rect 34352 3667 34364 3675
rect 34384 3667 34396 3675
rect 34416 3667 34428 3675
rect 34448 3667 34460 3675
rect 34472 3667 34476 3675
rect 34480 3667 34492 3675
rect 34496 3667 34500 3675
rect 34512 3667 34524 3675
rect 34544 3667 34556 3675
rect 34560 3667 34564 3675
rect 34576 3667 34588 3675
rect 34608 3667 34620 3675
rect 34628 3667 34660 3675
rect 34668 3667 34680 3675
rect 34700 3667 34712 3675
rect 34720 3667 34752 3675
rect 34760 3667 34776 3675
rect 34784 3667 34808 3675
rect 34824 3667 34828 3675
rect 34832 3667 34844 3675
rect 34852 3667 34868 3675
rect 34876 3667 34900 3675
rect 34912 3667 34936 3675
rect 34944 3667 34960 3675
rect 34968 3667 34992 3675
rect 35008 3667 35012 3675
rect 35016 3667 35028 3675
rect 35036 3667 35052 3675
rect 35060 3667 35072 3675
rect 35076 3667 35080 3675
rect 35100 3667 35104 3675
rect 35108 3667 35120 3675
rect 35132 3667 35136 3675
rect 35140 3667 35144 3675
rect 35164 3667 35168 3675
rect 35172 3667 35176 3675
rect 35240 3667 35244 3675
rect 35248 3667 35252 3675
rect 35272 3667 35276 3675
rect 35280 3667 35292 3675
rect 35296 3667 35308 3675
rect 35312 3667 35316 3675
rect 35332 3667 35356 3675
rect 35364 3667 35380 3675
rect 35388 3667 35412 3675
rect 35428 3667 35444 3675
rect 35460 3667 35472 3675
rect 35484 3667 35488 3675
rect 35492 3667 35504 3675
rect 35508 3667 35512 3675
rect 35524 3667 35536 3675
rect 35552 3667 35564 3675
rect 35576 3667 35580 3675
rect 35584 3667 35596 3675
rect 35600 3667 35604 3675
rect 35616 3667 35628 3675
rect 35740 3667 35752 3675
rect 35756 3667 35760 3675
rect 35772 3667 35784 3675
rect 35804 3667 35816 3675
rect 35828 3667 35832 3675
rect 35836 3667 35848 3675
rect 35868 3667 35880 3675
rect 35892 3667 35896 3675
rect 35900 3667 35912 3675
rect 35916 3667 35920 3675
rect 35932 3667 35944 3675
rect 35964 3667 35976 3675
rect 36000 3667 36016 3675
rect 36024 3667 36040 3675
rect 36048 3667 36080 3675
rect 36088 3667 36104 3675
rect 36120 3667 36144 3675
rect 36152 3667 36168 3675
rect 36184 3667 36200 3675
rect 36208 3667 36232 3675
rect 36248 3667 36260 3675
rect 36280 3667 36292 3675
rect 36296 3667 36308 3675
rect 36312 3667 36324 3675
rect 36340 3667 36356 3675
rect 36364 3667 36396 3675
rect 36404 3667 36416 3675
rect 36436 3667 36448 3675
rect 36456 3667 36488 3675
rect 36496 3667 36508 3675
rect 36524 3667 36540 3675
rect 36548 3667 36580 3675
rect 36588 3667 36604 3675
rect 36616 3667 36632 3675
rect 36640 3667 36672 3675
rect 36680 3667 36692 3675
rect 36708 3667 36724 3675
rect 36732 3667 36764 3675
rect 36772 3667 36788 3675
rect 36800 3667 36816 3675
rect 36824 3667 36856 3675
rect 36864 3667 36880 3675
rect 36896 3667 36912 3675
rect 36928 3667 36944 3675
rect 36960 3667 36976 3675
rect 36984 3667 37016 3675
rect 37024 3667 37040 3675
rect 37048 3667 37080 3675
rect 37088 3667 37100 3675
rect 37120 3667 37132 3675
rect 37136 3667 37148 3675
rect 37152 3667 37164 3675
rect 37184 3667 37196 3675
rect 37212 3667 37224 3675
rect 37228 3667 37240 3675
rect 37244 3667 37256 3675
rect 37272 3667 37284 3675
rect 37304 3667 37316 3675
rect 37320 3667 37332 3675
rect 37336 3667 37348 3675
rect 37364 3667 37380 3675
rect 37396 3667 37420 3675
rect 37428 3667 37444 3675
rect 37460 3667 37508 3675
rect 37524 3667 37540 3675
rect 37552 3667 37600 3675
rect 37612 3667 37628 3675
rect 37644 3667 37692 3675
rect 37704 3667 37720 3675
rect 37736 3667 37784 3675
rect 37800 3667 37804 3675
rect 37808 3667 37812 3675
rect 37828 3667 37876 3675
rect 37892 3667 37904 3675
rect 37920 3667 37968 3675
rect 37984 3667 37996 3675
rect 38000 3667 38004 3675
rect 38016 3667 38028 3675
rect 38040 3667 38044 3675
rect 38048 3667 38060 3675
rect 38076 3667 38100 3675
rect 38108 3667 38120 3675
rect 38132 3667 38136 3675
rect 38140 3667 38152 3675
rect 38156 3667 38160 3675
rect 38172 3667 38184 3675
rect 38196 3667 38200 3675
rect 38204 3667 38216 3675
rect 38220 3667 38224 3675
rect 38236 3667 38248 3675
rect 38288 3667 38292 3675
rect 38296 3667 38308 3675
rect 38312 3667 38316 3675
rect 38328 3667 38340 3675
rect 38352 3667 38356 3675
rect 38360 3667 38372 3675
rect 38392 3667 38400 3675
rect 38424 3667 38436 3675
rect 38456 3667 38468 3675
rect 38472 3667 38476 3675
rect 38488 3667 38500 3675
rect 38512 3667 38516 3675
rect 38520 3667 38532 3675
rect 38548 3667 38596 3675
rect 38612 3667 38616 3675
rect 38620 3667 38624 3675
rect 38644 3667 38648 3675
rect 38652 3667 38664 3675
rect 38676 3667 38680 3675
rect 38684 3667 38688 3675
rect 38708 3667 38712 3675
rect 38716 3667 38720 3675
rect 38784 3667 38788 3675
rect 38792 3667 38804 3675
rect 38816 3667 38820 3675
rect 38824 3667 38828 3675
rect 38840 3667 38852 3675
rect 38856 3667 38860 3675
rect 38908 3667 38912 3675
rect 38916 3667 38920 3675
rect 38932 3667 38944 3675
rect 38948 3667 38952 3675
rect 38972 3667 38976 3675
rect 38980 3667 38984 3675
rect 39004 3667 39008 3675
rect 39012 3667 39016 3675
rect 39036 3667 39040 3675
rect 39044 3667 39056 3675
rect 39068 3667 39072 3675
rect 39076 3667 39080 3675
rect 39092 3667 39104 3675
rect 39108 3667 39112 3675
rect 39192 3667 39196 3675
rect 39200 3667 39212 3675
rect 39224 3667 39228 3675
rect 39232 3667 39236 3675
rect 39332 3667 39336 3675
rect 39340 3667 39344 3675
rect 39364 3667 39368 3675
rect 39372 3667 39376 3675
rect 39388 3667 39400 3675
rect 39404 3667 39408 3675
rect 39428 3667 39432 3675
rect 39436 3667 39440 3675
rect 39456 3667 39504 3675
rect 39520 3667 39544 3675
rect 39552 3667 39564 3675
rect 39576 3667 39580 3675
rect 39584 3667 39596 3675
rect 39612 3667 39624 3675
rect 39628 3667 39632 3675
rect 39644 3667 39656 3675
rect 39668 3667 39672 3675
rect 39676 3667 39688 3675
rect 39704 3667 39752 3675
rect 39764 3667 39780 3675
rect 39796 3667 39844 3675
rect 39860 3667 39884 3675
rect 39892 3667 39904 3675
rect 39912 3667 39936 3675
rect 39952 3667 39964 3675
rect 39968 3667 39972 3675
rect 39984 3667 39996 3675
rect 40004 3667 40028 3675
rect 40044 3667 40056 3675
rect 40060 3667 40064 3675
rect 40076 3667 40088 3675
rect 40100 3667 40104 3675
rect 40108 3667 40120 3675
rect 40136 3667 40160 3675
rect 40168 3667 40180 3675
rect 40192 3667 40196 3675
rect 40200 3667 40212 3675
rect 40228 3667 40240 3675
rect 40244 3667 40248 3675
rect 40260 3667 40272 3675
rect 40280 3667 40304 3675
rect 40320 3667 40368 3675
rect 40384 3667 40388 3675
rect 40392 3667 40396 3675
rect 40412 3667 40460 3675
rect 40472 3667 40488 3675
rect 40504 3667 40552 3675
rect 40568 3667 40580 3675
rect 40596 3667 40644 3675
rect 40660 3667 40672 3675
rect 40688 3667 40736 3675
rect 40752 3667 40756 3675
rect 40760 3667 40764 3675
rect 40776 3667 40788 3675
rect 40792 3667 40800 3675
rect 8018 3653 8026 3661
rect 13178 3659 13186 3667
rect 17258 3659 17266 3667
rect 20294 3650 20298 3658
rect 20302 3650 20306 3658
rect 20912 3650 20924 3658
rect 21538 3650 21550 3658
rect 21614 3650 21626 3658
rect 21966 3650 21978 3658
rect 22042 3650 22054 3658
rect 22180 3650 22192 3658
rect 22256 3650 22268 3658
rect 22476 3650 22482 3658
rect 22484 3650 22490 3658
rect 22690 3650 22696 3658
rect 22698 3650 22704 3658
rect 23094 3650 23108 3658
rect 23400 3650 23414 3658
rect 24042 3650 24056 3658
rect 24890 3650 24896 3658
rect 24898 3650 24904 3658
rect 25112 3650 25124 3658
rect 25188 3650 25200 3658
rect 25852 3650 25858 3658
rect 25860 3650 25866 3658
rect 25928 3650 25934 3658
rect 25936 3650 25942 3658
rect 26174 3650 26178 3658
rect 26182 3650 26186 3658
rect 26250 3650 26254 3658
rect 26258 3650 26262 3658
rect 26494 3650 26500 3658
rect 26502 3650 26508 3658
rect 26570 3650 26576 3658
rect 26578 3650 26584 3658
rect 27022 3650 27034 3658
rect 27098 3650 27110 3658
rect 27556 3650 27570 3658
rect 27632 3650 27646 3658
rect 27878 3650 27890 3658
rect 27954 3650 27966 3658
rect 28198 3650 28212 3658
rect 28274 3650 28288 3658
rect 18480 3640 18488 3648
rect 24032 3640 24040 3648
rect 35600 3637 35608 3645
rect 39264 3637 39272 3645
rect 39424 3637 39432 3645
rect 6786 3613 6794 3621
rect 6898 3613 6906 3621
rect 12698 3619 12706 3627
rect 13962 3619 13970 3627
rect 31152 3617 31160 3625
rect 35296 3617 35304 3625
rect 37168 3617 37176 3625
rect 38288 3617 38296 3625
rect 38784 3617 38792 3625
rect 39136 3617 39144 3625
rect 39840 3617 39848 3625
rect 6482 3593 6490 3601
rect 6674 3593 6682 3601
rect 7778 3593 7786 3601
rect 14138 3599 14146 3607
rect 14538 3599 14546 3607
rect 16410 3599 16418 3607
rect 25296 3600 25304 3608
rect 27312 3600 27320 3608
rect 31536 3597 31544 3605
rect 6034 3573 6042 3581
rect 8178 3573 8186 3581
rect 8242 3573 8250 3581
rect 12506 3579 12514 3587
rect 12762 3579 12770 3587
rect 15066 3579 15074 3587
rect 15242 3579 15250 3587
rect 15370 3579 15378 3587
rect 15466 3579 15474 3587
rect 15946 3579 15954 3587
rect 15994 3579 16002 3587
rect 16218 3579 16226 3587
rect 16394 3579 16402 3587
rect 17434 3579 17442 3587
rect 19280 3580 19288 3588
rect 24224 3580 24232 3588
rect 24336 3580 24344 3588
rect 24416 3580 24424 3588
rect 24432 3580 24440 3588
rect 24928 3580 24936 3588
rect 28080 3580 28088 3588
rect 29984 3577 29992 3585
rect 30400 3577 30408 3585
rect 31312 3577 31320 3585
rect 32032 3577 32040 3585
rect 33424 3577 33432 3585
rect 33504 3577 33512 3585
rect 36368 3577 36376 3585
rect 36416 3577 36424 3585
rect 36576 3577 36584 3585
rect 36688 3577 36696 3585
rect 39968 3577 39976 3585
rect 40496 3577 40504 3585
rect 40672 3577 40680 3585
rect 6050 3553 6058 3561
rect 7666 3553 7674 3561
rect 7730 3553 7738 3561
rect 7826 3553 7834 3561
rect 7874 3553 7882 3561
rect 7938 3553 7946 3561
rect 8386 3553 8394 3561
rect 8450 3553 8458 3561
rect 8498 3553 8506 3561
rect 8642 3553 8650 3561
rect 9122 3553 9130 3561
rect 9186 3553 9194 3561
rect 10098 3553 10106 3561
rect 10130 3553 10138 3561
rect 10178 3553 10186 3561
rect 12282 3559 12290 3567
rect 12826 3559 12834 3567
rect 13354 3559 13362 3567
rect 14330 3559 14338 3567
rect 14442 3559 14450 3567
rect 14730 3559 14738 3567
rect 14778 3559 14786 3567
rect 14986 3559 14994 3567
rect 15050 3559 15058 3567
rect 16074 3559 16082 3567
rect 16106 3559 16114 3567
rect 16234 3559 16242 3567
rect 16266 3559 16274 3567
rect 16282 3559 16290 3567
rect 16442 3559 16450 3567
rect 16490 3559 16498 3567
rect 16714 3559 16722 3567
rect 16794 3559 16802 3567
rect 17066 3559 17074 3567
rect 17162 3559 17170 3567
rect 17242 3559 17250 3567
rect 17306 3559 17314 3567
rect 17370 3559 17378 3567
rect 17514 3559 17522 3567
rect 19072 3561 19082 3566
rect 19456 3560 19464 3568
rect 20080 3560 20088 3568
rect 20288 3560 20296 3568
rect 21298 3561 21308 3566
rect 21552 3560 21560 3568
rect 21984 3560 21992 3568
rect 22816 3560 22824 3568
rect 23424 3560 23432 3568
rect 23952 3560 23960 3568
rect 24064 3560 24072 3568
rect 25936 3560 25944 3568
rect 26560 3560 26568 3568
rect 27248 3560 27256 3568
rect 28256 3560 28264 3568
rect 36912 3557 36920 3565
rect 37008 3557 37016 3565
rect 37248 3557 37256 3565
rect 37280 3557 37288 3565
rect 6930 3533 6938 3541
rect 6962 3533 6970 3541
rect 6978 3533 6986 3541
rect 7154 3533 7162 3541
rect 10290 3533 10298 3541
rect 10434 3533 10442 3541
rect 10530 3533 10538 3541
rect 10546 3533 10554 3541
rect 13802 3539 13810 3547
rect 14058 3539 14066 3547
rect 15642 3539 15650 3547
rect 16010 3539 16018 3547
rect 17418 3539 17426 3547
rect 21472 3540 21480 3548
rect 22752 3540 22760 3548
rect 22832 3540 22840 3548
rect 22992 3540 23000 3548
rect 28080 3540 28088 3548
rect 28240 3540 28248 3548
rect 30080 3537 30088 3545
rect 30528 3537 30536 3545
rect 30608 3537 30616 3545
rect 31024 3537 31032 3545
rect 31232 3537 31240 3545
rect 31328 3537 31336 3545
rect 31824 3537 31832 3545
rect 32064 3537 32072 3545
rect 33248 3537 33256 3545
rect 34176 3537 34184 3545
rect 34992 3537 35000 3545
rect 35104 3537 35112 3545
rect 35984 3537 35992 3545
rect 36112 3537 36120 3545
rect 36432 3537 36440 3545
rect 36752 3537 36760 3545
rect 37504 3537 37512 3545
rect 38016 3537 38024 3545
rect 38816 3537 38824 3545
rect 39376 3537 39384 3545
rect 39472 3537 39480 3545
rect 39984 3537 39992 3545
rect 40608 3537 40616 3545
rect 5874 3513 5882 3521
rect 6066 3513 6074 3521
rect 6226 3513 6234 3521
rect 6434 3513 6442 3521
rect 7058 3513 7066 3521
rect 7106 3513 7114 3521
rect 7570 3513 7578 3521
rect 9170 3513 9178 3521
rect 9522 3513 9530 3521
rect 9666 3513 9674 3521
rect 9682 3513 9690 3521
rect 9698 3513 9706 3521
rect 10018 3513 10026 3521
rect 10722 3513 10730 3521
rect 10850 3513 10858 3521
rect 12010 3519 12018 3527
rect 12186 3519 12194 3527
rect 12426 3519 12434 3527
rect 13258 3519 13266 3527
rect 13338 3519 13346 3527
rect 14810 3519 14818 3527
rect 15114 3519 15122 3527
rect 17130 3519 17138 3527
rect 17146 3519 17154 3527
rect 17306 3519 17314 3527
rect 19056 3520 19064 3528
rect 19152 3520 19160 3528
rect 19904 3520 19912 3528
rect 20368 3520 20376 3528
rect 22208 3520 22216 3528
rect 22560 3520 22568 3528
rect 22736 3520 22744 3528
rect 23184 3520 23192 3528
rect 23616 3520 23624 3528
rect 23648 3520 23656 3528
rect 24400 3520 24408 3528
rect 24432 3520 24440 3528
rect 25904 3520 25912 3528
rect 26224 3520 26232 3528
rect 26400 3520 26408 3528
rect 26544 3520 26552 3528
rect 27264 3520 27272 3528
rect 27904 3520 27912 3528
rect 28336 3520 28344 3528
rect 29488 3517 29496 3525
rect 29904 3517 29912 3525
rect 30096 3517 30104 3525
rect 30432 3517 30440 3525
rect 33632 3517 33640 3525
rect 33728 3517 33736 3525
rect 33760 3517 33768 3525
rect 33952 3517 33960 3525
rect 33984 3517 33992 3525
rect 34240 3517 34248 3525
rect 34544 3517 34552 3525
rect 34560 3517 34568 3525
rect 34608 3517 34616 3525
rect 34624 3517 34632 3525
rect 34736 3517 34744 3525
rect 35456 3517 35464 3525
rect 35760 3517 35768 3525
rect 38688 3517 38696 3525
rect 38864 3517 38872 3525
rect 39184 3517 39192 3525
rect 39712 3517 39720 3525
rect 5938 3493 5946 3501
rect 5954 3493 5962 3501
rect 6498 3493 6506 3501
rect 6546 3493 6554 3501
rect 6642 3493 6650 3501
rect 6658 3493 6666 3501
rect 6802 3493 6810 3501
rect 6866 3493 6874 3501
rect 6914 3493 6922 3501
rect 7282 3493 7290 3501
rect 7346 3493 7354 3501
rect 7426 3493 7434 3501
rect 7794 3493 7802 3501
rect 7874 3493 7882 3501
rect 7938 3493 7946 3501
rect 8034 3493 8042 3501
rect 8210 3493 8218 3501
rect 8434 3493 8442 3501
rect 9154 3493 9162 3501
rect 9234 3493 9242 3501
rect 9250 3493 9258 3501
rect 9954 3493 9962 3501
rect 10274 3493 10282 3501
rect 10386 3493 10394 3501
rect 10418 3493 10426 3501
rect 10674 3493 10682 3501
rect 10882 3493 10890 3501
rect 12234 3499 12242 3507
rect 14282 3499 14290 3507
rect 14810 3499 14818 3507
rect 14938 3499 14946 3507
rect 15818 3499 15826 3507
rect 15834 3499 15842 3507
rect 15898 3499 15906 3507
rect 16074 3499 16082 3507
rect 16154 3499 16162 3507
rect 16170 3499 16178 3507
rect 16890 3499 16898 3507
rect 16906 3499 16914 3507
rect 19904 3500 19912 3508
rect 21760 3500 21768 3508
rect 22368 3500 22376 3508
rect 25264 3500 25272 3508
rect 25584 3500 25592 3508
rect 25744 3500 25752 3508
rect 27840 3500 27848 3508
rect 28480 3500 28488 3508
rect 38440 3505 38441 3510
rect 29856 3497 29864 3505
rect 30032 3497 30040 3505
rect 33056 3497 33064 3505
rect 33136 3497 33144 3505
rect 33168 3497 33176 3505
rect 33296 3497 33304 3505
rect 34400 3497 34408 3505
rect 35440 3497 35448 3505
rect 35728 3497 35736 3505
rect 36448 3497 36456 3505
rect 38144 3497 38152 3505
rect 38640 3497 38648 3505
rect 38688 3497 38696 3505
rect 5842 3473 5850 3481
rect 6354 3473 6362 3481
rect 6882 3473 6890 3481
rect 7442 3473 7450 3481
rect 7634 3473 7642 3481
rect 7794 3473 7802 3481
rect 8994 3473 9002 3481
rect 9042 3473 9050 3481
rect 9058 3473 9066 3481
rect 9762 3473 9770 3481
rect 9874 3473 9882 3481
rect 10114 3473 10122 3481
rect 10162 3473 10170 3481
rect 10210 3473 10218 3481
rect 10322 3473 10330 3481
rect 10402 3473 10410 3481
rect 10450 3473 10458 3481
rect 10658 3473 10666 3481
rect 10866 3473 10874 3481
rect 13450 3479 13458 3487
rect 13898 3479 13906 3487
rect 14602 3479 14610 3487
rect 16266 3479 16274 3487
rect 19296 3480 19304 3488
rect 21120 3480 21128 3488
rect 25952 3480 25960 3488
rect 28016 3480 28024 3488
rect 32944 3477 32952 3485
rect 6434 3453 6442 3461
rect 6754 3453 6762 3461
rect 6802 3453 6810 3461
rect 8018 3453 8026 3461
rect 8034 3453 8042 3461
rect 8514 3453 8522 3461
rect 8690 3453 8698 3461
rect 9618 3453 9626 3461
rect 9810 3453 9818 3461
rect 15338 3459 15346 3467
rect 15962 3459 15970 3467
rect 16026 3459 16034 3467
rect 16634 3459 16642 3467
rect 16650 3459 16658 3467
rect 17066 3459 17074 3467
rect 22976 3460 22984 3468
rect 23168 3460 23176 3468
rect 25504 3460 25512 3468
rect 25536 3460 25544 3468
rect 27424 3460 27432 3468
rect 27456 3460 27464 3468
rect 29428 3467 29440 3475
rect 29444 3467 29448 3475
rect 29460 3467 29472 3475
rect 29488 3467 29504 3475
rect 29512 3467 29544 3475
rect 29552 3467 29564 3475
rect 29584 3467 29596 3475
rect 29604 3467 29636 3475
rect 29644 3467 29660 3475
rect 29676 3467 29700 3475
rect 29708 3467 29724 3475
rect 29740 3467 29744 3475
rect 29748 3467 29752 3475
rect 29764 3467 29776 3475
rect 29780 3467 29792 3475
rect 29800 3467 29816 3475
rect 29832 3467 29880 3475
rect 29896 3467 29912 3475
rect 29920 3467 29944 3475
rect 29960 3467 29972 3475
rect 29992 3467 30004 3475
rect 30008 3467 30020 3475
rect 30024 3467 30036 3475
rect 30108 3467 30112 3475
rect 30116 3467 30128 3475
rect 30148 3467 30160 3475
rect 30164 3467 30168 3475
rect 30180 3467 30192 3475
rect 30208 3467 30224 3475
rect 30240 3467 30288 3475
rect 30304 3467 30316 3475
rect 30336 3467 30348 3475
rect 30360 3467 30364 3475
rect 30368 3467 30380 3475
rect 30400 3467 30412 3475
rect 30416 3467 30420 3475
rect 30452 3467 30456 3475
rect 30460 3467 30472 3475
rect 30544 3467 30548 3475
rect 30552 3467 30564 3475
rect 30708 3467 30720 3475
rect 30724 3467 30728 3475
rect 30740 3467 30752 3475
rect 30760 3467 30784 3475
rect 30800 3467 30824 3475
rect 30832 3467 30844 3475
rect 30856 3467 30860 3475
rect 30864 3467 30876 3475
rect 30892 3467 30916 3475
rect 30924 3467 30940 3475
rect 30956 3467 30972 3475
rect 30988 3467 30992 3475
rect 30996 3467 31008 3475
rect 31012 3467 31024 3475
rect 31028 3467 31032 3475
rect 31052 3467 31056 3475
rect 31060 3467 31064 3475
rect 31192 3467 31196 3475
rect 31200 3467 31204 3475
rect 31224 3467 31228 3475
rect 31232 3467 31244 3475
rect 31248 3467 31260 3475
rect 31264 3467 31268 3475
rect 31284 3467 31288 3475
rect 31292 3467 31296 3475
rect 31316 3467 31320 3475
rect 31324 3467 31336 3475
rect 31340 3467 31352 3475
rect 31356 3467 31360 3475
rect 31376 3467 31392 3475
rect 31408 3467 31424 3475
rect 31432 3467 31456 3475
rect 31472 3467 31496 3475
rect 31504 3467 31516 3475
rect 31528 3467 31532 3475
rect 31536 3467 31548 3475
rect 31552 3467 31556 3475
rect 31568 3467 31580 3475
rect 31660 3467 31672 3475
rect 31692 3467 31704 3475
rect 31708 3467 31720 3475
rect 31724 3467 31736 3475
rect 31752 3467 31764 3475
rect 31784 3467 31796 3475
rect 31800 3467 31812 3475
rect 31816 3467 31828 3475
rect 31848 3467 31860 3475
rect 31876 3467 31900 3475
rect 31908 3467 31924 3475
rect 31940 3467 31944 3475
rect 31948 3467 31952 3475
rect 31964 3467 31976 3475
rect 31980 3467 31992 3475
rect 32004 3467 32008 3475
rect 32012 3467 32016 3475
rect 32112 3467 32116 3475
rect 32120 3467 32132 3475
rect 32144 3467 32148 3475
rect 32152 3467 32156 3475
rect 32204 3467 32208 3475
rect 32212 3467 32224 3475
rect 32236 3467 32240 3475
rect 32244 3467 32248 3475
rect 32260 3467 32272 3475
rect 32276 3467 32280 3475
rect 32296 3467 32312 3475
rect 32328 3467 32344 3475
rect 32352 3467 32384 3475
rect 32392 3467 32404 3475
rect 32424 3467 32436 3475
rect 32440 3467 32452 3475
rect 32456 3467 32468 3475
rect 32488 3467 32500 3475
rect 32580 3467 32592 3475
rect 32604 3467 32608 3475
rect 32612 3467 32624 3475
rect 32628 3467 32632 3475
rect 32672 3467 32684 3475
rect 32696 3467 32700 3475
rect 32704 3467 32716 3475
rect 32720 3467 32724 3475
rect 32736 3467 32748 3475
rect 32760 3467 32764 3475
rect 32768 3467 32780 3475
rect 32784 3467 32788 3475
rect 32924 3467 32936 3475
rect 32940 3467 32944 3475
rect 32956 3467 32968 3475
rect 32984 3467 33000 3475
rect 33008 3467 33040 3475
rect 33048 3467 33064 3475
rect 33072 3467 33104 3475
rect 33112 3467 33128 3475
rect 33144 3467 33160 3475
rect 33176 3467 33180 3475
rect 33184 3467 33196 3475
rect 33208 3467 33212 3475
rect 33216 3467 33220 3475
rect 33332 3467 33336 3475
rect 33340 3467 33344 3475
rect 33456 3467 33460 3475
rect 33464 3467 33468 3475
rect 33480 3467 33492 3475
rect 33496 3467 33500 3475
rect 33520 3467 33524 3475
rect 33528 3467 33540 3475
rect 33552 3467 33556 3475
rect 33560 3467 33564 3475
rect 33660 3467 33664 3475
rect 33668 3467 33672 3475
rect 33692 3467 33696 3475
rect 33700 3467 33712 3475
rect 33716 3467 33728 3475
rect 33732 3467 33736 3475
rect 33752 3467 33776 3475
rect 33784 3467 33800 3475
rect 33808 3467 33832 3475
rect 33848 3467 33860 3475
rect 33880 3467 33892 3475
rect 33904 3467 33908 3475
rect 33912 3467 33924 3475
rect 33928 3467 33932 3475
rect 34036 3467 34048 3475
rect 34068 3467 34080 3475
rect 34084 3467 34088 3475
rect 34100 3467 34112 3475
rect 34132 3467 34144 3475
rect 34152 3467 34184 3475
rect 34192 3467 34208 3475
rect 34224 3467 34236 3475
rect 34244 3467 34276 3475
rect 34284 3467 34300 3475
rect 34308 3467 34332 3475
rect 34348 3467 34352 3475
rect 34356 3467 34368 3475
rect 34380 3467 34384 3475
rect 34388 3467 34392 3475
rect 34520 3467 34524 3475
rect 34528 3467 34532 3475
rect 34544 3467 34556 3475
rect 34560 3467 34564 3475
rect 34584 3467 34588 3475
rect 34592 3467 34596 3475
rect 34612 3467 34660 3475
rect 34676 3467 34680 3475
rect 34684 3467 34688 3475
rect 34704 3467 34752 3475
rect 34768 3467 34816 3475
rect 34832 3467 34848 3475
rect 34864 3467 34868 3475
rect 34872 3467 34884 3475
rect 34896 3467 34900 3475
rect 34904 3467 34908 3475
rect 35036 3467 35040 3475
rect 35044 3467 35048 3475
rect 35208 3467 35212 3475
rect 35216 3467 35228 3475
rect 35240 3467 35244 3475
rect 35248 3467 35252 3475
rect 35264 3467 35276 3475
rect 35280 3467 35292 3475
rect 35304 3467 35308 3475
rect 35312 3467 35316 3475
rect 35332 3467 35380 3475
rect 35396 3467 35408 3475
rect 35428 3467 35440 3475
rect 35452 3467 35456 3475
rect 35460 3467 35472 3475
rect 35544 3467 35548 3475
rect 35552 3467 35564 3475
rect 35584 3467 35596 3475
rect 35600 3467 35604 3475
rect 35708 3467 35720 3475
rect 35724 3467 35728 3475
rect 35740 3467 35752 3475
rect 35772 3467 35784 3475
rect 35800 3467 35848 3475
rect 35864 3467 35868 3475
rect 35872 3467 35876 3475
rect 35888 3467 35900 3475
rect 35904 3467 35916 3475
rect 35928 3467 35932 3475
rect 35936 3467 35940 3475
rect 35960 3467 35964 3475
rect 35968 3467 35972 3475
rect 36036 3467 36040 3475
rect 36044 3467 36056 3475
rect 36068 3467 36072 3475
rect 36076 3467 36080 3475
rect 36092 3467 36104 3475
rect 36108 3467 36112 3475
rect 36128 3467 36144 3475
rect 36160 3467 36176 3475
rect 36184 3467 36216 3475
rect 36224 3467 36236 3475
rect 36252 3467 36268 3475
rect 36276 3467 36308 3475
rect 36316 3467 36332 3475
rect 36348 3467 36372 3475
rect 36380 3467 36396 3475
rect 36412 3467 36416 3475
rect 36420 3467 36424 3475
rect 36436 3467 36448 3475
rect 36452 3467 36464 3475
rect 36472 3467 36488 3475
rect 36504 3467 36508 3475
rect 36512 3467 36516 3475
rect 36528 3467 36540 3475
rect 36544 3467 36556 3475
rect 36568 3467 36572 3475
rect 36576 3467 36580 3475
rect 36592 3467 36604 3475
rect 36608 3467 36612 3475
rect 36676 3467 36680 3475
rect 36684 3467 36688 3475
rect 36708 3467 36712 3475
rect 36716 3467 36720 3475
rect 36732 3467 36744 3475
rect 36748 3467 36760 3475
rect 36772 3467 36776 3475
rect 36780 3467 36784 3475
rect 36800 3467 36816 3475
rect 36824 3467 36836 3475
rect 36840 3467 36852 3475
rect 36864 3467 36868 3475
rect 36872 3467 36876 3475
rect 36896 3467 36900 3475
rect 36904 3467 36908 3475
rect 37004 3467 37008 3475
rect 37012 3467 37016 3475
rect 37028 3467 37040 3475
rect 37044 3467 37056 3475
rect 37068 3467 37072 3475
rect 37076 3467 37080 3475
rect 37208 3467 37212 3475
rect 37216 3467 37220 3475
rect 37268 3467 37272 3475
rect 37276 3467 37288 3475
rect 37300 3467 37304 3475
rect 37308 3467 37312 3475
rect 37324 3467 37336 3475
rect 37340 3467 37344 3475
rect 37504 3467 37508 3475
rect 37512 3467 37516 3475
rect 37528 3467 37540 3475
rect 37544 3467 37548 3475
rect 37612 3467 37616 3475
rect 37620 3467 37624 3475
rect 37644 3467 37648 3475
rect 37652 3467 37656 3475
rect 37668 3467 37680 3475
rect 37684 3467 37696 3475
rect 37704 3467 37720 3475
rect 37736 3467 37784 3475
rect 37800 3467 37816 3475
rect 37832 3467 37844 3475
rect 37856 3467 37860 3475
rect 37864 3467 37876 3475
rect 37980 3467 37984 3475
rect 37988 3467 38000 3475
rect 38020 3467 38032 3475
rect 38036 3467 38040 3475
rect 38112 3467 38124 3475
rect 38128 3467 38132 3475
rect 38144 3467 38156 3475
rect 38176 3467 38188 3475
rect 38192 3467 38196 3475
rect 38208 3467 38220 3475
rect 38232 3467 38236 3475
rect 38240 3467 38252 3475
rect 38268 3467 38280 3475
rect 38284 3467 38288 3475
rect 38300 3467 38312 3475
rect 38324 3467 38328 3475
rect 38332 3467 38344 3475
rect 38348 3467 38352 3475
rect 38364 3467 38376 3475
rect 38456 3467 38468 3475
rect 38488 3467 38500 3475
rect 38504 3467 38516 3475
rect 38520 3467 38532 3475
rect 38552 3467 38564 3475
rect 38572 3467 38604 3475
rect 38612 3467 38628 3475
rect 38644 3467 38660 3475
rect 38676 3467 38680 3475
rect 38684 3467 38696 3475
rect 38708 3467 38712 3475
rect 38716 3467 38720 3475
rect 38848 3467 38852 3475
rect 38856 3467 38860 3475
rect 38940 3467 38944 3475
rect 38948 3467 38952 3475
rect 38964 3467 38976 3475
rect 38980 3467 38984 3475
rect 39004 3467 39008 3475
rect 39012 3467 39016 3475
rect 39028 3467 39040 3475
rect 39044 3467 39056 3475
rect 39068 3467 39072 3475
rect 39076 3467 39080 3475
rect 39100 3467 39104 3475
rect 39108 3467 39112 3475
rect 39240 3467 39244 3475
rect 39248 3467 39260 3475
rect 39272 3467 39276 3475
rect 39280 3467 39284 3475
rect 39296 3467 39308 3475
rect 39312 3467 39324 3475
rect 39332 3467 39348 3475
rect 39364 3467 39368 3475
rect 39372 3467 39376 3475
rect 39388 3467 39400 3475
rect 39404 3467 39416 3475
rect 39428 3467 39432 3475
rect 39436 3467 39440 3475
rect 39456 3467 39472 3475
rect 39480 3467 39504 3475
rect 39520 3467 39536 3475
rect 39552 3467 39564 3475
rect 39568 3467 39580 3475
rect 39584 3467 39596 3475
rect 39772 3467 39784 3475
rect 39896 3467 39908 3475
rect 39912 3467 39916 3475
rect 39928 3467 39940 3475
rect 39956 3467 39972 3475
rect 39980 3467 40012 3475
rect 40020 3467 40036 3475
rect 40044 3467 40056 3475
rect 40060 3467 40064 3475
rect 40084 3467 40088 3475
rect 40092 3467 40104 3475
rect 40116 3467 40120 3475
rect 40124 3467 40128 3475
rect 40148 3467 40152 3475
rect 40156 3467 40160 3475
rect 40224 3467 40228 3475
rect 40232 3467 40236 3475
rect 40412 3467 40416 3475
rect 40420 3467 40424 3475
rect 40436 3467 40448 3475
rect 40452 3467 40456 3475
rect 40472 3467 40488 3475
rect 40504 3467 40552 3475
rect 40568 3467 40580 3475
rect 40584 3467 40588 3475
rect 40600 3467 40612 3475
rect 40624 3467 40628 3475
rect 40632 3467 40644 3475
rect 40780 3467 40784 3475
rect 40788 3467 40800 3475
rect 18740 3452 18742 3460
rect 19098 3450 19106 3458
rect 19248 3450 19254 3458
rect 19708 3450 19716 3458
rect 19858 3450 19864 3458
rect 20334 3450 20348 3458
rect 20858 3450 20872 3458
rect 21180 3452 21182 3460
rect 22844 3450 22848 3458
rect 22934 3450 22942 3458
rect 23052 3456 23054 3460
rect 23250 3456 23252 3460
rect 23058 3452 23060 3456
rect 23256 3452 23258 3456
rect 23454 3450 23458 3458
rect 23544 3450 23552 3458
rect 25022 3452 25024 3460
rect 25236 3452 25238 3460
rect 25326 3450 25334 3458
rect 25476 3450 25482 3458
rect 27022 3450 27030 3458
rect 27172 3450 27178 3458
rect 27236 3450 27244 3458
rect 27386 3450 27392 3458
rect 28306 3450 28314 3458
rect 28456 3450 28462 3458
rect 29936 3457 29944 3465
rect 32656 3457 32664 3465
rect 33040 3457 33048 3465
rect 36832 3457 36840 3465
rect 40432 3457 40440 3465
rect 6834 3433 6842 3441
rect 7010 3433 7018 3441
rect 7954 3433 7962 3441
rect 8626 3433 8634 3441
rect 8722 3433 8730 3441
rect 8738 3433 8746 3441
rect 8962 3433 8970 3441
rect 9106 3433 9114 3441
rect 9442 3433 9450 3441
rect 9522 3433 9530 3441
rect 9826 3433 9834 3441
rect 13002 3439 13010 3447
rect 13722 3439 13730 3447
rect 13786 3439 13794 3447
rect 14250 3439 14258 3447
rect 15482 3439 15490 3447
rect 16266 3439 16274 3447
rect 20704 3440 20712 3448
rect 23408 3440 23416 3448
rect 26560 3440 26568 3448
rect 27200 3440 27208 3448
rect 29904 3437 29912 3445
rect 30256 3437 30264 3445
rect 30400 3437 30408 3445
rect 30704 3437 30712 3445
rect 31104 3437 31112 3445
rect 31424 3437 31432 3445
rect 31648 3437 31656 3445
rect 32352 3437 32360 3445
rect 32960 3437 32968 3445
rect 33712 3437 33720 3445
rect 33984 3437 33992 3445
rect 34336 3437 34344 3445
rect 34608 3437 34616 3445
rect 34752 3437 34760 3445
rect 35008 3437 35016 3445
rect 35408 3437 35416 3445
rect 35424 3437 35432 3445
rect 36192 3437 36200 3445
rect 36432 3437 36440 3445
rect 36576 3437 36584 3445
rect 37168 3437 37176 3445
rect 37312 3437 37320 3445
rect 37360 3437 37368 3445
rect 37632 3437 37640 3445
rect 38096 3437 38104 3445
rect 38752 3437 38760 3445
rect 38960 3437 38968 3445
rect 39328 3437 39336 3445
rect 5874 3413 5882 3421
rect 6066 3413 6074 3421
rect 6306 3413 6314 3421
rect 6354 3413 6362 3421
rect 6674 3413 6682 3421
rect 7634 3413 7642 3421
rect 8034 3413 8042 3421
rect 8866 3413 8874 3421
rect 9202 3413 9210 3421
rect 9266 3413 9274 3421
rect 10178 3413 10186 3421
rect 10194 3413 10202 3421
rect 10482 3413 10490 3421
rect 10770 3413 10778 3421
rect 12314 3419 12322 3427
rect 12570 3419 12578 3427
rect 12618 3419 12626 3427
rect 12890 3419 12898 3427
rect 13034 3419 13042 3427
rect 13466 3419 13474 3427
rect 13914 3419 13922 3427
rect 14138 3419 14146 3427
rect 14234 3419 14242 3427
rect 14426 3419 14434 3427
rect 17226 3419 17234 3427
rect 19456 3420 19464 3428
rect 20080 3420 20088 3428
rect 21088 3420 21096 3428
rect 21744 3420 21752 3428
rect 22560 3420 22568 3428
rect 22768 3420 22776 3428
rect 23792 3420 23800 3428
rect 24464 3420 24472 3428
rect 24480 3420 24488 3428
rect 25296 3420 25304 3428
rect 25584 3420 25592 3428
rect 25712 3420 25720 3428
rect 26960 3420 26968 3428
rect 29680 3417 29688 3425
rect 30064 3417 30072 3425
rect 30368 3417 30376 3425
rect 30512 3417 30520 3425
rect 30544 3417 30552 3425
rect 31152 3417 31160 3425
rect 31296 3417 31304 3425
rect 31312 3417 31320 3425
rect 31728 3417 31736 3425
rect 32864 3417 32872 3425
rect 33008 3417 33016 3425
rect 37568 3417 37576 3425
rect 37920 3417 37928 3425
rect 38144 3417 38152 3425
rect 38432 3417 38440 3425
rect 39888 3417 39896 3425
rect 40320 3417 40328 3425
rect 40400 3417 40408 3425
rect 5730 3393 5738 3401
rect 5778 3393 5786 3401
rect 6018 3393 6026 3401
rect 6514 3393 6522 3401
rect 6690 3393 6698 3401
rect 6738 3393 6746 3401
rect 6834 3393 6842 3401
rect 7010 3393 7018 3401
rect 7026 3393 7034 3401
rect 7042 3393 7050 3401
rect 7090 3393 7098 3401
rect 7106 3393 7114 3401
rect 7138 3393 7146 3401
rect 7170 3393 7178 3401
rect 7330 3393 7338 3401
rect 7442 3393 7450 3401
rect 7602 3393 7610 3401
rect 7842 3393 7850 3401
rect 7874 3393 7882 3401
rect 8114 3393 8122 3401
rect 8162 3393 8170 3401
rect 8194 3393 8202 3401
rect 8226 3393 8234 3401
rect 8290 3393 8298 3401
rect 8386 3393 8394 3401
rect 8418 3393 8426 3401
rect 8562 3393 8570 3401
rect 8770 3393 8778 3401
rect 8914 3393 8922 3401
rect 9058 3393 9066 3401
rect 9106 3393 9114 3401
rect 9218 3393 9226 3401
rect 9282 3393 9290 3401
rect 9426 3393 9434 3401
rect 9506 3393 9514 3401
rect 9714 3393 9722 3401
rect 9970 3393 9978 3401
rect 10098 3393 10106 3401
rect 10114 3393 10122 3401
rect 10226 3393 10234 3401
rect 10562 3393 10570 3401
rect 10770 3393 10778 3401
rect 10850 3393 10858 3401
rect 12106 3399 12114 3407
rect 12234 3399 12242 3407
rect 14538 3399 14546 3407
rect 15002 3399 15010 3407
rect 15066 3399 15074 3407
rect 15562 3399 15570 3407
rect 15642 3399 15650 3407
rect 15690 3399 15698 3407
rect 16842 3399 16850 3407
rect 16986 3399 16994 3407
rect 18672 3400 18680 3408
rect 25536 3400 25544 3408
rect 27456 3400 27464 3408
rect 27504 3400 27512 3408
rect 30240 3397 30248 3405
rect 32864 3397 32872 3405
rect 33296 3397 33304 3405
rect 33600 3397 33608 3405
rect 36768 3397 36776 3405
rect 38304 3397 38312 3405
rect 38368 3397 38376 3405
rect 38544 3397 38552 3405
rect 38768 3397 38776 3405
rect 39264 3397 39272 3405
rect 39328 3397 39336 3405
rect 39632 3397 39640 3405
rect 39872 3397 39880 3405
rect 39920 3397 39928 3405
rect 40176 3397 40184 3405
rect 40688 3397 40696 3405
rect 6002 3373 6010 3381
rect 6082 3373 6090 3381
rect 6290 3373 6298 3381
rect 6482 3373 6490 3381
rect 6514 3373 6522 3381
rect 6530 3373 6538 3381
rect 6738 3373 6746 3381
rect 6866 3373 6874 3381
rect 6882 3373 6890 3381
rect 6994 3373 7002 3381
rect 7506 3373 7514 3381
rect 9090 3373 9098 3381
rect 9122 3373 9130 3381
rect 9154 3373 9162 3381
rect 9170 3373 9178 3381
rect 9682 3373 9690 3381
rect 9714 3373 9722 3381
rect 9794 3373 9802 3381
rect 9906 3373 9914 3381
rect 10002 3373 10010 3381
rect 10114 3373 10122 3381
rect 10834 3373 10842 3381
rect 10882 3373 10890 3381
rect 12362 3379 12370 3387
rect 12378 3379 12386 3387
rect 12554 3379 12562 3387
rect 12618 3379 12626 3387
rect 13610 3379 13618 3387
rect 13786 3379 13794 3387
rect 14090 3379 14098 3387
rect 14522 3379 14530 3387
rect 14682 3379 14690 3387
rect 14698 3379 14706 3387
rect 14938 3379 14946 3387
rect 15082 3379 15090 3387
rect 15306 3379 15314 3387
rect 15338 3379 15346 3387
rect 15626 3379 15634 3387
rect 16058 3379 16066 3387
rect 16618 3379 16626 3387
rect 16778 3379 16786 3387
rect 17066 3379 17074 3387
rect 17370 3379 17378 3387
rect 18512 3380 18520 3388
rect 19408 3380 19416 3388
rect 19824 3380 19832 3388
rect 20032 3380 20040 3388
rect 20240 3380 20248 3388
rect 20320 3380 20328 3388
rect 20928 3380 20936 3388
rect 21696 3380 21704 3388
rect 22336 3380 22344 3388
rect 22592 3380 22600 3388
rect 22960 3380 22968 3388
rect 23104 3380 23112 3388
rect 23344 3380 23352 3388
rect 24288 3380 24296 3388
rect 24624 3380 24632 3388
rect 26592 3380 26600 3388
rect 27872 3380 27880 3388
rect 28128 3380 28136 3388
rect 29920 3377 29928 3385
rect 30928 3377 30936 3385
rect 30992 3377 31000 3385
rect 31104 3377 31112 3385
rect 32144 3377 32152 3385
rect 32288 3377 32296 3385
rect 33136 3377 33144 3385
rect 33424 3377 33432 3385
rect 39488 3377 39496 3385
rect 8514 3353 8522 3361
rect 8546 3353 8554 3361
rect 8594 3353 8602 3361
rect 8802 3353 8810 3361
rect 9282 3353 9290 3361
rect 9458 3353 9466 3361
rect 9618 3353 9626 3361
rect 10034 3353 10042 3361
rect 10082 3353 10090 3361
rect 10450 3353 10458 3361
rect 10514 3353 10522 3361
rect 10626 3353 10634 3361
rect 10738 3353 10746 3361
rect 13242 3359 13250 3367
rect 13338 3359 13346 3367
rect 13738 3359 13746 3367
rect 13946 3359 13954 3367
rect 14666 3359 14674 3367
rect 14746 3359 14754 3367
rect 15306 3359 15314 3367
rect 15386 3359 15394 3367
rect 15786 3359 15794 3367
rect 15834 3359 15842 3367
rect 17306 3359 17314 3367
rect 19872 3360 19880 3368
rect 25120 3360 25128 3368
rect 25760 3360 25768 3368
rect 30224 3357 30232 3365
rect 30480 3357 30488 3365
rect 32816 3357 32824 3365
rect 32992 3357 33000 3365
rect 33584 3357 33592 3365
rect 36144 3357 36152 3365
rect 40160 3357 40168 3365
rect 40256 3357 40264 3365
rect 19040 3348 19044 3353
rect 22352 3348 22356 3353
rect 5810 3333 5818 3341
rect 5826 3333 5834 3341
rect 6066 3333 6074 3341
rect 6082 3333 6090 3341
rect 6114 3333 6122 3341
rect 6786 3333 6794 3341
rect 6850 3333 6858 3341
rect 8338 3333 8346 3341
rect 9522 3333 9530 3341
rect 9698 3333 9706 3341
rect 10898 3333 10906 3341
rect 12042 3339 12050 3347
rect 13498 3339 13506 3347
rect 14554 3339 14562 3347
rect 14650 3339 14658 3347
rect 15178 3339 15186 3347
rect 15242 3339 15250 3347
rect 15898 3339 15906 3347
rect 16042 3339 16050 3347
rect 16458 3339 16466 3347
rect 16570 3339 16578 3347
rect 16666 3339 16674 3347
rect 17034 3339 17042 3347
rect 17178 3339 17186 3347
rect 17258 3339 17266 3347
rect 17514 3339 17522 3347
rect 18496 3340 18504 3348
rect 18656 3340 18664 3348
rect 18832 3340 18840 3348
rect 19632 3340 19640 3348
rect 19840 3340 19848 3348
rect 20048 3340 20056 3348
rect 20656 3340 20664 3348
rect 20848 3340 20856 3348
rect 21488 3340 21496 3348
rect 22128 3340 22136 3348
rect 22608 3340 22616 3348
rect 23168 3340 23176 3348
rect 23840 3340 23848 3348
rect 24208 3340 24216 3348
rect 24272 3340 24280 3348
rect 24304 3340 24312 3348
rect 25456 3340 25464 3348
rect 26576 3340 26584 3348
rect 27152 3340 27160 3348
rect 28080 3340 28088 3348
rect 28224 3340 28232 3348
rect 31840 3337 31848 3345
rect 36048 3337 36056 3345
rect 37296 3337 37304 3345
rect 6002 3313 6010 3321
rect 7090 3313 7098 3321
rect 7314 3313 7322 3321
rect 7378 3313 7386 3321
rect 7410 3313 7418 3321
rect 7826 3313 7834 3321
rect 8210 3313 8218 3321
rect 10770 3313 10778 3321
rect 23008 3320 23016 3328
rect 23152 3320 23160 3328
rect 23632 3320 23640 3328
rect 25968 3320 25976 3328
rect 34192 3317 34200 3325
rect 34800 3317 34808 3325
rect 35664 3317 35672 3325
rect 35680 3317 35688 3325
rect 35952 3317 35960 3325
rect 36976 3317 36984 3325
rect 6562 3293 6570 3301
rect 7282 3293 7290 3301
rect 7762 3293 7770 3301
rect 7842 3293 7850 3301
rect 8706 3293 8714 3301
rect 9202 3293 9210 3301
rect 13322 3299 13330 3307
rect 15258 3299 15266 3307
rect 15866 3299 15874 3307
rect 16106 3299 16114 3307
rect 21696 3300 21704 3308
rect 6498 3273 6506 3281
rect 7122 3273 7130 3281
rect 7618 3273 7626 3281
rect 9954 3273 9962 3281
rect 10322 3273 10330 3281
rect 10354 3273 10362 3281
rect 10594 3273 10602 3281
rect 10754 3273 10762 3281
rect 10834 3273 10842 3281
rect 13898 3279 13906 3287
rect 17098 3279 17106 3287
rect 40480 3277 40488 3285
rect 29420 3267 29424 3275
rect 29428 3267 29440 3275
rect 29444 3267 29448 3275
rect 29488 3267 29500 3275
rect 29512 3267 29516 3275
rect 29520 3267 29532 3275
rect 29536 3267 29540 3275
rect 29604 3267 29608 3275
rect 29612 3267 29624 3275
rect 29628 3267 29632 3275
rect 29644 3267 29656 3275
rect 29668 3267 29672 3275
rect 29676 3267 29688 3275
rect 29692 3267 29696 3275
rect 29708 3267 29720 3275
rect 29736 3267 29752 3275
rect 29768 3267 29792 3275
rect 29800 3267 29816 3275
rect 29824 3267 29856 3275
rect 29864 3267 29880 3275
rect 29896 3267 29908 3275
rect 29920 3267 29924 3275
rect 29928 3267 29940 3275
rect 30052 3267 30064 3275
rect 30076 3267 30080 3275
rect 30084 3267 30096 3275
rect 30100 3267 30104 3275
rect 30208 3267 30220 3275
rect 30240 3267 30252 3275
rect 30256 3267 30268 3275
rect 30272 3267 30284 3275
rect 30460 3267 30472 3275
rect 30492 3267 30504 3275
rect 30508 3267 30520 3275
rect 30524 3267 30536 3275
rect 30552 3267 30568 3275
rect 30584 3267 30596 3275
rect 30600 3267 30612 3275
rect 30616 3267 30628 3275
rect 30648 3267 30660 3275
rect 30680 3267 30692 3275
rect 30712 3267 30724 3275
rect 30744 3267 30756 3275
rect 30760 3267 30772 3275
rect 30776 3267 30788 3275
rect 30808 3267 30820 3275
rect 30828 3267 30860 3275
rect 30868 3267 30884 3275
rect 30892 3267 30916 3275
rect 30932 3267 30948 3275
rect 30956 3267 30980 3275
rect 30996 3267 31008 3275
rect 31012 3267 31016 3275
rect 31028 3267 31040 3275
rect 31052 3267 31056 3275
rect 31060 3267 31072 3275
rect 31216 3267 31228 3275
rect 31232 3267 31244 3275
rect 31248 3267 31260 3275
rect 31276 3267 31288 3275
rect 31308 3267 31320 3275
rect 31324 3267 31336 3275
rect 31340 3267 31352 3275
rect 31372 3267 31384 3275
rect 31400 3267 31424 3275
rect 31432 3267 31448 3275
rect 31464 3267 31468 3275
rect 31472 3267 31476 3275
rect 31488 3267 31500 3275
rect 31504 3267 31516 3275
rect 31528 3267 31532 3275
rect 31536 3267 31540 3275
rect 31552 3267 31564 3275
rect 31568 3267 31580 3275
rect 31592 3267 31596 3275
rect 31600 3267 31604 3275
rect 31748 3267 31752 3275
rect 31756 3267 31760 3275
rect 31780 3267 31784 3275
rect 31788 3267 31792 3275
rect 31952 3267 31956 3275
rect 31960 3267 31972 3275
rect 31976 3267 31988 3275
rect 31992 3267 31996 3275
rect 32016 3267 32020 3275
rect 32024 3267 32028 3275
rect 32048 3267 32052 3275
rect 32056 3267 32060 3275
rect 32080 3267 32084 3275
rect 32088 3267 32092 3275
rect 32112 3267 32116 3275
rect 32120 3267 32132 3275
rect 32136 3267 32148 3275
rect 32152 3267 32156 3275
rect 32396 3267 32400 3275
rect 32404 3267 32408 3275
rect 32428 3267 32432 3275
rect 32436 3267 32448 3275
rect 32452 3267 32464 3275
rect 32468 3267 32472 3275
rect 32492 3267 32496 3275
rect 32500 3267 32504 3275
rect 32524 3267 32528 3275
rect 32532 3267 32536 3275
rect 32556 3267 32560 3275
rect 32564 3267 32568 3275
rect 32588 3267 32592 3275
rect 32596 3267 32608 3275
rect 32612 3267 32624 3275
rect 32628 3267 32632 3275
rect 32792 3267 32796 3275
rect 32800 3267 32804 3275
rect 32824 3267 32828 3275
rect 32832 3267 32844 3275
rect 32848 3267 32860 3275
rect 32864 3267 32868 3275
rect 32888 3267 32892 3275
rect 32896 3267 32900 3275
rect 32916 3267 32920 3275
rect 32924 3267 32936 3275
rect 32940 3267 32952 3275
rect 32956 3267 32960 3275
rect 32976 3267 33000 3275
rect 33008 3267 33024 3275
rect 33032 3267 33056 3275
rect 33072 3267 33076 3275
rect 33080 3267 33092 3275
rect 33096 3267 33108 3275
rect 33112 3267 33116 3275
rect 33136 3267 33140 3275
rect 33144 3267 33148 3275
rect 33164 3267 33168 3275
rect 33172 3267 33184 3275
rect 33188 3267 33200 3275
rect 33204 3267 33208 3275
rect 33224 3267 33228 3275
rect 33232 3267 33236 3275
rect 33256 3267 33260 3275
rect 33264 3267 33276 3275
rect 33280 3267 33292 3275
rect 33296 3267 33300 3275
rect 33320 3267 33324 3275
rect 33328 3267 33332 3275
rect 33348 3267 33364 3275
rect 33372 3267 33396 3275
rect 33412 3267 33436 3275
rect 33444 3267 33460 3275
rect 33476 3267 33500 3275
rect 33508 3267 33524 3275
rect 33532 3267 33544 3275
rect 33548 3267 33552 3275
rect 33568 3267 33592 3275
rect 33600 3267 33616 3275
rect 33624 3267 33656 3275
rect 33664 3267 33676 3275
rect 33696 3267 33708 3275
rect 33712 3267 33724 3275
rect 33728 3267 33740 3275
rect 33852 3267 33864 3275
rect 33876 3267 33880 3275
rect 33884 3267 33896 3275
rect 33900 3267 33904 3275
rect 33916 3267 33928 3275
rect 33944 3267 33956 3275
rect 33968 3267 33972 3275
rect 33976 3267 33988 3275
rect 33992 3267 33996 3275
rect 34008 3267 34020 3275
rect 34028 3267 34052 3275
rect 34068 3267 34080 3275
rect 34084 3267 34088 3275
rect 34100 3267 34112 3275
rect 34124 3267 34128 3275
rect 34132 3267 34144 3275
rect 34160 3267 34172 3275
rect 34176 3267 34180 3275
rect 34192 3267 34204 3275
rect 34216 3267 34220 3275
rect 34224 3267 34236 3275
rect 34252 3267 34276 3275
rect 34284 3267 34296 3275
rect 34308 3267 34312 3275
rect 34316 3267 34328 3275
rect 34344 3267 34356 3275
rect 34360 3267 34364 3275
rect 34376 3267 34388 3275
rect 34400 3267 34420 3275
rect 34436 3267 34460 3275
rect 34468 3267 34480 3275
rect 34492 3267 34496 3275
rect 34500 3267 34512 3275
rect 34528 3267 34540 3275
rect 34544 3267 34548 3275
rect 34560 3267 34572 3275
rect 34584 3267 34588 3275
rect 34592 3267 34604 3275
rect 34620 3267 34644 3275
rect 34652 3267 34668 3275
rect 34684 3267 34700 3275
rect 34716 3267 34720 3275
rect 34724 3267 34736 3275
rect 34740 3267 34752 3275
rect 34756 3267 34760 3275
rect 34780 3267 34784 3275
rect 34788 3267 34800 3275
rect 34812 3267 34816 3275
rect 34820 3267 34824 3275
rect 34844 3267 34848 3275
rect 34852 3267 34856 3275
rect 34876 3267 34880 3275
rect 34884 3267 34888 3275
rect 34900 3267 34912 3275
rect 34916 3267 34920 3275
rect 34936 3267 34960 3275
rect 34968 3267 34984 3275
rect 34992 3267 35024 3275
rect 35032 3267 35044 3275
rect 35060 3267 35076 3275
rect 35084 3267 35116 3275
rect 35124 3267 35140 3275
rect 35156 3267 35168 3275
rect 35172 3267 35184 3275
rect 35188 3267 35200 3275
rect 35216 3267 35228 3275
rect 35248 3267 35260 3275
rect 35264 3267 35276 3275
rect 35280 3267 35292 3275
rect 35340 3267 35352 3275
rect 35356 3267 35368 3275
rect 35372 3267 35384 3275
rect 35400 3267 35416 3275
rect 35424 3267 35456 3275
rect 35464 3267 35480 3275
rect 35492 3267 35508 3275
rect 35516 3267 35548 3275
rect 35556 3267 35568 3275
rect 35588 3267 35600 3275
rect 35608 3267 35640 3275
rect 35648 3267 35664 3275
rect 35672 3267 35696 3275
rect 35708 3267 35732 3275
rect 35740 3267 35756 3275
rect 35764 3267 35788 3275
rect 35804 3267 35808 3275
rect 35812 3267 35824 3275
rect 35832 3267 35848 3275
rect 35856 3267 35868 3275
rect 35872 3267 35876 3275
rect 35896 3267 35900 3275
rect 35904 3267 35916 3275
rect 35928 3267 35932 3275
rect 35936 3267 35940 3275
rect 35960 3267 35964 3275
rect 35968 3267 35972 3275
rect 36036 3267 36040 3275
rect 36044 3267 36048 3275
rect 36068 3267 36072 3275
rect 36076 3267 36088 3275
rect 36092 3267 36104 3275
rect 36108 3267 36112 3275
rect 36128 3267 36132 3275
rect 36136 3267 36140 3275
rect 36160 3267 36164 3275
rect 36168 3267 36180 3275
rect 36184 3267 36196 3275
rect 36200 3267 36204 3275
rect 36220 3267 36224 3275
rect 36228 3267 36232 3275
rect 36252 3267 36256 3275
rect 36260 3267 36272 3275
rect 36276 3267 36288 3275
rect 36292 3267 36296 3275
rect 36424 3267 36428 3275
rect 36432 3267 36444 3275
rect 36448 3267 36460 3275
rect 36464 3267 36468 3275
rect 36484 3267 36488 3275
rect 36492 3267 36496 3275
rect 36516 3267 36520 3275
rect 36524 3267 36536 3275
rect 36540 3267 36552 3275
rect 36556 3267 36560 3275
rect 36576 3267 36600 3275
rect 36608 3267 36624 3275
rect 36632 3267 36656 3275
rect 36672 3267 36688 3275
rect 36696 3267 36720 3275
rect 36736 3267 36748 3275
rect 36752 3267 36756 3275
rect 36768 3267 36780 3275
rect 36792 3267 36796 3275
rect 36800 3267 36812 3275
rect 36828 3267 36840 3275
rect 36844 3267 36848 3275
rect 36860 3267 36872 3275
rect 36884 3267 36888 3275
rect 36892 3267 36904 3275
rect 36920 3267 36968 3275
rect 36984 3267 37000 3275
rect 37012 3267 37060 3275
rect 37076 3267 37092 3275
rect 37108 3267 37124 3275
rect 37140 3267 37156 3275
rect 37172 3267 37220 3275
rect 37236 3267 37240 3275
rect 37244 3267 37248 3275
rect 37260 3267 37272 3275
rect 37276 3267 37288 3275
rect 37300 3267 37304 3275
rect 37308 3267 37312 3275
rect 37328 3267 37344 3275
rect 37352 3267 37364 3275
rect 37368 3267 37380 3275
rect 37392 3267 37396 3275
rect 37400 3267 37404 3275
rect 37420 3267 37468 3275
rect 37484 3267 37496 3275
rect 37512 3267 37560 3275
rect 37576 3267 37592 3275
rect 37608 3267 37620 3275
rect 37632 3267 37636 3275
rect 37640 3267 37652 3275
rect 37672 3267 37684 3275
rect 37688 3267 37692 3275
rect 37704 3267 37716 3275
rect 37736 3267 37748 3275
rect 37752 3267 37756 3275
rect 37768 3267 37780 3275
rect 37792 3267 37796 3275
rect 37800 3267 37812 3275
rect 37956 3267 37968 3275
rect 37972 3267 37984 3275
rect 37988 3267 38000 3275
rect 38020 3267 38032 3275
rect 38048 3267 38060 3275
rect 38064 3267 38076 3275
rect 38080 3267 38092 3275
rect 38108 3267 38124 3275
rect 38140 3267 38164 3275
rect 38172 3267 38188 3275
rect 38204 3267 38208 3275
rect 38212 3267 38216 3275
rect 38228 3267 38240 3275
rect 38244 3267 38256 3275
rect 38264 3267 38280 3275
rect 38296 3267 38300 3275
rect 38304 3267 38308 3275
rect 38320 3267 38332 3275
rect 38336 3267 38348 3275
rect 38360 3267 38364 3275
rect 38368 3267 38372 3275
rect 38388 3267 38400 3275
rect 38412 3267 38436 3275
rect 38452 3267 38464 3275
rect 38484 3267 38496 3275
rect 38500 3267 38512 3275
rect 38516 3267 38528 3275
rect 38544 3267 38560 3275
rect 38576 3267 38588 3275
rect 38592 3267 38604 3275
rect 38608 3267 38620 3275
rect 38636 3267 38652 3275
rect 38668 3267 38680 3275
rect 38684 3267 38696 3275
rect 38700 3267 38712 3275
rect 38728 3267 38740 3275
rect 38760 3267 38772 3275
rect 38776 3267 38788 3275
rect 38792 3267 38804 3275
rect 38820 3267 38836 3275
rect 38852 3267 38864 3275
rect 38868 3267 38880 3275
rect 38884 3267 38896 3275
rect 38912 3267 38928 3275
rect 38944 3267 38956 3275
rect 38960 3267 38972 3275
rect 38976 3267 38988 3275
rect 39004 3267 39020 3275
rect 39028 3267 39060 3275
rect 39068 3267 39084 3275
rect 39100 3267 39104 3275
rect 39108 3267 39112 3275
rect 39132 3267 39136 3275
rect 39140 3267 39152 3275
rect 39164 3267 39168 3275
rect 39172 3267 39176 3275
rect 39272 3267 39276 3275
rect 39280 3267 39284 3275
rect 39304 3267 39308 3275
rect 39312 3267 39324 3275
rect 39328 3267 39340 3275
rect 39344 3267 39348 3275
rect 39364 3267 39368 3275
rect 39372 3267 39376 3275
rect 39396 3267 39400 3275
rect 39404 3267 39416 3275
rect 39420 3267 39432 3275
rect 39436 3267 39440 3275
rect 39460 3267 39464 3275
rect 39468 3267 39472 3275
rect 39488 3267 39504 3275
rect 39512 3267 39536 3275
rect 39552 3267 39576 3275
rect 39584 3267 39600 3275
rect 39616 3267 39632 3275
rect 39648 3267 39664 3275
rect 39672 3267 39696 3275
rect 39712 3267 39724 3275
rect 39728 3267 39732 3275
rect 39744 3267 39756 3275
rect 39768 3267 39772 3275
rect 39776 3267 39788 3275
rect 39804 3267 39816 3275
rect 39820 3267 39824 3275
rect 39836 3267 39848 3275
rect 39860 3267 39864 3275
rect 39868 3267 39880 3275
rect 39900 3267 39912 3275
rect 40024 3267 40036 3275
rect 40040 3267 40052 3275
rect 40056 3267 40068 3275
rect 40084 3267 40100 3275
rect 40116 3267 40140 3275
rect 40148 3267 40164 3275
rect 40180 3267 40228 3275
rect 40240 3267 40256 3275
rect 40272 3267 40320 3275
rect 40336 3267 40340 3275
rect 40344 3267 40348 3275
rect 40360 3267 40372 3275
rect 40376 3267 40388 3275
rect 40400 3267 40404 3275
rect 40408 3267 40412 3275
rect 40432 3267 40436 3275
rect 40440 3267 40452 3275
rect 40464 3267 40468 3275
rect 40472 3267 40476 3275
rect 40496 3267 40500 3275
rect 40504 3267 40508 3275
rect 40604 3267 40608 3275
rect 40612 3267 40616 3275
rect 40628 3267 40640 3275
rect 40644 3267 40648 3275
rect 40668 3267 40672 3275
rect 40676 3267 40680 3275
rect 40696 3267 40712 3275
rect 40720 3267 40752 3275
rect 40760 3267 40772 3275
rect 40788 3267 40800 3275
rect 6050 3253 6058 3261
rect 7586 3253 7594 3261
rect 7698 3253 7706 3261
rect 8226 3253 8234 3261
rect 22460 3250 22462 3258
rect 22468 3250 22470 3258
rect 25392 3250 25394 3258
rect 25400 3250 25402 3258
rect 27310 3250 27320 3258
rect 28380 3250 28390 3258
rect 37952 3257 37960 3265
rect 6178 3233 6186 3241
rect 8834 3233 8842 3241
rect 8850 3233 8858 3241
rect 9490 3233 9498 3241
rect 10450 3233 10458 3241
rect 12058 3239 12066 3247
rect 16138 3239 16146 3247
rect 27200 3240 27208 3248
rect 32656 3237 32664 3245
rect 33664 3237 33672 3245
rect 40384 3237 40392 3245
rect 7794 3213 7802 3221
rect 8450 3213 8458 3221
rect 8850 3213 8858 3221
rect 9554 3213 9562 3221
rect 9570 3213 9578 3221
rect 10242 3213 10250 3221
rect 10274 3213 10282 3221
rect 12682 3219 12690 3227
rect 14346 3219 14354 3227
rect 15306 3219 15314 3227
rect 16266 3219 16274 3227
rect 28096 3220 28104 3228
rect 31056 3217 31064 3225
rect 35360 3217 35368 3225
rect 36320 3217 36328 3225
rect 6674 3193 6682 3201
rect 8034 3193 8042 3201
rect 8642 3193 8650 3201
rect 14922 3199 14930 3207
rect 15594 3199 15602 3207
rect 15626 3199 15634 3207
rect 16570 3199 16578 3207
rect 17290 3199 17298 3207
rect 17546 3199 17554 3207
rect 22944 3200 22952 3208
rect 24288 3200 24296 3208
rect 27600 3200 27608 3208
rect 6802 3173 6810 3181
rect 7026 3173 7034 3181
rect 8738 3173 8746 3181
rect 9170 3173 9178 3181
rect 9730 3173 9738 3181
rect 10034 3173 10042 3181
rect 10082 3173 10090 3181
rect 10482 3173 10490 3181
rect 13002 3179 13010 3187
rect 13242 3179 13250 3187
rect 13306 3179 13314 3187
rect 13338 3179 13346 3187
rect 14106 3179 14114 3187
rect 14794 3179 14802 3187
rect 15450 3179 15458 3187
rect 15834 3179 15842 3187
rect 21072 3180 21080 3188
rect 23296 3180 23304 3188
rect 24432 3180 24440 3188
rect 26336 3180 26344 3188
rect 27824 3180 27832 3188
rect 29856 3177 29864 3185
rect 31008 3177 31016 3185
rect 31360 3177 31368 3185
rect 32416 3177 32424 3185
rect 33120 3177 33128 3185
rect 34080 3177 34088 3185
rect 34208 3177 34216 3185
rect 34256 3177 34264 3185
rect 35936 3177 35944 3185
rect 36144 3177 36152 3185
rect 36224 3177 36232 3185
rect 36592 3177 36600 3185
rect 37056 3177 37064 3185
rect 37296 3177 37304 3185
rect 37504 3177 37512 3185
rect 37776 3177 37784 3185
rect 38128 3177 38136 3185
rect 38656 3177 38664 3185
rect 38832 3177 38840 3185
rect 38928 3177 38936 3185
rect 39104 3177 39112 3185
rect 39728 3177 39736 3185
rect 39888 3177 39896 3185
rect 39952 3177 39960 3185
rect 7106 3153 7114 3161
rect 7202 3153 7210 3161
rect 7378 3153 7386 3161
rect 9298 3153 9306 3161
rect 9458 3153 9466 3161
rect 9762 3153 9770 3161
rect 10018 3153 10026 3161
rect 12314 3159 12322 3167
rect 12506 3159 12514 3167
rect 12570 3159 12578 3167
rect 12698 3159 12706 3167
rect 12890 3159 12898 3167
rect 13498 3159 13506 3167
rect 13562 3159 13570 3167
rect 13770 3159 13778 3167
rect 14090 3159 14098 3167
rect 14442 3159 14450 3167
rect 14650 3159 14658 3167
rect 15322 3159 15330 3167
rect 15338 3159 15346 3167
rect 15434 3159 15442 3167
rect 15530 3159 15538 3167
rect 16906 3159 16914 3167
rect 17514 3159 17522 3167
rect 18640 3160 18648 3168
rect 19040 3161 19050 3166
rect 19424 3160 19432 3168
rect 20656 3160 20664 3168
rect 20880 3160 20888 3168
rect 22096 3160 22104 3168
rect 22320 3160 22328 3168
rect 22592 3160 22600 3168
rect 23008 3160 23016 3168
rect 23776 3160 23784 3168
rect 24272 3160 24280 3168
rect 24478 3161 24488 3166
rect 25040 3160 25048 3168
rect 25760 3160 25768 3168
rect 26160 3160 26168 3168
rect 26976 3160 26984 3168
rect 27886 3161 27896 3166
rect 28256 3160 28264 3168
rect 34352 3157 34360 3165
rect 5730 3133 5738 3141
rect 5874 3133 5882 3141
rect 5890 3133 5898 3141
rect 6034 3133 6042 3141
rect 6082 3133 6090 3141
rect 6114 3133 6122 3141
rect 6482 3133 6490 3141
rect 6498 3133 6506 3141
rect 6594 3133 6602 3141
rect 6626 3133 6634 3141
rect 6818 3133 6826 3141
rect 6866 3133 6874 3141
rect 6914 3133 6922 3141
rect 7682 3133 7690 3141
rect 7730 3133 7738 3141
rect 7746 3133 7754 3141
rect 8050 3133 8058 3141
rect 8130 3133 8138 3141
rect 8354 3133 8362 3141
rect 9074 3133 9082 3141
rect 9106 3133 9114 3141
rect 9778 3133 9786 3141
rect 9794 3133 9802 3141
rect 9858 3133 9866 3141
rect 10114 3133 10122 3141
rect 10162 3133 10170 3141
rect 10226 3133 10234 3141
rect 10354 3133 10362 3141
rect 10658 3133 10666 3141
rect 14682 3139 14690 3147
rect 14714 3139 14722 3147
rect 15050 3139 15058 3147
rect 15482 3139 15490 3147
rect 15530 3139 15538 3147
rect 16154 3139 16162 3147
rect 16234 3139 16242 3147
rect 16314 3139 16322 3147
rect 16330 3139 16338 3147
rect 16458 3139 16466 3147
rect 16522 3139 16530 3147
rect 16730 3139 16738 3147
rect 17114 3139 17122 3147
rect 17178 3139 17186 3147
rect 18464 3140 18472 3148
rect 25120 3140 25128 3148
rect 25344 3140 25352 3148
rect 25776 3140 25784 3148
rect 29424 3137 29432 3145
rect 29488 3137 29496 3145
rect 29584 3137 29592 3145
rect 29760 3137 29768 3145
rect 31024 3137 31032 3145
rect 31344 3137 31352 3145
rect 31824 3137 31832 3145
rect 31904 3137 31912 3145
rect 33008 3137 33016 3145
rect 33888 3137 33896 3145
rect 34224 3137 34232 3145
rect 35904 3137 35912 3145
rect 35936 3137 35944 3145
rect 36160 3137 36168 3145
rect 36368 3137 36376 3145
rect 36960 3137 36968 3145
rect 38320 3137 38328 3145
rect 38672 3137 38680 3145
rect 38848 3137 38856 3145
rect 40368 3137 40376 3145
rect 5986 3113 5994 3121
rect 6306 3113 6314 3121
rect 6658 3113 6666 3121
rect 6914 3113 6922 3121
rect 6978 3113 6986 3121
rect 8434 3113 8442 3121
rect 8466 3113 8474 3121
rect 8482 3113 8490 3121
rect 8674 3113 8682 3121
rect 9074 3113 9082 3121
rect 12234 3119 12242 3127
rect 12954 3119 12962 3127
rect 13594 3119 13602 3127
rect 13610 3119 13618 3127
rect 13834 3119 13842 3127
rect 14362 3119 14370 3127
rect 15882 3119 15890 3127
rect 17258 3119 17266 3127
rect 19216 3120 19224 3128
rect 19632 3120 19640 3128
rect 20240 3120 20248 3128
rect 21056 3120 21064 3128
rect 22080 3120 22088 3128
rect 23024 3120 23032 3128
rect 23312 3120 23320 3128
rect 23856 3120 23864 3128
rect 24192 3120 24200 3128
rect 24816 3120 24824 3128
rect 24848 3120 24856 3128
rect 26192 3120 26200 3128
rect 26400 3120 26408 3128
rect 26416 3120 26424 3128
rect 26960 3120 26968 3128
rect 27168 3120 27176 3128
rect 28336 3120 28344 3128
rect 29888 3117 29896 3125
rect 30224 3117 30232 3125
rect 30400 3117 30408 3125
rect 32912 3117 32920 3125
rect 33152 3117 33160 3125
rect 33200 3117 33208 3125
rect 33312 3117 33320 3125
rect 33632 3117 33640 3125
rect 34624 3117 34632 3125
rect 34784 3117 34792 3125
rect 38384 3117 38392 3125
rect 38448 3117 38456 3125
rect 38576 3117 38584 3125
rect 39056 3117 39064 3125
rect 5778 3093 5786 3101
rect 6018 3093 6026 3101
rect 6434 3093 6442 3101
rect 6546 3093 6554 3101
rect 6690 3093 6698 3101
rect 6818 3093 6826 3101
rect 7362 3093 7370 3101
rect 7410 3093 7418 3101
rect 7490 3093 7498 3101
rect 7634 3093 7642 3101
rect 7810 3093 7818 3101
rect 8466 3093 8474 3101
rect 8690 3093 8698 3101
rect 8994 3093 9002 3101
rect 9058 3093 9066 3101
rect 9138 3093 9146 3101
rect 9282 3093 9290 3101
rect 9714 3093 9722 3101
rect 10050 3093 10058 3101
rect 10178 3093 10186 3101
rect 10194 3093 10202 3101
rect 10610 3093 10618 3101
rect 10658 3093 10666 3101
rect 10802 3093 10810 3101
rect 12170 3099 12178 3107
rect 12186 3099 12194 3107
rect 12282 3099 12290 3107
rect 12298 3099 12306 3107
rect 14010 3099 14018 3107
rect 14746 3099 14754 3107
rect 15290 3099 15298 3107
rect 15338 3099 15346 3107
rect 15706 3099 15714 3107
rect 16778 3099 16786 3107
rect 16986 3099 16994 3107
rect 19488 3100 19496 3108
rect 20448 3100 20456 3108
rect 21280 3100 21288 3108
rect 21728 3100 21736 3108
rect 22096 3100 22104 3108
rect 23408 3100 23416 3108
rect 24624 3100 24632 3108
rect 24640 3100 24648 3108
rect 25312 3100 25320 3108
rect 30192 3097 30200 3105
rect 30496 3097 30504 3105
rect 31712 3097 31720 3105
rect 31872 3097 31880 3105
rect 35920 3097 35928 3105
rect 36096 3097 36104 3105
rect 36288 3097 36296 3105
rect 36800 3097 36808 3105
rect 37104 3097 37112 3105
rect 37120 3097 37128 3105
rect 37136 3097 37144 3105
rect 37168 3097 37176 3105
rect 38048 3097 38056 3105
rect 39232 3097 39240 3105
rect 39632 3097 39640 3105
rect 6786 3073 6794 3081
rect 6802 3073 6810 3081
rect 8210 3073 8218 3081
rect 8306 3073 8314 3081
rect 8802 3073 8810 3081
rect 8946 3073 8954 3081
rect 9698 3073 9706 3081
rect 9890 3073 9898 3081
rect 10018 3073 10026 3081
rect 10322 3073 10330 3081
rect 12618 3079 12626 3087
rect 12746 3079 12754 3087
rect 13754 3079 13762 3087
rect 13962 3079 13970 3087
rect 15338 3079 15346 3087
rect 16074 3079 16082 3087
rect 17034 3079 17042 3087
rect 17050 3079 17058 3087
rect 19248 3080 19256 3088
rect 22336 3080 22344 3088
rect 22784 3080 22792 3088
rect 24672 3080 24680 3088
rect 26560 3080 26568 3088
rect 28048 3080 28056 3088
rect 38976 3077 38984 3085
rect 39152 3077 39160 3085
rect 6258 3053 6266 3061
rect 8642 3053 8650 3061
rect 8818 3053 8826 3061
rect 9890 3053 9898 3061
rect 10370 3053 10378 3061
rect 10610 3053 10618 3061
rect 15642 3059 15650 3067
rect 16538 3059 16546 3067
rect 22768 3060 22776 3068
rect 27424 3060 27432 3068
rect 29460 3067 29472 3075
rect 29492 3067 29504 3075
rect 29508 3067 29520 3075
rect 29524 3067 29536 3075
rect 29552 3067 29564 3075
rect 29584 3067 29596 3075
rect 29600 3067 29612 3075
rect 29616 3067 29628 3075
rect 29648 3067 29660 3075
rect 29664 3067 29668 3075
rect 29772 3067 29784 3075
rect 29788 3067 29792 3075
rect 29804 3067 29816 3075
rect 29828 3067 29832 3075
rect 29836 3067 29848 3075
rect 29868 3067 29880 3075
rect 29952 3067 29956 3075
rect 29960 3067 29972 3075
rect 30044 3067 30048 3075
rect 30052 3067 30064 3075
rect 30084 3067 30096 3075
rect 30100 3067 30104 3075
rect 30176 3067 30188 3075
rect 30208 3067 30220 3075
rect 30224 3067 30228 3075
rect 30240 3067 30252 3075
rect 30260 3067 30284 3075
rect 30300 3067 30312 3075
rect 30316 3067 30320 3075
rect 30332 3067 30344 3075
rect 30352 3067 30376 3075
rect 30400 3067 30416 3075
rect 30424 3067 30440 3075
rect 30456 3067 30460 3075
rect 30464 3067 30468 3075
rect 30488 3067 30492 3075
rect 30496 3067 30508 3075
rect 30512 3067 30524 3075
rect 30528 3067 30532 3075
rect 30552 3067 30556 3075
rect 30560 3067 30564 3075
rect 30580 3067 30584 3075
rect 30588 3067 30600 3075
rect 30604 3067 30616 3075
rect 30620 3067 30624 3075
rect 30644 3067 30648 3075
rect 30652 3067 30656 3075
rect 30992 3067 30996 3075
rect 31000 3067 31004 3075
rect 31084 3067 31088 3075
rect 31092 3067 31096 3075
rect 31208 3067 31212 3075
rect 31216 3067 31220 3075
rect 31232 3067 31244 3075
rect 31248 3067 31252 3075
rect 31268 3067 31284 3075
rect 31300 3067 31348 3075
rect 31364 3067 31380 3075
rect 31396 3067 31408 3075
rect 31420 3067 31424 3075
rect 31428 3067 31440 3075
rect 31708 3067 31720 3075
rect 31724 3067 31736 3075
rect 31740 3067 31752 3075
rect 31772 3067 31784 3075
rect 31952 3067 31956 3075
rect 31960 3067 31972 3075
rect 31976 3067 31980 3075
rect 31992 3067 32000 3075
rect 32084 3067 32096 3075
rect 32116 3067 32128 3075
rect 32132 3067 32144 3075
rect 32148 3067 32160 3075
rect 32180 3067 32192 3075
rect 32200 3067 32232 3075
rect 32240 3067 32256 3075
rect 32272 3067 32296 3075
rect 32304 3067 32320 3075
rect 32336 3067 32340 3075
rect 32344 3067 32348 3075
rect 32360 3067 32372 3075
rect 32376 3067 32388 3075
rect 32396 3067 32412 3075
rect 32428 3067 32444 3075
rect 32452 3067 32464 3075
rect 32468 3067 32480 3075
rect 32492 3067 32496 3075
rect 32500 3067 32504 3075
rect 32632 3067 32636 3075
rect 32640 3067 32644 3075
rect 32656 3067 32668 3075
rect 32672 3067 32684 3075
rect 32696 3067 32700 3075
rect 32704 3067 32708 3075
rect 32724 3067 32740 3075
rect 32748 3067 32772 3075
rect 32788 3067 32800 3075
rect 32812 3067 32844 3075
rect 32852 3067 32868 3075
rect 32884 3067 32896 3075
rect 32904 3067 32936 3075
rect 32944 3067 32960 3075
rect 32976 3067 33000 3075
rect 33008 3067 33024 3075
rect 33040 3067 33056 3075
rect 33064 3067 33076 3075
rect 33080 3067 33092 3075
rect 33104 3067 33108 3075
rect 33112 3067 33116 3075
rect 33132 3067 33148 3075
rect 33156 3067 33168 3075
rect 33172 3067 33184 3075
rect 33192 3067 33208 3075
rect 33224 3067 33228 3075
rect 33232 3067 33236 3075
rect 33248 3067 33260 3075
rect 33264 3067 33276 3075
rect 33288 3067 33292 3075
rect 33296 3067 33300 3075
rect 33316 3067 33332 3075
rect 33340 3067 33364 3075
rect 33380 3067 33396 3075
rect 33412 3067 33424 3075
rect 33428 3067 33440 3075
rect 33444 3067 33456 3075
rect 33476 3067 33488 3075
rect 33492 3067 33496 3075
rect 33508 3067 33520 3075
rect 33536 3067 33552 3075
rect 33568 3067 33616 3075
rect 33632 3067 33644 3075
rect 33648 3067 33652 3075
rect 33664 3067 33676 3075
rect 33688 3067 33692 3075
rect 33696 3067 33708 3075
rect 33712 3067 33716 3075
rect 33820 3067 33832 3075
rect 33852 3067 33864 3075
rect 33868 3067 33880 3075
rect 33884 3067 33896 3075
rect 33912 3067 33928 3075
rect 33944 3067 33956 3075
rect 33960 3067 33972 3075
rect 33976 3067 33988 3075
rect 34008 3067 34020 3075
rect 34032 3067 34036 3075
rect 34040 3067 34052 3075
rect 34164 3067 34176 3075
rect 34188 3067 34192 3075
rect 34196 3067 34208 3075
rect 34212 3067 34216 3075
rect 34228 3067 34240 3075
rect 34252 3067 34256 3075
rect 34260 3067 34272 3075
rect 34288 3067 34312 3075
rect 34320 3067 34336 3075
rect 34352 3067 34356 3075
rect 34360 3067 34364 3075
rect 34384 3067 34388 3075
rect 34392 3067 34404 3075
rect 34408 3067 34420 3075
rect 34424 3067 34428 3075
rect 34448 3067 34452 3075
rect 34456 3067 34460 3075
rect 34508 3067 34512 3075
rect 34516 3067 34520 3075
rect 34632 3067 34636 3075
rect 34640 3067 34644 3075
rect 34656 3067 34668 3075
rect 34672 3067 34676 3075
rect 34696 3067 34700 3075
rect 34704 3067 34708 3075
rect 34724 3067 34772 3075
rect 34788 3067 34804 3075
rect 34820 3067 34832 3075
rect 34844 3067 34848 3075
rect 34852 3067 34864 3075
rect 34884 3067 34896 3075
rect 34900 3067 34904 3075
rect 34936 3067 34940 3075
rect 34944 3067 34956 3075
rect 34976 3067 34988 3075
rect 34992 3067 34996 3075
rect 35008 3067 35020 3075
rect 35036 3067 35052 3075
rect 35068 3067 35116 3075
rect 35132 3067 35148 3075
rect 35164 3067 35168 3075
rect 35172 3067 35184 3075
rect 35196 3067 35200 3075
rect 35204 3067 35208 3075
rect 35288 3067 35292 3075
rect 35296 3067 35300 3075
rect 35492 3067 35496 3075
rect 35500 3067 35504 3075
rect 35516 3067 35528 3075
rect 35532 3067 35536 3075
rect 35552 3067 35576 3075
rect 35584 3067 35600 3075
rect 35608 3067 35632 3075
rect 35648 3067 35664 3075
rect 35672 3067 35696 3075
rect 35712 3067 35724 3075
rect 35728 3067 35732 3075
rect 35744 3067 35756 3075
rect 35764 3067 35788 3075
rect 35804 3067 35828 3075
rect 35836 3067 35848 3075
rect 35856 3067 35880 3075
rect 35896 3067 35920 3075
rect 35928 3067 35944 3075
rect 35960 3067 35964 3075
rect 35968 3067 35972 3075
rect 35992 3067 35996 3075
rect 36000 3067 36012 3075
rect 36016 3067 36028 3075
rect 36032 3067 36036 3075
rect 36116 3067 36120 3075
rect 36124 3067 36128 3075
rect 36148 3067 36152 3075
rect 36156 3067 36160 3075
rect 36172 3067 36184 3075
rect 36188 3067 36192 3075
rect 36208 3067 36224 3075
rect 36240 3067 36288 3075
rect 36304 3067 36316 3075
rect 36332 3067 36380 3075
rect 36396 3067 36420 3075
rect 36428 3067 36440 3075
rect 36452 3067 36456 3075
rect 36460 3067 36472 3075
rect 36576 3067 36580 3075
rect 36584 3067 36596 3075
rect 36616 3067 36628 3075
rect 36632 3067 36636 3075
rect 36648 3067 36660 3075
rect 36680 3067 36692 3075
rect 36696 3067 36700 3075
rect 36712 3067 36724 3075
rect 36732 3067 36756 3075
rect 36772 3067 36784 3075
rect 36788 3067 36792 3075
rect 36804 3067 36816 3075
rect 36824 3067 36848 3075
rect 36864 3067 36888 3075
rect 36896 3067 36912 3075
rect 36928 3067 36952 3075
rect 36960 3067 36976 3075
rect 36984 3067 37008 3075
rect 37020 3067 37044 3075
rect 37052 3067 37068 3075
rect 37076 3067 37100 3075
rect 37116 3067 37128 3075
rect 37148 3067 37160 3075
rect 37172 3067 37176 3075
rect 37180 3067 37192 3075
rect 37196 3067 37200 3075
rect 37304 3067 37316 3075
rect 37428 3067 37440 3075
rect 37444 3067 37448 3075
rect 37460 3067 37472 3075
rect 37488 3067 37504 3075
rect 37512 3067 37544 3075
rect 37552 3067 37568 3075
rect 37576 3067 37600 3075
rect 37616 3067 37620 3075
rect 37624 3067 37636 3075
rect 37644 3067 37660 3075
rect 37668 3067 37692 3075
rect 37708 3067 37724 3075
rect 37732 3067 37756 3075
rect 37772 3067 37796 3075
rect 37804 3067 37816 3075
rect 37824 3067 37848 3075
rect 37864 3067 37888 3075
rect 37896 3067 37912 3075
rect 37928 3067 37944 3075
rect 37960 3067 37964 3075
rect 37968 3067 37980 3075
rect 37984 3067 37996 3075
rect 38000 3067 38004 3075
rect 38024 3067 38028 3075
rect 38032 3067 38036 3075
rect 38100 3067 38104 3075
rect 38108 3067 38112 3075
rect 38132 3067 38136 3075
rect 38140 3067 38144 3075
rect 38156 3067 38168 3075
rect 38172 3067 38176 3075
rect 38192 3067 38216 3075
rect 38224 3067 38240 3075
rect 38248 3067 38280 3075
rect 38288 3067 38300 3075
rect 38316 3067 38332 3075
rect 38340 3067 38372 3075
rect 38380 3067 38396 3075
rect 38412 3067 38416 3075
rect 38420 3067 38424 3075
rect 38444 3067 38448 3075
rect 38452 3067 38464 3075
rect 38476 3067 38480 3075
rect 38484 3067 38488 3075
rect 38500 3067 38512 3075
rect 38516 3067 38528 3075
rect 38536 3067 38552 3075
rect 38568 3067 38584 3075
rect 38592 3067 38616 3075
rect 38632 3067 38644 3075
rect 38664 3067 38676 3075
rect 38680 3067 38692 3075
rect 38696 3067 38708 3075
rect 38820 3067 38832 3075
rect 38844 3067 38848 3075
rect 38852 3067 38864 3075
rect 38868 3067 38872 3075
rect 38884 3067 38896 3075
rect 38912 3067 38928 3075
rect 38944 3067 38968 3075
rect 38976 3067 38992 3075
rect 39000 3067 39012 3075
rect 39016 3067 39020 3075
rect 39036 3067 39060 3075
rect 39068 3067 39084 3075
rect 39092 3067 39104 3075
rect 39108 3067 39112 3075
rect 39132 3067 39136 3075
rect 39140 3067 39152 3075
rect 39160 3067 39176 3075
rect 39184 3067 39196 3075
rect 39200 3067 39204 3075
rect 39224 3067 39228 3075
rect 39232 3067 39244 3075
rect 39256 3067 39260 3075
rect 39264 3067 39268 3075
rect 39364 3067 39368 3075
rect 39372 3067 39376 3075
rect 39488 3067 39492 3075
rect 39496 3067 39500 3075
rect 39596 3067 39600 3075
rect 39604 3067 39608 3075
rect 39620 3067 39632 3075
rect 39636 3067 39640 3075
rect 39660 3067 39664 3075
rect 39668 3067 39680 3075
rect 39692 3067 39696 3075
rect 39700 3067 39704 3075
rect 39800 3067 39804 3075
rect 39808 3067 39812 3075
rect 39832 3067 39836 3075
rect 39840 3067 39844 3075
rect 39924 3067 39928 3075
rect 39932 3067 39936 3075
rect 39948 3067 39960 3075
rect 39964 3067 39968 3075
rect 39988 3067 39992 3075
rect 39996 3067 40000 3075
rect 40016 3067 40064 3075
rect 40080 3067 40092 3075
rect 40108 3067 40156 3075
rect 40172 3067 40188 3075
rect 40196 3067 40220 3075
rect 40236 3067 40248 3075
rect 40268 3067 40280 3075
rect 40284 3067 40296 3075
rect 40300 3067 40312 3075
rect 40424 3067 40436 3075
rect 40440 3067 40452 3075
rect 40456 3067 40468 3075
rect 40488 3067 40500 3075
rect 40516 3067 40528 3075
rect 40532 3067 40544 3075
rect 40548 3067 40560 3075
rect 40580 3067 40592 3075
rect 40696 3067 40700 3075
rect 40704 3067 40716 3075
rect 40720 3067 40724 3075
rect 40736 3067 40748 3075
rect 40764 3067 40780 3075
rect 19944 3052 19946 3060
rect 21576 3050 21580 3058
rect 21666 3050 21674 3058
rect 22394 3050 22402 3058
rect 22544 3050 22550 3058
rect 23362 3050 23376 3058
rect 23432 3050 23440 3058
rect 23582 3050 23588 3058
rect 23882 3050 23886 3058
rect 23972 3050 23980 3058
rect 24390 3056 24392 3060
rect 24604 3056 24606 3060
rect 24396 3052 24398 3056
rect 24610 3052 24612 3056
rect 24700 3050 24708 3058
rect 24850 3050 24856 3058
rect 25364 3050 25368 3058
rect 25454 3050 25462 3058
rect 25658 3056 25660 3060
rect 25872 3056 25874 3060
rect 26086 3056 26088 3060
rect 26300 3056 26302 3060
rect 26514 3056 26516 3060
rect 26728 3056 26730 3060
rect 27086 3056 27088 3060
rect 25664 3052 25666 3056
rect 25878 3052 25880 3056
rect 26092 3052 26094 3056
rect 26306 3052 26308 3056
rect 26520 3052 26522 3056
rect 26734 3052 26736 3056
rect 27092 3052 27094 3056
rect 27290 3050 27294 3058
rect 27380 3050 27388 3058
rect 27798 3056 27800 3060
rect 28012 3056 28014 3060
rect 27804 3052 27806 3056
rect 28018 3052 28020 3056
rect 2936 3039 2944 3047
rect 6658 3033 6666 3041
rect 7858 3033 7866 3041
rect 7874 3033 7882 3041
rect 8626 3033 8634 3041
rect 8674 3033 8682 3041
rect 9250 3033 9258 3041
rect 9330 3033 9338 3041
rect 10290 3033 10298 3041
rect 13210 3039 13218 3047
rect 15194 3039 15202 3047
rect 15322 3039 15330 3047
rect 15962 3039 15970 3047
rect 17354 3039 17362 3047
rect 31632 3037 31640 3045
rect 31888 3037 31896 3045
rect 33872 3037 33880 3045
rect 33952 3037 33960 3045
rect 34336 3037 34344 3045
rect 34912 3037 34920 3045
rect 37584 3037 37592 3045
rect 37744 3037 37752 3045
rect 37856 3037 37864 3045
rect 38016 3037 38024 3045
rect 38096 3037 38104 3045
rect 40272 3037 40280 3045
rect 632 3019 640 3027
rect 936 3019 944 3027
rect 1272 3019 1280 3027
rect 2104 3019 2112 3027
rect 3144 3019 3152 3027
rect 3384 3019 3392 3027
rect 3800 3019 3808 3027
rect 4408 3019 4416 3027
rect 6002 3013 6010 3021
rect 6386 3013 6394 3021
rect 6722 3013 6730 3021
rect 6850 3013 6858 3021
rect 7170 3013 7178 3021
rect 9202 3013 9210 3021
rect 9906 3013 9914 3021
rect 12762 3019 12770 3027
rect 13498 3019 13506 3027
rect 13834 3019 13842 3027
rect 13882 3019 13890 3027
rect 14410 3019 14418 3027
rect 14666 3019 14674 3027
rect 14746 3019 14754 3027
rect 16538 3019 16546 3027
rect 16714 3019 16722 3027
rect 17162 3019 17170 3027
rect 17354 3019 17362 3027
rect 18464 3020 18472 3028
rect 18656 3020 18664 3028
rect 22160 3020 22168 3028
rect 22672 3020 22680 3028
rect 22800 3020 22808 3028
rect 25936 3020 25944 3028
rect 26176 3020 26184 3028
rect 28272 3020 28280 3028
rect 28656 3020 28664 3028
rect 29536 3017 29544 3025
rect 30928 3017 30936 3025
rect 32944 3017 32952 3025
rect 33936 3017 33944 3025
rect 34176 3017 34184 3025
rect 34448 3017 34456 3025
rect 35824 3017 35832 3025
rect 35904 3017 35912 3025
rect 36016 3017 36024 3025
rect 36320 3017 36328 3025
rect 37072 3017 37080 3025
rect 37264 3017 37272 3025
rect 37376 3017 37384 3025
rect 38592 3017 38600 3025
rect 38864 3017 38872 3025
rect 39024 3017 39032 3025
rect 40448 3017 40456 3025
rect 40512 3017 40520 3025
rect 40736 3017 40744 3025
rect 424 2999 432 3007
rect 552 2999 560 3007
rect 568 2999 576 3007
rect 648 2999 656 3007
rect 680 2999 688 3007
rect 840 2999 848 3007
rect 872 2999 880 3007
rect 952 2999 960 3007
rect 1112 2999 1120 3007
rect 1144 2999 1152 3007
rect 1368 2999 1376 3007
rect 1384 2999 1392 3007
rect 1512 2999 1520 3007
rect 1576 2999 1584 3007
rect 1784 2999 1792 3007
rect 1816 2999 1824 3007
rect 1848 2999 1856 3007
rect 1928 2999 1936 3007
rect 1944 2999 1952 3007
rect 2008 2999 2016 3007
rect 2120 2999 2128 3007
rect 2152 2999 2160 3007
rect 2184 2999 2192 3007
rect 2424 2999 2432 3007
rect 2536 2999 2544 3007
rect 2568 2999 2576 3007
rect 2632 2999 2640 3007
rect 2664 2999 2672 3007
rect 2776 2999 2784 3007
rect 2984 2999 2992 3007
rect 3080 2999 3088 3007
rect 3176 2999 3184 3007
rect 3240 2999 3248 3007
rect 3304 2999 3312 3007
rect 3400 2999 3408 3007
rect 3416 2999 3424 3007
rect 3576 2999 3584 3007
rect 3704 2999 3712 3007
rect 3944 2999 3952 3007
rect 3976 2999 3984 3007
rect 3992 2999 4000 3007
rect 4120 2999 4128 3007
rect 4248 2999 4256 3007
rect 4360 2999 4368 3007
rect 4376 2999 4384 3007
rect 4472 2999 4480 3007
rect 4552 2999 4560 3007
rect 4568 2999 4576 3007
rect 5890 2993 5898 3001
rect 6034 2993 6042 3001
rect 6162 2993 6170 3001
rect 6482 2993 6490 3001
rect 6706 2993 6714 3001
rect 6850 2993 6858 3001
rect 7154 2993 7162 3001
rect 7250 2993 7258 3001
rect 7970 2993 7978 3001
rect 8242 2993 8250 3001
rect 8338 2993 8346 3001
rect 8386 2993 8394 3001
rect 8434 2993 8442 3001
rect 8482 2993 8490 3001
rect 8498 2993 8506 3001
rect 8562 2993 8570 3001
rect 8610 2993 8618 3001
rect 9218 2993 9226 3001
rect 9618 2993 9626 3001
rect 10050 2993 10058 3001
rect 10210 2993 10218 3001
rect 10626 2993 10634 3001
rect 10770 2993 10778 3001
rect 13274 2999 13282 3007
rect 14986 2999 14994 3007
rect 16138 2999 16146 3007
rect 17146 2999 17154 3007
rect 19040 3000 19048 3008
rect 19680 3000 19688 3008
rect 21120 3000 21128 3008
rect 22592 3000 22600 3008
rect 26208 3000 26216 3008
rect 26352 3000 26360 3008
rect 26432 3000 26440 3008
rect 30384 2997 30392 3005
rect 30496 2997 30504 3005
rect 30608 2997 30616 3005
rect 30688 2997 30696 3005
rect 31216 2997 31224 3005
rect 31392 2997 31400 3005
rect 32144 2997 32152 3005
rect 32672 2997 32680 3005
rect 32832 2997 32840 3005
rect 33088 2997 33096 3005
rect 33360 2997 33368 3005
rect 33664 2997 33672 3005
rect 36080 2997 36088 3005
rect 36704 2997 36712 3005
rect 37152 2997 37160 3005
rect 37184 2997 37192 3005
rect 37248 2997 37256 3005
rect 37600 2997 37608 3005
rect 37744 2997 37752 3005
rect 37872 2997 37880 3005
rect 38224 2997 38232 3005
rect 38368 2997 38376 3005
rect 38432 2997 38440 3005
rect 39552 2997 39560 3005
rect 1176 2979 1184 2987
rect 1256 2979 1264 2987
rect 1560 2979 1568 2987
rect 2104 2979 2112 2987
rect 3368 2979 3376 2987
rect 3496 2979 3504 2987
rect 3640 2979 3648 2987
rect 3656 2979 3664 2987
rect 3704 2979 3712 2987
rect 3784 2979 3792 2987
rect 4040 2979 4048 2987
rect 5858 2973 5866 2981
rect 5970 2973 5978 2981
rect 6418 2973 6426 2981
rect 7346 2973 7354 2981
rect 7810 2973 7818 2981
rect 8226 2973 8234 2981
rect 8290 2973 8298 2981
rect 8338 2973 8346 2981
rect 8386 2973 8394 2981
rect 9042 2973 9050 2981
rect 9426 2973 9434 2981
rect 9810 2973 9818 2981
rect 9938 2973 9946 2981
rect 10450 2973 10458 2981
rect 10482 2973 10490 2981
rect 10578 2973 10586 2981
rect 12250 2979 12258 2987
rect 12394 2979 12402 2987
rect 12810 2979 12818 2987
rect 12938 2979 12946 2987
rect 13098 2979 13106 2987
rect 13338 2979 13346 2987
rect 13610 2979 13618 2987
rect 13770 2979 13778 2987
rect 13786 2979 13794 2987
rect 14058 2979 14066 2987
rect 14218 2979 14226 2987
rect 14714 2979 14722 2987
rect 16026 2979 16034 2987
rect 16522 2979 16530 2987
rect 16586 2979 16594 2987
rect 16618 2979 16626 2987
rect 16650 2979 16658 2987
rect 19216 2980 19224 2988
rect 19504 2980 19512 2988
rect 20032 2980 20040 2988
rect 20320 2980 20328 2988
rect 20864 2980 20872 2988
rect 23168 2980 23176 2988
rect 23392 2980 23400 2988
rect 24656 2980 24664 2988
rect 24736 2980 24744 2988
rect 26640 2980 26648 2988
rect 26848 2980 26856 2988
rect 27184 2980 27192 2988
rect 27408 2980 27416 2988
rect 33472 2977 33480 2985
rect 38128 2977 38136 2985
rect 39440 2977 39448 2985
rect 39536 2977 39544 2985
rect 39952 2977 39960 2985
rect 40064 2977 40072 2985
rect 40176 2977 40184 2985
rect 40208 2977 40216 2985
rect 872 2959 880 2967
rect 1176 2959 1184 2967
rect 2808 2959 2816 2967
rect 2824 2959 2832 2967
rect 3560 2959 3568 2967
rect 3688 2959 3696 2967
rect 3944 2959 3952 2967
rect 4152 2959 4160 2967
rect 5954 2953 5962 2961
rect 6258 2953 6266 2961
rect 6418 2953 6426 2961
rect 6530 2953 6538 2961
rect 7922 2953 7930 2961
rect 8002 2953 8010 2961
rect 8866 2953 8874 2961
rect 9250 2953 9258 2961
rect 9410 2953 9418 2961
rect 9426 2953 9434 2961
rect 9970 2953 9978 2961
rect 10066 2953 10074 2961
rect 10082 2953 10090 2961
rect 10274 2953 10282 2961
rect 10802 2953 10810 2961
rect 13322 2959 13330 2967
rect 15114 2959 15122 2967
rect 15578 2959 15586 2967
rect 15626 2959 15634 2967
rect 15674 2959 15682 2967
rect 16186 2959 16194 2967
rect 16202 2959 16210 2967
rect 16314 2959 16322 2967
rect 16330 2959 16338 2967
rect 16458 2959 16466 2967
rect 16858 2959 16866 2967
rect 16874 2959 16882 2967
rect 17034 2959 17042 2967
rect 17050 2959 17058 2967
rect 17226 2959 17234 2967
rect 25776 2960 25784 2968
rect 25792 2960 25800 2968
rect 30080 2957 30088 2965
rect 30192 2957 30200 2965
rect 31200 2957 31208 2965
rect 31984 2957 31992 2965
rect 32176 2957 32184 2965
rect 33104 2957 33112 2965
rect 33824 2957 33832 2965
rect 34048 2957 34056 2965
rect 37744 2957 37752 2965
rect 38272 2957 38280 2965
rect 38416 2957 38424 2965
rect 39280 2957 39288 2965
rect 19040 2948 19044 2953
rect 20672 2948 20676 2953
rect 26422 2948 26429 2953
rect 27195 2948 27202 2953
rect 504 2939 512 2947
rect 536 2939 544 2947
rect 664 2939 672 2947
rect 744 2939 752 2947
rect 888 2939 896 2947
rect 984 2939 992 2947
rect 1064 2939 1072 2947
rect 1320 2939 1328 2947
rect 1384 2939 1392 2947
rect 1528 2939 1536 2947
rect 2888 2939 2896 2947
rect 3016 2939 3024 2947
rect 4056 2939 4064 2947
rect 4248 2939 4256 2947
rect 4296 2939 4304 2947
rect 4568 2939 4576 2947
rect 6194 2933 6202 2941
rect 6386 2933 6394 2941
rect 6514 2933 6522 2941
rect 6578 2933 6586 2941
rect 6850 2933 6858 2941
rect 7170 2933 7178 2941
rect 7298 2933 7306 2941
rect 7314 2933 7322 2941
rect 7362 2933 7370 2941
rect 7586 2933 7594 2941
rect 8034 2933 8042 2941
rect 8866 2933 8874 2941
rect 8946 2933 8954 2941
rect 9042 2933 9050 2941
rect 9090 2933 9098 2941
rect 9842 2933 9850 2941
rect 9874 2933 9882 2941
rect 10018 2933 10026 2941
rect 10450 2933 10458 2941
rect 10850 2933 10858 2941
rect 11994 2939 12002 2947
rect 12010 2939 12018 2947
rect 12058 2939 12066 2947
rect 12330 2939 12338 2947
rect 13354 2939 13362 2947
rect 14090 2939 14098 2947
rect 14730 2939 14738 2947
rect 14874 2939 14882 2947
rect 15002 2939 15010 2947
rect 15098 2939 15106 2947
rect 15290 2939 15298 2947
rect 15370 2939 15378 2947
rect 15466 2939 15474 2947
rect 15594 2939 15602 2947
rect 15802 2939 15810 2947
rect 16042 2939 16050 2947
rect 16698 2939 16706 2947
rect 18832 2940 18840 2948
rect 19232 2940 19240 2948
rect 19424 2940 19432 2948
rect 19504 2940 19512 2948
rect 21072 2940 21080 2948
rect 21744 2940 21752 2948
rect 22368 2940 22376 2948
rect 23184 2940 23192 2948
rect 23808 2940 23816 2948
rect 24496 2940 24504 2948
rect 25072 2940 25080 2948
rect 25552 2940 25560 2948
rect 25776 2940 25784 2948
rect 25888 2940 25896 2948
rect 26208 2940 26216 2948
rect 26272 2940 26280 2948
rect 27440 2940 27448 2948
rect 27920 2940 27928 2948
rect 28112 2940 28120 2948
rect 35680 2937 35688 2945
rect 1096 2919 1104 2927
rect 1976 2919 1984 2927
rect 3544 2919 3552 2927
rect 4136 2919 4144 2927
rect 4168 2919 4176 2927
rect 7058 2913 7066 2921
rect 7122 2913 7130 2921
rect 7250 2913 7258 2921
rect 7346 2913 7354 2921
rect 7490 2913 7498 2921
rect 7522 2913 7530 2921
rect 7634 2913 7642 2921
rect 7714 2913 7722 2921
rect 7778 2913 7786 2921
rect 8146 2913 8154 2921
rect 8722 2913 8730 2921
rect 10162 2913 10170 2921
rect 10370 2913 10378 2921
rect 12426 2919 12434 2927
rect 14682 2919 14690 2927
rect 20256 2920 20264 2928
rect 25440 2920 25448 2928
rect 33920 2917 33928 2925
rect 35200 2917 35208 2925
rect 1688 2899 1696 2907
rect 1944 2899 1952 2907
rect 2328 2899 2336 2907
rect 2856 2899 2864 2907
rect 6434 2893 6442 2901
rect 6498 2893 6506 2901
rect 6994 2893 7002 2901
rect 7346 2893 7354 2901
rect 7474 2893 7482 2901
rect 7618 2893 7626 2901
rect 15754 2899 15762 2907
rect 22112 2900 22120 2908
rect 22144 2900 22152 2908
rect 23392 2900 23400 2908
rect 24912 2900 24920 2908
rect 38720 2897 38728 2905
rect 776 2879 784 2887
rect 1672 2879 1680 2887
rect 1800 2879 1808 2887
rect 2344 2879 2352 2887
rect 3064 2879 3072 2887
rect 3224 2879 3232 2887
rect 3432 2879 3440 2887
rect 3928 2879 3936 2887
rect 4232 2879 4240 2887
rect 6178 2873 6186 2881
rect 6722 2873 6730 2881
rect 6898 2873 6906 2881
rect 8402 2873 8410 2881
rect 8546 2873 8554 2881
rect 10034 2873 10042 2881
rect 10226 2873 10234 2881
rect 13146 2879 13154 2887
rect 14298 2879 14306 2887
rect 15770 2879 15778 2887
rect 516 2863 540 2867
rect 3832 2859 3840 2867
rect 7330 2853 7338 2861
rect 8482 2853 8490 2861
rect 10386 2853 10394 2861
rect 27888 2860 27896 2868
rect 29396 2867 29408 2875
rect 29428 2867 29440 2875
rect 29444 2867 29448 2875
rect 29460 2867 29472 2875
rect 29492 2867 29504 2875
rect 29512 2867 29544 2875
rect 29552 2867 29564 2875
rect 29584 2867 29596 2875
rect 29600 2867 29612 2875
rect 29616 2867 29628 2875
rect 29644 2867 29660 2875
rect 29676 2867 29688 2875
rect 29692 2867 29704 2875
rect 29708 2867 29720 2875
rect 29740 2867 29752 2875
rect 29896 2867 29908 2875
rect 29928 2867 29940 2875
rect 29944 2867 29956 2875
rect 29960 2867 29972 2875
rect 29988 2867 30000 2875
rect 30020 2867 30032 2875
rect 30036 2867 30048 2875
rect 30052 2867 30064 2875
rect 30084 2867 30096 2875
rect 30112 2867 30124 2875
rect 30128 2867 30140 2875
rect 30144 2867 30156 2875
rect 30204 2867 30216 2875
rect 30220 2867 30232 2875
rect 30236 2867 30248 2875
rect 30296 2867 30308 2875
rect 30312 2867 30324 2875
rect 30328 2867 30340 2875
rect 30412 2867 30416 2875
rect 30420 2867 30432 2875
rect 30668 2867 30680 2875
rect 30684 2867 30688 2875
rect 30792 2867 30804 2875
rect 30808 2867 30820 2875
rect 30824 2867 30836 2875
rect 30852 2867 30868 2875
rect 30884 2867 30908 2875
rect 30916 2867 30932 2875
rect 30948 2867 30964 2875
rect 30972 2867 30984 2875
rect 30988 2867 31000 2875
rect 31008 2867 31024 2875
rect 31040 2867 31056 2875
rect 31064 2867 31076 2875
rect 31080 2867 31092 2875
rect 31100 2867 31116 2875
rect 31132 2867 31148 2875
rect 31156 2867 31168 2875
rect 31172 2867 31184 2875
rect 31196 2867 31200 2875
rect 31204 2867 31208 2875
rect 31228 2867 31232 2875
rect 31236 2867 31240 2875
rect 31336 2867 31340 2875
rect 31344 2867 31348 2875
rect 31360 2867 31372 2875
rect 31376 2867 31380 2875
rect 31400 2867 31404 2875
rect 31408 2867 31412 2875
rect 31432 2867 31436 2875
rect 31440 2867 31444 2875
rect 31464 2867 31468 2875
rect 31472 2867 31484 2875
rect 31496 2867 31500 2875
rect 31504 2867 31508 2875
rect 31520 2867 31532 2875
rect 31536 2867 31548 2875
rect 31560 2867 31564 2875
rect 31568 2867 31572 2875
rect 31584 2867 31596 2875
rect 31600 2867 31604 2875
rect 31620 2867 31624 2875
rect 31628 2867 31640 2875
rect 31652 2867 31656 2875
rect 31660 2867 31664 2875
rect 31676 2867 31688 2875
rect 31692 2867 31696 2875
rect 31712 2867 31716 2875
rect 31720 2867 31732 2875
rect 31744 2867 31748 2875
rect 31752 2867 31756 2875
rect 31768 2867 31780 2875
rect 31784 2867 31788 2875
rect 31804 2867 31820 2875
rect 31836 2867 31852 2875
rect 31860 2867 31892 2875
rect 31900 2867 31916 2875
rect 31932 2867 31944 2875
rect 31948 2867 31960 2875
rect 31964 2867 31976 2875
rect 32000 2867 32008 2875
rect 32024 2867 32036 2875
rect 32040 2867 32052 2875
rect 32056 2867 32068 2875
rect 32084 2867 32100 2875
rect 32116 2867 32128 2875
rect 32132 2867 32144 2875
rect 32148 2867 32160 2875
rect 32208 2867 32220 2875
rect 32224 2867 32236 2875
rect 32240 2867 32252 2875
rect 32324 2867 32328 2875
rect 32332 2867 32344 2875
rect 32364 2867 32376 2875
rect 32380 2867 32384 2875
rect 32396 2867 32408 2875
rect 32428 2867 32440 2875
rect 32456 2867 32504 2875
rect 32520 2867 32524 2875
rect 32528 2867 32532 2875
rect 32548 2867 32596 2875
rect 32612 2867 32628 2875
rect 32644 2867 32648 2875
rect 32652 2867 32664 2875
rect 32676 2867 32680 2875
rect 32684 2867 32688 2875
rect 32708 2867 32712 2875
rect 32716 2867 32720 2875
rect 32768 2867 32772 2875
rect 32776 2867 32780 2875
rect 32800 2867 32804 2875
rect 32808 2867 32820 2875
rect 32824 2867 32836 2875
rect 32840 2867 32844 2875
rect 32860 2867 32876 2875
rect 32892 2867 32896 2875
rect 32900 2867 32912 2875
rect 32916 2867 32928 2875
rect 32932 2867 32936 2875
rect 32956 2867 32960 2875
rect 32964 2867 32968 2875
rect 32988 2867 32992 2875
rect 32996 2867 33000 2875
rect 33020 2867 33024 2875
rect 33028 2867 33032 2875
rect 33052 2867 33056 2875
rect 33060 2867 33072 2875
rect 33076 2867 33088 2875
rect 33092 2867 33096 2875
rect 33116 2867 33120 2875
rect 33124 2867 33128 2875
rect 33144 2867 33148 2875
rect 33152 2867 33164 2875
rect 33168 2867 33180 2875
rect 33184 2867 33188 2875
rect 33316 2867 33320 2875
rect 33324 2867 33336 2875
rect 33340 2867 33352 2875
rect 33356 2867 33360 2875
rect 33408 2867 33412 2875
rect 33416 2867 33428 2875
rect 33432 2867 33444 2875
rect 33448 2867 33452 2875
rect 33472 2867 33476 2875
rect 33480 2867 33492 2875
rect 33504 2867 33508 2875
rect 33512 2867 33516 2875
rect 33536 2867 33540 2875
rect 33544 2867 33548 2875
rect 33568 2867 33572 2875
rect 33576 2867 33580 2875
rect 33592 2867 33604 2875
rect 33608 2867 33612 2875
rect 33628 2867 33652 2875
rect 33660 2867 33676 2875
rect 33684 2867 33708 2875
rect 33724 2867 33736 2875
rect 33756 2867 33768 2875
rect 33780 2867 33784 2875
rect 33788 2867 33800 2875
rect 33804 2867 33808 2875
rect 33872 2867 33876 2875
rect 33880 2867 33892 2875
rect 33896 2867 33900 2875
rect 33940 2867 33952 2875
rect 33964 2867 33968 2875
rect 33972 2867 33984 2875
rect 33988 2867 33992 2875
rect 34004 2867 34016 2875
rect 34032 2867 34048 2875
rect 34064 2867 34088 2875
rect 34096 2867 34112 2875
rect 34120 2867 34132 2875
rect 34136 2867 34140 2875
rect 34160 2867 34164 2875
rect 34168 2867 34180 2875
rect 34184 2867 34196 2875
rect 34200 2867 34204 2875
rect 34300 2867 34304 2875
rect 34308 2867 34312 2875
rect 34332 2867 34336 2875
rect 34340 2867 34344 2875
rect 34356 2867 34368 2875
rect 34372 2867 34376 2875
rect 34400 2867 34416 2875
rect 34424 2867 34440 2875
rect 34448 2867 34480 2875
rect 34488 2867 34504 2875
rect 34520 2867 34524 2875
rect 34528 2867 34532 2875
rect 34552 2867 34556 2875
rect 34560 2867 34572 2875
rect 34584 2867 34588 2875
rect 34592 2867 34596 2875
rect 34608 2867 34620 2875
rect 34624 2867 34628 2875
rect 34644 2867 34648 2875
rect 34652 2867 34664 2875
rect 34676 2867 34680 2875
rect 34684 2867 34688 2875
rect 34700 2867 34712 2875
rect 34716 2867 34720 2875
rect 34736 2867 34740 2875
rect 34744 2867 34756 2875
rect 34768 2867 34772 2875
rect 34776 2867 34780 2875
rect 34792 2867 34804 2875
rect 34808 2867 34812 2875
rect 34908 2867 34912 2875
rect 34916 2867 34920 2875
rect 34932 2867 34944 2875
rect 34948 2867 34960 2875
rect 34972 2867 34976 2875
rect 34980 2867 34984 2875
rect 35080 2867 35084 2875
rect 35088 2867 35100 2875
rect 35112 2867 35116 2875
rect 35120 2867 35124 2875
rect 35136 2867 35148 2875
rect 35152 2867 35156 2875
rect 35172 2867 35188 2875
rect 35204 2867 35220 2875
rect 35228 2867 35260 2875
rect 35268 2867 35284 2875
rect 35300 2867 35304 2875
rect 35308 2867 35312 2875
rect 35332 2867 35336 2875
rect 35340 2867 35352 2875
rect 35364 2867 35368 2875
rect 35372 2867 35376 2875
rect 35388 2867 35400 2875
rect 35404 2867 35416 2875
rect 35428 2867 35432 2875
rect 35436 2867 35440 2875
rect 35460 2867 35464 2875
rect 35468 2867 35472 2875
rect 35492 2867 35496 2875
rect 35500 2867 35504 2875
rect 35524 2867 35528 2875
rect 35532 2867 35536 2875
rect 35548 2867 35560 2875
rect 35564 2867 35576 2875
rect 35588 2867 35592 2875
rect 35596 2867 35600 2875
rect 35612 2867 35624 2875
rect 35628 2867 35632 2875
rect 35652 2867 35656 2875
rect 35660 2867 35664 2875
rect 35676 2867 35688 2875
rect 35692 2867 35696 2875
rect 35716 2867 35720 2875
rect 35724 2867 35736 2875
rect 35748 2867 35752 2875
rect 35756 2867 35760 2875
rect 35856 2867 35860 2875
rect 35864 2867 35868 2875
rect 35888 2867 35892 2875
rect 35896 2867 35908 2875
rect 35912 2867 35924 2875
rect 35928 2867 35932 2875
rect 35948 2867 35952 2875
rect 35956 2867 35960 2875
rect 35980 2867 35984 2875
rect 35988 2867 36000 2875
rect 36004 2867 36016 2875
rect 36020 2867 36024 2875
rect 36040 2867 36064 2875
rect 36072 2867 36088 2875
rect 36096 2867 36120 2875
rect 36136 2867 36152 2875
rect 36168 2867 36184 2875
rect 36200 2867 36224 2875
rect 36232 2867 36248 2875
rect 36256 2867 36280 2875
rect 36296 2867 36300 2875
rect 36304 2867 36316 2875
rect 36324 2867 36340 2875
rect 36348 2867 36372 2875
rect 36388 2867 36392 2875
rect 36396 2867 36408 2875
rect 36412 2867 36424 2875
rect 36428 2867 36432 2875
rect 36452 2867 36456 2875
rect 36460 2867 36464 2875
rect 36484 2867 36488 2875
rect 36492 2867 36496 2875
rect 36516 2867 36520 2875
rect 36524 2867 36528 2875
rect 36548 2867 36552 2875
rect 36556 2867 36568 2875
rect 36572 2867 36584 2875
rect 36588 2867 36592 2875
rect 36720 2867 36724 2875
rect 36728 2867 36740 2875
rect 36744 2867 36756 2875
rect 36760 2867 36764 2875
rect 36780 2867 36784 2875
rect 36788 2867 36792 2875
rect 36812 2867 36816 2875
rect 36820 2867 36832 2875
rect 36836 2867 36848 2875
rect 36852 2867 36856 2875
rect 36872 2867 36888 2875
rect 36904 2867 36920 2875
rect 36928 2867 36952 2875
rect 36968 2867 36992 2875
rect 37000 2867 37012 2875
rect 37020 2867 37044 2875
rect 37060 2867 37084 2875
rect 37092 2867 37108 2875
rect 37124 2867 37128 2875
rect 37132 2867 37136 2875
rect 37156 2867 37160 2875
rect 37164 2867 37176 2875
rect 37180 2867 37192 2875
rect 37196 2867 37200 2875
rect 37248 2867 37252 2875
rect 37256 2867 37268 2875
rect 37272 2867 37284 2875
rect 37288 2867 37292 2875
rect 37340 2867 37344 2875
rect 37348 2867 37360 2875
rect 37364 2867 37376 2875
rect 37380 2867 37384 2875
rect 37404 2867 37408 2875
rect 37412 2867 37416 2875
rect 37436 2867 37440 2875
rect 37444 2867 37448 2875
rect 37468 2867 37472 2875
rect 37476 2867 37480 2875
rect 37500 2867 37504 2875
rect 37508 2867 37520 2875
rect 37524 2867 37536 2875
rect 37540 2867 37544 2875
rect 37564 2867 37568 2875
rect 37572 2867 37584 2875
rect 37616 2867 37640 2875
rect 37656 2867 37660 2875
rect 37664 2867 37676 2875
rect 37680 2867 37692 2875
rect 37696 2867 37700 2875
rect 37720 2867 37724 2875
rect 37728 2867 37740 2875
rect 37744 2867 37756 2875
rect 37760 2867 37764 2875
rect 37784 2867 37788 2875
rect 37792 2867 37796 2875
rect 38004 2867 38008 2875
rect 38012 2867 38016 2875
rect 38036 2867 38040 2875
rect 38044 2867 38056 2875
rect 38060 2867 38072 2875
rect 38076 2867 38080 2875
rect 38100 2867 38104 2875
rect 38108 2867 38112 2875
rect 38132 2867 38136 2875
rect 38140 2867 38144 2875
rect 38164 2867 38168 2875
rect 38172 2867 38176 2875
rect 38196 2867 38200 2875
rect 38204 2867 38216 2875
rect 38220 2867 38232 2875
rect 38236 2867 38240 2875
rect 38256 2867 38280 2875
rect 38288 2867 38304 2875
rect 38312 2867 38324 2875
rect 38328 2867 38332 2875
rect 38352 2867 38356 2875
rect 38360 2867 38372 2875
rect 38380 2867 38396 2875
rect 38404 2867 38416 2875
rect 38420 2867 38424 2875
rect 38444 2867 38448 2875
rect 38452 2867 38464 2875
rect 38468 2867 38480 2875
rect 38484 2867 38488 2875
rect 38508 2867 38512 2875
rect 38516 2867 38528 2875
rect 38536 2867 38552 2875
rect 38560 2867 38584 2875
rect 38600 2867 38616 2875
rect 38632 2867 38644 2875
rect 38656 2867 38660 2875
rect 38664 2867 38676 2875
rect 38680 2867 38684 2875
rect 38696 2867 38708 2875
rect 38728 2867 38740 2875
rect 38760 2867 38772 2875
rect 38792 2867 38804 2875
rect 38816 2867 38820 2875
rect 38824 2867 38836 2875
rect 38840 2867 38844 2875
rect 38856 2867 38868 2875
rect 38880 2867 38884 2875
rect 38888 2867 38900 2875
rect 39004 2867 39008 2875
rect 39012 2867 39024 2875
rect 39168 2867 39180 2875
rect 39184 2867 39188 2875
rect 39200 2867 39212 2875
rect 39224 2867 39228 2875
rect 39232 2867 39244 2875
rect 39264 2867 39276 2875
rect 39288 2867 39292 2875
rect 39296 2867 39308 2875
rect 39328 2867 39340 2875
rect 39344 2867 39348 2875
rect 39380 2867 39384 2875
rect 39388 2867 39400 2875
rect 39420 2867 39432 2875
rect 39436 2867 39448 2875
rect 39452 2867 39464 2875
rect 39512 2867 39524 2875
rect 39528 2867 39540 2875
rect 39544 2867 39556 2875
rect 39576 2867 39588 2875
rect 39604 2867 39616 2875
rect 39620 2867 39632 2875
rect 39636 2867 39648 2875
rect 39668 2867 39680 2875
rect 39784 2867 39788 2875
rect 39792 2867 39804 2875
rect 39808 2867 39812 2875
rect 39824 2867 39836 2875
rect 39852 2867 39864 2875
rect 39876 2867 39880 2875
rect 39884 2867 39896 2875
rect 39900 2867 39904 2875
rect 39916 2867 39928 2875
rect 39944 2867 39960 2875
rect 39976 2867 40000 2875
rect 40008 2867 40024 2875
rect 40032 2867 40064 2875
rect 40072 2867 40088 2875
rect 40104 2867 40116 2875
rect 40124 2867 40156 2875
rect 40164 2867 40180 2875
rect 40196 2867 40212 2875
rect 40228 2867 40244 2875
rect 40260 2867 40276 2875
rect 40284 2867 40316 2875
rect 40324 2867 40340 2875
rect 40348 2867 40360 2875
rect 40364 2867 40368 2875
rect 40388 2867 40392 2875
rect 40396 2867 40408 2875
rect 40416 2867 40432 2875
rect 40440 2867 40464 2875
rect 40480 2867 40484 2875
rect 40488 2867 40500 2875
rect 40508 2867 40524 2875
rect 40532 2867 40556 2875
rect 40572 2867 40588 2875
rect 40604 2867 40620 2875
rect 40636 2867 40660 2875
rect 40668 2867 40684 2875
rect 40692 2867 40724 2875
rect 40732 2867 40748 2875
rect 40764 2867 40780 2875
rect 18472 2848 18476 2860
rect 19560 2850 19562 2858
rect 19568 2850 19570 2858
rect 20598 2850 20600 2858
rect 20606 2850 20608 2858
rect 21216 2850 21226 2858
rect 21858 2850 21868 2858
rect 22286 2850 22296 2858
rect 22714 2850 22724 2858
rect 24126 2850 24130 2858
rect 24134 2850 24138 2858
rect 24554 2850 24558 2858
rect 24562 2850 24566 2858
rect 24768 2850 24772 2858
rect 24776 2850 24780 2858
rect 25196 2850 25200 2858
rect 25204 2850 25208 2858
rect 25830 2850 25842 2858
rect 26044 2850 26056 2858
rect 26686 2850 26698 2858
rect 26900 2850 26912 2858
rect 27220 2850 27232 2858
rect 27542 2850 27554 2858
rect 27962 2850 27966 2858
rect 27970 2850 27974 2858
rect 28168 2850 28180 2858
rect 28382 2850 28394 2858
rect 4616 2839 4624 2847
rect 8754 2833 8762 2841
rect 10898 2833 10906 2841
rect 12762 2839 12770 2847
rect 13786 2839 13794 2847
rect 14026 2839 14034 2847
rect 15850 2839 15858 2847
rect 28320 2840 28328 2848
rect 1064 2819 1072 2827
rect 1304 2819 1312 2827
rect 1592 2819 1600 2827
rect 1720 2819 1728 2827
rect 2200 2819 2208 2827
rect 2504 2819 2512 2827
rect 2632 2819 2640 2827
rect 3128 2819 3136 2827
rect 3160 2819 3168 2827
rect 4472 2819 4480 2827
rect 4504 2819 4512 2827
rect 4536 2819 4544 2827
rect 6530 2813 6538 2821
rect 7554 2813 7562 2821
rect 7634 2813 7642 2821
rect 7794 2813 7802 2821
rect 8674 2813 8682 2821
rect 8994 2813 9002 2821
rect 9362 2813 9370 2821
rect 14026 2819 14034 2827
rect 15050 2819 15058 2827
rect 26864 2820 26872 2828
rect 32736 2817 32744 2825
rect 37568 2817 37576 2825
rect 38416 2817 38424 2825
rect 1864 2799 1872 2807
rect 2824 2799 2832 2807
rect 4248 2799 4256 2807
rect 4568 2799 4576 2807
rect 9874 2793 9882 2801
rect 9906 2793 9914 2801
rect 12826 2799 12834 2807
rect 13178 2799 13186 2807
rect 13594 2799 13602 2807
rect 15434 2799 15442 2807
rect 15450 2799 15458 2807
rect 16138 2799 16146 2807
rect 16186 2799 16194 2807
rect 16410 2799 16418 2807
rect 23120 2800 23128 2808
rect 24592 2800 24600 2808
rect 25296 2800 25304 2808
rect 31424 2797 31432 2805
rect 34144 2797 34152 2805
rect 1432 2779 1440 2787
rect 2120 2779 2128 2787
rect 2856 2779 2864 2787
rect 6210 2773 6218 2781
rect 7506 2773 7514 2781
rect 7810 2773 7818 2781
rect 7906 2773 7914 2781
rect 8034 2773 8042 2781
rect 8658 2773 8666 2781
rect 8674 2773 8682 2781
rect 8738 2773 8746 2781
rect 10482 2773 10490 2781
rect 10626 2773 10634 2781
rect 10866 2773 10874 2781
rect 16266 2779 16274 2787
rect 16650 2779 16658 2787
rect 23264 2780 23272 2788
rect 26480 2780 26488 2788
rect 29488 2777 29496 2785
rect 33120 2777 33128 2785
rect 33376 2777 33384 2785
rect 34048 2777 34056 2785
rect 34144 2777 34152 2785
rect 34576 2777 34584 2785
rect 34752 2777 34760 2785
rect 35904 2777 35912 2785
rect 36352 2777 36360 2785
rect 36688 2777 36696 2785
rect 38224 2777 38232 2785
rect 38352 2777 38360 2785
rect 38592 2777 38600 2785
rect 39744 2777 39752 2785
rect 39872 2777 39880 2785
rect 40432 2777 40440 2785
rect 536 2759 544 2767
rect 824 2759 832 2767
rect 1128 2759 1136 2767
rect 1368 2759 1376 2767
rect 1768 2759 1776 2767
rect 1896 2759 1904 2767
rect 1944 2759 1952 2767
rect 2936 2759 2944 2767
rect 3048 2759 3056 2767
rect 3192 2759 3200 2767
rect 3288 2759 3296 2767
rect 3416 2759 3424 2767
rect 3640 2759 3648 2767
rect 3880 2759 3888 2767
rect 4008 2759 4016 2767
rect 4072 2759 4080 2767
rect 4136 2759 4144 2767
rect 4168 2759 4176 2767
rect 4264 2759 4272 2767
rect 4312 2759 4320 2767
rect 5730 2753 5738 2761
rect 5954 2753 5962 2761
rect 6626 2753 6634 2761
rect 6706 2753 6714 2761
rect 6802 2753 6810 2761
rect 7010 2753 7018 2761
rect 7074 2753 7082 2761
rect 8226 2753 8234 2761
rect 8818 2753 8826 2761
rect 8930 2753 8938 2761
rect 9026 2753 9034 2761
rect 9074 2753 9082 2761
rect 9106 2753 9114 2761
rect 9154 2753 9162 2761
rect 9266 2753 9274 2761
rect 9282 2753 9290 2761
rect 9634 2753 9642 2761
rect 9778 2753 9786 2761
rect 9810 2753 9818 2761
rect 10818 2753 10826 2761
rect 12138 2759 12146 2767
rect 13418 2759 13426 2767
rect 14218 2759 14226 2767
rect 14410 2759 14418 2767
rect 14826 2759 14834 2767
rect 14874 2759 14882 2767
rect 14986 2759 14994 2767
rect 15082 2759 15090 2767
rect 15210 2759 15218 2767
rect 15258 2759 15266 2767
rect 15402 2759 15410 2767
rect 15530 2759 15538 2767
rect 15578 2759 15586 2767
rect 16234 2759 16242 2767
rect 16778 2759 16786 2767
rect 16794 2759 16802 2767
rect 16810 2759 16818 2767
rect 16858 2759 16866 2767
rect 17434 2759 17442 2767
rect 17498 2759 17506 2767
rect 18832 2760 18840 2768
rect 18864 2760 18872 2768
rect 19040 2761 19050 2766
rect 19634 2761 19644 2766
rect 19888 2760 19896 2768
rect 20320 2760 20328 2768
rect 20528 2760 20536 2768
rect 21152 2760 21160 2768
rect 21520 2760 21528 2768
rect 21808 2760 21816 2768
rect 22448 2760 22456 2768
rect 22880 2760 22888 2768
rect 23424 2760 23432 2768
rect 24144 2760 24152 2768
rect 24496 2760 24504 2768
rect 24790 2761 24791 2766
rect 25216 2760 25224 2768
rect 26064 2760 26072 2768
rect 26704 2760 26712 2768
rect 27568 2760 27576 2768
rect 28192 2760 28200 2768
rect 32896 2757 32904 2765
rect 34176 2757 34184 2765
rect 34864 2757 34872 2765
rect 1416 2739 1424 2747
rect 6914 2733 6922 2741
rect 7218 2733 7226 2741
rect 7234 2733 7242 2741
rect 7330 2733 7338 2741
rect 9586 2733 9594 2741
rect 9602 2733 9610 2741
rect 10258 2733 10266 2741
rect 10386 2733 10394 2741
rect 10434 2733 10442 2741
rect 10626 2733 10634 2741
rect 12314 2739 12322 2747
rect 12538 2739 12546 2747
rect 12762 2739 12770 2747
rect 13914 2739 13922 2747
rect 13930 2739 13938 2747
rect 14010 2739 14018 2747
rect 14762 2739 14770 2747
rect 15594 2739 15602 2747
rect 15690 2739 15698 2747
rect 15722 2739 15730 2747
rect 15946 2739 15954 2747
rect 16042 2739 16050 2747
rect 16538 2739 16546 2747
rect 16602 2739 16610 2747
rect 17354 2739 17362 2747
rect 17466 2739 17474 2747
rect 19216 2740 19224 2748
rect 26864 2740 26872 2748
rect 26928 2740 26936 2748
rect 29680 2737 29688 2745
rect 30736 2737 30744 2745
rect 32064 2737 32072 2745
rect 32304 2737 32312 2745
rect 34336 2737 34344 2745
rect 34512 2737 34520 2745
rect 36816 2737 36824 2745
rect 36912 2737 36920 2745
rect 37536 2737 37544 2745
rect 38048 2737 38056 2745
rect 38560 2737 38568 2745
rect 39648 2737 39656 2745
rect 40496 2737 40504 2745
rect 792 2719 800 2727
rect 1240 2719 1248 2727
rect 1656 2719 1664 2727
rect 1848 2719 1856 2727
rect 2104 2719 2112 2727
rect 2504 2719 2512 2727
rect 2520 2719 2528 2727
rect 2616 2719 2624 2727
rect 3960 2719 3968 2727
rect 4056 2719 4064 2727
rect 4344 2719 4352 2727
rect 5826 2713 5834 2721
rect 6226 2713 6234 2721
rect 6418 2713 6426 2721
rect 6530 2713 6538 2721
rect 6658 2713 6666 2721
rect 6754 2713 6762 2721
rect 6866 2713 6874 2721
rect 7234 2713 7242 2721
rect 8098 2713 8106 2721
rect 8338 2713 8346 2721
rect 8562 2713 8570 2721
rect 8658 2713 8666 2721
rect 9874 2713 9882 2721
rect 9970 2713 9978 2721
rect 10018 2713 10026 2721
rect 10082 2713 10090 2721
rect 10098 2713 10106 2721
rect 10322 2713 10330 2721
rect 10690 2713 10698 2721
rect 10770 2713 10778 2721
rect 10802 2713 10810 2721
rect 10818 2713 10826 2721
rect 12074 2719 12082 2727
rect 12298 2719 12306 2727
rect 12634 2719 12642 2727
rect 13114 2719 13122 2727
rect 13466 2719 13474 2727
rect 13578 2719 13586 2727
rect 13626 2719 13634 2727
rect 13674 2719 13682 2727
rect 13770 2719 13778 2727
rect 14298 2719 14306 2727
rect 14346 2719 14354 2727
rect 14362 2719 14370 2727
rect 14490 2719 14498 2727
rect 14538 2719 14546 2727
rect 14554 2719 14562 2727
rect 14618 2719 14626 2727
rect 15482 2719 15490 2727
rect 15610 2719 15618 2727
rect 16394 2719 16402 2727
rect 16746 2719 16754 2727
rect 18816 2720 18824 2728
rect 19024 2720 19032 2728
rect 19248 2720 19256 2728
rect 19456 2720 19464 2728
rect 19616 2720 19624 2728
rect 20096 2720 20104 2728
rect 20544 2720 20552 2728
rect 21216 2720 21224 2728
rect 21504 2720 21512 2728
rect 21984 2720 21992 2728
rect 22368 2720 22376 2728
rect 22672 2720 22680 2728
rect 23728 2720 23736 2728
rect 23744 2720 23752 2728
rect 23840 2720 23848 2728
rect 24160 2720 24168 2728
rect 24800 2720 24808 2728
rect 25008 2720 25016 2728
rect 25232 2720 25240 2728
rect 25408 2720 25416 2728
rect 25440 2720 25448 2728
rect 26080 2720 26088 2728
rect 26416 2720 26424 2728
rect 27584 2720 27592 2728
rect 28320 2720 28328 2728
rect 29584 2717 29592 2725
rect 33072 2717 33080 2725
rect 33152 2717 33160 2725
rect 33296 2717 33304 2725
rect 33696 2717 33704 2725
rect 33728 2717 33736 2725
rect 34368 2717 34376 2725
rect 34528 2717 34536 2725
rect 34560 2717 34568 2725
rect 36096 2717 36104 2725
rect 36112 2717 36120 2725
rect 37056 2717 37064 2725
rect 37280 2717 37288 2725
rect 37472 2717 37480 2725
rect 37600 2717 37608 2725
rect 37792 2717 37800 2725
rect 37968 2717 37976 2725
rect 38448 2717 38456 2725
rect 39168 2717 39176 2725
rect 40032 2717 40040 2725
rect 40144 2717 40152 2725
rect 40304 2717 40312 2725
rect 40608 2717 40616 2725
rect 488 2699 496 2707
rect 504 2699 512 2707
rect 584 2699 592 2707
rect 904 2699 912 2707
rect 936 2699 944 2707
rect 1048 2699 1056 2707
rect 1288 2699 1296 2707
rect 1320 2699 1328 2707
rect 1384 2699 1392 2707
rect 1416 2699 1424 2707
rect 1576 2699 1584 2707
rect 1704 2699 1712 2707
rect 1880 2699 1888 2707
rect 1960 2699 1968 2707
rect 1976 2699 1984 2707
rect 2072 2699 2080 2707
rect 2088 2699 2096 2707
rect 2136 2699 2144 2707
rect 2216 2699 2224 2707
rect 2232 2699 2240 2707
rect 2328 2699 2336 2707
rect 2408 2699 2416 2707
rect 2424 2699 2432 2707
rect 2520 2699 2528 2707
rect 2648 2699 2656 2707
rect 2664 2699 2672 2707
rect 2760 2699 2768 2707
rect 2808 2699 2816 2707
rect 2840 2699 2848 2707
rect 2872 2699 2880 2707
rect 2952 2699 2960 2707
rect 2984 2699 2992 2707
rect 3032 2699 3040 2707
rect 3112 2699 3120 2707
rect 3144 2699 3152 2707
rect 3176 2699 3184 2707
rect 3352 2699 3360 2707
rect 3368 2699 3376 2707
rect 3464 2699 3472 2707
rect 3544 2699 3552 2707
rect 3736 2699 3744 2707
rect 3816 2699 3824 2707
rect 4136 2699 4144 2707
rect 4232 2699 4240 2707
rect 4520 2699 4528 2707
rect 4552 2699 4560 2707
rect 5874 2693 5882 2701
rect 5890 2693 5898 2701
rect 5922 2693 5930 2701
rect 6018 2693 6026 2701
rect 6066 2693 6074 2701
rect 6226 2693 6234 2701
rect 6594 2693 6602 2701
rect 6866 2693 6874 2701
rect 6962 2693 6970 2701
rect 6978 2693 6986 2701
rect 7026 2693 7034 2701
rect 7490 2693 7498 2701
rect 7570 2693 7578 2701
rect 7650 2693 7658 2701
rect 7778 2693 7786 2701
rect 7810 2693 7818 2701
rect 7986 2693 7994 2701
rect 8146 2693 8154 2701
rect 8370 2693 8378 2701
rect 8402 2693 8410 2701
rect 8626 2693 8634 2701
rect 8690 2693 8698 2701
rect 8722 2693 8730 2701
rect 8930 2693 8938 2701
rect 9042 2693 9050 2701
rect 9346 2693 9354 2701
rect 9378 2693 9386 2701
rect 9426 2693 9434 2701
rect 9458 2693 9466 2701
rect 9890 2693 9898 2701
rect 10594 2693 10602 2701
rect 10722 2693 10730 2701
rect 12826 2699 12834 2707
rect 13050 2699 13058 2707
rect 14106 2699 14114 2707
rect 14186 2699 14194 2707
rect 15626 2699 15634 2707
rect 16650 2699 16658 2707
rect 16682 2699 16690 2707
rect 16730 2699 16738 2707
rect 21568 2700 21576 2708
rect 21696 2700 21704 2708
rect 23520 2700 23528 2708
rect 35320 2705 35321 2710
rect 29760 2697 29768 2705
rect 31152 2697 31160 2705
rect 33424 2697 33432 2705
rect 33568 2697 33576 2705
rect 34256 2697 34264 2705
rect 34528 2697 34536 2705
rect 35008 2697 35016 2705
rect 35056 2697 35064 2705
rect 35456 2697 35464 2705
rect 36512 2697 36520 2705
rect 456 2679 464 2687
rect 680 2679 688 2687
rect 936 2679 944 2687
rect 968 2679 976 2687
rect 1064 2679 1072 2687
rect 1400 2679 1408 2687
rect 1608 2679 1616 2687
rect 2072 2679 2080 2687
rect 2168 2679 2176 2687
rect 2184 2679 2192 2687
rect 2344 2679 2352 2687
rect 2440 2679 2448 2687
rect 2456 2679 2464 2687
rect 3848 2679 3856 2687
rect 6114 2673 6122 2681
rect 6290 2673 6298 2681
rect 6418 2673 6426 2681
rect 7074 2673 7082 2681
rect 7426 2673 7434 2681
rect 7490 2673 7498 2681
rect 7762 2673 7770 2681
rect 8242 2673 8250 2681
rect 8818 2673 8826 2681
rect 8850 2673 8858 2681
rect 9378 2673 9386 2681
rect 9570 2673 9578 2681
rect 10610 2673 10618 2681
rect 10674 2673 10682 2681
rect 10818 2673 10826 2681
rect 12250 2679 12258 2687
rect 12442 2679 12450 2687
rect 13274 2679 13282 2687
rect 13322 2679 13330 2687
rect 13898 2679 13906 2687
rect 14106 2679 14114 2687
rect 15034 2679 15042 2687
rect 16522 2679 16530 2687
rect 20720 2680 20728 2688
rect 20896 2680 20904 2688
rect 23680 2680 23688 2688
rect 26224 2680 26232 2688
rect 28128 2680 28136 2688
rect 33776 2677 33784 2685
rect 33888 2677 33896 2685
rect 37424 2677 37432 2685
rect 40144 2677 40152 2685
rect 40768 2677 40776 2685
rect 696 2659 704 2667
rect 1224 2659 1232 2667
rect 1320 2659 1328 2667
rect 2648 2659 2656 2667
rect 2856 2659 2864 2667
rect 2968 2659 2976 2667
rect 3384 2659 3392 2667
rect 7026 2653 7034 2661
rect 7186 2653 7194 2661
rect 7298 2653 7306 2661
rect 7346 2653 7354 2661
rect 7650 2653 7658 2661
rect 7714 2653 7722 2661
rect 7906 2653 7914 2661
rect 8146 2653 8154 2661
rect 9714 2653 9722 2661
rect 10146 2653 10154 2661
rect 10162 2653 10170 2661
rect 10178 2653 10186 2661
rect 12250 2659 12258 2667
rect 12362 2659 12370 2667
rect 18880 2660 18888 2668
rect 20496 2660 20504 2668
rect 21328 2660 21336 2668
rect 21584 2660 21592 2668
rect 22816 2660 22824 2668
rect 23248 2660 23256 2668
rect 27520 2660 27528 2668
rect 28576 2660 28584 2668
rect 29520 2667 29532 2675
rect 29536 2667 29540 2675
rect 29552 2667 29564 2675
rect 29584 2667 29596 2675
rect 29600 2667 29612 2675
rect 29616 2667 29628 2675
rect 29644 2667 29660 2675
rect 29668 2667 29700 2675
rect 29708 2667 29724 2675
rect 29732 2667 29756 2675
rect 29772 2667 29784 2675
rect 29804 2667 29816 2675
rect 29828 2667 29832 2675
rect 29836 2667 29848 2675
rect 29852 2667 29856 2675
rect 29868 2667 29880 2675
rect 29896 2667 29912 2675
rect 29928 2667 29952 2675
rect 29960 2667 29976 2675
rect 29984 2667 29996 2675
rect 30000 2667 30004 2675
rect 30020 2667 30044 2675
rect 30052 2667 30068 2675
rect 30076 2667 30100 2675
rect 30116 2667 30120 2675
rect 30124 2667 30136 2675
rect 30144 2667 30160 2675
rect 30168 2667 30192 2675
rect 30208 2667 30212 2675
rect 30216 2667 30228 2675
rect 30240 2667 30244 2675
rect 30248 2667 30252 2675
rect 30272 2667 30276 2675
rect 30280 2667 30284 2675
rect 30412 2667 30416 2675
rect 30420 2667 30424 2675
rect 30444 2667 30448 2675
rect 30452 2667 30464 2675
rect 30468 2667 30480 2675
rect 30484 2667 30488 2675
rect 30508 2667 30512 2675
rect 30516 2667 30520 2675
rect 30532 2667 30544 2675
rect 30548 2667 30552 2675
rect 30568 2667 30584 2675
rect 30600 2667 30648 2675
rect 30664 2667 30668 2675
rect 30672 2667 30676 2675
rect 30692 2667 30740 2675
rect 30756 2667 30780 2675
rect 30788 2667 30800 2675
rect 30812 2667 30816 2675
rect 30820 2667 30832 2675
rect 30976 2667 30988 2675
rect 30992 2667 30996 2675
rect 31008 2667 31020 2675
rect 31040 2667 31052 2675
rect 31068 2667 31116 2675
rect 31132 2667 31148 2675
rect 31156 2667 31168 2675
rect 31172 2667 31184 2675
rect 31196 2667 31200 2675
rect 31204 2667 31208 2675
rect 31224 2667 31240 2675
rect 31248 2667 31260 2675
rect 31264 2667 31276 2675
rect 31288 2667 31292 2675
rect 31296 2667 31300 2675
rect 31320 2667 31324 2675
rect 31328 2667 31332 2675
rect 31444 2667 31448 2675
rect 31452 2667 31456 2675
rect 31476 2667 31480 2675
rect 31484 2667 31488 2675
rect 31500 2667 31512 2675
rect 31516 2667 31528 2675
rect 31536 2667 31552 2675
rect 31568 2667 31616 2675
rect 31632 2667 31636 2675
rect 31640 2667 31644 2675
rect 31656 2667 31668 2675
rect 31672 2667 31684 2675
rect 31696 2667 31700 2675
rect 31704 2667 31708 2675
rect 31804 2667 31808 2675
rect 31812 2667 31824 2675
rect 31836 2667 31840 2675
rect 31844 2667 31848 2675
rect 31860 2667 31872 2675
rect 31876 2667 31880 2675
rect 31928 2667 31932 2675
rect 31936 2667 31940 2675
rect 31952 2667 31964 2675
rect 31968 2667 31972 2675
rect 31992 2667 31996 2675
rect 32000 2667 32004 2675
rect 32020 2667 32036 2675
rect 32044 2667 32076 2675
rect 32084 2667 32100 2675
rect 32116 2667 32128 2675
rect 32140 2667 32144 2675
rect 32148 2667 32160 2675
rect 32272 2667 32284 2675
rect 32296 2667 32300 2675
rect 32304 2667 32316 2675
rect 32320 2667 32324 2675
rect 32336 2667 32348 2675
rect 32360 2667 32364 2675
rect 32368 2667 32380 2675
rect 32400 2667 32412 2675
rect 32484 2667 32488 2675
rect 32492 2667 32504 2675
rect 32524 2667 32536 2675
rect 32540 2667 32544 2675
rect 32576 2667 32580 2675
rect 32584 2667 32596 2675
rect 32616 2667 32628 2675
rect 32632 2667 32636 2675
rect 32648 2667 32660 2675
rect 32680 2667 32692 2675
rect 32696 2667 32700 2675
rect 32712 2667 32724 2675
rect 32736 2667 32740 2675
rect 32744 2667 32756 2675
rect 32760 2667 32764 2675
rect 32804 2667 32816 2675
rect 32828 2667 32832 2675
rect 32836 2667 32848 2675
rect 32852 2667 32856 2675
rect 32992 2667 33004 2675
rect 33008 2667 33012 2675
rect 33024 2667 33036 2675
rect 33052 2667 33068 2675
rect 33076 2667 33108 2675
rect 33116 2667 33132 2675
rect 33148 2667 33160 2675
rect 33168 2667 33200 2675
rect 33208 2667 33224 2675
rect 33240 2667 33264 2675
rect 33272 2667 33288 2675
rect 33304 2667 33352 2675
rect 33368 2667 33380 2675
rect 33396 2667 33444 2675
rect 33460 2667 33476 2675
rect 33484 2667 33496 2675
rect 33500 2667 33512 2675
rect 33524 2667 33528 2675
rect 33532 2667 33536 2675
rect 33664 2667 33668 2675
rect 33672 2667 33676 2675
rect 33688 2667 33700 2675
rect 33704 2667 33708 2675
rect 33728 2667 33732 2675
rect 33736 2667 33740 2675
rect 33760 2667 33764 2675
rect 33768 2667 33772 2675
rect 33792 2667 33796 2675
rect 33800 2667 33812 2675
rect 33824 2667 33828 2675
rect 33832 2667 33836 2675
rect 33848 2667 33860 2675
rect 33864 2667 33868 2675
rect 33932 2667 33936 2675
rect 33940 2667 33944 2675
rect 33964 2667 33968 2675
rect 33972 2667 33976 2675
rect 33988 2667 34000 2675
rect 34004 2667 34016 2675
rect 34024 2667 34040 2675
rect 34056 2667 34060 2675
rect 34064 2667 34068 2675
rect 34080 2667 34092 2675
rect 34096 2667 34108 2675
rect 34116 2667 34132 2675
rect 34148 2667 34196 2675
rect 34212 2667 34224 2675
rect 34228 2667 34232 2675
rect 34244 2667 34256 2675
rect 34268 2667 34272 2675
rect 34276 2667 34288 2675
rect 34292 2667 34296 2675
rect 34400 2667 34412 2675
rect 34524 2667 34536 2675
rect 34540 2667 34544 2675
rect 34556 2667 34568 2675
rect 34588 2667 34600 2675
rect 34612 2667 34616 2675
rect 34620 2667 34632 2675
rect 34836 2667 34848 2675
rect 34868 2667 34880 2675
rect 34884 2667 34888 2675
rect 34900 2667 34912 2675
rect 34932 2667 34944 2675
rect 34952 2667 34984 2675
rect 34992 2667 35004 2675
rect 35024 2667 35036 2675
rect 35044 2667 35076 2675
rect 35084 2667 35096 2675
rect 35116 2667 35128 2675
rect 35136 2667 35168 2675
rect 35176 2667 35188 2675
rect 35208 2667 35220 2675
rect 35228 2667 35260 2675
rect 35268 2667 35284 2675
rect 35300 2667 35324 2675
rect 35332 2667 35348 2675
rect 35364 2667 35380 2675
rect 35388 2667 35400 2675
rect 35404 2667 35416 2675
rect 35428 2667 35432 2675
rect 35436 2667 35440 2675
rect 35460 2667 35464 2675
rect 35468 2667 35472 2675
rect 35568 2667 35572 2675
rect 35576 2667 35580 2675
rect 35592 2667 35604 2675
rect 35608 2667 35620 2675
rect 35628 2667 35644 2675
rect 35660 2667 35708 2675
rect 35724 2667 35740 2675
rect 35756 2667 35768 2675
rect 35780 2667 35784 2675
rect 35788 2667 35800 2675
rect 35820 2667 35832 2675
rect 35836 2667 35840 2675
rect 36036 2667 36048 2675
rect 36052 2667 36064 2675
rect 36068 2667 36080 2675
rect 36096 2667 36112 2675
rect 36128 2667 36152 2675
rect 36160 2667 36176 2675
rect 36192 2667 36208 2675
rect 36216 2667 36228 2675
rect 36232 2667 36244 2675
rect 36256 2667 36260 2675
rect 36264 2667 36268 2675
rect 36284 2667 36300 2675
rect 36308 2667 36320 2675
rect 36324 2667 36336 2675
rect 36348 2667 36352 2675
rect 36356 2667 36360 2675
rect 36376 2667 36424 2675
rect 36440 2667 36456 2675
rect 36472 2667 36488 2675
rect 36504 2667 36520 2675
rect 36536 2667 36584 2675
rect 36600 2667 36612 2675
rect 36616 2667 36620 2675
rect 36632 2667 36644 2675
rect 36656 2667 36660 2675
rect 36664 2667 36676 2675
rect 36696 2667 36708 2675
rect 36780 2667 36784 2675
rect 36788 2667 36800 2675
rect 36820 2667 36832 2675
rect 36836 2667 36848 2675
rect 36852 2667 36864 2675
rect 36880 2667 36896 2675
rect 36912 2667 36924 2675
rect 36928 2667 36940 2675
rect 36944 2667 36956 2675
rect 36976 2667 36988 2675
rect 37004 2667 37016 2675
rect 37020 2667 37032 2675
rect 37036 2667 37048 2675
rect 37068 2667 37080 2675
rect 37160 2667 37172 2675
rect 37184 2667 37188 2675
rect 37192 2667 37204 2675
rect 37208 2667 37212 2675
rect 37224 2667 37236 2675
rect 37276 2667 37280 2675
rect 37284 2667 37296 2675
rect 37300 2667 37304 2675
rect 37316 2667 37328 2675
rect 37368 2667 37372 2675
rect 37376 2667 37388 2675
rect 37392 2667 37396 2675
rect 37408 2667 37420 2675
rect 37440 2667 37452 2675
rect 37472 2667 37484 2675
rect 37504 2667 37516 2675
rect 37528 2667 37532 2675
rect 37536 2667 37548 2675
rect 37552 2667 37556 2675
rect 37568 2667 37580 2675
rect 37684 2667 37688 2675
rect 37692 2667 37704 2675
rect 37708 2667 37712 2675
rect 37724 2667 37736 2675
rect 37744 2667 37768 2675
rect 37784 2667 37808 2675
rect 37816 2667 37832 2675
rect 37848 2667 37852 2675
rect 37856 2667 37860 2675
rect 37880 2667 37884 2675
rect 37888 2667 37900 2675
rect 37904 2667 37916 2675
rect 37920 2667 37924 2675
rect 38004 2667 38008 2675
rect 38012 2667 38016 2675
rect 38036 2667 38040 2675
rect 38044 2667 38048 2675
rect 38256 2667 38260 2675
rect 38264 2667 38276 2675
rect 38288 2667 38292 2675
rect 38296 2667 38300 2675
rect 38312 2667 38324 2675
rect 38328 2667 38332 2675
rect 38352 2667 38356 2675
rect 38360 2667 38364 2675
rect 38380 2667 38396 2675
rect 38404 2667 38436 2675
rect 38444 2667 38460 2675
rect 38468 2667 38480 2675
rect 38484 2667 38488 2675
rect 38508 2667 38512 2675
rect 38516 2667 38528 2675
rect 38536 2667 38552 2675
rect 38560 2667 38572 2675
rect 38576 2667 38580 2675
rect 38600 2667 38604 2675
rect 38608 2667 38620 2675
rect 38628 2667 38644 2675
rect 38652 2667 38664 2675
rect 38668 2667 38672 2675
rect 38692 2667 38696 2675
rect 38700 2667 38712 2675
rect 38724 2667 38728 2675
rect 38732 2667 38736 2675
rect 38756 2667 38760 2675
rect 38764 2667 38768 2675
rect 38788 2667 38792 2675
rect 38796 2667 38800 2675
rect 38812 2667 38824 2675
rect 38828 2667 38832 2675
rect 38852 2667 38856 2675
rect 38860 2667 38872 2675
rect 38876 2667 38888 2675
rect 38892 2667 38896 2675
rect 38912 2667 38928 2675
rect 38944 2667 38948 2675
rect 38952 2667 38964 2675
rect 38968 2667 38980 2675
rect 38984 2667 38988 2675
rect 39004 2667 39008 2675
rect 39012 2667 39016 2675
rect 39036 2667 39040 2675
rect 39044 2667 39056 2675
rect 39060 2667 39072 2675
rect 39076 2667 39080 2675
rect 39208 2667 39212 2675
rect 39216 2667 39228 2675
rect 39232 2667 39244 2675
rect 39248 2667 39252 2675
rect 39272 2667 39276 2675
rect 39280 2667 39292 2675
rect 39296 2667 39308 2675
rect 39312 2667 39316 2675
rect 39336 2667 39340 2675
rect 39344 2667 39348 2675
rect 39476 2667 39480 2675
rect 39484 2667 39488 2675
rect 39600 2667 39604 2675
rect 39608 2667 39612 2675
rect 39692 2667 39696 2675
rect 39700 2667 39704 2675
rect 39716 2667 39728 2675
rect 39732 2667 39736 2675
rect 39756 2667 39760 2675
rect 39764 2667 39768 2675
rect 39784 2667 39832 2675
rect 39848 2667 39860 2675
rect 39880 2667 39892 2675
rect 39904 2667 39908 2675
rect 39912 2667 39924 2675
rect 40036 2667 40048 2675
rect 40052 2667 40064 2675
rect 40068 2667 40080 2675
rect 40100 2667 40112 2675
rect 40256 2667 40268 2675
rect 40288 2667 40300 2675
rect 40304 2667 40316 2675
rect 40320 2667 40332 2675
rect 40404 2667 40408 2675
rect 40412 2667 40424 2675
rect 40444 2667 40456 2675
rect 40460 2667 40464 2675
rect 40496 2667 40500 2675
rect 40504 2667 40516 2675
rect 40536 2667 40548 2675
rect 40552 2667 40556 2675
rect 40568 2667 40580 2675
rect 40596 2667 40612 2675
rect 40628 2667 40676 2675
rect 40692 2667 40696 2675
rect 40700 2667 40704 2675
rect 40716 2667 40728 2675
rect 40732 2667 40744 2675
rect 40756 2667 40760 2675
rect 40764 2667 40768 2675
rect 18932 2656 18934 2660
rect 18938 2652 18940 2656
rect 19098 2650 19106 2658
rect 19248 2650 19254 2658
rect 19582 2650 19588 2658
rect 19590 2650 19596 2658
rect 19780 2650 19786 2658
rect 19788 2650 19794 2658
rect 19874 2650 19880 2658
rect 20746 2650 20754 2658
rect 20896 2650 20902 2658
rect 21388 2650 21396 2658
rect 21538 2650 21544 2658
rect 21602 2650 21610 2658
rect 21752 2650 21758 2658
rect 23442 2650 23456 2658
rect 23962 2650 23966 2658
rect 24052 2650 24060 2658
rect 24256 2656 24258 2660
rect 24400 2656 24402 2660
rect 24684 2656 24686 2660
rect 24898 2656 24900 2660
rect 24262 2652 24264 2656
rect 24406 2652 24408 2656
rect 24690 2652 24692 2656
rect 24904 2652 24906 2656
rect 25032 2650 25036 2658
rect 25122 2650 25130 2658
rect 25326 2656 25328 2660
rect 25540 2656 25542 2660
rect 25968 2656 25970 2660
rect 25332 2652 25334 2656
rect 25546 2652 25548 2656
rect 25974 2652 25976 2656
rect 26102 2650 26106 2658
rect 26192 2650 26200 2658
rect 26744 2650 26748 2658
rect 26834 2650 26842 2658
rect 26958 2650 26962 2658
rect 27048 2650 27056 2658
rect 27182 2656 27184 2660
rect 27188 2652 27190 2656
rect 27386 2650 27390 2658
rect 27476 2650 27484 2658
rect 27680 2656 27682 2660
rect 30544 2657 30552 2665
rect 30944 2657 30952 2665
rect 32784 2657 32792 2665
rect 35616 2657 35624 2665
rect 37904 2657 37912 2665
rect 27686 2652 27688 2656
rect 1064 2639 1072 2647
rect 1976 2639 1984 2647
rect 2280 2639 2288 2647
rect 3512 2639 3520 2647
rect 3576 2639 3584 2647
rect 3592 2639 3600 2647
rect 3912 2639 3920 2647
rect 3928 2639 3936 2647
rect 4328 2639 4336 2647
rect 6466 2633 6474 2641
rect 6674 2633 6682 2641
rect 7506 2633 7514 2641
rect 7954 2633 7962 2641
rect 8258 2633 8266 2641
rect 8898 2633 8906 2641
rect 9746 2633 9754 2641
rect 9858 2633 9866 2641
rect 10290 2633 10298 2641
rect 10610 2633 10618 2641
rect 12490 2639 12498 2647
rect 16058 2639 16066 2647
rect 23104 2640 23112 2648
rect 25600 2640 25608 2648
rect 26928 2640 26936 2648
rect 28384 2640 28392 2648
rect 30512 2637 30520 2645
rect 30864 2637 30872 2645
rect 31360 2637 31368 2645
rect 31504 2637 31512 2645
rect 31824 2637 31832 2645
rect 32544 2637 32552 2645
rect 33840 2637 33848 2645
rect 33872 2637 33880 2645
rect 34608 2637 34616 2645
rect 36160 2637 36168 2645
rect 36496 2637 36504 2645
rect 37600 2637 37608 2645
rect 38352 2643 38360 2645
rect 38346 2637 38360 2643
rect 39440 2637 39448 2645
rect 38344 2629 38352 2637
rect 488 2619 496 2627
rect 808 2619 816 2627
rect 1208 2619 1216 2627
rect 1672 2619 1680 2627
rect 1800 2619 1808 2627
rect 2152 2619 2160 2627
rect 3336 2619 3344 2627
rect 3944 2619 3952 2627
rect 4120 2619 4128 2627
rect 4216 2619 4224 2627
rect 4296 2619 4304 2627
rect 4504 2619 4512 2627
rect 5858 2613 5866 2621
rect 6082 2613 6090 2621
rect 6194 2613 6202 2621
rect 6226 2613 6234 2621
rect 6274 2613 6282 2621
rect 6482 2613 6490 2621
rect 6674 2613 6682 2621
rect 8226 2613 8234 2621
rect 9330 2613 9338 2621
rect 9362 2613 9370 2621
rect 9458 2613 9466 2621
rect 10450 2613 10458 2621
rect 12298 2619 12306 2627
rect 13338 2619 13346 2627
rect 13578 2619 13586 2627
rect 13994 2619 14002 2627
rect 14474 2619 14482 2627
rect 15306 2619 15314 2627
rect 15322 2619 15330 2627
rect 15498 2619 15506 2627
rect 16058 2619 16066 2627
rect 16458 2619 16466 2627
rect 16586 2619 16594 2627
rect 16650 2619 16658 2627
rect 16842 2619 16850 2627
rect 18672 2620 18680 2628
rect 19904 2620 19912 2628
rect 21216 2620 21224 2628
rect 21280 2620 21288 2628
rect 22016 2620 22024 2628
rect 22416 2620 22424 2628
rect 23936 2620 23944 2628
rect 24944 2620 24952 2628
rect 26032 2620 26040 2628
rect 27360 2620 27368 2628
rect 28320 2620 28328 2628
rect 29376 2617 29384 2625
rect 29488 2617 29496 2625
rect 29712 2617 29720 2625
rect 29888 2617 29896 2625
rect 30256 2617 30264 2625
rect 30320 2617 30328 2625
rect 30464 2617 30472 2625
rect 30576 2617 30584 2625
rect 30816 2617 30824 2625
rect 31024 2617 31032 2625
rect 31072 2617 31080 2625
rect 32000 2617 32008 2625
rect 32304 2617 32312 2625
rect 33184 2617 33192 2625
rect 33232 2617 33240 2625
rect 33248 2617 33256 2625
rect 34464 2617 34472 2625
rect 36080 2617 36088 2625
rect 36496 2617 36504 2625
rect 36704 2617 36712 2625
rect 36784 2617 36792 2625
rect 36848 2617 36856 2625
rect 37136 2617 37144 2625
rect 37168 2617 37176 2625
rect 37360 2617 37368 2625
rect 37824 2617 37832 2625
rect 38640 2617 38648 2625
rect 38816 2617 38824 2625
rect 40288 2617 40296 2625
rect 40304 2617 40312 2625
rect 40368 2617 40376 2625
rect 584 2599 592 2607
rect 664 2599 672 2607
rect 696 2599 704 2607
rect 824 2599 832 2607
rect 856 2599 864 2607
rect 888 2599 896 2607
rect 920 2599 928 2607
rect 968 2599 976 2607
rect 1048 2599 1056 2607
rect 1080 2599 1088 2607
rect 1160 2599 1168 2607
rect 1192 2599 1200 2607
rect 1256 2599 1264 2607
rect 1656 2599 1664 2607
rect 1688 2599 1696 2607
rect 1704 2599 1712 2607
rect 1736 2599 1744 2607
rect 1832 2599 1840 2607
rect 1848 2599 1856 2607
rect 2104 2599 2112 2607
rect 2136 2599 2144 2607
rect 2280 2599 2288 2607
rect 2408 2599 2416 2607
rect 2856 2599 2864 2607
rect 2936 2599 2944 2607
rect 3016 2599 3024 2607
rect 3032 2599 3040 2607
rect 3176 2599 3184 2607
rect 3352 2599 3360 2607
rect 3464 2599 3472 2607
rect 3560 2599 3568 2607
rect 3832 2599 3840 2607
rect 3960 2599 3968 2607
rect 4200 2599 4208 2607
rect 4280 2599 4288 2607
rect 4376 2599 4384 2607
rect 4456 2599 4464 2607
rect 4472 2599 4480 2607
rect 6082 2593 6090 2601
rect 6210 2593 6218 2601
rect 6626 2593 6634 2601
rect 6706 2593 6714 2601
rect 7218 2593 7226 2601
rect 7426 2593 7434 2601
rect 7842 2593 7850 2601
rect 8034 2593 8042 2601
rect 8338 2593 8346 2601
rect 8594 2593 8602 2601
rect 8626 2593 8634 2601
rect 8642 2593 8650 2601
rect 8658 2593 8666 2601
rect 8738 2593 8746 2601
rect 9202 2593 9210 2601
rect 9506 2593 9514 2601
rect 9842 2593 9850 2601
rect 10066 2593 10074 2601
rect 10514 2593 10522 2601
rect 10802 2593 10810 2601
rect 12042 2599 12050 2607
rect 12362 2599 12370 2607
rect 12426 2599 12434 2607
rect 12474 2599 12482 2607
rect 12618 2599 12626 2607
rect 12650 2599 12658 2607
rect 12746 2599 12754 2607
rect 13034 2599 13042 2607
rect 14666 2599 14674 2607
rect 14938 2599 14946 2607
rect 15066 2599 15074 2607
rect 16026 2599 16034 2607
rect 20064 2600 20072 2608
rect 29888 2597 29896 2605
rect 30192 2597 30200 2605
rect 30272 2597 30280 2605
rect 30688 2597 30696 2605
rect 31024 2597 31032 2605
rect 31680 2597 31688 2605
rect 31776 2597 31784 2605
rect 32000 2597 32008 2605
rect 32928 2597 32936 2605
rect 34368 2597 34376 2605
rect 34992 2597 35000 2605
rect 35328 2597 35336 2605
rect 38384 2597 38392 2605
rect 38480 2597 38488 2605
rect 39120 2597 39128 2605
rect 40288 2597 40296 2605
rect 40528 2597 40536 2605
rect 760 2579 768 2587
rect 1144 2579 1152 2587
rect 1304 2579 1312 2587
rect 1432 2579 1440 2587
rect 1528 2579 1536 2587
rect 2328 2579 2336 2587
rect 3288 2579 3296 2587
rect 3448 2579 3456 2587
rect 3464 2579 3472 2587
rect 3880 2579 3888 2587
rect 4168 2579 4176 2587
rect 4184 2579 4192 2587
rect 5826 2573 5834 2581
rect 6546 2573 6554 2581
rect 6642 2573 6650 2581
rect 6882 2573 6890 2581
rect 6914 2573 6922 2581
rect 6994 2573 7002 2581
rect 7026 2573 7034 2581
rect 7058 2573 7066 2581
rect 7154 2573 7162 2581
rect 8082 2573 8090 2581
rect 8162 2573 8170 2581
rect 8354 2573 8362 2581
rect 8386 2573 8394 2581
rect 9922 2573 9930 2581
rect 12106 2579 12114 2587
rect 12154 2579 12162 2587
rect 12442 2579 12450 2587
rect 12650 2579 12658 2587
rect 12746 2579 12754 2587
rect 13226 2579 13234 2587
rect 13386 2579 13394 2587
rect 13434 2579 13442 2587
rect 13498 2579 13506 2587
rect 13610 2579 13618 2587
rect 13882 2579 13890 2587
rect 14346 2579 14354 2587
rect 14426 2579 14434 2587
rect 15482 2579 15490 2587
rect 15626 2579 15634 2587
rect 15770 2579 15778 2587
rect 15866 2579 15874 2587
rect 16266 2579 16274 2587
rect 16714 2579 16722 2587
rect 16730 2579 16738 2587
rect 17114 2579 17122 2587
rect 17178 2579 17186 2587
rect 17370 2579 17378 2587
rect 17434 2579 17442 2587
rect 17498 2579 17506 2587
rect 19152 2580 19160 2588
rect 20496 2580 20504 2588
rect 21632 2580 21640 2588
rect 21840 2580 21848 2588
rect 22000 2580 22008 2588
rect 23040 2580 23048 2588
rect 23472 2580 23480 2588
rect 23840 2580 23848 2588
rect 23888 2580 23896 2588
rect 24176 2580 24184 2588
rect 24304 2580 24312 2588
rect 24320 2580 24328 2588
rect 25168 2580 25176 2588
rect 25504 2580 25512 2588
rect 25664 2580 25672 2588
rect 25888 2580 25896 2588
rect 27600 2580 27608 2588
rect 28240 2580 28248 2588
rect 29904 2577 29912 2585
rect 30384 2577 30392 2585
rect 30528 2577 30536 2585
rect 30848 2577 30856 2585
rect 31152 2577 31160 2585
rect 31728 2577 31736 2585
rect 31952 2577 31960 2585
rect 34272 2577 34280 2585
rect 34624 2577 34632 2585
rect 36352 2577 36360 2585
rect 36480 2577 36488 2585
rect 39712 2577 39720 2585
rect 39872 2577 39880 2585
rect 2248 2559 2256 2567
rect 2376 2559 2384 2567
rect 2520 2559 2528 2567
rect 2760 2559 2768 2567
rect 2952 2559 2960 2567
rect 3176 2559 3184 2567
rect 5874 2553 5882 2561
rect 6466 2553 6474 2561
rect 6498 2553 6506 2561
rect 6546 2553 6554 2561
rect 6930 2553 6938 2561
rect 7026 2553 7034 2561
rect 9202 2553 9210 2561
rect 9250 2553 9258 2561
rect 9266 2553 9274 2561
rect 9346 2553 9354 2561
rect 9378 2553 9386 2561
rect 9666 2553 9674 2561
rect 9874 2553 9882 2561
rect 9954 2553 9962 2561
rect 10242 2553 10250 2561
rect 10306 2553 10314 2561
rect 10754 2553 10762 2561
rect 12314 2559 12322 2567
rect 12890 2559 12898 2567
rect 14554 2559 14562 2567
rect 16058 2559 16066 2567
rect 16154 2559 16162 2567
rect 16714 2559 16722 2567
rect 16986 2559 16994 2567
rect 19040 2560 19048 2568
rect 24624 2560 24632 2568
rect 26832 2560 26840 2568
rect 30240 2557 30248 2565
rect 32592 2557 32600 2565
rect 32816 2557 32824 2565
rect 33056 2557 33064 2565
rect 33360 2557 33368 2565
rect 34400 2557 34408 2565
rect 35008 2557 35016 2565
rect 35440 2557 35448 2565
rect 35728 2557 35736 2565
rect 35808 2557 35816 2565
rect 36880 2557 36888 2565
rect 36976 2557 36984 2565
rect 37056 2557 37064 2565
rect 37312 2557 37320 2565
rect 37648 2557 37656 2565
rect 37760 2557 37768 2565
rect 38016 2557 38024 2565
rect 38032 2557 38040 2565
rect 38576 2557 38584 2565
rect 38896 2557 38904 2565
rect 39008 2557 39016 2565
rect 19056 2548 19060 2553
rect 20094 2548 20098 2553
rect 20720 2548 20724 2553
rect 21830 2548 21834 2553
rect 26292 2548 26296 2553
rect 456 2539 464 2547
rect 808 2539 816 2547
rect 904 2539 912 2547
rect 952 2539 960 2547
rect 1544 2539 1552 2547
rect 1816 2539 1824 2547
rect 1928 2539 1936 2547
rect 1992 2539 2000 2547
rect 2088 2539 2096 2547
rect 2648 2539 2656 2547
rect 2728 2539 2736 2547
rect 2776 2539 2784 2547
rect 3112 2539 3120 2547
rect 3128 2539 3136 2547
rect 3496 2539 3504 2547
rect 3608 2539 3616 2547
rect 3912 2539 3920 2547
rect 4024 2539 4032 2547
rect 4200 2539 4208 2547
rect 4232 2539 4240 2547
rect 4552 2539 4560 2547
rect 4632 2539 4640 2547
rect 6162 2533 6170 2541
rect 6226 2533 6234 2541
rect 6738 2533 6746 2541
rect 6754 2533 6762 2541
rect 6786 2533 6794 2541
rect 7106 2533 7114 2541
rect 7346 2533 7354 2541
rect 7426 2533 7434 2541
rect 7618 2533 7626 2541
rect 7634 2533 7642 2541
rect 7698 2533 7706 2541
rect 7714 2533 7722 2541
rect 7842 2533 7850 2541
rect 7906 2533 7914 2541
rect 8386 2533 8394 2541
rect 8466 2533 8474 2541
rect 8898 2533 8906 2541
rect 8914 2533 8922 2541
rect 9122 2533 9130 2541
rect 9186 2533 9194 2541
rect 9730 2533 9738 2541
rect 9858 2533 9866 2541
rect 9954 2533 9962 2541
rect 10194 2533 10202 2541
rect 10226 2533 10234 2541
rect 10418 2533 10426 2541
rect 10466 2533 10474 2541
rect 10514 2533 10522 2541
rect 10594 2533 10602 2541
rect 12570 2539 12578 2547
rect 12922 2539 12930 2547
rect 13370 2539 13378 2547
rect 13482 2539 13490 2547
rect 13658 2539 13666 2547
rect 14506 2539 14514 2547
rect 14762 2539 14770 2547
rect 14938 2539 14946 2547
rect 15114 2539 15122 2547
rect 15322 2539 15330 2547
rect 15418 2539 15426 2547
rect 15530 2539 15538 2547
rect 15610 2539 15618 2547
rect 15642 2539 15650 2547
rect 16074 2539 16082 2547
rect 16122 2539 16130 2547
rect 16266 2539 16274 2547
rect 16538 2539 16546 2547
rect 16570 2539 16578 2547
rect 16650 2539 16658 2547
rect 16698 2539 16706 2547
rect 16746 2539 16754 2547
rect 16762 2539 16770 2547
rect 16810 2539 16818 2547
rect 17130 2539 17138 2547
rect 17354 2539 17362 2547
rect 18496 2540 18504 2548
rect 20304 2540 20312 2548
rect 21120 2540 21128 2548
rect 21408 2540 21416 2548
rect 22256 2540 22264 2548
rect 22624 2540 22632 2548
rect 22656 2540 22664 2548
rect 23056 2540 23064 2548
rect 23344 2540 23352 2548
rect 23472 2540 23480 2548
rect 23696 2540 23704 2548
rect 23760 2540 23768 2548
rect 24800 2540 24808 2548
rect 26256 2540 26264 2548
rect 26512 2540 26520 2548
rect 27056 2540 27064 2548
rect 27520 2540 27528 2548
rect 27792 2540 27800 2548
rect 28208 2540 28216 2548
rect 28576 2540 28584 2548
rect 29664 2537 29672 2545
rect 33232 2537 33240 2545
rect 2216 2519 2224 2527
rect 6546 2513 6554 2521
rect 6578 2513 6586 2521
rect 6594 2513 6602 2521
rect 7410 2513 7418 2521
rect 8258 2513 8266 2521
rect 8578 2513 8586 2521
rect 8594 2513 8602 2521
rect 8770 2513 8778 2521
rect 8818 2513 8826 2521
rect 9490 2513 9498 2521
rect 9586 2513 9594 2521
rect 9602 2513 9610 2521
rect 9858 2513 9866 2521
rect 10114 2513 10122 2521
rect 10274 2513 10282 2521
rect 10530 2513 10538 2521
rect 13130 2519 13138 2527
rect 15386 2519 15394 2527
rect 15706 2519 15714 2527
rect 16394 2519 16402 2527
rect 17242 2519 17250 2527
rect 19552 2520 19560 2528
rect 20704 2520 20712 2528
rect 24976 2520 24984 2528
rect 25440 2520 25448 2528
rect 38960 2517 38968 2525
rect 2024 2499 2032 2507
rect 2232 2499 2240 2507
rect 3720 2499 3728 2507
rect 3736 2499 3744 2507
rect 8146 2493 8154 2501
rect 15050 2499 15058 2507
rect 15274 2499 15282 2507
rect 15674 2499 15682 2507
rect 32288 2497 32296 2505
rect 568 2479 576 2487
rect 680 2479 688 2487
rect 840 2479 848 2487
rect 872 2479 880 2487
rect 1032 2479 1040 2487
rect 1064 2479 1072 2487
rect 1080 2479 1088 2487
rect 1176 2479 1184 2487
rect 2264 2479 2272 2487
rect 2392 2479 2400 2487
rect 4264 2479 4272 2487
rect 4360 2479 4368 2487
rect 6066 2473 6074 2481
rect 6610 2473 6618 2481
rect 6690 2473 6698 2481
rect 7234 2473 7242 2481
rect 8146 2473 8154 2481
rect 8322 2473 8330 2481
rect 9058 2473 9066 2481
rect 10546 2473 10554 2481
rect 13850 2479 13858 2487
rect 24736 2480 24744 2488
rect 37920 2477 37928 2485
rect 572 2463 596 2467
rect 4452 2463 4476 2467
rect 6690 2453 6698 2461
rect 8322 2453 8330 2461
rect 9730 2453 9738 2461
rect 10050 2453 10058 2461
rect 28416 2460 28424 2468
rect 29396 2467 29408 2475
rect 29428 2467 29440 2475
rect 29444 2467 29448 2475
rect 29460 2467 29472 2475
rect 29492 2467 29504 2475
rect 29516 2467 29520 2475
rect 29524 2467 29536 2475
rect 29672 2467 29676 2475
rect 29680 2467 29692 2475
rect 29696 2467 29700 2475
rect 29712 2467 29724 2475
rect 29736 2467 29740 2475
rect 29744 2467 29756 2475
rect 29964 2467 29976 2475
rect 29988 2467 29992 2475
rect 29996 2467 30008 2475
rect 30012 2467 30016 2475
rect 30056 2467 30068 2475
rect 30080 2467 30084 2475
rect 30088 2467 30100 2475
rect 30104 2467 30108 2475
rect 30120 2467 30132 2475
rect 30172 2467 30176 2475
rect 30180 2467 30192 2475
rect 30196 2467 30200 2475
rect 30212 2467 30224 2475
rect 30244 2467 30256 2475
rect 30260 2467 30264 2475
rect 30276 2467 30288 2475
rect 30304 2467 30320 2475
rect 30328 2467 30360 2475
rect 30368 2467 30384 2475
rect 30400 2467 30416 2475
rect 30432 2467 30436 2475
rect 30440 2467 30452 2475
rect 30456 2467 30468 2475
rect 30472 2467 30476 2475
rect 30496 2467 30500 2475
rect 30504 2467 30508 2475
rect 30528 2467 30532 2475
rect 30536 2467 30540 2475
rect 30560 2467 30564 2475
rect 30568 2467 30572 2475
rect 30592 2467 30596 2475
rect 30600 2467 30612 2475
rect 30616 2467 30628 2475
rect 30632 2467 30636 2475
rect 30652 2467 30668 2475
rect 30684 2467 30688 2475
rect 30692 2467 30704 2475
rect 30708 2467 30720 2475
rect 30724 2467 30728 2475
rect 30748 2467 30752 2475
rect 30756 2467 30760 2475
rect 30772 2467 30784 2475
rect 30788 2467 30792 2475
rect 30812 2467 30816 2475
rect 30820 2467 30824 2475
rect 30844 2467 30848 2475
rect 30852 2467 30864 2475
rect 30876 2467 30880 2475
rect 30884 2467 30888 2475
rect 30908 2467 30912 2475
rect 30916 2467 30920 2475
rect 30932 2467 30944 2475
rect 30948 2467 30952 2475
rect 30972 2467 30976 2475
rect 30980 2467 30984 2475
rect 31004 2467 31008 2475
rect 31012 2467 31024 2475
rect 31036 2467 31040 2475
rect 31044 2467 31048 2475
rect 31224 2467 31228 2475
rect 31232 2467 31236 2475
rect 31300 2467 31304 2475
rect 31308 2467 31312 2475
rect 31332 2467 31336 2475
rect 31340 2467 31344 2475
rect 31356 2467 31368 2475
rect 31372 2467 31376 2475
rect 31392 2467 31416 2475
rect 31424 2467 31440 2475
rect 31448 2467 31460 2475
rect 31464 2467 31468 2475
rect 31488 2467 31492 2475
rect 31496 2467 31508 2475
rect 31520 2467 31524 2475
rect 31528 2467 31532 2475
rect 31708 2467 31712 2475
rect 31716 2467 31720 2475
rect 31740 2467 31744 2475
rect 31748 2467 31752 2475
rect 31764 2467 31776 2475
rect 31780 2467 31784 2475
rect 31800 2467 31824 2475
rect 31832 2467 31848 2475
rect 31856 2467 31880 2475
rect 31896 2467 31900 2475
rect 31904 2467 31916 2475
rect 31924 2467 31940 2475
rect 31948 2467 31972 2475
rect 31988 2467 32000 2475
rect 32012 2467 32036 2475
rect 32052 2467 32064 2475
rect 32068 2467 32072 2475
rect 32084 2467 32096 2475
rect 32108 2467 32112 2475
rect 32116 2467 32128 2475
rect 32148 2467 32160 2475
rect 32180 2467 32192 2475
rect 32212 2467 32224 2475
rect 32228 2467 32232 2475
rect 32244 2467 32256 2475
rect 32268 2467 32272 2475
rect 32276 2467 32288 2475
rect 32292 2467 32296 2475
rect 32492 2467 32504 2475
rect 32516 2467 32520 2475
rect 32524 2467 32536 2475
rect 32540 2467 32544 2475
rect 32584 2467 32596 2475
rect 32608 2467 32612 2475
rect 32616 2467 32628 2475
rect 32632 2467 32636 2475
rect 32648 2467 32660 2475
rect 32764 2467 32768 2475
rect 32772 2467 32784 2475
rect 32788 2467 32792 2475
rect 32896 2467 32908 2475
rect 32920 2467 32924 2475
rect 32928 2467 32940 2475
rect 32944 2467 32948 2475
rect 32960 2467 32972 2475
rect 33012 2467 33016 2475
rect 33020 2467 33032 2475
rect 33036 2467 33040 2475
rect 33080 2467 33092 2475
rect 33104 2467 33108 2475
rect 33112 2467 33124 2475
rect 33128 2467 33132 2475
rect 33144 2467 33156 2475
rect 33324 2467 33328 2475
rect 33332 2467 33344 2475
rect 33364 2467 33376 2475
rect 33380 2467 33384 2475
rect 33416 2467 33420 2475
rect 33424 2467 33436 2475
rect 33456 2467 33468 2475
rect 33472 2467 33476 2475
rect 33548 2467 33560 2475
rect 33580 2467 33592 2475
rect 33596 2467 33600 2475
rect 33612 2467 33624 2475
rect 33636 2467 33640 2475
rect 33644 2467 33656 2475
rect 33672 2467 33720 2475
rect 33736 2467 33748 2475
rect 33768 2467 33780 2475
rect 33792 2467 33796 2475
rect 33800 2467 33812 2475
rect 33924 2467 33936 2475
rect 33956 2467 33968 2475
rect 33972 2467 33976 2475
rect 33988 2467 34000 2475
rect 34012 2467 34016 2475
rect 34020 2467 34032 2475
rect 34048 2467 34060 2475
rect 34064 2467 34068 2475
rect 34080 2467 34092 2475
rect 34100 2467 34124 2475
rect 34140 2467 34188 2475
rect 34204 2467 34208 2475
rect 34212 2467 34216 2475
rect 34228 2467 34240 2475
rect 34244 2467 34256 2475
rect 34268 2467 34272 2475
rect 34276 2467 34280 2475
rect 34292 2467 34304 2475
rect 34308 2467 34320 2475
rect 34332 2467 34336 2475
rect 34340 2467 34344 2475
rect 34424 2467 34428 2475
rect 34432 2467 34436 2475
rect 34516 2467 34520 2475
rect 34524 2467 34528 2475
rect 34540 2467 34552 2475
rect 34556 2467 34568 2475
rect 34580 2467 34584 2475
rect 34588 2467 34592 2475
rect 34612 2467 34616 2475
rect 34620 2467 34624 2475
rect 34688 2467 34692 2475
rect 34696 2467 34708 2475
rect 34720 2467 34724 2475
rect 34728 2467 34732 2475
rect 34780 2467 34784 2475
rect 34788 2467 34800 2475
rect 34812 2467 34816 2475
rect 34820 2467 34824 2475
rect 34952 2467 34956 2475
rect 34960 2467 34964 2475
rect 34976 2467 34988 2475
rect 34992 2467 34996 2475
rect 35016 2467 35020 2475
rect 35024 2467 35028 2475
rect 35044 2467 35092 2475
rect 35108 2467 35112 2475
rect 35116 2467 35120 2475
rect 35136 2467 35184 2475
rect 35200 2467 35224 2475
rect 35232 2467 35244 2475
rect 35256 2467 35260 2475
rect 35264 2467 35276 2475
rect 35296 2467 35308 2475
rect 35320 2467 35324 2475
rect 35328 2467 35340 2475
rect 35360 2467 35372 2475
rect 35376 2467 35380 2475
rect 35452 2467 35464 2475
rect 35468 2467 35472 2475
rect 35576 2467 35588 2475
rect 35592 2467 35604 2475
rect 35608 2467 35620 2475
rect 35636 2467 35652 2475
rect 35668 2467 35692 2475
rect 35700 2467 35716 2475
rect 35732 2467 35748 2475
rect 35756 2467 35768 2475
rect 35772 2467 35784 2475
rect 35796 2467 35800 2475
rect 35804 2467 35808 2475
rect 35820 2467 35832 2475
rect 35836 2467 35840 2475
rect 35936 2467 35940 2475
rect 35944 2467 35948 2475
rect 35960 2467 35972 2475
rect 35976 2467 35988 2475
rect 36000 2467 36004 2475
rect 36008 2467 36012 2475
rect 36028 2467 36076 2475
rect 36088 2467 36104 2475
rect 36120 2467 36168 2475
rect 36184 2467 36200 2475
rect 36216 2467 36228 2475
rect 36240 2467 36244 2475
rect 36248 2467 36260 2475
rect 36280 2467 36292 2475
rect 36296 2467 36300 2475
rect 36532 2467 36544 2475
rect 36548 2467 36560 2475
rect 36564 2467 36576 2475
rect 36596 2467 36608 2475
rect 36620 2467 36624 2475
rect 36628 2467 36640 2475
rect 36660 2467 36672 2475
rect 36692 2467 36704 2475
rect 36708 2467 36712 2475
rect 36724 2467 36736 2475
rect 36756 2467 36768 2475
rect 36776 2467 36800 2475
rect 36816 2467 36832 2475
rect 36840 2467 36872 2475
rect 36880 2467 36896 2475
rect 36912 2467 36924 2475
rect 36928 2467 36940 2475
rect 36944 2467 36956 2475
rect 36976 2467 36988 2475
rect 37092 2467 37096 2475
rect 37100 2467 37112 2475
rect 37116 2467 37120 2475
rect 37132 2467 37144 2475
rect 37152 2467 37176 2475
rect 37192 2467 37240 2475
rect 37256 2467 37268 2475
rect 37284 2467 37332 2475
rect 37348 2467 37360 2475
rect 37376 2467 37424 2475
rect 37440 2467 37452 2475
rect 37472 2467 37484 2475
rect 37496 2467 37500 2475
rect 37504 2467 37516 2475
rect 37536 2467 37548 2475
rect 37552 2467 37556 2475
rect 37568 2467 37580 2475
rect 37600 2467 37612 2475
rect 37616 2467 37620 2475
rect 37632 2467 37644 2475
rect 37656 2467 37660 2475
rect 37664 2467 37676 2475
rect 37692 2467 37716 2475
rect 37724 2467 37736 2475
rect 37744 2467 37768 2475
rect 37784 2467 37808 2475
rect 37816 2467 37832 2475
rect 37848 2467 37852 2475
rect 37856 2467 37860 2475
rect 37880 2467 37884 2475
rect 37888 2467 37900 2475
rect 37904 2467 37916 2475
rect 37920 2467 37924 2475
rect 38052 2467 38056 2475
rect 38060 2467 38064 2475
rect 38160 2467 38164 2475
rect 38168 2467 38172 2475
rect 38192 2467 38196 2475
rect 38200 2467 38212 2475
rect 38216 2467 38228 2475
rect 38232 2467 38236 2475
rect 38256 2467 38260 2475
rect 38264 2467 38276 2475
rect 38288 2467 38292 2475
rect 38296 2467 38300 2475
rect 38320 2467 38324 2475
rect 38328 2467 38332 2475
rect 38352 2467 38356 2475
rect 38360 2467 38364 2475
rect 38376 2467 38388 2475
rect 38392 2467 38396 2475
rect 38412 2467 38436 2475
rect 38444 2467 38460 2475
rect 38468 2467 38480 2475
rect 38484 2467 38488 2475
rect 38504 2467 38528 2475
rect 38536 2467 38552 2475
rect 38560 2467 38572 2475
rect 38576 2467 38580 2475
rect 38596 2467 38620 2475
rect 38628 2467 38644 2475
rect 38652 2467 38664 2475
rect 38668 2467 38672 2475
rect 38692 2467 38696 2475
rect 38700 2467 38712 2475
rect 38720 2467 38736 2475
rect 38744 2467 38768 2475
rect 38784 2467 38796 2475
rect 38816 2467 38828 2475
rect 38840 2467 38844 2475
rect 38848 2467 38860 2475
rect 38864 2467 38868 2475
rect 38932 2467 38936 2475
rect 38940 2467 38952 2475
rect 38956 2467 38960 2475
rect 38972 2467 38984 2475
rect 38992 2467 39016 2475
rect 39032 2467 39056 2475
rect 39064 2467 39080 2475
rect 39096 2467 39100 2475
rect 39104 2467 39108 2475
rect 39128 2467 39132 2475
rect 39136 2467 39148 2475
rect 39152 2467 39164 2475
rect 39168 2467 39172 2475
rect 39188 2467 39200 2475
rect 39220 2467 39224 2475
rect 39228 2467 39240 2475
rect 39244 2467 39256 2475
rect 39260 2467 39264 2475
rect 39284 2467 39288 2475
rect 39292 2467 39304 2475
rect 39312 2467 39328 2475
rect 39336 2467 39360 2475
rect 39376 2467 39392 2475
rect 39400 2467 39424 2475
rect 39440 2467 39488 2475
rect 39504 2467 39508 2475
rect 39512 2467 39516 2475
rect 39532 2467 39580 2475
rect 39596 2467 39612 2475
rect 39628 2467 39632 2475
rect 39636 2467 39648 2475
rect 39660 2467 39664 2475
rect 39668 2467 39672 2475
rect 39692 2467 39696 2475
rect 39700 2467 39704 2475
rect 39716 2467 39728 2475
rect 39732 2467 39736 2475
rect 39752 2467 39768 2475
rect 39784 2467 39832 2475
rect 39848 2467 39864 2475
rect 39880 2467 39892 2475
rect 39904 2467 39908 2475
rect 39912 2467 39924 2475
rect 40036 2467 40048 2475
rect 40052 2467 40064 2475
rect 40068 2467 40080 2475
rect 40100 2467 40112 2475
rect 40256 2467 40268 2475
rect 40288 2467 40300 2475
rect 40304 2467 40316 2475
rect 40320 2467 40332 2475
rect 40404 2467 40408 2475
rect 40412 2467 40424 2475
rect 40444 2467 40456 2475
rect 40460 2467 40472 2475
rect 40476 2467 40488 2475
rect 40504 2467 40516 2475
rect 40536 2467 40548 2475
rect 40552 2467 40564 2475
rect 40568 2467 40580 2475
rect 40596 2467 40608 2475
rect 40628 2467 40640 2475
rect 40644 2467 40656 2475
rect 40660 2467 40672 2475
rect 40688 2467 40704 2475
rect 40720 2467 40732 2475
rect 40736 2467 40748 2475
rect 40752 2467 40764 2475
rect 40780 2467 40792 2475
rect 18776 2450 18786 2458
rect 18990 2450 19000 2458
rect 21280 2450 21290 2458
rect 23206 2450 23216 2458
rect 27644 2450 27646 2458
rect 27652 2450 27654 2458
rect 27858 2450 27860 2458
rect 27866 2450 27868 2458
rect 1176 2439 1184 2447
rect 5810 2433 5818 2441
rect 6306 2433 6314 2441
rect 8146 2433 8154 2441
rect 12234 2439 12242 2447
rect 16410 2439 16418 2447
rect 17098 2439 17106 2447
rect 26288 2440 26296 2448
rect 28560 2440 28568 2448
rect 35152 2437 35160 2445
rect 40032 2437 40040 2445
rect 1352 2419 1360 2427
rect 1560 2419 1568 2427
rect 2424 2419 2432 2427
rect 2648 2419 2656 2427
rect 3176 2419 3184 2427
rect 3320 2419 3328 2427
rect 3816 2419 3824 2427
rect 4024 2419 4032 2427
rect 4056 2419 4064 2427
rect 4392 2419 4400 2427
rect 4408 2419 4416 2427
rect 4456 2419 4464 2427
rect 6082 2413 6090 2421
rect 7378 2413 7386 2421
rect 7666 2413 7674 2421
rect 8050 2413 8058 2421
rect 8258 2413 8266 2421
rect 8466 2413 8474 2421
rect 9730 2413 9738 2421
rect 9778 2413 9786 2421
rect 12698 2419 12706 2427
rect 15626 2419 15634 2427
rect 19120 2420 19128 2428
rect 20784 2420 20792 2428
rect 38800 2417 38808 2425
rect 39376 2417 39384 2425
rect 680 2399 688 2407
rect 1032 2399 1040 2407
rect 1432 2399 1440 2407
rect 1848 2399 1856 2407
rect 2024 2399 2032 2407
rect 2296 2399 2304 2407
rect 2680 2399 2688 2407
rect 3304 2399 3312 2407
rect 3512 2399 3520 2407
rect 4088 2399 4096 2407
rect 8034 2393 8042 2401
rect 9650 2393 9658 2401
rect 10418 2393 10426 2401
rect 12890 2399 12898 2407
rect 13770 2399 13778 2407
rect 15882 2399 15890 2407
rect 16314 2399 16322 2407
rect 16330 2399 16338 2407
rect 17242 2399 17250 2407
rect 26512 2400 26520 2408
rect 27760 2400 27768 2408
rect 29408 2397 29416 2405
rect 34816 2397 34824 2405
rect 632 2379 640 2387
rect 1688 2379 1696 2387
rect 1736 2379 1744 2387
rect 2504 2379 2512 2387
rect 3272 2379 3280 2387
rect 3352 2379 3360 2387
rect 6290 2373 6298 2381
rect 6322 2373 6330 2381
rect 6338 2373 6346 2381
rect 6482 2373 6490 2381
rect 7218 2373 7226 2381
rect 7250 2373 7258 2381
rect 7266 2373 7274 2381
rect 8130 2373 8138 2381
rect 8402 2373 8410 2381
rect 8818 2373 8826 2381
rect 9218 2373 9226 2381
rect 9298 2373 9306 2381
rect 9714 2373 9722 2381
rect 10034 2373 10042 2381
rect 10146 2373 10154 2381
rect 10450 2373 10458 2381
rect 13930 2379 13938 2387
rect 13962 2379 13970 2387
rect 14858 2379 14866 2387
rect 14874 2379 14882 2387
rect 16314 2379 16322 2387
rect 16842 2379 16850 2387
rect 16858 2379 16866 2387
rect 24560 2380 24568 2388
rect 25424 2380 25432 2388
rect 30768 2377 30776 2385
rect 31200 2377 31208 2385
rect 32400 2377 32408 2385
rect 32448 2377 32456 2385
rect 33376 2377 33384 2385
rect 34464 2377 34472 2385
rect 34704 2377 34712 2385
rect 36096 2377 36104 2385
rect 36944 2377 36952 2385
rect 37456 2377 37464 2385
rect 40096 2377 40104 2385
rect 40368 2377 40376 2385
rect 488 2359 496 2367
rect 568 2359 576 2367
rect 776 2359 784 2367
rect 1000 2359 1008 2367
rect 1416 2359 1424 2367
rect 1496 2359 1504 2367
rect 1608 2359 1616 2367
rect 1960 2359 1968 2367
rect 3000 2359 3008 2367
rect 4280 2359 4288 2367
rect 4360 2359 4368 2367
rect 4520 2359 4528 2367
rect 6754 2353 6762 2361
rect 6946 2353 6954 2361
rect 7298 2353 7306 2361
rect 7346 2353 7354 2361
rect 7554 2353 7562 2361
rect 7634 2353 7642 2361
rect 7778 2353 7786 2361
rect 8690 2353 8698 2361
rect 8738 2353 8746 2361
rect 9346 2353 9354 2361
rect 9378 2353 9386 2361
rect 9634 2353 9642 2361
rect 9842 2353 9850 2361
rect 10514 2353 10522 2361
rect 10898 2353 10906 2361
rect 12570 2359 12578 2367
rect 12874 2359 12882 2367
rect 14762 2359 14770 2367
rect 14954 2359 14962 2367
rect 15002 2359 15010 2367
rect 15162 2359 15170 2367
rect 16394 2359 16402 2367
rect 16554 2359 16562 2367
rect 16586 2359 16594 2367
rect 16618 2359 16626 2367
rect 16938 2359 16946 2367
rect 16986 2359 16994 2367
rect 17306 2359 17314 2367
rect 17450 2359 17458 2367
rect 18720 2360 18728 2368
rect 18928 2360 18936 2368
rect 19296 2360 19304 2368
rect 20352 2360 20360 2368
rect 21216 2360 21224 2368
rect 21872 2360 21880 2368
rect 22448 2361 22458 2366
rect 22864 2360 22872 2368
rect 23264 2360 23272 2368
rect 23505 2361 23510 2366
rect 23984 2360 23992 2368
rect 24608 2360 24616 2368
rect 24960 2360 24968 2368
rect 26240 2360 26248 2368
rect 27932 2361 27942 2366
rect 27966 2361 27976 2366
rect 35312 2357 35320 2365
rect 35344 2357 35352 2365
rect 36064 2357 36072 2365
rect 36384 2357 36392 2365
rect 36608 2357 36616 2365
rect 632 2339 640 2347
rect 792 2339 800 2347
rect 6146 2333 6154 2341
rect 6226 2333 6234 2341
rect 6290 2333 6298 2341
rect 6498 2333 6506 2341
rect 6626 2333 6634 2341
rect 6770 2333 6778 2341
rect 6930 2333 6938 2341
rect 7122 2333 7130 2341
rect 7250 2333 7258 2341
rect 7314 2333 7322 2341
rect 7474 2333 7482 2341
rect 7794 2333 7802 2341
rect 7954 2333 7962 2341
rect 8194 2333 8202 2341
rect 8498 2333 8506 2341
rect 8738 2333 8746 2341
rect 8866 2333 8874 2341
rect 8946 2333 8954 2341
rect 9266 2333 9274 2341
rect 10562 2333 10570 2341
rect 10770 2333 10778 2341
rect 12554 2339 12562 2347
rect 13018 2339 13026 2347
rect 13786 2339 13794 2347
rect 14938 2339 14946 2347
rect 15066 2339 15074 2347
rect 15434 2339 15442 2347
rect 15482 2339 15490 2347
rect 15498 2339 15506 2347
rect 15706 2339 15714 2347
rect 15898 2339 15906 2347
rect 15962 2339 15970 2347
rect 19536 2340 19544 2348
rect 19664 2340 19672 2348
rect 20592 2340 20600 2348
rect 25472 2340 25480 2348
rect 26928 2340 26936 2348
rect 27968 2340 27976 2348
rect 31344 2337 31352 2345
rect 36352 2337 36360 2345
rect 36640 2337 36648 2345
rect 37024 2337 37032 2345
rect 37584 2337 37592 2345
rect 37808 2337 37816 2345
rect 38048 2337 38056 2345
rect 38144 2337 38152 2345
rect 38240 2337 38248 2345
rect 38256 2337 38264 2345
rect 38304 2337 38312 2345
rect 39968 2337 39976 2345
rect 40384 2337 40392 2345
rect 40672 2337 40680 2345
rect 744 2319 752 2327
rect 872 2319 880 2327
rect 1000 2319 1008 2327
rect 2504 2319 2512 2327
rect 2536 2319 2544 2327
rect 2552 2319 2560 2327
rect 2728 2319 2736 2327
rect 2760 2319 2768 2327
rect 2824 2319 2832 2327
rect 6514 2313 6522 2321
rect 6642 2313 6650 2321
rect 6706 2313 6714 2321
rect 6962 2313 6970 2321
rect 7026 2313 7034 2321
rect 7714 2313 7722 2321
rect 8114 2313 8122 2321
rect 8130 2313 8138 2321
rect 8242 2313 8250 2321
rect 8322 2313 8330 2321
rect 8482 2313 8490 2321
rect 8706 2313 8714 2321
rect 9458 2313 9466 2321
rect 9490 2313 9498 2321
rect 9554 2313 9562 2321
rect 9650 2313 9658 2321
rect 9874 2313 9882 2321
rect 9938 2313 9946 2321
rect 9986 2313 9994 2321
rect 10130 2313 10138 2321
rect 10146 2313 10154 2321
rect 10306 2313 10314 2321
rect 10450 2313 10458 2321
rect 10546 2313 10554 2321
rect 10610 2313 10618 2321
rect 10802 2313 10810 2321
rect 12122 2319 12130 2327
rect 12186 2319 12194 2327
rect 12922 2319 12930 2327
rect 13402 2319 13410 2327
rect 13418 2319 13426 2327
rect 13642 2319 13650 2327
rect 13850 2319 13858 2327
rect 14682 2319 14690 2327
rect 14906 2319 14914 2327
rect 15034 2319 15042 2327
rect 15258 2319 15266 2327
rect 15578 2319 15586 2327
rect 15770 2319 15778 2327
rect 16154 2319 16162 2327
rect 16538 2319 16546 2327
rect 17066 2319 17074 2327
rect 18528 2320 18536 2328
rect 18704 2320 18712 2328
rect 18736 2320 18744 2328
rect 18944 2320 18952 2328
rect 19280 2320 19288 2328
rect 19328 2320 19336 2328
rect 19360 2320 19368 2328
rect 19696 2320 19704 2328
rect 20624 2320 20632 2328
rect 20944 2320 20952 2328
rect 21456 2320 21464 2328
rect 22832 2320 22840 2328
rect 23072 2320 23080 2328
rect 23488 2320 23496 2328
rect 24000 2320 24008 2328
rect 26528 2320 26536 2328
rect 27264 2320 27272 2328
rect 27984 2320 27992 2328
rect 29792 2317 29800 2325
rect 29872 2317 29880 2325
rect 30176 2317 30184 2325
rect 30928 2317 30936 2325
rect 31120 2317 31128 2325
rect 31376 2317 31384 2325
rect 31440 2317 31448 2325
rect 31888 2317 31896 2325
rect 32000 2317 32008 2325
rect 35040 2317 35048 2325
rect 35616 2317 35624 2325
rect 35696 2317 35704 2325
rect 35776 2317 35784 2325
rect 36592 2317 36600 2325
rect 36640 2317 36648 2325
rect 36672 2317 36680 2325
rect 36816 2317 36824 2325
rect 37136 2317 37144 2325
rect 37184 2317 37192 2325
rect 37216 2317 37224 2325
rect 37952 2317 37960 2325
rect 37968 2317 37976 2325
rect 39312 2317 39320 2325
rect 39904 2317 39912 2325
rect 424 2299 432 2307
rect 504 2299 512 2307
rect 600 2299 608 2307
rect 616 2299 624 2307
rect 840 2299 848 2307
rect 904 2299 912 2307
rect 968 2299 976 2307
rect 1048 2299 1056 2307
rect 1144 2299 1152 2307
rect 1336 2299 1344 2307
rect 1432 2299 1440 2307
rect 1528 2299 1536 2307
rect 1544 2299 1552 2307
rect 1672 2299 1680 2307
rect 1864 2299 1872 2307
rect 1880 2299 1888 2307
rect 1896 2299 1904 2307
rect 2008 2299 2016 2307
rect 2088 2299 2096 2307
rect 2136 2299 2144 2307
rect 2248 2299 2256 2307
rect 2280 2299 2288 2307
rect 2312 2299 2320 2307
rect 2328 2299 2336 2307
rect 2408 2299 2416 2307
rect 3160 2299 3168 2307
rect 3480 2299 3488 2307
rect 3688 2299 3696 2307
rect 3912 2299 3920 2307
rect 4040 2299 4048 2307
rect 4360 2299 4368 2307
rect 4376 2299 4384 2307
rect 4424 2299 4432 2307
rect 4440 2299 4448 2307
rect 4568 2299 4576 2307
rect 4600 2299 4608 2307
rect 4664 2299 4672 2307
rect 5746 2293 5754 2301
rect 5778 2293 5786 2301
rect 5890 2293 5898 2301
rect 5906 2293 5914 2301
rect 5938 2293 5946 2301
rect 6018 2293 6026 2301
rect 6050 2293 6058 2301
rect 6066 2293 6074 2301
rect 6242 2293 6250 2301
rect 6258 2293 6266 2301
rect 6354 2293 6362 2301
rect 6386 2293 6394 2301
rect 6562 2293 6570 2301
rect 6610 2293 6618 2301
rect 7186 2293 7194 2301
rect 7250 2293 7258 2301
rect 7394 2293 7402 2301
rect 7522 2293 7530 2301
rect 7570 2293 7578 2301
rect 7650 2293 7658 2301
rect 7746 2293 7754 2301
rect 8066 2293 8074 2301
rect 8226 2293 8234 2301
rect 8274 2293 8282 2301
rect 8306 2293 8314 2301
rect 8450 2293 8458 2301
rect 8834 2293 8842 2301
rect 9186 2293 9194 2301
rect 9586 2293 9594 2301
rect 9666 2293 9674 2301
rect 9698 2293 9706 2301
rect 9746 2293 9754 2301
rect 9986 2293 9994 2301
rect 10114 2293 10122 2301
rect 10130 2293 10138 2301
rect 10162 2293 10170 2301
rect 10242 2293 10250 2301
rect 10498 2293 10506 2301
rect 10578 2293 10586 2301
rect 10642 2293 10650 2301
rect 12058 2299 12066 2307
rect 14922 2299 14930 2307
rect 15050 2299 15058 2307
rect 15562 2299 15570 2307
rect 17050 2299 17058 2307
rect 19760 2300 19768 2308
rect 21616 2300 21624 2308
rect 22048 2300 22056 2308
rect 22208 2300 22216 2308
rect 27280 2300 27288 2308
rect 27888 2300 27896 2308
rect 28208 2300 28216 2308
rect 31920 2297 31928 2305
rect 32032 2297 32040 2305
rect 32112 2297 32120 2305
rect 32160 2297 32168 2305
rect 32848 2297 32856 2305
rect 33392 2297 33400 2305
rect 33872 2297 33880 2305
rect 34368 2297 34376 2305
rect 35888 2297 35896 2305
rect 36464 2297 36472 2305
rect 40256 2297 40264 2305
rect 1704 2279 1712 2287
rect 1768 2279 1776 2287
rect 1928 2279 1936 2287
rect 2152 2279 2160 2287
rect 2168 2279 2176 2287
rect 2648 2279 2656 2287
rect 2968 2279 2976 2287
rect 3000 2279 3008 2287
rect 3096 2279 3104 2287
rect 3208 2279 3216 2287
rect 3640 2279 3648 2287
rect 3704 2279 3712 2287
rect 3960 2279 3968 2287
rect 3976 2279 3984 2287
rect 3992 2279 4000 2287
rect 6050 2273 6058 2281
rect 6546 2273 6554 2281
rect 7554 2273 7562 2281
rect 7618 2273 7626 2281
rect 7730 2273 7738 2281
rect 7746 2273 7754 2281
rect 8306 2273 8314 2281
rect 10082 2273 10090 2281
rect 10690 2273 10698 2281
rect 12890 2279 12898 2287
rect 13450 2279 13458 2287
rect 13722 2279 13730 2287
rect 13834 2279 13842 2287
rect 14026 2279 14034 2287
rect 14138 2279 14146 2287
rect 14282 2279 14290 2287
rect 14474 2279 14482 2287
rect 16154 2279 16162 2287
rect 16346 2279 16354 2287
rect 16778 2279 16786 2287
rect 20384 2280 20392 2288
rect 23760 2280 23768 2288
rect 24144 2280 24152 2288
rect 24320 2280 24328 2288
rect 24400 2280 24408 2288
rect 24768 2280 24776 2288
rect 25856 2280 25864 2288
rect 26272 2280 26280 2288
rect 38032 2277 38040 2285
rect 1752 2259 1760 2267
rect 2120 2259 2128 2267
rect 2712 2259 2720 2267
rect 7570 2253 7578 2261
rect 7650 2253 7658 2261
rect 8002 2253 8010 2261
rect 8130 2253 8138 2261
rect 8738 2253 8746 2261
rect 9362 2253 9370 2261
rect 9490 2253 9498 2261
rect 9906 2253 9914 2261
rect 10114 2253 10122 2261
rect 14746 2259 14754 2267
rect 14858 2259 14866 2267
rect 16762 2259 16770 2267
rect 17082 2259 17090 2267
rect 23760 2260 23768 2268
rect 25840 2260 25848 2268
rect 29460 2267 29472 2275
rect 29492 2267 29504 2275
rect 29508 2267 29520 2275
rect 29524 2267 29536 2275
rect 29552 2267 29564 2275
rect 29584 2267 29596 2275
rect 29600 2267 29612 2275
rect 29616 2267 29628 2275
rect 29648 2267 29660 2275
rect 29664 2267 29668 2275
rect 29740 2267 29752 2275
rect 29756 2267 29760 2275
rect 29772 2267 29784 2275
rect 29800 2267 29816 2275
rect 29832 2267 29880 2275
rect 29896 2267 29944 2275
rect 29960 2267 29972 2275
rect 29976 2267 29980 2275
rect 29992 2267 30004 2275
rect 30016 2267 30020 2275
rect 30024 2267 30036 2275
rect 30180 2267 30192 2275
rect 30196 2267 30200 2275
rect 30212 2267 30224 2275
rect 30244 2267 30256 2275
rect 30260 2267 30264 2275
rect 30276 2267 30288 2275
rect 30296 2267 30320 2275
rect 30336 2267 30348 2275
rect 30352 2267 30356 2275
rect 30368 2267 30380 2275
rect 30392 2267 30396 2275
rect 30400 2267 30412 2275
rect 30428 2267 30452 2275
rect 30460 2267 30472 2275
rect 30484 2267 30488 2275
rect 30492 2267 30504 2275
rect 30608 2267 30612 2275
rect 30616 2267 30628 2275
rect 30648 2267 30660 2275
rect 30664 2267 30668 2275
rect 30740 2267 30752 2275
rect 30756 2267 30760 2275
rect 30772 2267 30784 2275
rect 30800 2267 30816 2275
rect 30832 2267 30880 2275
rect 30896 2267 30912 2275
rect 30928 2267 30932 2275
rect 30936 2267 30948 2275
rect 30960 2267 30964 2275
rect 30968 2267 30972 2275
rect 31052 2267 31056 2275
rect 31060 2267 31064 2275
rect 31240 2267 31244 2275
rect 31248 2267 31252 2275
rect 31264 2267 31276 2275
rect 31280 2267 31292 2275
rect 31300 2267 31316 2275
rect 31332 2267 31336 2275
rect 31340 2267 31344 2275
rect 31356 2267 31368 2275
rect 31372 2267 31384 2275
rect 31392 2267 31408 2275
rect 31424 2267 31472 2275
rect 31488 2267 31504 2275
rect 31520 2267 31524 2275
rect 31528 2267 31540 2275
rect 31552 2267 31556 2275
rect 31560 2267 31564 2275
rect 31708 2267 31712 2275
rect 31716 2267 31720 2275
rect 31740 2267 31744 2275
rect 31748 2267 31752 2275
rect 31764 2267 31776 2275
rect 31780 2267 31784 2275
rect 31800 2267 31816 2275
rect 31832 2267 31864 2275
rect 31872 2267 31888 2275
rect 31904 2267 31920 2275
rect 31936 2267 31940 2275
rect 31944 2267 31956 2275
rect 31968 2267 31972 2275
rect 31976 2267 31980 2275
rect 31992 2267 32000 2275
rect 32012 2267 32036 2275
rect 32052 2267 32064 2275
rect 32068 2267 32072 2275
rect 32084 2267 32096 2275
rect 32108 2267 32112 2275
rect 32116 2267 32128 2275
rect 32144 2267 32168 2275
rect 32176 2267 32192 2275
rect 32208 2267 32212 2275
rect 32216 2267 32220 2275
rect 32240 2267 32244 2275
rect 32248 2267 32260 2275
rect 32264 2267 32276 2275
rect 32280 2267 32284 2275
rect 32300 2267 32324 2275
rect 32332 2267 32348 2275
rect 32356 2267 32380 2275
rect 32396 2267 32412 2275
rect 32428 2267 32440 2275
rect 32452 2267 32456 2275
rect 32460 2267 32472 2275
rect 32476 2267 32480 2275
rect 32492 2267 32504 2275
rect 32512 2267 32536 2275
rect 32552 2267 32564 2275
rect 32568 2267 32572 2275
rect 32584 2267 32596 2275
rect 32608 2267 32612 2275
rect 32616 2267 32628 2275
rect 32632 2267 32636 2275
rect 32648 2267 32660 2275
rect 32772 2267 32784 2275
rect 32788 2267 32792 2275
rect 32804 2267 32816 2275
rect 32836 2267 32848 2275
rect 32852 2267 32864 2275
rect 32868 2267 32880 2275
rect 32896 2267 32912 2275
rect 32928 2267 32940 2275
rect 32944 2267 32956 2275
rect 32960 2267 32972 2275
rect 32992 2267 33004 2275
rect 33020 2267 33044 2275
rect 33052 2267 33068 2275
rect 33084 2267 33088 2275
rect 33092 2267 33096 2275
rect 33108 2267 33120 2275
rect 33124 2267 33136 2275
rect 33148 2267 33152 2275
rect 33156 2267 33160 2275
rect 33172 2267 33184 2275
rect 33188 2267 33192 2275
rect 33208 2267 33224 2275
rect 33240 2267 33256 2275
rect 33264 2267 33296 2275
rect 33304 2267 33320 2275
rect 33328 2267 33340 2275
rect 33344 2267 33348 2275
rect 33368 2267 33372 2275
rect 33376 2267 33388 2275
rect 33396 2267 33412 2275
rect 33420 2267 33432 2275
rect 33436 2267 33440 2275
rect 33456 2267 33480 2275
rect 33488 2267 33504 2275
rect 33512 2267 33536 2275
rect 33552 2267 33564 2275
rect 33584 2267 33596 2275
rect 33608 2267 33612 2275
rect 33616 2267 33628 2275
rect 33632 2267 33636 2275
rect 33648 2267 33660 2275
rect 33680 2267 33692 2275
rect 33696 2267 33700 2275
rect 33712 2267 33724 2275
rect 33740 2267 33756 2275
rect 33764 2267 33796 2275
rect 33804 2267 33820 2275
rect 33832 2267 33848 2275
rect 33856 2267 33888 2275
rect 33896 2267 33912 2275
rect 33928 2267 33932 2275
rect 33936 2267 33940 2275
rect 33960 2267 33964 2275
rect 33968 2267 33980 2275
rect 33992 2267 33996 2275
rect 34000 2267 34004 2275
rect 34016 2267 34028 2275
rect 34032 2267 34036 2275
rect 34100 2267 34104 2275
rect 34108 2267 34112 2275
rect 34132 2267 34136 2275
rect 34140 2267 34144 2275
rect 34156 2267 34168 2275
rect 34172 2267 34184 2275
rect 34192 2267 34208 2275
rect 34224 2267 34240 2275
rect 34248 2267 34260 2275
rect 34264 2267 34276 2275
rect 34288 2267 34292 2275
rect 34296 2267 34300 2275
rect 34312 2267 34324 2275
rect 34328 2267 34332 2275
rect 34348 2267 34364 2275
rect 34380 2267 34396 2275
rect 34404 2267 34436 2275
rect 34444 2267 34456 2275
rect 34472 2267 34488 2275
rect 34496 2267 34528 2275
rect 34536 2267 34552 2275
rect 34560 2267 34592 2275
rect 34600 2267 34616 2275
rect 34632 2267 34644 2275
rect 34648 2267 34660 2275
rect 34664 2267 34676 2275
rect 34788 2267 34800 2275
rect 34812 2267 34816 2275
rect 34820 2267 34832 2275
rect 34836 2267 34840 2275
rect 34852 2267 34864 2275
rect 34876 2267 34880 2275
rect 34884 2267 34896 2275
rect 34900 2267 34904 2275
rect 34916 2267 34928 2275
rect 34940 2267 34944 2275
rect 34948 2267 34960 2275
rect 34980 2267 34992 2275
rect 35064 2267 35068 2275
rect 35072 2267 35084 2275
rect 35200 2267 35208 2275
rect 35212 2267 35224 2275
rect 35228 2267 35240 2275
rect 35260 2267 35272 2275
rect 35288 2267 35312 2275
rect 35320 2267 35336 2275
rect 35352 2267 35356 2275
rect 35360 2267 35364 2275
rect 35376 2267 35388 2275
rect 35392 2267 35404 2275
rect 35416 2267 35420 2275
rect 35424 2267 35428 2275
rect 35444 2267 35460 2275
rect 35468 2267 35492 2275
rect 35508 2267 35524 2275
rect 35532 2267 35564 2275
rect 35572 2267 35588 2275
rect 35596 2267 35620 2275
rect 35636 2267 35640 2275
rect 35644 2267 35656 2275
rect 35668 2267 35672 2275
rect 35676 2267 35680 2275
rect 35808 2267 35812 2275
rect 35816 2267 35828 2275
rect 35832 2267 35844 2275
rect 35848 2267 35852 2275
rect 35872 2267 35876 2275
rect 35880 2267 35884 2275
rect 35900 2267 35916 2275
rect 35924 2267 35948 2275
rect 35964 2267 35976 2275
rect 35980 2267 35984 2275
rect 36000 2267 36008 2275
rect 36020 2267 36024 2275
rect 36028 2267 36040 2275
rect 36044 2267 36048 2275
rect 36060 2267 36072 2275
rect 36088 2267 36100 2275
rect 36112 2267 36116 2275
rect 36120 2267 36132 2275
rect 36136 2267 36140 2275
rect 36152 2267 36164 2275
rect 36244 2267 36256 2275
rect 36276 2267 36288 2275
rect 36292 2267 36304 2275
rect 36308 2267 36320 2275
rect 36340 2267 36352 2275
rect 36368 2267 36392 2275
rect 36400 2267 36416 2275
rect 36432 2267 36436 2275
rect 36440 2267 36444 2275
rect 36456 2267 36468 2275
rect 36472 2267 36484 2275
rect 36496 2267 36500 2275
rect 36504 2267 36508 2275
rect 36524 2267 36540 2275
rect 36548 2267 36560 2275
rect 36564 2267 36576 2275
rect 36588 2267 36592 2275
rect 36596 2267 36600 2275
rect 36620 2267 36624 2275
rect 36628 2267 36632 2275
rect 36728 2267 36732 2275
rect 36736 2267 36740 2275
rect 36752 2267 36764 2275
rect 36768 2267 36772 2275
rect 36980 2267 36984 2275
rect 36988 2267 36992 2275
rect 37004 2267 37016 2275
rect 37020 2267 37024 2275
rect 37040 2267 37056 2275
rect 37072 2267 37120 2275
rect 37136 2267 37160 2275
rect 37168 2267 37180 2275
rect 37192 2267 37196 2275
rect 37200 2267 37212 2275
rect 37216 2267 37220 2275
rect 37232 2267 37244 2275
rect 37260 2267 37276 2275
rect 37292 2267 37316 2275
rect 37324 2267 37340 2275
rect 37348 2267 37360 2275
rect 37364 2267 37368 2275
rect 37388 2267 37392 2275
rect 37396 2267 37408 2275
rect 37416 2267 37432 2275
rect 37440 2267 37452 2275
rect 37456 2267 37460 2275
rect 37480 2267 37484 2275
rect 37488 2267 37500 2275
rect 37508 2267 37524 2275
rect 37532 2267 37556 2275
rect 37572 2267 37588 2275
rect 37604 2267 37616 2275
rect 37628 2267 37632 2275
rect 37636 2267 37648 2275
rect 37652 2267 37656 2275
rect 37668 2267 37680 2275
rect 37720 2267 37724 2275
rect 37728 2267 37740 2275
rect 37744 2267 37748 2275
rect 37760 2267 37772 2275
rect 38292 2267 38304 2275
rect 38308 2267 38312 2275
rect 38324 2267 38336 2275
rect 38356 2267 38368 2275
rect 38376 2267 38400 2275
rect 38416 2267 38428 2275
rect 38448 2267 38460 2275
rect 38472 2267 38476 2275
rect 38480 2267 38492 2275
rect 38604 2267 38616 2275
rect 38628 2267 38632 2275
rect 38636 2267 38648 2275
rect 38652 2267 38656 2275
rect 38668 2267 38680 2275
rect 38700 2267 38712 2275
rect 38728 2267 38752 2275
rect 38760 2267 38776 2275
rect 38784 2267 38796 2275
rect 38800 2267 38804 2275
rect 38824 2267 38828 2275
rect 38832 2267 38844 2275
rect 38848 2267 38860 2275
rect 38864 2267 38868 2275
rect 38884 2267 38888 2275
rect 38892 2267 38896 2275
rect 38916 2267 38920 2275
rect 38924 2267 38936 2275
rect 38940 2267 38952 2275
rect 38956 2267 38960 2275
rect 38980 2267 38984 2275
rect 38988 2267 39000 2275
rect 39004 2267 39016 2275
rect 39020 2267 39024 2275
rect 39044 2267 39048 2275
rect 39052 2267 39056 2275
rect 39076 2267 39080 2275
rect 39084 2267 39088 2275
rect 39108 2267 39112 2275
rect 39116 2267 39120 2275
rect 39140 2267 39144 2275
rect 39148 2267 39160 2275
rect 39164 2267 39176 2275
rect 39180 2267 39184 2275
rect 39232 2267 39236 2275
rect 39240 2267 39252 2275
rect 39256 2267 39268 2275
rect 39272 2267 39276 2275
rect 39296 2267 39300 2275
rect 39304 2267 39308 2275
rect 39484 2267 39488 2275
rect 39492 2267 39496 2275
rect 39508 2267 39520 2275
rect 39524 2267 39528 2275
rect 39576 2267 39580 2275
rect 39584 2267 39588 2275
rect 39600 2267 39612 2275
rect 39616 2267 39620 2275
rect 39636 2267 39652 2275
rect 39668 2267 39684 2275
rect 39692 2267 39724 2275
rect 39732 2267 39748 2275
rect 39756 2267 39768 2275
rect 39772 2267 39776 2275
rect 39796 2267 39800 2275
rect 39804 2267 39816 2275
rect 39824 2267 39840 2275
rect 39848 2267 39872 2275
rect 39888 2267 39892 2275
rect 39896 2267 39908 2275
rect 39920 2267 39924 2275
rect 39928 2267 39932 2275
rect 40076 2267 40080 2275
rect 40084 2267 40088 2275
rect 40100 2267 40112 2275
rect 40116 2267 40120 2275
rect 40168 2267 40172 2275
rect 40176 2267 40180 2275
rect 40192 2267 40204 2275
rect 40208 2267 40212 2275
rect 40232 2267 40236 2275
rect 40240 2267 40244 2275
rect 40264 2267 40268 2275
rect 40272 2267 40276 2275
rect 40296 2267 40300 2275
rect 40304 2267 40316 2275
rect 40328 2267 40332 2275
rect 40336 2267 40340 2275
rect 40500 2267 40504 2275
rect 40508 2267 40520 2275
rect 40532 2267 40536 2275
rect 40540 2267 40544 2275
rect 40592 2267 40596 2275
rect 40600 2267 40612 2275
rect 40624 2267 40628 2275
rect 40632 2267 40636 2275
rect 40648 2267 40660 2275
rect 40664 2267 40668 2275
rect 40716 2267 40720 2275
rect 40724 2267 40728 2275
rect 40740 2267 40752 2275
rect 40756 2267 40760 2275
rect 40776 2267 40792 2275
rect 19382 2250 19386 2258
rect 19472 2250 19480 2258
rect 19810 2252 19812 2260
rect 20024 2252 20026 2260
rect 20848 2252 20850 2260
rect 25572 2256 25574 2260
rect 25578 2252 25580 2256
rect 25706 2250 25710 2258
rect 25796 2250 25804 2258
rect 26626 2256 26628 2260
rect 27054 2256 27056 2260
rect 26632 2252 26634 2256
rect 27060 2252 27062 2256
rect 27150 2250 27158 2258
rect 27300 2250 27306 2258
rect 27364 2250 27372 2258
rect 27514 2250 27520 2258
rect 27578 2250 27586 2258
rect 27728 2250 27734 2258
rect 27792 2250 27800 2258
rect 27942 2250 27948 2258
rect 28006 2250 28020 2258
rect 28220 2250 28234 2258
rect 28434 2250 28448 2258
rect 32656 2257 32664 2265
rect 33936 2257 33944 2265
rect 34032 2257 34040 2265
rect 34112 2257 34120 2265
rect 34128 2257 34136 2265
rect 664 2239 672 2247
rect 2776 2239 2784 2247
rect 3256 2239 3264 2247
rect 4232 2239 4240 2247
rect 4424 2239 4432 2247
rect 7106 2233 7114 2241
rect 7906 2233 7914 2241
rect 8274 2233 8282 2241
rect 8626 2233 8634 2241
rect 16138 2239 16146 2247
rect 25648 2240 25656 2248
rect 27104 2240 27112 2248
rect 29648 2237 29656 2245
rect 30576 2237 30584 2245
rect 31968 2237 31976 2245
rect 37184 2237 37192 2245
rect 37264 2237 37272 2245
rect 37808 2237 37816 2245
rect 38032 2237 38040 2245
rect 38864 2237 38872 2245
rect 39904 2237 39912 2245
rect 568 2219 576 2227
rect 1080 2219 1088 2227
rect 1256 2219 1264 2227
rect 1400 2219 1408 2227
rect 1432 2219 1440 2227
rect 1496 2219 1504 2227
rect 1624 2219 1632 2227
rect 1720 2219 1728 2227
rect 1736 2219 1744 2227
rect 1768 2219 1776 2227
rect 1848 2219 1856 2227
rect 2168 2219 2176 2227
rect 2184 2219 2192 2227
rect 2264 2219 2272 2227
rect 2344 2219 2352 2227
rect 2376 2219 2384 2227
rect 3880 2219 3888 2227
rect 3976 2219 3984 2227
rect 4440 2219 4448 2227
rect 4504 2219 4512 2227
rect 6066 2213 6074 2221
rect 6402 2213 6410 2221
rect 6418 2213 6426 2221
rect 6434 2213 6442 2221
rect 6866 2213 6874 2221
rect 8210 2213 8218 2221
rect 8866 2213 8874 2221
rect 9074 2213 9082 2221
rect 12874 2219 12882 2227
rect 12938 2219 12946 2227
rect 13066 2219 13074 2227
rect 13962 2219 13970 2227
rect 14090 2219 14098 2227
rect 14362 2219 14370 2227
rect 14938 2219 14946 2227
rect 15754 2219 15762 2227
rect 16218 2219 16226 2227
rect 16602 2219 16610 2227
rect 17210 2219 17218 2227
rect 17546 2219 17554 2227
rect 19312 2220 19320 2228
rect 20768 2220 20776 2228
rect 23120 2220 23128 2228
rect 23952 2220 23960 2228
rect 24512 2220 24520 2228
rect 29984 2217 29992 2225
rect 30256 2217 30264 2225
rect 31440 2217 31448 2225
rect 32464 2217 32472 2225
rect 32704 2217 32712 2225
rect 33280 2217 33288 2225
rect 35440 2217 35448 2225
rect 38128 2217 38136 2225
rect 38480 2217 38488 2225
rect 38576 2217 38584 2225
rect 38688 2217 38696 2225
rect 38784 2217 38792 2225
rect 39296 2217 39304 2225
rect 40096 2217 40104 2225
rect 40304 2217 40312 2225
rect 440 2199 448 2207
rect 472 2199 480 2207
rect 520 2199 528 2207
rect 536 2199 544 2207
rect 584 2199 592 2207
rect 616 2199 624 2207
rect 632 2199 640 2207
rect 664 2199 672 2207
rect 760 2199 768 2207
rect 792 2199 800 2207
rect 952 2199 960 2207
rect 1160 2199 1168 2207
rect 1304 2199 1312 2207
rect 1368 2199 1376 2207
rect 1784 2199 1792 2207
rect 1816 2199 1824 2207
rect 2024 2199 2032 2207
rect 2056 2199 2064 2207
rect 2088 2199 2096 2207
rect 2120 2199 2128 2207
rect 2200 2199 2208 2207
rect 2216 2199 2224 2207
rect 2248 2199 2256 2207
rect 2312 2199 2320 2207
rect 2328 2199 2336 2207
rect 2440 2199 2448 2207
rect 2568 2199 2576 2207
rect 2648 2199 2656 2207
rect 2680 2199 2688 2207
rect 2808 2199 2816 2207
rect 2856 2199 2864 2207
rect 2888 2199 2896 2207
rect 2952 2199 2960 2207
rect 2968 2199 2976 2207
rect 3032 2199 3040 2207
rect 3144 2199 3152 2207
rect 3320 2199 3328 2207
rect 3352 2199 3360 2207
rect 3448 2199 3456 2207
rect 3464 2199 3472 2207
rect 3560 2199 3568 2207
rect 3720 2199 3728 2207
rect 3848 2199 3856 2207
rect 3976 2199 3984 2207
rect 4104 2199 4112 2207
rect 4184 2199 4192 2207
rect 4328 2199 4336 2207
rect 4344 2199 4352 2207
rect 4552 2199 4560 2207
rect 5890 2193 5898 2201
rect 6098 2193 6106 2201
rect 6178 2193 6186 2201
rect 6514 2193 6522 2201
rect 6882 2193 6890 2201
rect 7010 2193 7018 2201
rect 7042 2193 7050 2201
rect 7346 2193 7354 2201
rect 7378 2193 7386 2201
rect 7410 2193 7418 2201
rect 7778 2193 7786 2201
rect 7890 2193 7898 2201
rect 8226 2193 8234 2201
rect 8434 2193 8442 2201
rect 8530 2193 8538 2201
rect 8850 2193 8858 2201
rect 9058 2193 9066 2201
rect 9074 2193 9082 2201
rect 9426 2193 9434 2201
rect 9826 2193 9834 2201
rect 9842 2193 9850 2201
rect 9954 2193 9962 2201
rect 9970 2193 9978 2201
rect 10018 2193 10026 2201
rect 10098 2193 10106 2201
rect 10418 2193 10426 2201
rect 10466 2193 10474 2201
rect 10818 2193 10826 2201
rect 14490 2199 14498 2207
rect 14682 2199 14690 2207
rect 15498 2199 15506 2207
rect 18896 2200 18904 2208
rect 19472 2200 19480 2208
rect 20160 2200 20168 2208
rect 24768 2200 24776 2208
rect 24912 2200 24920 2208
rect 25488 2200 25496 2208
rect 26256 2200 26264 2208
rect 29504 2197 29512 2205
rect 30368 2197 30376 2205
rect 31600 2197 31608 2205
rect 32240 2197 32248 2205
rect 32544 2197 32552 2205
rect 32624 2197 32632 2205
rect 32880 2197 32888 2205
rect 33344 2197 33352 2205
rect 33776 2197 33784 2205
rect 34192 2197 34200 2205
rect 34560 2197 34568 2205
rect 34960 2197 34968 2205
rect 35136 2197 35144 2205
rect 35856 2197 35864 2205
rect 36304 2197 36312 2205
rect 37456 2197 37464 2205
rect 40032 2197 40040 2205
rect 472 2179 480 2187
rect 504 2179 512 2187
rect 840 2179 848 2187
rect 1480 2179 1488 2187
rect 1592 2179 1600 2187
rect 1704 2179 1712 2187
rect 1800 2179 1808 2187
rect 1912 2179 1920 2187
rect 3992 2179 4000 2187
rect 4008 2179 4016 2187
rect 4072 2179 4080 2187
rect 4216 2179 4224 2187
rect 4328 2179 4336 2187
rect 4376 2179 4384 2187
rect 4472 2179 4480 2187
rect 5730 2173 5738 2181
rect 6034 2173 6042 2181
rect 7026 2173 7034 2181
rect 7922 2173 7930 2181
rect 8946 2173 8954 2181
rect 10466 2173 10474 2181
rect 10578 2173 10586 2181
rect 12090 2179 12098 2187
rect 12154 2179 12162 2187
rect 12330 2179 12338 2187
rect 12426 2179 12434 2187
rect 12458 2179 12466 2187
rect 12474 2179 12482 2187
rect 12506 2179 12514 2187
rect 12842 2179 12850 2187
rect 12890 2179 12898 2187
rect 13498 2179 13506 2187
rect 13578 2179 13586 2187
rect 13594 2179 13602 2187
rect 14106 2179 14114 2187
rect 14426 2179 14434 2187
rect 14538 2179 14546 2187
rect 14618 2179 14626 2187
rect 14810 2179 14818 2187
rect 15034 2179 15042 2187
rect 15082 2179 15090 2187
rect 15962 2179 15970 2187
rect 16490 2179 16498 2187
rect 16730 2179 16738 2187
rect 16970 2179 16978 2187
rect 16986 2179 16994 2187
rect 17354 2179 17362 2187
rect 17434 2179 17442 2187
rect 17466 2179 17474 2187
rect 17498 2179 17506 2187
rect 19184 2180 19192 2188
rect 19696 2180 19704 2188
rect 19728 2180 19736 2188
rect 19888 2180 19896 2188
rect 19920 2180 19928 2188
rect 20304 2180 20312 2188
rect 20736 2180 20744 2188
rect 21136 2180 21144 2188
rect 21424 2180 21432 2188
rect 21456 2180 21464 2188
rect 23600 2180 23608 2188
rect 24400 2180 24408 2188
rect 24432 2180 24440 2188
rect 24624 2180 24632 2188
rect 25824 2180 25832 2188
rect 26112 2180 26120 2188
rect 26752 2180 26760 2188
rect 28224 2180 28232 2188
rect 28256 2180 28264 2188
rect 32768 2177 32776 2185
rect 32992 2177 33000 2185
rect 33248 2177 33256 2185
rect 36336 2177 36344 2185
rect 696 2159 704 2167
rect 760 2159 768 2167
rect 888 2159 896 2167
rect 1192 2159 1200 2167
rect 1240 2159 1248 2167
rect 1288 2159 1296 2167
rect 1464 2159 1472 2167
rect 1608 2159 1616 2167
rect 1720 2159 1728 2167
rect 1992 2159 2000 2167
rect 2552 2159 2560 2167
rect 2792 2159 2800 2167
rect 3992 2159 4000 2167
rect 4216 2159 4224 2167
rect 5810 2153 5818 2161
rect 6050 2153 6058 2161
rect 6082 2153 6090 2161
rect 6130 2153 6138 2161
rect 6162 2153 6170 2161
rect 6610 2153 6618 2161
rect 6770 2153 6778 2161
rect 6818 2153 6826 2161
rect 7906 2153 7914 2161
rect 8242 2153 8250 2161
rect 8386 2153 8394 2161
rect 8530 2153 8538 2161
rect 8722 2153 8730 2161
rect 8818 2153 8826 2161
rect 8866 2153 8874 2161
rect 9314 2153 9322 2161
rect 9970 2153 9978 2161
rect 10066 2153 10074 2161
rect 10146 2153 10154 2161
rect 10162 2153 10170 2161
rect 10226 2153 10234 2161
rect 10706 2153 10714 2161
rect 10834 2153 10842 2161
rect 13994 2159 14002 2167
rect 14010 2159 14018 2167
rect 14410 2159 14418 2167
rect 14714 2159 14722 2167
rect 14794 2159 14802 2167
rect 16394 2159 16402 2167
rect 16410 2159 16418 2167
rect 16586 2159 16594 2167
rect 16666 2159 16674 2167
rect 16842 2159 16850 2167
rect 16970 2159 16978 2167
rect 17050 2159 17058 2167
rect 23984 2160 23992 2168
rect 25456 2160 25464 2168
rect 29472 2157 29480 2165
rect 29696 2157 29704 2165
rect 29808 2157 29816 2165
rect 29904 2157 29912 2165
rect 30416 2157 30424 2165
rect 30880 2157 30888 2165
rect 31472 2157 31480 2165
rect 31920 2157 31928 2165
rect 33472 2157 33480 2165
rect 34976 2157 34984 2165
rect 35088 2157 35096 2165
rect 36048 2157 36056 2165
rect 36256 2157 36264 2165
rect 39936 2157 39944 2165
rect 40432 2157 40440 2165
rect 24838 2148 24845 2153
rect 696 2139 704 2147
rect 728 2139 736 2147
rect 968 2139 976 2147
rect 1224 2139 1232 2147
rect 1272 2139 1280 2147
rect 3208 2139 3216 2147
rect 3320 2139 3328 2147
rect 3368 2139 3376 2147
rect 3512 2139 3520 2147
rect 3912 2139 3920 2147
rect 4376 2139 4384 2147
rect 4408 2139 4416 2147
rect 4456 2139 4464 2147
rect 4584 2139 4592 2147
rect 4616 2139 4624 2147
rect 6002 2133 6010 2141
rect 6194 2133 6202 2141
rect 6306 2133 6314 2141
rect 7218 2133 7226 2141
rect 9106 2133 9114 2141
rect 10162 2133 10170 2141
rect 10418 2133 10426 2141
rect 10882 2133 10890 2141
rect 11994 2139 12002 2147
rect 12218 2139 12226 2147
rect 12442 2139 12450 2147
rect 12522 2139 12530 2147
rect 13322 2139 13330 2147
rect 13434 2139 13442 2147
rect 13770 2139 13778 2147
rect 13914 2139 13922 2147
rect 14442 2139 14450 2147
rect 15130 2139 15138 2147
rect 15530 2139 15538 2147
rect 15626 2139 15634 2147
rect 15722 2139 15730 2147
rect 15850 2139 15858 2147
rect 15930 2139 15938 2147
rect 16026 2139 16034 2147
rect 16170 2139 16178 2147
rect 16266 2139 16274 2147
rect 16602 2139 16610 2147
rect 16634 2139 16642 2147
rect 16906 2139 16914 2147
rect 17002 2139 17010 2147
rect 17018 2139 17026 2147
rect 17226 2139 17234 2147
rect 17498 2139 17506 2147
rect 19152 2140 19160 2148
rect 20112 2140 20120 2148
rect 22288 2140 22296 2148
rect 22864 2140 22872 2148
rect 23296 2140 23304 2148
rect 23360 2140 23368 2148
rect 23792 2140 23800 2148
rect 24208 2140 24216 2148
rect 24416 2140 24424 2148
rect 25648 2140 25656 2148
rect 25824 2140 25832 2148
rect 25904 2140 25912 2148
rect 26096 2140 26104 2148
rect 26960 2140 26968 2148
rect 27376 2140 27384 2148
rect 37680 2137 37688 2145
rect 38512 2137 38520 2145
rect 38896 2137 38904 2145
rect 1432 2119 1440 2127
rect 2152 2119 2160 2127
rect 2504 2119 2512 2127
rect 2648 2119 2656 2127
rect 3000 2119 3008 2127
rect 3064 2119 3072 2127
rect 7538 2113 7546 2121
rect 7666 2113 7674 2121
rect 7698 2113 7706 2121
rect 7778 2113 7786 2121
rect 8386 2113 8394 2121
rect 10562 2113 10570 2121
rect 10610 2113 10618 2121
rect 10834 2113 10842 2121
rect 13114 2119 13122 2127
rect 13130 2119 13138 2127
rect 15386 2119 15394 2127
rect 19328 2120 19336 2128
rect 23584 2120 23592 2128
rect 27392 2120 27400 2128
rect 1176 2099 1184 2107
rect 2120 2099 2128 2107
rect 3352 2099 3360 2107
rect 3992 2099 4000 2107
rect 7282 2093 7290 2101
rect 9698 2093 9706 2101
rect 9714 2093 9722 2101
rect 12730 2099 12738 2107
rect 14602 2099 14610 2107
rect 17130 2099 17138 2107
rect 18720 2100 18728 2108
rect 488 2079 496 2087
rect 552 2079 560 2087
rect 600 2079 608 2087
rect 648 2079 656 2087
rect 1288 2079 1296 2087
rect 1384 2079 1392 2087
rect 1896 2079 1904 2087
rect 1944 2079 1952 2087
rect 2040 2079 2048 2087
rect 2824 2079 2832 2087
rect 2840 2079 2848 2087
rect 2872 2079 2880 2087
rect 3048 2079 3056 2087
rect 3064 2079 3072 2087
rect 3160 2079 3168 2087
rect 3432 2079 3440 2087
rect 3752 2079 3760 2087
rect 3832 2079 3840 2087
rect 3864 2079 3872 2087
rect 4440 2079 4448 2087
rect 7858 2073 7866 2081
rect 9442 2073 9450 2081
rect 9490 2073 9498 2081
rect 9586 2073 9594 2081
rect 9778 2073 9786 2081
rect 9986 2073 9994 2081
rect 10498 2073 10506 2081
rect 12698 2079 12706 2087
rect 24368 2080 24376 2088
rect 32368 2077 32376 2085
rect 2104 2059 2112 2067
rect 2536 2059 2544 2067
rect 8018 2053 8026 2061
rect 8386 2053 8394 2061
rect 8402 2053 8410 2061
rect 9026 2053 9034 2061
rect 9186 2053 9194 2061
rect 14714 2059 14722 2067
rect 26912 2060 26920 2068
rect 29420 2067 29424 2075
rect 29428 2067 29440 2075
rect 29444 2067 29448 2075
rect 29488 2067 29500 2075
rect 29512 2067 29516 2075
rect 29520 2067 29532 2075
rect 29536 2067 29540 2075
rect 29604 2067 29608 2075
rect 29612 2067 29624 2075
rect 29628 2067 29632 2075
rect 29644 2067 29656 2075
rect 29668 2067 29672 2075
rect 29676 2067 29688 2075
rect 29704 2067 29728 2075
rect 29736 2067 29748 2075
rect 29760 2067 29764 2075
rect 29768 2067 29780 2075
rect 29796 2067 29808 2075
rect 29812 2067 29816 2075
rect 29828 2067 29840 2075
rect 29852 2067 29856 2075
rect 29860 2067 29872 2075
rect 29892 2067 29904 2075
rect 29916 2067 29920 2075
rect 29924 2067 29936 2075
rect 29956 2067 29968 2075
rect 29972 2067 29984 2075
rect 29988 2067 30000 2075
rect 30020 2067 30032 2075
rect 30036 2067 30040 2075
rect 30052 2067 30064 2075
rect 30084 2067 30096 2075
rect 30116 2067 30128 2075
rect 30140 2067 30144 2075
rect 30148 2067 30160 2075
rect 30180 2067 30192 2075
rect 30196 2067 30200 2075
rect 30212 2067 30224 2075
rect 30240 2067 30256 2075
rect 30272 2067 30320 2075
rect 30332 2067 30348 2075
rect 30364 2067 30412 2075
rect 30428 2067 30444 2075
rect 30456 2067 30504 2075
rect 30516 2067 30532 2075
rect 30548 2067 30596 2075
rect 30612 2067 30624 2075
rect 30640 2067 30688 2075
rect 30704 2067 30720 2075
rect 30732 2067 30780 2075
rect 30796 2067 30808 2075
rect 30824 2067 30872 2075
rect 30888 2067 30904 2075
rect 30920 2067 30932 2075
rect 30944 2067 30948 2075
rect 30952 2067 30964 2075
rect 31508 2067 31512 2075
rect 31516 2067 31520 2075
rect 31532 2067 31544 2075
rect 31548 2067 31552 2075
rect 31568 2067 31584 2075
rect 31600 2067 31616 2075
rect 31624 2067 31656 2075
rect 31672 2067 31684 2075
rect 31688 2067 31692 2075
rect 31704 2067 31716 2075
rect 31728 2067 31732 2075
rect 31736 2067 31740 2075
rect 31996 2067 32000 2075
rect 32004 2067 32008 2075
rect 32088 2067 32092 2075
rect 32096 2067 32100 2075
rect 32120 2067 32124 2075
rect 32128 2067 32132 2075
rect 32180 2067 32184 2075
rect 32188 2067 32192 2075
rect 32304 2067 32308 2075
rect 32312 2067 32324 2075
rect 32328 2067 32340 2075
rect 32344 2067 32348 2075
rect 32368 2067 32372 2075
rect 32376 2067 32380 2075
rect 32396 2067 32412 2075
rect 32420 2067 32444 2075
rect 32460 2067 32484 2075
rect 32492 2067 32504 2075
rect 32512 2067 32536 2075
rect 32552 2067 32576 2075
rect 32584 2067 32596 2075
rect 32608 2067 32612 2075
rect 32616 2067 32628 2075
rect 32632 2067 32636 2075
rect 32648 2067 32660 2075
rect 32740 2067 32752 2075
rect 32772 2067 32784 2075
rect 32788 2067 32792 2075
rect 32804 2067 32816 2075
rect 32836 2067 32848 2075
rect 32856 2067 32888 2075
rect 32896 2067 32912 2075
rect 32928 2067 32940 2075
rect 32948 2067 32980 2075
rect 32988 2067 33004 2075
rect 33020 2067 33036 2075
rect 33052 2067 33056 2075
rect 33060 2067 33072 2075
rect 33084 2067 33088 2075
rect 33092 2067 33096 2075
rect 33108 2067 33120 2075
rect 33124 2067 33128 2075
rect 33192 2067 33196 2075
rect 33200 2067 33204 2075
rect 33316 2067 33320 2075
rect 33324 2067 33336 2075
rect 33340 2067 33352 2075
rect 33356 2067 33360 2075
rect 33380 2067 33384 2075
rect 33388 2067 33392 2075
rect 33408 2067 33412 2075
rect 33416 2067 33428 2075
rect 33432 2067 33444 2075
rect 33448 2067 33452 2075
rect 33468 2067 33472 2075
rect 33476 2067 33480 2075
rect 33500 2067 33504 2075
rect 33508 2067 33520 2075
rect 33524 2067 33536 2075
rect 33540 2067 33544 2075
rect 33720 2067 33724 2075
rect 33728 2067 33732 2075
rect 33744 2067 33756 2075
rect 33760 2067 33772 2075
rect 33784 2067 33788 2075
rect 33792 2067 33796 2075
rect 33816 2067 33820 2075
rect 33824 2067 33828 2075
rect 34244 2067 34248 2075
rect 34252 2067 34256 2075
rect 34320 2067 34324 2075
rect 34328 2067 34332 2075
rect 34352 2067 34356 2075
rect 34360 2067 34364 2075
rect 34376 2067 34388 2075
rect 34392 2067 34396 2075
rect 34412 2067 34436 2075
rect 34444 2067 34460 2075
rect 34468 2067 34480 2075
rect 34484 2067 34488 2075
rect 34508 2067 34512 2075
rect 34516 2067 34528 2075
rect 34536 2067 34552 2075
rect 34560 2067 34592 2075
rect 34600 2067 34616 2075
rect 34632 2067 34656 2075
rect 34664 2067 34680 2075
rect 34696 2067 34712 2075
rect 34720 2067 34744 2075
rect 34760 2067 34776 2075
rect 34784 2067 34816 2075
rect 34824 2067 34840 2075
rect 34856 2067 34880 2075
rect 34888 2067 34904 2075
rect 34920 2067 34968 2075
rect 34984 2067 35000 2075
rect 35012 2067 35060 2075
rect 35076 2067 35080 2075
rect 35084 2067 35088 2075
rect 35104 2067 35152 2075
rect 35168 2067 35184 2075
rect 35200 2067 35204 2075
rect 35208 2067 35220 2075
rect 35232 2067 35236 2075
rect 35240 2067 35244 2075
rect 35264 2067 35268 2075
rect 35272 2067 35276 2075
rect 35340 2067 35344 2075
rect 35348 2067 35360 2075
rect 35372 2067 35376 2075
rect 35380 2067 35384 2075
rect 35396 2067 35408 2075
rect 35412 2067 35416 2075
rect 35436 2067 35440 2075
rect 35444 2067 35448 2075
rect 35468 2067 35472 2075
rect 35476 2067 35480 2075
rect 35500 2067 35504 2075
rect 35508 2067 35520 2075
rect 35532 2067 35536 2075
rect 35540 2067 35544 2075
rect 35556 2067 35568 2075
rect 35572 2067 35584 2075
rect 35596 2067 35600 2075
rect 35604 2067 35608 2075
rect 35624 2067 35628 2075
rect 35632 2067 35636 2075
rect 35648 2067 35660 2075
rect 35664 2067 35676 2075
rect 35684 2067 35700 2075
rect 35716 2067 35720 2075
rect 35724 2067 35728 2075
rect 35740 2067 35752 2075
rect 35756 2067 35768 2075
rect 35780 2067 35784 2075
rect 35788 2067 35792 2075
rect 35808 2067 35824 2075
rect 35832 2067 35856 2075
rect 35872 2067 35888 2075
rect 35904 2067 35916 2075
rect 35920 2067 35932 2075
rect 35936 2067 35948 2075
rect 36000 2067 36008 2075
rect 36012 2067 36024 2075
rect 36028 2067 36040 2075
rect 36060 2067 36072 2075
rect 36088 2067 36100 2075
rect 36104 2067 36116 2075
rect 36120 2067 36132 2075
rect 36152 2067 36164 2075
rect 36244 2067 36256 2075
rect 36268 2067 36272 2075
rect 36276 2067 36288 2075
rect 36292 2067 36296 2075
rect 36360 2067 36364 2075
rect 36368 2067 36380 2075
rect 36384 2067 36388 2075
rect 36428 2067 36440 2075
rect 36452 2067 36456 2075
rect 36460 2067 36472 2075
rect 36476 2067 36480 2075
rect 36492 2067 36504 2075
rect 36516 2067 36520 2075
rect 36524 2067 36536 2075
rect 36552 2067 36564 2075
rect 36568 2067 36572 2075
rect 36584 2067 36596 2075
rect 36608 2067 36612 2075
rect 36616 2067 36628 2075
rect 36644 2067 36656 2075
rect 36660 2067 36664 2075
rect 36676 2067 36688 2075
rect 36700 2067 36704 2075
rect 36708 2067 36720 2075
rect 36736 2067 36748 2075
rect 36752 2067 36756 2075
rect 36768 2067 36780 2075
rect 36792 2067 36796 2075
rect 36800 2067 36812 2075
rect 36956 2067 36968 2075
rect 36972 2067 36976 2075
rect 37048 2067 37060 2075
rect 37080 2067 37092 2075
rect 37096 2067 37100 2075
rect 37112 2067 37124 2075
rect 37136 2067 37140 2075
rect 37144 2067 37156 2075
rect 37172 2067 37196 2075
rect 37204 2067 37216 2075
rect 37228 2067 37232 2075
rect 37236 2067 37248 2075
rect 37268 2067 37280 2075
rect 37292 2067 37296 2075
rect 37300 2067 37312 2075
rect 37332 2067 37344 2075
rect 37348 2067 37360 2075
rect 37364 2067 37376 2075
rect 37396 2067 37408 2075
rect 37416 2067 37448 2075
rect 37456 2067 37472 2075
rect 37488 2067 37504 2075
rect 37520 2067 37524 2075
rect 37528 2067 37540 2075
rect 37552 2067 37556 2075
rect 37560 2067 37564 2075
rect 37576 2067 37588 2075
rect 37592 2067 37596 2075
rect 37692 2067 37696 2075
rect 37700 2067 37704 2075
rect 37716 2067 37728 2075
rect 37732 2067 37736 2075
rect 37756 2067 37760 2075
rect 37764 2067 37768 2075
rect 37784 2067 37832 2075
rect 37848 2067 37852 2075
rect 37856 2067 37860 2075
rect 37880 2067 37884 2075
rect 37888 2067 37900 2075
rect 37912 2067 37916 2075
rect 37920 2067 37924 2075
rect 37944 2067 37948 2075
rect 37952 2067 37956 2075
rect 38020 2067 38024 2075
rect 38028 2067 38040 2075
rect 38052 2067 38056 2075
rect 38060 2067 38064 2075
rect 38112 2067 38116 2075
rect 38120 2067 38132 2075
rect 38144 2067 38148 2075
rect 38152 2067 38156 2075
rect 38284 2067 38288 2075
rect 38292 2067 38296 2075
rect 38308 2067 38320 2075
rect 38324 2067 38336 2075
rect 38348 2067 38352 2075
rect 38356 2067 38360 2075
rect 38376 2067 38392 2075
rect 38400 2067 38424 2075
rect 38440 2067 38456 2075
rect 38472 2067 38496 2075
rect 38504 2067 38520 2075
rect 38536 2067 38584 2075
rect 38600 2067 38604 2075
rect 38608 2067 38612 2075
rect 38624 2067 38636 2075
rect 38640 2067 38652 2075
rect 38664 2067 38668 2075
rect 38672 2067 38676 2075
rect 38804 2067 38808 2075
rect 38812 2067 38816 2075
rect 38828 2067 38840 2075
rect 38844 2067 38856 2075
rect 38868 2067 38872 2075
rect 38876 2067 38880 2075
rect 38896 2067 38900 2075
rect 38904 2067 38908 2075
rect 38920 2067 38932 2075
rect 38936 2067 38948 2075
rect 38956 2067 38972 2075
rect 38988 2067 39036 2075
rect 39052 2067 39068 2075
rect 39084 2067 39096 2075
rect 39108 2067 39112 2075
rect 39116 2067 39128 2075
rect 39148 2067 39160 2075
rect 39164 2067 39168 2075
rect 39240 2067 39252 2075
rect 39256 2067 39260 2075
rect 39492 2067 39504 2075
rect 39508 2067 39520 2075
rect 39524 2067 39536 2075
rect 39556 2067 39568 2075
rect 39584 2067 39608 2075
rect 39616 2067 39632 2075
rect 39648 2067 39652 2075
rect 39656 2067 39660 2075
rect 39672 2067 39684 2075
rect 39688 2067 39700 2075
rect 39712 2067 39716 2075
rect 39720 2067 39724 2075
rect 39736 2067 39748 2075
rect 39752 2067 39764 2075
rect 39772 2067 39788 2075
rect 39804 2067 39820 2075
rect 39828 2067 39840 2075
rect 39844 2067 39856 2075
rect 39868 2067 39872 2075
rect 39876 2067 39880 2075
rect 39900 2067 39904 2075
rect 39908 2067 39912 2075
rect 39932 2067 39936 2075
rect 39940 2067 39944 2075
rect 39964 2067 39968 2075
rect 39972 2067 39976 2075
rect 39988 2067 40000 2075
rect 40004 2067 40016 2075
rect 40028 2067 40032 2075
rect 40036 2067 40040 2075
rect 40052 2067 40064 2075
rect 40068 2067 40072 2075
rect 40120 2067 40124 2075
rect 40128 2067 40132 2075
rect 40144 2067 40156 2075
rect 40160 2067 40164 2075
rect 40244 2067 40248 2075
rect 40252 2067 40256 2075
rect 40276 2067 40280 2075
rect 40284 2067 40288 2075
rect 40300 2067 40312 2075
rect 40316 2067 40320 2075
rect 40336 2067 40360 2075
rect 40368 2067 40384 2075
rect 40392 2067 40416 2075
rect 40432 2067 40448 2075
rect 40456 2067 40480 2075
rect 40496 2067 40544 2075
rect 40560 2067 40564 2075
rect 40568 2067 40572 2075
rect 40588 2067 40636 2075
rect 40652 2067 40664 2075
rect 40680 2067 40728 2075
rect 40744 2067 40760 2075
rect 40768 2067 40792 2075
rect 18784 2050 18786 2058
rect 18792 2050 18794 2058
rect 19212 2050 19214 2058
rect 19220 2050 19222 2058
rect 19838 2050 19840 2058
rect 19846 2050 19848 2058
rect 20258 2050 20268 2058
rect 20472 2050 20482 2058
rect 24254 2050 24258 2058
rect 24262 2050 24266 2058
rect 24468 2050 24472 2058
rect 24476 2050 24480 2058
rect 24674 2050 24686 2058
rect 24888 2050 24900 2058
rect 25102 2050 25114 2058
rect 25530 2050 25542 2058
rect 25850 2050 25862 2058
rect 26072 2050 26076 2058
rect 26080 2050 26084 2058
rect 26148 2050 26152 2058
rect 26156 2050 26160 2058
rect 26392 2050 26398 2058
rect 26400 2050 26406 2058
rect 26468 2050 26474 2058
rect 26476 2050 26482 2058
rect 27226 2050 27238 2058
rect 27440 2050 27452 2058
rect 27654 2050 27666 2058
rect 27868 2050 27880 2058
rect 28082 2050 28094 2058
rect 28296 2050 28308 2058
rect 648 2039 656 2047
rect 2824 2039 2832 2047
rect 23584 2040 23592 2048
rect 23776 2040 23784 2048
rect 31072 2037 31080 2045
rect 32192 2037 32200 2045
rect 33584 2037 33592 2045
rect 34192 2037 34200 2045
rect 35712 2037 35720 2045
rect 37424 2037 37432 2045
rect 39744 2037 39752 2045
rect 40304 2037 40312 2045
rect 760 2019 768 2027
rect 1144 2019 1152 2027
rect 1192 2019 1200 2027
rect 1512 2019 1520 2027
rect 1768 2019 1776 2027
rect 1880 2019 1888 2027
rect 2184 2019 2192 2027
rect 2216 2019 2224 2027
rect 3080 2019 3088 2027
rect 3480 2019 3488 2027
rect 3512 2019 3520 2027
rect 3768 2019 3776 2027
rect 4248 2019 4256 2027
rect 6146 2013 6154 2021
rect 6530 2013 6538 2021
rect 6562 2013 6570 2021
rect 7554 2013 7562 2021
rect 7842 2013 7850 2021
rect 8338 2013 8346 2021
rect 9122 2013 9130 2021
rect 9154 2013 9162 2021
rect 9330 2013 9338 2021
rect 10162 2013 10170 2021
rect 10306 2013 10314 2021
rect 10482 2013 10490 2021
rect 10802 2013 10810 2021
rect 12794 2019 12802 2027
rect 12810 2019 12818 2027
rect 13594 2019 13602 2027
rect 15178 2019 15186 2027
rect 16090 2019 16098 2027
rect 16970 2019 16978 2027
rect 22080 2020 22088 2028
rect 23136 2020 23144 2028
rect 31008 2017 31016 2025
rect 31728 2017 31736 2025
rect 32624 2017 32632 2025
rect 38864 2017 38872 2025
rect 728 1999 736 2007
rect 2152 1999 2160 2007
rect 2536 1999 2544 2007
rect 2568 1999 2576 2007
rect 2776 1999 2784 2007
rect 3864 1999 3872 2007
rect 4008 1999 4016 2007
rect 6642 1993 6650 2001
rect 6946 1993 6954 2001
rect 7074 1993 7082 2001
rect 8162 1993 8170 2001
rect 8194 1993 8202 2001
rect 8402 1993 8410 2001
rect 8466 1993 8474 2001
rect 8594 1993 8602 2001
rect 8770 1993 8778 2001
rect 9794 1993 9802 2001
rect 10274 1993 10282 2001
rect 12682 1999 12690 2007
rect 13194 1999 13202 2007
rect 13466 1999 13474 2007
rect 13706 1999 13714 2007
rect 14170 1999 14178 2007
rect 14426 1999 14434 2007
rect 16026 1999 16034 2007
rect 16266 1999 16274 2007
rect 16650 1999 16658 2007
rect 17114 1999 17122 2007
rect 17226 1999 17234 2007
rect 26624 2000 26632 2008
rect 32032 1997 32040 2005
rect 1320 1979 1328 1987
rect 1896 1979 1904 1987
rect 1976 1979 1984 1987
rect 3000 1979 3008 1987
rect 4136 1979 4144 1987
rect 7938 1973 7946 1981
rect 14666 1979 14674 1987
rect 14874 1979 14882 1987
rect 15370 1979 15378 1987
rect 16714 1979 16722 1987
rect 17034 1979 17042 1987
rect 25984 1980 25992 1988
rect 26416 1980 26424 1988
rect 29568 1977 29576 1985
rect 29632 1977 29640 1985
rect 30256 1977 30264 1985
rect 30528 1977 30536 1985
rect 30608 1977 30616 1985
rect 30688 1977 30696 1985
rect 30784 1977 30792 1985
rect 34704 1977 34712 1985
rect 34976 1977 34984 1985
rect 36320 1977 36328 1985
rect 36848 1977 36856 1985
rect 37168 1977 37176 1985
rect 37856 1977 37864 1985
rect 40128 1977 40136 1985
rect 952 1959 960 1967
rect 1128 1959 1136 1967
rect 1240 1959 1248 1967
rect 1288 1959 1296 1967
rect 2296 1959 2304 1967
rect 2824 1959 2832 1967
rect 2840 1959 2848 1967
rect 2872 1959 2880 1967
rect 2888 1959 2896 1967
rect 3720 1959 3728 1967
rect 3752 1959 3760 1967
rect 3960 1959 3968 1967
rect 4280 1959 4288 1967
rect 6274 1953 6282 1961
rect 6386 1953 6394 1961
rect 6402 1953 6410 1961
rect 6770 1953 6778 1961
rect 6882 1953 6890 1961
rect 6930 1953 6938 1961
rect 7522 1953 7530 1961
rect 7602 1953 7610 1961
rect 7762 1953 7770 1961
rect 8306 1953 8314 1961
rect 8434 1953 8442 1961
rect 8658 1953 8666 1961
rect 8690 1953 8698 1961
rect 9714 1953 9722 1961
rect 10338 1953 10346 1961
rect 10450 1953 10458 1961
rect 12426 1959 12434 1967
rect 12442 1959 12450 1967
rect 12474 1959 12482 1967
rect 12986 1959 12994 1967
rect 13274 1959 13282 1967
rect 13338 1959 13346 1967
rect 13834 1959 13842 1967
rect 14634 1959 14642 1967
rect 14666 1959 14674 1967
rect 14714 1959 14722 1967
rect 14858 1959 14866 1967
rect 15274 1959 15282 1967
rect 15562 1959 15570 1967
rect 15722 1959 15730 1967
rect 16186 1959 16194 1967
rect 16234 1959 16242 1967
rect 16282 1959 16290 1967
rect 16362 1959 16370 1967
rect 16410 1959 16418 1967
rect 16586 1959 16594 1967
rect 16826 1959 16834 1967
rect 17354 1959 17362 1967
rect 17450 1959 17458 1967
rect 18848 1960 18856 1968
rect 20128 1960 20136 1968
rect 20208 1960 20216 1968
rect 20416 1960 20424 1968
rect 20784 1961 20794 1966
rect 21696 1960 21704 1968
rect 21920 1960 21928 1968
rect 22272 1960 22280 1968
rect 22496 1960 22504 1968
rect 22768 1960 22776 1968
rect 22974 1961 22984 1966
rect 23184 1960 23192 1968
rect 23200 1960 23208 1968
rect 23616 1960 23624 1968
rect 23840 1960 23848 1968
rect 24048 1960 24056 1968
rect 24918 1961 24919 1966
rect 25920 1960 25928 1968
rect 27872 1960 27880 1968
rect 28320 1960 28328 1968
rect 31328 1957 31336 1965
rect 33824 1957 33832 1965
rect 34032 1957 34040 1965
rect 34880 1957 34888 1965
rect 34976 1957 34984 1965
rect 536 1939 544 1947
rect 552 1939 560 1947
rect 3672 1939 3680 1947
rect 5906 1933 5914 1941
rect 6370 1933 6378 1941
rect 6578 1933 6586 1941
rect 6642 1933 6650 1941
rect 6706 1933 6714 1941
rect 6754 1933 6762 1941
rect 6834 1933 6842 1941
rect 7218 1933 7226 1941
rect 7250 1933 7258 1941
rect 7330 1933 7338 1941
rect 7346 1933 7354 1941
rect 7442 1933 7450 1941
rect 7826 1933 7834 1941
rect 7906 1933 7914 1941
rect 8018 1933 8026 1941
rect 8226 1933 8234 1941
rect 8466 1933 8474 1941
rect 8482 1933 8490 1941
rect 8514 1933 8522 1941
rect 8674 1933 8682 1941
rect 8770 1933 8778 1941
rect 8898 1933 8906 1941
rect 8946 1933 8954 1941
rect 9202 1933 9210 1941
rect 9346 1933 9354 1941
rect 9362 1933 9370 1941
rect 10018 1933 10026 1941
rect 10690 1933 10698 1941
rect 12122 1939 12130 1947
rect 12922 1939 12930 1947
rect 12938 1939 12946 1947
rect 14602 1939 14610 1947
rect 15210 1939 15218 1947
rect 15498 1939 15506 1947
rect 15594 1939 15602 1947
rect 15818 1939 15826 1947
rect 16058 1939 16066 1947
rect 16474 1939 16482 1947
rect 16794 1939 16802 1947
rect 19296 1940 19304 1948
rect 19744 1940 19752 1948
rect 20048 1940 20056 1948
rect 20368 1940 20376 1948
rect 20576 1940 20584 1948
rect 21280 1940 21288 1948
rect 29376 1937 29384 1945
rect 29552 1937 29560 1945
rect 30400 1937 30408 1945
rect 30672 1937 30680 1945
rect 31184 1937 31192 1945
rect 31296 1937 31304 1945
rect 31376 1937 31384 1945
rect 31424 1937 31432 1945
rect 31616 1937 31624 1945
rect 31712 1937 31720 1945
rect 32032 1937 32040 1945
rect 32128 1937 32136 1945
rect 32240 1937 32248 1945
rect 32528 1937 32536 1945
rect 33088 1937 33096 1945
rect 33232 1937 33240 1945
rect 33808 1937 33816 1945
rect 34016 1937 34024 1945
rect 34272 1937 34280 1945
rect 34352 1937 34360 1945
rect 35056 1937 35064 1945
rect 35744 1937 35752 1945
rect 36032 1937 36040 1945
rect 36080 1937 36088 1945
rect 36672 1937 36680 1945
rect 36864 1937 36872 1945
rect 37072 1937 37080 1945
rect 38720 1937 38728 1945
rect 39024 1937 39032 1945
rect 39120 1937 39128 1945
rect 39280 1937 39288 1945
rect 39888 1937 39896 1945
rect 40368 1937 40376 1945
rect 424 1919 432 1927
rect 456 1919 464 1927
rect 920 1919 928 1927
rect 1352 1919 1360 1927
rect 1448 1919 1456 1927
rect 1576 1919 1584 1927
rect 1592 1919 1600 1927
rect 1608 1919 1616 1927
rect 1640 1919 1648 1927
rect 1720 1919 1728 1927
rect 1768 1919 1776 1927
rect 1800 1919 1808 1927
rect 2072 1919 2080 1927
rect 2232 1919 2240 1927
rect 2248 1919 2256 1927
rect 2312 1919 2320 1927
rect 2424 1919 2432 1927
rect 2904 1919 2912 1927
rect 3032 1919 3040 1927
rect 3048 1919 3056 1927
rect 3064 1919 3072 1927
rect 3416 1919 3424 1927
rect 3464 1919 3472 1927
rect 3928 1919 3936 1927
rect 3992 1919 4000 1927
rect 4568 1919 4576 1927
rect 4632 1919 4640 1927
rect 6066 1913 6074 1921
rect 6402 1913 6410 1921
rect 6706 1913 6714 1921
rect 8274 1913 8282 1921
rect 10546 1913 10554 1921
rect 12154 1919 12162 1927
rect 12186 1919 12194 1927
rect 12314 1919 12322 1927
rect 13658 1919 13666 1927
rect 14730 1919 14738 1927
rect 15834 1919 15842 1927
rect 16218 1919 16226 1927
rect 17386 1919 17394 1927
rect 18624 1920 18632 1928
rect 19264 1920 19272 1928
rect 21472 1920 21480 1928
rect 21504 1920 21512 1928
rect 21920 1920 21928 1928
rect 22096 1920 22104 1928
rect 22656 1920 22664 1928
rect 22880 1920 22888 1928
rect 24208 1920 24216 1928
rect 24496 1920 24504 1928
rect 24592 1920 24600 1928
rect 24704 1920 24712 1928
rect 25568 1920 25576 1928
rect 26112 1920 26120 1928
rect 26464 1920 26472 1928
rect 26608 1920 26616 1928
rect 26640 1920 26648 1928
rect 26960 1920 26968 1928
rect 27904 1920 27912 1928
rect 34832 1917 34840 1925
rect 35040 1917 35048 1925
rect 35152 1917 35160 1925
rect 35520 1917 35528 1925
rect 35568 1917 35576 1925
rect 35664 1917 35672 1925
rect 37312 1917 37320 1925
rect 37664 1917 37672 1925
rect 37728 1917 37736 1925
rect 38160 1917 38168 1925
rect 38256 1917 38264 1925
rect 38544 1917 38552 1925
rect 39104 1917 39112 1925
rect 39200 1917 39208 1925
rect 39312 1917 39320 1925
rect 39552 1917 39560 1925
rect 440 1899 448 1907
rect 600 1899 608 1907
rect 744 1899 752 1907
rect 776 1899 784 1907
rect 856 1899 864 1907
rect 968 1899 976 1907
rect 1160 1899 1168 1907
rect 1176 1899 1184 1907
rect 1304 1899 1312 1907
rect 1432 1899 1440 1907
rect 1528 1899 1536 1907
rect 1704 1899 1712 1907
rect 1784 1899 1792 1907
rect 1864 1899 1872 1907
rect 1896 1899 1904 1907
rect 2008 1899 2016 1907
rect 2088 1899 2096 1907
rect 2168 1899 2176 1907
rect 2200 1899 2208 1907
rect 2232 1899 2240 1907
rect 2456 1899 2464 1907
rect 2520 1899 2528 1907
rect 2552 1899 2560 1907
rect 2840 1899 2848 1907
rect 3048 1899 3056 1907
rect 3096 1899 3104 1907
rect 3176 1899 3184 1907
rect 3192 1899 3200 1907
rect 3336 1899 3344 1907
rect 3368 1899 3376 1907
rect 3448 1899 3456 1907
rect 3496 1899 3504 1907
rect 3528 1899 3536 1907
rect 3704 1899 3712 1907
rect 3720 1899 3728 1907
rect 3784 1899 3792 1907
rect 3816 1899 3824 1907
rect 4024 1899 4032 1907
rect 4056 1899 4064 1907
rect 4184 1899 4192 1907
rect 4392 1899 4400 1907
rect 4456 1899 4464 1907
rect 4536 1899 4544 1907
rect 4568 1899 4576 1907
rect 5794 1893 5802 1901
rect 6018 1893 6026 1901
rect 6034 1893 6042 1901
rect 6162 1893 6170 1901
rect 6418 1893 6426 1901
rect 6514 1893 6522 1901
rect 6562 1893 6570 1901
rect 6610 1893 6618 1901
rect 6626 1893 6634 1901
rect 6962 1893 6970 1901
rect 7090 1893 7098 1901
rect 7266 1893 7274 1901
rect 7346 1893 7354 1901
rect 7570 1893 7578 1901
rect 7650 1893 7658 1901
rect 7826 1893 7834 1901
rect 7858 1893 7866 1901
rect 7938 1893 7946 1901
rect 8322 1893 8330 1901
rect 9058 1893 9066 1901
rect 9394 1893 9402 1901
rect 9554 1893 9562 1901
rect 10034 1893 10042 1901
rect 10082 1893 10090 1901
rect 10258 1893 10266 1901
rect 10290 1893 10298 1901
rect 10658 1893 10666 1901
rect 10706 1893 10714 1901
rect 12378 1899 12386 1907
rect 12890 1899 12898 1907
rect 13210 1899 13218 1907
rect 13306 1899 13314 1907
rect 13578 1899 13586 1907
rect 13722 1899 13730 1907
rect 13978 1899 13986 1907
rect 14218 1899 14226 1907
rect 14522 1899 14530 1907
rect 15066 1899 15074 1907
rect 16666 1899 16674 1907
rect 23424 1900 23432 1908
rect 24304 1900 24312 1908
rect 25328 1900 25336 1908
rect 28352 1900 28360 1908
rect 30288 1897 30296 1905
rect 31600 1897 31608 1905
rect 31616 1897 31624 1905
rect 31920 1897 31928 1905
rect 32064 1897 32072 1905
rect 32496 1897 32504 1905
rect 35984 1897 35992 1905
rect 36352 1897 36360 1905
rect 37040 1897 37048 1905
rect 37472 1897 37480 1905
rect 37760 1897 37768 1905
rect 38528 1897 38536 1905
rect 40208 1897 40216 1905
rect 792 1879 800 1887
rect 1128 1879 1136 1887
rect 1656 1879 1664 1887
rect 1816 1879 1824 1887
rect 1864 1879 1872 1887
rect 1912 1879 1920 1887
rect 2552 1879 2560 1887
rect 2568 1879 2576 1887
rect 2632 1879 2640 1887
rect 2712 1879 2720 1887
rect 3144 1879 3152 1887
rect 3800 1879 3808 1887
rect 4072 1879 4080 1887
rect 4248 1879 4256 1887
rect 5778 1873 5786 1881
rect 6818 1873 6826 1881
rect 7266 1873 7274 1881
rect 7810 1873 7818 1881
rect 8978 1873 8986 1881
rect 9074 1873 9082 1881
rect 9186 1873 9194 1881
rect 9234 1873 9242 1881
rect 12698 1879 12706 1887
rect 13018 1879 13026 1887
rect 13130 1879 13138 1887
rect 13146 1879 13154 1887
rect 14442 1879 14450 1887
rect 15626 1879 15634 1887
rect 15754 1879 15762 1887
rect 16074 1879 16082 1887
rect 19312 1880 19320 1888
rect 19952 1880 19960 1888
rect 27616 1880 27624 1888
rect 31248 1877 31256 1885
rect 38800 1877 38808 1885
rect 1192 1859 1200 1867
rect 2104 1859 2112 1867
rect 2872 1859 2880 1867
rect 7090 1853 7098 1861
rect 7202 1853 7210 1861
rect 7218 1853 7226 1861
rect 7650 1853 7658 1861
rect 7714 1853 7722 1861
rect 7858 1853 7866 1861
rect 8418 1853 8426 1861
rect 8450 1853 8458 1861
rect 8738 1853 8746 1861
rect 15386 1859 15394 1867
rect 16858 1859 16866 1867
rect 22736 1860 22744 1868
rect 29428 1867 29440 1875
rect 29444 1867 29448 1875
rect 29460 1867 29472 1875
rect 29488 1867 29504 1875
rect 29512 1867 29544 1875
rect 29552 1867 29564 1875
rect 29584 1867 29596 1875
rect 29604 1867 29636 1875
rect 29644 1867 29660 1875
rect 29676 1867 29688 1875
rect 29696 1867 29728 1875
rect 29736 1867 29752 1875
rect 29768 1867 29784 1875
rect 29800 1867 29804 1875
rect 29808 1867 29820 1875
rect 29832 1867 29836 1875
rect 29840 1867 29844 1875
rect 29856 1867 29868 1875
rect 29872 1867 29876 1875
rect 29896 1867 29900 1875
rect 29904 1867 29908 1875
rect 29920 1867 29932 1875
rect 29936 1867 29940 1875
rect 29960 1867 29964 1875
rect 29968 1867 29980 1875
rect 29984 1867 29996 1875
rect 30000 1867 30004 1875
rect 30020 1867 30044 1875
rect 30052 1867 30068 1875
rect 30076 1867 30100 1875
rect 30116 1867 30128 1875
rect 30148 1867 30160 1875
rect 30172 1867 30176 1875
rect 30180 1867 30192 1875
rect 30196 1867 30200 1875
rect 30212 1867 30224 1875
rect 30240 1867 30252 1875
rect 30264 1867 30268 1875
rect 30272 1867 30284 1875
rect 30288 1867 30292 1875
rect 30332 1867 30344 1875
rect 30356 1867 30360 1875
rect 30364 1867 30376 1875
rect 30380 1867 30384 1875
rect 30400 1867 30408 1875
rect 30448 1867 30452 1875
rect 30456 1867 30468 1875
rect 30472 1867 30476 1875
rect 30488 1867 30500 1875
rect 30516 1867 30532 1875
rect 30548 1867 30572 1875
rect 30580 1867 30596 1875
rect 30604 1867 30628 1875
rect 30644 1867 30648 1875
rect 30652 1867 30664 1875
rect 30668 1867 30680 1875
rect 30684 1867 30688 1875
rect 30708 1867 30712 1875
rect 30716 1867 30720 1875
rect 30816 1867 30820 1875
rect 30824 1867 30836 1875
rect 30840 1867 30852 1875
rect 30856 1867 30860 1875
rect 30956 1867 30960 1875
rect 30964 1867 30968 1875
rect 30988 1867 30992 1875
rect 30996 1867 31008 1875
rect 31012 1867 31024 1875
rect 31028 1867 31032 1875
rect 31052 1867 31056 1875
rect 31060 1867 31064 1875
rect 31272 1867 31276 1875
rect 31280 1867 31284 1875
rect 31296 1867 31308 1875
rect 31312 1867 31316 1875
rect 31332 1867 31336 1875
rect 31340 1867 31352 1875
rect 31364 1867 31368 1875
rect 31372 1867 31376 1875
rect 31388 1867 31400 1875
rect 31404 1867 31408 1875
rect 31428 1867 31432 1875
rect 31436 1867 31440 1875
rect 31456 1867 31472 1875
rect 31480 1867 31512 1875
rect 31528 1867 31544 1875
rect 31560 1867 31564 1875
rect 31568 1867 31580 1875
rect 31592 1867 31596 1875
rect 31600 1867 31604 1875
rect 31624 1867 31628 1875
rect 31632 1867 31636 1875
rect 31668 1867 31672 1875
rect 31676 1867 31688 1875
rect 31708 1867 31720 1875
rect 31724 1867 31736 1875
rect 31752 1867 31764 1875
rect 31784 1867 31796 1875
rect 31800 1867 31812 1875
rect 31816 1867 31828 1875
rect 31848 1867 31860 1875
rect 31872 1867 31876 1875
rect 31880 1867 31884 1875
rect 31904 1867 31908 1875
rect 31912 1867 31916 1875
rect 31964 1867 31968 1875
rect 31972 1867 31984 1875
rect 32088 1867 32092 1875
rect 32096 1867 32108 1875
rect 32128 1867 32140 1875
rect 32144 1867 32148 1875
rect 32180 1867 32184 1875
rect 32188 1867 32200 1875
rect 32220 1867 32232 1875
rect 32236 1867 32240 1875
rect 32252 1867 32264 1875
rect 32284 1867 32296 1875
rect 32312 1867 32360 1875
rect 32376 1867 32388 1875
rect 32404 1867 32452 1875
rect 32468 1867 32484 1875
rect 32500 1867 32504 1875
rect 32508 1867 32520 1875
rect 32532 1867 32536 1875
rect 32540 1867 32544 1875
rect 32564 1867 32568 1875
rect 32572 1867 32576 1875
rect 32672 1867 32676 1875
rect 32680 1867 32684 1875
rect 32696 1867 32708 1875
rect 32712 1867 32716 1875
rect 32732 1867 32756 1875
rect 32764 1867 32780 1875
rect 32788 1867 32820 1875
rect 32828 1867 32844 1875
rect 32860 1867 32872 1875
rect 32880 1867 32912 1875
rect 32920 1867 32936 1875
rect 32952 1867 32964 1875
rect 32976 1867 32980 1875
rect 32984 1867 32996 1875
rect 33016 1867 33028 1875
rect 33132 1867 33136 1875
rect 33140 1867 33152 1875
rect 33156 1867 33160 1875
rect 33172 1867 33184 1875
rect 33200 1867 33216 1875
rect 33232 1867 33256 1875
rect 33264 1867 33280 1875
rect 33288 1867 33312 1875
rect 33328 1867 33332 1875
rect 33336 1867 33348 1875
rect 33352 1867 33364 1875
rect 33368 1867 33372 1875
rect 33392 1867 33396 1875
rect 33400 1867 33404 1875
rect 33468 1867 33472 1875
rect 33476 1867 33480 1875
rect 33500 1867 33504 1875
rect 33508 1867 33520 1875
rect 33524 1867 33536 1875
rect 33540 1867 33544 1875
rect 33564 1867 33568 1875
rect 33572 1867 33584 1875
rect 33588 1867 33600 1875
rect 33604 1867 33608 1875
rect 33628 1867 33632 1875
rect 33636 1867 33648 1875
rect 33652 1867 33664 1875
rect 33668 1867 33672 1875
rect 33720 1867 33724 1875
rect 33728 1867 33740 1875
rect 33744 1867 33756 1875
rect 33760 1867 33764 1875
rect 33784 1867 33788 1875
rect 33792 1867 33796 1875
rect 33860 1867 33864 1875
rect 33868 1867 33872 1875
rect 33892 1867 33896 1875
rect 33900 1867 33912 1875
rect 33916 1867 33928 1875
rect 33932 1867 33936 1875
rect 33956 1867 33960 1875
rect 33964 1867 33976 1875
rect 33984 1867 34000 1875
rect 34008 1867 34032 1875
rect 34048 1867 34064 1875
rect 34080 1867 34092 1875
rect 34104 1867 34108 1875
rect 34112 1867 34124 1875
rect 34128 1867 34132 1875
rect 34236 1867 34248 1875
rect 34328 1867 34340 1875
rect 34360 1867 34372 1875
rect 34376 1867 34380 1875
rect 34392 1867 34400 1875
rect 34420 1867 34436 1875
rect 34444 1867 34476 1875
rect 34484 1867 34500 1875
rect 34516 1867 34528 1875
rect 34536 1867 34568 1875
rect 34576 1867 34592 1875
rect 34608 1867 34620 1875
rect 34632 1867 34636 1875
rect 34640 1867 34652 1875
rect 34672 1867 34684 1875
rect 34860 1867 34872 1875
rect 34876 1867 34880 1875
rect 34892 1867 34904 1875
rect 34920 1867 34936 1875
rect 34944 1867 34976 1875
rect 34984 1867 35000 1875
rect 35016 1867 35028 1875
rect 35036 1867 35068 1875
rect 35076 1867 35092 1875
rect 35108 1867 35120 1875
rect 35128 1867 35160 1875
rect 35168 1867 35184 1875
rect 35200 1867 35216 1875
rect 35232 1867 35236 1875
rect 35240 1867 35252 1875
rect 35264 1867 35268 1875
rect 35272 1867 35276 1875
rect 35532 1867 35536 1875
rect 35540 1867 35544 1875
rect 35564 1867 35568 1875
rect 35572 1867 35584 1875
rect 35588 1867 35600 1875
rect 35604 1867 35608 1875
rect 35656 1867 35660 1875
rect 35664 1867 35676 1875
rect 35680 1867 35692 1875
rect 35696 1867 35700 1875
rect 35748 1867 35752 1875
rect 35756 1867 35768 1875
rect 35772 1867 35784 1875
rect 35788 1867 35792 1875
rect 35812 1867 35816 1875
rect 35820 1867 35824 1875
rect 35836 1867 35848 1875
rect 35852 1867 35856 1875
rect 35876 1867 35880 1875
rect 35884 1867 35888 1875
rect 35900 1867 35912 1875
rect 35916 1867 35928 1875
rect 35940 1867 35944 1875
rect 35948 1867 35952 1875
rect 35968 1867 35984 1875
rect 35992 1867 36004 1875
rect 36008 1867 36020 1875
rect 36032 1867 36036 1875
rect 36040 1867 36044 1875
rect 36060 1867 36076 1875
rect 36084 1867 36096 1875
rect 36100 1867 36112 1875
rect 36124 1867 36128 1875
rect 36132 1867 36136 1875
rect 36152 1867 36168 1875
rect 36176 1867 36200 1875
rect 36216 1867 36232 1875
rect 36240 1867 36272 1875
rect 36280 1867 36296 1875
rect 36312 1867 36316 1875
rect 36320 1867 36324 1875
rect 36344 1867 36348 1875
rect 36352 1867 36364 1875
rect 36376 1867 36380 1875
rect 36384 1867 36388 1875
rect 36468 1867 36472 1875
rect 36476 1867 36480 1875
rect 36492 1867 36504 1875
rect 36508 1867 36520 1875
rect 36532 1867 36536 1875
rect 36540 1867 36544 1875
rect 36560 1867 36564 1875
rect 36568 1867 36572 1875
rect 36584 1867 36596 1875
rect 36600 1867 36612 1875
rect 36624 1867 36628 1875
rect 36632 1867 36636 1875
rect 36732 1867 36736 1875
rect 36740 1867 36752 1875
rect 36764 1867 36768 1875
rect 36772 1867 36776 1875
rect 36788 1867 36800 1875
rect 36804 1867 36808 1875
rect 36824 1867 36828 1875
rect 36832 1867 36844 1875
rect 36856 1867 36860 1875
rect 36864 1867 36868 1875
rect 36880 1867 36892 1875
rect 36896 1867 36900 1875
rect 36948 1867 36952 1875
rect 36956 1867 36960 1875
rect 36972 1867 36984 1875
rect 36988 1867 36992 1875
rect 37088 1867 37092 1875
rect 37096 1867 37100 1875
rect 37112 1867 37124 1875
rect 37128 1867 37140 1875
rect 37152 1867 37156 1875
rect 37160 1867 37164 1875
rect 37184 1867 37188 1875
rect 37192 1867 37196 1875
rect 37340 1867 37344 1875
rect 37348 1867 37360 1875
rect 37364 1867 37376 1875
rect 37380 1867 37384 1875
rect 37404 1867 37408 1875
rect 37412 1867 37424 1875
rect 37432 1867 37448 1875
rect 37456 1867 37480 1875
rect 37496 1867 37512 1875
rect 37528 1867 37540 1875
rect 37552 1867 37556 1875
rect 37560 1867 37572 1875
rect 37576 1867 37580 1875
rect 37592 1867 37600 1875
rect 37616 1867 37620 1875
rect 37624 1867 37636 1875
rect 37640 1867 37644 1875
rect 37656 1867 37668 1875
rect 37748 1867 37760 1875
rect 37780 1867 37792 1875
rect 37796 1867 37808 1875
rect 37812 1867 37824 1875
rect 37968 1867 37980 1875
rect 37984 1867 37988 1875
rect 38000 1867 38012 1875
rect 38020 1867 38044 1875
rect 38060 1867 38072 1875
rect 38076 1867 38080 1875
rect 38092 1867 38104 1875
rect 38112 1867 38136 1875
rect 38152 1867 38176 1875
rect 38184 1867 38196 1875
rect 38208 1867 38212 1875
rect 38216 1867 38228 1875
rect 38372 1867 38384 1875
rect 38388 1867 38392 1875
rect 38404 1867 38416 1875
rect 38436 1867 38448 1875
rect 38464 1867 38512 1875
rect 38528 1867 38576 1875
rect 38592 1867 38604 1875
rect 38624 1867 38636 1875
rect 38648 1867 38652 1875
rect 38656 1867 38668 1875
rect 38740 1867 38744 1875
rect 38748 1867 38760 1875
rect 38780 1867 38792 1875
rect 38796 1867 38800 1875
rect 38872 1867 38884 1875
rect 38888 1867 38892 1875
rect 38964 1867 38976 1875
rect 38996 1867 39008 1875
rect 39012 1867 39016 1875
rect 39028 1867 39040 1875
rect 39052 1867 39056 1875
rect 39060 1867 39072 1875
rect 39088 1867 39136 1875
rect 39152 1867 39168 1875
rect 39176 1867 39188 1875
rect 39192 1867 39200 1875
rect 39216 1867 39220 1875
rect 39224 1867 39228 1875
rect 39240 1867 39252 1875
rect 39256 1867 39260 1875
rect 39404 1867 39408 1875
rect 39412 1867 39416 1875
rect 39436 1867 39440 1875
rect 39444 1867 39456 1875
rect 39460 1867 39472 1875
rect 39476 1867 39480 1875
rect 39500 1867 39504 1875
rect 39508 1867 39520 1875
rect 39528 1867 39544 1875
rect 39552 1867 39576 1875
rect 39592 1867 39604 1875
rect 39624 1867 39636 1875
rect 39648 1867 39652 1875
rect 39656 1867 39668 1875
rect 39672 1867 39676 1875
rect 39688 1867 39700 1875
rect 39780 1867 39792 1875
rect 39904 1867 39916 1875
rect 39920 1867 39924 1875
rect 39936 1867 39948 1875
rect 39968 1867 39980 1875
rect 39988 1867 40020 1875
rect 40028 1867 40044 1875
rect 40052 1867 40076 1875
rect 40092 1867 40108 1875
rect 40124 1867 40136 1875
rect 40148 1867 40152 1875
rect 40156 1867 40168 1875
rect 40172 1867 40176 1875
rect 40188 1867 40200 1875
rect 40212 1867 40216 1875
rect 40220 1867 40232 1875
rect 40248 1867 40260 1875
rect 40264 1867 40268 1875
rect 40280 1867 40292 1875
rect 40300 1867 40324 1875
rect 40340 1867 40352 1875
rect 40356 1867 40360 1875
rect 40372 1867 40384 1875
rect 40392 1867 40416 1875
rect 40432 1867 40480 1875
rect 40496 1867 40544 1875
rect 40560 1867 40576 1875
rect 40592 1867 40604 1875
rect 40616 1867 40620 1875
rect 40624 1867 40636 1875
rect 19152 1850 19156 1858
rect 19242 1850 19250 1858
rect 19366 1850 19370 1858
rect 19456 1850 19464 1858
rect 21524 1850 21530 1858
rect 21532 1850 21538 1858
rect 21730 1850 21744 1858
rect 21944 1850 21958 1858
rect 22586 1850 22600 1858
rect 23014 1850 23028 1858
rect 23228 1850 23242 1858
rect 23658 1856 23662 1858
rect 23736 1850 23750 1858
rect 23790 1850 23804 1858
rect 23970 1850 23982 1858
rect 24304 1850 24310 1858
rect 24518 1850 24524 1858
rect 24612 1850 24624 1858
rect 24946 1850 24952 1858
rect 25040 1850 25052 1858
rect 25262 1850 25264 1858
rect 25354 1850 25364 1858
rect 25456 1850 25458 1858
rect 25690 1850 25692 1858
rect 25782 1850 25792 1858
rect 25884 1850 25886 1858
rect 26098 1850 26100 1858
rect 26332 1850 26334 1858
rect 26538 1850 26540 1858
rect 26752 1850 26754 1858
rect 26834 1850 26842 1858
rect 26922 1850 26928 1858
rect 26930 1850 26936 1858
rect 26976 1850 26982 1858
rect 26984 1850 26990 1858
rect 27136 1850 27142 1858
rect 27144 1850 27150 1858
rect 27190 1850 27196 1858
rect 27198 1850 27204 1858
rect 27284 1850 27290 1858
rect 27498 1850 27504 1858
rect 27712 1850 27718 1858
rect 27806 1850 27808 1858
rect 28028 1850 28030 1858
rect 28242 1850 28244 1858
rect 28456 1850 28458 1858
rect 32672 1857 32680 1865
rect 33440 1857 33448 1865
rect 696 1839 704 1847
rect 2088 1839 2096 1847
rect 2792 1839 2800 1847
rect 3800 1839 3808 1847
rect 6466 1833 6474 1841
rect 6754 1833 6762 1841
rect 8322 1833 8330 1841
rect 8690 1833 8698 1841
rect 9042 1833 9050 1841
rect 9058 1833 9066 1841
rect 10066 1833 10074 1841
rect 14538 1839 14546 1847
rect 16602 1839 16610 1847
rect 22256 1840 22264 1848
rect 23408 1840 23416 1848
rect 29456 1837 29464 1845
rect 30080 1837 30088 1845
rect 30736 1837 30744 1845
rect 31056 1837 31064 1845
rect 31136 1837 31144 1845
rect 31296 1837 31304 1845
rect 32240 1837 32248 1845
rect 32624 1837 32632 1845
rect 33536 1837 33544 1845
rect 34816 1837 34824 1845
rect 35616 1837 35624 1845
rect 35840 1837 35848 1845
rect 37600 1837 37608 1845
rect 424 1819 432 1827
rect 1352 1819 1360 1827
rect 1768 1819 1776 1827
rect 1832 1819 1840 1827
rect 2152 1819 2160 1827
rect 2328 1819 2336 1827
rect 2856 1819 2864 1827
rect 3464 1819 3472 1827
rect 3512 1819 3520 1827
rect 3720 1819 3728 1827
rect 4024 1819 4032 1827
rect 5938 1813 5946 1821
rect 6242 1813 6250 1821
rect 6610 1813 6618 1821
rect 6642 1813 6650 1821
rect 6722 1813 6730 1821
rect 7362 1813 7370 1821
rect 8098 1813 8106 1821
rect 8114 1813 8122 1821
rect 8642 1813 8650 1821
rect 8722 1813 8730 1821
rect 8802 1813 8810 1821
rect 9218 1813 9226 1821
rect 9474 1813 9482 1821
rect 10210 1813 10218 1821
rect 10402 1813 10410 1821
rect 10818 1813 10826 1821
rect 12122 1819 12130 1827
rect 12298 1819 12306 1827
rect 12826 1819 12834 1827
rect 12874 1819 12882 1827
rect 12890 1819 12898 1827
rect 12954 1819 12962 1827
rect 13306 1819 13314 1827
rect 13530 1819 13538 1827
rect 13834 1819 13842 1827
rect 13866 1819 13874 1827
rect 14474 1819 14482 1827
rect 14506 1819 14514 1827
rect 14554 1819 14562 1827
rect 14730 1819 14738 1827
rect 14858 1819 14866 1827
rect 14938 1819 14946 1827
rect 15306 1819 15314 1827
rect 16074 1819 16082 1827
rect 18672 1820 18680 1828
rect 19520 1820 19528 1828
rect 22016 1820 22024 1828
rect 23920 1820 23928 1828
rect 24336 1820 24344 1828
rect 25760 1820 25768 1828
rect 26480 1820 26488 1828
rect 30240 1817 30248 1825
rect 30784 1817 30792 1825
rect 31136 1817 31144 1825
rect 32672 1817 32680 1825
rect 32736 1817 32744 1825
rect 33072 1817 33080 1825
rect 33104 1817 33112 1825
rect 34400 1817 34408 1825
rect 36832 1817 36840 1825
rect 36912 1817 36920 1825
rect 36928 1817 36936 1825
rect 37152 1817 37160 1825
rect 37280 1817 37288 1825
rect 37600 1817 37608 1825
rect 37856 1817 37864 1825
rect 38832 1817 38840 1825
rect 38864 1817 38872 1825
rect 38896 1817 38904 1825
rect 39024 1817 39032 1825
rect 39264 1817 39272 1825
rect 39344 1817 39352 1825
rect 40288 1817 40296 1825
rect 40720 1817 40728 1825
rect 40768 1817 40776 1825
rect 552 1799 560 1807
rect 648 1799 656 1807
rect 680 1799 688 1807
rect 712 1799 720 1807
rect 728 1799 736 1807
rect 744 1799 752 1807
rect 824 1799 832 1807
rect 840 1799 848 1807
rect 920 1799 928 1807
rect 1000 1799 1008 1807
rect 1112 1799 1120 1807
rect 1192 1799 1200 1807
rect 1208 1799 1216 1807
rect 1240 1799 1248 1807
rect 1272 1799 1280 1807
rect 1368 1799 1376 1807
rect 1384 1799 1392 1807
rect 1464 1799 1472 1807
rect 1496 1799 1504 1807
rect 1512 1799 1520 1807
rect 1576 1799 1584 1807
rect 1592 1799 1600 1807
rect 1608 1799 1616 1807
rect 1688 1799 1696 1807
rect 1704 1799 1712 1807
rect 1752 1799 1760 1807
rect 2040 1799 2048 1807
rect 2264 1799 2272 1807
rect 2296 1799 2304 1807
rect 2360 1799 2368 1807
rect 2712 1799 2720 1807
rect 2728 1799 2736 1807
rect 2760 1799 2768 1807
rect 2840 1799 2848 1807
rect 2872 1799 2880 1807
rect 2936 1799 2944 1807
rect 2968 1799 2976 1807
rect 3128 1799 3136 1807
rect 3208 1799 3216 1807
rect 3272 1799 3280 1807
rect 3432 1799 3440 1807
rect 3480 1799 3488 1807
rect 3544 1799 3552 1807
rect 3736 1799 3744 1807
rect 3800 1799 3808 1807
rect 3896 1799 3904 1807
rect 3912 1799 3920 1807
rect 3992 1799 4000 1807
rect 4040 1799 4048 1807
rect 4056 1799 4064 1807
rect 4088 1799 4096 1807
rect 4184 1799 4192 1807
rect 4280 1799 4288 1807
rect 4296 1799 4304 1807
rect 4392 1799 4400 1807
rect 4424 1799 4432 1807
rect 4456 1799 4464 1807
rect 4536 1799 4544 1807
rect 4584 1799 4592 1807
rect 5858 1793 5866 1801
rect 5890 1793 5898 1801
rect 5922 1793 5930 1801
rect 6562 1793 6570 1801
rect 7394 1793 7402 1801
rect 7410 1793 7418 1801
rect 7458 1793 7466 1801
rect 7474 1793 7482 1801
rect 7602 1793 7610 1801
rect 7682 1793 7690 1801
rect 7858 1793 7866 1801
rect 7874 1793 7882 1801
rect 7890 1793 7898 1801
rect 7906 1793 7914 1801
rect 8002 1793 8010 1801
rect 8578 1793 8586 1801
rect 8658 1793 8666 1801
rect 8946 1793 8954 1801
rect 9170 1793 9178 1801
rect 9202 1793 9210 1801
rect 9298 1793 9306 1801
rect 9346 1793 9354 1801
rect 9794 1793 9802 1801
rect 9842 1793 9850 1801
rect 10738 1793 10746 1801
rect 10834 1793 10842 1801
rect 12650 1799 12658 1807
rect 14074 1799 14082 1807
rect 16586 1799 16594 1807
rect 17034 1799 17042 1807
rect 17482 1799 17490 1807
rect 18896 1800 18904 1808
rect 22464 1800 22472 1808
rect 22880 1800 22888 1808
rect 23248 1800 23256 1808
rect 24544 1800 24552 1808
rect 25408 1800 25416 1808
rect 26656 1800 26664 1808
rect 27600 1800 27608 1808
rect 30064 1797 30072 1805
rect 30144 1797 30152 1805
rect 30336 1797 30344 1805
rect 30896 1797 30904 1805
rect 31504 1797 31512 1805
rect 31520 1797 31528 1805
rect 31552 1797 31560 1805
rect 31728 1797 31736 1805
rect 31872 1797 31880 1805
rect 32096 1797 32104 1805
rect 32480 1797 32488 1805
rect 34352 1797 34360 1805
rect 34560 1797 34568 1805
rect 34640 1797 34648 1805
rect 35264 1797 35272 1805
rect 36176 1797 36184 1805
rect 36320 1797 36328 1805
rect 36832 1797 36840 1805
rect 36944 1797 36952 1805
rect 37024 1797 37032 1805
rect 37376 1797 37384 1805
rect 37600 1797 37608 1805
rect 38320 1797 38328 1805
rect 38480 1797 38488 1805
rect 38672 1797 38680 1805
rect 40432 1797 40440 1805
rect 648 1779 656 1787
rect 904 1779 912 1787
rect 2008 1779 2016 1787
rect 2024 1779 2032 1787
rect 2264 1779 2272 1787
rect 2312 1779 2320 1787
rect 2616 1779 2624 1787
rect 3000 1779 3008 1787
rect 3160 1779 3168 1787
rect 3576 1779 3584 1787
rect 4392 1779 4400 1787
rect 4440 1779 4448 1787
rect 5970 1773 5978 1781
rect 6210 1773 6218 1781
rect 7218 1773 7226 1781
rect 7458 1773 7466 1781
rect 7474 1773 7482 1781
rect 7586 1773 7594 1781
rect 7634 1773 7642 1781
rect 7746 1773 7754 1781
rect 7810 1773 7818 1781
rect 7826 1773 7834 1781
rect 8306 1773 8314 1781
rect 8786 1773 8794 1781
rect 8898 1773 8906 1781
rect 9378 1773 9386 1781
rect 9554 1773 9562 1781
rect 9698 1773 9706 1781
rect 9746 1773 9754 1781
rect 9778 1773 9786 1781
rect 9890 1773 9898 1781
rect 10178 1773 10186 1781
rect 10386 1773 10394 1781
rect 10418 1773 10426 1781
rect 10738 1773 10746 1781
rect 12106 1779 12114 1787
rect 12506 1779 12514 1787
rect 13386 1779 13394 1787
rect 13930 1779 13938 1787
rect 14746 1779 14754 1787
rect 15066 1779 15074 1787
rect 15258 1779 15266 1787
rect 15658 1779 15666 1787
rect 16138 1779 16146 1787
rect 17130 1779 17138 1787
rect 19888 1780 19896 1788
rect 21360 1780 21368 1788
rect 21872 1780 21880 1788
rect 21968 1780 21976 1788
rect 22400 1780 22408 1788
rect 23568 1780 23576 1788
rect 23744 1780 23752 1788
rect 23776 1780 23784 1788
rect 24208 1780 24216 1788
rect 24736 1780 24744 1788
rect 25552 1780 25560 1788
rect 25664 1780 25672 1788
rect 26000 1780 26008 1788
rect 26208 1780 26216 1788
rect 26640 1780 26648 1788
rect 26784 1780 26792 1788
rect 26960 1780 26968 1788
rect 27808 1780 27816 1788
rect 28432 1780 28440 1788
rect 29776 1777 29784 1785
rect 30752 1777 30760 1785
rect 31088 1777 31096 1785
rect 32672 1777 32680 1785
rect 33136 1777 33144 1785
rect 33648 1777 33656 1785
rect 34208 1777 34216 1785
rect 34368 1777 34376 1785
rect 35616 1777 35624 1785
rect 36176 1777 36184 1785
rect 36496 1777 36504 1785
rect 40560 1777 40568 1785
rect 1336 1759 1344 1767
rect 2072 1759 2080 1767
rect 2568 1759 2576 1767
rect 3656 1759 3664 1767
rect 4264 1759 4272 1767
rect 5778 1753 5786 1761
rect 6386 1753 6394 1761
rect 6514 1753 6522 1761
rect 7074 1753 7082 1761
rect 7714 1753 7722 1761
rect 8258 1753 8266 1761
rect 8306 1753 8314 1761
rect 8402 1753 8410 1761
rect 8722 1753 8730 1761
rect 8882 1753 8890 1761
rect 9410 1753 9418 1761
rect 9458 1753 9466 1761
rect 10066 1753 10074 1761
rect 10370 1753 10378 1761
rect 10786 1753 10794 1761
rect 10802 1753 10810 1761
rect 12186 1759 12194 1767
rect 12554 1759 12562 1767
rect 12634 1759 12642 1767
rect 12746 1759 12754 1767
rect 13706 1759 13714 1767
rect 14106 1759 14114 1767
rect 14282 1759 14290 1767
rect 14986 1759 14994 1767
rect 15114 1759 15122 1767
rect 20928 1760 20936 1768
rect 21504 1760 21512 1768
rect 21760 1760 21768 1768
rect 27984 1760 27992 1768
rect 28224 1760 28232 1768
rect 30208 1757 30216 1765
rect 30320 1757 30328 1765
rect 32848 1757 32856 1765
rect 33600 1757 33608 1765
rect 33872 1757 33880 1765
rect 34256 1757 34264 1765
rect 34672 1757 34680 1765
rect 35008 1757 35016 1765
rect 35296 1757 35304 1765
rect 35632 1757 35640 1765
rect 35696 1757 35704 1765
rect 36000 1757 36008 1765
rect 36496 1757 36504 1765
rect 37056 1757 37064 1765
rect 37648 1757 37656 1765
rect 37760 1757 37768 1765
rect 38832 1757 38840 1765
rect 39216 1757 39224 1765
rect 39312 1757 39320 1765
rect 39616 1757 39624 1765
rect 39776 1757 39784 1765
rect 40032 1757 40040 1765
rect 40608 1757 40616 1765
rect 19112 1748 19116 1753
rect 23058 1748 23062 1753
rect 1624 1739 1632 1747
rect 2184 1739 2192 1747
rect 2584 1739 2592 1747
rect 2664 1739 2672 1747
rect 3032 1739 3040 1747
rect 3448 1739 3456 1747
rect 3528 1739 3536 1747
rect 4088 1739 4096 1747
rect 4120 1739 4128 1747
rect 4488 1739 4496 1747
rect 6002 1733 6010 1741
rect 6290 1733 6298 1741
rect 6418 1733 6426 1741
rect 6562 1733 6570 1741
rect 6834 1733 6842 1741
rect 6882 1733 6890 1741
rect 6946 1733 6954 1741
rect 7154 1733 7162 1741
rect 7506 1733 7514 1741
rect 7554 1733 7562 1741
rect 8098 1733 8106 1741
rect 8706 1733 8714 1741
rect 8738 1733 8746 1741
rect 8770 1733 8778 1741
rect 8930 1733 8938 1741
rect 8946 1733 8954 1741
rect 9042 1733 9050 1741
rect 9154 1733 9162 1741
rect 9634 1733 9642 1741
rect 9698 1733 9706 1741
rect 9938 1733 9946 1741
rect 10210 1733 10218 1741
rect 10738 1733 10746 1741
rect 10882 1733 10890 1741
rect 12362 1739 12370 1747
rect 12522 1739 12530 1747
rect 12778 1739 12786 1747
rect 12858 1739 12866 1747
rect 12938 1739 12946 1747
rect 13626 1739 13634 1747
rect 14218 1739 14226 1747
rect 14970 1739 14978 1747
rect 15514 1739 15522 1747
rect 15626 1739 15634 1747
rect 16922 1739 16930 1747
rect 16938 1739 16946 1747
rect 17034 1739 17042 1747
rect 17274 1739 17282 1747
rect 18848 1740 18856 1748
rect 19696 1740 19704 1748
rect 19904 1740 19912 1748
rect 19952 1740 19960 1748
rect 20576 1740 20584 1748
rect 21984 1740 21992 1748
rect 22192 1740 22200 1748
rect 22592 1740 22600 1748
rect 22688 1740 22696 1748
rect 23264 1740 23272 1748
rect 23552 1740 23560 1748
rect 23760 1740 23768 1748
rect 24096 1740 24104 1748
rect 24176 1740 24184 1748
rect 27360 1740 27368 1748
rect 27584 1740 27592 1748
rect 28416 1740 28424 1748
rect 34720 1737 34728 1745
rect 35392 1737 35400 1745
rect 36304 1737 36312 1745
rect 36432 1737 36440 1745
rect 1176 1719 1184 1727
rect 2344 1719 2352 1727
rect 2360 1719 2368 1727
rect 3752 1719 3760 1727
rect 10098 1713 10106 1721
rect 13658 1719 13666 1727
rect 13898 1719 13906 1727
rect 15322 1719 15330 1727
rect 15818 1719 15826 1727
rect 16330 1719 16338 1727
rect 16538 1719 16546 1727
rect 21568 1720 21576 1728
rect 26016 1720 26024 1728
rect 26944 1720 26952 1728
rect 27152 1720 27160 1728
rect 30000 1717 30008 1725
rect 39168 1717 39176 1725
rect 2696 1699 2704 1707
rect 3800 1699 3808 1707
rect 4200 1699 4208 1707
rect 7954 1693 7962 1701
rect 9714 1693 9722 1701
rect 10674 1693 10682 1701
rect 10722 1693 10730 1701
rect 13866 1699 13874 1707
rect 15706 1699 15714 1707
rect 18928 1700 18936 1708
rect 24736 1700 24744 1708
rect 39296 1697 39304 1705
rect 632 1679 640 1687
rect 1096 1679 1104 1687
rect 1224 1679 1232 1687
rect 1608 1679 1616 1687
rect 1976 1679 1984 1687
rect 2056 1679 2064 1687
rect 2248 1679 2256 1687
rect 2776 1679 2784 1687
rect 3560 1679 3568 1687
rect 4008 1679 4016 1687
rect 4104 1679 4112 1687
rect 4504 1679 4512 1687
rect 4552 1679 4560 1687
rect 4568 1679 4576 1687
rect 4600 1679 4608 1687
rect 5874 1673 5882 1681
rect 6578 1673 6586 1681
rect 6674 1673 6682 1681
rect 7362 1673 7370 1681
rect 7394 1673 7402 1681
rect 7618 1673 7626 1681
rect 7922 1673 7930 1681
rect 8562 1673 8570 1681
rect 8642 1673 8650 1681
rect 8802 1673 8810 1681
rect 8962 1673 8970 1681
rect 9762 1673 9770 1681
rect 9906 1673 9914 1681
rect 10002 1673 10010 1681
rect 13130 1679 13138 1687
rect 13818 1679 13826 1687
rect 14090 1679 14098 1687
rect 16714 1679 16722 1687
rect 22224 1680 22232 1688
rect 29396 1667 29408 1675
rect 29428 1667 29440 1675
rect 29444 1667 29448 1675
rect 29460 1667 29472 1675
rect 29488 1667 29504 1675
rect 29512 1667 29544 1675
rect 29552 1667 29564 1675
rect 29580 1667 29596 1675
rect 29604 1667 29636 1675
rect 29644 1667 29660 1675
rect 29676 1667 29688 1675
rect 29700 1667 29704 1675
rect 29708 1667 29720 1675
rect 29740 1667 29752 1675
rect 29772 1667 29784 1675
rect 29788 1667 29792 1675
rect 29804 1667 29816 1675
rect 29832 1667 29848 1675
rect 29856 1667 29888 1675
rect 29896 1667 29912 1675
rect 29920 1667 29944 1675
rect 29960 1667 29964 1675
rect 29968 1667 29980 1675
rect 29984 1667 29996 1675
rect 30000 1667 30004 1675
rect 30020 1667 30024 1675
rect 30028 1667 30032 1675
rect 30052 1667 30056 1675
rect 30060 1667 30072 1675
rect 30076 1667 30088 1675
rect 30092 1667 30096 1675
rect 30112 1667 30128 1675
rect 30144 1667 30148 1675
rect 30152 1667 30164 1675
rect 30168 1667 30180 1675
rect 30184 1667 30188 1675
rect 30236 1667 30240 1675
rect 30244 1667 30256 1675
rect 30260 1667 30272 1675
rect 30276 1667 30280 1675
rect 30296 1667 30312 1675
rect 30328 1667 30332 1675
rect 30336 1667 30348 1675
rect 30352 1667 30364 1675
rect 30368 1667 30372 1675
rect 30392 1667 30396 1675
rect 30400 1667 30404 1675
rect 30420 1667 30424 1675
rect 30428 1667 30440 1675
rect 30444 1667 30456 1675
rect 30460 1667 30464 1675
rect 30484 1667 30488 1675
rect 30492 1667 30504 1675
rect 30516 1667 30520 1675
rect 30524 1667 30528 1675
rect 30548 1667 30552 1675
rect 30556 1667 30568 1675
rect 30580 1667 30584 1675
rect 30588 1667 30592 1675
rect 30604 1667 30616 1675
rect 30620 1667 30624 1675
rect 30644 1667 30648 1675
rect 30652 1667 30656 1675
rect 30668 1667 30680 1675
rect 30684 1667 30688 1675
rect 30708 1667 30712 1675
rect 30716 1667 30728 1675
rect 30740 1667 30744 1675
rect 30748 1667 30752 1675
rect 30864 1667 30868 1675
rect 30872 1667 30876 1675
rect 30940 1667 30944 1675
rect 30948 1667 30952 1675
rect 31032 1667 31036 1675
rect 31040 1667 31044 1675
rect 31064 1667 31068 1675
rect 31072 1667 31084 1675
rect 31088 1667 31100 1675
rect 31104 1667 31108 1675
rect 31128 1667 31132 1675
rect 31136 1667 31148 1675
rect 31156 1667 31172 1675
rect 31180 1667 31212 1675
rect 31220 1667 31236 1675
rect 31252 1667 31264 1675
rect 31272 1667 31304 1675
rect 31312 1667 31324 1675
rect 31340 1667 31356 1675
rect 31364 1667 31396 1675
rect 31404 1667 31420 1675
rect 31428 1667 31452 1675
rect 31464 1667 31488 1675
rect 31496 1667 31512 1675
rect 31520 1667 31544 1675
rect 31556 1667 31580 1675
rect 31588 1667 31604 1675
rect 31612 1667 31636 1675
rect 31652 1667 31656 1675
rect 31660 1667 31672 1675
rect 31684 1667 31688 1675
rect 31692 1667 31696 1675
rect 31716 1667 31720 1675
rect 31724 1667 31736 1675
rect 31808 1667 31812 1675
rect 31816 1667 31828 1675
rect 31848 1667 31860 1675
rect 31864 1667 31876 1675
rect 31880 1667 31884 1675
rect 31904 1667 31908 1675
rect 31912 1667 31916 1675
rect 31932 1667 31936 1675
rect 31940 1667 31952 1675
rect 31956 1667 31960 1675
rect 32160 1667 32172 1675
rect 32176 1667 32188 1675
rect 32192 1667 32204 1675
rect 32224 1667 32236 1675
rect 32248 1667 32252 1675
rect 32256 1667 32268 1675
rect 32288 1667 32300 1675
rect 32380 1667 32392 1675
rect 32412 1667 32424 1675
rect 32428 1667 32432 1675
rect 32444 1667 32456 1675
rect 32476 1667 32488 1675
rect 32500 1667 32504 1675
rect 32508 1667 32520 1675
rect 32540 1667 32552 1675
rect 32572 1667 32584 1675
rect 32588 1667 32592 1675
rect 32604 1667 32616 1675
rect 32636 1667 32648 1675
rect 32660 1667 32664 1675
rect 32668 1667 32680 1675
rect 32856 1667 32868 1675
rect 32980 1667 32992 1675
rect 32996 1667 33000 1675
rect 33012 1667 33024 1675
rect 33040 1667 33056 1675
rect 33064 1667 33096 1675
rect 33104 1667 33120 1675
rect 33128 1667 33140 1675
rect 33144 1667 33148 1675
rect 33168 1667 33172 1675
rect 33176 1667 33188 1675
rect 33200 1667 33204 1675
rect 33208 1667 33212 1675
rect 33308 1667 33312 1675
rect 33316 1667 33320 1675
rect 33340 1667 33344 1675
rect 33348 1667 33360 1675
rect 33364 1667 33376 1675
rect 33380 1667 33384 1675
rect 33404 1667 33408 1675
rect 33412 1667 33416 1675
rect 33432 1667 33448 1675
rect 33456 1667 33480 1675
rect 33496 1667 33508 1675
rect 33512 1667 33516 1675
rect 33528 1667 33540 1675
rect 33552 1667 33556 1675
rect 33560 1667 33572 1675
rect 33576 1667 33580 1675
rect 33684 1667 33696 1675
rect 33808 1667 33820 1675
rect 33824 1667 33828 1675
rect 33840 1667 33852 1675
rect 33868 1667 33884 1675
rect 33892 1667 33924 1675
rect 33932 1667 33948 1675
rect 33964 1667 33980 1675
rect 33996 1667 34000 1675
rect 34004 1667 34016 1675
rect 34028 1667 34032 1675
rect 34036 1667 34040 1675
rect 34052 1667 34064 1675
rect 34068 1667 34072 1675
rect 34120 1667 34124 1675
rect 34128 1667 34132 1675
rect 34212 1667 34216 1675
rect 34220 1667 34224 1675
rect 34304 1667 34308 1675
rect 34312 1667 34316 1675
rect 34328 1667 34340 1675
rect 34344 1667 34348 1675
rect 34368 1667 34372 1675
rect 34376 1667 34380 1675
rect 34400 1667 34412 1675
rect 34420 1667 34452 1675
rect 34460 1667 34476 1675
rect 34492 1667 34508 1675
rect 34524 1667 34528 1675
rect 34532 1667 34544 1675
rect 34556 1667 34560 1675
rect 34564 1667 34568 1675
rect 34580 1667 34592 1675
rect 34596 1667 34600 1675
rect 34680 1667 34684 1675
rect 34688 1667 34692 1675
rect 34804 1667 34808 1675
rect 34812 1667 34816 1675
rect 34828 1667 34840 1675
rect 34844 1667 34848 1675
rect 34912 1667 34916 1675
rect 34920 1667 34924 1675
rect 34944 1667 34948 1675
rect 34952 1667 34956 1675
rect 34968 1667 34980 1675
rect 34984 1667 34996 1675
rect 35008 1667 35012 1675
rect 35016 1667 35020 1675
rect 35036 1667 35084 1675
rect 35100 1667 35104 1675
rect 35108 1667 35112 1675
rect 35128 1667 35176 1675
rect 35192 1667 35196 1675
rect 35200 1667 35204 1675
rect 35220 1667 35268 1675
rect 35284 1667 35296 1675
rect 35300 1667 35304 1675
rect 35316 1667 35328 1675
rect 35336 1667 35360 1675
rect 35376 1667 35400 1675
rect 35408 1667 35424 1675
rect 35440 1667 35444 1675
rect 35448 1667 35452 1675
rect 35472 1667 35476 1675
rect 35480 1667 35492 1675
rect 35496 1667 35508 1675
rect 35512 1667 35516 1675
rect 35532 1667 35548 1675
rect 35564 1667 35568 1675
rect 35572 1667 35584 1675
rect 35588 1667 35600 1675
rect 35604 1667 35608 1675
rect 35628 1667 35632 1675
rect 35636 1667 35640 1675
rect 35656 1667 35660 1675
rect 35664 1667 35676 1675
rect 35680 1667 35692 1675
rect 35696 1667 35700 1675
rect 35720 1667 35724 1675
rect 35728 1667 35732 1675
rect 35748 1667 35752 1675
rect 35756 1667 35768 1675
rect 35772 1667 35784 1675
rect 35788 1667 35792 1675
rect 35812 1667 35816 1675
rect 35820 1667 35824 1675
rect 35920 1667 35924 1675
rect 35928 1667 35932 1675
rect 35944 1667 35956 1675
rect 35960 1667 35964 1675
rect 36012 1667 36016 1675
rect 36020 1667 36024 1675
rect 36036 1667 36048 1675
rect 36052 1667 36056 1675
rect 36104 1667 36108 1675
rect 36112 1667 36116 1675
rect 36128 1667 36140 1675
rect 36144 1667 36148 1675
rect 36468 1667 36472 1675
rect 36476 1667 36480 1675
rect 36492 1667 36504 1675
rect 36508 1667 36512 1675
rect 36532 1667 36536 1675
rect 36540 1667 36544 1675
rect 36560 1667 36608 1675
rect 36624 1667 36640 1675
rect 36656 1667 36672 1675
rect 36688 1667 36704 1675
rect 36720 1667 36768 1675
rect 36784 1667 36788 1675
rect 36792 1667 36796 1675
rect 36812 1667 36860 1675
rect 36876 1667 36880 1675
rect 36884 1667 36888 1675
rect 36904 1667 36952 1675
rect 36968 1667 36972 1675
rect 36976 1667 36980 1675
rect 36996 1667 37044 1675
rect 37060 1667 37084 1675
rect 37092 1667 37104 1675
rect 37116 1667 37120 1675
rect 37124 1667 37136 1675
rect 37156 1667 37168 1675
rect 37188 1667 37200 1675
rect 37220 1667 37232 1675
rect 37236 1667 37240 1675
rect 37252 1667 37264 1675
rect 37272 1667 37296 1675
rect 37312 1667 37336 1675
rect 37344 1667 37356 1675
rect 37364 1667 37388 1675
rect 37404 1667 37428 1675
rect 37436 1667 37448 1675
rect 37460 1667 37464 1675
rect 37468 1667 37480 1675
rect 37496 1667 37520 1675
rect 37528 1667 37540 1675
rect 37552 1667 37556 1675
rect 37560 1667 37572 1675
rect 37588 1667 37636 1675
rect 37652 1667 37668 1675
rect 37684 1667 37696 1675
rect 37708 1667 37712 1675
rect 37716 1667 37728 1675
rect 37840 1667 37852 1675
rect 37856 1667 37868 1675
rect 37872 1667 37884 1675
rect 37900 1667 37916 1675
rect 37932 1667 37956 1675
rect 37964 1667 37980 1675
rect 37996 1667 38012 1675
rect 38020 1667 38032 1675
rect 38036 1667 38048 1675
rect 38056 1667 38072 1675
rect 38088 1667 38104 1675
rect 38112 1667 38124 1675
rect 38128 1667 38140 1675
rect 38152 1667 38156 1675
rect 38160 1667 38164 1675
rect 38180 1667 38196 1675
rect 38204 1667 38228 1675
rect 38244 1667 38256 1675
rect 38276 1667 38288 1675
rect 38292 1667 38304 1675
rect 38308 1667 38320 1675
rect 38336 1667 38352 1675
rect 38368 1667 38380 1675
rect 38384 1667 38396 1675
rect 38400 1667 38412 1675
rect 38432 1667 38444 1675
rect 38448 1667 38452 1675
rect 38484 1667 38488 1675
rect 38492 1667 38504 1675
rect 38524 1667 38536 1675
rect 38540 1667 38552 1675
rect 38556 1667 38568 1675
rect 38584 1667 38600 1675
rect 38616 1667 38640 1675
rect 38648 1667 38664 1675
rect 38680 1667 38684 1675
rect 38688 1667 38692 1675
rect 38704 1667 38716 1675
rect 38720 1667 38732 1675
rect 38740 1667 38756 1675
rect 38772 1667 38788 1675
rect 38796 1667 38820 1675
rect 38836 1667 38852 1675
rect 38868 1667 38880 1675
rect 38884 1667 38896 1675
rect 38900 1667 38912 1675
rect 38928 1667 38944 1675
rect 38960 1667 38984 1675
rect 38992 1667 39008 1675
rect 39024 1667 39040 1675
rect 39048 1667 39060 1675
rect 39064 1667 39076 1675
rect 39088 1667 39092 1675
rect 39096 1667 39100 1675
rect 39112 1667 39124 1675
rect 39128 1667 39132 1675
rect 39388 1667 39392 1675
rect 39396 1667 39400 1675
rect 39528 1667 39532 1675
rect 39536 1667 39540 1675
rect 39552 1667 39564 1675
rect 39568 1667 39580 1675
rect 39588 1667 39604 1675
rect 39620 1667 39668 1675
rect 39684 1667 39700 1675
rect 39712 1667 39760 1675
rect 39776 1667 39792 1675
rect 39808 1667 39820 1675
rect 39832 1667 39836 1675
rect 39840 1667 39852 1675
rect 39872 1667 39884 1675
rect 39888 1667 39892 1675
rect 40248 1667 40260 1675
rect 40264 1667 40268 1675
rect 40280 1667 40292 1675
rect 40308 1667 40324 1675
rect 40340 1667 40388 1675
rect 40404 1667 40408 1675
rect 40412 1667 40416 1675
rect 40436 1667 40440 1675
rect 40444 1667 40456 1675
rect 40468 1667 40472 1675
rect 40476 1667 40480 1675
rect 40500 1667 40504 1675
rect 40508 1667 40520 1675
rect 40524 1667 40536 1675
rect 40540 1667 40544 1675
rect 40564 1667 40568 1675
rect 40572 1667 40576 1675
rect 40592 1667 40608 1675
rect 40616 1667 40640 1675
rect 40656 1667 40680 1675
rect 40688 1667 40704 1675
rect 40720 1667 40736 1675
rect 40752 1667 40768 1675
rect 40776 1667 40800 1675
rect 820 1663 844 1667
rect 1192 1659 1200 1667
rect 1608 1659 1616 1667
rect 2776 1659 2784 1667
rect 3444 1663 3468 1667
rect 3928 1659 3936 1667
rect 4584 1659 4592 1667
rect 8002 1653 8010 1661
rect 9106 1653 9114 1661
rect 9234 1653 9242 1661
rect 19394 1650 19396 1658
rect 19402 1650 19404 1658
rect 20448 1650 20450 1658
rect 20456 1650 20458 1658
rect 22746 1650 22756 1658
rect 24792 1650 24800 1658
rect 25532 1650 25536 1658
rect 25540 1650 25544 1658
rect 25608 1650 25612 1658
rect 25616 1650 25620 1658
rect 25960 1650 25964 1658
rect 25968 1650 25972 1658
rect 26036 1650 26040 1658
rect 26044 1650 26048 1658
rect 26174 1650 26178 1658
rect 26182 1650 26186 1658
rect 26250 1650 26254 1658
rect 26258 1650 26262 1658
rect 26602 1650 26606 1658
rect 26610 1650 26614 1658
rect 26678 1650 26682 1658
rect 26686 1650 26690 1658
rect 26816 1650 26820 1658
rect 26824 1650 26828 1658
rect 26892 1650 26896 1658
rect 26900 1650 26904 1658
rect 27564 1650 27570 1658
rect 27572 1650 27578 1658
rect 27640 1650 27646 1658
rect 27648 1650 27654 1658
rect 27862 1650 27874 1658
rect 27976 1650 27982 1658
rect 27984 1650 27990 1658
rect 28052 1650 28058 1658
rect 28060 1650 28066 1658
rect 33344 1657 33352 1665
rect 2840 1639 2848 1647
rect 6402 1633 6410 1641
rect 8466 1633 8474 1641
rect 9202 1633 9210 1641
rect 9858 1633 9866 1641
rect 9906 1633 9914 1641
rect 10482 1633 10490 1641
rect 16026 1639 16034 1647
rect 25120 1640 25128 1648
rect 31824 1637 31832 1645
rect 36208 1637 36216 1645
rect 504 1619 512 1627
rect 584 1619 592 1627
rect 808 1619 816 1627
rect 1192 1619 1200 1627
rect 1736 1619 1744 1627
rect 1896 1619 1904 1627
rect 2616 1619 2624 1627
rect 2936 1619 2944 1627
rect 3080 1619 3088 1627
rect 3144 1619 3152 1627
rect 3336 1619 3344 1627
rect 3608 1619 3616 1627
rect 3768 1619 3776 1627
rect 4216 1619 4224 1627
rect 4536 1619 4544 1627
rect 6162 1613 6170 1621
rect 7282 1613 7290 1621
rect 8466 1613 8474 1621
rect 8642 1613 8650 1621
rect 8866 1613 8874 1621
rect 9042 1613 9050 1621
rect 9106 1613 9114 1621
rect 9506 1613 9514 1621
rect 9746 1613 9754 1621
rect 9922 1613 9930 1621
rect 10482 1613 10490 1621
rect 10530 1613 10538 1621
rect 10546 1613 10554 1621
rect 15690 1619 15698 1627
rect 15706 1619 15714 1627
rect 16506 1619 16514 1627
rect 16522 1619 16530 1627
rect 21584 1620 21592 1628
rect 648 1599 656 1607
rect 920 1599 928 1607
rect 1272 1599 1280 1607
rect 1752 1599 1760 1607
rect 2104 1599 2112 1607
rect 3480 1599 3488 1607
rect 4008 1599 4016 1607
rect 4040 1599 4048 1607
rect 6962 1593 6970 1601
rect 7906 1593 7914 1601
rect 8162 1593 8170 1601
rect 13018 1599 13026 1607
rect 13626 1599 13634 1607
rect 13642 1599 13650 1607
rect 14042 1599 14050 1607
rect 16714 1599 16722 1607
rect 19296 1600 19304 1608
rect 24480 1600 24488 1608
rect 25984 1600 25992 1608
rect 26144 1600 26152 1608
rect 26224 1600 26232 1608
rect 27632 1600 27640 1608
rect 31680 1597 31688 1605
rect 32032 1597 32040 1605
rect 36032 1597 36040 1605
rect 36048 1597 36056 1605
rect 36816 1597 36824 1605
rect 37376 1597 37384 1605
rect 2808 1579 2816 1587
rect 2984 1579 2992 1587
rect 4136 1579 4144 1587
rect 4376 1579 4384 1587
rect 6930 1573 6938 1581
rect 7506 1573 7514 1581
rect 8034 1573 8042 1581
rect 8850 1573 8858 1581
rect 8962 1573 8970 1581
rect 9058 1573 9066 1581
rect 9074 1573 9082 1581
rect 9218 1573 9226 1581
rect 9378 1573 9386 1581
rect 9986 1573 9994 1581
rect 10034 1573 10042 1581
rect 10114 1573 10122 1581
rect 10194 1573 10202 1581
rect 10594 1573 10602 1581
rect 13146 1579 13154 1587
rect 13210 1579 13218 1587
rect 13402 1579 13410 1587
rect 14026 1579 14034 1587
rect 14218 1579 14226 1587
rect 15450 1579 15458 1587
rect 16010 1579 16018 1587
rect 16106 1579 16114 1587
rect 16202 1579 16210 1587
rect 16954 1579 16962 1587
rect 17162 1579 17170 1587
rect 23888 1580 23896 1588
rect 27744 1580 27752 1588
rect 29840 1577 29848 1585
rect 30096 1577 30104 1585
rect 31120 1577 31128 1585
rect 31648 1577 31656 1585
rect 31664 1577 31672 1585
rect 32720 1577 32728 1585
rect 32864 1577 32872 1585
rect 36192 1577 36200 1585
rect 37456 1577 37464 1585
rect 37808 1577 37816 1585
rect 37984 1577 37992 1585
rect 38080 1577 38088 1585
rect 38144 1577 38152 1585
rect 38736 1577 38744 1585
rect 38816 1577 38824 1585
rect 39104 1577 39112 1585
rect 936 1559 944 1567
rect 1000 1559 1008 1567
rect 1032 1559 1040 1567
rect 1144 1559 1152 1567
rect 1304 1559 1312 1567
rect 1336 1559 1344 1567
rect 1608 1559 1616 1567
rect 1656 1559 1664 1567
rect 2744 1559 2752 1567
rect 2760 1559 2768 1567
rect 2808 1559 2816 1567
rect 3064 1559 3072 1567
rect 3304 1559 3312 1567
rect 3352 1559 3360 1567
rect 3576 1559 3584 1567
rect 3848 1559 3856 1567
rect 4472 1559 4480 1567
rect 4504 1559 4512 1567
rect 4584 1559 4592 1567
rect 4632 1559 4640 1567
rect 4664 1559 4672 1567
rect 5810 1553 5818 1561
rect 5826 1553 5834 1561
rect 6050 1553 6058 1561
rect 6306 1553 6314 1561
rect 6914 1553 6922 1561
rect 7426 1553 7434 1561
rect 8018 1553 8026 1561
rect 8050 1553 8058 1561
rect 8626 1553 8634 1561
rect 9058 1553 9066 1561
rect 9122 1553 9130 1561
rect 9202 1553 9210 1561
rect 9650 1553 9658 1561
rect 9730 1553 9738 1561
rect 10754 1553 10762 1561
rect 10834 1553 10842 1561
rect 13722 1559 13730 1567
rect 14154 1559 14162 1567
rect 14314 1559 14322 1567
rect 14410 1559 14418 1567
rect 14554 1559 14562 1567
rect 14666 1559 14674 1567
rect 14874 1559 14882 1567
rect 15034 1559 15042 1567
rect 15130 1559 15138 1567
rect 15162 1559 15170 1567
rect 15194 1559 15202 1567
rect 15882 1559 15890 1567
rect 16026 1559 16034 1567
rect 16122 1559 16130 1567
rect 16538 1559 16546 1567
rect 16634 1559 16642 1567
rect 16682 1559 16690 1567
rect 16730 1559 16738 1567
rect 17258 1559 17266 1567
rect 17306 1559 17314 1567
rect 17354 1559 17362 1567
rect 17434 1559 17442 1567
rect 18656 1560 18664 1568
rect 19072 1561 19082 1566
rect 19456 1560 19464 1568
rect 19468 1561 19478 1566
rect 19744 1560 19752 1568
rect 20160 1560 20168 1568
rect 20576 1560 20584 1568
rect 21378 1561 21388 1566
rect 21774 1561 21784 1566
rect 21968 1560 21976 1568
rect 23088 1560 23096 1568
rect 23520 1560 23528 1568
rect 23728 1560 23736 1568
rect 24272 1560 24280 1568
rect 24288 1560 24296 1568
rect 24544 1560 24552 1568
rect 24736 1560 24744 1568
rect 26416 1560 26424 1568
rect 26848 1560 26856 1568
rect 27056 1560 27064 1568
rect 28096 1560 28104 1568
rect 29792 1557 29800 1565
rect 30496 1557 30504 1565
rect 30640 1557 30648 1565
rect 32976 1557 32984 1565
rect 36128 1557 36136 1565
rect 36336 1557 36344 1565
rect 37776 1557 37784 1565
rect 39808 1557 39816 1565
rect 40688 1557 40696 1565
rect 1816 1539 1824 1547
rect 6578 1533 6586 1541
rect 6626 1533 6634 1541
rect 7378 1533 7386 1541
rect 7458 1533 7466 1541
rect 7682 1533 7690 1541
rect 7778 1533 7786 1541
rect 8226 1533 8234 1541
rect 8274 1533 8282 1541
rect 8498 1533 8506 1541
rect 8738 1533 8746 1541
rect 9906 1533 9914 1541
rect 10258 1533 10266 1541
rect 10850 1533 10858 1541
rect 12442 1539 12450 1547
rect 12682 1539 12690 1547
rect 13258 1539 13266 1547
rect 13466 1539 13474 1547
rect 13482 1539 13490 1547
rect 14426 1539 14434 1547
rect 14538 1539 14546 1547
rect 15322 1539 15330 1547
rect 15434 1539 15442 1547
rect 15834 1539 15842 1547
rect 17098 1539 17106 1547
rect 17226 1539 17234 1547
rect 19536 1540 19544 1548
rect 20592 1540 20600 1548
rect 20976 1540 20984 1548
rect 21200 1540 21208 1548
rect 21376 1540 21384 1548
rect 21392 1540 21400 1548
rect 21424 1540 21432 1548
rect 22432 1540 22440 1548
rect 26224 1540 26232 1548
rect 29616 1537 29624 1545
rect 29856 1537 29864 1545
rect 30496 1537 30504 1545
rect 30976 1537 30984 1545
rect 31344 1537 31352 1545
rect 31600 1537 31608 1545
rect 31840 1537 31848 1545
rect 32016 1537 32024 1545
rect 32128 1537 32136 1545
rect 32320 1537 32328 1545
rect 32608 1537 32616 1545
rect 32880 1537 32888 1545
rect 33248 1537 33256 1545
rect 33376 1537 33384 1545
rect 34720 1537 34728 1545
rect 35120 1537 35128 1545
rect 35680 1537 35688 1545
rect 36896 1537 36904 1545
rect 37440 1537 37448 1545
rect 37648 1537 37656 1545
rect 37696 1537 37704 1545
rect 38992 1537 39000 1545
rect 39088 1537 39096 1545
rect 40672 1537 40680 1545
rect 568 1519 576 1527
rect 600 1519 608 1527
rect 712 1519 720 1527
rect 1000 1519 1008 1527
rect 1096 1519 1104 1527
rect 1336 1519 1344 1527
rect 1368 1519 1376 1527
rect 1544 1519 1552 1527
rect 1992 1519 2000 1527
rect 2104 1519 2112 1527
rect 2424 1519 2432 1527
rect 2488 1519 2496 1527
rect 2680 1519 2688 1527
rect 2872 1519 2880 1527
rect 2920 1519 2928 1527
rect 3000 1519 3008 1527
rect 3016 1519 3024 1527
rect 3128 1519 3136 1527
rect 3928 1519 3936 1527
rect 3992 1519 4000 1527
rect 4168 1519 4176 1527
rect 4408 1519 4416 1527
rect 5730 1513 5738 1521
rect 5922 1513 5930 1521
rect 7474 1513 7482 1521
rect 7522 1513 7530 1521
rect 7586 1513 7594 1521
rect 7746 1513 7754 1521
rect 7810 1513 7818 1521
rect 7954 1513 7962 1521
rect 9874 1513 9882 1521
rect 10322 1513 10330 1521
rect 10370 1513 10378 1521
rect 10546 1513 10554 1521
rect 10706 1513 10714 1521
rect 12154 1519 12162 1527
rect 12170 1519 12178 1527
rect 12858 1519 12866 1527
rect 13098 1519 13106 1527
rect 13450 1519 13458 1527
rect 13498 1519 13506 1527
rect 13690 1519 13698 1527
rect 13722 1519 13730 1527
rect 13754 1519 13762 1527
rect 13946 1519 13954 1527
rect 14282 1519 14290 1527
rect 14490 1519 14498 1527
rect 14762 1519 14770 1527
rect 14938 1519 14946 1527
rect 14954 1519 14962 1527
rect 15658 1519 15666 1527
rect 18640 1520 18648 1528
rect 19728 1520 19736 1528
rect 19760 1520 19768 1528
rect 20496 1520 20504 1528
rect 21024 1520 21032 1528
rect 22480 1520 22488 1528
rect 22624 1520 22632 1528
rect 23104 1520 23112 1528
rect 23312 1520 23320 1528
rect 24256 1520 24264 1528
rect 24288 1520 24296 1528
rect 24752 1520 24760 1528
rect 25136 1520 25144 1528
rect 26208 1520 26216 1528
rect 28112 1520 28120 1528
rect 34992 1517 35000 1525
rect 35040 1517 35048 1525
rect 35296 1517 35304 1525
rect 35488 1517 35496 1525
rect 36560 1517 36568 1525
rect 37792 1517 37800 1525
rect 37872 1517 37880 1525
rect 38832 1517 38840 1525
rect 39072 1517 39080 1525
rect 39152 1517 39160 1525
rect 37688 1511 37696 1513
rect 40456 1511 40464 1513
rect 424 1499 432 1507
rect 488 1499 496 1507
rect 520 1499 528 1507
rect 600 1499 608 1507
rect 632 1499 640 1507
rect 664 1499 672 1507
rect 792 1499 800 1507
rect 824 1499 832 1507
rect 904 1499 912 1507
rect 936 1499 944 1507
rect 1032 1499 1040 1507
rect 1208 1499 1216 1507
rect 1288 1499 1296 1507
rect 1368 1499 1376 1507
rect 1400 1499 1408 1507
rect 1576 1499 1584 1507
rect 1720 1499 1728 1507
rect 1768 1499 1776 1507
rect 1880 1499 1888 1507
rect 1944 1499 1952 1507
rect 1960 1499 1968 1507
rect 2040 1499 2048 1507
rect 2184 1499 2192 1507
rect 2200 1499 2208 1507
rect 2600 1499 2608 1507
rect 2904 1499 2912 1507
rect 2952 1499 2960 1507
rect 3096 1499 3104 1507
rect 3160 1499 3168 1507
rect 3320 1499 3328 1507
rect 3400 1499 3408 1507
rect 3432 1499 3440 1507
rect 3512 1499 3520 1507
rect 3784 1499 3792 1507
rect 3992 1499 4000 1507
rect 4376 1499 4384 1507
rect 4440 1499 4448 1507
rect 4504 1499 4512 1507
rect 4520 1499 4528 1507
rect 4600 1499 4608 1507
rect 5874 1493 5882 1501
rect 5938 1493 5946 1501
rect 6066 1493 6074 1501
rect 6098 1493 6106 1501
rect 6178 1493 6186 1501
rect 6258 1493 6266 1501
rect 6594 1493 6602 1501
rect 7074 1493 7082 1501
rect 7090 1493 7098 1501
rect 7138 1493 7146 1501
rect 7266 1493 7274 1501
rect 7330 1493 7338 1501
rect 7842 1493 7850 1501
rect 7906 1493 7914 1501
rect 8050 1493 8058 1501
rect 8610 1493 8618 1501
rect 8802 1493 8810 1501
rect 8978 1493 8986 1501
rect 9058 1493 9066 1501
rect 9090 1493 9098 1501
rect 9122 1493 9130 1501
rect 9346 1493 9354 1501
rect 9474 1493 9482 1501
rect 9490 1493 9498 1501
rect 9938 1493 9946 1501
rect 9954 1493 9962 1501
rect 10098 1493 10106 1501
rect 10418 1493 10426 1501
rect 10434 1493 10442 1501
rect 10674 1493 10682 1501
rect 10866 1493 10874 1501
rect 12042 1499 12050 1507
rect 12170 1499 12178 1507
rect 12618 1499 12626 1507
rect 12746 1499 12754 1507
rect 13082 1499 13090 1507
rect 13146 1499 13154 1507
rect 13290 1499 13298 1507
rect 13322 1499 13330 1507
rect 13370 1499 13378 1507
rect 14730 1499 14738 1507
rect 14922 1499 14930 1507
rect 15146 1499 15154 1507
rect 15178 1499 15186 1507
rect 15626 1499 15634 1507
rect 15642 1499 15650 1507
rect 15898 1499 15906 1507
rect 16074 1499 16082 1507
rect 16138 1499 16146 1507
rect 16586 1499 16594 1507
rect 17178 1499 17186 1507
rect 21760 1500 21768 1508
rect 22160 1500 22168 1508
rect 22704 1500 22712 1508
rect 24080 1500 24088 1508
rect 24448 1500 24456 1508
rect 25776 1500 25784 1508
rect 37682 1505 37696 1511
rect 40450 1505 40464 1511
rect 30672 1497 30680 1505
rect 31776 1497 31784 1505
rect 33088 1497 33096 1505
rect 33568 1497 33576 1505
rect 34048 1497 34056 1505
rect 34640 1497 34648 1505
rect 36912 1497 36920 1505
rect 37120 1497 37128 1505
rect 37184 1497 37192 1505
rect 37680 1497 37688 1505
rect 37744 1497 37752 1505
rect 37840 1497 37848 1505
rect 38432 1497 38440 1505
rect 39952 1497 39960 1505
rect 40448 1497 40456 1505
rect 40784 1497 40792 1505
rect 744 1479 752 1487
rect 1064 1479 1072 1487
rect 1240 1479 1248 1487
rect 1528 1479 1536 1487
rect 1624 1479 1632 1487
rect 1784 1479 1792 1487
rect 2056 1479 2064 1487
rect 2504 1479 2512 1487
rect 2632 1479 2640 1487
rect 2808 1479 2816 1487
rect 3192 1479 3200 1487
rect 3240 1479 3248 1487
rect 4040 1479 4048 1487
rect 4120 1479 4128 1487
rect 4568 1479 4576 1487
rect 6658 1473 6666 1481
rect 8114 1473 8122 1481
rect 8402 1473 8410 1481
rect 9170 1473 9178 1481
rect 9330 1473 9338 1481
rect 10594 1473 10602 1481
rect 12762 1479 12770 1487
rect 12954 1479 12962 1487
rect 14794 1479 14802 1487
rect 17290 1479 17298 1487
rect 20112 1480 20120 1488
rect 20336 1480 20344 1488
rect 22832 1480 22840 1488
rect 24688 1480 24696 1488
rect 24816 1480 24824 1488
rect 27440 1480 27448 1488
rect 31728 1477 31736 1485
rect 34400 1477 34408 1485
rect 39712 1477 39720 1485
rect 1768 1459 1776 1467
rect 2136 1459 2144 1467
rect 2168 1459 2176 1467
rect 2984 1459 2992 1467
rect 3304 1459 3312 1467
rect 3992 1459 4000 1467
rect 6946 1453 6954 1461
rect 7858 1453 7866 1461
rect 8370 1453 8378 1461
rect 8610 1453 8618 1461
rect 8930 1453 8938 1461
rect 9970 1453 9978 1461
rect 10242 1453 10250 1461
rect 10386 1453 10394 1461
rect 10594 1453 10602 1461
rect 13370 1459 13378 1467
rect 14234 1459 14242 1467
rect 15370 1459 15378 1467
rect 15498 1459 15506 1467
rect 15530 1459 15538 1467
rect 16618 1459 16626 1467
rect 20768 1460 20776 1468
rect 27008 1460 27016 1468
rect 29396 1467 29408 1475
rect 29428 1467 29440 1475
rect 29444 1467 29448 1475
rect 29460 1467 29472 1475
rect 29488 1467 29504 1475
rect 29512 1467 29544 1475
rect 29552 1467 29568 1475
rect 29576 1467 29588 1475
rect 29592 1467 29596 1475
rect 29616 1467 29620 1475
rect 29624 1467 29636 1475
rect 29644 1467 29660 1475
rect 29668 1467 29692 1475
rect 29708 1467 29724 1475
rect 29732 1467 29756 1475
rect 29772 1467 29796 1475
rect 29804 1467 29816 1475
rect 29824 1467 29848 1475
rect 29864 1467 29888 1475
rect 29896 1467 29908 1475
rect 29920 1467 29924 1475
rect 29928 1467 29940 1475
rect 29956 1467 29980 1475
rect 29988 1467 30004 1475
rect 30020 1467 30024 1475
rect 30028 1467 30032 1475
rect 30052 1467 30056 1475
rect 30060 1467 30072 1475
rect 30076 1467 30088 1475
rect 30092 1467 30096 1475
rect 30116 1467 30120 1475
rect 30124 1467 30128 1475
rect 30192 1467 30196 1475
rect 30200 1467 30204 1475
rect 30224 1467 30228 1475
rect 30232 1467 30244 1475
rect 30248 1467 30260 1475
rect 30264 1467 30268 1475
rect 30288 1467 30292 1475
rect 30296 1467 30308 1475
rect 30316 1467 30332 1475
rect 30340 1467 30364 1475
rect 30380 1467 30396 1475
rect 30412 1467 30424 1475
rect 30436 1467 30440 1475
rect 30444 1467 30456 1475
rect 30460 1467 30464 1475
rect 30476 1467 30488 1475
rect 30500 1467 30504 1475
rect 30508 1467 30520 1475
rect 30536 1467 30584 1475
rect 30600 1467 30624 1475
rect 30632 1467 30648 1475
rect 30664 1467 30668 1475
rect 30672 1467 30676 1475
rect 30696 1467 30700 1475
rect 30704 1467 30716 1475
rect 30720 1467 30732 1475
rect 30736 1467 30740 1475
rect 30756 1467 30760 1475
rect 30764 1467 30768 1475
rect 30788 1467 30792 1475
rect 30796 1467 30808 1475
rect 30812 1467 30824 1475
rect 30828 1467 30832 1475
rect 30852 1467 30856 1475
rect 30860 1467 30872 1475
rect 30880 1467 30896 1475
rect 30904 1467 30928 1475
rect 30944 1467 30956 1475
rect 30976 1467 30988 1475
rect 31000 1467 31004 1475
rect 31008 1467 31020 1475
rect 31024 1467 31028 1475
rect 31156 1467 31160 1475
rect 31164 1467 31176 1475
rect 31180 1467 31184 1475
rect 31200 1467 31208 1475
rect 31228 1467 31240 1475
rect 31256 1467 31280 1475
rect 31288 1467 31304 1475
rect 31312 1467 31324 1475
rect 31328 1467 31332 1475
rect 31352 1467 31356 1475
rect 31360 1467 31372 1475
rect 31384 1467 31388 1475
rect 31392 1467 31396 1475
rect 31416 1467 31420 1475
rect 31424 1467 31436 1475
rect 31448 1467 31452 1475
rect 31456 1467 31460 1475
rect 31508 1467 31512 1475
rect 31516 1467 31528 1475
rect 31540 1467 31544 1475
rect 31548 1467 31552 1475
rect 31632 1467 31636 1475
rect 31640 1467 31644 1475
rect 31656 1467 31668 1475
rect 31672 1467 31676 1475
rect 31692 1467 31708 1475
rect 31724 1467 31740 1475
rect 31748 1467 31780 1475
rect 31788 1467 31804 1475
rect 31816 1467 31832 1475
rect 31840 1467 31872 1475
rect 31880 1467 31896 1475
rect 31912 1467 31924 1475
rect 31932 1467 31964 1475
rect 31972 1467 31988 1475
rect 32004 1467 32016 1475
rect 32028 1467 32032 1475
rect 32036 1467 32048 1475
rect 32068 1467 32080 1475
rect 32092 1467 32096 1475
rect 32100 1467 32112 1475
rect 32116 1467 32120 1475
rect 32132 1467 32144 1475
rect 32248 1467 32252 1475
rect 32256 1467 32268 1475
rect 32272 1467 32276 1475
rect 32288 1467 32300 1475
rect 32340 1467 32344 1475
rect 32348 1467 32360 1475
rect 32364 1467 32368 1475
rect 32380 1467 32392 1475
rect 32412 1467 32424 1475
rect 32440 1467 32464 1475
rect 32472 1467 32488 1475
rect 32496 1467 32528 1475
rect 32536 1467 32552 1475
rect 32568 1467 32584 1475
rect 32600 1467 32616 1475
rect 32632 1467 32648 1475
rect 32656 1467 32688 1475
rect 32696 1467 32708 1475
rect 32724 1467 32740 1475
rect 32748 1467 32780 1475
rect 32788 1467 32800 1475
rect 32812 1467 32836 1475
rect 32852 1467 32864 1475
rect 32884 1467 32896 1475
rect 32908 1467 32912 1475
rect 32916 1467 32928 1475
rect 32932 1467 32936 1475
rect 32948 1467 32960 1475
rect 33000 1467 33004 1475
rect 33008 1467 33020 1475
rect 33024 1467 33028 1475
rect 33132 1467 33144 1475
rect 33164 1467 33176 1475
rect 33180 1467 33192 1475
rect 33196 1467 33208 1475
rect 33224 1467 33240 1475
rect 33248 1467 33280 1475
rect 33288 1467 33304 1475
rect 33312 1467 33324 1475
rect 33328 1467 33332 1475
rect 33352 1467 33356 1475
rect 33360 1467 33372 1475
rect 33384 1467 33388 1475
rect 33392 1467 33396 1475
rect 33416 1467 33420 1475
rect 33424 1467 33428 1475
rect 33492 1467 33496 1475
rect 33500 1467 33504 1475
rect 33524 1467 33528 1475
rect 33532 1467 33536 1475
rect 33584 1467 33588 1475
rect 33592 1467 33596 1475
rect 33616 1467 33620 1475
rect 33624 1467 33636 1475
rect 33640 1467 33652 1475
rect 33656 1467 33660 1475
rect 33680 1467 33684 1475
rect 33688 1467 33692 1475
rect 33708 1467 33712 1475
rect 33716 1467 33728 1475
rect 33732 1467 33744 1475
rect 33748 1467 33752 1475
rect 33772 1467 33776 1475
rect 33780 1467 33792 1475
rect 33804 1467 33808 1475
rect 33812 1467 33816 1475
rect 33836 1467 33840 1475
rect 33844 1467 33856 1475
rect 33868 1467 33872 1475
rect 33876 1467 33880 1475
rect 33892 1467 33904 1475
rect 33908 1467 33912 1475
rect 34008 1467 34012 1475
rect 34016 1467 34020 1475
rect 34032 1467 34044 1475
rect 34048 1467 34060 1475
rect 34072 1467 34076 1475
rect 34080 1467 34084 1475
rect 34104 1467 34108 1475
rect 34112 1467 34116 1475
rect 34212 1467 34216 1475
rect 34220 1467 34224 1475
rect 34304 1467 34308 1475
rect 34312 1467 34316 1475
rect 34396 1467 34400 1475
rect 34404 1467 34408 1475
rect 34420 1467 34432 1475
rect 34436 1467 34448 1475
rect 34460 1467 34464 1475
rect 34468 1467 34472 1475
rect 34492 1467 34496 1475
rect 34500 1467 34504 1475
rect 34524 1467 34528 1475
rect 34532 1467 34536 1475
rect 34556 1467 34560 1475
rect 34564 1467 34568 1475
rect 34580 1467 34592 1475
rect 34596 1467 34608 1475
rect 34620 1467 34624 1475
rect 34628 1467 34632 1475
rect 34680 1467 34684 1475
rect 34688 1467 34700 1475
rect 34712 1467 34716 1475
rect 34720 1467 34724 1475
rect 34804 1467 34808 1475
rect 34812 1467 34816 1475
rect 34828 1467 34840 1475
rect 34844 1467 34848 1475
rect 34912 1467 34916 1475
rect 34920 1467 34924 1475
rect 34944 1467 34948 1475
rect 34952 1467 34956 1475
rect 34968 1467 34980 1475
rect 34984 1467 34996 1475
rect 35008 1467 35012 1475
rect 35016 1467 35020 1475
rect 35040 1467 35044 1475
rect 35048 1467 35060 1475
rect 35072 1467 35076 1475
rect 35080 1467 35084 1475
rect 35164 1467 35168 1475
rect 35172 1467 35176 1475
rect 35336 1467 35340 1475
rect 35344 1467 35348 1475
rect 35368 1467 35372 1475
rect 35376 1467 35380 1475
rect 35392 1467 35404 1475
rect 35408 1467 35412 1475
rect 35428 1467 35452 1475
rect 35460 1467 35476 1475
rect 35484 1467 35508 1475
rect 35524 1467 35528 1475
rect 35532 1467 35544 1475
rect 35552 1467 35568 1475
rect 35576 1467 35608 1475
rect 35616 1467 35632 1475
rect 35648 1467 35660 1475
rect 35672 1467 35676 1475
rect 35680 1467 35692 1475
rect 35712 1467 35724 1475
rect 35928 1467 35940 1475
rect 35944 1467 35948 1475
rect 35960 1467 35972 1475
rect 35992 1467 36000 1475
rect 36012 1467 36044 1475
rect 36052 1467 36068 1475
rect 36076 1467 36100 1475
rect 36116 1467 36120 1475
rect 36124 1467 36136 1475
rect 36144 1467 36160 1475
rect 36168 1467 36200 1475
rect 36208 1467 36224 1475
rect 36240 1467 36264 1475
rect 36272 1467 36288 1475
rect 36304 1467 36320 1475
rect 36328 1467 36352 1475
rect 36368 1467 36380 1475
rect 36400 1467 36412 1475
rect 36416 1467 36428 1475
rect 36432 1467 36444 1475
rect 36580 1467 36584 1475
rect 36588 1467 36600 1475
rect 36604 1467 36608 1475
rect 36620 1467 36632 1475
rect 36648 1467 36664 1475
rect 36680 1467 36704 1475
rect 36712 1467 36728 1475
rect 36736 1467 36748 1475
rect 36752 1467 36756 1475
rect 36772 1467 36796 1475
rect 36804 1467 36820 1475
rect 36828 1467 36860 1475
rect 36868 1467 36880 1475
rect 36900 1467 36912 1475
rect 36920 1467 36952 1475
rect 36960 1467 36972 1475
rect 36992 1467 37004 1475
rect 37012 1467 37044 1475
rect 37052 1467 37068 1475
rect 37076 1467 37100 1475
rect 37116 1467 37132 1475
rect 37148 1467 37164 1475
rect 37180 1467 37204 1475
rect 37212 1467 37228 1475
rect 37236 1467 37248 1475
rect 37252 1467 37256 1475
rect 37272 1467 37296 1475
rect 37304 1467 37320 1475
rect 37328 1467 37352 1475
rect 37364 1467 37388 1475
rect 37396 1467 37412 1475
rect 37420 1467 37452 1475
rect 37460 1467 37476 1475
rect 37492 1467 37504 1475
rect 37508 1467 37520 1475
rect 37524 1467 37536 1475
rect 37556 1467 37568 1475
rect 37712 1467 37724 1475
rect 37744 1467 37756 1475
rect 37760 1467 37772 1475
rect 37776 1467 37788 1475
rect 37808 1467 37820 1475
rect 37836 1467 37848 1475
rect 37852 1467 37864 1475
rect 37868 1467 37880 1475
rect 37928 1467 37940 1475
rect 37944 1467 37956 1475
rect 37960 1467 37972 1475
rect 37992 1467 38004 1475
rect 38108 1467 38112 1475
rect 38116 1467 38128 1475
rect 38132 1467 38136 1475
rect 38148 1467 38160 1475
rect 38172 1467 38176 1475
rect 38180 1467 38192 1475
rect 38212 1467 38224 1475
rect 38328 1467 38332 1475
rect 38336 1467 38348 1475
rect 38368 1467 38380 1475
rect 38384 1467 38396 1475
rect 38400 1467 38412 1475
rect 38432 1467 38444 1475
rect 38448 1467 38452 1475
rect 38464 1467 38476 1475
rect 38492 1467 38508 1475
rect 38524 1467 38572 1475
rect 38588 1467 38592 1475
rect 38596 1467 38600 1475
rect 38616 1467 38664 1475
rect 38680 1467 38684 1475
rect 38688 1467 38692 1475
rect 38708 1467 38756 1475
rect 38772 1467 38788 1475
rect 38804 1467 38816 1475
rect 38828 1467 38832 1475
rect 38836 1467 38848 1475
rect 38868 1467 38880 1475
rect 38884 1467 38888 1475
rect 38920 1467 38924 1475
rect 38928 1467 38940 1475
rect 39144 1467 39156 1475
rect 39160 1467 39164 1475
rect 39268 1467 39280 1475
rect 39284 1467 39288 1475
rect 39300 1467 39312 1475
rect 39324 1467 39328 1475
rect 39332 1467 39344 1475
rect 39364 1467 39376 1475
rect 39488 1467 39500 1475
rect 39520 1467 39532 1475
rect 39536 1467 39540 1475
rect 39552 1467 39564 1475
rect 39576 1467 39580 1475
rect 39584 1467 39596 1475
rect 39612 1467 39660 1475
rect 39676 1467 39692 1475
rect 39704 1467 39752 1475
rect 39768 1467 39784 1475
rect 39800 1467 39804 1475
rect 39808 1467 39820 1475
rect 39832 1467 39836 1475
rect 39840 1467 39844 1475
rect 39864 1467 39868 1475
rect 39872 1467 39876 1475
rect 39972 1467 39976 1475
rect 39980 1467 39984 1475
rect 40032 1467 40036 1475
rect 40040 1467 40052 1475
rect 40064 1467 40068 1475
rect 40072 1467 40076 1475
rect 40088 1467 40100 1475
rect 40104 1467 40108 1475
rect 40128 1467 40132 1475
rect 40136 1467 40140 1475
rect 40156 1467 40172 1475
rect 40180 1467 40212 1475
rect 40220 1467 40236 1475
rect 40252 1467 40264 1475
rect 40276 1467 40280 1475
rect 40284 1467 40296 1475
rect 40316 1467 40328 1475
rect 40440 1467 40452 1475
rect 40456 1467 40460 1475
rect 40472 1467 40484 1475
rect 40504 1467 40516 1475
rect 40520 1467 40532 1475
rect 40536 1467 40548 1475
rect 40568 1467 40580 1475
rect 40724 1467 40736 1475
rect 40756 1467 40768 1475
rect 40772 1467 40784 1475
rect 40788 1467 40800 1475
rect 19130 1450 19138 1458
rect 19280 1450 19286 1458
rect 19778 1450 19782 1458
rect 19868 1450 19876 1458
rect 19992 1450 19996 1458
rect 20082 1450 20090 1458
rect 20382 1450 20390 1458
rect 20532 1450 20538 1458
rect 21238 1450 21246 1458
rect 21388 1450 21394 1458
rect 21778 1450 21792 1458
rect 21832 1450 21840 1458
rect 21984 1450 21990 1458
rect 21992 1450 21998 1458
rect 22126 1450 22140 1458
rect 22348 1456 22352 1458
rect 22420 1450 22434 1458
rect 22474 1450 22488 1458
rect 22562 1456 22566 1458
rect 23062 1450 23076 1458
rect 23116 1450 23130 1458
rect 23204 1456 23208 1458
rect 23276 1450 23290 1458
rect 23330 1450 23344 1458
rect 23632 1456 23636 1458
rect 23704 1450 23718 1458
rect 23758 1450 23772 1458
rect 24140 1450 24142 1458
rect 24234 1450 24242 1458
rect 24572 1450 24574 1458
rect 24778 1450 24780 1458
rect 24992 1450 24994 1458
rect 25470 1450 25478 1458
rect 25684 1450 25692 1458
rect 26022 1450 26034 1458
rect 26236 1450 26248 1458
rect 26326 1450 26334 1458
rect 26540 1450 26548 1458
rect 26878 1450 26890 1458
rect 26968 1450 26976 1458
rect 27306 1450 27318 1458
rect 28060 1450 28064 1458
rect 36032 1457 36040 1465
rect 36800 1457 36808 1465
rect 2440 1439 2448 1447
rect 2488 1439 2496 1447
rect 3944 1439 3952 1447
rect 3960 1439 3968 1447
rect 6962 1433 6970 1441
rect 7122 1433 7130 1441
rect 7234 1433 7242 1441
rect 7346 1433 7354 1441
rect 7394 1433 7402 1441
rect 7410 1433 7418 1441
rect 7554 1433 7562 1441
rect 7570 1433 7578 1441
rect 8130 1433 8138 1441
rect 13738 1439 13746 1447
rect 13770 1439 13778 1447
rect 15258 1439 15266 1447
rect 16202 1439 16210 1447
rect 19296 1440 19304 1448
rect 19968 1440 19976 1448
rect 23536 1440 23544 1448
rect 29648 1437 29656 1445
rect 30528 1437 30536 1445
rect 30720 1437 30728 1445
rect 30960 1437 30968 1445
rect 31008 1437 31016 1445
rect 31088 1437 31096 1445
rect 32768 1437 32776 1445
rect 34704 1437 34712 1445
rect 35520 1437 35528 1445
rect 35824 1437 35832 1445
rect 36288 1437 36296 1445
rect 36576 1437 36584 1445
rect 40656 1437 40664 1445
rect 856 1419 864 1427
rect 984 1419 992 1427
rect 1256 1419 1264 1427
rect 1480 1419 1488 1427
rect 1720 1419 1728 1427
rect 1736 1419 1744 1427
rect 1864 1419 1872 1427
rect 1960 1419 1968 1427
rect 2552 1419 2560 1427
rect 2584 1419 2592 1427
rect 2728 1419 2736 1427
rect 2744 1419 2752 1427
rect 2760 1419 2768 1427
rect 2824 1419 2832 1427
rect 2920 1419 2928 1427
rect 2968 1419 2976 1427
rect 3224 1419 3232 1427
rect 3368 1419 3376 1427
rect 3416 1419 3424 1427
rect 3464 1419 3472 1427
rect 3512 1419 3520 1427
rect 3624 1419 3632 1427
rect 3640 1419 3648 1427
rect 3656 1419 3664 1427
rect 3752 1419 3760 1427
rect 4104 1419 4112 1427
rect 4264 1419 4272 1427
rect 4392 1419 4400 1427
rect 4456 1419 4464 1427
rect 5730 1413 5738 1421
rect 6098 1413 6106 1421
rect 6322 1413 6330 1421
rect 7266 1413 7274 1421
rect 7298 1413 7306 1421
rect 7362 1413 7370 1421
rect 8290 1413 8298 1421
rect 8322 1413 8330 1421
rect 9378 1413 9386 1421
rect 9458 1413 9466 1421
rect 12298 1419 12306 1427
rect 12762 1419 12770 1427
rect 13466 1419 13474 1427
rect 13642 1419 13650 1427
rect 15258 1419 15266 1427
rect 15370 1419 15378 1427
rect 15482 1419 15490 1427
rect 15514 1419 15522 1427
rect 16522 1419 16530 1427
rect 16906 1419 16914 1427
rect 17226 1419 17234 1427
rect 17338 1419 17346 1427
rect 17354 1419 17362 1427
rect 17434 1419 17442 1427
rect 18688 1420 18696 1428
rect 21840 1420 21848 1428
rect 22480 1420 22488 1428
rect 25024 1420 25032 1428
rect 26752 1420 26760 1428
rect 29504 1417 29512 1425
rect 30096 1417 30104 1425
rect 30240 1417 30248 1425
rect 30336 1417 30344 1425
rect 30384 1417 30392 1425
rect 30544 1417 30552 1425
rect 30592 1417 30600 1425
rect 31408 1417 31416 1425
rect 31488 1417 31496 1425
rect 31936 1417 31944 1425
rect 32304 1417 32312 1425
rect 32512 1417 32520 1425
rect 32752 1417 32760 1425
rect 33232 1417 33240 1425
rect 33392 1417 33400 1425
rect 33584 1417 33592 1425
rect 33824 1417 33832 1425
rect 34032 1417 34040 1425
rect 34208 1417 34216 1425
rect 35232 1417 35240 1425
rect 37616 1417 37624 1425
rect 38336 1417 38344 1425
rect 38384 1417 38392 1425
rect 38512 1417 38520 1425
rect 39024 1417 39032 1425
rect 40560 1417 40568 1425
rect 488 1399 496 1407
rect 520 1399 528 1407
rect 552 1399 560 1407
rect 776 1399 784 1407
rect 792 1399 800 1407
rect 808 1399 816 1407
rect 840 1399 848 1407
rect 872 1399 880 1407
rect 888 1399 896 1407
rect 904 1399 912 1407
rect 968 1399 976 1407
rect 1016 1399 1024 1407
rect 1144 1399 1152 1407
rect 1176 1399 1184 1407
rect 1432 1399 1440 1407
rect 1528 1399 1536 1407
rect 1640 1399 1648 1407
rect 1928 1399 1936 1407
rect 1976 1399 1984 1407
rect 1992 1399 2000 1407
rect 2008 1399 2016 1407
rect 2168 1399 2176 1407
rect 2232 1399 2240 1407
rect 2248 1399 2256 1407
rect 2408 1399 2416 1407
rect 2472 1399 2480 1407
rect 2616 1399 2624 1407
rect 2632 1399 2640 1407
rect 2680 1399 2688 1407
rect 2728 1399 2736 1407
rect 2760 1399 2768 1407
rect 2776 1399 2784 1407
rect 2952 1399 2960 1407
rect 3000 1399 3008 1407
rect 3288 1399 3296 1407
rect 3352 1399 3360 1407
rect 3368 1399 3376 1407
rect 3384 1399 3392 1407
rect 3480 1399 3488 1407
rect 3544 1399 3552 1407
rect 3640 1399 3648 1407
rect 3672 1399 3680 1407
rect 3752 1399 3760 1407
rect 3784 1399 3792 1407
rect 4088 1399 4096 1407
rect 4168 1399 4176 1407
rect 4184 1399 4192 1407
rect 4296 1399 4304 1407
rect 4488 1399 4496 1407
rect 4504 1399 4512 1407
rect 4536 1399 4544 1407
rect 4568 1399 4576 1407
rect 4616 1399 4624 1407
rect 6226 1393 6234 1401
rect 6242 1393 6250 1401
rect 6306 1393 6314 1401
rect 6338 1393 6346 1401
rect 6354 1393 6362 1401
rect 6514 1393 6522 1401
rect 6546 1393 6554 1401
rect 6594 1393 6602 1401
rect 6690 1393 6698 1401
rect 7346 1393 7354 1401
rect 7538 1393 7546 1401
rect 7618 1393 7626 1401
rect 7762 1393 7770 1401
rect 8050 1393 8058 1401
rect 8082 1393 8090 1401
rect 8386 1393 8394 1401
rect 8466 1393 8474 1401
rect 8498 1393 8506 1401
rect 8594 1393 8602 1401
rect 8626 1393 8634 1401
rect 8818 1393 8826 1401
rect 8914 1393 8922 1401
rect 9074 1393 9082 1401
rect 9442 1393 9450 1401
rect 9602 1393 9610 1401
rect 9650 1393 9658 1401
rect 9682 1393 9690 1401
rect 9858 1393 9866 1401
rect 9986 1393 9994 1401
rect 10018 1393 10026 1401
rect 10082 1393 10090 1401
rect 10162 1393 10170 1401
rect 10226 1393 10234 1401
rect 10322 1393 10330 1401
rect 10546 1393 10554 1401
rect 10690 1393 10698 1401
rect 12426 1399 12434 1407
rect 12490 1399 12498 1407
rect 13050 1399 13058 1407
rect 14074 1399 14082 1407
rect 15242 1399 15250 1407
rect 15322 1399 15330 1407
rect 15386 1399 15394 1407
rect 15866 1399 15874 1407
rect 15898 1399 15906 1407
rect 15962 1399 15970 1407
rect 15994 1399 16002 1407
rect 16938 1399 16946 1407
rect 17050 1399 17058 1407
rect 23584 1400 23592 1408
rect 25872 1400 25880 1408
rect 26368 1400 26376 1408
rect 28016 1400 28024 1408
rect 30480 1397 30488 1405
rect 33072 1397 33080 1405
rect 33104 1397 33112 1405
rect 33648 1397 33656 1405
rect 34800 1397 34808 1405
rect 35600 1397 35608 1405
rect 35856 1397 35864 1405
rect 36672 1397 36680 1405
rect 36768 1397 36776 1405
rect 38112 1397 38120 1405
rect 38560 1397 38568 1405
rect 40064 1397 40072 1405
rect 40384 1397 40392 1405
rect 40784 1397 40792 1405
rect 456 1379 464 1387
rect 776 1379 784 1387
rect 952 1379 960 1387
rect 1000 1379 1008 1387
rect 1160 1379 1168 1387
rect 1432 1379 1440 1387
rect 1816 1379 1824 1387
rect 2104 1379 2112 1387
rect 2216 1379 2224 1387
rect 2312 1379 2320 1387
rect 2600 1379 2608 1387
rect 2696 1379 2704 1387
rect 3288 1379 3296 1387
rect 4232 1379 4240 1387
rect 5794 1373 5802 1381
rect 6146 1373 6154 1381
rect 6210 1373 6218 1381
rect 6450 1373 6458 1381
rect 6690 1373 6698 1381
rect 6962 1373 6970 1381
rect 7010 1373 7018 1381
rect 8114 1373 8122 1381
rect 8130 1373 8138 1381
rect 8210 1373 8218 1381
rect 8322 1373 8330 1381
rect 8386 1373 8394 1381
rect 8482 1373 8490 1381
rect 8514 1373 8522 1381
rect 8690 1373 8698 1381
rect 8706 1373 8714 1381
rect 8946 1373 8954 1381
rect 9682 1373 9690 1381
rect 10098 1373 10106 1381
rect 10914 1373 10922 1381
rect 12202 1379 12210 1387
rect 12410 1379 12418 1387
rect 12442 1379 12450 1387
rect 12746 1379 12754 1387
rect 12810 1379 12818 1387
rect 13162 1379 13170 1387
rect 13274 1379 13282 1387
rect 14026 1379 14034 1387
rect 14618 1379 14626 1387
rect 14698 1379 14706 1387
rect 15402 1379 15410 1387
rect 15946 1379 15954 1387
rect 17482 1379 17490 1387
rect 18944 1380 18952 1388
rect 20848 1380 20856 1388
rect 21040 1380 21048 1388
rect 21056 1380 21064 1388
rect 21264 1380 21272 1388
rect 21440 1380 21448 1388
rect 21808 1380 21816 1388
rect 22112 1380 22120 1388
rect 22256 1380 22264 1388
rect 22384 1380 22392 1388
rect 22496 1380 22504 1388
rect 23392 1380 23400 1388
rect 23824 1380 23832 1388
rect 24656 1380 24664 1388
rect 24880 1380 24888 1388
rect 25504 1380 25512 1388
rect 26736 1380 26744 1388
rect 26896 1380 26904 1388
rect 27648 1380 27656 1388
rect 27840 1380 27848 1388
rect 29440 1377 29448 1385
rect 29824 1377 29832 1385
rect 30384 1377 30392 1385
rect 31232 1377 31240 1385
rect 31392 1377 31400 1385
rect 32064 1377 32072 1385
rect 37856 1377 37864 1385
rect 38000 1377 38008 1385
rect 38336 1377 38344 1385
rect 5810 1353 5818 1361
rect 5874 1353 5882 1361
rect 6050 1353 6058 1361
rect 6162 1353 6170 1361
rect 6306 1353 6314 1361
rect 6386 1353 6394 1361
rect 7186 1353 7194 1361
rect 7634 1353 7642 1361
rect 7986 1353 7994 1361
rect 9602 1353 9610 1361
rect 9746 1353 9754 1361
rect 9858 1353 9866 1361
rect 10578 1353 10586 1361
rect 10818 1353 10826 1361
rect 10834 1353 10842 1361
rect 14538 1359 14546 1367
rect 14602 1359 14610 1367
rect 15690 1359 15698 1367
rect 16266 1359 16274 1367
rect 19888 1360 19896 1368
rect 20416 1360 20424 1368
rect 29776 1357 29784 1365
rect 30688 1357 30696 1365
rect 31712 1357 31720 1365
rect 31872 1357 31880 1365
rect 32208 1357 32216 1365
rect 33664 1357 33672 1365
rect 33712 1357 33720 1365
rect 33888 1357 33896 1365
rect 34816 1357 34824 1365
rect 36384 1357 36392 1365
rect 36480 1357 36488 1365
rect 36896 1357 36904 1365
rect 37248 1357 37256 1365
rect 37328 1357 37336 1365
rect 37440 1357 37448 1365
rect 37792 1357 37800 1365
rect 37856 1357 37864 1365
rect 38208 1357 38216 1365
rect 38672 1357 38680 1365
rect 38976 1357 38984 1365
rect 39136 1357 39144 1365
rect 40048 1357 40056 1365
rect 40208 1357 40216 1365
rect 20126 1348 20130 1353
rect 21252 1348 21256 1353
rect 27339 1348 27346 1353
rect 1368 1339 1376 1347
rect 1416 1339 1424 1347
rect 1480 1339 1488 1347
rect 1800 1339 1808 1347
rect 2344 1339 2352 1347
rect 2424 1339 2432 1347
rect 2440 1339 2448 1347
rect 2952 1339 2960 1347
rect 3080 1339 3088 1347
rect 3208 1339 3216 1347
rect 3672 1339 3680 1347
rect 3880 1339 3888 1347
rect 4184 1339 4192 1347
rect 4200 1339 4208 1347
rect 4312 1339 4320 1347
rect 4360 1339 4368 1347
rect 4408 1339 4416 1347
rect 6002 1333 6010 1341
rect 7058 1333 7066 1341
rect 7106 1333 7114 1341
rect 7202 1333 7210 1341
rect 8162 1333 8170 1341
rect 8322 1333 8330 1341
rect 8706 1333 8714 1341
rect 8722 1333 8730 1341
rect 8930 1333 8938 1341
rect 9042 1333 9050 1341
rect 9090 1333 9098 1341
rect 9106 1333 9114 1341
rect 9154 1333 9162 1341
rect 9266 1333 9274 1341
rect 9698 1333 9706 1341
rect 10290 1333 10298 1341
rect 10418 1333 10426 1341
rect 10514 1333 10522 1341
rect 10594 1333 10602 1341
rect 10786 1333 10794 1341
rect 10818 1333 10826 1341
rect 12730 1339 12738 1347
rect 12922 1339 12930 1347
rect 13850 1339 13858 1347
rect 14026 1339 14034 1347
rect 14090 1339 14098 1347
rect 14154 1339 14162 1347
rect 14250 1339 14258 1347
rect 14634 1339 14642 1347
rect 14762 1339 14770 1347
rect 14890 1339 14898 1347
rect 14938 1339 14946 1347
rect 15098 1339 15106 1347
rect 16218 1339 16226 1347
rect 16490 1339 16498 1347
rect 16650 1339 16658 1347
rect 16730 1339 16738 1347
rect 17034 1339 17042 1347
rect 17178 1339 17186 1347
rect 17466 1339 17474 1347
rect 18512 1340 18520 1348
rect 18928 1340 18936 1348
rect 21808 1340 21816 1348
rect 23104 1340 23112 1348
rect 24368 1340 24376 1348
rect 24864 1340 24872 1348
rect 25072 1340 25080 1348
rect 25696 1340 25704 1348
rect 26992 1340 27000 1348
rect 28464 1340 28472 1348
rect 1992 1319 2000 1327
rect 9762 1313 9770 1321
rect 9794 1313 9802 1321
rect 10018 1313 10026 1321
rect 10178 1313 10186 1321
rect 10274 1313 10282 1321
rect 10530 1313 10538 1321
rect 10594 1313 10602 1321
rect 12442 1319 12450 1327
rect 13914 1319 13922 1327
rect 14218 1319 14226 1327
rect 14474 1319 14482 1327
rect 14586 1319 14594 1327
rect 14922 1319 14930 1327
rect 15146 1319 15154 1327
rect 15754 1319 15762 1327
rect 15882 1319 15890 1327
rect 16346 1319 16354 1327
rect 16954 1319 16962 1327
rect 25488 1320 25496 1328
rect 2664 1299 2672 1307
rect 3400 1299 3408 1307
rect 3576 1299 3584 1307
rect 6242 1293 6250 1301
rect 6498 1293 6506 1301
rect 6786 1293 6794 1301
rect 6850 1293 6858 1301
rect 7778 1293 7786 1301
rect 8594 1293 8602 1301
rect 9778 1293 9786 1301
rect 13578 1299 13586 1307
rect 26240 1300 26248 1308
rect 33744 1297 33752 1305
rect 35904 1297 35912 1305
rect 1192 1279 1200 1287
rect 1400 1279 1408 1287
rect 2024 1279 2032 1287
rect 2152 1279 2160 1287
rect 2392 1279 2400 1287
rect 2472 1279 2480 1287
rect 2648 1279 2656 1287
rect 2792 1279 2800 1287
rect 3272 1279 3280 1287
rect 3736 1279 3744 1287
rect 3768 1279 3776 1287
rect 4520 1279 4528 1287
rect 4552 1279 4560 1287
rect 6530 1273 6538 1281
rect 6914 1273 6922 1281
rect 7522 1273 7530 1281
rect 8114 1273 8122 1281
rect 8466 1273 8474 1281
rect 8754 1273 8762 1281
rect 9090 1273 9098 1281
rect 9234 1273 9242 1281
rect 9346 1273 9354 1281
rect 9586 1273 9594 1281
rect 9874 1273 9882 1281
rect 10242 1273 10250 1281
rect 10578 1273 10586 1281
rect 10722 1273 10730 1281
rect 13130 1279 13138 1287
rect 14362 1279 14370 1287
rect 15642 1279 15650 1287
rect 29396 1267 29408 1275
rect 29428 1267 29440 1275
rect 29444 1267 29448 1275
rect 29460 1267 29472 1275
rect 29488 1267 29504 1275
rect 29512 1267 29544 1275
rect 29552 1267 29568 1275
rect 29576 1267 29600 1275
rect 29616 1267 29620 1275
rect 29624 1267 29636 1275
rect 29644 1267 29660 1275
rect 29668 1267 29692 1275
rect 29708 1267 29712 1275
rect 29716 1267 29728 1275
rect 29732 1267 29744 1275
rect 29748 1267 29752 1275
rect 29772 1267 29776 1275
rect 29780 1267 29784 1275
rect 29800 1267 29804 1275
rect 29808 1267 29820 1275
rect 29824 1267 29836 1275
rect 29840 1267 29844 1275
rect 29892 1267 29896 1275
rect 29900 1267 29912 1275
rect 29916 1267 29928 1275
rect 29932 1267 29936 1275
rect 29956 1267 29960 1275
rect 29964 1267 29968 1275
rect 30032 1267 30036 1275
rect 30040 1267 30044 1275
rect 30064 1267 30068 1275
rect 30072 1267 30084 1275
rect 30088 1267 30100 1275
rect 30104 1267 30108 1275
rect 30128 1267 30132 1275
rect 30136 1267 30140 1275
rect 30152 1267 30164 1275
rect 30168 1267 30172 1275
rect 30192 1267 30196 1275
rect 30200 1267 30204 1275
rect 30220 1267 30268 1275
rect 30284 1267 30296 1275
rect 30300 1267 30304 1275
rect 30316 1267 30328 1275
rect 30340 1267 30344 1275
rect 30348 1267 30360 1275
rect 30536 1267 30548 1275
rect 30552 1267 30556 1275
rect 30568 1267 30580 1275
rect 30600 1267 30612 1275
rect 30616 1267 30620 1275
rect 30632 1267 30644 1275
rect 30652 1267 30676 1275
rect 30692 1267 30704 1275
rect 30708 1267 30712 1275
rect 30724 1267 30736 1275
rect 30744 1267 30768 1275
rect 30784 1267 30796 1275
rect 30800 1267 30804 1275
rect 30816 1267 30828 1275
rect 30840 1267 30844 1275
rect 30848 1267 30860 1275
rect 30864 1267 30868 1275
rect 30972 1267 30984 1275
rect 31004 1267 31016 1275
rect 31020 1267 31032 1275
rect 31036 1267 31048 1275
rect 31064 1267 31080 1275
rect 31088 1267 31120 1275
rect 31128 1267 31144 1275
rect 31152 1267 31184 1275
rect 31224 1267 31228 1275
rect 31232 1267 31236 1275
rect 31256 1267 31260 1275
rect 31264 1267 31276 1275
rect 31288 1267 31292 1275
rect 31296 1267 31300 1275
rect 31396 1267 31400 1275
rect 31404 1267 31408 1275
rect 31428 1267 31432 1275
rect 31436 1267 31440 1275
rect 31452 1267 31464 1275
rect 31468 1267 31480 1275
rect 31488 1267 31504 1275
rect 31520 1267 31524 1275
rect 31528 1267 31532 1275
rect 31544 1267 31556 1275
rect 31560 1267 31572 1275
rect 31580 1267 31596 1275
rect 31612 1267 31628 1275
rect 31636 1267 31648 1275
rect 31652 1267 31664 1275
rect 31676 1267 31680 1275
rect 31684 1267 31688 1275
rect 31704 1267 31708 1275
rect 31712 1267 31716 1275
rect 31728 1267 31740 1275
rect 31744 1267 31756 1275
rect 31768 1267 31772 1275
rect 31776 1267 31780 1275
rect 31796 1267 31812 1275
rect 31820 1267 31832 1275
rect 31836 1267 31848 1275
rect 31860 1267 31864 1275
rect 31868 1267 31872 1275
rect 31884 1267 31896 1275
rect 31900 1267 31904 1275
rect 31984 1267 31988 1275
rect 31992 1267 31996 1275
rect 32076 1267 32080 1275
rect 32084 1267 32096 1275
rect 32108 1267 32112 1275
rect 32116 1267 32120 1275
rect 32132 1267 32144 1275
rect 32148 1267 32152 1275
rect 32200 1267 32204 1275
rect 32208 1267 32212 1275
rect 32224 1267 32236 1275
rect 32240 1267 32244 1275
rect 32292 1267 32296 1275
rect 32300 1267 32304 1275
rect 32316 1267 32328 1275
rect 32332 1267 32336 1275
rect 32352 1267 32356 1275
rect 32360 1267 32372 1275
rect 32384 1267 32388 1275
rect 32392 1267 32396 1275
rect 32408 1267 32420 1275
rect 32424 1267 32428 1275
rect 32636 1267 32640 1275
rect 32644 1267 32648 1275
rect 32660 1267 32672 1275
rect 32676 1267 32688 1275
rect 32696 1267 32712 1275
rect 32728 1267 32732 1275
rect 32736 1267 32740 1275
rect 32752 1267 32764 1275
rect 32768 1267 32780 1275
rect 32792 1267 32796 1275
rect 32800 1267 32804 1275
rect 32824 1267 32828 1275
rect 32832 1267 32836 1275
rect 32856 1267 32860 1275
rect 32864 1267 32868 1275
rect 32888 1267 32892 1275
rect 32896 1267 32900 1275
rect 32912 1267 32924 1275
rect 32928 1267 32940 1275
rect 32952 1267 32956 1275
rect 32960 1267 32964 1275
rect 32980 1267 32996 1275
rect 33004 1267 33016 1275
rect 33020 1267 33032 1275
rect 33040 1267 33056 1275
rect 33072 1267 33088 1275
rect 33096 1267 33120 1275
rect 33136 1267 33152 1275
rect 33168 1267 33180 1275
rect 33184 1267 33196 1275
rect 33200 1267 33212 1275
rect 33316 1267 33320 1275
rect 33324 1267 33336 1275
rect 33356 1267 33368 1275
rect 33372 1267 33376 1275
rect 33388 1267 33400 1275
rect 33420 1267 33432 1275
rect 33448 1267 33496 1275
rect 33512 1267 33516 1275
rect 33520 1267 33524 1275
rect 33540 1267 33588 1275
rect 33604 1267 33620 1275
rect 33628 1267 33640 1275
rect 33644 1267 33656 1275
rect 33668 1267 33672 1275
rect 33676 1267 33680 1275
rect 33696 1267 33712 1275
rect 33720 1267 33732 1275
rect 33736 1267 33748 1275
rect 33760 1267 33764 1275
rect 33768 1267 33772 1275
rect 33784 1267 33796 1275
rect 33800 1267 33804 1275
rect 33824 1267 33828 1275
rect 33832 1267 33836 1275
rect 33848 1267 33860 1275
rect 33864 1267 33868 1275
rect 33888 1267 33892 1275
rect 33896 1267 33908 1275
rect 33916 1267 33932 1275
rect 33940 1267 33972 1275
rect 33980 1267 33996 1275
rect 34012 1267 34024 1275
rect 34028 1267 34040 1275
rect 34044 1267 34056 1275
rect 34072 1267 34088 1275
rect 34104 1267 34128 1275
rect 34136 1267 34152 1275
rect 34168 1267 34172 1275
rect 34176 1267 34180 1275
rect 34192 1267 34204 1275
rect 34208 1267 34220 1275
rect 34228 1267 34244 1275
rect 34260 1267 34264 1275
rect 34268 1267 34272 1275
rect 34284 1267 34296 1275
rect 34300 1267 34312 1275
rect 34320 1267 34336 1275
rect 34352 1267 34368 1275
rect 34376 1267 34388 1275
rect 34392 1267 34400 1275
rect 34416 1267 34420 1275
rect 34424 1267 34428 1275
rect 34524 1267 34528 1275
rect 34532 1267 34536 1275
rect 34556 1267 34560 1275
rect 34564 1267 34568 1275
rect 34580 1267 34592 1275
rect 34596 1267 34608 1275
rect 34616 1267 34632 1275
rect 34648 1267 34652 1275
rect 34656 1267 34660 1275
rect 34672 1267 34684 1275
rect 34688 1267 34700 1275
rect 34712 1267 34716 1275
rect 34720 1267 34724 1275
rect 34852 1267 34856 1275
rect 34860 1267 34864 1275
rect 34876 1267 34888 1275
rect 34892 1267 34896 1275
rect 34912 1267 34928 1275
rect 34944 1267 34960 1275
rect 34968 1267 35000 1275
rect 35008 1267 35024 1275
rect 35040 1267 35056 1275
rect 35072 1267 35076 1275
rect 35080 1267 35092 1275
rect 35104 1267 35108 1275
rect 35112 1267 35116 1275
rect 35128 1267 35140 1275
rect 35144 1267 35148 1275
rect 35164 1267 35180 1275
rect 35200 1267 35212 1275
rect 35220 1267 35252 1275
rect 35260 1267 35276 1275
rect 35284 1267 35316 1275
rect 35324 1267 35340 1275
rect 35356 1267 35360 1275
rect 35364 1267 35368 1275
rect 35388 1267 35392 1275
rect 35396 1267 35408 1275
rect 35420 1267 35424 1275
rect 35428 1267 35432 1275
rect 35444 1267 35456 1275
rect 35460 1267 35472 1275
rect 35484 1267 35488 1275
rect 35492 1267 35496 1275
rect 35512 1267 35560 1275
rect 35576 1267 35624 1275
rect 35640 1267 35656 1275
rect 35672 1267 35688 1275
rect 35704 1267 35720 1275
rect 35736 1267 35784 1275
rect 35800 1267 35804 1275
rect 35808 1267 35812 1275
rect 35828 1267 35876 1275
rect 35892 1267 35916 1275
rect 35924 1267 35940 1275
rect 35956 1267 35972 1275
rect 35988 1267 36000 1275
rect 36012 1267 36036 1275
rect 36052 1267 36100 1275
rect 36116 1267 36120 1275
rect 36124 1267 36128 1275
rect 36144 1267 36192 1275
rect 36208 1267 36232 1275
rect 36240 1267 36256 1275
rect 36272 1267 36276 1275
rect 36280 1267 36284 1275
rect 36304 1267 36308 1275
rect 36312 1267 36324 1275
rect 36328 1267 36340 1275
rect 36344 1267 36348 1275
rect 36364 1267 36368 1275
rect 36372 1267 36376 1275
rect 36396 1267 36400 1275
rect 36404 1267 36416 1275
rect 36420 1267 36432 1275
rect 36436 1267 36440 1275
rect 36456 1267 36460 1275
rect 36464 1267 36468 1275
rect 36488 1267 36492 1275
rect 36496 1267 36508 1275
rect 36512 1267 36524 1275
rect 36528 1267 36532 1275
rect 36580 1267 36584 1275
rect 36588 1267 36600 1275
rect 36604 1267 36616 1275
rect 36620 1267 36624 1275
rect 36640 1267 36664 1275
rect 36672 1267 36688 1275
rect 36696 1267 36720 1275
rect 36736 1267 36748 1275
rect 36768 1267 36780 1275
rect 36792 1267 36796 1275
rect 36800 1267 36812 1275
rect 36816 1267 36820 1275
rect 36832 1267 36844 1275
rect 36856 1267 36860 1275
rect 36864 1267 36876 1275
rect 36892 1267 36916 1275
rect 36924 1267 36936 1275
rect 36948 1267 36952 1275
rect 36956 1267 36968 1275
rect 36984 1267 37008 1275
rect 37016 1267 37028 1275
rect 37040 1267 37044 1275
rect 37048 1267 37060 1275
rect 37064 1267 37068 1275
rect 37080 1267 37092 1275
rect 37112 1267 37124 1275
rect 37144 1267 37156 1275
rect 37176 1267 37188 1275
rect 37200 1267 37204 1275
rect 37208 1267 37220 1275
rect 37224 1267 37228 1275
rect 37268 1267 37280 1275
rect 37292 1267 37296 1275
rect 37300 1267 37312 1275
rect 37316 1267 37320 1275
rect 37332 1267 37344 1275
rect 37488 1267 37500 1275
rect 37512 1267 37516 1275
rect 37520 1267 37532 1275
rect 37536 1267 37540 1275
rect 37552 1267 37564 1275
rect 37580 1267 37596 1275
rect 37612 1267 37636 1275
rect 37644 1267 37660 1275
rect 37668 1267 37680 1275
rect 37684 1267 37688 1275
rect 37704 1267 37728 1275
rect 37736 1267 37752 1275
rect 37760 1267 37792 1275
rect 37800 1267 37816 1275
rect 37832 1267 37844 1275
rect 37852 1267 37884 1275
rect 37892 1267 37908 1275
rect 37920 1267 37936 1275
rect 37944 1267 37976 1275
rect 37984 1267 38000 1275
rect 38016 1267 38032 1275
rect 38048 1267 38052 1275
rect 38056 1267 38068 1275
rect 38080 1267 38084 1275
rect 38088 1267 38092 1275
rect 38104 1267 38116 1275
rect 38120 1267 38132 1275
rect 38144 1267 38148 1275
rect 38152 1267 38156 1275
rect 38236 1267 38240 1275
rect 38244 1267 38248 1275
rect 38260 1267 38272 1275
rect 38276 1267 38280 1275
rect 38344 1267 38348 1275
rect 38352 1267 38356 1275
rect 38376 1267 38380 1275
rect 38384 1267 38396 1275
rect 38400 1267 38412 1275
rect 38416 1267 38420 1275
rect 38440 1267 38444 1275
rect 38448 1267 38452 1275
rect 38472 1267 38476 1275
rect 38480 1267 38484 1275
rect 38504 1267 38508 1275
rect 38512 1267 38516 1275
rect 38536 1267 38540 1275
rect 38544 1267 38556 1275
rect 38560 1267 38572 1275
rect 38576 1267 38580 1275
rect 38596 1267 38612 1275
rect 38628 1267 38632 1275
rect 38636 1267 38648 1275
rect 38652 1267 38664 1275
rect 38668 1267 38672 1275
rect 38688 1267 38704 1275
rect 38720 1267 38724 1275
rect 38728 1267 38740 1275
rect 38744 1267 38756 1275
rect 38760 1267 38764 1275
rect 38780 1267 38796 1275
rect 38812 1267 38816 1275
rect 38820 1267 38832 1275
rect 38836 1267 38848 1275
rect 38852 1267 38856 1275
rect 38876 1267 38880 1275
rect 38884 1267 38888 1275
rect 38936 1267 38940 1275
rect 38944 1267 38948 1275
rect 39028 1267 39032 1275
rect 39036 1267 39040 1275
rect 39120 1267 39124 1275
rect 39128 1267 39132 1275
rect 39152 1267 39156 1275
rect 39160 1267 39164 1275
rect 39244 1267 39248 1275
rect 39252 1267 39256 1275
rect 39336 1267 39340 1275
rect 39344 1267 39348 1275
rect 39360 1267 39372 1275
rect 39376 1267 39380 1275
rect 39400 1267 39404 1275
rect 39408 1267 39412 1275
rect 39424 1267 39436 1275
rect 39440 1267 39452 1275
rect 39460 1267 39476 1275
rect 39492 1267 39496 1275
rect 39500 1267 39504 1275
rect 39516 1267 39528 1275
rect 39532 1267 39544 1275
rect 39556 1267 39560 1275
rect 39564 1267 39568 1275
rect 39580 1267 39592 1275
rect 39596 1267 39600 1275
rect 39616 1267 39620 1275
rect 39624 1267 39636 1275
rect 39648 1267 39652 1275
rect 39656 1267 39660 1275
rect 39672 1267 39684 1275
rect 39688 1267 39692 1275
rect 39740 1267 39744 1275
rect 39748 1267 39752 1275
rect 39764 1267 39776 1275
rect 39780 1267 39784 1275
rect 39880 1267 39884 1275
rect 39888 1267 39892 1275
rect 39904 1267 39916 1275
rect 39920 1267 39924 1275
rect 39944 1267 39948 1275
rect 39952 1267 39956 1275
rect 39972 1267 40020 1275
rect 40036 1267 40048 1275
rect 40064 1267 40112 1275
rect 40128 1267 40144 1275
rect 40156 1267 40204 1275
rect 40220 1267 40224 1275
rect 40228 1267 40232 1275
rect 40248 1267 40296 1275
rect 40312 1267 40328 1275
rect 40344 1267 40356 1275
rect 40368 1267 40372 1275
rect 40376 1267 40388 1275
rect 40408 1267 40420 1275
rect 40424 1267 40428 1275
rect 40460 1267 40464 1275
rect 40468 1267 40480 1275
rect 40500 1267 40512 1275
rect 40516 1267 40528 1275
rect 40532 1267 40544 1275
rect 40560 1267 40576 1275
rect 40592 1267 40616 1275
rect 40624 1267 40640 1275
rect 40656 1267 40672 1275
rect 40680 1267 40692 1275
rect 40696 1267 40708 1275
rect 40716 1267 40732 1275
rect 40748 1267 40796 1275
rect 3636 1263 3660 1267
rect 4056 1259 4064 1267
rect 6578 1253 6586 1261
rect 7666 1253 7674 1261
rect 7682 1253 7690 1261
rect 7858 1253 7866 1261
rect 7890 1253 7898 1261
rect 8018 1253 8026 1261
rect 8114 1253 8122 1261
rect 8466 1253 8474 1261
rect 8514 1253 8522 1261
rect 9426 1253 9434 1261
rect 9506 1253 9514 1261
rect 16458 1259 16466 1267
rect 18472 1248 18476 1260
rect 18570 1250 18572 1258
rect 18578 1250 18580 1258
rect 18990 1250 19000 1258
rect 19204 1250 19214 1258
rect 21534 1250 21536 1258
rect 21542 1250 21544 1258
rect 21962 1250 21964 1258
rect 21970 1250 21972 1258
rect 22390 1250 22392 1258
rect 22398 1250 22400 1258
rect 24926 1250 24928 1258
rect 24934 1250 24936 1258
rect 25140 1250 25142 1258
rect 25148 1250 25150 1258
rect 28120 1250 28122 1258
rect 28128 1250 28130 1258
rect 36272 1257 36280 1265
rect 39280 1257 39288 1265
rect 39296 1257 39304 1265
rect 9554 1233 9562 1241
rect 12938 1239 12946 1247
rect 13066 1239 13074 1247
rect 13834 1239 13842 1247
rect 19536 1240 19544 1248
rect 20608 1240 20616 1248
rect 36224 1237 36232 1245
rect 39760 1237 39768 1245
rect 424 1219 432 1227
rect 632 1219 640 1227
rect 1192 1219 1200 1227
rect 1336 1219 1344 1227
rect 1400 1219 1408 1227
rect 1576 1219 1584 1227
rect 1592 1219 1600 1227
rect 1704 1219 1712 1227
rect 2168 1219 2176 1227
rect 2568 1219 2576 1227
rect 2728 1219 2736 1227
rect 2776 1219 2784 1227
rect 2984 1219 2992 1227
rect 3224 1219 3232 1227
rect 3304 1219 3312 1227
rect 3800 1219 3808 1227
rect 3944 1219 3952 1227
rect 4136 1219 4144 1227
rect 4168 1219 4176 1227
rect 4200 1219 4208 1227
rect 4440 1219 4448 1227
rect 4664 1219 4672 1227
rect 6418 1213 6426 1221
rect 6626 1213 6634 1221
rect 6754 1213 6762 1221
rect 7218 1213 7226 1221
rect 7538 1213 7546 1221
rect 7618 1213 7626 1221
rect 8754 1213 8762 1221
rect 8882 1213 8890 1221
rect 9346 1213 9354 1221
rect 10258 1213 10266 1221
rect 10818 1213 10826 1221
rect 12762 1219 12770 1227
rect 13658 1219 13666 1227
rect 14234 1219 14242 1227
rect 14426 1219 14434 1227
rect 15114 1219 15122 1227
rect 15882 1219 15890 1227
rect 30080 1217 30088 1225
rect 31024 1217 31032 1225
rect 32720 1217 32728 1225
rect 34416 1217 34424 1225
rect 35312 1217 35320 1225
rect 36992 1217 37000 1225
rect 37232 1217 37240 1225
rect 39520 1217 39528 1225
rect 39632 1217 39640 1225
rect 2008 1199 2016 1207
rect 2328 1199 2336 1207
rect 2504 1199 2512 1207
rect 3864 1199 3872 1207
rect 4264 1199 4272 1207
rect 4600 1199 4608 1207
rect 5746 1193 5754 1201
rect 6978 1193 6986 1201
rect 7586 1193 7594 1201
rect 9506 1193 9514 1201
rect 9698 1193 9706 1201
rect 9714 1193 9722 1201
rect 9938 1193 9946 1201
rect 10162 1193 10170 1201
rect 12234 1199 12242 1207
rect 13594 1199 13602 1207
rect 14346 1199 14354 1207
rect 16410 1199 16418 1207
rect 16570 1199 16578 1207
rect 16858 1199 16866 1207
rect 20144 1200 20152 1208
rect 21056 1200 21064 1208
rect 30656 1197 30664 1205
rect 37600 1197 37608 1205
rect 808 1179 816 1187
rect 1064 1179 1072 1187
rect 1128 1179 1136 1187
rect 1416 1179 1424 1187
rect 2072 1179 2080 1187
rect 2216 1179 2224 1187
rect 2424 1179 2432 1187
rect 2552 1179 2560 1187
rect 2808 1179 2816 1187
rect 4456 1179 4464 1187
rect 6978 1173 6986 1181
rect 7234 1173 7242 1181
rect 7634 1173 7642 1181
rect 8642 1173 8650 1181
rect 9154 1173 9162 1181
rect 9346 1173 9354 1181
rect 10322 1173 10330 1181
rect 10450 1173 10458 1181
rect 10834 1173 10842 1181
rect 12506 1179 12514 1187
rect 12602 1179 12610 1187
rect 14874 1179 14882 1187
rect 15962 1179 15970 1187
rect 17034 1179 17042 1187
rect 17290 1179 17298 1187
rect 29408 1177 29416 1185
rect 29568 1177 29576 1185
rect 29872 1177 29880 1185
rect 30400 1177 30408 1185
rect 30896 1177 30904 1185
rect 31664 1177 31672 1185
rect 32000 1177 32008 1185
rect 32608 1177 32616 1185
rect 34080 1177 34088 1185
rect 34448 1177 34456 1185
rect 35840 1177 35848 1185
rect 36464 1177 36472 1185
rect 36848 1177 36856 1185
rect 36944 1177 36952 1185
rect 37008 1177 37016 1185
rect 37680 1177 37688 1185
rect 37824 1177 37832 1185
rect 38176 1177 38184 1185
rect 38656 1177 38664 1185
rect 40112 1177 40120 1185
rect 40224 1177 40232 1185
rect 648 1159 656 1167
rect 744 1159 752 1167
rect 1512 1159 1520 1167
rect 1688 1159 1696 1167
rect 1736 1159 1744 1167
rect 2232 1159 2240 1167
rect 3048 1159 3056 1167
rect 3176 1159 3184 1167
rect 3208 1159 3216 1167
rect 3288 1159 3296 1167
rect 3352 1159 3360 1167
rect 3400 1159 3408 1167
rect 3496 1159 3504 1167
rect 3544 1159 3552 1167
rect 3592 1159 3600 1167
rect 3816 1159 3824 1167
rect 3848 1159 3856 1167
rect 4408 1159 4416 1167
rect 4632 1159 4640 1167
rect 6178 1153 6186 1161
rect 6194 1153 6202 1161
rect 6290 1153 6298 1161
rect 6482 1153 6490 1161
rect 6834 1153 6842 1161
rect 6882 1153 6890 1161
rect 7074 1153 7082 1161
rect 7474 1153 7482 1161
rect 7826 1153 7834 1161
rect 7842 1153 7850 1161
rect 8306 1153 8314 1161
rect 8578 1153 8586 1161
rect 8930 1153 8938 1161
rect 10018 1153 10026 1161
rect 10514 1153 10522 1161
rect 12250 1159 12258 1167
rect 13098 1159 13106 1167
rect 13178 1159 13186 1167
rect 13722 1159 13730 1167
rect 13770 1159 13778 1167
rect 13786 1159 13794 1167
rect 13930 1159 13938 1167
rect 14026 1159 14034 1167
rect 14314 1159 14322 1167
rect 14602 1159 14610 1167
rect 15002 1159 15010 1167
rect 15242 1159 15250 1167
rect 15290 1159 15298 1167
rect 15562 1159 15570 1167
rect 15786 1159 15794 1167
rect 15946 1159 15954 1167
rect 16074 1159 16082 1167
rect 16122 1159 16130 1167
rect 16346 1159 16354 1167
rect 16570 1159 16578 1167
rect 16634 1159 16642 1167
rect 16746 1159 16754 1167
rect 16794 1159 16802 1167
rect 16890 1159 16898 1167
rect 16954 1159 16962 1167
rect 18704 1160 18712 1168
rect 19040 1160 19048 1168
rect 19698 1161 19708 1166
rect 19904 1160 19912 1168
rect 20976 1160 20984 1168
rect 21040 1160 21048 1168
rect 21248 1160 21256 1168
rect 21472 1160 21480 1168
rect 21808 1160 21816 1168
rect 21904 1160 21912 1168
rect 22528 1160 22536 1168
rect 23088 1160 23096 1168
rect 23360 1160 23368 1168
rect 23792 1160 23800 1168
rect 24000 1160 24008 1168
rect 24992 1160 25000 1168
rect 25184 1160 25192 1168
rect 25201 1161 25206 1166
rect 25424 1160 25432 1168
rect 25696 1160 25704 1168
rect 26304 1160 26312 1168
rect 27776 1160 27784 1168
rect 28480 1160 28488 1168
rect 1016 1139 1024 1147
rect 1064 1139 1072 1147
rect 3368 1139 3376 1147
rect 6338 1133 6346 1141
rect 6434 1133 6442 1141
rect 6514 1133 6522 1141
rect 7458 1133 7466 1141
rect 7794 1133 7802 1141
rect 7890 1133 7898 1141
rect 7938 1133 7946 1141
rect 7954 1133 7962 1141
rect 8066 1133 8074 1141
rect 8114 1133 8122 1141
rect 8450 1133 8458 1141
rect 8802 1133 8810 1141
rect 8978 1133 8986 1141
rect 9250 1133 9258 1141
rect 9490 1133 9498 1141
rect 9730 1133 9738 1141
rect 9922 1133 9930 1141
rect 10082 1133 10090 1141
rect 10162 1133 10170 1141
rect 10226 1133 10234 1141
rect 10706 1133 10714 1141
rect 10866 1133 10874 1141
rect 14794 1139 14802 1147
rect 16138 1139 16146 1147
rect 16218 1139 16226 1147
rect 16842 1139 16850 1147
rect 16986 1139 16994 1147
rect 17162 1139 17170 1147
rect 17226 1139 17234 1147
rect 17242 1139 17250 1147
rect 17274 1139 17282 1147
rect 17418 1139 17426 1147
rect 18832 1140 18840 1148
rect 23648 1140 23656 1148
rect 24016 1140 24024 1148
rect 27376 1140 27384 1148
rect 28640 1140 28648 1148
rect 29552 1137 29560 1145
rect 29920 1137 29928 1145
rect 30416 1137 30424 1145
rect 30720 1137 30728 1145
rect 31344 1137 31352 1145
rect 31376 1137 31384 1145
rect 31440 1137 31448 1145
rect 31744 1137 31752 1145
rect 32112 1137 32120 1145
rect 32416 1137 32424 1145
rect 32592 1137 32600 1145
rect 33072 1137 33080 1145
rect 33664 1137 33672 1145
rect 33792 1137 33800 1145
rect 34464 1137 34472 1145
rect 34592 1137 34600 1145
rect 34768 1137 34776 1145
rect 35008 1137 35016 1145
rect 35376 1137 35384 1145
rect 36720 1137 36728 1145
rect 37616 1137 37624 1145
rect 37952 1137 37960 1145
rect 38240 1137 38248 1145
rect 38976 1137 38984 1145
rect 39744 1137 39752 1145
rect 40352 1137 40360 1145
rect 40624 1137 40632 1145
rect 488 1119 496 1127
rect 696 1119 704 1127
rect 728 1119 736 1127
rect 776 1119 784 1127
rect 1144 1119 1152 1127
rect 1224 1119 1232 1127
rect 1544 1119 1552 1127
rect 2072 1119 2080 1127
rect 2264 1119 2272 1127
rect 2376 1119 2384 1127
rect 3032 1119 3040 1127
rect 3080 1119 3088 1127
rect 3240 1119 3248 1127
rect 3496 1119 3504 1127
rect 4088 1119 4096 1127
rect 4232 1119 4240 1127
rect 4248 1119 4256 1127
rect 4424 1119 4432 1127
rect 4520 1119 4528 1127
rect 5794 1113 5802 1121
rect 6338 1113 6346 1121
rect 6866 1113 6874 1121
rect 6898 1113 6906 1121
rect 7170 1113 7178 1121
rect 7394 1113 7402 1121
rect 8178 1113 8186 1121
rect 8866 1113 8874 1121
rect 10322 1113 10330 1121
rect 10354 1113 10362 1121
rect 10482 1113 10490 1121
rect 12010 1119 12018 1127
rect 12746 1119 12754 1127
rect 13194 1119 13202 1127
rect 13626 1119 13634 1127
rect 14794 1119 14802 1127
rect 15034 1119 15042 1127
rect 15258 1119 15266 1127
rect 15354 1119 15362 1127
rect 16394 1119 16402 1127
rect 16474 1119 16482 1127
rect 17178 1119 17186 1127
rect 17450 1119 17458 1127
rect 19248 1120 19256 1128
rect 19344 1120 19352 1128
rect 19984 1120 19992 1128
rect 20320 1120 20328 1128
rect 21488 1120 21496 1128
rect 22240 1120 22248 1128
rect 22848 1120 22856 1128
rect 23808 1120 23816 1128
rect 26144 1120 26152 1128
rect 26336 1120 26344 1128
rect 26576 1120 26584 1128
rect 26784 1120 26792 1128
rect 27216 1120 27224 1128
rect 27760 1120 27768 1128
rect 28256 1120 28264 1128
rect 28288 1120 28296 1128
rect 33648 1117 33656 1125
rect 34032 1117 34040 1125
rect 39872 1117 39880 1125
rect 40064 1117 40072 1125
rect 40384 1117 40392 1125
rect 440 1099 448 1107
rect 504 1099 512 1107
rect 552 1099 560 1107
rect 600 1099 608 1107
rect 616 1099 624 1107
rect 792 1099 800 1107
rect 936 1099 944 1107
rect 1032 1099 1040 1107
rect 1208 1099 1216 1107
rect 1320 1099 1328 1107
rect 1416 1099 1424 1107
rect 1560 1099 1568 1107
rect 1608 1099 1616 1107
rect 1624 1099 1632 1107
rect 1656 1099 1664 1107
rect 1672 1099 1680 1107
rect 1880 1099 1888 1107
rect 1912 1099 1920 1107
rect 1928 1099 1936 1107
rect 2008 1099 2016 1107
rect 2136 1099 2144 1107
rect 2184 1099 2192 1107
rect 2200 1099 2208 1107
rect 2280 1099 2288 1107
rect 2344 1099 2352 1107
rect 2520 1099 2528 1107
rect 2536 1099 2544 1107
rect 2648 1099 2656 1107
rect 2760 1099 2768 1107
rect 2888 1099 2896 1107
rect 2984 1099 2992 1107
rect 3000 1099 3008 1107
rect 3064 1099 3072 1107
rect 3096 1099 3104 1107
rect 3240 1099 3248 1107
rect 3336 1099 3344 1107
rect 3480 1099 3488 1107
rect 3512 1099 3520 1107
rect 3608 1099 3616 1107
rect 3624 1099 3632 1107
rect 3704 1099 3712 1107
rect 3880 1099 3888 1107
rect 3960 1099 3968 1107
rect 4184 1099 4192 1107
rect 4216 1099 4224 1107
rect 4424 1099 4432 1107
rect 4488 1099 4496 1107
rect 4568 1099 4576 1107
rect 4648 1099 4656 1107
rect 6002 1093 6010 1101
rect 6082 1093 6090 1101
rect 6098 1093 6106 1101
rect 6642 1093 6650 1101
rect 6770 1093 6778 1101
rect 7106 1093 7114 1101
rect 7234 1093 7242 1101
rect 7298 1093 7306 1101
rect 7570 1093 7578 1101
rect 7602 1093 7610 1101
rect 7698 1093 7706 1101
rect 7794 1093 7802 1101
rect 7906 1093 7914 1101
rect 7970 1093 7978 1101
rect 8578 1093 8586 1101
rect 8674 1093 8682 1101
rect 8802 1093 8810 1101
rect 8850 1093 8858 1101
rect 8866 1093 8874 1101
rect 8898 1093 8906 1101
rect 9330 1093 9338 1101
rect 9474 1093 9482 1101
rect 9522 1093 9530 1101
rect 10754 1093 10762 1101
rect 10898 1093 10906 1101
rect 12922 1099 12930 1107
rect 13466 1099 13474 1107
rect 13642 1099 13650 1107
rect 14170 1099 14178 1107
rect 14986 1099 14994 1107
rect 15898 1099 15906 1107
rect 19520 1100 19528 1108
rect 22928 1100 22936 1108
rect 24080 1100 24088 1108
rect 24160 1100 24168 1108
rect 24416 1100 24424 1108
rect 24640 1100 24648 1108
rect 25952 1100 25960 1108
rect 27984 1100 27992 1108
rect 31264 1097 31272 1105
rect 31456 1097 31464 1105
rect 32048 1097 32056 1105
rect 32640 1097 32648 1105
rect 32656 1097 32664 1105
rect 33168 1097 33176 1105
rect 33824 1097 33832 1105
rect 35056 1097 35064 1105
rect 36032 1097 36040 1105
rect 36880 1097 36888 1105
rect 37072 1097 37080 1105
rect 37120 1097 37128 1105
rect 37440 1097 37448 1105
rect 38288 1097 38296 1105
rect 38560 1097 38568 1105
rect 38640 1097 38648 1105
rect 38912 1097 38920 1105
rect 39920 1097 39928 1105
rect 504 1079 512 1087
rect 840 1079 848 1087
rect 1128 1079 1136 1087
rect 1192 1079 1200 1087
rect 1208 1079 1216 1087
rect 1256 1079 1264 1087
rect 1368 1079 1376 1087
rect 1384 1079 1392 1087
rect 2488 1079 2496 1087
rect 3128 1079 3136 1087
rect 3560 1079 3568 1087
rect 3720 1079 3728 1087
rect 3896 1079 3904 1087
rect 3992 1079 4000 1087
rect 4408 1079 4416 1087
rect 4584 1079 4592 1087
rect 7314 1073 7322 1081
rect 7922 1073 7930 1081
rect 8418 1073 8426 1081
rect 8594 1073 8602 1081
rect 9042 1073 9050 1081
rect 9586 1073 9594 1081
rect 10914 1073 10922 1081
rect 12042 1079 12050 1087
rect 12762 1079 12770 1087
rect 13210 1079 13218 1087
rect 13530 1079 13538 1087
rect 13850 1079 13858 1087
rect 14682 1079 14690 1087
rect 16346 1079 16354 1087
rect 16922 1079 16930 1087
rect 17050 1079 17058 1087
rect 17130 1079 17138 1087
rect 20592 1080 20600 1088
rect 22080 1080 22088 1088
rect 23968 1080 23976 1088
rect 25264 1080 25272 1088
rect 27792 1080 27800 1088
rect 28448 1080 28456 1088
rect 30864 1077 30872 1085
rect 31504 1077 31512 1085
rect 32448 1077 32456 1085
rect 32640 1077 32648 1085
rect 33008 1077 33016 1085
rect 33024 1077 33032 1085
rect 33632 1077 33640 1085
rect 35520 1077 35528 1085
rect 35584 1077 35592 1085
rect 36240 1077 36248 1085
rect 36864 1077 36872 1085
rect 2056 1059 2064 1067
rect 6866 1053 6874 1061
rect 7650 1053 7658 1061
rect 8594 1053 8602 1061
rect 8722 1053 8730 1061
rect 9202 1053 9210 1061
rect 10354 1053 10362 1061
rect 10770 1053 10778 1061
rect 12618 1059 12626 1067
rect 12698 1059 12706 1067
rect 12826 1059 12834 1067
rect 13802 1059 13810 1067
rect 16074 1059 16082 1067
rect 22704 1060 22712 1068
rect 22912 1060 22920 1068
rect 29396 1067 29408 1075
rect 29428 1067 29440 1075
rect 29444 1067 29448 1075
rect 29460 1067 29472 1075
rect 29488 1067 29504 1075
rect 29512 1067 29544 1075
rect 29552 1067 29568 1075
rect 29576 1067 29600 1075
rect 29612 1067 29636 1075
rect 29644 1067 29660 1075
rect 29668 1067 29692 1075
rect 29708 1067 29712 1075
rect 29716 1067 29728 1075
rect 29740 1067 29744 1075
rect 29748 1067 29752 1075
rect 29772 1067 29776 1075
rect 29780 1067 29784 1075
rect 29848 1067 29852 1075
rect 29856 1067 29860 1075
rect 29880 1067 29884 1075
rect 29888 1067 29900 1075
rect 29904 1067 29916 1075
rect 29920 1067 29924 1075
rect 29944 1067 29948 1075
rect 29952 1067 29964 1075
rect 29972 1067 29988 1075
rect 29996 1067 30020 1075
rect 30036 1067 30048 1075
rect 30068 1067 30080 1075
rect 30092 1067 30096 1075
rect 30100 1067 30112 1075
rect 30116 1067 30120 1075
rect 30132 1067 30144 1075
rect 30152 1067 30176 1075
rect 30192 1067 30216 1075
rect 30224 1067 30236 1075
rect 30248 1067 30252 1075
rect 30256 1067 30268 1075
rect 30372 1067 30376 1075
rect 30380 1067 30392 1075
rect 30412 1067 30424 1075
rect 30428 1067 30432 1075
rect 30444 1067 30456 1075
rect 30476 1067 30488 1075
rect 30492 1067 30496 1075
rect 30508 1067 30520 1075
rect 30532 1067 30536 1075
rect 30540 1067 30552 1075
rect 30572 1067 30584 1075
rect 30596 1067 30600 1075
rect 30604 1067 30616 1075
rect 30636 1067 30648 1075
rect 30652 1067 30656 1075
rect 30668 1067 30680 1075
rect 30696 1067 30712 1075
rect 30728 1067 30776 1075
rect 30788 1067 30804 1075
rect 30820 1067 30868 1075
rect 30884 1067 30888 1075
rect 30892 1067 30896 1075
rect 30908 1067 30920 1075
rect 30924 1067 30936 1075
rect 30948 1067 30952 1075
rect 30956 1067 30960 1075
rect 30976 1067 30980 1075
rect 30984 1067 30988 1075
rect 31000 1067 31012 1075
rect 31016 1067 31028 1075
rect 31040 1067 31044 1075
rect 31048 1067 31052 1075
rect 31212 1067 31216 1075
rect 31220 1067 31224 1075
rect 31244 1067 31248 1075
rect 31252 1067 31256 1075
rect 31268 1067 31280 1075
rect 31284 1067 31288 1075
rect 31304 1067 31328 1075
rect 31336 1067 31352 1075
rect 31360 1067 31372 1075
rect 31376 1067 31380 1075
rect 31396 1067 31420 1075
rect 31428 1067 31444 1075
rect 31452 1067 31464 1075
rect 31468 1067 31472 1075
rect 31488 1067 31512 1075
rect 31520 1067 31536 1075
rect 31544 1067 31568 1075
rect 31584 1067 31596 1075
rect 31616 1067 31628 1075
rect 31640 1067 31644 1075
rect 31648 1067 31660 1075
rect 31664 1067 31668 1075
rect 31680 1067 31692 1075
rect 31732 1067 31736 1075
rect 31740 1067 31752 1075
rect 31756 1067 31760 1075
rect 31772 1067 31784 1075
rect 32208 1067 32220 1075
rect 32224 1067 32228 1075
rect 32240 1067 32252 1075
rect 32272 1067 32284 1075
rect 32300 1067 32348 1075
rect 32364 1067 32368 1075
rect 32372 1067 32376 1075
rect 32392 1067 32440 1075
rect 32456 1067 32472 1075
rect 32480 1067 32504 1075
rect 32520 1067 32536 1075
rect 32552 1067 32564 1075
rect 32568 1067 32580 1075
rect 32584 1067 32596 1075
rect 32616 1067 32628 1075
rect 32644 1067 32668 1075
rect 32676 1067 32692 1075
rect 32708 1067 32712 1075
rect 32716 1067 32720 1075
rect 32732 1067 32744 1075
rect 32748 1067 32760 1075
rect 32772 1067 32776 1075
rect 32780 1067 32784 1075
rect 32800 1067 32808 1075
rect 32812 1067 32816 1075
rect 32836 1067 32840 1075
rect 32844 1067 32848 1075
rect 32868 1067 32872 1075
rect 32876 1067 32880 1075
rect 32900 1067 32904 1075
rect 32908 1067 32920 1075
rect 32932 1067 32936 1075
rect 32940 1067 32944 1075
rect 32956 1067 32968 1075
rect 32972 1067 32976 1075
rect 32992 1067 32996 1075
rect 33000 1067 33012 1075
rect 33024 1067 33028 1075
rect 33032 1067 33036 1075
rect 33148 1067 33152 1075
rect 33156 1067 33160 1075
rect 33224 1067 33228 1075
rect 33232 1067 33236 1075
rect 33256 1067 33260 1075
rect 33264 1067 33268 1075
rect 33316 1067 33320 1075
rect 33324 1067 33328 1075
rect 33348 1067 33352 1075
rect 33356 1067 33360 1075
rect 33372 1067 33384 1075
rect 33388 1067 33392 1075
rect 33412 1067 33416 1075
rect 33420 1067 33424 1075
rect 33440 1067 33488 1075
rect 33504 1067 33516 1075
rect 33532 1067 33580 1075
rect 33600 1067 33612 1075
rect 33628 1067 33640 1075
rect 33652 1067 33656 1075
rect 33660 1067 33672 1075
rect 33692 1067 33704 1075
rect 33708 1067 33712 1075
rect 33944 1067 33956 1075
rect 33960 1067 33972 1075
rect 33976 1067 33988 1075
rect 34008 1067 34020 1075
rect 34028 1067 34060 1075
rect 34068 1067 34080 1075
rect 34100 1067 34112 1075
rect 34124 1067 34128 1075
rect 34132 1067 34144 1075
rect 34256 1067 34268 1075
rect 34280 1067 34284 1075
rect 34288 1067 34300 1075
rect 34304 1067 34308 1075
rect 34320 1067 34332 1075
rect 34372 1067 34376 1075
rect 34380 1067 34392 1075
rect 34396 1067 34400 1075
rect 34412 1067 34424 1075
rect 34440 1067 34452 1075
rect 34464 1067 34468 1075
rect 34472 1067 34484 1075
rect 34488 1067 34492 1075
rect 34504 1067 34516 1075
rect 34532 1067 34544 1075
rect 34556 1067 34560 1075
rect 34564 1067 34576 1075
rect 34580 1067 34584 1075
rect 34596 1067 34608 1075
rect 34616 1067 34640 1075
rect 34656 1067 34668 1075
rect 34672 1067 34676 1075
rect 34688 1067 34700 1075
rect 34712 1067 34716 1075
rect 34720 1067 34732 1075
rect 34876 1067 34888 1075
rect 34892 1067 34896 1075
rect 34908 1067 34920 1075
rect 34940 1067 34952 1075
rect 34968 1067 35016 1075
rect 35032 1067 35056 1075
rect 35064 1067 35076 1075
rect 35084 1067 35108 1075
rect 35124 1067 35148 1075
rect 35156 1067 35172 1075
rect 35188 1067 35200 1075
rect 35220 1067 35224 1075
rect 35228 1067 35240 1075
rect 35244 1067 35256 1075
rect 35260 1067 35264 1075
rect 35284 1067 35288 1075
rect 35292 1067 35296 1075
rect 35308 1067 35320 1075
rect 35324 1067 35328 1075
rect 35344 1067 35360 1075
rect 35376 1067 35424 1075
rect 35440 1067 35444 1075
rect 35448 1067 35452 1075
rect 35464 1067 35476 1075
rect 35480 1067 35492 1075
rect 35504 1067 35508 1075
rect 35512 1067 35516 1075
rect 35528 1067 35540 1075
rect 35544 1067 35548 1075
rect 35644 1067 35648 1075
rect 35652 1067 35656 1075
rect 35668 1067 35680 1075
rect 35684 1067 35688 1075
rect 35708 1067 35712 1075
rect 35716 1067 35720 1075
rect 35736 1067 35784 1075
rect 35800 1067 35804 1075
rect 35808 1067 35812 1075
rect 35824 1067 35836 1075
rect 35840 1067 35852 1075
rect 35864 1067 35868 1075
rect 35872 1067 35876 1075
rect 35896 1067 35900 1075
rect 35904 1067 35916 1075
rect 35928 1067 35932 1075
rect 35936 1067 35940 1075
rect 35960 1067 35964 1075
rect 35968 1067 35972 1075
rect 35984 1067 35996 1075
rect 36000 1067 36004 1075
rect 36024 1067 36028 1075
rect 36032 1067 36036 1075
rect 36052 1067 36100 1075
rect 36116 1067 36120 1075
rect 36124 1067 36128 1075
rect 36144 1067 36192 1075
rect 36208 1067 36232 1075
rect 36240 1067 36252 1075
rect 36260 1067 36284 1075
rect 36300 1067 36324 1075
rect 36332 1067 36348 1075
rect 36364 1067 36368 1075
rect 36372 1067 36376 1075
rect 36396 1067 36400 1075
rect 36404 1067 36416 1075
rect 36420 1067 36432 1075
rect 36436 1067 36440 1075
rect 36488 1067 36492 1075
rect 36496 1067 36508 1075
rect 36512 1067 36524 1075
rect 36528 1067 36532 1075
rect 36580 1067 36584 1075
rect 36588 1067 36600 1075
rect 36604 1067 36616 1075
rect 36620 1067 36624 1075
rect 36644 1067 36648 1075
rect 36652 1067 36664 1075
rect 36672 1067 36688 1075
rect 36696 1067 36720 1075
rect 36736 1067 36752 1075
rect 36768 1067 36780 1075
rect 36792 1067 36796 1075
rect 36800 1067 36812 1075
rect 36816 1067 36820 1075
rect 36832 1067 36844 1075
rect 36884 1067 36888 1075
rect 36892 1067 36904 1075
rect 36908 1067 36912 1075
rect 36924 1067 36936 1075
rect 36956 1067 36968 1075
rect 36984 1067 37008 1075
rect 37016 1067 37032 1075
rect 37040 1067 37072 1075
rect 37080 1067 37096 1075
rect 37112 1067 37124 1075
rect 37136 1067 37140 1075
rect 37144 1067 37156 1075
rect 37176 1067 37188 1075
rect 37268 1067 37280 1075
rect 37300 1067 37312 1075
rect 37316 1067 37320 1075
rect 37332 1067 37344 1075
rect 37364 1067 37376 1075
rect 37380 1067 37392 1075
rect 37396 1067 37408 1075
rect 37428 1067 37440 1075
rect 37444 1067 37448 1075
rect 37460 1067 37472 1075
rect 37488 1067 37504 1075
rect 37520 1067 37568 1075
rect 37580 1067 37596 1075
rect 37612 1067 37660 1075
rect 37676 1067 37680 1075
rect 37684 1067 37688 1075
rect 37700 1067 37712 1075
rect 37716 1067 37728 1075
rect 37740 1067 37744 1075
rect 37748 1067 37752 1075
rect 37768 1067 37816 1075
rect 37832 1067 37848 1075
rect 37864 1067 37868 1075
rect 37872 1067 37884 1075
rect 37896 1067 37900 1075
rect 37904 1067 37908 1075
rect 38020 1067 38024 1075
rect 38028 1067 38032 1075
rect 38160 1067 38164 1075
rect 38168 1067 38172 1075
rect 38192 1067 38196 1075
rect 38200 1067 38212 1075
rect 38216 1067 38228 1075
rect 38232 1067 38236 1075
rect 38256 1067 38260 1075
rect 38264 1067 38268 1075
rect 38284 1067 38288 1075
rect 38292 1067 38304 1075
rect 38308 1067 38320 1075
rect 38324 1067 38328 1075
rect 38344 1067 38360 1075
rect 38376 1067 38392 1075
rect 38400 1067 38424 1075
rect 38440 1067 38464 1075
rect 38472 1067 38488 1075
rect 38504 1067 38508 1075
rect 38512 1067 38516 1075
rect 38536 1067 38540 1075
rect 38544 1067 38556 1075
rect 38560 1067 38572 1075
rect 38576 1067 38580 1075
rect 38596 1067 38600 1075
rect 38604 1067 38608 1075
rect 38628 1067 38632 1075
rect 38636 1067 38648 1075
rect 38652 1067 38664 1075
rect 38668 1067 38672 1075
rect 38688 1067 38704 1075
rect 38720 1067 38724 1075
rect 38728 1067 38740 1075
rect 38744 1067 38756 1075
rect 38760 1067 38764 1075
rect 38780 1067 38796 1075
rect 38812 1067 38828 1075
rect 38836 1067 38860 1075
rect 38876 1067 38924 1075
rect 38940 1067 38952 1075
rect 38968 1067 39016 1075
rect 39032 1067 39044 1075
rect 39048 1067 39052 1075
rect 39064 1067 39076 1075
rect 39088 1067 39092 1075
rect 39096 1067 39108 1075
rect 39344 1067 39356 1075
rect 39360 1067 39364 1075
rect 39376 1067 39388 1075
rect 39408 1067 39420 1075
rect 39424 1067 39428 1075
rect 39440 1067 39452 1075
rect 39460 1067 39484 1075
rect 39500 1067 39524 1075
rect 39532 1067 39548 1075
rect 39564 1067 39588 1075
rect 39596 1067 39612 1075
rect 39620 1067 39632 1075
rect 39636 1067 39640 1075
rect 39656 1067 39680 1075
rect 39688 1067 39704 1075
rect 39712 1067 39736 1075
rect 39752 1067 39756 1075
rect 39760 1067 39772 1075
rect 39780 1067 39796 1075
rect 39804 1067 39836 1075
rect 39844 1067 39860 1075
rect 39876 1067 39888 1075
rect 39900 1067 39904 1075
rect 39908 1067 39920 1075
rect 39940 1067 39952 1075
rect 40064 1067 40076 1075
rect 40080 1067 40084 1075
rect 40096 1067 40108 1075
rect 40128 1067 40140 1075
rect 40148 1067 40180 1075
rect 40188 1067 40204 1075
rect 40212 1067 40224 1075
rect 40228 1067 40232 1075
rect 40252 1067 40256 1075
rect 40260 1067 40272 1075
rect 40276 1067 40288 1075
rect 40292 1067 40296 1075
rect 40312 1067 40328 1075
rect 40344 1067 40360 1075
rect 40368 1067 40392 1075
rect 40408 1067 40420 1075
rect 40424 1067 40428 1075
rect 40440 1067 40452 1075
rect 40460 1067 40484 1075
rect 40500 1067 40512 1075
rect 40516 1067 40520 1075
rect 40532 1067 40544 1075
rect 40552 1067 40576 1075
rect 40592 1067 40640 1075
rect 40656 1067 40672 1075
rect 40688 1067 40692 1075
rect 40696 1067 40708 1075
rect 40720 1067 40724 1075
rect 40728 1067 40732 1075
rect 40752 1067 40756 1075
rect 40760 1067 40772 1075
rect 40776 1067 40788 1075
rect 40792 1067 40796 1075
rect 20222 1052 20224 1060
rect 20436 1052 20438 1060
rect 20650 1052 20652 1060
rect 20864 1052 20866 1060
rect 21148 1052 21150 1060
rect 21452 1050 21460 1058
rect 21602 1050 21608 1058
rect 21848 1050 21856 1058
rect 21936 1050 21942 1058
rect 21944 1050 21950 1058
rect 22030 1050 22036 1058
rect 22356 1050 22370 1058
rect 22562 1050 22568 1058
rect 22570 1050 22576 1058
rect 22656 1050 22662 1058
rect 22712 1050 22718 1058
rect 22720 1050 22726 1058
rect 23046 1050 23060 1058
rect 23100 1050 23114 1058
rect 23394 1050 23408 1058
rect 23680 1050 23686 1058
rect 23688 1050 23694 1058
rect 23734 1050 23740 1058
rect 23742 1050 23748 1058
rect 23828 1050 23834 1058
rect 24042 1050 24048 1058
rect 24256 1050 24262 1058
rect 24470 1050 24476 1058
rect 24564 1050 24576 1058
rect 24662 1050 24670 1058
rect 24766 1050 24768 1058
rect 24860 1050 24868 1058
rect 25074 1050 25082 1058
rect 25288 1050 25296 1058
rect 25618 1050 25630 1058
rect 25832 1050 25844 1058
rect 26166 1050 26172 1058
rect 26260 1050 26272 1058
rect 26482 1050 26484 1058
rect 26696 1050 26698 1058
rect 26902 1050 26904 1058
rect 27116 1050 27118 1058
rect 27330 1050 27332 1058
rect 27528 1050 27532 1058
rect 27536 1050 27540 1058
rect 27742 1050 27746 1058
rect 27750 1050 27754 1058
rect 27948 1050 27960 1058
rect 28038 1050 28046 1058
rect 35968 1057 35976 1065
rect 36400 1057 36408 1065
rect 37296 1057 37304 1065
rect 1000 1039 1008 1047
rect 3272 1039 3280 1047
rect 3944 1039 3952 1047
rect 4584 1039 4592 1047
rect 7026 1033 7034 1041
rect 8898 1033 8906 1041
rect 10018 1033 10026 1041
rect 13354 1039 13362 1047
rect 13450 1039 13458 1047
rect 13514 1039 13522 1047
rect 13882 1039 13890 1047
rect 15082 1039 15090 1047
rect 15418 1039 15426 1047
rect 15818 1039 15826 1047
rect 16538 1039 16546 1047
rect 16714 1039 16722 1047
rect 18640 1040 18648 1048
rect 26304 1040 26312 1048
rect 29456 1037 29464 1045
rect 30304 1037 30312 1045
rect 31136 1037 31144 1045
rect 31824 1037 31832 1045
rect 32000 1037 32008 1045
rect 34192 1037 34200 1045
rect 35280 1037 35288 1045
rect 35504 1037 35512 1045
rect 35776 1037 35784 1045
rect 38400 1037 38408 1045
rect 38432 1037 38440 1045
rect 39008 1037 39016 1045
rect 536 1019 544 1027
rect 856 1019 864 1027
rect 1192 1019 1200 1027
rect 1240 1019 1248 1027
rect 1288 1019 1296 1027
rect 1400 1019 1408 1027
rect 1656 1019 1664 1027
rect 1768 1019 1776 1027
rect 2072 1019 2080 1027
rect 3384 1019 3392 1027
rect 3448 1019 3456 1027
rect 3496 1019 3504 1027
rect 3720 1019 3728 1027
rect 3736 1019 3744 1027
rect 4056 1019 4064 1027
rect 4248 1019 4256 1027
rect 4360 1019 4368 1027
rect 4456 1019 4464 1027
rect 4616 1019 4624 1027
rect 6450 1013 6458 1021
rect 6850 1013 6858 1021
rect 6930 1013 6938 1021
rect 7026 1013 7034 1021
rect 7218 1013 7226 1021
rect 7362 1013 7370 1021
rect 7570 1013 7578 1021
rect 7666 1013 7674 1021
rect 8194 1013 8202 1021
rect 8626 1013 8634 1021
rect 9090 1013 9098 1021
rect 9842 1013 9850 1021
rect 10050 1013 10058 1021
rect 10450 1013 10458 1021
rect 10498 1013 10506 1021
rect 10610 1013 10618 1021
rect 10850 1013 10858 1021
rect 10914 1013 10922 1021
rect 12362 1019 12370 1027
rect 13498 1019 13506 1027
rect 14234 1019 14242 1027
rect 14298 1019 14306 1027
rect 14554 1019 14562 1027
rect 14666 1019 14674 1027
rect 14810 1019 14818 1027
rect 15306 1019 15314 1027
rect 15514 1019 15522 1027
rect 17370 1019 17378 1027
rect 17434 1019 17442 1027
rect 23488 1020 23496 1028
rect 23856 1020 23864 1028
rect 27680 1020 27688 1028
rect 29568 1017 29576 1025
rect 29968 1017 29976 1025
rect 30048 1017 30056 1025
rect 31616 1017 31624 1025
rect 31728 1017 31736 1025
rect 31872 1017 31880 1025
rect 32480 1017 32488 1025
rect 32576 1017 32584 1025
rect 33056 1017 33064 1025
rect 33088 1017 33096 1025
rect 33552 1017 33560 1025
rect 34128 1017 34136 1025
rect 34352 1017 34360 1025
rect 35920 1017 35928 1025
rect 36704 1017 36712 1025
rect 37152 1017 37160 1025
rect 37264 1017 37272 1025
rect 37312 1017 37320 1025
rect 37632 1017 37640 1025
rect 37648 1017 37656 1025
rect 38128 1017 38136 1025
rect 39056 1017 39064 1025
rect 39120 1017 39128 1025
rect 39168 1017 39176 1025
rect 39632 1017 39640 1025
rect 40032 1017 40040 1025
rect 40208 1017 40216 1025
rect 40480 1017 40488 1025
rect 40608 1017 40616 1025
rect 536 999 544 1007
rect 568 999 576 1007
rect 600 999 608 1007
rect 664 999 672 1007
rect 712 999 720 1007
rect 760 999 768 1007
rect 776 999 784 1007
rect 840 999 848 1007
rect 872 999 880 1007
rect 904 999 912 1007
rect 920 999 928 1007
rect 1000 999 1008 1007
rect 1032 999 1040 1007
rect 1064 999 1072 1007
rect 1304 999 1312 1007
rect 1320 999 1328 1007
rect 1688 999 1696 1007
rect 1768 999 1776 1007
rect 1800 999 1808 1007
rect 1816 999 1824 1007
rect 1896 999 1904 1007
rect 2088 999 2096 1007
rect 2200 999 2208 1007
rect 2232 999 2240 1007
rect 2664 999 2672 1007
rect 2696 999 2704 1007
rect 2824 999 2832 1007
rect 2856 999 2864 1007
rect 2984 999 2992 1007
rect 3016 999 3024 1007
rect 3144 999 3152 1007
rect 3224 999 3232 1007
rect 3240 999 3248 1007
rect 3320 999 3328 1007
rect 3448 999 3456 1007
rect 3544 999 3552 1007
rect 3976 999 3984 1007
rect 4072 999 4080 1007
rect 4264 999 4272 1007
rect 4392 999 4400 1007
rect 4408 999 4416 1007
rect 4520 999 4528 1007
rect 4536 999 4544 1007
rect 4568 999 4576 1007
rect 5858 993 5866 1001
rect 6082 993 6090 1001
rect 6114 993 6122 1001
rect 6578 993 6586 1001
rect 6610 993 6618 1001
rect 6834 993 6842 1001
rect 7586 993 7594 1001
rect 7650 993 7658 1001
rect 7682 993 7690 1001
rect 7698 993 7706 1001
rect 8162 993 8170 1001
rect 8178 993 8186 1001
rect 8258 993 8266 1001
rect 8402 993 8410 1001
rect 8418 993 8426 1001
rect 8450 993 8458 1001
rect 8994 993 9002 1001
rect 9058 993 9066 1001
rect 9122 993 9130 1001
rect 9202 993 9210 1001
rect 9346 993 9354 1001
rect 9490 993 9498 1001
rect 9522 993 9530 1001
rect 9586 993 9594 1001
rect 9826 993 9834 1001
rect 9858 993 9866 1001
rect 10386 993 10394 1001
rect 10674 993 10682 1001
rect 10738 993 10746 1001
rect 10866 993 10874 1001
rect 12234 999 12242 1007
rect 13658 999 13666 1007
rect 15066 999 15074 1007
rect 15802 999 15810 1007
rect 21824 1000 21832 1008
rect 23632 1000 23640 1008
rect 24544 1000 24552 1008
rect 25168 1000 25176 1008
rect 26416 1000 26424 1008
rect 27152 1000 27160 1008
rect 29648 997 29656 1005
rect 29728 997 29736 1005
rect 30016 997 30024 1005
rect 31104 997 31112 1005
rect 31120 997 31128 1005
rect 31488 997 31496 1005
rect 31936 997 31944 1005
rect 32336 997 32344 1005
rect 32432 997 32440 1005
rect 32928 997 32936 1005
rect 33136 997 33144 1005
rect 33344 997 33352 1005
rect 33376 997 33384 1005
rect 33888 997 33896 1005
rect 34784 997 34792 1005
rect 37712 997 37720 1005
rect 38784 997 38792 1005
rect 38832 997 38840 1005
rect 39696 997 39704 1005
rect 39728 997 39736 1005
rect 648 979 656 987
rect 2152 979 2160 987
rect 2360 979 2368 987
rect 2504 979 2512 987
rect 2536 979 2544 987
rect 2600 979 2608 987
rect 2632 979 2640 987
rect 2712 979 2720 987
rect 2776 979 2784 987
rect 2872 979 2880 987
rect 3032 979 3040 987
rect 3272 979 3280 987
rect 4184 979 4192 987
rect 4216 979 4224 987
rect 4296 979 4304 987
rect 4440 979 4448 987
rect 4472 979 4480 987
rect 4504 979 4512 987
rect 6018 973 6026 981
rect 6034 973 6042 981
rect 6066 973 6074 981
rect 6914 973 6922 981
rect 6962 973 6970 981
rect 6994 973 7002 981
rect 7202 973 7210 981
rect 7714 973 7722 981
rect 7794 973 7802 981
rect 7842 973 7850 981
rect 8210 973 8218 981
rect 8290 973 8298 981
rect 8434 973 8442 981
rect 8658 973 8666 981
rect 8674 973 8682 981
rect 8882 973 8890 981
rect 9090 973 9098 981
rect 9154 973 9162 981
rect 9282 973 9290 981
rect 9794 973 9802 981
rect 9954 973 9962 981
rect 10178 973 10186 981
rect 10242 973 10250 981
rect 10322 973 10330 981
rect 10418 973 10426 981
rect 12442 979 12450 987
rect 12474 979 12482 987
rect 12682 979 12690 987
rect 12986 979 12994 987
rect 13130 979 13138 987
rect 13578 979 13586 987
rect 14330 979 14338 987
rect 14410 979 14418 987
rect 15370 979 15378 987
rect 16314 979 16322 987
rect 16522 979 16530 987
rect 17482 979 17490 987
rect 18512 980 18520 988
rect 19040 980 19048 988
rect 19312 980 19320 988
rect 19344 980 19352 988
rect 20144 980 20152 988
rect 20512 980 20520 988
rect 21024 980 21032 988
rect 22688 980 22696 988
rect 23056 980 23064 988
rect 23088 980 23096 988
rect 23712 980 23720 988
rect 23920 980 23928 988
rect 24688 980 24696 988
rect 25312 980 25320 988
rect 25328 980 25336 988
rect 25520 980 25528 988
rect 25552 980 25560 988
rect 25936 980 25944 988
rect 26208 980 26216 988
rect 26768 980 26776 988
rect 27520 980 27528 988
rect 27920 980 27928 988
rect 28480 980 28488 988
rect 29440 977 29448 985
rect 29744 977 29752 985
rect 32880 977 32888 985
rect 33248 977 33256 985
rect 33600 977 33608 985
rect 33632 977 33640 985
rect 33792 977 33800 985
rect 33904 977 33912 985
rect 34784 977 34792 985
rect 34944 977 34952 985
rect 35904 977 35912 985
rect 37136 977 37144 985
rect 38096 977 38104 985
rect 38128 977 38136 985
rect 40688 977 40696 985
rect 472 959 480 967
rect 1704 959 1712 967
rect 2456 959 2464 967
rect 2664 959 2672 967
rect 2840 959 2848 967
rect 3400 959 3408 967
rect 3768 959 3776 967
rect 6434 953 6442 961
rect 6482 953 6490 961
rect 7410 953 7418 961
rect 8146 953 8154 961
rect 8466 953 8474 961
rect 9634 953 9642 961
rect 9698 953 9706 961
rect 10322 953 10330 961
rect 10882 953 10890 961
rect 13850 959 13858 967
rect 14170 959 14178 967
rect 15690 959 15698 967
rect 15722 959 15730 967
rect 15898 959 15906 967
rect 15994 959 16002 967
rect 26608 960 26616 968
rect 27248 960 27256 968
rect 27728 960 27736 968
rect 30944 957 30952 965
rect 31424 957 31432 965
rect 32160 957 32168 965
rect 32352 957 32360 965
rect 33232 957 33240 965
rect 34384 957 34392 965
rect 39264 957 39272 965
rect 40512 957 40520 965
rect 19540 948 19544 953
rect 20752 948 20756 953
rect 21394 948 21398 953
rect 504 939 512 947
rect 808 939 816 947
rect 1080 939 1088 947
rect 1176 939 1184 947
rect 1384 939 1392 947
rect 1656 939 1664 947
rect 1672 939 1680 947
rect 1688 939 1696 947
rect 1896 939 1904 947
rect 2024 939 2032 947
rect 2392 939 2400 947
rect 2440 939 2448 947
rect 2984 939 2992 947
rect 3064 939 3072 947
rect 3096 939 3104 947
rect 3352 939 3360 947
rect 3432 939 3440 947
rect 3608 939 3616 947
rect 3832 939 3840 947
rect 4008 939 4016 947
rect 4024 939 4032 947
rect 4056 939 4064 947
rect 4440 939 4448 947
rect 5826 933 5834 941
rect 6674 933 6682 941
rect 7186 933 7194 941
rect 7698 933 7706 941
rect 7810 933 7818 941
rect 7906 933 7914 941
rect 7970 933 7978 941
rect 8706 933 8714 941
rect 8786 933 8794 941
rect 8898 933 8906 941
rect 8930 933 8938 941
rect 9474 933 9482 941
rect 9522 933 9530 941
rect 9666 933 9674 941
rect 10722 933 10730 941
rect 10786 933 10794 941
rect 10898 933 10906 941
rect 10914 933 10922 941
rect 12346 939 12354 947
rect 13914 939 13922 947
rect 14106 939 14114 947
rect 14730 939 14738 947
rect 14746 939 14754 947
rect 14890 939 14898 947
rect 14938 939 14946 947
rect 15210 939 15218 947
rect 15354 939 15362 947
rect 16938 939 16946 947
rect 16986 939 16994 947
rect 17098 939 17106 947
rect 17194 939 17202 947
rect 17290 939 17298 947
rect 17338 939 17346 947
rect 17466 939 17474 947
rect 19040 940 19048 948
rect 19904 940 19912 948
rect 20096 940 20104 948
rect 20528 940 20536 948
rect 20960 940 20968 948
rect 21424 940 21432 948
rect 21632 940 21640 948
rect 22048 940 22056 948
rect 22208 940 22216 948
rect 22384 940 22392 948
rect 22608 940 22616 948
rect 23424 940 23432 948
rect 23904 940 23912 948
rect 25760 940 25768 948
rect 27712 940 27720 948
rect 27904 940 27912 948
rect 38816 937 38824 945
rect 2104 919 2112 927
rect 3240 919 3248 927
rect 3864 919 3872 927
rect 4040 919 4048 927
rect 6546 913 6554 921
rect 6594 913 6602 921
rect 6946 913 6954 921
rect 7106 913 7114 921
rect 7522 913 7530 921
rect 7602 913 7610 921
rect 7650 913 7658 921
rect 8610 913 8618 921
rect 9010 913 9018 921
rect 9026 913 9034 921
rect 10322 913 10330 921
rect 10738 913 10746 921
rect 12442 919 12450 927
rect 12506 919 12514 927
rect 12922 919 12930 927
rect 15498 919 15506 927
rect 16426 919 16434 927
rect 17242 919 17250 927
rect 25104 920 25112 928
rect 25200 920 25208 928
rect 27888 920 27896 928
rect 32048 917 32056 925
rect 32512 917 32520 925
rect 33168 917 33176 925
rect 1928 899 1936 907
rect 6482 893 6490 901
rect 7122 893 7130 901
rect 7666 893 7674 901
rect 9442 893 9450 901
rect 9602 893 9610 901
rect 15706 899 15714 907
rect 26032 900 26040 908
rect 27312 900 27320 908
rect 520 879 528 887
rect 888 879 896 887
rect 1048 879 1056 887
rect 1336 879 1344 887
rect 1784 879 1792 887
rect 1832 879 1840 887
rect 2216 879 2224 887
rect 2680 879 2688 887
rect 2952 879 2960 887
rect 2968 879 2976 887
rect 3720 879 3728 887
rect 4552 879 4560 887
rect 7426 873 7434 881
rect 10018 873 10026 881
rect 12378 879 12386 887
rect 12474 879 12482 887
rect 16138 879 16146 887
rect 16154 879 16162 887
rect 19936 880 19944 888
rect 22224 880 22232 888
rect 34528 877 34536 885
rect 34960 877 34968 885
rect 29396 867 29408 875
rect 29428 867 29440 875
rect 29444 867 29448 875
rect 29460 867 29472 875
rect 29488 867 29504 875
rect 29512 867 29544 875
rect 29552 867 29568 875
rect 29576 867 29588 875
rect 29592 867 29596 875
rect 29612 867 29636 875
rect 29644 867 29660 875
rect 29668 867 29692 875
rect 29708 867 29712 875
rect 29716 867 29728 875
rect 29740 867 29744 875
rect 29748 867 29752 875
rect 29772 867 29776 875
rect 29780 867 29784 875
rect 29880 867 29884 875
rect 29888 867 29900 875
rect 29904 867 29916 875
rect 29920 867 29924 875
rect 29944 867 29948 875
rect 29952 867 29964 875
rect 29968 867 29980 875
rect 29984 867 29988 875
rect 30008 867 30012 875
rect 30016 867 30020 875
rect 30040 867 30044 875
rect 30048 867 30052 875
rect 30072 867 30076 875
rect 30080 867 30084 875
rect 30104 867 30108 875
rect 30112 867 30124 875
rect 30128 867 30140 875
rect 30144 867 30148 875
rect 30196 867 30200 875
rect 30204 867 30216 875
rect 30220 867 30232 875
rect 30236 867 30240 875
rect 30260 867 30264 875
rect 30268 867 30272 875
rect 30292 867 30296 875
rect 30300 867 30304 875
rect 30324 867 30328 875
rect 30332 867 30336 875
rect 30356 867 30360 875
rect 30364 867 30376 875
rect 30380 867 30392 875
rect 30396 867 30400 875
rect 30416 867 30432 875
rect 30448 867 30464 875
rect 30472 867 30496 875
rect 30512 867 30524 875
rect 30528 867 30532 875
rect 30544 867 30556 875
rect 30568 867 30572 875
rect 30576 867 30588 875
rect 30592 867 30596 875
rect 30700 867 30712 875
rect 30732 867 30744 875
rect 30748 867 30760 875
rect 30764 867 30776 875
rect 30824 867 30836 875
rect 30840 867 30852 875
rect 30856 867 30868 875
rect 30884 867 30900 875
rect 30908 867 30940 875
rect 30948 867 30964 875
rect 30980 867 30992 875
rect 31000 867 31032 875
rect 31040 867 31056 875
rect 31072 867 31076 875
rect 31080 867 31084 875
rect 31104 867 31108 875
rect 31112 867 31124 875
rect 31136 867 31140 875
rect 31144 867 31148 875
rect 31160 867 31172 875
rect 31176 867 31188 875
rect 31200 867 31204 875
rect 31208 867 31212 875
rect 31232 867 31236 875
rect 31240 867 31244 875
rect 31264 867 31268 875
rect 31272 867 31276 875
rect 31296 867 31300 875
rect 31304 867 31308 875
rect 31320 867 31332 875
rect 31336 867 31348 875
rect 31356 867 31372 875
rect 31388 867 31404 875
rect 31412 867 31436 875
rect 31452 867 31464 875
rect 31484 867 31496 875
rect 31500 867 31512 875
rect 31516 867 31528 875
rect 31544 867 31560 875
rect 31576 867 31600 875
rect 31608 867 31624 875
rect 31640 867 31688 875
rect 31704 867 31720 875
rect 31732 867 31780 875
rect 31796 867 31812 875
rect 31828 867 31844 875
rect 31860 867 31876 875
rect 31892 867 31940 875
rect 31956 867 31960 875
rect 31964 867 31968 875
rect 31984 867 32032 875
rect 32048 867 32052 875
rect 32056 867 32060 875
rect 32076 867 32124 875
rect 32140 867 32144 875
rect 32148 867 32152 875
rect 32164 867 32176 875
rect 32180 867 32192 875
rect 32204 867 32208 875
rect 32212 867 32216 875
rect 32312 867 32316 875
rect 32320 867 32332 875
rect 32344 867 32348 875
rect 32352 867 32356 875
rect 32368 867 32380 875
rect 32384 867 32388 875
rect 32436 867 32440 875
rect 32444 867 32448 875
rect 32460 867 32472 875
rect 32476 867 32488 875
rect 32500 867 32504 875
rect 32508 867 32512 875
rect 32524 867 32536 875
rect 32540 867 32544 875
rect 32592 867 32596 875
rect 32600 867 32604 875
rect 32616 867 32628 875
rect 32632 867 32636 875
rect 32652 867 32668 875
rect 32684 867 32700 875
rect 32708 867 32740 875
rect 32748 867 32764 875
rect 32780 867 32792 875
rect 32796 867 32808 875
rect 32812 867 32824 875
rect 32936 867 32948 875
rect 32960 867 32964 875
rect 32968 867 32980 875
rect 32984 867 32988 875
rect 33028 867 33040 875
rect 33052 867 33056 875
rect 33060 867 33072 875
rect 33076 867 33080 875
rect 33092 867 33104 875
rect 33116 867 33120 875
rect 33124 867 33136 875
rect 33140 867 33144 875
rect 33184 867 33196 875
rect 33208 867 33212 875
rect 33216 867 33228 875
rect 33232 867 33236 875
rect 33248 867 33260 875
rect 33532 867 33544 875
rect 33548 867 33552 875
rect 33564 867 33576 875
rect 33600 867 33608 875
rect 33620 867 33624 875
rect 33628 867 33640 875
rect 33660 867 33672 875
rect 33692 867 33704 875
rect 33708 867 33712 875
rect 33724 867 33736 875
rect 33756 867 33768 875
rect 33780 867 33784 875
rect 33788 867 33800 875
rect 34028 867 34032 875
rect 34036 867 34048 875
rect 34052 867 34056 875
rect 34160 867 34172 875
rect 34192 867 34204 875
rect 34208 867 34220 875
rect 34224 867 34236 875
rect 34252 867 34268 875
rect 34276 867 34308 875
rect 34316 867 34332 875
rect 34344 867 34360 875
rect 34368 867 34400 875
rect 34408 867 34424 875
rect 34436 867 34452 875
rect 34460 867 34492 875
rect 34500 867 34516 875
rect 34532 867 34544 875
rect 34548 867 34560 875
rect 34564 867 34576 875
rect 34596 867 34608 875
rect 34616 867 34648 875
rect 34656 867 34668 875
rect 34688 867 34700 875
rect 34708 867 34740 875
rect 34748 867 34760 875
rect 34780 867 34792 875
rect 34796 867 34808 875
rect 34812 867 34824 875
rect 34840 867 34856 875
rect 34872 867 34884 875
rect 34888 867 34900 875
rect 34904 867 34916 875
rect 34936 867 34948 875
rect 34952 867 34956 875
rect 35028 867 35040 875
rect 35044 867 35056 875
rect 35060 867 35072 875
rect 35088 867 35100 875
rect 35120 867 35132 875
rect 35136 867 35148 875
rect 35152 867 35164 875
rect 35184 867 35196 875
rect 35340 867 35352 875
rect 35372 867 35384 875
rect 35388 867 35400 875
rect 35404 867 35416 875
rect 35464 867 35476 875
rect 35480 867 35492 875
rect 35496 867 35508 875
rect 35528 867 35540 875
rect 35544 867 35548 875
rect 35580 867 35584 875
rect 35588 867 35600 875
rect 35620 867 35632 875
rect 35636 867 35640 875
rect 35712 867 35724 875
rect 35728 867 35732 875
rect 35804 867 35816 875
rect 35820 867 35832 875
rect 35836 867 35848 875
rect 35868 867 35880 875
rect 35896 867 35920 875
rect 35928 867 35944 875
rect 35960 867 35976 875
rect 35984 867 35996 875
rect 36000 867 36012 875
rect 36024 867 36028 875
rect 36032 867 36036 875
rect 36052 867 36100 875
rect 36116 867 36132 875
rect 36144 867 36192 875
rect 36208 867 36224 875
rect 36240 867 36252 875
rect 36264 867 36268 875
rect 36272 867 36284 875
rect 36304 867 36316 875
rect 36320 867 36324 875
rect 36336 867 36348 875
rect 36364 867 36380 875
rect 36396 867 36444 875
rect 36460 867 36464 875
rect 36468 867 36472 875
rect 36488 867 36536 875
rect 36552 867 36568 875
rect 36580 867 36628 875
rect 36644 867 36648 875
rect 36652 867 36656 875
rect 36672 867 36720 875
rect 36736 867 36752 875
rect 36768 867 36780 875
rect 36792 867 36796 875
rect 36800 867 36812 875
rect 36832 867 36844 875
rect 36848 867 36852 875
rect 36924 867 36936 875
rect 36940 867 36944 875
rect 36956 867 36968 875
rect 36988 867 37000 875
rect 37016 867 37064 875
rect 37080 867 37096 875
rect 37108 867 37156 875
rect 37172 867 37176 875
rect 37180 867 37184 875
rect 37200 867 37248 875
rect 37264 867 37268 875
rect 37272 867 37276 875
rect 37296 867 37300 875
rect 37304 867 37316 875
rect 37328 867 37332 875
rect 37336 867 37340 875
rect 37360 867 37364 875
rect 37368 867 37372 875
rect 37436 867 37440 875
rect 37444 867 37448 875
rect 37468 867 37472 875
rect 37476 867 37480 875
rect 37492 867 37504 875
rect 37508 867 37512 875
rect 37532 867 37536 875
rect 37540 867 37552 875
rect 37556 867 37568 875
rect 37572 867 37576 875
rect 37624 867 37628 875
rect 37632 867 37644 875
rect 37648 867 37660 875
rect 37664 867 37668 875
rect 37688 867 37692 875
rect 37696 867 37708 875
rect 37716 867 37732 875
rect 37740 867 37764 875
rect 37780 867 37784 875
rect 37788 867 37800 875
rect 37808 867 37824 875
rect 37832 867 37856 875
rect 37872 867 37888 875
rect 37904 867 37920 875
rect 37936 867 37960 875
rect 37968 867 37984 875
rect 37992 867 38016 875
rect 38028 867 38052 875
rect 38060 867 38076 875
rect 38084 867 38108 875
rect 38124 867 38136 875
rect 38156 867 38168 875
rect 38180 867 38184 875
rect 38188 867 38200 875
rect 38204 867 38208 875
rect 38220 867 38232 875
rect 38252 867 38264 875
rect 38280 867 38304 875
rect 38312 867 38328 875
rect 38336 867 38360 875
rect 38376 867 38392 875
rect 38400 867 38424 875
rect 38440 867 38452 875
rect 38456 867 38460 875
rect 38472 867 38484 875
rect 38492 867 38516 875
rect 38532 867 38544 875
rect 38548 867 38552 875
rect 38564 867 38576 875
rect 38584 867 38608 875
rect 38624 867 38672 875
rect 38688 867 38700 875
rect 38716 867 38764 875
rect 38780 867 38796 875
rect 38812 867 38824 875
rect 38836 867 38840 875
rect 38844 867 38856 875
rect 39052 867 39056 875
rect 39060 867 39072 875
rect 39092 867 39104 875
rect 39108 867 39112 875
rect 39124 867 39136 875
rect 39156 867 39168 875
rect 39184 867 39232 875
rect 39248 867 39260 875
rect 39276 867 39324 875
rect 39340 867 39356 875
rect 39372 867 39388 875
rect 39404 867 39420 875
rect 39436 867 39484 875
rect 39500 867 39516 875
rect 39532 867 39536 875
rect 39540 867 39552 875
rect 39564 867 39568 875
rect 39572 867 39576 875
rect 39596 867 39600 875
rect 39604 867 39616 875
rect 39620 867 39632 875
rect 39636 867 39640 875
rect 39656 867 39672 875
rect 39688 867 39692 875
rect 39696 867 39708 875
rect 39712 867 39724 875
rect 39728 867 39732 875
rect 39780 867 39784 875
rect 39788 867 39800 875
rect 39804 867 39816 875
rect 39820 867 39824 875
rect 39872 867 39876 875
rect 39880 867 39892 875
rect 39896 867 39908 875
rect 39912 867 39916 875
rect 39936 867 39940 875
rect 39944 867 39948 875
rect 39964 867 39968 875
rect 39972 867 39984 875
rect 39988 867 40000 875
rect 40004 867 40008 875
rect 40028 867 40032 875
rect 40036 867 40040 875
rect 40296 867 40300 875
rect 40304 867 40308 875
rect 40356 867 40360 875
rect 40364 867 40376 875
rect 40388 867 40392 875
rect 40396 867 40400 875
rect 40496 867 40500 875
rect 40504 867 40508 875
rect 40528 867 40532 875
rect 40536 867 40540 875
rect 40552 867 40564 875
rect 40568 867 40580 875
rect 40592 867 40596 875
rect 40600 867 40604 875
rect 40616 867 40628 875
rect 40632 867 40636 875
rect 40700 867 40704 875
rect 40708 867 40712 875
rect 40732 867 40736 875
rect 40740 867 40744 875
rect 40756 867 40768 875
rect 40772 867 40784 875
rect 40796 867 40800 875
rect 868 863 892 867
rect 1512 859 1520 867
rect 2936 859 2944 867
rect 7138 853 7146 861
rect 8738 853 8746 861
rect 8754 853 8762 861
rect 10418 853 10426 861
rect 10770 853 10778 861
rect 13050 859 13058 867
rect 13242 859 13250 867
rect 16810 859 16818 867
rect 19608 850 19610 858
rect 19616 850 19618 858
rect 21090 850 21092 858
rect 21098 850 21100 858
rect 22326 850 22328 858
rect 22334 850 22336 858
rect 22540 850 22542 858
rect 22548 850 22550 858
rect 23746 850 23750 858
rect 23754 850 23758 858
rect 24174 850 24178 858
rect 24182 850 24186 858
rect 25266 850 25276 858
rect 25472 850 25474 858
rect 25480 850 25482 858
rect 25686 850 25688 858
rect 25694 850 25696 858
rect 7458 833 7466 841
rect 7634 833 7642 841
rect 14138 839 14146 847
rect 23072 840 23080 848
rect 23712 840 23720 848
rect 24128 840 24136 848
rect 31168 837 31176 845
rect 33056 837 33064 845
rect 424 819 432 827
rect 552 819 560 827
rect 840 819 848 827
rect 1288 819 1296 827
rect 1304 819 1312 827
rect 1992 819 2000 827
rect 2088 819 2096 827
rect 2408 819 2416 827
rect 3256 819 3264 827
rect 3448 819 3456 827
rect 3576 819 3584 827
rect 3656 819 3664 827
rect 3976 819 3984 827
rect 4056 819 4064 827
rect 4072 819 4080 827
rect 4312 819 4320 827
rect 4376 819 4384 827
rect 4472 819 4480 827
rect 4632 819 4640 827
rect 6882 813 6890 821
rect 7842 813 7850 821
rect 7906 813 7914 821
rect 8946 813 8954 821
rect 9282 813 9290 821
rect 9378 813 9386 821
rect 10530 813 10538 821
rect 10882 813 10890 821
rect 13082 819 13090 827
rect 14170 819 14178 827
rect 14538 819 14546 827
rect 14618 819 14626 827
rect 14922 819 14930 827
rect 15498 819 15506 827
rect 16826 819 16834 827
rect 32096 817 32104 825
rect 32864 817 32872 825
rect 36544 817 36552 825
rect 40048 817 40056 825
rect 1080 799 1088 807
rect 1480 799 1488 807
rect 2104 799 2112 807
rect 2984 799 2992 807
rect 6834 793 6842 801
rect 7218 793 7226 801
rect 8914 793 8922 801
rect 9154 793 9162 801
rect 9762 793 9770 801
rect 10370 793 10378 801
rect 10610 793 10618 801
rect 13210 799 13218 807
rect 13834 799 13842 807
rect 13978 799 13986 807
rect 15882 799 15890 807
rect 16170 799 16178 807
rect 16602 799 16610 807
rect 16714 799 16722 807
rect 17242 799 17250 807
rect 24736 800 24744 808
rect 24816 800 24824 808
rect 25216 800 25224 808
rect 33360 800 33368 805
rect 33472 800 33480 805
rect 35024 800 35032 805
rect 40400 800 40408 805
rect 40720 800 40728 805
rect 1704 779 1712 787
rect 2184 779 2192 787
rect 2264 779 2272 787
rect 2344 779 2352 787
rect 2600 779 2608 787
rect 2648 779 2656 787
rect 2712 779 2720 787
rect 3912 779 3920 787
rect 6258 773 6266 781
rect 6482 773 6490 781
rect 6530 773 6538 781
rect 6802 773 6810 781
rect 7042 773 7050 781
rect 7506 773 7514 781
rect 8146 773 8154 781
rect 8194 773 8202 781
rect 8226 773 8234 781
rect 8274 773 8282 781
rect 8306 773 8314 781
rect 9730 773 9738 781
rect 9938 773 9946 781
rect 10114 773 10122 781
rect 10210 773 10218 781
rect 10450 773 10458 781
rect 10514 773 10522 781
rect 10546 773 10554 781
rect 10594 773 10602 781
rect 10674 773 10682 781
rect 12810 779 12818 787
rect 14858 779 14866 787
rect 14874 779 14882 787
rect 15370 779 15378 787
rect 16266 779 16274 787
rect 16730 779 16738 787
rect 16746 779 16754 787
rect 17226 779 17234 787
rect 17482 779 17490 787
rect 20720 780 20728 788
rect 26448 780 26456 788
rect 26496 780 26504 788
rect 26848 780 26856 788
rect 920 759 928 767
rect 1480 759 1488 767
rect 1528 759 1536 767
rect 2568 759 2576 767
rect 2824 759 2832 767
rect 2872 759 2880 767
rect 3176 759 3184 767
rect 3368 759 3376 767
rect 3400 759 3408 767
rect 3432 759 3440 767
rect 3464 759 3472 767
rect 4280 759 4288 767
rect 4360 759 4368 767
rect 4600 759 4608 767
rect 6322 753 6330 761
rect 7346 753 7354 761
rect 7746 753 7754 761
rect 8130 753 8138 761
rect 8434 753 8442 761
rect 8770 753 8778 761
rect 9682 753 9690 761
rect 9778 753 9786 761
rect 9794 753 9802 761
rect 9874 753 9882 761
rect 12170 759 12178 767
rect 12314 759 12322 767
rect 12570 759 12578 767
rect 13210 759 13218 767
rect 13258 759 13266 767
rect 13418 759 13426 767
rect 14394 759 14402 767
rect 15002 759 15010 767
rect 15690 759 15698 767
rect 15754 759 15762 767
rect 15802 759 15810 767
rect 16682 759 16690 767
rect 18848 760 18856 768
rect 19056 761 19066 766
rect 19328 760 19336 768
rect 19682 761 19692 766
rect 19888 760 19896 768
rect 20480 760 20488 768
rect 20804 761 20807 766
rect 21408 760 21416 768
rect 22048 760 22056 768
rect 22480 760 22488 768
rect 23472 760 23480 768
rect 24528 760 24536 768
rect 24800 760 24808 768
rect 25810 761 25820 766
rect 26448 760 26456 768
rect 27296 760 27304 768
rect 27504 760 27512 768
rect 27696 760 27704 768
rect 27888 760 27896 768
rect 776 739 784 747
rect 1144 739 1152 747
rect 1496 739 1504 747
rect 1672 739 1680 747
rect 3336 739 3344 747
rect 6578 733 6586 741
rect 6802 733 6810 741
rect 6866 733 6874 741
rect 7074 733 7082 741
rect 8482 733 8490 741
rect 8898 733 8906 741
rect 9426 733 9434 741
rect 9442 733 9450 741
rect 9458 733 9466 741
rect 10802 733 10810 741
rect 12186 739 12194 747
rect 14506 739 14514 747
rect 14554 739 14562 747
rect 17018 739 17026 747
rect 17274 739 17282 747
rect 17370 739 17378 747
rect 17434 739 17442 747
rect 19952 740 19960 748
rect 21392 740 21400 748
rect 22640 740 22648 748
rect 24352 740 24360 748
rect 24704 740 24712 748
rect 29424 737 29432 745
rect 568 719 576 727
rect 648 719 656 727
rect 1016 719 1024 727
rect 1864 719 1872 727
rect 2024 719 2032 727
rect 2248 719 2256 727
rect 2376 719 2384 727
rect 2600 719 2608 727
rect 3128 719 3136 727
rect 3544 719 3552 727
rect 3720 719 3728 727
rect 4040 719 4048 727
rect 4088 719 4096 727
rect 4520 719 4528 727
rect 4568 719 4576 727
rect 5938 713 5946 721
rect 6050 713 6058 721
rect 7170 713 7178 721
rect 7986 713 7994 721
rect 8050 713 8058 721
rect 8130 713 8138 721
rect 8578 713 8586 721
rect 8674 713 8682 721
rect 8770 713 8778 721
rect 9282 713 9290 721
rect 10354 713 10362 721
rect 12170 719 12178 727
rect 12234 719 12242 727
rect 12986 719 12994 727
rect 13386 719 13394 727
rect 14810 719 14818 727
rect 14874 719 14882 727
rect 15770 719 15778 727
rect 15786 719 15794 727
rect 15818 719 15826 727
rect 15850 719 15858 727
rect 15930 719 15938 727
rect 17034 719 17042 727
rect 17178 719 17186 727
rect 17290 719 17298 727
rect 18832 720 18840 728
rect 19152 720 19160 728
rect 19968 720 19976 728
rect 21568 720 21576 728
rect 22064 720 22072 728
rect 22272 720 22280 728
rect 23024 720 23032 728
rect 23472 720 23480 728
rect 23776 720 23784 728
rect 24512 720 24520 728
rect 25232 720 25240 728
rect 25424 720 25432 728
rect 27520 720 27528 728
rect 27824 720 27832 728
rect 520 699 528 707
rect 536 699 544 707
rect 632 699 640 707
rect 664 699 672 707
rect 760 699 768 707
rect 824 699 832 707
rect 856 699 864 707
rect 1064 699 1072 707
rect 1096 699 1104 707
rect 1176 699 1184 707
rect 1208 699 1216 707
rect 1272 699 1280 707
rect 1320 699 1328 707
rect 1384 699 1392 707
rect 1464 699 1472 707
rect 1512 699 1520 707
rect 1640 699 1648 707
rect 1720 699 1728 707
rect 1784 699 1792 707
rect 1800 699 1808 707
rect 1976 699 1984 707
rect 2008 699 2016 707
rect 2072 699 2080 707
rect 2248 699 2256 707
rect 2424 699 2432 707
rect 2440 699 2448 707
rect 2472 699 2480 707
rect 2648 699 2656 707
rect 2680 699 2688 707
rect 3000 699 3008 707
rect 3064 699 3072 707
rect 3080 699 3088 707
rect 3240 699 3248 707
rect 3272 699 3280 707
rect 3352 699 3360 707
rect 3592 699 3600 707
rect 3672 699 3680 707
rect 3928 699 3936 707
rect 3944 699 3952 707
rect 3960 699 3968 707
rect 4040 699 4048 707
rect 4088 699 4096 707
rect 4152 699 4160 707
rect 4264 699 4272 707
rect 4296 699 4304 707
rect 4392 699 4400 707
rect 4456 699 4464 707
rect 4488 699 4496 707
rect 4520 699 4528 707
rect 5778 693 5786 701
rect 5842 693 5850 701
rect 6050 693 6058 701
rect 6914 693 6922 701
rect 6930 693 6938 701
rect 7058 693 7066 701
rect 7474 693 7482 701
rect 7826 693 7834 701
rect 7922 693 7930 701
rect 8002 693 8010 701
rect 8018 693 8026 701
rect 8290 693 8298 701
rect 8530 693 8538 701
rect 8786 693 8794 701
rect 8850 693 8858 701
rect 8930 693 8938 701
rect 8962 693 8970 701
rect 9842 693 9850 701
rect 10402 693 10410 701
rect 10434 693 10442 701
rect 10514 693 10522 701
rect 10690 693 10698 701
rect 10722 693 10730 701
rect 10754 693 10762 701
rect 10866 693 10874 701
rect 12106 699 12114 707
rect 13546 699 13554 707
rect 15050 699 15058 707
rect 15130 699 15138 707
rect 15626 699 15634 707
rect 17082 699 17090 707
rect 25840 700 25848 708
rect 26160 700 26168 708
rect 28048 700 28056 708
rect 424 679 432 687
rect 1192 679 1200 687
rect 1944 679 1952 687
rect 2328 679 2336 687
rect 2456 679 2464 687
rect 2712 679 2720 687
rect 2872 679 2880 687
rect 3096 679 3104 687
rect 3144 679 3152 687
rect 3288 679 3296 687
rect 3768 679 3776 687
rect 3816 679 3824 687
rect 3944 679 3952 687
rect 6722 673 6730 681
rect 7042 673 7050 681
rect 7314 673 7322 681
rect 7346 673 7354 681
rect 7378 673 7386 681
rect 8946 673 8954 681
rect 9826 673 9834 681
rect 12298 679 12306 687
rect 13450 679 13458 687
rect 22784 680 22792 688
rect 23088 680 23096 688
rect 23920 680 23928 688
rect 25376 680 25384 688
rect 25792 680 25800 688
rect 25984 680 25992 688
rect 26384 680 26392 688
rect 1096 659 1104 667
rect 2328 659 2336 667
rect 6914 653 6922 661
rect 7394 653 7402 661
rect 7554 653 7562 661
rect 7634 653 7642 661
rect 7698 653 7706 661
rect 7986 653 7994 661
rect 8034 653 8042 661
rect 8706 653 8714 661
rect 12298 659 12306 667
rect 12874 659 12882 667
rect 12890 659 12898 667
rect 13482 659 13490 667
rect 15130 659 15138 667
rect 16138 659 16146 667
rect 17114 659 17122 667
rect 19968 660 19976 668
rect 20352 660 20360 668
rect 22416 660 22424 668
rect 24576 660 24584 668
rect 25568 660 25576 668
rect 27264 660 27272 668
rect 29396 667 29408 675
rect 29428 667 29440 675
rect 29444 667 29448 675
rect 29460 667 29472 675
rect 29488 667 29504 675
rect 29512 667 29544 675
rect 29552 667 29568 675
rect 29576 667 29588 675
rect 29592 667 29596 675
rect 20414 656 20416 660
rect 20628 656 20630 660
rect 20420 652 20422 656
rect 20634 652 20636 656
rect 21030 650 21034 658
rect 21120 650 21128 658
rect 21548 650 21562 658
rect 22030 650 22038 658
rect 22180 650 22186 658
rect 22458 650 22472 658
rect 22608 650 22614 658
rect 22664 650 22670 658
rect 22672 650 22678 658
rect 23442 650 23456 658
rect 23496 650 23510 658
rect 23796 650 23802 658
rect 23898 650 23900 658
rect 23990 650 24000 658
rect 24326 650 24328 658
rect 24488 650 24494 658
rect 24496 650 24502 658
rect 24542 650 24548 658
rect 24550 650 24556 658
rect 24616 656 24620 658
rect 24694 650 24708 658
rect 24748 650 24762 658
rect 25184 650 25190 658
rect 25192 650 25198 658
rect 25342 650 25348 658
rect 25390 650 25404 658
rect 25604 650 25618 658
rect 26766 652 26768 660
rect 26980 652 26982 660
rect 27284 650 27298 658
rect 28002 652 28004 660
rect 1752 639 1760 647
rect 1816 639 1824 647
rect 3144 639 3152 647
rect 4440 639 4448 647
rect 6818 633 6826 641
rect 7794 633 7802 641
rect 7874 633 7882 641
rect 8194 633 8202 641
rect 9154 633 9162 641
rect 9826 633 9834 641
rect 9938 633 9946 641
rect 9970 633 9978 641
rect 10050 633 10058 641
rect 10210 633 10218 641
rect 10642 633 10650 641
rect 12586 639 12594 647
rect 14362 639 14370 647
rect 15962 639 15970 647
rect 15978 639 15986 647
rect 16650 639 16658 647
rect 16986 639 16994 647
rect 17034 639 17042 647
rect 17050 639 17058 647
rect 24464 640 24472 648
rect 696 619 704 627
rect 1240 619 1248 627
rect 2248 619 2256 627
rect 2424 619 2432 627
rect 2632 619 2640 627
rect 2712 619 2720 627
rect 2856 619 2864 627
rect 3448 619 3456 627
rect 3672 619 3680 627
rect 3736 619 3744 627
rect 3768 619 3776 627
rect 3784 619 3792 627
rect 4360 619 4368 627
rect 4552 619 4560 627
rect 5922 613 5930 621
rect 6242 613 6250 621
rect 6482 613 6490 621
rect 6546 613 6554 621
rect 7186 613 7194 621
rect 7650 613 7658 621
rect 8194 613 8202 621
rect 8626 613 8634 621
rect 8770 613 8778 621
rect 8914 613 8922 621
rect 9058 613 9066 621
rect 9154 613 9162 621
rect 9778 613 9786 621
rect 10434 613 10442 621
rect 10450 613 10458 621
rect 10610 613 10618 621
rect 13466 619 13474 627
rect 14362 619 14370 627
rect 14410 619 14418 627
rect 14426 619 14434 627
rect 14474 619 14482 627
rect 14506 619 14514 627
rect 14938 619 14946 627
rect 15130 619 15138 627
rect 16170 619 16178 627
rect 16202 619 16210 627
rect 16330 619 16338 627
rect 16970 619 16978 627
rect 20368 620 20376 628
rect 20592 620 20600 628
rect 22000 620 22008 628
rect 24016 620 24024 628
rect 24880 620 24888 628
rect 27408 620 27416 628
rect 29504 617 29512 625
rect 29584 617 29592 625
rect 568 599 576 607
rect 584 599 592 607
rect 744 599 752 607
rect 776 599 784 607
rect 872 599 880 607
rect 904 599 912 607
rect 1016 599 1024 607
rect 1032 599 1040 607
rect 1112 599 1120 607
rect 1128 599 1136 607
rect 1192 599 1200 607
rect 1224 599 1232 607
rect 1256 599 1264 607
rect 1272 599 1280 607
rect 1352 599 1360 607
rect 1400 599 1408 607
rect 1416 599 1424 607
rect 1432 599 1440 607
rect 1800 599 1808 607
rect 1960 599 1968 607
rect 2056 599 2064 607
rect 2264 599 2272 607
rect 2328 599 2336 607
rect 2360 599 2368 607
rect 2392 599 2400 607
rect 2408 599 2416 607
rect 2600 599 2608 607
rect 2680 599 2688 607
rect 2696 599 2704 607
rect 2840 599 2848 607
rect 2920 599 2928 607
rect 3080 599 3088 607
rect 3160 599 3168 607
rect 3224 599 3232 607
rect 3368 599 3376 607
rect 3640 599 3648 607
rect 3672 599 3680 607
rect 3832 599 3840 607
rect 3928 599 3936 607
rect 3976 599 3984 607
rect 4200 599 4208 607
rect 4264 599 4272 607
rect 4376 599 4384 607
rect 4536 599 4544 607
rect 5762 593 5770 601
rect 5874 593 5882 601
rect 5938 593 5946 601
rect 6130 593 6138 601
rect 6258 593 6266 601
rect 6290 593 6298 601
rect 6466 593 6474 601
rect 6482 593 6490 601
rect 6786 593 6794 601
rect 6818 593 6826 601
rect 6850 593 6858 601
rect 7154 593 7162 601
rect 7426 593 7434 601
rect 7442 593 7450 601
rect 7506 593 7514 601
rect 7522 593 7530 601
rect 7602 593 7610 601
rect 7650 593 7658 601
rect 7666 593 7674 601
rect 7682 593 7690 601
rect 7762 593 7770 601
rect 8242 593 8250 601
rect 8402 593 8410 601
rect 8482 593 8490 601
rect 8530 593 8538 601
rect 8658 593 8666 601
rect 8738 593 8746 601
rect 8978 593 8986 601
rect 9506 593 9514 601
rect 9794 593 9802 601
rect 9858 593 9866 601
rect 9890 593 9898 601
rect 10034 593 10042 601
rect 10194 593 10202 601
rect 10306 593 10314 601
rect 10370 593 10378 601
rect 10594 593 10602 601
rect 10754 593 10762 601
rect 10770 593 10778 601
rect 10786 593 10794 601
rect 13834 599 13842 607
rect 14618 599 14626 607
rect 14730 599 14738 607
rect 15322 599 15330 607
rect 15434 599 15442 607
rect 16458 599 16466 607
rect 16714 599 16722 607
rect 17178 599 17186 607
rect 19536 600 19544 608
rect 19920 600 19928 608
rect 24944 600 24952 608
rect 25808 600 25816 608
rect 26864 600 26872 608
rect 27072 600 27080 608
rect 29456 597 29464 605
rect 504 579 512 587
rect 536 579 544 587
rect 680 579 688 587
rect 792 579 800 587
rect 840 579 848 587
rect 872 579 880 587
rect 1208 579 1216 587
rect 1256 579 1264 587
rect 1624 579 1632 587
rect 1736 579 1744 587
rect 1832 579 1840 587
rect 1944 579 1952 587
rect 2936 579 2944 587
rect 3080 579 3088 587
rect 3192 579 3200 587
rect 3992 579 4000 587
rect 4088 579 4096 587
rect 4280 579 4288 587
rect 4440 579 4448 587
rect 4472 579 4480 587
rect 4488 579 4496 587
rect 5810 573 5818 581
rect 5874 573 5882 581
rect 5890 573 5898 581
rect 6082 573 6090 581
rect 7090 573 7098 581
rect 7298 573 7306 581
rect 7314 573 7322 581
rect 7330 573 7338 581
rect 7586 573 7594 581
rect 9378 573 9386 581
rect 9474 573 9482 581
rect 10002 573 10010 581
rect 10370 573 10378 581
rect 10514 573 10522 581
rect 12106 579 12114 587
rect 12330 579 12338 587
rect 12698 579 12706 587
rect 14858 579 14866 587
rect 16506 579 16514 587
rect 16714 579 16722 587
rect 17066 579 17074 587
rect 17194 579 17202 587
rect 17386 579 17394 587
rect 19040 580 19048 588
rect 20512 580 20520 588
rect 20736 580 20744 588
rect 21264 580 21272 588
rect 23168 580 23176 588
rect 25376 580 25384 588
rect 25776 580 25784 588
rect 26016 580 26024 588
rect 26192 580 26200 588
rect 26560 580 26568 588
rect 26656 580 26664 588
rect 26880 580 26888 588
rect 2344 559 2352 567
rect 3256 559 3264 567
rect 3832 559 3840 567
rect 3880 559 3888 567
rect 3944 559 3952 567
rect 4168 559 4176 567
rect 6210 553 6218 561
rect 6226 553 6234 561
rect 6498 553 6506 561
rect 6594 553 6602 561
rect 6610 553 6618 561
rect 6754 553 6762 561
rect 6818 553 6826 561
rect 6946 553 6954 561
rect 7074 553 7082 561
rect 7090 553 7098 561
rect 7170 553 7178 561
rect 7218 553 7226 561
rect 8514 553 8522 561
rect 8674 553 8682 561
rect 8802 553 8810 561
rect 8994 553 9002 561
rect 9602 553 9610 561
rect 12826 559 12834 567
rect 13642 559 13650 567
rect 14682 559 14690 567
rect 15050 559 15058 567
rect 16042 559 16050 567
rect 16090 559 16098 567
rect 17242 559 17250 567
rect 17306 559 17314 567
rect 17434 559 17442 567
rect 21360 560 21368 568
rect 19524 548 19528 553
rect 20523 548 20530 553
rect 21188 548 21192 553
rect 22424 548 22428 553
rect 23462 548 23466 553
rect 27476 548 27485 553
rect 28102 548 28109 553
rect 600 539 608 547
rect 632 539 640 547
rect 696 539 704 547
rect 1352 539 1360 547
rect 1384 539 1392 547
rect 2008 539 2016 547
rect 2888 539 2896 547
rect 4488 539 4496 547
rect 5778 533 5786 541
rect 6050 533 6058 541
rect 6306 533 6314 541
rect 6370 533 6378 541
rect 7746 533 7754 541
rect 7810 533 7818 541
rect 7826 533 7834 541
rect 7842 533 7850 541
rect 8578 533 8586 541
rect 9650 533 9658 541
rect 9666 533 9674 541
rect 10146 533 10154 541
rect 10258 533 10266 541
rect 10802 533 10810 541
rect 11994 539 12002 547
rect 12090 539 12098 547
rect 12218 539 12226 547
rect 14170 539 14178 547
rect 14586 539 14594 547
rect 15290 539 15298 547
rect 16250 539 16258 547
rect 16474 539 16482 547
rect 16746 539 16754 547
rect 16794 539 16802 547
rect 16890 539 16898 547
rect 17098 539 17106 547
rect 17146 539 17154 547
rect 17434 539 17442 547
rect 19072 540 19080 548
rect 19488 540 19496 548
rect 19744 540 19752 548
rect 20096 540 20104 548
rect 20176 540 20184 548
rect 20736 540 20744 548
rect 23312 540 23320 548
rect 24496 540 24504 548
rect 24720 540 24728 548
rect 25152 540 25160 548
rect 25792 540 25800 548
rect 26000 540 26008 548
rect 27664 540 27672 548
rect 28304 540 28312 548
rect 776 519 784 527
rect 1080 519 1088 527
rect 1816 519 1824 527
rect 2696 519 2704 527
rect 2760 519 2768 527
rect 3736 519 3744 527
rect 6034 513 6042 521
rect 6354 513 6362 521
rect 9170 513 9178 521
rect 9410 513 9418 521
rect 9442 513 9450 521
rect 10402 513 10410 521
rect 10434 513 10442 521
rect 13194 519 13202 527
rect 14490 519 14498 527
rect 17226 519 17234 527
rect 18896 520 18904 528
rect 23472 520 23480 528
rect 25088 520 25096 528
rect 2504 499 2512 507
rect 3656 499 3664 507
rect 4184 499 4192 507
rect 6466 493 6474 501
rect 7362 493 7370 501
rect 7378 493 7386 501
rect 7410 493 7418 501
rect 8034 493 8042 501
rect 8178 493 8186 501
rect 8354 493 8362 501
rect 10210 493 10218 501
rect 13386 499 13394 507
rect 15114 499 15122 507
rect 22160 500 22168 508
rect 488 479 496 487
rect 616 479 624 487
rect 1176 479 1184 487
rect 1368 479 1376 487
rect 1608 479 1616 487
rect 2072 479 2080 487
rect 2088 479 2096 487
rect 2376 479 2384 487
rect 2584 479 2592 487
rect 3048 479 3056 487
rect 3064 479 3072 487
rect 3960 479 3968 487
rect 4632 479 4640 487
rect 5922 473 5930 481
rect 6834 473 6842 481
rect 7586 473 7594 481
rect 7762 473 7770 481
rect 8546 473 8554 481
rect 9010 473 9018 481
rect 9906 473 9914 481
rect 10018 473 10026 481
rect 10578 473 10586 481
rect 17418 479 17426 487
rect 20768 480 20776 488
rect 664 459 672 467
rect 1820 463 1844 467
rect 10882 453 10890 461
rect 13066 459 13074 467
rect 15386 459 15394 467
rect 23232 460 23240 468
rect 18784 450 18786 458
rect 18792 450 18794 458
rect 18990 450 19000 458
rect 19204 450 19214 458
rect 20234 450 20236 458
rect 20242 450 20244 458
rect 22104 450 22114 458
rect 23194 450 23198 458
rect 23202 450 23206 458
rect 23408 450 23412 458
rect 23416 450 23420 458
rect 26066 450 26068 458
rect 26074 450 26076 458
rect 27318 450 27320 458
rect 27326 450 27328 458
rect 27730 450 27732 458
rect 27738 450 27740 458
rect 28158 450 28160 458
rect 28166 450 28168 458
rect 8434 433 8442 441
rect 22256 440 22264 448
rect 712 419 720 427
rect 1448 419 1456 427
rect 1656 419 1664 427
rect 1768 419 1776 427
rect 1864 419 1872 427
rect 2152 419 2160 427
rect 2200 419 2208 427
rect 3144 419 3152 427
rect 3256 419 3264 427
rect 3560 419 3568 427
rect 3592 419 3600 427
rect 3832 419 3840 427
rect 3864 419 3872 427
rect 4280 419 4288 427
rect 4648 419 4656 427
rect 7554 413 7562 421
rect 7762 413 7770 421
rect 8098 413 8106 421
rect 8674 413 8682 421
rect 8898 413 8906 421
rect 9298 413 9306 421
rect 9570 413 9578 421
rect 9890 413 9898 421
rect 10050 413 10058 421
rect 14682 419 14690 427
rect 16202 419 16210 427
rect 16330 419 16338 427
rect 17114 419 17122 427
rect 19536 420 19544 428
rect 27632 420 27640 428
rect 27664 420 27672 428
rect 568 399 576 407
rect 776 399 784 407
rect 2136 399 2144 407
rect 2456 399 2464 407
rect 3480 399 3488 407
rect 3800 399 3808 407
rect 3912 399 3920 407
rect 4024 399 4032 407
rect 6546 393 6554 401
rect 6850 393 6858 401
rect 8834 393 8842 401
rect 14490 399 14498 407
rect 14794 399 14802 407
rect 16218 399 16226 407
rect 17354 399 17362 407
rect 27040 400 27048 408
rect 824 379 832 387
rect 1208 379 1216 387
rect 1224 379 1232 387
rect 1416 379 1424 387
rect 2216 379 2224 387
rect 2504 379 2512 387
rect 2984 379 2992 387
rect 3368 379 3376 387
rect 4184 379 4192 387
rect 6258 373 6266 381
rect 6322 373 6330 381
rect 6386 373 6394 381
rect 6962 373 6970 381
rect 7858 373 7866 381
rect 10034 373 10042 381
rect 10322 373 10330 381
rect 10354 373 10362 381
rect 10386 373 10394 381
rect 10738 373 10746 381
rect 12442 379 12450 387
rect 13306 379 13314 387
rect 13466 379 13474 387
rect 14666 379 14674 387
rect 14842 379 14850 387
rect 15898 379 15906 387
rect 17370 379 17378 387
rect 20128 380 20136 388
rect 22048 380 22056 388
rect 24752 380 24760 388
rect 26016 380 26024 388
rect 472 359 480 367
rect 1064 359 1072 367
rect 1368 359 1376 367
rect 1656 359 1664 367
rect 1672 359 1680 367
rect 2408 359 2416 367
rect 3176 359 3184 367
rect 3400 359 3408 367
rect 3624 359 3632 367
rect 3704 359 3712 367
rect 3848 359 3856 367
rect 4056 359 4064 367
rect 4120 359 4128 367
rect 5730 353 5738 361
rect 5762 353 5770 361
rect 5986 353 5994 361
rect 6146 353 6154 361
rect 6178 353 6186 361
rect 6530 353 6538 361
rect 6578 353 6586 361
rect 6658 353 6666 361
rect 6754 353 6762 361
rect 6786 353 6794 361
rect 6818 353 6826 361
rect 7058 353 7066 361
rect 7634 353 7642 361
rect 7906 353 7914 361
rect 7922 353 7930 361
rect 8290 353 8298 361
rect 8322 353 8330 361
rect 8354 353 8362 361
rect 8386 353 8394 361
rect 8434 353 8442 361
rect 8658 353 8666 361
rect 8722 353 8730 361
rect 9218 353 9226 361
rect 9410 353 9418 361
rect 9554 353 9562 361
rect 9682 353 9690 361
rect 9794 353 9802 361
rect 10130 353 10138 361
rect 10818 353 10826 361
rect 12010 359 12018 367
rect 12122 359 12130 367
rect 12362 359 12370 367
rect 12474 359 12482 367
rect 12538 359 12546 367
rect 13194 359 13202 367
rect 13338 359 13346 367
rect 14490 359 14498 367
rect 14602 359 14610 367
rect 14842 359 14850 367
rect 15770 359 15778 367
rect 15850 359 15858 367
rect 15946 359 15954 367
rect 16618 359 16626 367
rect 16666 359 16674 367
rect 16698 359 16706 367
rect 17210 359 17218 367
rect 17258 359 17266 367
rect 17274 359 17282 367
rect 19712 360 19720 368
rect 19760 360 19768 368
rect 19952 360 19960 368
rect 20304 360 20312 368
rect 21344 360 21352 368
rect 21552 360 21560 368
rect 22016 360 22024 368
rect 23248 360 23256 368
rect 23520 360 23528 368
rect 23712 360 23720 368
rect 23900 361 23910 366
rect 24496 360 24504 368
rect 24688 360 24696 368
rect 24944 360 24952 368
rect 25168 360 25176 368
rect 25936 360 25944 368
rect 26128 360 26136 368
rect 27440 360 27448 368
rect 27856 360 27864 368
rect 27872 360 27880 368
rect 28224 360 28232 368
rect 2008 339 2016 347
rect 2616 339 2624 347
rect 2664 339 2672 347
rect 4328 339 4336 347
rect 5810 333 5818 341
rect 5890 333 5898 341
rect 6050 333 6058 341
rect 6082 333 6090 341
rect 8818 333 8826 341
rect 9266 333 9274 341
rect 9330 333 9338 341
rect 9378 333 9386 341
rect 9586 333 9594 341
rect 9698 333 9706 341
rect 10050 333 10058 341
rect 10226 333 10234 341
rect 10466 333 10474 341
rect 10722 333 10730 341
rect 14218 339 14226 347
rect 15514 339 15522 347
rect 15706 339 15714 347
rect 15786 339 15794 347
rect 15818 339 15826 347
rect 15946 339 15954 347
rect 16042 339 16050 347
rect 16138 339 16146 347
rect 16458 339 16466 347
rect 16554 339 16562 347
rect 16794 339 16802 347
rect 16826 339 16834 347
rect 16906 339 16914 347
rect 17226 339 17234 347
rect 17274 339 17282 347
rect 21744 340 21752 348
rect 22688 340 22696 348
rect 23920 340 23928 348
rect 26560 340 26568 348
rect 27408 340 27416 348
rect 696 319 704 327
rect 744 319 752 327
rect 1112 319 1120 327
rect 1256 319 1264 327
rect 1592 319 1600 327
rect 3176 319 3184 327
rect 3224 319 3232 327
rect 3352 319 3360 327
rect 3384 319 3392 327
rect 4536 319 4544 327
rect 5762 313 5770 321
rect 5954 313 5962 321
rect 7074 313 7082 321
rect 7154 313 7162 321
rect 7186 313 7194 321
rect 7826 313 7834 321
rect 8098 313 8106 321
rect 8306 313 8314 321
rect 8578 313 8586 321
rect 8978 313 8986 321
rect 9890 313 9898 321
rect 10098 313 10106 321
rect 10130 313 10138 321
rect 10242 313 10250 321
rect 10274 313 10282 321
rect 10738 313 10746 321
rect 10770 313 10778 321
rect 12202 319 12210 327
rect 12282 319 12290 327
rect 12298 319 12306 327
rect 12554 319 12562 327
rect 12602 319 12610 327
rect 12682 319 12690 327
rect 12746 319 12754 327
rect 12858 319 12866 327
rect 13114 319 13122 327
rect 13258 319 13266 327
rect 13770 319 13778 327
rect 14234 319 14242 327
rect 14730 319 14738 327
rect 16026 319 16034 327
rect 16218 319 16226 327
rect 17306 319 17314 327
rect 18640 320 18648 328
rect 18736 320 18744 328
rect 18944 320 18952 328
rect 19696 320 19704 328
rect 19760 320 19768 328
rect 19776 320 19784 328
rect 20288 320 20296 328
rect 20816 320 20824 328
rect 21536 320 21544 328
rect 22064 320 22072 328
rect 22608 320 22616 328
rect 23024 320 23032 328
rect 23696 320 23704 328
rect 23728 320 23736 328
rect 24288 320 24296 328
rect 25760 320 25768 328
rect 27760 320 27768 328
rect 28304 320 28312 328
rect 29424 317 29432 325
rect 29488 317 29496 325
rect 728 299 736 307
rect 744 299 752 307
rect 808 299 816 307
rect 936 299 944 307
rect 1032 299 1040 307
rect 1112 299 1120 307
rect 1192 299 1200 307
rect 1528 299 1536 307
rect 1640 299 1648 307
rect 1720 299 1728 307
rect 1736 299 1744 307
rect 1752 299 1760 307
rect 1848 299 1856 307
rect 1880 299 1888 307
rect 1912 299 1920 307
rect 2008 299 2016 307
rect 2168 299 2176 307
rect 2184 299 2192 307
rect 2264 299 2272 307
rect 2344 299 2352 307
rect 2456 299 2464 307
rect 2568 299 2576 307
rect 2584 299 2592 307
rect 2760 299 2768 307
rect 2840 299 2848 307
rect 2856 299 2864 307
rect 2936 299 2944 307
rect 2952 299 2960 307
rect 3128 299 3136 307
rect 3240 299 3248 307
rect 3320 299 3328 307
rect 3576 299 3584 307
rect 3608 299 3616 307
rect 3880 299 3888 307
rect 3896 299 3904 307
rect 4008 299 4016 307
rect 4040 299 4048 307
rect 4152 299 4160 307
rect 4296 299 4304 307
rect 4312 299 4320 307
rect 4360 299 4368 307
rect 4488 299 4496 307
rect 4552 299 4560 307
rect 4632 299 4640 307
rect 5794 293 5802 301
rect 5906 293 5914 301
rect 6050 293 6058 301
rect 6370 293 6378 301
rect 6562 293 6570 301
rect 7202 293 7210 301
rect 7682 293 7690 301
rect 7746 293 7754 301
rect 7970 293 7978 301
rect 7986 293 7994 301
rect 8258 293 8266 301
rect 8322 293 8330 301
rect 8578 293 8586 301
rect 8610 293 8618 301
rect 8626 293 8634 301
rect 8658 293 8666 301
rect 8738 293 8746 301
rect 9042 293 9050 301
rect 9058 293 9066 301
rect 9186 293 9194 301
rect 9586 293 9594 301
rect 10018 293 10026 301
rect 10066 293 10074 301
rect 10194 293 10202 301
rect 10322 293 10330 301
rect 10546 293 10554 301
rect 10562 293 10570 301
rect 10658 293 10666 301
rect 10786 293 10794 301
rect 13530 299 13538 307
rect 13706 299 13714 307
rect 15066 299 15074 307
rect 15242 299 15250 307
rect 16026 299 16034 307
rect 16858 299 16866 307
rect 2040 279 2048 287
rect 2504 279 2512 287
rect 2792 279 2800 287
rect 3736 279 3744 287
rect 4056 279 4064 287
rect 6002 273 6010 281
rect 6194 273 6202 281
rect 6514 273 6522 281
rect 7170 273 7178 281
rect 7218 273 7226 281
rect 7666 273 7674 281
rect 7970 273 7978 281
rect 9634 273 9642 281
rect 10530 273 10538 281
rect 10802 273 10810 281
rect 12106 279 12114 287
rect 13578 279 13586 287
rect 13722 279 13730 287
rect 13898 279 13906 287
rect 14154 279 14162 287
rect 14346 279 14354 287
rect 15546 279 15554 287
rect 21184 280 21192 288
rect 22832 280 22840 288
rect 24912 280 24920 288
rect 25344 280 25352 288
rect 27184 280 27192 288
rect 27216 280 27224 288
rect 28656 280 28664 288
rect 1416 259 1424 267
rect 2840 259 2848 267
rect 3416 259 3424 267
rect 4152 259 4160 267
rect 4216 259 4224 267
rect 6674 253 6682 261
rect 6690 253 6698 261
rect 7442 253 7450 261
rect 7490 253 7498 261
rect 7522 253 7530 261
rect 8114 253 8122 261
rect 8162 253 8170 261
rect 8450 253 8458 261
rect 8610 253 8618 261
rect 8642 253 8650 261
rect 8722 253 8730 261
rect 8754 253 8762 261
rect 9410 253 9418 261
rect 9506 253 9514 261
rect 9522 253 9530 261
rect 9618 253 9626 261
rect 15258 259 15266 267
rect 15306 259 15314 267
rect 15610 259 15618 267
rect 19536 260 19544 268
rect 22944 260 22952 268
rect 24080 260 24088 268
rect 24320 260 24328 268
rect 29396 267 29408 275
rect 29428 267 29440 275
rect 29444 267 29448 275
rect 29460 267 29472 275
rect 29488 267 29504 275
rect 29512 267 29544 275
rect 29552 267 29568 275
rect 29576 267 29588 275
rect 29592 267 29596 275
rect 18542 252 18544 260
rect 18702 250 18710 258
rect 18852 250 18858 258
rect 18916 250 18924 258
rect 19066 250 19072 258
rect 19130 250 19144 258
rect 19494 250 19500 258
rect 19740 250 19754 258
rect 20264 250 20278 258
rect 20318 250 20326 258
rect 20676 250 20690 258
rect 20730 250 20738 258
rect 20818 250 20824 258
rect 20826 250 20832 258
rect 21024 250 21038 258
rect 21124 250 21136 258
rect 21634 250 21642 258
rect 21848 250 21856 258
rect 22178 250 22190 258
rect 22276 250 22284 258
rect 22380 250 22382 258
rect 22594 250 22596 258
rect 23116 250 23124 258
rect 23330 250 23338 258
rect 23544 250 23558 258
rect 23686 250 23692 258
rect 23694 250 23700 258
rect 23844 250 23850 258
rect 23892 250 23906 258
rect 24042 250 24048 258
rect 24098 250 24104 258
rect 24106 250 24112 258
rect 24256 250 24262 258
rect 24724 250 24730 258
rect 24732 250 24738 258
rect 24882 250 24888 258
rect 24930 250 24944 258
rect 25358 250 25372 258
rect 25556 250 25564 258
rect 25706 250 25712 258
rect 25898 250 25912 258
rect 25952 250 25960 258
rect 26096 250 26110 258
rect 26402 250 26406 258
rect 26492 250 26500 258
rect 26578 250 26586 258
rect 26728 250 26734 258
rect 26792 250 26800 258
rect 26942 250 26948 258
rect 27006 250 27014 258
rect 27156 250 27162 258
rect 27542 252 27544 260
rect 27686 252 27688 260
rect 1960 239 1968 247
rect 1992 239 2000 247
rect 2312 239 2320 247
rect 3096 239 3104 247
rect 4424 239 4432 247
rect 6706 233 6714 241
rect 6914 233 6922 241
rect 8194 233 8202 241
rect 8290 233 8298 241
rect 8594 233 8602 241
rect 8642 233 8650 241
rect 8994 233 9002 241
rect 9826 233 9834 241
rect 10130 233 10138 241
rect 10578 233 10586 241
rect 12938 239 12946 247
rect 15498 239 15506 247
rect 28032 240 28040 248
rect 424 219 432 227
rect 1784 219 1792 227
rect 2024 219 2032 227
rect 2072 219 2080 227
rect 2184 219 2192 227
rect 2232 219 2240 227
rect 2248 219 2256 227
rect 2296 219 2304 227
rect 2344 219 2352 227
rect 2456 219 2464 227
rect 2504 219 2512 227
rect 3048 219 3056 227
rect 3160 219 3168 227
rect 3992 219 4000 227
rect 4184 219 4192 227
rect 4520 219 4528 227
rect 4600 219 4608 227
rect 4616 219 4624 227
rect 6018 213 6026 221
rect 6322 213 6330 221
rect 6466 213 6474 221
rect 6690 213 6698 221
rect 6914 213 6922 221
rect 6978 213 6986 221
rect 7330 213 7338 221
rect 7490 213 7498 221
rect 7826 213 7834 221
rect 7954 213 7962 221
rect 8130 213 8138 221
rect 8994 213 9002 221
rect 9074 213 9082 221
rect 9314 213 9322 221
rect 9858 213 9866 221
rect 10130 213 10138 221
rect 12490 219 12498 227
rect 14170 219 14178 227
rect 14874 219 14882 227
rect 14922 219 14930 227
rect 15642 219 15650 227
rect 15738 219 15746 227
rect 17114 219 17122 227
rect 17290 219 17298 227
rect 17562 219 17570 227
rect 18656 220 18664 228
rect 19280 220 19288 228
rect 20688 220 20696 228
rect 24640 220 24648 228
rect 26112 220 26120 228
rect 26528 220 26536 228
rect 27616 220 27624 228
rect 28416 220 28424 228
rect 504 199 512 207
rect 584 199 592 207
rect 680 199 688 207
rect 712 199 720 207
rect 792 199 800 207
rect 840 199 848 207
rect 856 199 864 207
rect 952 199 960 207
rect 1032 199 1040 207
rect 1048 199 1056 207
rect 1144 199 1152 207
rect 1272 199 1280 207
rect 1288 199 1296 207
rect 1512 199 1520 207
rect 1624 199 1632 207
rect 1704 199 1712 207
rect 1800 199 1808 207
rect 1832 199 1840 207
rect 1960 199 1968 207
rect 2040 199 2048 207
rect 2120 199 2128 207
rect 2248 199 2256 207
rect 2280 199 2288 207
rect 2312 199 2320 207
rect 2440 199 2448 207
rect 2456 199 2464 207
rect 2536 199 2544 207
rect 2568 199 2576 207
rect 2664 199 2672 207
rect 2872 199 2880 207
rect 2936 199 2944 207
rect 3000 199 3008 207
rect 3032 199 3040 207
rect 3112 199 3120 207
rect 3256 199 3264 207
rect 3320 199 3328 207
rect 3352 199 3360 207
rect 3368 199 3376 207
rect 3416 199 3424 207
rect 3656 199 3664 207
rect 3672 199 3680 207
rect 3768 199 3776 207
rect 3832 199 3840 207
rect 3864 199 3872 207
rect 3928 199 3936 207
rect 3960 199 3968 207
rect 4024 199 4032 207
rect 4168 199 4176 207
rect 4200 199 4208 207
rect 4216 199 4224 207
rect 4248 199 4256 207
rect 4264 199 4272 207
rect 4344 199 4352 207
rect 4360 199 4368 207
rect 4440 199 4448 207
rect 4536 199 4544 207
rect 5986 193 5994 201
rect 6146 193 6154 201
rect 6162 193 6170 201
rect 6178 193 6186 201
rect 6274 193 6282 201
rect 6770 193 6778 201
rect 6802 193 6810 201
rect 6882 193 6890 201
rect 6930 193 6938 201
rect 6946 193 6954 201
rect 7058 193 7066 201
rect 7282 193 7290 201
rect 7810 193 7818 201
rect 7922 193 7930 201
rect 7938 193 7946 201
rect 8354 193 8362 201
rect 8370 193 8378 201
rect 8498 193 8506 201
rect 8562 193 8570 201
rect 9154 193 9162 201
rect 9458 193 9466 201
rect 9570 193 9578 201
rect 9586 193 9594 201
rect 9682 193 9690 201
rect 9762 193 9770 201
rect 9842 193 9850 201
rect 10050 193 10058 201
rect 10146 193 10154 201
rect 10162 193 10170 201
rect 10242 193 10250 201
rect 10482 193 10490 201
rect 10546 193 10554 201
rect 10562 193 10570 201
rect 10706 193 10714 201
rect 10786 193 10794 201
rect 15066 199 15074 207
rect 15290 199 15298 207
rect 15386 199 15394 207
rect 16970 199 16978 207
rect 17306 199 17314 207
rect 21728 200 21736 208
rect 24080 200 24088 208
rect 24496 200 24504 208
rect 24704 200 24712 208
rect 24720 200 24728 208
rect 28640 200 28648 208
rect 504 179 512 187
rect 552 179 560 187
rect 1192 179 1200 187
rect 1544 179 1552 187
rect 1560 179 1568 187
rect 1608 179 1616 187
rect 2216 179 2224 187
rect 2248 179 2256 187
rect 2520 179 2528 187
rect 2712 179 2720 187
rect 2968 179 2976 187
rect 3448 179 3456 187
rect 3560 179 3568 187
rect 3592 179 3600 187
rect 3880 179 3888 187
rect 4104 179 4112 187
rect 5842 173 5850 181
rect 5906 173 5914 181
rect 7170 173 7178 181
rect 7266 173 7274 181
rect 7586 173 7594 181
rect 9138 173 9146 181
rect 9618 173 9626 181
rect 10418 173 10426 181
rect 10626 173 10634 181
rect 12026 179 12034 187
rect 12202 179 12210 187
rect 12890 179 12898 187
rect 12954 179 12962 187
rect 13146 179 13154 187
rect 13194 179 13202 187
rect 13290 179 13298 187
rect 13306 179 13314 187
rect 13754 179 13762 187
rect 13866 179 13874 187
rect 13930 179 13938 187
rect 14154 179 14162 187
rect 14218 179 14226 187
rect 14730 179 14738 187
rect 14794 179 14802 187
rect 15594 179 15602 187
rect 16426 179 16434 187
rect 16954 179 16962 187
rect 16986 179 16994 187
rect 19280 180 19288 188
rect 19424 180 19432 188
rect 19456 180 19464 188
rect 19504 180 19512 188
rect 19872 180 19880 188
rect 20240 180 20248 188
rect 20656 180 20664 188
rect 21040 180 21048 188
rect 21456 180 21464 188
rect 22080 180 22088 188
rect 22800 180 22808 188
rect 23664 180 23672 188
rect 23872 180 23880 188
rect 27216 180 27224 188
rect 27440 180 27448 188
rect 27968 180 27976 188
rect 28176 180 28184 188
rect 28608 180 28616 188
rect 952 159 960 167
rect 2968 159 2976 167
rect 3864 159 3872 167
rect 4088 159 4096 167
rect 4600 159 4608 167
rect 5906 153 5914 161
rect 5938 153 5946 161
rect 7378 153 7386 161
rect 8274 153 8282 161
rect 8450 153 8458 161
rect 9618 153 9626 161
rect 9762 153 9770 161
rect 9794 153 9802 161
rect 10370 153 10378 161
rect 10450 153 10458 161
rect 10610 153 10618 161
rect 10866 153 10874 161
rect 12122 159 12130 167
rect 12426 159 12434 167
rect 12634 159 12642 167
rect 12666 159 12674 167
rect 12682 159 12690 167
rect 14922 159 14930 167
rect 15322 159 15330 167
rect 16570 159 16578 167
rect 16586 159 16594 167
rect 16730 159 16738 167
rect 16794 159 16802 167
rect 16826 159 16834 167
rect 16922 159 16930 167
rect 17002 159 17010 167
rect 19104 160 19112 168
rect 28224 160 28232 168
rect 29408 157 29416 165
rect 21068 148 21072 153
rect 22788 148 22792 153
rect 23858 148 23862 153
rect 27771 148 27780 153
rect 456 139 464 147
rect 536 139 544 147
rect 808 139 816 147
rect 1464 139 1472 147
rect 1512 139 1520 147
rect 1528 139 1536 147
rect 1976 139 1984 147
rect 2168 139 2176 147
rect 2408 139 2416 147
rect 2616 139 2624 147
rect 2664 139 2672 147
rect 3208 139 3216 147
rect 3368 139 3376 147
rect 3448 139 3456 147
rect 3496 139 3504 147
rect 3576 139 3584 147
rect 4232 139 4240 147
rect 4264 139 4272 147
rect 4552 139 4560 147
rect 5938 133 5946 141
rect 6098 133 6106 141
rect 7170 133 7178 141
rect 7282 133 7290 141
rect 7522 133 7530 141
rect 7922 133 7930 141
rect 9250 133 9258 141
rect 9314 133 9322 141
rect 9362 133 9370 141
rect 9778 133 9786 141
rect 10194 133 10202 141
rect 10226 133 10234 141
rect 10274 133 10282 141
rect 10306 133 10314 141
rect 12506 139 12514 147
rect 12906 139 12914 147
rect 12954 139 12962 147
rect 13050 139 13058 147
rect 13274 139 13282 147
rect 13354 139 13362 147
rect 13386 139 13394 147
rect 13530 139 13538 147
rect 13546 139 13554 147
rect 13658 139 13666 147
rect 14042 139 14050 147
rect 14362 139 14370 147
rect 15114 139 15122 147
rect 16010 139 16018 147
rect 16074 139 16082 147
rect 16154 139 16162 147
rect 16266 139 16274 147
rect 16346 139 16354 147
rect 16394 139 16402 147
rect 16506 139 16514 147
rect 16538 139 16546 147
rect 16634 139 16642 147
rect 17386 139 17394 147
rect 19040 140 19048 148
rect 21888 140 21896 148
rect 22512 140 22520 148
rect 22720 140 22728 148
rect 22800 140 22808 148
rect 23584 140 23592 148
rect 24272 140 24280 148
rect 24496 140 24504 148
rect 25088 140 25096 148
rect 25328 140 25336 148
rect 25504 140 25512 148
rect 1304 119 1312 127
rect 1576 119 1584 127
rect 1624 119 1632 127
rect 1944 119 1952 127
rect 2216 119 2224 127
rect 2424 119 2432 127
rect 2568 119 2576 127
rect 6194 113 6202 121
rect 6498 113 6506 121
rect 6530 113 6538 121
rect 8258 113 8266 121
rect 8578 113 8586 121
rect 8626 113 8634 121
rect 8914 113 8922 121
rect 8978 113 8986 121
rect 9490 113 9498 121
rect 9746 113 9754 121
rect 13418 119 13426 127
rect 13434 119 13442 127
rect 13898 119 13906 127
rect 15434 119 15442 127
rect 15626 119 15634 127
rect 15818 119 15826 127
rect 19680 120 19688 128
rect 3464 99 3472 107
rect 8866 93 8874 101
rect 16602 99 16610 107
rect 16538 79 16546 87
rect 3288 59 3296 67
rect 21744 60 21752 68
rect 22864 60 22872 68
use secLibDualRail  secLibDualRail_0
timestamp 1602346068
transform 1 0 29332 0 1 61
box -208 -43 15580 11283
use dualRail  dualRail_0
timestamp 1600868604
transform 1 0 11982 0 1 43
box -412 -43 5994 4083
use dualRailAS  dualRailAS_0
timestamp 1600868604
transform 1 0 5718 0 1 37
box -408 -43 5626 3740
use singleRail  singleRail_0
timestamp 1600868604
transform 1 0 412 0 1 43
box -412 -43 4682 3083
use pDualRail  pDualRail_0
timestamp 1600868604
transform 1 0 18452 0 1 44
box -208 -43 10406 7283
<< end >>
