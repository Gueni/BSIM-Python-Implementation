*** TEST 005 partitioning ***
*
* ngSPICE test for PLS experiments
*
* AES SBOX PLS test init file generator - protected dualRail SBOX area illuminated
*
* Author: Jan Belohoubek, 08/2020
* jan.belohoubek@fit.cvut.cz
*
* https://users.fit.cvut.cz/~belohja4/
*
*
* **************************************

.include ../../models.lib
.include ../../tsmc180nmcmos.lib
.include secLibDualRail.spice

* **************************************
* --- Test ---
* **************************************

* --- Settings
.param showPlots = 0
.param writeFile = 1
.param run_inputSet = 0

* redefine defaults ...
.include test00X_settings.inc

.csparam showPlots = {showPlots}
.csparam writeFile = {writeFile}
.csparam run_inputSet = {run_inputSet}

.global showPlots writeFile run_inputSet

* --- End of Settins

Vtrig LaserTrig 0 0 PWL(0ns 0V 40ns 0V 41ns SUPP)

.param beamDistanceTop = 0
.param beamDistanceBot = 0

.global LaserTrig beamDistanceTop beamDistanceBot

* --- inputs
Vvin0 INPUT_0 0 0 PWL(0ns 0V 5ns  0V 7ns  0V)
Vvin1 INPUT_1 0 0 PWL(0ns 0V 6ns  0V 8ns  0V)
Vvin2 INPUT_2 0 0 PWL(0ns 0V 7ns  0V 9ns  0V)
Vvin3 INPUT_3 0 0 PWL(0ns 0V 8ns  0V 10ns 0V)
Vvin4 INPUT_4 0 0 PWL(0ns 0V 9ns  0V 11ns 0V)
Vvin5 INPUT_5 0 0 PWL(0ns 0V 10ns 0V 12ns 0V)
Vvin6 INPUT_6 0 0 PWL(0ns 0V 11ns 0V 13ns 0V)
Vvin7 INPUT_7 0 0 PWL(0ns 0V 12ns 0V 14ns 0V)

Vvin0D D_INPUT_0 0 0 PWL(0ns 0V 5ns  0V 7ns  0V)
Vvin1D D_INPUT_1 0 0 PWL(0ns 0V 6ns  0V 8ns  0V)
Vvin2D D_INPUT_2 0 0 PWL(0ns 0V 7ns  0V 9ns  0V)
Vvin3D D_INPUT_3 0 0 PWL(0ns 0V 8ns  0V 10ns 0V)
Vvin4D D_INPUT_4 0 0 PWL(0ns 0V 9ns  0V 11ns 0V)
Vvin5D D_INPUT_5 0 0 PWL(0ns 0V 10ns 0V 12ns 0V)
Vvin6D D_INPUT_6 0 0 PWL(0ns 0V 11ns 0V 13ns 0V)
Vvin7D D_INPUT_7 0 0 PWL(0ns 0V 12ns 0V 14ns 0V)


* --- outputs
C0 VSS GATE_222 10fF
C1 VSS GATE_366 10fF
C2 VSS GATE_479 10fF
C3 VSS GATE_579 10fF
C4 VSS GATE_662 10fF
C5 VSS GATE_741 10fF
C6 VSS GATE_811 10fF
C7 VSS GATE_865 10fF

C0d VSS D_GATE_222 10fF
C1d VSS D_GATE_366 10fF
C2d VSS D_GATE_479 10fF
C3d VSS D_GATE_579 10fF
C4d VSS D_GATE_662 10fF
C5d VSS D_GATE_741 10fF
C6d VSS D_GATE_811 10fF
C7d VSS D_GATE_865 10fF

* --- circuit layout model

Xsbox1 
+ INVX1_1624/A INVX1_732/A INVX1_957/A INVX1_731/A INVX1_1150/A INVX1_1726/A INVX1_1149/A INVX1_1447/A INVX1_1477/A INVX1_1725/A INVX1_1623/A INVX1_1448/A INVX1_1315/A INVX1_1724/A INVX1_1723/A INVX1_1136/A INVX1_1135/A INVX1_1474/A INVX1_958/A INVX1_1461/A INVX1_954/A INVX1_953/A INVX1_1316/A INVX1_1722/A INVX1_1721/A INVX1_428/A INVX1_427/A INVX1_730/A INVX1_729/A INVX1_1449/A INVX1_1472/A INVX1_1471/A INVX1_1473/A INVX1_1143/A INVX1_436/A INVX1_1320/A INVX1_435/A INVX1_1319/A INVX1_1142/A INVX1_1141/A INVX1_937/A INVX1_938/A INVX1_1144/A INVX1_1124/A INVX1_1123/A INVX1_1125/A INVX1_411/A INVX1_409/A INVX1_412/A INVX1_1450/A INVX1_1138/A 
+ INVX1_1137/A INVX1_1462/A INVX1_1126/A INVX1_410/A INVX1_1322/A INVX1_1321/A INVX1_1478/A INVX1_442/A INVX1_441/A INVX1_1548/Y INVX1_1547/Y INVX1_1019/Y INVX1_1020/Y INVX1_909/Y INVX1_910/Y INVX1_439/Y INVX1_440/Y INVX1_1308/Y INVX1_1307/Y INVX1_932/Y INVX1_931/Y INVX1_1127/Y INVX1_1128/Y INVX1_488/Y INVX1_487/Y INVX1_1111/Y INVX1_1112/Y INVX1_281/Y INVX1_282/Y INVX1_935/Y INVX1_936/Y INVX1_1120/Y INVX1_1119/Y INVX1_1310/Y INVX1_1309/Y INVX1_434/Y INVX1_433/Y INVX1_1465/Y INVX1_1466/Y 
+ INVX1_1470/Y INVX1_1469/Y INVX1_681/Y INVX1_682/Y INVX1_1299/Y INVX1_1300/Y INVX1_1289/Y INVX1_1290/Y INVX1_727/Y INVX1_728/Y INVX1_363/Y INVX1_364/Y INVX1_413/Y INVX1_414/Y INVX1_1719/Y INVX1_1720/Y INVX1_939/Y INVX1_940/Y INVX1_703/Y INVX1_704/Y INVX1_1705/Y INVX1_1706/Y INVX1_1132/Y INVX1_1131/Y INVX1_399/Y INVX1_400/Y INVX1_1715/Y INVX1_1716/Y INVX1_1702/Y INVX1_1701/Y INVX1_1101/Y INVX1_1102/Y INVX1_1621/Y INVX1_1622/Y INVX1_1714/Y INVX1_1713/Y INVX1_1146/Y INVX1_1145/Y INVX1_726/Y INVX1_725/Y INVX1_439/A INVX1_440/A INVX1_1310/A INVX1_1309/A INVX1_1465/A INVX1_1466/A INVX1_727/A INVX1_728/A INVX1_1621/A INVX1_1622/A INVX1_726/A 
+ INVX1_725/A NOR3X1_439/A NOR3X1_439/B NOR3X1_439/C NOR3X1_440/A NOR3X1_440/B NOR3X1_440/C NOR3X1_1310/A NOR3X1_1310/B NOR3X1_1310/C NOR3X1_1309/A NOR3X1_1309/B NOR3X1_1309/C NOR3X1_1465/A NOR3X1_1465/B NOR3X1_1465/C NOR3X1_1466/A NOR3X1_1466/B NOR3X1_1466/C NOR3X1_727/A NOR3X1_727/B NOR3X1_727/C NOR3X1_728/A NOR3X1_728/B NOR3X1_728/C NOR3X1_1621/A NOR3X1_1621/B NOR3X1_1621/C NOR3X1_1622/A NOR3X1_1622/B NOR3X1_1622/C NOR3X1_726/A NOR3X1_726/B NOR3X1_726/C NOR3X1_725/A NOR3X1_725/B NOR3X1_725/C INVX1_424/Y INVX1_426/Y INVX1_425/Y INVX1_423/Y INVX1_1297/Y INVX1_1295/Y INVX1_1298/Y INVX1_1296/Y INVX1_1444/Y INVX1_1446/Y INVX1_1445/Y INVX1_1443/Y INVX1_714/Y INVX1_716/Y 
+ INVX1_715/Y INVX1_713/Y INVX1_1614/Y INVX1_1616/Y INVX1_1615/Y INVX1_1613/Y INVX1_719/Y INVX1_717/Y INVX1_720/Y INVX1_718/Y INVX1_424/A INVX1_423/A INVX1_716/A INVX1_715/A INVX1_1614/A INVX1_1616/A INVX1_1615/A INVX1_1613/A NOR3X1_424/A NOR3X1_424/B NOR3X1_424/C NOR3X1_423/A NOR3X1_423/B NOR3X1_423/C NOR3X1_716/A NOR3X1_716/B NOR3X1_716/C NOR3X1_715/A NOR3X1_715/B NOR3X1_715/C NOR3X1_1614/A NOR3X1_1614/B NOR3X1_1614/C NOR3X1_1616/A NOR3X1_1616/B NOR3X1_1616/C NOR3X1_1615/A NOR3X1_1615/B NOR3X1_1615/C NOR3X1_1613/A NOR3X1_1613/B NOR3X1_1613/C INVX1_421/Y INVX1_422/Y INVX1_701/Y INVX1_699/Y INVX1_702/Y INVX1_700/Y INVX1_1611/Y INVX1_1609/Y INVX1_1612/Y 
+ INVX1_1610/Y INVX1_1607/Y INVX1_1605/Y INVX1_1608/Y INVX1_1606/Y INVX1_1607/A INVX1_1605/A INVX1_1608/A INVX1_1606/A NOR3X1_1607/A NOR3X1_1607/B NOR3X1_1607/C NOR3X1_1605/A NOR3X1_1605/B NOR3X1_1605/C NOR3X1_1608/A NOR3X1_1608/B NOR3X1_1608/C NOR3X1_1606/A NOR3X1_1606/B NOR3X1_1606/C INVX1_1588/Y INVX1_1590/Y INVX1_1589/Y INVX1_1587/Y INVX1_1592/Y INVX1_1594/Y INVX1_1593/Y INVX1_1591/Y INVX1_638/Y INVX1_637/Y INVX1_232/Y INVX1_231/Y INVX1_70/Y INVX1_69/Y INVX1_1077/Y INVX1_1078/Y INVX1_807/Y INVX1_808/Y 
+ VSS VDD 
+ GATE_222 GATE_366 GATE_479 GATE_579 GATE_662 GATE_741 GATE_811 GATE_865 D_GATE_222 D_GATE_366 D_GATE_479 D_GATE_579 D_GATE_662 D_GATE_741 D_GATE_811 D_GATE_865 
+ AES_SBOX_4

.include outputs_3.plw

* **************************************
* --- Simulation Settings ---
* **************************************

.param SIM_LEN = 50ns
.csparam SIM_LEN = {SIM_LEN}

.tran 0.1ns 'SIM_LEN'
.param SIMSTEP = 'SIM_LEN/0.1ns'
.csparam SIMSTEP = {SIMSTEP}

* **************************************
* --- Simulation Control ---
* **************************************

.control
    .include ../inputsD.inc

    run
    
    if ('writeFile' > 0)   
      wrdata ivdd_4.out i(vvdd)
      wrdata ivss_4.out i(vvss)
      *snsave sim_4.snap
    end
    
    set wr_vecnames
    set wr_singlescale
    wrdata outputs_4.out V("GATE_222") V("GATE_366") V("GATE_479") V("GATE_579") V("GATE_662") V("GATE_741") V("GATE_811") V("GATE_865") V("D_GATE_222") V("D_GATE_366") V("D_GATE_479") V("D_GATE_579") V("D_GATE_662") V("D_GATE_741") V("D_GATE_811") V("D_GATE_865") 
    
    if ('showPlots' < 1)
        quit
    end
       
.endc

.end
