* SUBCKT HEAD: NAME;  INPUTS; POWER; OUTPUTS
.subckt AES_SBOX_0
+ INPUT_0 INPUT_1 INPUT_2 INPUT_3 INPUT_4 INPUT_5 INPUT_6 INPUT_7 D_INPUT_0 D_INPUT_1 D_INPUT_2 D_INPUT_3 D_INPUT_4 D_INPUT_5 D_INPUT_6 D_INPUT_7 
+ VSS VDD 
+ OR2X1_LOC_515/Y OR2X1_LOC_751/A OR2X1_LOC_334/A OR2X1_LOC_836/A OR2X1_LOC_240/A OR2X1_LOC_461/Y AND2X1_LOC_809/A AND2X1_LOC_276/Y OR2X1_LOC_100/Y OR2X1_LOC_516/B AND2X1_LOC_729/B OR2X1_LOC_527/Y OR2X1_LOC_111/Y OR2X1_LOC_323/Y AND2X1_LOC_155/Y OR2X1_LOC_273/Y OR2X1_LOC_433/Y OR2X1_LOC_743/Y OR2X1_LOC_409/B AND2X1_LOC_458/Y OR2X1_LOC_519/Y OR2X1_LOC_692/Y OR2X1_LOC_599/A OR2X1_LOC_763/Y OR2X1_LOC_48/Y OR2X1_LOC_406/A OR2X1_LOC_511/Y OR2X1_LOC_604/A OR2X1_LOC_235/B OR2X1_LOC_246/Y OR2X1_LOC_74/A OR2X1_LOC_13/B OR2X1_LOC_16/A OR2X1_LOC_287/B OR2X1_LOC_637/B OR2X1_LOC_294/Y OR2X1_LOC_415/Y OR2X1_LOC_631/A OR2X1_LOC_598/Y OR2X1_LOC_398/Y OR2X1_LOC_309/Y OR2X1_LOC_283/Y OR2X1_LOC_488/Y OR2X1_LOC_289/Y OR2X1_LOC_417/Y OR2X1_LOC_226/Y OR2X1_LOC_815/A OR2X1_LOC_121/Y OR2X1_LOC_831/A OR2X1_LOC_543/A OR2X1_LOC_606/Y 
+ OR2X1_LOC_302/A OR2X1_LOC_450/B AND2X1_LOC_847/Y AND2X1_LOC_91/B OR2X1_LOC_611/Y AND2X1_LOC_56/B OR2X1_LOC_78/A OR2X1_LOC_532/B OR2X1_LOC_96/B OR2X1_LOC_71/A OR2X1_LOC_535/A OR2X1_LOC_195/A OR2X1_LOC_296/Y OR2X1_LOC_138/A OR2X1_LOC_541/A OR2X1_LOC_838/B OR2X1_LOC_506/A OR2X1_LOC_378/Y OR2X1_LOC_98/B OR2X1_LOC_389/A OR2X1_LOC_448/A OR2X1_LOC_630/B OR2X1_LOC_144/Y OR2X1_LOC_306/Y OR2X1_LOC_503/A OR2X1_LOC_696/Y OR2X1_LOC_588/Y OR2X1_LOC_376/Y OR2X1_LOC_322/Y OR2X1_LOC_164/Y OR2X1_LOC_673/A OR2X1_LOC_693/Y AND2X1_LOC_377/Y OR2X1_LOC_748/A OR2X1_LOC_83/A OR2X1_LOC_89/A OR2X1_LOC_45/B OR2X1_LOC_52/B OR2X1_LOC_619/Y OR2X1_LOC_151/A OR2X1_LOC_185/A AND2X1_LOC_86/B OR2X1_LOC_160/A OR2X1_LOC_154/A OR2X1_LOC_130/A OR2X1_LOC_266/A OR2X1_LOC_634/A OR2X1_LOC_541/B OR2X1_LOC_633/A OR2X1_LOC_777/B OR2X1_LOC_549/A 
+ OR2X1_LOC_391/B OR2X1_LOC_387/Y OR2X1_LOC_597/A OR2X1_LOC_329/Y OR2X1_LOC_421/Y OR2X1_LOC_304/Y OR2X1_LOC_56/Y OR2X1_LOC_158/A OR2X1_LOC_70/Y OR2X1_LOC_3/Y OR2X1_LOC_40/Y OR2X1_LOC_694/Y OR2X1_LOC_426/Y AND2X1_LOC_51/Y AND2X1_LOC_31/Y AND2X1_LOC_44/Y AND2X1_LOC_47/Y OR2X1_LOC_790/B OR2X1_LOC_635/A OR2X1_LOC_769/B OR2X1_LOC_409/Y OR2X1_LOC_430/Y OR2X1_LOC_51/Y OR2X1_LOC_95/Y OR2X1_LOC_64/Y OR2X1_LOC_375/A AND2X1_LOC_36/Y AND2X1_LOC_18/Y OR2X1_LOC_809/B OR2X1_LOC_513/Y OR2X1_LOC_473/A AND2X1_LOC_101/B OR2X1_LOC_600/A OR2X1_LOC_744/A OR2X1_LOC_557/A AND2X1_LOC_19/Y OR2X1_LOC_7/A OR2X1_LOC_344/A OR2X1_LOC_748/Y OR2X1_LOC_589/A OR2X1_LOC_161/B OR2X1_LOC_80/Y OR2X1_LOC_87/A OR2X1_LOC_32/B OR2X1_LOC_269/B OR2X1_LOC_291/Y OR2X1_LOC_824/Y OR2X1_LOC_234/Y AND2X1_LOC_462/B OR2X1_LOC_691/Y OR2X1_LOC_325/A 
+ OR2X1_LOC_547/B OR2X1_LOC_112/A OR2X1_LOC_516/A OR2X1_LOC_750/Y OR2X1_LOC_814/Y OR2X1_LOC_335/B OR2X1_LOC_286/B OR2X1_LOC_489/A OR2X1_LOC_333/A OR2X1_LOC_446/B OR2X1_LOC_227/A OR2X1_LOC_427/A AND2X1_LOC_81/B AND2X1_LOC_82/Y OR2X1_LOC_87/B OR2X1_LOC_428/A OR2X1_LOC_382/Y OR2X1_LOC_39/A OR2X1_LOC_848/A AND2X1_LOC_41/A OR2X1_LOC_161/A OR2X1_LOC_78/B OR2X1_LOC_278/Y OR2X1_LOC_342/B OR2X1_LOC_485/A AND2X1_LOC_94/Y OR2X1_LOC_91/A AND2X1_LOC_612/B OR2X1_LOC_56/A OR2X1_LOC_136/Y OR2X1_LOC_459/A OR2X1_LOC_272/Y OR2X1_LOC_827/Y OR2X1_LOC_419/Y OR2X1_LOC_43/Y OR2X1_LOC_297/A OR2X1_LOC_534/Y OR2X1_LOC_490/Y OR2X1_LOC_789/B OR2X1_LOC_160/B OR2X1_LOC_756/B OR2X1_LOC_256/Y AND2X1_LOC_7/B OR2X1_LOC_20/A OR2X1_LOC_422/Y OR2X1_LOC_628/Y OR2X1_LOC_93/Y OR2X1_LOC_779/B OR2X1_LOC_520/A OR2X1_LOC_706/B AND2X1_LOC_48/Y 
+ OR2X1_LOC_405/Y OR2X1_LOC_399/A OR2X1_LOC_625/Y OR2X1_LOC_481/A OR2X1_LOC_585/Y OR2X1_LOC_416/A OR2X1_LOC_638/B OR2X1_LOC_459/B OR2X1_LOC_325/B OR2X1_LOC_168/B OR2X1_LOC_147/A OR2X1_LOC_512/A OR2X1_LOC_708/B OR2X1_LOC_502/Y OR2X1_LOC_156/A OR2X1_LOC_780/B OR2X1_LOC_828/B OR2X1_LOC_831/B OR2X1_LOC_435/A OR2X1_LOC_369/Y OR2X1_LOC_122/A OR2X1_LOC_299/Y OR2X1_LOC_607/A OR2X1_LOC_300/Y OR2X1_LOC_464/A OR2X1_LOC_65/B OR2X1_LOC_778/B AND2X1_LOC_72/B OR2X1_LOC_335/A AND2X1_LOC_57/Y OR2X1_LOC_68/Y OR2X1_LOC_672/Y OR2X1_LOC_622/B OR2X1_LOC_813/A OR2X1_LOC_690/A OR2X1_LOC_256/A OR2X1_LOC_278/A OR2X1_LOC_246/A OR2X1_LOC_86/A OR2X1_LOC_437/A AND2X1_LOC_65/A OR2X1_LOC_69/A OR2X1_LOC_71/Y OR2X1_LOC_57/Y OR2X1_LOC_371/Y OR2X1_LOC_310/Y OR2X1_LOC_706/A OR2X1_LOC_709/A OR2X1_LOC_378/A AND2X1_LOC_548/Y OR2X1_LOC_22/Y 
+ OR2X1_LOC_36/Y OR2X1_LOC_26/Y OR2X1_LOC_355/B OR2X1_LOC_448/B OR2X1_LOC_596/Y AND2X1_LOC_95/Y AND2X1_LOC_12/Y AND2X1_LOC_59/Y OR2X1_LOC_707/B OR2X1_LOC_753/Y OR2X1_LOC_12/Y OR2X1_LOC_59/Y OR2X1_LOC_18/Y OR2X1_LOC_31/Y OR2X1_LOC_44/Y OR2X1_LOC_47/Y AND2X1_LOC_70/Y AND2X1_LOC_40/Y AND2X1_LOC_3/Y AND2X1_LOC_64/Y AND2X1_LOC_22/Y OR2X1_LOC_66/A OR2X1_LOC_307/B OR2X1_LOC_197/A OR2X1_LOC_460/A OR2X1_LOC_582/Y OR2X1_LOC_451/A OR2X1_LOC_329/B OR2X1_LOC_66/Y OR2X1_LOC_121/A OR2X1_LOC_185/Y OR2X1_LOC_405/A OR2X1_LOC_67/A OR2X1_LOC_666/A OR2X1_LOC_816/A OR2X1_LOC_410/Y AND2X1_LOC_687/Y OR2X1_LOC_368/A OR2X1_LOC_87/Y OR2X1_LOC_373/Y OR2X1_LOC_517/A OR2X1_LOC_687/Y OR2X1_LOC_270/Y OR2X1_LOC_88/A OR2X1_LOC_411/A OR2X1_LOC_264/Y OR2X1_LOC_544/B OR2X1_LOC_682/Y OR2X1_LOC_683/Y OR2X1_LOC_686/B OR2X1_LOC_685/A 
+ OR2X1_LOC_88/Y AND2X1_LOC_374/Y OR2X1_LOC_599/Y OR2X1_LOC_644/A AND2X1_LOC_88/Y OR2X1_LOC_374/Y 

* NETLIST 
XAND2X1_LOC_587 AND2X1_LOC_587/a_36_24# AND2X1_LOC_588/B AND2X1_LOC_587/a_8_24# VSS VDD D_INPUT_7 AND2X1_LOC_51/A AND2X1_LOC

XAND2X1_LOC_50 AND2X1_LOC_50/a_36_24# AND2X1_LOC_50/Y AND2X1_LOC_50/a_8_24# VSS VDD D_INPUT_6 D_INPUT_7 AND2X1_LOC

XAND2X1_LOC_25 AND2X1_LOC_25/a_36_24# AND2X1_LOC_25/Y AND2X1_LOC_25/a_8_24# VSS VDD INPUT_6 D_INPUT_7 AND2X1_LOC

XOR2X1_LOC_1 OR2X1_LOC_1/a_8_216# OR2X1_LOC_1/a_36_216# OR2X1_LOC_3/B VSS VDD D_INPUT_7 INPUT_6 OR2X1_LOC

XOR2X1_LOC_17 OR2X1_LOC_17/a_8_216# OR2X1_LOC_17/a_36_216# OR2X1_LOC_17/Y VSS VDD D_INPUT_7 D_INPUT_6 OR2X1_LOC

XAND2X1_LOC_429 AND2X1_LOC_429/a_36_24# AND2X1_LOC_430/B AND2X1_LOC_429/a_8_24# VSS VDD D_INPUT_7 AND2X1_LOC_11/Y AND2X1_LOC

XAND2X1_LOC_1 AND2X1_LOC_1/a_36_24# AND2X1_LOC_1/Y AND2X1_LOC_1/a_8_24# VSS VDD D_INPUT_6 INPUT_7 AND2X1_LOC

XOR2X1_LOC_762 OR2X1_LOC_762/a_8_216# OR2X1_LOC_762/a_36_216# OR2X1_LOC_762/Y VSS VDD OR2X1_LOC_11/Y D_INPUT_6 OR2X1_LOC

XOR2X1_LOC_581 OR2X1_LOC_581/a_8_216# OR2X1_LOC_581/a_36_216# OR2X1_LOC_581/Y VSS VDD OR2X1_LOC_2/Y D_INPUT_6 OR2X1_LOC

XOR2X1_LOC_25 OR2X1_LOC_25/a_8_216# OR2X1_LOC_25/a_36_216# OR2X1_LOC_25/Y VSS VDD INPUT_7 D_INPUT_6 OR2X1_LOC

XAND2X1_LOC_408 AND2X1_LOC_408/a_36_24# AND2X1_LOC_409/B AND2X1_LOC_408/a_8_24# VSS VDD D_INPUT_6 AND2X1_LOC_21/Y AND2X1_LOC

XAND2X1_LOC_53 AND2X1_LOC_53/a_36_24# AND2X1_LOC_53/Y AND2X1_LOC_53/a_8_24# VSS VDD D_INPUT_5 AND2X1_LOC_50/Y AND2X1_LOC

XAND2X1_LOC_21 AND2X1_LOC_21/a_36_24# AND2X1_LOC_21/Y AND2X1_LOC_21/a_8_24# VSS VDD INPUT_4 D_INPUT_5 AND2X1_LOC

XAND2X1_LOC_2 AND2X1_LOC_2/a_36_24# AND2X1_LOC_2/Y AND2X1_LOC_2/a_8_24# VSS VDD D_INPUT_4 D_INPUT_5 AND2X1_LOC

XOR2X1_LOC_30 OR2X1_LOC_30/a_8_216# OR2X1_LOC_30/a_36_216# OR2X1_LOC_51/B VSS VDD D_INPUT_5 D_INPUT_4 OR2X1_LOC

XOR2X1_LOC_11 OR2X1_LOC_11/a_8_216# OR2X1_LOC_11/a_36_216# OR2X1_LOC_11/Y VSS VDD D_INPUT_5 INPUT_4 OR2X1_LOC

XOR2X1_LOC_752 OR2X1_LOC_752/a_8_216# OR2X1_LOC_752/a_36_216# OR2X1_LOC_753/A VSS VDD OR2X1_LOC_70/A D_INPUT_5 OR2X1_LOC

XAND2X1_LOC_425 AND2X1_LOC_425/a_36_24# AND2X1_LOC_425/Y AND2X1_LOC_425/a_8_24# VSS VDD D_INPUT_5 AND2X1_LOC_17/Y AND2X1_LOC

XAND2X1_LOC_386 AND2X1_LOC_386/a_36_24# AND2X1_LOC_387/B AND2X1_LOC_386/a_8_24# VSS VDD D_INPUT_4 AND2X1_LOC_17/Y AND2X1_LOC

XAND2X1_LOC_11 AND2X1_LOC_11/a_36_24# AND2X1_LOC_11/Y AND2X1_LOC_11/a_8_24# VSS VDD D_INPUT_4 INPUT_5 AND2X1_LOC

XAND2X1_LOC_328 AND2X1_LOC_328/a_36_24# OR2X1_LOC_596/A AND2X1_LOC_328/a_8_24# VSS VDD D_INPUT_4 AND2X1_LOC_50/Y AND2X1_LOC

XOR2X1_LOC_21 OR2X1_LOC_21/a_8_216# OR2X1_LOC_21/a_36_216# OR2X1_LOC_22/A VSS VDD INPUT_5 D_INPUT_4 OR2X1_LOC

XOR2X1_LOC_529 OR2X1_LOC_529/a_8_216# OR2X1_LOC_529/a_36_216# OR2X1_LOC_529/Y VSS VDD OR2X1_LOC_26/Y D_INPUT_3 OR2X1_LOC

XAND2X1_LOC_14 AND2X1_LOC_14/a_36_24# OR2X1_LOC_377/A AND2X1_LOC_14/a_8_24# VSS VDD D_INPUT_2 D_INPUT_3 AND2X1_LOC

XOR2X1_LOC_414 OR2X1_LOC_414/a_8_216# OR2X1_LOC_414/a_36_216# OR2X1_LOC_414/Y VSS VDD OR2X1_LOC_6/B D_INPUT_3 OR2X1_LOC

XOR2X1_LOC_5 OR2X1_LOC_5/a_8_216# OR2X1_LOC_5/a_36_216# OR2X1_LOC_6/A VSS VDD D_INPUT_3 INPUT_2 OR2X1_LOC

XAND2X1_LOC_8 AND2X1_LOC_8/a_36_24# AND2X1_LOC_8/Y AND2X1_LOC_8/a_8_24# VSS VDD INPUT_2 D_INPUT_3 AND2X1_LOC

XOR2X1_LOC_381 OR2X1_LOC_381/a_8_216# OR2X1_LOC_381/a_36_216# OR2X1_LOC_382/A VSS VDD OR2X1_LOC_12/Y D_INPUT_3 OR2X1_LOC

XOR2X1_LOC_37 OR2X1_LOC_37/a_8_216# OR2X1_LOC_37/a_36_216# OR2X1_LOC_85/A VSS VDD D_INPUT_3 D_INPUT_2 OR2X1_LOC

XAND2X1_LOC_618 AND2X1_LOC_618/a_36_24# AND2X1_LOC_619/B AND2X1_LOC_618/a_8_24# VSS VDD D_INPUT_3 OR2X1_LOC_80/A AND2X1_LOC

XOR2X1_LOC_671 OR2X1_LOC_671/a_8_216# OR2X1_LOC_671/a_36_216# OR2X1_LOC_671/Y VSS VDD OR2X1_LOC_6/B D_INPUT_2 OR2X1_LOC

XAND2X1_LOC_5 AND2X1_LOC_5/a_36_24# OR2X1_LOC_68/B AND2X1_LOC_5/a_8_24# VSS VDD D_INPUT_2 INPUT_3 AND2X1_LOC

XOR2X1_LOC_8 OR2X1_LOC_8/a_8_216# OR2X1_LOC_8/a_36_216# OR2X1_LOC_8/Y VSS VDD INPUT_3 D_INPUT_2 OR2X1_LOC

XAND2X1_LOC_372 AND2X1_LOC_372/a_36_24# OR2X1_LOC_458/B AND2X1_LOC_372/a_8_24# VSS VDD D_INPUT_1 OR2X1_LOC_778/B AND2X1_LOC

XOR2X1_LOC_119 OR2X1_LOC_119/a_8_216# OR2X1_LOC_119/a_36_216# OR2X1_LOC_426/B VSS VDD OR2X1_LOC_46/A D_INPUT_1 OR2X1_LOC

XAND2X1_LOC_153 AND2X1_LOC_153/a_36_24# OR2X1_LOC_155/A AND2X1_LOC_153/a_8_24# VSS VDD D_INPUT_1 AND2X1_LOC_42/B AND2X1_LOC

XAND2X1_LOC_143 AND2X1_LOC_143/a_36_24# OR2X1_LOC_502/A AND2X1_LOC_143/a_8_24# VSS VDD D_INPUT_1 AND2X1_LOC_8/Y AND2X1_LOC

XOR2X1_LOC_293 OR2X1_LOC_293/a_8_216# OR2X1_LOC_293/a_36_216# OR2X1_LOC_585/A VSS VDD OR2X1_LOC_6/A D_INPUT_1 OR2X1_LOC

XAND2X1_LOC_46 AND2X1_LOC_46/a_36_24# AND2X1_LOC_48/A AND2X1_LOC_46/a_8_24# VSS VDD D_INPUT_1 OR2X1_LOC_377/A AND2X1_LOC

XOR2X1_LOC_92 OR2X1_LOC_92/a_8_216# OR2X1_LOC_92/a_36_216# OR2X1_LOC_92/Y VSS VDD OR2X1_LOC_8/Y D_INPUT_1 OR2X1_LOC

XAND2X1_LOC_4 AND2X1_LOC_4/a_36_24# OR2X1_LOC_19/B AND2X1_LOC_4/a_8_24# VSS VDD INPUT_0 D_INPUT_1 AND2X1_LOC

XOR2X1_LOC_42 OR2X1_LOC_42/a_8_216# OR2X1_LOC_42/a_36_216# OR2X1_LOC_43/A VSS VDD OR2X1_LOC_85/A D_INPUT_1 OR2X1_LOC

XOR2X1_LOC_54 OR2X1_LOC_54/a_8_216# OR2X1_LOC_54/a_36_216# OR2X1_LOC_54/Y VSS VDD D_INPUT_1 D_INPUT_0 OR2X1_LOC

XAND2X1_LOC_9 AND2X1_LOC_9/a_36_24# OR2X1_LOC_62/B AND2X1_LOC_9/a_8_24# VSS VDD D_INPUT_0 D_INPUT_1 AND2X1_LOC

XAND2X1_LOC_817 AND2X1_LOC_817/a_36_24# OR2X1_LOC_847/B AND2X1_LOC_817/a_8_24# VSS VDD D_INPUT_1 AND2X1_LOC_817/B AND2X1_LOC

XOR2X1_LOC_28 OR2X1_LOC_28/a_8_216# OR2X1_LOC_28/a_36_216# OR2X1_LOC_49/A VSS VDD D_INPUT_1 INPUT_0 OR2X1_LOC

XAND2X1_LOC_225 AND2X1_LOC_225/a_36_24# OR2X1_LOC_814/A AND2X1_LOC_225/a_8_24# VSS VDD D_INPUT_1 OR2X1_LOC_68/B AND2X1_LOC

XAND2X1_LOC_749 AND2X1_LOC_749/a_36_24# OR2X1_LOC_750/A AND2X1_LOC_749/a_8_24# VSS VDD D_INPUT_0 AND2X1_LOC_8/Y AND2X1_LOC

XAND2X1_LOC_514 AND2X1_LOC_514/a_36_24# AND2X1_LOC_514/Y AND2X1_LOC_514/a_8_24# VSS VDD D_INPUT_0 OR2X1_LOC_136/Y AND2X1_LOC

XAND2X1_LOC_110 AND2X1_LOC_110/a_36_24# AND2X1_LOC_110/Y AND2X1_LOC_110/a_8_24# VSS VDD D_INPUT_0 OR2X1_LOC_377/A AND2X1_LOC

XAND2X1_LOC_690 AND2X1_LOC_690/a_36_24# OR2X1_LOC_691/A AND2X1_LOC_690/a_8_24# VSS VDD D_INPUT_0 OR2X1_LOC_634/A AND2X1_LOC

XOR2X1_LOC_413 OR2X1_LOC_413/a_8_216# OR2X1_LOC_413/a_36_216# OR2X1_LOC_413/Y VSS VDD OR2X1_LOC_690/A D_INPUT_0 OR2X1_LOC

XOR2X1_LOC_233 OR2X1_LOC_233/a_8_216# OR2X1_LOC_233/a_36_216# OR2X1_LOC_291/A VSS VDD OR2X1_LOC_46/A D_INPUT_0 OR2X1_LOC

XAND2X1_LOC_28 AND2X1_LOC_28/a_36_24# OR2X1_LOC_80/A AND2X1_LOC_28/a_8_24# VSS VDD D_INPUT_0 INPUT_1 AND2X1_LOC

XOR2X1_LOC_4 OR2X1_LOC_4/a_8_216# OR2X1_LOC_4/a_36_216# OR2X1_LOC_6/B VSS VDD INPUT_1 D_INPUT_0 OR2X1_LOC

XOR2X1_LOC_86 OR2X1_LOC_86/a_8_216# OR2X1_LOC_86/a_36_216# OR2X1_LOC_86/Y VSS VDD OR2X1_LOC_86/A D_INPUT_0 OR2X1_LOC

XAND2X1_LOC_275 AND2X1_LOC_275/a_36_24# OR2X1_LOC_276/A AND2X1_LOC_275/a_8_24# VSS VDD D_INPUT_0 OR2X1_LOC_274/Y AND2X1_LOC

XOR2X1_LOC_512 OR2X1_LOC_512/a_8_216# OR2X1_LOC_512/a_36_216# OR2X1_LOC_512/Y VSS VDD OR2X1_LOC_512/A D_INPUT_0 OR2X1_LOC

XAND2X1_LOC_761 AND2X1_LOC_761/a_36_24# OR2X1_LOC_801/B AND2X1_LOC_761/a_8_24# VSS VDD D_INPUT_0 OR2X1_LOC_644/A AND2X1_LOC

XAND2X1_LOC_17 AND2X1_LOC_17/a_36_24# AND2X1_LOC_17/Y AND2X1_LOC_17/a_8_24# VSS VDD INPUT_6 INPUT_7 AND2X1_LOC

XOR2X1_LOC_50 OR2X1_LOC_50/a_8_216# OR2X1_LOC_50/a_36_216# OR2X1_LOC_70/A VSS VDD INPUT_7 INPUT_6 OR2X1_LOC

XOR2X1_LOC_429 OR2X1_LOC_429/a_8_216# OR2X1_LOC_429/a_36_216# OR2X1_LOC_429/Y VSS VDD OR2X1_LOC_11/Y INPUT_7 OR2X1_LOC

XOR2X1_LOC_587 OR2X1_LOC_587/a_8_216# OR2X1_LOC_587/a_36_216# OR2X1_LOC_588/A VSS VDD OR2X1_LOC_51/B INPUT_7 OR2X1_LOC

XOR2X1_LOC_408 OR2X1_LOC_408/a_8_216# OR2X1_LOC_408/a_36_216# OR2X1_LOC_408/Y VSS VDD OR2X1_LOC_22/A INPUT_6 OR2X1_LOC

XAND2X1_LOC_762 AND2X1_LOC_762/a_36_24# AND2X1_LOC_763/B AND2X1_LOC_762/a_8_24# VSS VDD INPUT_6 AND2X1_LOC_11/Y AND2X1_LOC

XAND2X1_LOC_581 AND2X1_LOC_581/a_36_24# AND2X1_LOC_582/B AND2X1_LOC_581/a_8_24# VSS VDD INPUT_6 AND2X1_LOC_2/Y AND2X1_LOC

XAND2X1_LOC_752 AND2X1_LOC_752/a_36_24# AND2X1_LOC_753/B AND2X1_LOC_752/a_8_24# VSS VDD INPUT_5 AND2X1_LOC_50/Y AND2X1_LOC

XAND2X1_LOC_30 AND2X1_LOC_30/a_36_24# AND2X1_LOC_51/A AND2X1_LOC_30/a_8_24# VSS VDD INPUT_4 INPUT_5 AND2X1_LOC

XOR2X1_LOC_425 OR2X1_LOC_425/a_8_216# OR2X1_LOC_425/a_36_216# OR2X1_LOC_426/A VSS VDD OR2X1_LOC_17/Y INPUT_5 OR2X1_LOC

XOR2X1_LOC_2 OR2X1_LOC_2/a_8_216# OR2X1_LOC_2/a_36_216# OR2X1_LOC_2/Y VSS VDD INPUT_5 INPUT_4 OR2X1_LOC

XOR2X1_LOC_53 OR2X1_LOC_53/a_8_216# OR2X1_LOC_53/a_36_216# OR2X1_LOC_53/Y VSS VDD OR2X1_LOC_70/A INPUT_5 OR2X1_LOC

XOR2X1_LOC_328 OR2X1_LOC_328/a_8_216# OR2X1_LOC_328/a_36_216# OR2X1_LOC_421/A VSS VDD OR2X1_LOC_70/A INPUT_4 OR2X1_LOC

XOR2X1_LOC_386 OR2X1_LOC_386/a_8_216# OR2X1_LOC_386/a_36_216# OR2X1_LOC_387/A VSS VDD OR2X1_LOC_17/Y INPUT_4 OR2X1_LOC

XAND2X1_LOC_381 AND2X1_LOC_381/a_36_24# AND2X1_LOC_817/B AND2X1_LOC_381/a_8_24# VSS VDD INPUT_3 AND2X1_LOC_12/Y AND2X1_LOC

XAND2X1_LOC_529 AND2X1_LOC_529/a_36_24# OR2X1_LOC_548/B AND2X1_LOC_529/a_8_24# VSS VDD INPUT_3 OR2X1_LOC_66/A AND2X1_LOC

XAND2X1_LOC_37 AND2X1_LOC_37/a_36_24# AND2X1_LOC_42/B AND2X1_LOC_37/a_8_24# VSS VDD INPUT_2 INPUT_3 AND2X1_LOC

XOR2X1_LOC_618 OR2X1_LOC_618/a_8_216# OR2X1_LOC_618/a_36_216# OR2X1_LOC_618/Y VSS VDD OR2X1_LOC_49/A INPUT_3 OR2X1_LOC

XOR2X1_LOC_14 OR2X1_LOC_14/a_8_216# OR2X1_LOC_14/a_36_216# OR2X1_LOC_46/A VSS VDD INPUT_3 INPUT_2 OR2X1_LOC

XAND2X1_LOC_414 AND2X1_LOC_414/a_36_24# OR2X1_LOC_415/A AND2X1_LOC_414/a_8_24# VSS VDD INPUT_3 OR2X1_LOC_19/B AND2X1_LOC

XAND2X1_LOC_671 AND2X1_LOC_671/a_36_24# AND2X1_LOC_672/B AND2X1_LOC_671/a_8_24# VSS VDD INPUT_2 OR2X1_LOC_19/B AND2X1_LOC

XOR2X1_LOC_143 OR2X1_LOC_143/a_8_216# OR2X1_LOC_143/a_36_216# OR2X1_LOC_696/A VSS VDD OR2X1_LOC_8/Y INPUT_1 OR2X1_LOC

XAND2X1_LOC_92 AND2X1_LOC_92/a_36_24# AND2X1_LOC_92/Y AND2X1_LOC_92/a_8_24# VSS VDD INPUT_1 AND2X1_LOC_8/Y AND2X1_LOC

XAND2X1_LOC_42 AND2X1_LOC_42/a_36_24# AND2X1_LOC_43/B AND2X1_LOC_42/a_8_24# VSS VDD INPUT_1 AND2X1_LOC_42/B AND2X1_LOC

XAND2X1_LOC_54 AND2X1_LOC_54/a_36_24# OR2X1_LOC_62/A AND2X1_LOC_54/a_8_24# VSS VDD INPUT_0 INPUT_1 AND2X1_LOC

XOR2X1_LOC_817 OR2X1_LOC_817/a_8_216# OR2X1_LOC_817/a_36_216# OR2X1_LOC_817/Y VSS VDD OR2X1_LOC_382/A INPUT_1 OR2X1_LOC

XAND2X1_LOC_119 AND2X1_LOC_119/a_36_24# OR2X1_LOC_121/B AND2X1_LOC_119/a_8_24# VSS VDD INPUT_1 OR2X1_LOC_377/A AND2X1_LOC

XOR2X1_LOC_225 OR2X1_LOC_225/a_8_216# OR2X1_LOC_225/a_36_216# OR2X1_LOC_417/A VSS VDD OR2X1_LOC_6/A INPUT_1 OR2X1_LOC

XAND2X1_LOC_293 AND2X1_LOC_293/a_36_24# OR2X1_LOC_598/A AND2X1_LOC_293/a_8_24# VSS VDD INPUT_1 OR2X1_LOC_68/B AND2X1_LOC

XOR2X1_LOC_9 OR2X1_LOC_9/a_8_216# OR2X1_LOC_9/a_36_216# OR2X1_LOC_9/Y VSS VDD INPUT_1 INPUT_0 OR2X1_LOC

XOR2X1_LOC_46 OR2X1_LOC_46/a_8_216# OR2X1_LOC_46/a_36_216# OR2X1_LOC_48/B VSS VDD OR2X1_LOC_46/A INPUT_1 OR2X1_LOC

XOR2X1_LOC_372 OR2X1_LOC_372/a_8_216# OR2X1_LOC_372/a_36_216# OR2X1_LOC_372/Y VSS VDD OR2X1_LOC_371/Y INPUT_1 OR2X1_LOC

XOR2X1_LOC_153 OR2X1_LOC_153/a_8_216# OR2X1_LOC_153/a_36_216# OR2X1_LOC_743/A VSS VDD OR2X1_LOC_85/A INPUT_1 OR2X1_LOC

XOR2X1_LOC_110 OR2X1_LOC_110/a_8_216# OR2X1_LOC_110/a_36_216# OR2X1_LOC_323/A VSS VDD OR2X1_LOC_46/A INPUT_0 OR2X1_LOC

XOR2X1_LOC_690 OR2X1_LOC_690/a_8_216# OR2X1_LOC_690/a_36_216# OR2X1_LOC_690/Y VSS VDD OR2X1_LOC_690/A INPUT_0 OR2X1_LOC

XAND2X1_LOC_512 AND2X1_LOC_512/a_36_24# AND2X1_LOC_512/Y AND2X1_LOC_512/a_8_24# VSS VDD INPUT_0 OR2X1_LOC_306/Y AND2X1_LOC

XAND2X1_LOC_86 AND2X1_LOC_86/a_36_24# AND2X1_LOC_86/Y AND2X1_LOC_86/a_8_24# VSS VDD INPUT_0 AND2X1_LOC_86/B AND2X1_LOC

XOR2X1_LOC_275 OR2X1_LOC_275/a_8_216# OR2X1_LOC_275/a_36_216# OR2X1_LOC_275/Y VSS VDD OR2X1_LOC_275/A INPUT_0 OR2X1_LOC

XOR2X1_LOC_761 OR2X1_LOC_761/a_8_216# OR2X1_LOC_761/a_36_216# OR2X1_LOC_761/Y VSS VDD OR2X1_LOC_599/Y INPUT_0 OR2X1_LOC

XAND2X1_LOC_413 AND2X1_LOC_413/a_36_24# OR2X1_LOC_461/A AND2X1_LOC_413/a_8_24# VSS VDD INPUT_0 OR2X1_LOC_634/A AND2X1_LOC

XAND2X1_LOC_233 AND2X1_LOC_233/a_36_24# AND2X1_LOC_824/B AND2X1_LOC_233/a_8_24# VSS VDD INPUT_0 OR2X1_LOC_377/A AND2X1_LOC

XOR2X1_LOC_749 OR2X1_LOC_749/a_8_216# OR2X1_LOC_749/a_36_216# OR2X1_LOC_749/Y VSS VDD OR2X1_LOC_8/Y INPUT_0 OR2X1_LOC

XOR2X1_LOC_514 OR2X1_LOC_514/a_8_216# OR2X1_LOC_514/a_36_216# OR2X1_LOC_515/A VSS VDD OR2X1_LOC_138/A INPUT_0 OR2X1_LOC

XOR2X1_LOC_515 OR2X1_LOC_515/a_8_216# OR2X1_LOC_515/a_36_216# OR2X1_LOC_515/Y VSS VDD OR2X1_LOC_515/A OR2X1_LOC_446/B OR2X1_LOC

XAND2X1_LOC_750 AND2X1_LOC_750/a_36_24# OR2X1_LOC_751/A AND2X1_LOC_750/a_8_24# VSS VDD OR2X1_LOC_604/A OR2X1_LOC_749/Y AND2X1_LOC

XAND2X1_LOC_291 AND2X1_LOC_291/a_36_24# OR2X1_LOC_334/A AND2X1_LOC_291/a_8_24# VSS VDD AND2X1_LOC_36/Y AND2X1_LOC_824/B AND2X1_LOC

XAND2X1_LOC_824 AND2X1_LOC_824/a_36_24# OR2X1_LOC_836/A AND2X1_LOC_824/a_8_24# VSS VDD OR2X1_LOC_66/A AND2X1_LOC_824/B AND2X1_LOC

XAND2X1_LOC_234 AND2X1_LOC_234/a_36_24# OR2X1_LOC_240/A AND2X1_LOC_234/a_8_24# VSS VDD AND2X1_LOC_47/Y AND2X1_LOC_824/B AND2X1_LOC

XOR2X1_LOC_461 OR2X1_LOC_461/a_8_216# OR2X1_LOC_461/a_36_216# OR2X1_LOC_461/Y VSS VDD OR2X1_LOC_461/A OR2X1_LOC_461/B OR2X1_LOC

XAND2X1_LOC_801 AND2X1_LOC_801/a_36_24# AND2X1_LOC_809/A AND2X1_LOC_801/a_8_24# VSS VDD OR2X1_LOC_761/Y AND2X1_LOC_801/B AND2X1_LOC

XAND2X1_LOC_276 AND2X1_LOC_276/a_36_24# AND2X1_LOC_276/Y AND2X1_LOC_276/a_8_24# VSS VDD OR2X1_LOC_271/Y OR2X1_LOC_275/Y AND2X1_LOC

XOR2X1_LOC_100 OR2X1_LOC_100/a_8_216# OR2X1_LOC_100/a_36_216# OR2X1_LOC_100/Y VSS VDD AND2X1_LOC_88/Y AND2X1_LOC_86/Y OR2X1_LOC

XAND2X1_LOC_513 AND2X1_LOC_513/a_36_24# OR2X1_LOC_516/B AND2X1_LOC_513/a_8_24# VSS VDD OR2X1_LOC_511/Y AND2X1_LOC_512/Y AND2X1_LOC

XAND2X1_LOC_691 AND2X1_LOC_691/a_36_24# AND2X1_LOC_729/B AND2X1_LOC_691/a_8_24# VSS VDD OR2X1_LOC_689/Y OR2X1_LOC_690/Y AND2X1_LOC

XOR2X1_LOC_527 OR2X1_LOC_527/a_8_216# OR2X1_LOC_527/a_36_216# OR2X1_LOC_527/Y VSS VDD OR2X1_LOC_323/A OR2X1_LOC_64/Y OR2X1_LOC

XOR2X1_LOC_111 OR2X1_LOC_111/a_8_216# OR2X1_LOC_111/a_36_216# OR2X1_LOC_111/Y VSS VDD OR2X1_LOC_323/A OR2X1_LOC_31/Y OR2X1_LOC

XOR2X1_LOC_323 OR2X1_LOC_323/a_8_216# OR2X1_LOC_323/a_36_216# OR2X1_LOC_323/Y VSS VDD OR2X1_LOC_323/A OR2X1_LOC_95/Y OR2X1_LOC

XOR2X1_LOC_681 OR2X1_LOC_681/a_8_216# OR2X1_LOC_681/a_36_216# OR2X1_LOC_681/Y VSS VDD OR2X1_LOC_743/A OR2X1_LOC_31/Y OR2X1_LOC

XAND2X1_LOC_155 AND2X1_LOC_155/a_36_24# AND2X1_LOC_155/Y AND2X1_LOC_155/a_8_24# VSS VDD OR2X1_LOC_52/B OR2X1_LOC_743/A AND2X1_LOC

XOR2X1_LOC_273 OR2X1_LOC_273/a_8_216# OR2X1_LOC_273/a_36_216# OR2X1_LOC_273/Y VSS VDD OR2X1_LOC_743/A OR2X1_LOC_36/Y OR2X1_LOC

XOR2X1_LOC_433 OR2X1_LOC_433/a_8_216# OR2X1_LOC_433/a_36_216# OR2X1_LOC_433/Y VSS VDD OR2X1_LOC_743/A OR2X1_LOC_70/Y OR2X1_LOC

XOR2X1_LOC_743 OR2X1_LOC_743/a_8_216# OR2X1_LOC_743/a_36_216# OR2X1_LOC_743/Y VSS VDD OR2X1_LOC_743/A OR2X1_LOC_3/Y OR2X1_LOC

XAND2X1_LOC_407 AND2X1_LOC_407/a_36_24# OR2X1_LOC_409/B AND2X1_LOC_407/a_8_24# VSS VDD OR2X1_LOC_56/A OR2X1_LOC_743/A AND2X1_LOC

XAND2X1_LOC_458 AND2X1_LOC_458/a_36_24# AND2X1_LOC_458/Y AND2X1_LOC_458/a_8_24# VSS VDD OR2X1_LOC_372/Y AND2X1_LOC_374/Y AND2X1_LOC

XOR2X1_LOC_519 OR2X1_LOC_519/a_8_216# OR2X1_LOC_519/a_36_216# OR2X1_LOC_519/Y VSS VDD OR2X1_LOC_158/A OR2X1_LOC_48/B OR2X1_LOC

XOR2X1_LOC_692 OR2X1_LOC_692/a_8_216# OR2X1_LOC_692/a_36_216# OR2X1_LOC_692/Y VSS VDD OR2X1_LOC_48/B OR2X1_LOC_18/Y OR2X1_LOC

XAND2X1_LOC_598 AND2X1_LOC_598/a_36_24# OR2X1_LOC_599/A AND2X1_LOC_598/a_8_24# VSS VDD OR2X1_LOC_48/B OR2X1_LOC_585/A AND2X1_LOC

XOR2X1_LOC_763 OR2X1_LOC_763/a_8_216# OR2X1_LOC_763/a_36_216# OR2X1_LOC_763/Y VSS VDD OR2X1_LOC_762/Y OR2X1_LOC_48/B OR2X1_LOC

XOR2X1_LOC_48 OR2X1_LOC_48/a_8_216# OR2X1_LOC_48/a_36_216# OR2X1_LOC_48/Y VSS VDD OR2X1_LOC_47/Y OR2X1_LOC_48/B OR2X1_LOC

XAND2X1_LOC_405 AND2X1_LOC_405/a_36_24# OR2X1_LOC_406/A AND2X1_LOC_405/a_8_24# VSS VDD OR2X1_LOC_48/B OR2X1_LOC_329/B AND2X1_LOC

XOR2X1_LOC_511 OR2X1_LOC_511/a_8_216# OR2X1_LOC_511/a_36_216# OR2X1_LOC_511/Y VSS VDD OR2X1_LOC_48/B OR2X1_LOC_31/Y OR2X1_LOC

XOR2X1_LOC_159 OR2X1_LOC_159/a_8_216# OR2X1_LOC_159/a_36_216# OR2X1_LOC_604/A VSS VDD OR2X1_LOC_9/Y OR2X1_LOC_6/A OR2X1_LOC

XAND2X1_LOC_62 AND2X1_LOC_62/a_36_24# OR2X1_LOC_235/B AND2X1_LOC_62/a_8_24# VSS VDD OR2X1_LOC_9/Y OR2X1_LOC_54/Y AND2X1_LOC

XOR2X1_LOC_246 OR2X1_LOC_246/a_8_216# OR2X1_LOC_246/a_36_216# OR2X1_LOC_246/Y VSS VDD OR2X1_LOC_246/A OR2X1_LOC_9/Y OR2X1_LOC

XOR2X1_LOC_73 OR2X1_LOC_73/a_8_216# OR2X1_LOC_73/a_36_216# OR2X1_LOC_74/A VSS VDD OR2X1_LOC_85/A OR2X1_LOC_9/Y OR2X1_LOC

XOR2X1_LOC_10 OR2X1_LOC_10/a_8_216# OR2X1_LOC_10/a_36_216# OR2X1_LOC_13/B VSS VDD OR2X1_LOC_9/Y OR2X1_LOC_8/Y OR2X1_LOC

XOR2X1_LOC_15 OR2X1_LOC_15/a_8_216# OR2X1_LOC_15/a_36_216# OR2X1_LOC_16/A VSS VDD OR2X1_LOC_46/A OR2X1_LOC_9/Y OR2X1_LOC

XAND2X1_LOC_278 AND2X1_LOC_278/a_36_24# OR2X1_LOC_287/B AND2X1_LOC_278/a_8_24# VSS VDD OR2X1_LOC_9/Y OR2X1_LOC_633/A AND2X1_LOC

XAND2X1_LOC_585 AND2X1_LOC_585/a_36_24# OR2X1_LOC_637/B AND2X1_LOC_585/a_8_24# VSS VDD AND2X1_LOC_22/Y OR2X1_LOC_598/A AND2X1_LOC

XOR2X1_LOC_688 OR2X1_LOC_688/a_8_216# OR2X1_LOC_688/a_36_216# OR2X1_LOC_688/Y VSS VDD OR2X1_LOC_598/A OR2X1_LOC_154/A OR2X1_LOC

XOR2X1_LOC_294 OR2X1_LOC_294/a_8_216# OR2X1_LOC_294/a_36_216# OR2X1_LOC_294/Y VSS VDD OR2X1_LOC_598/A AND2X1_LOC_41/A OR2X1_LOC

XOR2X1_LOC_415 OR2X1_LOC_415/a_8_216# OR2X1_LOC_415/a_36_216# OR2X1_LOC_415/Y VSS VDD OR2X1_LOC_415/A OR2X1_LOC_598/A OR2X1_LOC

XAND2X1_LOC_625 AND2X1_LOC_625/a_36_24# OR2X1_LOC_631/A AND2X1_LOC_625/a_8_24# VSS VDD OR2X1_LOC_66/Y OR2X1_LOC_598/A AND2X1_LOC

XOR2X1_LOC_598 OR2X1_LOC_598/a_8_216# OR2X1_LOC_598/a_36_216# OR2X1_LOC_598/Y VSS VDD OR2X1_LOC_598/A AND2X1_LOC_48/A OR2X1_LOC

XOR2X1_LOC_398 OR2X1_LOC_398/a_8_216# OR2X1_LOC_398/a_36_216# OR2X1_LOC_398/Y VSS VDD OR2X1_LOC_598/A OR2X1_LOC_78/B OR2X1_LOC

XOR2X1_LOC_309 OR2X1_LOC_309/a_8_216# OR2X1_LOC_309/a_36_216# OR2X1_LOC_309/Y VSS VDD OR2X1_LOC_417/A OR2X1_LOC_22/Y OR2X1_LOC

XOR2X1_LOC_283 OR2X1_LOC_283/a_8_216# OR2X1_LOC_283/a_36_216# OR2X1_LOC_283/Y VSS VDD OR2X1_LOC_417/A OR2X1_LOC_26/Y OR2X1_LOC

XOR2X1_LOC_488 OR2X1_LOC_488/a_8_216# OR2X1_LOC_488/a_36_216# OR2X1_LOC_488/Y VSS VDD OR2X1_LOC_417/A OR2X1_LOC_158/A OR2X1_LOC

XOR2X1_LOC_289 OR2X1_LOC_289/a_8_216# OR2X1_LOC_289/a_36_216# OR2X1_LOC_289/Y VSS VDD OR2X1_LOC_417/A OR2X1_LOC_51/Y OR2X1_LOC

XOR2X1_LOC_417 OR2X1_LOC_417/a_8_216# OR2X1_LOC_417/a_36_216# OR2X1_LOC_417/Y VSS VDD OR2X1_LOC_417/A OR2X1_LOC_47/Y OR2X1_LOC

XOR2X1_LOC_226 OR2X1_LOC_226/a_8_216# OR2X1_LOC_226/a_36_216# OR2X1_LOC_226/Y VSS VDD OR2X1_LOC_417/A OR2X1_LOC_18/Y OR2X1_LOC

XAND2X1_LOC_814 AND2X1_LOC_814/a_36_24# OR2X1_LOC_815/A AND2X1_LOC_814/a_8_24# VSS VDD OR2X1_LOC_600/A OR2X1_LOC_417/A AND2X1_LOC

XOR2X1_LOC_121 OR2X1_LOC_121/a_8_216# OR2X1_LOC_121/a_36_216# OR2X1_LOC_121/Y VSS VDD OR2X1_LOC_121/A OR2X1_LOC_121/B OR2X1_LOC

XAND2X1_LOC_300 AND2X1_LOC_300/a_36_24# OR2X1_LOC_831/A AND2X1_LOC_300/a_8_24# VSS VDD AND2X1_LOC_59/Y OR2X1_LOC_121/B AND2X1_LOC

XAND2X1_LOC_369 AND2X1_LOC_369/a_36_24# OR2X1_LOC_543/A AND2X1_LOC_369/a_8_24# VSS VDD AND2X1_LOC_22/Y OR2X1_LOC_121/B AND2X1_LOC

XOR2X1_LOC_606 OR2X1_LOC_606/a_8_216# OR2X1_LOC_606/a_36_216# OR2X1_LOC_606/Y VSS VDD OR2X1_LOC_121/B OR2X1_LOC_532/B OR2X1_LOC

XAND2X1_LOC_299 AND2X1_LOC_299/a_36_24# OR2X1_LOC_302/A AND2X1_LOC_299/a_8_24# VSS VDD AND2X1_LOC_12/Y OR2X1_LOC_121/B AND2X1_LOC

XAND2X1_LOC_426 AND2X1_LOC_426/a_36_24# OR2X1_LOC_450/B AND2X1_LOC_426/a_8_24# VSS VDD OR2X1_LOC_121/B AND2X1_LOC_425/Y AND2X1_LOC

XAND2X1_LOC_847 AND2X1_LOC_847/a_36_24# AND2X1_LOC_847/Y AND2X1_LOC_847/a_8_24# VSS VDD OR2X1_LOC_817/Y OR2X1_LOC_820/Y AND2X1_LOC

XAND2X1_LOC_90 AND2X1_LOC_90/a_36_24# AND2X1_LOC_91/B AND2X1_LOC_90/a_8_24# VSS VDD AND2X1_LOC_42/B OR2X1_LOC_62/A AND2X1_LOC

XOR2X1_LOC_611 OR2X1_LOC_611/a_8_216# OR2X1_LOC_611/a_36_216# OR2X1_LOC_611/Y VSS VDD OR2X1_LOC_62/A OR2X1_LOC_6/A OR2X1_LOC

XAND2X1_LOC_55 AND2X1_LOC_55/a_36_24# AND2X1_LOC_56/B AND2X1_LOC_55/a_8_24# VSS VDD OR2X1_LOC_68/B OR2X1_LOC_62/A AND2X1_LOC

XAND2X1_LOC_77 AND2X1_LOC_77/a_36_24# OR2X1_LOC_78/A AND2X1_LOC_77/a_8_24# VSS VDD OR2X1_LOC_377/A OR2X1_LOC_62/A AND2X1_LOC

XAND2X1_LOC_102 AND2X1_LOC_102/a_36_24# OR2X1_LOC_532/B AND2X1_LOC_102/a_8_24# VSS VDD AND2X1_LOC_8/Y OR2X1_LOC_62/A AND2X1_LOC

XOR2X1_LOC_819 OR2X1_LOC_819/a_8_216# OR2X1_LOC_819/a_36_216# OR2X1_LOC_820/A VSS VDD OR2X1_LOC_62/A OR2X1_LOC_47/Y OR2X1_LOC

XOR2X1_LOC_94 OR2X1_LOC_94/a_8_216# OR2X1_LOC_94/a_36_216# OR2X1_LOC_96/B VSS VDD OR2X1_LOC_62/A OR2X1_LOC_46/A OR2X1_LOC

XOR2X1_LOC_62 OR2X1_LOC_62/a_8_216# OR2X1_LOC_62/a_36_216# OR2X1_LOC_71/A VSS VDD OR2X1_LOC_62/A OR2X1_LOC_62/B OR2X1_LOC

XAND2X1_LOC_534 AND2X1_LOC_534/a_36_24# OR2X1_LOC_535/A AND2X1_LOC_534/a_8_24# VSS VDD AND2X1_LOC_43/B AND2X1_LOC_59/Y AND2X1_LOC

XAND2X1_LOC_43 AND2X1_LOC_43/a_36_24# OR2X1_LOC_195/A AND2X1_LOC_43/a_8_24# VSS VDD AND2X1_LOC_22/Y AND2X1_LOC_43/B AND2X1_LOC

XOR2X1_LOC_296 OR2X1_LOC_296/a_8_216# OR2X1_LOC_296/a_36_216# OR2X1_LOC_296/Y VSS VDD AND2X1_LOC_56/B AND2X1_LOC_43/B OR2X1_LOC

XAND2X1_LOC_136 AND2X1_LOC_136/a_36_24# OR2X1_LOC_138/A AND2X1_LOC_136/a_8_24# VSS VDD AND2X1_LOC_3/Y AND2X1_LOC_43/B AND2X1_LOC

XAND2X1_LOC_684 AND2X1_LOC_684/a_36_24# OR2X1_LOC_686/A AND2X1_LOC_684/a_8_24# VSS VDD AND2X1_LOC_12/Y AND2X1_LOC_43/B AND2X1_LOC

XAND2X1_LOC_272 AND2X1_LOC_272/a_36_24# OR2X1_LOC_541/A AND2X1_LOC_272/a_8_24# VSS VDD AND2X1_LOC_31/Y AND2X1_LOC_43/B AND2X1_LOC

XAND2X1_LOC_827 AND2X1_LOC_827/a_36_24# OR2X1_LOC_838/B AND2X1_LOC_827/a_8_24# VSS VDD AND2X1_LOC_43/B OR2X1_LOC_375/A AND2X1_LOC

XAND2X1_LOC_419 AND2X1_LOC_419/a_36_24# OR2X1_LOC_506/A AND2X1_LOC_419/a_8_24# VSS VDD AND2X1_LOC_36/Y AND2X1_LOC_43/B AND2X1_LOC

XOR2X1_LOC_378 OR2X1_LOC_378/a_8_216# OR2X1_LOC_378/a_36_216# OR2X1_LOC_378/Y VSS VDD OR2X1_LOC_378/A AND2X1_LOC_43/B OR2X1_LOC

XAND2X1_LOC_93 AND2X1_LOC_93/a_36_24# OR2X1_LOC_98/B AND2X1_LOC_93/a_8_24# VSS VDD OR2X1_LOC_66/A AND2X1_LOC_92/Y AND2X1_LOC

XAND2X1_LOC_387 AND2X1_LOC_387/a_36_24# OR2X1_LOC_389/A AND2X1_LOC_387/a_8_24# VSS VDD AND2X1_LOC_92/Y AND2X1_LOC_387/B AND2X1_LOC

XAND2X1_LOC_422 AND2X1_LOC_422/a_36_24# OR2X1_LOC_448/A AND2X1_LOC_422/a_8_24# VSS VDD AND2X1_LOC_12/Y AND2X1_LOC_92/Y AND2X1_LOC

XAND2X1_LOC_628 AND2X1_LOC_628/a_36_24# OR2X1_LOC_630/B AND2X1_LOC_628/a_8_24# VSS VDD AND2X1_LOC_47/Y AND2X1_LOC_92/Y AND2X1_LOC

XAND2X1_LOC_268 AND2X1_LOC_268/a_36_24# OR2X1_LOC_269/A AND2X1_LOC_268/a_8_24# VSS VDD AND2X1_LOC_36/Y AND2X1_LOC_92/Y AND2X1_LOC

XOR2X1_LOC_144 OR2X1_LOC_144/a_8_216# OR2X1_LOC_144/a_36_216# OR2X1_LOC_144/Y VSS VDD OR2X1_LOC_696/A OR2X1_LOC_59/Y OR2X1_LOC

XOR2X1_LOC_306 OR2X1_LOC_306/a_8_216# OR2X1_LOC_306/a_36_216# OR2X1_LOC_306/Y VSS VDD OR2X1_LOC_696/A OR2X1_LOC_22/Y OR2X1_LOC

XAND2X1_LOC_502 AND2X1_LOC_502/a_36_24# OR2X1_LOC_503/A AND2X1_LOC_502/a_8_24# VSS VDD OR2X1_LOC_89/A OR2X1_LOC_696/A AND2X1_LOC

XOR2X1_LOC_696 OR2X1_LOC_696/a_8_216# OR2X1_LOC_696/a_36_216# OR2X1_LOC_696/Y VSS VDD OR2X1_LOC_696/A OR2X1_LOC_26/Y OR2X1_LOC

XAND2X1_LOC_818 AND2X1_LOC_818/a_36_24# OR2X1_LOC_820/B AND2X1_LOC_818/a_8_24# VSS VDD OR2X1_LOC_6/A OR2X1_LOC_696/A AND2X1_LOC

XOR2X1_LOC_588 OR2X1_LOC_588/a_8_216# OR2X1_LOC_588/a_36_216# OR2X1_LOC_588/Y VSS VDD OR2X1_LOC_588/A OR2X1_LOC_696/A OR2X1_LOC

XOR2X1_LOC_376 OR2X1_LOC_376/a_8_216# OR2X1_LOC_376/a_36_216# OR2X1_LOC_376/Y VSS VDD OR2X1_LOC_376/A OR2X1_LOC_696/A OR2X1_LOC

XOR2X1_LOC_322 OR2X1_LOC_322/a_8_216# OR2X1_LOC_322/a_36_216# OR2X1_LOC_322/Y VSS VDD OR2X1_LOC_696/A OR2X1_LOC_44/Y OR2X1_LOC

XOR2X1_LOC_164 OR2X1_LOC_164/a_8_216# OR2X1_LOC_164/a_36_216# OR2X1_LOC_164/Y VSS VDD OR2X1_LOC_696/A OR2X1_LOC_18/Y OR2X1_LOC

XAND2X1_LOC_672 AND2X1_LOC_672/a_36_24# OR2X1_LOC_673/A AND2X1_LOC_672/a_8_24# VSS VDD OR2X1_LOC_375/A AND2X1_LOC_672/B AND2X1_LOC

XOR2X1_LOC_693 OR2X1_LOC_693/a_8_216# OR2X1_LOC_693/a_36_216# OR2X1_LOC_693/Y VSS VDD OR2X1_LOC_36/Y OR2X1_LOC_46/A OR2X1_LOC

XAND2X1_LOC_377 AND2X1_LOC_377/a_36_24# AND2X1_LOC_377/Y AND2X1_LOC_377/a_8_24# VSS VDD AND2X1_LOC_3/Y OR2X1_LOC_46/A AND2X1_LOC

XOR2X1_LOC_699 OR2X1_LOC_699/a_8_216# OR2X1_LOC_699/a_36_216# OR2X1_LOC_748/A VSS VDD OR2X1_LOC_158/A OR2X1_LOC_46/A OR2X1_LOC

XOR2X1_LOC_82 OR2X1_LOC_82/a_8_216# OR2X1_LOC_82/a_36_216# OR2X1_LOC_83/A VSS VDD OR2X1_LOC_80/A OR2X1_LOC_46/A OR2X1_LOC

XOR2X1_LOC_77 OR2X1_LOC_77/a_8_216# OR2X1_LOC_77/a_36_216# OR2X1_LOC_89/A VSS VDD OR2X1_LOC_54/Y OR2X1_LOC_46/A OR2X1_LOC

XOR2X1_LOC_23 OR2X1_LOC_23/a_8_216# OR2X1_LOC_23/a_36_216# OR2X1_LOC_45/B VSS VDD OR2X1_LOC_46/A OR2X1_LOC_6/B OR2X1_LOC

XOR2X1_LOC_49 OR2X1_LOC_49/a_8_216# OR2X1_LOC_49/a_36_216# OR2X1_LOC_52/B VSS VDD OR2X1_LOC_49/A OR2X1_LOC_46/A OR2X1_LOC

XOR2X1_LOC_619 OR2X1_LOC_619/a_8_216# OR2X1_LOC_619/a_36_216# OR2X1_LOC_619/Y VSS VDD OR2X1_LOC_618/Y OR2X1_LOC_36/Y OR2X1_LOC

XAND2X1_LOC_150 AND2X1_LOC_150/a_36_24# OR2X1_LOC_151/A AND2X1_LOC_150/a_8_24# VSS VDD AND2X1_LOC_42/B OR2X1_LOC_235/B AND2X1_LOC

XAND2X1_LOC_73 AND2X1_LOC_73/a_36_24# OR2X1_LOC_185/A AND2X1_LOC_73/a_8_24# VSS VDD OR2X1_LOC_62/B AND2X1_LOC_42/B AND2X1_LOC

XAND2X1_LOC_85 AND2X1_LOC_85/a_36_24# AND2X1_LOC_86/B AND2X1_LOC_85/a_8_24# VSS VDD AND2X1_LOC_18/Y AND2X1_LOC_42/B AND2X1_LOC

XAND2X1_LOC_126 AND2X1_LOC_126/a_36_24# OR2X1_LOC_160/A AND2X1_LOC_126/a_8_24# VSS VDD OR2X1_LOC_19/B AND2X1_LOC_42/B AND2X1_LOC

XAND2X1_LOC_38 AND2X1_LOC_38/a_36_24# OR2X1_LOC_154/A AND2X1_LOC_38/a_8_24# VSS VDD OR2X1_LOC_80/A AND2X1_LOC_42/B AND2X1_LOC

XAND2X1_LOC_129 AND2X1_LOC_129/a_36_24# OR2X1_LOC_130/A AND2X1_LOC_129/a_8_24# VSS VDD OR2X1_LOC_49/A AND2X1_LOC_42/B AND2X1_LOC

XAND2X1_LOC_263 AND2X1_LOC_263/a_36_24# OR2X1_LOC_266/A AND2X1_LOC_263/a_8_24# VSS VDD AND2X1_LOC_22/Y AND2X1_LOC_42/B AND2X1_LOC

XAND2X1_LOC_412 AND2X1_LOC_412/a_36_24# OR2X1_LOC_634/A AND2X1_LOC_412/a_8_24# VSS VDD AND2X1_LOC_42/B AND2X1_LOC_44/Y AND2X1_LOC

XAND2X1_LOC_255 AND2X1_LOC_255/a_36_24# OR2X1_LOC_541/B AND2X1_LOC_255/a_8_24# VSS VDD AND2X1_LOC_42/B OR2X1_LOC_375/A AND2X1_LOC

XAND2X1_LOC_277 AND2X1_LOC_277/a_36_24# OR2X1_LOC_633/A AND2X1_LOC_277/a_8_24# VSS VDD AND2X1_LOC_42/B AND2X1_LOC_47/Y AND2X1_LOC

XAND2X1_LOC_245 AND2X1_LOC_245/a_36_24# OR2X1_LOC_777/B AND2X1_LOC_245/a_8_24# VSS VDD OR2X1_LOC_66/A AND2X1_LOC_42/B AND2X1_LOC

XOR2X1_LOC_548 OR2X1_LOC_548/a_8_216# OR2X1_LOC_548/a_36_216# OR2X1_LOC_549/A VSS VDD OR2X1_LOC_548/A OR2X1_LOC_548/B OR2X1_LOC

XAND2X1_LOC_382 AND2X1_LOC_382/a_36_24# OR2X1_LOC_391/B AND2X1_LOC_382/a_8_24# VSS VDD OR2X1_LOC_80/A AND2X1_LOC_817/B AND2X1_LOC

XOR2X1_LOC_387 OR2X1_LOC_387/a_8_216# OR2X1_LOC_387/a_36_216# OR2X1_LOC_387/Y VSS VDD OR2X1_LOC_387/A OR2X1_LOC_92/Y OR2X1_LOC

XAND2X1_LOC_596 AND2X1_LOC_596/a_36_24# OR2X1_LOC_597/A AND2X1_LOC_596/a_8_24# VSS VDD OR2X1_LOC_44/Y OR2X1_LOC_421/A AND2X1_LOC

XOR2X1_LOC_329 OR2X1_LOC_329/a_8_216# OR2X1_LOC_329/a_36_216# OR2X1_LOC_329/Y VSS VDD OR2X1_LOC_421/A OR2X1_LOC_329/B OR2X1_LOC

XOR2X1_LOC_421 OR2X1_LOC_421/a_8_216# OR2X1_LOC_421/a_36_216# OR2X1_LOC_421/Y VSS VDD OR2X1_LOC_421/A OR2X1_LOC_91/A OR2X1_LOC

XOR2X1_LOC_304 OR2X1_LOC_304/a_8_216# OR2X1_LOC_304/a_36_216# OR2X1_LOC_304/Y VSS VDD OR2X1_LOC_428/A OR2X1_LOC_53/Y OR2X1_LOC

XOR2X1_LOC_56 OR2X1_LOC_56/a_8_216# OR2X1_LOC_56/a_36_216# OR2X1_LOC_56/Y VSS VDD OR2X1_LOC_56/A OR2X1_LOC_53/Y OR2X1_LOC

XOR2X1_LOC_157 OR2X1_LOC_157/a_8_216# OR2X1_LOC_157/a_36_216# OR2X1_LOC_158/A VSS VDD OR2X1_LOC_17/Y OR2X1_LOC_2/Y OR2X1_LOC

XOR2X1_LOC_70 OR2X1_LOC_70/a_8_216# OR2X1_LOC_70/a_36_216# OR2X1_LOC_70/Y VSS VDD OR2X1_LOC_70/A OR2X1_LOC_2/Y OR2X1_LOC

XOR2X1_LOC_3 OR2X1_LOC_3/a_8_216# OR2X1_LOC_3/a_36_216# OR2X1_LOC_3/Y VSS VDD OR2X1_LOC_2/Y OR2X1_LOC_3/B OR2X1_LOC

XOR2X1_LOC_40 OR2X1_LOC_40/a_8_216# OR2X1_LOC_40/a_36_216# OR2X1_LOC_40/Y VSS VDD OR2X1_LOC_25/Y OR2X1_LOC_2/Y OR2X1_LOC

XOR2X1_LOC_694 OR2X1_LOC_694/a_8_216# OR2X1_LOC_694/a_36_216# OR2X1_LOC_694/Y VSS VDD OR2X1_LOC_426/A OR2X1_LOC_427/A OR2X1_LOC

XOR2X1_LOC_426 OR2X1_LOC_426/a_8_216# OR2X1_LOC_426/a_36_216# OR2X1_LOC_426/Y VSS VDD OR2X1_LOC_426/A OR2X1_LOC_426/B OR2X1_LOC

XAND2X1_LOC_51 AND2X1_LOC_51/a_36_24# AND2X1_LOC_51/Y AND2X1_LOC_51/a_8_24# VSS VDD AND2X1_LOC_51/A AND2X1_LOC_50/Y AND2X1_LOC

XAND2X1_LOC_31 AND2X1_LOC_31/a_36_24# AND2X1_LOC_31/Y AND2X1_LOC_31/a_8_24# VSS VDD AND2X1_LOC_1/Y AND2X1_LOC_51/A AND2X1_LOC

XAND2X1_LOC_44 AND2X1_LOC_44/a_36_24# AND2X1_LOC_44/Y AND2X1_LOC_44/a_8_24# VSS VDD AND2X1_LOC_17/Y AND2X1_LOC_51/A AND2X1_LOC

XAND2X1_LOC_47 AND2X1_LOC_47/a_36_24# AND2X1_LOC_47/Y AND2X1_LOC_47/a_8_24# VSS VDD AND2X1_LOC_25/Y AND2X1_LOC_51/A AND2X1_LOC

XAND2X1_LOC_753 AND2X1_LOC_753/a_36_24# OR2X1_LOC_790/B AND2X1_LOC_753/a_8_24# VSS VDD OR2X1_LOC_185/Y AND2X1_LOC_753/B AND2X1_LOC

XAND2X1_LOC_582 AND2X1_LOC_582/a_36_24# OR2X1_LOC_635/A AND2X1_LOC_582/a_8_24# VSS VDD OR2X1_LOC_161/B AND2X1_LOC_582/B AND2X1_LOC

XAND2X1_LOC_763 AND2X1_LOC_763/a_36_24# OR2X1_LOC_769/B AND2X1_LOC_763/a_8_24# VSS VDD AND2X1_LOC_48/A AND2X1_LOC_763/B AND2X1_LOC

XOR2X1_LOC_409 OR2X1_LOC_409/a_8_216# OR2X1_LOC_409/a_36_216# OR2X1_LOC_409/Y VSS VDD OR2X1_LOC_408/Y OR2X1_LOC_409/B OR2X1_LOC

XOR2X1_LOC_430 OR2X1_LOC_430/a_8_216# OR2X1_LOC_430/a_36_216# OR2X1_LOC_430/Y VSS VDD OR2X1_LOC_429/Y OR2X1_LOC_604/A OR2X1_LOC

XOR2X1_LOC_51 OR2X1_LOC_51/a_8_216# OR2X1_LOC_51/a_36_216# OR2X1_LOC_51/Y VSS VDD OR2X1_LOC_70/A OR2X1_LOC_51/B OR2X1_LOC

XOR2X1_LOC_95 OR2X1_LOC_95/a_8_216# OR2X1_LOC_95/a_36_216# OR2X1_LOC_95/Y VSS VDD OR2X1_LOC_70/A OR2X1_LOC_11/Y OR2X1_LOC

XOR2X1_LOC_64 OR2X1_LOC_64/a_8_216# OR2X1_LOC_64/a_36_216# OR2X1_LOC_64/Y VSS VDD OR2X1_LOC_70/A OR2X1_LOC_22/A OR2X1_LOC

XAND2X1_LOC_157 AND2X1_LOC_157/a_36_24# OR2X1_LOC_375/A AND2X1_LOC_157/a_8_24# VSS VDD AND2X1_LOC_2/Y AND2X1_LOC_17/Y AND2X1_LOC

XAND2X1_LOC_36 AND2X1_LOC_36/a_36_24# AND2X1_LOC_36/Y AND2X1_LOC_36/a_8_24# VSS VDD AND2X1_LOC_17/Y AND2X1_LOC_21/Y AND2X1_LOC

XAND2X1_LOC_18 AND2X1_LOC_18/a_36_24# AND2X1_LOC_18/Y AND2X1_LOC_18/a_8_24# VSS VDD AND2X1_LOC_11/Y AND2X1_LOC_17/Y AND2X1_LOC

XOR2X1_LOC_801 OR2X1_LOC_801/a_8_216# OR2X1_LOC_801/a_36_216# OR2X1_LOC_809/B VSS VDD OR2X1_LOC_800/Y OR2X1_LOC_801/B OR2X1_LOC

XOR2X1_LOC_513 OR2X1_LOC_513/a_8_216# OR2X1_LOC_513/a_36_216# OR2X1_LOC_513/Y VSS VDD OR2X1_LOC_512/Y OR2X1_LOC_779/B OR2X1_LOC

XOR2X1_LOC_276 OR2X1_LOC_276/a_8_216# OR2X1_LOC_276/a_36_216# OR2X1_LOC_473/A VSS VDD OR2X1_LOC_276/A OR2X1_LOC_276/B OR2X1_LOC

XAND2X1_LOC_100 AND2X1_LOC_100/a_36_24# AND2X1_LOC_101/B AND2X1_LOC_100/a_8_24# VSS VDD OR2X1_LOC_86/Y OR2X1_LOC_88/Y AND2X1_LOC

XOR2X1_LOC_104 OR2X1_LOC_104/a_8_216# OR2X1_LOC_104/a_36_216# OR2X1_LOC_600/A VSS VDD OR2X1_LOC_8/Y OR2X1_LOC_6/B OR2X1_LOC

XOR2X1_LOC_126 OR2X1_LOC_126/a_8_216# OR2X1_LOC_126/a_36_216# OR2X1_LOC_744/A VSS VDD OR2X1_LOC_85/A OR2X1_LOC_6/B OR2X1_LOC

XAND2X1_LOC_490 AND2X1_LOC_490/a_36_24# OR2X1_LOC_557/A AND2X1_LOC_490/a_8_24# VSS VDD OR2X1_LOC_6/B AND2X1_LOC_86/B AND2X1_LOC

XAND2X1_LOC_19 AND2X1_LOC_19/a_36_24# AND2X1_LOC_19/Y AND2X1_LOC_19/a_8_24# VSS VDD OR2X1_LOC_6/B OR2X1_LOC_68/B AND2X1_LOC

XOR2X1_LOC_6 OR2X1_LOC_6/a_8_216# OR2X1_LOC_6/a_36_216# OR2X1_LOC_7/A VSS VDD OR2X1_LOC_6/A OR2X1_LOC_6/B OR2X1_LOC

XAND2X1_LOC_256 AND2X1_LOC_256/a_36_24# OR2X1_LOC_344/A AND2X1_LOC_256/a_8_24# VSS VDD OR2X1_LOC_6/B OR2X1_LOC_541/B AND2X1_LOC

XOR2X1_LOC_748 OR2X1_LOC_748/a_8_216# OR2X1_LOC_748/a_36_216# OR2X1_LOC_748/Y VSS VDD OR2X1_LOC_748/A OR2X1_LOC_6/B OR2X1_LOC

XOR2X1_LOC_129 OR2X1_LOC_129/a_8_216# OR2X1_LOC_129/a_36_216# OR2X1_LOC_589/A VSS VDD OR2X1_LOC_85/A OR2X1_LOC_80/A OR2X1_LOC

XAND2X1_LOC_133 AND2X1_LOC_133/a_36_24# OR2X1_LOC_161/B AND2X1_LOC_133/a_8_24# VSS VDD AND2X1_LOC_8/Y OR2X1_LOC_80/A AND2X1_LOC

XOR2X1_LOC_80 OR2X1_LOC_80/a_8_216# OR2X1_LOC_80/a_36_216# OR2X1_LOC_80/Y VSS VDD OR2X1_LOC_80/A OR2X1_LOC_6/A OR2X1_LOC

XAND2X1_LOC_49 AND2X1_LOC_49/a_36_24# OR2X1_LOC_87/A AND2X1_LOC_49/a_8_24# VSS VDD OR2X1_LOC_377/A OR2X1_LOC_80/A AND2X1_LOC

XOR2X1_LOC_29 OR2X1_LOC_29/a_8_216# OR2X1_LOC_29/a_36_216# OR2X1_LOC_32/B VSS VDD OR2X1_LOC_80/A OR2X1_LOC_8/Y OR2X1_LOC

XAND2X1_LOC_236 AND2X1_LOC_236/a_36_24# OR2X1_LOC_269/B AND2X1_LOC_236/a_8_24# VSS VDD OR2X1_LOC_68/B OR2X1_LOC_80/A AND2X1_LOC

XOR2X1_LOC_291 OR2X1_LOC_291/a_8_216# OR2X1_LOC_291/a_36_216# OR2X1_LOC_291/Y VSS VDD OR2X1_LOC_291/A OR2X1_LOC_36/Y OR2X1_LOC

XOR2X1_LOC_824 OR2X1_LOC_824/a_8_216# OR2X1_LOC_824/a_36_216# OR2X1_LOC_824/Y VSS VDD OR2X1_LOC_291/A OR2X1_LOC_26/Y OR2X1_LOC

XOR2X1_LOC_234 OR2X1_LOC_234/a_8_216# OR2X1_LOC_234/a_36_216# OR2X1_LOC_234/Y VSS VDD OR2X1_LOC_291/A OR2X1_LOC_47/Y OR2X1_LOC

XAND2X1_LOC_461 AND2X1_LOC_461/a_36_24# AND2X1_LOC_462/B AND2X1_LOC_461/a_8_24# VSS VDD OR2X1_LOC_411/Y OR2X1_LOC_413/Y AND2X1_LOC

XOR2X1_LOC_691 OR2X1_LOC_691/a_8_216# OR2X1_LOC_691/a_36_216# OR2X1_LOC_691/Y VSS VDD OR2X1_LOC_691/A OR2X1_LOC_691/B OR2X1_LOC

XAND2X1_LOC_323 AND2X1_LOC_323/a_36_24# OR2X1_LOC_325/A AND2X1_LOC_323/a_8_24# VSS VDD AND2X1_LOC_95/Y AND2X1_LOC_110/Y AND2X1_LOC

XAND2X1_LOC_527 AND2X1_LOC_527/a_36_24# OR2X1_LOC_547/B AND2X1_LOC_527/a_8_24# VSS VDD AND2X1_LOC_64/Y AND2X1_LOC_110/Y AND2X1_LOC

XAND2X1_LOC_111 AND2X1_LOC_111/a_36_24# OR2X1_LOC_112/A AND2X1_LOC_111/a_8_24# VSS VDD AND2X1_LOC_31/Y AND2X1_LOC_110/Y AND2X1_LOC

XAND2X1_LOC_515 AND2X1_LOC_515/a_36_24# OR2X1_LOC_516/A AND2X1_LOC_515/a_8_24# VSS VDD OR2X1_LOC_417/Y AND2X1_LOC_514/Y AND2X1_LOC

XOR2X1_LOC_750 OR2X1_LOC_750/a_8_216# OR2X1_LOC_750/a_36_216# OR2X1_LOC_750/Y VSS VDD OR2X1_LOC_750/A OR2X1_LOC_161/A OR2X1_LOC

XOR2X1_LOC_814 OR2X1_LOC_814/a_8_216# OR2X1_LOC_814/a_36_216# OR2X1_LOC_814/Y VSS VDD OR2X1_LOC_814/A OR2X1_LOC_756/B OR2X1_LOC

XAND2X1_LOC_309 AND2X1_LOC_309/a_36_24# OR2X1_LOC_335/B AND2X1_LOC_309/a_8_24# VSS VDD AND2X1_LOC_22/Y OR2X1_LOC_814/A AND2X1_LOC

XAND2X1_LOC_283 AND2X1_LOC_283/a_36_24# OR2X1_LOC_286/B AND2X1_LOC_283/a_8_24# VSS VDD OR2X1_LOC_66/A OR2X1_LOC_814/A AND2X1_LOC

XAND2X1_LOC_488 AND2X1_LOC_488/a_36_24# OR2X1_LOC_489/A AND2X1_LOC_488/a_8_24# VSS VDD OR2X1_LOC_375/A OR2X1_LOC_814/A AND2X1_LOC

XAND2X1_LOC_289 AND2X1_LOC_289/a_36_24# OR2X1_LOC_333/A AND2X1_LOC_289/a_8_24# VSS VDD AND2X1_LOC_51/Y OR2X1_LOC_814/A AND2X1_LOC

XAND2X1_LOC_417 AND2X1_LOC_417/a_36_24# OR2X1_LOC_446/B AND2X1_LOC_417/a_8_24# VSS VDD AND2X1_LOC_47/Y OR2X1_LOC_814/A AND2X1_LOC

XAND2X1_LOC_226 AND2X1_LOC_226/a_36_24# OR2X1_LOC_227/A AND2X1_LOC_226/a_8_24# VSS VDD AND2X1_LOC_18/Y OR2X1_LOC_814/A AND2X1_LOC

XOR2X1_LOC_133 OR2X1_LOC_133/a_8_216# OR2X1_LOC_133/a_36_216# OR2X1_LOC_427/A VSS VDD OR2X1_LOC_49/A OR2X1_LOC_8/Y OR2X1_LOC

XAND2X1_LOC_80 AND2X1_LOC_80/a_36_24# AND2X1_LOC_81/B AND2X1_LOC_80/a_8_24# VSS VDD OR2X1_LOC_68/B OR2X1_LOC_49/A AND2X1_LOC

XAND2X1_LOC_82 AND2X1_LOC_82/a_36_24# AND2X1_LOC_82/Y AND2X1_LOC_82/a_8_24# VSS VDD OR2X1_LOC_377/A OR2X1_LOC_49/A AND2X1_LOC

XAND2X1_LOC_29 AND2X1_LOC_29/a_36_24# OR2X1_LOC_87/B AND2X1_LOC_29/a_8_24# VSS VDD AND2X1_LOC_8/Y OR2X1_LOC_49/A AND2X1_LOC

XOR2X1_LOC_236 OR2X1_LOC_236/a_8_216# OR2X1_LOC_236/a_36_216# OR2X1_LOC_428/A VSS VDD OR2X1_LOC_49/A OR2X1_LOC_6/A OR2X1_LOC

XOR2X1_LOC_382 OR2X1_LOC_382/a_8_216# OR2X1_LOC_382/a_36_216# OR2X1_LOC_382/Y VSS VDD OR2X1_LOC_382/A OR2X1_LOC_49/A OR2X1_LOC

XOR2X1_LOC_38 OR2X1_LOC_38/a_8_216# OR2X1_LOC_38/a_36_216# OR2X1_LOC_39/A VSS VDD OR2X1_LOC_85/A OR2X1_LOC_49/A OR2X1_LOC

XOR2X1_LOC_847 OR2X1_LOC_847/a_8_216# OR2X1_LOC_847/a_36_216# OR2X1_LOC_848/A VSS VDD OR2X1_LOC_847/A OR2X1_LOC_847/B OR2X1_LOC

XAND2X1_LOC_10 AND2X1_LOC_10/a_36_24# AND2X1_LOC_41/A AND2X1_LOC_10/a_8_24# VSS VDD AND2X1_LOC_8/Y OR2X1_LOC_62/B AND2X1_LOC

XAND2X1_LOC_159 AND2X1_LOC_159/a_36_24# OR2X1_LOC_161/A AND2X1_LOC_159/a_8_24# VSS VDD OR2X1_LOC_68/B OR2X1_LOC_62/B AND2X1_LOC

XAND2X1_LOC_15 AND2X1_LOC_15/a_36_24# OR2X1_LOC_78/B AND2X1_LOC_15/a_8_24# VSS VDD OR2X1_LOC_62/B OR2X1_LOC_377/A AND2X1_LOC

XOR2X1_LOC_278 OR2X1_LOC_278/a_8_216# OR2X1_LOC_278/a_36_216# OR2X1_LOC_278/Y VSS VDD OR2X1_LOC_278/A OR2X1_LOC_62/B OR2X1_LOC

XAND2X1_LOC_246 AND2X1_LOC_246/a_36_24# OR2X1_LOC_342/B AND2X1_LOC_246/a_8_24# VSS VDD OR2X1_LOC_62/B OR2X1_LOC_777/B AND2X1_LOC

XOR2X1_LOC_102 OR2X1_LOC_102/a_8_216# OR2X1_LOC_102/a_36_216# OR2X1_LOC_485/A VSS VDD OR2X1_LOC_54/Y OR2X1_LOC_8/Y OR2X1_LOC

XAND2X1_LOC_94 AND2X1_LOC_94/a_36_24# AND2X1_LOC_94/Y AND2X1_LOC_94/a_8_24# VSS VDD OR2X1_LOC_377/A OR2X1_LOC_54/Y AND2X1_LOC

XOR2X1_LOC_90 OR2X1_LOC_90/a_8_216# OR2X1_LOC_90/a_36_216# OR2X1_LOC_91/A VSS VDD OR2X1_LOC_54/Y OR2X1_LOC_85/A OR2X1_LOC

XAND2X1_LOC_611 AND2X1_LOC_611/a_36_24# AND2X1_LOC_612/B AND2X1_LOC_611/a_8_24# VSS VDD OR2X1_LOC_68/B OR2X1_LOC_54/Y AND2X1_LOC

XOR2X1_LOC_55 OR2X1_LOC_55/a_8_216# OR2X1_LOC_55/a_36_216# OR2X1_LOC_56/A VSS VDD OR2X1_LOC_54/Y OR2X1_LOC_6/A OR2X1_LOC

XAND2X1_LOC_819 AND2X1_LOC_819/a_36_24# AND2X1_LOC_820/B AND2X1_LOC_819/a_8_24# VSS VDD AND2X1_LOC_47/Y OR2X1_LOC_54/Y AND2X1_LOC

XOR2X1_LOC_136 OR2X1_LOC_136/a_8_216# OR2X1_LOC_136/a_36_216# OR2X1_LOC_136/Y VSS VDD OR2X1_LOC_43/A OR2X1_LOC_3/Y OR2X1_LOC

XOR2X1_LOC_684 OR2X1_LOC_684/a_8_216# OR2X1_LOC_684/a_36_216# OR2X1_LOC_684/Y VSS VDD OR2X1_LOC_43/A OR2X1_LOC_12/Y OR2X1_LOC

XAND2X1_LOC_378 AND2X1_LOC_378/a_36_24# OR2X1_LOC_459/A AND2X1_LOC_378/a_8_24# VSS VDD OR2X1_LOC_43/A AND2X1_LOC_377/Y AND2X1_LOC

XOR2X1_LOC_272 OR2X1_LOC_272/a_8_216# OR2X1_LOC_272/a_36_216# OR2X1_LOC_272/Y VSS VDD OR2X1_LOC_43/A OR2X1_LOC_31/Y OR2X1_LOC

XOR2X1_LOC_827 OR2X1_LOC_827/a_8_216# OR2X1_LOC_827/a_36_216# OR2X1_LOC_827/Y VSS VDD OR2X1_LOC_158/A OR2X1_LOC_43/A OR2X1_LOC

XOR2X1_LOC_419 OR2X1_LOC_419/a_8_216# OR2X1_LOC_419/a_36_216# OR2X1_LOC_419/Y VSS VDD OR2X1_LOC_43/A OR2X1_LOC_36/Y OR2X1_LOC

XOR2X1_LOC_43 OR2X1_LOC_43/a_8_216# OR2X1_LOC_43/a_36_216# OR2X1_LOC_43/Y VSS VDD OR2X1_LOC_43/A OR2X1_LOC_22/Y OR2X1_LOC

XAND2X1_LOC_296 AND2X1_LOC_296/a_36_24# OR2X1_LOC_297/A AND2X1_LOC_296/a_8_24# VSS VDD OR2X1_LOC_43/A OR2X1_LOC_56/A AND2X1_LOC

XOR2X1_LOC_534 OR2X1_LOC_534/a_8_216# OR2X1_LOC_534/a_36_216# OR2X1_LOC_534/Y VSS VDD OR2X1_LOC_59/Y OR2X1_LOC_43/A OR2X1_LOC

XOR2X1_LOC_490 OR2X1_LOC_490/a_8_216# OR2X1_LOC_490/a_36_216# OR2X1_LOC_490/Y VSS VDD OR2X1_LOC_86/A OR2X1_LOC_19/B OR2X1_LOC

XAND2X1_LOC_748 AND2X1_LOC_748/a_36_24# OR2X1_LOC_789/B AND2X1_LOC_748/a_8_24# VSS VDD OR2X1_LOC_19/B OR2X1_LOC_709/A AND2X1_LOC

XAND2X1_LOC_23 AND2X1_LOC_23/a_36_24# OR2X1_LOC_160/B AND2X1_LOC_23/a_8_24# VSS VDD OR2X1_LOC_19/B OR2X1_LOC_377/A AND2X1_LOC

XAND2X1_LOC_104 AND2X1_LOC_104/a_36_24# OR2X1_LOC_756/B AND2X1_LOC_104/a_8_24# VSS VDD OR2X1_LOC_19/B AND2X1_LOC_8/Y AND2X1_LOC

XOR2X1_LOC_256 OR2X1_LOC_256/a_8_216# OR2X1_LOC_256/a_36_216# OR2X1_LOC_256/Y VSS VDD OR2X1_LOC_256/A OR2X1_LOC_19/B OR2X1_LOC

XAND2X1_LOC_6 AND2X1_LOC_6/a_36_24# AND2X1_LOC_7/B AND2X1_LOC_6/a_8_24# VSS VDD OR2X1_LOC_19/B OR2X1_LOC_68/B AND2X1_LOC

XOR2X1_LOC_19 OR2X1_LOC_19/a_8_216# OR2X1_LOC_19/a_36_216# OR2X1_LOC_20/A VSS VDD OR2X1_LOC_6/A OR2X1_LOC_19/B OR2X1_LOC

XOR2X1_LOC_422 OR2X1_LOC_422/a_8_216# OR2X1_LOC_422/a_36_216# OR2X1_LOC_422/Y VSS VDD OR2X1_LOC_92/Y OR2X1_LOC_12/Y OR2X1_LOC

XOR2X1_LOC_628 OR2X1_LOC_628/a_8_216# OR2X1_LOC_628/a_36_216# OR2X1_LOC_628/Y VSS VDD OR2X1_LOC_92/Y OR2X1_LOC_47/Y OR2X1_LOC

XOR2X1_LOC_93 OR2X1_LOC_93/a_8_216# OR2X1_LOC_93/a_36_216# OR2X1_LOC_93/Y VSS VDD OR2X1_LOC_92/Y OR2X1_LOC_26/Y OR2X1_LOC

XOR2X1_LOC_268 OR2X1_LOC_268/a_8_216# OR2X1_LOC_268/a_36_216# OR2X1_LOC_268/Y VSS VDD OR2X1_LOC_92/Y OR2X1_LOC_36/Y OR2X1_LOC

XAND2X1_LOC_511 AND2X1_LOC_511/a_36_24# OR2X1_LOC_779/B AND2X1_LOC_511/a_8_24# VSS VDD AND2X1_LOC_31/Y AND2X1_LOC_48/A AND2X1_LOC

XAND2X1_LOC_519 AND2X1_LOC_519/a_36_24# OR2X1_LOC_520/A AND2X1_LOC_519/a_8_24# VSS VDD AND2X1_LOC_48/A OR2X1_LOC_375/A AND2X1_LOC

XAND2X1_LOC_692 AND2X1_LOC_692/a_36_24# OR2X1_LOC_706/B AND2X1_LOC_692/a_8_24# VSS VDD AND2X1_LOC_18/Y AND2X1_LOC_48/A AND2X1_LOC

XAND2X1_LOC_48 AND2X1_LOC_48/a_36_24# AND2X1_LOC_48/Y AND2X1_LOC_48/a_8_24# VSS VDD AND2X1_LOC_48/A AND2X1_LOC_47/Y AND2X1_LOC

XOR2X1_LOC_405 OR2X1_LOC_405/a_8_216# OR2X1_LOC_405/a_36_216# OR2X1_LOC_405/Y VSS VDD OR2X1_LOC_405/A AND2X1_LOC_48/A OR2X1_LOC

XAND2X1_LOC_398 AND2X1_LOC_398/a_36_24# OR2X1_LOC_399/A AND2X1_LOC_398/a_8_24# VSS VDD OR2X1_LOC_16/A OR2X1_LOC_585/A AND2X1_LOC

XOR2X1_LOC_625 OR2X1_LOC_625/a_8_216# OR2X1_LOC_625/a_36_216# OR2X1_LOC_625/Y VSS VDD OR2X1_LOC_585/A OR2X1_LOC_67/A OR2X1_LOC

XAND2X1_LOC_688 AND2X1_LOC_688/a_36_24# OR2X1_LOC_689/A AND2X1_LOC_688/a_8_24# VSS VDD OR2X1_LOC_39/A OR2X1_LOC_585/A AND2X1_LOC

XAND2X1_LOC_294 AND2X1_LOC_294/a_36_24# OR2X1_LOC_481/A AND2X1_LOC_294/a_8_24# VSS VDD OR2X1_LOC_13/B OR2X1_LOC_585/A AND2X1_LOC

XOR2X1_LOC_585 OR2X1_LOC_585/a_8_216# OR2X1_LOC_585/a_36_216# OR2X1_LOC_585/Y VSS VDD OR2X1_LOC_585/A OR2X1_LOC_22/Y OR2X1_LOC

XAND2X1_LOC_415 AND2X1_LOC_415/a_36_24# OR2X1_LOC_416/A AND2X1_LOC_415/a_8_24# VSS VDD OR2X1_LOC_585/A OR2X1_LOC_414/Y AND2X1_LOC

XAND2X1_LOC_588 AND2X1_LOC_588/a_36_24# OR2X1_LOC_638/B AND2X1_LOC_588/a_8_24# VSS VDD OR2X1_LOC_502/A AND2X1_LOC_588/B AND2X1_LOC

XAND2X1_LOC_376 AND2X1_LOC_376/a_36_24# OR2X1_LOC_459/B AND2X1_LOC_376/a_8_24# VSS VDD OR2X1_LOC_502/A OR2X1_LOC_375/Y AND2X1_LOC

XAND2X1_LOC_322 AND2X1_LOC_322/a_36_24# OR2X1_LOC_325/B AND2X1_LOC_322/a_8_24# VSS VDD AND2X1_LOC_44/Y OR2X1_LOC_502/A AND2X1_LOC

XAND2X1_LOC_164 AND2X1_LOC_164/a_36_24# OR2X1_LOC_168/B AND2X1_LOC_164/a_8_24# VSS VDD AND2X1_LOC_18/Y OR2X1_LOC_502/A AND2X1_LOC

XAND2X1_LOC_144 AND2X1_LOC_144/a_36_24# OR2X1_LOC_147/A AND2X1_LOC_144/a_8_24# VSS VDD AND2X1_LOC_59/Y OR2X1_LOC_502/A AND2X1_LOC

XOR2X1_LOC_818 OR2X1_LOC_818/a_8_216# OR2X1_LOC_818/a_36_216# OR2X1_LOC_818/Y VSS VDD OR2X1_LOC_502/A OR2X1_LOC_68/B OR2X1_LOC

XAND2X1_LOC_306 AND2X1_LOC_306/a_36_24# OR2X1_LOC_512/A AND2X1_LOC_306/a_8_24# VSS VDD AND2X1_LOC_22/Y OR2X1_LOC_502/A AND2X1_LOC

XAND2X1_LOC_696 AND2X1_LOC_696/a_36_24# OR2X1_LOC_708/B AND2X1_LOC_696/a_8_24# VSS VDD OR2X1_LOC_66/A OR2X1_LOC_502/A AND2X1_LOC

XOR2X1_LOC_502 OR2X1_LOC_502/a_8_216# OR2X1_LOC_502/a_36_216# OR2X1_LOC_502/Y VSS VDD OR2X1_LOC_502/A OR2X1_LOC_78/A OR2X1_LOC

XOR2X1_LOC_155 OR2X1_LOC_155/a_8_216# OR2X1_LOC_155/a_36_216# OR2X1_LOC_156/A VSS VDD OR2X1_LOC_155/A OR2X1_LOC_87/A OR2X1_LOC

XAND2X1_LOC_743 AND2X1_LOC_743/a_36_24# OR2X1_LOC_780/B AND2X1_LOC_743/a_8_24# VSS VDD AND2X1_LOC_3/Y OR2X1_LOC_155/A AND2X1_LOC

XAND2X1_LOC_681 AND2X1_LOC_681/a_36_24# OR2X1_LOC_685/B AND2X1_LOC_681/a_8_24# VSS VDD AND2X1_LOC_31/Y OR2X1_LOC_155/A AND2X1_LOC

XOR2X1_LOC_407 OR2X1_LOC_407/a_8_216# OR2X1_LOC_407/a_36_216# OR2X1_LOC_828/B VSS VDD OR2X1_LOC_155/A AND2X1_LOC_56/B OR2X1_LOC

XAND2X1_LOC_273 AND2X1_LOC_273/a_36_24# OR2X1_LOC_831/B AND2X1_LOC_273/a_8_24# VSS VDD AND2X1_LOC_36/Y OR2X1_LOC_155/A AND2X1_LOC

XAND2X1_LOC_433 AND2X1_LOC_433/a_36_24# OR2X1_LOC_435/A AND2X1_LOC_433/a_8_24# VSS VDD AND2X1_LOC_70/Y OR2X1_LOC_155/A AND2X1_LOC

XOR2X1_LOC_369 OR2X1_LOC_369/a_8_216# OR2X1_LOC_369/a_36_216# OR2X1_LOC_369/Y VSS VDD OR2X1_LOC_426/B OR2X1_LOC_22/Y OR2X1_LOC

XAND2X1_LOC_121 AND2X1_LOC_121/a_36_24# OR2X1_LOC_122/A AND2X1_LOC_121/a_8_24# VSS VDD OR2X1_LOC_426/B OR2X1_LOC_666/A AND2X1_LOC

XOR2X1_LOC_299 OR2X1_LOC_299/a_8_216# OR2X1_LOC_299/a_36_216# OR2X1_LOC_299/Y VSS VDD OR2X1_LOC_426/B OR2X1_LOC_12/Y OR2X1_LOC

XAND2X1_LOC_606 AND2X1_LOC_606/a_36_24# OR2X1_LOC_607/A AND2X1_LOC_606/a_8_24# VSS VDD OR2X1_LOC_485/A OR2X1_LOC_426/B AND2X1_LOC

XOR2X1_LOC_300 OR2X1_LOC_300/a_8_216# OR2X1_LOC_300/a_36_216# OR2X1_LOC_300/Y VSS VDD OR2X1_LOC_426/B OR2X1_LOC_59/Y OR2X1_LOC

XOR2X1_LOC_458 OR2X1_LOC_458/a_8_216# OR2X1_LOC_458/a_36_216# OR2X1_LOC_464/A VSS VDD OR2X1_LOC_374/Y OR2X1_LOC_458/B OR2X1_LOC

XOR2X1_LOC_63 OR2X1_LOC_63/a_8_216# OR2X1_LOC_63/a_36_216# OR2X1_LOC_65/B VSS VDD OR2X1_LOC_71/A OR2X1_LOC_8/Y OR2X1_LOC

XAND2X1_LOC_371 AND2X1_LOC_371/a_36_24# OR2X1_LOC_778/B AND2X1_LOC_371/a_8_24# VSS VDD OR2X1_LOC_68/B AND2X1_LOC_31/Y AND2X1_LOC

XAND2X1_LOC_71 AND2X1_LOC_71/a_36_24# AND2X1_LOC_72/B AND2X1_LOC_71/a_8_24# VSS VDD OR2X1_LOC_68/B OR2X1_LOC_235/B AND2X1_LOC

XAND2X1_LOC_310 AND2X1_LOC_310/a_36_24# OR2X1_LOC_335/A AND2X1_LOC_310/a_8_24# VSS VDD OR2X1_LOC_68/B AND2X1_LOC_40/Y AND2X1_LOC

XAND2X1_LOC_57 AND2X1_LOC_57/a_36_24# AND2X1_LOC_57/Y AND2X1_LOC_57/a_8_24# VSS VDD OR2X1_LOC_68/B AND2X1_LOC_44/Y AND2X1_LOC

XOR2X1_LOC_68 OR2X1_LOC_68/a_8_216# OR2X1_LOC_68/a_36_216# OR2X1_LOC_68/Y VSS VDD OR2X1_LOC_87/A OR2X1_LOC_68/B OR2X1_LOC

XOR2X1_LOC_672 OR2X1_LOC_672/a_8_216# OR2X1_LOC_672/a_36_216# OR2X1_LOC_672/Y VSS VDD OR2X1_LOC_671/Y OR2X1_LOC_158/A OR2X1_LOC

XAND2X1_LOC_619 AND2X1_LOC_619/a_36_24# OR2X1_LOC_622/B AND2X1_LOC_619/a_8_24# VSS VDD AND2X1_LOC_36/Y AND2X1_LOC_619/B AND2X1_LOC

XOR2X1_LOC_263 OR2X1_LOC_263/a_8_216# OR2X1_LOC_263/a_36_216# OR2X1_LOC_813/A VSS VDD OR2X1_LOC_85/A OR2X1_LOC_22/Y OR2X1_LOC

XOR2X1_LOC_412 OR2X1_LOC_412/a_8_216# OR2X1_LOC_412/a_36_216# OR2X1_LOC_690/A VSS VDD OR2X1_LOC_44/Y OR2X1_LOC_85/A OR2X1_LOC

XOR2X1_LOC_255 OR2X1_LOC_255/a_8_216# OR2X1_LOC_255/a_36_216# OR2X1_LOC_256/A VSS VDD OR2X1_LOC_158/A OR2X1_LOC_85/A OR2X1_LOC

XOR2X1_LOC_277 OR2X1_LOC_277/a_8_216# OR2X1_LOC_277/a_36_216# OR2X1_LOC_278/A VSS VDD OR2X1_LOC_47/Y OR2X1_LOC_85/A OR2X1_LOC

XOR2X1_LOC_245 OR2X1_LOC_245/a_8_216# OR2X1_LOC_245/a_36_216# OR2X1_LOC_246/A VSS VDD OR2X1_LOC_85/A OR2X1_LOC_26/Y OR2X1_LOC

XOR2X1_LOC_85 OR2X1_LOC_85/a_8_216# OR2X1_LOC_85/a_36_216# OR2X1_LOC_86/A VSS VDD OR2X1_LOC_85/A OR2X1_LOC_18/Y OR2X1_LOC

XOR2X1_LOC_150 OR2X1_LOC_150/a_8_216# OR2X1_LOC_150/a_36_216# OR2X1_LOC_437/A VSS VDD OR2X1_LOC_71/A OR2X1_LOC_85/A OR2X1_LOC

XAND2X1_LOC_63 AND2X1_LOC_63/a_36_24# AND2X1_LOC_65/A AND2X1_LOC_63/a_8_24# VSS VDD AND2X1_LOC_8/Y OR2X1_LOC_235/B AND2X1_LOC

XAND2X1_LOC_68 AND2X1_LOC_68/a_36_24# OR2X1_LOC_69/A AND2X1_LOC_68/a_8_24# VSS VDD OR2X1_LOC_6/A OR2X1_LOC_52/B AND2X1_LOC

XOR2X1_LOC_71 OR2X1_LOC_71/a_8_216# OR2X1_LOC_71/a_36_216# OR2X1_LOC_71/Y VSS VDD OR2X1_LOC_71/A OR2X1_LOC_6/A OR2X1_LOC

XOR2X1_LOC_57 OR2X1_LOC_57/a_8_216# OR2X1_LOC_57/a_36_216# OR2X1_LOC_57/Y VSS VDD OR2X1_LOC_44/Y OR2X1_LOC_6/A OR2X1_LOC

XOR2X1_LOC_371 OR2X1_LOC_371/a_8_216# OR2X1_LOC_371/a_36_216# OR2X1_LOC_371/Y VSS VDD OR2X1_LOC_31/Y OR2X1_LOC_6/A OR2X1_LOC

XOR2X1_LOC_310 OR2X1_LOC_310/a_8_216# OR2X1_LOC_310/a_36_216# OR2X1_LOC_310/Y VSS VDD OR2X1_LOC_40/Y OR2X1_LOC_6/A OR2X1_LOC

XAND2X1_LOC_693 AND2X1_LOC_693/a_36_24# OR2X1_LOC_706/A AND2X1_LOC_693/a_8_24# VSS VDD OR2X1_LOC_377/A AND2X1_LOC_36/Y AND2X1_LOC

XAND2X1_LOC_699 AND2X1_LOC_699/a_36_24# OR2X1_LOC_709/A AND2X1_LOC_699/a_8_24# VSS VDD OR2X1_LOC_377/A OR2X1_LOC_375/A AND2X1_LOC

XOR2X1_LOC_377 OR2X1_LOC_377/a_8_216# OR2X1_LOC_377/a_36_216# OR2X1_LOC_378/A VSS VDD OR2X1_LOC_377/A OR2X1_LOC_3/Y OR2X1_LOC

XAND2X1_LOC_548 AND2X1_LOC_548/a_36_24# AND2X1_LOC_548/Y AND2X1_LOC_548/a_8_24# VSS VDD OR2X1_LOC_529/Y OR2X1_LOC_530/Y AND2X1_LOC

XOR2X1_LOC_22 OR2X1_LOC_22/a_8_216# OR2X1_LOC_22/a_36_216# OR2X1_LOC_22/Y VSS VDD OR2X1_LOC_22/A OR2X1_LOC_3/B OR2X1_LOC

XOR2X1_LOC_36 OR2X1_LOC_36/a_8_216# OR2X1_LOC_36/a_36_216# OR2X1_LOC_36/Y VSS VDD OR2X1_LOC_22/A OR2X1_LOC_17/Y OR2X1_LOC

XOR2X1_LOC_26 OR2X1_LOC_26/a_8_216# OR2X1_LOC_26/a_36_216# OR2X1_LOC_26/Y VSS VDD OR2X1_LOC_25/Y OR2X1_LOC_22/A OR2X1_LOC

XAND2X1_LOC_329 AND2X1_LOC_329/a_36_24# OR2X1_LOC_355/B AND2X1_LOC_329/a_8_24# VSS VDD OR2X1_LOC_405/A OR2X1_LOC_596/A AND2X1_LOC

XAND2X1_LOC_421 AND2X1_LOC_421/a_36_24# OR2X1_LOC_448/B AND2X1_LOC_421/a_8_24# VSS VDD AND2X1_LOC_91/B OR2X1_LOC_596/A AND2X1_LOC

XOR2X1_LOC_596 OR2X1_LOC_596/a_8_216# OR2X1_LOC_596/a_36_216# OR2X1_LOC_596/Y VSS VDD OR2X1_LOC_596/A AND2X1_LOC_44/Y OR2X1_LOC

XAND2X1_LOC_95 AND2X1_LOC_95/a_36_24# AND2X1_LOC_95/Y AND2X1_LOC_95/a_8_24# VSS VDD AND2X1_LOC_11/Y AND2X1_LOC_50/Y AND2X1_LOC

XAND2X1_LOC_12 AND2X1_LOC_12/a_36_24# AND2X1_LOC_12/Y AND2X1_LOC_12/a_8_24# VSS VDD AND2X1_LOC_1/Y AND2X1_LOC_11/Y AND2X1_LOC

XAND2X1_LOC_59 AND2X1_LOC_59/a_36_24# AND2X1_LOC_59/Y AND2X1_LOC_59/a_8_24# VSS VDD AND2X1_LOC_11/Y AND2X1_LOC_25/Y AND2X1_LOC

XAND2X1_LOC_694 AND2X1_LOC_694/a_36_24# OR2X1_LOC_707/B AND2X1_LOC_694/a_8_24# VSS VDD OR2X1_LOC_161/B AND2X1_LOC_425/Y AND2X1_LOC

XOR2X1_LOC_753 OR2X1_LOC_753/a_8_216# OR2X1_LOC_753/a_36_216# OR2X1_LOC_753/Y VSS VDD OR2X1_LOC_753/A OR2X1_LOC_816/A OR2X1_LOC

XOR2X1_LOC_12 OR2X1_LOC_12/a_8_216# OR2X1_LOC_12/a_36_216# OR2X1_LOC_12/Y VSS VDD OR2X1_LOC_11/Y OR2X1_LOC_3/B OR2X1_LOC

XOR2X1_LOC_59 OR2X1_LOC_59/a_8_216# OR2X1_LOC_59/a_36_216# OR2X1_LOC_59/Y VSS VDD OR2X1_LOC_25/Y OR2X1_LOC_11/Y OR2X1_LOC

XOR2X1_LOC_18 OR2X1_LOC_18/a_8_216# OR2X1_LOC_18/a_36_216# OR2X1_LOC_18/Y VSS VDD OR2X1_LOC_17/Y OR2X1_LOC_11/Y OR2X1_LOC

XOR2X1_LOC_31 OR2X1_LOC_31/a_8_216# OR2X1_LOC_31/a_36_216# OR2X1_LOC_31/Y VSS VDD OR2X1_LOC_51/B OR2X1_LOC_3/B OR2X1_LOC

XOR2X1_LOC_44 OR2X1_LOC_44/a_8_216# OR2X1_LOC_44/a_36_216# OR2X1_LOC_44/Y VSS VDD OR2X1_LOC_51/B OR2X1_LOC_17/Y OR2X1_LOC

XOR2X1_LOC_47 OR2X1_LOC_47/a_8_216# OR2X1_LOC_47/a_36_216# OR2X1_LOC_47/Y VSS VDD OR2X1_LOC_51/B OR2X1_LOC_25/Y OR2X1_LOC

XAND2X1_LOC_70 AND2X1_LOC_70/a_36_24# AND2X1_LOC_70/Y AND2X1_LOC_70/a_8_24# VSS VDD AND2X1_LOC_2/Y AND2X1_LOC_50/Y AND2X1_LOC

XAND2X1_LOC_40 AND2X1_LOC_40/a_36_24# AND2X1_LOC_40/Y AND2X1_LOC_40/a_8_24# VSS VDD AND2X1_LOC_2/Y AND2X1_LOC_25/Y AND2X1_LOC

XAND2X1_LOC_3 AND2X1_LOC_3/a_36_24# AND2X1_LOC_3/Y AND2X1_LOC_3/a_8_24# VSS VDD AND2X1_LOC_1/Y AND2X1_LOC_2/Y AND2X1_LOC

XAND2X1_LOC_64 AND2X1_LOC_64/a_36_24# AND2X1_LOC_64/Y AND2X1_LOC_64/a_8_24# VSS VDD AND2X1_LOC_21/Y AND2X1_LOC_50/Y AND2X1_LOC

XAND2X1_LOC_22 AND2X1_LOC_22/a_36_24# AND2X1_LOC_22/Y AND2X1_LOC_22/a_8_24# VSS VDD AND2X1_LOC_1/Y AND2X1_LOC_21/Y AND2X1_LOC

XAND2X1_LOC_26 AND2X1_LOC_26/a_36_24# OR2X1_LOC_66/A AND2X1_LOC_26/a_8_24# VSS VDD AND2X1_LOC_21/Y AND2X1_LOC_25/Y AND2X1_LOC

XAND2X1_LOC_304 AND2X1_LOC_304/a_36_24# OR2X1_LOC_307/B AND2X1_LOC_304/a_8_24# VSS VDD AND2X1_LOC_53/Y OR2X1_LOC_269/B AND2X1_LOC

XAND2X1_LOC_56 AND2X1_LOC_56/a_36_24# OR2X1_LOC_197/A AND2X1_LOC_56/a_8_24# VSS VDD AND2X1_LOC_53/Y AND2X1_LOC_56/B AND2X1_LOC

XAND2X1_LOC_409 AND2X1_LOC_409/a_36_24# OR2X1_LOC_460/A AND2X1_LOC_409/a_8_24# VSS VDD OR2X1_LOC_828/B AND2X1_LOC_409/B AND2X1_LOC

XOR2X1_LOC_582 OR2X1_LOC_582/a_8_216# OR2X1_LOC_582/a_36_216# OR2X1_LOC_582/Y VSS VDD OR2X1_LOC_581/Y OR2X1_LOC_427/A OR2X1_LOC

XAND2X1_LOC_430 AND2X1_LOC_430/a_36_24# OR2X1_LOC_451/A AND2X1_LOC_430/a_8_24# VSS VDD OR2X1_LOC_161/A AND2X1_LOC_430/B AND2X1_LOC

XOR2X1_LOC_274 OR2X1_LOC_274/a_8_216# OR2X1_LOC_274/a_36_216# OR2X1_LOC_274/Y VSS VDD OR2X1_LOC_831/B OR2X1_LOC_541/A OR2X1_LOC

XAND2X1_LOC_599 AND2X1_LOC_599/a_36_24# OR2X1_LOC_644/A AND2X1_LOC_599/a_8_24# VSS VDD AND2X1_LOC_36/Y OR2X1_LOC_598/Y AND2X1_LOC

XAND2X1_LOC_274 AND2X1_LOC_274/a_36_24# OR2X1_LOC_275/A AND2X1_LOC_274/a_8_24# VSS VDD OR2X1_LOC_272/Y OR2X1_LOC_273/Y AND2X1_LOC

XOR2X1_LOC_599 OR2X1_LOC_599/a_8_216# OR2X1_LOC_599/a_36_216# OR2X1_LOC_599/Y VSS VDD OR2X1_LOC_599/A OR2X1_LOC_36/Y OR2X1_LOC

XAND2X1_LOC_411 AND2X1_LOC_411/a_36_24# OR2X1_LOC_461/B AND2X1_LOC_411/a_8_24# VSS VDD OR2X1_LOC_756/B OR2X1_LOC_410/Y AND2X1_LOC

XAND2X1_LOC_800 AND2X1_LOC_800/a_36_24# AND2X1_LOC_801/B AND2X1_LOC_800/a_8_24# VSS VDD AND2X1_LOC_687/Y OR2X1_LOC_760/Y AND2X1_LOC

XOR2X1_LOC_271 OR2X1_LOC_271/a_8_216# OR2X1_LOC_271/a_36_216# OR2X1_LOC_271/Y VSS VDD OR2X1_LOC_368/A OR2X1_LOC_271/B OR2X1_LOC

XAND2X1_LOC_88 AND2X1_LOC_88/a_36_24# AND2X1_LOC_88/Y AND2X1_LOC_88/a_8_24# VSS VDD AND2X1_LOC_3/Y OR2X1_LOC_87/Y AND2X1_LOC

XOR2X1_LOC_689 OR2X1_LOC_689/a_8_216# OR2X1_LOC_689/a_36_216# OR2X1_LOC_689/Y VSS VDD OR2X1_LOC_689/A OR2X1_LOC_31/Y OR2X1_LOC

XAND2X1_LOC_374 AND2X1_LOC_374/a_36_24# AND2X1_LOC_374/Y AND2X1_LOC_374/a_8_24# VSS VDD OR2X1_LOC_322/Y OR2X1_LOC_373/Y AND2X1_LOC

XAND2X1_LOC_327 AND2X1_LOC_327/a_36_24# OR2X1_LOC_329/B AND2X1_LOC_327/a_8_24# VSS VDD OR2X1_LOC_65/B OR2X1_LOC_517/A AND2X1_LOC

XOR2X1_LOC_66 OR2X1_LOC_66/a_8_216# OR2X1_LOC_66/a_36_216# OR2X1_LOC_66/Y VSS VDD OR2X1_LOC_66/A AND2X1_LOC_3/Y OR2X1_LOC

XOR2X1_LOC_120 OR2X1_LOC_120/a_8_216# OR2X1_LOC_120/a_36_216# OR2X1_LOC_121/A VSS VDD OR2X1_LOC_154/A AND2X1_LOC_41/A OR2X1_LOC

XOR2X1_LOC_820 OR2X1_LOC_820/a_8_216# OR2X1_LOC_820/a_36_216# OR2X1_LOC_820/Y VSS VDD OR2X1_LOC_820/A OR2X1_LOC_820/B OR2X1_LOC

XAND2X1_LOC_375 AND2X1_LOC_375/a_36_24# OR2X1_LOC_376/A AND2X1_LOC_375/a_8_24# VSS VDD OR2X1_LOC_31/Y OR2X1_LOC_158/A AND2X1_LOC

XAND2X1_LOC_530 AND2X1_LOC_530/a_36_24# OR2X1_LOC_548/A AND2X1_LOC_530/a_8_24# VSS VDD AND2X1_LOC_36/Y OR2X1_LOC_532/B AND2X1_LOC

XOR2X1_LOC_185 OR2X1_LOC_185/a_8_216# OR2X1_LOC_185/a_36_216# OR2X1_LOC_185/Y VSS VDD OR2X1_LOC_185/A AND2X1_LOC_56/B OR2X1_LOC

XOR2X1_LOC_800 OR2X1_LOC_800/a_8_216# OR2X1_LOC_800/a_36_216# OR2X1_LOC_800/Y VSS VDD OR2X1_LOC_800/A OR2X1_LOC_687/Y OR2X1_LOC

XAND2X1_LOC_271 AND2X1_LOC_271/a_36_24# OR2X1_LOC_276/B AND2X1_LOC_271/a_8_24# VSS VDD OR2X1_LOC_269/Y OR2X1_LOC_270/Y AND2X1_LOC

XOR2X1_LOC_88 OR2X1_LOC_88/a_8_216# OR2X1_LOC_88/a_36_216# OR2X1_LOC_88/Y VSS VDD OR2X1_LOC_88/A OR2X1_LOC_3/Y OR2X1_LOC

XOR2X1_LOC_411 OR2X1_LOC_411/a_8_216# OR2X1_LOC_411/a_36_216# OR2X1_LOC_411/Y VSS VDD OR2X1_LOC_411/A OR2X1_LOC_600/A OR2X1_LOC

XAND2X1_LOC_689 AND2X1_LOC_689/a_36_24# OR2X1_LOC_691/B AND2X1_LOC_689/a_8_24# VSS VDD AND2X1_LOC_31/Y OR2X1_LOC_688/Y AND2X1_LOC

XAND2X1_LOC_820 AND2X1_LOC_820/a_36_24# OR2X1_LOC_847/A AND2X1_LOC_820/a_8_24# VSS VDD OR2X1_LOC_818/Y AND2X1_LOC_820/B AND2X1_LOC

XOR2X1_LOC_327 OR2X1_LOC_327/a_8_216# OR2X1_LOC_327/a_36_216# OR2X1_LOC_405/A VSS VDD OR2X1_LOC_264/Y AND2X1_LOC_65/A OR2X1_LOC

XAND2X1_LOC_66 AND2X1_LOC_66/a_36_24# OR2X1_LOC_67/A AND2X1_LOC_66/a_8_24# VSS VDD OR2X1_LOC_3/Y OR2X1_LOC_26/Y AND2X1_LOC

XOR2X1_LOC_375 OR2X1_LOC_375/a_8_216# OR2X1_LOC_375/a_36_216# OR2X1_LOC_375/Y VSS VDD OR2X1_LOC_375/A AND2X1_LOC_31/Y OR2X1_LOC

XAND2X1_LOC_120 AND2X1_LOC_120/a_36_24# OR2X1_LOC_666/A AND2X1_LOC_120/a_8_24# VSS VDD OR2X1_LOC_13/B OR2X1_LOC_39/A AND2X1_LOC

XOR2X1_LOC_374 OR2X1_LOC_374/a_8_216# OR2X1_LOC_374/a_36_216# OR2X1_LOC_374/Y VSS VDD OR2X1_LOC_544/B OR2X1_LOC_325/B OR2X1_LOC

XOR2X1_LOC_530 OR2X1_LOC_530/a_8_216# OR2X1_LOC_530/a_36_216# OR2X1_LOC_530/Y VSS VDD OR2X1_LOC_485/A OR2X1_LOC_36/Y OR2X1_LOC

XAND2X1_LOC_185 AND2X1_LOC_185/a_36_24# OR2X1_LOC_816/A AND2X1_LOC_185/a_8_24# VSS VDD OR2X1_LOC_56/A OR2X1_LOC_74/A AND2X1_LOC

XOR2X1_LOC_410 OR2X1_LOC_410/a_8_216# OR2X1_LOC_410/a_36_216# OR2X1_LOC_410/Y VSS VDD AND2X1_LOC_51/Y AND2X1_LOC_12/Y OR2X1_LOC

XAND2X1_LOC_687 AND2X1_LOC_687/a_36_24# AND2X1_LOC_687/Y AND2X1_LOC_687/a_8_24# VSS VDD AND2X1_LOC_687/A AND2X1_LOC_687/B AND2X1_LOC

XOR2X1_LOC_760 OR2X1_LOC_760/a_8_216# OR2X1_LOC_760/a_36_216# OR2X1_LOC_760/Y VSS VDD OR2X1_LOC_329/B OR2X1_LOC_64/Y OR2X1_LOC

XAND2X1_LOC_270 AND2X1_LOC_270/a_36_24# OR2X1_LOC_368/A AND2X1_LOC_270/a_8_24# VSS VDD OR2X1_LOC_18/Y OR2X1_LOC_36/Y AND2X1_LOC

XAND2X1_LOC_269 AND2X1_LOC_269/a_36_24# OR2X1_LOC_271/B AND2X1_LOC_269/a_8_24# VSS VDD OR2X1_LOC_428/A OR2X1_LOC_268/Y AND2X1_LOC

XOR2X1_LOC_87 OR2X1_LOC_87/a_8_216# OR2X1_LOC_87/a_36_216# OR2X1_LOC_87/Y VSS VDD OR2X1_LOC_87/A OR2X1_LOC_87/B OR2X1_LOC

XOR2X1_LOC_373 OR2X1_LOC_373/a_8_216# OR2X1_LOC_373/a_36_216# OR2X1_LOC_373/Y VSS VDD OR2X1_LOC_89/A OR2X1_LOC_26/Y OR2X1_LOC

XAND2X1_LOC_264 AND2X1_LOC_264/a_36_24# OR2X1_LOC_517/A AND2X1_LOC_264/a_8_24# VSS VDD OR2X1_LOC_13/B OR2X1_LOC_89/A AND2X1_LOC

XAND2X1_LOC_760 AND2X1_LOC_760/a_36_24# OR2X1_LOC_800/A AND2X1_LOC_760/a_8_24# VSS VDD AND2X1_LOC_64/Y OR2X1_LOC_405/A AND2X1_LOC

XOR2X1_LOC_687 OR2X1_LOC_687/a_8_216# OR2X1_LOC_687/a_36_216# OR2X1_LOC_687/Y VSS VDD OR2X1_LOC_687/A OR2X1_LOC_687/B OR2X1_LOC

XOR2X1_LOC_269 OR2X1_LOC_269/a_8_216# OR2X1_LOC_269/a_36_216# OR2X1_LOC_269/Y VSS VDD OR2X1_LOC_269/A OR2X1_LOC_269/B OR2X1_LOC

XOR2X1_LOC_270 OR2X1_LOC_270/a_8_216# OR2X1_LOC_270/a_36_216# OR2X1_LOC_270/Y VSS VDD AND2X1_LOC_36/Y AND2X1_LOC_18/Y OR2X1_LOC

XAND2X1_LOC_87 AND2X1_LOC_87/a_36_24# OR2X1_LOC_88/A AND2X1_LOC_87/a_8_24# VSS VDD OR2X1_LOC_32/B OR2X1_LOC_52/B AND2X1_LOC

XAND2X1_LOC_410 AND2X1_LOC_410/a_36_24# OR2X1_LOC_411/A AND2X1_LOC_410/a_8_24# VSS VDD OR2X1_LOC_12/Y OR2X1_LOC_51/Y AND2X1_LOC

XOR2X1_LOC_264 OR2X1_LOC_264/a_8_216# OR2X1_LOC_264/a_36_216# OR2X1_LOC_264/Y VSS VDD OR2X1_LOC_78/A AND2X1_LOC_41/A OR2X1_LOC

XAND2X1_LOC_373 AND2X1_LOC_373/a_36_24# OR2X1_LOC_544/B AND2X1_LOC_373/a_8_24# VSS VDD OR2X1_LOC_66/A OR2X1_LOC_78/A AND2X1_LOC

XAND2X1_LOC_685 AND2X1_LOC_685/a_36_24# AND2X1_LOC_687/A AND2X1_LOC_685/a_8_24# VSS VDD OR2X1_LOC_681/Y OR2X1_LOC_682/Y AND2X1_LOC

XAND2X1_LOC_686 AND2X1_LOC_686/a_36_24# AND2X1_LOC_687/B AND2X1_LOC_686/a_8_24# VSS VDD OR2X1_LOC_683/Y OR2X1_LOC_684/Y AND2X1_LOC

XOR2X1_LOC_686 OR2X1_LOC_686/a_8_216# OR2X1_LOC_686/a_36_216# OR2X1_LOC_687/A VSS VDD OR2X1_LOC_686/A OR2X1_LOC_686/B OR2X1_LOC

XOR2X1_LOC_685 OR2X1_LOC_685/a_8_216# OR2X1_LOC_685/a_36_216# OR2X1_LOC_687/B VSS VDD OR2X1_LOC_685/A OR2X1_LOC_685/B OR2X1_LOC

XOR2X1_LOC_682 OR2X1_LOC_682/a_8_216# OR2X1_LOC_682/a_36_216# OR2X1_LOC_682/Y VSS VDD OR2X1_LOC_604/A OR2X1_LOC_36/Y OR2X1_LOC

XOR2X1_LOC_683 OR2X1_LOC_683/a_8_216# OR2X1_LOC_683/a_36_216# OR2X1_LOC_683/Y VSS VDD OR2X1_LOC_22/Y OR2X1_LOC_16/A OR2X1_LOC

XAND2X1_LOC_683 AND2X1_LOC_683/a_36_24# OR2X1_LOC_686/B AND2X1_LOC_683/a_8_24# VSS VDD OR2X1_LOC_78/B AND2X1_LOC_22/Y AND2X1_LOC

XAND2X1_LOC_682 AND2X1_LOC_682/a_36_24# OR2X1_LOC_685/A AND2X1_LOC_682/a_8_24# VSS VDD AND2X1_LOC_36/Y OR2X1_LOC_161/A AND2X1_LOC

C769 D_INPUT_7 VDD 0.36fF
C984 D_INPUT_7 AND2X1_LOC_25/a_8_24# 0.09fF
C3521 D_INPUT_7 AND2X1_LOC_1/Y 0.01fF
C5902 D_INPUT_7 AND2X1_LOC_50/a_8_24# 0.12fF
C7191 D_INPUT_7 AND2X1_LOC_12/a_8_24# 0.01fF
C8183 D_INPUT_7 AND2X1_LOC_21/Y 0.01fF
C8946 D_INPUT_7 AND2X1_LOC_51/a_8_24# 0.02fF
C11954 D_INPUT_7 AND2X1_LOC_17/Y 0.01fF
C12795 D_INPUT_7 AND2X1_LOC_11/Y 0.27fF
C14591 D_INPUT_7 AND2X1_LOC_11/a_8_24# 0.01fF
C15045 D_INPUT_7 OR2X1_LOC_51/B 0.05fF
C17454 D_INPUT_7 AND2X1_LOC_25/Y 0.01fF
C17508 D_INPUT_7 AND2X1_LOC_51/Y 0.09fF
C17926 D_INPUT_7 OR2X1_LOC_17/Y 0.01fF
C18536 D_INPUT_7 INPUT_6 0.61fF
C21624 D_INPUT_7 INPUT_7 0.85fF
C21773 D_INPUT_7 INPUT_4 0.29fF
C21799 D_INPUT_7 AND2X1_LOC_51/A 0.34fF
C22978 D_INPUT_7 AND2X1_LOC_2/Y 0.98fF
C24090 D_INPUT_7 D_INPUT_6 1.00fF
C27606 D_INPUT_7 OR2X1_LOC_2/Y 0.20fF
C28495 D_INPUT_7 AND2X1_LOC_1/a_8_24# 0.01fF
C28913 D_INPUT_7 AND2X1_LOC_17/a_8_24# 0.01fF
C29273 INPUT_5 D_INPUT_7 0.40fF
C29430 D_INPUT_7 OR2X1_LOC_17/a_8_216# 0.14fF
C33694 D_INPUT_7 OR2X1_LOC_2/a_8_216# 0.01fF
C34778 AND2X1_LOC_50/Y D_INPUT_7 0.01fF
C39851 D_INPUT_7 D_INPUT_5 0.08fF
C39891 AND2X1_LOC_12/Y D_INPUT_7 0.24fF
C39946 D_INPUT_7 AND2X1_LOC_21/a_8_24# 0.01fF
C41426 D_INPUT_7 AND2X1_LOC_587/a_8_24# 0.10fF
C43811 D_INPUT_7 AND2X1_LOC_30/a_8_24# 0.10fF
C46371 D_INPUT_7 D_INPUT_4 0.08fF
C55317 D_INPUT_7 AND2X1_LOC_2/a_8_24# 0.01fF
C57911 D_INPUT_7 VSS 0.12fF
C85 OR2X1_LOC_12/Y D_INPUT_6 0.41fF
C1058 OR2X1_LOC_30/a_8_216# D_INPUT_6 0.03fF
C2073 OR2X1_LOC_50/a_8_216# D_INPUT_6 0.01fF
C2326 D_INPUT_5 D_INPUT_6 1.12fF
C2443 AND2X1_LOC_21/a_8_24# D_INPUT_6 0.01fF
C2791 OR2X1_LOC_18/Y D_INPUT_6 1.63fF
C3943 AND2X1_LOC_587/a_8_24# D_INPUT_6 0.01fF
C4466 OR2X1_LOC_3/a_8_216# D_INPUT_6 0.01fF
C5711 OR2X1_LOC_429/Y D_INPUT_6 0.04fF
C6464 OR2X1_LOC_51/Y D_INPUT_6 0.90fF
C8730 D_INPUT_4 D_INPUT_6 1.24fF
C10491 OR2X1_LOC_762/a_36_216# D_INPUT_6 0.01fF
C10996 OR2X1_LOC_581/a_8_216# D_INPUT_6 0.07fF
C12095 OR2X1_LOC_30/a_36_216# D_INPUT_6 0.03fF
C18925 OR2X1_LOC_25/a_8_216# D_INPUT_6 0.01fF
C19284 VDD D_INPUT_6 0.24fF
C21946 OR2X1_LOC_44/Y D_INPUT_6 0.02fF
C21990 AND2X1_LOC_1/Y D_INPUT_6 0.01fF
C22742 OR2X1_LOC_158/A D_INPUT_6 0.37fF
C25391 OR2X1_LOC_31/Y D_INPUT_6 0.03fF
C26568 AND2X1_LOC_21/Y D_INPUT_6 0.07fF
C27189 OR2X1_LOC_11/a_8_216# D_INPUT_6 0.01fF
C27514 OR2X1_LOC_51/a_8_216# D_INPUT_6 0.01fF
C29015 OR2X1_LOC_12/a_8_216# D_INPUT_6 0.01fF
C29031 OR2X1_LOC_425/a_8_216# D_INPUT_6 0.01fF
C29870 OR2X1_LOC_638/B D_INPUT_6 0.08fF
C30374 AND2X1_LOC_17/Y D_INPUT_6 0.09fF
C31693 OR2X1_LOC_429/a_8_216# D_INPUT_6 0.01fF
C33446 OR2X1_LOC_51/B D_INPUT_6 0.01fF
C34916 OR2X1_LOC_428/A D_INPUT_6 0.07fF
C35884 AND2X1_LOC_51/Y D_INPUT_6 0.37fF
C36282 OR2X1_LOC_17/Y D_INPUT_6 1.09fF
C36905 D_INPUT_6 INPUT_6 0.72fF
C38091 OR2X1_LOC_70/A D_INPUT_6 1.10fF
C38492 OR2X1_LOC_47/Y D_INPUT_6 0.03fF
C38955 OR2X1_LOC_3/B D_INPUT_6 0.01fF
C39958 INPUT_7 D_INPUT_6 0.25fF
C40010 OR2X1_LOC_426/A D_INPUT_6 0.21fF
C40036 INPUT_4 D_INPUT_6 0.97fF
C40051 AND2X1_LOC_51/A D_INPUT_6 0.18fF
C41723 OR2X1_LOC_40/Y D_INPUT_6 0.04fF
C42699 OR2X1_LOC_22/a_8_216# D_INPUT_6 0.02fF
C43998 OR2X1_LOC_3/Y D_INPUT_6 0.08fF
C45262 OR2X1_LOC_11/Y D_INPUT_6 0.70fF
C45329 OR2X1_LOC_64/Y D_INPUT_6 0.11fF
C46113 OR2X1_LOC_2/Y D_INPUT_6 0.59fF
C46546 OR2X1_LOC_25/Y D_INPUT_6 0.01fF
C47065 AND2X1_LOC_1/a_8_24# D_INPUT_6 0.01fF
C47529 AND2X1_LOC_17/a_8_24# D_INPUT_6 0.01fF
C47902 INPUT_5 D_INPUT_6 0.08fF
C48085 OR2X1_LOC_17/a_8_216# D_INPUT_6 0.08fF
C52296 OR2X1_LOC_2/a_8_216# D_INPUT_6 0.01fF
C55525 OR2X1_LOC_157/a_8_216# D_INPUT_6 0.01fF
C55571 OR2X1_LOC_762/a_8_216# D_INPUT_6 0.05fF
C56330 D_INPUT_6 VSS 0.19fF
C1143 AND2X1_LOC_2/Y D_INPUT_5 0.03fF
C2264 D_INPUT_5 OR2X1_LOC_378/a_8_216# 0.02fF
C4129 D_INPUT_5 OR2X1_LOC_502/A 0.06fF
C4636 D_INPUT_5 AND2X1_LOC_3/Y 0.09fF
C5817 D_INPUT_5 OR2X1_LOC_2/Y 0.02fF
C6194 D_INPUT_5 OR2X1_LOC_25/Y 0.05fF
C6719 D_INPUT_5 AND2X1_LOC_1/a_8_24# 0.01fF
C7177 D_INPUT_5 AND2X1_LOC_17/a_8_24# 0.01fF
C7551 INPUT_5 D_INPUT_5 1.38fF
C7742 D_INPUT_5 OR2X1_LOC_17/a_8_216# 0.01fF
C8934 D_INPUT_5 OR2X1_LOC_752/a_8_216# 0.03fF
C9392 D_INPUT_5 OR2X1_LOC_378/Y 0.15fF
C9539 D_INPUT_5 OR2X1_LOC_378/A 0.30fF
C11713 D_INPUT_5 OR2X1_LOC_375/a_8_216# 0.01fF
C11999 D_INPUT_5 OR2X1_LOC_2/a_8_216# 0.01fF
C12313 D_INPUT_5 OR2X1_LOC_36/Y 0.03fF
C13131 AND2X1_LOC_50/Y D_INPUT_5 1.38fF
C13983 AND2X1_LOC_375/a_8_24# D_INPUT_5 0.02fF
C14222 D_INPUT_5 OR2X1_LOC_376/a_8_216# 0.01fF
C14422 D_INPUT_5 AND2X1_LOC_43/B 0.93fF
C16527 D_INPUT_5 AND2X1_LOC_64/a_8_24# 0.09fF
C16942 D_INPUT_5 OR2X1_LOC_30/a_8_216# 0.01fF
C17936 D_INPUT_5 OR2X1_LOC_50/a_8_216# 0.01fF
C18230 AND2X1_LOC_12/Y D_INPUT_5 0.01fF
C18317 D_INPUT_5 AND2X1_LOC_21/a_8_24# 0.19fF
C18624 AND2X1_LOC_752/a_8_24# D_INPUT_5 0.01fF
C19991 D_INPUT_5 OR2X1_LOC_753/A 0.01fF
C22094 OR2X1_LOC_377/A D_INPUT_5 0.06fF
C22547 D_INPUT_5 OR2X1_LOC_375/A 0.06fF
C24186 AND2X1_LOC_753/B D_INPUT_5 0.03fF
C24572 D_INPUT_5 D_INPUT_4 0.95fF
C25004 OR2X1_LOC_376/A D_INPUT_5 0.04fF
C28264 D_INPUT_5 OR2X1_LOC_375/Y 0.01fF
C29902 D_INPUT_5 AND2X1_LOC_409/B 0.03fF
C30696 D_INPUT_5 OR2X1_LOC_376/Y 0.01fF
C30737 OR2X1_LOC_696/A D_INPUT_5 0.25fF
C33412 D_INPUT_5 AND2X1_LOC_2/a_8_24# 0.05fF
C34671 D_INPUT_5 AND2X1_LOC_53/a_8_24# 0.10fF
C35051 VDD D_INPUT_5 0.13fF
C35230 D_INPUT_5 AND2X1_LOC_25/a_8_24# 0.01fF
C37735 D_INPUT_5 AND2X1_LOC_1/Y 0.01fF
C38375 OR2X1_LOC_158/A D_INPUT_5 0.03fF
C40121 AND2X1_LOC_50/a_8_24# D_INPUT_5 0.01fF
C40392 D_INPUT_5 AND2X1_LOC_429/a_8_24# 0.01fF
C41193 D_INPUT_5 OR2X1_LOC_31/Y 0.03fF
C41461 D_INPUT_5 AND2X1_LOC_12/a_8_24# 0.01fF
C42332 D_INPUT_5 AND2X1_LOC_3/a_8_24# 0.01fF
C42466 D_INPUT_5 AND2X1_LOC_21/Y 0.18fF
C46062 D_INPUT_5 AND2X1_LOC_430/B 0.01fF
C46355 AND2X1_LOC_17/Y D_INPUT_5 0.18fF
C47211 D_INPUT_5 AND2X1_LOC_11/Y 0.65fF
C47952 D_INPUT_5 AND2X1_LOC_44/Y 0.03fF
C49031 D_INPUT_5 AND2X1_LOC_11/a_8_24# 0.01fF
C49107 D_INPUT_5 OR2X1_LOC_377/a_8_216# 0.02fF
C49526 D_INPUT_5 OR2X1_LOC_51/B 0.01fF
C51901 D_INPUT_5 AND2X1_LOC_25/Y 0.01fF
C51955 D_INPUT_5 AND2X1_LOC_51/Y 0.03fF
C52370 D_INPUT_5 OR2X1_LOC_17/Y 0.40fF
C52978 D_INPUT_5 INPUT_6 0.06fF
C54154 D_INPUT_5 OR2X1_LOC_70/A 0.09fF
C54166 D_INPUT_5 AND2X1_LOC_31/Y 4.74fF
C55049 D_INPUT_5 AND2X1_LOC_36/Y 0.06fF
C55986 D_INPUT_5 INPUT_7 0.06fF
C56147 INPUT_4 D_INPUT_5 1.01fF
C56191 D_INPUT_5 AND2X1_LOC_51/A 0.19fF
C57531 D_INPUT_5 VSS 0.10fF
C2103 D_INPUT_4 AND2X1_LOC_25/Y 0.01fF
C2178 D_INPUT_4 AND2X1_LOC_51/Y 0.02fF
C2612 D_INPUT_4 OR2X1_LOC_17/Y 0.01fF
C3199 D_INPUT_4 INPUT_6 0.90fF
C4353 D_INPUT_4 AND2X1_LOC_31/Y 0.02fF
C5214 D_INPUT_4 AND2X1_LOC_36/Y 0.48fF
C6142 D_INPUT_4 INPUT_7 0.02fF
C6274 INPUT_4 D_INPUT_4 0.06fF
C6292 AND2X1_LOC_51/A D_INPUT_4 0.05fF
C7521 AND2X1_LOC_2/Y D_INPUT_4 0.04fF
C10553 OR2X1_LOC_502/A D_INPUT_4 0.11fF
C12261 D_INPUT_4 OR2X1_LOC_2/Y 0.09fF
C13190 D_INPUT_4 AND2X1_LOC_1/a_8_24# 0.02fF
C13220 AND2X1_LOC_386/a_8_24# D_INPUT_4 0.01fF
C13612 D_INPUT_4 AND2X1_LOC_17/a_8_24# 0.02fF
C13962 INPUT_5 D_INPUT_4 1.83fF
C14159 D_INPUT_4 OR2X1_LOC_17/a_8_216# 0.02fF
C15748 AND2X1_LOC_11/a_36_24# D_INPUT_4 0.01fF
C18400 D_INPUT_4 OR2X1_LOC_2/a_8_216# 0.02fF
C19468 AND2X1_LOC_50/Y D_INPUT_4 0.36fF
C20326 AND2X1_LOC_40/Y D_INPUT_4 0.07fF
C23375 D_INPUT_4 OR2X1_LOC_30/a_8_216# 0.07fF
C24274 AND2X1_LOC_387/B D_INPUT_4 0.01fF
C24710 AND2X1_LOC_21/a_8_24# D_INPUT_4 0.02fF
C25031 AND2X1_LOC_59/Y D_INPUT_4 0.08fF
C28432 AND2X1_LOC_30/a_8_24# D_INPUT_4 0.04fF
C33522 D_INPUT_4 OR2X1_LOC_21/a_8_216# 0.02fF
C38838 D_INPUT_4 OR2X1_LOC_596/A 0.01fF
C39025 D_INPUT_4 OR2X1_LOC_21/a_36_216# 0.03fF
C41420 VDD D_INPUT_4 0.53fF
C41644 D_INPUT_4 AND2X1_LOC_25/a_8_24# 0.01fF
C41926 D_INPUT_4 AND2X1_LOC_328/a_8_24# 0.10fF
C44210 AND2X1_LOC_1/Y D_INPUT_4 0.03fF
C46712 AND2X1_LOC_50/a_8_24# D_INPUT_4 0.02fF
C48988 D_INPUT_4 AND2X1_LOC_21/Y 0.01fF
C49745 AND2X1_LOC_51/a_8_24# D_INPUT_4 0.16fF
C50361 D_INPUT_4 AND2X1_LOC_47/Y 0.44fF
C52650 AND2X1_LOC_70/Y D_INPUT_4 0.02fF
C52774 AND2X1_LOC_17/Y D_INPUT_4 0.04fF
C53570 D_INPUT_4 AND2X1_LOC_11/Y 0.16fF
C54251 D_INPUT_4 AND2X1_LOC_44/Y 0.04fF
C55375 AND2X1_LOC_11/a_8_24# D_INPUT_4 0.04fF
C57301 D_INPUT_4 VSS -1.44fF
C87 AND2X1_LOC_55/a_8_24# D_INPUT_3 0.26fF
C1281 OR2X1_LOC_49/A D_INPUT_3 0.04fF
C1303 D_INPUT_3 OR2X1_LOC_381/a_36_216# 0.03fF
C1802 D_INPUT_3 AND2X1_LOC_820/a_8_24# 0.01fF
C2730 D_INPUT_3 AND2X1_LOC_42/B 0.03fF
C3880 VDD D_INPUT_3 1.12fF
C4350 D_INPUT_3 OR2X1_LOC_6/a_8_216# 0.01fF
C5123 D_INPUT_3 AND2X1_LOC_820/B 0.03fF
C5141 D_INPUT_3 OR2X1_LOC_427/A 0.02fF
C5743 D_INPUT_3 OR2X1_LOC_80/A 0.23fF
C6030 D_INPUT_3 OR2X1_LOC_6/A 0.08fF
C6108 D_INPUT_2 D_INPUT_3 0.28fF
C6771 D_INPUT_3 OR2X1_LOC_382/A 0.02fF
C7223 OR2X1_LOC_158/A D_INPUT_3 0.04fF
C7318 D_INPUT_3 OR2X1_LOC_847/A 0.54fF
C9508 OR2X1_LOC_529/a_8_216# D_INPUT_3 0.06fF
C9548 OR2X1_LOC_824/a_8_216# D_INPUT_3 0.01fF
C9611 D_INPUT_3 AND2X1_LOC_8/a_36_24# 0.01fF
C9874 OR2X1_LOC_744/A D_INPUT_3 0.09fF
C10722 D_INPUT_3 AND2X1_LOC_819/a_36_24# 0.01fF
C11106 D_INPUT_3 OR2X1_LOC_56/A 0.10fF
C11156 D_INPUT_3 AND2X1_LOC_9/a_8_24# 0.01fF
C11172 AND2X1_LOC_56/B D_INPUT_3 0.04fF
C11181 AND2X1_LOC_8/Y D_INPUT_3 0.02fF
C12033 D_INPUT_3 OR2X1_LOC_83/A 0.02fF
C12359 OR2X1_LOC_6/B D_INPUT_3 0.92fF
C12530 D_INPUT_3 AND2X1_LOC_47/Y 0.81fF
C12570 D_INPUT_3 OR2X1_LOC_598/A 0.02fF
C12979 D_INPUT_3 OR2X1_LOC_71/Y 0.17fF
C13004 D_INPUT_3 D_INPUT_1 0.04fF
C13270 OR2X1_LOC_426/B D_INPUT_3 0.07fF
C13404 D_INPUT_3 OR2X1_LOC_225/a_8_216# 0.01fF
C14533 OR2X1_LOC_235/B D_INPUT_3 0.01fF
C15294 OR2X1_LOC_9/Y D_INPUT_3 0.90fF
C16220 D_INPUT_3 OR2X1_LOC_92/Y 0.03fF
C16591 OR2X1_LOC_600/A D_INPUT_3 11.43fF
C17597 D_INPUT_3 AND2X1_LOC_672/a_8_24# 0.07fF
C18465 D_INPUT_3 OR2X1_LOC_62/B 0.03fF
C19013 D_INPUT_3 OR2X1_LOC_13/B 0.05fF
C19559 D_INPUT_3 OR2X1_LOC_428/A 0.03fF
C20183 D_INPUT_3 OR2X1_LOC_54/Y 0.16fF
C20568 D_INPUT_3 OR2X1_LOC_26/Y 0.08fF
C20578 D_INPUT_3 OR2X1_LOC_89/A 0.04fF
C21432 D_INPUT_3 OR2X1_LOC_824/Y 0.01fF
C21507 D_INPUT_3 OR2X1_LOC_95/Y 0.02fF
C22743 D_INPUT_3 OR2X1_LOC_820/B 0.02fF
C23226 D_INPUT_3 OR2X1_LOC_47/Y 0.08fF
C23533 OR2X1_LOC_625/Y D_INPUT_3 0.07fF
C25115 OR2X1_LOC_93/Y D_INPUT_3 0.01fF
C25670 D_INPUT_3 OR2X1_LOC_46/A 0.08fF
C25928 D_INPUT_3 INPUT_2 0.09fF
C26039 D_INPUT_3 OR2X1_LOC_93/a_8_216# 0.01fF
C26344 OR2X1_LOC_40/Y D_INPUT_3 0.03fF
C26447 D_INPUT_3 OR2X1_LOC_618/a_8_216# 0.01fF
C26466 D_INPUT_3 OR2X1_LOC_7/A 0.24fF
C27732 OR2X1_LOC_43/A D_INPUT_3 0.05fF
C28595 OR2X1_LOC_3/Y D_INPUT_3 0.91fF
C28639 D_INPUT_3 OR2X1_LOC_673/A 0.15fF
C28948 OR2X1_LOC_502/A D_INPUT_3 3.76fF
C29056 D_INPUT_3 OR2X1_LOC_618/Y 0.01fF
C29783 INPUT_0 D_INPUT_3 0.07fF
C29879 OR2X1_LOC_64/Y D_INPUT_3 0.03fF
C29905 D_INPUT_3 OR2X1_LOC_417/A 0.08fF
C31906 INPUT_3 D_INPUT_3 1.09fF
C32394 D_INPUT_3 AND2X1_LOC_28/a_8_24# 0.01fF
C32838 D_INPUT_3 INPUT_1 0.35fF
C33160 D_INPUT_3 OR2X1_LOC_517/A 0.03fF
C33631 AND2X1_LOC_62/a_8_24# D_INPUT_3 0.01fF
C33906 D_INPUT_3 OR2X1_LOC_415/Y 0.02fF
C34512 OR2X1_LOC_818/a_8_216# D_INPUT_3 0.08fF
C35264 D_INPUT_3 OR2X1_LOC_278/Y 0.03fF
C35336 D_INPUT_3 OR2X1_LOC_19/B 0.04fF
C37317 OR2X1_LOC_604/A D_INPUT_3 0.04fF
C38315 D_INPUT_3 D_INPUT_0 0.18fF
C38941 OR2X1_LOC_143/a_8_216# D_INPUT_3 0.01fF
C40035 D_INPUT_3 OR2X1_LOC_619/a_8_216# 0.01fF
C40687 D_INPUT_3 OR2X1_LOC_12/Y 0.23fF
C40759 AND2X1_LOC_54/a_8_24# D_INPUT_3 0.01fF
C42540 OR2X1_LOC_256/Y D_INPUT_3 0.03fF
C43889 D_INPUT_3 OR2X1_LOC_585/A 0.03fF
C44478 D_INPUT_3 OR2X1_LOC_437/A 0.07fF
C44734 D_INPUT_3 OR2X1_LOC_753/A 0.07fF
C45192 D_INPUT_3 OR2X1_LOC_37/a_8_216# 0.04fF
C45256 OR2X1_LOC_62/A D_INPUT_3 1.06fF
C45526 OR2X1_LOC_8/Y D_INPUT_3 0.24fF
C45600 D_INPUT_3 OR2X1_LOC_67/A 0.03fF
C45624 D_INPUT_3 OR2X1_LOC_672/Y 0.02fF
C46564 D_INPUT_3 AND2X1_LOC_672/B 0.54fF
C46920 D_INPUT_3 OR2X1_LOC_818/Y 0.01fF
C46947 D_INPUT_3 OR2X1_LOC_85/A 0.06fF
C47346 OR2X1_LOC_51/Y D_INPUT_3 0.03fF
C49193 D_INPUT_3 AND2X1_LOC_8/a_8_24# 0.07fF
C49535 D_INPUT_3 OR2X1_LOC_414/a_8_216# 0.07fF
C50345 OR2X1_LOC_91/A D_INPUT_3 0.13fF
C50953 D_INPUT_3 OR2X1_LOC_68/B 4.00fF
C51234 OR2X1_LOC_490/Y D_INPUT_3 0.04fF
C51235 D_INPUT_3 OR2X1_LOC_74/A 0.02fF
C51936 D_INPUT_3 OR2X1_LOC_381/a_8_216# 0.02fF
C53341 D_INPUT_3 AND2X1_LOC_37/a_8_24# 0.01fF
C55011 OR2X1_LOC_485/A D_INPUT_3 0.10fF
C55676 OR2X1_LOC_696/A D_INPUT_3 0.11fF
C55837 D_INPUT_3 AND2X1_LOC_819/a_8_24# 0.05fF
C57246 D_INPUT_3 VSS 0.73fF
C250 D_INPUT_2 OR2X1_LOC_80/A 0.16fF
C6784 OR2X1_LOC_6/B D_INPUT_2 0.05fF
C17210 D_INPUT_2 AND2X1_LOC_14/a_8_24# 0.02fF
C17988 D_INPUT_2 OR2X1_LOC_8/a_8_216# 0.03fF
C23460 OR2X1_LOC_671/a_8_216# D_INPUT_2 0.03fF
C23572 D_INPUT_2 OR2X1_LOC_8/a_36_216# 0.03fF
C24319 INPUT_0 D_INPUT_2 0.02fF
C26425 INPUT_3 D_INPUT_2 0.76fF
C26943 D_INPUT_2 AND2X1_LOC_28/a_8_24# 0.01fF
C27359 D_INPUT_2 INPUT_1 0.12fF
C32839 D_INPUT_2 D_INPUT_0 0.38fF
C34365 OR2X1_LOC_671/a_36_216# D_INPUT_2 0.03fF
C35241 AND2X1_LOC_54/a_8_24# D_INPUT_2 0.01fF
C39586 D_INPUT_2 OR2X1_LOC_37/a_8_216# 0.03fF
C39637 OR2X1_LOC_62/A D_INPUT_2 0.09fF
C39897 OR2X1_LOC_8/Y D_INPUT_2 0.01fF
C41231 OR2X1_LOC_377/A D_INPUT_2 0.10fF
C41243 D_INPUT_2 OR2X1_LOC_85/A 0.05fF
C45191 D_INPUT_2 OR2X1_LOC_37/a_36_216# 0.03fF
C54483 VDD D_INPUT_2 0.26fF
C57247 D_INPUT_2 VSS 0.50fF
C93 OR2X1_LOC_94/a_8_216# D_INPUT_1 0.01fF
C121 OR2X1_LOC_485/A D_INPUT_1 0.02fF
C418 OR2X1_LOC_633/A D_INPUT_1 0.04fF
C554 OR2X1_LOC_827/Y D_INPUT_1 0.04fF
C792 OR2X1_LOC_696/A D_INPUT_1 0.95fF
C808 AND2X1_LOC_64/Y D_INPUT_1 0.05fF
C854 AND2X1_LOC_82/Y D_INPUT_1 0.03fF
C890 AND2X1_LOC_86/a_8_24# D_INPUT_1 0.05fF
C1381 OR2X1_LOC_756/B D_INPUT_1 0.22fF
C2607 OR2X1_LOC_49/A D_INPUT_1 0.47fF
C2725 OR2X1_LOC_87/B D_INPUT_1 0.18fF
C2741 AND2X1_LOC_85/a_8_24# D_INPUT_1 0.02fF
C3050 OR2X1_LOC_671/Y D_INPUT_1 0.25fF
C3152 OR2X1_LOC_42/a_8_216# D_INPUT_1 0.07fF
C3212 OR2X1_LOC_532/B D_INPUT_1 0.11fF
C4007 AND2X1_LOC_42/B D_INPUT_1 0.67fF
C4354 OR2X1_LOC_185/Y D_INPUT_1 0.07fF
C4770 AND2X1_LOC_817/B D_INPUT_1 0.26fF
C5104 VDD D_INPUT_1 1.93fF
C6444 OR2X1_LOC_63/a_8_216# D_INPUT_1 0.01fF
C7075 D_INPUT_1 OR2X1_LOC_80/A 0.34fF
C7351 OR2X1_LOC_6/A D_INPUT_1 0.13fF
C8092 OR2X1_LOC_45/B D_INPUT_1 0.02fF
C8239 OR2X1_LOC_160/A D_INPUT_1 0.10fF
C8279 AND2X1_LOC_86/B D_INPUT_1 4.06fF
C8598 OR2X1_LOC_158/A D_INPUT_1 0.81fF
C8672 OR2X1_LOC_847/A D_INPUT_1 0.20fF
C8700 OR2X1_LOC_42/a_36_216# D_INPUT_1 0.03fF
C8723 AND2X1_LOC_46/a_8_24# D_INPUT_1 0.03fF
C9034 OR2X1_LOC_274/a_8_216# D_INPUT_1 0.04fF
C9521 OR2X1_LOC_185/A D_INPUT_1 0.07fF
C10418 OR2X1_LOC_293/a_8_216# D_INPUT_1 0.10fF
C11126 OR2X1_LOC_744/A D_INPUT_1 0.02fF
C11888 AND2X1_LOC_91/B D_INPUT_1 0.51fF
C12406 OR2X1_LOC_56/A D_INPUT_1 0.04fF
C12460 AND2X1_LOC_9/a_8_24# D_INPUT_1 0.07fF
C12471 AND2X1_LOC_56/B D_INPUT_1 0.03fF
C12478 AND2X1_LOC_8/Y D_INPUT_1 13.54fF
C12495 OR2X1_LOC_291/A D_INPUT_1 0.04fF
C12630 D_INPUT_1 AND2X1_LOC_236/a_8_24# 0.02fF
C13676 OR2X1_LOC_6/B D_INPUT_1 0.25fF
C13840 AND2X1_LOC_47/Y D_INPUT_1 12.92fF
C13891 D_INPUT_1 OR2X1_LOC_598/A 1.05fF
C14477 OR2X1_LOC_15/a_8_216# D_INPUT_1 0.01fF
C14529 OR2X1_LOC_426/B D_INPUT_1 0.21fF
C14589 AND2X1_LOC_95/Y D_INPUT_1 0.03fF
C15415 AND2X1_LOC_817/a_8_24# D_INPUT_1 0.07fF
C15432 AND2X1_LOC_490/a_8_24# D_INPUT_1 0.02fF
C15767 OR2X1_LOC_235/B D_INPUT_1 1.10fF
C15884 OR2X1_LOC_293/a_36_216# D_INPUT_1 0.03fF
C15916 OR2X1_LOC_276/B D_INPUT_1 0.07fF
C16197 AND2X1_LOC_70/Y D_INPUT_1 0.03fF
C16593 OR2X1_LOC_9/Y D_INPUT_1 0.71fF
C16691 OR2X1_LOC_96/B D_INPUT_1 0.33fF
C17523 OR2X1_LOC_65/B D_INPUT_1 0.01fF
C17586 OR2X1_LOC_62/a_8_216# D_INPUT_1 0.01fF
C17819 AND2X1_LOC_44/Y D_INPUT_1 0.15fF
C17885 OR2X1_LOC_600/A D_INPUT_1 0.06fF
C17958 OR2X1_LOC_619/Y D_INPUT_1 0.14fF
C18792 AND2X1_LOC_18/Y D_INPUT_1 5.02fF
C19182 AND2X1_LOC_606/a_8_24# D_INPUT_1 0.01fF
C19766 OR2X1_LOC_62/B D_INPUT_1 0.11fF
C20190 OR2X1_LOC_121/B D_INPUT_1 0.01fF
C21496 OR2X1_LOC_54/Y D_INPUT_1 0.34fF
C21845 OR2X1_LOC_161/A D_INPUT_1 0.13fF
C21941 OR2X1_LOC_92/a_8_216# D_INPUT_1 0.07fF
C22691 AND2X1_LOC_41/A D_INPUT_1 0.03fF
C23547 OR2X1_LOC_847/a_8_216# D_INPUT_1 0.02fF
C23566 AND2X1_LOC_102/a_8_24# D_INPUT_1 0.01fF
C23733 D_INPUT_1 OR2X1_LOC_71/A 0.26fF
C24125 AND2X1_LOC_31/Y D_INPUT_1 0.02fF
C24468 OR2X1_LOC_47/Y D_INPUT_1 0.07fF
C24658 D_INPUT_1 OR2X1_LOC_121/A 0.03fF
C24730 OR2X1_LOC_607/A D_INPUT_1 0.01fF
C24912 AND2X1_LOC_72/B D_INPUT_1 0.03fF
C25008 AND2X1_LOC_36/Y D_INPUT_1 8.61fF
C25513 OR2X1_LOC_16/A D_INPUT_1 0.19fF
C26468 OR2X1_LOC_847/B D_INPUT_1 0.01fF
C26485 OR2X1_LOC_557/A D_INPUT_1 0.03fF
C26947 OR2X1_LOC_46/A D_INPUT_1 0.18fF
C27253 INPUT_2 D_INPUT_1 0.10fF
C27334 OR2X1_LOC_269/B D_INPUT_1 3.89fF
C27647 OR2X1_LOC_40/Y D_INPUT_1 0.02fF
C27737 OR2X1_LOC_618/a_8_216# D_INPUT_1 0.01fF
C28437 OR2X1_LOC_831/B D_INPUT_1 0.06fF
C28871 OR2X1_LOC_161/B D_INPUT_1 0.07fF
C29003 OR2X1_LOC_43/A D_INPUT_1 0.12fF
C29873 OR2X1_LOC_3/Y D_INPUT_1 0.03fF
C29934 OR2X1_LOC_673/A D_INPUT_1 0.01fF
C30231 OR2X1_LOC_502/A D_INPUT_1 0.09fF
C30362 OR2X1_LOC_618/Y D_INPUT_1 0.01fF
C30557 OR2X1_LOC_489/A D_INPUT_1 0.04fF
C30661 AND2X1_LOC_104/a_8_24# D_INPUT_1 0.01fF
C30686 AND2X1_LOC_3/Y D_INPUT_1 0.06fF
C30804 D_INPUT_1 AND2X1_LOC_225/a_8_24# 0.03fF
C31072 INPUT_0 D_INPUT_1 0.25fF
C31395 AND2X1_LOC_7/B D_INPUT_1 0.07fF
C32805 OR2X1_LOC_287/B D_INPUT_1 0.06fF
C32910 OR2X1_LOC_28/a_8_216# D_INPUT_1 0.01fF
C33132 OR2X1_LOC_160/B D_INPUT_1 0.72fF
C33207 INPUT_3 D_INPUT_1 0.04fF
C33969 OR2X1_LOC_151/A D_INPUT_1 0.07fF
C34122 INPUT_1 D_INPUT_1 0.44fF
C34469 OR2X1_LOC_827/a_8_216# D_INPUT_1 0.01fF
C34913 AND2X1_LOC_62/a_8_24# D_INPUT_1 0.01fF
C35396 OR2X1_LOC_234/a_8_216# D_INPUT_1 0.01fF
C36465 AND2X1_LOC_90/a_8_24# D_INPUT_1 0.01fF
C36553 OR2X1_LOC_278/Y D_INPUT_1 0.02fF
C36611 OR2X1_LOC_19/B D_INPUT_1 0.17fF
C38268 AND2X1_LOC_382/a_8_24# D_INPUT_1 0.02fF
C38270 OR2X1_LOC_36/Y D_INPUT_1 0.05fF
C38637 OR2X1_LOC_66/A D_INPUT_1 0.10fF
C39633 D_INPUT_0 D_INPUT_1 0.18fF
C39942 AND2X1_LOC_40/Y D_INPUT_1 0.06fF
C39963 OR2X1_LOC_848/A D_INPUT_1 0.03fF
C40181 OR2X1_LOC_143/a_8_216# D_INPUT_1 0.12fF
C40855 OR2X1_LOC_119/a_8_216# D_INPUT_1 0.02fF
C42548 OR2X1_LOC_234/Y D_INPUT_1 -0.00fF
C42952 OR2X1_LOC_78/A D_INPUT_1 0.10fF
C43506 OR2X1_LOC_814/A D_INPUT_1 0.07fF
C44301 AND2X1_LOC_12/Y D_INPUT_1 0.11fF
C44718 OR2X1_LOC_18/Y D_INPUT_1 0.67fF
C44725 AND2X1_LOC_59/Y D_INPUT_1 0.03fF
C45198 OR2X1_LOC_585/A D_INPUT_1 0.06fF
C46076 OR2X1_LOC_753/A D_INPUT_1 0.03fF
C46565 OR2X1_LOC_119/a_36_216# D_INPUT_1 0.03fF
C46607 OR2X1_LOC_62/A D_INPUT_1 0.17fF
C46882 OR2X1_LOC_8/Y D_INPUT_1 0.13fF
C47318 OR2X1_LOC_9/a_8_216# D_INPUT_1 0.01fF
C47850 OR2X1_LOC_39/A D_INPUT_1 0.13fF
C47915 AND2X1_LOC_672/B D_INPUT_1 0.46fF
C48307 OR2X1_LOC_377/A D_INPUT_1 0.22fF
C48312 OR2X1_LOC_85/A D_INPUT_1 0.26fF
C48645 OR2X1_LOC_78/B D_INPUT_1 0.10fF
C48698 OR2X1_LOC_375/A D_INPUT_1 0.10fF
C49011 D_INPUT_1 OR2X1_LOC_549/A 0.14fF
C49573 OR2X1_LOC_391/B D_INPUT_1 0.82fF
C50405 OR2X1_LOC_405/A D_INPUT_1 0.01fF
C50488 AND2X1_LOC_8/a_8_24# D_INPUT_1 0.01fF
C51107 AND2X1_LOC_277/a_8_24# D_INPUT_1 0.01fF
C52078 OR2X1_LOC_233/a_8_216# D_INPUT_1 0.01fF
C52205 D_INPUT_1 OR2X1_LOC_68/B 1.05fF
C52522 OR2X1_LOC_74/A D_INPUT_1 0.05fF
C52937 OR2X1_LOC_87/A D_INPUT_1 0.04fF
C54100 OR2X1_LOC_541/A D_INPUT_1 0.03fF
C54948 OR2X1_LOC_778/B D_INPUT_1 0.16fF
C55447 OR2X1_LOC_154/A D_INPUT_1 0.87fF
C56411 D_INPUT_1 VSS 0.74fF
C90 D_INPUT_0 AND2X1_LOC_3/Y 0.54fF
C440 INPUT_0 D_INPUT_0 0.59fF
C514 D_INPUT_0 OR2X1_LOC_690/A 0.11fF
C548 OR2X1_LOC_64/Y D_INPUT_0 0.07fF
C567 D_INPUT_0 OR2X1_LOC_417/A 0.07fF
C771 D_INPUT_0 AND2X1_LOC_7/B 0.04fF
C955 OR2X1_LOC_836/A D_INPUT_0 0.01fF
C1892 OR2X1_LOC_473/A D_INPUT_0 0.15fF
C2603 OR2X1_LOC_160/B D_INPUT_0 0.14fF
C2677 AND2X1_LOC_86/Y D_INPUT_0 0.02fF
C2683 INPUT_3 D_INPUT_0 4.74fF
C3180 AND2X1_LOC_28/a_8_24# D_INPUT_0 0.04fF
C3417 OR2X1_LOC_151/A D_INPUT_0 0.27fF
C3596 INPUT_1 D_INPUT_0 1.88fF
C3900 OR2X1_LOC_517/A D_INPUT_0 0.22fF
C4299 AND2X1_LOC_62/a_8_24# D_INPUT_0 0.01fF
C5440 OR2X1_LOC_548/A D_INPUT_0 0.01fF
C5682 D_INPUT_0 OR2X1_LOC_66/a_8_216# 0.02fF
C6050 OR2X1_LOC_19/B D_INPUT_0 0.81fF
C6095 D_INPUT_0 OR2X1_LOC_838/B 0.03fF
C6305 AND2X1_LOC_110/Y D_INPUT_0 0.03fF
C6456 OR2X1_LOC_275/A D_INPUT_0 0.03fF
C6691 OR2X1_LOC_136/a_8_216# D_INPUT_0 0.01fF
C7384 D_INPUT_0 OR2X1_LOC_750/A 0.43fF
C7757 OR2X1_LOC_36/Y D_INPUT_0 0.37fF
C8106 D_INPUT_0 OR2X1_LOC_66/A 0.51fF
C8635 OR2X1_LOC_413/a_8_216# D_INPUT_0 0.06fF
C9459 AND2X1_LOC_40/Y D_INPUT_0 0.10fF
C9711 OR2X1_LOC_143/a_8_216# D_INPUT_0 0.01fF
C9910 D_INPUT_0 AND2X1_LOC_43/B 0.05fF
C10826 OR2X1_LOC_619/a_8_216# D_INPUT_0 0.01fF
C11458 D_INPUT_0 OR2X1_LOC_12/Y 2.67fF
C11537 AND2X1_LOC_54/a_8_24# D_INPUT_0 0.02fF
C11618 OR2X1_LOC_272/Y D_INPUT_0 0.03fF
C11701 D_INPUT_0 OR2X1_LOC_644/A 0.17fF
C11941 D_INPUT_0 OR2X1_LOC_234/Y 0.03fF
C12370 D_INPUT_0 OR2X1_LOC_78/A 0.16fF
C12458 D_INPUT_0 OR2X1_LOC_155/A 0.19fF
C12945 D_INPUT_0 OR2X1_LOC_814/A 0.16fF
C13344 AND2X1_LOC_387/B D_INPUT_0 2.06fF
C13605 OR2X1_LOC_121/Y D_INPUT_0 0.01fF
C13723 AND2X1_LOC_12/Y D_INPUT_0 0.35fF
C14140 D_INPUT_0 OR2X1_LOC_48/B 0.07fF
C14147 OR2X1_LOC_18/Y D_INPUT_0 1.81fF
C14154 AND2X1_LOC_59/Y D_INPUT_0 0.61fF
C14593 D_INPUT_0 OR2X1_LOC_585/A 0.11fF
C15147 D_INPUT_0 OR2X1_LOC_437/A 0.01fF
C15306 OR2X1_LOC_411/Y D_INPUT_0 0.12fF
C15388 D_INPUT_0 OR2X1_LOC_753/A 0.27fF
C15811 D_INPUT_0 OR2X1_LOC_37/a_8_216# 0.02fF
C15886 OR2X1_LOC_62/A D_INPUT_0 0.11fF
C15938 D_INPUT_0 OR2X1_LOC_88/Y 0.03fF
C16152 OR2X1_LOC_8/Y D_INPUT_0 0.26fF
C16255 D_INPUT_0 OR2X1_LOC_52/B 3.70fF
C16657 AND2X1_LOC_81/B D_INPUT_0 0.01fF
C16661 AND2X1_LOC_49/a_8_24# D_INPUT_0 0.03fF
C16712 OR2X1_LOC_22/Y D_INPUT_0 0.23fF
C16779 D_INPUT_0 OR2X1_LOC_66/Y 0.06fF
C17014 AND2X1_LOC_387/a_8_24# D_INPUT_0 0.01fF
C17088 D_INPUT_0 OR2X1_LOC_39/A 0.10fF
C17159 AND2X1_LOC_672/B D_INPUT_0 0.15fF
C17475 OR2X1_LOC_818/Y D_INPUT_0 0.02fF
C17494 OR2X1_LOC_377/A D_INPUT_0 0.39fF
C17514 D_INPUT_0 OR2X1_LOC_85/A 0.22fF
C17757 OR2X1_LOC_136/Y D_INPUT_0 0.07fF
C17846 OR2X1_LOC_51/Y D_INPUT_0 0.04fF
C17863 D_INPUT_0 OR2X1_LOC_78/B 0.54fF
C17933 D_INPUT_0 OR2X1_LOC_375/A 0.27fF
C18262 D_INPUT_0 OR2X1_LOC_549/A 0.26fF
C18921 D_INPUT_0 OR2X1_LOC_86/A 0.19fF
C19119 D_INPUT_0 AND2X1_LOC_65/A 0.09fF
C19656 OR2X1_LOC_405/A D_INPUT_0 0.05fF
C20181 D_INPUT_0 OR2X1_LOC_4/a_8_216# 0.01fF
C21428 OR2X1_LOC_233/a_8_216# D_INPUT_0 0.08fF
C21546 D_INPUT_0 OR2X1_LOC_68/B 0.33fF
C21854 D_INPUT_0 OR2X1_LOC_74/A 0.10fF
C22257 OR2X1_LOC_87/A D_INPUT_0 0.10fF
C22316 OR2X1_LOC_263/a_8_216# D_INPUT_0 0.06fF
C22610 OR2X1_LOC_389/A D_INPUT_0 0.01fF
C23088 OR2X1_LOC_71/a_8_216# D_INPUT_0 0.02fF
C23164 AND2X1_LOC_5/a_8_24# D_INPUT_0 0.02fF
C23565 OR2X1_LOC_415/A D_INPUT_0 0.01fF
C23811 OR2X1_LOC_691/Y D_INPUT_0 0.03fF
C23973 AND2X1_LOC_37/a_8_24# D_INPUT_0 0.01fF
C24377 OR2X1_LOC_278/a_8_216# D_INPUT_0 0.03fF
C24770 OR2X1_LOC_154/A D_INPUT_0 0.59fF
C24863 D_INPUT_0 AND2X1_LOC_6/a_8_24# 0.01fF
C25628 OR2X1_LOC_485/A D_INPUT_0 0.17fF
C25636 AND2X1_LOC_111/a_8_24# D_INPUT_0 0.02fF
C25869 D_INPUT_0 OR2X1_LOC_633/A 0.01fF
C25918 AND2X1_LOC_110/a_8_24# D_INPUT_0 0.04fF
C26239 OR2X1_LOC_696/A D_INPUT_0 0.94fF
C26253 AND2X1_LOC_64/Y D_INPUT_0 0.93fF
C26373 OR2X1_LOC_512/A D_INPUT_0 0.06fF
C26510 D_INPUT_0 OR2X1_LOC_54/a_8_216# 0.02fF
C26802 OR2X1_LOC_756/B D_INPUT_0 0.14fF
C27995 OR2X1_LOC_49/A D_INPUT_0 0.14fF
C28024 D_INPUT_0 OR2X1_LOC_596/A 0.02fF
C28525 AND2X1_LOC_820/a_8_24# D_INPUT_0 0.03fF
C28608 D_INPUT_0 OR2X1_LOC_532/B 0.54fF
C29415 AND2X1_LOC_42/B D_INPUT_0 0.20fF
C29820 OR2X1_LOC_185/Y D_INPUT_0 0.43fF
C29845 OR2X1_LOC_278/a_36_216# D_INPUT_0 0.01fF
C30552 VDD D_INPUT_0 0.94fF
C31847 D_INPUT_0 AND2X1_LOC_820/B 0.04fF
C31885 D_INPUT_0 OR2X1_LOC_63/a_8_216# 0.02fF
C31953 D_INPUT_0 OR2X1_LOC_54/a_36_216# 0.03fF
C32456 D_INPUT_0 OR2X1_LOC_80/A 0.89fF
C32764 D_INPUT_0 OR2X1_LOC_6/A 0.36fF
C33193 D_INPUT_0 OR2X1_LOC_44/Y 0.03fF
C33314 D_INPUT_0 OR2X1_LOC_750/Y 0.79fF
C33480 OR2X1_LOC_45/B D_INPUT_0 0.11fF
C33551 OR2X1_LOC_809/B D_INPUT_0 0.12fF
C33620 OR2X1_LOC_160/A D_INPUT_0 0.22fF
C33938 OR2X1_LOC_158/A D_INPUT_0 0.12fF
C34011 OR2X1_LOC_847/A D_INPUT_0 0.03fF
C34880 OR2X1_LOC_185/A D_INPUT_0 0.75fF
C35794 OR2X1_LOC_276/A D_INPUT_0 0.05fF
C36158 OR2X1_LOC_824/a_8_216# D_INPUT_0 0.01fF
C36482 OR2X1_LOC_744/A D_INPUT_0 0.03fF
C36604 OR2X1_LOC_31/Y D_INPUT_0 0.10fF
C37549 D_INPUT_0 OR2X1_LOC_446/B 0.05fF
C37736 D_INPUT_0 OR2X1_LOC_56/A 0.03fF
C37796 D_INPUT_0 AND2X1_LOC_9/a_8_24# 0.10fF
C37807 AND2X1_LOC_56/B D_INPUT_0 0.03fF
C37816 AND2X1_LOC_8/Y D_INPUT_0 1.53fF
C37840 OR2X1_LOC_291/A D_INPUT_0 0.02fF
C38158 D_INPUT_0 AND2X1_LOC_92/Y 6.40fF
C39021 OR2X1_LOC_6/B D_INPUT_0 2.28fF
C39193 AND2X1_LOC_47/Y D_INPUT_0 0.10fF
C39226 D_INPUT_0 OR2X1_LOC_598/A 7.74fF
C39611 OR2X1_LOC_71/Y D_INPUT_0 0.04fF
C39878 OR2X1_LOC_426/B D_INPUT_0 0.18fF
C39919 AND2X1_LOC_95/Y D_INPUT_0 0.11fF
C39962 OR2X1_LOC_743/A D_INPUT_0 0.07fF
C39982 OR2X1_LOC_415/a_8_216# D_INPUT_0 0.01fF
C39986 OR2X1_LOC_246/A D_INPUT_0 1.93fF
C40183 AND2X1_LOC_22/Y D_INPUT_0 0.16fF
C41166 OR2X1_LOC_235/B D_INPUT_0 0.11fF
C41307 OR2X1_LOC_276/B D_INPUT_0 0.48fF
C41368 D_INPUT_0 OR2X1_LOC_779/B 0.02fF
C41546 OR2X1_LOC_709/A D_INPUT_0 0.02fF
C41596 AND2X1_LOC_70/Y D_INPUT_0 0.23fF
C41992 OR2X1_LOC_9/Y D_INPUT_0 0.10fF
C42935 OR2X1_LOC_92/Y D_INPUT_0 0.03fF
C42973 D_INPUT_0 OR2X1_LOC_65/B 0.03fF
C43270 D_INPUT_0 AND2X1_LOC_44/Y 0.31fF
C43316 OR2X1_LOC_600/A D_INPUT_0 0.10fF
C43397 D_INPUT_0 OR2X1_LOC_619/Y 0.08fF
C44182 D_INPUT_0 AND2X1_LOC_18/Y 0.83fF
C44355 OR2X1_LOC_813/A D_INPUT_0 0.03fF
C44825 D_INPUT_0 OR2X1_LOC_512/a_8_216# 0.02fF
C45150 OR2X1_LOC_130/A D_INPUT_0 0.02fF
C45208 OR2X1_LOC_62/B D_INPUT_0 0.23fF
C45765 D_INPUT_0 OR2X1_LOC_13/B 13.90fF
C46796 D_INPUT_0 OR2X1_LOC_548/B 0.01fF
C46986 D_INPUT_0 OR2X1_LOC_54/Y 0.41fF
C47020 OR2X1_LOC_276/a_8_216# D_INPUT_0 0.03fF
C47389 D_INPUT_0 OR2X1_LOC_161/A 0.53fF
C47410 OR2X1_LOC_26/Y D_INPUT_0 0.35fF
C47418 D_INPUT_0 OR2X1_LOC_89/A 1.72fF
C47445 D_INPUT_0 AND2X1_LOC_51/Y 0.12fF
C47482 OR2X1_LOC_92/a_8_216# D_INPUT_0 0.03fF
C48218 AND2X1_LOC_41/A D_INPUT_0 0.19fF
C48281 D_INPUT_0 OR2X1_LOC_824/Y 0.34fF
C48306 OR2X1_LOC_688/a_8_216# D_INPUT_0 0.06fF
C48840 D_INPUT_0 OR2X1_LOC_112/A 0.01fF
C49233 D_INPUT_0 OR2X1_LOC_71/A 0.23fF
C49454 D_INPUT_0 OR2X1_LOC_59/Y 0.10fF
C49482 AND2X1_LOC_749/a_8_24# D_INPUT_0 0.05fF
C49567 OR2X1_LOC_70/Y D_INPUT_0 0.30fF
C49629 AND2X1_LOC_14/a_8_24# D_INPUT_0 0.02fF
C49667 D_INPUT_0 AND2X1_LOC_31/Y 0.59fF
C49972 D_INPUT_0 OR2X1_LOC_240/A 0.01fF
C50045 OR2X1_LOC_47/Y D_INPUT_0 2.28fF
C50426 D_INPUT_0 OR2X1_LOC_8/a_8_216# 0.06fF
C50478 D_INPUT_0 OR2X1_LOC_512/a_36_216# 0.03fF
C50567 D_INPUT_0 AND2X1_LOC_36/Y 0.95fF
C51068 D_INPUT_0 OR2X1_LOC_16/A 0.14fF
C52325 D_INPUT_0 OR2X1_LOC_548/a_8_216# 0.01fF
C52516 D_INPUT_0 OR2X1_LOC_46/A 0.43fF
C52794 D_INPUT_0 INPUT_2 0.06fF
C52906 D_INPUT_0 OR2X1_LOC_269/B 0.45fF
C53207 OR2X1_LOC_40/Y D_INPUT_0 0.13fF
C53269 AND2X1_LOC_690/a_8_24# D_INPUT_0 0.01fF
C53297 OR2X1_LOC_618/a_8_216# D_INPUT_0 0.01fF
C53320 D_INPUT_0 OR2X1_LOC_7/A 0.05fF
C53611 OR2X1_LOC_691/A D_INPUT_0 0.01fF
C53765 D_INPUT_0 OR2X1_LOC_86/a_8_216# 0.07fF
C54123 D_INPUT_0 AND2X1_LOC_824/a_8_24# 0.01fF
C54431 D_INPUT_0 OR2X1_LOC_161/B 0.02fF
C54444 OR2X1_LOC_589/A D_INPUT_0 0.02fF
C54564 OR2X1_LOC_43/A D_INPUT_0 13.82fF
C55322 D_INPUT_0 AND2X1_LOC_625/a_8_24# 0.01fF
C55442 OR2X1_LOC_3/Y D_INPUT_0 0.14fF
C55825 OR2X1_LOC_502/A D_INPUT_0 0.10fF
C55917 AND2X1_LOC_48/A D_INPUT_0 0.05fF
C55950 OR2X1_LOC_618/Y D_INPUT_0 0.40fF
C56171 AND2X1_LOC_530/a_8_24# D_INPUT_0 0.01fF
C57034 D_INPUT_0 VSS 0.77fF
C3331 OR2X1_LOC_429/Y INPUT_7 0.17fF
C11905 INPUT_7 OR2X1_LOC_587/a_8_216# 0.05fF
C16399 OR2X1_LOC_25/a_8_216# INPUT_7 0.08fF
C16762 VDD INPUT_7 0.23fF
C19477 AND2X1_LOC_1/Y INPUT_7 0.01fF
C24163 AND2X1_LOC_21/Y INPUT_7 0.01fF
C24739 OR2X1_LOC_11/a_8_216# INPUT_7 0.01fF
C29243 OR2X1_LOC_429/a_8_216# INPUT_7 0.03fF
C31008 OR2X1_LOC_51/B INPUT_7 0.18fF
C33850 OR2X1_LOC_17/Y INPUT_7 0.35fF
C34445 INPUT_7 INPUT_6 0.16fF
C35662 OR2X1_LOC_70/A INPUT_7 0.58fF
C37557 INPUT_4 INPUT_7 0.06fF
C40203 OR2X1_LOC_429/a_36_216# INPUT_7 0.01fF
C42740 OR2X1_LOC_11/Y INPUT_7 0.07fF
C43565 OR2X1_LOC_2/Y INPUT_7 0.07fF
C44461 AND2X1_LOC_1/a_8_24# INPUT_7 0.01fF
C44898 AND2X1_LOC_17/a_8_24# INPUT_7 0.11fF
C45285 INPUT_5 INPUT_7 0.70fF
C49871 OR2X1_LOC_2/a_8_216# INPUT_7 0.01fF
C54707 OR2X1_LOC_30/a_8_216# INPUT_7 0.01fF
C55775 OR2X1_LOC_50/a_8_216# INPUT_7 0.09fF
C56108 AND2X1_LOC_21/a_8_24# INPUT_7 0.01fF
C56497 INPUT_7 VSS 0.16fF
C627 AND2X1_LOC_30/a_8_24# INPUT_6 0.02fF
C1074 OR2X1_LOC_375/A INPUT_6 0.09fF
C3311 AND2X1_LOC_425/Y INPUT_6 0.03fF
C3951 AND2X1_LOC_588/B INPUT_6 -0.01fF
C7863 AND2X1_LOC_157/a_8_24# INPUT_6 0.01fF
C12078 AND2X1_LOC_2/a_8_24# INPUT_6 0.02fF
C13776 VDD INPUT_6 0.46fF
C13952 AND2X1_LOC_25/a_8_24# INPUT_6 0.04fF
C16385 AND2X1_LOC_1/Y INPUT_6 0.29fF
C18894 AND2X1_LOC_50/a_8_24# INPUT_6 0.02fF
C19788 OR2X1_LOC_1/a_8_216# INPUT_6 0.07fF
C20187 AND2X1_LOC_12/a_8_24# INPUT_6 0.01fF
C21023 AND2X1_LOC_3/a_8_24# INPUT_6 0.01fF
C21100 AND2X1_LOC_21/Y INPUT_6 1.02fF
C21897 AND2X1_LOC_51/a_8_24# INPUT_6 0.01fF
C22493 AND2X1_LOC_47/Y INPUT_6 0.03fF
C24456 AND2X1_LOC_157/a_36_24# INPUT_6 -0.00fF
C24660 AND2X1_LOC_430/B INPUT_6 0.03fF
C24903 AND2X1_LOC_17/Y INPUT_6 0.06fF
C25692 AND2X1_LOC_11/Y INPUT_6 0.84fF
C26442 AND2X1_LOC_44/Y INPUT_6 0.54fF
C26629 OR2X1_LOC_22/A INPUT_6 0.08fF
C27967 OR2X1_LOC_51/B INPUT_6 0.49fF
C30363 AND2X1_LOC_25/Y INPUT_6 0.03fF
C30416 AND2X1_LOC_51/Y INPUT_6 0.07fF
C30760 OR2X1_LOC_1/a_36_216# INPUT_6 0.03fF
C30825 OR2X1_LOC_17/Y INPUT_6 0.03fF
C32652 AND2X1_LOC_31/Y INPUT_6 0.04fF
C32942 AND2X1_LOC_31/a_8_24# INPUT_6 0.01fF
C33603 AND2X1_LOC_36/Y INPUT_6 0.03fF
C34546 INPUT_4 INPUT_6 0.04fF
C34568 AND2X1_LOC_51/A INPUT_6 0.03fF
C35761 AND2X1_LOC_2/Y INPUT_6 0.20fF
C38770 OR2X1_LOC_502/A INPUT_6 0.02fF
C39252 AND2X1_LOC_3/Y INPUT_6 0.01fF
C40061 AND2X1_LOC_44/a_8_24# INPUT_6 0.01fF
C40462 OR2X1_LOC_2/Y INPUT_6 0.01fF
C40532 AND2X1_LOC_425/a_8_24# INPUT_6 0.02fF
C41349 AND2X1_LOC_1/a_8_24# INPUT_6 0.04fF
C41815 AND2X1_LOC_17/a_8_24# INPUT_6 0.04fF
C42184 INPUT_5 INPUT_6 0.06fF
C42539 INPUT_6 AND2X1_LOC_581/a_8_24# 0.03fF
C43191 OR2X1_LOC_408/a_8_216# INPUT_6 0.02fF
C47909 AND2X1_LOC_50/Y INPUT_6 0.03fF
C52729 OR2X1_LOC_50/a_8_216# INPUT_6 0.07fF
C52998 AND2X1_LOC_12/Y INPUT_6 0.03fF
C54341 OR2X1_LOC_408/a_36_216# INPUT_6 0.03fF
C54559 AND2X1_LOC_587/a_8_24# INPUT_6 0.01fF
C55964 AND2X1_LOC_47/a_8_24# INPUT_6 0.04fF
C56264 INPUT_6 VSS 0.26fF
C1390 INPUT_5 OR2X1_LOC_2/a_8_216# 0.06fF
C1674 INPUT_5 OR2X1_LOC_36/Y 0.01fF
C2494 INPUT_5 AND2X1_LOC_50/Y 0.87fF
C3787 INPUT_5 AND2X1_LOC_43/B 0.02fF
C7670 INPUT_5 AND2X1_LOC_21/a_8_24# 0.09fF
C8004 INPUT_5 AND2X1_LOC_752/a_8_24# 0.10fF
C9164 INPUT_5 AND2X1_LOC_587/a_8_24# 0.01fF
C11048 INPUT_5 OR2X1_LOC_429/Y 0.02fF
C11455 INPUT_5 AND2X1_LOC_30/a_8_24# 0.01fF
C11775 INPUT_5 OR2X1_LOC_51/Y 0.05fF
C11857 INPUT_5 OR2X1_LOC_375/A 0.02fF
C12738 INPUT_5 OR2X1_LOC_588/Y 0.03fF
C14683 INPUT_5 AND2X1_LOC_588/B 0.01fF
C16545 INPUT_5 OR2X1_LOC_21/a_8_216# 0.18fF
C17626 INPUT_5 OR2X1_LOC_375/Y 0.09fF
C19329 INPUT_5 AND2X1_LOC_409/B 0.26fF
C19657 INPUT_5 OR2X1_LOC_587/a_8_216# 0.01fF
C20204 INPUT_5 OR2X1_LOC_696/A 0.20fF
C23367 INPUT_5 OR2X1_LOC_53/a_8_216# -0.00fF
C23428 INPUT_5 OR2X1_LOC_47/a_8_216# 0.09fF
C24510 INPUT_5 VDD 0.49fF
C24735 INPUT_5 AND2X1_LOC_25/a_8_24# 0.01fF
C27175 INPUT_5 OR2X1_LOC_44/Y 0.04fF
C27219 INPUT_5 AND2X1_LOC_1/Y 0.01fF
C27844 INPUT_5 OR2X1_LOC_158/A 0.03fF
C28854 INPUT_5 OR2X1_LOC_47/a_36_216# 0.02fF
C29595 INPUT_5 AND2X1_LOC_50/a_8_24# 0.01fF
C30485 INPUT_5 OR2X1_LOC_1/a_8_216# 0.01fF
C30613 INPUT_5 OR2X1_LOC_31/Y 0.42fF
C31792 INPUT_5 AND2X1_LOC_21/Y 0.01fF
C32543 INPUT_5 AND2X1_LOC_51/a_8_24# 0.01fF
C34007 INPUT_5 OR2X1_LOC_409/B 0.03fF
C34230 INPUT_5 OR2X1_LOC_425/a_8_216# 0.07fF
C35596 INPUT_5 AND2X1_LOC_17/Y 0.20fF
C37331 INPUT_5 OR2X1_LOC_22/A 0.05fF
C38180 INPUT_5 AND2X1_LOC_11/a_8_24# 0.11fF
C38674 INPUT_5 OR2X1_LOC_51/B 0.02fF
C41085 INPUT_5 AND2X1_LOC_25/Y 0.01fF
C41151 INPUT_5 AND2X1_LOC_51/Y 0.37fF
C41509 INPUT_5 OR2X1_LOC_1/a_36_216# -0.00fF
C41584 INPUT_5 OR2X1_LOC_17/Y 0.35fF
C41675 INPUT_5 OR2X1_LOC_588/A 0.01fF
C43421 INPUT_5 OR2X1_LOC_70/A 0.10fF
C43429 INPUT_5 AND2X1_LOC_31/Y 0.67fF
C44282 INPUT_5 OR2X1_LOC_3/B 0.77fF
C45431 INPUT_5 INPUT_4 0.29fF
C45460 INPUT_5 AND2X1_LOC_51/A 1.17fF
C46663 INPUT_5 AND2X1_LOC_2/Y 0.04fF
C47311 INPUT_5 OR2X1_LOC_44/a_8_216# 0.01fF
C49948 INPUT_5 OR2X1_LOC_31/a_8_216# 0.01fF
C50643 INPUT_5 OR2X1_LOC_11/Y 0.06fF
C51083 INPUT_5 AND2X1_LOC_44/a_8_24# 0.05fF
C51422 INPUT_5 OR2X1_LOC_2/Y 0.02fF
C51813 INPUT_5 OR2X1_LOC_25/Y 4.36fF
C52319 INPUT_5 AND2X1_LOC_1/a_8_24# 0.01fF
C52755 INPUT_5 AND2X1_LOC_17/a_8_24# 0.01fF
C53029 INPUT_5 OR2X1_LOC_36/a_8_216# 0.01fF
C54434 INPUT_5 OR2X1_LOC_752/a_8_216# 0.02fF
C58119 INPUT_5 VSS 0.22fF
C3466 INPUT_4 OR2X1_LOC_429/Y 0.01fF
C3865 INPUT_4 AND2X1_LOC_30/a_8_24# 0.10fF
C4133 INPUT_4 OR2X1_LOC_51/Y 0.06fF
C6121 INPUT_4 OR2X1_LOC_386/a_8_216# 0.07fF
C16027 INPUT_4 OR2X1_LOC_581/Y 0.01fF
C16572 INPUT_4 OR2X1_LOC_25/a_8_216# 0.01fF
C16905 VDD INPUT_4 0.04fF
C18260 INPUT_4 OR2X1_LOC_427/A 1.20fF
C20051 INPUT_4 OR2X1_LOC_430/a_8_216# 0.01fF
C20288 OR2X1_LOC_158/A INPUT_4 0.04fF
C23114 INPUT_4 OR2X1_LOC_31/Y 0.03fF
C24833 INPUT_4 OR2X1_LOC_11/a_8_216# 0.26fF
C27099 INPUT_4 OR2X1_LOC_582/a_8_216# 0.01fF
C28171 INPUT_4 OR2X1_LOC_430/Y 0.01fF
C31116 INPUT_4 OR2X1_LOC_51/B 0.10fF
C32476 INPUT_4 OR2X1_LOC_428/A 0.02fF
C33990 INPUT_4 OR2X1_LOC_17/Y 2.19fF
C35677 OR2X1_LOC_70/Y INPUT_4 0.01fF
C35756 INPUT_4 OR2X1_LOC_70/A 0.33fF
C36152 INPUT_4 OR2X1_LOC_47/Y 0.06fF
C41635 OR2X1_LOC_3/Y INPUT_4 0.06fF
C41663 INPUT_4 OR2X1_LOC_582/Y 0.01fF
C42877 INPUT_4 OR2X1_LOC_11/Y 0.05fF
C43726 INPUT_4 OR2X1_LOC_2/Y 1.11fF
C44098 INPUT_4 OR2X1_LOC_25/Y 0.04fF
C45612 INPUT_4 OR2X1_LOC_17/a_8_216# 0.01fF
C46754 OR2X1_LOC_328/a_8_216# INPUT_4 0.07fF
C49985 INPUT_4 OR2X1_LOC_2/a_8_216# 0.05fF
C53214 OR2X1_LOC_157/a_8_216# INPUT_4 0.01fF
C54844 INPUT_4 OR2X1_LOC_30/a_8_216# 0.01fF
C55894 INPUT_4 OR2X1_LOC_50/a_8_216# 0.01fF
C57597 INPUT_4 VSS 0.40fF
C1594 INPUT_3 OR2X1_LOC_66/A 0.50fF
C3220 OR2X1_LOC_143/a_8_216# INPUT_3 0.01fF
C4957 INPUT_3 AND2X1_LOC_54/a_8_24# 0.01fF
C7180 INPUT_3 AND2X1_LOC_12/Y 0.10fF
C9423 INPUT_3 OR2X1_LOC_37/a_8_216# 0.02fF
C9510 INPUT_3 OR2X1_LOC_62/A 0.53fF
C9696 INPUT_3 OR2X1_LOC_8/Y 0.05fF
C10719 INPUT_3 AND2X1_LOC_672/B 0.02fF
C11015 INPUT_3 OR2X1_LOC_377/A 0.01fF
C11042 INPUT_3 OR2X1_LOC_85/A 0.10fF
C13332 INPUT_3 AND2X1_LOC_8/a_8_24# 0.02fF
C13725 INPUT_3 OR2X1_LOC_4/a_8_216# 0.01fF
C14946 INPUT_3 OR2X1_LOC_5/a_8_216# 0.02fF
C15047 INPUT_3 OR2X1_LOC_68/B 3.84fF
C16642 INPUT_3 AND2X1_LOC_5/a_8_24# 0.11fF
C17431 INPUT_3 AND2X1_LOC_37/a_8_24# 0.14fF
C19803 OR2X1_LOC_696/A INPUT_3 0.01fF
C19929 INPUT_3 AND2X1_LOC_819/a_8_24# 0.03fF
C20416 INPUT_3 AND2X1_LOC_55/a_8_24# 0.03fF
C21560 OR2X1_LOC_49/A INPUT_3 0.41fF
C22004 INPUT_3 OR2X1_LOC_671/Y 0.09fF
C22114 INPUT_3 AND2X1_LOC_820/a_8_24# 0.06fF
C22240 INPUT_3 OR2X1_LOC_532/B 0.57fF
C23056 INPUT_3 AND2X1_LOC_42/B 0.34fF
C24153 INPUT_3 VDD 0.49fF
C25411 INPUT_3 AND2X1_LOC_820/B 0.05fF
C26077 INPUT_3 OR2X1_LOC_80/A 0.23fF
C26316 INPUT_3 OR2X1_LOC_6/A 0.21fF
C27553 INPUT_3 OR2X1_LOC_847/A 0.25fF
C28425 INPUT_3 OR2X1_LOC_185/A 0.03fF
C31399 INPUT_3 AND2X1_LOC_56/B 0.01fF
C31409 INPUT_3 AND2X1_LOC_8/Y 0.02fF
C32520 INPUT_3 OR2X1_LOC_6/B 0.27fF
C32564 INPUT_3 AND2X1_LOC_73/a_8_24# 0.03fF
C32752 INPUT_3 AND2X1_LOC_47/Y 0.09fF
C33046 INPUT_3 AND2X1_LOC_820/a_36_24# 0.01fF
C34675 INPUT_3 OR2X1_LOC_235/B 0.01fF
C35459 INPUT_3 OR2X1_LOC_9/Y 0.21fF
C36726 INPUT_3 OR2X1_LOC_600/A 0.03fF
C38651 INPUT_3 OR2X1_LOC_62/B 0.17fF
C40322 INPUT_3 OR2X1_LOC_54/Y 0.18fF
C42635 INPUT_3 OR2X1_LOC_71/A 0.01fF
C42996 INPUT_3 AND2X1_LOC_14/a_8_24# 0.01fF
C43798 INPUT_3 OR2X1_LOC_8/a_8_216# 0.03fF
C43959 INPUT_3 AND2X1_LOC_36/Y 0.07fF
C45997 INPUT_3 OR2X1_LOC_46/A 0.03fF
C46229 INPUT_3 INPUT_2 0.52fF
C46820 INPUT_3 OR2X1_LOC_618/a_8_216# 0.01fF
C49084 INPUT_3 OR2X1_LOC_673/A 0.10fF
C49370 INPUT_3 OR2X1_LOC_502/A 2.49fF
C50169 INPUT_3 INPUT_0 0.33fF
C52881 INPUT_3 AND2X1_LOC_28/a_8_24# 0.01fF
C53280 INPUT_3 INPUT_1 1.06fF
C53992 INPUT_3 AND2X1_LOC_62/a_8_24# 0.01fF
C55832 INPUT_3 OR2X1_LOC_19/B 0.36fF
C58021 INPUT_3 VSS 0.35fF
C2063 OR2X1_LOC_585/A INPUT_2 0.08fF
C2937 OR2X1_LOC_753/A INPUT_2 0.02fF
C3652 OR2X1_LOC_8/Y INPUT_2 1.74fF
C4628 AND2X1_LOC_672/B INPUT_2 0.01fF
C4938 OR2X1_LOC_85/A INPUT_2 0.02fF
C7255 AND2X1_LOC_8/a_8_24# INPUT_2 0.01fF
C8275 OR2X1_LOC_143/a_36_216# INPUT_2 0.03fF
C8927 OR2X1_LOC_5/a_8_216# INPUT_2 0.05fF
C11427 AND2X1_LOC_37/a_8_24# INPUT_2 0.09fF
C14449 OR2X1_LOC_5/a_36_216# INPUT_2 0.03fF
C15465 OR2X1_LOC_49/A INPUT_2 0.01fF
C15908 OR2X1_LOC_671/Y INPUT_2 0.02fF
C18070 VDD INPUT_2 0.23fF
C20244 OR2X1_LOC_104/a_8_216# INPUT_2 0.14fF
C20316 OR2X1_LOC_6/A INPUT_2 0.18fF
C25408 AND2X1_LOC_8/Y INPUT_2 0.01fF
C26549 OR2X1_LOC_6/B INPUT_2 0.29fF
C26774 AND2X1_LOC_47/Y INPUT_2 0.06fF
C28687 OR2X1_LOC_235/B INPUT_2 0.01fF
C29503 OR2X1_LOC_9/Y INPUT_2 0.02fF
C30775 OR2X1_LOC_600/A INPUT_2 0.10fF
C34305 OR2X1_LOC_54/Y INPUT_2 0.23fF
C42914 OR2X1_LOC_673/A INPUT_2 0.08fF
C43161 OR2X1_LOC_502/A INPUT_2 0.03fF
C43997 INPUT_0 INPUT_2 0.02fF
C45703 INPUT_2 OR2X1_LOC_14/a_8_216# 0.05fF
C47298 INPUT_1 INPUT_2 0.26fF
C55305 AND2X1_LOC_671/a_8_24# INPUT_2 0.10fF
C56646 INPUT_2 VSS 0.21fF
C536 OR2X1_LOC_273/Y INPUT_1 0.03fF
C550 OR2X1_LOC_19/B INPUT_1 0.08fF
C735 OR2X1_LOC_323/A INPUT_1 0.03fF
C1552 INPUT_1 OR2X1_LOC_300/a_8_216# 0.01fF
C2066 INPUT_1 OR2X1_LOC_748/Y 0.01fF
C2250 OR2X1_LOC_36/Y INPUT_1 0.22fF
C2595 OR2X1_LOC_604/A INPUT_1 0.09fF
C2608 INPUT_1 OR2X1_LOC_66/A 5.99fF
C2746 OR2X1_LOC_412/a_36_216# INPUT_1 0.02fF
C2800 INPUT_1 OR2X1_LOC_98/B 0.10fF
C3047 AND2X1_LOC_94/Y INPUT_1 0.17fF
C4313 INPUT_1 AND2X1_LOC_43/B 0.04fF
C5264 INPUT_1 OR2X1_LOC_749/a_8_216# 0.01fF
C5439 AND2X1_LOC_530/a_36_24# INPUT_1 0.01fF
C5887 INPUT_1 OR2X1_LOC_12/Y 0.17fF
C5958 AND2X1_LOC_54/a_8_24# INPUT_1 0.08fF
C8632 OR2X1_LOC_18/Y INPUT_1 0.21fF
C9065 INPUT_1 OR2X1_LOC_585/A 0.03fF
C9661 INPUT_1 OR2X1_LOC_437/A 0.39fF
C9928 INPUT_1 OR2X1_LOC_753/A 0.01fF
C10338 INPUT_1 OR2X1_LOC_37/a_8_216# 0.01fF
C10419 OR2X1_LOC_62/A INPUT_1 2.58fF
C10665 OR2X1_LOC_8/Y INPUT_1 1.48fF
C10769 INPUT_1 OR2X1_LOC_52/B 0.50fF
C11200 OR2X1_LOC_22/Y INPUT_1 3.08fF
C11475 OR2X1_LOC_820/a_8_216# INPUT_1 0.01fF
C11574 INPUT_1 OR2X1_LOC_39/A 0.06fF
C11643 AND2X1_LOC_672/B INPUT_1 0.10fF
C11970 INPUT_1 AND2X1_LOC_278/a_8_24# 0.17fF
C11975 OR2X1_LOC_377/A INPUT_1 0.27fF
C11987 INPUT_1 AND2X1_LOC_824/B 0.01fF
C12001 INPUT_1 OR2X1_LOC_85/A 1.41fF
C12355 OR2X1_LOC_51/Y INPUT_1 0.15fF
C12438 INPUT_1 OR2X1_LOC_375/A 0.58fF
C14237 AND2X1_LOC_28/a_36_24# INPUT_1 0.01fF
C14239 OR2X1_LOC_416/A INPUT_1 0.03fF
C14356 INPUT_1 OR2X1_LOC_268/Y 0.01fF
C15026 OR2X1_LOC_817/a_8_216# INPUT_1 0.05fF
C15314 OR2X1_LOC_91/A INPUT_1 0.15fF
C15776 OR2X1_LOC_32/B INPUT_1 0.24fF
C15817 INPUT_1 OR2X1_LOC_371/Y 0.38fF
C15939 INPUT_1 OR2X1_LOC_68/B 0.35fF
C16268 INPUT_1 OR2X1_LOC_74/A 0.09fF
C17048 AND2X1_LOC_54/a_36_24# INPUT_1 0.01fF
C17558 AND2X1_LOC_5/a_8_24# INPUT_1 0.01fF
C18129 INPUT_1 OR2X1_LOC_300/Y 0.54fF
C18381 INPUT_1 AND2X1_LOC_847/Y 0.03fF
C18415 AND2X1_LOC_37/a_8_24# INPUT_1 0.01fF
C20038 OR2X1_LOC_634/A INPUT_1 0.53fF
C20386 INPUT_1 OR2X1_LOC_633/A 0.09fF
C20562 OR2X1_LOC_827/Y INPUT_1 0.03fF
C20752 OR2X1_LOC_696/A INPUT_1 0.03fF
C20910 INPUT_1 AND2X1_LOC_819/a_8_24# 0.01fF
C20974 OR2X1_LOC_271/B INPUT_1 0.05fF
C21406 AND2X1_LOC_55/a_8_24# INPUT_1 0.03fF
C22557 OR2X1_LOC_49/A INPUT_1 0.14fF
C23004 OR2X1_LOC_671/Y INPUT_1 0.01fF
C23167 INPUT_1 OR2X1_LOC_532/B 1.02fF
C23972 AND2X1_LOC_42/B INPUT_1 0.32fF
C25088 VDD INPUT_1 0.98fF
C25382 INPUT_1 AND2X1_LOC_269/a_8_24# 0.02fF
C26203 INPUT_1 OR2X1_LOC_749/Y 0.13fF
C26364 INPUT_1 AND2X1_LOC_820/B 0.01fF
C26392 OR2X1_LOC_427/A INPUT_1 0.16fF
C26427 OR2X1_LOC_271/a_8_216# INPUT_1 0.02fF
C27001 INPUT_1 OR2X1_LOC_80/A 1.42fF
C27221 OR2X1_LOC_104/a_8_216# INPUT_1 0.01fF
C27295 INPUT_1 OR2X1_LOC_6/A 0.57fF
C27703 INPUT_1 OR2X1_LOC_44/Y 3.92fF
C27982 OR2X1_LOC_45/B INPUT_1 1.11fF
C28018 INPUT_1 OR2X1_LOC_382/A 0.05fF
C28441 OR2X1_LOC_158/A INPUT_1 0.30fF
C28524 OR2X1_LOC_847/A INPUT_1 0.02fF
C28975 OR2X1_LOC_748/A INPUT_1 0.06fF
C29231 AND2X1_LOC_92/a_8_24# INPUT_1 0.02fF
C29367 OR2X1_LOC_185/A INPUT_1 0.39fF
C29427 INPUT_1 AND2X1_LOC_119/a_8_24# 0.10fF
C30790 INPUT_1 OR2X1_LOC_153/a_8_216# 0.18fF
C31026 OR2X1_LOC_744/A INPUT_1 0.14fF
C31161 OR2X1_LOC_31/Y INPUT_1 0.42fF
C31584 INPUT_1 AND2X1_LOC_270/a_8_24# 0.01fF
C31955 INPUT_1 OR2X1_LOC_751/A 0.29fF
C32226 INPUT_1 OR2X1_LOC_56/A 0.21fF
C32230 OR2X1_LOC_819/a_8_216# INPUT_1 0.02fF
C32296 AND2X1_LOC_56/B INPUT_1 2.51fF
C32308 AND2X1_LOC_8/Y INPUT_1 0.04fF
C32689 INPUT_1 AND2X1_LOC_92/Y 0.01fF
C32773 INPUT_1 OR2X1_LOC_371/a_8_216# 0.03fF
C33200 OR2X1_LOC_83/A INPUT_1 0.03fF
C33518 OR2X1_LOC_6/B INPUT_1 0.44fF
C33703 AND2X1_LOC_47/Y INPUT_1 0.55fF
C33741 INPUT_1 OR2X1_LOC_598/A 0.10fF
C34341 OR2X1_LOC_426/B INPUT_1 0.07fF
C34409 AND2X1_LOC_95/Y INPUT_1 0.02fF
C34452 OR2X1_LOC_743/A INPUT_1 0.48fF
C34477 OR2X1_LOC_246/A INPUT_1 0.10fF
C34489 INPUT_1 OR2X1_LOC_225/a_8_216# 0.06fF
C35651 OR2X1_LOC_235/B INPUT_1 0.07fF
C36535 OR2X1_LOC_96/B INPUT_1 0.02fF
C36985 OR2X1_LOC_817/Y INPUT_1 0.01fF
C37349 OR2X1_LOC_92/Y INPUT_1 0.15fF
C37663 INPUT_1 AND2X1_LOC_44/Y 0.03fF
C37714 OR2X1_LOC_600/A INPUT_1 0.73fF
C37788 INPUT_1 OR2X1_LOC_619/Y 0.03fF
C38694 INPUT_1 AND2X1_LOC_234/a_8_24# 0.02fF
C38765 AND2X1_LOC_672/a_8_24# INPUT_1 0.03fF
C39605 OR2X1_LOC_62/B INPUT_1 0.03fF
C40094 INPUT_1 OR2X1_LOC_13/B 0.07fF
C40640 INPUT_1 OR2X1_LOC_428/A 0.60fF
C41279 INPUT_1 OR2X1_LOC_54/Y 0.25fF
C41688 OR2X1_LOC_26/Y INPUT_1 0.09fF
C41711 INPUT_1 OR2X1_LOC_820/Y 0.01fF
C42644 INPUT_1 OR2X1_LOC_95/Y 0.80fF
C42647 INPUT_1 OR2X1_LOC_368/A 0.01fF
C43064 INPUT_1 AND2X1_LOC_293/a_8_24# 0.03fF
C43352 OR2X1_LOC_820/A INPUT_1 0.12fF
C43582 INPUT_1 OR2X1_LOC_71/A 0.07fF
C43779 INPUT_1 OR2X1_LOC_59/Y 0.09fF
C43867 INPUT_1 OR2X1_LOC_820/B 0.42fF
C43887 OR2X1_LOC_70/Y INPUT_1 0.03fF
C43947 AND2X1_LOC_14/a_8_24# INPUT_1 0.01fF
C44295 INPUT_1 OR2X1_LOC_240/A 0.04fF
C44374 OR2X1_LOC_47/Y INPUT_1 0.25fF
C44744 INPUT_1 OR2X1_LOC_8/a_8_216# 0.01fF
C44909 INPUT_1 AND2X1_LOC_36/Y 0.12fF
C45445 INPUT_1 OR2X1_LOC_16/A 2.12fF
C45618 OR2X1_LOC_273/a_8_216# INPUT_1 0.03fF
C45819 OR2X1_LOC_110/a_8_216# INPUT_1 0.03fF
C46086 OR2X1_LOC_268/a_8_216# INPUT_1 0.03fF
C46795 INPUT_1 OR2X1_LOC_548/a_8_216# 0.06fF
C46984 INPUT_1 OR2X1_LOC_46/A 1.18fF
C47205 INPUT_1 OR2X1_LOC_748/a_8_216# 0.01fF
C47428 INPUT_1 AND2X1_LOC_847/a_8_24# 0.02fF
C47725 OR2X1_LOC_40/Y INPUT_1 0.06fF
C47846 INPUT_1 OR2X1_LOC_7/A 0.22fF
C48233 INPUT_1 OR2X1_LOC_46/a_8_216# 0.07fF
C48303 AND2X1_LOC_42/a_8_24# INPUT_1 0.06fF
C48969 OR2X1_LOC_589/A INPUT_1 0.02fF
C49040 INPUT_1 AND2X1_LOC_618/a_8_24# 0.14fF
C49083 OR2X1_LOC_43/A INPUT_1 0.17fF
C49981 OR2X1_LOC_3/Y INPUT_1 1.38fF
C50035 OR2X1_LOC_673/A INPUT_1 0.03fF
C50057 INPUT_1 AND2X1_LOC_462/B 0.09fF
C50277 OR2X1_LOC_671/a_8_216# INPUT_1 0.01fF
C50308 OR2X1_LOC_329/B INPUT_1 0.07fF
C50340 OR2X1_LOC_502/A INPUT_1 0.06fF
C50667 AND2X1_LOC_530/a_8_24# INPUT_1 0.03fF
C51124 INPUT_0 INPUT_1 7.14fF
C51211 INPUT_1 OR2X1_LOC_690/A 0.63fF
C51256 INPUT_1 OR2X1_LOC_417/A 0.45fF
C52519 INPUT_1 OR2X1_LOC_77/a_8_216# 0.05fF
C52916 OR2X1_LOC_287/B INPUT_1 0.14fF
C53361 OR2X1_LOC_412/a_8_216# INPUT_1 0.02fF
C53813 AND2X1_LOC_28/a_8_24# INPUT_1 0.09fF
C55253 INPUT_1 OR2X1_LOC_415/Y 0.05fF
C55508 AND2X1_LOC_672/a_36_24# INPUT_1 0.01fF
C56170 OR2X1_LOC_548/A INPUT_1 0.07fF
C57035 INPUT_1 VSS 0.98fF
C639 OR2X1_LOC_598/Y INPUT_0 0.03fF
C703 AND2X1_LOC_40/Y INPUT_0 0.07fF
C1213 INPUT_0 AND2X1_LOC_43/B 0.29fF
C2256 INPUT_0 OR2X1_LOC_749/a_8_216# 0.06fF
C2452 AND2X1_LOC_377/Y INPUT_0 0.06fF
C2810 INPUT_0 OR2X1_LOC_12/Y 0.02fF
C2880 INPUT_0 AND2X1_LOC_54/a_8_24# 0.14fF
C2939 INPUT_0 OR2X1_LOC_459/B 0.40fF
C3359 INPUT_0 OR2X1_LOC_828/B 0.07fF
C3699 INPUT_0 OR2X1_LOC_78/A 0.03fF
C3813 INPUT_0 OR2X1_LOC_155/A 0.02fF
C4613 AND2X1_LOC_387/B INPUT_0 0.07fF
C4956 AND2X1_LOC_12/Y INPUT_0 0.04fF
C5008 AND2X1_LOC_376/a_8_24# INPUT_0 0.01fF
C5355 INPUT_0 OR2X1_LOC_48/B 4.08fF
C5364 INPUT_0 OR2X1_LOC_18/Y 0.06fF
C5376 AND2X1_LOC_59/Y INPUT_0 0.07fF
C5878 INPUT_0 OR2X1_LOC_585/A 0.03fF
C6168 AND2X1_LOC_763/a_8_24# INPUT_0 0.04fF
C6460 INPUT_0 OR2X1_LOC_437/A 0.07fF
C6714 INPUT_0 OR2X1_LOC_753/A 0.08fF
C7276 INPUT_0 OR2X1_LOC_62/A 0.06fF
C7484 OR2X1_LOC_8/Y INPUT_0 0.02fF
C7611 INPUT_0 OR2X1_LOC_52/B 0.04fF
C7876 INPUT_0 OR2X1_LOC_9/a_8_216# 0.08fF
C7960 AND2X1_LOC_378/a_8_24# INPUT_0 0.01fF
C8112 INPUT_0 OR2X1_LOC_22/Y 1.46fF
C8471 INPUT_0 OR2X1_LOC_39/A 0.40fF
C8846 INPUT_0 OR2X1_LOC_818/Y 0.02fF
C8859 INPUT_0 AND2X1_LOC_278/a_8_24# 0.01fF
C8866 OR2X1_LOC_377/A INPUT_0 0.25fF
C8884 INPUT_0 AND2X1_LOC_824/B 0.04fF
C8900 INPUT_0 OR2X1_LOC_85/A 0.03fF
C9222 INPUT_0 OR2X1_LOC_51/Y 0.03fF
C9237 INPUT_0 OR2X1_LOC_78/B 0.08fF
C9297 AND2X1_LOC_94/a_8_24# INPUT_0 0.04fF
C9324 INPUT_0 OR2X1_LOC_375/A 0.12fF
C10741 INPUT_0 OR2X1_LOC_599/Y 0.11fF
C11767 OR2X1_LOC_769/B INPUT_0 0.03fF
C12183 INPUT_0 OR2X1_LOC_91/A 0.13fF
C12551 INPUT_0 OR2X1_LOC_138/A 0.04fF
C12745 INPUT_0 AND2X1_LOC_4/a_8_24# 0.04fF
C12771 INPUT_0 OR2X1_LOC_5/a_8_216# 0.01fF
C12899 INPUT_0 OR2X1_LOC_68/B 1.35fF
C13204 INPUT_0 OR2X1_LOC_74/A 0.01fF
C13492 OR2X1_LOC_459/A INPUT_0 0.34fF
C14473 INPUT_0 OR2X1_LOC_275/a_8_216# 0.02fF
C14900 INPUT_0 OR2X1_LOC_415/A 0.01fF
C15096 OR2X1_LOC_43/Y INPUT_0 0.01fF
C15142 INPUT_0 OR2X1_LOC_690/Y 0.01fF
C15532 INPUT_0 OR2X1_LOC_461/B 0.13fF
C16070 OR2X1_LOC_154/A INPUT_0 0.35fF
C16745 INPUT_0 AND2X1_LOC_763/B 0.02fF
C16830 OR2X1_LOC_461/a_8_216# INPUT_0 0.01fF
C16862 INPUT_0 OR2X1_LOC_634/A 0.09fF
C16936 INPUT_0 OR2X1_LOC_94/a_8_216# 0.01fF
C16987 OR2X1_LOC_485/A INPUT_0 1.06fF
C17217 INPUT_0 OR2X1_LOC_633/A 0.58fF
C17379 INPUT_0 OR2X1_LOC_827/Y 0.01fF
C17572 OR2X1_LOC_696/A INPUT_0 0.11fF
C17581 AND2X1_LOC_64/Y INPUT_0 0.16fF
C17636 AND2X1_LOC_86/a_8_24# INPUT_0 0.03fF
C18217 INPUT_0 AND2X1_LOC_55/a_8_24# 0.02fF
C18737 INPUT_0 OR2X1_LOC_43/a_8_216# 0.01fF
C18830 INPUT_0 AND2X1_LOC_699/a_8_24# 0.02fF
C19087 INPUT_0 OR2X1_LOC_82/a_8_216# 0.03fF
C19362 OR2X1_LOC_49/A INPUT_0 0.22fF
C19378 INPUT_0 OR2X1_LOC_596/A 0.03fF
C19814 OR2X1_LOC_671/Y INPUT_0 0.05fF
C19862 INPUT_0 AND2X1_LOC_529/a_8_24# 0.02fF
C19913 INPUT_0 AND2X1_LOC_820/a_8_24# 0.01fF
C19958 INPUT_0 OR2X1_LOC_42/a_8_216# 0.01fF
C20037 INPUT_0 OR2X1_LOC_532/B 2.01fF
C20694 INPUT_0 AND2X1_LOC_691/a_8_24# 0.01fF
C20838 INPUT_0 AND2X1_LOC_42/B 0.08fF
C21226 OR2X1_LOC_185/Y INPUT_0 0.07fF
C21970 VDD INPUT_0 0.83fF
C22036 INPUT_0 OR2X1_LOC_689/A 0.03fF
C23321 INPUT_0 OR2X1_LOC_427/A 0.03fF
C23970 INPUT_0 OR2X1_LOC_80/A 0.35fF
C24215 INPUT_0 OR2X1_LOC_6/A 1.54fF
C24610 INPUT_0 OR2X1_LOC_44/Y 0.18fF
C24616 INPUT_0 OR2X1_LOC_82/a_36_216# 0.02fF
C24875 OR2X1_LOC_45/B INPUT_0 0.05fF
C24992 OR2X1_LOC_160/A INPUT_0 0.36fF
C25052 AND2X1_LOC_86/B INPUT_0 0.02fF
C25316 OR2X1_LOC_158/A INPUT_0 0.33fF
C25396 INPUT_0 OR2X1_LOC_847/A 0.04fF
C25505 INPUT_0 OR2X1_LOC_275/a_36_216# 0.03fF
C25815 AND2X1_LOC_94/a_36_24# INPUT_0 0.01fF
C26242 OR2X1_LOC_185/A INPUT_0 0.17fF
C26804 INPUT_0 OR2X1_LOC_111/Y 0.03fF
C28092 INPUT_0 OR2X1_LOC_31/Y 2.10fF
C29128 INPUT_0 OR2X1_LOC_56/A 0.09fF
C29223 INPUT_0 AND2X1_LOC_56/B 13.29fF
C29239 INPUT_0 AND2X1_LOC_8/Y 0.08fF
C30096 INPUT_0 OR2X1_LOC_83/A 0.05fF
C30375 INPUT_0 OR2X1_LOC_596/a_8_216# 0.01fF
C30379 OR2X1_LOC_6/B INPUT_0 0.17fF
C30411 AND2X1_LOC_73/a_8_24# INPUT_0 0.02fF
C30596 INPUT_0 AND2X1_LOC_47/Y 0.06fF
C30641 INPUT_0 OR2X1_LOC_598/A 0.11fF
C31248 OR2X1_LOC_426/B INPUT_0 0.10fF
C31304 INPUT_0 AND2X1_LOC_414/a_8_24# 0.02fF
C31319 AND2X1_LOC_95/Y INPUT_0 0.17fF
C31377 INPUT_0 OR2X1_LOC_743/A 0.04fF
C31609 AND2X1_LOC_22/Y INPUT_0 0.07fF
C32496 OR2X1_LOC_235/B INPUT_0 0.07fF
C32886 INPUT_0 OR2X1_LOC_57/a_8_216# 0.05fF
C32915 AND2X1_LOC_70/Y INPUT_0 0.07fF
C33311 OR2X1_LOC_9/Y INPUT_0 0.03fF
C33448 INPUT_0 OR2X1_LOC_96/B 0.03fF
C33824 INPUT_0 OR2X1_LOC_637/B 0.01fF
C34535 INPUT_0 AND2X1_LOC_44/Y 0.09fF
C34578 INPUT_0 OR2X1_LOC_600/A 0.07fF
C34667 INPUT_0 OR2X1_LOC_619/Y 0.07fF
C35130 OR2X1_LOC_690/a_8_216# INPUT_0 0.08fF
C35420 INPUT_0 AND2X1_LOC_18/Y 0.07fF
C35555 OR2X1_LOC_596/Y INPUT_0 0.03fF
C35558 INPUT_0 AND2X1_LOC_413/a_8_24# 0.01fF
C35682 INPUT_0 AND2X1_LOC_672/a_8_24# 0.03fF
C36400 INPUT_0 AND2X1_LOC_688/a_8_24# 0.01fF
C36474 INPUT_0 OR2X1_LOC_62/B 0.04fF
C37002 INPUT_0 OR2X1_LOC_13/B 0.50fF
C37504 INPUT_0 OR2X1_LOC_428/A 0.10fF
C37914 INPUT_0 OR2X1_LOC_548/B 0.01fF
C37989 AND2X1_LOC_512/Y INPUT_0 0.01fF
C38144 INPUT_0 OR2X1_LOC_54/Y 4.71fF
C38358 INPUT_0 OR2X1_LOC_57/a_36_216# 0.03fF
C38460 INPUT_0 OR2X1_LOC_689/a_8_216# 0.01fF
C38512 INPUT_0 OR2X1_LOC_26/Y 0.50fF
C38555 OR2X1_LOC_461/Y INPUT_0 0.01fF
C38563 INPUT_0 AND2X1_LOC_51/Y 0.02fF
C38927 OR2X1_LOC_306/a_8_216# INPUT_0 0.01fF
C39300 INPUT_0 AND2X1_LOC_41/A 0.10fF
C39500 INPUT_0 OR2X1_LOC_95/Y 0.02fF
C39846 INPUT_0 AND2X1_LOC_136/a_8_24# 0.04fF
C40401 INPUT_0 OR2X1_LOC_71/A 0.19fF
C40546 INPUT_0 OR2X1_LOC_59/Y 0.03fF
C40677 OR2X1_LOC_70/Y INPUT_0 0.02fF
C40704 AND2X1_LOC_514/Y INPUT_0 0.03fF
C40791 INPUT_0 AND2X1_LOC_31/Y 0.07fF
C41070 INPUT_0 OR2X1_LOC_461/A 0.15fF
C41194 INPUT_0 OR2X1_LOC_47/Y 0.02fF
C41414 AND2X1_LOC_73/a_36_24# INPUT_0 0.01fF
C41747 INPUT_0 AND2X1_LOC_36/Y 5.83fF
C42224 INPUT_0 OR2X1_LOC_16/A 0.03fF
C42755 INPUT_0 AND2X1_LOC_126/a_8_24# 0.02fF
C43307 INPUT_0 AND2X1_LOC_729/B 0.04fF
C43772 INPUT_0 OR2X1_LOC_46/A 1.42fF
C44128 INPUT_0 OR2X1_LOC_269/B 0.07fF
C44413 OR2X1_LOC_40/Y INPUT_0 0.15fF
C44577 INPUT_0 OR2X1_LOC_7/A 0.03fF
C45699 INPUT_0 OR2X1_LOC_161/B 0.47fF
C45711 OR2X1_LOC_589/A INPUT_0 0.03fF
C45853 INPUT_0 OR2X1_LOC_43/A 0.63fF
C46809 OR2X1_LOC_3/Y INPUT_0 0.10fF
C46891 INPUT_0 OR2X1_LOC_673/A 0.03fF
C46949 INPUT_0 AND2X1_LOC_409/a_8_24# 0.01fF
C47153 OR2X1_LOC_502/A INPUT_0 1.47fF
C47321 INPUT_0 AND2X1_LOC_48/A 0.09fF
C47524 AND2X1_LOC_530/a_8_24# INPUT_0 0.03fF
C47694 INPUT_0 AND2X1_LOC_3/Y 0.23fF
C48126 INPUT_0 OR2X1_LOC_690/A 0.82fF
C48182 INPUT_0 OR2X1_LOC_64/Y 0.07fF
C48217 INPUT_0 OR2X1_LOC_417/A 0.07fF
C48371 INPUT_0 AND2X1_LOC_7/B 0.45fF
C48516 INPUT_0 OR2X1_LOC_407/a_8_216# 0.03fF
C49678 INPUT_0 OR2X1_LOC_14/a_8_216# 0.01fF
C49818 AND2X1_LOC_512/a_8_24# INPUT_0 0.03fF
C49821 OR2X1_LOC_287/B INPUT_0 0.16fF
C49946 INPUT_0 OR2X1_LOC_28/a_8_216# 0.01fF
C50089 OR2X1_LOC_160/B INPUT_0 0.07fF
C50602 INPUT_0 AND2X1_LOC_233/a_8_24# 0.01fF
C50745 INPUT_0 AND2X1_LOC_28/a_8_24# 0.03fF
C50893 OR2X1_LOC_53/Y INPUT_0 0.02fF
C51404 INPUT_0 AND2X1_LOC_619/B 0.10fF
C51463 INPUT_0 OR2X1_LOC_827/a_8_216# 0.01fF
C52109 INPUT_0 OR2X1_LOC_415/Y 0.03fF
C52485 INPUT_0 OR2X1_LOC_460/A 0.01fF
C52828 INPUT_0 OR2X1_LOC_818/a_8_216# 0.01fF
C53673 INPUT_0 OR2X1_LOC_19/B 0.20fF
C54927 INPUT_0 OR2X1_LOC_689/Y 0.02fF
C55261 INPUT_0 OR2X1_LOC_36/Y 6.37fF
C55559 INPUT_0 OR2X1_LOC_66/A 0.11fF
C55658 OR2X1_LOC_306/Y INPUT_0 0.07fF
C56025 AND2X1_LOC_94/Y INPUT_0 0.53fF
C57468 INPUT_0 VSS -4.74fF
C1039 AND2X1_LOC_7/B OR2X1_LOC_515/A 0.03fF
C7337 OR2X1_LOC_515/A OR2X1_LOC_515/a_8_216# 0.39fF
C10101 AND2X1_LOC_43/B OR2X1_LOC_515/A 0.01fF
C12681 OR2X1_LOC_155/A OR2X1_LOC_515/A 0.03fF
C24964 OR2X1_LOC_154/A OR2X1_LOC_515/A 0.01fF
C28232 OR2X1_LOC_596/A OR2X1_LOC_515/A 0.02fF
C30766 VDD OR2X1_LOC_515/A -0.00fF
C37810 OR2X1_LOC_446/B OR2X1_LOC_515/A 0.06fF
C38012 AND2X1_LOC_56/B OR2X1_LOC_515/A 0.02fF
C41763 OR2X1_LOC_709/A OR2X1_LOC_515/A 0.01fF
C43508 OR2X1_LOC_514/a_8_216# OR2X1_LOC_515/A -0.00fF
C50832 AND2X1_LOC_36/Y OR2X1_LOC_515/A 0.01fF
C56316 OR2X1_LOC_515/A VSS 0.18fF
C3882 OR2X1_LOC_749/Y AND2X1_LOC_750/a_8_24# 0.01fF
C4121 OR2X1_LOC_751/A OR2X1_LOC_749/Y 0.01fF
C4373 OR2X1_LOC_819/a_8_216# OR2X1_LOC_749/Y 0.40fF
C5608 OR2X1_LOC_6/B OR2X1_LOC_749/Y 0.01fF
C9948 OR2X1_LOC_600/A OR2X1_LOC_749/Y 0.46fF
C14774 OR2X1_LOC_95/Y OR2X1_LOC_749/Y 0.01fF
C15441 OR2X1_LOC_820/A OR2X1_LOC_749/Y 0.01fF
C16464 OR2X1_LOC_47/Y OR2X1_LOC_749/Y 0.04fF
C38471 OR2X1_LOC_62/A OR2X1_LOC_749/Y 0.09fF
C53336 VDD OR2X1_LOC_749/Y 0.08fF
C55969 OR2X1_LOC_44/Y OR2X1_LOC_749/Y 0.01fF
C56315 OR2X1_LOC_749/Y VSS 0.23fF
C2188 AND2X1_LOC_824/B OR2X1_LOC_240/A 0.02fF
C2827 AND2X1_LOC_824/B OR2X1_LOC_334/A 0.01fF
C4720 AND2X1_LOC_824/B OR2X1_LOC_46/A 0.10fF
C6299 AND2X1_LOC_824/B AND2X1_LOC_824/a_8_24# 0.01fF
C9215 AND2X1_LOC_824/B AND2X1_LOC_7/B 0.03fF
C9414 OR2X1_LOC_836/A AND2X1_LOC_824/B 0.01fF
C14541 OR2X1_LOC_19/B AND2X1_LOC_824/B 1.76fF
C18276 AND2X1_LOC_824/B AND2X1_LOC_43/B 0.07fF
C21616 AND2X1_LOC_824/B OR2X1_LOC_410/Y 0.11fF
C25488 AND2X1_LOC_824/B OR2X1_LOC_39/A 0.14fF
C25891 OR2X1_LOC_377/A AND2X1_LOC_824/B 3.84fF
C26317 AND2X1_LOC_824/B OR2X1_LOC_375/A 0.06fF
C29881 AND2X1_LOC_824/B OR2X1_LOC_68/B 2.67fF
C31401 AND2X1_LOC_824/B AND2X1_LOC_291/a_8_24# 0.01fF
C32549 AND2X1_LOC_824/B OR2X1_LOC_461/B 0.05fF
C33851 OR2X1_LOC_461/a_8_216# AND2X1_LOC_824/B 0.04fF
C33888 OR2X1_LOC_634/A AND2X1_LOC_824/B 0.17fF
C35126 OR2X1_LOC_756/B AND2X1_LOC_824/B 0.46fF
C38910 VDD AND2X1_LOC_824/B 0.51fF
C43155 AND2X1_LOC_92/a_8_24# AND2X1_LOC_824/B 0.01fF
C44948 OR2X1_LOC_461/a_36_216# AND2X1_LOC_824/B 0.02fF
C46388 AND2X1_LOC_56/B AND2X1_LOC_824/B 0.26fF
C46406 AND2X1_LOC_8/Y AND2X1_LOC_824/B 0.01fF
C46742 AND2X1_LOC_824/B AND2X1_LOC_92/Y 0.09fF
C47869 AND2X1_LOC_824/B OR2X1_LOC_598/A 0.21fF
C48564 AND2X1_LOC_95/Y AND2X1_LOC_824/B 0.04fF
C52825 AND2X1_LOC_824/B AND2X1_LOC_234/a_8_24# 0.06fF
C55827 OR2X1_LOC_461/Y AND2X1_LOC_824/B 0.01fF
C56986 AND2X1_LOC_824/B VSS 0.22fF
C2146 OR2X1_LOC_377/A OR2X1_LOC_461/A 0.70fF
C6073 OR2X1_LOC_461/A OR2X1_LOC_68/B 0.04fF
C8863 OR2X1_LOC_461/B OR2X1_LOC_461/A 0.32fF
C10154 OR2X1_LOC_461/a_8_216# OR2X1_LOC_461/A 0.47fF
C15199 VDD OR2X1_LOC_461/A 0.01fF
C24002 OR2X1_LOC_461/A OR2X1_LOC_598/A 0.10fF
C24668 AND2X1_LOC_95/Y OR2X1_LOC_461/A 0.14fF
C28886 AND2X1_LOC_413/a_8_24# OR2X1_LOC_461/A 0.01fF
C36939 OR2X1_LOC_46/A OR2X1_LOC_461/A 0.65fF
C56633 OR2X1_LOC_461/A VSS 0.17fF
C4625 OR2X1_LOC_43/A OR2X1_LOC_761/Y 0.01fF
C32410 OR2X1_LOC_696/A OR2X1_LOC_761/Y 0.02fF
C36711 VDD OR2X1_LOC_761/Y 0.12fF
C38057 OR2X1_LOC_761/Y AND2X1_LOC_801/a_8_24# 0.23fF
C46387 OR2X1_LOC_743/A OR2X1_LOC_761/Y 0.01fF
C52088 OR2X1_LOC_761/Y OR2X1_LOC_13/B 0.06fF
C53121 AND2X1_LOC_512/Y OR2X1_LOC_761/Y 0.01fF
C57025 OR2X1_LOC_761/Y VSS 0.06fF
C5437 OR2X1_LOC_275/Y OR2X1_LOC_52/B 0.03fF
C5957 OR2X1_LOC_22/Y OR2X1_LOC_275/Y 0.14fF
C6254 OR2X1_LOC_275/Y OR2X1_LOC_39/A 0.04fF
C10094 OR2X1_LOC_91/A OR2X1_LOC_275/Y 0.03fF
C11041 OR2X1_LOC_74/A OR2X1_LOC_275/Y 0.06fF
C23262 OR2X1_LOC_158/A OR2X1_LOC_275/Y 0.02fF
C25958 OR2X1_LOC_31/Y OR2X1_LOC_275/Y 0.28fF
C28034 AND2X1_LOC_276/Y OR2X1_LOC_275/Y 0.01fF
C44897 OR2X1_LOC_329/B OR2X1_LOC_275/Y 0.08fF
C49298 OR2X1_LOC_517/A OR2X1_LOC_275/Y 0.09fF
C54768 OR2X1_LOC_275/Y AND2X1_LOC_276/a_8_24# 0.05fF
C56598 OR2X1_LOC_275/Y VSS 0.27fF
C1585 AND2X1_LOC_86/Y OR2X1_LOC_66/A 0.01fF
C2951 AND2X1_LOC_86/Y AND2X1_LOC_40/Y 0.09fF
C4363 AND2X1_LOC_86/Y OR2X1_LOC_398/Y 0.03fF
C5798 AND2X1_LOC_86/Y OR2X1_LOC_78/A 0.02fF
C7168 AND2X1_LOC_86/Y OR2X1_LOC_100/a_8_216# 0.18fF
C7617 AND2X1_LOC_86/Y AND2X1_LOC_59/Y 0.13fF
C10215 AND2X1_LOC_86/Y AND2X1_LOC_81/B 0.02fF
C11376 AND2X1_LOC_86/Y OR2X1_LOC_78/B 0.32fF
C11463 AND2X1_LOC_86/Y OR2X1_LOC_375/A 0.02fF
C11762 AND2X1_LOC_86/Y OR2X1_LOC_549/A 0.02fF
C19809 AND2X1_LOC_86/Y AND2X1_LOC_64/Y 0.11fF
C19869 AND2X1_LOC_86/Y AND2X1_LOC_86/a_8_24# 0.01fF
C22083 AND2X1_LOC_86/Y OR2X1_LOC_100/Y 0.02fF
C24148 AND2X1_LOC_86/Y VDD 0.05fF
C26071 AND2X1_LOC_86/Y OR2X1_LOC_80/A 0.16fF
C27173 AND2X1_LOC_86/Y OR2X1_LOC_160/A 0.08fF
C28419 AND2X1_LOC_86/Y OR2X1_LOC_185/A 0.10fF
C31402 AND2X1_LOC_86/Y AND2X1_LOC_8/Y 0.18fF
C32505 AND2X1_LOC_86/Y OR2X1_LOC_6/B 0.20fF
C32789 AND2X1_LOC_86/Y OR2X1_LOC_598/A 0.12fF
C35074 AND2X1_LOC_86/Y AND2X1_LOC_70/Y 0.02fF
C36673 AND2X1_LOC_86/Y AND2X1_LOC_44/Y 0.12fF
C38643 AND2X1_LOC_86/Y OR2X1_LOC_62/B 0.01fF
C38688 AND2X1_LOC_86/Y AND2X1_LOC_88/Y 0.07fF
C42627 AND2X1_LOC_86/Y OR2X1_LOC_71/A 0.01fF
C47983 AND2X1_LOC_86/Y OR2X1_LOC_161/B 0.06fF
C49048 AND2X1_LOC_86/Y AND2X1_LOC_133/a_8_24# 0.03fF
C49572 AND2X1_LOC_86/Y OR2X1_LOC_398/a_8_216# 0.50fF
C58063 AND2X1_LOC_86/Y VSS -0.44fF
C948 AND2X1_LOC_512/Y OR2X1_LOC_599/Y 0.13fF
C1648 AND2X1_LOC_512/Y OR2X1_LOC_511/Y 0.10fF
C7197 AND2X1_LOC_512/Y OR2X1_LOC_485/A 0.02fF
C7838 OR2X1_LOC_696/A AND2X1_LOC_512/Y 0.07fF
C11601 AND2X1_LOC_512/Y OR2X1_LOC_761/a_8_216# 0.01fF
C12173 VDD AND2X1_LOC_512/Y 0.85fF
C13542 AND2X1_LOC_512/Y AND2X1_LOC_801/a_8_24# 0.01fF
C14838 AND2X1_LOC_512/Y OR2X1_LOC_44/Y 0.07fF
C15097 OR2X1_LOC_45/B AND2X1_LOC_512/Y 0.03fF
C15527 OR2X1_LOC_158/A AND2X1_LOC_512/Y 0.07fF
C18133 AND2X1_LOC_512/Y OR2X1_LOC_744/A 0.07fF
C19056 AND2X1_LOC_512/Y AND2X1_LOC_809/A 0.07fF
C19424 AND2X1_LOC_512/Y OR2X1_LOC_56/A 0.07fF
C20025 AND2X1_LOC_512/Y OR2X1_LOC_417/Y 0.07fF
C24555 AND2X1_LOC_512/Y OR2X1_LOC_92/Y 0.07fF
C24928 AND2X1_LOC_512/Y OR2X1_LOC_600/A 0.07fF
C24998 AND2X1_LOC_512/Y OR2X1_LOC_619/Y 0.43fF
C25631 AND2X1_LOC_512/Y OR2X1_LOC_534/a_8_216# 0.03fF
C26160 OR2X1_LOC_329/Y AND2X1_LOC_512/Y 0.02fF
C27346 AND2X1_LOC_512/Y OR2X1_LOC_13/B 0.04fF
C27819 AND2X1_LOC_512/Y OR2X1_LOC_428/A 0.07fF
C28821 AND2X1_LOC_512/Y OR2X1_LOC_26/Y 0.07fF
C29784 AND2X1_LOC_512/Y OR2X1_LOC_95/Y 0.01fF
C30847 AND2X1_LOC_512/Y OR2X1_LOC_59/Y 0.08fF
C30994 OR2X1_LOC_70/Y AND2X1_LOC_512/Y 0.27fF
C31113 AND2X1_LOC_512/Y OR2X1_LOC_534/a_36_216# 0.01fF
C31471 AND2X1_LOC_512/Y OR2X1_LOC_47/Y 0.07fF
C33533 AND2X1_LOC_512/Y AND2X1_LOC_729/B 0.01fF
C33825 AND2X1_LOC_512/Y AND2X1_LOC_513/a_8_24# 0.03fF
C33970 AND2X1_LOC_512/Y OR2X1_LOC_46/A 0.06fF
C34583 OR2X1_LOC_40/Y AND2X1_LOC_512/Y 0.01fF
C34752 AND2X1_LOC_512/Y OR2X1_LOC_7/A 0.07fF
C35993 AND2X1_LOC_512/Y OR2X1_LOC_43/A 0.02fF
C36571 AND2X1_LOC_512/Y OR2X1_LOC_534/Y 0.02fF
C37141 AND2X1_LOC_512/Y OR2X1_LOC_329/B 0.07fF
C38141 AND2X1_LOC_512/Y OR2X1_LOC_64/Y 0.07fF
C39318 AND2X1_LOC_512/Y OR2X1_LOC_516/B 0.02fF
C39835 AND2X1_LOC_512/a_8_24# AND2X1_LOC_512/Y 0.01fF
C45433 AND2X1_LOC_512/Y OR2X1_LOC_36/Y 0.42fF
C45595 AND2X1_LOC_512/Y OR2X1_LOC_419/Y 0.10fF
C45740 OR2X1_LOC_604/A AND2X1_LOC_512/Y 0.07fF
C49475 AND2X1_LOC_512/Y AND2X1_LOC_801/B 0.02fF
C51859 AND2X1_LOC_512/Y OR2X1_LOC_48/B 0.46fF
C54482 AND2X1_LOC_512/Y OR2X1_LOC_22/Y 0.11fF
C54808 AND2X1_LOC_512/Y OR2X1_LOC_39/A 0.10fF
C55576 AND2X1_LOC_512/Y OR2X1_LOC_51/Y 0.01fF
C57751 AND2X1_LOC_512/Y VSS 0.14fF
C5776 OR2X1_LOC_689/a_8_216# OR2X1_LOC_690/Y 0.40fF
C13164 OR2X1_LOC_43/A OR2X1_LOC_690/Y 0.01fF
C15221 OR2X1_LOC_690/Y OR2X1_LOC_690/A 0.01fF
C22201 OR2X1_LOC_689/Y OR2X1_LOC_690/Y 0.09fF
C29228 OR2X1_LOC_690/Y OR2X1_LOC_585/A 0.35fF
C30084 OR2X1_LOC_690/Y OR2X1_LOC_753/A 0.09fF
C45294 VDD OR2X1_LOC_690/Y 0.10fF
C45343 OR2X1_LOC_689/A OR2X1_LOC_690/Y 0.09fF
C48780 OR2X1_LOC_158/A OR2X1_LOC_690/Y 0.03fF
C51545 OR2X1_LOC_690/Y OR2X1_LOC_31/Y 0.02fF
C57318 OR2X1_LOC_690/Y VSS 0.24fF
C4880 OR2X1_LOC_323/A OR2X1_LOC_36/Y 0.04fF
C5201 OR2X1_LOC_323/A OR2X1_LOC_604/A 0.03fF
C6104 OR2X1_LOC_323/A OR2X1_LOC_164/Y 0.02fF
C7924 OR2X1_LOC_323/A OR2X1_LOC_372/Y 0.01fF
C11276 OR2X1_LOC_323/A OR2X1_LOC_18/Y 0.05fF
C12401 OR2X1_LOC_323/A OR2X1_LOC_437/A 0.05fF
C12924 OR2X1_LOC_323/A OR2X1_LOC_323/Y 0.02fF
C13464 OR2X1_LOC_323/A AND2X1_LOC_374/Y 0.02fF
C15065 OR2X1_LOC_323/A OR2X1_LOC_51/Y 0.03fF
C17083 OR2X1_LOC_323/A OR2X1_LOC_268/Y 0.70fF
C18563 OR2X1_LOC_323/A OR2X1_LOC_371/Y 0.02fF
C18989 OR2X1_LOC_323/A OR2X1_LOC_74/A 0.15fF
C22891 OR2X1_LOC_323/A OR2X1_LOC_485/A 0.06fF
C23537 OR2X1_LOC_323/A OR2X1_LOC_696/A 0.15fF
C23660 OR2X1_LOC_323/A AND2X1_LOC_458/Y 0.01fF
C29073 OR2X1_LOC_323/A OR2X1_LOC_427/A 0.05fF
C29112 OR2X1_LOC_323/A OR2X1_LOC_271/a_8_216# 0.01fF
C29957 OR2X1_LOC_323/A OR2X1_LOC_6/A 0.02fF
C30389 OR2X1_LOC_323/A OR2X1_LOC_44/Y 0.03fF
C30672 OR2X1_LOC_45/B OR2X1_LOC_323/A 0.01fF
C31140 OR2X1_LOC_323/A OR2X1_LOC_158/A 0.03fF
C32595 OR2X1_LOC_323/A OR2X1_LOC_111/Y 0.01fF
C33711 OR2X1_LOC_323/A OR2X1_LOC_744/A 0.03fF
C33889 OR2X1_LOC_323/A OR2X1_LOC_31/Y 0.22fF
C34267 OR2X1_LOC_323/A AND2X1_LOC_270/a_8_24# 0.01fF
C34977 OR2X1_LOC_323/A OR2X1_LOC_56/A 0.69fF
C35442 OR2X1_LOC_323/A OR2X1_LOC_371/a_8_216# 0.01fF
C40031 OR2X1_LOC_323/A OR2X1_LOC_92/Y 0.03fF
C40078 OR2X1_LOC_323/A OR2X1_LOC_271/Y 0.01fF
C40435 OR2X1_LOC_323/A OR2X1_LOC_600/A 0.03fF
C40564 OR2X1_LOC_323/A OR2X1_LOC_372/a_8_216# 0.01fF
C43000 OR2X1_LOC_323/A OR2X1_LOC_111/a_8_216# 0.01fF
C43438 OR2X1_LOC_323/A OR2X1_LOC_428/A 0.24fF
C44432 OR2X1_LOC_323/A OR2X1_LOC_26/Y 0.03fF
C45415 OR2X1_LOC_323/A OR2X1_LOC_95/Y 0.06fF
C45420 OR2X1_LOC_323/A OR2X1_LOC_368/A 0.50fF
C47253 OR2X1_LOC_323/A OR2X1_LOC_47/Y 0.02fF
C50536 OR2X1_LOC_323/A OR2X1_LOC_7/A 0.10fF
C51674 OR2X1_LOC_323/A OR2X1_LOC_322/Y 0.02fF
C52980 OR2X1_LOC_323/A OR2X1_LOC_329/B 0.03fF
C53925 OR2X1_LOC_323/A OR2X1_LOC_64/Y 0.24fF
C53974 OR2X1_LOC_323/A OR2X1_LOC_417/A 0.13fF
C58105 OR2X1_LOC_323/A VSS 0.79fF
C475 OR2X1_LOC_485/A OR2X1_LOC_743/A 2.04fF
C1126 OR2X1_LOC_696/A OR2X1_LOC_743/A 2.59fF
C2436 OR2X1_LOC_743/A OR2X1_LOC_743/Y 0.02fF
C3033 OR2X1_LOC_743/A OR2X1_LOC_422/Y 0.21fF
C3163 OR2X1_LOC_743/A OR2X1_LOC_760/Y 0.09fF
C4826 OR2X1_LOC_743/A OR2X1_LOC_761/a_8_216# 0.01fF
C5114 OR2X1_LOC_682/a_8_216# OR2X1_LOC_743/A 0.01fF
C5410 VDD OR2X1_LOC_743/A 0.87fF
C5503 OR2X1_LOC_743/A AND2X1_LOC_274/a_8_24# 0.24fF
C6783 OR2X1_LOC_743/A OR2X1_LOC_427/A 0.13fF
C6787 OR2X1_LOC_743/A AND2X1_LOC_801/a_8_24# 0.01fF
C7316 OR2X1_LOC_743/A OR2X1_LOC_681/Y 0.02fF
C7704 OR2X1_LOC_743/A OR2X1_LOC_6/A 0.03fF
C8165 OR2X1_LOC_743/A OR2X1_LOC_44/Y 0.21fF
C8448 OR2X1_LOC_45/B OR2X1_LOC_743/A 0.29fF
C8878 OR2X1_LOC_158/A OR2X1_LOC_743/A 0.10fF
C11461 OR2X1_LOC_744/A OR2X1_LOC_743/A 0.14fF
C11620 OR2X1_LOC_743/A OR2X1_LOC_31/Y 1.42fF
C12729 OR2X1_LOC_743/A OR2X1_LOC_56/A 0.06fF
C13322 OR2X1_LOC_417/Y OR2X1_LOC_743/A 0.03fF
C14842 OR2X1_LOC_426/B OR2X1_LOC_743/A 6.55fF
C15022 OR2X1_LOC_743/A OR2X1_LOC_246/A 2.92fF
C15658 OR2X1_LOC_743/A OR2X1_LOC_743/a_8_216# 0.09fF
C17824 OR2X1_LOC_743/A OR2X1_LOC_92/Y 0.12fF
C18319 OR2X1_LOC_743/A OR2X1_LOC_619/Y 0.10fF
C20663 OR2X1_LOC_743/A OR2X1_LOC_13/B 0.18fF
C21184 OR2X1_LOC_743/A OR2X1_LOC_428/A 0.11fF
C21803 OR2X1_LOC_682/Y OR2X1_LOC_743/A 0.38fF
C22632 OR2X1_LOC_306/a_8_216# OR2X1_LOC_743/A 0.03fF
C23143 OR2X1_LOC_743/A OR2X1_LOC_95/Y 0.06fF
C24321 OR2X1_LOC_743/A OR2X1_LOC_433/a_8_216# 0.01fF
C24349 OR2X1_LOC_70/Y OR2X1_LOC_743/A 0.35fF
C24824 OR2X1_LOC_743/A OR2X1_LOC_47/Y 0.03fF
C25801 OR2X1_LOC_743/A OR2X1_LOC_16/A 0.08fF
C25991 OR2X1_LOC_743/A OR2X1_LOC_273/a_8_216# 0.01fF
C26857 OR2X1_LOC_743/A AND2X1_LOC_729/B 0.62fF
C27308 OR2X1_LOC_743/A OR2X1_LOC_46/A 0.14fF
C27664 OR2X1_LOC_599/A OR2X1_LOC_743/A 0.10fF
C27963 OR2X1_LOC_40/Y OR2X1_LOC_743/A 0.03fF
C28115 OR2X1_LOC_743/A OR2X1_LOC_7/A 0.16fF
C29203 OR2X1_LOC_589/A OR2X1_LOC_743/A 0.12fF
C29352 OR2X1_LOC_43/A OR2X1_LOC_743/A 0.10fF
C29402 OR2X1_LOC_743/A AND2X1_LOC_685/a_8_24# 0.19fF
C30219 OR2X1_LOC_3/Y OR2X1_LOC_743/A 13.39fF
C31487 OR2X1_LOC_743/A OR2X1_LOC_273/a_36_216# 0.01fF
C31506 OR2X1_LOC_743/A OR2X1_LOC_64/Y 0.15fF
C31535 OR2X1_LOC_743/A OR2X1_LOC_417/A 0.03fF
C33023 OR2X1_LOC_421/A OR2X1_LOC_743/A 0.04fF
C33159 AND2X1_LOC_512/a_8_24# OR2X1_LOC_743/A 0.01fF
C33571 OR2X1_LOC_306/a_36_216# OR2X1_LOC_743/A 0.02fF
C33692 OR2X1_LOC_743/A AND2X1_LOC_687/a_8_24# 0.08fF
C35244 OR2X1_LOC_743/A OR2X1_LOC_433/a_36_216# 0.03fF
C35973 OR2X1_LOC_681/a_8_216# OR2X1_LOC_743/A 0.07fF
C36766 OR2X1_LOC_743/A OR2X1_LOC_421/Y 1.01fF
C36941 OR2X1_LOC_743/A OR2X1_LOC_273/Y 0.27fF
C37394 OR2X1_LOC_743/A OR2X1_LOC_275/A 0.01fF
C37573 OR2X1_LOC_136/a_8_216# OR2X1_LOC_743/A 0.04fF
C38007 OR2X1_LOC_743/A AND2X1_LOC_407/a_8_24# 0.11fF
C38638 OR2X1_LOC_743/A OR2X1_LOC_36/Y 0.25fF
C38959 OR2X1_LOC_604/A OR2X1_LOC_743/A 0.61fF
C39066 OR2X1_LOC_306/Y OR2X1_LOC_743/A 0.01fF
C39931 AND2X1_LOC_155/Y OR2X1_LOC_743/A 0.01fF
C40376 OR2X1_LOC_743/A AND2X1_LOC_687/A 0.07fF
C41512 OR2X1_LOC_681/a_36_216# OR2X1_LOC_743/A 0.03fF
C42344 OR2X1_LOC_743/A OR2X1_LOC_12/Y 0.12fF
C42472 OR2X1_LOC_743/A OR2X1_LOC_422/a_8_216# 0.01fF
C42555 OR2X1_LOC_272/Y OR2X1_LOC_743/A 0.09fF
C42595 OR2X1_LOC_743/A AND2X1_LOC_801/B 0.03fF
C45070 OR2X1_LOC_743/A OR2X1_LOC_48/B 0.11fF
C45077 OR2X1_LOC_743/A OR2X1_LOC_18/Y 0.14fF
C45559 OR2X1_LOC_743/A OR2X1_LOC_585/A 0.05fF
C46157 OR2X1_LOC_743/A OR2X1_LOC_437/A 0.07fF
C47369 OR2X1_LOC_743/A OR2X1_LOC_52/B 0.08fF
C47844 OR2X1_LOC_743/A OR2X1_LOC_22/Y 0.28fF
C48212 OR2X1_LOC_743/A OR2X1_LOC_39/A 1.05fF
C48567 OR2X1_LOC_421/a_8_216# OR2X1_LOC_743/A 0.01fF
C48859 OR2X1_LOC_136/Y OR2X1_LOC_743/A 0.03fF
C48951 OR2X1_LOC_51/Y OR2X1_LOC_743/A 0.06fF
C50449 OR2X1_LOC_743/A OR2X1_LOC_599/Y 0.03fF
C51910 OR2X1_LOC_743/A OR2X1_LOC_91/A 0.07fF
C52879 OR2X1_LOC_743/A OR2X1_LOC_74/A -0.01fF
C53218 AND2X1_LOC_155/a_8_24# OR2X1_LOC_743/A 0.05fF
C54682 OR2X1_LOC_743/A OR2X1_LOC_300/Y 0.12fF
C55866 OR2X1_LOC_696/Y OR2X1_LOC_743/A 0.02fF
C57367 OR2X1_LOC_743/A VSS 0.42fF
C15693 OR2X1_LOC_18/Y OR2X1_LOC_372/Y 0.01fF
C17872 OR2X1_LOC_372/Y AND2X1_LOC_374/Y 0.21fF
C19483 OR2X1_LOC_51/Y OR2X1_LOC_372/Y 0.06fF
C23078 OR2X1_LOC_372/Y OR2X1_LOC_371/Y 0.12fF
C35054 OR2X1_LOC_45/B OR2X1_LOC_372/Y 0.01fF
C44950 OR2X1_LOC_600/A OR2X1_LOC_372/Y 0.06fF
C49020 OR2X1_LOC_26/Y OR2X1_LOC_372/Y 0.03fF
C49970 OR2X1_LOC_95/Y OR2X1_LOC_372/Y 0.02fF
C56576 OR2X1_LOC_372/Y VSS -0.02fF
C37 AND2X1_LOC_687/Y OR2X1_LOC_48/B 0.02fF
C229 OR2X1_LOC_48/B OR2X1_LOC_373/Y 0.02fF
C881 AND2X1_LOC_729/B OR2X1_LOC_48/B 0.03fF
C1208 AND2X1_LOC_513/a_8_24# OR2X1_LOC_48/B 0.03fF
C1351 OR2X1_LOC_46/A OR2X1_LOC_48/B 0.04fF
C1703 OR2X1_LOC_599/A OR2X1_LOC_48/B 0.79fF
C1996 OR2X1_LOC_40/Y OR2X1_LOC_48/B 6.64fF
C2162 OR2X1_LOC_7/A OR2X1_LOC_48/B 0.91fF
C2271 OR2X1_LOC_48/B OR2X1_LOC_511/a_8_216# 0.02fF
C3278 OR2X1_LOC_589/A OR2X1_LOC_48/B 0.35fF
C3426 OR2X1_LOC_43/A OR2X1_LOC_48/B 0.32fF
C4244 OR2X1_LOC_3/Y OR2X1_LOC_48/B 0.15fF
C4532 OR2X1_LOC_329/B OR2X1_LOC_48/B 0.14fF
C5526 OR2X1_LOC_64/Y OR2X1_LOC_48/B 0.26fF
C6680 OR2X1_LOC_516/B OR2X1_LOC_48/B 0.03fF
C7065 OR2X1_LOC_421/A OR2X1_LOC_48/B 0.09fF
C9821 OR2X1_LOC_763/Y OR2X1_LOC_48/B 0.01fF
C10254 OR2X1_LOC_48/Y OR2X1_LOC_48/B 0.28fF
C10961 OR2X1_LOC_763/a_8_216# OR2X1_LOC_48/B 0.10fF
C12621 AND2X1_LOC_596/a_8_24# OR2X1_LOC_48/B 0.02fF
C12757 OR2X1_LOC_36/Y OR2X1_LOC_48/B 0.15fF
C13090 OR2X1_LOC_604/A OR2X1_LOC_48/B 0.05fF
C13870 OR2X1_LOC_304/a_8_216# OR2X1_LOC_48/B 0.04fF
C16366 OR2X1_LOC_48/B OR2X1_LOC_12/Y 3.68fF
C18141 OR2X1_LOC_597/A OR2X1_LOC_48/B 0.12fF
C19100 OR2X1_LOC_18/Y OR2X1_LOC_48/B 1.89fF
C19584 OR2X1_LOC_585/A OR2X1_LOC_48/B 0.10fF
C20185 OR2X1_LOC_48/B OR2X1_LOC_437/A 0.04fF
C21300 OR2X1_LOC_48/B OR2X1_LOC_52/B 0.20fF
C21702 OR2X1_LOC_48/B OR2X1_LOC_48/a_8_216# 0.03fF
C21795 OR2X1_LOC_22/Y OR2X1_LOC_48/B 0.37fF
C21858 OR2X1_LOC_48/B OR2X1_LOC_387/a_8_216# 0.05fF
C22130 OR2X1_LOC_48/B OR2X1_LOC_39/A 0.07fF
C22916 OR2X1_LOC_51/Y OR2X1_LOC_48/B 0.07fF
C23721 AND2X1_LOC_596/a_36_24# OR2X1_LOC_48/B 0.01fF
C25798 OR2X1_LOC_91/A OR2X1_LOC_48/B 0.21fF
C26781 OR2X1_LOC_74/A OR2X1_LOC_48/B 0.07fF
C27186 OR2X1_LOC_48/B OR2X1_LOC_48/a_36_216# 0.01fF
C29756 OR2X1_LOC_696/Y OR2X1_LOC_48/B 0.02fF
C30562 OR2X1_LOC_485/A OR2X1_LOC_48/B 0.09fF
C31197 OR2X1_LOC_696/A OR2X1_LOC_48/B 3.00fF
C33029 OR2X1_LOC_519/a_8_216# OR2X1_LOC_48/B 0.05fF
C33041 OR2X1_LOC_48/B OR2X1_LOC_433/Y 0.03fF
C35480 VDD OR2X1_LOC_48/B 1.05fF
C36800 OR2X1_LOC_427/A OR2X1_LOC_48/B 0.09fF
C37692 OR2X1_LOC_6/A OR2X1_LOC_48/B 0.01fF
C38109 OR2X1_LOC_48/B OR2X1_LOC_44/Y 2.73fF
C38364 OR2X1_LOC_45/B OR2X1_LOC_48/B 0.30fF
C38425 AND2X1_LOC_410/a_8_24# OR2X1_LOC_48/B 0.23fF
C38864 OR2X1_LOC_158/A OR2X1_LOC_48/B 0.25fF
C39484 OR2X1_LOC_304/Y OR2X1_LOC_48/B 0.21fF
C41463 OR2X1_LOC_744/A OR2X1_LOC_48/B 1.17fF
C41670 OR2X1_LOC_31/Y OR2X1_LOC_48/B 0.38fF
C42770 OR2X1_LOC_56/A OR2X1_LOC_48/B 0.15fF
C43364 OR2X1_LOC_417/Y OR2X1_LOC_48/B 0.07fF
C43770 OR2X1_LOC_696/a_8_216# OR2X1_LOC_48/B 0.02fF
C44910 OR2X1_LOC_426/B OR2X1_LOC_48/B 0.24fF
C45146 OR2X1_LOC_409/B OR2X1_LOC_48/B 0.12fF
C47045 OR2X1_LOC_48/B OR2X1_LOC_387/A 0.05fF
C47566 OR2X1_LOC_693/a_8_216# OR2X1_LOC_48/B 0.02fF
C48086 OR2X1_LOC_692/a_8_216# OR2X1_LOC_48/B 0.03fF
C48092 OR2X1_LOC_92/Y OR2X1_LOC_48/B 0.13fF
C48432 OR2X1_LOC_692/Y OR2X1_LOC_48/B 0.02fF
C48467 OR2X1_LOC_600/A OR2X1_LOC_48/B 0.07fF
C48550 OR2X1_LOC_619/Y OR2X1_LOC_48/B 0.14fF
C50595 OR2X1_LOC_762/Y OR2X1_LOC_48/B 0.29fF
C50874 OR2X1_LOC_48/B OR2X1_LOC_13/B 0.57fF
C51342 OR2X1_LOC_48/B OR2X1_LOC_428/A 0.53fF
C51904 OR2X1_LOC_516/A OR2X1_LOC_48/B 0.03fF
C52346 AND2X1_LOC_598/a_8_24# OR2X1_LOC_48/B 0.10fF
C52358 OR2X1_LOC_26/Y OR2X1_LOC_48/B 0.17fF
C52382 OR2X1_LOC_89/A OR2X1_LOC_48/B 0.32fF
C53289 OR2X1_LOC_95/Y OR2X1_LOC_48/B 0.03fF
C53883 OR2X1_LOC_693/Y OR2X1_LOC_48/B 0.01fF
C54340 OR2X1_LOC_48/B OR2X1_LOC_59/Y 11.05fF
C54449 OR2X1_LOC_433/a_8_216# OR2X1_LOC_48/B 0.02fF
C54481 OR2X1_LOC_70/Y OR2X1_LOC_48/B 0.17fF
C54506 AND2X1_LOC_514/Y OR2X1_LOC_48/B 0.03fF
C54979 OR2X1_LOC_47/Y OR2X1_LOC_48/B 0.18fF
C56000 OR2X1_LOC_48/B OR2X1_LOC_16/A 0.11fF
C56694 OR2X1_LOC_48/B VSS 0.90fF
C2513 OR2X1_LOC_9/Y OR2X1_LOC_485/A 0.11fF
C2776 OR2X1_LOC_9/Y OR2X1_LOC_633/A 0.04fF
C3162 OR2X1_LOC_696/A OR2X1_LOC_9/Y 1.74fF
C3256 OR2X1_LOC_9/Y AND2X1_LOC_819/a_8_24# 0.01fF
C4820 OR2X1_LOC_49/A OR2X1_LOC_9/Y 0.06fF
C5228 OR2X1_LOC_9/Y OR2X1_LOC_671/Y 0.02fF
C6246 OR2X1_LOC_9/Y AND2X1_LOC_42/B 0.01fF
C7446 OR2X1_LOC_9/Y VDD 0.72fF
C8002 OR2X1_LOC_9/Y OR2X1_LOC_6/a_8_216# 0.03fF
C8782 OR2X1_LOC_9/Y AND2X1_LOC_820/B 0.01fF
C9494 OR2X1_LOC_9/Y OR2X1_LOC_80/A 0.61fF
C9702 OR2X1_LOC_9/Y OR2X1_LOC_6/A 0.48fF
C10835 OR2X1_LOC_9/Y OR2X1_LOC_158/A 0.29fF
C10911 OR2X1_LOC_9/Y OR2X1_LOC_847/A 0.02fF
C13161 OR2X1_LOC_9/Y OR2X1_LOC_824/a_8_216# 0.01fF
C14701 OR2X1_LOC_9/Y OR2X1_LOC_56/A 0.07fF
C14754 OR2X1_LOC_9/Y AND2X1_LOC_9/a_8_24# 0.01fF
C15909 OR2X1_LOC_9/Y OR2X1_LOC_6/B 0.18fF
C16744 OR2X1_LOC_9/Y OR2X1_LOC_15/a_8_216# 0.05fF
C16990 OR2X1_LOC_9/Y OR2X1_LOC_246/A 0.14fF
C18082 OR2X1_LOC_9/Y OR2X1_LOC_235/B 0.34fF
C19015 OR2X1_LOC_9/Y OR2X1_LOC_96/B 0.73fF
C20224 OR2X1_LOC_9/Y OR2X1_LOC_600/A 0.08fF
C20280 OR2X1_LOC_9/Y OR2X1_LOC_619/Y 0.01fF
C22145 OR2X1_LOC_9/Y OR2X1_LOC_62/B 0.01fF
C23181 OR2X1_LOC_9/Y OR2X1_LOC_428/A 0.09fF
C23824 OR2X1_LOC_9/Y OR2X1_LOC_54/Y 3.68fF
C24179 OR2X1_LOC_9/Y OR2X1_LOC_26/Y 0.05fF
C24553 OR2X1_LOC_9/Y OR2X1_LOC_246/a_8_216# 0.07fF
C24975 OR2X1_LOC_9/Y OR2X1_LOC_824/Y 0.04fF
C25089 OR2X1_LOC_9/Y OR2X1_LOC_95/Y 0.03fF
C26788 OR2X1_LOC_9/Y OR2X1_LOC_47/Y 0.07fF
C27481 OR2X1_LOC_9/Y OR2X1_LOC_246/Y 0.35fF
C29257 OR2X1_LOC_9/Y OR2X1_LOC_46/A 0.39fF
C29917 OR2X1_LOC_9/Y OR2X1_LOC_159/a_8_216# 0.06fF
C29919 OR2X1_LOC_9/Y OR2X1_LOC_40/Y 0.76fF
C30024 OR2X1_LOC_9/Y OR2X1_LOC_618/a_8_216# 0.01fF
C31311 OR2X1_LOC_9/Y OR2X1_LOC_43/A 2.80fF
C32467 OR2X1_LOC_9/Y OR2X1_LOC_502/A 0.08fF
C32683 OR2X1_LOC_9/Y OR2X1_LOC_618/Y 0.01fF
C37132 OR2X1_LOC_9/Y AND2X1_LOC_62/a_8_24# 0.25fF
C40881 OR2X1_LOC_9/Y OR2X1_LOC_604/A 0.04fF
C42607 OR2X1_LOC_143/a_8_216# OR2X1_LOC_9/Y 0.01fF
C43684 OR2X1_LOC_9/Y OR2X1_LOC_73/a_8_216# 0.02fF
C43780 OR2X1_LOC_9/Y OR2X1_LOC_619/a_8_216# 0.01fF
C47643 OR2X1_LOC_9/Y OR2X1_LOC_585/A 0.01fF
C48290 OR2X1_LOC_9/Y OR2X1_LOC_437/A 0.09fF
C48502 OR2X1_LOC_9/Y OR2X1_LOC_753/A 0.03fF
C49006 OR2X1_LOC_9/Y OR2X1_LOC_62/A 0.83fF
C49196 OR2X1_LOC_8/Y OR2X1_LOC_9/Y 2.63fF
C49324 OR2X1_LOC_9/Y OR2X1_LOC_672/Y 0.53fF
C49346 OR2X1_LOC_9/Y OR2X1_LOC_73/a_36_216# 0.03fF
C50570 OR2X1_LOC_9/Y OR2X1_LOC_85/A 0.36fF
C50912 OR2X1_LOC_9/Y OR2X1_LOC_51/Y 0.05fF
C54537 OR2X1_LOC_9/Y OR2X1_LOC_68/B 0.10fF
C54801 OR2X1_LOC_9/Y OR2X1_LOC_74/A 0.53fF
C57896 OR2X1_LOC_9/Y VSS 0.52fF
C5 OR2X1_LOC_633/A OR2X1_LOC_598/A 0.32fF
C407 AND2X1_LOC_64/Y OR2X1_LOC_598/A 0.15fF
C962 OR2X1_LOC_756/B OR2X1_LOC_598/A 0.07fF
C2189 OR2X1_LOC_49/A OR2X1_LOC_598/A 0.03fF
C2815 OR2X1_LOC_532/B OR2X1_LOC_598/A 0.31fF
C3615 AND2X1_LOC_42/B OR2X1_LOC_598/A 0.14fF
C3998 OR2X1_LOC_185/Y OR2X1_LOC_598/A 0.10fF
C4718 VDD OR2X1_LOC_598/A 0.98fF
C6650 OR2X1_LOC_80/A OR2X1_LOC_598/A 0.17fF
C6931 OR2X1_LOC_6/A OR2X1_LOC_598/A 0.12fF
C7793 OR2X1_LOC_160/A OR2X1_LOC_598/A 0.30fF
C8158 OR2X1_LOC_158/A OR2X1_LOC_598/A 0.10fF
C9094 OR2X1_LOC_185/A OR2X1_LOC_598/A 0.10fF
C10752 OR2X1_LOC_744/A OR2X1_LOC_598/A 0.04fF
C10864 OR2X1_LOC_31/Y OR2X1_LOC_598/A 0.06fF
C11164 OR2X1_LOC_264/Y OR2X1_LOC_598/A 0.01fF
C11502 AND2X1_LOC_91/B OR2X1_LOC_598/A 0.10fF
C12051 AND2X1_LOC_56/B OR2X1_LOC_598/A 0.08fF
C12057 AND2X1_LOC_8/Y OR2X1_LOC_598/A 0.10fF
C12951 OR2X1_LOC_83/A OR2X1_LOC_598/A 0.02fF
C13300 OR2X1_LOC_6/B OR2X1_LOC_598/A 0.26fF
C13448 AND2X1_LOC_47/Y OR2X1_LOC_598/A 0.14fF
C14199 AND2X1_LOC_95/Y OR2X1_LOC_598/A 0.22fF
C14255 OR2X1_LOC_415/a_8_216# OR2X1_LOC_598/A 0.03fF
C14493 AND2X1_LOC_22/Y OR2X1_LOC_598/A 0.11fF
C14648 OR2X1_LOC_296/a_8_216# OR2X1_LOC_598/A -0.02fF
C15777 AND2X1_LOC_70/Y OR2X1_LOC_598/A 1.43fF
C17039 AND2X1_LOC_256/a_8_24# OR2X1_LOC_598/A 0.01fF
C17433 AND2X1_LOC_44/Y OR2X1_LOC_598/A 0.08fF
C18370 AND2X1_LOC_18/Y OR2X1_LOC_598/A 0.14fF
C18444 AND2X1_LOC_413/a_8_24# OR2X1_LOC_598/A 0.01fF
C19791 OR2X1_LOC_415/a_36_216# OR2X1_LOC_598/A 0.03fF
C21052 OR2X1_LOC_54/Y OR2X1_LOC_598/A 0.19fF
C21449 OR2X1_LOC_161/A OR2X1_LOC_598/A 0.02fF
C21499 OR2X1_LOC_461/Y OR2X1_LOC_598/A 0.01fF
C21502 AND2X1_LOC_51/Y OR2X1_LOC_598/A 2.38fF
C22261 AND2X1_LOC_41/A OR2X1_LOC_598/A 0.78fF
C22325 OR2X1_LOC_688/a_8_216# OR2X1_LOC_598/A 0.05fF
C23734 AND2X1_LOC_31/Y OR2X1_LOC_598/A 0.03fF
C24024 OR2X1_LOC_240/A OR2X1_LOC_598/A 0.01fF
C24099 OR2X1_LOC_47/Y OR2X1_LOC_598/A 0.09fF
C24634 AND2X1_LOC_36/Y OR2X1_LOC_598/A 0.35fF
C24672 OR2X1_LOC_598/A OR2X1_LOC_334/A 0.03fF
C26352 OR2X1_LOC_598/A OR2X1_LOC_548/a_8_216# 0.01fF
C26542 OR2X1_LOC_46/A OR2X1_LOC_598/A 1.33fF
C26920 OR2X1_LOC_269/B OR2X1_LOC_598/A 0.03fF
C27312 AND2X1_LOC_690/a_8_24# OR2X1_LOC_598/A 0.08fF
C27642 OR2X1_LOC_691/A OR2X1_LOC_598/A 0.03fF
C27707 OR2X1_LOC_294/a_8_216# OR2X1_LOC_598/A 0.01fF
C27972 OR2X1_LOC_777/B OR2X1_LOC_598/A 0.07fF
C28491 OR2X1_LOC_161/B OR2X1_LOC_598/A 0.88fF
C28971 OR2X1_LOC_630/B OR2X1_LOC_598/A 0.02fF
C29354 AND2X1_LOC_625/a_8_24# OR2X1_LOC_598/A -0.00fF
C29464 OR2X1_LOC_3/Y OR2X1_LOC_598/A 0.02fF
C29560 AND2X1_LOC_462/B OR2X1_LOC_598/A 0.02fF
C29830 OR2X1_LOC_502/A OR2X1_LOC_598/A 0.03fF
C29920 AND2X1_LOC_48/A OR2X1_LOC_598/A 0.04fF
C30181 AND2X1_LOC_530/a_8_24# OR2X1_LOC_598/A 0.01fF
C30311 AND2X1_LOC_3/Y OR2X1_LOC_598/A 0.70fF
C30691 OR2X1_LOC_690/A OR2X1_LOC_598/A 0.31fF
C31015 AND2X1_LOC_7/B OR2X1_LOC_598/A 0.27fF
C32031 OR2X1_LOC_473/A OR2X1_LOC_598/A 0.75fF
C32741 OR2X1_LOC_160/B OR2X1_LOC_598/A 0.14fF
C33592 OR2X1_LOC_151/A OR2X1_LOC_598/A 0.84fF
C34793 OR2X1_LOC_415/Y OR2X1_LOC_598/A 0.20fF
C34862 OR2X1_LOC_631/A OR2X1_LOC_598/A 0.03fF
C35324 OR2X1_LOC_49/a_8_216# OR2X1_LOC_598/A 0.11fF
C35665 OR2X1_LOC_548/A OR2X1_LOC_598/A 0.01fF
C35885 OR2X1_LOC_66/a_8_216# OR2X1_LOC_598/A 0.02fF
C36230 OR2X1_LOC_19/B OR2X1_LOC_598/A 0.09fF
C38221 OR2X1_LOC_66/A OR2X1_LOC_598/A 0.11fF
C38619 AND2X1_LOC_585/a_8_24# OR2X1_LOC_598/A 0.06fF
C39571 AND2X1_LOC_40/Y OR2X1_LOC_598/A 0.08fF
C39972 AND2X1_LOC_43/B OR2X1_LOC_598/A 0.11fF
C40331 AND2X1_LOC_625/a_36_24# OR2X1_LOC_598/A 0.01fF
C42556 OR2X1_LOC_78/A OR2X1_LOC_598/A 0.25fF
C43099 OR2X1_LOC_814/A OR2X1_LOC_598/A 0.07fF
C43799 OR2X1_LOC_121/Y OR2X1_LOC_598/A 0.03fF
C43897 AND2X1_LOC_12/Y OR2X1_LOC_598/A 0.22fF
C44333 AND2X1_LOC_59/Y OR2X1_LOC_598/A 0.01fF
C44774 OR2X1_LOC_585/A OR2X1_LOC_598/A 0.02fF
C45649 OR2X1_LOC_753/A OR2X1_LOC_598/A 1.12fF
C46553 OR2X1_LOC_52/B OR2X1_LOC_598/A 0.34fF
C46978 AND2X1_LOC_81/B OR2X1_LOC_598/A 0.01fF
C46980 AND2X1_LOC_49/a_8_24# OR2X1_LOC_598/A 0.04fF
C47054 OR2X1_LOC_22/Y OR2X1_LOC_598/A 0.03fF
C47130 OR2X1_LOC_66/Y OR2X1_LOC_598/A 0.09fF
C47446 OR2X1_LOC_39/A OR2X1_LOC_598/A 0.06fF
C47864 OR2X1_LOC_377/A OR2X1_LOC_598/A 0.49fF
C48267 OR2X1_LOC_78/B OR2X1_LOC_598/A 0.23fF
C48323 OR2X1_LOC_375/A OR2X1_LOC_598/A 0.25fF
C48623 OR2X1_LOC_598/A OR2X1_LOC_549/A 1.50fF
C49479 AND2X1_LOC_65/A OR2X1_LOC_598/A 0.09fF
C50794 OR2X1_LOC_769/B OR2X1_LOC_598/A 0.03fF
C51657 OR2X1_LOC_32/B OR2X1_LOC_598/A 0.46fF
C51840 OR2X1_LOC_68/B OR2X1_LOC_598/A 0.08fF
C52342 OR2X1_LOC_598/a_8_216# OR2X1_LOC_598/A 0.04fF
C52511 OR2X1_LOC_87/A OR2X1_LOC_598/A 0.10fF
C53344 AND2X1_LOC_291/a_8_24# OR2X1_LOC_598/A 0.02fF
C54525 OR2X1_LOC_461/B OR2X1_LOC_598/A 0.02fF
C55016 OR2X1_LOC_154/A OR2X1_LOC_598/A 0.29fF
C55136 AND2X1_LOC_6/a_8_24# OR2X1_LOC_598/A 0.02fF
C55852 OR2X1_LOC_461/a_8_216# OR2X1_LOC_598/A 0.01fF
C55871 OR2X1_LOC_634/A OR2X1_LOC_598/A 0.56fF
C56342 OR2X1_LOC_598/A VSS -4.30fF
C456 OR2X1_LOC_164/Y OR2X1_LOC_417/A 0.07fF
C2994 OR2X1_LOC_417/A OR2X1_LOC_12/Y 0.07fF
C3961 OR2X1_LOC_283/Y OR2X1_LOC_417/A 0.07fF
C5561 OR2X1_LOC_18/Y OR2X1_LOC_417/A 1.28fF
C6609 OR2X1_LOC_417/A OR2X1_LOC_437/A 1.39fF
C6905 OR2X1_LOC_417/A OR2X1_LOC_753/A 0.07fF
C8289 OR2X1_LOC_22/Y OR2X1_LOC_417/A 0.31fF
C8652 OR2X1_LOC_417/A OR2X1_LOC_39/A 0.07fF
C9135 OR2X1_LOC_417/A OR2X1_LOC_226/Y 0.05fF
C9432 OR2X1_LOC_51/Y OR2X1_LOC_417/A 1.54fF
C12385 OR2X1_LOC_91/A OR2X1_LOC_417/A 0.77fF
C12916 OR2X1_LOC_417/A OR2X1_LOC_371/Y 0.07fF
C13357 OR2X1_LOC_74/A OR2X1_LOC_417/A 0.75fF
C15444 OR2X1_LOC_417/A AND2X1_LOC_814/a_8_24# 0.11fF
C15834 OR2X1_LOC_417/a_8_216# OR2X1_LOC_417/A 0.02fF
C17136 OR2X1_LOC_485/A OR2X1_LOC_417/A 0.12fF
C17736 OR2X1_LOC_696/A OR2X1_LOC_417/A 0.41fF
C17943 OR2X1_LOC_417/A AND2X1_LOC_458/Y 0.03fF
C20894 OR2X1_LOC_369/Y OR2X1_LOC_417/A -0.00fF
C22179 VDD OR2X1_LOC_417/A 1.16fF
C23070 OR2X1_LOC_382/Y OR2X1_LOC_417/A 0.01fF
C23515 OR2X1_LOC_427/A OR2X1_LOC_417/A 0.17fF
C24783 OR2X1_LOC_417/A OR2X1_LOC_44/Y 0.17fF
C25040 OR2X1_LOC_45/B OR2X1_LOC_417/A 0.06fF
C25489 OR2X1_LOC_158/A OR2X1_LOC_417/A 0.20fF
C26079 OR2X1_LOC_628/Y OR2X1_LOC_417/A 0.04fF
C26932 OR2X1_LOC_111/Y OR2X1_LOC_417/A 0.03fF
C28044 OR2X1_LOC_309/Y OR2X1_LOC_417/A 0.19fF
C28075 OR2X1_LOC_744/A OR2X1_LOC_417/A 4.19fF
C28218 OR2X1_LOC_31/Y OR2X1_LOC_417/A 0.17fF
C28591 OR2X1_LOC_488/a_8_216# OR2X1_LOC_417/A 0.01fF
C29318 OR2X1_LOC_417/A OR2X1_LOC_56/A 0.28fF
C30633 OR2X1_LOC_519/Y OR2X1_LOC_417/A 0.01fF
C30668 OR2X1_LOC_529/Y OR2X1_LOC_417/A 0.03fF
C31162 OR2X1_LOC_71/Y OR2X1_LOC_417/A 0.03fF
C31422 OR2X1_LOC_426/B OR2X1_LOC_417/A 0.20fF
C31564 OR2X1_LOC_246/A OR2X1_LOC_417/A 0.03fF
C31577 OR2X1_LOC_225/a_8_216# OR2X1_LOC_417/A 0.05fF
C34396 OR2X1_LOC_92/Y OR2X1_LOC_417/A 0.10fF
C34803 OR2X1_LOC_600/A OR2X1_LOC_417/A 0.42fF
C36878 OR2X1_LOC_666/A OR2X1_LOC_417/A 0.24fF
C37142 OR2X1_LOC_417/A OR2X1_LOC_13/B 0.14fF
C37211 OR2X1_LOC_111/a_8_216# OR2X1_LOC_417/A 0.02fF
C37674 OR2X1_LOC_417/A OR2X1_LOC_428/A 1.09fF
C38698 OR2X1_LOC_26/Y OR2X1_LOC_417/A 2.10fF
C38710 OR2X1_LOC_89/A OR2X1_LOC_417/A 0.30fF
C39407 OR2X1_LOC_417/A OR2X1_LOC_816/A 0.02fF
C39597 OR2X1_LOC_488/Y OR2X1_LOC_417/A 0.01fF
C39622 OR2X1_LOC_417/A OR2X1_LOC_95/Y 0.63fF
C40727 OR2X1_LOC_417/A OR2X1_LOC_59/Y 0.30fF
C40841 AND2X1_LOC_514/Y OR2X1_LOC_417/A 0.01fF
C41324 OR2X1_LOC_47/Y OR2X1_LOC_417/A 5.23fF
C41669 OR2X1_LOC_625/Y OR2X1_LOC_417/A 0.09fF
C42441 OR2X1_LOC_417/A OR2X1_LOC_16/A 0.03fF
C42859 OR2X1_LOC_417/A OR2X1_LOC_373/Y 0.03fF
C43925 OR2X1_LOC_417/A OR2X1_LOC_46/A 0.67fF
C44620 OR2X1_LOC_40/Y OR2X1_LOC_417/A 0.27fF
C44730 OR2X1_LOC_417/A OR2X1_LOC_7/A 0.45fF
C46045 OR2X1_LOC_43/A OR2X1_LOC_417/A 0.07fF
C46963 OR2X1_LOC_3/Y OR2X1_LOC_417/A 0.49fF
C47338 OR2X1_LOC_329/B OR2X1_LOC_417/A 0.14fF
C48326 OR2X1_LOC_64/Y OR2X1_LOC_417/A 3.41fF
C48744 OR2X1_LOC_417/A OR2X1_LOC_226/a_8_216# 0.06fF
C49087 OR2X1_LOC_283/a_8_216# OR2X1_LOC_417/A 0.01fF
C51163 OR2X1_LOC_628/a_8_216# OR2X1_LOC_417/A 0.14fF
C53737 OR2X1_LOC_417/A OR2X1_LOC_278/Y 0.04fF
C54877 OR2X1_LOC_369/a_8_216# OR2X1_LOC_417/A 0.09fF
C55418 OR2X1_LOC_36/Y OR2X1_LOC_417/A 0.15fF
C55776 OR2X1_LOC_604/A OR2X1_LOC_417/A 0.17fF
C56996 OR2X1_LOC_417/A VSS -3.77fF
C23 OR2X1_LOC_405/A OR2X1_LOC_121/B 0.11fF
C1931 OR2X1_LOC_121/B OR2X1_LOC_68/B 0.06fF
C2685 OR2X1_LOC_121/B OR2X1_LOC_87/A 0.23fF
C3095 OR2X1_LOC_121/B AND2X1_LOC_29/a_8_24# 0.05fF
C3480 OR2X1_LOC_121/B AND2X1_LOC_426/a_8_24# 0.03fF
C5127 OR2X1_LOC_154/A OR2X1_LOC_121/B 0.14fF
C5433 OR2X1_LOC_121/B AND2X1_LOC_299/a_8_24# 0.03fF
C6643 AND2X1_LOC_64/Y OR2X1_LOC_121/B 2.88fF
C6871 AND2X1_LOC_369/a_8_24# OR2X1_LOC_121/B 0.04fF
C7229 OR2X1_LOC_756/B OR2X1_LOC_121/B 0.03fF
C8486 OR2X1_LOC_49/A OR2X1_LOC_121/B 0.18fF
C8511 OR2X1_LOC_121/B OR2X1_LOC_596/A 2.49fF
C8642 OR2X1_LOC_121/B OR2X1_LOC_87/B 0.72fF
C8737 OR2X1_LOC_121/B OR2X1_LOC_374/Y 0.03fF
C8988 OR2X1_LOC_100/Y OR2X1_LOC_121/B 0.16fF
C9110 OR2X1_LOC_121/B OR2X1_LOC_532/B 0.30fF
C9930 AND2X1_LOC_42/B OR2X1_LOC_121/B 0.04fF
C10305 OR2X1_LOC_185/Y OR2X1_LOC_121/B 0.09fF
C11030 VDD OR2X1_LOC_121/B 0.60fF
C14130 OR2X1_LOC_160/A OR2X1_LOC_121/B 0.17fF
C14501 OR2X1_LOC_325/A OR2X1_LOC_121/B 0.01fF
C14601 AND2X1_LOC_46/a_8_24# OR2X1_LOC_121/B 0.01fF
C14731 OR2X1_LOC_121/B OR2X1_LOC_544/B 0.27fF
C15343 OR2X1_LOC_185/A OR2X1_LOC_121/B 1.76fF
C16217 OR2X1_LOC_264/a_8_216# OR2X1_LOC_121/B 0.01fF
C16535 OR2X1_LOC_121/B AND2X1_LOC_299/a_36_24# 0.01fF
C17439 OR2X1_LOC_264/Y OR2X1_LOC_121/B 1.38fF
C17718 AND2X1_LOC_91/B OR2X1_LOC_121/B 0.06fF
C18382 AND2X1_LOC_56/B OR2X1_LOC_121/B 0.10fF
C18390 AND2X1_LOC_8/Y OR2X1_LOC_121/B 0.46fF
C18732 OR2X1_LOC_121/B AND2X1_LOC_92/Y 0.10fF
C19532 OR2X1_LOC_6/B OR2X1_LOC_121/B 0.03fF
C19730 OR2X1_LOC_121/B AND2X1_LOC_47/Y 0.25fF
C20058 OR2X1_LOC_121/B OR2X1_LOC_506/A 0.47fF
C20476 AND2X1_LOC_95/Y OR2X1_LOC_121/B 0.04fF
C20765 AND2X1_LOC_22/Y OR2X1_LOC_121/B 0.07fF
C21942 OR2X1_LOC_121/B OR2X1_LOC_779/B 0.03fF
C22099 OR2X1_LOC_709/A OR2X1_LOC_121/B 0.07fF
C22160 AND2X1_LOC_70/Y OR2X1_LOC_121/B 0.09fF
C23312 OR2X1_LOC_121/B AND2X1_LOC_273/a_8_24# 0.01fF
C23772 OR2X1_LOC_121/B AND2X1_LOC_44/Y 0.18fF
C24648 OR2X1_LOC_121/B AND2X1_LOC_18/Y 1.53fF
C25570 OR2X1_LOC_121/B OR2X1_LOC_130/A 0.03fF
C25655 OR2X1_LOC_121/B OR2X1_LOC_780/B 0.17fF
C25668 OR2X1_LOC_121/B AND2X1_LOC_88/Y 0.03fF
C26014 AND2X1_LOC_88/a_8_24# OR2X1_LOC_121/B 0.01fF
C27669 OR2X1_LOC_121/B OR2X1_LOC_161/A 0.99fF
C27724 OR2X1_LOC_121/B AND2X1_LOC_51/Y 0.16fF
C27955 OR2X1_LOC_121/a_8_216# OR2X1_LOC_121/B 0.07fF
C28472 AND2X1_LOC_41/A OR2X1_LOC_121/B 0.11fF
C29928 OR2X1_LOC_121/B AND2X1_LOC_31/Y 0.10fF
C30463 OR2X1_LOC_121/B OR2X1_LOC_121/A 0.14fF
C30845 OR2X1_LOC_121/B AND2X1_LOC_36/Y 0.11fF
C31121 AND2X1_LOC_46/a_36_24# OR2X1_LOC_121/B 0.01fF
C33175 OR2X1_LOC_121/B OR2X1_LOC_269/B 0.10fF
C34181 OR2X1_LOC_121/B OR2X1_LOC_777/B 0.03fF
C34236 OR2X1_LOC_121/B OR2X1_LOC_831/B 0.01fF
C34699 OR2X1_LOC_121/B OR2X1_LOC_161/B 0.19fF
C36068 OR2X1_LOC_502/A OR2X1_LOC_121/B 0.07fF
C36171 AND2X1_LOC_48/A OR2X1_LOC_121/B 0.08fF
C36546 OR2X1_LOC_121/B AND2X1_LOC_3/Y 0.03fF
C37196 OR2X1_LOC_121/B AND2X1_LOC_7/B 0.16fF
C38305 OR2X1_LOC_473/A OR2X1_LOC_121/B 0.03fF
C38999 OR2X1_LOC_160/B OR2X1_LOC_121/B 0.10fF
C39494 OR2X1_LOC_327/a_8_216# OR2X1_LOC_121/B 0.01fF
C39824 OR2X1_LOC_151/A OR2X1_LOC_121/B 0.10fF
C39833 AND2X1_LOC_322/a_8_24# OR2X1_LOC_121/B 0.01fF
C42603 OR2X1_LOC_121/B OR2X1_LOC_606/a_36_216# 0.02fF
C42860 AND2X1_LOC_110/Y OR2X1_LOC_121/B 0.06fF
C43347 OR2X1_LOC_121/B OR2X1_LOC_448/A 0.11fF
C44599 OR2X1_LOC_121/B OR2X1_LOC_66/A 0.15fF
C45457 OR2X1_LOC_325/B OR2X1_LOC_121/B 0.01fF
C45864 OR2X1_LOC_831/A OR2X1_LOC_121/B 0.02fF
C45955 AND2X1_LOC_40/Y OR2X1_LOC_121/B 0.09fF
C46465 OR2X1_LOC_121/B AND2X1_LOC_43/B 0.07fF
C48319 OR2X1_LOC_121/B OR2X1_LOC_606/Y 0.04fF
C48561 AND2X1_LOC_323/a_8_24# OR2X1_LOC_121/B 0.01fF
C48990 OR2X1_LOC_121/B OR2X1_LOC_78/A 1.47fF
C49016 OR2X1_LOC_121/B OR2X1_LOC_448/B 0.03fF
C49073 OR2X1_LOC_121/B OR2X1_LOC_155/A 1.92fF
C49581 OR2X1_LOC_121/B OR2X1_LOC_814/A 0.10fF
C50350 AND2X1_LOC_12/Y OR2X1_LOC_121/B 8.95fF
C50715 OR2X1_LOC_168/B OR2X1_LOC_121/B 0.03fF
C50767 AND2X1_LOC_59/Y OR2X1_LOC_121/B 1.87fF
C53275 AND2X1_LOC_81/B OR2X1_LOC_121/B 0.05fF
C54093 OR2X1_LOC_377/A OR2X1_LOC_121/B 0.02fF
C54462 OR2X1_LOC_121/B OR2X1_LOC_78/B 0.05fF
C54522 OR2X1_LOC_121/B OR2X1_LOC_375/A 0.30fF
C55695 OR2X1_LOC_121/B AND2X1_LOC_65/A 0.03fF
C57184 OR2X1_LOC_121/B VSS 0.70fF
C1334 OR2X1_LOC_817/Y AND2X1_LOC_847/Y 0.05fF
C8059 VDD OR2X1_LOC_817/Y 0.12fF
C10714 OR2X1_LOC_817/Y OR2X1_LOC_44/Y 0.02fF
C11960 OR2X1_LOC_748/A OR2X1_LOC_817/Y 0.01fF
C20809 OR2X1_LOC_600/A OR2X1_LOC_817/Y 0.01fF
C30234 OR2X1_LOC_817/Y AND2X1_LOC_847/a_8_24# 0.23fF
C32754 OR2X1_LOC_3/Y OR2X1_LOC_817/Y 0.02fF
C54122 OR2X1_LOC_817/a_8_216# OR2X1_LOC_817/Y -0.00fF
C57360 OR2X1_LOC_817/Y VSS 0.06fF
C184 OR2X1_LOC_62/A AND2X1_LOC_14/a_8_24# 0.20fF
C610 OR2X1_LOC_62/A OR2X1_LOC_47/Y 3.63fF
C932 AND2X1_LOC_143/a_8_24# OR2X1_LOC_62/A 0.09fF
C1204 OR2X1_LOC_62/A AND2X1_LOC_36/Y 0.09fF
C1711 OR2X1_LOC_62/A OR2X1_LOC_16/A 0.23fF
C3182 OR2X1_LOC_62/A OR2X1_LOC_46/A 0.50fF
C5177 OR2X1_LOC_43/A OR2X1_LOC_62/A 0.18fF
C6117 OR2X1_LOC_62/A OR2X1_LOC_673/A 0.04fF
C6408 OR2X1_LOC_502/A OR2X1_LOC_62/A 0.31fF
C6530 OR2X1_LOC_62/A OR2X1_LOC_618/Y 0.12fF
C9098 OR2X1_LOC_287/B OR2X1_LOC_62/A 0.02fF
C10743 OR2X1_LOC_62/A AND2X1_LOC_619/B 0.03fF
C10794 AND2X1_LOC_102/a_36_24# OR2X1_LOC_62/A 0.01fF
C12890 OR2X1_LOC_62/A OR2X1_LOC_38/a_8_216# -0.03fF
C12961 OR2X1_LOC_62/A OR2X1_LOC_19/B 0.08fF
C17606 OR2X1_LOC_62/A OR2X1_LOC_619/a_8_216# 0.09fF
C17748 OR2X1_LOC_62/A AND2X1_LOC_619/a_8_24# 0.15fF
C19196 OR2X1_LOC_62/A OR2X1_LOC_78/A 0.02fF
C21444 OR2X1_LOC_62/A OR2X1_LOC_585/A 1.25fF
C22290 OR2X1_LOC_62/A OR2X1_LOC_753/A 0.20fF
C23060 OR2X1_LOC_8/Y OR2X1_LOC_62/A 0.06fF
C23366 OR2X1_LOC_62/A OR2X1_LOC_622/B 0.13fF
C23433 OR2X1_LOC_62/A OR2X1_LOC_9/a_8_216# 0.06fF
C24031 OR2X1_LOC_62/A AND2X1_LOC_672/B 0.04fF
C24355 OR2X1_LOC_377/A OR2X1_LOC_62/A 0.13fF
C24368 OR2X1_LOC_62/A OR2X1_LOC_85/A 3.25fF
C24784 OR2X1_LOC_62/A OR2X1_LOC_375/A 0.61fF
C26497 AND2X1_LOC_77/a_8_24# OR2X1_LOC_62/A 0.19fF
C27193 OR2X1_LOC_62/A AND2X1_LOC_277/a_8_24# 0.01fF
C28191 OR2X1_LOC_62/A AND2X1_LOC_4/a_8_24# 0.02fF
C28314 OR2X1_LOC_62/A OR2X1_LOC_68/B 2.41fF
C28794 OR2X1_LOC_62/A AND2X1_LOC_619/a_36_24# 0.01fF
C30305 OR2X1_LOC_62/A OR2X1_LOC_415/A 0.01fF
C32313 OR2X1_LOC_62/A OR2X1_LOC_94/a_8_216# 0.18fF
C32653 OR2X1_LOC_62/A OR2X1_LOC_633/A 0.09fF
C33024 OR2X1_LOC_696/A OR2X1_LOC_62/A 0.03fF
C33660 AND2X1_LOC_55/a_8_24# OR2X1_LOC_62/A 0.03fF
C34097 OR2X1_LOC_611/a_8_216# OR2X1_LOC_62/A 0.02fF
C34768 OR2X1_LOC_49/A OR2X1_LOC_62/A 0.51fF
C35191 OR2X1_LOC_671/Y OR2X1_LOC_62/A 0.09fF
C35351 OR2X1_LOC_62/A OR2X1_LOC_532/B 0.01fF
C36181 OR2X1_LOC_62/A AND2X1_LOC_42/B 0.78fF
C37328 VDD OR2X1_LOC_62/A 1.20fF
C39290 OR2X1_LOC_62/A OR2X1_LOC_80/A 0.09fF
C39578 OR2X1_LOC_62/A OR2X1_LOC_6/A 0.58fF
C39615 OR2X1_LOC_611/a_36_216# OR2X1_LOC_62/A 0.11fF
C40707 OR2X1_LOC_158/A OR2X1_LOC_62/A 0.08fF
C40776 OR2X1_LOC_62/A OR2X1_LOC_847/A 0.02fF
C43038 OR2X1_LOC_824/a_8_216# OR2X1_LOC_62/A 0.03fF
C44669 OR2X1_LOC_62/A OR2X1_LOC_56/A 0.10fF
C44709 OR2X1_LOC_62/A AND2X1_LOC_9/a_8_24# 0.01fF
C44739 AND2X1_LOC_8/Y OR2X1_LOC_62/A 1.05fF
C45945 OR2X1_LOC_6/B OR2X1_LOC_62/A 0.73fF
C46129 OR2X1_LOC_62/A AND2X1_LOC_47/Y 0.04fF
C46819 OR2X1_LOC_62/A OR2X1_LOC_15/a_8_216# 0.11fF
C46921 OR2X1_LOC_62/A AND2X1_LOC_414/a_8_24# 0.04fF
C48237 OR2X1_LOC_235/B OR2X1_LOC_62/A 0.18fF
C49097 OR2X1_LOC_62/A OR2X1_LOC_96/B 0.12fF
C50024 OR2X1_LOC_62/A OR2X1_LOC_62/a_8_216# 0.05fF
C50322 OR2X1_LOC_600/A OR2X1_LOC_62/A 0.07fF
C50390 OR2X1_LOC_62/A OR2X1_LOC_619/Y -0.01fF
C51290 OR2X1_LOC_62/A AND2X1_LOC_672/a_8_24# 0.02fF
C52101 OR2X1_LOC_62/A OR2X1_LOC_62/B 0.42fF
C53821 OR2X1_LOC_62/A OR2X1_LOC_54/Y 0.17fF
C54998 OR2X1_LOC_62/A OR2X1_LOC_824/Y 0.01fF
C55069 OR2X1_LOC_62/A OR2X1_LOC_95/Y 0.11fF
C55903 AND2X1_LOC_102/a_8_24# OR2X1_LOC_62/A 0.04fF
C56043 OR2X1_LOC_62/A OR2X1_LOC_71/A 0.24fF
C57256 OR2X1_LOC_62/A VSS 0.23fF
C63 AND2X1_LOC_53/Y AND2X1_LOC_43/B 1.01fF
C355 OR2X1_LOC_502/A AND2X1_LOC_43/B 0.26fF
C472 AND2X1_LOC_48/A AND2X1_LOC_43/B 0.13fF
C873 AND2X1_LOC_3/Y AND2X1_LOC_43/B 0.35fF
C1536 AND2X1_LOC_43/B AND2X1_LOC_7/B 0.37fF
C2750 AND2X1_LOC_43/B OR2X1_LOC_513/Y 0.02fF
C3326 OR2X1_LOC_160/B AND2X1_LOC_43/B 0.14fF
C4108 OR2X1_LOC_151/A AND2X1_LOC_43/B 4.32fF
C4497 AND2X1_LOC_300/a_8_24# AND2X1_LOC_43/B 0.04fF
C5274 AND2X1_LOC_43/B OR2X1_LOC_415/Y 0.08fF
C5482 AND2X1_LOC_43/B AND2X1_LOC_413/a_36_24# 0.01fF
C5510 AND2X1_LOC_43/B OR2X1_LOC_378/Y 0.06fF
C5637 AND2X1_LOC_43/B OR2X1_LOC_378/A 0.50fF
C6848 OR2X1_LOC_19/B AND2X1_LOC_43/B 0.18fF
C7057 AND2X1_LOC_534/a_8_24# AND2X1_LOC_43/B 0.22fF
C7097 AND2X1_LOC_110/Y AND2X1_LOC_43/B 0.02fF
C7837 AND2X1_LOC_43/B OR2X1_LOC_515/a_8_216# 0.01fF
C7927 AND2X1_LOC_43/B OR2X1_LOC_375/a_8_216# 0.04fF
C8848 AND2X1_LOC_43/B OR2X1_LOC_66/A 0.11fF
C9304 AND2X1_LOC_94/Y AND2X1_LOC_43/B 0.09fF
C9346 AND2X1_LOC_50/Y AND2X1_LOC_43/B 0.02fF
C9694 OR2X1_LOC_686/B AND2X1_LOC_43/B 0.01fF
C10090 OR2X1_LOC_831/A AND2X1_LOC_43/B 0.03fF
C10183 AND2X1_LOC_40/Y AND2X1_LOC_43/B 0.10fF
C11151 AND2X1_LOC_56/a_8_24# AND2X1_LOC_43/B 0.04fF
C12342 OR2X1_LOC_687/Y AND2X1_LOC_43/B 0.03fF
C12461 AND2X1_LOC_43/B AND2X1_LOC_827/a_36_24# 0.01fF
C12611 OR2X1_LOC_535/A AND2X1_LOC_43/B 0.05fF
C13143 AND2X1_LOC_43/B OR2X1_LOC_78/A 0.23fF
C13165 OR2X1_LOC_458/B AND2X1_LOC_43/B 0.12fF
C13248 AND2X1_LOC_43/B OR2X1_LOC_155/A 0.04fF
C13719 AND2X1_LOC_43/B OR2X1_LOC_814/A 0.07fF
C13945 AND2X1_LOC_43/B OR2X1_LOC_410/Y 0.03fF
C14110 AND2X1_LOC_387/B AND2X1_LOC_43/B 0.07fF
C14462 AND2X1_LOC_12/Y AND2X1_LOC_43/B 0.41fF
C14831 AND2X1_LOC_752/a_8_24# AND2X1_LOC_43/B 0.04fF
C14875 AND2X1_LOC_59/Y AND2X1_LOC_43/B 5.75fF
C15315 AND2X1_LOC_43/a_8_24# AND2X1_LOC_43/B 0.10fF
C16116 AND2X1_LOC_43/B AND2X1_LOC_272/a_8_24# 0.06fF
C16660 OR2X1_LOC_197/A AND2X1_LOC_43/B 0.05fF
C17492 AND2X1_LOC_692/a_8_24# AND2X1_LOC_43/B 0.04fF
C18132 AND2X1_LOC_534/a_36_24# AND2X1_LOC_43/B 0.01fF
C18263 OR2X1_LOC_377/A AND2X1_LOC_43/B 0.24fF
C18633 AND2X1_LOC_43/B OR2X1_LOC_78/B 0.11fF
C18720 OR2X1_LOC_375/A AND2X1_LOC_43/B 0.54fF
C18904 AND2X1_LOC_43/B OR2X1_LOC_515/Y 0.20fF
C18995 AND2X1_LOC_43/B OR2X1_LOC_549/A 0.07fF
C19444 AND2X1_LOC_43/B AND2X1_LOC_411/a_8_24# 0.05fF
C20377 AND2X1_LOC_753/B AND2X1_LOC_43/B 0.91fF
C20401 OR2X1_LOC_405/A AND2X1_LOC_43/B 0.12fF
C20906 OR2X1_LOC_195/A AND2X1_LOC_43/B 0.14fF
C21161 AND2X1_LOC_300/a_36_24# AND2X1_LOC_43/B 0.01fF
C21991 AND2X1_LOC_43/B OR2X1_LOC_138/A 0.01fF
C22256 AND2X1_LOC_56/a_36_24# AND2X1_LOC_43/B 0.01fF
C22319 AND2X1_LOC_43/B OR2X1_LOC_68/B 6.42fF
C22956 OR2X1_LOC_459/A AND2X1_LOC_43/B 0.07fF
C23035 OR2X1_LOC_87/A AND2X1_LOC_43/B 0.10fF
C24202 OR2X1_LOC_541/A AND2X1_LOC_43/B 0.03fF
C24500 AND2X1_LOC_43/B OR2X1_LOC_375/Y 0.01fF
C25496 OR2X1_LOC_154/A AND2X1_LOC_43/B 3.15fF
C25621 AND2X1_LOC_684/a_8_24# AND2X1_LOC_43/B 0.06fF
C26143 AND2X1_LOC_43/B AND2X1_LOC_409/B 0.07fF
C26256 OR2X1_LOC_634/A AND2X1_LOC_43/B 0.11fF
C26354 AND2X1_LOC_43/a_36_24# AND2X1_LOC_43/B 0.01fF
C26986 AND2X1_LOC_64/Y AND2X1_LOC_43/B 0.26fF
C27513 OR2X1_LOC_756/B AND2X1_LOC_43/B 0.42fF
C28541 AND2X1_LOC_692/a_36_24# AND2X1_LOC_43/B 0.01fF
C28707 OR2X1_LOC_49/A AND2X1_LOC_43/B 0.07fF
C28728 AND2X1_LOC_43/B OR2X1_LOC_596/A 0.11fF
C29382 OR2X1_LOC_532/B AND2X1_LOC_43/B 0.05fF
C30178 AND2X1_LOC_42/B AND2X1_LOC_43/B 0.20fF
C30442 AND2X1_LOC_43/B AND2X1_LOC_411/a_36_24# 0.01fF
C30548 OR2X1_LOC_185/Y AND2X1_LOC_43/B 0.45fF
C30952 AND2X1_LOC_53/a_8_24# AND2X1_LOC_43/B 0.03fF
C31306 VDD AND2X1_LOC_43/B 1.38fF
C33253 AND2X1_LOC_43/B OR2X1_LOC_80/A 0.01fF
C33264 AND2X1_LOC_43/B AND2X1_LOC_419/a_8_24# 0.04fF
C34304 OR2X1_LOC_160/A AND2X1_LOC_43/B 0.02fF
C35426 AND2X1_LOC_92/a_8_24# AND2X1_LOC_43/B 0.04fF
C35593 OR2X1_LOC_185/A AND2X1_LOC_43/B 0.03fF
C36816 AND2X1_LOC_753/a_8_24# AND2X1_LOC_43/B 0.05fF
C37942 AND2X1_LOC_91/B AND2X1_LOC_43/B 0.07fF
C38310 AND2X1_LOC_43/B OR2X1_LOC_446/B 0.75fF
C38569 AND2X1_LOC_56/B AND2X1_LOC_43/B 0.12fF
C38585 AND2X1_LOC_8/Y AND2X1_LOC_43/B 0.07fF
C38926 AND2X1_LOC_43/B AND2X1_LOC_92/Y 0.13fF
C39463 OR2X1_LOC_83/A AND2X1_LOC_43/B 0.01fF
C39735 OR2X1_LOC_6/B AND2X1_LOC_43/B 0.07fF
C39945 AND2X1_LOC_47/Y AND2X1_LOC_43/B 0.19fF
C40215 OR2X1_LOC_506/A AND2X1_LOC_43/B 0.15fF
C40665 AND2X1_LOC_95/Y AND2X1_LOC_43/B 0.14fF
C40935 AND2X1_LOC_22/Y AND2X1_LOC_43/B 0.42fF
C41055 OR2X1_LOC_706/A AND2X1_LOC_43/B 0.03fF
C41918 OR2X1_LOC_638/B AND2X1_LOC_43/B 0.02fF
C42120 OR2X1_LOC_276/B AND2X1_LOC_43/B 0.07fF
C42297 OR2X1_LOC_709/A AND2X1_LOC_43/B 0.02fF
C42343 AND2X1_LOC_70/Y AND2X1_LOC_43/B 0.22fF
C44005 AND2X1_LOC_43/B AND2X1_LOC_44/Y 0.08fF
C44028 AND2X1_LOC_43/B OR2X1_LOC_514/a_8_216# 0.01fF
C44922 AND2X1_LOC_43/B AND2X1_LOC_18/Y 0.10fF
C45058 AND2X1_LOC_43/B AND2X1_LOC_413/a_8_24# 0.05fF
C48154 AND2X1_LOC_43/B OR2X1_LOC_161/A 0.22fF
C48229 AND2X1_LOC_43/B AND2X1_LOC_51/Y 0.21fF
C48919 AND2X1_LOC_41/A AND2X1_LOC_43/B 0.40fF
C49472 AND2X1_LOC_136/a_8_24# AND2X1_LOC_43/B 0.01fF
C50025 AND2X1_LOC_43/B AND2X1_LOC_419/a_36_24# 0.01fF
C50439 AND2X1_LOC_31/Y AND2X1_LOC_43/B 0.38fF
C50937 AND2X1_LOC_43/B OR2X1_LOC_121/A 0.03fF
C51292 AND2X1_LOC_43/B AND2X1_LOC_36/Y 0.19fF
C52041 AND2X1_LOC_43/B AND2X1_LOC_827/a_8_24# 0.01fF
C52181 AND2X1_LOC_92/a_36_24# AND2X1_LOC_43/B 0.01fF
C53276 AND2X1_LOC_43/B OR2X1_LOC_46/A 12.07fF
C53631 AND2X1_LOC_753/a_36_24# AND2X1_LOC_43/B 0.01fF
C53675 AND2X1_LOC_43/B OR2X1_LOC_269/B 2.72fF
C54598 AND2X1_LOC_43/B OR2X1_LOC_378/a_8_216# 0.08fF
C55145 AND2X1_LOC_43/B OR2X1_LOC_161/B 8.08fF
C55177 AND2X1_LOC_43/B OR2X1_LOC_514/a_36_216# 0.02fF
C56837 AND2X1_LOC_43/B VSS -4.45fF
C1047 AND2X1_LOC_92/Y OR2X1_LOC_120/a_8_216# 0.05fF
C1086 OR2X1_LOC_596/A AND2X1_LOC_92/Y 0.03fF
C1228 OR2X1_LOC_87/B AND2X1_LOC_92/Y 0.03fF
C1749 OR2X1_LOC_532/B AND2X1_LOC_92/Y 0.14fF
C2566 AND2X1_LOC_42/B AND2X1_LOC_92/Y 0.15fF
C2952 OR2X1_LOC_185/Y AND2X1_LOC_92/Y 0.53fF
C3671 VDD AND2X1_LOC_92/Y 1.85fF
C6435 AND2X1_LOC_92/Y OR2X1_LOC_750/Y 0.10fF
C6668 OR2X1_LOC_160/A AND2X1_LOC_92/Y 0.17fF
C7847 AND2X1_LOC_92/a_8_24# AND2X1_LOC_92/Y 0.01fF
C8001 OR2X1_LOC_185/A AND2X1_LOC_92/Y 0.11fF
C9722 OR2X1_LOC_541/B AND2X1_LOC_92/Y 0.02fF
C10422 AND2X1_LOC_91/B AND2X1_LOC_92/Y 0.20fF
C10974 AND2X1_LOC_56/B AND2X1_LOC_92/Y 1.27fF
C10987 AND2X1_LOC_8/Y AND2X1_LOC_92/Y 2.07fF
C12139 OR2X1_LOC_6/B AND2X1_LOC_92/Y 0.01fF
C12377 AND2X1_LOC_47/Y AND2X1_LOC_92/Y 0.26fF
C12666 OR2X1_LOC_506/A AND2X1_LOC_92/Y 0.03fF
C13124 AND2X1_LOC_95/Y AND2X1_LOC_92/Y 0.22fF
C13422 AND2X1_LOC_22/Y AND2X1_LOC_92/Y 0.17fF
C13544 AND2X1_LOC_153/a_8_24# AND2X1_LOC_92/Y 0.06fF
C14520 OR2X1_LOC_276/B AND2X1_LOC_92/Y 0.02fF
C14687 OR2X1_LOC_709/A AND2X1_LOC_92/Y 0.07fF
C14725 AND2X1_LOC_70/Y AND2X1_LOC_92/Y 0.07fF
C15880 AND2X1_LOC_273/a_8_24# AND2X1_LOC_92/Y 0.06fF
C15911 AND2X1_LOC_92/Y AND2X1_LOC_256/a_8_24# 0.01fF
C16325 AND2X1_LOC_92/Y AND2X1_LOC_44/Y 1.81fF
C16833 AND2X1_LOC_92/Y AND2X1_LOC_628/a_8_24# 0.02fF
C17246 AND2X1_LOC_18/Y AND2X1_LOC_92/Y 0.17fF
C18198 OR2X1_LOC_130/A AND2X1_LOC_92/Y 0.18fF
C20318 OR2X1_LOC_161/A AND2X1_LOC_92/Y 9.54fF
C20417 AND2X1_LOC_51/Y AND2X1_LOC_92/Y 0.13fF
C21134 AND2X1_LOC_41/A AND2X1_LOC_92/Y 0.33fF
C22721 AND2X1_LOC_31/Y AND2X1_LOC_92/Y 0.10fF
C22982 AND2X1_LOC_92/Y OR2X1_LOC_240/A 0.82fF
C23206 AND2X1_LOC_92/Y OR2X1_LOC_121/A 0.03fF
C23579 AND2X1_LOC_92/Y AND2X1_LOC_36/Y 0.08fF
C25509 OR2X1_LOC_46/A AND2X1_LOC_92/Y 0.03fF
C25845 AND2X1_LOC_92/Y OR2X1_LOC_269/B 0.13fF
C26902 AND2X1_LOC_92/Y OR2X1_LOC_777/B 0.10fF
C26945 OR2X1_LOC_831/B AND2X1_LOC_92/Y 5.64fF
C26968 AND2X1_LOC_92/Y OR2X1_LOC_344/A 0.01fF
C27386 AND2X1_LOC_92/Y OR2X1_LOC_161/B 0.07fF
C27868 AND2X1_LOC_92/Y OR2X1_LOC_630/B 0.01fF
C28733 OR2X1_LOC_502/A AND2X1_LOC_92/Y 0.14fF
C28875 AND2X1_LOC_48/A AND2X1_LOC_92/Y 0.07fF
C29245 AND2X1_LOC_3/Y AND2X1_LOC_92/Y 0.07fF
C29907 AND2X1_LOC_7/B AND2X1_LOC_92/Y 0.29fF
C30417 AND2X1_LOC_372/a_8_24# AND2X1_LOC_92/Y 0.03fF
C31646 OR2X1_LOC_160/B AND2X1_LOC_92/Y 0.11fF
C32436 OR2X1_LOC_151/A AND2X1_LOC_92/Y 0.17fF
C35403 AND2X1_LOC_110/Y AND2X1_LOC_92/Y 0.03fF
C37108 AND2X1_LOC_92/Y OR2X1_LOC_66/A 0.09fF
C37929 AND2X1_LOC_93/a_8_24# AND2X1_LOC_92/Y 0.11fF
C38034 OR2X1_LOC_405/Y AND2X1_LOC_92/Y 0.04fF
C38351 OR2X1_LOC_831/A AND2X1_LOC_92/Y 0.07fF
C38432 AND2X1_LOC_40/Y AND2X1_LOC_92/Y 0.10fF
C39880 AND2X1_LOC_519/a_8_24# AND2X1_LOC_92/Y 0.01fF
C41397 OR2X1_LOC_78/A AND2X1_LOC_92/Y 0.14fF
C41523 OR2X1_LOC_155/A AND2X1_LOC_92/Y 0.20fF
C42027 OR2X1_LOC_814/A AND2X1_LOC_92/Y 0.26fF
C42797 AND2X1_LOC_12/Y AND2X1_LOC_92/Y 0.14fF
C43159 OR2X1_LOC_168/B AND2X1_LOC_92/Y 0.08fF
C43218 AND2X1_LOC_59/Y AND2X1_LOC_92/Y 0.31fF
C45507 OR2X1_LOC_520/A AND2X1_LOC_92/Y 0.01fF
C46177 AND2X1_LOC_387/a_8_24# AND2X1_LOC_92/Y 0.08fF
C46728 OR2X1_LOC_377/A AND2X1_LOC_92/Y 0.04fF
C47119 OR2X1_LOC_78/B AND2X1_LOC_92/Y 0.17fF
C47198 OR2X1_LOC_375/A AND2X1_LOC_92/Y 0.09fF
C47525 AND2X1_LOC_92/Y OR2X1_LOC_549/A 0.05fF
C48884 OR2X1_LOC_405/A AND2X1_LOC_92/Y 0.20fF
C49234 AND2X1_LOC_19/Y AND2X1_LOC_92/Y 0.12fF
C50813 AND2X1_LOC_92/Y OR2X1_LOC_68/B 0.10fF
C51440 OR2X1_LOC_87/A AND2X1_LOC_92/Y 0.09fF
C51771 OR2X1_LOC_389/A AND2X1_LOC_92/Y 0.06fF
C51825 AND2X1_LOC_422/a_8_24# AND2X1_LOC_92/Y 0.04fF
C52632 OR2X1_LOC_541/A AND2X1_LOC_92/Y 0.03fF
C53964 OR2X1_LOC_154/A AND2X1_LOC_92/Y 0.37fF
C54723 OR2X1_LOC_634/A AND2X1_LOC_92/Y 0.02fF
C55496 AND2X1_LOC_64/Y AND2X1_LOC_92/Y 0.19fF
C56035 OR2X1_LOC_756/B AND2X1_LOC_92/Y 0.10fF
C56580 AND2X1_LOC_92/Y VSS 0.47fF
C112 OR2X1_LOC_696/A OR2X1_LOC_6/B 0.07fF
C238 OR2X1_LOC_696/A OR2X1_LOC_529/Y 0.03fF
C687 OR2X1_LOC_696/A OR2X1_LOC_481/A 0.02fF
C731 OR2X1_LOC_696/A OR2X1_LOC_71/Y 0.04fF
C991 OR2X1_LOC_696/A OR2X1_LOC_585/a_8_216# 0.02fF
C1034 OR2X1_LOC_696/A OR2X1_LOC_426/B 0.17fF
C1192 OR2X1_LOC_696/A OR2X1_LOC_225/a_8_216# 0.01fF
C1221 OR2X1_LOC_696/A OR2X1_LOC_409/B 0.05fF
C1492 OR2X1_LOC_696/A AND2X1_LOC_374/a_8_24# 0.02fF
C2332 OR2X1_LOC_696/A OR2X1_LOC_235/B 0.79fF
C3103 OR2X1_LOC_696/A OR2X1_LOC_387/A 0.02fF
C4043 OR2X1_LOC_696/A OR2X1_LOC_92/Y 14.46fF
C4055 OR2X1_LOC_696/A AND2X1_LOC_801/a_36_24# 0.01fF
C4379 OR2X1_LOC_696/A OR2X1_LOC_600/A 10.88fF
C4430 OR2X1_LOC_696/A OR2X1_LOC_619/Y 0.15fF
C4875 OR2X1_LOC_696/A AND2X1_LOC_818/a_8_24# 0.06fF
C6216 OR2X1_LOC_696/A OR2X1_LOC_62/B 0.01fF
C6828 OR2X1_LOC_696/A OR2X1_LOC_13/B 1.19fF
C6889 OR2X1_LOC_696/A OR2X1_LOC_111/a_8_216# 0.01fF
C7344 OR2X1_LOC_696/A OR2X1_LOC_428/A 0.50fF
C7987 OR2X1_LOC_696/A OR2X1_LOC_54/Y 0.14fF
C8381 OR2X1_LOC_696/A OR2X1_LOC_26/Y 2.03fF
C8394 OR2X1_LOC_696/A OR2X1_LOC_89/A 0.28fF
C8761 OR2X1_LOC_696/A OR2X1_LOC_306/a_8_216# 0.09fF
C8916 OR2X1_LOC_696/A OR2X1_LOC_588/A 0.04fF
C9200 OR2X1_LOC_696/A OR2X1_LOC_824/Y 0.16fF
C9327 OR2X1_LOC_696/A OR2X1_LOC_95/Y 1.22fF
C9334 OR2X1_LOC_696/A OR2X1_LOC_368/A 0.01fF
C10408 OR2X1_LOC_696/A OR2X1_LOC_59/Y 0.04fF
C10478 OR2X1_LOC_696/A OR2X1_LOC_820/B 0.04fF
C10500 OR2X1_LOC_696/A OR2X1_LOC_70/Y 0.05fF
C10525 OR2X1_LOC_696/A AND2X1_LOC_514/Y 0.07fF
C10647 OR2X1_LOC_696/A OR2X1_LOC_70/A 0.02fF
C10991 OR2X1_LOC_696/A OR2X1_LOC_47/Y 0.26fF
C11261 OR2X1_LOC_696/A OR2X1_LOC_625/Y 0.07fF
C12035 OR2X1_LOC_696/A OR2X1_LOC_16/A 4.44fF
C12247 OR2X1_LOC_696/A OR2X1_LOC_225/a_36_216# -0.00fF
C12941 OR2X1_LOC_696/A OR2X1_LOC_93/Y 0.01fF
C13089 OR2X1_LOC_696/A AND2X1_LOC_729/B 0.08fF
C13521 OR2X1_LOC_696/A OR2X1_LOC_46/A 0.03fF
C13875 OR2X1_LOC_696/A OR2X1_LOC_599/A 0.12fF
C13889 OR2X1_LOC_696/A OR2X1_LOC_93/a_8_216# 0.01fF
C14214 OR2X1_LOC_696/A OR2X1_LOC_40/Y 0.16fF
C14281 OR2X1_LOC_696/A OR2X1_LOC_618/a_8_216# 0.01fF
C14307 OR2X1_LOC_696/A OR2X1_LOC_7/A 0.36fF
C15421 OR2X1_LOC_696/A OR2X1_LOC_589/A 0.36fF
C15424 OR2X1_LOC_696/A OR2X1_LOC_322/Y 0.16fF
C15530 OR2X1_LOC_696/A OR2X1_LOC_43/A 0.61fF
C15869 OR2X1_LOC_696/A OR2X1_LOC_585/Y 0.04fF
C16383 OR2X1_LOC_696/A OR2X1_LOC_3/Y 0.56fF
C16740 OR2X1_LOC_696/A OR2X1_LOC_329/B 0.21fF
C16959 OR2X1_LOC_696/A OR2X1_LOC_618/Y 0.01fF
C17620 OR2X1_LOC_696/A OR2X1_LOC_11/Y 0.05fF
C17688 OR2X1_LOC_696/A OR2X1_LOC_64/Y 0.41fF
C18187 OR2X1_LOC_696/A OR2X1_LOC_226/a_8_216# 0.04fF
C18895 OR2X1_LOC_696/A OR2X1_LOC_25/Y 0.01fF
C19294 OR2X1_LOC_696/A OR2X1_LOC_421/A 0.07fF
C19401 OR2X1_LOC_696/A AND2X1_LOC_512/a_8_24# 0.02fF
C21035 OR2X1_LOC_696/A OR2X1_LOC_517/A 0.03fF
C21525 OR2X1_LOC_696/A AND2X1_LOC_62/a_8_24# 0.01fF
C21545 OR2X1_LOC_696/A OR2X1_LOC_752/a_8_216# 0.03fF
C21859 OR2X1_LOC_696/A OR2X1_LOC_323/a_8_216# 0.01fF
C23220 OR2X1_LOC_696/A OR2X1_LOC_278/Y 0.03fF
C23240 OR2X1_LOC_696/A OR2X1_LOC_95/a_8_216# 0.02fF
C24373 OR2X1_LOC_696/A AND2X1_LOC_407/a_8_24# 0.04fF
C24905 OR2X1_LOC_696/A OR2X1_LOC_36/Y 0.30fF
C25062 OR2X1_LOC_696/A OR2X1_LOC_419/Y 0.02fF
C25236 OR2X1_LOC_696/A OR2X1_LOC_604/A 0.29fF
C26544 OR2X1_LOC_696/A AND2X1_LOC_375/a_8_24# 0.08fF
C27977 OR2X1_LOC_696/A OR2X1_LOC_619/a_8_216# 0.01fF
C28584 OR2X1_LOC_696/A OR2X1_LOC_12/Y 0.72fF
C28764 OR2X1_LOC_696/A AND2X1_LOC_801/B 0.01fF
C29053 OR2X1_LOC_696/A OR2X1_LOC_59/a_8_216# 0.01fF
C29198 OR2X1_LOC_696/A OR2X1_LOC_226/a_36_216# -0.00fF
C30335 OR2X1_LOC_696/A OR2X1_LOC_256/Y 0.12fF
C31202 OR2X1_LOC_696/A OR2X1_LOC_18/Y 4.93fF
C31660 OR2X1_LOC_696/A OR2X1_LOC_585/A 0.89fF
C32251 OR2X1_LOC_696/A OR2X1_LOC_437/A 0.41fF
C32454 OR2X1_LOC_696/A OR2X1_LOC_753/A 0.10fF
C32792 OR2X1_LOC_696/A OR2X1_LOC_323/Y 0.29fF
C33251 OR2X1_LOC_696/A OR2X1_LOC_8/Y 0.03fF
C33300 OR2X1_LOC_696/A OR2X1_LOC_67/A 0.03fF
C33322 OR2X1_LOC_696/A AND2X1_LOC_374/Y 0.01fF
C33329 OR2X1_LOC_696/A OR2X1_LOC_52/B 0.14fF
C33330 OR2X1_LOC_696/A OR2X1_LOC_672/Y 0.04fF
C33841 OR2X1_LOC_696/A OR2X1_LOC_22/Y 0.59fF
C33940 OR2X1_LOC_696/A OR2X1_LOC_387/a_8_216# 0.01fF
C34148 OR2X1_LOC_696/A OR2X1_LOC_39/A 1.36fF
C34563 OR2X1_LOC_696/A OR2X1_LOC_85/A 0.06fF
C34680 OR2X1_LOC_696/A OR2X1_LOC_226/Y 0.21fF
C34968 OR2X1_LOC_696/A OR2X1_LOC_51/Y 0.21fF
C36414 OR2X1_LOC_696/A OR2X1_LOC_599/Y 0.10fF
C36686 OR2X1_LOC_696/A OR2X1_LOC_387/Y 0.01fF
C37095 OR2X1_LOC_696/A OR2X1_LOC_511/Y 0.07fF
C37512 OR2X1_LOC_696/A OR2X1_LOC_376/A 0.20fF
C37878 OR2X1_LOC_696/A OR2X1_LOC_91/A 0.22fF
C38399 OR2X1_LOC_696/A OR2X1_LOC_371/Y 0.07fF
C38861 OR2X1_LOC_696/A OR2X1_LOC_74/A 0.76fF
C41875 OR2X1_LOC_696/A OR2X1_LOC_696/Y 0.03fF
C42730 OR2X1_LOC_696/A OR2X1_LOC_485/A 0.27fF
C45182 OR2X1_LOC_696/A OR2X1_LOC_49/A 0.02fF
C45227 OR2X1_LOC_696/A OR2X1_LOC_310/Y 0.03fF
C45270 OR2X1_LOC_696/A OR2X1_LOC_433/Y 0.02fF
C46559 OR2X1_LOC_696/A OR2X1_LOC_369/Y -0.01fF
C46603 OR2X1_LOC_696/A OR2X1_LOC_53/a_8_216# 0.05fF
C47295 OR2X1_LOC_696/A OR2X1_LOC_761/a_8_216# 0.04fF
C47884 OR2X1_LOC_696/A VDD 1.03fF
C48420 OR2X1_LOC_696/A OR2X1_LOC_6/a_8_216# 0.01fF
C48754 OR2X1_LOC_696/A OR2X1_LOC_382/Y 0.02fF
C49187 OR2X1_LOC_696/A OR2X1_LOC_427/A 0.91fF
C49191 OR2X1_LOC_696/A AND2X1_LOC_801/a_8_24# -0.07fF
C49571 OR2X1_LOC_696/A OR2X1_LOC_322/a_8_216# 0.05fF
C50081 OR2X1_LOC_696/A OR2X1_LOC_6/A 0.17fF
C50493 OR2X1_LOC_696/A OR2X1_LOC_44/Y 0.66fF
C50823 OR2X1_LOC_45/B OR2X1_LOC_696/A 0.12fF
C51233 OR2X1_LOC_696/A OR2X1_LOC_158/A 0.32fF
C52705 OR2X1_LOC_696/A OR2X1_LOC_111/Y 0.07fF
C52807 OR2X1_LOC_696/A OR2X1_LOC_588/a_8_216# 0.07fF
C53428 OR2X1_LOC_696/A OR2X1_LOC_529/a_8_216# 0.03fF
C53491 OR2X1_LOC_696/A OR2X1_LOC_824/a_8_216# 0.01fF
C53825 OR2X1_LOC_696/A OR2X1_LOC_744/A 0.87fF
C53961 OR2X1_LOC_696/A OR2X1_LOC_31/Y 0.56fF
C54670 OR2X1_LOC_696/A AND2X1_LOC_809/A 0.02fF
C55038 OR2X1_LOC_696/A OR2X1_LOC_56/A 13.19fF
C55089 OR2X1_LOC_696/A AND2X1_LOC_9/a_8_24# 0.01fF
C55602 OR2X1_LOC_696/A OR2X1_LOC_417/Y 0.07fF
C56019 OR2X1_LOC_696/A OR2X1_LOC_696/a_8_216# 0.07fF
C58100 OR2X1_LOC_696/A VSS -7.03fF
C7411 AND2X1_LOC_672/B OR2X1_LOC_673/A 0.02fF
C7695 OR2X1_LOC_502/A AND2X1_LOC_672/B 0.03fF
C14207 OR2X1_LOC_19/B AND2X1_LOC_672/B 0.02fF
C23534 AND2X1_LOC_672/B OR2X1_LOC_753/A 0.04fF
C29525 AND2X1_LOC_672/B OR2X1_LOC_68/B 0.03fF
C35976 OR2X1_LOC_49/A AND2X1_LOC_672/B 0.08fF
C38559 VDD AND2X1_LOC_672/B 0.16fF
C46035 AND2X1_LOC_8/Y AND2X1_LOC_672/B 0.90fF
C48224 AND2X1_LOC_672/B AND2X1_LOC_414/a_8_24# 0.01fF
C49447 OR2X1_LOC_235/B AND2X1_LOC_672/B 0.01fF
C52539 AND2X1_LOC_672/B AND2X1_LOC_672/a_8_24# 0.11fF
C53345 AND2X1_LOC_672/B OR2X1_LOC_62/B 0.42fF
C55012 AND2X1_LOC_672/B OR2X1_LOC_54/Y 0.03fF
C57217 AND2X1_LOC_672/B VSS 0.19fF
C3572 OR2X1_LOC_62/B OR2X1_LOC_415/A 0.01fF
C7472 OR2X1_LOC_415/A OR2X1_LOC_71/A 0.01fF
C14106 OR2X1_LOC_502/A OR2X1_LOC_415/A 0.01fF
C20571 OR2X1_LOC_19/B OR2X1_LOC_415/A 0.83fF
C29804 OR2X1_LOC_415/A OR2X1_LOC_753/A 0.60fF
C47074 OR2X1_LOC_415/A OR2X1_LOC_80/A 0.07fF
C52453 AND2X1_LOC_8/Y OR2X1_LOC_415/A 0.04fF
C57107 OR2X1_LOC_415/A VSS 0.13fF
C1363 OR2X1_LOC_18/Y OR2X1_LOC_46/A 0.04fF
C1813 OR2X1_LOC_585/A OR2X1_LOC_46/A 0.27fF
C2423 OR2X1_LOC_46/A OR2X1_LOC_437/A 0.07fF
C2610 OR2X1_LOC_411/Y OR2X1_LOC_46/A 0.01fF
C2695 OR2X1_LOC_46/A OR2X1_LOC_753/A 0.18fF
C3431 OR2X1_LOC_8/Y OR2X1_LOC_46/A 0.23fF
C3535 OR2X1_LOC_46/A OR2X1_LOC_52/B 0.03fF
C3536 OR2X1_LOC_672/Y OR2X1_LOC_46/A 0.01fF
C3804 OR2X1_LOC_46/A OR2X1_LOC_9/a_8_216# 0.01fF
C3994 OR2X1_LOC_22/Y OR2X1_LOC_46/A 0.05fF
C4305 OR2X1_LOC_46/A OR2X1_LOC_39/A 0.19fF
C4712 OR2X1_LOC_377/A OR2X1_LOC_46/A 0.14fF
C4730 OR2X1_LOC_85/A OR2X1_LOC_46/A 1.17fF
C5051 OR2X1_LOC_51/Y OR2X1_LOC_46/A 0.01fF
C5132 OR2X1_LOC_375/A OR2X1_LOC_46/A 0.07fF
C5908 OR2X1_LOC_46/A AND2X1_LOC_411/a_8_24# 0.04fF
C6506 OR2X1_LOC_599/Y OR2X1_LOC_46/A 0.06fF
C6854 OR2X1_LOC_413/Y OR2X1_LOC_46/A 0.01fF
C6952 OR2X1_LOC_416/A OR2X1_LOC_46/A 0.26fF
C7282 OR2X1_LOC_414/a_8_216# OR2X1_LOC_46/A 0.01fF
C8111 OR2X1_LOC_91/A OR2X1_LOC_46/A 0.11fF
C8630 OR2X1_LOC_32/B OR2X1_LOC_46/A 0.51fF
C8674 OR2X1_LOC_233/a_8_216# OR2X1_LOC_46/A 0.01fF
C8771 OR2X1_LOC_46/A OR2X1_LOC_68/B 0.03fF
C9069 OR2X1_LOC_74/A OR2X1_LOC_46/A 0.01fF
C9869 OR2X1_LOC_46/A OR2X1_LOC_23/a_8_216# 0.01fF
C10748 OR2X1_LOC_699/a_8_216# OR2X1_LOC_46/A 0.01fF
C11479 OR2X1_LOC_46/A OR2X1_LOC_461/B 0.03fF
C12806 OR2X1_LOC_634/A OR2X1_LOC_46/A 0.35fF
C12851 OR2X1_LOC_94/a_8_216# OR2X1_LOC_46/A 0.03fF
C12897 OR2X1_LOC_485/A OR2X1_LOC_46/A 0.02fF
C13324 OR2X1_LOC_827/Y OR2X1_LOC_46/A 0.01fF
C13788 OR2X1_LOC_54/a_8_216# OR2X1_LOC_46/A 0.01fF
C14996 OR2X1_LOC_82/a_8_216# OR2X1_LOC_46/A 0.01fF
C15054 OR2X1_LOC_80/a_8_216# OR2X1_LOC_46/A 0.02fF
C15226 OR2X1_LOC_49/A OR2X1_LOC_46/A 0.38fF
C15661 OR2X1_LOC_671/Y OR2X1_LOC_46/A 0.06fF
C15787 OR2X1_LOC_42/a_8_216# OR2X1_LOC_46/A 0.01fF
C17098 OR2X1_LOC_46/A AND2X1_LOC_412/a_8_24# 0.02fF
C17808 VDD OR2X1_LOC_46/A 1.61fF
C19199 OR2X1_LOC_427/A OR2X1_LOC_46/A 0.27fF
C19818 OR2X1_LOC_46/A OR2X1_LOC_80/A 0.56fF
C20093 OR2X1_LOC_46/A OR2X1_LOC_6/A 0.16fF
C20200 OR2X1_LOC_289/a_8_216# OR2X1_LOC_46/A 0.01fF
C20528 OR2X1_LOC_46/A OR2X1_LOC_44/Y 0.03fF
C20786 OR2X1_LOC_45/B OR2X1_LOC_46/A 0.24fF
C20849 AND2X1_LOC_410/a_8_24# OR2X1_LOC_46/A 0.01fF
C21254 OR2X1_LOC_158/A OR2X1_LOC_46/A 0.25fF
C22087 AND2X1_LOC_92/a_8_24# OR2X1_LOC_46/A 0.03fF
C22782 OR2X1_LOC_111/Y OR2X1_LOC_46/A 0.18fF
C22791 OR2X1_LOC_411/a_8_216# OR2X1_LOC_46/A 0.01fF
C23867 OR2X1_LOC_744/A OR2X1_LOC_46/A 0.15fF
C24018 OR2X1_LOC_31/Y OR2X1_LOC_46/A 0.77fF
C24258 OR2X1_LOC_129/a_8_216# OR2X1_LOC_46/A 0.01fF
C25094 OR2X1_LOC_46/A OR2X1_LOC_56/A 0.49fF
C25174 AND2X1_LOC_56/B OR2X1_LOC_46/A 0.48fF
C25203 OR2X1_LOC_291/A OR2X1_LOC_46/A 0.15fF
C25643 OR2X1_LOC_291/Y OR2X1_LOC_46/A 0.17fF
C26009 OR2X1_LOC_83/A OR2X1_LOC_46/A 0.03fF
C26300 OR2X1_LOC_6/B OR2X1_LOC_46/A 0.30fF
C26503 AND2X1_LOC_47/Y OR2X1_LOC_46/A 0.03fF
C26724 OR2X1_LOC_672/a_8_216# OR2X1_LOC_46/A 0.01fF
C27202 OR2X1_LOC_426/B OR2X1_LOC_46/A 0.10fF
C27268 AND2X1_LOC_95/Y OR2X1_LOC_46/A 0.20fF
C27336 OR2X1_LOC_246/A OR2X1_LOC_46/A 0.03fF
C27431 OR2X1_LOC_46/A OR2X1_LOC_599/a_8_216# 0.14fF
C28483 OR2X1_LOC_235/B OR2X1_LOC_46/A 0.08fF
C29377 OR2X1_LOC_96/B OR2X1_LOC_46/A 0.01fF
C29667 OR2X1_LOC_693/a_8_216# OR2X1_LOC_46/A 0.07fF
C30090 OR2X1_LOC_46/A OR2X1_LOC_414/Y 0.01fF
C30184 OR2X1_LOC_92/Y OR2X1_LOC_46/A 0.02fF
C30288 OR2X1_LOC_62/a_8_216# OR2X1_LOC_46/A 0.01fF
C30487 OR2X1_LOC_46/A AND2X1_LOC_44/Y 0.37fF
C30499 OR2X1_LOC_692/Y OR2X1_LOC_46/A 0.03fF
C30534 OR2X1_LOC_600/A OR2X1_LOC_46/A 3.25fF
C30615 OR2X1_LOC_619/Y OR2X1_LOC_46/A 0.10fF
C31181 OR2X1_LOC_289/Y OR2X1_LOC_46/A 0.01fF
C31486 OR2X1_LOC_46/A AND2X1_LOC_413/a_8_24# 0.03fF
C31774 OR2X1_LOC_133/a_8_216# OR2X1_LOC_46/A 0.06fF
C31795 OR2X1_LOC_411/A OR2X1_LOC_46/A 0.03fF
C32344 OR2X1_LOC_62/B OR2X1_LOC_46/A 0.23fF
C32921 OR2X1_LOC_46/A OR2X1_LOC_13/B 0.03fF
C33452 OR2X1_LOC_46/A OR2X1_LOC_428/A 0.02fF
C34069 OR2X1_LOC_54/Y OR2X1_LOC_46/A 1.17fF
C34431 OR2X1_LOC_26/Y OR2X1_LOC_46/A 0.33fF
C34441 OR2X1_LOC_89/A OR2X1_LOC_46/A 0.05fF
C35334 OR2X1_LOC_95/Y OR2X1_LOC_46/A 0.08fF
C36276 OR2X1_LOC_46/A OR2X1_LOC_71/A 0.08fF
C36463 OR2X1_LOC_46/A OR2X1_LOC_59/Y 0.04fF
C36537 OR2X1_LOC_46/A OR2X1_LOC_820/B 0.04fF
C36565 OR2X1_LOC_70/Y OR2X1_LOC_46/A 0.03fF
C36575 AND2X1_LOC_514/Y OR2X1_LOC_46/A 0.03fF
C36958 OR2X1_LOC_46/A OR2X1_LOC_240/A 0.03fF
C37046 OR2X1_LOC_47/Y OR2X1_LOC_46/A 0.26fF
C37055 AND2X1_LOC_461/a_8_24# OR2X1_LOC_46/A 0.01fF
C38069 OR2X1_LOC_46/A OR2X1_LOC_16/A 0.18fF
C38311 AND2X1_LOC_827/a_8_24# OR2X1_LOC_46/A 0.17fF
C39151 AND2X1_LOC_729/B OR2X1_LOC_46/A 0.02fF
C39938 OR2X1_LOC_599/A OR2X1_LOC_46/A 0.02fF
C40221 OR2X1_LOC_159/a_8_216# OR2X1_LOC_46/A 0.01fF
C40224 OR2X1_LOC_40/Y OR2X1_LOC_46/A 0.22fF
C40371 OR2X1_LOC_7/A OR2X1_LOC_46/A 0.03fF
C40740 OR2X1_LOC_46/A OR2X1_LOC_46/a_8_216# 0.01fF
C41077 OR2X1_LOC_46/A AND2X1_LOC_415/a_8_24# 0.02fF
C41538 OR2X1_LOC_589/A OR2X1_LOC_46/A 0.03fF
C41680 OR2X1_LOC_43/A OR2X1_LOC_46/A 0.56fF
C42586 OR2X1_LOC_3/Y OR2X1_LOC_46/A 0.15fF
C42669 AND2X1_LOC_462/B OR2X1_LOC_46/A 0.03fF
C43861 OR2X1_LOC_690/A OR2X1_LOC_46/A 0.39fF
C43892 OR2X1_LOC_64/Y OR2X1_LOC_46/A 0.05fF
C45202 OR2X1_LOC_46/A OR2X1_LOC_77/a_8_216# 0.07fF
C45598 AND2X1_LOC_512/a_8_24# OR2X1_LOC_46/A 0.17fF
C45687 OR2X1_LOC_46/A OR2X1_LOC_28/a_8_216# 0.42fF
C46475 OR2X1_LOC_46/A AND2X1_LOC_233/a_8_24# 0.01fF
C47402 OR2X1_LOC_827/a_8_216# OR2X1_LOC_46/A 0.01fF
C47786 AND2X1_LOC_62/a_8_24# OR2X1_LOC_46/A 0.02fF
C48674 OR2X1_LOC_46/A OR2X1_LOC_49/a_8_216# 0.03fF
C49507 OR2X1_LOC_46/A OR2X1_LOC_38/a_8_216# 0.01fF
C49578 OR2X1_LOC_19/B OR2X1_LOC_46/A 0.25fF
C49624 OR2X1_LOC_838/B OR2X1_LOC_46/A 0.06fF
C50754 AND2X1_LOC_377/a_8_24# OR2X1_LOC_46/A 0.11fF
C50847 OR2X1_LOC_46/A OR2X1_LOC_77/a_36_216# 0.01fF
C51185 OR2X1_LOC_36/Y OR2X1_LOC_46/A 3.86fF
C51495 OR2X1_LOC_604/A OR2X1_LOC_46/A 0.04fF
C51585 OR2X1_LOC_306/Y OR2X1_LOC_46/A 0.63fF
C51947 AND2X1_LOC_94/Y OR2X1_LOC_46/A 0.10fF
C52007 OR2X1_LOC_413/a_8_216# OR2X1_LOC_46/A 0.01fF
C53223 OR2X1_LOC_90/a_8_216# OR2X1_LOC_46/A 0.03fF
C54133 OR2X1_LOC_46/A OR2X1_LOC_49/a_36_216# 0.03fF
C54145 OR2X1_LOC_73/a_8_216# OR2X1_LOC_46/A 0.01fF
C54824 OR2X1_LOC_46/A OR2X1_LOC_12/Y 0.25fF
C55458 OR2X1_LOC_278/A OR2X1_LOC_46/A 3.80fF
C56819 OR2X1_LOC_46/A VSS 1.13fF
C6821 OR2X1_LOC_8/Y OR2X1_LOC_618/Y 0.01fF
C8240 OR2X1_LOC_618/Y OR2X1_LOC_85/A 0.03fF
C28571 OR2X1_LOC_618/Y AND2X1_LOC_9/a_8_24# 0.10fF
C35788 OR2X1_LOC_62/B OR2X1_LOC_618/Y 0.81fF
C54585 OR2X1_LOC_36/Y OR2X1_LOC_618/Y 0.10fF
C57082 OR2X1_LOC_618/Y VSS 0.12fF
C1577 AND2X1_LOC_91/B AND2X1_LOC_42/B 0.11fF
C2212 AND2X1_LOC_56/B AND2X1_LOC_42/B 0.05fF
C2223 AND2X1_LOC_8/Y AND2X1_LOC_42/B 0.43fF
C3086 AND2X1_LOC_42/B OR2X1_LOC_83/A 0.02fF
C3376 OR2X1_LOC_6/B AND2X1_LOC_42/B 1.13fF
C3411 AND2X1_LOC_73/a_8_24# AND2X1_LOC_42/B 0.09fF
C3571 AND2X1_LOC_42/B AND2X1_LOC_47/Y 1.43fF
C4256 AND2X1_LOC_95/Y AND2X1_LOC_42/B 0.08fF
C4524 AND2X1_LOC_22/Y AND2X1_LOC_42/B 0.52fF
C4692 AND2X1_LOC_153/a_8_24# AND2X1_LOC_42/B 0.11fF
C5451 OR2X1_LOC_235/B AND2X1_LOC_42/B 0.15fF
C5625 OR2X1_LOC_276/B AND2X1_LOC_42/B 0.07fF
C5886 AND2X1_LOC_70/Y AND2X1_LOC_42/B 0.03fF
C7547 AND2X1_LOC_42/B AND2X1_LOC_44/Y 0.45fF
C8507 AND2X1_LOC_42/B AND2X1_LOC_18/Y 2.19fF
C9526 AND2X1_LOC_42/B OR2X1_LOC_62/B 0.22fF
C10946 AND2X1_LOC_42/B OR2X1_LOC_548/B 0.04fF
C11165 AND2X1_LOC_42/B OR2X1_LOC_54/Y 0.03fF
C11530 AND2X1_LOC_42/B OR2X1_LOC_161/A 0.06fF
C11593 AND2X1_LOC_42/B AND2X1_LOC_51/Y 0.03fF
C12332 AND2X1_LOC_41/A AND2X1_LOC_42/B 0.74fF
C13306 AND2X1_LOC_102/a_8_24# AND2X1_LOC_42/B 0.17fF
C13437 AND2X1_LOC_42/B OR2X1_LOC_71/A 1.29fF
C13825 AND2X1_LOC_42/B AND2X1_LOC_31/Y 0.02fF
C14143 AND2X1_LOC_42/B OR2X1_LOC_240/A 0.16fF
C14357 AND2X1_LOC_42/B OR2X1_LOC_121/A 0.03fF
C14650 AND2X1_LOC_42/B AND2X1_LOC_72/B 0.03fF
C14723 AND2X1_LOC_42/B AND2X1_LOC_36/Y 0.16fF
C16455 AND2X1_LOC_42/B OR2X1_LOC_548/a_8_216# 0.05fF
C17918 AND2X1_LOC_42/a_8_24# AND2X1_LOC_42/B 0.06fF
C18139 AND2X1_LOC_42/B OR2X1_LOC_831/B 0.06fF
C18200 AND2X1_LOC_150/a_8_24# AND2X1_LOC_42/B 0.03fF
C18618 AND2X1_LOC_42/B OR2X1_LOC_161/B 0.05fF
C18741 AND2X1_LOC_42/B AND2X1_LOC_618/a_8_24# 0.01fF
C18787 AND2X1_LOC_42/B OR2X1_LOC_87/a_8_216# 0.01fF
C19666 OR2X1_LOC_3/Y AND2X1_LOC_42/B 0.08fF
C19728 AND2X1_LOC_42/B OR2X1_LOC_673/A 0.02fF
C20011 OR2X1_LOC_502/A AND2X1_LOC_42/B 0.05fF
C20126 AND2X1_LOC_48/A AND2X1_LOC_42/B 0.01fF
C20508 AND2X1_LOC_42/B AND2X1_LOC_3/Y 0.06fF
C21175 AND2X1_LOC_42/B AND2X1_LOC_7/B 0.06fF
C21403 OR2X1_LOC_296/Y AND2X1_LOC_42/B 0.03fF
C21711 AND2X1_LOC_372/a_8_24# AND2X1_LOC_42/B 0.17fF
C22975 OR2X1_LOC_160/B AND2X1_LOC_42/B 0.21fF
C23771 OR2X1_LOC_151/A AND2X1_LOC_42/B 0.07fF
C24277 AND2X1_LOC_42/B AND2X1_LOC_619/B 0.01fF
C24955 AND2X1_LOC_42/B OR2X1_LOC_415/Y 0.06fF
C26444 OR2X1_LOC_19/B AND2X1_LOC_42/B 0.13fF
C28411 AND2X1_LOC_42/B OR2X1_LOC_66/A 6.03fF
C28831 AND2X1_LOC_94/Y AND2X1_LOC_42/B 0.02fF
C28955 AND2X1_LOC_42/a_36_24# AND2X1_LOC_42/B 0.01fF
C29714 AND2X1_LOC_40/Y AND2X1_LOC_42/B 0.03fF
C29774 AND2X1_LOC_42/B OR2X1_LOC_87/Y 0.01fF
C31179 AND2X1_LOC_42/B OR2X1_LOC_398/Y 0.03fF
C31251 AND2X1_LOC_42/B AND2X1_LOC_619/a_8_24# 0.02fF
C32113 AND2X1_LOC_42/B AND2X1_LOC_255/a_8_24# 0.03fF
C32634 AND2X1_LOC_42/B OR2X1_LOC_78/A 0.10fF
C32651 OR2X1_LOC_458/B AND2X1_LOC_42/B 0.04fF
C33214 AND2X1_LOC_42/B OR2X1_LOC_814/A 0.07fF
C33977 AND2X1_LOC_12/Y AND2X1_LOC_42/B 0.03fF
C34371 AND2X1_LOC_59/Y AND2X1_LOC_42/B 0.07fF
C36688 AND2X1_LOC_42/B OR2X1_LOC_622/B 0.02fF
C37751 OR2X1_LOC_377/A AND2X1_LOC_42/B 5.91fF
C38095 AND2X1_LOC_42/B OR2X1_LOC_78/B 0.07fF
C38183 AND2X1_LOC_42/B OR2X1_LOC_375/A 0.29fF
C38485 AND2X1_LOC_42/B OR2X1_LOC_549/A 0.07fF
C39358 AND2X1_LOC_42/B AND2X1_LOC_65/A 0.01fF
C39944 AND2X1_LOC_10/a_8_24# AND2X1_LOC_42/B 0.01fF
C40211 AND2X1_LOC_19/Y AND2X1_LOC_42/B 0.06fF
C40595 AND2X1_LOC_42/B AND2X1_LOC_277/a_8_24# 0.09fF
C41672 AND2X1_LOC_42/B AND2X1_LOC_38/a_8_24# 0.01fF
C41772 AND2X1_LOC_42/B OR2X1_LOC_68/B 0.17fF
C42518 AND2X1_LOC_42/B OR2X1_LOC_87/A 2.63fF
C42545 AND2X1_LOC_42/B AND2X1_LOC_19/a_8_24# 0.01fF
C42934 AND2X1_LOC_42/B AND2X1_LOC_29/a_8_24# 0.01fF
C43740 OR2X1_LOC_541/A AND2X1_LOC_42/B 0.02fF
C43807 AND2X1_LOC_63/a_8_24# AND2X1_LOC_42/B 0.01fF
C44587 AND2X1_LOC_42/B OR2X1_LOC_778/B 0.14fF
C45018 AND2X1_LOC_42/B AND2X1_LOC_245/a_8_24# 0.02fF
C45102 OR2X1_LOC_154/A AND2X1_LOC_42/B 0.38fF
C46266 AND2X1_LOC_42/B OR2X1_LOC_633/A 0.15fF
C46669 AND2X1_LOC_64/Y AND2X1_LOC_42/B 0.14fF
C46821 AND2X1_LOC_42/B AND2X1_LOC_819/a_8_24# 0.01fF
C47292 OR2X1_LOC_756/B AND2X1_LOC_42/B 0.04fF
C48464 AND2X1_LOC_42/B OR2X1_LOC_120/a_8_216# 0.04fF
C48498 OR2X1_LOC_49/A AND2X1_LOC_42/B 0.38fF
C48634 AND2X1_LOC_42/B OR2X1_LOC_87/B 0.10fF
C48651 AND2X1_LOC_85/a_8_24# AND2X1_LOC_42/B 0.01fF
C48875 AND2X1_LOC_42/B AND2X1_LOC_263/a_8_24# 0.11fF
C48975 AND2X1_LOC_529/a_8_24# AND2X1_LOC_42/B 0.06fF
C49111 AND2X1_LOC_42/B OR2X1_LOC_532/B 0.86fF
C50344 OR2X1_LOC_185/Y AND2X1_LOC_42/B 0.07fF
C50355 AND2X1_LOC_42/B AND2X1_LOC_412/a_8_24# 0.10fF
C51055 VDD AND2X1_LOC_42/B 1.64fF
C52353 AND2X1_LOC_42/B AND2X1_LOC_820/B 0.83fF
C52992 AND2X1_LOC_42/B OR2X1_LOC_80/A 0.32fF
C54068 OR2X1_LOC_160/A AND2X1_LOC_42/B 0.71fF
C54109 AND2X1_LOC_86/B AND2X1_LOC_42/B 0.01fF
C54339 AND2X1_LOC_42/B OR2X1_LOC_266/A 0.23fF
C54562 AND2X1_LOC_46/a_8_24# AND2X1_LOC_42/B 0.01fF
C55362 OR2X1_LOC_185/A AND2X1_LOC_42/B 0.06fF
C57189 AND2X1_LOC_42/B VSS 0.72fF
C3081 OR2X1_LOC_68/B OR2X1_LOC_548/B 0.01fF
C7393 OR2X1_LOC_633/A OR2X1_LOC_548/B 0.01fF
C14133 OR2X1_LOC_80/A OR2X1_LOC_548/B 0.03fF
C16370 OR2X1_LOC_185/A OR2X1_LOC_548/B 0.05fF
C26703 OR2X1_LOC_62/B OR2X1_LOC_548/B 0.01fF
C30629 OR2X1_LOC_71/A OR2X1_LOC_548/B 0.01fF
C31913 AND2X1_LOC_36/Y OR2X1_LOC_548/B 0.03fF
C33700 OR2X1_LOC_548/B OR2X1_LOC_548/a_8_216# 0.07fF
C43063 OR2X1_LOC_548/A OR2X1_LOC_548/B 0.04fF
C43699 OR2X1_LOC_19/B OR2X1_LOC_548/B 0.01fF
C45676 OR2X1_LOC_66/A OR2X1_LOC_548/B 0.11fF
C55141 OR2X1_LOC_377/A OR2X1_LOC_548/B 0.13fF
C56262 OR2X1_LOC_548/B VSS 0.11fF
C3181 AND2X1_LOC_817/B AND2X1_LOC_236/a_8_24# 0.01fF
C5937 AND2X1_LOC_817/B AND2X1_LOC_817/a_8_24# 0.20fF
C14075 AND2X1_LOC_817/B OR2X1_LOC_847/a_8_216# 0.01fF
C17026 AND2X1_LOC_817/B OR2X1_LOC_847/B 0.01fF
C17850 AND2X1_LOC_817/B OR2X1_LOC_269/B 0.05fF
C30551 AND2X1_LOC_817/B OR2X1_LOC_848/A 0.16fF
C34774 AND2X1_LOC_12/Y AND2X1_LOC_817/B 0.01fF
C42631 AND2X1_LOC_817/B OR2X1_LOC_68/B 0.01fF
C51850 AND2X1_LOC_817/B VDD 0.37fF
C53817 AND2X1_LOC_817/B OR2X1_LOC_80/A 0.46fF
C58019 AND2X1_LOC_817/B VSS 0.16fF
C7387 VDD OR2X1_LOC_387/A 0.06fF
C10035 OR2X1_LOC_44/Y OR2X1_LOC_387/A 0.02fF
C13391 OR2X1_LOC_744/A OR2X1_LOC_387/A 0.18fF
C13546 OR2X1_LOC_31/Y OR2X1_LOC_387/A 0.01fF
C16931 OR2X1_LOC_409/B OR2X1_LOC_387/A 0.16fF
C23125 OR2X1_LOC_428/A OR2X1_LOC_387/A 0.06fF
C26310 OR2X1_LOC_70/A OR2X1_LOC_387/A 0.32fF
C26698 OR2X1_LOC_47/Y OR2X1_LOC_387/A 0.01fF
C29864 OR2X1_LOC_40/Y OR2X1_LOC_387/A 0.83fF
C32049 OR2X1_LOC_3/Y OR2X1_LOC_387/A 0.01fF
C33373 OR2X1_LOC_64/Y OR2X1_LOC_387/A 0.02fF
C34947 OR2X1_LOC_421/A OR2X1_LOC_387/A 0.02fF
C37029 OR2X1_LOC_328/a_8_216# OR2X1_LOC_387/A 0.40fF
C37546 OR2X1_LOC_763/Y OR2X1_LOC_387/A 0.18fF
C44313 OR2X1_LOC_12/Y OR2X1_LOC_387/A 0.03fF
C47061 OR2X1_LOC_18/Y OR2X1_LOC_387/A 0.02fF
C47559 OR2X1_LOC_585/A OR2X1_LOC_387/A 0.06fF
C49837 OR2X1_LOC_387/A OR2X1_LOC_387/a_8_216# 0.01fF
C50863 OR2X1_LOC_51/Y OR2X1_LOC_387/A 0.01fF
C52617 OR2X1_LOC_387/Y OR2X1_LOC_387/A 0.05fF
C56389 OR2X1_LOC_387/A VSS 0.17fF
C619 OR2X1_LOC_421/A AND2X1_LOC_596/a_8_24# 0.01fF
C725 OR2X1_LOC_421/A OR2X1_LOC_36/Y 0.05fF
C4414 OR2X1_LOC_421/A OR2X1_LOC_12/Y 0.02fF
C6128 OR2X1_LOC_421/A OR2X1_LOC_597/A 0.01fF
C7078 OR2X1_LOC_421/A OR2X1_LOC_18/Y 0.01fF
C9313 OR2X1_LOC_421/A OR2X1_LOC_52/B 0.04fF
C9800 OR2X1_LOC_421/A OR2X1_LOC_22/Y 0.11fF
C10480 OR2X1_LOC_421/A OR2X1_LOC_421/a_8_216# 0.18fF
C10865 OR2X1_LOC_421/A OR2X1_LOC_51/Y 0.01fF
C13881 OR2X1_LOC_421/A OR2X1_LOC_91/A 0.10fF
C18652 OR2X1_LOC_421/A OR2X1_LOC_485/A 0.03fF
C21164 OR2X1_LOC_421/A OR2X1_LOC_433/Y 0.04fF
C23642 OR2X1_LOC_421/A VDD 0.63fF
C24947 OR2X1_LOC_421/A OR2X1_LOC_427/A 0.03fF
C26237 OR2X1_LOC_421/A OR2X1_LOC_44/Y 0.15fF
C26518 OR2X1_LOC_45/B OR2X1_LOC_421/A 0.04fF
C26958 OR2X1_LOC_421/A OR2X1_LOC_158/A 2.52fF
C29534 OR2X1_LOC_421/A OR2X1_LOC_744/A 0.04fF
C29723 OR2X1_LOC_421/A OR2X1_LOC_31/Y 0.06fF
C32884 OR2X1_LOC_421/A OR2X1_LOC_426/B 0.02fF
C35357 OR2X1_LOC_421/A OR2X1_LOC_693/a_8_216# 0.01fF
C35881 OR2X1_LOC_421/A OR2X1_LOC_692/a_8_216# 0.01fF
C35887 OR2X1_LOC_421/A OR2X1_LOC_92/Y 0.07fF
C36220 OR2X1_LOC_421/A OR2X1_LOC_692/Y 0.01fF
C39200 OR2X1_LOC_421/A OR2X1_LOC_428/A 2.69fF
C39782 OR2X1_LOC_421/A OR2X1_LOC_682/Y 0.12fF
C41769 OR2X1_LOC_421/A OR2X1_LOC_693/Y 0.01fF
C42349 OR2X1_LOC_421/A OR2X1_LOC_433/a_8_216# 0.01fF
C42412 OR2X1_LOC_421/A OR2X1_LOC_70/Y 0.05fF
C42543 OR2X1_LOC_421/A OR2X1_LOC_70/A 0.22fF
C42917 OR2X1_LOC_421/A OR2X1_LOC_47/Y 0.14fF
C43951 OR2X1_LOC_421/A OR2X1_LOC_16/A 0.03fF
C44173 OR2X1_LOC_421/A AND2X1_LOC_687/Y 0.02fF
C45812 OR2X1_LOC_421/A OR2X1_LOC_599/A 0.12fF
C46148 OR2X1_LOC_421/A OR2X1_LOC_40/Y 0.03fF
C46301 OR2X1_LOC_421/A OR2X1_LOC_7/A 0.05fF
C47502 OR2X1_LOC_421/A OR2X1_LOC_589/A 0.04fF
C47644 OR2X1_LOC_421/A OR2X1_LOC_43/A 0.03fF
C48536 OR2X1_LOC_421/A OR2X1_LOC_3/Y 0.01fF
C48805 OR2X1_LOC_421/A OR2X1_LOC_329/B 0.01fF
C49824 OR2X1_LOC_421/A OR2X1_LOC_64/Y 0.09fF
C55137 OR2X1_LOC_421/A OR2X1_LOC_763/a_8_216# 0.05fF
C57990 OR2X1_LOC_421/A VSS 0.14fF
C1669 OR2X1_LOC_53/Y OR2X1_LOC_689/Y 0.01fF
C1979 OR2X1_LOC_53/Y OR2X1_LOC_36/Y 0.06fF
C3150 OR2X1_LOC_53/Y OR2X1_LOC_304/a_8_216# 0.07fF
C6131 OR2X1_LOC_53/Y OR2X1_LOC_59/a_8_216# 0.40fF
C8370 OR2X1_LOC_53/Y OR2X1_LOC_18/Y 0.03fF
C8817 OR2X1_LOC_53/Y OR2X1_LOC_585/A 0.05fF
C9668 OR2X1_LOC_53/Y OR2X1_LOC_753/A 0.03fF
C10966 OR2X1_LOC_53/Y OR2X1_LOC_22/Y 0.07fF
C12079 OR2X1_LOC_53/Y OR2X1_LOC_51/Y 0.03fF
C14606 OR2X1_LOC_53/Y OR2X1_LOC_56/a_8_216# 0.07fF
C19882 OR2X1_LOC_53/Y OR2X1_LOC_485/A 0.02fF
C21634 OR2X1_LOC_53/Y OR2X1_LOC_43/a_8_216# 0.01fF
C23619 OR2X1_LOC_53/Y AND2X1_LOC_691/a_8_24# 0.01fF
C24843 OR2X1_LOC_53/Y VDD 0.17fF
C27445 OR2X1_LOC_53/Y OR2X1_LOC_44/Y 0.06fF
C27745 OR2X1_LOC_45/B OR2X1_LOC_53/Y 0.03fF
C30948 OR2X1_LOC_53/Y OR2X1_LOC_31/Y 0.42fF
C31965 OR2X1_LOC_53/Y OR2X1_LOC_56/A 0.06fF
C37481 OR2X1_LOC_53/Y OR2X1_LOC_600/A 0.03fF
C40414 OR2X1_LOC_53/Y OR2X1_LOC_428/A 0.32fF
C43509 OR2X1_LOC_53/Y OR2X1_LOC_59/Y 0.05fF
C43778 OR2X1_LOC_53/Y OR2X1_LOC_70/A 0.01fF
C44160 OR2X1_LOC_53/Y OR2X1_LOC_47/Y 0.02fF
C46255 OR2X1_LOC_53/Y AND2X1_LOC_729/B 0.02fF
C48835 OR2X1_LOC_53/Y OR2X1_LOC_43/A 1.78fF
C49723 OR2X1_LOC_53/Y OR2X1_LOC_3/Y 0.04fF
C50962 OR2X1_LOC_53/Y OR2X1_LOC_690/A 0.25fF
C52115 OR2X1_LOC_53/Y OR2X1_LOC_25/Y 0.09fF
C58039 OR2X1_LOC_53/Y VSS 0.55fF
C2983 OR2X1_LOC_157/a_8_216# OR2X1_LOC_2/Y 0.04fF
C4584 OR2X1_LOC_2/Y OR2X1_LOC_30/a_8_216# 0.02fF
C5576 OR2X1_LOC_50/a_8_216# OR2X1_LOC_2/Y 0.02fF
C9412 OR2X1_LOC_429/Y OR2X1_LOC_2/Y 0.29fF
C10102 OR2X1_LOC_51/Y OR2X1_LOC_2/Y 0.07fF
C14596 OR2X1_LOC_2/Y OR2X1_LOC_581/a_8_216# 0.01fF
C22007 OR2X1_LOC_2/Y OR2X1_LOC_581/Y 0.04fF
C22576 OR2X1_LOC_2/Y OR2X1_LOC_25/a_8_216# 0.02fF
C24209 OR2X1_LOC_427/A OR2X1_LOC_2/Y 0.10fF
C26172 OR2X1_LOC_158/A OR2X1_LOC_2/Y 0.14fF
C28942 OR2X1_LOC_31/Y OR2X1_LOC_2/Y 0.01fF
C30675 OR2X1_LOC_2/Y OR2X1_LOC_11/a_8_216# 0.02fF
C31096 OR2X1_LOC_51/a_8_216# OR2X1_LOC_2/Y 0.01fF
C32576 OR2X1_LOC_425/a_8_216# OR2X1_LOC_2/Y 0.01fF
C35242 OR2X1_LOC_2/Y OR2X1_LOC_429/a_8_216# 0.02fF
C36951 OR2X1_LOC_2/Y OR2X1_LOC_51/B 0.03fF
C39879 OR2X1_LOC_2/Y OR2X1_LOC_17/Y 0.22fF
C41602 OR2X1_LOC_70/Y OR2X1_LOC_2/Y 0.10fF
C41712 OR2X1_LOC_2/Y OR2X1_LOC_70/A 0.83fF
C42105 OR2X1_LOC_47/Y OR2X1_LOC_2/Y 0.08fF
C42576 OR2X1_LOC_2/Y OR2X1_LOC_3/B 0.12fF
C43683 OR2X1_LOC_426/A OR2X1_LOC_2/Y 0.18fF
C45330 OR2X1_LOC_40/Y OR2X1_LOC_2/Y 0.09fF
C48957 OR2X1_LOC_2/Y OR2X1_LOC_11/Y 0.03fF
C50148 OR2X1_LOC_2/Y OR2X1_LOC_25/Y 0.38fF
C51161 OR2X1_LOC_70/a_8_216# OR2X1_LOC_2/Y 0.08fF
C51608 OR2X1_LOC_2/Y OR2X1_LOC_17/a_8_216# 0.41fF
C55256 OR2X1_LOC_2/Y OR2X1_LOC_40/a_8_216# 0.07fF
C57017 OR2X1_LOC_2/Y VSS 0.49fF
C1752 OR2X1_LOC_426/A OR2X1_LOC_684/Y 0.16fF
C2581 OR2X1_LOC_426/A OR2X1_LOC_52/B 0.01fF
C3435 OR2X1_LOC_429/Y OR2X1_LOC_426/A 0.05fF
C4107 OR2X1_LOC_51/Y OR2X1_LOC_426/A 0.02fF
C7093 OR2X1_LOC_91/A OR2X1_LOC_426/A 0.16fF
C8667 OR2X1_LOC_426/A OR2X1_LOC_581/a_8_216# 0.40fF
C15966 OR2X1_LOC_426/A OR2X1_LOC_581/Y 0.34fF
C16849 VDD OR2X1_LOC_426/A 0.08fF
C18205 OR2X1_LOC_426/A OR2X1_LOC_427/A 0.42fF
C18341 OR2X1_LOC_426/A AND2X1_LOC_687/B 1.00fF
C19854 OR2X1_LOC_684/a_8_216# OR2X1_LOC_426/A 0.01fF
C20019 OR2X1_LOC_430/a_8_216# OR2X1_LOC_426/A 0.01fF
C23085 OR2X1_LOC_426/A OR2X1_LOC_31/Y 0.03fF
C24195 OR2X1_LOC_426/A OR2X1_LOC_426/Y 0.01fF
C26197 OR2X1_LOC_426/B OR2X1_LOC_426/A 0.15fF
C26660 OR2X1_LOC_425/a_8_216# OR2X1_LOC_426/A -0.00fF
C27040 OR2X1_LOC_426/A OR2X1_LOC_582/a_8_216# 0.01fF
C28134 OR2X1_LOC_426/A OR2X1_LOC_430/Y 0.01fF
C33618 OR2X1_LOC_426/A OR2X1_LOC_426/a_8_216# 0.04fF
C35631 OR2X1_LOC_70/Y OR2X1_LOC_426/A 1.53fF
C35736 OR2X1_LOC_426/A OR2X1_LOC_70/A 0.26fF
C37104 OR2X1_LOC_426/A OR2X1_LOC_16/A 0.33fF
C39440 OR2X1_LOC_426/A OR2X1_LOC_7/A 0.01fF
C40667 OR2X1_LOC_43/A OR2X1_LOC_426/A 0.30fF
C41585 OR2X1_LOC_3/Y OR2X1_LOC_426/A 0.01fF
C41625 OR2X1_LOC_426/A OR2X1_LOC_582/Y 0.01fF
C42907 OR2X1_LOC_64/Y OR2X1_LOC_426/A 0.03fF
C45120 OR2X1_LOC_70/a_8_216# OR2X1_LOC_426/A 0.01fF
C50531 OR2X1_LOC_604/A OR2X1_LOC_426/A 0.03fF
C53868 OR2X1_LOC_426/A OR2X1_LOC_12/Y 0.18fF
C57165 OR2X1_LOC_426/A VSS 0.36fF
C1560 AND2X1_LOC_587/a_8_24# AND2X1_LOC_51/A 0.01fF
C3041 AND2X1_LOC_51/A AND2X1_LOC_47/a_8_24# 0.01fF
C7059 AND2X1_LOC_588/B AND2X1_LOC_51/A 0.01fF
C16943 VDD AND2X1_LOC_51/A 0.37fF
C19664 AND2X1_LOC_1/Y AND2X1_LOC_51/A 0.01fF
C24325 AND2X1_LOC_51/A AND2X1_LOC_21/Y 0.07fF
C25050 AND2X1_LOC_51/a_8_24# AND2X1_LOC_51/A 0.20fF
C25630 AND2X1_LOC_51/A AND2X1_LOC_47/Y 0.04fF
C28095 AND2X1_LOC_17/Y AND2X1_LOC_51/A 0.73fF
C28860 AND2X1_LOC_51/A AND2X1_LOC_11/Y 0.12fF
C29582 AND2X1_LOC_51/A AND2X1_LOC_44/Y 0.01fF
C33623 AND2X1_LOC_51/A AND2X1_LOC_51/Y 0.43fF
C35793 AND2X1_LOC_51/A AND2X1_LOC_31/Y 0.09fF
C36124 AND2X1_LOC_31/a_8_24# AND2X1_LOC_51/A 0.03fF
C43375 AND2X1_LOC_51/A AND2X1_LOC_44/a_8_24# 0.04fF
C51082 AND2X1_LOC_50/Y AND2X1_LOC_51/A 0.01fF
C57403 AND2X1_LOC_51/A VSS -0.04fF
C2486 AND2X1_LOC_753/B AND2X1_LOC_41/A 0.91fF
C3985 AND2X1_LOC_753/B AND2X1_LOC_31/Y 0.04fF
C7193 AND2X1_LOC_753/B OR2X1_LOC_269/B 0.16fF
C9884 AND2X1_LOC_753/B AND2X1_LOC_53/Y 0.12fF
C10136 AND2X1_LOC_753/B OR2X1_LOC_502/A 0.03fF
C10282 AND2X1_LOC_753/B AND2X1_LOC_48/A 0.15fF
C10658 AND2X1_LOC_753/B AND2X1_LOC_3/Y 0.04fF
C11275 AND2X1_LOC_753/B AND2X1_LOC_7/B 0.04fF
C18564 AND2X1_LOC_753/B OR2X1_LOC_66/A 0.07fF
C19050 AND2X1_LOC_50/Y AND2X1_LOC_753/B 0.03fF
C19923 AND2X1_LOC_753/B AND2X1_LOC_40/Y 0.07fF
C20949 AND2X1_LOC_753/B AND2X1_LOC_56/a_8_24# 0.04fF
C23854 AND2X1_LOC_753/B AND2X1_LOC_387/B 0.07fF
C24619 AND2X1_LOC_753/B AND2X1_LOC_59/Y 0.07fF
C26398 AND2X1_LOC_753/B OR2X1_LOC_197/A 0.05fF
C28418 AND2X1_LOC_753/B OR2X1_LOC_375/A 0.68fF
C32635 AND2X1_LOC_753/B OR2X1_LOC_87/A 0.20fF
C35823 AND2X1_LOC_753/B AND2X1_LOC_763/B 0.02fF
C36638 AND2X1_LOC_753/B AND2X1_LOC_64/Y 0.07fF
C38382 AND2X1_LOC_753/B OR2X1_LOC_596/A 0.07fF
C40210 AND2X1_LOC_753/B OR2X1_LOC_185/Y 0.21fF
C40621 AND2X1_LOC_753/B AND2X1_LOC_53/a_8_24# 0.06fF
C40966 AND2X1_LOC_753/B VDD 0.15fF
C46768 AND2X1_LOC_753/B AND2X1_LOC_753/a_8_24# 0.02fF
C48558 AND2X1_LOC_753/B AND2X1_LOC_56/B 0.02fF
C50627 AND2X1_LOC_753/B AND2X1_LOC_95/Y 0.07fF
C50915 AND2X1_LOC_753/B AND2X1_LOC_22/Y 0.07fF
C51820 AND2X1_LOC_753/B OR2X1_LOC_638/B 0.07fF
C52209 AND2X1_LOC_753/B AND2X1_LOC_70/Y 0.07fF
C53863 AND2X1_LOC_753/B AND2X1_LOC_44/Y 0.02fF
C54726 AND2X1_LOC_753/B AND2X1_LOC_18/Y 0.33fF
C58117 AND2X1_LOC_753/B VSS 0.46fF
C8644 AND2X1_LOC_581/a_8_24# AND2X1_LOC_582/B 0.01fF
C18927 AND2X1_LOC_12/Y AND2X1_LOC_582/B 0.14fF
C25388 AND2X1_LOC_425/Y AND2X1_LOC_582/B 0.01fF
C35764 VDD AND2X1_LOC_582/B 0.02fF
C44802 AND2X1_LOC_582/a_8_24# AND2X1_LOC_582/B 0.01fF
C46841 AND2X1_LOC_430/B AND2X1_LOC_582/B 0.01fF
C55958 OR2X1_LOC_635/A AND2X1_LOC_582/B 0.83fF
C56247 AND2X1_LOC_582/B VSS 0.08fF
C10732 AND2X1_LOC_36/Y AND2X1_LOC_763/B 0.01fF
C15618 AND2X1_LOC_53/Y AND2X1_LOC_763/B 0.12fF
C15902 OR2X1_LOC_502/A AND2X1_LOC_763/B 0.01fF
C16032 AND2X1_LOC_48/A AND2X1_LOC_763/B 0.04fF
C24861 AND2X1_LOC_50/Y AND2X1_LOC_763/B 0.01fF
C26680 AND2X1_LOC_56/a_8_24# AND2X1_LOC_763/B 0.09fF
C28260 OR2X1_LOC_828/B AND2X1_LOC_763/B 0.04fF
C34151 OR2X1_LOC_375/A AND2X1_LOC_763/B 0.02fF
C42575 AND2X1_LOC_64/Y AND2X1_LOC_763/B 1.15fF
C46999 VDD AND2X1_LOC_763/B 0.30fF
C54260 AND2X1_LOC_56/B AND2X1_LOC_763/B 0.51fF
C54287 AND2X1_LOC_21/Y AND2X1_LOC_763/B 0.01fF
C55661 AND2X1_LOC_47/Y AND2X1_LOC_763/B 0.01fF
C56263 AND2X1_LOC_763/B VSS 0.19fF
C4029 OR2X1_LOC_408/Y OR2X1_LOC_409/B 0.14fF
C7395 OR2X1_LOC_22/A OR2X1_LOC_408/Y 0.02fF
C20545 OR2X1_LOC_11/Y OR2X1_LOC_408/Y 0.02fF
C27716 OR2X1_LOC_36/Y OR2X1_LOC_408/Y 0.03fF
C50731 VDD OR2X1_LOC_408/Y 0.12fF
C56874 OR2X1_LOC_408/Y VSS 0.13fF
C13285 VDD OR2X1_LOC_588/A 0.09fF
C26109 OR2X1_LOC_22/A OR2X1_LOC_588/A 0.02fF
C27410 OR2X1_LOC_51/B OR2X1_LOC_588/A 0.09fF
C32888 OR2X1_LOC_3/B OR2X1_LOC_588/A 0.01fF
C38362 OR2X1_LOC_31/a_8_216# OR2X1_LOC_588/A 0.40fF
C39150 OR2X1_LOC_11/Y OR2X1_LOC_588/A 0.02fF
C49655 OR2X1_LOC_409/Y OR2X1_LOC_588/A 0.19fF
C56496 OR2X1_LOC_588/A VSS 0.17fF
C1384 OR2X1_LOC_70/Y OR2X1_LOC_429/Y 0.06fF
C1474 OR2X1_LOC_429/Y OR2X1_LOC_70/A 0.17fF
C7330 OR2X1_LOC_429/Y OR2X1_LOC_582/Y 0.13fF
C9788 OR2X1_LOC_429/Y OR2X1_LOC_25/Y 0.01fF
C10784 OR2X1_LOC_429/Y OR2X1_LOC_70/a_8_216# 0.05fF
C16078 OR2X1_LOC_604/A OR2X1_LOC_429/Y 0.23fF
C18786 OR2X1_LOC_157/a_8_216# OR2X1_LOC_429/Y 0.03fF
C21866 OR2X1_LOC_429/Y OR2X1_LOC_70/a_36_216# 0.01fF
C24309 OR2X1_LOC_157/a_36_216# OR2X1_LOC_429/Y 0.01fF
C25864 OR2X1_LOC_429/Y OR2X1_LOC_51/Y 0.03fF
C30307 OR2X1_LOC_429/Y OR2X1_LOC_581/a_8_216# 0.05fF
C35781 OR2X1_LOC_429/Y OR2X1_LOC_581/a_36_216# 0.01fF
C37643 OR2X1_LOC_429/Y OR2X1_LOC_581/Y 0.05fF
C38195 OR2X1_LOC_429/Y OR2X1_LOC_25/a_8_216# 0.41fF
C38508 VDD OR2X1_LOC_429/Y 0.66fF
C39877 OR2X1_LOC_429/Y OR2X1_LOC_427/A 0.02fF
C41674 OR2X1_LOC_429/Y OR2X1_LOC_430/a_8_216# 0.06fF
C41923 OR2X1_LOC_158/A OR2X1_LOC_429/Y 0.01fF
C43815 OR2X1_LOC_429/Y OR2X1_LOC_25/a_36_216# 0.01fF
C44745 OR2X1_LOC_429/Y OR2X1_LOC_31/Y 0.02fF
C46990 OR2X1_LOC_429/Y OR2X1_LOC_51/a_8_216# 0.03fF
C48575 OR2X1_LOC_429/Y OR2X1_LOC_425/a_8_216# 0.05fF
C48940 OR2X1_LOC_429/Y OR2X1_LOC_582/a_8_216# 0.05fF
C52521 OR2X1_LOC_429/Y OR2X1_LOC_51/a_36_216# 0.01fF
C52951 OR2X1_LOC_429/Y OR2X1_LOC_51/B 0.02fF
C54032 OR2X1_LOC_429/Y OR2X1_LOC_425/a_36_216# 0.01fF
C54338 OR2X1_LOC_429/Y OR2X1_LOC_428/A 0.02fF
C54412 OR2X1_LOC_429/Y OR2X1_LOC_582/a_36_216# 0.01fF
C55857 OR2X1_LOC_429/Y OR2X1_LOC_17/Y 0.03fF
C57506 OR2X1_LOC_429/Y VSS -1.29fF
C1076 OR2X1_LOC_22/Y OR2X1_LOC_70/A 0.97fF
C2242 OR2X1_LOC_51/Y OR2X1_LOC_70/A 0.10fF
C3177 OR2X1_LOC_70/A OR2X1_LOC_588/Y 0.02fF
C6611 OR2X1_LOC_70/A OR2X1_LOC_581/a_8_216# 0.01fF
C13768 OR2X1_LOC_70/A OR2X1_LOC_53/a_8_216# 0.08fF
C14145 OR2X1_LOC_70/A OR2X1_LOC_581/Y 0.09fF
C14636 OR2X1_LOC_70/A OR2X1_LOC_25/a_8_216# 0.01fF
C14981 VDD OR2X1_LOC_70/A 0.27fF
C17559 OR2X1_LOC_70/A OR2X1_LOC_44/Y 0.09fF
C18359 OR2X1_LOC_158/A OR2X1_LOC_70/A 0.20fF
C20976 OR2X1_LOC_744/A OR2X1_LOC_70/A 0.28fF
C21091 OR2X1_LOC_31/Y OR2X1_LOC_70/A 0.05fF
C22926 OR2X1_LOC_70/A OR2X1_LOC_11/a_8_216# 0.39fF
C23277 OR2X1_LOC_51/a_8_216# OR2X1_LOC_70/A 0.06fF
C24300 OR2X1_LOC_70/A OR2X1_LOC_585/a_8_216# 0.01fF
C24480 OR2X1_LOC_70/A OR2X1_LOC_409/B 0.89fF
C24789 OR2X1_LOC_425/a_8_216# OR2X1_LOC_70/A 0.01fF
C27397 OR2X1_LOC_429/a_8_216# OR2X1_LOC_70/A 0.01fF
C27814 OR2X1_LOC_70/A OR2X1_LOC_22/A 0.10fF
C29132 OR2X1_LOC_51/B OR2X1_LOC_70/A 0.16fF
C29827 OR2X1_LOC_70/A OR2X1_LOC_762/Y 0.01fF
C30585 OR2X1_LOC_70/A OR2X1_LOC_428/A 0.03fF
C31572 OR2X1_LOC_26/Y OR2X1_LOC_70/A 0.68fF
C31964 OR2X1_LOC_70/A OR2X1_LOC_17/Y 0.26fF
C33640 OR2X1_LOC_70/A OR2X1_LOC_59/Y 0.01fF
C33845 OR2X1_LOC_70/A OR2X1_LOC_11/a_36_216# -0.00fF
C34180 OR2X1_LOC_47/Y OR2X1_LOC_70/A 0.13fF
C34605 OR2X1_LOC_3/B OR2X1_LOC_70/A 0.22fF
C37367 OR2X1_LOC_40/Y OR2X1_LOC_70/A 0.02fF
C39107 OR2X1_LOC_70/A OR2X1_LOC_585/Y 0.01fF
C39623 OR2X1_LOC_3/Y OR2X1_LOC_70/A 0.12fF
C40836 OR2X1_LOC_11/Y OR2X1_LOC_70/A 1.07fF
C40924 OR2X1_LOC_64/a_8_216# OR2X1_LOC_70/A 0.07fF
C42109 OR2X1_LOC_70/A OR2X1_LOC_25/Y 1.12fF
C44704 OR2X1_LOC_328/a_8_216# OR2X1_LOC_70/A 0.18fF
C47433 OR2X1_LOC_40/a_8_216# OR2X1_LOC_70/A 0.06fF
C51242 OR2X1_LOC_157/a_8_216# OR2X1_LOC_70/A 0.01fF
C51984 OR2X1_LOC_70/A OR2X1_LOC_12/Y 0.02fF
C52487 OR2X1_LOC_70/A OR2X1_LOC_59/a_8_216# 0.01fF
C53302 OR2X1_LOC_70/A OR2X1_LOC_26/a_8_216# 0.08fF
C54603 OR2X1_LOC_18/Y OR2X1_LOC_70/A 0.03fF
C55044 OR2X1_LOC_70/A OR2X1_LOC_585/A 0.10fF
C56928 OR2X1_LOC_70/A VSS 0.35fF
C3925 AND2X1_LOC_17/Y AND2X1_LOC_18/a_8_24# 0.06fF
C7138 VDD AND2X1_LOC_17/Y 0.93fF
C9907 AND2X1_LOC_17/Y AND2X1_LOC_1/Y 0.02fF
C11372 AND2X1_LOC_17/Y AND2X1_LOC_40/a_8_24# 0.01fF
C12314 AND2X1_LOC_17/Y AND2X1_LOC_50/a_8_24# 0.20fF
C14531 AND2X1_LOC_17/Y AND2X1_LOC_21/Y 0.09fF
C15812 AND2X1_LOC_17/Y AND2X1_LOC_47/Y 0.08fF
C16867 AND2X1_LOC_22/Y AND2X1_LOC_17/Y 0.29fF
C18015 AND2X1_LOC_17/Y AND2X1_LOC_430/B 0.01fF
C18224 AND2X1_LOC_70/Y AND2X1_LOC_17/Y 0.42fF
C19146 AND2X1_LOC_17/Y AND2X1_LOC_11/Y 0.98fF
C19439 AND2X1_LOC_17/Y AND2X1_LOC_425/a_36_24# 0.01fF
C19883 AND2X1_LOC_17/Y AND2X1_LOC_44/Y 0.75fF
C23885 AND2X1_LOC_17/Y AND2X1_LOC_25/Y 0.13fF
C23931 AND2X1_LOC_17/Y AND2X1_LOC_51/Y 1.81fF
C26102 AND2X1_LOC_17/Y AND2X1_LOC_31/Y 0.80fF
C26419 AND2X1_LOC_17/Y AND2X1_LOC_31/a_8_24# 0.01fF
C26985 AND2X1_LOC_17/Y AND2X1_LOC_36/Y 0.01fF
C29224 AND2X1_LOC_2/Y AND2X1_LOC_17/Y 0.33fF
C29341 AND2X1_LOC_17/Y OR2X1_LOC_269/B 0.02fF
C32189 AND2X1_LOC_17/Y OR2X1_LOC_502/A 0.29fF
C32730 AND2X1_LOC_17/Y AND2X1_LOC_3/Y 0.05fF
C33366 AND2X1_LOC_17/Y AND2X1_LOC_7/B 0.65fF
C33595 AND2X1_LOC_17/Y AND2X1_LOC_44/a_8_24# 0.01fF
C34010 AND2X1_LOC_17/Y AND2X1_LOC_425/a_8_24# 0.04fF
C34858 AND2X1_LOC_17/Y AND2X1_LOC_386/a_8_24# 0.11fF
C40185 AND2X1_LOC_70/a_8_24# AND2X1_LOC_17/Y 0.01fF
C41109 AND2X1_LOC_50/Y AND2X1_LOC_17/Y 0.02fF
C41987 AND2X1_LOC_40/Y AND2X1_LOC_17/Y 0.01fF
C46376 AND2X1_LOC_17/Y AND2X1_LOC_22/a_8_24# 0.01fF
C46400 AND2X1_LOC_12/Y AND2X1_LOC_17/Y 0.01fF
C49439 AND2X1_LOC_17/Y AND2X1_LOC_47/a_8_24# 0.01fF
C52900 AND2X1_LOC_17/Y AND2X1_LOC_425/Y 0.01fF
C53501 AND2X1_LOC_588/B AND2X1_LOC_17/Y 0.69fF
C54909 AND2X1_LOC_17/Y OR2X1_LOC_87/A 0.04fF
C57781 AND2X1_LOC_17/Y VSS -0.81fF
C1782 AND2X1_LOC_18/Y OR2X1_LOC_801/B 0.07fF
C5574 AND2X1_LOC_41/A OR2X1_LOC_801/B 0.07fF
C8056 AND2X1_LOC_36/Y OR2X1_LOC_801/B 0.10fF
C8694 AND2X1_LOC_748/a_8_24# OR2X1_LOC_801/B -0.01fF
C10388 OR2X1_LOC_269/B OR2X1_LOC_801/B 0.07fF
C11937 OR2X1_LOC_161/B OR2X1_LOC_801/B 0.07fF
C13429 AND2X1_LOC_48/A OR2X1_LOC_801/B 0.39fF
C13796 AND2X1_LOC_3/Y OR2X1_LOC_801/B 0.09fF
C14201 OR2X1_LOC_789/B OR2X1_LOC_801/B 0.04fF
C14483 AND2X1_LOC_7/B OR2X1_LOC_801/B 0.07fF
C16207 OR2X1_LOC_160/B OR2X1_LOC_801/B 0.07fF
C19652 OR2X1_LOC_800/Y OR2X1_LOC_801/B 0.06fF
C19716 AND2X1_LOC_748/a_36_24# OR2X1_LOC_801/B 0.01fF
C19782 OR2X1_LOC_19/B OR2X1_LOC_801/B 0.02fF
C23119 AND2X1_LOC_40/Y OR2X1_LOC_801/B 0.14fF
C27323 AND2X1_LOC_12/Y OR2X1_LOC_801/B 0.01fF
C31489 OR2X1_LOC_78/B OR2X1_LOC_801/B 0.07fF
C34822 OR2X1_LOC_138/A OR2X1_LOC_801/B 0.13fF
C36108 OR2X1_LOC_801/a_8_216# OR2X1_LOC_801/B 0.07fF
C37314 OR2X1_LOC_691/Y OR2X1_LOC_801/B 0.01fF
C38282 OR2X1_LOC_154/A OR2X1_LOC_801/B 0.07fF
C43457 OR2X1_LOC_185/Y OR2X1_LOC_801/B 0.07fF
C47388 OR2X1_LOC_809/B OR2X1_LOC_801/B 0.03fF
C56311 OR2X1_LOC_801/B VSS 0.33fF
C12245 OR2X1_LOC_512/Y OR2X1_LOC_779/B 0.08fF
C14119 AND2X1_LOC_44/Y OR2X1_LOC_512/Y 0.01fF
C17732 OR2X1_LOC_512/Y OR2X1_LOC_513/a_8_216# 0.39fF
C18847 AND2X1_LOC_41/A OR2X1_LOC_512/Y 0.03fF
C26155 AND2X1_LOC_53/Y OR2X1_LOC_512/Y 0.02fF
C29378 OR2X1_LOC_160/B OR2X1_LOC_512/Y 0.04fF
C40419 AND2X1_LOC_12/Y OR2X1_LOC_512/Y 0.02fF
C44768 OR2X1_LOC_375/A OR2X1_LOC_512/Y 0.01fF
C56362 OR2X1_LOC_512/Y VSS 0.18fF
C1329 VDD OR2X1_LOC_276/A 0.21fF
C9833 OR2X1_LOC_6/B OR2X1_LOC_276/A 0.04fF
C12097 OR2X1_LOC_276/A OR2X1_LOC_276/B 0.01fF
C12383 AND2X1_LOC_70/Y OR2X1_LOC_276/A 0.01fF
C15287 OR2X1_LOC_276/A AND2X1_LOC_275/a_8_24# 0.09fF
C21204 OR2X1_LOC_276/A AND2X1_LOC_36/Y 0.16fF
C21805 OR2X1_LOC_274/Y OR2X1_LOC_276/A 0.01fF
C40245 OR2X1_LOC_121/Y OR2X1_LOC_276/A 0.02fF
C40366 AND2X1_LOC_12/Y OR2X1_LOC_276/A 0.29fF
C45055 OR2X1_LOC_276/A OR2X1_LOC_549/A 0.03fF
C57204 OR2X1_LOC_276/A VSS 0.14fF
C5820 VDD OR2X1_LOC_86/Y 0.12fF
C15208 OR2X1_LOC_426/B OR2X1_LOC_86/Y 0.05fF
C18261 OR2X1_LOC_86/Y OR2X1_LOC_92/Y 0.01fF
C24749 OR2X1_LOC_70/Y OR2X1_LOC_86/Y 0.01fF
C26797 OR2X1_LOC_86/Y AND2X1_LOC_100/a_8_24# 0.23fF
C29747 OR2X1_LOC_86/Y OR2X1_LOC_43/A 0.09fF
C37389 OR2X1_LOC_86/Y OR2X1_LOC_19/B 0.03fF
C45477 OR2X1_LOC_86/Y OR2X1_LOC_18/Y 0.02fF
C47472 OR2X1_LOC_86/Y OR2X1_LOC_88/Y 0.08fF
C50437 OR2X1_LOC_86/Y OR2X1_LOC_86/A 0.01fF
C57450 OR2X1_LOC_86/Y VSS -0.09fF
C129 AND2X1_LOC_64/Y OR2X1_LOC_6/B 0.16fF
C154 OR2X1_LOC_6/B AND2X1_LOC_82/Y 0.02fF
C185 OR2X1_LOC_6/B AND2X1_LOC_86/a_8_24# 0.11fF
C648 OR2X1_LOC_6/B OR2X1_LOC_756/B 0.02fF
C1886 OR2X1_LOC_49/A OR2X1_LOC_6/B 0.21fF
C2038 OR2X1_LOC_6/B OR2X1_LOC_87/B 0.10fF
C2068 OR2X1_LOC_6/B AND2X1_LOC_85/a_8_24# 0.14fF
C2354 OR2X1_LOC_6/B OR2X1_LOC_671/Y 0.06fF
C2596 OR2X1_LOC_6/B OR2X1_LOC_532/B 0.09fF
C3253 OR2X1_LOC_6/B AND2X1_LOC_14/a_36_24# 0.01fF
C3738 OR2X1_LOC_185/Y OR2X1_LOC_6/B 0.10fF
C4434 OR2X1_LOC_6/B VDD 0.85fF
C4950 OR2X1_LOC_6/B OR2X1_LOC_6/a_8_216# 0.08fF
C6417 OR2X1_LOC_6/B OR2X1_LOC_80/A 0.29fF
C6556 OR2X1_LOC_104/a_8_216# OR2X1_LOC_6/B 0.09fF
C6649 OR2X1_LOC_6/B OR2X1_LOC_6/A 0.56fF
C6735 OR2X1_LOC_6/B OR2X1_LOC_611/a_36_216# 0.01fF
C7112 OR2X1_LOC_6/B OR2X1_LOC_44/Y 0.01fF
C7414 OR2X1_LOC_45/B OR2X1_LOC_6/B 1.16fF
C7527 OR2X1_LOC_160/A OR2X1_LOC_6/B 0.14fF
C7586 OR2X1_LOC_6/B AND2X1_LOC_86/B 0.61fF
C7852 OR2X1_LOC_6/B OR2X1_LOC_158/A 0.03fF
C7964 OR2X1_LOC_6/B OR2X1_LOC_847/A 0.02fF
C8457 OR2X1_LOC_6/B OR2X1_LOC_748/A 0.14fF
C8826 OR2X1_LOC_6/B OR2X1_LOC_185/A 0.14fF
C10473 OR2X1_LOC_6/B OR2X1_LOC_744/A 0.19fF
C10516 OR2X1_LOC_6/B OR2X1_LOC_541/B 0.01fF
C11184 OR2X1_LOC_6/B AND2X1_LOC_750/a_8_24# -0.03fF
C11213 AND2X1_LOC_91/B OR2X1_LOC_6/B 0.11fF
C11506 OR2X1_LOC_6/B OR2X1_LOC_751/A 0.04fF
C11724 OR2X1_LOC_6/B OR2X1_LOC_56/A 0.21fF
C11729 OR2X1_LOC_6/B OR2X1_LOC_819/a_8_216# 0.04fF
C11815 OR2X1_LOC_6/B AND2X1_LOC_56/B 0.03fF
C11827 OR2X1_LOC_6/B AND2X1_LOC_8/Y 0.12fF
C12678 OR2X1_LOC_6/B OR2X1_LOC_83/A 0.02fF
C13166 OR2X1_LOC_6/B AND2X1_LOC_85/a_36_24# 0.01fF
C13230 OR2X1_LOC_6/B AND2X1_LOC_47/Y 0.09fF
C13637 OR2X1_LOC_6/B AND2X1_LOC_5/a_36_24# 0.01fF
C13816 OR2X1_LOC_6/B OR2X1_LOC_15/a_8_216# 0.02fF
C13930 OR2X1_LOC_6/B AND2X1_LOC_95/Y 0.51fF
C14240 OR2X1_LOC_6/B AND2X1_LOC_22/Y 0.07fF
C14808 OR2X1_LOC_6/B AND2X1_LOC_490/a_8_24# 0.11fF
C15127 OR2X1_LOC_6/B OR2X1_LOC_235/B 0.07fF
C15304 OR2X1_LOC_6/B OR2X1_LOC_276/B 0.02fF
C15505 OR2X1_LOC_6/B AND2X1_LOC_70/Y 0.50fF
C16031 OR2X1_LOC_6/B OR2X1_LOC_96/B 0.03fF
C16752 OR2X1_LOC_6/B AND2X1_LOC_256/a_8_24# 0.07fF
C17178 OR2X1_LOC_6/B AND2X1_LOC_44/Y 11.35fF
C17218 OR2X1_LOC_6/B OR2X1_LOC_600/A 9.11fF
C17631 OR2X1_LOC_6/B AND2X1_LOC_628/a_8_24# 0.03fF
C18063 OR2X1_LOC_6/B AND2X1_LOC_18/Y 0.64fF
C18494 OR2X1_LOC_6/B AND2X1_LOC_275/a_8_24# 0.04fF
C19126 OR2X1_LOC_6/B OR2X1_LOC_62/B 0.30fF
C20195 OR2X1_LOC_6/B OR2X1_LOC_428/A 0.08fF
C20835 OR2X1_LOC_6/B OR2X1_LOC_54/Y 0.30fF
C20892 OR2X1_LOC_6/B OR2X1_LOC_276/a_8_216# 0.04fF
C21163 OR2X1_LOC_6/B OR2X1_LOC_161/A 0.04fF
C21205 OR2X1_LOC_6/B OR2X1_LOC_26/Y 0.03fF
C21244 OR2X1_LOC_6/B AND2X1_LOC_51/Y 0.21fF
C21966 OR2X1_LOC_6/B AND2X1_LOC_41/A 0.07fF
C22177 OR2X1_LOC_6/B OR2X1_LOC_95/Y 0.07fF
C22856 OR2X1_LOC_6/B OR2X1_LOC_820/A 0.80fF
C23116 OR2X1_LOC_6/B OR2X1_LOC_71/A 0.91fF
C23250 OR2X1_LOC_6/B OR2X1_LOC_59/Y 0.05fF
C23459 OR2X1_LOC_6/B AND2X1_LOC_14/a_8_24# 0.03fF
C23883 OR2X1_LOC_6/B OR2X1_LOC_47/Y 0.07fF
C24225 OR2X1_LOC_6/B OR2X1_LOC_8/a_8_216# 0.01fF
C24389 OR2X1_LOC_6/B AND2X1_LOC_36/Y 0.05fF
C24854 OR2X1_LOC_6/B OR2X1_LOC_16/A 0.97fF
C24925 OR2X1_LOC_6/B OR2X1_LOC_274/Y 0.01fF
C26496 OR2X1_LOC_6/B OR2X1_LOC_748/a_8_216# 0.10fF
C26965 OR2X1_LOC_6/B OR2X1_LOC_40/Y 0.06fF
C27723 OR2X1_LOC_6/B OR2X1_LOC_777/B 0.07fF
C28326 OR2X1_LOC_6/B AND2X1_LOC_398/a_8_24# 0.01fF
C28368 OR2X1_LOC_6/B OR2X1_LOC_43/A 4.64fF
C28678 OR2X1_LOC_6/B OR2X1_LOC_630/B 0.01fF
C29060 OR2X1_LOC_6/B AND2X1_LOC_625/a_8_24# 0.02fF
C29221 OR2X1_LOC_6/B OR2X1_LOC_3/Y 1.16fF
C29267 OR2X1_LOC_6/B AND2X1_LOC_133/a_8_24# 0.01fF
C29502 OR2X1_LOC_6/B AND2X1_LOC_275/a_36_24# 0.01fF
C29512 OR2X1_LOC_6/B OR2X1_LOC_671/a_8_216# 0.01fF
C29556 OR2X1_LOC_6/B OR2X1_LOC_502/A 0.08fF
C29797 OR2X1_LOC_6/B OR2X1_LOC_398/a_8_216# 0.01fF
C30071 OR2X1_LOC_6/B AND2X1_LOC_3/Y 0.49fF
C30711 OR2X1_LOC_6/B AND2X1_LOC_7/B 0.65fF
C31832 OR2X1_LOC_6/B OR2X1_LOC_473/A 0.16fF
C31996 OR2X1_LOC_6/B OR2X1_LOC_14/a_8_216# 0.03fF
C32145 OR2X1_LOC_6/B OR2X1_LOC_287/B 0.02fF
C32424 OR2X1_LOC_6/B OR2X1_LOC_160/B 0.14fF
C33071 OR2X1_LOC_6/B AND2X1_LOC_28/a_8_24# 0.03fF
C33234 OR2X1_LOC_6/B AND2X1_LOC_750/a_36_24# 0.01fF
C33282 OR2X1_LOC_6/B OR2X1_LOC_151/A 0.07fF
C34164 OR2X1_LOC_6/B AND2X1_LOC_628/a_36_24# 0.01fF
C34199 OR2X1_LOC_6/B AND2X1_LOC_62/a_8_24# 0.02fF
C35670 OR2X1_LOC_6/B OR2X1_LOC_66/a_8_216# 0.04fF
C36010 OR2X1_LOC_6/B OR2X1_LOC_19/B 0.08fF
C37214 OR2X1_LOC_126/a_8_216# OR2X1_LOC_6/B 0.03fF
C37281 OR2X1_LOC_6/B OR2X1_LOC_611/Y 0.01fF
C37468 OR2X1_LOC_6/B OR2X1_LOC_748/Y 0.02fF
C37517 OR2X1_LOC_6/B OR2X1_LOC_14/a_36_216# 0.02fF
C37603 OR2X1_LOC_6/B OR2X1_LOC_36/Y 0.04fF
C37915 OR2X1_LOC_604/A OR2X1_LOC_6/B 0.09fF
C37925 OR2X1_LOC_6/B OR2X1_LOC_66/A 0.35fF
C39277 AND2X1_LOC_40/Y OR2X1_LOC_6/B 0.10fF
C39305 OR2X1_LOC_6/B OR2X1_LOC_399/A 0.01fF
C39323 OR2X1_LOC_6/B OR2X1_LOC_87/Y 0.03fF
C40235 OR2X1_LOC_6/B AND2X1_LOC_133/a_36_24# 0.01fF
C40624 OR2X1_LOC_6/B OR2X1_LOC_73/a_8_216# 0.05fF
C40766 OR2X1_LOC_6/B OR2X1_LOC_749/a_8_216# 0.06fF
C40767 OR2X1_LOC_6/B OR2X1_LOC_398/Y 0.01fF
C41381 OR2X1_LOC_6/B AND2X1_LOC_54/a_8_24# 0.04fF
C42238 OR2X1_LOC_6/B OR2X1_LOC_78/A 0.12fF
C42869 OR2X1_LOC_6/B OR2X1_LOC_814/A 0.07fF
C43507 OR2X1_LOC_121/Y OR2X1_LOC_6/B 0.01fF
C43629 AND2X1_LOC_12/Y OR2X1_LOC_6/B 0.22fF
C44058 AND2X1_LOC_59/Y OR2X1_LOC_6/B 0.08fF
C44525 OR2X1_LOC_6/B OR2X1_LOC_585/A 0.38fF
C45387 OR2X1_LOC_6/B OR2X1_LOC_753/A 0.12fF
C45830 OR2X1_LOC_6/B OR2X1_LOC_37/a_8_216# 0.06fF
C46159 OR2X1_LOC_8/Y OR2X1_LOC_6/B 3.36fF
C46708 AND2X1_LOC_81/B OR2X1_LOC_6/B 0.04fF
C46884 OR2X1_LOC_6/B OR2X1_LOC_66/Y 0.01fF
C47151 OR2X1_LOC_6/B OR2X1_LOC_39/A 2.65fF
C47604 OR2X1_LOC_6/B OR2X1_LOC_377/A 0.05fF
C47626 OR2X1_LOC_6/B OR2X1_LOC_85/A 0.19fF
C47954 OR2X1_LOC_6/B OR2X1_LOC_51/Y 0.05fF
C47968 OR2X1_LOC_6/B OR2X1_LOC_78/B 0.13fF
C48051 OR2X1_LOC_6/B OR2X1_LOC_375/A 0.17fF
C48369 OR2X1_LOC_6/B OR2X1_LOC_549/A 0.89fF
C49178 OR2X1_LOC_6/B AND2X1_LOC_65/A 0.16fF
C49286 AND2X1_LOC_381/a_8_24# OR2X1_LOC_6/B 0.26fF
C49868 OR2X1_LOC_6/B AND2X1_LOC_28/a_36_24# 0.01fF
C50276 OR2X1_LOC_6/B OR2X1_LOC_4/a_8_216# 0.06fF
C51395 OR2X1_LOC_6/B OR2X1_LOC_32/B 0.03fF
C51598 OR2X1_LOC_6/B OR2X1_LOC_68/B 2.20fF
C51885 OR2X1_LOC_6/B OR2X1_LOC_74/A 0.07fF
C52250 OR2X1_LOC_6/B OR2X1_LOC_87/A 0.07fF
C52278 OR2X1_LOC_6/B AND2X1_LOC_19/a_8_24# 0.03fF
C52631 OR2X1_LOC_6/B OR2X1_LOC_23/a_8_216# 0.22fF
C53203 OR2X1_LOC_6/B AND2X1_LOC_5/a_8_24# 0.02fF
C53812 OR2X1_LOC_126/a_36_216# OR2X1_LOC_6/B 0.03fF
C54765 OR2X1_LOC_154/A OR2X1_LOC_6/B 0.10fF
C56106 OR2X1_LOC_6/B OR2X1_LOC_827/Y 0.02fF
C57890 OR2X1_LOC_6/B VSS 1.05fF
C144 OR2X1_LOC_6/A OR2X1_LOC_80/A 0.14fF
C915 OR2X1_LOC_45/B OR2X1_LOC_80/A 0.05fF
C1030 OR2X1_LOC_160/A OR2X1_LOC_80/A 0.06fF
C1061 AND2X1_LOC_86/B OR2X1_LOC_80/A 0.27fF
C1449 OR2X1_LOC_847/A OR2X1_LOC_80/A 0.03fF
C1462 AND2X1_LOC_278/a_36_24# OR2X1_LOC_80/A 0.01fF
C2310 OR2X1_LOC_185/A OR2X1_LOC_80/A 0.15fF
C3969 OR2X1_LOC_744/A OR2X1_LOC_80/A 0.23fF
C4319 OR2X1_LOC_129/a_8_216# OR2X1_LOC_80/A 0.01fF
C4687 AND2X1_LOC_91/B OR2X1_LOC_80/A 0.12fF
C5209 AND2X1_LOC_56/B OR2X1_LOC_80/A 0.08fF
C5217 AND2X1_LOC_8/Y OR2X1_LOC_80/A 0.07fF
C5401 OR2X1_LOC_80/A AND2X1_LOC_236/a_8_24# 0.02fF
C5694 OR2X1_LOC_291/Y OR2X1_LOC_80/A 0.07fF
C6088 OR2X1_LOC_83/A OR2X1_LOC_80/A 0.29fF
C6589 AND2X1_LOC_47/Y OR2X1_LOC_80/A 0.23fF
C7463 OR2X1_LOC_415/a_8_216# OR2X1_LOC_80/A 0.06fF
C8309 AND2X1_LOC_817/a_8_24# OR2X1_LOC_80/A 0.02fF
C8687 OR2X1_LOC_235/B OR2X1_LOC_80/A 0.11fF
C10757 OR2X1_LOC_600/A OR2X1_LOC_80/A 0.50fF
C11591 AND2X1_LOC_18/Y OR2X1_LOC_80/A 0.06fF
C12568 OR2X1_LOC_62/B OR2X1_LOC_80/A 0.05fF
C14280 OR2X1_LOC_54/Y OR2X1_LOC_80/A 0.10fF
C14662 OR2X1_LOC_26/Y OR2X1_LOC_80/A 0.72fF
C16304 OR2X1_LOC_847/a_8_216# OR2X1_LOC_80/A 0.02fF
C16501 OR2X1_LOC_80/A OR2X1_LOC_71/A 0.05fF
C16679 OR2X1_LOC_59/Y OR2X1_LOC_80/A 0.04fF
C16853 AND2X1_LOC_14/a_8_24# OR2X1_LOC_80/A 0.02fF
C17192 OR2X1_LOC_240/A OR2X1_LOC_80/A 0.08fF
C17285 OR2X1_LOC_47/Y OR2X1_LOC_80/A 0.40fF
C17818 AND2X1_LOC_36/Y OR2X1_LOC_80/A 0.15fF
C18368 OR2X1_LOC_16/A OR2X1_LOC_80/A 5.77fF
C19326 OR2X1_LOC_847/B OR2X1_LOC_80/A 0.05fF
C19653 OR2X1_LOC_80/A OR2X1_LOC_548/a_8_216# 0.05fF
C20198 OR2X1_LOC_269/B OR2X1_LOC_80/A 0.09fF
C20533 OR2X1_LOC_40/Y OR2X1_LOC_80/A 0.01fF
C21041 AND2X1_LOC_42/a_8_24# OR2X1_LOC_80/A 0.09fF
C21813 OR2X1_LOC_589/A OR2X1_LOC_80/A 0.11fF
C21872 AND2X1_LOC_618/a_8_24# OR2X1_LOC_80/A 0.11fF
C22823 OR2X1_LOC_3/Y OR2X1_LOC_80/A 0.03fF
C22892 OR2X1_LOC_673/A OR2X1_LOC_80/A 0.05fF
C23145 OR2X1_LOC_502/A OR2X1_LOC_80/A 0.10fF
C23338 OR2X1_LOC_80/A OR2X1_LOC_398/a_8_216# 0.21fF
C23506 AND2X1_LOC_530/a_8_24# OR2X1_LOC_80/A 0.05fF
C23581 AND2X1_LOC_104/a_8_24# OR2X1_LOC_80/A 0.04fF
C26575 AND2X1_LOC_28/a_8_24# OR2X1_LOC_80/A 0.04fF
C27335 AND2X1_LOC_619/B OR2X1_LOC_80/A 0.02fF
C28080 OR2X1_LOC_415/Y OR2X1_LOC_80/A 0.04fF
C28943 OR2X1_LOC_548/A OR2X1_LOC_80/A 0.05fF
C29362 AND2X1_LOC_90/a_8_24# OR2X1_LOC_80/A 0.06fF
C29524 OR2X1_LOC_19/B OR2X1_LOC_80/A 0.37fF
C31167 OR2X1_LOC_36/Y OR2X1_LOC_80/A 0.16fF
C31511 OR2X1_LOC_66/A OR2X1_LOC_80/A 1.47fF
C31920 AND2X1_LOC_94/Y OR2X1_LOC_80/A 0.02fF
C32796 AND2X1_LOC_40/Y OR2X1_LOC_80/A 0.03fF
C32810 OR2X1_LOC_399/A OR2X1_LOC_80/A 0.02fF
C32832 OR2X1_LOC_848/A OR2X1_LOC_80/A 0.61fF
C34337 AND2X1_LOC_619/a_8_24# OR2X1_LOC_80/A 0.01fF
C34927 AND2X1_LOC_54/a_8_24# OR2X1_LOC_80/A 0.03fF
C35734 OR2X1_LOC_78/A OR2X1_LOC_80/A 0.10fF
C37020 AND2X1_LOC_12/Y OR2X1_LOC_80/A 0.75fF
C37893 OR2X1_LOC_585/A OR2X1_LOC_80/A 0.10fF
C38771 OR2X1_LOC_753/A OR2X1_LOC_80/A 0.10fF
C39210 OR2X1_LOC_37/a_8_216# OR2X1_LOC_80/A 0.47fF
C39875 OR2X1_LOC_622/B OR2X1_LOC_80/A 0.01fF
C40003 AND2X1_LOC_49/a_8_24# OR2X1_LOC_80/A 0.05fF
C40343 AND2X1_LOC_90/a_36_24# OR2X1_LOC_80/A 0.01fF
C40434 OR2X1_LOC_39/A OR2X1_LOC_80/A 0.76fF
C40842 AND2X1_LOC_278/a_8_24# OR2X1_LOC_80/A 0.17fF
C40845 OR2X1_LOC_377/A OR2X1_LOC_80/A 12.76fF
C40857 OR2X1_LOC_85/A OR2X1_LOC_80/A 0.09fF
C41247 OR2X1_LOC_78/B OR2X1_LOC_80/A 2.46fF
C41297 OR2X1_LOC_375/A OR2X1_LOC_80/A 0.03fF
C41667 OR2X1_LOC_80/A OR2X1_LOC_549/A 0.05fF
C42632 AND2X1_LOC_381/a_8_24# OR2X1_LOC_80/A 0.02fF
C43575 OR2X1_LOC_4/a_8_216# OR2X1_LOC_80/A -0.03fF
C44773 OR2X1_LOC_32/B OR2X1_LOC_80/A 1.04fF
C44971 OR2X1_LOC_68/B OR2X1_LOC_80/A 1.66fF
C46629 AND2X1_LOC_5/a_8_24# OR2X1_LOC_80/A 0.01fF
C49506 OR2X1_LOC_633/A OR2X1_LOC_80/A 1.43fF
C51352 OR2X1_LOC_80/a_8_216# OR2X1_LOC_80/A 0.02fF
C51573 OR2X1_LOC_49/A OR2X1_LOC_80/A 0.10fF
C51713 AND2X1_LOC_612/B OR2X1_LOC_80/A 0.15fF
C51722 AND2X1_LOC_85/a_8_24# OR2X1_LOC_80/A 0.02fF
C52171 OR2X1_LOC_532/B OR2X1_LOC_80/A 0.46fF
C54137 VDD OR2X1_LOC_80/A 0.47fF
C56408 OR2X1_LOC_80/A VSS -3.61fF
C3395 VDD OR2X1_LOC_291/A 0.03fF
C6687 OR2X1_LOC_158/A OR2X1_LOC_291/A 0.02fF
C9046 OR2X1_LOC_824/a_8_216# OR2X1_LOC_291/A 0.01fF
C14064 OR2X1_LOC_235/B OR2X1_LOC_291/A 0.05fF
C16173 OR2X1_LOC_291/A OR2X1_LOC_619/Y 0.40fF
C17965 OR2X1_LOC_62/B OR2X1_LOC_291/A 0.03fF
C19699 OR2X1_LOC_291/A OR2X1_LOC_54/Y 0.11fF
C20075 OR2X1_LOC_291/A OR2X1_LOC_26/Y 0.01fF
C20943 OR2X1_LOC_291/A OR2X1_LOC_824/Y 0.02fF
C21944 OR2X1_LOC_291/A OR2X1_LOC_71/A 0.08fF
C22777 OR2X1_LOC_291/A OR2X1_LOC_47/Y 1.93fF
C25846 OR2X1_LOC_40/Y OR2X1_LOC_291/A 0.06fF
C33697 OR2X1_LOC_291/A OR2X1_LOC_234/a_8_216# 0.39fF
C36511 OR2X1_LOC_36/Y OR2X1_LOC_291/A 0.56fF
C40683 OR2X1_LOC_291/A OR2X1_LOC_234/Y 0.03fF
C40792 OR2X1_LOC_291/A OR2X1_LOC_278/A 0.19fF
C41609 OR2X1_LOC_291/a_8_216# OR2X1_LOC_291/A 0.05fF
C43390 OR2X1_LOC_291/A OR2X1_LOC_585/A 0.04fF
C44260 OR2X1_LOC_291/A OR2X1_LOC_753/A 0.08fF
C45010 OR2X1_LOC_8/Y OR2X1_LOC_291/A 0.36fF
C46452 OR2X1_LOC_291/A OR2X1_LOC_85/A 0.05fF
C50376 OR2X1_LOC_233/a_8_216# OR2X1_LOC_291/A -0.00fF
C50785 OR2X1_LOC_291/A OR2X1_LOC_74/A 0.03fF
C57145 OR2X1_LOC_291/A VSS 0.75fF
C4347 OR2X1_LOC_413/Y AND2X1_LOC_461/a_8_24# 0.01fF
C7671 OR2X1_LOC_413/Y OR2X1_LOC_7/A 0.14fF
C9944 OR2X1_LOC_413/Y AND2X1_LOC_462/B 0.79fF
C11067 OR2X1_LOC_413/Y OR2X1_LOC_690/A 0.09fF
C25804 OR2X1_LOC_411/Y OR2X1_LOC_413/Y 0.21fF
C27273 OR2X1_LOC_22/Y OR2X1_LOC_413/Y 0.06fF
C41006 VDD OR2X1_LOC_413/Y 0.04fF
C43755 OR2X1_LOC_413/Y OR2X1_LOC_44/Y 0.03fF
C57219 OR2X1_LOC_413/Y VSS 0.02fF
C5731 OR2X1_LOC_691/A OR2X1_LOC_377/A 0.01fF
C18912 OR2X1_LOC_691/A VDD 0.21fF
C21986 OR2X1_LOC_691/A OR2X1_LOC_160/A 0.03fF
C36344 OR2X1_LOC_691/A OR2X1_LOC_688/a_8_216# 0.01fF
C37770 OR2X1_LOC_691/A AND2X1_LOC_31/Y 0.03fF
C38699 OR2X1_LOC_691/A AND2X1_LOC_36/Y 0.07fF
C40986 OR2X1_LOC_691/A OR2X1_LOC_269/B 0.02fF
C41379 OR2X1_LOC_691/A AND2X1_LOC_690/a_8_24# 0.01fF
C42290 OR2X1_LOC_691/A AND2X1_LOC_824/a_8_24# 0.20fF
C47467 OR2X1_LOC_691/A OR2X1_LOC_691/B 0.61fF
C50629 OR2X1_LOC_691/A OR2X1_LOC_19/B 0.03fF
C52565 OR2X1_LOC_691/A OR2X1_LOC_66/A 0.79fF
C55249 OR2X1_LOC_691/A AND2X1_LOC_689/a_8_24# 0.01fF
C57978 OR2X1_LOC_691/A VSS 0.30fF
C606 OR2X1_LOC_151/A AND2X1_LOC_110/Y 0.05fF
C611 AND2X1_LOC_322/a_8_24# AND2X1_LOC_110/Y 0.01fF
C3632 AND2X1_LOC_534/a_8_24# AND2X1_LOC_110/Y 0.01fF
C5266 AND2X1_LOC_110/Y OR2X1_LOC_66/A 0.03fF
C6125 OR2X1_LOC_325/B AND2X1_LOC_110/Y 0.01fF
C9155 OR2X1_LOC_535/A AND2X1_LOC_110/Y 0.01fF
C9171 AND2X1_LOC_110/Y AND2X1_LOC_323/a_8_24# 0.09fF
C9624 AND2X1_LOC_110/Y OR2X1_LOC_78/A 0.03fF
C9738 AND2X1_LOC_110/Y OR2X1_LOC_155/A 0.03fF
C11359 AND2X1_LOC_59/Y AND2X1_LOC_110/Y 0.03fF
C15122 AND2X1_LOC_110/Y OR2X1_LOC_78/B 0.03fF
C16874 OR2X1_LOC_405/A AND2X1_LOC_110/Y 0.03fF
C21589 AND2X1_LOC_110/Y AND2X1_LOC_527/a_8_24# 0.08fF
C22050 OR2X1_LOC_154/A AND2X1_LOC_110/Y 0.03fF
C22374 AND2X1_LOC_110/Y AND2X1_LOC_299/a_8_24# 0.01fF
C22970 AND2X1_LOC_110/Y AND2X1_LOC_111/a_8_24# 0.09fF
C23586 AND2X1_LOC_64/Y AND2X1_LOC_110/Y 0.39fF
C25909 AND2X1_LOC_110/Y OR2X1_LOC_532/B 0.03fF
C27105 OR2X1_LOC_185/Y AND2X1_LOC_110/Y 0.02fF
C27817 AND2X1_LOC_110/Y OR2X1_LOC_302/A 0.01fF
C27827 VDD AND2X1_LOC_110/Y 0.39fF
C30798 OR2X1_LOC_809/B AND2X1_LOC_110/Y 0.02fF
C30875 OR2X1_LOC_160/A AND2X1_LOC_110/Y 0.03fF
C31255 OR2X1_LOC_325/A AND2X1_LOC_110/Y 0.01fF
C32078 OR2X1_LOC_185/A AND2X1_LOC_110/Y 0.03fF
C34499 AND2X1_LOC_91/B AND2X1_LOC_110/Y 0.03fF
C34918 AND2X1_LOC_110/Y OR2X1_LOC_446/B 0.03fF
C35092 AND2X1_LOC_110/Y AND2X1_LOC_56/B 0.05fF
C36461 AND2X1_LOC_110/Y AND2X1_LOC_47/Y 0.03fF
C36718 AND2X1_LOC_110/Y OR2X1_LOC_506/A 0.03fF
C37155 AND2X1_LOC_95/Y AND2X1_LOC_110/Y 0.07fF
C38822 AND2X1_LOC_70/Y AND2X1_LOC_110/Y 0.04fF
C40454 AND2X1_LOC_110/Y AND2X1_LOC_44/Y 0.03fF
C44477 AND2X1_LOC_110/Y OR2X1_LOC_161/A 0.06fF
C44574 AND2X1_LOC_110/Y AND2X1_LOC_51/Y 0.03fF
C46919 AND2X1_LOC_110/Y AND2X1_LOC_31/Y 0.04fF
C50176 AND2X1_LOC_110/Y OR2X1_LOC_269/B 0.03fF
C51225 AND2X1_LOC_110/Y OR2X1_LOC_777/B 0.02fF
C51710 AND2X1_LOC_110/Y OR2X1_LOC_161/B 0.48fF
C53066 AND2X1_LOC_110/Y OR2X1_LOC_502/A 0.07fF
C55977 OR2X1_LOC_160/B AND2X1_LOC_110/Y 0.26fF
C57606 AND2X1_LOC_110/Y VSS 0.19fF
C1005 AND2X1_LOC_514/Y OR2X1_LOC_22/Y 0.07fF
C2136 AND2X1_LOC_514/Y OR2X1_LOC_51/Y 0.02fF
C5058 AND2X1_LOC_514/Y OR2X1_LOC_91/A 0.02fF
C8677 AND2X1_LOC_514/Y OR2X1_LOC_417/a_8_216# 0.03fF
C14873 VDD AND2X1_LOC_514/Y 0.72fF
C17081 AND2X1_LOC_514/Y OR2X1_LOC_6/A 0.01fF
C17495 AND2X1_LOC_514/Y OR2X1_LOC_44/Y 0.07fF
C18251 OR2X1_LOC_158/A AND2X1_LOC_514/Y 0.07fF
C19707 AND2X1_LOC_514/Y OR2X1_LOC_417/a_36_216# 0.01fF
C20867 AND2X1_LOC_514/Y OR2X1_LOC_744/A 0.07fF
C22166 AND2X1_LOC_514/Y OR2X1_LOC_56/A 0.09fF
C22745 OR2X1_LOC_417/Y AND2X1_LOC_514/Y 0.23fF
C24270 AND2X1_LOC_514/Y OR2X1_LOC_426/B 0.07fF
C27241 AND2X1_LOC_514/Y OR2X1_LOC_92/Y 0.07fF
C27585 AND2X1_LOC_514/Y OR2X1_LOC_600/A 0.07fF
C30476 AND2X1_LOC_514/Y OR2X1_LOC_428/A 0.07fF
C32362 AND2X1_LOC_514/Y OR2X1_LOC_95/Y 0.19fF
C34106 AND2X1_LOC_514/Y OR2X1_LOC_47/Y 0.08fF
C37261 OR2X1_LOC_40/Y AND2X1_LOC_514/Y 0.08fF
C37406 AND2X1_LOC_514/Y OR2X1_LOC_7/A 0.07fF
C39871 OR2X1_LOC_329/B AND2X1_LOC_514/Y 0.46fF
C40806 AND2X1_LOC_514/Y OR2X1_LOC_64/Y 0.02fF
C48257 AND2X1_LOC_514/Y OR2X1_LOC_36/Y 0.05fF
C48563 OR2X1_LOC_604/A AND2X1_LOC_514/Y 0.10fF
C55555 AND2X1_LOC_514/Y OR2X1_LOC_437/A 0.01fF
C57620 AND2X1_LOC_514/Y VSS -1.44fF
C821 OR2X1_LOC_160/B OR2X1_LOC_750/A 0.03fF
C4360 OR2X1_LOC_19/B OR2X1_LOC_750/A 0.05fF
C6296 OR2X1_LOC_750/A OR2X1_LOC_66/A 0.03fF
C11197 OR2X1_LOC_750/A OR2X1_LOC_814/A 0.09fF
C11961 AND2X1_LOC_12/Y OR2X1_LOC_750/A 0.03fF
C12413 AND2X1_LOC_59/Y OR2X1_LOC_750/A 5.93fF
C15759 OR2X1_LOC_377/A OR2X1_LOC_750/A 0.02fF
C16147 OR2X1_LOC_750/A OR2X1_LOC_78/B 0.01fF
C17542 AND2X1_LOC_23/a_8_24# OR2X1_LOC_750/A 0.08fF
C19812 OR2X1_LOC_750/A OR2X1_LOC_68/B 0.04fF
C22301 OR2X1_LOC_750/A OR2X1_LOC_750/a_8_216# 0.02fF
C23092 OR2X1_LOC_154/A OR2X1_LOC_750/A 0.07fF
C25111 OR2X1_LOC_756/B OR2X1_LOC_750/A 0.07fF
C26627 OR2X1_LOC_750/A OR2X1_LOC_333/A 0.03fF
C28843 VDD OR2X1_LOC_750/A 0.25fF
C38202 AND2X1_LOC_95/Y OR2X1_LOC_750/A 0.03fF
C38491 AND2X1_LOC_22/Y OR2X1_LOC_750/A 0.03fF
C41503 OR2X1_LOC_750/A AND2X1_LOC_44/Y 0.06fF
C42456 OR2X1_LOC_750/A AND2X1_LOC_18/Y 0.09fF
C45558 OR2X1_LOC_750/A OR2X1_LOC_161/A 0.17fF
C46405 AND2X1_LOC_41/A OR2X1_LOC_750/A 0.01fF
C47765 AND2X1_LOC_749/a_8_24# OR2X1_LOC_750/A 0.01fF
C51191 OR2X1_LOC_750/A OR2X1_LOC_269/B 0.01fF
C55243 OR2X1_LOC_750/A AND2X1_LOC_7/B 0.01fF
C56893 OR2X1_LOC_750/A VSS -0.10fF
C35 OR2X1_LOC_814/Y OR2X1_LOC_814/A 0.01fF
C323 OR2X1_LOC_814/A OR2X1_LOC_227/A 0.01fF
C503 OR2X1_LOC_814/A OR2X1_LOC_269/B 0.11fF
C1562 OR2X1_LOC_814/A OR2X1_LOC_777/B 0.07fF
C1630 OR2X1_LOC_814/A OR2X1_LOC_831/B 0.07fF
C2087 OR2X1_LOC_814/A OR2X1_LOC_161/B 0.03fF
C3473 OR2X1_LOC_502/A OR2X1_LOC_814/A 0.13fF
C3583 AND2X1_LOC_48/A OR2X1_LOC_814/A 0.09fF
C3809 OR2X1_LOC_814/A OR2X1_LOC_489/A 0.01fF
C3966 AND2X1_LOC_3/Y OR2X1_LOC_814/A 0.22fF
C4574 OR2X1_LOC_814/A AND2X1_LOC_7/B 0.45fF
C6023 OR2X1_LOC_287/B OR2X1_LOC_814/A 0.06fF
C6303 OR2X1_LOC_160/B OR2X1_LOC_814/A 17.61fF
C7183 OR2X1_LOC_151/A OR2X1_LOC_814/A 0.07fF
C11914 OR2X1_LOC_814/A OR2X1_LOC_66/A 2.38fF
C13283 AND2X1_LOC_40/Y OR2X1_LOC_814/A 2.78fF
C16158 OR2X1_LOC_814/A OR2X1_LOC_78/A 0.15fF
C16248 OR2X1_LOC_814/A OR2X1_LOC_155/A 0.03fF
C16668 OR2X1_LOC_814/A OR2X1_LOC_68/a_8_216# 0.03fF
C17488 AND2X1_LOC_12/Y OR2X1_LOC_814/A 1.72fF
C17924 AND2X1_LOC_59/Y OR2X1_LOC_814/A 0.17fF
C20439 AND2X1_LOC_310/a_8_24# OR2X1_LOC_814/A 0.01fF
C20522 AND2X1_LOC_81/B OR2X1_LOC_814/A 0.03fF
C21751 OR2X1_LOC_814/A OR2X1_LOC_78/B 0.33fF
C21819 OR2X1_LOC_375/A OR2X1_LOC_814/A 0.51fF
C22133 OR2X1_LOC_814/A OR2X1_LOC_549/A 0.15fF
C22268 OR2X1_LOC_814/A OR2X1_LOC_68/a_36_216# 0.01fF
C22995 OR2X1_LOC_814/A AND2X1_LOC_65/A 0.07fF
C23501 OR2X1_LOC_405/A OR2X1_LOC_814/A 0.01fF
C25321 OR2X1_LOC_814/A OR2X1_LOC_68/B 0.09fF
C26005 OR2X1_LOC_87/A OR2X1_LOC_814/A 0.82fF
C27535 OR2X1_LOC_814/A AND2X1_LOC_417/a_8_24# -0.01fF
C28548 OR2X1_LOC_154/A OR2X1_LOC_814/A 0.32fF
C28818 OR2X1_LOC_814/A OR2X1_LOC_435/A 0.04fF
C30060 AND2X1_LOC_64/Y OR2X1_LOC_814/A 0.18fF
C30583 OR2X1_LOC_756/B OR2X1_LOC_814/A 2.44fF
C31606 OR2X1_LOC_814/A AND2X1_LOC_289/a_8_24# 0.11fF
C31986 OR2X1_LOC_814/A OR2X1_LOC_374/Y 0.07fF
C32097 OR2X1_LOC_814/A OR2X1_LOC_333/A 0.37fF
C32367 OR2X1_LOC_532/B OR2X1_LOC_814/A 0.13fF
C33637 OR2X1_LOC_185/Y OR2X1_LOC_814/A 2.28fF
C33994 OR2X1_LOC_814/a_8_216# OR2X1_LOC_814/A 0.07fF
C34326 VDD OR2X1_LOC_814/A 2.61fF
C37377 OR2X1_LOC_160/A OR2X1_LOC_814/A 0.10fF
C38654 OR2X1_LOC_185/A OR2X1_LOC_814/A 0.05fF
C40741 OR2X1_LOC_264/Y OR2X1_LOC_814/A 0.06fF
C41043 AND2X1_LOC_91/B OR2X1_LOC_814/A 0.46fF
C42678 OR2X1_LOC_814/A AND2X1_LOC_289/a_36_24# 0.02fF
C43046 OR2X1_LOC_68/Y OR2X1_LOC_814/A 0.01fF
C43059 AND2X1_LOC_47/Y OR2X1_LOC_814/A 0.25fF
C43830 AND2X1_LOC_95/Y OR2X1_LOC_814/A 0.17fF
C44115 AND2X1_LOC_22/Y OR2X1_LOC_814/A 0.28fF
C44272 AND2X1_LOC_153/a_8_24# OR2X1_LOC_814/A 0.03fF
C45082 OR2X1_LOC_235/B OR2X1_LOC_814/A 0.03fF
C45391 OR2X1_LOC_814/A AND2X1_LOC_226/a_8_24# 0.07fF
C45495 AND2X1_LOC_70/Y OR2X1_LOC_814/A 0.14fF
C47240 OR2X1_LOC_814/A AND2X1_LOC_44/Y 0.03fF
C48173 OR2X1_LOC_814/A AND2X1_LOC_18/Y 0.67fF
C49068 OR2X1_LOC_130/A OR2X1_LOC_814/A 0.19fF
C49126 OR2X1_LOC_62/B OR2X1_LOC_814/A 0.03fF
C51167 OR2X1_LOC_814/A OR2X1_LOC_161/A 0.02fF
C51227 OR2X1_LOC_814/A AND2X1_LOC_51/Y 2.15fF
C51968 AND2X1_LOC_41/A OR2X1_LOC_814/A 0.10fF
C53447 AND2X1_LOC_31/Y OR2X1_LOC_814/A 0.77fF
C54325 OR2X1_LOC_814/A AND2X1_LOC_36/Y 0.02fF
C54417 OR2X1_LOC_814/A AND2X1_LOC_488/a_8_24# 0.01fF
C55888 OR2X1_LOC_557/A OR2X1_LOC_814/A 0.06fF
C56834 OR2X1_LOC_814/A VSS 0.82fF
C605 OR2X1_LOC_49/A OR2X1_LOC_56/A 1.94fF
C688 OR2X1_LOC_49/A AND2X1_LOC_56/B 0.07fF
C697 OR2X1_LOC_49/A AND2X1_LOC_8/Y 0.62fF
C1582 OR2X1_LOC_49/A OR2X1_LOC_83/A 0.03fF
C2111 OR2X1_LOC_49/A AND2X1_LOC_47/Y 0.10fF
C2328 OR2X1_LOC_49/A OR2X1_LOC_672/a_8_216# 0.01fF
C2434 OR2X1_LOC_49/A AND2X1_LOC_129/a_8_24# 0.03fF
C2504 OR2X1_LOC_49/A OR2X1_LOC_481/A 0.42fF
C2745 OR2X1_LOC_49/A OR2X1_LOC_15/a_8_216# 0.01fF
C2834 OR2X1_LOC_49/A AND2X1_LOC_414/a_8_24# 0.03fF
C2844 OR2X1_LOC_49/A AND2X1_LOC_95/Y 0.02fF
C4059 OR2X1_LOC_49/A OR2X1_LOC_235/B 0.11fF
C4904 OR2X1_LOC_49/A OR2X1_LOC_96/B 0.21fF
C5633 OR2X1_LOC_49/A OR2X1_LOC_414/Y 0.01fF
C6057 OR2X1_LOC_49/A AND2X1_LOC_44/Y 0.84fF
C6094 OR2X1_LOC_49/A OR2X1_LOC_600/A 0.59fF
C6616 OR2X1_LOC_49/A AND2X1_LOC_818/a_8_24# 0.03fF
C7200 OR2X1_LOC_49/A AND2X1_LOC_672/a_8_24# 0.04fF
C7396 OR2X1_LOC_49/A OR2X1_LOC_133/a_8_216# 0.01fF
C8043 OR2X1_LOC_49/A OR2X1_LOC_62/B 0.03fF
C9118 OR2X1_LOC_49/A OR2X1_LOC_428/A 0.22fF
C9759 OR2X1_LOC_49/A OR2X1_LOC_54/Y 0.60fF
C10117 OR2X1_LOC_49/A OR2X1_LOC_89/A 0.07fF
C11026 OR2X1_LOC_49/A OR2X1_LOC_95/Y 0.02fF
C11800 OR2X1_LOC_49/A AND2X1_LOC_102/a_8_24# 0.04fF
C11973 OR2X1_LOC_49/A OR2X1_LOC_71/A 0.19fF
C12198 OR2X1_LOC_49/A OR2X1_LOC_820/B 0.03fF
C12647 OR2X1_LOC_49/A OR2X1_LOC_240/A 0.07fF
C12773 OR2X1_LOC_49/A OR2X1_LOC_47/Y 0.07fF
C13330 OR2X1_LOC_49/A AND2X1_LOC_36/Y 0.17fF
C13793 OR2X1_LOC_49/A OR2X1_LOC_16/A 0.10fF
C15882 OR2X1_LOC_49/A OR2X1_LOC_159/a_8_216# 0.04fF
C15978 OR2X1_LOC_49/A OR2X1_LOC_618/a_8_216# 0.18fF
C16393 OR2X1_LOC_49/A OR2X1_LOC_236/a_8_216# 0.13fF
C16727 OR2X1_LOC_49/A AND2X1_LOC_415/a_8_24# 0.04fF
C17267 OR2X1_LOC_49/A OR2X1_LOC_87/a_8_216# 0.02fF
C17290 OR2X1_LOC_49/A OR2X1_LOC_43/A 0.91fF
C18177 OR2X1_LOC_49/A OR2X1_LOC_3/Y 0.32fF
C18280 OR2X1_LOC_49/A OR2X1_LOC_673/A 0.05fF
C18527 OR2X1_LOC_49/A OR2X1_LOC_502/A 8.26fF
C19497 OR2X1_LOC_49/A OR2X1_LOC_606/a_8_216# 0.11fF
C19726 OR2X1_LOC_49/A AND2X1_LOC_7/B 0.07fF
C19998 OR2X1_LOC_49/A OR2X1_LOC_55/a_8_216# 0.03fF
C20799 OR2X1_LOC_49/A OR2X1_LOC_77/a_8_216# 0.01fF
C21176 OR2X1_LOC_49/A OR2X1_LOC_287/B 0.03fF
C22911 OR2X1_LOC_49/A OR2X1_LOC_827/a_8_216# 0.04fF
C23558 OR2X1_LOC_49/A OR2X1_LOC_415/Y 0.14fF
C24139 OR2X1_LOC_49/A OR2X1_LOC_49/a_8_216# 0.06fF
C24505 OR2X1_LOC_49/A AND2X1_LOC_80/a_8_24# 0.03fF
C24927 OR2X1_LOC_49/A OR2X1_LOC_38/a_8_216# 0.03fF
C25013 OR2X1_LOC_49/A OR2X1_LOC_19/B 0.20fF
C25019 OR2X1_LOC_49/A OR2X1_LOC_606/a_36_216# 0.03fF
C26948 OR2X1_LOC_49/A OR2X1_LOC_604/A 0.09fF
C26953 OR2X1_LOC_49/A OR2X1_LOC_66/A 0.05fF
C27388 OR2X1_LOC_49/A AND2X1_LOC_94/Y -0.01fF
C28266 OR2X1_LOC_49/A AND2X1_LOC_40/Y 0.02fF
C28324 OR2X1_LOC_49/A OR2X1_LOC_87/Y 0.01fF
C28638 OR2X1_LOC_49/A OR2X1_LOC_90/a_8_216# 0.01fF
C29601 OR2X1_LOC_49/A OR2X1_LOC_73/a_8_216# 0.01fF
C30303 OR2X1_LOC_49/A OR2X1_LOC_12/Y 0.01fF
C30402 OR2X1_LOC_49/A OR2X1_LOC_38/a_36_216# 0.02fF
C30494 OR2X1_LOC_49/A OR2X1_LOC_606/Y 0.02fF
C31195 OR2X1_LOC_49/A OR2X1_LOC_78/A 0.07fF
C32923 OR2X1_LOC_49/A AND2X1_LOC_59/Y 0.03fF
C33389 OR2X1_LOC_49/A OR2X1_LOC_585/A 0.45fF
C34208 OR2X1_LOC_49/A OR2X1_LOC_753/A 0.06fF
C34988 OR2X1_LOC_49/A OR2X1_LOC_8/Y 0.19fF
C35067 OR2X1_LOC_49/A OR2X1_LOC_672/Y 0.01fF
C35289 OR2X1_LOC_49/A OR2X1_LOC_622/B 0.01fF
C35333 OR2X1_LOC_49/A OR2X1_LOC_9/a_8_216# 0.02fF
C35882 OR2X1_LOC_49/A OR2X1_LOC_39/A 0.01fF
C36289 OR2X1_LOC_49/A OR2X1_LOC_377/A 0.10fF
C36312 OR2X1_LOC_49/A OR2X1_LOC_85/A 0.33fF
C36639 OR2X1_LOC_49/A OR2X1_LOC_78/B 0.05fF
C36693 OR2X1_LOC_49/A OR2X1_LOC_375/A 0.14fF
C38313 OR2X1_LOC_49/A OR2X1_LOC_382/a_8_216# 0.05fF
C38539 OR2X1_LOC_49/A OR2X1_LOC_416/A 0.09fF
C38568 OR2X1_LOC_49/A AND2X1_LOC_8/a_8_24# 0.01fF
C38798 OR2X1_LOC_49/A AND2X1_LOC_19/Y 0.10fF
C39650 OR2X1_LOC_49/A OR2X1_LOC_91/A 0.13fF
C40315 OR2X1_LOC_49/A OR2X1_LOC_68/B 2.63fF
C40591 OR2X1_LOC_49/A OR2X1_LOC_74/A 0.09fF
C40963 OR2X1_LOC_49/A AND2X1_LOC_80/a_36_24# 0.01fF
C40968 OR2X1_LOC_49/A OR2X1_LOC_87/A 0.71fF
C41000 OR2X1_LOC_49/A AND2X1_LOC_19/a_8_24# 0.02fF
C41298 OR2X1_LOC_49/A OR2X1_LOC_381/a_8_216# 0.01fF
C41422 OR2X1_LOC_49/A AND2X1_LOC_29/a_8_24# 0.12fF
C42307 OR2X1_LOC_49/A OR2X1_LOC_699/a_8_216# 0.01fF
C44400 OR2X1_LOC_49/A OR2X1_LOC_634/A 0.01fF
C44449 OR2X1_LOC_49/A OR2X1_LOC_94/a_8_216# 0.03fF
C44772 OR2X1_LOC_49/A OR2X1_LOC_633/A 0.27fF
C44920 OR2X1_LOC_49/A OR2X1_LOC_827/Y 0.81fF
C45190 OR2X1_LOC_49/A AND2X1_LOC_64/Y 0.06fF
C45446 OR2X1_LOC_49/A OR2X1_LOC_54/a_8_216# 0.06fF
C47140 OR2X1_LOC_49/A OR2X1_LOC_87/B 0.23fF
C47476 OR2X1_LOC_49/A OR2X1_LOC_671/Y 0.81fF
C47596 OR2X1_LOC_49/A OR2X1_LOC_42/a_8_216# 0.01fF
C47690 OR2X1_LOC_49/A OR2X1_LOC_532/B 1.08fF
C48855 OR2X1_LOC_49/A AND2X1_LOC_412/a_8_24# 0.01fF
C49634 OR2X1_LOC_49/A VDD 0.69fF
C50485 OR2X1_LOC_49/A OR2X1_LOC_382/Y 0.01fF
C50935 OR2X1_LOC_49/A OR2X1_LOC_427/A 0.10fF
C51804 OR2X1_LOC_49/A OR2X1_LOC_6/A 0.62fF
C52540 OR2X1_LOC_49/A OR2X1_LOC_382/A 0.11fF
C52623 OR2X1_LOC_49/A OR2X1_LOC_160/A 0.11fF
C52970 OR2X1_LOC_49/A OR2X1_LOC_158/A 2.63fF
C53054 OR2X1_LOC_49/A OR2X1_LOC_847/A 0.03fF
C53136 OR2X1_LOC_49/A AND2X1_LOC_46/a_8_24# 0.01fF
C53513 OR2X1_LOC_49/A OR2X1_LOC_748/A 0.03fF
C53978 OR2X1_LOC_49/A AND2X1_LOC_119/a_8_24# -0.01fF
C54814 OR2X1_LOC_49/A OR2X1_LOC_293/a_8_216# 0.01fF
C58065 OR2X1_LOC_49/A VSS 0.78fF
C419 AND2X1_LOC_12/Y OR2X1_LOC_847/B 0.04fF
C8310 OR2X1_LOC_847/B OR2X1_LOC_68/B 0.05fF
C20860 OR2X1_LOC_847/A OR2X1_LOC_847/B 0.17fF
C27640 AND2X1_LOC_817/a_8_24# OR2X1_LOC_847/B 0.01fF
C35637 OR2X1_LOC_847/a_8_216# OR2X1_LOC_847/B 0.47fF
C56761 OR2X1_LOC_847/B VSS 0.16fF
C1409 OR2X1_LOC_62/B AND2X1_LOC_4/a_8_24# 0.01fF
C1519 OR2X1_LOC_62/B OR2X1_LOC_68/B 0.08fF
C1821 OR2X1_LOC_62/B OR2X1_LOC_74/A 0.02fF
C2245 OR2X1_LOC_62/B OR2X1_LOC_87/A 0.03fF
C2314 OR2X1_LOC_62/B AND2X1_LOC_15/a_36_24# 0.01fF
C3511 AND2X1_LOC_63/a_8_24# OR2X1_LOC_62/B 0.01fF
C4337 OR2X1_LOC_62/B OR2X1_LOC_278/a_8_216# 0.03fF
C4731 OR2X1_LOC_154/A OR2X1_LOC_62/B 0.08fF
C5867 OR2X1_LOC_62/B OR2X1_LOC_633/A 0.03fF
C6224 AND2X1_LOC_64/Y OR2X1_LOC_62/B 0.10fF
C6289 AND2X1_LOC_86/a_8_24# OR2X1_LOC_62/B 0.01fF
C6878 AND2X1_LOC_55/a_8_24# OR2X1_LOC_62/B 0.01fF
C7366 OR2X1_LOC_611/a_8_216# OR2X1_LOC_62/B 0.01fF
C8597 AND2X1_LOC_529/a_8_24# OR2X1_LOC_62/B 0.01fF
C8713 OR2X1_LOC_62/B OR2X1_LOC_532/B 0.34fF
C9917 OR2X1_LOC_185/Y OR2X1_LOC_62/B 0.05fF
C9937 OR2X1_LOC_62/B OR2X1_LOC_278/a_36_216# 0.03fF
C10653 VDD OR2X1_LOC_62/B 1.24fF
C12872 OR2X1_LOC_62/B OR2X1_LOC_6/A 0.02fF
C13715 OR2X1_LOC_160/A OR2X1_LOC_62/B 0.16fF
C13743 AND2X1_LOC_86/B OR2X1_LOC_62/B 0.02fF
C14006 OR2X1_LOC_62/B OR2X1_LOC_266/A 0.02fF
C14969 OR2X1_LOC_185/A OR2X1_LOC_62/B 0.03fF
C17331 AND2X1_LOC_91/B OR2X1_LOC_62/B 0.03fF
C17937 AND2X1_LOC_56/B OR2X1_LOC_62/B 0.01fF
C17946 AND2X1_LOC_8/Y OR2X1_LOC_62/B 0.21fF
C18429 OR2X1_LOC_291/Y OR2X1_LOC_62/B 0.01fF
C19307 OR2X1_LOC_62/B AND2X1_LOC_47/Y 0.27fF
C20057 OR2X1_LOC_62/B AND2X1_LOC_414/a_8_24# 0.01fF
C20074 AND2X1_LOC_95/Y OR2X1_LOC_62/B 0.21fF
C20354 AND2X1_LOC_22/Y OR2X1_LOC_62/B 0.05fF
C20557 OR2X1_LOC_296/a_8_216# OR2X1_LOC_62/B 0.01fF
C21337 OR2X1_LOC_235/B OR2X1_LOC_62/B 0.45fF
C23158 OR2X1_LOC_62/B OR2X1_LOC_62/a_8_216# 0.10fF
C23383 OR2X1_LOC_62/B AND2X1_LOC_44/Y 0.19fF
C23423 OR2X1_LOC_600/A OR2X1_LOC_62/B 0.03fF
C23497 OR2X1_LOC_62/B OR2X1_LOC_619/Y 0.03fF
C24271 OR2X1_LOC_62/B AND2X1_LOC_18/Y 0.09fF
C26904 OR2X1_LOC_62/B OR2X1_LOC_54/Y 0.13fF
C27274 OR2X1_LOC_62/B OR2X1_LOC_161/A 0.29fF
C27321 OR2X1_LOC_62/B AND2X1_LOC_51/Y 0.03fF
C28068 AND2X1_LOC_41/A OR2X1_LOC_62/B 0.01fF
C29114 OR2X1_LOC_62/B OR2X1_LOC_71/A 2.24fF
C29899 OR2X1_LOC_62/B OR2X1_LOC_47/Y 0.02fF
C30182 AND2X1_LOC_143/a_8_24# OR2X1_LOC_62/B 0.01fF
C30343 OR2X1_LOC_62/B AND2X1_LOC_72/B 0.05fF
C30434 OR2X1_LOC_62/B AND2X1_LOC_36/Y 0.03fF
C30949 OR2X1_LOC_62/B OR2X1_LOC_16/A 0.05fF
C31435 AND2X1_LOC_126/a_8_24# OR2X1_LOC_62/B 0.01fF
C33061 OR2X1_LOC_40/Y OR2X1_LOC_62/B 0.02fF
C33797 OR2X1_LOC_62/B OR2X1_LOC_777/B 3.41fF
C34081 OR2X1_LOC_62/B OR2X1_LOC_62/a_36_216# 0.03fF
C34281 OR2X1_LOC_62/B OR2X1_LOC_161/B 0.03fF
C35316 AND2X1_LOC_133/a_8_24# OR2X1_LOC_62/B 0.01fF
C35666 OR2X1_LOC_502/A OR2X1_LOC_62/B 0.04fF
C35841 OR2X1_LOC_62/B OR2X1_LOC_398/a_8_216# 0.01fF
C36146 OR2X1_LOC_62/B AND2X1_LOC_3/Y 0.03fF
C36976 OR2X1_LOC_296/Y OR2X1_LOC_62/B 0.37fF
C38560 OR2X1_LOC_160/B OR2X1_LOC_62/B 0.12fF
C39293 OR2X1_LOC_62/B AND2X1_LOC_246/a_8_24# 0.09fF
C39419 OR2X1_LOC_151/A OR2X1_LOC_62/B 0.11fF
C41742 OR2X1_LOC_62/B AND2X1_LOC_15/a_8_24# 0.03fF
C42156 OR2X1_LOC_19/B OR2X1_LOC_62/B 0.08fF
C43466 OR2X1_LOC_611/Y OR2X1_LOC_62/B 0.01fF
C43857 OR2X1_LOC_36/Y OR2X1_LOC_62/B 0.02fF
C44180 OR2X1_LOC_62/B OR2X1_LOC_66/A 0.09fF
C45537 AND2X1_LOC_40/Y OR2X1_LOC_62/B 0.03fF
C46501 AND2X1_LOC_159/a_8_24# OR2X1_LOC_62/B 0.11fF
C47072 OR2X1_LOC_62/B OR2X1_LOC_398/Y 0.03fF
C48586 OR2X1_LOC_62/B OR2X1_LOC_78/A 0.05fF
C49046 OR2X1_LOC_291/a_8_216# OR2X1_LOC_62/B 0.01fF
C49925 AND2X1_LOC_12/Y OR2X1_LOC_62/B 0.03fF
C50369 AND2X1_LOC_59/Y OR2X1_LOC_62/B 0.02fF
C50809 OR2X1_LOC_62/B OR2X1_LOC_585/A 0.05fF
C51614 OR2X1_LOC_62/B OR2X1_LOC_753/A 0.03fF
C52365 OR2X1_LOC_8/Y OR2X1_LOC_62/B 0.70fF
C53286 OR2X1_LOC_62/B OR2X1_LOC_39/A 0.03fF
C53729 OR2X1_LOC_377/A OR2X1_LOC_62/B 0.06fF
C53751 OR2X1_LOC_62/B OR2X1_LOC_85/A 0.15fF
C54049 OR2X1_LOC_62/B OR2X1_LOC_78/B 0.03fF
C54105 OR2X1_LOC_62/B OR2X1_LOC_375/A 0.10fF
C55287 OR2X1_LOC_62/B AND2X1_LOC_65/A 0.01fF
C55895 AND2X1_LOC_10/a_8_24# OR2X1_LOC_62/B 0.09fF
C57188 OR2X1_LOC_62/B VSS 0.42fF
C1263 OR2X1_LOC_54/Y OR2X1_LOC_382/a_8_216# -0.03fF
C1475 AND2X1_LOC_8/a_8_24# OR2X1_LOC_54/Y 0.03fF
C2617 OR2X1_LOC_91/A OR2X1_LOC_54/Y 3.49fF
C2668 AND2X1_LOC_62/a_36_24# OR2X1_LOC_54/Y 0.01fF
C3130 OR2X1_LOC_233/a_8_216# OR2X1_LOC_54/Y 0.01fF
C3241 OR2X1_LOC_54/Y OR2X1_LOC_68/B 0.10fF
C3548 OR2X1_LOC_74/A OR2X1_LOC_54/Y 0.02fF
C4188 OR2X1_LOC_54/Y OR2X1_LOC_381/a_8_216# 0.03fF
C4327 AND2X1_LOC_611/a_8_24# OR2X1_LOC_54/Y 0.01fF
C4366 AND2X1_LOC_671/a_36_24# OR2X1_LOC_54/Y 0.01fF
C5138 OR2X1_LOC_699/a_8_216# OR2X1_LOC_54/Y 0.03fF
C5593 AND2X1_LOC_37/a_8_24# OR2X1_LOC_54/Y 0.01fF
C7331 OR2X1_LOC_485/A OR2X1_LOC_54/Y 0.05fF
C7408 OR2X1_LOC_10/a_8_216# OR2X1_LOC_54/Y 0.01fF
C8122 OR2X1_LOC_54/Y AND2X1_LOC_819/a_8_24# 0.01fF
C8278 OR2X1_LOC_54/a_8_216# OR2X1_LOC_54/Y 0.01fF
C9924 AND2X1_LOC_612/B OR2X1_LOC_54/Y 0.01fF
C10195 OR2X1_LOC_671/Y OR2X1_LOC_54/Y 0.01fF
C10386 OR2X1_LOC_532/B OR2X1_LOC_54/Y 0.07fF
C12335 VDD OR2X1_LOC_54/Y 0.48fF
C13255 OR2X1_LOC_382/Y OR2X1_LOC_54/Y 0.01fF
C13661 OR2X1_LOC_54/Y AND2X1_LOC_820/B 0.01fF
C13696 OR2X1_LOC_427/A OR2X1_LOC_54/Y 0.41fF
C14558 OR2X1_LOC_54/Y OR2X1_LOC_6/A 0.48fF
C15245 OR2X1_LOC_54/Y OR2X1_LOC_382/A 0.10fF
C15659 OR2X1_LOC_158/A OR2X1_LOC_54/Y 0.36fF
C16232 OR2X1_LOC_748/A OR2X1_LOC_54/Y 0.01fF
C16624 OR2X1_LOC_185/A OR2X1_LOC_54/Y 0.07fF
C17538 OR2X1_LOC_293/a_8_216# OR2X1_LOC_54/Y 0.01fF
C19587 OR2X1_LOC_54/Y OR2X1_LOC_56/A 0.29fF
C19669 AND2X1_LOC_56/B OR2X1_LOC_54/Y 0.18fF
C19683 AND2X1_LOC_8/Y OR2X1_LOC_54/Y 0.07fF
C20874 AND2X1_LOC_73/a_8_24# OR2X1_LOC_54/Y 0.06fF
C21015 AND2X1_LOC_47/Y OR2X1_LOC_54/Y 0.05fF
C21429 OR2X1_LOC_481/A OR2X1_LOC_54/Y 0.07fF
C21661 OR2X1_LOC_54/Y OR2X1_LOC_15/a_8_216# 0.04fF
C23044 OR2X1_LOC_235/B OR2X1_LOC_54/Y 0.08fF
C24725 OR2X1_LOC_92/Y OR2X1_LOC_54/Y 0.04fF
C24819 OR2X1_LOC_62/a_8_216# OR2X1_LOC_54/Y 0.02fF
C25073 OR2X1_LOC_600/A OR2X1_LOC_54/Y 1.06fF
C25154 OR2X1_LOC_619/Y OR2X1_LOC_54/Y 0.15fF
C25589 OR2X1_LOC_54/Y AND2X1_LOC_818/a_8_24# 0.10fF
C26090 AND2X1_LOC_672/a_8_24# OR2X1_LOC_54/Y 0.03fF
C27436 OR2X1_LOC_54/Y OR2X1_LOC_13/B 0.01fF
C27960 OR2X1_LOC_54/Y OR2X1_LOC_428/A 0.14fF
C28966 OR2X1_LOC_26/Y OR2X1_LOC_54/Y 0.08fF
C28982 OR2X1_LOC_89/A OR2X1_LOC_54/Y 0.02fF
C29807 OR2X1_LOC_824/Y OR2X1_LOC_54/Y 0.42fF
C29882 OR2X1_LOC_95/Y OR2X1_LOC_54/Y 0.08fF
C30647 AND2X1_LOC_102/a_8_24# OR2X1_LOC_54/Y 0.04fF
C30807 OR2X1_LOC_54/Y OR2X1_LOC_71/A 0.47fF
C31084 OR2X1_LOC_54/Y OR2X1_LOC_820/B 0.53fF
C31509 OR2X1_LOC_54/Y OR2X1_LOC_240/A 0.12fF
C31590 OR2X1_LOC_47/Y OR2X1_LOC_54/Y 0.08fF
C32071 OR2X1_LOC_54/Y AND2X1_LOC_36/Y 6.20fF
C32609 OR2X1_LOC_54/Y OR2X1_LOC_16/A 0.02fF
C33505 OR2X1_LOC_93/Y OR2X1_LOC_54/Y 0.02fF
C34749 OR2X1_LOC_159/a_8_216# OR2X1_LOC_54/Y 0.40fF
C34753 OR2X1_LOC_40/Y OR2X1_LOC_54/Y 0.08fF
C34912 OR2X1_LOC_7/A OR2X1_LOC_54/Y 0.65fF
C36123 OR2X1_LOC_43/A OR2X1_LOC_54/Y 0.28fF
C36538 OR2X1_LOC_54/Y AND2X1_LOC_818/a_36_24# 0.01fF
C36970 OR2X1_LOC_3/Y OR2X1_LOC_54/Y 0.02fF
C37038 OR2X1_LOC_673/A OR2X1_LOC_54/Y 0.05fF
C37330 OR2X1_LOC_502/A OR2X1_LOC_54/Y 0.14fF
C37664 AND2X1_LOC_530/a_8_24# OR2X1_LOC_54/Y 0.04fF
C39596 OR2X1_LOC_54/Y OR2X1_LOC_77/a_8_216# 0.14fF
C41691 AND2X1_LOC_102/a_36_24# OR2X1_LOC_54/Y 0.01fF
C41836 OR2X1_LOC_54/Y OR2X1_LOC_150/a_8_216# 0.01fF
C42070 AND2X1_LOC_62/a_8_24# OR2X1_LOC_54/Y 0.04fF
C42352 OR2X1_LOC_54/Y OR2X1_LOC_415/Y 0.16fF
C42655 OR2X1_LOC_234/a_8_216# OR2X1_LOC_54/Y 0.01fF
C43826 OR2X1_LOC_54/Y OR2X1_LOC_38/a_8_216# 0.04fF
C43898 OR2X1_LOC_19/B OR2X1_LOC_54/Y 0.05fF
C45576 OR2X1_LOC_36/Y OR2X1_LOC_54/Y 0.03fF
C45898 OR2X1_LOC_604/A OR2X1_LOC_54/Y 0.20fF
C45913 OR2X1_LOC_54/Y OR2X1_LOC_66/A 0.03fF
C47612 OR2X1_LOC_143/a_8_216# OR2X1_LOC_54/Y 0.01fF
C47740 OR2X1_LOC_90/a_8_216# OR2X1_LOC_54/Y 0.07fF
C48952 AND2X1_LOC_530/a_36_24# OR2X1_LOC_54/Y 0.01fF
C49374 OR2X1_LOC_54/Y OR2X1_LOC_12/Y 0.02fF
C49579 AND2X1_LOC_671/a_8_24# OR2X1_LOC_54/Y 0.03fF
C49882 OR2X1_LOC_54/Y OR2X1_LOC_234/Y -0.01fF
C52466 OR2X1_LOC_585/A OR2X1_LOC_54/Y 0.01fF
C53057 OR2X1_LOC_54/Y OR2X1_LOC_437/A 0.01fF
C54029 OR2X1_LOC_8/Y OR2X1_LOC_54/Y 1.99fF
C54950 OR2X1_LOC_54/Y OR2X1_LOC_39/A 0.01fF
C55393 OR2X1_LOC_377/A OR2X1_LOC_54/Y 0.29fF
C55405 OR2X1_LOC_85/A OR2X1_LOC_54/Y 0.54fF
C55765 OR2X1_LOC_51/Y OR2X1_LOC_54/Y 0.06fF
C55829 AND2X1_LOC_94/a_8_24# OR2X1_LOC_54/Y 0.02fF
C55848 OR2X1_LOC_375/A OR2X1_LOC_54/Y 0.05fF
C56820 OR2X1_LOC_54/Y VSS 1.08fF
C25 OR2X1_LOC_43/A OR2X1_LOC_73/a_8_216# 0.03fF
C359 AND2X1_LOC_377/Y OR2X1_LOC_43/A 0.10fF
C701 OR2X1_LOC_43/A OR2X1_LOC_12/Y 0.41fF
C846 OR2X1_LOC_694/a_8_216# OR2X1_LOC_43/A 0.06fF
C923 OR2X1_LOC_272/Y OR2X1_LOC_43/A 0.03fF
C3437 OR2X1_LOC_43/A OR2X1_LOC_18/Y 0.25fF
C3896 OR2X1_LOC_43/A OR2X1_LOC_585/A 0.10fF
C4271 OR2X1_LOC_43/A OR2X1_LOC_827/a_36_216# 0.01fF
C4420 OR2X1_LOC_43/A OR2X1_LOC_437/A 0.22fF
C4684 OR2X1_LOC_43/A OR2X1_LOC_753/A 0.10fF
C4732 OR2X1_LOC_43/A OR2X1_LOC_684/Y 0.01fF
C5206 OR2X1_LOC_43/A OR2X1_LOC_88/Y 0.03fF
C5386 OR2X1_LOC_8/Y OR2X1_LOC_43/A 0.04fF
C5525 OR2X1_LOC_43/A OR2X1_LOC_52/B 0.21fF
C5528 OR2X1_LOC_43/A OR2X1_LOC_672/Y 0.01fF
C5780 OR2X1_LOC_43/A OR2X1_LOC_9/a_8_216# 0.02fF
C5858 AND2X1_LOC_514/a_8_24# OR2X1_LOC_43/A 0.03fF
C5872 AND2X1_LOC_378/a_8_24# OR2X1_LOC_43/A 0.04fF
C6007 OR2X1_LOC_43/A OR2X1_LOC_22/Y 0.21fF
C6323 OR2X1_LOC_43/A OR2X1_LOC_39/A 0.37fF
C6800 OR2X1_LOC_43/A OR2X1_LOC_85/A 1.61fF
C7048 OR2X1_LOC_136/Y OR2X1_LOC_43/A 0.07fF
C7140 OR2X1_LOC_43/A OR2X1_LOC_51/Y 0.19fF
C8276 OR2X1_LOC_43/A OR2X1_LOC_86/A 0.03fF
C8707 OR2X1_LOC_43/A OR2X1_LOC_599/Y 0.31fF
C8852 OR2X1_LOC_43/A OR2X1_LOC_382/a_8_216# 0.01fF
C10185 OR2X1_LOC_43/A OR2X1_LOC_91/A 10.31fF
C11117 OR2X1_LOC_43/A OR2X1_LOC_74/A 0.17fF
C11803 OR2X1_LOC_43/A OR2X1_LOC_381/a_8_216# 0.01fF
C12425 OR2X1_LOC_43/A OR2X1_LOC_275/a_8_216# 0.06fF
C12810 OR2X1_LOC_699/a_8_216# OR2X1_LOC_43/A 0.03fF
C13098 OR2X1_LOC_43/Y OR2X1_LOC_43/A 0.01fF
C14378 OR2X1_LOC_43/A OR2X1_LOC_382/a_36_216# -0.01fF
C14910 OR2X1_LOC_43/A OR2X1_LOC_94/a_8_216# 0.43fF
C14954 OR2X1_LOC_485/A OR2X1_LOC_43/A 0.53fF
C15806 OR2X1_LOC_43/A OR2X1_LOC_54/a_8_216# 0.04fF
C16649 OR2X1_LOC_43/A OR2X1_LOC_43/a_8_216# 0.01fF
C16976 AND2X1_LOC_378/a_36_24# OR2X1_LOC_43/A 0.01fF
C17707 OR2X1_LOC_671/Y OR2X1_LOC_43/A 0.43fF
C17869 OR2X1_LOC_43/A OR2X1_LOC_42/a_8_216# 0.03fF
C18329 OR2X1_LOC_699/a_36_216# OR2X1_LOC_43/A 0.01fF
C18653 OR2X1_LOC_43/A AND2X1_LOC_691/a_8_24# 0.01fF
C19306 OR2X1_LOC_43/A OR2X1_LOC_761/a_8_216# 0.02fF
C19932 VDD OR2X1_LOC_43/A 1.08fF
C19993 OR2X1_LOC_689/A OR2X1_LOC_43/A 0.39fF
C21277 OR2X1_LOC_43/A OR2X1_LOC_427/A 1.26fF
C21280 OR2X1_LOC_43/A AND2X1_LOC_801/a_8_24# -0.00fF
C21411 OR2X1_LOC_43/A AND2X1_LOC_687/B 1.51fF
C22191 OR2X1_LOC_43/A OR2X1_LOC_6/A 0.19fF
C22635 OR2X1_LOC_43/A OR2X1_LOC_44/Y 0.13fF
C22896 OR2X1_LOC_45/B OR2X1_LOC_43/A 0.13fF
C22924 OR2X1_LOC_43/A OR2X1_LOC_382/A 0.02fF
C23318 OR2X1_LOC_158/A OR2X1_LOC_43/A 0.53fF
C23886 OR2X1_LOC_748/A OR2X1_LOC_43/A 0.01fF
C25844 OR2X1_LOC_744/A OR2X1_LOC_43/A 0.10fF
C26029 OR2X1_LOC_43/A OR2X1_LOC_31/Y 0.38fF
C26756 OR2X1_LOC_43/A AND2X1_LOC_809/A 0.01fF
C27142 OR2X1_LOC_43/A OR2X1_LOC_56/A 2.31fF
C27691 OR2X1_LOC_417/Y OR2X1_LOC_43/A 0.03fF
C28754 OR2X1_LOC_672/a_8_216# OR2X1_LOC_43/A 0.03fF
C28940 OR2X1_LOC_43/A OR2X1_LOC_481/A 0.07fF
C28985 OR2X1_LOC_43/A OR2X1_LOC_71/Y 0.03fF
C29208 OR2X1_LOC_426/B OR2X1_LOC_43/A 0.28fF
C31426 OR2X1_LOC_43/A OR2X1_LOC_96/B 0.03fF
C32185 OR2X1_LOC_43/A OR2X1_LOC_92/Y 0.13fF
C32213 OR2X1_LOC_43/A OR2X1_LOC_65/B 0.03fF
C32528 OR2X1_LOC_692/Y OR2X1_LOC_43/A 0.01fF
C32582 OR2X1_LOC_600/A OR2X1_LOC_43/A 0.18fF
C32605 OR2X1_LOC_43/A AND2X1_LOC_296/a_8_24# 0.01fF
C32661 OR2X1_LOC_43/A OR2X1_LOC_619/Y 0.10fF
C33108 OR2X1_LOC_690/a_8_216# OR2X1_LOC_43/A -0.01fF
C33111 OR2X1_LOC_43/A AND2X1_LOC_818/a_8_24# 0.01fF
C33267 OR2X1_LOC_43/A OR2X1_LOC_534/a_8_216# 0.02fF
C33823 OR2X1_LOC_133/a_8_216# OR2X1_LOC_43/A 0.04fF
C33848 OR2X1_LOC_329/Y OR2X1_LOC_43/A 0.01fF
C35002 OR2X1_LOC_43/A OR2X1_LOC_13/B 7.97fF
C35466 OR2X1_LOC_43/A OR2X1_LOC_428/A 0.43fF
C36434 OR2X1_LOC_689/a_8_216# OR2X1_LOC_43/A 0.01fF
C36489 OR2X1_LOC_43/A OR2X1_LOC_26/Y 0.13fF
C36505 OR2X1_LOC_43/A OR2X1_LOC_89/A 0.53fF
C36585 OR2X1_LOC_43/A OR2X1_LOC_419/a_8_216# 0.01fF
C36851 OR2X1_LOC_306/a_8_216# OR2X1_LOC_43/A 0.03fF
C37426 OR2X1_LOC_43/A OR2X1_LOC_95/Y 0.15fF
C38505 OR2X1_LOC_43/A OR2X1_LOC_59/Y 0.07fF
C38617 OR2X1_LOC_43/A OR2X1_LOC_820/B 0.02fF
C38650 OR2X1_LOC_70/Y OR2X1_LOC_43/A 0.13fF
C38763 OR2X1_LOC_43/A OR2X1_LOC_534/a_36_216# 0.03fF
C39156 OR2X1_LOC_43/A OR2X1_LOC_47/Y 0.18fF
C39886 OR2X1_LOC_246/Y OR2X1_LOC_43/A 0.07fF
C40113 OR2X1_LOC_43/A OR2X1_LOC_16/A 0.15fF
C41202 OR2X1_LOC_43/A AND2X1_LOC_729/B 0.80fF
C42045 OR2X1_LOC_599/A OR2X1_LOC_43/A 0.03fF
C42351 OR2X1_LOC_159/a_8_216# OR2X1_LOC_43/A 0.04fF
C42354 OR2X1_LOC_40/Y OR2X1_LOC_43/A 0.52fF
C42509 OR2X1_LOC_43/A OR2X1_LOC_7/A 0.22fF
C42908 OR2X1_LOC_43/A OR2X1_LOC_236/a_8_216# 0.03fF
C43650 OR2X1_LOC_589/A OR2X1_LOC_43/A 1.11fF
C43706 OR2X1_LOC_43/A OR2X1_LOC_297/A 0.01fF
C44366 OR2X1_LOC_43/A OR2X1_LOC_534/Y 0.44fF
C44681 OR2X1_LOC_3/Y OR2X1_LOC_43/A 0.48fF
C44996 OR2X1_LOC_329/B OR2X1_LOC_43/A 0.03fF
C45966 OR2X1_LOC_43/A OR2X1_LOC_690/A 0.77fF
C45990 OR2X1_LOC_272/a_8_216# OR2X1_LOC_43/A 0.06fF
C46015 OR2X1_LOC_43/A OR2X1_LOC_64/Y 0.19fF
C46515 OR2X1_LOC_43/A OR2X1_LOC_55/a_8_216# 0.03fF
C47401 OR2X1_LOC_43/A OR2X1_LOC_77/a_8_216# 0.04fF
C47779 AND2X1_LOC_512/a_8_24# OR2X1_LOC_43/A 0.01fF
C48600 OR2X1_LOC_43/A OR2X1_LOC_236/a_36_216# 0.01fF
C49387 OR2X1_LOC_43/A OR2X1_LOC_517/A 0.10fF
C49468 OR2X1_LOC_43/A OR2X1_LOC_827/a_8_216# 0.05fF
C51510 OR2X1_LOC_43/A OR2X1_LOC_278/Y 0.03fF
C51601 OR2X1_LOC_43/A OR2X1_LOC_19/B 0.07fF
C52017 OR2X1_LOC_43/A OR2X1_LOC_275/A 0.06fF
C52924 OR2X1_LOC_43/A OR2X1_LOC_689/Y 0.01fF
C53239 OR2X1_LOC_43/A OR2X1_LOC_36/Y 0.29fF
C53354 OR2X1_LOC_43/A OR2X1_LOC_419/Y 0.01fF
C53557 OR2X1_LOC_604/A OR2X1_LOC_43/A 0.10fF
C53680 OR2X1_LOC_306/Y OR2X1_LOC_43/A 0.09fF
C55262 OR2X1_LOC_43/A OR2X1_LOC_90/a_8_216# 0.07fF
C57423 OR2X1_LOC_43/A VSS 1.00fF
C38 OR2X1_LOC_19/B AND2X1_LOC_233/a_8_24# 0.17fF
C872 OR2X1_LOC_19/B OR2X1_LOC_517/A 0.05fF
C3072 OR2X1_LOC_19/B OR2X1_LOC_278/Y 0.02fF
C3183 OR2X1_LOC_19/B OR2X1_LOC_838/B 0.01fF
C4729 OR2X1_LOC_36/Y OR2X1_LOC_19/B 0.08fF
C4934 OR2X1_LOC_19/B OR2X1_LOC_19/a_8_216# 0.09fF
C5035 OR2X1_LOC_19/B OR2X1_LOC_66/A 0.86fF
C5411 OR2X1_LOC_691/a_8_216# OR2X1_LOC_19/B 0.01fF
C5472 AND2X1_LOC_94/Y OR2X1_LOC_19/B 0.03fF
C5863 OR2X1_LOC_490/a_8_216# OR2X1_LOC_19/B 0.01fF
C8699 OR2X1_LOC_19/B AND2X1_LOC_671/a_8_24# 0.09fF
C8734 OR2X1_LOC_19/B OR2X1_LOC_644/A -0.01fF
C9093 OR2X1_LOC_19/B OR2X1_LOC_278/A 0.07fF
C9407 OR2X1_LOC_19/B OR2X1_LOC_78/A 1.94fF
C10332 AND2X1_LOC_387/B OR2X1_LOC_19/B 0.07fF
C10716 AND2X1_LOC_12/Y OR2X1_LOC_19/B 0.10fF
C11116 OR2X1_LOC_18/Y OR2X1_LOC_19/B 0.89fF
C11124 AND2X1_LOC_59/Y OR2X1_LOC_19/B 3.84fF
C11589 OR2X1_LOC_19/B OR2X1_LOC_585/A 0.09fF
C12444 OR2X1_LOC_19/B OR2X1_LOC_753/A 0.20fF
C13009 OR2X1_LOC_19/B OR2X1_LOC_88/Y 0.01fF
C13214 OR2X1_LOC_8/Y OR2X1_LOC_19/B 0.06fF
C13772 OR2X1_LOC_22/Y OR2X1_LOC_19/B 0.03fF
C14137 OR2X1_LOC_19/B OR2X1_LOC_39/A 0.98fF
C14252 OR2X1_LOC_19/B AND2X1_LOC_761/a_8_24# 0.01fF
C14535 OR2X1_LOC_377/A OR2X1_LOC_19/B 0.32fF
C14553 OR2X1_LOC_19/B OR2X1_LOC_85/A 0.04fF
C14903 OR2X1_LOC_19/B OR2X1_LOC_78/B 0.01fF
C14971 OR2X1_LOC_19/B OR2X1_LOC_375/A 0.07fF
C15240 OR2X1_LOC_19/B OR2X1_LOC_549/A 0.02fF
C15900 OR2X1_LOC_19/B OR2X1_LOC_86/A 0.01fF
C16038 OR2X1_LOC_19/B OR2X1_LOC_20/A 0.01fF
C16288 AND2X1_LOC_23/a_8_24# OR2X1_LOC_19/B 0.04fF
C17059 OR2X1_LOC_19/B OR2X1_LOC_414/a_8_216# 0.06fF
C17839 OR2X1_LOC_91/A OR2X1_LOC_19/B 0.03fF
C18365 OR2X1_LOC_32/B OR2X1_LOC_19/B 0.01fF
C18411 OR2X1_LOC_19/B AND2X1_LOC_4/a_8_24# 0.14fF
C18516 OR2X1_LOC_19/B OR2X1_LOC_68/B 1.64fF
C18840 OR2X1_LOC_490/Y OR2X1_LOC_19/B 0.01fF
C18841 OR2X1_LOC_19/B OR2X1_LOC_74/A 0.07fF
C19283 OR2X1_LOC_263/a_8_216# OR2X1_LOC_19/B 0.01fF
C19629 OR2X1_LOC_19/B OR2X1_LOC_23/a_8_216# -0.04fF
C20062 OR2X1_LOC_19/B OR2X1_LOC_71/a_8_216# 0.02fF
C20783 OR2X1_LOC_691/Y OR2X1_LOC_19/B 0.04fF
C21904 OR2X1_LOC_19/B AND2X1_LOC_6/a_8_24# 0.09fF
C22598 OR2X1_LOC_461/a_8_216# OR2X1_LOC_19/B 0.14fF
C22621 OR2X1_LOC_634/A OR2X1_LOC_19/B 0.03fF
C22666 OR2X1_LOC_19/B OR2X1_LOC_414/a_36_216# 0.01fF
C22722 OR2X1_LOC_485/A OR2X1_LOC_19/B 0.06fF
C22966 OR2X1_LOC_19/B OR2X1_LOC_633/A 0.05fF
C23075 OR2X1_LOC_19/B OR2X1_LOC_256/a_8_216# 0.02fF
C23325 AND2X1_LOC_64/Y OR2X1_LOC_19/B 0.34fF
C23358 AND2X1_LOC_599/a_8_24# OR2X1_LOC_19/B 0.02fF
C23925 AND2X1_LOC_55/a_8_24# OR2X1_LOC_19/B 0.01fF
C24766 OR2X1_LOC_19/B OR2X1_LOC_82/a_8_216# 0.03fF
C25516 AND2X1_LOC_529/a_8_24# OR2X1_LOC_19/B 0.01fF
C25652 OR2X1_LOC_19/B OR2X1_LOC_532/B 0.14fF
C26854 OR2X1_LOC_19/B AND2X1_LOC_412/a_8_24# 0.07fF
C27592 VDD OR2X1_LOC_19/B 1.34fF
C27758 OR2X1_LOC_19/B OR2X1_LOC_256/A 0.08fF
C28516 OR2X1_LOC_19/B OR2X1_LOC_256/a_36_216# 0.03fF
C28930 OR2X1_LOC_19/B OR2X1_LOC_63/a_8_216# 0.02fF
C29803 OR2X1_LOC_19/B OR2X1_LOC_6/A 0.17fF
C30227 OR2X1_LOC_19/B OR2X1_LOC_82/a_36_216# 0.01fF
C30361 OR2X1_LOC_19/B OR2X1_LOC_750/Y 0.01fF
C30478 OR2X1_LOC_45/B OR2X1_LOC_19/B 0.10fF
C30619 OR2X1_LOC_160/A OR2X1_LOC_19/B 0.10fF
C31860 OR2X1_LOC_185/A OR2X1_LOC_19/B 0.03fF
C33537 OR2X1_LOC_744/A OR2X1_LOC_19/B 0.05fF
C34244 AND2X1_LOC_91/B OR2X1_LOC_19/B 0.09fF
C34789 OR2X1_LOC_19/B OR2X1_LOC_56/A 0.24fF
C34889 AND2X1_LOC_56/B OR2X1_LOC_19/B 0.24fF
C34903 AND2X1_LOC_8/Y OR2X1_LOC_19/B 0.63fF
C35299 OR2X1_LOC_291/Y OR2X1_LOC_19/B 0.07fF
C35712 OR2X1_LOC_19/B OR2X1_LOC_83/A 0.07fF
C36046 AND2X1_LOC_73/a_8_24# OR2X1_LOC_19/B 0.01fF
C36189 OR2X1_LOC_19/B AND2X1_LOC_47/Y 0.03fF
C36589 OR2X1_LOC_19/B OR2X1_LOC_71/Y 0.01fF
C36841 OR2X1_LOC_426/B OR2X1_LOC_19/B 0.84fF
C36892 OR2X1_LOC_19/B AND2X1_LOC_414/a_8_24# 0.01fF
C36907 AND2X1_LOC_95/Y OR2X1_LOC_19/B 0.05fF
C36995 OR2X1_LOC_19/B OR2X1_LOC_246/A 0.07fF
C37210 AND2X1_LOC_22/Y OR2X1_LOC_19/B 0.19fF
C38147 OR2X1_LOC_235/B OR2X1_LOC_19/B 0.10fF
C38509 OR2X1_LOC_709/A OR2X1_LOC_19/B 0.04fF
C38562 AND2X1_LOC_70/Y OR2X1_LOC_19/B 0.04fF
C39801 OR2X1_LOC_19/B OR2X1_LOC_414/Y 0.05fF
C39900 OR2X1_LOC_19/B OR2X1_LOC_92/Y 0.13fF
C39913 OR2X1_LOC_19/B OR2X1_LOC_65/B 0.03fF
C40167 OR2X1_LOC_19/B AND2X1_LOC_44/Y 0.10fF
C40227 OR2X1_LOC_600/A OR2X1_LOC_19/B 0.08fF
C40320 OR2X1_LOC_19/B OR2X1_LOC_619/Y 0.07fF
C40388 OR2X1_LOC_19/B AND2X1_LOC_4/a_36_24# 0.01fF
C41229 OR2X1_LOC_19/B AND2X1_LOC_234/a_8_24# 0.04fF
C41281 OR2X1_LOC_813/A OR2X1_LOC_19/B 0.01fF
C41552 OR2X1_LOC_19/B AND2X1_LOC_606/a_8_24# 0.02fF
C42092 OR2X1_LOC_19/B OR2X1_LOC_130/A 0.04fF
C42725 OR2X1_LOC_19/B OR2X1_LOC_13/B 0.09fF
C44281 OR2X1_LOC_19/B OR2X1_LOC_26/Y 0.14fF
C44310 OR2X1_LOC_19/B AND2X1_LOC_51/Y 0.03fF
C44349 OR2X1_LOC_19/B OR2X1_LOC_92/a_8_216# 0.01fF
C45071 AND2X1_LOC_41/A OR2X1_LOC_19/B 0.46fF
C45215 OR2X1_LOC_19/B OR2X1_LOC_95/Y 0.14fF
C45791 AND2X1_LOC_57/Y OR2X1_LOC_19/B 0.02fF
C46176 OR2X1_LOC_19/B OR2X1_LOC_71/A 0.08fF
C46384 OR2X1_LOC_19/B OR2X1_LOC_59/Y 0.16fF
C46511 OR2X1_LOC_70/Y OR2X1_LOC_19/B 0.01fF
C46608 OR2X1_LOC_19/B AND2X1_LOC_31/Y 0.03fF
C46930 OR2X1_LOC_19/B OR2X1_LOC_240/A 3.24fF
C47010 OR2X1_LOC_19/B OR2X1_LOC_47/Y 0.08fF
C47274 OR2X1_LOC_19/B OR2X1_LOC_607/A 0.01fF
C47594 OR2X1_LOC_19/B AND2X1_LOC_36/Y 0.19fF
C47913 OR2X1_LOC_19/B OR2X1_LOC_29/a_8_216# 0.01fF
C48106 OR2X1_LOC_19/B OR2X1_LOC_16/A 0.07fF
C48348 OR2X1_LOC_19/B AND2X1_LOC_827/a_8_24# 0.02fF
C48671 AND2X1_LOC_100/a_8_24# OR2X1_LOC_19/B 0.02fF
C49942 OR2X1_LOC_19/B OR2X1_LOC_269/B 0.08fF
C50242 OR2X1_LOC_40/Y OR2X1_LOC_19/B 0.07fF
C50392 OR2X1_LOC_19/B OR2X1_LOC_7/A 0.03fF
C50793 OR2X1_LOC_19/B OR2X1_LOC_86/a_8_216# 0.01fF
C50807 AND2X1_LOC_42/a_8_24# OR2X1_LOC_19/B 0.06fF
C51447 OR2X1_LOC_19/B OR2X1_LOC_161/B 0.17fF
C52467 OR2X1_LOC_19/B AND2X1_LOC_234/a_36_24# 0.01fF
C52475 OR2X1_LOC_3/Y OR2X1_LOC_19/B 0.70fF
C52835 OR2X1_LOC_502/A OR2X1_LOC_19/B 0.11fF
C52940 AND2X1_LOC_48/A OR2X1_LOC_19/B 0.37fF
C53306 OR2X1_LOC_19/B AND2X1_LOC_3/Y 0.32fF
C53785 OR2X1_LOC_64/Y OR2X1_LOC_19/B 0.09fF
C53959 OR2X1_LOC_19/B AND2X1_LOC_7/B 0.19fF
C54113 OR2X1_LOC_836/A OR2X1_LOC_19/B 0.03fF
C54131 AND2X1_LOC_101/B OR2X1_LOC_19/B 0.01fF
C55741 OR2X1_LOC_160/B OR2X1_LOC_19/B 0.04fF
C56132 OR2X1_LOC_691/B OR2X1_LOC_19/B 0.02fF
C57218 OR2X1_LOC_19/B VSS -4.13fF
C16 OR2X1_LOC_263/a_8_216# OR2X1_LOC_92/Y 0.01fF
C762 OR2X1_LOC_92/Y OR2X1_LOC_71/a_8_216# 0.01fF
C3434 OR2X1_LOC_485/A OR2X1_LOC_92/Y 0.24fF
C5789 OR2X1_LOC_310/Y OR2X1_LOC_92/Y 0.13fF
C5836 OR2X1_LOC_422/Y OR2X1_LOC_92/Y 0.01fF
C5856 OR2X1_LOC_92/Y OR2X1_LOC_433/Y 0.20fF
C5999 OR2X1_LOC_92/Y OR2X1_LOC_760/Y 0.03fF
C8075 OR2X1_LOC_682/a_8_216# OR2X1_LOC_92/Y 0.03fF
C8412 VDD OR2X1_LOC_92/Y 3.25fF
C8628 OR2X1_LOC_92/Y OR2X1_LOC_256/A 0.07fF
C9748 OR2X1_LOC_92/Y OR2X1_LOC_427/A 0.69fF
C10619 OR2X1_LOC_92/Y OR2X1_LOC_6/A 0.14fF
C11016 OR2X1_LOC_92/Y OR2X1_LOC_44/Y 0.13fF
C11279 OR2X1_LOC_45/B OR2X1_LOC_92/Y 0.96fF
C11750 OR2X1_LOC_158/A OR2X1_LOC_92/Y 0.24fF
C14350 OR2X1_LOC_744/A OR2X1_LOC_92/Y 0.17fF
C14540 OR2X1_LOC_92/Y OR2X1_LOC_31/Y 0.06fF
C15577 OR2X1_LOC_92/Y OR2X1_LOC_56/A 0.54fF
C16170 OR2X1_LOC_417/Y OR2X1_LOC_92/Y 0.07fF
C16569 OR2X1_LOC_92/Y AND2X1_LOC_276/Y 0.05fF
C16940 OR2X1_LOC_625/a_8_216# OR2X1_LOC_92/Y 0.02fF
C17421 OR2X1_LOC_481/A OR2X1_LOC_92/Y 0.03fF
C17470 OR2X1_LOC_92/Y OR2X1_LOC_71/Y 0.76fF
C17681 OR2X1_LOC_426/B OR2X1_LOC_92/Y 1.38fF
C17880 OR2X1_LOC_92/Y OR2X1_LOC_246/A 0.03fF
C17915 OR2X1_LOC_92/Y OR2X1_LOC_409/B 0.03fF
C17996 OR2X1_LOC_92/Y OR2X1_LOC_599/a_8_216# 0.03fF
C20801 OR2X1_LOC_92/Y OR2X1_LOC_65/B 0.02fF
C20836 OR2X1_LOC_271/Y OR2X1_LOC_92/Y 0.06fF
C21132 OR2X1_LOC_600/A OR2X1_LOC_92/Y 0.03fF
C21227 OR2X1_LOC_92/Y OR2X1_LOC_619/Y 0.14fF
C22222 OR2X1_LOC_813/A OR2X1_LOC_92/Y 0.01fF
C22524 OR2X1_LOC_625/a_36_216# OR2X1_LOC_92/Y 0.02fF
C23585 OR2X1_LOC_92/Y OR2X1_LOC_13/B 0.87fF
C24080 OR2X1_LOC_92/Y OR2X1_LOC_428/A 0.32fF
C24659 OR2X1_LOC_682/Y OR2X1_LOC_92/Y 0.14fF
C25065 OR2X1_LOC_92/Y OR2X1_LOC_26/Y 0.44fF
C25081 OR2X1_LOC_92/Y OR2X1_LOC_89/A 0.11fF
C25722 OR2X1_LOC_92/Y OR2X1_LOC_816/A 0.04fF
C25977 OR2X1_LOC_92/Y OR2X1_LOC_95/Y 0.35fF
C26911 OR2X1_LOC_92/Y OR2X1_LOC_71/A -0.00fF
C27067 OR2X1_LOC_92/Y OR2X1_LOC_59/Y 0.08fF
C27216 OR2X1_LOC_70/Y OR2X1_LOC_92/Y 0.47fF
C27696 OR2X1_LOC_92/Y OR2X1_LOC_47/Y 3.24fF
C28423 OR2X1_LOC_246/Y OR2X1_LOC_92/Y 0.13fF
C28675 OR2X1_LOC_92/Y OR2X1_LOC_16/A 0.10fF
C28915 OR2X1_LOC_92/Y AND2X1_LOC_687/Y 0.02fF
C29261 AND2X1_LOC_100/a_8_24# OR2X1_LOC_92/Y 0.03fF
C29331 OR2X1_LOC_92/Y OR2X1_LOC_268/a_8_216# 0.28fF
C29731 OR2X1_LOC_92/Y AND2X1_LOC_729/B 0.01fF
C30258 OR2X1_LOC_92/Y OR2X1_LOC_753/Y 0.01fF
C30515 OR2X1_LOC_599/A OR2X1_LOC_92/Y 0.07fF
C30830 OR2X1_LOC_40/Y OR2X1_LOC_92/Y 0.21fF
C30986 OR2X1_LOC_92/Y OR2X1_LOC_7/A 2.74fF
C31219 OR2X1_LOC_92/Y OR2X1_LOC_753/a_8_216# 0.01fF
C31388 OR2X1_LOC_92/Y OR2X1_LOC_86/a_8_216# 0.01fF
C32033 OR2X1_LOC_589/A OR2X1_LOC_92/Y 0.12fF
C32237 OR2X1_LOC_92/Y AND2X1_LOC_685/a_8_24# 0.35fF
C33074 OR2X1_LOC_3/Y OR2X1_LOC_92/Y 2.08fF
C33388 OR2X1_LOC_329/B OR2X1_LOC_92/Y 15.03fF
C34359 OR2X1_LOC_64/Y OR2X1_LOC_92/Y 0.28fF
C34761 AND2X1_LOC_101/B OR2X1_LOC_92/Y 0.51fF
C37604 OR2X1_LOC_517/A OR2X1_LOC_92/Y 0.10fF
C39695 OR2X1_LOC_92/Y OR2X1_LOC_421/Y 0.04fF
C39791 OR2X1_LOC_92/Y OR2X1_LOC_278/Y 0.08fF
C39908 OR2X1_LOC_92/Y AND2X1_LOC_800/a_8_24# 0.02fF
C40909 OR2X1_LOC_92/Y AND2X1_LOC_407/a_8_24# 0.04fF
C41544 OR2X1_LOC_36/Y OR2X1_LOC_92/Y 0.39fF
C41690 OR2X1_LOC_92/Y OR2X1_LOC_85/a_8_216# 0.33fF
C41859 OR2X1_LOC_604/A OR2X1_LOC_92/Y 0.06fF
C42716 OR2X1_LOC_490/a_8_216# OR2X1_LOC_92/Y 0.04fF
C43211 OR2X1_LOC_92/Y AND2X1_LOC_276/a_8_24# 0.17fF
C43357 OR2X1_LOC_92/Y AND2X1_LOC_687/A 0.02fF
C45295 OR2X1_LOC_92/Y OR2X1_LOC_12/Y 7.34fF
C45389 OR2X1_LOC_422/a_8_216# OR2X1_LOC_92/Y 0.02fF
C45550 OR2X1_LOC_92/Y AND2X1_LOC_801/B 0.01fF
C47131 OR2X1_LOC_597/A OR2X1_LOC_92/Y 0.02fF
C47186 OR2X1_LOC_256/Y OR2X1_LOC_92/Y 0.07fF
C48101 OR2X1_LOC_18/Y OR2X1_LOC_92/Y 0.30fF
C48569 OR2X1_LOC_92/Y OR2X1_LOC_585/A 0.14fF
C49142 OR2X1_LOC_92/Y OR2X1_LOC_437/A 0.41fF
C49403 OR2X1_LOC_92/Y OR2X1_LOC_753/A 0.17fF
C49989 OR2X1_LOC_92/Y OR2X1_LOC_88/Y 0.06fF
C50124 OR2X1_LOC_8/Y OR2X1_LOC_92/Y 0.02fF
C50226 OR2X1_LOC_92/Y OR2X1_LOC_67/A 0.12fF
C50250 OR2X1_LOC_92/Y OR2X1_LOC_52/B 0.27fF
C50752 OR2X1_LOC_22/Y OR2X1_LOC_92/Y 0.39fF
C50820 OR2X1_LOC_92/Y OR2X1_LOC_387/a_8_216# 0.01fF
C51048 OR2X1_LOC_92/Y OR2X1_LOC_39/A 0.10fF
C51171 OR2X1_LOC_92/Y OR2X1_LOC_760/a_8_216# 0.06fF
C51407 OR2X1_LOC_421/a_8_216# OR2X1_LOC_92/Y 0.03fF
C51475 OR2X1_LOC_92/Y OR2X1_LOC_85/A 0.18fF
C51808 OR2X1_LOC_51/Y OR2X1_LOC_92/Y 0.06fF
C52909 OR2X1_LOC_92/Y OR2X1_LOC_86/A 0.07fF
C53305 OR2X1_LOC_92/Y OR2X1_LOC_599/Y 0.18fF
C53656 OR2X1_LOC_387/Y OR2X1_LOC_92/Y 0.01fF
C53830 OR2X1_LOC_92/Y OR2X1_LOC_268/Y 0.05fF
C54026 OR2X1_LOC_92/Y AND2X1_LOC_294/a_8_24# 0.01fF
C54753 OR2X1_LOC_91/A OR2X1_LOC_92/Y 0.64fF
C55769 OR2X1_LOC_490/Y OR2X1_LOC_92/Y 0.10fF
C55770 OR2X1_LOC_92/Y OR2X1_LOC_74/A 0.07fF
C57173 OR2X1_LOC_92/Y VSS 0.90fF
C11 AND2X1_LOC_40/Y AND2X1_LOC_48/A 0.42fF
C1440 AND2X1_LOC_48/A AND2X1_LOC_519/a_8_24# 0.10fF
C2239 OR2X1_LOC_687/Y AND2X1_LOC_48/A 0.03fF
C3032 AND2X1_LOC_48/A OR2X1_LOC_78/A 0.01fF
C3117 AND2X1_LOC_48/A OR2X1_LOC_155/A 0.07fF
C3963 AND2X1_LOC_387/B AND2X1_LOC_48/A 0.08fF
C4301 AND2X1_LOC_12/Y AND2X1_LOC_48/A 0.22fF
C4717 AND2X1_LOC_59/Y AND2X1_LOC_48/A 2.09fF
C5481 AND2X1_LOC_763/a_8_24# AND2X1_LOC_48/A 0.03fF
C6930 AND2X1_LOC_48/A OR2X1_LOC_520/A 0.01fF
C7382 AND2X1_LOC_48/A AND2X1_LOC_692/a_8_24# 0.04fF
C7637 AND2X1_LOC_387/a_8_24# AND2X1_LOC_48/A 0.03fF
C7850 AND2X1_LOC_48/A AND2X1_LOC_761/a_8_24# 0.03fF
C8182 OR2X1_LOC_377/A AND2X1_LOC_48/A 0.10fF
C8580 AND2X1_LOC_48/A OR2X1_LOC_78/B 0.40fF
C8634 AND2X1_LOC_48/A OR2X1_LOC_375/A 0.87fF
C10294 OR2X1_LOC_405/A AND2X1_LOC_48/A 0.22fF
C10667 AND2X1_LOC_19/Y AND2X1_LOC_48/A 0.03fF
C12137 AND2X1_LOC_48/A OR2X1_LOC_68/B 0.03fF
C12645 AND2X1_LOC_48/A OR2X1_LOC_598/a_8_216# 0.09fF
C12866 AND2X1_LOC_48/A OR2X1_LOC_87/A 0.02fF
C12939 AND2X1_LOC_48/A OR2X1_LOC_706/B 0.01fF
C13216 OR2X1_LOC_389/A AND2X1_LOC_48/A 0.03fF
C14415 OR2X1_LOC_691/Y AND2X1_LOC_48/A 0.05fF
C15367 OR2X1_LOC_154/A AND2X1_LOC_48/A 0.19fF
C16096 AND2X1_LOC_511/a_8_24# AND2X1_LOC_48/A 0.03fF
C16583 AND2X1_LOC_763/a_36_24# AND2X1_LOC_48/A 0.01fF
C16912 AND2X1_LOC_64/Y AND2X1_LOC_48/A 0.13fF
C16944 AND2X1_LOC_599/a_8_24# AND2X1_LOC_48/A 0.02fF
C17429 OR2X1_LOC_756/B AND2X1_LOC_48/A 0.07fF
C18448 AND2X1_LOC_48/A AND2X1_LOC_692/a_36_24# 0.01fF
C18694 AND2X1_LOC_48/A OR2X1_LOC_596/A 0.03fF
C18827 AND2X1_LOC_48/A OR2X1_LOC_87/B 0.21fF
C19297 AND2X1_LOC_48/A OR2X1_LOC_532/B 0.04fF
C20519 OR2X1_LOC_185/Y AND2X1_LOC_48/A 0.02fF
C21278 VDD AND2X1_LOC_48/A 0.42fF
C24074 AND2X1_LOC_48/A OR2X1_LOC_750/Y 0.04fF
C24335 OR2X1_LOC_160/A AND2X1_LOC_48/A 0.03fF
C24805 AND2X1_LOC_48/A AND2X1_LOC_46/a_8_24# 0.01fF
C25527 AND2X1_LOC_48/A AND2X1_LOC_693/a_8_24# 0.01fF
C25567 OR2X1_LOC_185/A AND2X1_LOC_48/A 0.02fF
C26820 AND2X1_LOC_753/a_8_24# AND2X1_LOC_48/A 0.01fF
C28547 AND2X1_LOC_56/B AND2X1_LOC_48/A 0.10fF
C28559 AND2X1_LOC_48/A AND2X1_LOC_8/Y 0.03fF
C29687 AND2X1_LOC_48/A OR2X1_LOC_596/a_8_216# 0.02fF
C29880 AND2X1_LOC_48/A AND2X1_LOC_47/Y 0.10fF
C30341 AND2X1_LOC_48/A AND2X1_LOC_48/Y 0.01fF
C30612 AND2X1_LOC_95/Y AND2X1_LOC_48/A 0.10fF
C30927 AND2X1_LOC_22/Y AND2X1_LOC_48/A 1.14fF
C31032 AND2X1_LOC_48/A OR2X1_LOC_706/A 0.03fF
C32003 AND2X1_LOC_48/A OR2X1_LOC_779/B 0.32fF
C32205 AND2X1_LOC_70/Y AND2X1_LOC_48/A 0.17fF
C32642 AND2X1_LOC_511/a_36_24# AND2X1_LOC_48/A 0.01fF
C33892 AND2X1_LOC_48/A AND2X1_LOC_44/Y 8.45fF
C34767 AND2X1_LOC_48/A AND2X1_LOC_18/Y 0.60fF
C35165 AND2X1_LOC_48/A OR2X1_LOC_596/a_36_216# 0.02fF
C35700 AND2X1_LOC_48/A OR2X1_LOC_130/A 0.03fF
C37524 AND2X1_LOC_48/A OR2X1_LOC_513/a_8_216# 0.12fF
C37777 OR2X1_LOC_790/B AND2X1_LOC_48/A 0.01fF
C37781 AND2X1_LOC_48/A OR2X1_LOC_161/A 0.13fF
C38604 AND2X1_LOC_41/A AND2X1_LOC_48/A 0.22fF
C40047 AND2X1_LOC_48/A AND2X1_LOC_31/Y 0.14fF
C40977 AND2X1_LOC_48/A AND2X1_LOC_36/Y 0.59fF
C43409 AND2X1_LOC_48/A OR2X1_LOC_269/B 0.49fF
C44995 AND2X1_LOC_48/A OR2X1_LOC_161/B 0.07fF
C45090 AND2X1_LOC_48/A AND2X1_LOC_48/a_8_24# 0.01fF
C46095 AND2X1_LOC_48/A AND2X1_LOC_53/Y 0.02fF
C46424 OR2X1_LOC_502/A AND2X1_LOC_48/A 0.03fF
C46937 AND2X1_LOC_48/A AND2X1_LOC_3/Y 0.29fF
C47655 AND2X1_LOC_48/A AND2X1_LOC_7/B 0.28fF
C48796 AND2X1_LOC_48/A OR2X1_LOC_513/Y 0.01fF
C49407 OR2X1_LOC_160/B AND2X1_LOC_48/A 4.50fF
C54856 AND2X1_LOC_48/A OR2X1_LOC_66/A 0.13fF
C56187 OR2X1_LOC_598/Y AND2X1_LOC_48/A 0.17fF
C57365 AND2X1_LOC_48/A VSS 0.55fF
C1 OR2X1_LOC_246/Y OR2X1_LOC_585/A 0.09fF
C288 OR2X1_LOC_585/A OR2X1_LOC_16/A 0.21fF
C511 AND2X1_LOC_687/Y OR2X1_LOC_585/A 0.01fF
C1382 AND2X1_LOC_729/B OR2X1_LOC_585/A 0.06fF
C2200 OR2X1_LOC_599/A OR2X1_LOC_585/A 0.01fF
C2507 OR2X1_LOC_40/Y OR2X1_LOC_585/A 0.20fF
C2666 OR2X1_LOC_7/A OR2X1_LOC_585/A 0.15fF
C3325 OR2X1_LOC_585/A AND2X1_LOC_415/a_8_24# 0.03fF
C3743 OR2X1_LOC_589/A OR2X1_LOC_585/A 0.03fF
C3856 AND2X1_LOC_398/a_8_24# OR2X1_LOC_585/A 0.01fF
C4180 OR2X1_LOC_585/A OR2X1_LOC_585/Y 0.01fF
C4714 OR2X1_LOC_3/Y OR2X1_LOC_585/A 0.21fF
C5001 OR2X1_LOC_329/B OR2X1_LOC_585/A 0.21fF
C5032 OR2X1_LOC_502/A OR2X1_LOC_585/A 0.03fF
C5945 OR2X1_LOC_11/Y OR2X1_LOC_585/A 0.04fF
C5967 OR2X1_LOC_690/A OR2X1_LOC_585/A 0.03fF
C6001 OR2X1_LOC_64/Y OR2X1_LOC_585/A 0.88fF
C9380 OR2X1_LOC_517/A OR2X1_LOC_585/A 0.75fF
C9596 OR2X1_LOC_585/A OR2X1_LOC_150/a_8_216# 0.01fF
C10371 OR2X1_LOC_234/a_8_216# OR2X1_LOC_585/A 0.01fF
C10641 AND2X1_LOC_143/a_36_24# OR2X1_LOC_585/A 0.01fF
C10704 OR2X1_LOC_585/A OR2X1_LOC_49/a_8_216# 0.01fF
C10726 OR2X1_LOC_48/Y OR2X1_LOC_585/A 0.03fF
C11499 OR2X1_LOC_585/A OR2X1_LOC_278/Y 0.04fF
C11510 OR2X1_LOC_585/A OR2X1_LOC_38/a_8_216# 0.01fF
C11523 OR2X1_LOC_95/a_8_216# OR2X1_LOC_585/A 0.03fF
C11603 AND2X1_LOC_800/a_8_24# OR2X1_LOC_585/A 0.01fF
C12627 OR2X1_LOC_585/A AND2X1_LOC_407/a_8_24# 0.01fF
C12913 OR2X1_LOC_689/Y OR2X1_LOC_585/A 0.01fF
C13268 OR2X1_LOC_36/Y OR2X1_LOC_585/A 0.16fF
C13668 OR2X1_LOC_80/Y OR2X1_LOC_585/A 0.02fF
C14179 OR2X1_LOC_255/a_8_216# OR2X1_LOC_585/A 0.01fF
C14905 OR2X1_LOC_399/A OR2X1_LOC_585/A 0.01fF
C16511 AND2X1_LOC_377/Y OR2X1_LOC_585/A 0.06fF
C16885 OR2X1_LOC_585/A OR2X1_LOC_12/Y 0.19fF
C17105 AND2X1_LOC_671/a_8_24# OR2X1_LOC_585/A 0.23fF
C17125 AND2X1_LOC_801/B OR2X1_LOC_585/A 0.01fF
C17378 OR2X1_LOC_585/A OR2X1_LOC_234/Y 0.35fF
C18705 OR2X1_LOC_256/Y OR2X1_LOC_585/A 0.13fF
C19596 OR2X1_LOC_18/Y OR2X1_LOC_585/A 0.10fF
C20646 OR2X1_LOC_585/A OR2X1_LOC_437/A 0.26fF
C20922 OR2X1_LOC_585/A OR2X1_LOC_753/A 0.45fF
C21659 OR2X1_LOC_8/Y OR2X1_LOC_585/A 0.21fF
C21752 OR2X1_LOC_585/A OR2X1_LOC_67/A 0.16fF
C21793 OR2X1_LOC_585/A OR2X1_LOC_52/B 0.62fF
C22121 AND2X1_LOC_378/a_8_24# OR2X1_LOC_585/A 0.01fF
C22263 OR2X1_LOC_22/Y OR2X1_LOC_585/A 0.40fF
C22321 OR2X1_LOC_585/A OR2X1_LOC_387/a_8_216# 0.06fF
C22624 OR2X1_LOC_585/A OR2X1_LOC_39/A 0.10fF
C22748 OR2X1_LOC_760/a_8_216# OR2X1_LOC_585/A 0.01fF
C23042 OR2X1_LOC_377/A OR2X1_LOC_585/A 0.03fF
C23058 OR2X1_LOC_85/A OR2X1_LOC_585/A 0.06fF
C23381 OR2X1_LOC_51/Y OR2X1_LOC_585/A 0.14fF
C24828 OR2X1_LOC_599/Y OR2X1_LOC_585/A 0.04fF
C25157 OR2X1_LOC_387/Y OR2X1_LOC_585/A 0.01fF
C25214 OR2X1_LOC_416/A OR2X1_LOC_585/A 0.02fF
C25559 OR2X1_LOC_585/A AND2X1_LOC_294/a_8_24# 0.11fF
C26286 OR2X1_LOC_91/A OR2X1_LOC_585/A 0.06fF
C26783 OR2X1_LOC_32/B OR2X1_LOC_585/A 0.07fF
C26826 OR2X1_LOC_233/a_8_216# OR2X1_LOC_585/A 0.01fF
C27270 OR2X1_LOC_74/A OR2X1_LOC_585/A 0.02fF
C27565 OR2X1_LOC_459/A OR2X1_LOC_585/A 0.15fF
C27927 OR2X1_LOC_329/a_8_216# OR2X1_LOC_585/A 0.01fF
C31069 OR2X1_LOC_485/A OR2X1_LOC_585/A 0.08fF
C31128 OR2X1_LOC_10/a_8_216# OR2X1_LOC_585/A 0.01fF
C31411 OR2X1_LOC_256/a_8_216# OR2X1_LOC_585/A 0.01fF
C33680 OR2X1_LOC_760/Y OR2X1_LOC_585/A 0.01fF
C34717 AND2X1_LOC_691/a_8_24# OR2X1_LOC_585/A 0.01fF
C35963 VDD OR2X1_LOC_585/A 1.48fF
C36027 OR2X1_LOC_689/A OR2X1_LOC_585/A 0.01fF
C36153 OR2X1_LOC_256/A OR2X1_LOC_585/A 0.04fF
C37288 OR2X1_LOC_427/A OR2X1_LOC_585/A 0.03fF
C38176 OR2X1_LOC_585/A OR2X1_LOC_6/A 0.45fF
C38621 OR2X1_LOC_585/A OR2X1_LOC_44/Y 0.20fF
C38889 OR2X1_LOC_45/B OR2X1_LOC_585/A 0.19fF
C38911 OR2X1_LOC_102/a_8_216# OR2X1_LOC_585/A 0.01fF
C39342 OR2X1_LOC_158/A OR2X1_LOC_585/A 0.14fF
C40810 OR2X1_LOC_411/a_8_216# OR2X1_LOC_585/A 0.06fF
C41228 OR2X1_LOC_293/a_8_216# OR2X1_LOC_585/A 0.03fF
C41956 OR2X1_LOC_744/A OR2X1_LOC_585/A 0.14fF
C42133 OR2X1_LOC_31/Y OR2X1_LOC_585/A 0.08fF
C43257 OR2X1_LOC_585/A OR2X1_LOC_56/A 0.16fF
C43369 AND2X1_LOC_8/Y OR2X1_LOC_585/A 0.08fF
C44296 AND2X1_LOC_68/a_8_24# OR2X1_LOC_585/A 0.02fF
C44617 OR2X1_LOC_625/a_8_216# OR2X1_LOC_585/A 0.19fF
C45351 OR2X1_LOC_585/A OR2X1_LOC_585/a_8_216# 0.05fF
C45352 OR2X1_LOC_585/A OR2X1_LOC_15/a_8_216# 0.01fF
C45416 OR2X1_LOC_426/B OR2X1_LOC_585/A 0.03fF
C45597 OR2X1_LOC_246/A OR2X1_LOC_585/A 0.06fF
C45620 OR2X1_LOC_409/B OR2X1_LOC_585/A 0.01fF
C45689 OR2X1_LOC_585/A OR2X1_LOC_599/a_8_216# 0.01fF
C46797 OR2X1_LOC_235/B OR2X1_LOC_585/A 0.11fF
C48483 OR2X1_LOC_585/A OR2X1_LOC_414/Y 0.03fF
C48682 OR2X1_LOC_62/a_8_216# OR2X1_LOC_585/A 0.01fF
C48920 OR2X1_LOC_600/A OR2X1_LOC_585/A 7.57fF
C49001 OR2X1_LOC_619/Y OR2X1_LOC_585/A 0.03fF
C49471 OR2X1_LOC_690/a_8_216# OR2X1_LOC_585/A 0.01fF
C50178 OR2X1_LOC_329/Y OR2X1_LOC_585/A 0.01fF
C50304 OR2X1_LOC_585/A OR2X1_LOC_69/A 0.04fF
C50982 OR2X1_LOC_585/A OR2X1_LOC_585/a_36_216# 0.02fF
C51303 OR2X1_LOC_585/A OR2X1_LOC_13/B 1.20fF
C51818 OR2X1_LOC_585/A OR2X1_LOC_428/A 0.10fF
C52786 OR2X1_LOC_689/a_8_216# OR2X1_LOC_585/A 0.01fF
C52836 AND2X1_LOC_598/a_8_24# OR2X1_LOC_585/A 0.01fF
C52847 OR2X1_LOC_26/Y OR2X1_LOC_585/A 6.19fF
C53249 OR2X1_LOC_246/a_8_216# OR2X1_LOC_585/A 0.01fF
C53782 OR2X1_LOC_95/Y OR2X1_LOC_585/A 1.71fF
C54664 OR2X1_LOC_585/A OR2X1_LOC_71/A 0.10fF
C54827 OR2X1_LOC_585/A OR2X1_LOC_59/Y 3.43fF
C54955 OR2X1_LOC_70/Y OR2X1_LOC_585/A 0.09fF
C55462 OR2X1_LOC_47/Y OR2X1_LOC_585/A 0.79fF
C55739 AND2X1_LOC_143/a_8_24# OR2X1_LOC_585/A 0.05fF
C55773 OR2X1_LOC_625/Y OR2X1_LOC_585/A 0.01fF
C56836 OR2X1_LOC_585/A VSS 0.37fF
C2077 OR2X1_LOC_502/A OR2X1_LOC_459/B 0.01fF
C2095 OR2X1_LOC_687/Y OR2X1_LOC_502/A 0.07fF
C2545 OR2X1_LOC_502/A OR2X1_LOC_828/B 0.31fF
C2571 AND2X1_LOC_64/a_8_24# OR2X1_LOC_502/A 0.01fF
C2890 OR2X1_LOC_502/A OR2X1_LOC_78/A 1.30fF
C3010 OR2X1_LOC_502/A OR2X1_LOC_155/A 0.20fF
C3849 AND2X1_LOC_387/B OR2X1_LOC_502/A 0.01fF
C4172 OR2X1_LOC_100/a_8_216# OR2X1_LOC_502/A 0.01fF
C4182 AND2X1_LOC_12/Y OR2X1_LOC_502/A 0.16fF
C4217 AND2X1_LOC_376/a_8_24# OR2X1_LOC_502/A 0.01fF
C4589 AND2X1_LOC_59/Y OR2X1_LOC_502/A 0.62fF
C4835 OR2X1_LOC_502/A AND2X1_LOC_762/a_8_24# 0.01fF
C5046 OR2X1_LOC_502/A AND2X1_LOC_43/a_8_24# 0.01fF
C5903 OR2X1_LOC_502/A OR2X1_LOC_753/A 0.05fF
C6837 OR2X1_LOC_502/A OR2X1_LOC_818/a_36_216# 0.02fF
C7169 AND2X1_LOC_81/B OR2X1_LOC_502/A -0.01fF
C8031 OR2X1_LOC_502/A AND2X1_LOC_278/a_8_24# 0.08fF
C8036 OR2X1_LOC_377/A OR2X1_LOC_502/A 0.07fF
C8435 OR2X1_LOC_502/A OR2X1_LOC_78/B 1.39fF
C8491 AND2X1_LOC_94/a_8_24# OR2X1_LOC_502/A 0.01fF
C8510 OR2X1_LOC_502/A OR2X1_LOC_375/A 0.20fF
C9635 OR2X1_LOC_502/A AND2X1_LOC_65/A 0.06fF
C10040 OR2X1_LOC_502/A AND2X1_LOC_433/a_8_24# 0.01fF
C10109 AND2X1_LOC_164/a_36_24# OR2X1_LOC_502/A 0.01fF
C10168 OR2X1_LOC_405/A OR2X1_LOC_502/A 3.75fF
C10320 OR2X1_LOC_502/A AND2X1_LOC_8/a_8_24# 0.03fF
C10655 OR2X1_LOC_502/A OR2X1_LOC_195/A 0.02fF
C11267 AND2X1_LOC_588/B OR2X1_LOC_502/A 0.05fF
C11917 OR2X1_LOC_502/A AND2X1_LOC_4/a_8_24# 0.01fF
C12039 OR2X1_LOC_502/A OR2X1_LOC_68/B 0.43fF
C12733 OR2X1_LOC_502/A OR2X1_LOC_87/A 0.14fF
C12742 OR2X1_LOC_502/A AND2X1_LOC_696/a_8_24# 0.03fF
C13210 OR2X1_LOC_502/A AND2X1_LOC_611/a_8_24# 0.01fF
C13506 OR2X1_LOC_502/A AND2X1_LOC_144/a_8_24# 0.07fF
C15243 OR2X1_LOC_154/A OR2X1_LOC_502/A 0.21fF
C15526 OR2X1_LOC_502/A OR2X1_LOC_435/A 0.01fF
C15894 OR2X1_LOC_502/A AND2X1_LOC_409/B 0.09fF
C15949 AND2X1_LOC_511/a_8_24# OR2X1_LOC_502/A 0.01fF
C16772 AND2X1_LOC_64/Y OR2X1_LOC_502/A 0.39fF
C16892 OR2X1_LOC_502/A AND2X1_LOC_819/a_8_24# 0.03fF
C17306 OR2X1_LOC_756/B OR2X1_LOC_502/A 0.03fF
C17823 OR2X1_LOC_502/A AND2X1_LOC_18/a_8_24# 0.02fF
C17874 OR2X1_LOC_611/a_8_216# OR2X1_LOC_502/A 0.47fF
C18542 OR2X1_LOC_502/A OR2X1_LOC_596/A 0.04fF
C18719 OR2X1_LOC_502/A AND2X1_LOC_612/B 0.40fF
C19047 OR2X1_LOC_100/Y OR2X1_LOC_502/A 0.04fF
C19203 OR2X1_LOC_502/A OR2X1_LOC_532/B 0.18fF
C20392 OR2X1_LOC_185/Y OR2X1_LOC_502/A 0.07fF
C21050 OR2X1_LOC_502/A OR2X1_LOC_502/Y 0.01fF
C21135 VDD OR2X1_LOC_502/A 1.23fF
C21643 OR2X1_LOC_502/A AND2X1_LOC_328/a_8_24# 0.02fF
C22469 OR2X1_LOC_502/A AND2X1_LOC_306/a_8_24# 0.05fF
C23842 OR2X1_LOC_502/A AND2X1_LOC_696/a_36_24# 0.01fF
C24221 OR2X1_LOC_160/A OR2X1_LOC_502/A 0.45fF
C24514 AND2X1_LOC_95/a_8_24# OR2X1_LOC_502/A 0.01fF
C24548 OR2X1_LOC_502/A AND2X1_LOC_144/a_36_24# 0.01fF
C24569 OR2X1_LOC_325/A OR2X1_LOC_502/A 0.11fF
C24597 OR2X1_LOC_502/A OR2X1_LOC_847/A 0.03fF
C25426 OR2X1_LOC_185/A OR2X1_LOC_502/A 0.31fF
C26205 AND2X1_LOC_588/a_8_24# OR2X1_LOC_502/A 0.03fF
C26863 OR2X1_LOC_502/A AND2X1_LOC_8/a_36_24# 0.01fF
C27499 OR2X1_LOC_264/Y OR2X1_LOC_502/A 0.03fF
C27810 AND2X1_LOC_91/B OR2X1_LOC_502/A 3.91fF
C27921 OR2X1_LOC_502/A AND2X1_LOC_819/a_36_24# 0.01fF
C28198 OR2X1_LOC_502/A OR2X1_LOC_446/B 0.10fF
C28426 OR2X1_LOC_502/A AND2X1_LOC_56/B 0.17fF
C28442 OR2X1_LOC_502/A AND2X1_LOC_8/Y 0.07fF
C28458 OR2X1_LOC_502/A AND2X1_LOC_21/Y 0.50fF
C29260 OR2X1_LOC_502/A OR2X1_LOC_83/A 0.02fF
C29795 OR2X1_LOC_502/A AND2X1_LOC_47/Y 0.87fF
C30087 OR2X1_LOC_502/A OR2X1_LOC_506/A 6.75fF
C30247 OR2X1_LOC_502/A AND2X1_LOC_48/Y 0.02fF
C30470 OR2X1_LOC_502/A AND2X1_LOC_414/a_8_24# 0.05fF
C30484 AND2X1_LOC_95/Y OR2X1_LOC_502/A 0.24fF
C30587 OR2X1_LOC_502/A OR2X1_LOC_415/a_8_216# 0.05fF
C30778 AND2X1_LOC_22/Y OR2X1_LOC_502/A 0.33fF
C31707 OR2X1_LOC_235/B OR2X1_LOC_502/A 0.07fF
C31927 OR2X1_LOC_502/A OR2X1_LOC_779/B 1.53fF
C32024 OR2X1_LOC_709/A OR2X1_LOC_502/A 0.14fF
C32070 AND2X1_LOC_70/Y OR2X1_LOC_502/A 0.32fF
C33008 OR2X1_LOC_502/A AND2X1_LOC_11/Y 0.08fF
C33399 OR2X1_LOC_502/A AND2X1_LOC_306/a_36_24# 0.02fF
C33750 OR2X1_LOC_502/A AND2X1_LOC_44/Y 7.63fF
C33945 OR2X1_LOC_502/A AND2X1_LOC_36/a_8_24# 0.01fF
C34615 OR2X1_LOC_502/A AND2X1_LOC_18/Y 2.19fF
C35576 OR2X1_LOC_502/A OR2X1_LOC_130/A 0.87fF
C35708 OR2X1_LOC_502/A AND2X1_LOC_88/Y 0.02fF
C37649 OR2X1_LOC_502/A OR2X1_LOC_161/A 0.18fF
C37676 OR2X1_LOC_502/A AND2X1_LOC_25/Y 0.02fF
C37738 OR2X1_LOC_502/A AND2X1_LOC_51/Y 1.81fF
C38456 OR2X1_LOC_502/A AND2X1_LOC_41/A 0.13fF
C38951 OR2X1_LOC_502/A OR2X1_LOC_405/a_8_216# 0.03fF
C39602 OR2X1_LOC_502/A OR2X1_LOC_71/A 0.11fF
C39964 OR2X1_LOC_502/A AND2X1_LOC_31/Y 0.36fF
C40237 OR2X1_LOC_502/A OR2X1_LOC_240/A 0.03fF
C40599 AND2X1_LOC_143/a_8_24# OR2X1_LOC_502/A 0.02fF
C40860 OR2X1_LOC_502/A AND2X1_LOC_36/Y 0.99fF
C41369 OR2X1_LOC_502/A OR2X1_LOC_16/A 0.05fF
C43284 OR2X1_LOC_502/A AND2X1_LOC_26/a_8_24# 0.01fF
C43290 OR2X1_LOC_502/A OR2X1_LOC_269/B 0.50fF
C44078 OR2X1_LOC_502/A AND2X1_LOC_304/a_8_24# 0.03fF
C44108 OR2X1_LOC_502/A AND2X1_LOC_59/a_8_24# 0.04fF
C44354 OR2X1_LOC_502/A OR2X1_LOC_777/B 0.12fF
C44845 OR2X1_LOC_502/A OR2X1_LOC_161/B 0.23fF
C44932 OR2X1_LOC_502/A AND2X1_LOC_48/a_8_24# 0.01fF
C45925 OR2X1_LOC_3/Y OR2X1_LOC_502/A 0.03fF
C45989 OR2X1_LOC_502/A AND2X1_LOC_53/Y 0.01fF
C46074 OR2X1_LOC_502/A AND2X1_LOC_409/a_8_24# 0.01fF
C46830 OR2X1_LOC_502/A AND2X1_LOC_3/Y 0.37fF
C47523 OR2X1_LOC_502/A AND2X1_LOC_7/B 4.98fF
C48982 AND2X1_LOC_386/a_8_24# OR2X1_LOC_502/A 0.01fF
C49246 OR2X1_LOC_160/B OR2X1_LOC_502/A 0.10fF
C49748 OR2X1_LOC_502/A OR2X1_LOC_307/B 0.04fF
C49787 OR2X1_LOC_327/a_8_216# OR2X1_LOC_502/A 0.05fF
C50094 OR2X1_LOC_151/A OR2X1_LOC_502/A 0.57fF
C50108 AND2X1_LOC_322/a_8_24# OR2X1_LOC_502/A 0.04fF
C51298 OR2X1_LOC_502/A OR2X1_LOC_415/Y 0.02fF
C51661 OR2X1_LOC_502/A OR2X1_LOC_460/A 0.01fF
C51995 OR2X1_LOC_502/A OR2X1_LOC_818/a_8_216# 0.01fF
C52317 AND2X1_LOC_80/a_8_24# OR2X1_LOC_502/A 0.01fF
C52723 OR2X1_LOC_502/A AND2X1_LOC_414/a_36_24# 0.01fF
C53040 AND2X1_LOC_534/a_8_24# OR2X1_LOC_502/A -0.01fF
C54728 OR2X1_LOC_502/A OR2X1_LOC_66/A 0.28fF
C55065 OR2X1_LOC_502/A OR2X1_LOC_502/a_8_216# 0.01fF
C55191 AND2X1_LOC_94/Y OR2X1_LOC_502/A 0.03fF
C55193 AND2X1_LOC_164/a_8_24# OR2X1_LOC_502/A 0.01fF
C55227 AND2X1_LOC_50/Y OR2X1_LOC_502/A 0.06fF
C55574 OR2X1_LOC_325/B OR2X1_LOC_502/A 0.06fF
C55689 OR2X1_LOC_502/A OR2X1_LOC_405/Y 0.03fF
C56082 AND2X1_LOC_40/Y OR2X1_LOC_502/A 0.16fF
C57516 OR2X1_LOC_502/A VSS 0.69fF
C14 OR2X1_LOC_155/A OR2X1_LOC_269/B 0.10fF
C810 AND2X1_LOC_304/a_8_24# OR2X1_LOC_155/A 0.06fF
C1130 OR2X1_LOC_155/A OR2X1_LOC_831/B 0.11fF
C1591 OR2X1_LOC_155/A OR2X1_LOC_161/B 0.15fF
C3491 AND2X1_LOC_3/Y OR2X1_LOC_155/A 0.15fF
C4106 OR2X1_LOC_155/A AND2X1_LOC_7/B 0.14fF
C5220 OR2X1_LOC_155/A OR2X1_LOC_513/Y 0.02fF
C5841 OR2X1_LOC_160/B OR2X1_LOC_155/A 0.21fF
C6664 OR2X1_LOC_151/A OR2X1_LOC_155/A 0.07fF
C10455 OR2X1_LOC_155/A OR2X1_LOC_515/a_8_216# -0.02fF
C11415 OR2X1_LOC_155/A OR2X1_LOC_66/A 0.03fF
C12437 AND2X1_LOC_136/a_36_24# OR2X1_LOC_155/A 0.01fF
C12672 OR2X1_LOC_831/A OR2X1_LOC_155/A 0.17fF
C12685 OR2X1_LOC_598/Y OR2X1_LOC_155/A 0.30fF
C12752 AND2X1_LOC_40/Y OR2X1_LOC_155/A 2.28fF
C14933 OR2X1_LOC_687/Y OR2X1_LOC_155/A 0.53fF
C15650 OR2X1_LOC_155/A OR2X1_LOC_78/A 0.54fF
C16632 AND2X1_LOC_387/B OR2X1_LOC_155/A 0.07fF
C17022 AND2X1_LOC_12/Y OR2X1_LOC_155/A 0.06fF
C17367 OR2X1_LOC_168/B OR2X1_LOC_155/A 0.03fF
C17425 AND2X1_LOC_59/Y OR2X1_LOC_155/A 0.09fF
C20882 OR2X1_LOC_377/A OR2X1_LOC_155/A 0.01fF
C21243 OR2X1_LOC_155/A OR2X1_LOC_78/B 0.19fF
C21336 OR2X1_LOC_375/A OR2X1_LOC_155/A 0.04fF
C21529 OR2X1_LOC_155/A OR2X1_LOC_515/Y 0.04fF
C23038 OR2X1_LOC_405/A OR2X1_LOC_155/A 0.03fF
C24546 OR2X1_LOC_155/A OR2X1_LOC_138/A 0.05fF
C24812 AND2X1_LOC_681/a_8_24# OR2X1_LOC_155/A 0.06fF
C24848 OR2X1_LOC_155/A OR2X1_LOC_68/B 0.01fF
C25535 OR2X1_LOC_87/A OR2X1_LOC_155/A 0.15fF
C27210 AND2X1_LOC_699/a_36_24# OR2X1_LOC_155/A -0.01fF
C28071 OR2X1_LOC_154/A OR2X1_LOC_155/A 0.24fF
C28359 OR2X1_LOC_155/A OR2X1_LOC_435/A 0.01fF
C29558 AND2X1_LOC_64/Y OR2X1_LOC_155/A 0.11fF
C30112 OR2X1_LOC_756/B OR2X1_LOC_155/A 0.03fF
C30694 AND2X1_LOC_699/a_8_24# OR2X1_LOC_155/A 0.01fF
C31317 OR2X1_LOC_155/A OR2X1_LOC_596/A 0.05fF
C31919 OR2X1_LOC_532/B OR2X1_LOC_155/A 0.03fF
C33120 OR2X1_LOC_185/Y OR2X1_LOC_155/A 0.07fF
C33887 VDD OR2X1_LOC_155/A 0.67fF
C36867 OR2X1_LOC_160/A OR2X1_LOC_155/A 1.05fF
C37152 AND2X1_LOC_743/a_8_24# OR2X1_LOC_155/A 0.01fF
C37327 OR2X1_LOC_685/B OR2X1_LOC_155/A 0.02fF
C38140 OR2X1_LOC_185/A OR2X1_LOC_155/A 0.05fF
C40547 AND2X1_LOC_91/B OR2X1_LOC_155/A 0.15fF
C40880 OR2X1_LOC_155/A OR2X1_LOC_446/B 7.07fF
C41171 AND2X1_LOC_56/B OR2X1_LOC_155/A 0.26fF
C42358 OR2X1_LOC_155/A OR2X1_LOC_596/a_8_216# 0.04fF
C42589 AND2X1_LOC_47/Y OR2X1_LOC_155/A 0.19fF
C42885 OR2X1_LOC_506/A OR2X1_LOC_155/A 0.17fF
C43321 AND2X1_LOC_95/Y OR2X1_LOC_155/A 0.03fF
C43620 AND2X1_LOC_22/Y OR2X1_LOC_155/A 0.05fF
C44789 OR2X1_LOC_155/A OR2X1_LOC_779/B 0.03fF
C44925 OR2X1_LOC_709/A OR2X1_LOC_155/A 0.48fF
C44982 AND2X1_LOC_70/Y OR2X1_LOC_155/A 0.29fF
C46202 OR2X1_LOC_155/A AND2X1_LOC_273/a_8_24# 0.12fF
C46685 OR2X1_LOC_155/A AND2X1_LOC_44/Y 0.94fF
C46717 OR2X1_LOC_155/A OR2X1_LOC_514/a_8_216# 0.03fF
C47656 OR2X1_LOC_155/A AND2X1_LOC_18/Y 0.15fF
C47774 OR2X1_LOC_596/Y OR2X1_LOC_155/A 0.04fF
C48335 OR2X1_LOC_155/A OR2X1_LOC_512/a_8_216# 0.02fF
C48691 OR2X1_LOC_780/B OR2X1_LOC_155/A 0.50fF
C50724 OR2X1_LOC_155/A OR2X1_LOC_161/A 0.31fF
C50784 AND2X1_LOC_51/Y OR2X1_LOC_155/A 0.38fF
C51477 AND2X1_LOC_41/A OR2X1_LOC_155/A 0.18fF
C52024 AND2X1_LOC_136/a_8_24# OR2X1_LOC_155/A 0.03fF
C52976 AND2X1_LOC_31/Y OR2X1_LOC_155/A 3.29fF
C53808 OR2X1_LOC_155/A OR2X1_LOC_512/a_36_216# 0.01fF
C53865 OR2X1_LOC_155/A AND2X1_LOC_36/Y 0.11fF
C56778 OR2X1_LOC_155/A VSS -8.81fF
C366 OR2X1_LOC_426/B OR2X1_LOC_485/A 0.06fF
C2853 OR2X1_LOC_310/Y OR2X1_LOC_426/B 0.01fF
C2899 OR2X1_LOC_519/a_8_216# OR2X1_LOC_426/B 0.03fF
C5272 VDD OR2X1_LOC_426/B 2.02fF
C5504 OR2X1_LOC_426/B OR2X1_LOC_256/A 0.07fF
C6625 OR2X1_LOC_426/B OR2X1_LOC_427/A 0.02fF
C6641 OR2X1_LOC_426/B OR2X1_LOC_63/a_8_216# 0.02fF
C7577 OR2X1_LOC_426/B OR2X1_LOC_6/A 0.17fF
C7600 OR2X1_LOC_426/B OR2X1_LOC_299/a_8_216# 0.03fF
C7934 AND2X1_LOC_514/a_36_24# OR2X1_LOC_426/B 0.01fF
C8023 OR2X1_LOC_426/B OR2X1_LOC_44/Y 0.24fF
C8321 OR2X1_LOC_45/B OR2X1_LOC_426/B 0.13fF
C8757 OR2X1_LOC_158/A OR2X1_LOC_426/B 0.14fF
C9378 OR2X1_LOC_426/B OR2X1_LOC_304/Y 0.45fF
C11278 OR2X1_LOC_309/Y OR2X1_LOC_426/B 0.01fF
C11304 OR2X1_LOC_744/A OR2X1_LOC_426/B 0.17fF
C11521 OR2X1_LOC_426/B OR2X1_LOC_31/Y 0.13fF
C12576 OR2X1_LOC_426/B OR2X1_LOC_56/A 0.48fF
C13955 OR2X1_LOC_519/Y OR2X1_LOC_426/B 0.02fF
C14490 OR2X1_LOC_426/B OR2X1_LOC_71/Y 0.08fF
C14893 OR2X1_LOC_426/B OR2X1_LOC_246/A 0.97fF
C14931 OR2X1_LOC_426/B OR2X1_LOC_409/B 0.03fF
C17716 OR2X1_LOC_426/B OR2X1_LOC_65/B 0.28fF
C18078 OR2X1_LOC_426/B OR2X1_LOC_600/A 0.07fF
C18171 OR2X1_LOC_426/B OR2X1_LOC_619/Y 0.08fF
C18194 OR2X1_LOC_426/B OR2X1_LOC_88/A 0.25fF
C19160 OR2X1_LOC_426/B OR2X1_LOC_813/A 0.03fF
C19372 OR2X1_LOC_426/B AND2X1_LOC_606/a_8_24# 0.11fF
C20252 OR2X1_LOC_426/B OR2X1_LOC_666/A 0.18fF
C20572 OR2X1_LOC_426/B OR2X1_LOC_13/B 0.67fF
C21043 OR2X1_LOC_426/B OR2X1_LOC_428/A 0.10fF
C22085 OR2X1_LOC_426/B OR2X1_LOC_26/Y 0.10fF
C22105 OR2X1_LOC_426/B OR2X1_LOC_89/A 1.36fF
C22198 OR2X1_LOC_426/B OR2X1_LOC_92/a_8_216# 0.03fF
C22205 OR2X1_LOC_426/B OR2X1_LOC_426/a_8_216# 0.07fF
C23057 OR2X1_LOC_426/B OR2X1_LOC_95/Y 0.10fF
C23968 OR2X1_LOC_426/B OR2X1_LOC_71/A 0.03fF
C24104 OR2X1_LOC_426/B OR2X1_LOC_59/Y 0.30fF
C24250 OR2X1_LOC_70/Y OR2X1_LOC_426/B 5.79fF
C24741 OR2X1_LOC_426/B OR2X1_LOC_47/Y 0.04fF
C25700 OR2X1_LOC_426/B OR2X1_LOC_16/A 6.52fF
C25738 OR2X1_LOC_426/B AND2X1_LOC_121/a_8_24# 0.02fF
C25867 OR2X1_LOC_426/B OR2X1_LOC_273/a_8_216# 0.01fF
C26260 OR2X1_LOC_426/B AND2X1_LOC_100/a_8_24# 0.01fF
C26729 OR2X1_LOC_426/B AND2X1_LOC_729/B 0.03fF
C27828 OR2X1_LOC_40/Y OR2X1_LOC_426/B 0.67fF
C27978 OR2X1_LOC_426/B OR2X1_LOC_7/A 0.14fF
C28395 OR2X1_LOC_426/B OR2X1_LOC_86/a_8_216# 0.03fF
C29072 OR2X1_LOC_589/A OR2X1_LOC_426/B 0.03fF
C29668 OR2X1_LOC_426/B OR2X1_LOC_299/Y 0.02fF
C30101 OR2X1_LOC_3/Y OR2X1_LOC_426/B 1.56fF
C30393 OR2X1_LOC_329/B OR2X1_LOC_426/B 0.16fF
C31244 OR2X1_LOC_426/B OR2X1_LOC_122/A 0.02fF
C31392 OR2X1_LOC_426/B OR2X1_LOC_64/Y 0.16fF
C34618 OR2X1_LOC_426/B OR2X1_LOC_517/A 0.17fF
C35563 OR2X1_LOC_763/Y OR2X1_LOC_426/B 0.10fF
C35716 OR2X1_LOC_426/B OR2X1_LOC_88/a_8_216# 0.54fF
C36819 OR2X1_LOC_426/B OR2X1_LOC_273/Y 0.15fF
C37258 OR2X1_LOC_426/B OR2X1_LOC_275/A 0.03fF
C37836 OR2X1_LOC_426/B OR2X1_LOC_300/a_8_216# 0.01fF
C38489 OR2X1_LOC_426/B OR2X1_LOC_36/Y 0.68fF
C39642 OR2X1_LOC_490/a_8_216# OR2X1_LOC_426/B 0.02fF
C40871 OR2X1_LOC_426/B OR2X1_LOC_310/a_8_216# 0.02fF
C42210 OR2X1_LOC_426/B OR2X1_LOC_12/Y 5.42fF
C42425 OR2X1_LOC_426/B OR2X1_LOC_272/Y 0.03fF
C44924 OR2X1_LOC_426/B OR2X1_LOC_18/Y 0.20fF
C46063 OR2X1_LOC_426/B OR2X1_LOC_437/A 0.75fF
C46928 OR2X1_LOC_426/B OR2X1_LOC_88/Y 0.19fF
C47093 OR2X1_LOC_8/Y OR2X1_LOC_426/B 0.02fF
C47183 OR2X1_LOC_426/B OR2X1_LOC_67/A 0.17fF
C47222 OR2X1_LOC_426/B OR2X1_LOC_52/B 0.36fF
C47564 AND2X1_LOC_514/a_8_24# OR2X1_LOC_426/B 0.03fF
C47729 OR2X1_LOC_426/B OR2X1_LOC_22/Y 0.37fF
C48069 OR2X1_LOC_426/B OR2X1_LOC_39/A 0.12fF
C48518 OR2X1_LOC_426/B OR2X1_LOC_85/A 0.02fF
C48753 OR2X1_LOC_136/Y OR2X1_LOC_426/B 0.16fF
C48811 OR2X1_LOC_426/B OR2X1_LOC_51/Y 0.02fF
C49927 OR2X1_LOC_426/B OR2X1_LOC_86/A 0.03fF
C50906 OR2X1_LOC_309/a_8_216# OR2X1_LOC_426/B 0.01fF
C51783 OR2X1_LOC_426/B OR2X1_LOC_91/A 0.20fF
C52747 OR2X1_LOC_426/B OR2X1_LOC_74/A 0.13fF
C53217 OR2X1_LOC_426/B OR2X1_LOC_263/a_8_216# 0.31fF
C53926 OR2X1_LOC_426/B OR2X1_LOC_71/a_8_216# 0.05fF
C54597 OR2X1_LOC_426/B OR2X1_LOC_300/Y 0.09fF
C57519 OR2X1_LOC_426/B VSS -6.72fF
C1022 OR2X1_LOC_458/B OR2X1_LOC_777/B 0.03fF
C18591 OR2X1_LOC_458/B OR2X1_LOC_458/a_8_216# 0.13fF
C18654 OR2X1_LOC_458/B AND2X1_LOC_272/a_8_24# 0.20fF
C21225 OR2X1_LOC_458/B OR2X1_LOC_375/A 0.03fF
C22945 OR2X1_LOC_405/A OR2X1_LOC_458/B 0.16fF
C26611 OR2X1_LOC_458/B OR2X1_LOC_541/A 0.02fF
C27975 OR2X1_LOC_154/A OR2X1_LOC_458/B 0.03fF
C31505 OR2X1_LOC_458/B OR2X1_LOC_374/Y 0.11fF
C31851 OR2X1_LOC_458/B OR2X1_LOC_532/B 0.01fF
C33785 OR2X1_LOC_458/B VDD 0.29fF
C44877 OR2X1_LOC_458/B AND2X1_LOC_70/Y 0.03fF
C50615 OR2X1_LOC_458/B OR2X1_LOC_161/A 0.02fF
C52925 OR2X1_LOC_458/B AND2X1_LOC_31/Y 0.11fF
C56161 OR2X1_LOC_458/B OR2X1_LOC_269/B 0.03fF
C57942 OR2X1_LOC_458/B VSS 0.24fF
C88 OR2X1_LOC_8/Y OR2X1_LOC_71/A 0.32fF
C227 OR2X1_LOC_8/Y OR2X1_LOC_59/Y 0.04fF
C902 OR2X1_LOC_8/Y OR2X1_LOC_47/Y 0.06fF
C1619 OR2X1_LOC_8/Y OR2X1_LOC_246/Y 0.10fF
C1772 OR2X1_LOC_8/Y OR2X1_LOC_29/a_8_216# 0.06fF
C1911 OR2X1_LOC_8/Y OR2X1_LOC_16/A 0.08fF
C4064 OR2X1_LOC_8/Y OR2X1_LOC_40/Y 0.07fF
C4136 OR2X1_LOC_8/Y OR2X1_LOC_618/a_8_216# 0.01fF
C4179 OR2X1_LOC_8/Y OR2X1_LOC_7/A 0.03fF
C6532 OR2X1_LOC_133/a_36_216# OR2X1_LOC_8/Y 0.02fF
C6555 OR2X1_LOC_8/Y OR2X1_LOC_671/a_8_216# 0.40fF
C11175 OR2X1_LOC_8/Y OR2X1_LOC_150/a_8_216# 0.01fF
C11351 OR2X1_LOC_8/Y AND2X1_LOC_62/a_8_24# 0.01fF
C13107 OR2X1_LOC_8/Y OR2X1_LOC_278/Y 0.04fF
C14797 OR2X1_LOC_8/Y OR2X1_LOC_36/Y 0.04fF
C15110 OR2X1_LOC_8/Y OR2X1_LOC_604/A 0.08fF
C16716 OR2X1_LOC_143/a_8_216# OR2X1_LOC_8/Y 0.18fF
C17884 OR2X1_LOC_8/Y OR2X1_LOC_619/a_8_216# 0.01fF
C21178 OR2X1_LOC_8/Y OR2X1_LOC_18/Y 0.04fF
C22286 OR2X1_LOC_8/Y OR2X1_LOC_437/A 0.01fF
C22521 OR2X1_LOC_8/Y OR2X1_LOC_753/A 0.23fF
C24577 OR2X1_LOC_8/Y OR2X1_LOC_85/A 0.32fF
C24908 OR2X1_LOC_8/Y OR2X1_LOC_51/Y 0.03fF
C27852 OR2X1_LOC_8/Y OR2X1_LOC_91/A 0.03fF
C28440 OR2X1_LOC_8/Y OR2X1_LOC_5/a_8_216# 0.18fF
C28815 OR2X1_LOC_8/Y OR2X1_LOC_74/A 0.04fF
C30951 OR2X1_LOC_8/Y AND2X1_LOC_37/a_8_24# 0.08fF
C31361 OR2X1_LOC_8/Y OR2X1_LOC_278/a_8_216# 0.14fF
C32614 OR2X1_LOC_8/Y OR2X1_LOC_485/A 1.19fF
C32717 OR2X1_LOC_8/Y OR2X1_LOC_10/a_8_216# 0.06fF
C33026 OR2X1_LOC_8/Y OR2X1_LOC_827/Y 0.02fF
C34314 OR2X1_LOC_8/Y OR2X1_LOC_611/a_8_216# 0.14fF
C35371 OR2X1_LOC_8/Y OR2X1_LOC_671/Y 0.09fF
C37532 OR2X1_LOC_8/Y VDD 0.52fF
C38049 OR2X1_LOC_8/Y OR2X1_LOC_6/a_8_216# 0.02fF
C38902 OR2X1_LOC_8/Y OR2X1_LOC_63/a_8_216# 0.07fF
C39687 OR2X1_LOC_8/Y OR2X1_LOC_104/a_8_216# 0.01fF
C39775 OR2X1_LOC_8/Y OR2X1_LOC_6/A 2.38fF
C40157 OR2X1_LOC_8/Y OR2X1_LOC_44/Y 0.06fF
C40489 OR2X1_LOC_102/a_8_216# OR2X1_LOC_8/Y 0.05fF
C40889 OR2X1_LOC_8/Y OR2X1_LOC_158/A 0.02fF
C40997 OR2X1_LOC_8/Y OR2X1_LOC_847/A 0.34fF
C44855 OR2X1_LOC_8/Y OR2X1_LOC_56/A 0.24fF
C48438 OR2X1_LOC_8/Y OR2X1_LOC_235/B 1.03fF
C49331 OR2X1_LOC_8/Y OR2X1_LOC_96/B 0.18fF
C49369 OR2X1_LOC_8/Y OR2X1_LOC_6/a_36_216# 0.02fF
C50489 OR2X1_LOC_8/Y OR2X1_LOC_600/A 0.21fF
C50571 OR2X1_LOC_8/Y OR2X1_LOC_619/Y 0.16fF
C51736 OR2X1_LOC_133/a_8_216# OR2X1_LOC_8/Y 0.01fF
C52566 OR2X1_LOC_8/Y OR2X1_LOC_15/a_36_216# 0.02fF
C52932 OR2X1_LOC_8/Y OR2X1_LOC_13/B 0.01fF
C53398 OR2X1_LOC_8/Y OR2X1_LOC_428/A 0.07fF
C54387 OR2X1_LOC_8/Y OR2X1_LOC_26/Y 0.05fF
C54797 OR2X1_LOC_8/Y OR2X1_LOC_246/a_8_216# 0.01fF
C55360 OR2X1_LOC_8/Y OR2X1_LOC_95/Y 0.40fF
C57903 OR2X1_LOC_8/Y VSS 0.94fF
C491 AND2X1_LOC_371/a_8_24# OR2X1_LOC_68/B 0.11fF
C493 AND2X1_LOC_18/Y OR2X1_LOC_68/B 0.61fF
C571 AND2X1_LOC_413/a_8_24# OR2X1_LOC_68/B 0.01fF
C1464 OR2X1_LOC_130/A OR2X1_LOC_68/B 0.25fF
C3592 OR2X1_LOC_161/A OR2X1_LOC_68/B 0.04fF
C3640 OR2X1_LOC_461/Y OR2X1_LOC_68/B 0.01fF
C3642 AND2X1_LOC_51/Y OR2X1_LOC_68/B 3.59fF
C4343 AND2X1_LOC_41/A OR2X1_LOC_68/B 0.06fF
C4881 AND2X1_LOC_293/a_8_24# OR2X1_LOC_68/B -0.01fF
C5200 OR2X1_LOC_847/a_8_216# OR2X1_LOC_68/B 0.01fF
C5408 OR2X1_LOC_68/B OR2X1_LOC_71/A 0.08fF
C5613 AND2X1_LOC_749/a_8_24# OR2X1_LOC_68/B 0.03fF
C5825 AND2X1_LOC_31/Y OR2X1_LOC_68/B 0.71fF
C6358 OR2X1_LOC_68/B OR2X1_LOC_121/A 0.03fF
C6627 AND2X1_LOC_72/B OR2X1_LOC_68/B 0.05fF
C6758 AND2X1_LOC_36/Y OR2X1_LOC_68/B 0.25fF
C6798 OR2X1_LOC_68/B OR2X1_LOC_334/A 0.01fF
C7349 OR2X1_LOC_274/Y OR2X1_LOC_68/B 1.56fF
C8688 AND2X1_LOC_71/a_8_24# OR2X1_LOC_68/B 0.02fF
C8990 OR2X1_LOC_68/B OR2X1_LOC_227/A 0.04fF
C9140 OR2X1_LOC_269/B OR2X1_LOC_68/B 0.03fF
C10206 OR2X1_LOC_777/B OR2X1_LOC_68/B 0.03fF
C10264 OR2X1_LOC_831/B OR2X1_LOC_68/B 0.03fF
C10711 OR2X1_LOC_161/B OR2X1_LOC_68/B 0.07fF
C10791 AND2X1_LOC_618/a_8_24# OR2X1_LOC_68/B 0.03fF
C10807 OR2X1_LOC_87/a_8_216# OR2X1_LOC_68/B 0.04fF
C11766 OR2X1_LOC_673/A OR2X1_LOC_68/B 0.14fF
C11792 AND2X1_LOC_462/B OR2X1_LOC_68/B 0.05fF
C12526 AND2X1_LOC_3/Y OR2X1_LOC_68/B 0.11fF
C12973 OR2X1_LOC_690/A OR2X1_LOC_68/B 0.28fF
C13274 AND2X1_LOC_7/B OR2X1_LOC_68/B 0.29fF
C14664 OR2X1_LOC_287/B OR2X1_LOC_68/B 0.04fF
C15000 OR2X1_LOC_160/B OR2X1_LOC_68/B 12.78fF
C15770 OR2X1_LOC_151/A OR2X1_LOC_68/B 0.10fF
C17034 OR2X1_LOC_415/Y OR2X1_LOC_68/B 0.04fF
C17633 OR2X1_LOC_818/a_8_216# OR2X1_LOC_68/B 0.01fF
C18001 AND2X1_LOC_80/a_8_24# OR2X1_LOC_68/B 0.01fF
C20541 OR2X1_LOC_66/A OR2X1_LOC_68/B 0.21fF
C21867 AND2X1_LOC_40/Y OR2X1_LOC_68/B 0.77fF
C21889 OR2X1_LOC_87/Y OR2X1_LOC_68/B 0.02fF
C21893 OR2X1_LOC_848/A OR2X1_LOC_68/B 0.01fF
C22799 AND2X1_LOC_159/a_8_24# OR2X1_LOC_68/B 0.03fF
C23985 AND2X1_LOC_57/a_8_24# OR2X1_LOC_68/B 0.01fF
C24786 OR2X1_LOC_78/A OR2X1_LOC_68/B 0.30fF
C25268 OR2X1_LOC_68/a_8_216# OR2X1_LOC_68/B 0.04fF
C26076 AND2X1_LOC_12/Y OR2X1_LOC_68/B 5.00fF
C26495 AND2X1_LOC_59/Y OR2X1_LOC_68/B 0.20fF
C27781 OR2X1_LOC_753/A OR2X1_LOC_68/B 0.05fF
C28981 AND2X1_LOC_310/a_8_24# OR2X1_LOC_68/B 0.03fF
C29084 OR2X1_LOC_22/Y OR2X1_LOC_68/B 0.03fF
C29452 OR2X1_LOC_39/A OR2X1_LOC_68/B 0.03fF
C29869 AND2X1_LOC_278/a_8_24# OR2X1_LOC_68/B 0.02fF
C29871 OR2X1_LOC_377/A OR2X1_LOC_68/B 0.35fF
C30253 OR2X1_LOC_78/B OR2X1_LOC_68/B 0.55fF
C30302 OR2X1_LOC_375/A OR2X1_LOC_68/B 0.26fF
C30624 OR2X1_LOC_68/B OR2X1_LOC_549/A 0.09fF
C30728 OR2X1_LOC_68/a_36_216# OR2X1_LOC_68/B 0.03fF
C31566 AND2X1_LOC_381/a_8_24# OR2X1_LOC_68/B 0.01fF
C31942 OR2X1_LOC_405/A OR2X1_LOC_68/B 0.02fF
C31992 AND2X1_LOC_77/a_8_24# OR2X1_LOC_68/B 0.01fF
C32312 AND2X1_LOC_19/Y OR2X1_LOC_68/B 0.02fF
C32457 OR2X1_LOC_4/a_8_216# OR2X1_LOC_68/B 0.47fF
C34503 OR2X1_LOC_87/A OR2X1_LOC_68/B 3.45fF
C34979 AND2X1_LOC_611/a_8_24# OR2X1_LOC_68/B 0.02fF
C35332 AND2X1_LOC_291/a_8_24# OR2X1_LOC_68/B 0.01fF
C35404 AND2X1_LOC_5/a_8_24# OR2X1_LOC_68/B 0.05fF
C36559 OR2X1_LOC_778/B OR2X1_LOC_68/B 0.05fF
C37026 OR2X1_LOC_154/A OR2X1_LOC_68/B 0.31fF
C37143 AND2X1_LOC_6/a_8_24# OR2X1_LOC_68/B 0.14fF
C37811 OR2X1_LOC_461/a_8_216# OR2X1_LOC_68/B 0.01fF
C37830 OR2X1_LOC_634/A OR2X1_LOC_68/B 0.06fF
C38205 OR2X1_LOC_633/A OR2X1_LOC_68/B 0.04fF
C38605 AND2X1_LOC_64/Y OR2X1_LOC_68/B 0.22fF
C38649 AND2X1_LOC_82/Y OR2X1_LOC_68/B 0.02fF
C39148 OR2X1_LOC_756/B OR2X1_LOC_68/B 0.10fF
C39189 AND2X1_LOC_55/a_8_24# OR2X1_LOC_68/B 0.01fF
C40443 OR2X1_LOC_87/B OR2X1_LOC_68/B 0.07fF
C40458 AND2X1_LOC_612/B OR2X1_LOC_68/B 0.25fF
C40700 OR2X1_LOC_68/B OR2X1_LOC_333/A 0.17fF
C40797 AND2X1_LOC_529/a_8_24# OR2X1_LOC_68/B 0.01fF
C40929 OR2X1_LOC_532/B OR2X1_LOC_68/B 0.13fF
C42176 OR2X1_LOC_185/Y OR2X1_LOC_68/B 0.11fF
C42989 VDD OR2X1_LOC_68/B 1.42fF
C45220 OR2X1_LOC_6/A OR2X1_LOC_68/B 0.02fF
C46096 OR2X1_LOC_160/A OR2X1_LOC_68/B 0.62fF
C46482 OR2X1_LOC_158/A OR2X1_LOC_68/B 0.03fF
C46536 OR2X1_LOC_847/A OR2X1_LOC_68/B 0.03fF
C47351 AND2X1_LOC_92/a_8_24# OR2X1_LOC_68/B 0.03fF
C47452 OR2X1_LOC_185/A OR2X1_LOC_68/B 0.04fF
C48469 AND2X1_LOC_6/a_36_24# OR2X1_LOC_68/B 0.01fF
C49890 AND2X1_LOC_91/B OR2X1_LOC_68/B 0.31fF
C50451 AND2X1_LOC_56/B OR2X1_LOC_68/B 0.07fF
C50457 AND2X1_LOC_8/Y OR2X1_LOC_68/B 0.12fF
C51627 AND2X1_LOC_73/a_8_24# OR2X1_LOC_68/B 0.01fF
C51761 OR2X1_LOC_68/Y OR2X1_LOC_68/B 0.01fF
C51776 AND2X1_LOC_47/Y OR2X1_LOC_68/B 0.28fF
C52077 OR2X1_LOC_506/A OR2X1_LOC_68/B 0.02fF
C52084 AND2X1_LOC_82/a_8_24# OR2X1_LOC_68/B 0.02fF
C52509 AND2X1_LOC_95/Y OR2X1_LOC_68/B 0.12fF
C52850 AND2X1_LOC_22/Y OR2X1_LOC_68/B 0.68fF
C52962 AND2X1_LOC_153/a_8_24# OR2X1_LOC_68/B 0.02fF
C53380 AND2X1_LOC_817/a_8_24# OR2X1_LOC_68/B 0.01fF
C53774 OR2X1_LOC_235/B OR2X1_LOC_68/B 0.13fF
C53893 OR2X1_LOC_276/B OR2X1_LOC_68/B 0.07fF
C54056 OR2X1_LOC_68/B AND2X1_LOC_226/a_8_24# 0.02fF
C54140 AND2X1_LOC_70/Y OR2X1_LOC_68/B 0.03fF
C55824 AND2X1_LOC_44/Y OR2X1_LOC_68/B 10.49fF
C56409 OR2X1_LOC_68/B VSS 0.66fF
C1079 OR2X1_LOC_671/Y OR2X1_LOC_56/A 0.11fF
C5326 OR2X1_LOC_671/Y OR2X1_LOC_96/B 0.19fF
C6527 OR2X1_LOC_671/Y OR2X1_LOC_600/A 0.68fF
C11495 OR2X1_LOC_671/Y OR2X1_LOC_95/Y 0.02fF
C13246 OR2X1_LOC_671/Y OR2X1_LOC_47/Y 0.07fF
C16321 OR2X1_LOC_159/a_8_216# OR2X1_LOC_671/Y 0.02fF
C21522 OR2X1_LOC_671/Y OR2X1_LOC_14/a_8_216# 0.01fF
C21787 OR2X1_LOC_671/Y OR2X1_LOC_28/a_8_216# -0.04fF
C23319 OR2X1_LOC_671/Y OR2X1_LOC_827/a_8_216# 0.02fF
C35791 OR2X1_LOC_671/Y OR2X1_LOC_9/a_8_216# 0.01fF
C36725 OR2X1_LOC_671/Y OR2X1_LOC_85/A 0.09fF
C44899 OR2X1_LOC_671/Y OR2X1_LOC_94/a_8_216# 0.04fF
C45385 OR2X1_LOC_671/Y OR2X1_LOC_827/Y 0.01fF
C45899 OR2X1_LOC_671/Y OR2X1_LOC_54/a_8_216# 0.02fF
C48055 OR2X1_LOC_671/Y OR2X1_LOC_42/a_8_216# 0.15fF
C52142 OR2X1_LOC_104/a_8_216# OR2X1_LOC_671/Y 0.39fF
C52227 OR2X1_LOC_671/Y OR2X1_LOC_6/A 0.19fF
C53393 OR2X1_LOC_671/Y OR2X1_LOC_158/A 0.11fF
C57840 OR2X1_LOC_671/Y VSS 0.63fF
C5664 AND2X1_LOC_619/B AND2X1_LOC_619/a_8_24# 0.19fF
C25362 VDD AND2X1_LOC_619/B 0.24fF
C28799 OR2X1_LOC_847/A AND2X1_LOC_619/B 0.01fF
C45232 AND2X1_LOC_619/B AND2X1_LOC_36/Y 0.10fF
C56525 AND2X1_LOC_619/B VSS -0.09fF
C516 OR2X1_LOC_95/Y OR2X1_LOC_85/A 0.15fF
C1479 OR2X1_LOC_85/A OR2X1_LOC_71/A 0.85fF
C1639 OR2X1_LOC_85/A OR2X1_LOC_59/Y 2.47fF
C1774 OR2X1_LOC_70/Y OR2X1_LOC_85/A 0.35fF
C2285 OR2X1_LOC_47/Y OR2X1_LOC_85/A 1.67fF
C2669 OR2X1_LOC_85/A OR2X1_LOC_8/a_8_216# 0.40fF
C3035 OR2X1_LOC_246/Y OR2X1_LOC_85/A 0.40fF
C3306 OR2X1_LOC_85/A OR2X1_LOC_16/A 0.06fF
C3929 OR2X1_LOC_277/a_8_216# OR2X1_LOC_85/A 0.08fF
C5352 OR2X1_LOC_40/Y OR2X1_LOC_85/A 1.52fF
C5519 OR2X1_LOC_7/A OR2X1_LOC_85/A 0.08fF
C6626 OR2X1_LOC_589/A OR2X1_LOC_85/A 0.02fF
C7703 OR2X1_LOC_3/Y OR2X1_LOC_85/A 0.05fF
C8006 OR2X1_LOC_671/a_8_216# OR2X1_LOC_85/A 0.01fF
C9029 OR2X1_LOC_64/Y OR2X1_LOC_85/A 0.11fF
C9438 AND2X1_LOC_101/B OR2X1_LOC_85/A 0.21fF
C11150 OR2X1_LOC_412/a_8_216# OR2X1_LOC_85/A 0.05fF
C12300 OR2X1_LOC_517/A OR2X1_LOC_85/A 0.29fF
C12524 OR2X1_LOC_85/A OR2X1_LOC_150/a_8_216# 0.05fF
C13359 OR2X1_LOC_234/a_8_216# OR2X1_LOC_85/A 0.01fF
C14464 OR2X1_LOC_85/A OR2X1_LOC_278/Y 0.02fF
C16159 OR2X1_LOC_36/Y OR2X1_LOC_85/A 0.07fF
C16286 OR2X1_LOC_85/a_8_216# OR2X1_LOC_85/A 0.01fF
C16450 OR2X1_LOC_604/A OR2X1_LOC_85/A 0.11fF
C16578 OR2X1_LOC_80/Y OR2X1_LOC_85/A 0.02fF
C17100 OR2X1_LOC_255/a_8_216# OR2X1_LOC_85/A 0.02fF
C18035 OR2X1_LOC_85/A OR2X1_LOC_150/a_36_216# 0.03fF
C18210 OR2X1_LOC_90/a_8_216# OR2X1_LOC_85/A 0.02fF
C19189 OR2X1_LOC_73/a_8_216# OR2X1_LOC_85/A 0.08fF
C20364 OR2X1_LOC_85/A OR2X1_LOC_234/Y 0.01fF
C20509 OR2X1_LOC_278/A OR2X1_LOC_85/A 0.10fF
C21680 OR2X1_LOC_256/Y OR2X1_LOC_85/A 0.05fF
C22591 OR2X1_LOC_18/Y OR2X1_LOC_85/A 0.37fF
C23624 OR2X1_LOC_85/A OR2X1_LOC_437/A 0.01fF
C23781 OR2X1_LOC_90/a_36_216# OR2X1_LOC_85/A 0.01fF
C23880 OR2X1_LOC_85/A OR2X1_LOC_753/A 0.05fF
C24422 OR2X1_LOC_85/A OR2X1_LOC_88/Y 0.02fF
C24714 OR2X1_LOC_85/A OR2X1_LOC_52/B 0.15fF
C24717 OR2X1_LOC_672/Y OR2X1_LOC_85/A 0.12fF
C25170 OR2X1_LOC_22/Y OR2X1_LOC_85/A 0.30fF
C25499 OR2X1_LOC_85/A OR2X1_LOC_39/A 0.07fF
C26250 OR2X1_LOC_51/Y OR2X1_LOC_85/A 0.10fF
C27341 OR2X1_LOC_86/A OR2X1_LOC_85/A 0.71fF
C29220 OR2X1_LOC_91/A OR2X1_LOC_85/A 0.07fF
C29709 OR2X1_LOC_32/B OR2X1_LOC_85/A 0.05fF
C29769 OR2X1_LOC_233/a_8_216# OR2X1_LOC_85/A 0.01fF
C30192 OR2X1_LOC_74/A OR2X1_LOC_85/A 1.26fF
C30635 OR2X1_LOC_263/a_8_216# OR2X1_LOC_85/A 0.14fF
C33988 OR2X1_LOC_485/A OR2X1_LOC_85/A 0.70fF
C34050 OR2X1_LOC_85/A OR2X1_LOC_10/a_8_216# 0.03fF
C34310 OR2X1_LOC_256/a_8_216# OR2X1_LOC_85/A 0.05fF
C36872 OR2X1_LOC_85/A OR2X1_LOC_42/a_8_216# 0.06fF
C37379 OR2X1_LOC_245/a_8_216# OR2X1_LOC_85/A 0.08fF
C38924 VDD OR2X1_LOC_85/A 0.82fF
C39128 OR2X1_LOC_256/A OR2X1_LOC_85/A 0.34fF
C40222 OR2X1_LOC_427/A OR2X1_LOC_85/A 0.14fF
C41044 OR2X1_LOC_104/a_8_216# OR2X1_LOC_85/A 0.01fF
C41153 OR2X1_LOC_85/A OR2X1_LOC_6/A 0.09fF
C41604 OR2X1_LOC_85/A OR2X1_LOC_44/Y 0.21fF
C41864 OR2X1_LOC_45/B OR2X1_LOC_85/A 0.12fF
C41887 OR2X1_LOC_102/a_8_216# OR2X1_LOC_85/A 0.03fF
C42326 OR2X1_LOC_158/A OR2X1_LOC_85/A 0.36fF
C44776 OR2X1_LOC_85/A OR2X1_LOC_153/a_8_216# 0.08fF
C44970 OR2X1_LOC_744/A OR2X1_LOC_85/A 0.02fF
C45168 OR2X1_LOC_31/Y OR2X1_LOC_85/A 0.03fF
C45369 OR2X1_LOC_129/a_8_216# OR2X1_LOC_85/A 0.05fF
C46295 OR2X1_LOC_85/A OR2X1_LOC_56/A 0.34fF
C46390 AND2X1_LOC_87/a_8_24# OR2X1_LOC_85/A 0.01fF
C46900 OR2X1_LOC_291/Y OR2X1_LOC_85/A 0.06fF
C48279 OR2X1_LOC_71/Y OR2X1_LOC_85/A 0.07fF
C48661 OR2X1_LOC_246/A OR2X1_LOC_85/A 0.09fF
C49803 OR2X1_LOC_235/B OR2X1_LOC_85/A 0.01fF
C51514 OR2X1_LOC_65/B OR2X1_LOC_85/A 0.06fF
C51599 OR2X1_LOC_62/a_8_216# OR2X1_LOC_85/A 0.01fF
C51854 OR2X1_LOC_600/A OR2X1_LOC_85/A 0.66fF
C51927 OR2X1_LOC_85/A OR2X1_LOC_619/Y 0.10fF
C51948 OR2X1_LOC_88/A OR2X1_LOC_85/A 0.05fF
C52895 OR2X1_LOC_813/A OR2X1_LOC_85/A 0.47fF
C53088 OR2X1_LOC_133/a_8_216# OR2X1_LOC_85/A 0.05fF
C54216 OR2X1_LOC_85/A OR2X1_LOC_13/B 0.04fF
C54722 OR2X1_LOC_85/A OR2X1_LOC_428/A 0.07fF
C55794 OR2X1_LOC_26/Y OR2X1_LOC_85/A 0.13fF
C56231 OR2X1_LOC_246/a_8_216# OR2X1_LOC_85/A 0.01fF
C56927 OR2X1_LOC_85/A VSS 0.98fF
C242 OR2X1_LOC_427/A OR2X1_LOC_382/A 0.17fF
C1160 OR2X1_LOC_6/A OR2X1_LOC_382/A 0.10fF
C2343 OR2X1_LOC_158/A OR2X1_LOC_382/A 0.05fF
C2908 OR2X1_LOC_748/A OR2X1_LOC_382/A 0.57fF
C6127 OR2X1_LOC_56/A OR2X1_LOC_382/A 0.10fF
C11699 OR2X1_LOC_600/A OR2X1_LOC_382/A 0.13fF
C15617 OR2X1_LOC_89/A OR2X1_LOC_382/A 0.26fF
C17709 OR2X1_LOC_820/B OR2X1_LOC_382/A 0.02fF
C23764 OR2X1_LOC_3/Y OR2X1_LOC_382/A 0.17fF
C32412 OR2X1_LOC_604/A OR2X1_LOC_382/A 0.06fF
C35789 OR2X1_LOC_12/Y OR2X1_LOC_382/A 0.54fF
C43953 OR2X1_LOC_382/A OR2X1_LOC_382/a_8_216# 0.39fF
C47017 OR2X1_LOC_381/a_8_216# OR2X1_LOC_382/A 0.01fF
C48455 AND2X1_LOC_847/Y OR2X1_LOC_382/A 0.02fF
C55079 VDD OR2X1_LOC_382/A -0.00fF
C56652 OR2X1_LOC_382/A VSS 0.31fF
C879 AND2X1_LOC_8/Y OR2X1_LOC_87/B 0.11fF
C914 AND2X1_LOC_85/a_8_24# AND2X1_LOC_8/Y 0.01fF
C1405 AND2X1_LOC_8/Y OR2X1_LOC_532/B 0.07fF
C3361 VDD AND2X1_LOC_8/Y 0.62fF
C6322 OR2X1_LOC_160/A AND2X1_LOC_8/Y 0.63fF
C6352 AND2X1_LOC_8/Y AND2X1_LOC_29/a_36_24# 0.01fF
C6383 AND2X1_LOC_86/B AND2X1_LOC_8/Y 0.04fF
C6614 AND2X1_LOC_8/Y OR2X1_LOC_266/A 0.03fF
C6874 AND2X1_LOC_8/Y AND2X1_LOC_46/a_8_24# 0.10fF
C7655 OR2X1_LOC_185/A AND2X1_LOC_8/Y 0.11fF
C10072 AND2X1_LOC_91/B AND2X1_LOC_8/Y 0.28fF
C10144 AND2X1_LOC_86/a_36_24# AND2X1_LOC_8/Y 0.01fF
C12022 AND2X1_LOC_8/Y AND2X1_LOC_47/Y 0.07fF
C12779 AND2X1_LOC_95/Y AND2X1_LOC_8/Y 0.04fF
C13083 AND2X1_LOC_22/Y AND2X1_LOC_8/Y 0.06fF
C14025 OR2X1_LOC_235/B AND2X1_LOC_8/Y 0.16fF
C15994 AND2X1_LOC_8/Y AND2X1_LOC_44/Y 0.29fF
C16928 AND2X1_LOC_8/Y AND2X1_LOC_18/Y 0.04fF
C17137 AND2X1_LOC_8/Y AND2X1_LOC_672/a_8_24# 0.01fF
C17853 AND2X1_LOC_8/Y OR2X1_LOC_130/A 0.02fF
C21790 AND2X1_LOC_8/Y AND2X1_LOC_102/a_8_24# 0.01fF
C21919 AND2X1_LOC_8/Y OR2X1_LOC_71/A 0.13fF
C22138 AND2X1_LOC_749/a_8_24# AND2X1_LOC_8/Y 0.11fF
C23241 AND2X1_LOC_8/Y AND2X1_LOC_36/Y 0.24fF
C23527 AND2X1_LOC_8/Y AND2X1_LOC_46/a_36_24# 0.01fF
C27069 AND2X1_LOC_8/Y OR2X1_LOC_161/B 0.71fF
C28138 AND2X1_LOC_133/a_8_24# AND2X1_LOC_8/Y 0.05fF
C28175 AND2X1_LOC_8/Y OR2X1_LOC_673/A 0.75fF
C28607 AND2X1_LOC_8/Y OR2X1_LOC_398/a_8_216# 0.02fF
C28866 AND2X1_LOC_8/Y AND2X1_LOC_104/a_8_24# 0.09fF
C29570 AND2X1_LOC_8/Y AND2X1_LOC_7/B 8.23fF
C34645 AND2X1_LOC_90/a_8_24# AND2X1_LOC_8/Y 0.01fF
C36776 AND2X1_LOC_8/Y OR2X1_LOC_66/A 0.08fF
C38099 AND2X1_LOC_40/Y AND2X1_LOC_8/Y 0.06fF
C38159 AND2X1_LOC_8/Y OR2X1_LOC_87/Y 0.08fF
C39556 AND2X1_LOC_519/a_8_24# AND2X1_LOC_8/Y 0.01fF
C39616 AND2X1_LOC_8/Y OR2X1_LOC_398/Y 0.01fF
C41073 AND2X1_LOC_8/Y OR2X1_LOC_78/A 0.18fF
C42890 AND2X1_LOC_59/Y AND2X1_LOC_8/Y 1.81fF
C44232 AND2X1_LOC_8/Y OR2X1_LOC_753/A 0.70fF
C45163 OR2X1_LOC_520/A AND2X1_LOC_8/Y 0.01fF
C46392 OR2X1_LOC_377/A AND2X1_LOC_8/Y 0.10fF
C46782 AND2X1_LOC_8/Y OR2X1_LOC_78/B 0.20fF
C46855 AND2X1_LOC_8/Y OR2X1_LOC_375/A 0.45fF
C47173 AND2X1_LOC_8/Y OR2X1_LOC_549/A 0.07fF
C48057 AND2X1_LOC_8/Y AND2X1_LOC_65/A 0.01fF
C48712 AND2X1_LOC_8/Y AND2X1_LOC_8/a_8_24# 0.01fF
C48937 AND2X1_LOC_19/Y AND2X1_LOC_8/Y 0.03fF
C49281 AND2X1_LOC_8/Y AND2X1_LOC_277/a_8_24# 0.01fF
C50359 AND2X1_LOC_8/Y AND2X1_LOC_4/a_8_24# 0.01fF
C51547 AND2X1_LOC_8/Y AND2X1_LOC_29/a_8_24# 0.05fF
C52392 AND2X1_LOC_63/a_8_24# AND2X1_LOC_8/Y 0.04fF
C54430 OR2X1_LOC_634/A AND2X1_LOC_8/Y 0.02fF
C54751 AND2X1_LOC_8/Y OR2X1_LOC_633/A 0.42fF
C55139 AND2X1_LOC_64/Y AND2X1_LOC_8/Y 0.09fF
C55233 AND2X1_LOC_86/a_8_24# AND2X1_LOC_8/Y 0.04fF
C55714 OR2X1_LOC_756/B AND2X1_LOC_8/Y 0.01fF
C57328 AND2X1_LOC_8/Y VSS 0.59fF
C446 OR2X1_LOC_299/a_8_216# OR2X1_LOC_6/A 0.01fF
C483 OR2X1_LOC_611/a_36_216# OR2X1_LOC_6/A 0.03fF
C866 OR2X1_LOC_6/A OR2X1_LOC_44/Y 1.81fF
C966 OR2X1_LOC_80/a_36_216# OR2X1_LOC_6/A 0.03fF
C1137 OR2X1_LOC_45/B OR2X1_LOC_6/A 0.09fF
C1596 OR2X1_LOC_158/A OR2X1_LOC_6/A 1.94fF
C3124 OR2X1_LOC_111/Y OR2X1_LOC_6/A 0.16fF
C4167 OR2X1_LOC_744/A OR2X1_LOC_6/A 0.33fF
C4333 OR2X1_LOC_31/Y OR2X1_LOC_6/A 0.83fF
C4751 AND2X1_LOC_270/a_8_24# OR2X1_LOC_6/A 0.01fF
C5388 OR2X1_LOC_56/A OR2X1_LOC_6/A 0.77fF
C6429 AND2X1_LOC_68/a_8_24# OR2X1_LOC_6/A 0.01fF
C6760 OR2X1_LOC_519/Y OR2X1_LOC_6/A 0.01fF
C7286 OR2X1_LOC_481/A OR2X1_LOC_6/A 0.04fF
C7516 OR2X1_LOC_6/A OR2X1_LOC_15/a_8_216# 0.14fF
C7641 AND2X1_LOC_95/Y OR2X1_LOC_6/A 0.04fF
C7743 OR2X1_LOC_246/A OR2X1_LOC_6/A 0.01fF
C7755 OR2X1_LOC_225/a_8_216# OR2X1_LOC_6/A 0.18fF
C8908 OR2X1_LOC_235/B OR2X1_LOC_6/A 1.01fF
C9278 OR2X1_LOC_6/A OR2X1_LOC_57/a_8_216# 0.07fF
C9834 OR2X1_LOC_96/B OR2X1_LOC_6/A 0.01fF
C10684 OR2X1_LOC_271/Y OR2X1_LOC_6/A 0.01fF
C10949 OR2X1_LOC_600/A OR2X1_LOC_6/A 5.32fF
C11043 OR2X1_LOC_619/Y OR2X1_LOC_6/A 0.03fF
C11520 OR2X1_LOC_6/A AND2X1_LOC_818/a_8_24# 0.01fF
C12349 OR2X1_LOC_6/A OR2X1_LOC_69/A 0.01fF
C13424 OR2X1_LOC_6/A OR2X1_LOC_13/B 0.03fF
C13924 OR2X1_LOC_6/A OR2X1_LOC_428/A 0.23fF
C14926 OR2X1_LOC_26/Y OR2X1_LOC_6/A 0.14fF
C14944 OR2X1_LOC_89/A OR2X1_LOC_6/A 0.78fF
C15720 OR2X1_LOC_824/Y OR2X1_LOC_6/A 0.16fF
C15808 OR2X1_LOC_95/Y OR2X1_LOC_6/A 0.06fF
C15809 OR2X1_LOC_368/A OR2X1_LOC_6/A 0.01fF
C16751 OR2X1_LOC_6/A OR2X1_LOC_71/A 0.04fF
C16946 OR2X1_LOC_6/A OR2X1_LOC_59/Y 0.07fF
C17031 OR2X1_LOC_6/A OR2X1_LOC_820/B 0.03fF
C17063 OR2X1_LOC_70/Y OR2X1_LOC_6/A 0.03fF
C17532 OR2X1_LOC_47/Y OR2X1_LOC_6/A 0.11fF
C18426 OR2X1_LOC_6/A OR2X1_LOC_29/a_8_216# 0.03fF
C18571 OR2X1_LOC_6/A OR2X1_LOC_16/A 5.46fF
C19228 OR2X1_LOC_268/a_8_216# OR2X1_LOC_6/A 0.06fF
C19463 OR2X1_LOC_93/Y OR2X1_LOC_6/A 0.01fF
C20462 OR2X1_LOC_93/a_8_216# OR2X1_LOC_6/A 0.01fF
C20745 OR2X1_LOC_159/a_8_216# OR2X1_LOC_6/A 0.02fF
C20748 OR2X1_LOC_40/Y OR2X1_LOC_6/A 0.13fF
C20917 OR2X1_LOC_7/A OR2X1_LOC_6/A 0.26fF
C21597 OR2X1_LOC_6/A AND2X1_LOC_415/a_8_24# 0.01fF
C22037 OR2X1_LOC_589/A OR2X1_LOC_6/A 0.02fF
C22153 AND2X1_LOC_398/a_8_24# OR2X1_LOC_6/A 0.06fF
C22660 OR2X1_LOC_299/Y OR2X1_LOC_6/A 0.01fF
C23071 OR2X1_LOC_3/Y OR2X1_LOC_6/A 0.36fF
C23376 OR2X1_LOC_329/B OR2X1_LOC_6/A 0.23fF
C23984 OR2X1_LOC_6/A OR2X1_LOC_29/a_36_216# 0.02fF
C24297 OR2X1_LOC_690/A OR2X1_LOC_6/A 0.02fF
C24336 OR2X1_LOC_64/Y OR2X1_LOC_6/A 0.02fF
C24788 OR2X1_LOC_55/a_8_216# OR2X1_LOC_6/A 0.01fF
C25808 OR2X1_LOC_6/A OR2X1_LOC_14/a_8_216# 0.41fF
C26067 OR2X1_LOC_6/A OR2X1_LOC_28/a_8_216# -0.00fF
C26232 OR2X1_LOC_159/a_36_216# OR2X1_LOC_6/A 0.03fF
C27635 OR2X1_LOC_827/a_8_216# OR2X1_LOC_6/A 0.01fF
C28896 OR2X1_LOC_6/A OR2X1_LOC_49/a_8_216# 0.01fF
C29698 OR2X1_LOC_6/A OR2X1_LOC_278/Y 0.02fF
C30395 OR2X1_LOC_136/a_8_216# OR2X1_LOC_6/A 0.01fF
C31421 OR2X1_LOC_36/Y OR2X1_LOC_6/A 1.29fF
C31728 OR2X1_LOC_604/A OR2X1_LOC_6/A 0.05fF
C31817 OR2X1_LOC_80/Y OR2X1_LOC_6/A 0.02fF
C33798 OR2X1_LOC_6/A OR2X1_LOC_310/a_8_216# 0.02fF
C35060 OR2X1_LOC_6/A OR2X1_LOC_12/Y 0.46fF
C37661 OR2X1_LOC_57/Y OR2X1_LOC_6/A 0.01fF
C37701 OR2X1_LOC_18/Y OR2X1_LOC_6/A 1.02fF
C38561 AND2X1_LOC_398/a_36_24# OR2X1_LOC_6/A 0.02fF
C38787 OR2X1_LOC_6/A OR2X1_LOC_437/A 0.07fF
C39061 OR2X1_LOC_753/A OR2X1_LOC_6/A 0.10fF
C39294 OR2X1_LOC_6/A OR2X1_LOC_310/a_36_216# 0.03fF
C39898 OR2X1_LOC_6/A OR2X1_LOC_52/B 1.10fF
C40107 OR2X1_LOC_9/a_8_216# OR2X1_LOC_6/A 0.01fF
C40168 AND2X1_LOC_514/a_8_24# OR2X1_LOC_6/A 0.01fF
C40353 OR2X1_LOC_22/Y OR2X1_LOC_6/A 0.03fF
C40698 OR2X1_LOC_6/A OR2X1_LOC_39/A 0.04fF
C41399 OR2X1_LOC_136/Y OR2X1_LOC_6/A 0.54fF
C41493 OR2X1_LOC_51/Y OR2X1_LOC_6/A 1.45fF
C43194 OR2X1_LOC_6/A OR2X1_LOC_382/a_8_216# 0.19fF
C43418 OR2X1_LOC_416/A OR2X1_LOC_6/A 0.43fF
C44550 OR2X1_LOC_91/A OR2X1_LOC_6/A 0.15fF
C45132 OR2X1_LOC_5/a_8_216# OR2X1_LOC_6/A 0.01fF
C45539 OR2X1_LOC_74/A OR2X1_LOC_6/A 0.10fF
C46825 OR2X1_LOC_71/a_8_216# OR2X1_LOC_6/A 0.06fF
C49430 OR2X1_LOC_94/a_8_216# OR2X1_LOC_6/A 0.01fF
C49481 OR2X1_LOC_485/A OR2X1_LOC_6/A 0.04fF
C49901 OR2X1_LOC_827/Y OR2X1_LOC_6/A 0.01fF
C50300 OR2X1_LOC_271/B OR2X1_LOC_6/A 0.19fF
C50391 OR2X1_LOC_54/a_8_216# OR2X1_LOC_6/A 0.01fF
C51176 OR2X1_LOC_611/a_8_216# OR2X1_LOC_6/A 0.10fF
C51622 OR2X1_LOC_80/a_8_216# OR2X1_LOC_6/A 0.09fF
C51923 OR2X1_LOC_519/a_8_216# OR2X1_LOC_6/A 0.01fF
C52393 OR2X1_LOC_42/a_8_216# OR2X1_LOC_6/A 0.01fF
C54365 VDD OR2X1_LOC_6/A 1.48fF
C54679 OR2X1_LOC_6/A AND2X1_LOC_269/a_8_24# 0.01fF
C54899 OR2X1_LOC_6/a_8_216# OR2X1_LOC_6/A 0.01fF
C55274 OR2X1_LOC_382/Y OR2X1_LOC_6/A 0.01fF
C55743 OR2X1_LOC_427/A OR2X1_LOC_6/A 0.16fF
C55786 OR2X1_LOC_271/a_8_216# OR2X1_LOC_6/A 0.01fF
C56702 OR2X1_LOC_6/A VSS 1.62fF
C8323 VDD OR2X1_LOC_414/Y 0.19fF
C16418 OR2X1_LOC_83/A OR2X1_LOC_414/Y 0.73fF
C56524 OR2X1_LOC_414/Y VSS 0.16fF
C324 OR2X1_LOC_377/A AND2X1_LOC_41/A 0.84fF
C1466 OR2X1_LOC_377/A OR2X1_LOC_71/A 0.03fF
C1850 OR2X1_LOC_377/A AND2X1_LOC_31/Y 0.07fF
C2170 OR2X1_LOC_377/A OR2X1_LOC_240/A 7.16fF
C2796 OR2X1_LOC_377/A AND2X1_LOC_36/Y 8.97fF
C3545 OR2X1_LOC_377/A AND2X1_LOC_827/a_8_24# 0.03fF
C5056 OR2X1_LOC_377/A OR2X1_LOC_269/B 1.58fF
C6595 OR2X1_LOC_377/A OR2X1_LOC_161/B 0.03fF
C7679 OR2X1_LOC_377/A OR2X1_LOC_3/Y 0.28fF
C7741 OR2X1_LOC_377/A AND2X1_LOC_53/Y 0.01fF
C7762 OR2X1_LOC_377/A OR2X1_LOC_673/A 0.03fF
C8592 OR2X1_LOC_377/A AND2X1_LOC_3/Y 0.48fF
C9202 OR2X1_LOC_377/A AND2X1_LOC_7/B 0.12fF
C9402 OR2X1_LOC_377/A OR2X1_LOC_836/A 0.02fF
C10680 OR2X1_LOC_287/B OR2X1_LOC_377/A 0.04fF
C10933 OR2X1_LOC_160/B OR2X1_LOC_377/A 0.02fF
C11469 OR2X1_LOC_377/A AND2X1_LOC_233/a_8_24# 0.02fF
C13023 OR2X1_LOC_377/A OR2X1_LOC_415/Y 0.03fF
C13381 OR2X1_LOC_377/A OR2X1_LOC_378/A 0.32fF
C14062 AND2X1_LOC_80/a_8_24# OR2X1_LOC_377/A 0.03fF
C14150 OR2X1_LOC_377/A AND2X1_LOC_15/a_8_24# 0.05fF
C14592 OR2X1_LOC_377/A OR2X1_LOC_838/B 0.01fF
C16132 OR2X1_LOC_377/A OR2X1_LOC_36/Y 5.35fF
C16437 OR2X1_LOC_377/A OR2X1_LOC_66/A 0.22fF
C16840 OR2X1_LOC_691/a_8_216# OR2X1_LOC_377/A 0.02fF
C16914 OR2X1_LOC_377/A AND2X1_LOC_94/Y 0.46fF
C17760 AND2X1_LOC_40/Y OR2X1_LOC_377/A 0.23fF
C19475 OR2X1_LOC_377/A AND2X1_LOC_377/Y 0.03fF
C20079 OR2X1_LOC_377/A OR2X1_LOC_606/Y 0.15fF
C20754 OR2X1_LOC_377/A OR2X1_LOC_78/A 0.33fF
C21761 AND2X1_LOC_387/B OR2X1_LOC_377/A 0.02fF
C22147 AND2X1_LOC_12/Y OR2X1_LOC_377/A 0.12fF
C22581 AND2X1_LOC_59/Y OR2X1_LOC_377/A 0.11fF
C25079 OR2X1_LOC_377/A AND2X1_LOC_49/a_8_24# 0.04fF
C25381 OR2X1_LOC_377/A AND2X1_LOC_387/a_8_24# 0.03fF
C25479 OR2X1_LOC_377/A OR2X1_LOC_39/A 0.03fF
C26243 OR2X1_LOC_377/A OR2X1_LOC_78/B 4.27fF
C26306 OR2X1_LOC_377/A OR2X1_LOC_375/A 0.49fF
C26600 OR2X1_LOC_377/A OR2X1_LOC_549/A 0.90fF
C27409 OR2X1_LOC_377/A OR2X1_LOC_20/A 0.14fF
C27680 OR2X1_LOC_377/A AND2X1_LOC_23/a_8_24# 0.05fF
C28702 OR2X1_LOC_377/A AND2X1_LOC_277/a_8_24# 0.02fF
C30472 OR2X1_LOC_377/A OR2X1_LOC_459/A 0.14fF
C30877 OR2X1_LOC_377/A OR2X1_LOC_389/A 0.03fF
C31475 OR2X1_LOC_377/A AND2X1_LOC_5/a_8_24# 0.20fF
C32043 OR2X1_LOC_377/A OR2X1_LOC_691/Y 0.02fF
C32276 OR2X1_LOC_377/A OR2X1_LOC_750/a_8_216# 0.03fF
C32537 OR2X1_LOC_377/A OR2X1_LOC_461/B 0.01fF
C33067 OR2X1_LOC_154/A OR2X1_LOC_377/A 0.22fF
C33211 OR2X1_LOC_377/A AND2X1_LOC_6/a_8_24# 0.01fF
C33842 OR2X1_LOC_377/A OR2X1_LOC_461/a_8_216# 0.06fF
C33871 OR2X1_LOC_377/A OR2X1_LOC_634/A 0.05fF
C34184 OR2X1_LOC_377/A OR2X1_LOC_633/A 7.06fF
C34231 OR2X1_LOC_377/A AND2X1_LOC_110/a_8_24# 0.12fF
C34516 OR2X1_LOC_377/A OR2X1_LOC_376/Y 0.06fF
C34560 AND2X1_LOC_64/Y OR2X1_LOC_377/A 0.15fF
C34608 OR2X1_LOC_377/A AND2X1_LOC_82/Y 0.27fF
C35119 OR2X1_LOC_756/B OR2X1_LOC_377/A 0.66fF
C35747 OR2X1_LOC_377/A AND2X1_LOC_699/a_8_24# 0.09fF
C36315 OR2X1_LOC_377/A OR2X1_LOC_596/A 0.02fF
C36448 OR2X1_LOC_377/A OR2X1_LOC_87/B 0.04fF
C36937 OR2X1_LOC_377/A OR2X1_LOC_532/B 0.54fF
C38121 OR2X1_LOC_185/Y OR2X1_LOC_377/A 0.02fF
C38133 OR2X1_LOC_377/A AND2X1_LOC_412/a_8_24# 0.02fF
C38899 VDD OR2X1_LOC_377/A 2.16fF
C38963 OR2X1_LOC_377/A OR2X1_LOC_689/A 0.03fF
C41739 OR2X1_LOC_377/A OR2X1_LOC_750/Y 0.82fF
C41979 OR2X1_LOC_160/A OR2X1_LOC_377/A 0.07fF
C42040 OR2X1_LOC_377/A AND2X1_LOC_86/B 0.07fF
C42426 OR2X1_LOC_377/A OR2X1_LOC_847/A 0.03fF
C42513 OR2X1_LOC_377/A AND2X1_LOC_46/a_8_24# 0.01fF
C43285 OR2X1_LOC_377/A OR2X1_LOC_185/A 0.07fF
C45720 AND2X1_LOC_91/B OR2X1_LOC_377/A 0.07fF
C46375 OR2X1_LOC_377/A AND2X1_LOC_56/B 0.18fF
C47314 OR2X1_LOC_377/A OR2X1_LOC_83/A 0.07fF
C47818 OR2X1_LOC_377/A AND2X1_LOC_47/Y 0.13fF
C48164 OR2X1_LOC_377/A AND2X1_LOC_82/a_8_24# 0.01fF
C48556 AND2X1_LOC_95/Y OR2X1_LOC_377/A 0.22fF
C48816 AND2X1_LOC_22/Y OR2X1_LOC_377/A 0.07fF
C49777 OR2X1_LOC_235/B OR2X1_LOC_377/A 0.07fF
C50113 OR2X1_LOC_709/A OR2X1_LOC_377/A 0.25fF
C50159 AND2X1_LOC_70/Y OR2X1_LOC_377/A 0.23fF
C51780 OR2X1_LOC_377/A AND2X1_LOC_44/Y 0.11fF
C52660 OR2X1_LOC_377/A AND2X1_LOC_18/Y 0.12fF
C52949 OR2X1_LOC_377/A OR2X1_LOC_377/a_8_216# 0.06fF
C53644 OR2X1_LOC_377/A OR2X1_LOC_130/A 0.01fF
C55729 OR2X1_LOC_377/A OR2X1_LOC_161/A 0.03fF
C55820 OR2X1_LOC_377/A AND2X1_LOC_51/Y 0.57fF
C57776 OR2X1_LOC_377/A VSS -5.63fF
C4585 VDD OR2X1_LOC_529/Y 0.57fF
C5931 OR2X1_LOC_529/Y OR2X1_LOC_427/A 0.04fF
C7267 OR2X1_LOC_529/Y OR2X1_LOC_44/Y 0.03fF
C7533 OR2X1_LOC_45/B OR2X1_LOC_529/Y 0.02fF
C8013 OR2X1_LOC_158/A OR2X1_LOC_529/Y 0.03fF
C10618 OR2X1_LOC_529/Y OR2X1_LOC_744/A 0.04fF
C10787 OR2X1_LOC_529/Y OR2X1_LOC_31/Y 0.01fF
C18816 OR2X1_LOC_529/Y OR2X1_LOC_530/Y 0.21fF
C20298 OR2X1_LOC_529/Y OR2X1_LOC_428/A 0.02fF
C21372 OR2X1_LOC_529/Y OR2X1_LOC_26/Y 0.04fF
C21388 OR2X1_LOC_529/Y OR2X1_LOC_89/A 0.03fF
C22038 OR2X1_LOC_529/Y OR2X1_LOC_816/A 0.05fF
C22294 OR2X1_LOC_529/Y OR2X1_LOC_95/Y 0.03fF
C23403 OR2X1_LOC_529/Y OR2X1_LOC_59/Y 0.04fF
C23995 OR2X1_LOC_529/Y OR2X1_LOC_47/Y 0.06fF
C27271 OR2X1_LOC_529/Y OR2X1_LOC_7/A 0.06fF
C30646 OR2X1_LOC_529/Y OR2X1_LOC_64/Y 0.03fF
C37763 OR2X1_LOC_529/Y OR2X1_LOC_36/Y 0.04fF
C37870 OR2X1_LOC_529/Y OR2X1_LOC_419/Y 0.03fF
C38055 OR2X1_LOC_604/A OR2X1_LOC_529/Y 0.03fF
C44206 OR2X1_LOC_529/Y OR2X1_LOC_18/Y 0.02fF
C45273 OR2X1_LOC_529/Y OR2X1_LOC_437/A 0.07fF
C46940 OR2X1_LOC_529/Y OR2X1_LOC_22/Y 0.03fF
C47336 OR2X1_LOC_529/Y OR2X1_LOC_39/A 0.05fF
C48124 OR2X1_LOC_529/Y OR2X1_LOC_51/Y 0.54fF
C55847 OR2X1_LOC_529/Y OR2X1_LOC_485/A 0.04fF
C57623 OR2X1_LOC_529/Y VSS -0.01fF
C970 OR2X1_LOC_22/A OR2X1_LOC_21/a_8_216# -0.00fF
C8962 VDD OR2X1_LOC_22/A 0.27fF
C11584 OR2X1_LOC_22/A OR2X1_LOC_44/Y 0.06fF
C12318 OR2X1_LOC_158/A OR2X1_LOC_22/A 0.03fF
C13859 OR2X1_LOC_22/A OR2X1_LOC_588/a_8_216# 0.01fF
C14909 OR2X1_LOC_744/A OR2X1_LOC_22/A 0.01fF
C15059 OR2X1_LOC_31/Y OR2X1_LOC_22/A 0.05fF
C23198 OR2X1_LOC_51/B OR2X1_LOC_22/A 0.03fF
C24026 OR2X1_LOC_22/A OR2X1_LOC_409/a_8_216# 0.01fF
C25603 OR2X1_LOC_26/Y OR2X1_LOC_22/A 0.04fF
C26032 OR2X1_LOC_22/A OR2X1_LOC_17/Y 0.16fF
C28223 OR2X1_LOC_47/Y OR2X1_LOC_22/A 0.63fF
C28626 OR2X1_LOC_3/B OR2X1_LOC_22/A 0.44fF
C32299 OR2X1_LOC_22/A OR2X1_LOC_22/a_8_216# 0.08fF
C34883 OR2X1_LOC_11/Y OR2X1_LOC_22/A 1.53fF
C34971 OR2X1_LOC_64/a_8_216# OR2X1_LOC_22/A 0.03fF
C36054 OR2X1_LOC_22/A OR2X1_LOC_25/Y 0.11fF
C37247 OR2X1_LOC_22/A OR2X1_LOC_36/a_8_216# 0.18fF
C38291 OR2X1_LOC_22/A OR2X1_LOC_408/a_8_216# 0.41fF
C40442 OR2X1_LOC_64/a_36_216# OR2X1_LOC_22/A 0.02fF
C42102 OR2X1_LOC_36/Y OR2X1_LOC_22/A 0.03fF
C45233 OR2X1_LOC_409/Y OR2X1_LOC_22/A 0.01fF
C47326 OR2X1_LOC_22/A OR2X1_LOC_26/a_8_216# 0.06fF
C49596 OR2X1_LOC_22/A OR2X1_LOC_408/a_36_216# -0.00fF
C51237 OR2X1_LOC_22/Y OR2X1_LOC_22/A 0.02fF
C52369 OR2X1_LOC_51/Y OR2X1_LOC_22/A 0.09fF
C52822 OR2X1_LOC_22/A OR2X1_LOC_26/a_36_216# 0.02fF
C53299 OR2X1_LOC_22/A OR2X1_LOC_588/Y 0.02fF
C56926 OR2X1_LOC_22/A VSS -0.02fF
C123 AND2X1_LOC_91/B OR2X1_LOC_596/A 0.56fF
C495 OR2X1_LOC_596/A OR2X1_LOC_446/B 0.04fF
C707 AND2X1_LOC_56/B OR2X1_LOC_596/A 0.02fF
C1902 OR2X1_LOC_596/A OR2X1_LOC_596/a_8_216# 0.13fF
C2137 AND2X1_LOC_47/Y OR2X1_LOC_596/A 0.04fF
C2453 OR2X1_LOC_506/A OR2X1_LOC_596/A 0.29fF
C3179 AND2X1_LOC_22/Y OR2X1_LOC_596/A 0.01fF
C3748 AND2X1_LOC_329/a_8_24# OR2X1_LOC_596/A 0.06fF
C4407 OR2X1_LOC_709/A OR2X1_LOC_596/A 0.08fF
C6069 OR2X1_LOC_596/A AND2X1_LOC_44/Y 0.20fF
C6089 OR2X1_LOC_596/A OR2X1_LOC_514/a_8_216# 0.01fF
C6984 AND2X1_LOC_18/Y OR2X1_LOC_596/A 0.03fF
C7099 OR2X1_LOC_596/Y OR2X1_LOC_596/A 0.04fF
C10082 OR2X1_LOC_161/A OR2X1_LOC_596/A 0.03fF
C10178 AND2X1_LOC_51/Y OR2X1_LOC_596/A 0.14fF
C10872 AND2X1_LOC_41/A OR2X1_LOC_596/A 0.11fF
C11410 AND2X1_LOC_136/a_8_24# OR2X1_LOC_596/A 0.01fF
C12417 AND2X1_LOC_31/Y OR2X1_LOC_596/A 0.03fF
C13350 OR2X1_LOC_596/A AND2X1_LOC_36/Y 0.08fF
C15603 OR2X1_LOC_596/A OR2X1_LOC_269/B 0.05fF
C16673 OR2X1_LOC_596/A OR2X1_LOC_777/B 0.72fF
C17173 OR2X1_LOC_596/A OR2X1_LOC_161/B 0.06fF
C18272 AND2X1_LOC_53/Y OR2X1_LOC_596/A 0.07fF
C19054 AND2X1_LOC_3/Y OR2X1_LOC_596/A 0.04fF
C19735 AND2X1_LOC_7/B OR2X1_LOC_596/A 0.07fF
C20333 AND2X1_LOC_329/a_36_24# OR2X1_LOC_596/A 0.01fF
C20967 OR2X1_LOC_596/A OR2X1_LOC_513/Y 0.02fF
C21526 OR2X1_LOC_160/B OR2X1_LOC_596/A 0.03fF
C22354 OR2X1_LOC_151/A OR2X1_LOC_596/A 0.13fF
C26019 OR2X1_LOC_596/A OR2X1_LOC_515/a_8_216# 0.01fF
C26967 OR2X1_LOC_596/A OR2X1_LOC_66/A 0.03fF
C28289 AND2X1_LOC_40/Y OR2X1_LOC_596/A 0.05fF
C30437 OR2X1_LOC_687/Y OR2X1_LOC_596/A 0.03fF
C31212 OR2X1_LOC_78/A OR2X1_LOC_596/A 2.54fF
C32144 AND2X1_LOC_387/B OR2X1_LOC_596/A 4.20fF
C32509 AND2X1_LOC_12/Y OR2X1_LOC_596/A 1.29fF
C34172 AND2X1_LOC_421/a_8_24# OR2X1_LOC_596/A 0.11fF
C36652 OR2X1_LOC_78/B OR2X1_LOC_596/A 0.03fF
C36716 OR2X1_LOC_375/A OR2X1_LOC_596/A 0.07fF
C36969 OR2X1_LOC_596/A OR2X1_LOC_515/Y 0.13fF
C38407 OR2X1_LOC_405/A OR2X1_LOC_596/A 0.04fF
C40009 OR2X1_LOC_596/A OR2X1_LOC_138/A 0.01fF
C41002 OR2X1_LOC_87/A OR2X1_LOC_596/A 0.03fF
C43632 OR2X1_LOC_154/A OR2X1_LOC_596/A 0.07fF
C45205 AND2X1_LOC_64/Y OR2X1_LOC_596/A 0.03fF
C47718 OR2X1_LOC_532/B OR2X1_LOC_596/A 0.03fF
C48868 OR2X1_LOC_185/Y OR2X1_LOC_596/A 0.03fF
C49646 VDD OR2X1_LOC_596/A 0.41fF
C51604 OR2X1_LOC_596/A AND2X1_LOC_419/a_8_24# 0.01fF
C52646 OR2X1_LOC_160/A OR2X1_LOC_596/A 0.02fF
C56595 OR2X1_LOC_596/A VSS 0.25fF
C4664 AND2X1_LOC_11/Y AND2X1_LOC_18/a_8_24# 0.11fF
C6238 AND2X1_LOC_2/a_8_24# AND2X1_LOC_11/Y 0.22fF
C7977 VDD AND2X1_LOC_11/Y 0.90fF
C10696 AND2X1_LOC_1/Y AND2X1_LOC_11/Y 0.07fF
C12171 AND2X1_LOC_40/a_8_24# AND2X1_LOC_11/Y 0.01fF
C13367 AND2X1_LOC_11/Y AND2X1_LOC_429/a_8_24# 0.03fF
C14389 AND2X1_LOC_12/a_8_24# AND2X1_LOC_11/Y 0.01fF
C15290 AND2X1_LOC_21/Y AND2X1_LOC_11/Y 0.17fF
C16647 AND2X1_LOC_11/Y AND2X1_LOC_47/Y 0.08fF
C17632 AND2X1_LOC_22/Y AND2X1_LOC_11/Y 0.01fF
C19010 AND2X1_LOC_70/Y AND2X1_LOC_11/Y 0.77fF
C20674 AND2X1_LOC_11/Y AND2X1_LOC_44/Y 0.03fF
C24398 AND2X1_LOC_11/Y AND2X1_LOC_429/a_36_24# 0.01fF
C24654 AND2X1_LOC_11/Y AND2X1_LOC_25/Y 1.05fF
C24722 AND2X1_LOC_11/Y AND2X1_LOC_51/Y 1.18fF
C26899 AND2X1_LOC_11/Y AND2X1_LOC_31/Y 0.05fF
C27791 AND2X1_LOC_11/Y AND2X1_LOC_36/Y 0.07fF
C30023 AND2X1_LOC_2/Y AND2X1_LOC_11/Y 0.44fF
C33542 AND2X1_LOC_11/Y AND2X1_LOC_3/Y 0.29fF
C34156 AND2X1_LOC_11/Y AND2X1_LOC_7/B 0.03fF
C41010 AND2X1_LOC_70/a_8_24# AND2X1_LOC_11/Y 0.01fF
C41927 AND2X1_LOC_50/Y AND2X1_LOC_11/Y 0.08fF
C42817 AND2X1_LOC_40/Y AND2X1_LOC_11/Y 0.01fF
C47235 AND2X1_LOC_22/a_8_24# AND2X1_LOC_11/Y 0.01fF
C47255 AND2X1_LOC_12/Y AND2X1_LOC_11/Y 0.01fF
C47933 AND2X1_LOC_11/Y AND2X1_LOC_762/a_8_24# 0.11fF
C50232 AND2X1_LOC_47/a_8_24# AND2X1_LOC_11/Y 0.11fF
C55745 AND2X1_LOC_11/Y OR2X1_LOC_87/A 0.02fF
C57187 AND2X1_LOC_11/Y VSS -0.50fF
C916 AND2X1_LOC_387/B OR2X1_LOC_269/B 0.02fF
C2490 AND2X1_LOC_387/B OR2X1_LOC_161/B 0.07fF
C3561 AND2X1_LOC_387/B AND2X1_LOC_53/Y 0.07fF
C4304 AND2X1_LOC_387/B AND2X1_LOC_3/Y 0.04fF
C6708 OR2X1_LOC_160/B AND2X1_LOC_387/B 0.12fF
C13636 AND2X1_LOC_40/Y AND2X1_LOC_387/B 0.27fF
C15864 AND2X1_LOC_387/B OR2X1_LOC_644/A 0.03fF
C17868 AND2X1_LOC_12/Y AND2X1_LOC_387/B 0.03fF
C21230 AND2X1_LOC_387/B AND2X1_LOC_387/a_8_24# 0.04fF
C22200 AND2X1_LOC_387/B OR2X1_LOC_375/A 0.03fF
C26371 AND2X1_LOC_387/B OR2X1_LOC_87/A 0.03fF
C27913 AND2X1_LOC_387/B OR2X1_LOC_691/Y 0.03fF
C30439 AND2X1_LOC_599/a_8_24# AND2X1_LOC_387/B 0.03fF
C32787 AND2X1_LOC_387/B OR2X1_LOC_532/B 0.11fF
C34718 VDD AND2X1_LOC_387/B 0.18fF
C37488 AND2X1_LOC_387/B OR2X1_LOC_750/Y 0.10fF
C42068 AND2X1_LOC_387/B AND2X1_LOC_56/B 0.03fF
C43439 AND2X1_LOC_387/B AND2X1_LOC_47/Y 0.01fF
C44482 AND2X1_LOC_22/Y AND2X1_LOC_387/B 0.09fF
C45866 AND2X1_LOC_70/Y AND2X1_LOC_387/B 0.03fF
C47622 AND2X1_LOC_387/B AND2X1_LOC_44/Y 2.30fF
C52344 AND2X1_LOC_387/B AND2X1_LOC_41/A 0.11fF
C54701 AND2X1_LOC_387/B AND2X1_LOC_36/Y 0.06fF
C57780 AND2X1_LOC_387/B VSS 0.20fF
C5527 OR2X1_LOC_635/A AND2X1_LOC_425/Y 0.01fF
C5573 OR2X1_LOC_687/B AND2X1_LOC_425/Y 0.01fF
C7654 AND2X1_LOC_2/Y AND2X1_LOC_425/Y 0.10fF
C9349 AND2X1_LOC_425/Y OR2X1_LOC_161/B 0.01fF
C9953 AND2X1_LOC_425/Y OR2X1_LOC_451/A 0.01fF
C14366 AND2X1_LOC_425/Y AND2X1_LOC_581/a_8_24# 0.01fF
C15829 OR2X1_LOC_687/a_8_216# AND2X1_LOC_425/Y 0.01fF
C22698 OR2X1_LOC_687/Y AND2X1_LOC_425/Y 0.01fF
C24757 AND2X1_LOC_12/Y AND2X1_LOC_425/Y 0.48fF
C25493 OR2X1_LOC_686/a_8_216# AND2X1_LOC_425/Y 0.01fF
C28950 AND2X1_LOC_425/Y OR2X1_LOC_375/A 0.01fF
C34004 AND2X1_LOC_425/Y AND2X1_LOC_426/a_8_24# 0.05fF
C35693 AND2X1_LOC_157/a_8_24# AND2X1_LOC_425/Y 0.19fF
C36447 OR2X1_LOC_687/A AND2X1_LOC_425/Y 0.01fF
C36586 AND2X1_LOC_425/Y AND2X1_LOC_694/a_8_24# 0.05fF
C41576 VDD AND2X1_LOC_425/Y 0.46fF
C45051 OR2X1_LOC_450/B AND2X1_LOC_425/Y 0.01fF
C47875 AND2X1_LOC_425/Y OR2X1_LOC_707/B 0.01fF
C50746 AND2X1_LOC_582/a_8_24# AND2X1_LOC_425/Y 0.01fF
C50791 OR2X1_LOC_685/a_8_216# AND2X1_LOC_425/Y 0.01fF
C52589 AND2X1_LOC_425/Y AND2X1_LOC_430/B 1.50fF
C55008 AND2X1_LOC_425/Y AND2X1_LOC_430/a_8_24# 0.01fF
C57152 AND2X1_LOC_425/Y VSS 0.39fF
C105 OR2X1_LOC_47/Y OR2X1_LOC_753/A 0.05fF
C408 OR2X1_LOC_625/Y OR2X1_LOC_753/A 0.17fF
C870 OR2X1_LOC_246/Y OR2X1_LOC_753/A 0.08fF
C1154 OR2X1_LOC_753/A OR2X1_LOC_16/A 0.59fF
C3345 OR2X1_LOC_40/Y OR2X1_LOC_753/A 0.03fF
C3465 OR2X1_LOC_246/a_36_216# OR2X1_LOC_753/A 0.01fF
C3482 OR2X1_LOC_7/A OR2X1_LOC_753/A 0.10fF
C3719 OR2X1_LOC_753/A OR2X1_LOC_753/a_8_216# 0.12fF
C5542 OR2X1_LOC_3/Y OR2X1_LOC_753/A 0.13fF
C5628 AND2X1_LOC_462/B OR2X1_LOC_753/A 0.10fF
C6824 OR2X1_LOC_690/A OR2X1_LOC_753/A 0.03fF
C6875 OR2X1_LOC_64/Y OR2X1_LOC_753/A 0.02fF
C10440 OR2X1_LOC_753/A OR2X1_LOC_150/a_8_216# 0.04fF
C11195 OR2X1_LOC_234/a_8_216# OR2X1_LOC_753/A 0.03fF
C12353 OR2X1_LOC_753/A OR2X1_LOC_38/a_8_216# 0.03fF
C14109 OR2X1_LOC_36/Y OR2X1_LOC_753/A 0.06fF
C14394 OR2X1_LOC_604/A OR2X1_LOC_753/A 0.10fF
C15013 OR2X1_LOC_255/a_8_216# OR2X1_LOC_753/A 0.01fF
C15685 AND2X1_LOC_375/a_8_24# OR2X1_LOC_753/A 0.23fF
C17695 OR2X1_LOC_753/A OR2X1_LOC_12/Y 0.04fF
C17940 AND2X1_LOC_671/a_8_24# OR2X1_LOC_753/A 0.04fF
C18250 OR2X1_LOC_753/A OR2X1_LOC_234/Y 0.05fF
C19541 OR2X1_LOC_256/Y OR2X1_LOC_753/A 0.01fF
C20433 OR2X1_LOC_18/Y OR2X1_LOC_753/A 0.06fF
C21521 OR2X1_LOC_753/A OR2X1_LOC_437/A 0.19fF
C22657 OR2X1_LOC_753/A OR2X1_LOC_52/B 0.72fF
C23108 OR2X1_LOC_22/Y OR2X1_LOC_753/A 0.03fF
C23454 OR2X1_LOC_753/A OR2X1_LOC_39/A 0.03fF
C24206 OR2X1_LOC_51/Y OR2X1_LOC_753/A 0.07fF
C26027 OR2X1_LOC_255/a_36_216# OR2X1_LOC_753/A 0.01fF
C26372 AND2X1_LOC_294/a_8_24# OR2X1_LOC_753/A 0.01fF
C27161 OR2X1_LOC_91/A OR2X1_LOC_753/A 0.07fF
C27616 OR2X1_LOC_32/B OR2X1_LOC_753/A 0.10fF
C27670 OR2X1_LOC_233/a_8_216# OR2X1_LOC_753/A 0.03fF
C28105 OR2X1_LOC_74/A OR2X1_LOC_753/A 0.03fF
C31858 OR2X1_LOC_485/A OR2X1_LOC_753/A 0.11fF
C31931 OR2X1_LOC_10/a_8_216# OR2X1_LOC_753/A 0.01fF
C32201 OR2X1_LOC_256/a_8_216# OR2X1_LOC_753/A -0.03fF
C33151 OR2X1_LOC_233/a_36_216# OR2X1_LOC_753/A 0.01fF
C35556 AND2X1_LOC_691/a_8_24# OR2X1_LOC_753/A 0.03fF
C36771 VDD OR2X1_LOC_753/A 6.11fF
C36973 OR2X1_LOC_256/A OR2X1_LOC_753/A 0.09fF
C37441 OR2X1_LOC_10/a_36_216# OR2X1_LOC_753/A 0.17fF
C38117 OR2X1_LOC_427/A OR2X1_LOC_753/A 0.14fF
C39488 OR2X1_LOC_753/A OR2X1_LOC_44/Y 0.12fF
C39747 OR2X1_LOC_102/a_8_216# OR2X1_LOC_753/A 0.01fF
C40135 OR2X1_LOC_158/A OR2X1_LOC_753/A 0.14fF
C42103 OR2X1_LOC_293/a_8_216# OR2X1_LOC_753/A 0.01fF
C42840 OR2X1_LOC_744/A OR2X1_LOC_753/A 0.21fF
C43012 OR2X1_LOC_31/Y OR2X1_LOC_753/A 0.29fF
C44114 OR2X1_LOC_753/A OR2X1_LOC_56/A 0.17fF
C45097 OR2X1_LOC_83/A OR2X1_LOC_753/A 0.05fF
C45372 OR2X1_LOC_102/a_36_216# OR2X1_LOC_753/A 0.01fF
C46009 OR2X1_LOC_481/A OR2X1_LOC_753/A 0.01fF
C46226 OR2X1_LOC_753/A OR2X1_LOC_15/a_8_216# 0.03fF
C46489 OR2X1_LOC_415/a_8_216# OR2X1_LOC_753/A 0.35fF
C46496 OR2X1_LOC_246/A OR2X1_LOC_753/A 0.14fF
C46779 AND2X1_LOC_691/a_36_24# OR2X1_LOC_753/A 0.01fF
C47684 OR2X1_LOC_235/B OR2X1_LOC_753/A 0.17fF
C49537 OR2X1_LOC_62/a_8_216# OR2X1_LOC_753/A 0.03fF
C49782 OR2X1_LOC_600/A OR2X1_LOC_753/A 0.14fF
C49864 OR2X1_LOC_619/Y OR2X1_LOC_753/A 0.07fF
C52130 OR2X1_LOC_753/A OR2X1_LOC_13/B 0.10fF
C52651 OR2X1_LOC_753/A OR2X1_LOC_428/A 0.03fF
C53702 OR2X1_LOC_26/Y OR2X1_LOC_753/A 0.07fF
C53719 OR2X1_LOC_89/A OR2X1_LOC_753/A 0.11fF
C54069 OR2X1_LOC_246/a_8_216# OR2X1_LOC_753/A 0.04fF
C54307 OR2X1_LOC_753/A OR2X1_LOC_816/A 0.51fF
C54580 OR2X1_LOC_95/Y OR2X1_LOC_753/A 0.07fF
C55516 OR2X1_LOC_753/A OR2X1_LOC_71/A 0.16fF
C55691 OR2X1_LOC_753/A OR2X1_LOC_59/Y 0.07fF
C56784 OR2X1_LOC_753/A VSS 0.74fF
C2218 OR2X1_LOC_11/Y OR2X1_LOC_762/a_8_216# 0.02fF
C2278 OR2X1_LOC_409/Y OR2X1_LOC_11/Y 0.01fF
C2875 OR2X1_LOC_11/Y OR2X1_LOC_12/Y 0.18fF
C3405 OR2X1_LOC_11/Y OR2X1_LOC_59/a_8_216# 0.01fF
C4158 OR2X1_LOC_11/Y OR2X1_LOC_26/a_8_216# 0.01fF
C5446 OR2X1_LOC_18/Y OR2X1_LOC_11/Y 0.17fF
C8193 OR2X1_LOC_22/Y OR2X1_LOC_11/Y 0.78fF
C9300 OR2X1_LOC_51/Y OR2X1_LOC_11/Y 0.07fF
C10251 OR2X1_LOC_11/Y OR2X1_LOC_588/Y 0.01fF
C18113 OR2X1_LOC_11/Y OR2X1_LOC_18/a_8_216# 0.02fF
C22053 VDD OR2X1_LOC_11/Y 0.35fF
C23690 OR2X1_LOC_11/Y OR2X1_LOC_18/a_36_216# 0.03fF
C24691 OR2X1_LOC_11/Y OR2X1_LOC_44/Y 0.79fF
C25372 OR2X1_LOC_158/A OR2X1_LOC_11/Y 0.03fF
C26923 OR2X1_LOC_11/Y OR2X1_LOC_588/a_8_216# 0.01fF
C27948 OR2X1_LOC_744/A OR2X1_LOC_11/Y 0.11fF
C28139 OR2X1_LOC_31/Y OR2X1_LOC_11/Y 0.20fF
C29872 OR2X1_LOC_11/Y OR2X1_LOC_11/a_8_216# -0.00fF
C31259 OR2X1_LOC_11/Y OR2X1_LOC_585/a_8_216# 0.01fF
C31514 OR2X1_LOC_11/Y OR2X1_LOC_409/B 0.04fF
C31739 OR2X1_LOC_11/Y OR2X1_LOC_12/a_8_216# 0.18fF
C34423 OR2X1_LOC_11/Y OR2X1_LOC_429/a_8_216# 0.39fF
C36155 OR2X1_LOC_11/Y OR2X1_LOC_51/B 0.03fF
C36964 OR2X1_LOC_11/Y OR2X1_LOC_409/a_8_216# 0.01fF
C38594 OR2X1_LOC_26/Y OR2X1_LOC_11/Y 0.03fF
C39072 OR2X1_LOC_11/Y OR2X1_LOC_17/Y 0.13fF
C40618 OR2X1_LOC_11/Y OR2X1_LOC_59/Y 0.01fF
C41248 OR2X1_LOC_47/Y OR2X1_LOC_11/Y 0.23fF
C41713 OR2X1_LOC_11/Y OR2X1_LOC_3/B 0.33fF
C44486 OR2X1_LOC_40/Y OR2X1_LOC_11/Y 0.04fF
C46278 OR2X1_LOC_11/Y OR2X1_LOC_585/Y 0.01fF
C46876 OR2X1_LOC_3/Y OR2X1_LOC_11/Y 0.34fF
C48241 OR2X1_LOC_64/Y OR2X1_LOC_11/Y 0.04fF
C48285 OR2X1_LOC_11/Y OR2X1_LOC_64/a_8_216# 0.01fF
C49342 OR2X1_LOC_11/Y OR2X1_LOC_25/Y 0.03fF
C53660 OR2X1_LOC_11/Y OR2X1_LOC_95/a_8_216# 0.08fF
C55344 OR2X1_LOC_36/Y OR2X1_LOC_11/Y 0.03fF
C57016 OR2X1_LOC_11/Y VSS 0.81fF
C5261 OR2X1_LOC_51/B OR2X1_LOC_587/a_8_216# 0.01fF
C12920 OR2X1_LOC_51/B OR2X1_LOC_44/Y 0.01fF
C13663 OR2X1_LOC_158/A OR2X1_LOC_51/B 0.06fF
C16260 OR2X1_LOC_1/a_8_216# OR2X1_LOC_51/B 0.03fF
C16329 OR2X1_LOC_31/Y OR2X1_LOC_51/B 0.01fF
C18384 AND2X1_LOC_51/a_8_24# OR2X1_LOC_51/B 0.01fF
C18525 OR2X1_LOC_51/a_8_216# OR2X1_LOC_51/B 0.07fF
C27350 OR2X1_LOC_51/B OR2X1_LOC_17/Y 0.38fF
C29946 OR2X1_LOC_51/B OR2X1_LOC_3/B 0.21fF
C32818 OR2X1_LOC_51/B OR2X1_LOC_44/a_8_216# 0.04fF
C35405 OR2X1_LOC_51/B OR2X1_LOC_31/a_8_216# 0.02fF
C37361 OR2X1_LOC_51/B OR2X1_LOC_25/Y 0.03fF
C38589 OR2X1_LOC_51/B OR2X1_LOC_36/a_8_216# 0.01fF
C43444 OR2X1_LOC_36/Y OR2X1_LOC_51/B 0.09fF
C49212 OR2X1_LOC_50/a_8_216# OR2X1_LOC_51/B 0.39fF
C53723 OR2X1_LOC_51/Y OR2X1_LOC_51/B 0.07fF
C56930 OR2X1_LOC_51/B VSS 0.39fF
C1186 AND2X1_LOC_12/Y AND2X1_LOC_2/Y 1.05fF
C5365 AND2X1_LOC_2/Y OR2X1_LOC_375/A 0.01fF
C12238 AND2X1_LOC_2/Y AND2X1_LOC_157/a_8_24# 0.01fF
C16400 AND2X1_LOC_2/Y AND2X1_LOC_2/a_8_24# 0.01fF
C18085 AND2X1_LOC_2/Y VDD 0.52fF
C18310 AND2X1_LOC_2/Y AND2X1_LOC_25/a_8_24# 0.18fF
C20844 AND2X1_LOC_2/Y AND2X1_LOC_1/Y 0.11fF
C22371 AND2X1_LOC_2/Y AND2X1_LOC_40/a_8_24# 0.06fF
C23535 AND2X1_LOC_2/Y AND2X1_LOC_429/a_8_24# 0.01fF
C24513 AND2X1_LOC_2/Y AND2X1_LOC_12/a_8_24# 0.20fF
C25354 AND2X1_LOC_2/Y AND2X1_LOC_3/a_8_24# 0.01fF
C28973 AND2X1_LOC_2/Y AND2X1_LOC_430/B 0.02fF
C29107 AND2X1_LOC_2/Y AND2X1_LOC_70/Y 0.01fF
C30744 AND2X1_LOC_2/Y AND2X1_LOC_44/Y 0.03fF
C31807 AND2X1_LOC_2/Y AND2X1_LOC_11/a_8_24# 0.01fF
C33294 AND2X1_LOC_2/Y AND2X1_LOC_40/a_36_24# 0.01fF
C34687 AND2X1_LOC_2/Y AND2X1_LOC_25/Y 0.20fF
C34758 AND2X1_LOC_2/Y AND2X1_LOC_51/Y 0.01fF
C36952 AND2X1_LOC_2/Y AND2X1_LOC_31/Y 0.04fF
C43713 AND2X1_LOC_2/Y AND2X1_LOC_3/Y 0.01fF
C45022 AND2X1_LOC_2/Y AND2X1_LOC_425/a_8_24# 0.01fF
C52204 AND2X1_LOC_50/Y AND2X1_LOC_2/Y 0.03fF
C57842 AND2X1_LOC_2/Y VSS 0.18fF
C3119 AND2X1_LOC_21/a_36_24# AND2X1_LOC_21/Y 0.01fF
C3381 VDD AND2X1_LOC_21/Y 0.53fF
C6006 AND2X1_LOC_1/Y AND2X1_LOC_21/Y 0.90fF
C8512 AND2X1_LOC_588/a_8_24# AND2X1_LOC_21/Y 0.01fF
C12032 AND2X1_LOC_21/Y AND2X1_LOC_47/Y 0.07fF
C14029 OR2X1_LOC_638/B AND2X1_LOC_21/Y 0.01fF
C16013 AND2X1_LOC_21/Y AND2X1_LOC_44/Y 0.02fF
C16212 AND2X1_LOC_21/Y AND2X1_LOC_36/a_8_24# 0.01fF
C20046 AND2X1_LOC_21/Y AND2X1_LOC_25/Y 0.96fF
C20102 AND2X1_LOC_21/Y AND2X1_LOC_51/Y 0.04fF
C22348 AND2X1_LOC_21/Y AND2X1_LOC_31/Y 0.19fF
C22711 AND2X1_LOC_31/a_8_24# AND2X1_LOC_21/Y 0.17fF
C23258 AND2X1_LOC_21/Y AND2X1_LOC_36/Y 0.69fF
C25547 AND2X1_LOC_21/Y AND2X1_LOC_26/a_8_24# 0.03fF
C37277 AND2X1_LOC_50/Y AND2X1_LOC_21/Y 0.54fF
C40746 AND2X1_LOC_64/a_8_24# AND2X1_LOC_21/Y 0.13fF
C43151 AND2X1_LOC_21/Y AND2X1_LOC_762/a_8_24# 0.02fF
C49707 AND2X1_LOC_588/B AND2X1_LOC_21/Y 0.04fF
C55154 AND2X1_LOC_64/Y AND2X1_LOC_21/Y 0.01fF
C57244 AND2X1_LOC_21/Y VSS 0.28fF
C573 AND2X1_LOC_53/Y AND2X1_LOC_56/a_8_24# 0.21fF
C1812 OR2X1_LOC_687/Y AND2X1_LOC_53/Y 0.46fF
C3940 AND2X1_LOC_12/Y AND2X1_LOC_53/Y 0.09fF
C4318 AND2X1_LOC_59/Y AND2X1_LOC_53/Y 0.07fF
C6080 AND2X1_LOC_53/Y OR2X1_LOC_197/A 0.03fF
C6943 AND2X1_LOC_53/Y AND2X1_LOC_692/a_8_24# 0.02fF
C8130 AND2X1_LOC_53/Y OR2X1_LOC_78/B 0.07fF
C8208 AND2X1_LOC_53/Y OR2X1_LOC_375/A 0.44fF
C12454 AND2X1_LOC_53/Y OR2X1_LOC_87/A 0.02fF
C12501 AND2X1_LOC_53/Y OR2X1_LOC_706/B 0.04fF
C16480 AND2X1_LOC_64/Y AND2X1_LOC_53/Y 0.17fF
C18005 AND2X1_LOC_53/Y AND2X1_LOC_692/a_36_24# 0.01fF
C20111 OR2X1_LOC_185/Y AND2X1_LOC_53/Y 0.01fF
C20879 VDD AND2X1_LOC_53/Y 0.21fF
C25136 AND2X1_LOC_53/Y AND2X1_LOC_693/a_8_24# 0.02fF
C26404 AND2X1_LOC_753/a_8_24# AND2X1_LOC_53/Y 0.02fF
C29467 AND2X1_LOC_53/Y AND2X1_LOC_47/Y 0.07fF
C30216 AND2X1_LOC_95/Y AND2X1_LOC_53/Y 0.12fF
C30500 AND2X1_LOC_22/Y AND2X1_LOC_53/Y 0.21fF
C30600 AND2X1_LOC_53/Y OR2X1_LOC_706/A 0.09fF
C31643 AND2X1_LOC_53/Y OR2X1_LOC_779/B 0.34fF
C31822 AND2X1_LOC_70/Y AND2X1_LOC_53/Y 0.07fF
C33490 AND2X1_LOC_53/Y AND2X1_LOC_44/Y 0.02fF
C34335 AND2X1_LOC_53/Y AND2X1_LOC_18/Y 0.08fF
C37106 AND2X1_LOC_53/Y OR2X1_LOC_513/a_8_216# 0.01fF
C37383 OR2X1_LOC_790/B AND2X1_LOC_53/Y 0.05fF
C37388 AND2X1_LOC_53/Y OR2X1_LOC_161/A 0.08fF
C37447 AND2X1_LOC_53/Y AND2X1_LOC_51/Y 0.04fF
C38186 AND2X1_LOC_41/A AND2X1_LOC_53/Y 0.02fF
C39684 AND2X1_LOC_53/Y AND2X1_LOC_31/Y 0.10fF
C40580 AND2X1_LOC_53/Y AND2X1_LOC_36/Y 0.02fF
C41643 AND2X1_LOC_53/Y AND2X1_LOC_693/a_36_24# -0.01fF
C42974 AND2X1_LOC_753/a_36_24# AND2X1_LOC_53/Y 0.01fF
C43004 AND2X1_LOC_53/Y OR2X1_LOC_269/B 0.50fF
C43812 AND2X1_LOC_304/a_8_24# AND2X1_LOC_53/Y 0.09fF
C46517 AND2X1_LOC_53/Y AND2X1_LOC_3/Y 0.07fF
C47242 AND2X1_LOC_53/Y AND2X1_LOC_7/B 0.07fF
C48997 OR2X1_LOC_160/B AND2X1_LOC_53/Y 0.52fF
C54469 AND2X1_LOC_53/Y OR2X1_LOC_66/A 0.07fF
C55830 AND2X1_LOC_40/Y AND2X1_LOC_53/Y 0.08fF
C57340 AND2X1_LOC_53/Y VSS 0.86fF
C9816 AND2X1_LOC_31/Y AND2X1_LOC_409/B 0.03fF
C15707 AND2X1_LOC_409/B AND2X1_LOC_409/a_8_24# 0.03fF
C24856 AND2X1_LOC_50/Y AND2X1_LOC_409/B 0.24fF
C28255 OR2X1_LOC_828/B AND2X1_LOC_409/B 0.10fF
C30337 AND2X1_LOC_752/a_8_24# AND2X1_LOC_409/B 0.04fF
C34147 OR2X1_LOC_375/A AND2X1_LOC_409/B 0.03fF
C38837 OR2X1_LOC_21/a_8_216# AND2X1_LOC_409/B 0.47fF
C41323 AND2X1_LOC_752/a_36_24# AND2X1_LOC_409/B 0.01fF
C46992 VDD AND2X1_LOC_409/B 0.08fF
C56329 AND2X1_LOC_409/B VSS 0.28fF
C3360 OR2X1_LOC_157/a_8_216# OR2X1_LOC_25/Y 0.02fF
C9417 OR2X1_LOC_22/Y OR2X1_LOC_25/Y 0.24fF
C10484 OR2X1_LOC_51/Y OR2X1_LOC_25/Y 0.07fF
C11432 OR2X1_LOC_588/Y OR2X1_LOC_25/Y 0.03fF
C22054 OR2X1_LOC_53/a_8_216# OR2X1_LOC_25/Y 0.01fF
C22129 OR2X1_LOC_47/a_8_216# OR2X1_LOC_25/Y 0.09fF
C23263 VDD OR2X1_LOC_25/Y 0.09fF
C25838 OR2X1_LOC_25/Y OR2X1_LOC_44/Y 0.03fF
C26554 OR2X1_LOC_158/A OR2X1_LOC_25/Y 0.89fF
C29131 OR2X1_LOC_744/A OR2X1_LOC_25/Y 0.26fF
C29330 OR2X1_LOC_31/Y OR2X1_LOC_25/Y 0.26fF
C31459 OR2X1_LOC_51/a_8_216# OR2X1_LOC_25/Y 0.03fF
C32718 OR2X1_LOC_409/B OR2X1_LOC_25/Y 0.03fF
C32954 OR2X1_LOC_425/a_8_216# OR2X1_LOC_25/Y 0.04fF
C40217 OR2X1_LOC_17/Y OR2X1_LOC_25/Y 0.07fF
C42528 OR2X1_LOC_47/Y OR2X1_LOC_25/Y 0.18fF
C42953 OR2X1_LOC_3/B OR2X1_LOC_25/Y 0.33fF
C46776 OR2X1_LOC_22/a_8_216# OR2X1_LOC_25/Y 0.02fF
C55622 OR2X1_LOC_40/a_8_216# OR2X1_LOC_25/Y 0.04fF
C56583 OR2X1_LOC_25/Y VSS 0.25fF
C14020 OR2X1_LOC_70/Y OR2X1_LOC_581/Y 0.28fF
C23447 OR2X1_LOC_70/a_8_216# OR2X1_LOC_581/Y 0.40fF
C51318 VDD OR2X1_LOC_581/Y -0.00fF
C52648 OR2X1_LOC_427/A OR2X1_LOC_581/Y 0.14fF
C56768 OR2X1_LOC_581/Y VSS 0.08fF
C10895 VDD OR2X1_LOC_762/Y 0.17fF
C13582 OR2X1_LOC_762/Y OR2X1_LOC_44/Y 0.04fF
C16854 OR2X1_LOC_744/A OR2X1_LOC_762/Y 0.26fF
C20482 OR2X1_LOC_409/B OR2X1_LOC_762/Y 0.20fF
C26550 OR2X1_LOC_762/Y OR2X1_LOC_428/A 0.06fF
C36857 OR2X1_LOC_64/Y OR2X1_LOC_762/Y 0.18fF
C47950 OR2X1_LOC_762/Y OR2X1_LOC_12/Y 0.04fF
C50608 OR2X1_LOC_18/Y OR2X1_LOC_762/Y 0.07fF
C56787 OR2X1_LOC_762/Y VSS 0.24fF
C2957 AND2X1_LOC_40/a_8_24# AND2X1_LOC_1/Y 0.01fF
C5057 AND2X1_LOC_1/Y AND2X1_LOC_12/a_8_24# 0.09fF
C5929 AND2X1_LOC_1/Y AND2X1_LOC_3/a_8_24# 0.09fF
C7379 AND2X1_LOC_1/Y AND2X1_LOC_47/Y 0.20fF
C9598 AND2X1_LOC_1/Y AND2X1_LOC_430/B 0.09fF
C11389 AND2X1_LOC_1/Y AND2X1_LOC_44/Y 0.04fF
C15353 AND2X1_LOC_1/Y AND2X1_LOC_25/Y 0.31fF
C15393 AND2X1_LOC_1/Y AND2X1_LOC_51/Y 0.01fF
C17601 AND2X1_LOC_1/Y AND2X1_LOC_31/Y 0.07fF
C17964 AND2X1_LOC_1/Y AND2X1_LOC_31/a_8_24# -0.00fF
C32685 AND2X1_LOC_50/Y AND2X1_LOC_1/Y 0.02fF
C37753 AND2X1_LOC_1/Y AND2X1_LOC_22/a_8_24# 0.10fF
C40747 AND2X1_LOC_1/Y AND2X1_LOC_47/a_8_24# 0.01fF
C57529 AND2X1_LOC_1/Y VSS 0.46fF
C1807 OR2X1_LOC_687/A AND2X1_LOC_430/B 0.01fF
C6883 VDD AND2X1_LOC_430/B 0.47fF
C14186 AND2X1_LOC_3/a_8_24# AND2X1_LOC_430/B 0.19fF
C15819 AND2X1_LOC_582/a_8_24# AND2X1_LOC_430/B 0.01fF
C15865 OR2X1_LOC_685/a_8_216# AND2X1_LOC_430/B 0.01fF
C20225 AND2X1_LOC_430/a_8_24# AND2X1_LOC_430/B 0.10fF
C26927 OR2X1_LOC_687/B AND2X1_LOC_430/B 0.01fF
C33723 AND2X1_LOC_425/a_8_24# AND2X1_LOC_430/B 0.01fF
C35618 AND2X1_LOC_430/B AND2X1_LOC_581/a_8_24# 0.01fF
C37072 OR2X1_LOC_687/a_8_216# AND2X1_LOC_430/B 0.01fF
C46088 AND2X1_LOC_12/Y AND2X1_LOC_430/B 0.01fF
C46922 OR2X1_LOC_686/a_8_216# AND2X1_LOC_430/B 0.01fF
C56375 AND2X1_LOC_430/B VSS -0.26fF
C379 OR2X1_LOC_51/Y OR2X1_LOC_17/Y 1.58fF
C8274 OR2X1_LOC_17/Y OR2X1_LOC_587/a_8_216# 0.01fF
C9285 OR2X1_LOC_17/Y OR2X1_LOC_18/a_8_216# 0.03fF
C13181 VDD OR2X1_LOC_17/Y 0.05fF
C16481 OR2X1_LOC_158/A OR2X1_LOC_17/Y 0.10fF
C19278 OR2X1_LOC_31/Y OR2X1_LOC_17/Y 0.06fF
C21040 OR2X1_LOC_11/a_8_216# OR2X1_LOC_17/Y 0.01fF
C23000 OR2X1_LOC_17/Y OR2X1_LOC_12/a_8_216# 0.01fF
C25635 OR2X1_LOC_429/a_8_216# OR2X1_LOC_17/Y 0.05fF
C28755 OR2X1_LOC_17/Y OR2X1_LOC_428/A 0.03fF
C32356 OR2X1_LOC_47/Y OR2X1_LOC_17/Y 0.01fF
C32817 OR2X1_LOC_3/B OR2X1_LOC_17/Y 0.02fF
C35562 OR2X1_LOC_40/Y OR2X1_LOC_17/Y 0.01fF
C35713 OR2X1_LOC_17/Y OR2X1_LOC_44/a_8_216# 0.08fF
C36515 OR2X1_LOC_22/a_8_216# OR2X1_LOC_17/Y 0.01fF
C37798 OR2X1_LOC_3/Y OR2X1_LOC_17/Y 0.03fF
C41487 OR2X1_LOC_17/Y OR2X1_LOC_36/a_8_216# 0.08fF
C45505 OR2X1_LOC_40/a_8_216# OR2X1_LOC_17/Y 0.01fF
C50172 OR2X1_LOC_17/Y OR2X1_LOC_12/Y 0.01fF
C51125 OR2X1_LOC_30/a_8_216# OR2X1_LOC_17/Y 0.40fF
C52081 OR2X1_LOC_50/a_8_216# OR2X1_LOC_17/Y 0.01fF
C54551 OR2X1_LOC_3/a_8_216# OR2X1_LOC_17/Y 0.02fF
C55437 OR2X1_LOC_22/Y OR2X1_LOC_17/Y 0.01fF
C56821 OR2X1_LOC_17/Y VSS 0.84fF
C1029 OR2X1_LOC_3/a_8_216# OR2X1_LOC_3/B 0.03fF
C1893 OR2X1_LOC_22/Y OR2X1_LOC_3/B 0.02fF
C3082 OR2X1_LOC_51/Y OR2X1_LOC_3/B 0.69fF
C10860 OR2X1_LOC_3/B OR2X1_LOC_587/a_8_216# 0.01fF
C14635 OR2X1_LOC_3/B OR2X1_LOC_47/a_8_216# 0.05fF
C18427 OR2X1_LOC_3/B OR2X1_LOC_44/Y 0.01fF
C19174 OR2X1_LOC_158/A OR2X1_LOC_3/B 0.07fF
C21939 OR2X1_LOC_31/Y OR2X1_LOC_3/B 0.07fF
C25569 OR2X1_LOC_3/B OR2X1_LOC_12/a_8_216# 0.01fF
C35019 OR2X1_LOC_47/Y OR2X1_LOC_3/B 0.77fF
C38187 OR2X1_LOC_40/Y OR2X1_LOC_3/B 0.01fF
C38301 OR2X1_LOC_3/B OR2X1_LOC_44/a_8_216# 0.02fF
C39173 OR2X1_LOC_3/B OR2X1_LOC_22/a_8_216# 0.04fF
C40429 OR2X1_LOC_3/Y OR2X1_LOC_3/B 0.04fF
C40925 OR2X1_LOC_3/B OR2X1_LOC_31/a_8_216# 0.06fF
C44203 OR2X1_LOC_3/B OR2X1_LOC_36/a_8_216# 0.40fF
C48286 OR2X1_LOC_40/a_8_216# OR2X1_LOC_3/B 0.02fF
C49114 OR2X1_LOC_36/Y OR2X1_LOC_3/B 0.01fF
C56929 OR2X1_LOC_3/B VSS 0.31fF
C12677 VDD AND2X1_LOC_25/Y 0.33fF
C16050 AND2X1_LOC_95/a_8_24# AND2X1_LOC_25/Y 0.01fF
C16879 AND2X1_LOC_40/a_8_24# AND2X1_LOC_25/Y 0.14fF
C21419 AND2X1_LOC_25/Y AND2X1_LOC_47/Y 0.06fF
C22159 AND2X1_LOC_95/Y AND2X1_LOC_25/Y 0.02fF
C23765 AND2X1_LOC_70/Y AND2X1_LOC_25/Y 0.11fF
C25358 AND2X1_LOC_25/Y AND2X1_LOC_44/Y 0.04fF
C27901 AND2X1_LOC_40/a_36_24# AND2X1_LOC_25/Y 0.01fF
C29361 AND2X1_LOC_25/Y AND2X1_LOC_51/Y 0.09fF
C31574 AND2X1_LOC_25/Y AND2X1_LOC_31/Y 0.06fF
C32429 AND2X1_LOC_25/Y AND2X1_LOC_36/Y 0.01fF
C34808 AND2X1_LOC_25/Y AND2X1_LOC_26/a_8_24# 0.13fF
C35611 AND2X1_LOC_59/a_8_24# AND2X1_LOC_25/Y 0.13fF
C46798 AND2X1_LOC_50/Y AND2X1_LOC_25/Y 1.21fF
C51917 AND2X1_LOC_22/a_8_24# AND2X1_LOC_25/Y 0.11fF
C57186 AND2X1_LOC_25/Y VSS 0.21fF
C7076 AND2X1_LOC_50/Y AND2X1_LOC_70/a_8_24# 0.24fF
C8861 AND2X1_LOC_50/Y AND2X1_LOC_40/Y 0.07fF
C11465 AND2X1_LOC_50/Y AND2X1_LOC_64/a_8_24# 0.04fF
C13537 AND2X1_LOC_50/Y AND2X1_LOC_752/a_8_24# 0.04fF
C13577 AND2X1_LOC_50/Y AND2X1_LOC_59/Y 0.01fF
C13817 AND2X1_LOC_50/Y AND2X1_LOC_408/a_8_24# 0.17fF
C13822 AND2X1_LOC_50/Y AND2X1_LOC_762/a_8_24# 0.01fF
C17364 AND2X1_LOC_50/Y OR2X1_LOC_375/A 0.04fF
C24580 AND2X1_LOC_50/Y AND2X1_LOC_752/a_36_24# 0.01fF
C28025 AND2X1_LOC_50/Y AND2X1_LOC_64/a_36_24# 0.01fF
C29628 AND2X1_LOC_50/Y AND2X1_LOC_53/a_8_24# 0.03fF
C29992 AND2X1_LOC_50/Y VDD 0.40fF
C33354 AND2X1_LOC_50/Y AND2X1_LOC_95/a_8_24# 0.11fF
C38009 AND2X1_LOC_50/Y AND2X1_LOC_51/a_8_24# 0.11fF
C38645 AND2X1_LOC_50/Y AND2X1_LOC_47/Y 1.11fF
C39372 AND2X1_LOC_50/Y AND2X1_LOC_95/Y 0.01fF
C39662 AND2X1_LOC_50/Y AND2X1_LOC_22/Y 0.02fF
C40971 AND2X1_LOC_50/Y AND2X1_LOC_70/Y 0.05fF
C42700 AND2X1_LOC_50/Y AND2X1_LOC_44/Y 0.03fF
C46298 AND2X1_LOC_50/Y AND2X1_LOC_53/a_36_24# 0.01fF
C46857 AND2X1_LOC_50/Y AND2X1_LOC_51/Y 0.84fF
C49109 AND2X1_LOC_50/Y AND2X1_LOC_31/Y 0.07fF
C50026 AND2X1_LOC_50/Y AND2X1_LOC_36/Y 0.03fF
C52326 AND2X1_LOC_50/Y AND2X1_LOC_26/a_8_24# 0.01fF
C53141 AND2X1_LOC_50/Y AND2X1_LOC_59/a_8_24# 0.01fF
C58118 AND2X1_LOC_50/Y VSS 0.34fF
C12616 AND2X1_LOC_588/B AND2X1_LOC_44/a_8_24# 0.19fF
C42181 AND2X1_LOC_588/B VDD 0.38fF
C57910 AND2X1_LOC_588/B VSS -0.04fF
C56128 AND2X1_LOC_59/Y OR2X1_LOC_274/Y 0.01fF
C33827 AND2X1_LOC_41/A OR2X1_LOC_274/Y 0.01fF
C36208 OR2X1_LOC_274/Y AND2X1_LOC_36/Y 0.03fF
C3792 OR2X1_LOC_274/Y OR2X1_LOC_375/A 0.01fF
C4078 OR2X1_LOC_274/Y OR2X1_LOC_549/A 0.07fF
C23818 AND2X1_LOC_56/B OR2X1_LOC_274/Y 0.18fF
C23218 AND2X1_LOC_91/B OR2X1_LOC_274/Y 0.05fF
C55546 OR2X1_LOC_121/Y OR2X1_LOC_274/Y 0.10fF
C2751 AND2X1_LOC_3/Y OR2X1_LOC_644/A 0.02fF
C12014 AND2X1_LOC_40/Y OR2X1_LOC_644/A 0.14fF
C16692 AND2X1_LOC_59/Y OR2X1_LOC_644/A 0.13fF
C16277 AND2X1_LOC_12/Y OR2X1_LOC_644/A 0.02fF
C26341 OR2X1_LOC_691/Y OR2X1_LOC_644/A 0.31fF
C53158 AND2X1_LOC_36/Y OR2X1_LOC_644/A 0.05fF
C45939 AND2X1_LOC_44/Y OR2X1_LOC_644/A 0.09fF
C11950 OR2X1_LOC_598/Y OR2X1_LOC_644/A 0.01fF
C34071 OR2X1_LOC_275/A OR2X1_LOC_31/Y 0.25fF
C8875 OR2X1_LOC_275/A OR2X1_LOC_12/Y 0.03fF
C44687 OR2X1_LOC_275/A OR2X1_LOC_26/Y 0.04fF
C5121 OR2X1_LOC_275/A OR2X1_LOC_36/Y 0.02fF
C14195 OR2X1_LOC_22/Y OR2X1_LOC_275/A 0.07fF
C37427 OR2X1_LOC_275/A OR2X1_LOC_246/A 0.01fF
C14518 OR2X1_LOC_275/A OR2X1_LOC_39/A 0.04fF
C51883 OR2X1_LOC_589/A OR2X1_LOC_275/A 0.02fF
C52888 OR2X1_LOC_3/Y OR2X1_LOC_275/A 0.05fF
C31347 OR2X1_LOC_158/A OR2X1_LOC_275/A 0.02fF
C13717 OR2X1_LOC_275/A OR2X1_LOC_52/B 0.10fF
C44698 OR2X1_LOC_275/A OR2X1_LOC_89/A 0.03fF
C48519 OR2X1_LOC_275/A OR2X1_LOC_16/A 0.08fF
C43133 OR2X1_LOC_275/A OR2X1_LOC_13/B 0.03fF
C19235 OR2X1_LOC_275/A OR2X1_LOC_74/A 0.08fF
C3538 OR2X1_LOC_273/Y OR2X1_LOC_275/A 0.01fF
C4073 OR2X1_LOC_47/Y OR2X1_LOC_599/Y 0.02fF
C17980 OR2X1_LOC_36/Y OR2X1_LOC_599/Y 0.03fF
C26954 OR2X1_LOC_22/Y OR2X1_LOC_599/Y 0.03fF
C35771 OR2X1_LOC_485/A OR2X1_LOC_599/Y 0.01fF
C8605 OR2X1_LOC_589/A OR2X1_LOC_599/Y 0.03fF
C10819 OR2X1_LOC_64/Y OR2X1_LOC_599/Y 0.21fF
C2374 OR2X1_LOC_95/Y OR2X1_LOC_599/Y 0.25fF
C43766 OR2X1_LOC_45/B OR2X1_LOC_599/Y 3.79fF
C18422 OR2X1_LOC_306/Y OR2X1_LOC_599/Y 0.02fF
C5072 OR2X1_LOC_599/Y OR2X1_LOC_16/A 0.04fF
C56098 OR2X1_LOC_599/Y OR2X1_LOC_13/B 0.08fF
C6924 OR2X1_LOC_599/A OR2X1_LOC_599/Y 0.01fF
C6077 AND2X1_LOC_729/B OR2X1_LOC_599/Y 0.03fF
C55188 AND2X1_LOC_95/Y OR2X1_LOC_461/B 0.51fF
C53124 AND2X1_LOC_56/B OR2X1_LOC_461/B 0.01fF
C30734 AND2X1_LOC_801/B OR2X1_LOC_760/Y 0.81fF
C4255 OR2X1_LOC_271/B OR2X1_LOC_271/Y 0.02fF
C20412 AND2X1_LOC_22/Y AND2X1_LOC_88/Y 0.03fF
C36180 AND2X1_LOC_3/Y AND2X1_LOC_88/Y 0.81fF
C54095 OR2X1_LOC_78/B AND2X1_LOC_88/Y 0.03fF
C24302 AND2X1_LOC_18/Y AND2X1_LOC_88/Y 0.83fF
C29564 AND2X1_LOC_31/Y AND2X1_LOC_88/Y 0.03fF
C15016 OR2X1_LOC_185/A AND2X1_LOC_88/Y 0.03fF
C8648 OR2X1_LOC_100/Y AND2X1_LOC_88/Y 0.01fF
C54997 OR2X1_LOC_689/Y OR2X1_LOC_690/A 0.01fF
C1004 OR2X1_LOC_47/Y AND2X1_LOC_374/Y 0.01fF
C43876 OR2X1_LOC_31/Y AND2X1_LOC_374/Y 0.01fF
C21302 OR2X1_LOC_18/Y AND2X1_LOC_374/Y 0.02fF
C54491 OR2X1_LOC_26/Y AND2X1_LOC_374/Y 0.01fF
C28518 AND2X1_LOC_374/Y OR2X1_LOC_371/Y 0.03fF
C44977 OR2X1_LOC_56/A AND2X1_LOC_374/Y 0.02fF
C39017 OR2X1_LOC_427/A AND2X1_LOC_374/Y 0.03fF
C55436 OR2X1_LOC_95/Y AND2X1_LOC_374/Y 0.01fF
C40553 OR2X1_LOC_45/B AND2X1_LOC_374/Y 0.01fF
C40326 OR2X1_LOC_329/B OR2X1_LOC_47/Y 0.05fF
C23795 OR2X1_LOC_329/B OR2X1_LOC_44/Y 1.24fF
C27249 OR2X1_LOC_329/B OR2X1_LOC_31/Y 0.05fF
C4545 OR2X1_LOC_329/B OR2X1_LOC_18/Y 0.12fF
C39712 OR2X1_LOC_329/B OR2X1_LOC_59/Y 0.04fF
C37659 OR2X1_LOC_329/B OR2X1_LOC_26/Y 0.11fF
C54395 OR2X1_LOC_329/B OR2X1_LOC_36/Y 0.06fF
C7230 OR2X1_LOC_329/B OR2X1_LOC_22/Y 0.94fF
C11883 OR2X1_LOC_329/B OR2X1_LOC_371/Y 0.09fF
C5620 OR2X1_LOC_329/B OR2X1_LOC_437/A 0.11fF
C10391 OR2X1_LOC_329/B OR2X1_LOC_268/Y 0.03fF
C54546 OR2X1_LOC_329/B OR2X1_LOC_419/Y 0.10fF
C28303 OR2X1_LOC_329/B OR2X1_LOC_56/A 0.20fF
C11322 OR2X1_LOC_329/B OR2X1_LOC_91/A 0.07fF
C16098 OR2X1_LOC_329/B OR2X1_LOC_485/A 0.19fF
C7573 OR2X1_LOC_329/B OR2X1_LOC_39/A 0.12fF
C36634 OR2X1_LOC_329/B OR2X1_LOC_428/A 0.31fF
C22483 OR2X1_LOC_329/B OR2X1_LOC_427/A 0.09fF
C43722 OR2X1_LOC_329/B OR2X1_LOC_7/A 0.46fF
C27038 OR2X1_LOC_329/B OR2X1_LOC_744/A 0.57fF
C33765 OR2X1_LOC_329/B OR2X1_LOC_600/A 0.07fF
C47301 OR2X1_LOC_329/B OR2X1_LOC_64/Y 0.61fF
C38628 OR2X1_LOC_329/B OR2X1_LOC_95/Y 0.74fF
C8390 OR2X1_LOC_329/B OR2X1_LOC_51/Y 0.14fF
C43561 OR2X1_LOC_40/Y OR2X1_LOC_329/B 0.46fF
C39845 OR2X1_LOC_70/Y OR2X1_LOC_329/B 0.15fF
C24470 OR2X1_LOC_158/A OR2X1_LOC_329/B 0.88fF
C33852 OR2X1_LOC_329/B OR2X1_LOC_619/Y 0.07fF
C6717 OR2X1_LOC_329/B OR2X1_LOC_52/B 0.19fF
C24054 OR2X1_LOC_45/B OR2X1_LOC_329/B 0.26fF
C37677 OR2X1_LOC_329/B OR2X1_LOC_89/A 0.74fF
C55597 OR2X1_LOC_329/B OR2X1_LOC_164/Y 0.02fF
C41341 OR2X1_LOC_329/B OR2X1_LOC_16/A 0.04fF
C36177 OR2X1_LOC_329/B OR2X1_LOC_13/B 0.07fF
C12321 OR2X1_LOC_329/B OR2X1_LOC_74/A 0.07fF
C54696 OR2X1_LOC_604/A OR2X1_LOC_329/B 0.10fF
C25946 OR2X1_LOC_329/B OR2X1_LOC_111/Y 0.08fF
C28848 OR2X1_LOC_329/B OR2X1_LOC_527/Y 0.02fF
C29259 OR2X1_LOC_329/B AND2X1_LOC_276/Y 0.05fF
C33942 AND2X1_LOC_64/Y OR2X1_LOC_66/Y 0.05fF
C7820 AND2X1_LOC_3/Y OR2X1_LOC_66/Y 0.01fF
C49513 AND2X1_LOC_70/Y OR2X1_LOC_66/Y 0.04fF
C21441 AND2X1_LOC_12/Y OR2X1_LOC_66/Y 0.21fF
C8571 OR2X1_LOC_66/Y AND2X1_LOC_7/B 0.02fF
C29860 OR2X1_LOC_87/A OR2X1_LOC_66/Y 0.03fF
C9627 OR2X1_LOC_473/A OR2X1_LOC_66/Y 0.02fF
C25644 OR2X1_LOC_375/A OR2X1_LOC_66/Y 0.20fF
C55053 AND2X1_LOC_51/Y OR2X1_LOC_66/Y 0.05fF
C25948 OR2X1_LOC_66/Y OR2X1_LOC_549/A 0.04fF
C41257 OR2X1_LOC_160/A OR2X1_LOC_66/Y 0.03fF
C11103 OR2X1_LOC_151/A OR2X1_LOC_66/Y 0.03fF
C36241 OR2X1_LOC_532/B OR2X1_LOC_66/Y 0.03fF
C20089 OR2X1_LOC_66/Y OR2X1_LOC_78/A 0.03fF
C21343 OR2X1_LOC_121/Y OR2X1_LOC_66/Y 0.01fF
C12402 OR2X1_LOC_66/Y OR2X1_LOC_631/A 0.01fF
C26523 AND2X1_LOC_70/Y OR2X1_LOC_121/A 0.03fF
C55120 AND2X1_LOC_59/Y OR2X1_LOC_121/A 0.01fF
C41724 AND2X1_LOC_7/B OR2X1_LOC_121/A 0.05fF
C43493 OR2X1_LOC_160/B OR2X1_LOC_121/A 0.06fF
C32025 OR2X1_LOC_161/A OR2X1_LOC_121/A 0.02fF
C32856 AND2X1_LOC_41/A OR2X1_LOC_121/A 0.05fF
C37562 OR2X1_LOC_269/B OR2X1_LOC_121/A 0.03fF
C29034 AND2X1_LOC_18/Y OR2X1_LOC_121/A 0.09fF
C35267 AND2X1_LOC_36/Y OR2X1_LOC_121/A 0.06fF
C2842 OR2X1_LOC_375/A OR2X1_LOC_121/A 0.73fF
C24227 AND2X1_LOC_47/Y OR2X1_LOC_121/A 0.03fF
C38662 OR2X1_LOC_777/B OR2X1_LOC_121/A 0.03fF
C21549 OR2X1_LOC_541/B OR2X1_LOC_121/A 0.48fF
C9649 OR2X1_LOC_154/A OR2X1_LOC_121/A 0.03fF
C8329 OR2X1_LOC_541/A OR2X1_LOC_121/A 0.01fF
C22882 AND2X1_LOC_56/B OR2X1_LOC_121/A 0.05fF
C22288 AND2X1_LOC_91/B OR2X1_LOC_121/A 0.05fF
C15349 OR2X1_LOC_820/Y OR2X1_LOC_44/Y 0.01fF
C25444 OR2X1_LOC_600/A OR2X1_LOC_820/Y 0.23fF
C37390 OR2X1_LOC_3/Y OR2X1_LOC_820/Y 0.01fF
C16627 OR2X1_LOC_748/A OR2X1_LOC_820/Y 0.01fF
C31457 OR2X1_LOC_820/Y OR2X1_LOC_820/B 0.01fF
C5956 OR2X1_LOC_820/Y AND2X1_LOC_847/Y 0.92fF
C51603 OR2X1_LOC_376/A OR2X1_LOC_409/B 0.01fF
C46950 OR2X1_LOC_548/A AND2X1_LOC_36/Y 0.01fF
C25063 OR2X1_LOC_548/A OR2X1_LOC_532/B 0.06fF
C34210 OR2X1_LOC_548/A AND2X1_LOC_56/B 0.13fF
C1013 OR2X1_LOC_548/A OR2X1_LOC_415/Y 0.01fF
C28769 OR2X1_LOC_185/Y OR2X1_LOC_66/A 0.08fF
C4895 OR2X1_LOC_185/Y AND2X1_LOC_22/Y 5.21fF
C47104 OR2X1_LOC_185/Y AND2X1_LOC_64/Y 0.24fF
C20921 OR2X1_LOC_185/Y AND2X1_LOC_3/Y 0.09fF
C30109 OR2X1_LOC_185/Y AND2X1_LOC_40/Y 0.03fF
C6236 OR2X1_LOC_185/Y AND2X1_LOC_70/Y 0.04fF
C34794 OR2X1_LOC_185/Y AND2X1_LOC_59/Y 0.14fF
C34329 OR2X1_LOC_185/Y AND2X1_LOC_12/Y 6.10fF
C4635 OR2X1_LOC_185/Y AND2X1_LOC_95/Y 0.08fF
C6196 OR2X1_LOC_709/A OR2X1_LOC_185/Y 0.03fF
C45779 OR2X1_LOC_185/Y OR2X1_LOC_435/A 0.05fF
C18543 OR2X1_LOC_185/Y OR2X1_LOC_831/B 0.04fF
C21568 OR2X1_LOC_185/Y AND2X1_LOC_7/B 0.19fF
C47674 OR2X1_LOC_185/Y OR2X1_LOC_756/B 1.09fF
C23335 OR2X1_LOC_185/Y OR2X1_LOC_160/B 0.21fF
C21290 OR2X1_LOC_185/Y OR2X1_LOC_789/B 0.02fF
C38499 OR2X1_LOC_185/Y OR2X1_LOC_78/B 0.10fF
C11910 OR2X1_LOC_185/Y OR2X1_LOC_161/A 0.07fF
C12719 OR2X1_LOC_185/Y AND2X1_LOC_41/A 0.16fF
C37303 OR2X1_LOC_185/Y AND2X1_LOC_81/B 0.10fF
C44463 OR2X1_LOC_185/Y OR2X1_LOC_691/Y 0.03fF
C17437 OR2X1_LOC_185/Y OR2X1_LOC_269/B 3.79fF
C42899 OR2X1_LOC_185/Y OR2X1_LOC_87/A 0.07fF
C18997 OR2X1_LOC_185/Y OR2X1_LOC_161/B 0.12fF
C22741 OR2X1_LOC_185/Y OR2X1_LOC_473/A 0.11fF
C54384 OR2X1_LOC_185/Y OR2X1_LOC_809/B 1.02fF
C8860 OR2X1_LOC_185/Y AND2X1_LOC_18/Y 0.20fF
C15103 OR2X1_LOC_185/Y AND2X1_LOC_36/Y 0.10fF
C38572 OR2X1_LOC_185/Y OR2X1_LOC_375/A 0.03fF
C3958 OR2X1_LOC_185/Y AND2X1_LOC_47/Y 0.16fF
C7955 OR2X1_LOC_185/Y AND2X1_LOC_44/Y 0.12fF
C14231 OR2X1_LOC_185/Y AND2X1_LOC_31/Y 0.22fF
C11967 OR2X1_LOC_185/Y AND2X1_LOC_51/Y 4.12fF
C38893 OR2X1_LOC_185/Y OR2X1_LOC_549/A 0.10fF
C9823 OR2X1_LOC_185/Y OR2X1_LOC_130/A 0.08fF
C45498 OR2X1_LOC_185/Y OR2X1_LOC_154/A 0.54fF
C54459 OR2X1_LOC_185/Y OR2X1_LOC_160/A 0.24fF
C55760 OR2X1_LOC_185/Y OR2X1_LOC_185/A 0.03fF
C24157 OR2X1_LOC_185/Y OR2X1_LOC_151/A 0.25fF
C4218 OR2X1_LOC_185/Y OR2X1_LOC_506/A 0.15fF
C44121 OR2X1_LOC_185/Y OR2X1_LOC_541/A 0.05fF
C49543 OR2X1_LOC_185/Y OR2X1_LOC_532/B 11.79fF
C33017 OR2X1_LOC_185/Y OR2X1_LOC_78/A 0.13fF
C2627 OR2X1_LOC_185/Y AND2X1_LOC_56/B 0.04fF
C1973 OR2X1_LOC_185/Y AND2X1_LOC_91/B 0.10fF
C34207 OR2X1_LOC_121/Y OR2X1_LOC_185/Y 0.11fF
C23065 OR2X1_LOC_185/Y OR2X1_LOC_287/B 0.05fF
C5859 OR2X1_LOC_185/Y OR2X1_LOC_235/B 0.05fF
C26666 OR2X1_LOC_185/Y OR2X1_LOC_800/Y 0.01fF
C32422 OR2X1_LOC_276/B OR2X1_LOC_270/Y 0.10fF
C26966 OR2X1_LOC_276/B OR2X1_LOC_269/Y 0.02fF
C27276 OR2X1_LOC_274/Y OR2X1_LOC_276/B 0.01fF
C49208 OR2X1_LOC_276/B OR2X1_LOC_66/Y 0.03fF
C23647 OR2X1_LOC_22/Y OR2X1_LOC_88/Y 0.03fF
C46627 OR2X1_LOC_71/Y OR2X1_LOC_88/Y 0.07fF
C47076 OR2X1_LOC_246/A OR2X1_LOC_88/Y 0.02fF
C51338 OR2X1_LOC_813/A OR2X1_LOC_88/Y 0.22fF
C50013 OR2X1_LOC_65/B OR2X1_LOC_88/Y 0.03fF
C24009 OR2X1_LOC_88/Y OR2X1_LOC_39/A 0.03fF
C43415 OR2X1_LOC_744/A OR2X1_LOC_88/Y 0.03fF
C7441 OR2X1_LOC_64/Y OR2X1_LOC_88/Y 0.03fF
C6100 OR2X1_LOC_3/Y OR2X1_LOC_88/Y 0.03fF
C173 OR2X1_LOC_70/Y OR2X1_LOC_88/Y 0.02fF
C40299 OR2X1_LOC_45/B OR2X1_LOC_88/Y 0.03fF
C52750 OR2X1_LOC_88/Y OR2X1_LOC_13/B 0.03fF
C39371 OR2X1_LOC_411/Y OR2X1_LOC_44/Y 0.03fF
C23037 OR2X1_LOC_411/Y OR2X1_LOC_22/Y 0.03fF
C6709 OR2X1_LOC_411/Y OR2X1_LOC_690/A 0.10fF
C5554 OR2X1_LOC_411/Y AND2X1_LOC_462/B 0.01fF
C3392 OR2X1_LOC_411/Y OR2X1_LOC_7/A 0.03fF
C24098 OR2X1_LOC_51/Y OR2X1_LOC_411/Y 0.20fF
C22544 OR2X1_LOC_411/Y OR2X1_LOC_52/B 0.03fF
C1908 OR2X1_LOC_691/B OR2X1_LOC_66/A 0.01fF
C20151 AND2X1_LOC_64/Y OR2X1_LOC_691/B 0.03fF
C46689 OR2X1_LOC_691/B OR2X1_LOC_269/B 0.01fF
C44298 OR2X1_LOC_691/B AND2X1_LOC_36/Y 0.03fF
C43378 OR2X1_LOC_691/B AND2X1_LOC_31/Y 0.08fF
C18565 OR2X1_LOC_154/A OR2X1_LOC_691/B 0.01fF
C25101 OR2X1_LOC_847/A AND2X1_LOC_3/Y 0.03fF
C38524 AND2X1_LOC_12/Y OR2X1_LOC_847/A 0.05fF
C41332 OR2X1_LOC_847/A OR2X1_LOC_622/B 0.01fF
C736 OR2X1_LOC_847/A AND2X1_LOC_820/B 0.02fF
C42784 OR2X1_LOC_847/A OR2X1_LOC_78/B 0.03fF
C51359 AND2X1_LOC_82/Y OR2X1_LOC_847/A 0.03fF
C20885 OR2X1_LOC_557/A OR2X1_LOC_847/A 0.05fF
C50941 OR2X1_LOC_847/A OR2X1_LOC_633/A 0.03fF
C2621 AND2X1_LOC_86/B OR2X1_LOC_847/A 1.50fF
C37183 OR2X1_LOC_847/A OR2X1_LOC_78/A 0.03fF
C27213 OR2X1_LOC_287/B OR2X1_LOC_847/A 1.34fF
C18593 OR2X1_LOC_405/A OR2X1_LOC_66/A 0.10fF
C50932 OR2X1_LOC_405/A AND2X1_LOC_22/Y 0.03fF
C36649 AND2X1_LOC_64/Y OR2X1_LOC_405/A 0.11fF
C10676 OR2X1_LOC_405/A AND2X1_LOC_3/Y 2.06fF
C19949 OR2X1_LOC_405/A AND2X1_LOC_40/Y 0.03fF
C52235 OR2X1_LOC_405/A AND2X1_LOC_70/Y 0.54fF
C24643 OR2X1_LOC_405/A AND2X1_LOC_59/Y 0.10fF
C24252 AND2X1_LOC_12/Y OR2X1_LOC_405/A 0.08fF
C50654 OR2X1_LOC_405/A AND2X1_LOC_95/Y 8.69fF
C29562 OR2X1_LOC_405/A AND2X1_LOC_65/A 0.02fF
C34663 OR2X1_LOC_405/A OR2X1_LOC_778/B 0.05fF
C35434 OR2X1_LOC_405/A OR2X1_LOC_435/A 0.08fF
C8356 OR2X1_LOC_405/A OR2X1_LOC_831/B 0.07fF
C19538 OR2X1_LOC_405/A OR2X1_LOC_405/Y 0.14fF
C11289 OR2X1_LOC_405/A AND2X1_LOC_7/B 0.10fF
C37202 OR2X1_LOC_405/A OR2X1_LOC_756/B 0.05fF
C13104 OR2X1_LOC_405/A OR2X1_LOC_160/B 0.07fF
C28364 OR2X1_LOC_405/A OR2X1_LOC_78/B 0.11fF
C1675 OR2X1_LOC_405/A OR2X1_LOC_161/A 0.19fF
C48342 OR2X1_LOC_405/A OR2X1_LOC_446/B 0.06fF
C34168 OR2X1_LOC_405/A OR2X1_LOC_691/Y 0.06fF
C7212 OR2X1_LOC_405/A OR2X1_LOC_269/B 0.42fF
C32649 OR2X1_LOC_405/A OR2X1_LOC_87/A 0.17fF
C8792 OR2X1_LOC_405/A OR2X1_LOC_161/B 0.10fF
C12456 OR2X1_LOC_405/A OR2X1_LOC_473/A 0.01fF
C54746 OR2X1_LOC_405/A AND2X1_LOC_18/Y 0.13fF
C4841 OR2X1_LOC_405/A AND2X1_LOC_36/Y 0.07fF
C28438 OR2X1_LOC_405/A OR2X1_LOC_375/A 0.07fF
C49938 OR2X1_LOC_405/A AND2X1_LOC_47/Y 0.10fF
C3996 OR2X1_LOC_405/A AND2X1_LOC_31/Y 0.57fF
C1759 OR2X1_LOC_405/A AND2X1_LOC_51/Y 0.45fF
C8314 OR2X1_LOC_405/A OR2X1_LOC_777/B 0.11fF
C55736 OR2X1_LOC_405/A OR2X1_LOC_130/A 0.19fF
C35175 OR2X1_LOC_405/A OR2X1_LOC_154/A 0.69fF
C44147 OR2X1_LOC_405/A OR2X1_LOC_160/A 0.90fF
C45447 OR2X1_LOC_405/A OR2X1_LOC_185/A 9.54fF
C13918 OR2X1_LOC_405/A OR2X1_LOC_151/A 0.25fF
C50231 OR2X1_LOC_405/A OR2X1_LOC_506/A 0.03fF
C39094 OR2X1_LOC_405/A OR2X1_LOC_532/B 0.30fF
C22933 OR2X1_LOC_405/A OR2X1_LOC_78/A 0.18fF
C48573 OR2X1_LOC_405/A AND2X1_LOC_56/B 0.01fF
C47957 AND2X1_LOC_91/B OR2X1_LOC_405/A 0.55fF
C983 OR2X1_LOC_47/Y OR2X1_LOC_67/A 0.02fF
C40259 OR2X1_LOC_67/A OR2X1_LOC_44/Y 0.01fF
C18556 OR2X1_LOC_67/A OR2X1_LOC_12/Y 0.03fF
C7568 OR2X1_LOC_122/A OR2X1_LOC_67/A 0.03fF
C44942 OR2X1_LOC_67/A OR2X1_LOC_56/A 1.34fF
C43681 OR2X1_LOC_744/A OR2X1_LOC_67/A 0.03fF
C50576 OR2X1_LOC_600/A OR2X1_LOC_67/A 0.03fF
C7714 OR2X1_LOC_64/Y OR2X1_LOC_67/A 0.03fF
C6353 OR2X1_LOC_3/Y OR2X1_LOC_67/A 0.55fF
C52982 OR2X1_LOC_67/A OR2X1_LOC_13/B 0.03fF
C32486 OR2X1_LOC_375/A OR2X1_LOC_375/Y 0.01fF
C8166 AND2X1_LOC_31/Y OR2X1_LOC_375/Y 0.01fF
C13561 OR2X1_LOC_666/A OR2X1_LOC_44/Y 0.05fF
C50580 OR2X1_LOC_666/A OR2X1_LOC_18/Y 0.17fF
C29548 OR2X1_LOC_666/A OR2X1_LOC_59/Y 0.07fF
C27523 OR2X1_LOC_666/A OR2X1_LOC_26/Y 0.02fF
C44102 OR2X1_LOC_666/A OR2X1_LOC_36/Y 0.03fF
C53216 OR2X1_LOC_666/A OR2X1_LOC_22/Y 0.03fF
C51642 OR2X1_LOC_666/A OR2X1_LOC_437/A 0.03fF
C5875 OR2X1_LOC_666/A OR2X1_LOC_485/A 0.03fF
C53548 OR2X1_LOC_666/A OR2X1_LOC_39/A 0.17fF
C26528 OR2X1_LOC_666/A OR2X1_LOC_428/A 0.02fF
C12215 OR2X1_LOC_666/A OR2X1_LOC_427/A 0.07fF
C16829 OR2X1_LOC_744/A OR2X1_LOC_666/A 0.03fF
C36836 OR2X1_LOC_666/A OR2X1_LOC_64/Y 0.05fF
C35584 OR2X1_LOC_3/Y OR2X1_LOC_666/A 0.01fF
C14269 OR2X1_LOC_158/A OR2X1_LOC_666/A 0.06fF
C27543 OR2X1_LOC_666/A OR2X1_LOC_89/A 0.03fF
C26042 OR2X1_LOC_666/A OR2X1_LOC_13/B 0.02fF
C44408 OR2X1_LOC_604/A OR2X1_LOC_666/A 0.05fF
C3444 AND2X1_LOC_22/Y OR2X1_LOC_374/Y 0.03fF
C45474 AND2X1_LOC_64/Y OR2X1_LOC_374/Y 0.05fF
C4722 AND2X1_LOC_70/Y OR2X1_LOC_374/Y 0.56fF
C32793 AND2X1_LOC_12/Y OR2X1_LOC_374/Y 0.03fF
C39439 OR2X1_LOC_335/A OR2X1_LOC_374/Y 0.03fF
C46036 OR2X1_LOC_756/B OR2X1_LOC_374/Y 0.04fF
C10354 OR2X1_LOC_161/A OR2X1_LOC_374/Y 0.05fF
C15853 OR2X1_LOC_269/B OR2X1_LOC_374/Y 4.83fF
C41277 OR2X1_LOC_87/A OR2X1_LOC_374/Y 0.15fF
C17435 OR2X1_LOC_161/B OR2X1_LOC_374/Y 0.19fF
C36994 OR2X1_LOC_375/A OR2X1_LOC_374/Y 0.06fF
C2377 AND2X1_LOC_47/Y OR2X1_LOC_374/Y 0.25fF
C12643 AND2X1_LOC_31/Y OR2X1_LOC_374/Y 0.04fF
C10426 AND2X1_LOC_51/Y OR2X1_LOC_374/Y 0.01fF
C16954 OR2X1_LOC_777/B OR2X1_LOC_374/Y 0.03fF
C43907 OR2X1_LOC_154/A OR2X1_LOC_374/Y 0.19fF
C54169 OR2X1_LOC_185/A OR2X1_LOC_374/Y 0.03fF
C42562 OR2X1_LOC_541/A OR2X1_LOC_374/Y 0.20fF
C47944 OR2X1_LOC_532/B OR2X1_LOC_374/Y 0.04fF
C410 AND2X1_LOC_91/B OR2X1_LOC_374/Y 0.08fF
C28499 OR2X1_LOC_831/A OR2X1_LOC_374/Y 0.03fF
C50910 OR2X1_LOC_530/Y OR2X1_LOC_437/A -0.00fF
C53602 OR2X1_LOC_530/Y OR2X1_LOC_51/Y 0.31fF
C32650 OR2X1_LOC_47/Y OR2X1_LOC_816/A 0.04fF
C15979 OR2X1_LOC_816/A OR2X1_LOC_44/Y 0.03fF
C53051 OR2X1_LOC_18/Y OR2X1_LOC_816/A 0.03fF
C31977 OR2X1_LOC_816/A OR2X1_LOC_59/Y 0.03fF
C35213 OR2X1_LOC_816/A OR2X1_LOC_753/Y 0.21fF
C46654 OR2X1_LOC_36/Y OR2X1_LOC_816/A 0.19fF
C55675 OR2X1_LOC_22/Y OR2X1_LOC_816/A 0.03fF
C41780 AND2X1_LOC_548/Y OR2X1_LOC_816/A 0.01fF
C54108 OR2X1_LOC_816/A OR2X1_LOC_437/A 0.02fF
C32897 OR2X1_LOC_625/Y OR2X1_LOC_816/A 1.03fF
C17347 OR2X1_LOC_628/Y OR2X1_LOC_816/A 0.04fF
C46854 OR2X1_LOC_419/Y OR2X1_LOC_816/A 0.03fF
C20630 OR2X1_LOC_816/A OR2X1_LOC_56/A 0.01fF
C8443 OR2X1_LOC_485/A OR2X1_LOC_816/A 3.42fF
C56012 OR2X1_LOC_816/A OR2X1_LOC_39/A 0.69fF
C14712 OR2X1_LOC_427/A OR2X1_LOC_816/A 2.22fF
C35917 OR2X1_LOC_7/A OR2X1_LOC_816/A 0.80fF
C19346 OR2X1_LOC_744/A OR2X1_LOC_816/A 0.07fF
C39353 OR2X1_LOC_64/Y OR2X1_LOC_816/A 0.04fF
C592 OR2X1_LOC_51/Y OR2X1_LOC_816/A 0.26fF
C35790 OR2X1_LOC_40/Y OR2X1_LOC_816/A 0.02fF
C16735 OR2X1_LOC_158/A OR2X1_LOC_816/A 0.03fF
C16295 OR2X1_LOC_45/B OR2X1_LOC_816/A 0.03fF
C30020 OR2X1_LOC_89/A OR2X1_LOC_816/A 0.12fF
C28540 OR2X1_LOC_816/A OR2X1_LOC_13/B 0.03fF
C4523 OR2X1_LOC_74/A OR2X1_LOC_816/A 0.04fF
C47016 OR2X1_LOC_604/A OR2X1_LOC_816/A 0.03fF
C44037 AND2X1_LOC_95/Y OR2X1_LOC_410/Y 0.02fF
C30813 OR2X1_LOC_756/B OR2X1_LOC_410/Y 0.11fF
C41907 AND2X1_LOC_56/B OR2X1_LOC_410/Y 0.01fF
C17985 AND2X1_LOC_687/Y AND2X1_LOC_687/B 0.01fF
C13005 OR2X1_LOC_47/Y OR2X1_LOC_760/Y 0.01fF
C44760 OR2X1_LOC_485/A OR2X1_LOC_760/Y 0.01fF
C19736 OR2X1_LOC_64/Y OR2X1_LOC_760/Y 0.06fF
C11251 OR2X1_LOC_95/Y OR2X1_LOC_760/Y 0.04fF
C12491 OR2X1_LOC_70/Y OR2X1_LOC_760/Y 0.04fF
C14078 OR2X1_LOC_760/Y OR2X1_LOC_16/A 0.01fF
C15820 OR2X1_LOC_599/A OR2X1_LOC_760/Y 0.01fF
C16265 OR2X1_LOC_368/A OR2X1_LOC_44/Y 0.03fF
C19768 OR2X1_LOC_31/Y OR2X1_LOC_368/A 0.11fF
C53296 OR2X1_LOC_18/Y OR2X1_LOC_368/A 0.52fF
C46948 OR2X1_LOC_36/Y OR2X1_LOC_368/A 0.01fF
C14987 OR2X1_LOC_427/A OR2X1_LOC_368/A 0.40fF
C31180 OR2X1_LOC_95/Y OR2X1_LOC_368/A 0.05fF
C16531 OR2X1_LOC_45/B OR2X1_LOC_368/A 0.01fF
C37295 OR2X1_LOC_368/A OR2X1_LOC_322/Y 0.01fF
C31396 OR2X1_LOC_271/B OR2X1_LOC_18/Y 0.11fF
C25108 OR2X1_LOC_271/B OR2X1_LOC_36/Y 0.01fF
C14513 OR2X1_LOC_271/B OR2X1_LOC_7/A 0.01fF
C53977 OR2X1_LOC_744/A OR2X1_LOC_271/B 0.04fF
C50960 OR2X1_LOC_45/B OR2X1_LOC_271/B 0.01fF
C8458 OR2X1_LOC_87/Y OR2X1_LOC_66/A 0.16fF
C26571 AND2X1_LOC_64/Y OR2X1_LOC_87/Y 0.03fF
C14472 AND2X1_LOC_59/Y OR2X1_LOC_87/Y 0.03fF
C28474 OR2X1_LOC_87/B OR2X1_LOC_87/Y 0.01fF
C22615 OR2X1_LOC_87/A OR2X1_LOC_87/Y 0.03fF
C43595 OR2X1_LOC_87/Y AND2X1_LOC_44/Y 0.04fF
C33943 OR2X1_LOC_160/A OR2X1_LOC_87/Y 0.15fF
C36040 OR2X1_LOC_47/Y OR2X1_LOC_373/Y 1.57fF
C23006 OR2X1_LOC_31/Y OR2X1_LOC_373/Y 0.01fF
C35370 OR2X1_LOC_59/Y OR2X1_LOC_373/Y 0.15fF
C33384 OR2X1_LOC_26/Y OR2X1_LOC_373/Y 0.31fF
C50318 OR2X1_LOC_419/Y OR2X1_LOC_373/Y 0.03fF
C24057 OR2X1_LOC_56/A OR2X1_LOC_373/Y 0.15fF
C11816 OR2X1_LOC_485/A OR2X1_LOC_373/Y 0.03fF
C3288 OR2X1_LOC_39/A OR2X1_LOC_373/Y 0.05fF
C18102 OR2X1_LOC_427/A OR2X1_LOC_373/Y 0.03fF
C29491 OR2X1_LOC_600/A OR2X1_LOC_373/Y 0.03fF
C42823 OR2X1_LOC_64/Y OR2X1_LOC_373/Y 0.02fF
C34303 OR2X1_LOC_95/Y OR2X1_LOC_373/Y 0.03fF
C35523 OR2X1_LOC_70/Y OR2X1_LOC_373/Y 0.04fF
C33403 OR2X1_LOC_89/A OR2X1_LOC_373/Y 0.06fF
C51325 OR2X1_LOC_164/Y OR2X1_LOC_373/Y 0.03fF
C50464 OR2X1_LOC_604/A OR2X1_LOC_373/Y 0.03fF
C30584 OR2X1_LOC_373/Y OR2X1_LOC_406/A 0.03fF
C44693 OR2X1_LOC_517/A OR2X1_LOC_47/Y 0.02fF
C31453 OR2X1_LOC_517/A OR2X1_LOC_31/Y 0.13fF
C8887 OR2X1_LOC_18/Y OR2X1_LOC_517/A 0.15fF
C44036 OR2X1_LOC_517/A OR2X1_LOC_59/Y 0.03fF
C6138 OR2X1_LOC_517/A OR2X1_LOC_12/Y 0.13fF
C41972 OR2X1_LOC_517/A OR2X1_LOC_26/Y 0.40fF
C11531 OR2X1_LOC_22/Y OR2X1_LOC_517/A 0.20fF
C34387 OR2X1_LOC_517/A OR2X1_LOC_71/Y 0.03fF
C25560 OR2X1_LOC_517/A OR2X1_LOC_256/A 5.09fF
C37641 OR2X1_LOC_517/A OR2X1_LOC_65/B 0.19fF
C44959 OR2X1_LOC_625/Y OR2X1_LOC_517/A 0.01fF
C16553 OR2X1_LOC_490/Y OR2X1_LOC_517/A 1.24fF
C6304 OR2X1_LOC_272/Y OR2X1_LOC_517/A 0.18fF
C32500 OR2X1_LOC_517/A OR2X1_LOC_56/A 0.28fF
C15579 OR2X1_LOC_91/A OR2X1_LOC_517/A 4.66fF
C11851 OR2X1_LOC_517/A OR2X1_LOC_39/A 0.03fF
C49223 OR2X1_LOC_589/A OR2X1_LOC_517/A 0.05fF
C48158 OR2X1_LOC_517/A OR2X1_LOC_7/A 0.15fF
C31277 OR2X1_LOC_744/A OR2X1_LOC_517/A 0.06fF
C37964 OR2X1_LOC_600/A OR2X1_LOC_517/A 0.03fF
C51532 OR2X1_LOC_64/Y OR2X1_LOC_517/A 0.31fF
C42945 OR2X1_LOC_517/A OR2X1_LOC_95/Y 0.13fF
C12608 OR2X1_LOC_51/Y OR2X1_LOC_517/A 0.01fF
C47987 OR2X1_LOC_40/Y OR2X1_LOC_517/A 0.10fF
C50265 OR2X1_LOC_3/Y OR2X1_LOC_517/A 0.12fF
C44184 OR2X1_LOC_70/Y OR2X1_LOC_517/A 0.07fF
C28682 OR2X1_LOC_158/A OR2X1_LOC_517/A 0.01fF
C11020 OR2X1_LOC_517/A OR2X1_LOC_52/B 0.19fF
C41990 OR2X1_LOC_517/A OR2X1_LOC_89/A 0.26fF
C40425 OR2X1_LOC_517/A OR2X1_LOC_13/B 0.10fF
C16555 OR2X1_LOC_517/A OR2X1_LOC_74/A 0.06fF
C20703 OR2X1_LOC_800/A OR2X1_LOC_691/Y 0.01fF
C27939 OR2X1_LOC_687/Y OR2X1_LOC_687/A 0.18fF
C32223 OR2X1_LOC_185/Y OR2X1_LOC_687/Y 0.01fF
C53233 OR2X1_LOC_687/Y OR2X1_LOC_687/B 0.01fF
C22156 OR2X1_LOC_405/A OR2X1_LOC_687/Y 0.01fF
C8573 OR2X1_LOC_800/A OR2X1_LOC_687/Y 0.09fF
C49903 OR2X1_LOC_269/Y OR2X1_LOC_66/A 0.09fF
C42457 OR2X1_LOC_269/Y AND2X1_LOC_7/B 0.01fF
C38272 OR2X1_LOC_269/Y OR2X1_LOC_269/B 0.03fF
C39455 OR2X1_LOC_269/Y OR2X1_LOC_344/A 0.01fF
C29760 OR2X1_LOC_269/Y AND2X1_LOC_18/Y 0.02fF
C35959 OR2X1_LOC_269/Y AND2X1_LOC_36/Y 0.02fF
C3868 OR2X1_LOC_269/Y OR2X1_LOC_549/A 0.01fF
C23551 AND2X1_LOC_56/B OR2X1_LOC_269/Y 0.01fF
C5168 AND2X1_LOC_59/Y OR2X1_LOC_270/Y 0.28fF
C31104 AND2X1_LOC_95/Y OR2X1_LOC_270/Y 0.03fF
C48162 OR2X1_LOC_270/Y AND2X1_LOC_7/B 0.04fF
C17921 OR2X1_LOC_756/B OR2X1_LOC_270/Y 0.10fF
C43900 OR2X1_LOC_270/Y OR2X1_LOC_269/B 0.01fF
C45483 OR2X1_LOC_270/Y OR2X1_LOC_161/B 0.03fF
C45065 OR2X1_LOC_270/Y OR2X1_LOC_344/A 1.08fF
C35224 OR2X1_LOC_270/Y AND2X1_LOC_18/Y 0.01fF
C41500 OR2X1_LOC_270/Y AND2X1_LOC_36/Y 0.01fF
C9429 OR2X1_LOC_270/Y OR2X1_LOC_549/A 0.05fF
C26023 OR2X1_LOC_185/A OR2X1_LOC_270/Y 0.02fF
C19784 OR2X1_LOC_532/B OR2X1_LOC_270/Y 0.03fF
C28997 AND2X1_LOC_56/B OR2X1_LOC_270/Y 0.06fF
C25528 OR2X1_LOC_88/A OR2X1_LOC_26/Y 0.01fF
C21283 OR2X1_LOC_88/A OR2X1_LOC_65/B 0.43fF
C32529 OR2X1_LOC_589/A OR2X1_LOC_88/A 0.01fF
C31307 OR2X1_LOC_40/Y OR2X1_LOC_88/A 0.01fF
C33585 OR2X1_LOC_3/Y OR2X1_LOC_88/A 0.09fF
C15 OR2X1_LOC_88/A OR2X1_LOC_74/A 0.96fF
C22849 OR2X1_LOC_411/A OR2X1_LOC_600/A 0.09fF
C53453 OR2X1_LOC_411/A OR2X1_LOC_51/Y 0.01fF
C30340 OR2X1_LOC_411/A OR2X1_LOC_16/A 0.02fF
C54231 AND2X1_LOC_64/Y OR2X1_LOC_264/Y 0.10fF
C28036 OR2X1_LOC_264/Y AND2X1_LOC_3/Y 0.30fF
C37190 OR2X1_LOC_264/Y AND2X1_LOC_40/Y 0.18fF
C13495 OR2X1_LOC_264/Y AND2X1_LOC_70/Y 0.09fF
C47101 OR2X1_LOC_264/Y AND2X1_LOC_65/A 4.16fF
C30418 OR2X1_LOC_264/Y OR2X1_LOC_160/B 0.03fF
C45789 OR2X1_LOC_264/Y OR2X1_LOC_78/B 0.23fF
C19903 OR2X1_LOC_264/Y AND2X1_LOC_41/A 0.17fF
C44572 OR2X1_LOC_264/Y AND2X1_LOC_81/B 0.03fF
C15973 OR2X1_LOC_264/Y AND2X1_LOC_18/Y 0.22fF
C45860 OR2X1_LOC_264/Y OR2X1_LOC_375/A 0.12fF
C21440 OR2X1_LOC_264/Y AND2X1_LOC_31/Y 0.26fF
C46187 OR2X1_LOC_264/Y OR2X1_LOC_549/A 0.14fF
C40112 OR2X1_LOC_264/Y OR2X1_LOC_78/A 0.11fF
C34494 AND2X1_LOC_40/Y OR2X1_LOC_544/B 0.01fF
C10793 AND2X1_LOC_70/Y OR2X1_LOC_544/B 0.01fF
C38780 AND2X1_LOC_12/Y OR2X1_LOC_544/B 0.07fF
C9141 AND2X1_LOC_95/Y OR2X1_LOC_544/B 0.07fF
C34052 OR2X1_LOC_325/B OR2X1_LOC_544/B 0.23fF
C52079 OR2X1_LOC_756/B OR2X1_LOC_544/B 0.01fF
C27735 OR2X1_LOC_160/B OR2X1_LOC_544/B 0.14fF
C47509 OR2X1_LOC_87/A OR2X1_LOC_544/B 0.08fF
C23536 OR2X1_LOC_161/B OR2X1_LOC_544/B 0.02fF
C8433 AND2X1_LOC_47/Y OR2X1_LOC_544/B 0.09fF
C37016 AND2X1_LOC_687/A OR2X1_LOC_31/Y 0.11fF
C8200 OR2X1_LOC_36/Y AND2X1_LOC_687/A 0.04fF
C21320 OR2X1_LOC_91/A AND2X1_LOC_687/A 0.03fF
C53759 AND2X1_LOC_687/A OR2X1_LOC_7/A 0.03fF
C1000 OR2X1_LOC_64/Y AND2X1_LOC_687/A 0.03fF
C18282 OR2X1_LOC_51/Y AND2X1_LOC_687/A 0.19fF
C55879 OR2X1_LOC_3/Y AND2X1_LOC_687/A 0.04fF
C34291 OR2X1_LOC_158/A AND2X1_LOC_687/A 0.01fF
C16658 AND2X1_LOC_687/A OR2X1_LOC_52/B 0.26fF
C33882 OR2X1_LOC_45/B AND2X1_LOC_687/A 0.02fF
C51452 AND2X1_LOC_687/A OR2X1_LOC_16/A 0.03fF
C8547 OR2X1_LOC_604/A AND2X1_LOC_687/A 0.22fF
C32782 OR2X1_LOC_681/Y AND2X1_LOC_687/A 0.01fF
C16747 OR2X1_LOC_47/Y AND2X1_LOC_687/B 0.07fF
C3597 OR2X1_LOC_31/Y AND2X1_LOC_687/B 0.79fF
C34279 AND2X1_LOC_687/B OR2X1_LOC_12/Y 0.11fF
C39598 OR2X1_LOC_22/Y AND2X1_LOC_687/B 0.03fF
C38273 OR2X1_LOC_684/Y AND2X1_LOC_687/B 0.01fF
C43771 OR2X1_LOC_91/A AND2X1_LOC_687/B 0.07fF
C54934 OR2X1_LOC_427/A AND2X1_LOC_687/B 0.09fF
C20114 AND2X1_LOC_687/B OR2X1_LOC_7/A 0.08fF
C23554 OR2X1_LOC_64/Y AND2X1_LOC_687/B 0.03fF
C40695 OR2X1_LOC_51/Y AND2X1_LOC_687/B 0.03fF
C3839 OR2X1_LOC_694/Y AND2X1_LOC_687/B 0.01fF
C22275 OR2X1_LOC_3/Y AND2X1_LOC_687/B 0.08fF
C16266 OR2X1_LOC_70/Y AND2X1_LOC_687/B 0.22fF
C39119 AND2X1_LOC_687/B OR2X1_LOC_52/B 0.08fF
C342 OR2X1_LOC_45/B AND2X1_LOC_687/B 0.04fF
C17765 AND2X1_LOC_687/B OR2X1_LOC_16/A 0.13fF
C30979 OR2X1_LOC_604/A AND2X1_LOC_687/B 0.01fF
C50597 OR2X1_LOC_685/B OR2X1_LOC_687/A 0.12fF
C45533 OR2X1_LOC_682/Y OR2X1_LOC_36/Y 0.02fF
C2552 OR2X1_LOC_682/Y OR2X1_LOC_91/A 0.01fF
C27896 OR2X1_LOC_682/Y OR2X1_LOC_428/A 0.04fF
C34860 OR2X1_LOC_682/Y OR2X1_LOC_7/A 0.02fF
C38233 OR2X1_LOC_682/Y OR2X1_LOC_64/Y 0.01fF
C36915 OR2X1_LOC_682/Y OR2X1_LOC_3/Y 0.02fF
C15612 OR2X1_LOC_682/Y OR2X1_LOC_158/A 0.35fF
C54085 OR2X1_LOC_682/Y OR2X1_LOC_52/B 0.04fF
C15170 OR2X1_LOC_45/B OR2X1_LOC_682/Y 0.04fF
C12280 OR2X1_LOC_683/Y OR2X1_LOC_12/Y 0.02fF
C16273 OR2X1_LOC_683/Y OR2X1_LOC_684/Y 0.01fF
C32715 OR2X1_LOC_427/A OR2X1_LOC_683/Y 0.01fF
C50404 OR2X1_LOC_70/Y OR2X1_LOC_683/Y 0.01fF
C51884 OR2X1_LOC_683/Y OR2X1_LOC_16/A 0.08fF
C8936 OR2X1_LOC_604/A OR2X1_LOC_683/Y 0.02fF
C56115 OR2X1_LOC_686/B AND2X1_LOC_3/Y 0.12fF
C41365 AND2X1_LOC_70/Y OR2X1_LOC_686/B 0.01fF
C13509 AND2X1_LOC_12/Y OR2X1_LOC_686/B 0.94fF
C17642 OR2X1_LOC_686/B OR2X1_LOC_78/B 0.20fF
C54214 OR2X1_LOC_686/B OR2X1_LOC_161/B 0.27fF
C50534 OR2X1_LOC_635/A OR2X1_LOC_686/B 0.26fF
C49524 OR2X1_LOC_686/B AND2X1_LOC_31/Y 0.01fF
C47262 OR2X1_LOC_686/B AND2X1_LOC_51/Y 0.01fF
C53852 OR2X1_LOC_686/A OR2X1_LOC_686/B 0.13fF
C19626 OR2X1_LOC_685/A AND2X1_LOC_3/Y 0.01fF
C4954 AND2X1_LOC_70/Y OR2X1_LOC_685/A 0.01fF
C53671 OR2X1_LOC_685/A OR2X1_LOC_685/B 0.23fF
C37215 OR2X1_LOC_685/A OR2X1_LOC_78/B 0.01fF
C10644 OR2X1_LOC_685/A OR2X1_LOC_161/A 0.01fF
C41595 OR2X1_LOC_685/A OR2X1_LOC_87/A 0.01fF
C17677 OR2X1_LOC_685/A OR2X1_LOC_161/B 0.03fF
C12957 OR2X1_LOC_685/A AND2X1_LOC_31/Y 0.09fF
C10715 OR2X1_LOC_685/A AND2X1_LOC_51/Y 0.01fF
C393 VDD AND2X1_LOC_119/a_8_24# -0.00fF
C952 VDD OR2X1_LOC_588/a_8_216# 0.21fF
C981 VDD OR2X1_LOC_164/a_8_216# 0.21fF
C1197 VDD OR2X1_LOC_264/a_8_216# 0.21fF
C1679 AND2X1_LOC_55/a_8_24# AND2X1_LOC_414/a_8_24# 0.23fF
C1952 AND2X1_LOC_26/a_8_24# AND2X1_LOC_762/a_8_24# 0.23fF
C2021 VDD OR2X1_LOC_1/a_8_216# 0.21fF
C2372 VDD OR2X1_LOC_129/a_8_216# 0.21fF
C2445 AND2X1_LOC_73/a_8_24# AND2X1_LOC_529/a_8_24# 0.23fF
C2558 VDD OR2X1_LOC_488/a_8_216# 0.21fF
C2631 VDD AND2X1_LOC_270/a_8_24# -0.00fF
C4376 OR2X1_LOC_820/a_8_216# OR2X1_LOC_748/a_8_216# 0.47fF
C4431 VDD OR2X1_LOC_596/a_8_216# 0.21fF
C4935 VDD AND2X1_LOC_129/a_8_24# -0.00fF
C5524 AND2X1_LOC_54/a_8_24# AND2X1_LOC_28/a_8_24# 0.23fF
C5800 VDD AND2X1_LOC_153/a_8_24# -0.00fF
C6146 VDD OR2X1_LOC_743/a_8_216# 0.21fF
C6231 VDD AND2X1_LOC_817/a_8_24# -0.00fF
C6314 AND2X1_LOC_143/a_8_24# AND2X1_LOC_4/a_8_24# 0.23fF
C7856 OR2X1_LOC_693/a_8_216# VDD 0.21fF
C9312 OR2X1_LOC_690/a_8_216# VDD 0.21fF
C9505 VDD OR2X1_LOC_534/a_8_216# 0.21fF
C9919 VDD OR2X1_LOC_377/a_8_216# 0.21fF
C9967 AND2X1_LOC_11/a_8_24# AND2X1_LOC_25/a_8_24# 0.23fF
C10759 OR2X1_LOC_263/a_8_216# OR2X1_LOC_86/a_8_216# 0.47fF
C11216 OR2X1_LOC_111/a_8_216# VDD 0.21fF
C12378 VDD OR2X1_LOC_276/a_8_216# 0.21fF
C13573 VDD OR2X1_LOC_688/a_8_216# 0.21fF
C14028 AND2X1_LOC_588/a_8_24# AND2X1_LOC_36/a_8_24# 0.23fF
C14162 OR2X1_LOC_92/a_8_216# OR2X1_LOC_63/a_8_216# 0.47fF
C15450 VDD AND2X1_LOC_760/a_8_24# -0.00fF
C15600 AND2X1_LOC_819/a_8_24# AND2X1_LOC_618/a_8_24# 0.23fF
C16426 VDD AND2X1_LOC_748/a_8_24# -0.00fF
C16723 OR2X1_LOC_110/a_8_216# VDD 0.21fF
C17002 VDD OR2X1_LOC_268/a_8_216# 0.21fF
C17164 AND2X1_LOC_90/a_8_24# AND2X1_LOC_277/a_8_24# 0.23fF
C17498 OR2X1_LOC_44/a_8_216# OR2X1_LOC_47/a_8_216# 0.47fF
C18056 OR2X1_LOC_369/a_8_216# OR2X1_LOC_309/a_8_216# 0.47fF
C18623 VDD OR2X1_LOC_618/a_8_216# 0.21fF
C18963 VDD OR2X1_LOC_294/a_8_216# 0.21fF
C18999 VDD OR2X1_LOC_46/a_8_216# 0.21fF
C19844 VDD AND2X1_LOC_48/a_8_24# -0.00fF
C19884 VDD AND2X1_LOC_398/a_8_24# -0.00fF
C19911 VDD OR2X1_LOC_87/a_8_216# 0.21fF
C20857 VDD AND2X1_LOC_133/a_8_24# -0.00fF
C21250 AND2X1_LOC_22/a_8_24# AND2X1_LOC_47/a_8_24# 0.23fF
C22467 AND2X1_LOC_95/a_8_24# AND2X1_LOC_59/a_8_24# 0.23fF
C22630 VDD OR2X1_LOC_55/a_8_216# 0.21fF
C23464 OR2X1_LOC_827/a_8_216# OR2X1_LOC_42/a_8_216# 0.47fF
C24670 OR2X1_LOC_53/a_8_216# OR2X1_LOC_752/a_8_216# 0.47fF
C24953 VDD OR2X1_LOC_628/a_8_216# 0.21fF
C26115 VDD OR2X1_LOC_323/a_8_216# 0.21fF
C26553 OR2X1_LOC_681/a_8_216# VDD 0.21fF
C26767 VDD OR2X1_LOC_818/a_8_216# 0.21fF
C26925 OR2X1_LOC_696/a_8_216# OR2X1_LOC_511/a_8_216# 0.47fF
C27094 AND2X1_LOC_80/a_8_24# VDD -0.00fF
C27495 VDD OR2X1_LOC_95/a_8_216# 0.21fF
C27818 AND2X1_LOC_323/a_8_24# AND2X1_LOC_299/a_8_24# 0.23fF
C28058 OR2X1_LOC_291/a_8_216# OR2X1_LOC_278/a_8_216# 0.47fF
C28176 AND2X1_LOC_102/a_8_24# AND2X1_LOC_672/a_8_24# 0.23fF
C28213 OR2X1_LOC_136/a_8_216# VDD 0.21fF
C28625 VDD AND2X1_LOC_407/a_8_24# -0.00fF
C28920 VDD OR2X1_LOC_2/a_8_216# 0.21fF
C29194 AND2X1_LOC_382/a_8_24# VDD -0.00fF
C29874 VDD OR2X1_LOC_502/a_8_216# 0.21fF
C29915 OR2X1_LOC_691/a_8_216# VDD 0.21fF
C30323 OR2X1_LOC_304/a_8_216# VDD 0.21fF
C30868 VDD AND2X1_LOC_375/a_8_24# -0.00fF
C31143 OR2X1_LOC_143/a_8_216# VDD 0.21fF
C31598 VDD OR2X1_LOC_310/a_8_216# 0.21fF
C31784 VDD OR2X1_LOC_119/a_8_216# 0.21fF
C31820 VDD AND2X1_LOC_56/a_8_24# -0.00fF
C32247 VDD OR2X1_LOC_619/a_8_216# 0.21fF
C32348 VDD AND2X1_LOC_619/a_8_24# -0.00fF
C33278 VDD AND2X1_LOC_255/a_8_24# -0.00fF
C33295 AND2X1_LOC_70/a_8_24# AND2X1_LOC_40/a_8_24# 0.23fF
C33922 OR2X1_LOC_54/a_8_216# OR2X1_LOC_9/a_8_216# 0.47fF
C33996 AND2X1_LOC_63/a_8_24# AND2X1_LOC_10/a_8_24# 0.23fF
C34346 AND2X1_LOC_599/a_8_24# AND2X1_LOC_761/a_8_24# 0.23fF
C35454 AND2X1_LOC_752/a_8_24# VDD -0.00fF
C35852 VDD OR2X1_LOC_686/a_8_216# 0.21fF
C36681 OR2X1_LOC_15/a_8_216# OR2X1_LOC_38/a_8_216# 0.47fF
C38124 VDD AND2X1_LOC_692/a_8_24# -0.00fF
C40393 OR2X1_LOC_157/a_8_216# OR2X1_LOC_51/a_8_216# 0.47fF
C40420 OR2X1_LOC_57/a_8_216# OR2X1_LOC_19/a_8_216# 0.47fF
C41086 VDD AND2X1_LOC_10/a_8_24# -0.00fF
C41579 VDD AND2X1_LOC_309/a_8_24# -0.00fF
C42666 OR2X1_LOC_246/a_8_216# OR2X1_LOC_150/a_8_216# 0.47fF
C43613 VDD AND2X1_LOC_155/a_8_24# -0.00fF
C44426 VDD AND2X1_LOC_144/a_8_24# -0.00fF
C44623 VDD AND2X1_LOC_5/a_8_24# -0.00fF
C44947 VDD OR2X1_LOC_699/a_8_216# 0.21fF
C45476 VDD OR2X1_LOC_750/a_8_216# 0.21fF
C47948 VDD AND2X1_LOC_86/a_8_24# -0.00fF
C49338 VDD OR2X1_LOC_82/a_8_216# 0.21fF
C49720 OR2X1_LOC_519/a_8_216# VDD 0.21fF
C50139 VDD AND2X1_LOC_820/a_8_24# -0.00fF
C50354 AND2X1_LOC_82/a_8_24# AND2X1_LOC_77/a_8_24# 0.23fF
C51591 VDD OR2X1_LOC_761/a_8_216# 0.21fF
C51803 VDD OR2X1_LOC_814/a_8_216# 0.21fF
C51956 AND2X1_LOC_1/a_8_24# AND2X1_LOC_17/a_8_24# 0.23fF
C53403 OR2X1_LOC_274/a_8_216# OR2X1_LOC_120/a_8_216# 0.47fF
C54508 VDD OR2X1_LOC_289/a_8_216# 0.21fF
C55431 OR2X1_LOC_233/a_8_216# OR2X1_LOC_62/a_8_216# 0.47fF
C56314 AND2X1_LOC_750/a_8_24# VSS 0.10fF
C56331 AND2X1_LOC_419/a_8_24# VSS 0.10fF
C56410 AND2X1_LOC_225/a_8_24# VSS 0.10fF
C56467 AND2X1_LOC_405/a_8_24# VSS 0.10fF
C56501 AND2X1_LOC_289/a_8_24# VSS 0.10fF
C56503 AND2X1_LOC_278/a_8_24# VSS 0.10fF
C56504 AND2X1_LOC_245/a_8_24# VSS 0.10fF
C56523 AND2X1_LOC_426/a_8_24# VSS 0.10fF
C56597 AND2X1_LOC_276/a_8_24# VSS 0.10fF
C56662 AND2X1_LOC_264/a_8_24# VSS 0.10fF
C56666 AND2X1_LOC_275/a_8_24# VSS 0.10fF
C56701 AND2X1_LOC_818/a_8_24# VSS 0.10fF
C56715 AND2X1_LOC_296/a_8_24# VSS 0.10fF
C56720 AND2X1_LOC_263/a_8_24# VSS 0.10fF
C56741 AND2X1_LOC_433/a_8_24# VSS 0.10fF
C56777 AND2X1_LOC_273/a_8_24# VSS 0.10fF
C56858 AND2X1_LOC_9/a_8_24# VSS 0.10fF
C56963 AND2X1_LOC_687/a_8_24# VSS 0.10fF
C56985 AND2X1_LOC_19/a_8_24# VSS 0.10fF
C56989 AND2X1_LOC_461/a_8_24# VSS 0.10fF
C57064 AND2X1_LOC_696/a_8_24# VSS 0.10fF
C57190 AND2X1_LOC_37/a_8_24# VSS 0.10fF
C57215 AND2X1_LOC_693/a_8_24# VSS 0.10fF
C57225 AND2X1_LOC_126/a_8_24# VSS 0.10fF
C57296 AND2X1_LOC_57/a_8_24# VSS 0.10fF
C57350 AND2X1_LOC_23/a_8_24# VSS 0.10fF
C57377 AND2X1_LOC_690/a_8_24# VSS 0.10fF
C57463 AND2X1_LOC_21/a_8_24# VSS 0.10fF
C57465 AND2X1_LOC_43/a_8_24# VSS 0.10fF
C57511 AND2X1_LOC_110/a_8_24# VSS 0.10fF
C57530 AND2X1_LOC_53/a_8_24# VSS 0.10fF
C57535 AND2X1_LOC_42/a_8_24# VSS 0.10fF
C57596 AND2X1_LOC_30/a_8_24# VSS 0.10fF
C57604 AND2X1_LOC_378/a_8_24# VSS 0.10fF
C57750 AND2X1_LOC_513/a_8_24# VSS 0.10fF
C57777 AND2X1_LOC_71/a_8_24# VSS 0.10fF
C57779 AND2X1_LOC_93/a_8_24# VSS 0.10fF
C57816 AND2X1_LOC_512/a_8_24# VSS 0.10fF
C57828 VDD VSS 2.10fF
C57893 AND2X1_LOC_80/a_8_24# VSS 0.10fF
C57943 AND2X1_LOC_372/a_8_24# VSS 0.10fF
C57991 AND2X1_LOC_585/a_8_24# VSS 0.10fF
C58113 AND2X1_LOC_582/a_8_24# VSS 0.10fF
C2296 OR2X1_LOC_66/A AND2X1_LOC_246/a_8_24# 0.02fF
C4707 OR2X1_LOC_66/a_8_216# OR2X1_LOC_66/A 0.04fF
C6111 OR2X1_LOC_66/A OR2X1_LOC_548/a_36_216# 0.02fF
C7603 AND2X1_LOC_42/a_36_24# OR2X1_LOC_66/A 0.01fF
C7870 AND2X1_LOC_93/a_8_24# OR2X1_LOC_66/A 0.01fF
C9789 AND2X1_LOC_689/a_8_24# OR2X1_LOC_66/A 0.17fF
C10506 AND2X1_LOC_57/a_8_24# OR2X1_LOC_66/A 0.02fF
C13179 OR2X1_LOC_688/Y OR2X1_LOC_66/A 0.01fF
C14332 AND2X1_LOC_421/a_8_24# OR2X1_LOC_66/A 0.03fF
C20376 AND2X1_LOC_38/a_8_24# OR2X1_LOC_66/A 0.04fF
C21215 AND2X1_LOC_696/a_8_24# OR2X1_LOC_66/A 0.03fF
C22816 OR2X1_LOC_66/A AND2X1_LOC_417/a_8_24# 0.02fF
C23662 OR2X1_LOC_66/A AND2X1_LOC_245/a_8_24# 0.05fF
C25310 AND2X1_LOC_86/a_8_24# OR2X1_LOC_66/A 0.01fF
C27364 AND2X1_LOC_263/a_8_24# OR2X1_LOC_66/A 0.01fF
C27435 AND2X1_LOC_529/a_8_24# OR2X1_LOC_66/A 0.04fF
C38393 AND2X1_LOC_529/a_36_24# OR2X1_LOC_66/A 0.01fF
C40287 OR2X1_LOC_276/B OR2X1_LOC_66/A 0.07fF
C47227 OR2X1_LOC_688/a_8_216# OR2X1_LOC_66/A 0.02fF
C50533 AND2X1_LOC_126/a_8_24# OR2X1_LOC_66/A -0.00fF
C51282 OR2X1_LOC_66/A OR2X1_LOC_548/a_8_216# 0.02fF
C52208 AND2X1_LOC_690/a_8_24# OR2X1_LOC_66/A 0.17fF
C52732 AND2X1_LOC_42/a_8_24# OR2X1_LOC_66/A 0.02fF
C53118 AND2X1_LOC_824/a_8_24# OR2X1_LOC_66/A 0.03fF
C53543 OR2X1_LOC_87/a_8_216# OR2X1_LOC_66/A 0.22fF
C54963 OR2X1_LOC_66/A OR2X1_LOC_398/a_8_216# 0.03fF
C55754 OR2X1_LOC_606/a_8_216# OR2X1_LOC_66/A 0.01fF
C565 AND2X1_LOC_22/Y AND2X1_LOC_511/a_8_24# 0.02fF
C1555 AND2X1_LOC_22/Y AND2X1_LOC_369/a_8_24# 0.09fF
C2479 AND2X1_LOC_22/Y AND2X1_LOC_18/a_8_24# 0.01fF
C3030 AND2X1_LOC_22/Y AND2X1_LOC_289/a_8_24# 0.02fF
C3579 AND2X1_LOC_22/Y AND2X1_LOC_263/a_8_24# 0.05fF
C6137 AND2X1_LOC_22/Y AND2X1_LOC_328/a_8_24# 0.01fF
C6982 AND2X1_LOC_22/Y AND2X1_LOC_306/a_8_24# 0.04fF
C9142 AND2X1_LOC_22/Y AND2X1_LOC_95/a_8_24# 0.02fF
C14626 AND2X1_LOC_22/Y AND2X1_LOC_263/a_36_24# 0.01fF
C17969 AND2X1_LOC_22/Y AND2X1_LOC_273/a_8_24# 0.01fF
C19006 AND2X1_LOC_22/Y AND2X1_LOC_683/a_8_24# 0.11fF
C27394 AND2X1_LOC_22/Y AND2X1_LOC_71/a_8_24# 0.03fF
C27872 AND2X1_LOC_22/Y AND2X1_LOC_26/a_8_24# 0.02fF
C28647 AND2X1_LOC_22/Y AND2X1_LOC_304/a_8_24# 0.01fF
C28679 AND2X1_LOC_22/Y AND2X1_LOC_59/a_8_24# 0.02fF
C29510 AND2X1_LOC_22/Y AND2X1_LOC_48/a_8_24# 0.02fF
C33380 AND2X1_LOC_22/Y AND2X1_LOC_386/a_8_24# 0.02fF
C43975 AND2X1_LOC_22/Y AND2X1_LOC_71/a_36_24# 0.01fF
C45790 AND2X1_LOC_22/Y AND2X1_LOC_43/a_8_24# 0.04fF
C51445 AND2X1_LOC_22/Y AND2X1_LOC_309/a_8_24# 0.10fF
C53313 AND2X1_LOC_22/Y OR2X1_LOC_598/a_8_216# 0.03fF
C637 AND2X1_LOC_64/Y AND2X1_LOC_129/a_8_24# 0.02fF
C1525 AND2X1_LOC_64/Y AND2X1_LOC_153/a_8_24# 0.01fF
C1559 AND2X1_LOC_64/Y OR2X1_LOC_296/a_8_216# 0.01fF
C6606 AND2X1_LOC_64/Y AND2X1_LOC_88/a_8_24# 0.02fF
C10288 AND2X1_LOC_64/Y AND2X1_LOC_419/a_36_24# -0.00fF
C13417 AND2X1_LOC_64/Y AND2X1_LOC_71/a_8_24# 0.01fF
C14673 AND2X1_LOC_64/Y OR2X1_LOC_294/a_8_216# 0.01fF
C25604 AND2X1_LOC_64/Y OR2X1_LOC_502/a_8_216# 0.01fF
C25650 AND2X1_LOC_64/Y OR2X1_LOC_691/a_8_216# 0.01fF
C27519 AND2X1_LOC_64/Y AND2X1_LOC_56/a_8_24# 0.02fF
C29978 AND2X1_LOC_64/Y OR2X1_LOC_68/a_8_216# 0.01fF
C30783 OR2X1_LOC_100/a_8_216# AND2X1_LOC_64/Y 0.01fF
C33706 AND2X1_LOC_64/Y AND2X1_LOC_310/a_8_24# 0.01fF
C36576 AND2X1_LOC_64/Y AND2X1_LOC_433/a_8_24# 0.04fF
C41347 AND2X1_LOC_64/Y AND2X1_LOC_527/a_8_24# 0.18fF
C43909 AND2X1_LOC_64/Y OR2X1_LOC_185/a_8_216# 0.01fF
C47870 AND2X1_LOC_64/Y AND2X1_LOC_433/a_36_24# 0.01fF
C5553 AND2X1_LOC_43/a_8_24# AND2X1_LOC_3/Y 0.01fF
C8294 AND2X1_LOC_3/Y AND2X1_LOC_761/a_8_24# 0.01fF
C12476 AND2X1_LOC_681/a_8_24# AND2X1_LOC_3/Y 0.02fF
C13048 AND2X1_LOC_3/Y OR2X1_LOC_598/a_8_216# 0.01fF
C15836 AND2X1_LOC_684/a_8_24# AND2X1_LOC_3/Y 0.02fF
C16966 AND2X1_LOC_110/a_8_24# AND2X1_LOC_3/Y 0.02fF
C17295 AND2X1_LOC_599/a_8_24# AND2X1_LOC_3/Y 0.01fF
C18380 AND2X1_LOC_18/a_8_24# AND2X1_LOC_3/Y 0.03fF
C18456 AND2X1_LOC_699/a_8_24# AND2X1_LOC_3/Y 0.01fF
C21291 OR2X1_LOC_814/a_8_216# AND2X1_LOC_3/Y 0.02fF
C24960 AND2X1_LOC_743/a_8_24# AND2X1_LOC_3/Y 0.03fF
C25134 OR2X1_LOC_685/B AND2X1_LOC_3/Y 0.01fF
C26806 OR2X1_LOC_264/a_8_216# AND2X1_LOC_3/Y 0.01fF
C30560 AND2X1_LOC_682/a_8_24# AND2X1_LOC_3/Y 0.02fF
C31460 OR2X1_LOC_296/a_8_216# AND2X1_LOC_3/Y 0.01fF
C31874 AND2X1_LOC_490/a_8_24# AND2X1_LOC_3/Y 0.02fF
C34867 AND2X1_LOC_683/a_8_24# AND2X1_LOC_3/Y 0.02fF
C41459 AND2X1_LOC_3/Y AND2X1_LOC_488/a_8_24# 0.02fF
C42031 AND2X1_LOC_748/a_8_24# AND2X1_LOC_3/Y 0.08fF
C44592 OR2X1_LOC_294/a_8_216# AND2X1_LOC_3/Y 0.15fF
C44966 OR2X1_LOC_686/A AND2X1_LOC_3/Y 0.03fF
C48660 AND2X1_LOC_3/Y AND2X1_LOC_425/a_8_24# 0.20fF
C50282 OR2X1_LOC_327/a_8_216# AND2X1_LOC_3/Y 0.01fF
C52956 AND2X1_LOC_3/Y OR2X1_LOC_66/a_8_216# 0.07fF
C55631 AND2X1_LOC_585/a_8_24# AND2X1_LOC_3/Y 0.01fF
C1243 AND2X1_LOC_40/Y OR2X1_LOC_407/a_8_216# 0.01fF
C5870 AND2X1_LOC_40/Y AND2X1_LOC_80/a_8_24# 0.01fF
C8735 AND2X1_LOC_40/Y OR2X1_LOC_502/a_8_216# 0.01fF
C14002 OR2X1_LOC_100/a_8_216# AND2X1_LOC_40/Y 0.01fF
C15169 AND2X1_LOC_763/a_8_24# AND2X1_LOC_40/Y 0.01fF
C17271 AND2X1_LOC_40/Y AND2X1_LOC_387/a_8_24# 0.17fF
C17518 AND2X1_LOC_40/Y AND2X1_LOC_761/a_8_24# 0.17fF
C24661 AND2X1_LOC_40/Y AND2X1_LOC_373/a_8_24# 0.01fF
C31329 AND2X1_LOC_40/Y AND2X1_LOC_328/a_8_24# 0.04fF
C39271 AND2X1_LOC_40/Y OR2X1_LOC_596/a_8_216# 0.09fF
C41788 AND2X1_LOC_40/Y AND2X1_LOC_226/a_8_24# 0.03fF
C42375 AND2X1_LOC_40/Y AND2X1_LOC_328/a_36_24# 0.01fF
C1339 AND2X1_LOC_70/Y AND2X1_LOC_684/a_8_24# 0.01fF
C2408 AND2X1_LOC_70/Y AND2X1_LOC_110/a_8_24# 0.01fF
C10565 AND2X1_LOC_70/Y OR2X1_LOC_685/B 0.01fF
C11263 AND2X1_LOC_70/Y AND2X1_LOC_40/a_8_24# 0.01fF
C16012 AND2X1_LOC_70/Y AND2X1_LOC_682/a_8_24# 0.01fF
C17879 AND2X1_LOC_70/Y OR2X1_LOC_276/B 0.36fF
C19349 AND2X1_LOC_70/Y AND2X1_LOC_256/a_8_24# 0.02fF
C20260 AND2X1_LOC_70/Y AND2X1_LOC_628/a_8_24# 0.01fF
C20373 AND2X1_LOC_70/Y AND2X1_LOC_683/a_8_24# 0.01fF
C21068 AND2X1_LOC_70/Y AND2X1_LOC_275/a_8_24# 0.01fF
C23478 AND2X1_LOC_70/Y OR2X1_LOC_276/a_8_216# 0.01fF
C24971 AND2X1_LOC_70/Y OR2X1_LOC_405/a_8_216# 0.01fF
C27339 AND2X1_LOC_70/Y OR2X1_LOC_374/a_8_216# 0.17fF
C29988 AND2X1_LOC_70/Y OR2X1_LOC_294/a_8_216# 0.01fF
C30370 AND2X1_LOC_70/Y OR2X1_LOC_686/A 0.03fF
C31632 AND2X1_LOC_70/Y AND2X1_LOC_625/a_8_24# 0.01fF
C38214 AND2X1_LOC_70/Y OR2X1_LOC_66/a_8_216# 0.01fF
C40076 AND2X1_LOC_70/a_8_24# AND2X1_LOC_70/Y 0.01fF
C40938 AND2X1_LOC_70/Y AND2X1_LOC_164/a_8_24# 0.01fF
C49665 AND2X1_LOC_70/Y AND2X1_LOC_387/a_8_24# 0.01fF
C51944 AND2X1_LOC_70/Y AND2X1_LOC_23/a_8_24# 0.01fF
C52125 AND2X1_LOC_70/Y AND2X1_LOC_433/a_8_24# 0.04fF
C54077 AND2X1_LOC_70/Y AND2X1_LOC_681/a_8_24# 0.01fF
C555 OR2X1_LOC_47/Y OR2X1_LOC_3/a_8_216# 0.01fF
C634 OR2X1_LOC_47/Y OR2X1_LOC_234/a_36_216# 0.03fF
C1410 OR2X1_LOC_47/Y OR2X1_LOC_48/a_8_216# 0.07fF
C1924 OR2X1_LOC_47/Y OR2X1_LOC_760/a_8_216# 0.01fF
C4567 OR2X1_LOC_47/Y OR2X1_LOC_386/a_8_216# 0.01fF
C4796 OR2X1_LOC_47/Y AND2X1_LOC_294/a_8_24# 0.02fF
C7231 OR2X1_LOC_329/a_8_216# OR2X1_LOC_47/Y 0.01fF
C10763 OR2X1_LOC_47/Y OR2X1_LOC_256/a_8_216# 0.01fF
C11244 OR2X1_LOC_47/Y OR2X1_LOC_54/a_8_216# 0.06fF
C11484 OR2X1_LOC_47/Y OR2X1_LOC_18/a_8_216# 0.01fF
C12535 OR2X1_LOC_80/a_8_216# OR2X1_LOC_47/Y 0.01fF
C14067 OR2X1_LOC_47/Y OR2X1_LOC_373/a_8_216# 0.01fF
C17019 OR2X1_LOC_47/Y OR2X1_LOC_322/a_8_216# 0.01fF
C18311 OR2X1_LOC_102/a_8_216# OR2X1_LOC_47/Y 0.01fF
C20292 OR2X1_LOC_47/Y OR2X1_LOC_164/a_8_216# 0.01fF
C20982 OR2X1_LOC_529/a_8_216# OR2X1_LOC_47/Y 0.01fF
C21765 OR2X1_LOC_129/a_8_216# OR2X1_LOC_47/Y 0.02fF
C23146 OR2X1_LOC_47/Y OR2X1_LOC_371/a_8_216# 0.14fF
C23670 OR2X1_LOC_47/Y AND2X1_LOC_405/a_8_24# 0.01fF
C24970 OR2X1_LOC_47/Y OR2X1_LOC_599/a_8_216# 0.01fF
C25150 OR2X1_LOC_47/Y OR2X1_LOC_12/a_8_216# -0.00fF
C25175 AND2X1_LOC_374/a_8_24# OR2X1_LOC_47/Y 0.01fF
C27214 OR2X1_LOC_693/a_8_216# OR2X1_LOC_47/Y 0.06fF
C31926 AND2X1_LOC_598/a_8_24# OR2X1_LOC_47/Y 0.01fF
C32329 OR2X1_LOC_47/Y OR2X1_LOC_246/a_8_216# 0.01fF
C36198 OR2X1_LOC_277/a_8_216# OR2X1_LOC_47/Y 0.01fF
C38724 OR2X1_LOC_47/Y OR2X1_LOC_22/a_8_216# 0.39fF
C41336 OR2X1_LOC_47/Y OR2X1_LOC_64/a_8_216# 0.14fF
C44287 OR2X1_LOC_628/a_8_216# OR2X1_LOC_47/Y 0.01fF
C44916 OR2X1_LOC_47/Y OR2X1_LOC_150/a_8_216# 0.01fF
C45709 OR2X1_LOC_47/Y OR2X1_LOC_234/a_8_216# 0.05fF
C47028 OR2X1_LOC_47/Y AND2X1_LOC_800/a_8_24# 0.01fF
C47824 OR2X1_LOC_47/Y OR2X1_LOC_40/a_8_216# 0.11fF
C49632 OR2X1_LOC_255/a_8_216# OR2X1_LOC_47/Y 0.01fF
C52480 OR2X1_LOC_694/a_8_216# OR2X1_LOC_47/Y 0.01fF
C52561 OR2X1_LOC_47/Y AND2X1_LOC_801/B 0.01fF
C52889 OR2X1_LOC_47/Y OR2X1_LOC_59/a_8_216# 0.14fF
C3605 OR2X1_LOC_44/Y OR2X1_LOC_588/a_8_216# 0.19fF
C5253 OR2X1_LOC_44/Y AND2X1_LOC_750/a_8_24# 0.01fF
C5854 OR2X1_LOC_819/a_8_216# OR2X1_LOC_44/Y 0.01fF
C6830 OR2X1_LOC_696/a_8_216# OR2X1_LOC_44/Y 0.02fF
C9706 OR2X1_LOC_57/a_8_216# OR2X1_LOC_44/Y 0.01fF
C11012 OR2X1_LOC_692/a_8_216# OR2X1_LOC_44/Y 0.01fF
C11414 AND2X1_LOC_296/a_8_24# OR2X1_LOC_44/Y 0.04fF
C16672 AND2X1_LOC_293/a_8_24# OR2X1_LOC_44/Y 0.02fF
C16964 OR2X1_LOC_820/A OR2X1_LOC_44/Y 0.01fF
C17430 OR2X1_LOC_433/a_8_216# OR2X1_LOC_44/Y 0.01fF
C19073 AND2X1_LOC_121/a_8_24# OR2X1_LOC_44/Y 0.01fF
C20680 OR2X1_LOC_44/Y OR2X1_LOC_748/a_8_216# 0.01fF
C20940 AND2X1_LOC_847/a_8_24# OR2X1_LOC_44/Y 0.01fF
C21452 OR2X1_LOC_44/Y OR2X1_LOC_511/a_8_216# 0.05fF
C24791 OR2X1_LOC_64/a_8_216# OR2X1_LOC_44/Y 0.01fF
C26859 OR2X1_LOC_412/a_8_216# OR2X1_LOC_44/Y 0.06fF
C27976 AND2X1_LOC_296/a_36_24# OR2X1_LOC_44/Y 0.01fF
C30105 OR2X1_LOC_763/a_8_216# OR2X1_LOC_44/Y 0.01fF
C30164 OR2X1_LOC_95/a_8_216# OR2X1_LOC_44/Y 0.06fF
C31731 AND2X1_LOC_596/a_8_24# OR2X1_LOC_44/Y 0.01fF
C34876 OR2X1_LOC_762/a_8_216# OR2X1_LOC_44/Y 0.01fF
C34959 OR2X1_LOC_44/Y OR2X1_LOC_749/a_8_216# 0.01fF
C36795 OR2X1_LOC_26/a_8_216# OR2X1_LOC_44/Y 0.01fF
C41014 OR2X1_LOC_820/a_8_216# OR2X1_LOC_44/Y 0.01fF
C44673 OR2X1_LOC_817/a_8_216# OR2X1_LOC_44/Y 0.01fF
C51612 AND2X1_LOC_66/a_8_24# OR2X1_LOC_44/Y 0.01fF
C1003 OR2X1_LOC_31/Y OR2X1_LOC_47/a_8_216# 0.01fF
C2224 OR2X1_LOC_689/A OR2X1_LOC_31/Y 0.23fF
C2241 OR2X1_LOC_31/Y AND2X1_LOC_274/a_8_24# 0.01fF
C3835 OR2X1_LOC_31/Y OR2X1_LOC_322/a_8_216# 0.01fF
C7021 OR2X1_LOC_31/Y OR2X1_LOC_588/a_8_216# 0.03fF
C7058 OR2X1_LOC_31/Y OR2X1_LOC_164/a_8_216# 0.01fF
C7910 OR2X1_LOC_31/Y OR2X1_LOC_153/a_8_216# 0.01fF
C10355 OR2X1_LOC_696/a_8_216# OR2X1_LOC_31/Y 0.01fF
C11940 OR2X1_LOC_31/Y OR2X1_LOC_12/a_8_216# 0.01fF
C11962 AND2X1_LOC_374/a_8_24# OR2X1_LOC_31/Y 0.02fF
C15285 OR2X1_LOC_527/a_8_216# OR2X1_LOC_31/Y 0.14fF
C17345 OR2X1_LOC_111/a_8_216# OR2X1_LOC_31/Y 0.02fF
C18818 OR2X1_LOC_689/a_8_216# OR2X1_LOC_31/Y 0.09fF
C20986 OR2X1_LOC_433/a_8_216# OR2X1_LOC_31/Y 0.19fF
C23963 OR2X1_LOC_31/Y AND2X1_LOC_264/a_8_24# 0.01fF
C24343 OR2X1_LOC_689/a_36_216# OR2X1_LOC_31/Y 0.03fF
C24817 OR2X1_LOC_31/Y OR2X1_LOC_44/a_8_216# 0.01fF
C24885 OR2X1_LOC_31/Y OR2X1_LOC_511/a_8_216# 0.07fF
C25624 OR2X1_LOC_31/Y OR2X1_LOC_22/a_8_216# 0.01fF
C28177 OR2X1_LOC_272/a_8_216# OR2X1_LOC_31/Y 0.07fF
C30308 OR2X1_LOC_412/a_8_216# OR2X1_LOC_31/Y 0.01fF
C30345 OR2X1_LOC_31/Y AND2X1_LOC_687/a_8_24# 0.01fF
C31844 OR2X1_LOC_328/a_8_216# OR2X1_LOC_31/Y 0.01fF
C32186 OR2X1_LOC_31/Y OR2X1_LOC_323/a_8_216# 0.01fF
C32677 OR2X1_LOC_681/a_8_216# OR2X1_LOC_31/Y 0.18fF
C34413 OR2X1_LOC_31/Y OR2X1_LOC_40/a_8_216# 0.01fF
C36931 AND2X1_LOC_375/a_8_24# OR2X1_LOC_31/Y 0.08fF
C39113 OR2X1_LOC_694/a_8_216# OR2X1_LOC_31/Y 0.01fF
C43447 OR2X1_LOC_3/a_8_216# OR2X1_LOC_31/Y 0.01fF
C47630 OR2X1_LOC_31/Y OR2X1_LOC_386/a_8_216# 0.01fF
C48107 OR2X1_LOC_31/Y OR2X1_LOC_56/a_8_216# 0.14fF
C50850 OR2X1_LOC_275/a_8_216# OR2X1_LOC_31/Y 0.09fF
C54432 OR2X1_LOC_31/Y OR2X1_LOC_18/a_8_216# 0.10fF
C414 AND2X1_LOC_100/a_8_24# OR2X1_LOC_18/Y 0.03fF
C2605 OR2X1_LOC_18/Y OR2X1_LOC_86/a_8_216# 0.01fF
C5506 OR2X1_LOC_272/a_8_216# OR2X1_LOC_18/Y 0.10fF
C5994 OR2X1_LOC_18/Y OR2X1_LOC_226/a_8_216# 0.09fF
C10971 OR2X1_LOC_18/Y OR2X1_LOC_763/a_8_216# 0.01fF
C11033 OR2X1_LOC_18/Y OR2X1_LOC_95/a_8_216# 0.02fF
C12631 AND2X1_LOC_596/a_8_24# OR2X1_LOC_18/Y 0.02fF
C12906 OR2X1_LOC_18/Y OR2X1_LOC_85/a_8_216# 0.03fF
C15740 OR2X1_LOC_18/Y OR2X1_LOC_762/a_8_216# 0.04fF
C16547 OR2X1_LOC_18/Y OR2X1_LOC_95/a_36_216# 0.02fF
C17082 OR2X1_LOC_18/Y OR2X1_LOC_226/a_36_216# 0.03fF
C26814 OR2X1_LOC_18/Y OR2X1_LOC_762/a_36_216# 0.02fF
C27272 OR2X1_LOC_263/a_8_216# OR2X1_LOC_18/Y 0.01fF
C27998 OR2X1_LOC_18/Y OR2X1_LOC_71/a_8_216# 0.01fF
C31652 OR2X1_LOC_18/Y OR2X1_LOC_18/a_8_216# 0.01fF
C32211 OR2X1_LOC_18/Y AND2X1_LOC_458/a_8_24# 0.02fF
C32708 AND2X1_LOC_120/a_8_24# OR2X1_LOC_18/Y 0.02fF
C36814 OR2X1_LOC_18/Y OR2X1_LOC_63/a_8_216# 0.01fF
C36840 OR2X1_LOC_271/a_8_216# OR2X1_LOC_18/Y 0.01fF
C37820 OR2X1_LOC_18/Y OR2X1_LOC_289/a_8_216# 0.06fF
C40440 OR2X1_LOC_18/Y OR2X1_LOC_164/a_8_216# 0.07fF
C42056 OR2X1_LOC_488/a_8_216# OR2X1_LOC_18/Y 0.13fF
C42101 OR2X1_LOC_18/Y AND2X1_LOC_270/a_8_24# 0.05fF
C43328 OR2X1_LOC_18/Y OR2X1_LOC_371/a_8_216# 0.01fF
C47573 OR2X1_LOC_693/a_8_216# OR2X1_LOC_18/Y 0.04fF
C48095 OR2X1_LOC_692/a_8_216# OR2X1_LOC_18/Y 0.02fF
C48184 OR2X1_LOC_271/Y OR2X1_LOC_18/Y 0.26fF
C48845 OR2X1_LOC_527/a_8_216# OR2X1_LOC_18/Y 0.01fF
C49713 OR2X1_LOC_18/Y AND2X1_LOC_606/a_8_24# 0.01fF
C52461 OR2X1_LOC_18/Y OR2X1_LOC_92/a_8_216# 0.01fF
C55816 AND2X1_LOC_327/a_8_24# OR2X1_LOC_18/Y 0.09fF
C6629 OR2X1_LOC_23/a_8_216# OR2X1_LOC_59/Y -0.00fF
C11891 AND2X1_LOC_120/a_8_24# OR2X1_LOC_59/Y 0.03fF
C17067 OR2X1_LOC_289/a_8_216# OR2X1_LOC_59/Y 0.06fF
C20554 OR2X1_LOC_59/Y OR2X1_LOC_153/a_8_216# 0.02fF
C21084 OR2X1_LOC_129/a_8_216# OR2X1_LOC_59/Y 0.14fF
C23104 OR2X1_LOC_59/Y AND2X1_LOC_405/a_8_24# 0.02fF
C24053 OR2X1_LOC_59/Y OR2X1_LOC_585/a_8_216# 0.40fF
C26021 OR2X1_LOC_59/Y OR2X1_LOC_153/a_36_216# 0.02fF
C28148 OR2X1_LOC_59/Y OR2X1_LOC_534/a_8_216# 0.01fF
C34781 AND2X1_LOC_327/a_8_24# OR2X1_LOC_59/Y 0.01fF
C34874 OR2X1_LOC_59/Y OR2X1_LOC_29/a_8_216# 0.01fF
C35615 OR2X1_LOC_277/a_8_216# OR2X1_LOC_59/Y 0.14fF
C40661 OR2X1_LOC_272/a_8_216# OR2X1_LOC_59/Y 0.01fF
C41504 OR2X1_LOC_283/a_8_216# OR2X1_LOC_59/Y 0.01fF
C47441 OR2X1_LOC_59/Y OR2X1_LOC_300/a_8_216# 0.01fF
C48034 AND2X1_LOC_185/a_8_24# OR2X1_LOC_59/Y 0.02fF
C49176 OR2X1_LOC_304/a_8_216# OR2X1_LOC_59/Y 0.01fF
C3566 OR2X1_LOC_144/a_8_216# OR2X1_LOC_12/Y 0.06fF
C8363 OR2X1_LOC_763/a_8_216# OR2X1_LOC_12/Y 0.01fF
C9194 OR2X1_LOC_683/a_8_216# OR2X1_LOC_12/Y 0.01fF
C9692 AND2X1_LOC_264/a_36_24# OR2X1_LOC_12/Y 0.01fF
C9996 AND2X1_LOC_596/a_8_24# OR2X1_LOC_12/Y 0.18fF
C13157 OR2X1_LOC_762/a_8_216# OR2X1_LOC_12/Y 0.19fF
C13872 OR2X1_LOC_422/a_8_216# OR2X1_LOC_12/Y 0.04fF
C17756 OR2X1_LOC_684/Y OR2X1_LOC_12/Y 0.39fF
C19389 OR2X1_LOC_422/a_36_216# OR2X1_LOC_12/Y 0.02fF
C22478 AND2X1_LOC_294/a_8_24# OR2X1_LOC_12/Y 0.04fF
C24841 OR2X1_LOC_12/Y OR2X1_LOC_381/a_8_216# 0.06fF
C25771 OR2X1_LOC_699/a_8_216# OR2X1_LOC_12/Y 0.01fF
C28809 AND2X1_LOC_686/a_8_24# OR2X1_LOC_12/Y 0.01fF
C33408 AND2X1_LOC_294/a_36_24# OR2X1_LOC_12/Y 0.01fF
C35080 OR2X1_LOC_299/a_8_216# OR2X1_LOC_12/Y 0.01fF
C35814 AND2X1_LOC_410/a_8_24# OR2X1_LOC_12/Y 0.02fF
C35818 OR2X1_LOC_684/a_8_216# OR2X1_LOC_12/Y 0.01fF
C41386 OR2X1_LOC_625/a_8_216# OR2X1_LOC_12/Y 0.04fF
C49883 OR2X1_LOC_419/a_8_216# OR2X1_LOC_12/Y 0.01fF
C50107 OR2X1_LOC_306/a_8_216# OR2X1_LOC_12/Y 0.15fF
C51822 OR2X1_LOC_820/B OR2X1_LOC_12/Y 0.04fF
C54750 AND2X1_LOC_264/a_8_24# OR2X1_LOC_12/Y 0.04fF
C40729 OR2X1_LOC_753/a_8_216# OR2X1_LOC_753/Y 0.01fF
C5406 AND2X1_LOC_743/a_8_24# OR2X1_LOC_707/B 0.03fF
C8823 AND2X1_LOC_59/Y AND2X1_LOC_300/a_8_24# 0.03fF
C11327 AND2X1_LOC_59/Y AND2X1_LOC_534/a_8_24# 0.03fF
C15773 AND2X1_LOC_59/Y AND2X1_LOC_519/a_8_24# 0.01fF
C16272 AND2X1_LOC_59/Y AND2X1_LOC_271/a_8_24# 0.17fF
C16839 AND2X1_LOC_59/Y AND2X1_LOC_255/a_8_24# 0.01fF
C22047 AND2X1_LOC_59/Y AND2X1_LOC_387/a_8_24# 0.01fF
C22446 AND2X1_LOC_59/Y AND2X1_LOC_534/a_36_24# 0.01fF
C28947 AND2X1_LOC_59/Y OR2X1_LOC_750/a_8_216# 0.06fF
C32890 AND2X1_LOC_59/Y OR2X1_LOC_120/a_8_216# 0.01fF
C35989 AND2X1_LOC_59/Y AND2X1_LOC_328/a_8_24# 0.20fF
C39370 AND2X1_LOC_59/Y OR2X1_LOC_274/a_8_216# 0.01fF
C46506 AND2X1_LOC_59/Y OR2X1_LOC_276/B 0.09fF
C47962 AND2X1_LOC_59/Y AND2X1_LOC_273/a_8_24# 0.01fF
C49292 AND2X1_LOC_371/a_8_24# AND2X1_LOC_59/Y 0.03fF
C3721 AND2X1_LOC_12/Y AND2X1_LOC_625/a_8_24# 0.02fF
C4771 AND2X1_LOC_12/Y AND2X1_LOC_225/a_8_24# 0.01fF
C5962 AND2X1_LOC_12/Y AND2X1_LOC_425/a_8_24# 0.01fF
C7871 AND2X1_LOC_12/Y AND2X1_LOC_581/a_8_24# 0.01fF
C12341 AND2X1_LOC_12/Y AND2X1_LOC_382/a_8_24# 0.01fF
C17420 AND2X1_LOC_12/Y OR2X1_LOC_68/a_8_216# 0.01fF
C19960 AND2X1_LOC_12/Y AND2X1_LOC_421/a_8_24# 0.02fF
C21194 AND2X1_LOC_12/Y AND2X1_LOC_310/a_8_24# 0.01fF
C21393 AND2X1_LOC_12/Y AND2X1_LOC_692/a_8_24# 0.02fF
C21863 AND2X1_LOC_12/Y AND2X1_LOC_761/a_8_24# 0.01fF
C23839 AND2X1_LOC_12/Y AND2X1_LOC_381/a_8_24# 0.01fF
C24759 AND2X1_LOC_12/Y AND2X1_LOC_309/a_8_24# 0.02fF
C27164 AND2X1_LOC_12/Y AND2X1_LOC_422/a_8_24# 0.03fF
C28539 AND2X1_LOC_12/Y AND2X1_LOC_283/a_8_24# 0.01fF
C29585 AND2X1_LOC_12/Y AND2X1_LOC_299/a_8_24# 0.09fF
C30814 AND2X1_LOC_12/Y AND2X1_LOC_599/a_8_24# 0.01fF
C30999 AND2X1_LOC_12/Y AND2X1_LOC_369/a_8_24# 0.02fF
C31934 AND2X1_LOC_12/Y AND2X1_LOC_699/a_8_24# 0.01fF
C32321 AND2X1_LOC_12/Y AND2X1_LOC_289/a_8_24# 0.01fF
C40416 AND2X1_LOC_12/Y AND2X1_LOC_429/a_8_24# 0.20fF
C42381 AND2X1_LOC_12/Y AND2X1_LOC_3/a_8_24# 0.01fF
C42633 AND2X1_LOC_12/Y AND2X1_LOC_236/a_8_24# 0.01fF
C45041 AND2X1_LOC_12/Y AND2X1_LOC_153/a_8_24# 0.01fF
C45076 AND2X1_LOC_12/Y OR2X1_LOC_296/a_8_216# 0.03fF
C45487 AND2X1_LOC_12/Y AND2X1_LOC_817/a_8_24# 0.01fF
C46041 AND2X1_LOC_12/Y OR2X1_LOC_276/B 0.09fF
C48513 AND2X1_LOC_12/Y AND2X1_LOC_628/a_8_24# 0.02fF
C49265 AND2X1_LOC_12/Y AND2X1_LOC_275/a_8_24# 0.02fF
C49569 AND2X1_LOC_12/Y OR2X1_LOC_512/a_8_216# 0.01fF
C51623 AND2X1_LOC_12/Y OR2X1_LOC_276/a_8_216# 0.02fF
C51675 AND2X1_LOC_12/Y OR2X1_LOC_513/a_8_216# 0.01fF
C53248 AND2X1_LOC_12/Y AND2X1_LOC_136/a_8_24# 0.01fF
C53640 AND2X1_LOC_12/Y OR2X1_LOC_847/a_8_216# 0.01fF
C1549 AND2X1_LOC_95/Y OR2X1_LOC_185/a_8_216# 0.01fF
C2710 AND2X1_LOC_95/Y AND2X1_LOC_289/a_8_24# 0.01fF
C7042 AND2X1_LOC_95/Y OR2X1_LOC_185/a_36_216# 0.02fF
C9633 AND2X1_LOC_92/a_8_24# AND2X1_LOC_95/Y 0.17fF
C16236 AND2X1_LOC_95/Y OR2X1_LOC_276/B 0.01fF
C19135 AND2X1_LOC_95/Y AND2X1_LOC_413/a_8_24# 0.17fF
C23333 AND2X1_LOC_95/Y OR2X1_LOC_410/a_8_216# 0.01fF
C27122 AND2X1_LOC_95/Y AND2X1_LOC_71/a_8_24# 0.01fF
C28765 AND2X1_LOC_95/Y OR2X1_LOC_410/a_36_216# -0.00fF
C31782 AND2X1_LOC_95/Y OR2X1_LOC_407/a_8_216# 0.02fF
C33919 AND2X1_LOC_95/Y AND2X1_LOC_233/a_8_24# 0.01fF
C34203 AND2X1_LOC_95/Y AND2X1_LOC_322/a_8_24# 0.02fF
C37126 AND2X1_LOC_95/Y AND2X1_LOC_534/a_8_24# 0.04fF
C41139 AND2X1_LOC_95/Y AND2X1_LOC_159/a_8_24# 0.01fF
C42398 AND2X1_LOC_95/Y AND2X1_LOC_57/a_8_24# 0.07fF
C42762 AND2X1_LOC_95/Y AND2X1_LOC_323/a_8_24# 0.07fF
C49714 AND2X1_LOC_95/Y AND2X1_LOC_411/a_8_24# 0.13fF
C51159 AND2X1_LOC_95/Y AND2X1_LOC_309/a_8_24# 0.02fF
C25820 OR2X1_LOC_448/B AND2X1_LOC_422/a_8_24# 0.21fF
C5833 AND2X1_LOC_66/a_36_24# OR2X1_LOC_26/Y 0.01fF
C9491 OR2X1_LOC_26/Y OR2X1_LOC_43/a_8_216# 0.06fF
C9513 AND2X1_LOC_66/a_8_24# OR2X1_LOC_26/Y 0.17fF
C9935 OR2X1_LOC_80/a_8_216# OR2X1_LOC_26/Y 0.01fF
C11149 OR2X1_LOC_26/Y OR2X1_LOC_245/a_8_216# 0.11fF
C11336 OR2X1_LOC_26/Y OR2X1_LOC_373/a_8_216# 0.04fF
C13272 OR2X1_LOC_26/Y OR2X1_LOC_6/a_8_216# 0.01fF
C17592 OR2X1_LOC_26/Y OR2X1_LOC_164/a_8_216# 0.01fF
C18293 OR2X1_LOC_529/a_8_216# OR2X1_LOC_26/Y 0.01fF
C19045 OR2X1_LOC_129/a_8_216# OR2X1_LOC_26/Y 0.01fF
C20028 AND2X1_LOC_87/a_8_24# OR2X1_LOC_26/Y 0.01fF
C20930 OR2X1_LOC_696/a_8_216# OR2X1_LOC_26/Y 0.03fF
C21011 OR2X1_LOC_26/Y AND2X1_LOC_405/a_8_24# 0.01fF
C22026 OR2X1_LOC_26/Y OR2X1_LOC_585/a_8_216# 0.04fF
C22580 AND2X1_LOC_374/a_8_24# OR2X1_LOC_26/Y 0.05fF
C34294 AND2X1_LOC_513/a_8_24# OR2X1_LOC_26/Y 0.01fF
C34842 OR2X1_LOC_26/Y OR2X1_LOC_93/a_8_216# 0.07fF
C38706 OR2X1_LOC_26/Y OR2X1_LOC_64/a_8_216# 0.39fF
C39482 OR2X1_LOC_283/a_8_216# OR2X1_LOC_26/Y 0.03fF
C44208 OR2X1_LOC_26/Y OR2X1_LOC_95/a_8_216# 0.01fF
C44609 AND2X1_LOC_374/a_36_24# OR2X1_LOC_26/Y 0.01fF
C47158 OR2X1_LOC_490/a_8_216# OR2X1_LOC_26/Y 0.03fF
C51052 OR2X1_LOC_26/Y OR2X1_LOC_26/a_8_216# -0.00fF
C52664 OR2X1_LOC_490/a_36_216# OR2X1_LOC_26/Y 0.02fF
C891 AND2X1_LOC_512/a_8_24# OR2X1_LOC_36/Y 0.03fF
C3599 OR2X1_LOC_36/Y OR2X1_LOC_88/a_8_216# 0.02fF
C3616 OR2X1_LOC_36/Y OR2X1_LOC_378/A 0.07fF
C4660 AND2X1_LOC_502/a_36_24# OR2X1_LOC_36/Y 0.01fF
C7498 OR2X1_LOC_304/a_8_216# OR2X1_LOC_36/Y 0.01fF
C8812 OR2X1_LOC_36/Y OR2X1_LOC_310/a_8_216# 0.04fF
C9533 OR2X1_LOC_36/Y OR2X1_LOC_619/a_8_216# 0.03fF
C9765 AND2X1_LOC_377/Y OR2X1_LOC_36/Y 0.08fF
C11477 OR2X1_LOC_291/a_8_216# OR2X1_LOC_36/Y 0.10fF
C15293 OR2X1_LOC_36/Y OR2X1_LOC_48/a_8_216# 0.01fF
C18514 OR2X1_LOC_36/Y OR2X1_LOC_268/Y 0.60fF
C18958 OR2X1_LOC_36/Y OR2X1_LOC_56/a_8_216# 0.01fF
C21262 OR2X1_LOC_36/Y OR2X1_LOC_23/a_8_216# -0.00fF
C22593 OR2X1_LOC_291/a_36_216# OR2X1_LOC_36/Y 0.03fF
C23072 AND2X1_LOC_512/a_36_24# OR2X1_LOC_36/Y 0.01fF
C24378 OR2X1_LOC_36/Y OR2X1_LOC_587/a_8_216# 0.43fF
C28902 OR2X1_LOC_682/a_8_216# OR2X1_LOC_36/Y 0.18fF
C29253 OR2X1_LOC_689/A OR2X1_LOC_36/Y 0.03fF
C29523 OR2X1_LOC_36/Y AND2X1_LOC_269/a_8_24# 0.01fF
C30571 OR2X1_LOC_271/a_8_216# OR2X1_LOC_36/Y 0.01fF
C34853 OR2X1_LOC_824/a_8_216# OR2X1_LOC_36/Y 0.09fF
C35730 OR2X1_LOC_36/Y AND2X1_LOC_270/a_8_24# 0.15fF
C37347 OR2X1_LOC_696/a_8_216# OR2X1_LOC_36/Y 0.01fF
C38785 OR2X1_LOC_36/Y OR2X1_LOC_599/a_8_216# 0.09fF
C40984 OR2X1_LOC_693/a_8_216# OR2X1_LOC_36/Y 0.08fF
C41614 OR2X1_LOC_271/Y OR2X1_LOC_36/Y 0.01fF
C43203 OR2X1_LOC_36/Y AND2X1_LOC_606/a_8_24# 0.04fF
C43797 OR2X1_LOC_36/Y AND2X1_LOC_688/a_8_24# 0.02fF
C44183 AND2X1_LOC_502/a_8_24# OR2X1_LOC_36/Y 0.04fF
C44382 OR2X1_LOC_36/Y OR2X1_LOC_599/a_36_216# 0.03fF
C46077 OR2X1_LOC_36/Y OR2X1_LOC_419/a_8_216# 0.07fF
C48205 OR2X1_LOC_433/a_8_216# OR2X1_LOC_36/Y 0.01fF
C49575 OR2X1_LOC_36/Y OR2X1_LOC_29/a_8_216# 0.01fF
C49915 OR2X1_LOC_273/a_8_216# OR2X1_LOC_36/Y 0.03fF
C50086 OR2X1_LOC_110/a_8_216# OR2X1_LOC_36/Y 0.01fF
C50377 OR2X1_LOC_36/Y OR2X1_LOC_268/a_8_216# 0.01fF
C51058 AND2X1_LOC_513/a_8_24# OR2X1_LOC_36/Y 0.03fF
C52064 OR2X1_LOC_36/Y OR2X1_LOC_511/a_8_216# 0.01fF
C54360 OR2X1_LOC_36/Y AND2X1_LOC_606/a_36_24# 0.01fF
C55388 OR2X1_LOC_273/a_36_216# OR2X1_LOC_36/Y 0.03fF
C131 OR2X1_LOC_22/Y AND2X1_LOC_293/a_8_24# 0.03fF
C949 OR2X1_LOC_433/a_8_216# OR2X1_LOC_22/Y 0.01fF
C1489 OR2X1_LOC_22/Y AND2X1_LOC_461/a_8_24# 0.05fF
C3950 OR2X1_LOC_22/Y AND2X1_LOC_264/a_8_24# 0.03fF
C8710 OR2X1_LOC_22/Y OR2X1_LOC_226/a_8_216# 0.02fF
C9929 AND2X1_LOC_512/a_8_24# OR2X1_LOC_22/Y 0.01fF
C10379 OR2X1_LOC_22/Y OR2X1_LOC_412/a_8_216# 0.04fF
C13722 OR2X1_LOC_22/Y OR2X1_LOC_95/a_8_216# 0.01fF
C14527 OR2X1_LOC_22/Y OR2X1_LOC_40/a_8_216# 0.40fF
C17046 OR2X1_LOC_22/Y AND2X1_LOC_276/a_8_24# 0.01fF
C18044 OR2X1_LOC_22/Y AND2X1_LOC_461/a_36_24# 0.01fF
C19637 OR2X1_LOC_22/Y OR2X1_LOC_59/a_8_216# 0.01fF
C27571 OR2X1_LOC_309/a_8_216# OR2X1_LOC_22/Y 0.07fF
C29865 OR2X1_LOC_22/Y OR2X1_LOC_263/a_8_216# 0.01fF
C30108 OR2X1_LOC_329/a_8_216# OR2X1_LOC_22/Y 0.02fF
C30674 OR2X1_LOC_22/Y OR2X1_LOC_275/a_8_216# 0.05fF
C34934 OR2X1_LOC_22/Y OR2X1_LOC_43/a_8_216# 0.03fF
C36577 OR2X1_LOC_22/Y OR2X1_LOC_245/a_8_216# 0.02fF
C38212 OR2X1_LOC_22/Y AND2X1_LOC_274/a_8_24# 0.01fF
C40408 OR2X1_LOC_22/Y OR2X1_LOC_43/a_36_216# 0.03fF
C41096 OR2X1_LOC_329/a_36_216# OR2X1_LOC_22/Y 0.02fF
C42155 OR2X1_LOC_22/Y OR2X1_LOC_245/a_36_216# 0.02fF
C43979 OR2X1_LOC_22/Y OR2X1_LOC_153/a_8_216# 0.03fF
C47670 OR2X1_LOC_22/Y OR2X1_LOC_585/a_8_216# 0.01fF
C47988 OR2X1_LOC_22/Y OR2X1_LOC_599/a_8_216# 0.05fF
C50797 OR2X1_LOC_271/Y OR2X1_LOC_22/Y 0.02fF
C53277 AND2X1_LOC_502/a_8_24# OR2X1_LOC_22/Y 0.02fF
C55397 OR2X1_LOC_306/a_8_216# OR2X1_LOC_22/Y 0.01fF
C594 OR2X1_LOC_378/Y OR2X1_LOC_378/A 0.01fF
C22148 OR2X1_LOC_376/Y OR2X1_LOC_378/A 0.88fF
C40162 OR2X1_LOC_377/a_8_216# OR2X1_LOC_378/A 0.01fF
C51288 OR2X1_LOC_3/Y OR2X1_LOC_378/A 0.05fF
C56299 OR2X1_LOC_378/A VSS 0.02fF
C9038 OR2X1_LOC_709/A AND2X1_LOC_419/a_8_24# 0.02fF
C19754 OR2X1_LOC_709/A OR2X1_LOC_514/a_8_216# 0.01fF
C24997 OR2X1_LOC_709/A AND2X1_LOC_136/a_8_24# 0.21fF
C25591 OR2X1_LOC_709/A AND2X1_LOC_419/a_36_24# -0.01fF
C27447 OR2X1_LOC_709/A AND2X1_LOC_748/a_8_24# 0.03fF
C38408 OR2X1_LOC_709/A AND2X1_LOC_748/a_36_24# 0.01fF
C39548 OR2X1_LOC_709/A OR2X1_LOC_515/a_8_216# 0.01fF
C48213 AND2X1_LOC_692/a_8_24# OR2X1_LOC_706/A 0.01fF
C39516 AND2X1_LOC_458/a_8_24# OR2X1_LOC_371/Y 0.04fF
C55864 OR2X1_LOC_371/Y OR2X1_LOC_372/a_8_216# 0.43fF
C56113 OR2X1_LOC_527/a_8_216# OR2X1_LOC_371/Y 0.01fF
C11623 OR2X1_LOC_488/a_8_216# OR2X1_LOC_71/Y 0.01fF
C17144 OR2X1_LOC_488/a_36_216# OR2X1_LOC_71/Y -0.00fF
C20092 AND2X1_LOC_502/a_8_24# OR2X1_LOC_71/Y 0.01fF
C18388 AND2X1_LOC_68/a_8_24# OR2X1_LOC_69/A 0.01fF
C13055 OR2X1_LOC_327/a_8_216# AND2X1_LOC_65/A 0.01fF
C45787 OR2X1_LOC_264/a_8_216# AND2X1_LOC_65/A 0.05fF
C199 AND2X1_LOC_548/a_8_24# OR2X1_LOC_437/A 0.03fF
C4454 OR2X1_LOC_372/a_36_216# OR2X1_LOC_437/A 0.15fF
C12839 OR2X1_LOC_136/a_8_216# OR2X1_LOC_437/A 0.03fF
C13337 OR2X1_LOC_369/a_8_216# OR2X1_LOC_437/A 0.03fF
C14738 OR2X1_LOC_255/a_8_216# OR2X1_LOC_437/A 0.03fF
C16221 OR2X1_LOC_437/A OR2X1_LOC_310/a_8_216# 0.03fF
C20965 OR2X1_LOC_530/a_8_216# OR2X1_LOC_437/A 0.05fF
C22751 AND2X1_LOC_514/a_8_24# OR2X1_LOC_437/A 0.04fF
C25761 OR2X1_LOC_255/a_36_216# OR2X1_LOC_437/A 0.01fF
C26020 OR2X1_LOC_309/a_8_216# OR2X1_LOC_437/A -0.01fF
C26135 AND2X1_LOC_294/a_8_24# OR2X1_LOC_437/A 0.04fF
C31711 OR2X1_LOC_10/a_8_216# OR2X1_LOC_437/A 0.41fF
C31958 OR2X1_LOC_256/a_8_216# OR2X1_LOC_437/A -0.06fF
C34100 OR2X1_LOC_519/a_8_216# OR2X1_LOC_437/A 0.03fF
C38241 OR2X1_LOC_437/A OR2X1_LOC_322/a_8_216# 0.15fF
C39174 AND2X1_LOC_514/a_36_24# OR2X1_LOC_437/A 0.01fF
C39552 OR2X1_LOC_102/a_8_216# OR2X1_LOC_437/A 0.03fF
C49542 OR2X1_LOC_437/A OR2X1_LOC_322/a_36_216# 0.14fF
C49663 OR2X1_LOC_372/a_8_216# OR2X1_LOC_437/A 0.18fF
C5197 AND2X1_LOC_100/a_8_24# OR2X1_LOC_86/A 0.05fF
C7386 OR2X1_LOC_86/A OR2X1_LOC_86/a_8_216# 0.01fF
C3989 OR2X1_LOC_245/a_8_216# OR2X1_LOC_246/A 0.01fF
C9544 OR2X1_LOC_245/a_36_216# OR2X1_LOC_246/A 0.07fF
C22703 OR2X1_LOC_246/A OR2X1_LOC_246/a_8_216# 0.09fF
C26031 OR2X1_LOC_273/a_8_216# OR2X1_LOC_246/A 0.13fF
C28558 OR2X1_LOC_246/A OR2X1_LOC_86/a_8_216# 0.05fF
C31529 OR2X1_LOC_273/a_36_216# OR2X1_LOC_246/A 0.13fF
C37617 OR2X1_LOC_136/a_8_216# OR2X1_LOC_246/A 0.12fF
C53348 OR2X1_LOC_263/a_8_216# OR2X1_LOC_246/A 0.05fF
C3977 OR2X1_LOC_277/a_36_216# OR2X1_LOC_278/A 0.01fF
C10327 OR2X1_LOC_126/a_8_216# OR2X1_LOC_278/A 0.40fF
C13345 OR2X1_LOC_119/a_8_216# OR2X1_LOC_278/A 0.03fF
C15743 OR2X1_LOC_291/a_8_216# OR2X1_LOC_278/A 0.01fF
C54589 OR2X1_LOC_277/a_8_216# OR2X1_LOC_278/A 0.01fF
C30314 OR2X1_LOC_255/a_8_216# OR2X1_LOC_256/A 0.01fF
C47809 OR2X1_LOC_256/A OR2X1_LOC_256/a_8_216# 0.08fF
C1856 AND2X1_LOC_461/a_36_24# OR2X1_LOC_690/A 0.02fF
C8060 AND2X1_LOC_378/a_8_24# OR2X1_LOC_690/A 0.08fF
C20791 AND2X1_LOC_691/a_8_24# OR2X1_LOC_690/A 0.02fF
C22151 OR2X1_LOC_689/A OR2X1_LOC_690/A 0.03fF
C35217 OR2X1_LOC_690/a_8_216# OR2X1_LOC_690/A 0.01fF
C38557 OR2X1_LOC_689/a_8_216# OR2X1_LOC_690/A 0.01fF
C39960 AND2X1_LOC_293/a_8_24# OR2X1_LOC_690/A 0.18fF
C41278 AND2X1_LOC_461/a_8_24# OR2X1_LOC_690/A 0.16fF
C50396 OR2X1_LOC_412/a_8_216# OR2X1_LOC_690/A 0.02fF
C56211 OR2X1_LOC_413/a_8_216# OR2X1_LOC_690/A 0.02fF
C2231 OR2X1_LOC_813/A OR2X1_LOC_71/a_8_216# 0.41fF
C18376 AND2X1_LOC_619/a_8_24# OR2X1_LOC_622/B 0.01fF
C17898 OR2X1_LOC_672/Y OR2X1_LOC_73/a_8_216# 0.45fF
C51673 AND2X1_LOC_159/a_8_24# AND2X1_LOC_72/B 0.01fF
C9792 OR2X1_LOC_63/a_8_216# OR2X1_LOC_65/B 0.02fF
C15684 AND2X1_LOC_87/a_8_24# OR2X1_LOC_65/B 0.17fF
C22464 OR2X1_LOC_65/B AND2X1_LOC_606/a_8_24# 0.23fF
C28511 AND2X1_LOC_327/a_8_24# OR2X1_LOC_65/B -0.00fF
C38736 OR2X1_LOC_65/B OR2X1_LOC_88/a_8_216# 0.01fF
C32544 OR2X1_LOC_458/a_8_216# OR2X1_LOC_464/A -0.00fF
C9621 OR2X1_LOC_273/a_8_216# OR2X1_LOC_300/Y 0.39fF
C21727 OR2X1_LOC_300/a_8_216# OR2X1_LOC_300/Y 0.01fF
C35338 AND2X1_LOC_433/a_8_24# OR2X1_LOC_435/A 0.09fF
C12099 AND2X1_LOC_372/a_36_24# OR2X1_LOC_831/B 0.01fF
C29098 AND2X1_LOC_153/a_8_24# OR2X1_LOC_831/B 0.03fF
C31523 AND2X1_LOC_273/a_8_24# OR2X1_LOC_831/B 0.01fF
C45734 AND2X1_LOC_153/a_36_24# OR2X1_LOC_831/B 0.01fF
C46128 AND2X1_LOC_372/a_8_24# OR2X1_LOC_831/B 0.05fF
C48727 AND2X1_LOC_300/a_8_24# OR2X1_LOC_831/B 0.20fF
C53780 OR2X1_LOC_831/B AND2X1_LOC_273/a_36_24# 0.01fF
C17739 AND2X1_LOC_763/a_8_24# OR2X1_LOC_828/B 0.01fF
C8585 OR2X1_LOC_685/B OR2X1_LOC_685/a_8_216# 0.07fF
C16121 OR2X1_LOC_685/B OR2X1_LOC_161/A 0.01fF
C16208 OR2X1_LOC_685/B AND2X1_LOC_51/Y 0.01fF
C23289 OR2X1_LOC_685/B OR2X1_LOC_161/B 0.17fF
C36464 OR2X1_LOC_687/Y OR2X1_LOC_685/B 0.03fF
C42825 OR2X1_LOC_685/B OR2X1_LOC_78/B 0.11fF
C47323 OR2X1_LOC_685/B OR2X1_LOC_87/A 0.01fF
C55642 VDD OR2X1_LOC_685/B 0.21fF
C57713 OR2X1_LOC_685/B VSS 0.11fF
C14033 AND2X1_LOC_743/a_8_24# OR2X1_LOC_780/B 0.01fF
C34128 OR2X1_LOC_155/a_8_216# OR2X1_LOC_156/A 0.01fF
C29817 OR2X1_LOC_502/a_8_216# OR2X1_LOC_502/Y 0.05fF
C40736 AND2X1_LOC_696/a_8_24# OR2X1_LOC_708/B 0.01fF
C36788 OR2X1_LOC_818/Y AND2X1_LOC_820/a_8_24# 0.23fF
C38880 VDD OR2X1_LOC_818/Y 0.12fF
C40141 OR2X1_LOC_818/Y AND2X1_LOC_820/B 0.08fF
C57178 OR2X1_LOC_818/Y VSS 0.06fF
C42301 AND2X1_LOC_144/a_8_24# OR2X1_LOC_147/A 0.01fF
C13480 AND2X1_LOC_164/a_8_24# OR2X1_LOC_168/B 0.01fF
C3233 AND2X1_LOC_322/a_8_24# OR2X1_LOC_325/B 0.01fF
C16167 AND2X1_LOC_376/a_8_24# OR2X1_LOC_459/B 0.02fF
C46552 OR2X1_LOC_638/B AND2X1_LOC_408/a_8_24# 0.20fF
C8550 OR2X1_LOC_416/A AND2X1_LOC_415/a_8_24# 0.01fF
C15814 OR2X1_LOC_416/A OR2X1_LOC_49/a_8_216# 0.47fF
C18371 OR2X1_LOC_481/A AND2X1_LOC_818/a_8_24# 0.01fF
C23921 OR2X1_LOC_481/A OR2X1_LOC_820/B 0.04fF
C28108 OR2X1_LOC_481/A OR2X1_LOC_236/a_8_216# 0.01fF
C31551 OR2X1_LOC_481/A OR2X1_LOC_55/a_8_216# 0.01fF
C9379 OR2X1_LOC_690/a_8_216# OR2X1_LOC_689/A -0.00fF
C10635 OR2X1_LOC_689/A AND2X1_LOC_688/a_8_24# 0.01fF
C20862 OR2X1_LOC_3/Y OR2X1_LOC_689/A 0.02fF
C32539 AND2X1_LOC_377/Y OR2X1_LOC_689/A 0.03fF
C38511 OR2X1_LOC_689/A OR2X1_LOC_39/A 0.02fF
C43648 OR2X1_LOC_459/A OR2X1_LOC_689/A 0.09fF
C57459 OR2X1_LOC_689/A VSS 0.35fF
C5060 OR2X1_LOC_625/Y AND2X1_LOC_294/a_8_24# 0.02fF
C38372 OR2X1_LOC_625/Y OR2X1_LOC_753/a_8_216# -0.02fF
C44000 OR2X1_LOC_625/Y OR2X1_LOC_753/a_36_216# 0.01fF
C44556 OR2X1_LOC_625/Y OR2X1_LOC_628/a_8_216# 0.08fF
C29875 AND2X1_LOC_692/a_8_24# OR2X1_LOC_706/B 0.01fF
C8233 AND2X1_LOC_306/a_8_24# OR2X1_LOC_779/B 0.01fF
C21171 OR2X1_LOC_512/a_8_216# OR2X1_LOC_779/B 0.01fF
C23344 OR2X1_LOC_779/B OR2X1_LOC_513/a_8_216# 0.05fF
C29841 AND2X1_LOC_304/a_8_24# OR2X1_LOC_779/B 0.20fF
C968 OR2X1_LOC_428/A OR2X1_LOC_268/Y 0.06fF
C6188 OR2X1_LOC_268/a_8_216# OR2X1_LOC_268/Y 0.01fF
C41273 VDD OR2X1_LOC_268/Y 0.07fF
C44289 OR2X1_LOC_45/B OR2X1_LOC_268/Y 0.54fF
C44735 OR2X1_LOC_158/A OR2X1_LOC_268/Y 0.03fF
C48728 OR2X1_LOC_56/A OR2X1_LOC_268/Y 0.03fF
C56407 OR2X1_LOC_268/Y VSS -0.13fF
C33118 AND2X1_LOC_185/a_8_24# OR2X1_LOC_628/Y 0.01fF
C3022 AND2X1_LOC_271/a_8_24# AND2X1_LOC_7/B 0.02fF
C3586 AND2X1_LOC_7/B AND2X1_LOC_255/a_8_24# 0.01fF
C14730 AND2X1_LOC_291/a_8_24# AND2X1_LOC_7/B 0.01fF
C15124 OR2X1_LOC_269/a_8_216# AND2X1_LOC_7/B 0.01fF
C19009 AND2X1_LOC_18/a_8_24# AND2X1_LOC_7/B 0.01fF
C19158 AND2X1_LOC_699/a_8_24# AND2X1_LOC_7/B 0.02fF
C19712 AND2X1_LOC_7/B OR2X1_LOC_120/a_8_216# 0.01fF
C20944 AND2X1_LOC_7/B AND2X1_LOC_268/a_8_24# 0.02fF
C24326 AND2X1_LOC_7/B AND2X1_LOC_419/a_8_24# 0.01fF
C26128 OR2X1_LOC_274/a_8_216# AND2X1_LOC_7/B 0.03fF
C31875 AND2X1_LOC_7/B OR2X1_LOC_269/A 0.15fF
C33048 OR2X1_LOC_276/B AND2X1_LOC_7/B 0.08fF
C34479 AND2X1_LOC_7/B AND2X1_LOC_256/a_8_24# 0.01fF
C34957 AND2X1_LOC_7/B OR2X1_LOC_514/a_8_216# 0.02fF
C37369 AND2X1_LOC_7/B AND2X1_LOC_268/a_36_24# 0.02fF
C39178 OR2X1_LOC_121/a_8_216# AND2X1_LOC_7/B 0.02fF
C40058 OR2X1_LOC_405/a_8_216# AND2X1_LOC_7/B 0.01fF
C40124 AND2X1_LOC_136/a_8_24# AND2X1_LOC_7/B 0.02fF
C40893 AND2X1_LOC_749/a_8_24# AND2X1_LOC_7/B 0.01fF
C54954 AND2X1_LOC_7/B OR2X1_LOC_515/a_8_216# 0.01fF
C12827 OR2X1_LOC_256/Y OR2X1_LOC_255/a_8_216# 0.48fF
C23909 OR2X1_LOC_256/Y OR2X1_LOC_255/a_36_216# 0.01fF
C24263 OR2X1_LOC_256/Y AND2X1_LOC_294/a_8_24# 0.01fF
C10088 OR2X1_LOC_756/B OR2X1_LOC_410/a_8_216# 0.03fF
C12121 OR2X1_LOC_756/B AND2X1_LOC_488/a_8_24# 0.01fF
C12496 OR2X1_LOC_756/B OR2X1_LOC_374/a_8_216# 0.01fF
C41631 OR2X1_LOC_756/B AND2X1_LOC_283/a_8_24# 0.02fF
C45583 OR2X1_LOC_756/B AND2X1_LOC_289/a_8_24# 0.01fF
C45892 OR2X1_LOC_756/B AND2X1_LOC_85/a_8_24# 0.20fF
C48061 OR2X1_LOC_756/B OR2X1_LOC_814/a_8_216# 0.03fF
C55269 OR2X1_LOC_756/B OR2X1_LOC_270/a_8_216# 0.04fF
C3766 OR2X1_LOC_160/B AND2X1_LOC_159/a_8_24# 0.03fF
C5227 OR2X1_LOC_160/B AND2X1_LOC_255/a_8_24# 0.01fF
C10234 OR2X1_LOC_160/B AND2X1_LOC_692/a_8_24# 0.05fF
C10463 OR2X1_LOC_160/B AND2X1_LOC_387/a_8_24# 0.01fF
C12764 OR2X1_LOC_160/B AND2X1_LOC_23/a_8_24# 0.01fF
C17405 OR2X1_LOC_160/B OR2X1_LOC_750/a_8_216# 0.01fF
C19380 OR2X1_LOC_160/B AND2X1_LOC_110/a_8_24# 0.01fF
C20350 OR2X1_LOC_160/B AND2X1_LOC_159/a_36_24# 0.01fF
C21375 OR2X1_LOC_160/B AND2X1_LOC_289/a_8_24# 0.04fF
C21480 OR2X1_LOC_160/B OR2X1_LOC_120/a_8_216# 0.01fF
C27363 AND2X1_LOC_743/a_8_24# OR2X1_LOC_160/B 0.01fF
C27856 OR2X1_LOC_160/B OR2X1_LOC_274/a_8_216# 0.03fF
C34824 OR2X1_LOC_160/B OR2X1_LOC_276/B 0.07fF
C34969 OR2X1_LOC_160/B AND2X1_LOC_226/a_8_24# 0.01fF
C37509 OR2X1_LOC_155/a_8_216# OR2X1_LOC_160/B 0.01fF
C40355 OR2X1_LOC_160/B OR2X1_LOC_513/a_8_216# 0.03fF
C43952 OR2X1_LOC_160/B AND2X1_LOC_488/a_8_24# 0.04fF
C42440 AND2X1_LOC_748/a_8_24# OR2X1_LOC_789/B 0.01fF
C33876 OR2X1_LOC_534/a_8_216# OR2X1_LOC_534/Y 0.01fF
C42519 OR2X1_LOC_527/a_8_216# OR2X1_LOC_419/Y 0.13fF
C44324 AND2X1_LOC_502/a_8_24# OR2X1_LOC_419/Y 0.07fF
C46197 OR2X1_LOC_419/a_8_216# OR2X1_LOC_419/Y 0.01fF
C48234 OR2X1_LOC_527/a_36_216# OR2X1_LOC_419/Y 0.15fF
C3104 OR2X1_LOC_272/a_8_216# OR2X1_LOC_272/Y 0.01fF
C33102 OR2X1_LOC_272/Y AND2X1_LOC_274/a_8_24# 0.09fF
C2099 OR2X1_LOC_459/A AND2X1_LOC_688/a_8_24# 0.20fF
C29578 AND2X1_LOC_378/a_8_24# OR2X1_LOC_459/A 0.01fF
C1232 OR2X1_LOC_684/Y OR2X1_LOC_16/A 0.39fF
C14452 OR2X1_LOC_604/A OR2X1_LOC_684/Y 0.02fF
C32794 OR2X1_LOC_684/Y AND2X1_LOC_686/a_8_24# 0.02fF
C36833 VDD OR2X1_LOC_684/Y 0.03fF
C38192 OR2X1_LOC_427/A OR2X1_LOC_684/Y 0.01fF
C39843 OR2X1_LOC_684/a_8_216# OR2X1_LOC_684/Y 0.04fF
C55884 OR2X1_LOC_70/Y OR2X1_LOC_684/Y 0.01fF
C57004 OR2X1_LOC_684/Y VSS 0.34fF
C15404 OR2X1_LOC_136/a_8_216# OR2X1_LOC_136/Y 0.01fF
C51424 AND2X1_LOC_820/a_8_24# AND2X1_LOC_820/B -0.00fF
C53481 VDD AND2X1_LOC_820/B 0.19fF
C56649 AND2X1_LOC_820/B VSS 0.05fF
C1224 OR2X1_LOC_42/a_8_216# OR2X1_LOC_56/A 0.04fF
C5413 OR2X1_LOC_299/a_8_216# OR2X1_LOC_56/A 0.01fF
C12125 OR2X1_LOC_672/a_8_216# OR2X1_LOC_56/A 0.02fF
C15635 OR2X1_LOC_271/Y OR2X1_LOC_56/A 0.03fF
C15953 OR2X1_LOC_56/A AND2X1_LOC_296/a_8_24# 0.01fF
C16343 OR2X1_LOC_527/a_8_216# OR2X1_LOC_56/A 0.01fF
C16488 OR2X1_LOC_56/A AND2X1_LOC_818/a_8_24# 0.03fF
C16503 OR2X1_LOC_56/A AND2X1_LOC_458/a_36_24# 0.01fF
C17215 OR2X1_LOC_133/a_8_216# OR2X1_LOC_56/A 0.02fF
C18461 OR2X1_LOC_111/a_8_216# OR2X1_LOC_56/A 0.02fF
C22093 OR2X1_LOC_56/A OR2X1_LOC_820/B 0.02fF
C23417 AND2X1_LOC_327/a_8_24# OR2X1_LOC_56/A 0.01fF
C23681 AND2X1_LOC_121/a_8_24# OR2X1_LOC_56/A 0.02fF
C25727 OR2X1_LOC_159/a_8_216# OR2X1_LOC_56/A 0.05fF
C26254 OR2X1_LOC_236/a_8_216# OR2X1_LOC_56/A 0.46fF
C29762 OR2X1_LOC_55/a_8_216# OR2X1_LOC_56/A 0.05fF
C30556 OR2X1_LOC_77/a_8_216# OR2X1_LOC_56/A 0.01fF
C36318 AND2X1_LOC_185/a_8_24# OR2X1_LOC_56/A 0.04fF
C37489 OR2X1_LOC_304/a_8_216# OR2X1_LOC_56/A 0.03fF
C38386 OR2X1_LOC_90/a_8_216# OR2X1_LOC_56/A 0.01fF
C39405 OR2X1_LOC_73/a_8_216# OR2X1_LOC_56/A 0.01fF
C45263 OR2X1_LOC_9/a_8_216# OR2X1_LOC_56/A 0.01fF
C45393 OR2X1_LOC_56/A OR2X1_LOC_48/a_8_216# 0.07fF
C47600 AND2X1_LOC_185/a_36_24# OR2X1_LOC_56/A 0.01fF
C48387 OR2X1_LOC_56/A OR2X1_LOC_382/a_8_216# 0.03fF
C51304 OR2X1_LOC_56/A OR2X1_LOC_381/a_8_216# 0.01fF
C52286 OR2X1_LOC_699/a_8_216# OR2X1_LOC_56/A 0.02fF
C54370 OR2X1_LOC_94/a_8_216# OR2X1_LOC_56/A 0.02fF
C55356 OR2X1_LOC_54/a_8_216# OR2X1_LOC_56/A 0.02fF
C56131 OR2X1_LOC_56/A AND2X1_LOC_458/a_8_24# 0.05fF
C41647 AND2X1_LOC_611/a_8_24# AND2X1_LOC_612/B 0.02fF
C4996 OR2X1_LOC_91/A OR2X1_LOC_820/B 0.61fF
C10240 OR2X1_LOC_91/A AND2X1_LOC_685/a_8_24# 0.01fF
C13648 OR2X1_LOC_91/A OR2X1_LOC_77/a_8_216# 0.43fF
C14538 OR2X1_LOC_91/A AND2X1_LOC_687/a_8_24# 0.01fF
C16815 OR2X1_LOC_681/a_8_216# OR2X1_LOC_91/A 0.01fF
C23355 OR2X1_LOC_694/a_8_216# OR2X1_LOC_91/A 0.02fF
C41953 OR2X1_LOC_682/a_8_216# OR2X1_LOC_91/A 0.01fF
C44174 OR2X1_LOC_91/A OR2X1_LOC_681/Y 0.02fF
C51966 OR2X1_LOC_91/A OR2X1_LOC_225/a_8_216# 0.01fF
C27147 AND2X1_LOC_94/Y OR2X1_LOC_82/a_8_216# 0.13fF
C32608 AND2X1_LOC_94/Y OR2X1_LOC_82/a_36_216# 0.02fF
C53169 AND2X1_LOC_94/Y AND2X1_LOC_42/a_8_24# 0.01fF
C616 OR2X1_LOC_485/A OR2X1_LOC_599/a_8_216# 0.01fF
C4160 OR2X1_LOC_527/a_8_216# OR2X1_LOC_485/A 0.06fF
C4976 OR2X1_LOC_485/A AND2X1_LOC_606/a_8_24# 0.03fF
C5953 AND2X1_LOC_502/a_8_24# OR2X1_LOC_485/A 0.02fF
C7702 AND2X1_LOC_598/a_8_24# OR2X1_LOC_485/A 0.02fF
C7791 OR2X1_LOC_485/A OR2X1_LOC_92/a_8_216# 0.01fF
C7818 OR2X1_LOC_485/A OR2X1_LOC_419/a_8_216# 0.01fF
C8128 OR2X1_LOC_306/a_8_216# OR2X1_LOC_485/A 0.03fF
C8162 OR2X1_LOC_485/A OR2X1_LOC_246/a_8_216# 0.01fF
C13953 OR2X1_LOC_485/A OR2X1_LOC_753/a_8_216# -0.00fF
C17527 OR2X1_LOC_485/A OR2X1_LOC_226/a_8_216# 0.01fF
C20653 OR2X1_LOC_485/A OR2X1_LOC_150/a_8_216# 0.01fF
C25206 OR2X1_LOC_485/A OR2X1_LOC_255/a_8_216# 0.01fF
C25376 OR2X1_LOC_304/a_8_216# OR2X1_LOC_485/A 0.01fF
C28166 OR2X1_LOC_485/A AND2X1_LOC_801/B 0.01fF
C31294 OR2X1_LOC_485/A OR2X1_LOC_530/a_8_216# 0.04fF
C33683 OR2X1_LOC_485/A OR2X1_LOC_760/a_8_216# 0.01fF
C36518 OR2X1_LOC_485/A AND2X1_LOC_294/a_8_24# 0.01fF
C38930 OR2X1_LOC_329/a_8_216# OR2X1_LOC_485/A 0.02fF
C39468 OR2X1_LOC_485/A OR2X1_LOC_71/a_8_216# 0.03fF
C42163 OR2X1_LOC_485/A OR2X1_LOC_10/a_8_216# 0.01fF
C42485 OR2X1_LOC_485/A OR2X1_LOC_256/a_8_216# 0.40fF
C48596 OR2X1_LOC_485/A OR2X1_LOC_63/a_8_216# 0.01fF
C50174 OR2X1_LOC_102/a_8_216# OR2X1_LOC_485/A 0.01fF
C8599 AND2X1_LOC_246/a_8_24# OR2X1_LOC_342/B 0.01fF
C4761 OR2X1_LOC_85/a_8_216# OR2X1_LOC_278/Y 0.01fF
C35979 OR2X1_LOC_625/a_8_216# OR2X1_LOC_278/Y 0.01fF
C1275 AND2X1_LOC_136/a_8_24# OR2X1_LOC_78/B 0.03fF
C2009 AND2X1_LOC_749/a_8_24# OR2X1_LOC_78/B 0.01fF
C3750 AND2X1_LOC_748/a_8_24# OR2X1_LOC_78/B 0.04fF
C6564 OR2X1_LOC_686/A OR2X1_LOC_78/B 0.02fF
C8660 OR2X1_LOC_78/B OR2X1_LOC_398/a_8_216# 0.05fF
C14166 OR2X1_LOC_78/B OR2X1_LOC_398/a_36_216# 0.02fF
C14398 AND2X1_LOC_80/a_8_24# OR2X1_LOC_78/B 0.05fF
C14792 AND2X1_LOC_748/a_36_24# OR2X1_LOC_78/B 0.01fF
C17168 OR2X1_LOC_78/B OR2X1_LOC_502/a_8_216# 0.05fF
C22497 OR2X1_LOC_100/a_8_216# OR2X1_LOC_78/B 0.02fF
C25423 AND2X1_LOC_49/a_8_24# OR2X1_LOC_78/B 0.04fF
C30117 AND2X1_LOC_38/a_8_24# OR2X1_LOC_78/B 0.04fF
C30193 AND2X1_LOC_681/a_8_24# OR2X1_LOC_78/B 0.03fF
C32416 OR2X1_LOC_78/B AND2X1_LOC_417/a_8_24# 0.01fF
C33598 AND2X1_LOC_684/a_8_24# OR2X1_LOC_78/B 0.02fF
C33613 AND2X1_LOC_6/a_8_24# OR2X1_LOC_78/B 0.01fF
C36120 AND2X1_LOC_699/a_8_24# OR2X1_LOC_78/B 0.01fF
C41103 AND2X1_LOC_38/a_36_24# OR2X1_LOC_78/B 0.01fF
C41946 AND2X1_LOC_49/a_36_24# OR2X1_LOC_78/B 0.01fF
C44542 OR2X1_LOC_264/a_8_216# OR2X1_LOC_78/B 0.35fF
C48495 AND2X1_LOC_682/a_8_24# OR2X1_LOC_78/B 0.02fF
C49822 AND2X1_LOC_490/a_8_24# OR2X1_LOC_78/B 0.01fF
C52753 AND2X1_LOC_683/a_8_24# OR2X1_LOC_78/B 0.06fF
C1905 OR2X1_LOC_161/A AND2X1_LOC_246/a_36_24# 0.01fF
C3543 AND2X1_LOC_681/a_8_24# OR2X1_LOC_161/A 0.01fF
C4234 AND2X1_LOC_696/a_8_24# OR2X1_LOC_161/A 0.02fF
C5988 OR2X1_LOC_750/a_8_216# OR2X1_LOC_161/A 0.07fF
C7683 AND2X1_LOC_111/a_8_24# OR2X1_LOC_161/A 0.03fF
C7997 AND2X1_LOC_110/a_8_24# OR2X1_LOC_161/A 0.02fF
C13976 AND2X1_LOC_306/a_8_24# OR2X1_LOC_161/A 0.01fF
C19041 AND2X1_LOC_110/a_36_24# OR2X1_LOC_161/A 0.01fF
C21687 AND2X1_LOC_682/a_8_24# OR2X1_LOC_161/A 0.01fF
C23540 OR2X1_LOC_276/B OR2X1_LOC_161/A 0.02fF
C24307 AND2X1_LOC_111/a_36_24# OR2X1_LOC_161/A 0.01fF
C25960 AND2X1_LOC_430/a_8_24# OR2X1_LOC_161/A 0.05fF
C32011 OR2X1_LOC_161/A AND2X1_LOC_760/a_8_24# 0.04fF
C34256 AND2X1_LOC_71/a_8_24# OR2X1_LOC_161/A 0.01fF
C35542 AND2X1_LOC_304/a_8_24# OR2X1_LOC_161/A 0.01fF
C36381 AND2X1_LOC_48/a_8_24# OR2X1_LOC_161/A 0.04fF
C44452 AND2X1_LOC_534/a_8_24# OR2X1_LOC_161/A 0.01fF
C45229 OR2X1_LOC_161/A OR2X1_LOC_515/a_8_216# 0.05fF
C47668 AND2X1_LOC_48/a_36_24# OR2X1_LOC_161/A 0.01fF
C48584 AND2X1_LOC_159/a_8_24# OR2X1_LOC_161/A 0.01fF
C48800 OR2X1_LOC_161/A AND2X1_LOC_760/a_36_24# 0.01fF
C54776 AND2X1_LOC_310/a_8_24# OR2X1_LOC_161/A 0.17fF
C55202 AND2X1_LOC_387/a_8_24# OR2X1_LOC_161/A 0.02fF
C2186 AND2X1_LOC_41/A AND2X1_LOC_23/a_8_24# 0.04fF
C5356 AND2X1_LOC_41/A AND2X1_LOC_422/a_8_24# 0.02fF
C5697 AND2X1_LOC_41/A AND2X1_LOC_255/a_36_24# 0.01fF
C5755 AND2X1_LOC_144/a_8_24# AND2X1_LOC_41/A 0.04fF
C6805 AND2X1_LOC_41/A OR2X1_LOC_750/a_8_216# 0.01fF
C10832 AND2X1_LOC_41/A OR2X1_LOC_120/a_8_216# 0.05fF
C17293 AND2X1_LOC_41/A OR2X1_LOC_274/a_8_216# 0.01fF
C17686 AND2X1_LOC_41/A AND2X1_LOC_693/a_8_24# 0.01fF
C18669 AND2X1_LOC_41/A OR2X1_LOC_264/a_8_216# 0.09fF
C19048 AND2X1_LOC_753/a_8_24# AND2X1_LOC_41/A 0.03fF
C21960 AND2X1_LOC_41/A OR2X1_LOC_596/a_8_216# 0.01fF
C24327 AND2X1_LOC_41/A OR2X1_LOC_276/B 0.07fF
C25716 AND2X1_LOC_41/A AND2X1_LOC_256/a_8_24# 0.06fF
C27700 AND2X1_LOC_41/A OR2X1_LOC_512/a_8_216# 0.01fF
C29665 AND2X1_LOC_41/A OR2X1_LOC_264/a_36_216# 0.03fF
C29836 AND2X1_LOC_41/A OR2X1_LOC_513/a_8_216# 0.01fF
C30356 OR2X1_LOC_121/a_8_216# AND2X1_LOC_41/A 0.01fF
C36335 AND2X1_LOC_41/A OR2X1_LOC_294/a_8_216# 0.08fF
C50911 AND2X1_LOC_41/A AND2X1_LOC_255/a_8_24# 0.06fF
C54337 AND2X1_LOC_421/a_8_24# AND2X1_LOC_41/A 0.01fF
C55803 AND2X1_LOC_41/A AND2X1_LOC_692/a_8_24# 0.02fF
C56003 AND2X1_LOC_387/a_8_24# AND2X1_LOC_41/A 0.01fF
C8108 AND2X1_LOC_382/a_8_24# OR2X1_LOC_848/A 0.02fF
C38309 OR2X1_LOC_848/A AND2X1_LOC_236/a_8_24# 0.02fF
C2196 AND2X1_LOC_548/a_8_24# OR2X1_LOC_39/A 0.01fF
C3488 OR2X1_LOC_277/a_8_216# OR2X1_LOC_39/A 0.01fF
C4237 AND2X1_LOC_264/a_8_24# OR2X1_LOC_39/A 0.03fF
C10740 OR2X1_LOC_412/a_8_216# OR2X1_LOC_39/A 0.01fF
C12942 OR2X1_LOC_88/a_8_216# OR2X1_LOC_39/A 0.01fF
C15318 OR2X1_LOC_126/a_8_216# OR2X1_LOC_39/A 0.03fF
C15932 OR2X1_LOC_39/A OR2X1_LOC_19/a_8_216# 0.06fF
C17359 AND2X1_LOC_276/a_8_24# OR2X1_LOC_39/A 0.03fF
C18354 OR2X1_LOC_119/a_8_216# OR2X1_LOC_39/A 0.01fF
C19064 AND2X1_LOC_377/Y OR2X1_LOC_39/A 0.03fF
C22872 OR2X1_LOC_530/a_8_216# OR2X1_LOC_39/A 0.01fF
C24591 AND2X1_LOC_378/a_8_24# OR2X1_LOC_39/A 0.09fF
C30099 AND2X1_LOC_155/a_8_24# OR2X1_LOC_39/A 0.01fF
C30505 OR2X1_LOC_23/a_8_216# OR2X1_LOC_39/A 0.02fF
C31056 OR2X1_LOC_275/a_8_216# OR2X1_LOC_39/A 0.03fF
C31647 OR2X1_LOC_126/a_36_216# OR2X1_LOC_39/A 0.02fF
C35667 AND2X1_LOC_120/a_8_24# OR2X1_LOC_39/A 0.11fF
C38532 AND2X1_LOC_274/a_8_24# OR2X1_LOC_39/A 0.04fF
C44342 OR2X1_LOC_39/A OR2X1_LOC_153/a_8_216# 0.02fF
C46871 OR2X1_LOC_696/a_8_216# OR2X1_LOC_39/A 0.06fF
C48892 OR2X1_LOC_743/a_8_216# OR2X1_LOC_39/A 0.01fF
C51112 OR2X1_LOC_271/Y OR2X1_LOC_39/A 0.13fF
C53230 AND2X1_LOC_688/a_8_24# OR2X1_LOC_39/A 0.03fF
C10194 OR2X1_LOC_382/Y AND2X1_LOC_818/a_8_24# 0.01fF
C15660 OR2X1_LOC_382/Y OR2X1_LOC_820/B 0.90fF
C3604 OR2X1_LOC_329/a_8_216# OR2X1_LOC_428/A 0.04fF
C7810 OR2X1_LOC_18/a_8_216# OR2X1_LOC_428/A 0.01fF
C11341 OR2X1_LOC_682/a_8_216# OR2X1_LOC_428/A 0.05fF
C12020 OR2X1_LOC_428/A AND2X1_LOC_269/a_8_24# 0.10fF
C12197 OR2X1_LOC_6/a_8_216# OR2X1_LOC_428/A 0.02fF
C21239 OR2X1_LOC_225/a_8_216# OR2X1_LOC_428/A 0.01fF
C24131 OR2X1_LOC_271/Y OR2X1_LOC_428/A 0.03fF
C33816 OR2X1_LOC_93/a_8_216# OR2X1_LOC_428/A 0.02fF
C34619 OR2X1_LOC_236/a_8_216# OR2X1_LOC_428/A 0.01fF
C43119 OR2X1_LOC_763/a_8_216# OR2X1_LOC_428/A 0.05fF
C46079 OR2X1_LOC_304/a_8_216# OR2X1_LOC_428/A 0.02fF
C48792 OR2X1_LOC_422/a_8_216# OR2X1_LOC_428/A 0.01fF
C54058 OR2X1_LOC_428/A OR2X1_LOC_387/a_8_216# 0.06fF
C54671 OR2X1_LOC_421/a_8_216# OR2X1_LOC_428/A 0.01fF
C29813 AND2X1_LOC_519/a_8_24# OR2X1_LOC_87/B 0.02fF
C41179 OR2X1_LOC_87/B AND2X1_LOC_19/a_8_24# 0.04fF
C41607 AND2X1_LOC_29/a_8_24# OR2X1_LOC_87/B 0.04fF
C52420 OR2X1_LOC_87/B AND2X1_LOC_19/a_36_24# 0.01fF
C53278 AND2X1_LOC_46/a_8_24# OR2X1_LOC_87/B 0.19fF
C2039 AND2X1_LOC_82/Y AND2X1_LOC_490/a_8_24# 0.01fF
C15929 AND2X1_LOC_81/B OR2X1_LOC_502/a_8_216# 0.01fF
C21271 OR2X1_LOC_100/a_8_216# AND2X1_LOC_81/B 0.02fF
C277 OR2X1_LOC_684/a_8_216# OR2X1_LOC_427/A 0.01fF
C434 OR2X1_LOC_430/a_8_216# OR2X1_LOC_427/A 0.01fF
C2313 OR2X1_LOC_427/A OR2X1_LOC_164/a_8_216# 0.04fF
C2974 OR2X1_LOC_529/a_8_216# OR2X1_LOC_427/A 0.03fF
C5488 OR2X1_LOC_696/a_8_216# OR2X1_LOC_427/A 0.02fF
C5604 OR2X1_LOC_427/A AND2X1_LOC_405/a_8_24# 0.01fF
C7134 AND2X1_LOC_374/a_8_24# OR2X1_LOC_427/A 0.01fF
C7523 OR2X1_LOC_427/A OR2X1_LOC_582/a_8_216# 0.05fF
C10116 OR2X1_LOC_427/A AND2X1_LOC_296/a_8_24# 0.10fF
C10643 OR2X1_LOC_427/A AND2X1_LOC_818/a_8_24# 0.01fF
C14158 OR2X1_LOC_426/a_8_216# OR2X1_LOC_427/A 0.01fF
C16120 OR2X1_LOC_427/A OR2X1_LOC_820/B 0.02fF
C16690 OR2X1_LOC_427/A AND2X1_LOC_405/a_36_24# 0.01fF
C20120 OR2X1_LOC_427/A OR2X1_LOC_511/a_8_216# 0.02fF
C20249 OR2X1_LOC_427/A OR2X1_LOC_753/a_8_216# 0.01fF
C20410 OR2X1_LOC_427/A OR2X1_LOC_236/a_8_216# 0.01fF
C23933 OR2X1_LOC_427/A OR2X1_LOC_55/a_8_216# 0.02fF
C24745 OR2X1_LOC_427/A OR2X1_LOC_77/a_8_216# 0.01fF
C26265 OR2X1_LOC_628/a_8_216# OR2X1_LOC_427/A 0.02fF
C29641 OR2X1_LOC_683/a_8_216# OR2X1_LOC_427/A 0.01fF
C29950 OR2X1_LOC_427/A AND2X1_LOC_407/a_8_24# 0.04fF
C32547 OR2X1_LOC_90/a_8_216# OR2X1_LOC_427/A 0.40fF
C34292 OR2X1_LOC_694/a_8_216# OR2X1_LOC_427/A 0.07fF
C40930 OR2X1_LOC_427/A AND2X1_LOC_407/a_36_24# 0.01fF
C42293 OR2X1_LOC_427/A OR2X1_LOC_382/a_8_216# 0.02fF
C45314 OR2X1_LOC_427/A OR2X1_LOC_381/a_8_216# 0.01fF
C46363 OR2X1_LOC_699/a_8_216# OR2X1_LOC_427/A 0.05fF
C49492 OR2X1_LOC_427/A AND2X1_LOC_686/a_8_24# 0.02fF
C52160 OR2X1_LOC_427/A OR2X1_LOC_373/a_8_216# 0.02fF
C55134 OR2X1_LOC_427/A OR2X1_LOC_322/a_8_216# 0.01fF
C5015 OR2X1_LOC_446/B AND2X1_LOC_419/a_8_24# 0.01fF
C17326 OR2X1_LOC_446/B OR2X1_LOC_512/a_8_216# 0.03fF
C21706 OR2X1_LOC_446/B AND2X1_LOC_419/a_36_24# -0.00fF
C26056 AND2X1_LOC_304/a_8_24# OR2X1_LOC_446/B 0.04fF
C35610 OR2X1_LOC_446/B OR2X1_LOC_515/a_8_216# 0.01fF
C37006 AND2X1_LOC_304/a_36_24# OR2X1_LOC_446/B 0.01fF
C47250 AND2X1_LOC_289/a_8_24# OR2X1_LOC_333/A 0.13fF
C36588 AND2X1_LOC_309/a_8_24# OR2X1_LOC_335/B 0.02fF
C41222 AND2X1_LOC_387/a_8_24# OR2X1_LOC_750/Y 0.25fF
C5313 OR2X1_LOC_516/A AND2X1_LOC_515/a_8_24# 0.01fF
C28304 OR2X1_LOC_325/A AND2X1_LOC_322/a_8_24# 0.23fF
C36692 OR2X1_LOC_325/A AND2X1_LOC_323/a_8_24# 0.01fF
C8695 OR2X1_LOC_691/Y AND2X1_LOC_760/a_8_24# 0.01fF
C9646 AND2X1_LOC_748/a_8_24# OR2X1_LOC_691/Y 0.01fF
C20618 OR2X1_LOC_691/Y OR2X1_LOC_800/Y 0.01fF
C31823 OR2X1_LOC_691/Y AND2X1_LOC_761/a_8_24# 0.01fF
C37058 OR2X1_LOC_691/Y OR2X1_LOC_801/a_8_216# 0.01fF
C37139 OR2X1_LOC_800/a_8_216# OR2X1_LOC_691/Y 0.01fF
C40837 AND2X1_LOC_599/a_8_24# OR2X1_LOC_691/Y 0.01fF
C41295 OR2X1_LOC_691/Y OR2X1_LOC_185/a_8_216# 0.01fF
C10468 AND2X1_LOC_462/B AND2X1_LOC_293/a_36_24# 0.01fF
C38806 AND2X1_LOC_462/B AND2X1_LOC_293/a_8_24# 0.08fF
C19202 OR2X1_LOC_824/a_8_216# OR2X1_LOC_824/Y 0.01fF
C10197 OR2X1_LOC_129/a_8_216# OR2X1_LOC_291/Y 0.02fF
C24799 OR2X1_LOC_291/Y OR2X1_LOC_277/a_8_216# 0.02fF
C3001 AND2X1_LOC_421/a_8_24# OR2X1_LOC_269/B 0.01fF
C4558 AND2X1_LOC_387/a_8_24# OR2X1_LOC_269/B 0.01fF
C6890 AND2X1_LOC_23/a_8_24# OR2X1_LOC_269/B 0.02fF
C10221 AND2X1_LOC_422/a_8_24# OR2X1_LOC_269/B 0.01fF
C10602 AND2X1_LOC_144/a_8_24# OR2X1_LOC_269/B 0.01fF
C11059 OR2X1_LOC_269/a_8_216# OR2X1_LOC_269/B 0.04fF
C11592 OR2X1_LOC_750/a_8_216# OR2X1_LOC_269/B -0.06fF
C13120 AND2X1_LOC_511/a_8_24# OR2X1_LOC_269/B 0.01fF
C13298 AND2X1_LOC_43/a_36_24# OR2X1_LOC_269/B 0.01fF
C16571 OR2X1_LOC_269/a_36_216# OR2X1_LOC_269/B 0.03fF
C22718 OR2X1_LOC_750/a_36_216# OR2X1_LOC_269/B 0.01fF
C23850 AND2X1_LOC_753/a_8_24# OR2X1_LOC_269/B 0.06fF
C28500 AND2X1_LOC_329/a_8_24# OR2X1_LOC_269/B 0.03fF
C28992 OR2X1_LOC_276/B OR2X1_LOC_269/B 0.25fF
C32354 OR2X1_LOC_269/B OR2X1_LOC_512/a_8_216# 0.12fF
C41087 AND2X1_LOC_304/a_8_24# OR2X1_LOC_269/B 0.03fF
C41971 AND2X1_LOC_48/a_8_24# OR2X1_LOC_269/B 0.01fF
C43915 OR2X1_LOC_269/B AND2X1_LOC_225/a_8_24# 0.01fF
C51543 AND2X1_LOC_382/a_8_24# OR2X1_LOC_269/B 0.21fF
C52229 OR2X1_LOC_691/a_8_216# OR2X1_LOC_269/B 0.04fF
C52336 AND2X1_LOC_304/a_36_24# OR2X1_LOC_269/B 0.01fF
C55013 AND2X1_LOC_271/a_8_24# OR2X1_LOC_269/B 0.01fF
C14978 OR2X1_LOC_32/B OR2X1_LOC_412/a_8_216# -0.01fF
C34728 OR2X1_LOC_32/B OR2X1_LOC_23/a_8_216# 0.43fF
C49280 OR2X1_LOC_129/a_8_216# OR2X1_LOC_32/B 0.03fF
C897 AND2X1_LOC_683/a_8_24# OR2X1_LOC_87/A 0.02fF
C1172 OR2X1_LOC_155/a_8_216# OR2X1_LOC_87/A 0.04fF
C10931 AND2X1_LOC_150/a_8_24# OR2X1_LOC_87/A 0.03fF
C10944 OR2X1_LOC_686/A OR2X1_LOC_87/A 0.02fF
C11503 OR2X1_LOC_87/A OR2X1_LOC_87/a_8_216# 0.05fF
C20693 OR2X1_LOC_87/A AND2X1_LOC_226/a_36_24# 0.02fF
C25942 OR2X1_LOC_87/A OR2X1_LOC_68/a_8_216# 0.01fF
C29642 AND2X1_LOC_310/a_8_24# OR2X1_LOC_87/A 0.03fF
C34451 AND2X1_LOC_681/a_8_24# OR2X1_LOC_87/A 0.01fF
C35223 OR2X1_LOC_87/A AND2X1_LOC_19/a_8_24# 0.15fF
C37271 AND2X1_LOC_527/a_8_24# OR2X1_LOC_87/A 0.03fF
C37337 AND2X1_LOC_373/a_8_24# OR2X1_LOC_87/A 0.01fF
C37829 OR2X1_LOC_87/A AND2X1_LOC_684/a_8_24# 0.02fF
C47129 AND2X1_LOC_743/a_8_24# OR2X1_LOC_87/A 0.04fF
C52777 AND2X1_LOC_682/a_8_24# OR2X1_LOC_87/A 0.02fF
C52806 OR2X1_LOC_87/A AND2X1_LOC_129/a_8_24# 0.01fF
C53668 AND2X1_LOC_153/a_8_24# OR2X1_LOC_87/A 0.03fF
C54703 OR2X1_LOC_87/A AND2X1_LOC_226/a_8_24# 0.02fF
C8868 AND2X1_LOC_10/a_8_24# OR2X1_LOC_161/B 0.01fF
C10645 AND2X1_LOC_681/a_8_24# OR2X1_LOC_161/B 0.01fF
C12164 AND2X1_LOC_426/a_8_24# OR2X1_LOC_161/B 0.01fF
C12607 AND2X1_LOC_63/a_8_24# OR2X1_LOC_161/B 0.01fF
C14070 AND2X1_LOC_684/a_8_24# OR2X1_LOC_161/B 0.01fF
C14785 AND2X1_LOC_111/a_8_24# OR2X1_LOC_161/B 0.01fF
C14834 AND2X1_LOC_694/a_8_24# OR2X1_LOC_161/B 0.10fF
C15086 AND2X1_LOC_110/a_8_24# OR2X1_LOC_161/B 0.01fF
C21066 AND2X1_LOC_306/a_8_24# OR2X1_LOC_161/B 0.01fF
C23160 AND2X1_LOC_743/a_8_24# OR2X1_LOC_161/B 0.01fF
C28221 OR2X1_LOC_596/a_8_216# OR2X1_LOC_161/B 0.01fF
C28659 AND2X1_LOC_582/a_8_24# OR2X1_LOC_161/B 0.09fF
C28695 AND2X1_LOC_682/a_8_24# OR2X1_LOC_161/B 0.01fF
C29600 OR2X1_LOC_296/a_8_216# OR2X1_LOC_161/B 0.02fF
C32975 AND2X1_LOC_683/a_8_24# OR2X1_LOC_161/B 0.01fF
C39952 OR2X1_LOC_161/B OR2X1_LOC_374/a_8_216# 0.01fF
C40083 AND2X1_LOC_748/a_8_24# OR2X1_LOC_161/B 0.02fF
C42697 OR2X1_LOC_294/a_8_216# OR2X1_LOC_161/B 0.01fF
C43068 AND2X1_LOC_150/a_8_24# OR2X1_LOC_161/B 0.01fF
C43079 OR2X1_LOC_686/A OR2X1_LOC_161/B 0.52fF
C51212 OR2X1_LOC_161/B OR2X1_LOC_374/a_36_216# 0.01fF
C51689 AND2X1_LOC_534/a_8_24# OR2X1_LOC_161/B 0.02fF
C18249 OR2X1_LOC_589/A OR2X1_LOC_245/a_8_216# 0.01fF
C26117 OR2X1_LOC_129/a_8_216# OR2X1_LOC_589/A 0.01fF
C27064 OR2X1_LOC_589/A AND2X1_LOC_87/a_8_24# 0.01fF
C29399 OR2X1_LOC_589/A OR2X1_LOC_599/a_8_216# 0.02fF
C38450 OR2X1_LOC_589/A OR2X1_LOC_433/a_8_216# 0.05fF
C41462 OR2X1_LOC_589/A AND2X1_LOC_264/a_8_24# 0.17fF
C51488 OR2X1_LOC_589/A AND2X1_LOC_800/a_8_24# 0.03fF
C47494 OR2X1_LOC_820/A OR2X1_LOC_748/Y 0.05fF
C51220 OR2X1_LOC_748/a_8_216# OR2X1_LOC_748/Y -0.00fF
C12177 OR2X1_LOC_269/a_8_216# OR2X1_LOC_344/A 0.01fF
C17932 OR2X1_LOC_344/A AND2X1_LOC_268/a_8_24# 0.20fF
C28963 OR2X1_LOC_344/A OR2X1_LOC_269/A 0.01fF
C30142 OR2X1_LOC_276/B OR2X1_LOC_344/A 0.02fF
C56223 AND2X1_LOC_271/a_8_24# OR2X1_LOC_344/A 0.01fF
C3121 AND2X1_LOC_685/a_36_24# OR2X1_LOC_7/A 0.01fF
C5436 OR2X1_LOC_421/a_8_216# OR2X1_LOC_7/A 0.04fF
C7385 AND2X1_LOC_687/a_36_24# OR2X1_LOC_7/A 0.01fF
C8171 OR2X1_LOC_7/A AND2X1_LOC_294/a_8_24# 0.04fF
C10236 AND2X1_LOC_155/a_8_24# OR2X1_LOC_7/A -0.00fF
C14092 OR2X1_LOC_256/a_8_216# OR2X1_LOC_7/A 0.01fF
C18350 OR2X1_LOC_682/a_8_216# OR2X1_LOC_7/A 0.04fF
C20520 OR2X1_LOC_681/Y OR2X1_LOC_7/A 0.02fF
C20942 OR2X1_LOC_299/a_8_216# OR2X1_LOC_7/A 0.02fF
C21307 AND2X1_LOC_155/a_36_24# OR2X1_LOC_7/A 0.01fF
C21636 OR2X1_LOC_102/a_8_216# OR2X1_LOC_7/A 0.01fF
C25169 OR2X1_LOC_488/a_8_216# OR2X1_LOC_7/A 0.01fF
C28816 OR2X1_LOC_7/A OR2X1_LOC_743/a_8_216# 0.04fF
C31053 OR2X1_LOC_271/Y OR2X1_LOC_7/A 0.15fF
C31872 OR2X1_LOC_299/a_36_216# OR2X1_LOC_7/A 0.02fF
C40753 OR2X1_LOC_93/a_8_216# OR2X1_LOC_7/A 0.39fF
C41448 OR2X1_LOC_7/A OR2X1_LOC_753/a_8_216# -0.01fF
C42569 AND2X1_LOC_685/a_8_24# OR2X1_LOC_7/A 0.05fF
C46977 AND2X1_LOC_687/a_8_24# OR2X1_LOC_7/A 0.03fF
C47732 OR2X1_LOC_628/a_8_216# OR2X1_LOC_7/A 0.01fF
C48877 OR2X1_LOC_7/A OR2X1_LOC_323/a_8_216# 0.07fF
C49363 OR2X1_LOC_681/a_8_216# OR2X1_LOC_7/A 0.03fF
C52920 OR2X1_LOC_255/a_8_216# OR2X1_LOC_7/A 0.01fF
C53119 OR2X1_LOC_490/a_8_216# OR2X1_LOC_7/A 0.06fF
C55759 OR2X1_LOC_422/a_8_216# OR2X1_LOC_7/A 0.03fF
C55793 OR2X1_LOC_694/a_8_216# OR2X1_LOC_7/A 0.03fF
C5380 AND2X1_LOC_19/Y AND2X1_LOC_129/a_36_24# 0.01fF
C33036 AND2X1_LOC_19/Y AND2X1_LOC_19/a_8_24# 0.01fF
C50604 AND2X1_LOC_19/Y AND2X1_LOC_129/a_8_24# 0.22fF
C48695 OR2X1_LOC_557/A AND2X1_LOC_15/a_8_24# 0.01fF
C7558 OR2X1_LOC_529/a_8_216# OR2X1_LOC_744/A 0.05fF
C12170 OR2X1_LOC_744/A OR2X1_LOC_743/a_8_216# 0.02fF
C13848 OR2X1_LOC_693/a_8_216# OR2X1_LOC_744/A 0.01fF
C14345 OR2X1_LOC_692/a_8_216# OR2X1_LOC_744/A 0.01fF
C14421 OR2X1_LOC_744/A OR2X1_LOC_271/Y 0.03fF
C18651 AND2X1_LOC_598/a_8_24# OR2X1_LOC_744/A 0.04fF
C20787 OR2X1_LOC_744/A OR2X1_LOC_433/a_8_216# 0.01fF
C23025 OR2X1_LOC_744/A OR2X1_LOC_277/a_8_216# 0.01fF
C25793 AND2X1_LOC_398/a_8_24# OR2X1_LOC_744/A 0.23fF
C28093 OR2X1_LOC_744/A OR2X1_LOC_64/a_8_216# 0.01fF
C29658 AND2X1_LOC_598/a_36_24# OR2X1_LOC_744/A 0.01fF
C32305 OR2X1_LOC_744/A OR2X1_LOC_88/a_8_216# 0.01fF
C33375 OR2X1_LOC_744/A OR2X1_LOC_763/a_8_216# 0.01fF
C34573 OR2X1_LOC_369/a_8_216# OR2X1_LOC_744/A 0.03fF
C34739 OR2X1_LOC_126/a_8_216# OR2X1_LOC_744/A 0.01fF
C35033 AND2X1_LOC_596/a_8_24# OR2X1_LOC_744/A 0.01fF
C37702 OR2X1_LOC_119/a_8_216# OR2X1_LOC_744/A 0.01fF
C38114 OR2X1_LOC_744/A OR2X1_LOC_762/a_8_216# 0.01fF
C40091 OR2X1_LOC_744/A OR2X1_LOC_26/a_8_216# 0.01fF
C45738 OR2X1_LOC_369/a_36_216# OR2X1_LOC_744/A 0.02fF
C51274 OR2X1_LOC_126/a_36_216# OR2X1_LOC_744/A -0.00fF
C55367 OR2X1_LOC_744/A OR2X1_LOC_80/a_8_216# 0.01fF
C1912 AND2X1_LOC_515/a_8_24# OR2X1_LOC_600/A 0.01fF
C2131 OR2X1_LOC_600/A AND2X1_LOC_814/a_8_24# 0.07fF
C2551 OR2X1_LOC_600/A OR2X1_LOC_417/a_8_216# 0.01fF
C5384 OR2X1_LOC_600/A AND2X1_LOC_458/a_8_24# 0.02fF
C5450 OR2X1_LOC_611/a_8_216# OR2X1_LOC_600/A 0.02fF
C5932 OR2X1_LOC_600/A OR2X1_LOC_80/a_8_216# 0.01fF
C10876 OR2X1_LOC_104/a_8_216# OR2X1_LOC_600/A 0.02fF
C11509 OR2X1_LOC_600/A OR2X1_LOC_80/a_36_216# 0.02fF
C11715 AND2X1_LOC_410/a_8_24# OR2X1_LOC_600/A 0.01fF
C13658 OR2X1_LOC_600/A OR2X1_LOC_411/a_8_216# 0.03fF
C14354 OR2X1_LOC_529/a_8_216# OR2X1_LOC_600/A 0.03fF
C15416 OR2X1_LOC_600/A AND2X1_LOC_750/a_8_24# 0.01fF
C15946 OR2X1_LOC_600/A OR2X1_LOC_819/a_8_216# 0.01fF
C18031 OR2X1_LOC_600/A OR2X1_LOC_15/a_8_216# 0.02fF
C18289 OR2X1_LOC_600/A OR2X1_LOC_225/a_8_216# -0.01fF
C19890 OR2X1_LOC_529/a_36_216# OR2X1_LOC_600/A 0.02fF
C21550 OR2X1_LOC_600/A AND2X1_LOC_296/a_8_24# 0.01fF
C22069 OR2X1_LOC_600/A AND2X1_LOC_818/a_8_24# 0.06fF
C23623 OR2X1_LOC_600/A OR2X1_LOC_15/a_36_216# 0.01fF
C27018 OR2X1_LOC_600/A OR2X1_LOC_820/A 0.01fF
C27508 OR2X1_LOC_600/A OR2X1_LOC_820/B 0.04fF
C28262 AND2X1_LOC_410/a_36_24# OR2X1_LOC_600/A -0.00fF
C28919 OR2X1_LOC_600/A OR2X1_LOC_29/a_8_216# 0.05fF
C30704 OR2X1_LOC_600/A OR2X1_LOC_748/a_8_216# 0.01fF
C30953 OR2X1_LOC_600/A AND2X1_LOC_847/a_8_24# 0.01fF
C31680 OR2X1_LOC_600/A OR2X1_LOC_46/a_8_216# 0.01fF
C31729 OR2X1_LOC_600/A OR2X1_LOC_236/a_8_216# -0.00fF
C32521 AND2X1_LOC_398/a_8_24# OR2X1_LOC_600/A 0.05fF
C35206 OR2X1_LOC_600/A OR2X1_LOC_55/a_8_216# 0.01fF
C36250 OR2X1_LOC_600/A OR2X1_LOC_14/a_8_216# 0.05fF
C38422 AND2X1_LOC_62/a_8_24# OR2X1_LOC_600/A 0.04fF
C45137 OR2X1_LOC_600/A OR2X1_LOC_749/a_8_216# 0.01fF
C49289 AND2X1_LOC_398/a_36_24# OR2X1_LOC_600/A 0.01fF
C51301 OR2X1_LOC_820/a_8_216# OR2X1_LOC_600/A 0.01fF
C54819 OR2X1_LOC_600/A OR2X1_LOC_817/a_8_216# 0.01fF
C55195 AND2X1_LOC_62/a_36_24# OR2X1_LOC_600/A 0.01fF
C709 OR2X1_LOC_490/a_8_216# AND2X1_LOC_101/B 0.47fF
C3055 OR2X1_LOC_473/A AND2X1_LOC_625/a_36_24# 0.01fF
C34134 OR2X1_LOC_276/B OR2X1_LOC_473/A 0.10fF
C39651 OR2X1_LOC_276/a_8_216# OR2X1_LOC_473/A -0.00fF
C48208 OR2X1_LOC_473/A AND2X1_LOC_625/a_8_24# 0.12fF
C50235 OR2X1_LOC_809/B AND2X1_LOC_111/a_8_24# 0.04fF
C352 AND2X1_LOC_38/a_8_24# AND2X1_LOC_18/Y 0.01fF
C2471 OR2X1_LOC_269/a_8_216# AND2X1_LOC_18/Y 0.01fF
C6953 AND2X1_LOC_18/Y OR2X1_LOC_120/a_8_216# 0.01fF
C7147 AND2X1_LOC_85/a_8_24# AND2X1_LOC_18/Y 0.10fF
C7420 AND2X1_LOC_263/a_8_24# AND2X1_LOC_18/Y 0.03fF
C8230 AND2X1_LOC_18/Y AND2X1_LOC_268/a_8_24# 0.01fF
C13466 OR2X1_LOC_274/a_8_216# AND2X1_LOC_18/Y 0.18fF
C13892 AND2X1_LOC_693/a_8_24# AND2X1_LOC_18/Y 0.01fF
C15167 AND2X1_LOC_753/a_8_24# AND2X1_LOC_18/Y 0.01fF
C16451 OR2X1_LOC_270/a_8_216# AND2X1_LOC_18/Y 0.08fF
C19255 AND2X1_LOC_18/Y OR2X1_LOC_269/A 0.01fF
C20459 OR2X1_LOC_276/B AND2X1_LOC_18/Y 0.21fF
C21915 AND2X1_LOC_18/Y AND2X1_LOC_256/a_8_24# 0.05fF
C24608 AND2X1_LOC_88/a_8_24# AND2X1_LOC_18/Y 0.02fF
C27470 OR2X1_LOC_405/a_8_216# AND2X1_LOC_18/Y 0.02fF
C28311 AND2X1_LOC_749/a_8_24# AND2X1_LOC_18/Y 0.01fF
C31247 AND2X1_LOC_71/a_8_24# AND2X1_LOC_18/Y 0.02fF
C45401 AND2X1_LOC_159/a_8_24# AND2X1_LOC_18/Y 0.06fF
C46442 AND2X1_LOC_271/a_8_24# AND2X1_LOC_18/Y 0.01fF
C47030 AND2X1_LOC_18/Y AND2X1_LOC_255/a_8_24# 0.01fF
C54660 AND2X1_LOC_433/a_8_24# AND2X1_LOC_18/Y 0.01fF
C2549 AND2X1_LOC_36/Y AND2X1_LOC_761/a_8_24# 0.02fF
C7290 OR2X1_LOC_598/a_8_216# AND2X1_LOC_36/Y 0.06fF
C8741 OR2X1_LOC_269/a_8_216# AND2X1_LOC_36/Y 0.01fF
C10170 AND2X1_LOC_6/a_8_24# AND2X1_LOC_36/Y 0.01fF
C11595 AND2X1_LOC_599/a_8_24# AND2X1_LOC_36/Y 0.04fF
C12578 AND2X1_LOC_18/a_8_24# AND2X1_LOC_36/Y 0.01fF
C12728 AND2X1_LOC_699/a_8_24# AND2X1_LOC_36/Y 0.02fF
C14485 AND2X1_LOC_36/Y AND2X1_LOC_268/a_8_24# 0.01fF
C16312 AND2X1_LOC_328/a_8_24# AND2X1_LOC_36/Y 0.01fF
C17837 AND2X1_LOC_36/Y AND2X1_LOC_419/a_8_24# 0.01fF
C19287 AND2X1_LOC_95/a_8_24# AND2X1_LOC_36/Y 0.01fF
C19415 AND2X1_LOC_46/a_8_24# AND2X1_LOC_36/Y 0.03fF
C20180 AND2X1_LOC_693/a_8_24# AND2X1_LOC_36/Y 0.14fF
C22839 OR2X1_LOC_270/a_8_216# AND2X1_LOC_36/Y 0.06fF
C25522 AND2X1_LOC_36/Y OR2X1_LOC_269/A 0.01fF
C26673 OR2X1_LOC_276/B AND2X1_LOC_36/Y 0.09fF
C28126 AND2X1_LOC_273/a_8_24# AND2X1_LOC_36/Y 0.03fF
C28152 AND2X1_LOC_256/a_8_24# AND2X1_LOC_36/Y 0.01fF
C28575 AND2X1_LOC_36/Y OR2X1_LOC_514/a_8_216# 0.01fF
C28681 AND2X1_LOC_36/a_8_24# AND2X1_LOC_36/Y 0.01fF
C29018 AND2X1_LOC_628/a_8_24# AND2X1_LOC_36/Y 0.01fF
C32770 OR2X1_LOC_121/a_8_216# AND2X1_LOC_36/Y 0.05fF
C33776 AND2X1_LOC_136/a_8_24# AND2X1_LOC_36/Y 0.01fF
C34158 AND2X1_LOC_102/a_8_24# AND2X1_LOC_36/Y 0.03fF
C36229 AND2X1_LOC_748/a_8_24# AND2X1_LOC_36/Y -0.00fF
C36606 AND2X1_LOC_693/a_36_24# AND2X1_LOC_36/Y 0.01fF
C37423 AND2X1_LOC_36/Y OR2X1_LOC_548/a_8_216# 0.01fF
C37927 AND2X1_LOC_26/a_8_24# AND2X1_LOC_36/Y 0.01fF
C38789 AND2X1_LOC_59/a_8_24# AND2X1_LOC_36/Y 0.01fF
C39161 OR2X1_LOC_686/A AND2X1_LOC_36/Y 0.25fF
C41246 AND2X1_LOC_530/a_8_24# AND2X1_LOC_36/Y 0.04fF
C43564 AND2X1_LOC_386/a_8_24# AND2X1_LOC_36/Y 0.01fF
C48599 AND2X1_LOC_36/Y OR2X1_LOC_515/a_8_216# 0.01fF
C49973 OR2X1_LOC_691/a_8_216# AND2X1_LOC_36/Y 0.06fF
C52432 AND2X1_LOC_36/Y AND2X1_LOC_619/a_8_24# 0.06fF
C52726 AND2X1_LOC_271/a_8_24# AND2X1_LOC_36/Y 0.01fF
C53443 AND2X1_LOC_64/a_8_24# AND2X1_LOC_36/Y 0.20fF
C55842 AND2X1_LOC_36/Y AND2X1_LOC_762/a_8_24# 0.01fF
C55993 AND2X1_LOC_43/a_8_24# AND2X1_LOC_36/Y 0.01fF
C246 OR2X1_LOC_121/a_8_216# OR2X1_LOC_375/A 0.01fF
C1220 OR2X1_LOC_410/a_8_216# OR2X1_LOC_375/A 0.06fF
C1741 AND2X1_LOC_102/a_8_24# OR2X1_LOC_375/A 0.01fF
C4178 AND2X1_LOC_126/a_8_24# OR2X1_LOC_375/A 0.04fF
C12118 OR2X1_LOC_375/A AND2X1_LOC_581/a_8_24# 0.20fF
C14612 OR2X1_LOC_375/A OR2X1_LOC_66/a_8_216# 0.01fF
C14741 AND2X1_LOC_90/a_8_24# OR2X1_LOC_375/A 0.01fF
C15231 AND2X1_LOC_126/a_36_24# OR2X1_LOC_375/A 0.01fF
C15959 OR2X1_LOC_375/A OR2X1_LOC_375/a_8_216# 0.02fF
C19240 AND2X1_LOC_56/a_8_24# OR2X1_LOC_375/A 0.02fF
C19661 AND2X1_LOC_519/a_8_24# OR2X1_LOC_375/A 0.03fF
C20702 OR2X1_LOC_375/A AND2X1_LOC_255/a_8_24# 0.02fF
C22979 AND2X1_LOC_752/a_8_24# OR2X1_LOC_375/A 0.01fF
C24228 AND2X1_LOC_421/a_8_24# OR2X1_LOC_375/A 0.01fF
C25400 AND2X1_LOC_310/a_8_24# OR2X1_LOC_375/A 0.01fF
C25503 AND2X1_LOC_49/a_8_24# OR2X1_LOC_375/A 0.01fF
C25584 AND2X1_LOC_692/a_8_24# OR2X1_LOC_375/A 0.01fF
C28508 AND2X1_LOC_10/a_8_24# OR2X1_LOC_375/A 0.03fF
C28954 AND2X1_LOC_309/a_8_24# OR2X1_LOC_375/A 0.01fF
C29138 OR2X1_LOC_375/A AND2X1_LOC_277/a_8_24# 0.01fF
C30634 AND2X1_LOC_519/a_36_24# OR2X1_LOC_375/A 0.01fF
C31365 OR2X1_LOC_375/A AND2X1_LOC_422/a_8_24# 0.01fF
C31410 AND2X1_LOC_29/a_8_24# OR2X1_LOC_375/A 0.03fF
C31745 AND2X1_LOC_144/a_8_24# OR2X1_LOC_375/A 0.01fF
C33667 AND2X1_LOC_6/a_8_24# OR2X1_LOC_375/A 0.01fF
C36176 AND2X1_LOC_699/a_8_24# OR2X1_LOC_375/A 0.03fF
C36668 OR2X1_LOC_375/A OR2X1_LOC_120/a_8_216# 0.01fF
C38982 AND2X1_LOC_53/a_8_24# OR2X1_LOC_375/A 0.01fF
C42941 AND2X1_LOC_46/a_8_24# OR2X1_LOC_375/A 0.02fF
C43244 OR2X1_LOC_274/a_8_216# OR2X1_LOC_375/A 0.01fF
C43584 AND2X1_LOC_92/a_8_24# OR2X1_LOC_375/A 0.01fF
C43696 AND2X1_LOC_693/a_8_24# OR2X1_LOC_375/A 0.09fF
C43827 AND2X1_LOC_119/a_8_24# OR2X1_LOC_375/A 0.06fF
C45027 AND2X1_LOC_753/a_8_24# OR2X1_LOC_375/A 0.02fF
C46383 OR2X1_LOC_270/a_8_216# OR2X1_LOC_375/A 0.02fF
C51943 OR2X1_LOC_270/a_36_216# OR2X1_LOC_375/A 0.02fF
C53790 OR2X1_LOC_375/A OR2X1_LOC_512/a_8_216# 0.01fF
C55928 OR2X1_LOC_375/A OR2X1_LOC_513/a_8_216# 0.01fF
C2275 OR2X1_LOC_64/Y OR2X1_LOC_762/a_8_216# 0.01fF
C3079 OR2X1_LOC_694/a_8_216# OR2X1_LOC_64/Y 0.01fF
C8714 OR2X1_LOC_64/Y OR2X1_LOC_760/a_8_216# 0.01fF
C8972 OR2X1_LOC_421/a_8_216# OR2X1_LOC_64/Y 0.02fF
C11440 OR2X1_LOC_309/a_8_216# OR2X1_LOC_64/Y 0.06fF
C14014 OR2X1_LOC_329/a_8_216# OR2X1_LOC_64/Y 0.01fF
C14517 OR2X1_LOC_64/Y OR2X1_LOC_71/a_8_216# 0.05fF
C15223 AND2X1_LOC_515/a_8_24# OR2X1_LOC_64/Y 0.07fF
C21816 OR2X1_LOC_682/a_8_216# OR2X1_LOC_64/Y 0.02fF
C30590 OR2X1_LOC_625/a_8_216# OR2X1_LOC_64/Y 0.01fF
C31642 OR2X1_LOC_64/Y OR2X1_LOC_599/a_8_216# 0.01fF
C34356 OR2X1_LOC_692/a_8_216# OR2X1_LOC_64/Y 0.15fF
C35146 OR2X1_LOC_527/a_8_216# OR2X1_LOC_64/Y 0.08fF
C37165 OR2X1_LOC_111/a_8_216# OR2X1_LOC_64/Y 0.01fF
C38656 AND2X1_LOC_598/a_8_24# OR2X1_LOC_64/Y 0.01fF
C46061 OR2X1_LOC_64/Y AND2X1_LOC_685/a_8_24# 0.01fF
C48717 OR2X1_LOC_64/Y OR2X1_LOC_226/a_8_216# 0.01fF
C50450 OR2X1_LOC_64/Y AND2X1_LOC_687/a_8_24# 0.01fF
C52758 OR2X1_LOC_681/a_8_216# OR2X1_LOC_64/Y 0.01fF
C53683 OR2X1_LOC_64/Y OR2X1_LOC_763/a_8_216# 0.01fF
C55292 AND2X1_LOC_596/a_8_24# OR2X1_LOC_64/Y 0.01fF
C55505 OR2X1_LOC_64/Y OR2X1_LOC_85/a_8_216# 0.01fF
C163 OR2X1_LOC_95/Y OR2X1_LOC_760/a_8_216# 0.01fF
C5466 OR2X1_LOC_329/a_8_216# OR2X1_LOC_95/Y 0.01fF
C6753 AND2X1_LOC_515/a_8_24# OR2X1_LOC_95/Y 0.05fF
C9044 OR2X1_LOC_256/a_8_216# OR2X1_LOC_95/Y 0.03fF
C10346 OR2X1_LOC_95/Y AND2X1_LOC_458/a_8_24# 0.04fF
C14569 OR2X1_LOC_256/a_36_216# OR2X1_LOC_95/Y 0.01fF
C17816 AND2X1_LOC_515/a_36_24# OR2X1_LOC_95/Y 0.01fF
C18562 OR2X1_LOC_95/Y OR2X1_LOC_164/a_8_216# 0.02fF
C19233 OR2X1_LOC_529/a_8_216# OR2X1_LOC_95/Y 0.01fF
C20919 OR2X1_LOC_819/a_8_216# OR2X1_LOC_95/Y 0.01fF
C21435 OR2X1_LOC_95/Y OR2X1_LOC_371/a_8_216# 0.03fF
C22604 OR2X1_LOC_672/a_8_216# OR2X1_LOC_95/Y 0.01fF
C23292 OR2X1_LOC_95/Y OR2X1_LOC_599/a_8_216# 0.02fF
C24130 OR2X1_LOC_95/Y OR2X1_LOC_164/a_36_216# 0.02fF
C26476 OR2X1_LOC_95/Y OR2X1_LOC_372/a_8_216# -0.01fF
C27594 OR2X1_LOC_133/a_8_216# OR2X1_LOC_95/Y 0.01fF
C30250 AND2X1_LOC_598/a_8_24# OR2X1_LOC_95/Y 0.01fF
C30359 OR2X1_LOC_95/Y OR2X1_LOC_419/a_8_216# 0.01fF
C31854 OR2X1_LOC_820/A OR2X1_LOC_95/Y 0.17fF
C32317 OR2X1_LOC_95/Y OR2X1_LOC_820/B 0.04fF
C40006 OR2X1_LOC_95/Y OR2X1_LOC_226/a_8_216# -0.00fF
C40852 OR2X1_LOC_95/Y OR2X1_LOC_77/a_8_216# 0.01fF
C43738 OR2X1_LOC_95/Y OR2X1_LOC_323/a_8_216# 0.01fF
C45225 AND2X1_LOC_800/a_8_24# OR2X1_LOC_95/Y 0.01fF
C46345 OR2X1_LOC_95/Y AND2X1_LOC_407/a_8_24# 0.01fF
C49030 OR2X1_LOC_90/a_8_216# OR2X1_LOC_95/Y 0.01fF
C49990 OR2X1_LOC_73/a_8_216# OR2X1_LOC_95/Y 0.01fF
C50083 OR2X1_LOC_95/Y OR2X1_LOC_749/a_8_216# 0.01fF
C50877 AND2X1_LOC_801/B OR2X1_LOC_95/Y 0.01fF
C55987 OR2X1_LOC_95/Y OR2X1_LOC_387/a_8_216# 0.01fF
C4900 AND2X1_LOC_513/a_8_24# OR2X1_LOC_51/Y 0.08fF
C5395 OR2X1_LOC_51/Y OR2X1_LOC_93/a_8_216# 0.01fF
C6195 OR2X1_LOC_51/Y OR2X1_LOC_46/a_8_216# 0.01fF
C6694 OR2X1_LOC_51/Y OR2X1_LOC_22/a_8_216# 0.01fF
C7202 OR2X1_LOC_51/Y AND2X1_LOC_685/a_8_24# 0.05fF
C9973 OR2X1_LOC_144/a_8_216# OR2X1_LOC_51/Y 0.14fF
C10147 OR2X1_LOC_283/a_8_216# OR2X1_LOC_51/Y 0.01fF
C11547 OR2X1_LOC_51/Y AND2X1_LOC_687/a_8_24# 0.01fF
C13049 OR2X1_LOC_328/a_8_216# OR2X1_LOC_51/Y 0.01fF
C13869 OR2X1_LOC_681/a_8_216# OR2X1_LOC_51/Y 0.01fF
C15586 OR2X1_LOC_51/Y OR2X1_LOC_40/a_8_216# 0.01fF
C20314 OR2X1_LOC_694/a_8_216# OR2X1_LOC_51/Y 0.01fF
C24632 OR2X1_LOC_51/Y OR2X1_LOC_3/a_8_216# 0.01fF
C25401 OR2X1_LOC_51/Y OR2X1_LOC_48/a_8_216# 0.06fF
C28600 OR2X1_LOC_51/Y OR2X1_LOC_386/a_8_216# 0.01fF
C30866 AND2X1_LOC_155/a_8_24# OR2X1_LOC_51/Y 0.06fF
C34647 OR2X1_LOC_51/Y OR2X1_LOC_256/a_8_216# 0.05fF
C35354 OR2X1_LOC_51/Y OR2X1_LOC_18/a_8_216# 0.01fF
C38075 OR2X1_LOC_51/Y OR2X1_LOC_47/a_8_216# 0.01fF
C39798 OR2X1_LOC_51/Y OR2X1_LOC_6/a_8_216# 0.01fF
C41097 OR2X1_LOC_51/Y OR2X1_LOC_681/Y 0.01fF
C41651 OR2X1_LOC_51/Y OR2X1_LOC_289/a_8_216# 0.02fF
C42234 AND2X1_LOC_410/a_8_24# OR2X1_LOC_51/Y 0.01fF
C44221 OR2X1_LOC_51/Y OR2X1_LOC_411/a_8_216# 0.01fF
C48048 OR2X1_LOC_51/Y OR2X1_LOC_625/a_8_216# 0.01fF
C49228 OR2X1_LOC_51/Y OR2X1_LOC_12/a_8_216# 0.01fF
C49253 OR2X1_LOC_51/Y OR2X1_LOC_425/a_8_216# 0.39fF
C49267 AND2X1_LOC_374/a_8_24# OR2X1_LOC_51/Y 0.02fF
C49680 OR2X1_LOC_51/Y OR2X1_LOC_743/a_8_216# 0.01fF
C52899 OR2X1_LOC_51/Y OR2X1_LOC_534/a_8_216# 0.02fF
C10307 OR2X1_LOC_635/A AND2X1_LOC_684/a_8_24# 0.04fF
C29281 OR2X1_LOC_635/A AND2X1_LOC_683/a_8_24# 0.02fF
C45924 OR2X1_LOC_635/A AND2X1_LOC_683/a_36_24# 0.01fF
C18246 AND2X1_LOC_753/a_8_24# OR2X1_LOC_790/B 0.01fF
C455 AND2X1_LOC_47/Y AND2X1_LOC_819/a_8_24# 0.10fF
C1422 AND2X1_LOC_47/Y AND2X1_LOC_18/a_8_24# 0.01fF
C2075 AND2X1_LOC_47/Y OR2X1_LOC_120/a_8_216# 0.04fF
C2287 AND2X1_LOC_85/a_8_24# AND2X1_LOC_47/Y 0.01fF
C2555 AND2X1_LOC_47/Y AND2X1_LOC_263/a_8_24# 0.01fF
C5128 AND2X1_LOC_328/a_8_24# AND2X1_LOC_47/Y 0.01fF
C5965 AND2X1_LOC_306/a_8_24# AND2X1_LOC_47/Y 0.07fF
C8114 AND2X1_LOC_95/a_8_24# AND2X1_LOC_47/Y 0.01fF
C8920 AND2X1_LOC_92/a_8_24# AND2X1_LOC_47/Y 0.01fF
C14460 AND2X1_LOC_47/Y AND2X1_LOC_417/a_36_24# 0.01fF
C14579 AND2X1_LOC_153/a_8_24# AND2X1_LOC_47/Y 0.03fF
C15471 OR2X1_LOC_276/B AND2X1_LOC_47/Y 0.08fF
C16948 AND2X1_LOC_47/Y AND2X1_LOC_273/a_8_24# 0.02fF
C17878 AND2X1_LOC_47/Y AND2X1_LOC_628/a_8_24# 0.03fF
C18416 AND2X1_LOC_47/Y AND2X1_LOC_234/a_8_24# 0.01fF
C18481 AND2X1_LOC_672/a_8_24# AND2X1_LOC_47/Y 0.02fF
C23128 AND2X1_LOC_102/a_8_24# AND2X1_LOC_47/Y 0.01fF
C24001 AND2X1_LOC_31/a_8_24# AND2X1_LOC_47/Y 0.19fF
C24208 AND2X1_LOC_47/Y AND2X1_LOC_760/a_8_24# 0.07fF
C24967 AND2X1_LOC_47/Y OR2X1_LOC_374/a_8_216# 0.01fF
C26374 AND2X1_LOC_71/a_8_24# AND2X1_LOC_47/Y 0.10fF
C26868 AND2X1_LOC_26/a_8_24# AND2X1_LOC_47/Y 0.01fF
C27666 AND2X1_LOC_304/a_8_24# AND2X1_LOC_47/Y 0.01fF
C27692 AND2X1_LOC_59/a_8_24# AND2X1_LOC_47/Y 0.01fF
C28515 AND2X1_LOC_48/a_8_24# AND2X1_LOC_47/Y 0.05fF
C30225 AND2X1_LOC_104/a_8_24# AND2X1_LOC_47/Y 0.02fF
C31447 AND2X1_LOC_372/a_8_24# AND2X1_LOC_47/Y 0.03fF
C32322 AND2X1_LOC_386/a_8_24# AND2X1_LOC_47/Y 0.01fF
C36021 AND2X1_LOC_90/a_8_24# AND2X1_LOC_47/Y 0.02fF
C37145 AND2X1_LOC_47/Y OR2X1_LOC_515/a_8_216# 0.02fF
C38620 AND2X1_LOC_164/a_8_24# AND2X1_LOC_47/Y 0.01fF
C39022 AND2X1_LOC_93/a_8_24# AND2X1_LOC_47/Y 0.03fF
C40385 AND2X1_LOC_159/a_8_24# AND2X1_LOC_47/Y 0.02fF
C42754 AND2X1_LOC_47/Y OR2X1_LOC_515/a_36_216# 0.02fF
C44523 AND2X1_LOC_47/Y AND2X1_LOC_762/a_8_24# 0.01fF
C44738 AND2X1_LOC_43/a_8_24# AND2X1_LOC_47/Y 0.01fF
C49833 AND2X1_LOC_47/Y AND2X1_LOC_433/a_8_24# 0.01fF
C50058 AND2X1_LOC_47/Y AND2X1_LOC_8/a_8_24# 0.09fF
C50675 AND2X1_LOC_47/Y AND2X1_LOC_277/a_8_24# 0.04fF
C51647 AND2X1_LOC_38/a_8_24# AND2X1_LOC_47/Y 0.02fF
C54011 AND2X1_LOC_47/Y AND2X1_LOC_417/a_8_24# 0.04fF
C55761 AND2X1_LOC_511/a_8_24# AND2X1_LOC_47/Y 0.01fF
C272 AND2X1_LOC_696/a_8_24# AND2X1_LOC_44/Y 0.01fF
C284 AND2X1_LOC_19/a_8_24# AND2X1_LOC_44/Y 0.05fF
C678 AND2X1_LOC_29/a_8_24# AND2X1_LOC_44/Y 0.01fF
C1965 AND2X1_LOC_699/a_36_24# AND2X1_LOC_44/Y -0.02fF
C5505 AND2X1_LOC_699/a_8_24# AND2X1_LOC_44/Y -0.01fF
C6096 AND2X1_LOC_387/a_36_24# AND2X1_LOC_44/Y 0.01fF
C6341 AND2X1_LOC_44/Y AND2X1_LOC_761/a_36_24# 0.02fF
C7971 AND2X1_LOC_412/a_8_24# AND2X1_LOC_44/Y 0.02fF
C12254 AND2X1_LOC_46/a_8_24# AND2X1_LOC_44/Y 0.01fF
C12960 AND2X1_LOC_40/a_8_24# AND2X1_LOC_44/Y 0.01fF
C17174 OR2X1_LOC_596/a_8_216# AND2X1_LOC_44/Y 0.16fF
C17666 AND2X1_LOC_129/a_8_24# AND2X1_LOC_44/Y 0.01fF
C23047 AND2X1_LOC_44/Y OR2X1_LOC_512/a_8_216# 0.01fF
C25139 AND2X1_LOC_44/Y OR2X1_LOC_513/a_8_216# 0.01fF
C26661 AND2X1_LOC_136/a_8_24# AND2X1_LOC_44/Y 0.02fF
C27399 AND2X1_LOC_749/a_8_24# AND2X1_LOC_44/Y 0.03fF
C27951 AND2X1_LOC_31/a_8_24# AND2X1_LOC_44/Y 0.02fF
C30358 AND2X1_LOC_71/a_8_24# AND2X1_LOC_44/Y 0.01fF
C32474 OR2X1_LOC_87/a_8_216# AND2X1_LOC_44/Y 0.01fF
C33459 AND2X1_LOC_133/a_8_24# AND2X1_LOC_44/Y 0.07fF
C36340 AND2X1_LOC_386/a_8_24# AND2X1_LOC_44/Y 0.17fF
C41779 AND2X1_LOC_70/a_8_24# AND2X1_LOC_44/Y 0.01fF
C43988 AND2X1_LOC_749/a_36_24# AND2X1_LOC_44/Y 0.01fF
C44468 AND2X1_LOC_159/a_8_24# AND2X1_LOC_44/Y 0.01fF
C45718 AND2X1_LOC_57/a_8_24# AND2X1_LOC_44/Y 0.03fF
C47975 AND2X1_LOC_22/a_8_24# AND2X1_LOC_44/Y 0.02fF
C49657 AND2X1_LOC_421/a_8_24# AND2X1_LOC_44/Y 0.01fF
C50944 AND2X1_LOC_47/a_8_24# AND2X1_LOC_44/Y 0.02fF
C51044 AND2X1_LOC_692/a_8_24# AND2X1_LOC_44/Y 0.01fF
C51270 AND2X1_LOC_387/a_8_24# AND2X1_LOC_44/Y 0.03fF
C51536 AND2X1_LOC_44/Y AND2X1_LOC_761/a_8_24# 0.04fF
C1021 AND2X1_LOC_47/a_8_24# AND2X1_LOC_31/Y 0.01fF
C3917 AND2X1_LOC_31/Y AND2X1_LOC_433/a_8_24# 0.01fF
C6492 AND2X1_LOC_696/a_8_24# AND2X1_LOC_31/Y 0.01fF
C9231 AND2X1_LOC_684/a_8_24# AND2X1_LOC_31/Y 0.01fF
C9897 AND2X1_LOC_511/a_8_24# AND2X1_LOC_31/Y 0.01fF
C16257 AND2X1_LOC_306/a_8_24# AND2X1_LOC_31/Y 0.01fF
C19210 AND2X1_LOC_40/a_8_24# AND2X1_LOC_31/Y 0.01fF
C23989 AND2X1_LOC_682/a_8_24# AND2X1_LOC_31/Y 0.01fF
C25926 AND2X1_LOC_31/Y AND2X1_LOC_226/a_8_24# 0.01fF
C28226 AND2X1_LOC_683/a_8_24# AND2X1_LOC_31/Y 0.01fF
C28544 AND2X1_LOC_371/a_8_24# AND2X1_LOC_31/Y 0.04fF
C32389 OR2X1_LOC_688/a_8_216# AND2X1_LOC_31/Y 0.11fF
C34143 AND2X1_LOC_31/a_8_24# AND2X1_LOC_31/Y 0.02fF
C37828 AND2X1_LOC_304/a_8_24# AND2X1_LOC_31/Y 0.01fF
C38227 OR2X1_LOC_686/A AND2X1_LOC_31/Y 0.02fF
C41703 AND2X1_LOC_372/a_8_24# AND2X1_LOC_31/Y 0.01fF
C47776 AND2X1_LOC_31/Y OR2X1_LOC_375/a_8_216# 0.01fF
C48287 AND2X1_LOC_70/a_8_24# AND2X1_LOC_31/Y 0.01fF
C49093 AND2X1_LOC_164/a_8_24# AND2X1_LOC_31/Y 0.01fF
C51294 AND2X1_LOC_689/a_8_24# AND2X1_LOC_31/Y 0.01fF
C53382 AND2X1_LOC_31/Y OR2X1_LOC_68/a_8_216# 0.03fF
C54175 AND2X1_LOC_22/a_8_24# AND2X1_LOC_31/Y 0.01fF
C54592 AND2X1_LOC_752/a_8_24# AND2X1_LOC_31/Y 0.01fF
C54657 OR2X1_LOC_688/Y AND2X1_LOC_31/Y 0.11fF
C55890 OR2X1_LOC_458/a_8_216# AND2X1_LOC_31/Y 0.01fF
C3594 AND2X1_LOC_681/a_8_24# AND2X1_LOC_51/Y 0.01fF
C5047 AND2X1_LOC_144/a_8_24# AND2X1_LOC_51/Y 0.01fF
C6938 AND2X1_LOC_684/a_8_24# AND2X1_LOC_51/Y 0.01fF
C7599 AND2X1_LOC_511/a_8_24# AND2X1_LOC_51/Y 0.06fF
C16100 AND2X1_LOC_95/a_8_24# AND2X1_LOC_51/Y 0.17fF
C16955 AND2X1_LOC_40/a_8_24# AND2X1_LOC_51/Y 0.01fF
C21777 AND2X1_LOC_682/a_8_24# AND2X1_LOC_51/Y 0.01fF
C23102 AND2X1_LOC_329/a_8_24# AND2X1_LOC_51/Y 0.02fF
C26002 AND2X1_LOC_683/a_8_24# AND2X1_LOC_51/Y 0.01fF
C29064 AND2X1_LOC_51/Y OR2X1_LOC_513/a_8_216# 0.02fF
C31924 AND2X1_LOC_31/a_8_24# AND2X1_LOC_51/Y 0.01fF
C34541 AND2X1_LOC_51/Y OR2X1_LOC_513/a_36_216# 0.02fF
C35991 OR2X1_LOC_686/A AND2X1_LOC_51/Y 0.01fF
C37248 AND2X1_LOC_51/Y AND2X1_LOC_625/a_8_24# 0.02fF
C39080 OR2X1_LOC_407/a_8_216# AND2X1_LOC_51/Y 0.14fF
C39101 AND2X1_LOC_44/a_8_24# AND2X1_LOC_51/Y 0.01fF
C43901 AND2X1_LOC_15/a_8_24# AND2X1_LOC_51/Y 0.01fF
C45911 AND2X1_LOC_70/a_8_24# AND2X1_LOC_51/Y 0.04fF
C46762 OR2X1_LOC_691/a_8_216# AND2X1_LOC_51/Y 0.01fF
C46831 AND2X1_LOC_164/a_8_24# AND2X1_LOC_51/Y 0.15fF
C51178 AND2X1_LOC_51/Y OR2X1_LOC_68/a_8_216# 0.01fF
C51973 AND2X1_LOC_22/a_8_24# AND2X1_LOC_51/Y 0.01fF
C53541 AND2X1_LOC_587/a_8_24# AND2X1_LOC_51/Y 0.20fF
C54930 AND2X1_LOC_47/a_8_24# AND2X1_LOC_51/Y 0.01fF
C682 OR2X1_LOC_40/Y OR2X1_LOC_291/a_8_216# 0.01fF
C3785 OR2X1_LOC_40/Y OR2X1_LOC_3/a_8_216# 0.40fF
C4451 OR2X1_LOC_40/Y AND2X1_LOC_514/a_8_24# 0.02fF
C7797 OR2X1_LOC_40/Y OR2X1_LOC_386/a_8_216# 0.03fF
C7857 OR2X1_LOC_40/Y OR2X1_LOC_309/a_8_216# 0.01fF
C11890 OR2X1_LOC_40/Y AND2X1_LOC_814/a_8_24# 0.01fF
C12281 OR2X1_LOC_40/Y OR2X1_LOC_278/a_8_216# 0.01fF
C14657 OR2X1_LOC_40/Y OR2X1_LOC_18/a_8_216# 0.01fF
C15988 OR2X1_LOC_519/a_8_216# OR2X1_LOC_40/Y 0.01fF
C19051 OR2X1_LOC_40/Y OR2X1_LOC_6/a_8_216# 0.01fF
C24881 OR2X1_LOC_40/Y OR2X1_LOC_129/a_8_216# 0.01fF
C25789 OR2X1_LOC_40/Y AND2X1_LOC_87/a_8_24# 0.02fF
C28037 OR2X1_LOC_40/Y OR2X1_LOC_225/a_8_216# 0.01fF
C28268 OR2X1_LOC_40/Y OR2X1_LOC_12/a_8_216# 0.01fF
C35511 OR2X1_LOC_40/Y OR2X1_LOC_246/a_8_216# 0.14fF
C38059 OR2X1_LOC_40/Y AND2X1_LOC_548/a_8_24# 0.17fF
C39413 OR2X1_LOC_40/Y OR2X1_LOC_277/a_8_216# 0.06fF
C40611 OR2X1_LOC_40/Y OR2X1_LOC_93/a_8_216# 0.01fF
C50869 OR2X1_LOC_136/a_8_216# OR2X1_LOC_40/Y 0.01fF
C51312 OR2X1_LOC_369/a_8_216# OR2X1_LOC_40/Y 0.02fF
C54203 OR2X1_LOC_40/Y OR2X1_LOC_310/a_8_216# 0.01fF
C498 OR2X1_LOC_3/Y OR2X1_LOC_119/a_8_216# 0.01fF
C1272 OR2X1_LOC_3/Y AND2X1_LOC_377/Y 0.16fF
C1754 OR2X1_LOC_694/a_8_216# OR2X1_LOC_3/Y 0.02fF
C2466 OR2X1_LOC_136/a_36_216# OR2X1_LOC_3/Y 0.04fF
C6743 OR2X1_LOC_3/Y AND2X1_LOC_378/a_8_24# 0.17fF
C6826 OR2X1_LOC_3/Y OR2X1_LOC_48/a_8_216# 0.05fF
C7133 OR2X1_LOC_820/a_8_216# OR2X1_LOC_3/Y 0.01fF
C7629 OR2X1_LOC_3/Y OR2X1_LOC_421/a_8_216# 0.05fF
C8125 OR2X1_LOC_3/Y AND2X1_LOC_94/a_8_24# 0.01fF
C9749 OR2X1_LOC_3/Y OR2X1_LOC_382/a_8_216# 0.06fF
C10048 OR2X1_LOC_3/Y OR2X1_LOC_386/a_8_216# 0.02fF
C10512 OR2X1_LOC_3/Y OR2X1_LOC_56/a_8_216# 0.01fF
C10736 OR2X1_LOC_3/Y OR2X1_LOC_817/a_8_216# 0.01fF
C12682 OR2X1_LOC_3/Y OR2X1_LOC_381/a_8_216# 0.11fF
C14180 OR2X1_LOC_3/Y AND2X1_LOC_814/a_8_24# 0.01fF
C16888 OR2X1_LOC_3/Y OR2X1_LOC_18/a_8_216# 0.01fF
C17526 OR2X1_LOC_3/Y AND2X1_LOC_66/a_8_24# 0.01fF
C20495 OR2X1_LOC_682/a_8_216# OR2X1_LOC_3/Y 0.02fF
C22708 OR2X1_LOC_3/Y OR2X1_LOC_681/Y 0.04fF
C29307 OR2X1_LOC_3/Y OR2X1_LOC_625/a_8_216# 0.14fF
C30262 OR2X1_LOC_3/Y OR2X1_LOC_225/a_8_216# 0.01fF
C30512 OR2X1_LOC_3/Y OR2X1_LOC_12/a_8_216# 0.37fF
C34522 OR2X1_LOC_3/Y OR2X1_LOC_377/a_8_216# 0.02fF
C39003 OR2X1_LOC_3/Y OR2X1_LOC_820/A 0.02fF
C39513 OR2X1_LOC_3/Y OR2X1_LOC_820/B 0.05fF
C41088 OR2X1_LOC_3/Y AND2X1_LOC_121/a_8_24# 0.01fF
C41218 OR2X1_LOC_3/Y OR2X1_LOC_273/a_8_216# 0.05fF
C41682 OR2X1_LOC_3/Y OR2X1_LOC_277/a_8_216# 0.01fF
C42745 OR2X1_LOC_3/Y OR2X1_LOC_748/a_8_216# 0.01fF
C42980 OR2X1_LOC_3/Y AND2X1_LOC_847/a_8_24# 0.01fF
C44638 OR2X1_LOC_3/Y AND2X1_LOC_398/a_8_24# 0.01fF
C44710 OR2X1_LOC_3/Y AND2X1_LOC_685/a_8_24# 0.01fF
C45681 OR2X1_LOC_3/Y OR2X1_LOC_377/a_36_216# 0.03fF
C46913 OR2X1_LOC_3/Y OR2X1_LOC_272/a_8_216# 0.01fF
C49131 OR2X1_LOC_3/Y AND2X1_LOC_687/a_8_24# 0.01fF
C50673 OR2X1_LOC_328/a_8_216# OR2X1_LOC_3/Y 0.02fF
C51273 OR2X1_LOC_3/Y OR2X1_LOC_88/a_8_216# 0.01fF
C51451 OR2X1_LOC_681/a_8_216# OR2X1_LOC_3/Y 0.01fF
C53090 OR2X1_LOC_136/a_8_216# OR2X1_LOC_3/Y 0.04fF
C53733 OR2X1_LOC_126/a_8_216# OR2X1_LOC_3/Y 0.01fF
C55197 OR2X1_LOC_304/a_8_216# OR2X1_LOC_3/Y 0.01fF
C55231 OR2X1_LOC_490/a_8_216# OR2X1_LOC_3/Y 0.01fF
C1445 OR2X1_LOC_70/Y OR2X1_LOC_760/a_8_216# 0.14fF
C10777 OR2X1_LOC_70/Y AND2X1_LOC_686/a_8_24# 0.02fF
C13334 OR2X1_LOC_70/Y OR2X1_LOC_245/a_8_216# 0.01fF
C13530 OR2X1_LOC_70/Y OR2X1_LOC_373/a_8_216# 0.01fF
C17772 OR2X1_LOC_70/Y OR2X1_LOC_684/a_8_216# 0.02fF
C17941 OR2X1_LOC_70/Y OR2X1_LOC_430/a_8_216# 0.02fF
C23186 OR2X1_LOC_70/Y AND2X1_LOC_405/a_8_24# 0.01fF
C25037 OR2X1_LOC_70/Y OR2X1_LOC_582/a_8_216# 0.40fF
C28238 OR2X1_LOC_70/Y OR2X1_LOC_534/a_8_216# 0.01fF
C31552 OR2X1_LOC_70/Y OR2X1_LOC_426/a_8_216# 0.02fF
C33609 OR2X1_LOC_70/Y OR2X1_LOC_433/a_8_216# 0.08fF
C35689 OR2X1_LOC_70/Y AND2X1_LOC_100/a_8_24# 0.02fF
C37786 OR2X1_LOC_70/Y OR2X1_LOC_86/a_8_216# 0.15fF
C43030 OR2X1_LOC_70/Y OR2X1_LOC_70/a_8_216# -0.00fF
C43048 OR2X1_LOC_70/Y AND2X1_LOC_687/a_8_24# 0.26fF
C47315 OR2X1_LOC_683/a_8_216# OR2X1_LOC_70/Y 0.02fF
C49305 OR2X1_LOC_304/a_8_216# OR2X1_LOC_70/Y 0.01fF
C49340 OR2X1_LOC_490/a_8_216# OR2X1_LOC_70/Y 0.02fF
C263 OR2X1_LOC_158/A AND2X1_LOC_375/a_36_24# 0.01fF
C4303 OR2X1_LOC_158/A OR2X1_LOC_588/a_8_216# 0.05fF
C4964 OR2X1_LOC_158/A OR2X1_LOC_824/a_8_216# 0.14fF
C5126 OR2X1_LOC_158/A OR2X1_LOC_153/a_8_216# 0.01fF
C5853 OR2X1_LOC_158/A OR2X1_LOC_488/a_8_216# 0.02fF
C7674 OR2X1_LOC_158/A OR2X1_LOC_51/a_8_216# 0.02fF
C8322 OR2X1_LOC_158/A OR2X1_LOC_672/a_8_216# 0.03fF
C9609 OR2X1_LOC_158/A OR2X1_LOC_743/a_8_216# 0.01fF
C11426 OR2X1_LOC_158/A OR2X1_LOC_488/a_36_216# 0.03fF
C11813 OR2X1_LOC_158/A OR2X1_LOC_271/Y 0.11fF
C12124 OR2X1_LOC_158/A AND2X1_LOC_296/a_8_24# 0.02fF
C12660 OR2X1_LOC_158/A AND2X1_LOC_818/a_8_24# 0.02fF
C13405 OR2X1_LOC_133/a_8_216# OR2X1_LOC_158/A 0.02fF
C14625 OR2X1_LOC_111/a_8_216# OR2X1_LOC_158/A 0.03fF
C15962 OR2X1_LOC_158/A OR2X1_LOC_689/a_8_216# 0.01fF
C18173 OR2X1_LOC_158/A OR2X1_LOC_820/B 0.05fF
C20161 OR2X1_LOC_111/a_36_216# OR2X1_LOC_158/A 0.02fF
C21188 OR2X1_LOC_158/A AND2X1_LOC_264/a_8_24# 0.01fF
C21567 OR2X1_LOC_158/A OR2X1_LOC_689/a_36_216# 0.01fF
C21922 OR2X1_LOC_159/a_8_216# OR2X1_LOC_158/A 0.02fF
C22086 OR2X1_LOC_158/A OR2X1_LOC_44/a_8_216# 0.02fF
C22471 OR2X1_LOC_158/A OR2X1_LOC_236/a_8_216# 0.01fF
C23397 OR2X1_LOC_158/A AND2X1_LOC_685/a_8_24# 0.02fF
C25910 OR2X1_LOC_158/A OR2X1_LOC_55/a_8_216# 0.02fF
C26723 OR2X1_LOC_158/A OR2X1_LOC_77/a_8_216# 0.02fF
C27521 OR2X1_LOC_158/A OR2X1_LOC_44/a_36_216# 0.02fF
C27581 OR2X1_LOC_158/A OR2X1_LOC_412/a_8_216# 0.02fF
C34166 OR2X1_LOC_158/A AND2X1_LOC_276/a_8_24# 0.03fF
C34187 OR2X1_LOC_158/A AND2X1_LOC_375/a_8_24# 0.06fF
C34557 OR2X1_LOC_158/A OR2X1_LOC_90/a_8_216# 0.02fF
C34972 OR2X1_LOC_158/A OR2X1_LOC_310/a_8_216# 0.01fF
C35481 OR2X1_LOC_157/a_8_216# OR2X1_LOC_158/A 0.01fF
C35529 OR2X1_LOC_158/A OR2X1_LOC_73/a_8_216# 0.02fF
C36284 OR2X1_LOC_158/A OR2X1_LOC_422/a_8_216# 0.01fF
C41304 OR2X1_LOC_158/A OR2X1_LOC_9/a_8_216# 0.15fF
C42240 OR2X1_LOC_158/A OR2X1_LOC_421/a_8_216# 0.01fF
C44380 OR2X1_LOC_158/A OR2X1_LOC_382/a_8_216# 0.01fF
C45207 OR2X1_LOC_158/A OR2X1_LOC_56/a_8_216# 0.02fF
C47111 OR2X1_LOC_158/A AND2X1_LOC_155/a_8_24# 0.01fF
C47489 OR2X1_LOC_158/A OR2X1_LOC_381/a_8_216# 0.02fF
C48121 OR2X1_LOC_158/A OR2X1_LOC_275/a_8_216# 0.02fF
C48485 OR2X1_LOC_158/A OR2X1_LOC_699/a_8_216# 0.02fF
C50557 OR2X1_LOC_158/A OR2X1_LOC_94/a_8_216# 0.02fF
C51496 OR2X1_LOC_158/A OR2X1_LOC_54/a_8_216# 0.02fF
C52722 OR2X1_LOC_158/A AND2X1_LOC_120/a_8_24# 0.01fF
C53069 OR2X1_LOC_519/a_8_216# OR2X1_LOC_158/A 0.01fF
C53536 OR2X1_LOC_158/A OR2X1_LOC_42/a_8_216# 0.01fF
C55217 OR2X1_LOC_682/a_8_216# OR2X1_LOC_158/A 0.01fF
C55586 OR2X1_LOC_158/A AND2X1_LOC_274/a_8_24# 0.01fF
C47127 OR2X1_LOC_597/A OR2X1_LOC_692/a_8_216# 0.47fF
C17428 AND2X1_LOC_382/a_8_24# OR2X1_LOC_391/B 0.01fF
C5479 OR2X1_LOC_276/a_36_216# OR2X1_LOC_549/A 0.01fF
C8325 AND2X1_LOC_625/a_8_24# OR2X1_LOC_549/A 0.04fF
C14932 OR2X1_LOC_66/a_8_216# OR2X1_LOC_549/A 0.06fF
C20456 AND2X1_LOC_271/a_8_24# OR2X1_LOC_549/A 0.01fF
C25779 AND2X1_LOC_49/a_8_24# OR2X1_LOC_549/A 0.01fF
C32490 OR2X1_LOC_269/a_8_216# OR2X1_LOC_549/A 0.01fF
C33966 AND2X1_LOC_6/a_8_24# OR2X1_LOC_549/A 0.06fF
C38236 AND2X1_LOC_268/a_8_24# OR2X1_LOC_549/A 0.02fF
C46683 OR2X1_LOC_270/a_8_216# OR2X1_LOC_549/A 0.01fF
C49533 OR2X1_LOC_269/A OR2X1_LOC_549/A 0.02fF
C50713 OR2X1_LOC_276/B OR2X1_LOC_549/A 1.56fF
C52097 AND2X1_LOC_256/a_8_24# OR2X1_LOC_549/A 0.01fF
C53015 AND2X1_LOC_628/a_8_24# OR2X1_LOC_549/A 0.02fF
C53834 AND2X1_LOC_275/a_8_24# OR2X1_LOC_549/A 0.04fF
C56213 OR2X1_LOC_276/a_8_216# OR2X1_LOC_549/A 0.05fF
C4014 AND2X1_LOC_421/a_8_24# OR2X1_LOC_777/B 0.17fF
C30034 OR2X1_LOC_276/B OR2X1_LOC_777/B 0.07fF
C48200 OR2X1_LOC_777/B AND2X1_LOC_246/a_8_24# 0.20fF
C259 AND2X1_LOC_82/a_8_24# OR2X1_LOC_633/A 0.03fF
C34179 OR2X1_LOC_633/A AND2X1_LOC_278/a_8_24# 0.04fF
C36377 AND2X1_LOC_77/a_8_24# OR2X1_LOC_633/A 0.04fF
C37022 AND2X1_LOC_277/a_8_24# OR2X1_LOC_633/A 0.04fF
C41592 AND2X1_LOC_6/a_8_24# OR2X1_LOC_633/A 0.01fF
C45274 AND2X1_LOC_529/a_8_24# OR2X1_LOC_633/A 0.01fF
C48343 OR2X1_LOC_633/A AND2X1_LOC_277/a_36_24# 0.01fF
C52815 AND2X1_LOC_6/a_36_24# OR2X1_LOC_633/A 0.01fF
C12887 OR2X1_LOC_276/B OR2X1_LOC_541/B 0.01fF
C39273 OR2X1_LOC_541/B AND2X1_LOC_255/a_8_24# 0.01fF
C6336 OR2X1_LOC_634/A AND2X1_LOC_119/a_36_24# 0.01fF
C13532 OR2X1_LOC_634/A AND2X1_LOC_690/a_8_24# 0.11fF
C39377 OR2X1_LOC_634/A AND2X1_LOC_291/a_8_24# 0.02fF
C46326 OR2X1_LOC_634/A AND2X1_LOC_412/a_8_24# 0.01fF
C50635 OR2X1_LOC_634/A AND2X1_LOC_291/a_36_24# 0.02fF
C21547 OR2X1_LOC_130/A AND2X1_LOC_226/a_8_24# 0.03fF
C43574 OR2X1_LOC_130/A AND2X1_LOC_226/a_36_24# 0.01fF
C980 OR2X1_LOC_154/A OR2X1_LOC_276/B 0.10fF
C2886 OR2X1_LOC_154/A OR2X1_LOC_514/a_8_216# 0.03fF
C7687 OR2X1_LOC_154/A OR2X1_LOC_688/a_8_216# 0.01fF
C8080 OR2X1_LOC_154/A OR2X1_LOC_405/a_8_216# 0.02fF
C8164 OR2X1_LOC_154/A AND2X1_LOC_136/a_8_24# 0.02fF
C21409 OR2X1_LOC_154/A AND2X1_LOC_15/a_8_24# 0.07fF
C22814 OR2X1_LOC_154/A OR2X1_LOC_515/a_8_216# 0.03fF
C25929 OR2X1_LOC_154/A AND2X1_LOC_159/a_8_24# 0.16fF
C26385 OR2X1_LOC_154/A AND2X1_LOC_689/a_8_24# 0.01fF
C27176 OR2X1_LOC_154/A AND2X1_LOC_57/a_8_24# 0.03fF
C28489 OR2X1_LOC_154/A OR2X1_LOC_68/a_8_216# 0.01fF
C29773 OR2X1_LOC_154/A OR2X1_LOC_688/Y 0.01fF
C30996 OR2X1_LOC_154/A AND2X1_LOC_272/a_8_24# 0.05fF
C32140 OR2X1_LOC_154/A AND2X1_LOC_310/a_8_24# 0.01fF
C39432 OR2X1_LOC_154/A AND2X1_LOC_699/a_36_24# 0.01fF
C43037 OR2X1_LOC_154/A AND2X1_LOC_699/a_8_24# 0.04fF
C43567 OR2X1_LOC_154/A OR2X1_LOC_120/a_8_216# 0.20fF
C48355 OR2X1_LOC_154/A AND2X1_LOC_419/a_8_24# 0.02fF
C55693 OR2X1_LOC_154/A OR2X1_LOC_274/a_36_216# 0.03fF
C56206 OR2X1_LOC_154/A AND2X1_LOC_153/a_8_24# 0.01fF
C8083 OR2X1_LOC_160/A AND2X1_LOC_129/a_8_24# 0.01fF
C9425 OR2X1_LOC_160/A AND2X1_LOC_329/a_8_24# 0.03fF
C10031 OR2X1_LOC_160/A AND2X1_LOC_226/a_8_24# 0.03fF
C12622 OR2X1_LOC_155/a_8_216# OR2X1_LOC_160/A 0.02fF
C20775 OR2X1_LOC_160/A AND2X1_LOC_71/a_8_24# 0.04fF
C23014 OR2X1_LOC_160/A OR2X1_LOC_87/a_8_216# 0.01fF
C24401 OR2X1_LOC_160/A OR2X1_LOC_398/a_8_216# 0.01fF
C32930 AND2X1_LOC_585/a_8_24# OR2X1_LOC_160/A -0.00fF
C34802 OR2X1_LOC_160/A AND2X1_LOC_159/a_8_24# 0.01fF
C38613 OR2X1_LOC_160/A OR2X1_LOC_688/Y 0.10fF
C44024 AND2X1_LOC_585/a_36_24# OR2X1_LOC_160/A 0.02fF
C46859 OR2X1_LOC_160/A AND2X1_LOC_19/a_8_24# 0.01fF
C50977 OR2X1_LOC_160/A AND2X1_LOC_86/a_8_24# 0.01fF
C51373 OR2X1_LOC_160/A OR2X1_LOC_185/a_8_216# 0.02fF
C9480 AND2X1_LOC_86/B AND2X1_LOC_490/a_8_24# 0.04fF
C46014 AND2X1_LOC_86/B AND2X1_LOC_38/a_8_24# 0.20fF
C51030 AND2X1_LOC_86/B AND2X1_LOC_86/a_8_24# 0.06fF
C52868 AND2X1_LOC_85/a_8_24# AND2X1_LOC_86/B 0.01fF
C7091 OR2X1_LOC_185/A AND2X1_LOC_86/a_36_24# 0.01fF
C8855 AND2X1_LOC_73/a_8_24# OR2X1_LOC_185/A 0.02fF
C9323 OR2X1_LOC_185/A AND2X1_LOC_529/a_36_24# 0.01fF
C10213 OR2X1_LOC_185/A AND2X1_LOC_153/a_8_24# 0.01fF
C21216 OR2X1_LOC_185/A AND2X1_LOC_126/a_8_24# 0.03fF
C25161 OR2X1_LOC_185/A AND2X1_LOC_133/a_8_24# 0.02fF
C25646 OR2X1_LOC_185/A OR2X1_LOC_398/a_8_216# 0.02fF
C32153 OR2X1_LOC_185/A AND2X1_LOC_126/a_36_24# 0.01fF
C42337 AND2X1_LOC_310/a_8_24# OR2X1_LOC_185/A 0.01fF
C52213 OR2X1_LOC_185/A AND2X1_LOC_86/a_8_24# 0.02fF
C54374 OR2X1_LOC_185/A AND2X1_LOC_529/a_8_24# 0.04fF
C580 AND2X1_LOC_534/a_8_24# OR2X1_LOC_151/A 0.02fF
C19940 OR2X1_LOC_151/A AND2X1_LOC_111/a_8_24# 0.02fF
C34672 OR2X1_LOC_151/A OR2X1_LOC_296/a_8_216# -0.01fF
C35094 OR2X1_LOC_151/A AND2X1_LOC_329/a_8_24# 0.02fF
C11073 OR2X1_LOC_299/a_8_216# OR2X1_LOC_619/Y 0.01fF
C16113 AND2X1_LOC_87/a_8_24# OR2X1_LOC_619/Y 0.03fF
C22185 OR2X1_LOC_299/a_36_216# OR2X1_LOC_619/Y 0.01fF
C32654 AND2X1_LOC_87/a_36_24# OR2X1_LOC_619/Y 0.01fF
C39140 OR2X1_LOC_234/a_8_216# OR2X1_LOC_619/Y 0.03fF
C44667 OR2X1_LOC_119/a_8_216# OR2X1_LOC_619/Y 0.03fF
C50335 OR2X1_LOC_119/a_36_216# OR2X1_LOC_619/Y 0.01fF
C50412 OR2X1_LOC_234/a_36_216# OR2X1_LOC_619/Y 0.01fF
C3469 AND2X1_LOC_264/a_8_24# OR2X1_LOC_52/B 0.03fF
C5569 AND2X1_LOC_685/a_8_24# OR2X1_LOC_52/B 0.03fF
C9952 AND2X1_LOC_687/a_8_24# OR2X1_LOC_52/B 0.01fF
C12260 OR2X1_LOC_681/a_8_216# OR2X1_LOC_52/B 0.03fF
C14522 AND2X1_LOC_264/a_36_24# OR2X1_LOC_52/B 0.01fF
C15701 OR2X1_LOC_413/a_8_216# OR2X1_LOC_52/B 0.03fF
C16536 AND2X1_LOC_276/a_8_24# OR2X1_LOC_52/B 0.13fF
C18712 OR2X1_LOC_422/a_8_216# OR2X1_LOC_52/B 0.03fF
C18756 OR2X1_LOC_694/a_8_216# OR2X1_LOC_52/B 0.02fF
C21319 OR2X1_LOC_413/a_36_216# OR2X1_LOC_52/B 0.02fF
C22254 AND2X1_LOC_685/a_36_24# OR2X1_LOC_52/B 0.01fF
C24633 OR2X1_LOC_421/a_8_216# OR2X1_LOC_52/B 0.03fF
C26477 AND2X1_LOC_687/a_36_24# OR2X1_LOC_52/B 0.01fF
C29276 AND2X1_LOC_155/a_8_24# OR2X1_LOC_52/B 0.06fF
C30223 OR2X1_LOC_275/a_8_216# OR2X1_LOC_52/B 0.02fF
C33065 AND2X1_LOC_276/a_36_24# OR2X1_LOC_52/B 0.01fF
C37340 OR2X1_LOC_682/a_8_216# OR2X1_LOC_52/B -0.01fF
C37725 AND2X1_LOC_274/a_8_24# OR2X1_LOC_52/B 0.03fF
C39530 OR2X1_LOC_681/Y OR2X1_LOC_52/B 0.04fF
C40247 AND2X1_LOC_155/a_36_24# OR2X1_LOC_52/B 0.01fF
C43492 OR2X1_LOC_52/B OR2X1_LOC_153/a_8_216# 0.03fF
C45081 AND2X1_LOC_87/a_8_24# OR2X1_LOC_52/B 0.11fF
C46048 AND2X1_LOC_68/a_8_24# OR2X1_LOC_52/B -0.00fF
C48111 OR2X1_LOC_743/a_8_216# OR2X1_LOC_52/B 0.03fF
C50330 OR2X1_LOC_271/Y OR2X1_LOC_52/B 0.08fF
C54473 AND2X1_LOC_274/a_36_24# OR2X1_LOC_52/B 0.01fF
C258 OR2X1_LOC_45/B OR2X1_LOC_271/a_8_216# 0.01fF
C730 OR2X1_LOC_45/B OR2X1_LOC_681/Y 0.06fF
C4693 OR2X1_LOC_45/B OR2X1_LOC_153/a_8_216# 0.06fF
C5428 OR2X1_LOC_45/B AND2X1_LOC_270/a_8_24# 0.01fF
C6620 OR2X1_LOC_45/B OR2X1_LOC_371/a_8_216# 0.01fF
C8639 OR2X1_LOC_45/B OR2X1_LOC_599/a_8_216# 0.02fF
C10808 OR2X1_LOC_45/B OR2X1_LOC_693/a_8_216# 0.02fF
C11334 OR2X1_LOC_45/B OR2X1_LOC_271/Y 0.01fF
C11822 OR2X1_LOC_45/B OR2X1_LOC_372/a_8_216# 0.01fF
C12073 OR2X1_LOC_45/B OR2X1_LOC_527/a_8_216# 0.01fF
C19148 OR2X1_LOC_45/B OR2X1_LOC_29/a_8_216# 0.01fF
C19460 OR2X1_LOC_45/B OR2X1_LOC_273/a_8_216# 0.01fF
C19710 OR2X1_LOC_45/B OR2X1_LOC_110/a_8_216# 0.01fF
C19925 OR2X1_LOC_45/B OR2X1_LOC_277/a_8_216# 0.01fF
C19948 OR2X1_LOC_45/B OR2X1_LOC_268/a_8_216# 0.01fF
C21891 OR2X1_LOC_45/B OR2X1_LOC_693/a_36_216# 0.02fF
C21955 OR2X1_LOC_45/B OR2X1_LOC_46/a_8_216# 0.02fF
C22949 OR2X1_LOC_45/B AND2X1_LOC_685/a_8_24# 0.01fF
C26628 OR2X1_LOC_45/B AND2X1_LOC_512/a_8_24# 0.03fF
C27198 OR2X1_LOC_45/B AND2X1_LOC_687/a_8_24# 0.01fF
C27411 OR2X1_LOC_45/B OR2X1_LOC_46/a_36_216# 0.02fF
C29334 OR2X1_LOC_45/B OR2X1_LOC_88/a_8_216# 0.01fF
C29476 OR2X1_LOC_45/B OR2X1_LOC_681/a_8_216# 0.03fF
C31476 OR2X1_LOC_45/B OR2X1_LOC_300/a_8_216# 0.01fF
C31705 OR2X1_LOC_45/B OR2X1_LOC_126/a_8_216# 0.18fF
C33238 OR2X1_LOC_45/B OR2X1_LOC_304/a_8_216# 0.01fF
C34674 OR2X1_LOC_45/B OR2X1_LOC_119/a_8_216# 0.01fF
C35853 OR2X1_LOC_45/B OR2X1_LOC_422/a_8_216# 0.01fF
C41792 OR2X1_LOC_45/B OR2X1_LOC_421/a_8_216# 0.02fF
C51814 OR2X1_LOC_45/B AND2X1_LOC_458/a_8_24# 0.01fF
C54735 OR2X1_LOC_45/B OR2X1_LOC_682/a_8_216# 0.02fF
C55424 OR2X1_LOC_45/B AND2X1_LOC_269/a_8_24# 0.01fF
C1629 OR2X1_LOC_89/A OR2X1_LOC_382/a_8_216# 0.01fF
C4539 OR2X1_LOC_89/A OR2X1_LOC_381/a_8_216# 0.01fF
C5530 OR2X1_LOC_699/a_8_216# OR2X1_LOC_89/A 0.01fF
C6021 OR2X1_LOC_89/A AND2X1_LOC_814/a_8_24# 0.01fF
C7131 OR2X1_LOC_89/A OR2X1_LOC_382/a_36_216# -0.00fF
C9524 AND2X1_LOC_66/a_8_24# OR2X1_LOC_89/A 0.09fF
C11355 OR2X1_LOC_89/A OR2X1_LOC_373/a_8_216# 0.01fF
C20958 OR2X1_LOC_696/a_8_216# OR2X1_LOC_89/A 0.01fF
C21021 OR2X1_LOC_89/A AND2X1_LOC_405/a_8_24# 0.12fF
C25457 OR2X1_LOC_89/A AND2X1_LOC_296/a_8_24# 0.01fF
C25955 OR2X1_LOC_89/A AND2X1_LOC_818/a_8_24# 0.01fF
C27632 AND2X1_LOC_502/a_8_24# OR2X1_LOC_89/A 0.01fF
C31451 OR2X1_LOC_89/A OR2X1_LOC_820/B 0.02fF
C34390 OR2X1_LOC_89/A AND2X1_LOC_264/a_8_24# 0.02fF
C35326 OR2X1_LOC_89/A OR2X1_LOC_511/a_8_216# 0.01fF
C35492 OR2X1_LOC_89/A OR2X1_LOC_753/a_8_216# 0.01fF
C35664 OR2X1_LOC_236/a_8_216# OR2X1_LOC_89/A 0.01fF
C39146 OR2X1_LOC_89/A OR2X1_LOC_226/a_8_216# 0.01fF
C39157 OR2X1_LOC_89/A OR2X1_LOC_55/a_8_216# 0.01fF
C1333 OR2X1_LOC_82/a_8_216# OR2X1_LOC_83/A 0.02fF
C27259 AND2X1_LOC_42/a_8_24# OR2X1_LOC_83/A 0.01fF
C49862 OR2X1_LOC_414/a_8_216# OR2X1_LOC_83/A 0.01fF
C18236 OR2X1_LOC_748/A OR2X1_LOC_820/A 0.39fF
C18778 OR2X1_LOC_748/A OR2X1_LOC_820/B 0.40fF
C42338 OR2X1_LOC_820/a_8_216# OR2X1_LOC_748/A 0.01fF
C45987 OR2X1_LOC_748/A OR2X1_LOC_817/a_8_216# 0.01fF
C48050 OR2X1_LOC_748/A OR2X1_LOC_381/a_8_216# 0.39fF
C29579 AND2X1_LOC_377/Y AND2X1_LOC_378/a_36_24# 0.01fF
C32465 VDD AND2X1_LOC_377/Y 0.01fF
C57605 AND2X1_LOC_377/Y VSS 0.07fF
C10019 OR2X1_LOC_673/A AND2X1_LOC_8/a_8_24# 0.19fF
C10648 OR2X1_LOC_673/A AND2X1_LOC_277/a_8_24# 0.01fF
C34533 AND2X1_LOC_672/a_8_24# OR2X1_LOC_673/A 0.01fF
C39162 AND2X1_LOC_102/a_8_24# OR2X1_LOC_673/A 0.01fF
C52366 AND2X1_LOC_90/a_8_24# OR2X1_LOC_673/A 0.01fF
C35309 OR2X1_LOC_164/Y OR2X1_LOC_164/a_8_216# 0.14fF
C43576 OR2X1_LOC_527/a_8_216# OR2X1_LOC_164/Y 0.01fF
C21498 OR2X1_LOC_322/a_8_216# OR2X1_LOC_322/Y 0.01fF
C29547 AND2X1_LOC_374/a_8_24# OR2X1_LOC_322/Y 0.23fF
C32400 OR2X1_LOC_322/a_36_216# OR2X1_LOC_322/Y 0.01fF
C50028 OR2X1_LOC_322/Y OR2X1_LOC_323/a_8_216# 0.04fF
C5429 OR2X1_LOC_376/Y OR2X1_LOC_377/a_8_216# 0.01fF
C10343 OR2X1_LOC_64/a_8_216# OR2X1_LOC_588/Y 0.01fF
C1184 OR2X1_LOC_820/a_8_216# OR2X1_LOC_820/B 0.05fF
C3742 OR2X1_LOC_820/B OR2X1_LOC_382/a_8_216# 0.01fF
C6633 OR2X1_LOC_820/B OR2X1_LOC_381/a_8_216# 0.01fF
C7678 OR2X1_LOC_699/a_8_216# OR2X1_LOC_820/B 0.01fF
C8099 AND2X1_LOC_847/Y OR2X1_LOC_820/B 0.01fF
C14801 VDD OR2X1_LOC_820/B 0.11fF
C33031 OR2X1_LOC_820/A OR2X1_LOC_820/B 0.19fF
C36914 AND2X1_LOC_847/a_8_24# OR2X1_LOC_820/B 0.05fF
C42110 OR2X1_LOC_77/a_8_216# OR2X1_LOC_820/B 0.01fF
C48515 OR2X1_LOC_604/A OR2X1_LOC_820/B 0.01fF
C56700 OR2X1_LOC_820/B VSS -0.11fF
C54558 OR2X1_LOC_696/a_8_216# OR2X1_LOC_696/Y -0.00fF
C1327 OR2X1_LOC_306/Y AND2X1_LOC_512/a_8_24# 0.03fF
C23469 OR2X1_LOC_306/Y AND2X1_LOC_512/a_36_24# 0.01fF
C5602 VDD OR2X1_LOC_269/A -0.00fF
C12982 AND2X1_LOC_56/B OR2X1_LOC_269/A 0.01fF
C16411 OR2X1_LOC_276/B OR2X1_LOC_269/A 0.02fF
C56457 OR2X1_LOC_269/A VSS 0.38fF
C31058 OR2X1_LOC_276/B OR2X1_LOC_630/B 0.01fF
C8145 AND2X1_LOC_93/a_8_24# OR2X1_LOC_98/B 0.01fF
C2895 OR2X1_LOC_378/Y OR2X1_LOC_375/a_8_216# 0.39fF
C49605 OR2X1_LOC_378/Y OR2X1_LOC_378/a_8_216# 0.01fF
C6947 OR2X1_LOC_506/A AND2X1_LOC_419/a_8_24# 0.01fF
C50103 OR2X1_LOC_506/A AND2X1_LOC_433/a_8_24# 0.18fF
C15568 AND2X1_LOC_372/a_8_24# OR2X1_LOC_541/A 0.01fF
C29644 OR2X1_LOC_541/A AND2X1_LOC_272/a_8_24# 0.01fF
C48849 OR2X1_LOC_541/A OR2X1_LOC_274/a_8_216# 0.07fF
C13657 OR2X1_LOC_686/A AND2X1_LOC_684/a_8_24# 0.01fF
C19366 VDD OR2X1_LOC_686/A 0.21fF
C28294 AND2X1_LOC_582/a_8_24# OR2X1_LOC_686/A 0.08fF
C28331 OR2X1_LOC_686/A AND2X1_LOC_682/a_8_24# 0.27fF
C57651 OR2X1_LOC_686/A VSS -0.19fF
C34525 OR2X1_LOC_801/a_8_216# OR2X1_LOC_138/A 0.01fF
C55486 OR2X1_LOC_138/A OR2X1_LOC_514/a_8_216# 0.47fF
C45471 OR2X1_LOC_294/a_8_216# OR2X1_LOC_296/Y 0.01fF
C25575 AND2X1_LOC_43/a_8_24# OR2X1_LOC_195/A 0.09fF
C6948 OR2X1_LOC_71/a_8_216# OR2X1_LOC_71/A 0.01fF
C7821 OR2X1_LOC_291/a_36_216# OR2X1_LOC_71/A 0.01fF
C8341 OR2X1_LOC_278/a_8_216# OR2X1_LOC_71/A 0.03fF
C10330 AND2X1_LOC_86/a_8_24# OR2X1_LOC_71/A 0.01fF
C10818 AND2X1_LOC_55/a_8_24# OR2X1_LOC_71/A 0.02fF
C11290 OR2X1_LOC_611/a_8_216# OR2X1_LOC_71/A 0.02fF
C12472 AND2X1_LOC_529/a_8_24# OR2X1_LOC_71/A 0.01fF
C23134 AND2X1_LOC_73/a_8_24# OR2X1_LOC_71/A 0.04fF
C24007 AND2X1_LOC_414/a_8_24# OR2X1_LOC_71/A 0.02fF
C27013 OR2X1_LOC_62/a_8_216# OR2X1_LOC_71/A 0.01fF
C31269 OR2X1_LOC_92/a_8_216# OR2X1_LOC_71/A 0.01fF
C34073 AND2X1_LOC_143/a_8_24# OR2X1_LOC_71/A 0.05fF
C35307 AND2X1_LOC_126/a_8_24# OR2X1_LOC_71/A 0.01fF
C39260 AND2X1_LOC_133/a_8_24# OR2X1_LOC_71/A 0.01fF
C39787 OR2X1_LOC_71/A OR2X1_LOC_398/a_8_216# 0.01fF
C44156 OR2X1_LOC_71/A OR2X1_LOC_150/a_8_216# 0.18fF
C52957 OR2X1_LOC_291/a_8_216# OR2X1_LOC_71/A 0.01fF
C3534 OR2X1_LOC_96/B OR2X1_LOC_54/a_8_216# 0.01fF
C25840 OR2X1_LOC_820/A OR2X1_LOC_96/B 0.03fF
C30037 OR2X1_LOC_159/a_8_216# OR2X1_LOC_96/B 0.01fF
C21012 OR2X1_LOC_820/A AND2X1_LOC_750/a_8_24# -0.02fF
C21359 OR2X1_LOC_820/A OR2X1_LOC_751/A 0.82fF
C36217 OR2X1_LOC_820/A OR2X1_LOC_748/a_8_216# 0.04fF
C43058 OR2X1_LOC_820/A AND2X1_LOC_750/a_36_24# 0.01fF
C47980 OR2X1_LOC_604/A OR2X1_LOC_820/A 0.02fF
C57255 OR2X1_LOC_820/A VSS 0.29fF
C2637 AND2X1_LOC_73/a_8_24# OR2X1_LOC_532/B 0.03fF
C4339 AND2X1_LOC_329/a_8_24# OR2X1_LOC_532/B 0.01fF
C7652 AND2X1_LOC_371/a_8_24# OR2X1_LOC_532/B 0.01fF
C11977 OR2X1_LOC_405/a_8_216# OR2X1_LOC_532/B 0.01fF
C15664 OR2X1_LOC_532/B OR2X1_LOC_548/a_8_216# 0.01fF
C19545 AND2X1_LOC_530/a_8_24# OR2X1_LOC_532/B 0.01fF
C20166 OR2X1_LOC_606/a_8_216# OR2X1_LOC_532/B 0.07fF
C20916 AND2X1_LOC_372/a_8_24# OR2X1_LOC_532/B 0.01fF
C25178 AND2X1_LOC_80/a_8_24# OR2X1_LOC_532/B 0.17fF
C25248 AND2X1_LOC_15/a_8_24# OR2X1_LOC_532/B 0.01fF
C25471 AND2X1_LOC_90/a_8_24# OR2X1_LOC_532/B 0.01fF
C28015 OR2X1_LOC_691/a_8_216# OR2X1_LOC_532/B 0.01fF
C34845 OR2X1_LOC_458/a_8_216# OR2X1_LOC_532/B 0.01fF
C34901 OR2X1_LOC_532/B AND2X1_LOC_272/a_8_24# 0.01fF
C36135 AND2X1_LOC_49/a_8_24# OR2X1_LOC_532/B 0.10fF
C36458 AND2X1_LOC_387/a_8_24# OR2X1_LOC_532/B 0.01fF
C38747 AND2X1_LOC_23/a_8_24# OR2X1_LOC_532/B 0.01fF
C39827 OR2X1_LOC_532/B AND2X1_LOC_277/a_8_24# 0.01fF
C43472 OR2X1_LOC_532/B OR2X1_LOC_750/a_8_216# 0.01fF
C44389 OR2X1_LOC_532/B AND2X1_LOC_6/a_8_24# 0.01fF
C45186 AND2X1_LOC_111/a_8_24# OR2X1_LOC_532/B 0.01fF
C45510 AND2X1_LOC_110/a_8_24# OR2X1_LOC_532/B 0.01fF
C685 OR2X1_LOC_294/a_8_216# OR2X1_LOC_78/A 0.01fF
C686 AND2X1_LOC_304/a_8_24# OR2X1_LOC_78/A 0.01fF
C1570 AND2X1_LOC_48/a_8_24# OR2X1_LOC_78/A 0.01fF
C3335 AND2X1_LOC_104/a_8_24# OR2X1_LOC_78/A 0.03fF
C4599 AND2X1_LOC_329/a_36_24# OR2X1_LOC_78/A 0.01fF
C6210 OR2X1_LOC_327/a_8_216# OR2X1_LOC_78/A 0.02fF
C11658 OR2X1_LOC_78/A OR2X1_LOC_502/a_8_216# 0.03fF
C12130 AND2X1_LOC_93/a_8_24# OR2X1_LOC_78/A 0.07fF
C14384 AND2X1_LOC_104/a_36_24# OR2X1_LOC_78/A 0.01fF
C19943 AND2X1_LOC_49/a_8_24# OR2X1_LOC_78/A 0.01fF
C22792 OR2X1_LOC_78/A OR2X1_LOC_502/a_36_216# 0.03fF
C23022 AND2X1_LOC_77/a_8_24# OR2X1_LOC_78/A -0.01fF
C25439 AND2X1_LOC_696/a_8_24# OR2X1_LOC_78/A 0.01fF
C28112 AND2X1_LOC_6/a_8_24# OR2X1_LOC_78/A 0.04fF
C28653 AND2X1_LOC_511/a_8_24# OR2X1_LOC_78/A 0.01fF
C35049 AND2X1_LOC_306/a_8_24# OR2X1_LOC_78/A 0.01fF
C38126 AND2X1_LOC_119/a_8_24# OR2X1_LOC_78/A 0.17fF
C38946 OR2X1_LOC_264/a_8_216# OR2X1_LOC_78/A 0.01fF
C39088 AND2X1_LOC_6/a_36_24# OR2X1_LOC_78/A 0.01fF
C42808 AND2X1_LOC_82/a_8_24# OR2X1_LOC_78/A 0.01fF
C43721 OR2X1_LOC_296/a_8_216# OR2X1_LOC_78/A 0.01fF
C44129 AND2X1_LOC_329/a_8_24# OR2X1_LOC_78/A 0.04fF
C116 AND2X1_LOC_56/B AND2X1_LOC_699/a_8_24# 0.01fF
C435 AND2X1_LOC_56/B OR2X1_LOC_82/a_8_216# 0.06fF
C1891 AND2X1_LOC_56/B AND2X1_LOC_268/a_8_24# 0.01fF
C11812 AND2X1_LOC_56/B OR2X1_LOC_596/a_8_216# 0.01fF
C13276 AND2X1_LOC_56/B OR2X1_LOC_296/a_8_216# 0.07fF
C13677 AND2X1_LOC_56/B AND2X1_LOC_329/a_8_24# 0.04fF
C14188 AND2X1_LOC_56/B OR2X1_LOC_276/B 0.16fF
C15572 AND2X1_LOC_56/B AND2X1_LOC_256/a_8_24# 0.01fF
C16008 AND2X1_LOC_56/B OR2X1_LOC_514/a_8_216# 0.02fF
C16490 AND2X1_LOC_56/B AND2X1_LOC_628/a_8_24# 0.01fF
C20277 OR2X1_LOC_121/a_8_216# AND2X1_LOC_56/B 0.01fF
C21228 AND2X1_LOC_56/B OR2X1_LOC_410/a_8_216# 0.02fF
C21378 AND2X1_LOC_56/B AND2X1_LOC_136/a_8_24# 0.02fF
C22965 AND2X1_LOC_73/a_36_24# AND2X1_LOC_56/B 0.01fF
C28734 AND2X1_LOC_530/a_8_24# AND2X1_LOC_56/B 0.17fF
C29711 AND2X1_LOC_56/B OR2X1_LOC_407/a_8_216# 0.02fF
C31801 AND2X1_LOC_56/B AND2X1_LOC_233/a_8_24# 0.02fF
C35819 AND2X1_LOC_56/B OR2X1_LOC_515/a_8_216# 0.01fF
C39131 AND2X1_LOC_56/B AND2X1_LOC_56/a_8_24# 0.11fF
C39967 AND2X1_LOC_56/B AND2X1_LOC_271/a_8_24# 0.01fF
C46824 AND2X1_LOC_94/a_8_24# AND2X1_LOC_56/B 0.13fF
C47633 AND2X1_LOC_56/B AND2X1_LOC_411/a_8_24# 0.02fF
C52357 AND2X1_LOC_56/B OR2X1_LOC_269/a_8_216# 0.01fF
C52782 AND2X1_LOC_56/B AND2X1_LOC_699/a_36_24# -0.00fF
C53194 AND2X1_LOC_527/a_8_24# AND2X1_LOC_56/B 0.01fF
C55600 AND2X1_LOC_56/B OR2X1_LOC_185/a_8_216# 0.07fF
C264 AND2X1_LOC_91/B AND2X1_LOC_85/a_8_24# 0.01fF
C538 AND2X1_LOC_91/B AND2X1_LOC_263/a_8_24# 0.01fF
C2369 AND2X1_LOC_91/B OR2X1_LOC_814/a_8_216# 0.02fF
C13588 AND2X1_LOC_91/B OR2X1_LOC_276/B 0.10fF
C16305 AND2X1_LOC_91/B AND2X1_LOC_371/a_8_24# 0.15fF
C22758 AND2X1_LOC_91/B AND2X1_LOC_488/a_8_24# 0.02fF
C28263 AND2X1_LOC_91/B AND2X1_LOC_104/a_8_24# 0.01fF
C28451 AND2X1_LOC_91/B AND2X1_LOC_225/a_8_24# 0.05fF
C36621 AND2X1_LOC_91/B AND2X1_LOC_164/a_8_24# 0.03fF
C43530 AND2X1_LOC_91/B AND2X1_LOC_421/a_8_24# 0.03fF
C49710 AND2X1_LOC_91/B AND2X1_LOC_38/a_8_24# 0.01fF
C11534 AND2X1_LOC_847/a_8_24# AND2X1_LOC_847/Y 0.02fF
C35207 OR2X1_LOC_817/a_8_216# AND2X1_LOC_847/Y 0.06fF
C46421 OR2X1_LOC_817/a_36_216# AND2X1_LOC_847/Y 0.01fF
C48053 OR2X1_LOC_450/B AND2X1_LOC_426/a_8_24# 0.01fF
C50709 OR2X1_LOC_450/B AND2X1_LOC_694/a_8_24# 0.20fF
C4034 AND2X1_LOC_300/a_8_24# OR2X1_LOC_831/A 0.02fF
C9120 OR2X1_LOC_831/A AND2X1_LOC_273/a_36_24# 0.01fF
C43040 OR2X1_LOC_831/A AND2X1_LOC_273/a_8_24# 0.12fF
C843 OR2X1_LOC_121/Y OR2X1_LOC_276/a_36_216# 0.01fF
C3628 OR2X1_LOC_121/Y AND2X1_LOC_625/a_8_24# 0.04fF
C10259 OR2X1_LOC_121/Y OR2X1_LOC_66/a_8_216# 0.02fF
C15724 OR2X1_LOC_121/Y OR2X1_LOC_66/a_36_216# 0.01fF
C45918 OR2X1_LOC_121/Y OR2X1_LOC_276/B 0.02fF
C51516 OR2X1_LOC_121/Y OR2X1_LOC_276/a_8_216# 0.05fF
C53151 OR2X1_LOC_417/Y AND2X1_LOC_515/a_8_24# 0.23fF
C53767 OR2X1_LOC_417/Y OR2X1_LOC_417/a_8_216# 0.01fF
C11734 OR2X1_LOC_289/a_8_216# OR2X1_LOC_289/Y -0.00fF
C34552 OR2X1_LOC_369/a_8_216# OR2X1_LOC_309/Y 0.01fF
C47508 OR2X1_LOC_309/a_8_216# OR2X1_LOC_309/Y 0.01fF
C26514 AND2X1_LOC_599/a_8_24# OR2X1_LOC_598/Y 0.08fF
C37482 AND2X1_LOC_599/a_36_24# OR2X1_LOC_598/Y 0.01fF
C18121 AND2X1_LOC_611/a_8_24# OR2X1_LOC_415/Y 0.13fF
C29146 AND2X1_LOC_611/a_36_24# OR2X1_LOC_415/Y 0.01fF
C47868 OR2X1_LOC_415/Y OR2X1_LOC_548/a_8_216# 0.01fF
C51665 AND2X1_LOC_530/a_8_24# OR2X1_LOC_415/Y 0.01fF
C15793 OR2X1_LOC_688/Y AND2X1_LOC_689/a_8_24# 0.23fF
C35569 VDD OR2X1_LOC_688/Y 0.16fF
C57521 OR2X1_LOC_688/Y VSS 0.07fF
C41827 AND2X1_LOC_585/a_8_24# OR2X1_LOC_637/B 0.01fF
C12873 OR2X1_LOC_287/B AND2X1_LOC_77/a_8_24# -0.00fF
C17128 OR2X1_LOC_287/B AND2X1_LOC_283/a_8_24# 0.01fF
C23431 OR2X1_LOC_287/B OR2X1_LOC_814/a_8_216# 0.01fF
C32701 OR2X1_LOC_287/B AND2X1_LOC_82/a_8_24# 0.01fF
C43643 OR2X1_LOC_287/B AND2X1_LOC_488/a_8_24# 0.01fF
C3021 OR2X1_LOC_760/a_8_216# OR2X1_LOC_16/A 0.01fF
C8306 OR2X1_LOC_329/a_8_216# OR2X1_LOC_16/A 0.01fF
C12289 AND2X1_LOC_686/a_8_24# OR2X1_LOC_16/A 0.01fF
C13171 OR2X1_LOC_611/a_8_216# OR2X1_LOC_16/A 0.07fF
C13610 OR2X1_LOC_80/a_8_216# OR2X1_LOC_16/A 0.07fF
C16375 AND2X1_LOC_274/a_8_24# OR2X1_LOC_16/A 0.17fF
C18601 OR2X1_LOC_299/a_8_216# OR2X1_LOC_16/A 0.06fF
C19339 OR2X1_LOC_684/a_8_216# OR2X1_LOC_16/A 0.02fF
C21272 OR2X1_LOC_411/a_8_216# OR2X1_LOC_16/A 0.06fF
C21670 OR2X1_LOC_293/a_8_216# OR2X1_LOC_16/A 0.43fF
C25996 OR2X1_LOC_16/A OR2X1_LOC_599/a_8_216# 0.01fF
C32951 AND2X1_LOC_598/a_8_24# OR2X1_LOC_16/A 0.01fF
C36469 OR2X1_LOC_16/A OR2X1_LOC_29/a_8_216# 0.06fF
C40077 AND2X1_LOC_398/a_8_24# OR2X1_LOC_16/A 0.09fF
C48137 AND2X1_LOC_800/a_8_24# OR2X1_LOC_16/A 0.01fF
C48801 OR2X1_LOC_683/a_8_216# OR2X1_LOC_16/A 0.05fF
C49071 OR2X1_LOC_16/A OR2X1_LOC_300/a_8_216# 0.11fF
C53618 AND2X1_LOC_801/B OR2X1_LOC_16/A 0.03fF
C54705 OR2X1_LOC_291/a_8_216# OR2X1_LOC_16/A 0.11fF
C615 AND2X1_LOC_294/a_8_24# OR2X1_LOC_13/B 0.02fF
C7948 AND2X1_LOC_66/a_8_24# OR2X1_LOC_13/B 0.04fF
C8365 AND2X1_LOC_120/a_8_24# OR2X1_LOC_13/B 0.01fF
C10594 OR2X1_LOC_761/a_8_216# OR2X1_LOC_13/B 0.05fF
C12509 AND2X1_LOC_801/a_8_24# OR2X1_LOC_13/B 0.04fF
C14168 OR2X1_LOC_102/a_8_216# OR2X1_LOC_13/B 0.01fF
C24635 OR2X1_LOC_13/B OR2X1_LOC_534/a_8_216# 0.03fF
C28222 OR2X1_LOC_306/a_8_216# OR2X1_LOC_13/B 0.01fF
C31541 AND2X1_LOC_121/a_8_24# OR2X1_LOC_13/B 0.04fF
C32808 AND2X1_LOC_513/a_8_24# OR2X1_LOC_13/B 0.01fF
C32865 AND2X1_LOC_264/a_8_24# OR2X1_LOC_13/B 0.06fF
C34133 OR2X1_LOC_86/a_8_216# OR2X1_LOC_13/B 0.02fF
C38805 AND2X1_LOC_512/a_8_24# OR2X1_LOC_13/B 0.01fF
C42609 AND2X1_LOC_121/a_36_24# OR2X1_LOC_13/B 0.01fF
C44527 OR2X1_LOC_85/a_8_216# OR2X1_LOC_13/B 0.19fF
C45336 OR2X1_LOC_255/a_8_216# OR2X1_LOC_13/B 0.01fF
C48457 AND2X1_LOC_801/B OR2X1_LOC_13/B 0.02fF
C1194 OR2X1_LOC_133/a_8_216# OR2X1_LOC_74/A 0.40fF
C2454 OR2X1_LOC_111/a_8_216# OR2X1_LOC_74/A 0.05fF
C3881 OR2X1_LOC_74/A AND2X1_LOC_274/a_36_24# 0.01fF
C7949 OR2X1_LOC_110/a_8_216# OR2X1_LOC_74/A 0.06fF
C9019 OR2X1_LOC_74/A AND2X1_LOC_264/a_8_24# 0.02fF
C16784 OR2X1_LOC_74/A OR2X1_LOC_150/a_8_216# 0.14fF
C17315 OR2X1_LOC_74/A OR2X1_LOC_323/a_8_216# 0.03fF
C17583 OR2X1_LOC_74/A OR2X1_LOC_88/a_8_216# 0.05fF
C20423 AND2X1_LOC_185/a_8_24# OR2X1_LOC_74/A 0.08fF
C23514 OR2X1_LOC_73/a_8_216# OR2X1_LOC_74/A 0.02fF
C25515 OR2X1_LOC_291/a_8_216# OR2X1_LOC_74/A 0.01fF
C35720 OR2X1_LOC_275/a_8_216# OR2X1_LOC_74/A 0.07fF
C36930 OR2X1_LOC_278/a_8_216# OR2X1_LOC_74/A 0.01fF
C43340 OR2X1_LOC_74/A AND2X1_LOC_274/a_8_24# 0.05fF
C49169 OR2X1_LOC_74/A OR2X1_LOC_153/a_8_216# 0.05fF
C11176 OR2X1_LOC_246/Y OR2X1_LOC_10/a_8_216# 0.06fF
C33094 OR2X1_LOC_246/Y OR2X1_LOC_246/a_8_216# 0.01fF
C45668 OR2X1_LOC_246/Y OR2X1_LOC_150/a_8_216# 0.03fF
C389 OR2X1_LOC_235/B OR2X1_LOC_278/a_8_216# 0.01fF
C3004 OR2X1_LOC_235/B OR2X1_LOC_233/a_36_216# 0.01fF
C4200 OR2X1_LOC_235/B AND2X1_LOC_85/a_8_24# 0.01fF
C4424 OR2X1_LOC_235/B AND2X1_LOC_263/a_8_24# 0.02fF
C11926 OR2X1_LOC_235/B OR2X1_LOC_293/a_8_216# 0.05fF
C15914 OR2X1_LOC_235/B OR2X1_LOC_15/a_8_216# 0.01fF
C19168 OR2X1_LOC_235/B OR2X1_LOC_62/a_8_216# 0.02fF
C20491 OR2X1_LOC_235/B AND2X1_LOC_672/a_8_24# 0.01fF
C25042 OR2X1_LOC_235/B AND2X1_LOC_102/a_8_24# 0.01fF
C28338 OR2X1_LOC_235/B AND2X1_LOC_71/a_8_24# 0.11fF
C29941 OR2X1_LOC_235/B AND2X1_LOC_150/a_8_24# 0.11fF
C32130 OR2X1_LOC_235/B AND2X1_LOC_104/a_8_24# 0.01fF
C36923 OR2X1_LOC_235/B OR2X1_LOC_234/a_8_216# 0.02fF
C37926 AND2X1_LOC_90/a_8_24# OR2X1_LOC_235/B 0.02fF
C38038 OR2X1_LOC_235/B OR2X1_LOC_38/a_8_216# -0.02fF
C43686 OR2X1_LOC_235/B OR2X1_LOC_38/a_36_216# 0.01fF
C43773 OR2X1_LOC_235/B AND2X1_LOC_671/a_8_24# -0.01fF
C44937 OR2X1_LOC_235/B OR2X1_LOC_291/a_8_216# 0.01fF
C52022 OR2X1_LOC_235/B AND2X1_LOC_8/a_8_24# 0.01fF
C52583 OR2X1_LOC_235/B AND2X1_LOC_277/a_8_24# 0.01fF
C53626 OR2X1_LOC_235/B OR2X1_LOC_233/a_8_216# 0.02fF
C53633 OR2X1_LOC_235/B AND2X1_LOC_38/a_8_24# 0.03fF
C55674 OR2X1_LOC_235/B AND2X1_LOC_63/a_8_24# 0.11fF
C827 OR2X1_LOC_604/A OR2X1_LOC_77/a_8_216# 0.02fF
C2044 OR2X1_LOC_604/A OR2X1_LOC_236/a_36_216# 0.01fF
C5501 OR2X1_LOC_604/A OR2X1_LOC_55/a_36_216# 0.01fF
C5739 OR2X1_LOC_604/A OR2X1_LOC_683/a_8_216# 0.01fF
C6298 OR2X1_LOC_604/A OR2X1_LOC_77/a_36_216# 0.01fF
C8779 OR2X1_LOC_604/A OR2X1_LOC_90/a_8_216# 0.06fF
C9754 OR2X1_LOC_604/A OR2X1_LOC_73/a_8_216# 0.02fF
C14289 OR2X1_LOC_604/A OR2X1_LOC_90/a_36_216# 0.01fF
C15220 OR2X1_LOC_604/A OR2X1_LOC_73/a_36_216# 0.01fF
C18504 OR2X1_LOC_604/A OR2X1_LOC_382/a_8_216# 0.04fF
C21136 OR2X1_LOC_604/A AND2X1_LOC_155/a_8_24# 0.01fF
C21511 OR2X1_LOC_604/A OR2X1_LOC_381/a_8_216# 0.03fF
C22495 OR2X1_LOC_604/A OR2X1_LOC_699/a_8_216# 0.06fF
C24061 OR2X1_LOC_604/A OR2X1_LOC_382/a_36_216# -0.00fF
C25480 OR2X1_LOC_604/A AND2X1_LOC_686/a_8_24# 0.01fF
C26957 OR2X1_LOC_604/A OR2X1_LOC_381/a_36_216# 0.01fF
C27934 OR2X1_LOC_604/A OR2X1_LOC_699/a_36_216# 0.01fF
C32437 OR2X1_LOC_604/A OR2X1_LOC_684/a_8_216# 0.01fF
C32613 OR2X1_LOC_604/A OR2X1_LOC_430/a_8_216# 0.02fF
C36170 OR2X1_LOC_604/A AND2X1_LOC_750/a_8_24# 0.09fF
C38337 OR2X1_LOC_604/A OR2X1_LOC_672/a_8_216# 0.06fF
C39675 OR2X1_LOC_604/A OR2X1_LOC_743/a_8_216# 0.01fF
C42248 OR2X1_LOC_604/A AND2X1_LOC_296/a_8_24# 0.04fF
C42801 OR2X1_LOC_604/A AND2X1_LOC_818/a_8_24# 0.03fF
C43512 OR2X1_LOC_133/a_8_216# OR2X1_LOC_604/A 0.06fF
C43716 OR2X1_LOC_604/A OR2X1_LOC_430/a_36_216# 0.02fF
C43968 OR2X1_LOC_604/A OR2X1_LOC_672/a_36_216# 0.01fF
C46413 OR2X1_LOC_604/A OR2X1_LOC_426/a_8_216# 0.01fF
C46449 OR2X1_LOC_604/A OR2X1_LOC_419/a_8_216# 0.04fF
C52680 OR2X1_LOC_604/A OR2X1_LOC_236/a_8_216# 0.03fF
C54665 OR2X1_LOC_133/a_36_216# OR2X1_LOC_604/A 0.01fF
C56227 OR2X1_LOC_604/A OR2X1_LOC_55/a_8_216# 0.06fF
C8254 OR2X1_LOC_511/Y OR2X1_LOC_511/a_8_216# -0.00fF
C12828 OR2X1_LOC_48/Y OR2X1_LOC_48/a_8_216# 0.01fF
C26375 OR2X1_LOC_599/A OR2X1_LOC_696/a_8_216# 0.03fF
C40828 OR2X1_LOC_599/A OR2X1_LOC_511/a_8_216# 0.02fF
C20604 OR2X1_LOC_693/a_8_216# OR2X1_LOC_692/Y 0.02fF
C14864 OR2X1_LOC_409/B OR2X1_LOC_585/a_8_216# 0.01fF
C19402 OR2X1_LOC_409/B OR2X1_LOC_377/a_8_216# 0.02fF
C20625 OR2X1_LOC_409/B OR2X1_LOC_409/a_8_216# 0.07fF
C35282 OR2X1_LOC_409/B OR2X1_LOC_752/a_8_216# 0.01fF
C40351 AND2X1_LOC_375/a_8_24# OR2X1_LOC_409/B 0.01fF
C40562 OR2X1_LOC_409/B OR2X1_LOC_376/a_8_216# 0.01fF
C42966 OR2X1_LOC_409/B OR2X1_LOC_59/a_8_216# 0.01fF
C27645 OR2X1_LOC_273/Y AND2X1_LOC_274/a_8_24# 0.05fF
C48273 OR2X1_LOC_273/a_8_216# OR2X1_LOC_273/Y 0.02fF
C21846 OR2X1_LOC_681/Y AND2X1_LOC_685/a_8_24# 0.23fF
C54007 VDD OR2X1_LOC_681/Y 0.12fF
C57062 OR2X1_LOC_681/Y VSS 0.06fF
C11219 OR2X1_LOC_323/a_8_216# OR2X1_LOC_323/Y 0.02fF
C16968 OR2X1_LOC_527/a_8_216# OR2X1_LOC_527/Y 0.03fF
C14183 AND2X1_LOC_729/B OR2X1_LOC_43/a_8_216# 0.01fF
C16763 AND2X1_LOC_729/B OR2X1_LOC_761/a_8_216# 0.02fF
C34378 OR2X1_LOC_306/a_8_216# AND2X1_LOC_729/B 0.01fF
C45143 AND2X1_LOC_512/a_8_24# AND2X1_LOC_729/B 0.01fF
C45540 OR2X1_LOC_306/a_36_216# AND2X1_LOC_729/B 0.01fF
C33022 OR2X1_LOC_100/a_8_216# OR2X1_LOC_100/Y 0.01fF
C16625 OR2X1_LOC_271/Y AND2X1_LOC_276/Y 0.02fF
C39029 AND2X1_LOC_276/Y AND2X1_LOC_276/a_8_24# 0.01fF
C39922 AND2X1_LOC_801/B AND2X1_LOC_809/A 0.01fF
C14523 AND2X1_LOC_412/a_8_24# OR2X1_LOC_240/A 0.05fF
C36513 AND2X1_LOC_412/a_36_24# OR2X1_LOC_240/A 0.01fF
C38207 AND2X1_LOC_42/a_8_24# OR2X1_LOC_240/A 0.06fF
C45928 OR2X1_LOC_836/A AND2X1_LOC_824/a_8_24# 0.02fF
C9703 OR2X1_LOC_751/A AND2X1_LOC_750/a_8_24# 0.10fF
C16143 OR2X1_LOC_515/a_8_216# OR2X1_LOC_515/Y 0.01fF
C3188 AND2X1_LOC_687/A AND2X1_LOC_687/a_8_24# 0.10fF
C5443 OR2X1_LOC_681/a_8_216# AND2X1_LOC_687/A 0.03fF
C30638 OR2X1_LOC_682/a_8_216# AND2X1_LOC_687/A 0.47fF
C30981 VDD AND2X1_LOC_687/A -0.00fF
C47405 OR2X1_LOC_682/Y AND2X1_LOC_687/A 0.01fF
C55004 AND2X1_LOC_685/a_8_24# AND2X1_LOC_687/A 0.01fF
C57061 AND2X1_LOC_687/A VSS 0.38fF
C10967 OR2X1_LOC_687/B OR2X1_LOC_687/A 0.15fF
C30792 OR2X1_LOC_686/a_8_216# OR2X1_LOC_687/A -0.00fF
C44943 OR2X1_LOC_685/A OR2X1_LOC_687/A 0.15fF
C47088 VDD OR2X1_LOC_687/A -0.00fF
C56095 OR2X1_LOC_685/a_8_216# OR2X1_LOC_687/A 0.40fF
C57649 OR2X1_LOC_687/A VSS 0.22fF
C12723 VDD OR2X1_LOC_820/Y 0.06fF
C34902 OR2X1_LOC_820/Y AND2X1_LOC_847/a_8_24# 0.01fF
C56931 OR2X1_LOC_820/Y VSS 0.10fF
C1305 OR2X1_LOC_275/A OR2X1_LOC_517/A 0.24fF
C10984 OR2X1_LOC_517/A OR2X1_LOC_67/A 0.02fF
C17848 OR2X1_LOC_275/a_8_216# OR2X1_LOC_517/A 0.48fF
C23879 OR2X1_LOC_517/A OR2X1_LOC_245/a_8_216# 0.03fF
C25350 VDD OR2X1_LOC_517/A 0.15fF
C33860 OR2X1_LOC_625/a_8_216# OR2X1_LOC_517/A 0.01fF
C57201 OR2X1_LOC_517/A VSS 0.72fF
C12188 OR2X1_LOC_121/a_8_216# OR2X1_LOC_185/Y 0.03fF
C14719 OR2X1_LOC_185/Y AND2X1_LOC_760/a_8_24# 0.24fF
C14735 OR2X1_LOC_185/Y OR2X1_LOC_121/A 0.13fF
C15657 OR2X1_LOC_185/Y OR2X1_LOC_274/Y 0.02fF
C26777 OR2X1_LOC_185/Y OR2X1_LOC_800/A 0.01fF
C37450 OR2X1_LOC_185/Y OR2X1_LOC_66/Y 0.03fF
C40239 OR2X1_LOC_185/Y OR2X1_LOC_405/A 0.25fF
C43231 OR2X1_LOC_185/Y OR2X1_LOC_801/a_8_216# 0.01fF
C43338 OR2X1_LOC_185/Y OR2X1_LOC_800/a_8_216# 0.01fF
C48820 OR2X1_LOC_185/Y OR2X1_LOC_120/a_8_216# 0.03fF
C51419 OR2X1_LOC_185/Y VDD 2.10fF
C55272 OR2X1_LOC_185/Y OR2X1_LOC_274/a_8_216# 0.04fF
C58055 OR2X1_LOC_185/Y VSS -4.38fF
C2321 OR2X1_LOC_691/B OR2X1_LOC_691/a_8_216# 0.07fF
C57977 OR2X1_LOC_691/B VSS 0.20fF
C25275 AND2X1_LOC_800/a_8_24# OR2X1_LOC_760/Y 0.06fF
C56946 OR2X1_LOC_760/Y VSS -0.07fF
C21882 OR2X1_LOC_375/a_8_216# OR2X1_LOC_375/Y 0.02fF
C28357 AND2X1_LOC_376/a_8_24# OR2X1_LOC_375/Y 0.03fF
C28671 AND2X1_LOC_752/a_8_24# OR2X1_LOC_375/Y 0.23fF
C45246 VDD OR2X1_LOC_375/Y 0.33fF
C56388 OR2X1_LOC_375/Y VSS 0.07fF
C28874 AND2X1_LOC_599/a_8_24# OR2X1_LOC_644/A 0.01fF
C26959 OR2X1_LOC_548/A VDD -0.00fF
C48746 OR2X1_LOC_548/A OR2X1_LOC_548/a_8_216# 0.47fF
C57999 OR2X1_LOC_548/A VSS 0.15fF
C2387 OR2X1_LOC_270/Y AND2X1_LOC_271/a_8_24# 0.05fF
C21786 VDD OR2X1_LOC_270/Y 0.24fF
C56891 OR2X1_LOC_270/Y VSS -0.04fF
C45 OR2X1_LOC_411/Y AND2X1_LOC_461/a_8_24# 0.01fF
C14781 OR2X1_LOC_411/Y OR2X1_LOC_413/a_8_216# 0.40fF
C57310 OR2X1_LOC_411/Y VSS 0.22fF
C57471 OR2X1_LOC_88/A VSS 0.02fF
C9063 OR2X1_LOC_269/a_8_216# OR2X1_LOC_269/Y -0.00fF
C16187 VDD OR2X1_LOC_269/Y 0.12fF
C53021 OR2X1_LOC_269/Y AND2X1_LOC_271/a_8_24# 0.23fF
C56892 OR2X1_LOC_269/Y VSS 0.06fF
C22643 AND2X1_LOC_19/a_8_24# OR2X1_LOC_87/Y 0.01fF
C23039 AND2X1_LOC_29/a_8_24# OR2X1_LOC_87/Y 0.23fF
C30894 VDD OR2X1_LOC_87/Y 0.29fF
C39864 AND2X1_LOC_129/a_8_24# OR2X1_LOC_87/Y 0.02fF
C45970 AND2X1_LOC_88/a_8_24# OR2X1_LOC_87/Y 0.11fF
C54865 OR2X1_LOC_87/a_8_216# OR2X1_LOC_87/Y 0.01fF
C56876 OR2X1_LOC_87/Y VSS 0.19fF
C7661 OR2X1_LOC_666/A AND2X1_LOC_66/a_8_24# 0.01fF
C8070 AND2X1_LOC_120/a_8_24# OR2X1_LOC_666/A 0.01fF
C10875 VDD OR2X1_LOC_666/A 0.37fF
C52686 OR2X1_LOC_666/A OR2X1_LOC_67/A 0.01fF
C57518 OR2X1_LOC_666/A VSS 0.41fF
C12907 OR2X1_LOC_120/a_8_216# OR2X1_LOC_121/A 0.01fF
C15459 VDD OR2X1_LOC_121/A 0.12fF
C19351 OR2X1_LOC_274/a_8_216# OR2X1_LOC_121/A 0.01fF
C32341 OR2X1_LOC_121/a_8_216# OR2X1_LOC_121/A 0.08fF
C35839 OR2X1_LOC_274/Y OR2X1_LOC_121/A 0.01fF
C52947 AND2X1_LOC_255/a_8_24# OR2X1_LOC_121/A 0.01fF
C56242 OR2X1_LOC_121/A VSS 0.27fF
C2451 OR2X1_LOC_264/Y VDD 0.12fF
C7616 OR2X1_LOC_264/Y OR2X1_LOC_264/a_8_216# 0.05fF
C17091 OR2X1_LOC_264/Y AND2X1_LOC_88/Y 0.02fF
C57997 OR2X1_LOC_264/Y VSS 0.59fF
C40795 OR2X1_LOC_685/A AND2X1_LOC_681/a_8_24# 0.20fF
C50167 VDD OR2X1_LOC_685/A 0.21fF
C57714 OR2X1_LOC_685/A VSS 0.21fF
C13410 VDD OR2X1_LOC_816/A 0.32fF
C27483 OR2X1_LOC_530/Y OR2X1_LOC_816/A 0.02fF
C32974 AND2X1_LOC_548/a_8_24# OR2X1_LOC_816/A 0.01fF
C36184 OR2X1_LOC_816/A OR2X1_LOC_753/a_8_216# 0.02fF
C41740 OR2X1_LOC_816/A OR2X1_LOC_753/a_36_216# 0.02fF
C42242 OR2X1_LOC_628/a_8_216# OR2X1_LOC_816/A 0.01fF
C53797 OR2X1_LOC_816/A OR2X1_LOC_530/a_8_216# 0.01fF
C56724 OR2X1_LOC_816/A VSS 0.44fF
C400 OR2X1_LOC_684/a_8_216# AND2X1_LOC_687/B 0.47fF
C25677 AND2X1_LOC_687/B AND2X1_LOC_687/a_8_24# 0.01fF
C34408 OR2X1_LOC_694/a_8_216# AND2X1_LOC_687/B 0.02fF
C49582 AND2X1_LOC_686/a_8_24# AND2X1_LOC_687/B 0.04fF
C53649 VDD AND2X1_LOC_687/B 0.06fF
C57003 AND2X1_LOC_687/B VSS 0.06fF
C49923 OR2X1_LOC_275/A AND2X1_LOC_264/a_8_24# 0.01fF
C57257 OR2X1_LOC_275/A VSS 0.06fF
C18160 OR2X1_LOC_461/B AND2X1_LOC_233/a_8_24# 0.20fF
C45707 VDD OR2X1_LOC_461/B 0.21fF
C56738 OR2X1_LOC_461/B VSS 0.19fF
C49445 OR2X1_LOC_271/B OR2X1_LOC_271/a_8_216# 0.06fF
C57498 OR2X1_LOC_271/B VSS 0.06fF
C9808 OR2X1_LOC_847/A AND2X1_LOC_817/a_8_24# 0.01fF
C9828 AND2X1_LOC_490/a_8_24# OR2X1_LOC_847/A 0.06fF
C35827 OR2X1_LOC_847/A AND2X1_LOC_619/a_8_24# 0.01fF
C46427 OR2X1_LOC_847/A OR2X1_LOC_5/a_8_216# 0.47fF
C51423 OR2X1_LOC_847/A AND2X1_LOC_819/a_8_24# 0.01fF
C55604 VDD OR2X1_LOC_847/A 0.28fF
C16061 VDD OR2X1_LOC_687/B -0.00fF
C25119 OR2X1_LOC_685/a_8_216# OR2X1_LOC_687/B -0.00fF
C46485 OR2X1_LOC_687/B OR2X1_LOC_687/a_8_216# 0.39fF
C57712 OR2X1_LOC_687/B VSS 0.17fF
C16384 VDD OR2X1_LOC_274/Y 0.09fF
C30385 OR2X1_LOC_274/Y AND2X1_LOC_275/a_8_24# 0.01fF
C57304 OR2X1_LOC_274/Y VSS 0.07fF
C607 OR2X1_LOC_329/B OR2X1_LOC_310/a_8_216# 0.12fF
C7708 OR2X1_LOC_329/B OR2X1_LOC_760/a_8_216# 0.05fF
C13017 OR2X1_LOC_329/a_8_216# OR2X1_LOC_329/B 0.04fF
C13293 OR2X1_LOC_329/B OR2X1_LOC_760/a_36_216# 0.02fF
C16428 OR2X1_LOC_329/B AND2X1_LOC_276/a_36_24# 0.01fF
C21103 VDD OR2X1_LOC_329/B 0.42fF
C29384 OR2X1_LOC_329/B AND2X1_LOC_405/a_8_24# 0.03fF
C40358 OR2X1_LOC_329/B AND2X1_LOC_405/a_36_24# 0.01fF
C41128 OR2X1_LOC_329/B AND2X1_LOC_327/a_8_24# 0.01fF
C41796 OR2X1_LOC_329/B OR2X1_LOC_373/Y 0.07fF
C42024 OR2X1_LOC_329/B OR2X1_LOC_268/a_8_216# 0.02fF
C47747 OR2X1_LOC_329/B OR2X1_LOC_268/a_36_216# 0.01fF
C56049 OR2X1_LOC_329/B AND2X1_LOC_276/a_8_24# 0.03fF
C57709 OR2X1_LOC_329/B VSS -2.21fF
C2979 OR2X1_LOC_405/A OR2X1_LOC_405/a_8_216# 0.16fF
C11829 OR2X1_LOC_405/A AND2X1_LOC_372/a_8_24# 0.01fF
C25883 OR2X1_LOC_405/A AND2X1_LOC_272/a_8_24# -0.01fF
C37125 OR2X1_LOC_405/A OR2X1_LOC_185/a_8_216# 0.06fF
C40990 OR2X1_LOC_405/A VDD 1.35fF
C54740 OR2X1_LOC_405/A AND2X1_LOC_371/a_8_24# 0.01fF
C57996 OR2X1_LOC_405/A VSS 0.50fF
C7676 OR2X1_LOC_683/a_8_216# OR2X1_LOC_683/Y -0.00fF
C27320 OR2X1_LOC_683/Y AND2X1_LOC_686/a_8_24# 0.23fF
C31386 VDD OR2X1_LOC_683/Y 0.12fF
C57005 OR2X1_LOC_683/Y VSS 0.06fF
C12492 AND2X1_LOC_512/a_8_24# OR2X1_LOC_599/Y 0.09fF
C10180 VDD OR2X1_LOC_530/Y 0.16fF
C29801 OR2X1_LOC_530/Y AND2X1_LOC_548/a_8_24# 0.23fF
C57622 OR2X1_LOC_530/Y VSS 0.07fF
C11947 OR2X1_LOC_682/a_8_216# OR2X1_LOC_682/Y 0.01fF
C12279 OR2X1_LOC_682/Y VDD 0.05fF
C23074 OR2X1_LOC_682/a_36_216# OR2X1_LOC_682/Y -0.00fF
C36127 OR2X1_LOC_682/Y AND2X1_LOC_685/a_8_24# 0.01fF
C55288 OR2X1_LOC_682/Y OR2X1_LOC_421/a_8_216# 0.39fF
C57888 OR2X1_LOC_682/Y VSS 0.20fF
C15442 OR2X1_LOC_373/a_8_216# OR2X1_LOC_373/Y 0.03fF
C21820 OR2X1_LOC_373/Y OR2X1_LOC_164/a_8_216# 0.01fF
C25123 OR2X1_LOC_373/Y AND2X1_LOC_405/a_8_24# 0.03fF
C2048 AND2X1_LOC_121/a_8_24# OR2X1_LOC_67/A 0.21fF
C37597 VDD OR2X1_LOC_67/A 0.21fF
C46336 OR2X1_LOC_625/a_8_216# OR2X1_LOC_67/A 0.07fF
C56755 OR2X1_LOC_67/A VSS 0.43fF
C22835 OR2X1_LOC_410/Y AND2X1_LOC_411/a_8_24# 0.23fF
C34554 VDD OR2X1_LOC_410/Y 0.16fF
C56739 OR2X1_LOC_410/Y VSS 0.07fF
C10030 VDD OR2X1_LOC_411/A -0.00fF
C14924 OR2X1_LOC_411/A OR2X1_LOC_411/a_8_216# 0.47fF
C56800 OR2X1_LOC_411/A VSS 0.15fF
C15025 OR2X1_LOC_271/a_8_216# OR2X1_LOC_368/A 0.47fF
C20203 AND2X1_LOC_270/a_8_24# OR2X1_LOC_368/A 0.01fF
C56940 OR2X1_LOC_368/A VSS 0.28fF
C27649 OR2X1_LOC_689/Y AND2X1_LOC_691/a_8_24# 0.23fF
C28892 VDD OR2X1_LOC_689/Y 0.12fF
C57319 OR2X1_LOC_689/Y VSS 0.06fF
C21026 OR2X1_LOC_376/A OR2X1_LOC_376/a_8_216# 0.47fF
C57782 OR2X1_LOC_376/A VSS 0.15fF
C19600 OR2X1_LOC_800/A OR2X1_LOC_800/a_8_216# 0.47fF
C57734 OR2X1_LOC_800/A VSS -0.07fF
C24713 OR2X1_LOC_686/B AND2X1_LOC_684/a_8_24# 0.25fF
C30367 VDD OR2X1_LOC_686/B 0.21fF
C35658 OR2X1_LOC_686/B AND2X1_LOC_684/a_36_24# 0.01fF
C39310 OR2X1_LOC_686/B AND2X1_LOC_682/a_8_24# 0.04fF
C43697 OR2X1_LOC_686/B AND2X1_LOC_683/a_8_24# 0.03fF
C57650 OR2X1_LOC_686/B VSS 0.20fF
C4074 OR2X1_LOC_276/a_36_216# OR2X1_LOC_66/Y 0.02fF
C6832 OR2X1_LOC_66/Y AND2X1_LOC_625/a_8_24# 0.01fF
C38213 VDD OR2X1_LOC_66/Y 0.19fF
C56818 OR2X1_LOC_66/Y VSS 0.16fF
C19381 OR2X1_LOC_800/Y OR2X1_LOC_801/a_8_216# 0.39fF
C57677 OR2X1_LOC_800/Y VSS 0.18fF
C8472 VDD OR2X1_LOC_271/Y 0.28fF
C57497 OR2X1_LOC_271/Y VSS 0.26fF
C5317 OR2X1_LOC_276/B AND2X1_LOC_268/a_8_24# 0.02fF
C6813 VDD OR2X1_LOC_276/B 0.02fF
C19134 OR2X1_LOC_276/B AND2X1_LOC_256/a_8_24# 0.01fF
C20054 OR2X1_LOC_276/B AND2X1_LOC_628/a_8_24# 0.02fF
C20877 OR2X1_LOC_276/B AND2X1_LOC_275/a_8_24# 0.02fF
C23215 OR2X1_LOC_276/B OR2X1_LOC_276/a_8_216# 0.02fF
C43537 OR2X1_LOC_276/B AND2X1_LOC_271/a_8_24# 0.02fF
C55870 OR2X1_LOC_276/B OR2X1_LOC_269/a_8_216# 0.01fF
C57203 OR2X1_LOC_276/B VSS 0.21fF
C33082 VDD AND2X1_LOC_801/B 0.16fF
C34410 AND2X1_LOC_801/B AND2X1_LOC_801/a_8_24# 0.07fF
C57083 AND2X1_LOC_801/B VSS -0.07fF
C7295 OR2X1_LOC_687/Y OR2X1_LOC_687/a_8_216# 0.01fF
C23966 OR2X1_LOC_687/Y AND2X1_LOC_681/a_8_24# 0.06fF
C25105 OR2X1_LOC_687/Y OR2X1_LOC_800/a_8_216# 0.01fF
C29156 OR2X1_LOC_687/Y OR2X1_LOC_185/a_8_216# 0.03fF
C32989 VDD OR2X1_LOC_687/Y 0.28fF
C42026 OR2X1_LOC_687/Y OR2X1_LOC_685/a_8_216# 0.04fF
C46481 OR2X1_LOC_687/Y AND2X1_LOC_430/a_8_24# 0.23fF
C52604 OR2X1_LOC_687/Y AND2X1_LOC_760/a_8_24# 0.02fF
C57733 OR2X1_LOC_687/Y VSS 0.27fF
C16565 VDD AND2X1_LOC_687/Y 0.04fF
C57084 AND2X1_LOC_687/Y VSS 0.29fF

.ends

* wrdata outputs.out V("OR2X1_LOC_515/Y") V("OR2X1_LOC_751/A") V("OR2X1_LOC_334/A") V("OR2X1_LOC_836/A") V("OR2X1_LOC_240/A") V("OR2X1_LOC_461/Y") V("AND2X1_LOC_809/A") V("AND2X1_LOC_276/Y") V("OR2X1_LOC_100/Y") V("OR2X1_LOC_516/B") V("AND2X1_LOC_729/B") V("OR2X1_LOC_527/Y") V("OR2X1_LOC_111/Y") V("OR2X1_LOC_323/Y") V("AND2X1_LOC_155/Y") V("OR2X1_LOC_273/Y") V("OR2X1_LOC_433/Y") V("OR2X1_LOC_743/Y") V("OR2X1_LOC_409/B") V("AND2X1_LOC_458/Y") V("OR2X1_LOC_519/Y") V("OR2X1_LOC_692/Y") V("OR2X1_LOC_599/A") V("OR2X1_LOC_763/Y") V("OR2X1_LOC_48/Y") V("OR2X1_LOC_406/A") V("OR2X1_LOC_511/Y") V("OR2X1_LOC_604/A") V("OR2X1_LOC_235/B") V("OR2X1_LOC_246/Y") V("OR2X1_LOC_74/A") V("OR2X1_LOC_13/B") V("OR2X1_LOC_16/A") V("OR2X1_LOC_287/B") V("OR2X1_LOC_637/B") V("OR2X1_LOC_294/Y") V("OR2X1_LOC_415/Y") V("OR2X1_LOC_631/A") V("OR2X1_LOC_598/Y") V("OR2X1_LOC_398/Y") V("OR2X1_LOC_309/Y") V("OR2X1_LOC_283/Y") V("OR2X1_LOC_488/Y") V("OR2X1_LOC_289/Y") V("OR2X1_LOC_417/Y") V("OR2X1_LOC_226/Y") V("OR2X1_LOC_815/A") V("OR2X1_LOC_121/Y") V("OR2X1_LOC_831/A") V("OR2X1_LOC_543/A") V("OR2X1_LOC_606/Y") V("OR2X1_LOC_302/A") V("OR2X1_LOC_450/B") V("AND2X1_LOC_847/Y") V("AND2X1_LOC_91/B") V("OR2X1_LOC_611/Y") V("AND2X1_LOC_56/B") V("OR2X1_LOC_78/A") V("OR2X1_LOC_532/B") V("OR2X1_LOC_96/B") V("OR2X1_LOC_71/A") V("OR2X1_LOC_535/A") V("OR2X1_LOC_195/A") V("OR2X1_LOC_296/Y") V("OR2X1_LOC_138/A") V("OR2X1_LOC_541/A") V("OR2X1_LOC_838/B") V("OR2X1_LOC_506/A") V("OR2X1_LOC_378/Y") V("OR2X1_LOC_98/B") V("OR2X1_LOC_389/A") V("OR2X1_LOC_448/A") V("OR2X1_LOC_630/B") V("OR2X1_LOC_144/Y") V("OR2X1_LOC_306/Y") V("OR2X1_LOC_503/A") V("OR2X1_LOC_696/Y") V("OR2X1_LOC_588/Y") V("OR2X1_LOC_376/Y") V("OR2X1_LOC_322/Y") V("OR2X1_LOC_164/Y") V("OR2X1_LOC_673/A") V("OR2X1_LOC_693/Y") V("AND2X1_LOC_377/Y") V("OR2X1_LOC_748/A") V("OR2X1_LOC_83/A") V("OR2X1_LOC_89/A") V("OR2X1_LOC_45/B") V("OR2X1_LOC_52/B") V("OR2X1_LOC_619/Y") V("OR2X1_LOC_151/A") V("OR2X1_LOC_185/A") V("AND2X1_LOC_86/B") V("OR2X1_LOC_160/A") V("OR2X1_LOC_154/A") V("OR2X1_LOC_130/A") V("OR2X1_LOC_266/A") V("OR2X1_LOC_634/A") V("OR2X1_LOC_541/B") V("OR2X1_LOC_633/A") V("OR2X1_LOC_777/B") V("OR2X1_LOC_549/A") V("OR2X1_LOC_391/B") V("OR2X1_LOC_387/Y") V("OR2X1_LOC_597/A") V("OR2X1_LOC_329/Y") V("OR2X1_LOC_421/Y") V("OR2X1_LOC_304/Y") V("OR2X1_LOC_56/Y") V("OR2X1_LOC_158/A") V("OR2X1_LOC_70/Y") V("OR2X1_LOC_3/Y") V("OR2X1_LOC_40/Y") V("OR2X1_LOC_694/Y") V("OR2X1_LOC_426/Y") V("AND2X1_LOC_51/Y") V("AND2X1_LOC_31/Y") V("AND2X1_LOC_44/Y") V("AND2X1_LOC_47/Y") V("OR2X1_LOC_790/B") V("OR2X1_LOC_635/A") V("OR2X1_LOC_769/B") V("OR2X1_LOC_409/Y") V("OR2X1_LOC_430/Y") V("OR2X1_LOC_51/Y") V("OR2X1_LOC_95/Y") V("OR2X1_LOC_64/Y") V("OR2X1_LOC_375/A") V("AND2X1_LOC_36/Y") V("AND2X1_LOC_18/Y") V("OR2X1_LOC_809/B") V("OR2X1_LOC_513/Y") V("OR2X1_LOC_473/A") V("AND2X1_LOC_101/B") V("OR2X1_LOC_600/A") V("OR2X1_LOC_744/A") V("OR2X1_LOC_557/A") V("AND2X1_LOC_19/Y") V("OR2X1_LOC_7/A") V("OR2X1_LOC_344/A") V("OR2X1_LOC_748/Y") V("OR2X1_LOC_589/A") V("OR2X1_LOC_161/B") V("OR2X1_LOC_80/Y") V("OR2X1_LOC_87/A") V("OR2X1_LOC_32/B") V("OR2X1_LOC_269/B") V("OR2X1_LOC_291/Y") V("OR2X1_LOC_824/Y") V("OR2X1_LOC_234/Y") V("AND2X1_LOC_462/B") V("OR2X1_LOC_691/Y") V("OR2X1_LOC_325/A") V("OR2X1_LOC_547/B") V("OR2X1_LOC_112/A") V("OR2X1_LOC_516/A") V("OR2X1_LOC_750/Y") V("OR2X1_LOC_814/Y") V("OR2X1_LOC_335/B") V("OR2X1_LOC_286/B") V("OR2X1_LOC_489/A") V("OR2X1_LOC_333/A") V("OR2X1_LOC_446/B") V("OR2X1_LOC_227/A") V("OR2X1_LOC_427/A") V("AND2X1_LOC_81/B") V("AND2X1_LOC_82/Y") V("OR2X1_LOC_87/B") V("OR2X1_LOC_428/A") V("OR2X1_LOC_382/Y") V("OR2X1_LOC_39/A") V("OR2X1_LOC_848/A") V("AND2X1_LOC_41/A") V("OR2X1_LOC_161/A") V("OR2X1_LOC_78/B") V("OR2X1_LOC_278/Y") V("OR2X1_LOC_342/B") V("OR2X1_LOC_485/A") V("AND2X1_LOC_94/Y") V("OR2X1_LOC_91/A") V("AND2X1_LOC_612/B") V("OR2X1_LOC_56/A") V("OR2X1_LOC_136/Y") V("OR2X1_LOC_459/A") V("OR2X1_LOC_272/Y") V("OR2X1_LOC_827/Y") V("OR2X1_LOC_419/Y") V("OR2X1_LOC_43/Y") V("OR2X1_LOC_297/A") V("OR2X1_LOC_534/Y") V("OR2X1_LOC_490/Y") V("OR2X1_LOC_789/B") V("OR2X1_LOC_160/B") V("OR2X1_LOC_756/B") V("OR2X1_LOC_256/Y") V("AND2X1_LOC_7/B") V("OR2X1_LOC_20/A") V("OR2X1_LOC_422/Y") V("OR2X1_LOC_628/Y") V("OR2X1_LOC_93/Y") V("OR2X1_LOC_779/B") V("OR2X1_LOC_520/A") V("OR2X1_LOC_706/B") V("AND2X1_LOC_48/Y") V("OR2X1_LOC_405/Y") V("OR2X1_LOC_399/A") V("OR2X1_LOC_625/Y") V("OR2X1_LOC_481/A") V("OR2X1_LOC_585/Y") V("OR2X1_LOC_416/A") V("OR2X1_LOC_638/B") V("OR2X1_LOC_459/B") V("OR2X1_LOC_325/B") V("OR2X1_LOC_168/B") V("OR2X1_LOC_147/A") V("OR2X1_LOC_512/A") V("OR2X1_LOC_708/B") V("OR2X1_LOC_502/Y") V("OR2X1_LOC_156/A") V("OR2X1_LOC_780/B") V("OR2X1_LOC_828/B") V("OR2X1_LOC_831/B") V("OR2X1_LOC_435/A") V("OR2X1_LOC_369/Y") V("OR2X1_LOC_122/A") V("OR2X1_LOC_299/Y") V("OR2X1_LOC_607/A") V("OR2X1_LOC_300/Y") V("OR2X1_LOC_464/A") V("OR2X1_LOC_65/B") V("OR2X1_LOC_778/B") V("AND2X1_LOC_72/B") V("OR2X1_LOC_335/A") V("AND2X1_LOC_57/Y") V("OR2X1_LOC_68/Y") V("OR2X1_LOC_672/Y") V("OR2X1_LOC_622/B") V("OR2X1_LOC_813/A") V("OR2X1_LOC_690/A") V("OR2X1_LOC_256/A") V("OR2X1_LOC_278/A") V("OR2X1_LOC_246/A") V("OR2X1_LOC_86/A") V("OR2X1_LOC_437/A") V("AND2X1_LOC_65/A") V("OR2X1_LOC_69/A") V("OR2X1_LOC_71/Y") V("OR2X1_LOC_57/Y") V("OR2X1_LOC_371/Y") V("OR2X1_LOC_310/Y") V("OR2X1_LOC_706/A") V("OR2X1_LOC_709/A") V("OR2X1_LOC_378/A") V("AND2X1_LOC_548/Y") V("OR2X1_LOC_22/Y") V("OR2X1_LOC_36/Y") V("OR2X1_LOC_26/Y") V("OR2X1_LOC_355/B") V("OR2X1_LOC_448/B") V("OR2X1_LOC_596/Y") V("AND2X1_LOC_95/Y") V("AND2X1_LOC_12/Y") V("AND2X1_LOC_59/Y") V("OR2X1_LOC_707/B") V("OR2X1_LOC_753/Y") V("OR2X1_LOC_12/Y") V("OR2X1_LOC_59/Y") V("OR2X1_LOC_18/Y") V("OR2X1_LOC_31/Y") V("OR2X1_LOC_44/Y") V("OR2X1_LOC_47/Y") V("AND2X1_LOC_70/Y") V("AND2X1_LOC_40/Y") V("AND2X1_LOC_3/Y") V("AND2X1_LOC_64/Y") V("AND2X1_LOC_22/Y") V("OR2X1_LOC_66/A") V("OR2X1_LOC_307/B") V("OR2X1_LOC_197/A") V("OR2X1_LOC_460/A") V("OR2X1_LOC_582/Y") V("OR2X1_LOC_451/A") V("OR2X1_LOC_329/B") V("OR2X1_LOC_66/Y") V("OR2X1_LOC_121/A") V("OR2X1_LOC_185/Y") V("OR2X1_LOC_405/A") V("OR2X1_LOC_67/A") V("OR2X1_LOC_666/A") V("OR2X1_LOC_816/A") V("OR2X1_LOC_410/Y") V("AND2X1_LOC_687/Y") V("OR2X1_LOC_368/A") V("OR2X1_LOC_87/Y") V("OR2X1_LOC_373/Y") V("OR2X1_LOC_517/A") V("OR2X1_LOC_687/Y") V("OR2X1_LOC_270/Y") V("OR2X1_LOC_88/A") V("OR2X1_LOC_411/A") V("OR2X1_LOC_264/Y") V("OR2X1_LOC_544/B") V("OR2X1_LOC_682/Y") V("OR2X1_LOC_683/Y") V("OR2X1_LOC_686/B") V("OR2X1_LOC_685/A") V("OR2X1_LOC_88/Y") V("AND2X1_LOC_374/Y") V("OR2X1_LOC_599/Y") V("OR2X1_LOC_644/A") V("AND2X1_LOC_88/Y") V("OR2X1_LOC_374/Y") 

* SUBCKT HEAD: NAME;  INPUTS; POWER; OUTPUTS
.subckt AES_SBOX_1
+ OR2X1_LOC_515/Y OR2X1_LOC_751/A OR2X1_LOC_334/A OR2X1_LOC_836/A OR2X1_LOC_240/A OR2X1_LOC_461/Y AND2X1_LOC_809/A AND2X1_LOC_276/Y OR2X1_LOC_100/Y OR2X1_LOC_516/B AND2X1_LOC_729/B OR2X1_LOC_527/Y OR2X1_LOC_111/Y OR2X1_LOC_323/Y AND2X1_LOC_155/Y OR2X1_LOC_273/Y OR2X1_LOC_433/Y OR2X1_LOC_743/Y OR2X1_LOC_409/B AND2X1_LOC_458/Y OR2X1_LOC_519/Y OR2X1_LOC_692/Y OR2X1_LOC_599/A OR2X1_LOC_763/Y OR2X1_LOC_48/Y OR2X1_LOC_406/A OR2X1_LOC_511/Y OR2X1_LOC_604/A OR2X1_LOC_235/B OR2X1_LOC_246/Y OR2X1_LOC_74/A OR2X1_LOC_13/B OR2X1_LOC_16/A OR2X1_LOC_287/B OR2X1_LOC_637/B OR2X1_LOC_294/Y OR2X1_LOC_415/Y OR2X1_LOC_631/A OR2X1_LOC_598/Y OR2X1_LOC_398/Y OR2X1_LOC_309/Y OR2X1_LOC_283/Y OR2X1_LOC_488/Y OR2X1_LOC_289/Y OR2X1_LOC_417/Y OR2X1_LOC_226/Y OR2X1_LOC_815/A OR2X1_LOC_121/Y OR2X1_LOC_831/A OR2X1_LOC_543/A OR2X1_LOC_606/Y 
+ OR2X1_LOC_302/A OR2X1_LOC_450/B AND2X1_LOC_847/Y AND2X1_LOC_91/B OR2X1_LOC_611/Y AND2X1_LOC_56/B OR2X1_LOC_78/A OR2X1_LOC_532/B OR2X1_LOC_96/B OR2X1_LOC_71/A OR2X1_LOC_535/A OR2X1_LOC_195/A OR2X1_LOC_296/Y OR2X1_LOC_138/A OR2X1_LOC_541/A OR2X1_LOC_838/B OR2X1_LOC_506/A OR2X1_LOC_378/Y OR2X1_LOC_98/B OR2X1_LOC_389/A OR2X1_LOC_448/A OR2X1_LOC_630/B OR2X1_LOC_144/Y OR2X1_LOC_306/Y OR2X1_LOC_503/A OR2X1_LOC_696/Y OR2X1_LOC_588/Y OR2X1_LOC_376/Y OR2X1_LOC_322/Y OR2X1_LOC_164/Y OR2X1_LOC_673/A OR2X1_LOC_693/Y AND2X1_LOC_377/Y OR2X1_LOC_748/A OR2X1_LOC_83/A OR2X1_LOC_89/A OR2X1_LOC_45/B OR2X1_LOC_52/B OR2X1_LOC_619/Y OR2X1_LOC_151/A OR2X1_LOC_185/A AND2X1_LOC_86/B OR2X1_LOC_160/A OR2X1_LOC_154/A OR2X1_LOC_130/A OR2X1_LOC_266/A OR2X1_LOC_634/A OR2X1_LOC_541/B OR2X1_LOC_633/A OR2X1_LOC_777/B OR2X1_LOC_549/A 
+ OR2X1_LOC_391/B OR2X1_LOC_387/Y OR2X1_LOC_597/A OR2X1_LOC_329/Y OR2X1_LOC_421/Y OR2X1_LOC_304/Y OR2X1_LOC_56/Y OR2X1_LOC_158/A OR2X1_LOC_70/Y OR2X1_LOC_3/Y OR2X1_LOC_40/Y OR2X1_LOC_694/Y OR2X1_LOC_426/Y AND2X1_LOC_51/Y AND2X1_LOC_31/Y AND2X1_LOC_44/Y AND2X1_LOC_47/Y OR2X1_LOC_790/B OR2X1_LOC_635/A OR2X1_LOC_769/B OR2X1_LOC_409/Y OR2X1_LOC_430/Y OR2X1_LOC_51/Y OR2X1_LOC_95/Y OR2X1_LOC_64/Y OR2X1_LOC_375/A AND2X1_LOC_36/Y AND2X1_LOC_18/Y OR2X1_LOC_809/B OR2X1_LOC_513/Y OR2X1_LOC_473/A AND2X1_LOC_101/B OR2X1_LOC_600/A OR2X1_LOC_744/A OR2X1_LOC_557/A AND2X1_LOC_19/Y OR2X1_LOC_7/A OR2X1_LOC_344/A OR2X1_LOC_748/Y OR2X1_LOC_589/A OR2X1_LOC_161/B OR2X1_LOC_80/Y OR2X1_LOC_87/A OR2X1_LOC_32/B OR2X1_LOC_269/B OR2X1_LOC_291/Y OR2X1_LOC_824/Y OR2X1_LOC_234/Y AND2X1_LOC_462/B OR2X1_LOC_691/Y OR2X1_LOC_325/A 
+ OR2X1_LOC_547/B OR2X1_LOC_112/A OR2X1_LOC_516/A OR2X1_LOC_750/Y OR2X1_LOC_814/Y OR2X1_LOC_335/B OR2X1_LOC_286/B OR2X1_LOC_489/A OR2X1_LOC_333/A OR2X1_LOC_446/B OR2X1_LOC_227/A OR2X1_LOC_427/A AND2X1_LOC_81/B AND2X1_LOC_82/Y OR2X1_LOC_87/B OR2X1_LOC_428/A OR2X1_LOC_382/Y OR2X1_LOC_39/A OR2X1_LOC_848/A AND2X1_LOC_41/A OR2X1_LOC_161/A OR2X1_LOC_78/B OR2X1_LOC_278/Y OR2X1_LOC_342/B OR2X1_LOC_485/A AND2X1_LOC_94/Y OR2X1_LOC_91/A AND2X1_LOC_612/B OR2X1_LOC_56/A OR2X1_LOC_136/Y OR2X1_LOC_459/A OR2X1_LOC_272/Y OR2X1_LOC_827/Y OR2X1_LOC_419/Y OR2X1_LOC_43/Y OR2X1_LOC_297/A OR2X1_LOC_534/Y OR2X1_LOC_490/Y OR2X1_LOC_789/B OR2X1_LOC_160/B OR2X1_LOC_756/B OR2X1_LOC_256/Y AND2X1_LOC_7/B OR2X1_LOC_20/A OR2X1_LOC_422/Y OR2X1_LOC_628/Y OR2X1_LOC_93/Y OR2X1_LOC_779/B OR2X1_LOC_520/A OR2X1_LOC_706/B AND2X1_LOC_48/Y 
+ OR2X1_LOC_405/Y OR2X1_LOC_399/A OR2X1_LOC_625/Y OR2X1_LOC_481/A OR2X1_LOC_585/Y OR2X1_LOC_416/A OR2X1_LOC_638/B OR2X1_LOC_459/B OR2X1_LOC_325/B OR2X1_LOC_168/B OR2X1_LOC_147/A OR2X1_LOC_512/A OR2X1_LOC_708/B OR2X1_LOC_502/Y OR2X1_LOC_156/A OR2X1_LOC_780/B OR2X1_LOC_828/B OR2X1_LOC_831/B OR2X1_LOC_435/A OR2X1_LOC_369/Y OR2X1_LOC_122/A OR2X1_LOC_299/Y OR2X1_LOC_607/A OR2X1_LOC_300/Y OR2X1_LOC_464/A OR2X1_LOC_65/B OR2X1_LOC_778/B AND2X1_LOC_72/B OR2X1_LOC_335/A AND2X1_LOC_57/Y OR2X1_LOC_68/Y OR2X1_LOC_672/Y OR2X1_LOC_622/B OR2X1_LOC_813/A OR2X1_LOC_690/A OR2X1_LOC_256/A OR2X1_LOC_278/A OR2X1_LOC_246/A OR2X1_LOC_86/A OR2X1_LOC_437/A AND2X1_LOC_65/A OR2X1_LOC_69/A OR2X1_LOC_71/Y OR2X1_LOC_57/Y OR2X1_LOC_371/Y OR2X1_LOC_310/Y OR2X1_LOC_706/A OR2X1_LOC_709/A OR2X1_LOC_378/A AND2X1_LOC_548/Y OR2X1_LOC_22/Y 
+ OR2X1_LOC_36/Y OR2X1_LOC_26/Y OR2X1_LOC_355/B OR2X1_LOC_448/B OR2X1_LOC_596/Y AND2X1_LOC_95/Y AND2X1_LOC_12/Y AND2X1_LOC_59/Y OR2X1_LOC_707/B OR2X1_LOC_753/Y OR2X1_LOC_12/Y OR2X1_LOC_59/Y OR2X1_LOC_18/Y OR2X1_LOC_31/Y OR2X1_LOC_44/Y OR2X1_LOC_47/Y AND2X1_LOC_70/Y AND2X1_LOC_40/Y AND2X1_LOC_3/Y AND2X1_LOC_64/Y AND2X1_LOC_22/Y OR2X1_LOC_66/A OR2X1_LOC_307/B OR2X1_LOC_197/A OR2X1_LOC_460/A OR2X1_LOC_582/Y OR2X1_LOC_451/A OR2X1_LOC_329/B OR2X1_LOC_66/Y OR2X1_LOC_121/A OR2X1_LOC_185/Y OR2X1_LOC_405/A OR2X1_LOC_67/A OR2X1_LOC_666/A OR2X1_LOC_816/A OR2X1_LOC_410/Y AND2X1_LOC_687/Y OR2X1_LOC_368/A OR2X1_LOC_87/Y OR2X1_LOC_373/Y OR2X1_LOC_517/A OR2X1_LOC_687/Y OR2X1_LOC_270/Y OR2X1_LOC_88/A OR2X1_LOC_411/A OR2X1_LOC_264/Y OR2X1_LOC_544/B OR2X1_LOC_682/Y OR2X1_LOC_683/Y OR2X1_LOC_686/B OR2X1_LOC_685/A 
+ OR2X1_LOC_88/Y AND2X1_LOC_374/Y OR2X1_LOC_599/Y OR2X1_LOC_644/A AND2X1_LOC_88/Y OR2X1_LOC_374/Y 
+ VSS VDD 
+ OR2X1_LOC_452/A AND2X1_LOC_639/A OR2X1_LOC_460/Y OR2X1_LOC_198/A OR2X1_LOC_308/A OR2X1_LOC_379/Y OR2X1_LOC_643/A OR2X1_LOC_84/A OR2X1_LOC_538/A OR2X1_LOC_180/B OR2X1_LOC_668/Y OR2X1_LOC_34/B OR2X1_LOC_334/B OR2X1_LOC_834/A OR2X1_LOC_241/B OR2X1_LOC_523/A OR2X1_LOC_33/A OR2X1_LOC_61/B OR2X1_LOC_844/B OR2X1_LOC_623/B OR2X1_LOC_770/A OR2X1_LOC_324/A OR2X1_LOC_509/A OR2X1_LOC_703/A OR2X1_LOC_147/B OR2X1_LOC_201/A OR2X1_LOC_520/B OR2X1_LOC_703/B OR2X1_LOC_835/A OR2X1_LOC_709/B OR2X1_LOC_720/B OR2X1_LOC_343/B OR2X1_LOC_855/A OR2X1_LOC_449/B OR2X1_LOC_593/B OR2X1_LOC_773/B OR2X1_LOC_402/B OR2X1_LOC_307/A OR2X1_LOC_128/A OR2X1_LOC_194/B OR2X1_LOC_555/A OR2X1_LOC_719/B AND2X1_LOC_7/Y OR2X1_LOC_789/A OR2X1_LOC_769/A OR2X1_LOC_400/B OR2X1_LOC_781/B OR2X1_LOC_549/B OR2X1_LOC_391/A OR2X1_LOC_333/B OR2X1_LOC_190/B 
+ AND2X1_LOC_41/Y OR2X1_LOC_610/Y OR2X1_LOC_191/B OR2X1_LOC_169/B OR2X1_LOC_673/B OR2X1_LOC_346/B OR2X1_LOC_545/B OR2X1_LOC_444/B OR2X1_LOC_620/A OR2X1_LOC_786/A OR2X1_LOC_641/A OR2X1_LOC_758/Y OR2X1_LOC_637/A OR2X1_LOC_174/A AND2X1_LOC_72/Y OR2X1_LOC_175/B OR2X1_LOC_439/B OR2X1_LOC_835/B OR2X1_LOC_123/B OR2X1_LOC_633/B OR2X1_LOC_675/A OR2X1_LOC_501/B OR2X1_LOC_605/A OR2X1_LOC_544/A OR2X1_LOC_450/A OR2X1_LOC_103/Y OR2X1_LOC_106/Y OR2X1_LOC_695/Y OR2X1_LOC_280/Y OR2X1_LOC_601/Y OR2X1_LOC_612/B OR2X1_LOC_248/Y OR2X1_LOC_394/Y OR2X1_LOC_747/Y OR2X1_LOC_524/Y OR2X1_LOC_152/Y OR2X1_LOC_528/Y OR2X1_LOC_122/Y OR2X1_LOC_485/Y OR2X1_LOC_297/Y OR2X1_LOC_424/Y OR2X1_LOC_45/Y OR2X1_LOC_744/Y OR2X1_LOC_701/Y OR2X1_LOC_757/Y OR2X1_LOC_399/Y OR2X1_LOC_517/Y OR2X1_LOC_315/Y OR2X1_LOC_491/Y OR2X1_LOC_109/Y OR2X1_LOC_600/Y 
+ OR2X1_LOC_230/Y OR2X1_LOC_298/Y OR2X1_LOC_224/Y OR2X1_LOC_428/Y OR2X1_LOC_74/Y OR2X1_LOC_32/Y OR2X1_LOC_583/Y OR2X1_LOC_526/Y OR2X1_LOC_505/Y OR2X1_LOC_666/Y OR2X1_LOC_496/Y OR2X1_LOC_432/Y OR2X1_LOC_607/Y OR2X1_LOC_257/Y OR2X1_LOC_20/Y OR2X1_LOC_79/Y OR2X1_LOC_521/Y OR2X1_LOC_135/Y OR2X1_LOC_492/Y OR2X1_LOC_482/Y OR2X1_LOC_108/Y OR2X1_LOC_295/Y OR2X1_LOC_81/Y OR2X1_LOC_60/Y OR2X1_LOC_437/Y OR2X1_LOC_609/Y OR2X1_LOC_75/Y OR2X1_LOC_700/Y OR2X1_LOC_755/Y OR2X1_LOC_395/Y OR2X1_LOC_494/Y OR2X1_LOC_380/A OR2X1_LOC_603/Y OR2X1_LOC_261/A OR2X1_LOC_679/A OR2X1_LOC_229/Y OR2X1_LOC_13/Y OR2X1_LOC_765/Y OR2X1_LOC_131/Y AND2X1_LOC_793/B OR2X1_LOC_712/B OR2X1_LOC_791/B OR2X1_LOC_710/B OR2X1_LOC_401/B OR2X1_LOC_84/B OR2X1_LOC_61/A OR2X1_LOC_76/A OR2X1_LOC_702/A OR2X1_LOC_493/A OR2X1_LOC_833/B OR2X1_LOC_114/B 
+ OR2X1_LOC_346/A OR2X1_LOC_440/B OR2X1_LOC_646/A OR2X1_LOC_231/B OR2X1_LOC_770/B OR2X1_LOC_140/A OR2X1_LOC_260/Y OR2X1_LOC_678/Y OR2X1_LOC_193/A OR2X1_LOC_558/A OR2X1_LOC_605/B OR2X1_LOC_653/B OR2X1_LOC_788/B OR2X1_LOC_190/A OR2X1_LOC_98/A OR2X1_LOC_137/B OR2X1_LOC_192/B OR2X1_LOC_768/A OR2X1_LOC_128/B OR2X1_LOC_447/A OR2X1_LOC_489/B OR2X1_LOC_475/B OR2X1_LOC_644/B OR2X1_LOC_448/Y OR2X1_LOC_356/A OR2X1_LOC_176/Y OR2X1_LOC_290/Y OR2X1_LOC_677/Y OR2X1_LOC_83/Y OR2X1_LOC_237/Y OR2X1_LOC_669/A OR2X1_LOC_595/Y OR2X1_LOC_27/Y OR2X1_LOC_311/Y OR2X1_LOC_146/Y OR2X1_LOC_179/Y OR2X1_LOC_484/Y OR2X1_LOC_495/Y OR2X1_LOC_754/Y OR2X1_LOC_69/Y OR2X1_LOC_39/Y OR2X1_LOC_396/Y OR2X1_LOC_320/Y OR2X1_LOC_497/Y OR2X1_LOC_615/Y OR2X1_LOC_24/Y OR2X1_LOC_58/Y OR2X1_LOC_522/Y AND2X1_LOC_549/Y OR2X1_LOC_711/B OR2X1_LOC_713/A 
+ AND2X1_LOC_335/Y AND2X1_LOC_778/Y AND2X1_LOC_208/B OR2X1_LOC_72/Y OR2X1_LOC_184/Y OR2X1_LOC_152/A OR2X1_LOC_292/Y OR2X1_LOC_173/Y OR2X1_LOC_235/Y AND2X1_LOC_784/A AND2X1_LOC_633/Y AND2X1_LOC_541/Y AND2X1_LOC_634/Y OR2X1_LOC_813/Y OR2X1_LOC_624/B AND2X1_LOC_721/A AND2X1_LOC_69/Y OR2X1_LOC_208/A OR2X1_LOC_335/Y OR2X1_LOC_778/Y OR2X1_LOC_117/Y OR2X1_LOC_262/Y OR2X1_LOC_65/Y OR2X1_LOC_471/B AND2X1_LOC_303/A AND2X1_LOC_831/Y AND2X1_LOC_303/B AND2X1_LOC_787/A AND2X1_LOC_543/Y OR2X1_LOC_841/A OR2X1_LOC_841/B OR2X1_LOC_828/Y OR2X1_LOC_783/A OR2X1_LOC_156/Y OR2X1_LOC_708/Y OR2X1_LOC_308/Y OR2X1_LOC_149/B OR2X1_LOC_168/Y OR2X1_LOC_776/Y OR2X1_LOC_325/Y OR2X1_LOC_463/B OR2X1_LOC_651/B OR2X1_LOC_416/Y AND2X1_LOC_637/Y OR2X1_LOC_481/Y AND2X1_LOC_631/Y OR2X1_LOC_196/Y OR2X1_LOC_520/Y OR2X1_LOC_840/A OR2X1_LOC_779/Y AND2X1_LOC_632/A 
+ AND2X1_LOC_448/Y OR2X1_LOC_156/B OR2X1_LOC_636/A OR2X1_LOC_620/B OR2X1_LOC_247/Y OR2X1_LOC_231/A OR2X1_LOC_130/Y AND2X1_LOC_348/A OR2X1_LOC_105/Y OR2X1_LOC_181/A OR2X1_LOC_602/B OR2X1_LOC_345/A OR2X1_LOC_756/Y OR2X1_LOC_401/A OR2X1_LOC_507/A OR2X1_LOC_196/B OR2X1_LOC_707/A OR2X1_LOC_249/Y OR2X1_LOC_776/A OR2X1_LOC_793/B AND2X1_LOC_557/Y AND2X1_LOC_535/Y AND2X1_LOC_199/A AND2X1_LOC_508/A AND2X1_LOC_447/Y AND2X1_LOC_838/Y AND2X1_LOC_139/B OR2X1_LOC_178/Y OR2X1_LOC_613/Y OR2X1_LOC_67/Y OR2X1_LOC_312/Y OR2X1_LOC_647/B OR2X1_LOC_132/Y OR2X1_LOC_305/Y OR2X1_LOC_494/A OR2X1_LOC_91/Y OR2X1_LOC_766/Y OR2X1_LOC_670/Y OR2X1_LOC_533/A OR2X1_LOC_822/Y OR2X1_LOC_420/Y OR2X1_LOC_239/Y OR2X1_LOC_172/Y OR2X1_LOC_591/A OR2X1_LOC_349/B AND2X1_LOC_843/Y AND2X1_LOC_287/Y OR2X1_LOC_608/Y OR2X1_LOC_602/A OR2X1_LOC_78/Y OR2X1_LOC_240/B 
+ OR2X1_LOC_446/A OR2X1_LOC_546/A OR2X1_LOC_720/A OR2X1_LOC_546/B OR2X1_LOC_507/B OR2X1_LOC_486/B OR2X1_LOC_859/B AND2X1_LOC_154/Y OR2X1_LOC_189/A OR2X1_LOC_393/Y OR2X1_LOC_595/A AND2X1_LOC_391/Y OR2X1_LOC_823/Y OR2X1_LOC_697/Y OR2X1_LOC_759/Y OR2X1_LOC_34/A OR2X1_LOC_134/Y OR2X1_LOC_427/Y OR2X1_LOC_679/B OR2X1_LOC_754/A OR2X1_LOC_227/Y OR2X1_LOC_446/Y OR2X1_LOC_714/A OR2X1_LOC_338/B OR2X1_LOC_772/B OR2X1_LOC_286/Y OR2X1_LOC_787/B OR2X1_LOC_516/Y OR2X1_LOC_715/B OR2X1_LOC_339/A OR2X1_LOC_550/A OR2X1_LOC_856/A OR2X1_LOC_730/A AND2X1_LOC_462/Y AND2X1_LOC_240/Y AND2X1_LOC_839/B AND2X1_LOC_334/Y OR2X1_LOC_710/A OR2X1_LOC_792/B OR2X1_LOC_836/B OR2X1_LOC_779/A OR2X1_LOC_542/B OR2X1_LOC_383/Y OR2X1_LOC_451/B OR2X1_LOC_636/B OR2X1_LOC_523/B OR2X1_LOC_782/B AND2X1_LOC_52/Y OR2X1_LOC_545/A OR2X1_LOC_676/Y OR2X1_LOC_318/B 
+ OR2X1_LOC_614/Y OR2X1_LOC_259/B OR2X1_LOC_131/A OR2X1_LOC_586/Y AND2X1_LOC_789/Y OR2X1_LOC_348/B OR2X1_LOC_423/Y OR2X1_LOC_7/Y OR2X1_LOC_584/Y OR2X1_LOC_248/A OR2X1_LOC_183/Y OR2X1_LOC_33/B OR2X1_LOC_561/B OR2X1_LOC_127/Y OR2X1_LOC_698/Y OR2X1_LOC_764/Y OR2X1_LOC_380/Y OR2X1_LOC_757/A OR2X1_LOC_125/Y OR2X1_LOC_442/Y OR2X1_LOC_261/Y OR2X1_LOC_106/A AND2X1_LOC_216/A OR2X1_LOC_473/Y OR2X1_LOC_362/A OR2X1_LOC_574/A OR2X1_LOC_810/A AND2X1_LOC_79/Y OR2X1_LOC_719/A OR2X1_LOC_778/A OR2X1_LOC_435/B OR2X1_LOC_646/B OR2X1_LOC_790/A OR2X1_LOC_324/B OR2X1_LOC_148/A AND2X1_LOC_39/Y OR2X1_LOC_499/B OR2X1_LOC_781/A OR2X1_LOC_181/B OR2X1_LOC_210/B OR2X1_LOC_462/B OR2X1_LOC_259/A OR2X1_LOC_518/Y OR2X1_LOC_167/Y OR2X1_LOC_667/Y OR2X1_LOC_250/Y OR2X1_LOC_829/Y OR2X1_LOC_591/Y OR2X1_LOC_321/Y OR2X1_LOC_503/Y OR2X1_LOC_142/Y 
+ OR2X1_LOC_189/Y OR2X1_LOC_759/A OR2X1_LOC_487/Y OR2X1_LOC_406/Y OR2X1_LOC_96/Y OR2X1_LOC_594/Y OR2X1_LOC_533/Y OR2X1_LOC_165/Y OR2X1_LOC_145/Y OR2X1_LOC_680/Y OR2X1_LOC_251/Y OR2X1_LOC_418/Y OR2X1_LOC_52/Y OR2X1_LOC_238/Y OR2X1_LOC_525/Y OR2X1_LOC_163/Y AND2X1_LOC_451/Y AND2X1_LOC_463/B OR2X1_LOC_771/B OR2X1_LOC_639/B OR2X1_LOC_793/A OR2X1_LOC_400/A OR2X1_LOC_209/A OR2X1_LOC_113/B OR2X1_LOC_115/B OR2X1_LOC_342/A OR2X1_LOC_780/A OR2X1_LOC_791/A OR2X1_LOC_403/B OR2X1_LOC_124/B OR2X1_LOC_705/B OR2X1_LOC_347/B OR2X1_LOC_449/A OR2X1_LOC_76/B OR2X1_LOC_559/B OR2X1_LOC_493/B OR2X1_LOC_112/B OR2X1_LOC_302/B OR2X1_LOC_227/B OR2X1_LOC_97/A OR2X1_LOC_467/B OR2X1_LOC_168/A OR2X1_LOC_148/B OR2X1_LOC_728/A OR2X1_LOC_843/B OR2X1_LOC_506/B AND2X1_LOC_450/Y AND2X1_LOC_707/Y OR2X1_LOC_187/Y OR2X1_LOC_166/Y OR2X1_LOC_441/Y 
+ OR2X1_LOC_265/Y OR2X1_LOC_41/Y OR2X1_LOC_745/Y OR2X1_LOC_531/Y OR2X1_LOC_384/Y OR2X1_LOC_171/Y OR2X1_LOC_665/Y OR2X1_LOC_751/Y OR2X1_LOC_767/Y OR2X1_LOC_16/Y OR2X1_LOC_397/Y OR2X1_LOC_177/Y OR2X1_LOC_821/Y OR2X1_LOC_118/Y OR2X1_LOC_674/Y OR2X1_LOC_498/Y OR2X1_LOC_604/Y OR2X1_LOC_438/Y OR2X1_LOC_158/Y OR2X1_LOC_232/Y OR2X1_LOC_258/Y OR2X1_LOC_746/Y OR2X1_LOC_504/Y AND2X1_LOC_197/Y AND2X1_LOC_307/Y AND2X1_LOC_356/B OR2X1_LOC_597/Y AND2X1_LOC_390/B OR2X1_LOC_392/A OR2X1_LOC_549/Y OR2X1_LOC_784/B OR2X1_LOC_633/Y OR2X1_LOC_553/A OR2X1_LOC_640/A OR2X1_LOC_845/A OR2X1_LOC_188/Y OR2X1_LOC_590/Y OR2X1_LOC_460/B OR2X1_LOC_532/Y OR2X1_LOC_243/B OR2X1_LOC_664/Y OR2X1_LOC_151/Y AND2X1_LOC_624/A OR2X1_LOC_79/A OR2X1_LOC_755/A AND2X1_LOC_711/A AND2X1_LOC_706/Y OR2X1_LOC_673/Y AND2X1_LOC_776/Y AND2X1_LOC_168/Y AND2X1_LOC_326/B 
+ AND2X1_LOC_459/Y AND2X1_LOC_638/Y AND2X1_LOC_712/B AND2X1_LOC_727/A AND2X1_LOC_147/Y OR2X1_LOC_630/Y OR2X1_LOC_390/A OR2X1_LOC_506/Y OR2X1_LOC_447/Y OR2X1_LOC_852/B OR2X1_LOC_139/A OR2X1_LOC_199/B OR2X1_LOC_854/A AND2X1_LOC_67/Y OR2X1_LOC_612/Y AND2X1_LOC_848/Y OR2X1_LOC_450/Y OR2X1_LOC_303/A OR2X1_LOC_552/A OR2X1_LOC_303/B AND2X1_LOC_227/Y AND2X1_LOC_714/B AND2X1_LOC_454/A AND2X1_LOC_338/A AND2X1_LOC_489/Y AND2X1_LOC_286/Y OR2X1_LOC_632/A OR2X1_LOC_637/Y OR2X1_LOC_850/A OR2X1_LOC_288/A OR2X1_LOC_609/A AND2X1_LOC_342/Y OR2X1_LOC_669/Y AND2X1_LOC_779/Y AND2X1_LOC_840/B AND2X1_LOC_196/Y AND2X1_LOC_769/Y OR2X1_LOC_829/A AND2X1_LOC_520/Y AND2X1_LOC_464/Y AND2X1_LOC_783/B AND2X1_LOC_841/B OR2X1_LOC_158/B AND2X1_LOC_339/B AND2X1_LOC_715/A AND2X1_LOC_547/Y AND2X1_LOC_729/Y AND2X1_LOC_856/B OR2X1_LOC_656/B AND2X1_LOC_362/B AND2X1_LOC_473/Y 
+ AND2X1_LOC_810/B OR2X1_LOC_472/B OR2X1_LOC_243/A OR2X1_LOC_836/Y OR2X1_LOC_338/A AND2X1_LOC_687/Y OR2X1_LOC_687/Y AND2X1_LOC_456/B OR2X1_LOC_456/A AND2X1_LOC_99/A OR2X1_LOC_802/A OR2X1_LOC_798/Y OR2X1_LOC_99/B AND2X1_LOC_798/Y AND2X1_LOC_802/B OR2X1_LOC_113/Y OR2X1_LOC_539/Y OR2X1_LOC_319/Y AND2X1_LOC_113/Y AND2X1_LOC_798/A AND2X1_LOC_539/Y OR2X1_LOC_593/A OR2X1_LOC_539/B OR2X1_LOC_436/B AND2X1_LOC_434/Y AND2X1_LOC_537/Y AND2X1_LOC_592/Y AND2X1_LOC_593/Y OR2X1_LOC_799/A OR2X1_LOC_216/A OR2X1_LOC_88/Y AND2X1_LOC_374/Y OR2X1_LOC_599/Y OR2X1_LOC_373/Y OR2X1_LOC_644/A AND2X1_LOC_116/Y AND2X1_LOC_88/Y OR2X1_LOC_374/Y OR2X1_LOC_254/B OR2X1_LOC_252/Y OR2X1_LOC_544/B AND2X1_LOC_361/A AND2X1_LOC_483/Y AND2X1_LOC_436/Y OR2X1_LOC_631/B OR2X1_LOC_436/Y OR2X1_LOC_267/Y 

* NETLIST 
XOR2X1_LOC_451 OR2X1_LOC_451/a_8_216# OR2X1_LOC_451/a_36_216# OR2X1_LOC_452/A VSS VDD OR2X1_LOC_451/A OR2X1_LOC_451/B OR2X1_LOC

XAND2X1_LOC_635 AND2X1_LOC_635/a_36_24# AND2X1_LOC_639/A AND2X1_LOC_635/a_8_24# VSS VDD OR2X1_LOC_428/Y OR2X1_LOC_582/Y AND2X1_LOC

XOR2X1_LOC_460 OR2X1_LOC_460/a_8_216# OR2X1_LOC_460/a_36_216# OR2X1_LOC_460/Y VSS VDD OR2X1_LOC_460/A OR2X1_LOC_460/B OR2X1_LOC

XOR2X1_LOC_197 OR2X1_LOC_197/a_8_216# OR2X1_LOC_197/a_36_216# OR2X1_LOC_198/A VSS VDD OR2X1_LOC_197/A AND2X1_LOC_52/Y OR2X1_LOC

XOR2X1_LOC_307 OR2X1_LOC_307/a_8_216# OR2X1_LOC_307/a_36_216# OR2X1_LOC_308/A VSS VDD OR2X1_LOC_307/A OR2X1_LOC_307/B OR2X1_LOC

XOR2X1_LOC_379 OR2X1_LOC_379/a_8_216# OR2X1_LOC_379/a_36_216# OR2X1_LOC_379/Y VSS VDD OR2X1_LOC_66/A AND2X1_LOC_12/Y OR2X1_LOC

XAND2X1_LOC_595 AND2X1_LOC_595/a_36_24# OR2X1_LOC_643/A AND2X1_LOC_595/a_8_24# VSS VDD OR2X1_LOC_66/A OR2X1_LOC_249/Y AND2X1_LOC

XAND2X1_LOC_385 AND2X1_LOC_385/a_36_24# OR2X1_LOC_389/B AND2X1_LOC_385/a_8_24# VSS VDD OR2X1_LOC_66/A OR2X1_LOC_756/B AND2X1_LOC

XAND2X1_LOC_83 AND2X1_LOC_83/a_36_24# OR2X1_LOC_84/A AND2X1_LOC_83/a_8_24# VSS VDD OR2X1_LOC_66/A AND2X1_LOC_82/Y AND2X1_LOC

XAND2X1_LOC_311 AND2X1_LOC_311/a_36_24# OR2X1_LOC_538/A AND2X1_LOC_311/a_8_24# VSS VDD OR2X1_LOC_66/A OR2X1_LOC_532/B AND2X1_LOC

XAND2X1_LOC_176 AND2X1_LOC_176/a_36_24# OR2X1_LOC_180/B AND2X1_LOC_176/a_8_24# VSS VDD OR2X1_LOC_66/A AND2X1_LOC_91/B AND2X1_LOC

XOR2X1_LOC_668 OR2X1_LOC_668/a_8_216# OR2X1_LOC_668/a_36_216# OR2X1_LOC_668/Y VSS VDD OR2X1_LOC_375/A OR2X1_LOC_66/A OR2X1_LOC

XAND2X1_LOC_27 AND2X1_LOC_27/a_36_24# OR2X1_LOC_34/B AND2X1_LOC_27/a_8_24# VSS VDD AND2X1_LOC_7/B OR2X1_LOC_66/A AND2X1_LOC

XAND2X1_LOC_290 AND2X1_LOC_290/a_36_24# OR2X1_LOC_334/B AND2X1_LOC_290/a_8_24# VSS VDD OR2X1_LOC_78/B OR2X1_LOC_66/A AND2X1_LOC

XAND2X1_LOC_677 AND2X1_LOC_677/a_36_24# OR2X1_LOC_834/A AND2X1_LOC_677/a_8_24# VSS VDD OR2X1_LOC_66/A OR2X1_LOC_161/B AND2X1_LOC

XAND2X1_LOC_237 AND2X1_LOC_237/a_36_24# OR2X1_LOC_241/B AND2X1_LOC_237/a_8_24# VSS VDD OR2X1_LOC_66/A OR2X1_LOC_269/B AND2X1_LOC

XAND2X1_LOC_522 AND2X1_LOC_522/a_36_24# OR2X1_LOC_523/A AND2X1_LOC_522/a_8_24# VSS VDD AND2X1_LOC_22/Y OR2X1_LOC_532/B AND2X1_LOC

XAND2X1_LOC_589 AND2X1_LOC_589/a_36_24# OR2X1_LOC_592/A AND2X1_LOC_589/a_8_24# VSS VDD AND2X1_LOC_22/Y OR2X1_LOC_130/A AND2X1_LOC

XAND2X1_LOC_24 AND2X1_LOC_24/a_36_24# OR2X1_LOC_33/A AND2X1_LOC_24/a_8_24# VSS VDD AND2X1_LOC_22/Y OR2X1_LOC_160/B AND2X1_LOC

XAND2X1_LOC_58 AND2X1_LOC_58/a_36_24# OR2X1_LOC_61/B AND2X1_LOC_58/a_8_24# VSS VDD AND2X1_LOC_22/Y OR2X1_LOC_87/A AND2X1_LOC

XAND2X1_LOC_497 AND2X1_LOC_497/a_36_24# OR2X1_LOC_844/B AND2X1_LOC_497/a_8_24# VSS VDD AND2X1_LOC_22/Y AND2X1_LOC_72/B AND2X1_LOC

XAND2X1_LOC_615 AND2X1_LOC_615/a_36_24# OR2X1_LOC_623/B AND2X1_LOC_615/a_8_24# VSS VDD AND2X1_LOC_22/Y OR2X1_LOC_614/Y AND2X1_LOC

XAND2X1_LOC_766 AND2X1_LOC_766/a_36_24# OR2X1_LOC_770/A AND2X1_LOC_766/a_8_24# VSS VDD AND2X1_LOC_64/Y AND2X1_LOC_91/B AND2X1_LOC

XAND2X1_LOC_321 AND2X1_LOC_321/a_36_24# OR2X1_LOC_324/A AND2X1_LOC_321/a_8_24# VSS VDD AND2X1_LOC_41/A AND2X1_LOC_64/Y AND2X1_LOC

XAND2X1_LOC_503 AND2X1_LOC_503/a_36_24# OR2X1_LOC_509/A AND2X1_LOC_503/a_8_24# VSS VDD AND2X1_LOC_64/Y OR2X1_LOC_502/Y AND2X1_LOC

XAND2X1_LOC_312 AND2X1_LOC_312/a_36_24# OR2X1_LOC_703/A AND2X1_LOC_312/a_8_24# VSS VDD AND2X1_LOC_56/B AND2X1_LOC_64/Y AND2X1_LOC

XAND2X1_LOC_142 AND2X1_LOC_142/a_36_24# OR2X1_LOC_147/B AND2X1_LOC_142/a_8_24# VSS VDD OR2X1_LOC_87/A AND2X1_LOC_64/Y AND2X1_LOC

XAND2X1_LOC_314 AND2X1_LOC_314/a_36_24# OR2X1_LOC_317/A AND2X1_LOC_314/a_8_24# VSS VDD OR2X1_LOC_78/B AND2X1_LOC_64/Y AND2X1_LOC

XAND2X1_LOC_65 AND2X1_LOC_65/a_36_24# OR2X1_LOC_201/A AND2X1_LOC_65/a_8_24# VSS VDD AND2X1_LOC_65/A AND2X1_LOC_64/Y AND2X1_LOC

XAND2X1_LOC_518 AND2X1_LOC_518/a_36_24# OR2X1_LOC_520/B AND2X1_LOC_518/a_8_24# VSS VDD AND2X1_LOC_64/Y OR2X1_LOC_185/A AND2X1_LOC

XAND2X1_LOC_167 AND2X1_LOC_167/a_36_24# OR2X1_LOC_703/B AND2X1_LOC_167/a_8_24# VSS VDD AND2X1_LOC_64/Y OR2X1_LOC_161/A AND2X1_LOC

XAND2X1_LOC_822 AND2X1_LOC_822/a_36_24# OR2X1_LOC_835/A AND2X1_LOC_822/a_8_24# VSS VDD AND2X1_LOC_64/Y OR2X1_LOC_532/B AND2X1_LOC

XAND2X1_LOC_107 AND2X1_LOC_107/a_36_24# OR2X1_LOC_113/A AND2X1_LOC_107/a_8_24# VSS VDD AND2X1_LOC_64/Y OR2X1_LOC_78/A AND2X1_LOC

XAND2X1_LOC_698 AND2X1_LOC_698/a_36_24# OR2X1_LOC_709/B AND2X1_LOC_698/a_8_24# VSS VDD AND2X1_LOC_64/Y OR2X1_LOC_160/A AND2X1_LOC

XAND2X1_LOC_667 AND2X1_LOC_667/a_36_24# OR2X1_LOC_720/B AND2X1_LOC_667/a_8_24# VSS VDD AND2X1_LOC_64/Y OR2X1_LOC_264/Y AND2X1_LOC

XAND2X1_LOC_250 AND2X1_LOC_250/a_36_24# OR2X1_LOC_343/B AND2X1_LOC_250/a_8_24# VSS VDD AND2X1_LOC_64/Y OR2X1_LOC_249/Y AND2X1_LOC

XAND2X1_LOC_829 AND2X1_LOC_829/a_36_24# OR2X1_LOC_855/A AND2X1_LOC_829/a_8_24# VSS VDD AND2X1_LOC_64/Y OR2X1_LOC_828/Y AND2X1_LOC

XAND2X1_LOC_423 AND2X1_LOC_423/a_36_24# OR2X1_LOC_449/B AND2X1_LOC_423/a_8_24# VSS VDD AND2X1_LOC_7/B AND2X1_LOC_64/Y AND2X1_LOC

XAND2X1_LOC_253 AND2X1_LOC_253/a_36_24# OR2X1_LOC_254/A AND2X1_LOC_253/a_8_24# VSS VDD AND2X1_LOC_64/Y OR2X1_LOC_161/B AND2X1_LOC

XAND2X1_LOC_591 AND2X1_LOC_591/a_36_24# OR2X1_LOC_593/B AND2X1_LOC_591/a_8_24# VSS VDD AND2X1_LOC_64/Y OR2X1_LOC_590/Y AND2X1_LOC

XAND2X1_LOC_767 AND2X1_LOC_767/a_36_24# OR2X1_LOC_773/B AND2X1_LOC_767/a_8_24# VSS VDD AND2X1_LOC_3/Y OR2X1_LOC_78/Y AND2X1_LOC

XAND2X1_LOC_397 AND2X1_LOC_397/a_36_24# OR2X1_LOC_402/B AND2X1_LOC_397/a_8_24# VSS VDD AND2X1_LOC_3/Y AND2X1_LOC_82/Y AND2X1_LOC

XAND2X1_LOC_305 AND2X1_LOC_305/a_36_24# OR2X1_LOC_307/A AND2X1_LOC_305/a_8_24# VSS VDD AND2X1_LOC_3/Y AND2X1_LOC_91/B AND2X1_LOC

XAND2X1_LOC_127 AND2X1_LOC_127/a_36_24# OR2X1_LOC_128/A AND2X1_LOC_127/a_8_24# VSS VDD AND2X1_LOC_3/Y OR2X1_LOC_160/A AND2X1_LOC

XAND2X1_LOC_16 AND2X1_LOC_16/a_36_24# OR2X1_LOC_194/B AND2X1_LOC_16/a_8_24# VSS VDD AND2X1_LOC_3/Y OR2X1_LOC_78/B AND2X1_LOC

XAND2X1_LOC_481 AND2X1_LOC_481/a_36_24# OR2X1_LOC_555/A AND2X1_LOC_481/a_8_24# VSS VDD AND2X1_LOC_3/Y OR2X1_LOC_294/Y AND2X1_LOC

XAND2X1_LOC_665 AND2X1_LOC_665/a_36_24# OR2X1_LOC_719/B AND2X1_LOC_665/a_8_24# VSS VDD AND2X1_LOC_3/Y OR2X1_LOC_664/Y AND2X1_LOC

XAND2X1_LOC_7 AND2X1_LOC_7/a_36_24# AND2X1_LOC_7/Y AND2X1_LOC_7/a_8_24# VSS VDD AND2X1_LOC_3/Y AND2X1_LOC_7/B AND2X1_LOC

XAND2X1_LOC_281 AND2X1_LOC_281/a_36_24# OR2X1_LOC_285/B AND2X1_LOC_281/a_8_24# VSS VDD AND2X1_LOC_3/Y OR2X1_LOC_269/B AND2X1_LOC

XAND2X1_LOC_815 AND2X1_LOC_815/a_36_24# OR2X1_LOC_846/B AND2X1_LOC_815/a_8_24# VSS VDD AND2X1_LOC_3/Y OR2X1_LOC_814/Y AND2X1_LOC

XAND2X1_LOC_751 AND2X1_LOC_751/a_36_24# OR2X1_LOC_789/A AND2X1_LOC_751/a_8_24# VSS VDD AND2X1_LOC_3/Y OR2X1_LOC_750/Y AND2X1_LOC

XAND2X1_LOC_764 AND2X1_LOC_764/a_36_24# OR2X1_LOC_769/A AND2X1_LOC_764/a_8_24# VSS VDD AND2X1_LOC_40/Y OR2X1_LOC_160/A AND2X1_LOC

XAND2X1_LOC_393 AND2X1_LOC_393/a_36_24# OR2X1_LOC_400/B AND2X1_LOC_393/a_8_24# VSS VDD OR2X1_LOC_154/A AND2X1_LOC_40/Y AND2X1_LOC

XAND2X1_LOC_745 AND2X1_LOC_745/a_36_24# OR2X1_LOC_781/B AND2X1_LOC_745/a_8_24# VSS VDD AND2X1_LOC_40/Y OR2X1_LOC_161/A AND2X1_LOC

XAND2X1_LOC_531 AND2X1_LOC_531/a_36_24# OR2X1_LOC_549/B AND2X1_LOC_531/a_8_24# VSS VDD AND2X1_LOC_40/Y OR2X1_LOC_185/A AND2X1_LOC

XAND2X1_LOC_384 AND2X1_LOC_384/a_36_24# OR2X1_LOC_391/A AND2X1_LOC_384/a_8_24# VSS VDD AND2X1_LOC_40/Y OR2X1_LOC_383/Y AND2X1_LOC

XAND2X1_LOC_171 AND2X1_LOC_171/a_36_24# OR2X1_LOC_333/B AND2X1_LOC_171/a_8_24# VSS VDD OR2X1_LOC_160/B AND2X1_LOC_40/Y AND2X1_LOC

XAND2X1_LOC_183 AND2X1_LOC_183/a_36_24# OR2X1_LOC_190/B AND2X1_LOC_183/a_8_24# VSS VDD AND2X1_LOC_7/B AND2X1_LOC_40/Y AND2X1_LOC

XAND2X1_LOC_41 AND2X1_LOC_41/a_36_24# AND2X1_LOC_41/Y AND2X1_LOC_41/a_8_24# VSS VDD AND2X1_LOC_41/A AND2X1_LOC_40/Y AND2X1_LOC

XOR2X1_LOC_610 OR2X1_LOC_610/a_8_216# OR2X1_LOC_610/a_36_216# OR2X1_LOC_610/Y VSS VDD AND2X1_LOC_47/Y AND2X1_LOC_40/Y OR2X1_LOC

XAND2X1_LOC_187 AND2X1_LOC_187/a_36_24# OR2X1_LOC_191/B AND2X1_LOC_187/a_8_24# VSS VDD AND2X1_LOC_40/Y OR2X1_LOC_186/Y AND2X1_LOC

XAND2X1_LOC_166 AND2X1_LOC_166/a_36_24# OR2X1_LOC_169/B AND2X1_LOC_166/a_8_24# VSS VDD OR2X1_LOC_78/B AND2X1_LOC_40/Y AND2X1_LOC

XAND2X1_LOC_670 AND2X1_LOC_670/a_36_24# OR2X1_LOC_673/B AND2X1_LOC_670/a_8_24# VSS VDD AND2X1_LOC_40/Y OR2X1_LOC_532/B AND2X1_LOC

XAND2X1_LOC_292 AND2X1_LOC_292/a_36_24# OR2X1_LOC_346/B AND2X1_LOC_292/a_8_24# VSS VDD AND2X1_LOC_40/Y OR2X1_LOC_151/A AND2X1_LOC

XAND2X1_LOC_441 AND2X1_LOC_441/a_36_24# OR2X1_LOC_545/B AND2X1_LOC_441/a_8_24# VSS VDD AND2X1_LOC_40/Y OR2X1_LOC_87/A AND2X1_LOC

XAND2X1_LOC_442 AND2X1_LOC_442/a_36_24# OR2X1_LOC_444/B AND2X1_LOC_442/a_8_24# VSS VDD AND2X1_LOC_40/Y OR2X1_LOC_756/B AND2X1_LOC

XAND2X1_LOC_613 AND2X1_LOC_613/a_36_24# OR2X1_LOC_620/A AND2X1_LOC_613/a_8_24# VSS VDD AND2X1_LOC_40/Y AND2X1_LOC_56/B AND2X1_LOC

XAND2X1_LOC_262 AND2X1_LOC_262/a_36_24# OR2X1_LOC_786/A AND2X1_LOC_262/a_8_24# VSS VDD AND2X1_LOC_40/Y AND2X1_LOC_65/A AND2X1_LOC

XAND2X1_LOC_265 AND2X1_LOC_265/a_36_24# OR2X1_LOC_641/A AND2X1_LOC_265/a_8_24# VSS VDD AND2X1_LOC_40/Y OR2X1_LOC_264/Y AND2X1_LOC

XOR2X1_LOC_758 OR2X1_LOC_758/a_8_216# OR2X1_LOC_758/a_36_216# OR2X1_LOC_758/Y VSS VDD AND2X1_LOC_95/Y AND2X1_LOC_40/Y OR2X1_LOC

XAND2X1_LOC_586 AND2X1_LOC_586/a_36_24# OR2X1_LOC_637/A AND2X1_LOC_586/a_8_24# VSS VDD AND2X1_LOC_70/Y OR2X1_LOC_130/A AND2X1_LOC

XAND2X1_LOC_172 AND2X1_LOC_172/a_36_24# OR2X1_LOC_174/A AND2X1_LOC_172/a_8_24# VSS VDD AND2X1_LOC_70/Y OR2X1_LOC_532/B AND2X1_LOC

XAND2X1_LOC_72 AND2X1_LOC_72/a_36_24# AND2X1_LOC_72/Y AND2X1_LOC_72/a_8_24# VSS VDD AND2X1_LOC_70/Y AND2X1_LOC_72/B AND2X1_LOC

XAND2X1_LOC_173 AND2X1_LOC_173/a_36_24# OR2X1_LOC_175/B AND2X1_LOC_173/a_8_24# VSS VDD AND2X1_LOC_70/Y OR2X1_LOC_151/A AND2X1_LOC

XAND2X1_LOC_313 AND2X1_LOC_313/a_36_24# OR2X1_LOC_317/B AND2X1_LOC_313/a_8_24# VSS VDD AND2X1_LOC_70/Y AND2X1_LOC_91/B AND2X1_LOC

XAND2X1_LOC_177 AND2X1_LOC_177/a_36_24# OR2X1_LOC_439/B AND2X1_LOC_177/a_8_24# VSS VDD OR2X1_LOC_87/A AND2X1_LOC_70/Y AND2X1_LOC

XAND2X1_LOC_821 AND2X1_LOC_821/a_36_24# OR2X1_LOC_835/B AND2X1_LOC_821/a_8_24# VSS VDD AND2X1_LOC_41/A AND2X1_LOC_70/Y AND2X1_LOC

XAND2X1_LOC_117 AND2X1_LOC_117/a_36_24# OR2X1_LOC_123/B AND2X1_LOC_117/a_8_24# VSS VDD AND2X1_LOC_65/A AND2X1_LOC_70/Y AND2X1_LOC

XAND2X1_LOC_118 AND2X1_LOC_118/a_36_24# OR2X1_LOC_633/B AND2X1_LOC_118/a_8_24# VSS VDD AND2X1_LOC_70/Y OR2X1_LOC_78/A AND2X1_LOC

XAND2X1_LOC_674 AND2X1_LOC_674/a_36_24# OR2X1_LOC_675/A AND2X1_LOC_674/a_8_24# VSS VDD AND2X1_LOC_70/Y OR2X1_LOC_405/A AND2X1_LOC

XAND2X1_LOC_431 AND2X1_LOC_431/a_36_24# OR2X1_LOC_434/A AND2X1_LOC_431/a_8_24# VSS VDD AND2X1_LOC_70/Y OR2X1_LOC_269/B AND2X1_LOC

XAND2X1_LOC_498 AND2X1_LOC_498/a_36_24# OR2X1_LOC_501/B AND2X1_LOC_498/a_8_24# VSS VDD AND2X1_LOC_70/Y OR2X1_LOC_188/Y AND2X1_LOC

XAND2X1_LOC_604 AND2X1_LOC_604/a_36_24# OR2X1_LOC_605/A AND2X1_LOC_604/a_8_24# VSS VDD AND2X1_LOC_70/Y OR2X1_LOC_161/A AND2X1_LOC

XAND2X1_LOC_438 AND2X1_LOC_438/a_36_24# OR2X1_LOC_544/A AND2X1_LOC_438/a_8_24# VSS VDD OR2X1_LOC_160/B AND2X1_LOC_70/Y AND2X1_LOC

XAND2X1_LOC_427 AND2X1_LOC_427/a_36_24# OR2X1_LOC_450/A AND2X1_LOC_427/a_8_24# VSS VDD AND2X1_LOC_70/Y OR2X1_LOC_161/B AND2X1_LOC

XOR2X1_LOC_330 OR2X1_LOC_330/a_8_216# OR2X1_LOC_330/a_36_216# OR2X1_LOC_330/Y VSS VDD AND2X1_LOC_70/Y AND2X1_LOC_51/Y OR2X1_LOC

XOR2X1_LOC_103 OR2X1_LOC_103/a_8_216# OR2X1_LOC_103/a_36_216# OR2X1_LOC_103/Y VSS VDD OR2X1_LOC_485/A OR2X1_LOC_47/Y OR2X1_LOC

XOR2X1_LOC_106 OR2X1_LOC_106/a_8_216# OR2X1_LOC_106/a_36_216# OR2X1_LOC_106/Y VSS VDD OR2X1_LOC_106/A OR2X1_LOC_47/Y OR2X1_LOC

XOR2X1_LOC_695 OR2X1_LOC_695/a_8_216# OR2X1_LOC_695/a_36_216# OR2X1_LOC_695/Y VSS VDD OR2X1_LOC_47/Y OR2X1_LOC_45/B OR2X1_LOC

XOR2X1_LOC_280 OR2X1_LOC_280/a_8_216# OR2X1_LOC_280/a_36_216# OR2X1_LOC_280/Y VSS VDD OR2X1_LOC_428/A OR2X1_LOC_47/Y OR2X1_LOC

XOR2X1_LOC_601 OR2X1_LOC_601/a_8_216# OR2X1_LOC_601/a_36_216# OR2X1_LOC_601/Y VSS VDD OR2X1_LOC_47/Y OR2X1_LOC_16/A OR2X1_LOC

XAND2X1_LOC_610 AND2X1_LOC_610/a_36_24# OR2X1_LOC_612/B AND2X1_LOC_610/a_8_24# VSS VDD OR2X1_LOC_40/Y OR2X1_LOC_47/Y AND2X1_LOC

XOR2X1_LOC_248 OR2X1_LOC_248/a_8_216# OR2X1_LOC_248/a_36_216# OR2X1_LOC_248/Y VSS VDD OR2X1_LOC_248/A OR2X1_LOC_47/Y OR2X1_LOC

XOR2X1_LOC_394 OR2X1_LOC_394/a_8_216# OR2X1_LOC_394/a_36_216# OR2X1_LOC_394/Y VSS VDD OR2X1_LOC_744/A OR2X1_LOC_47/Y OR2X1_LOC

XOR2X1_LOC_747 OR2X1_LOC_747/a_8_216# OR2X1_LOC_747/a_36_216# OR2X1_LOC_747/Y VSS VDD OR2X1_LOC_52/B OR2X1_LOC_47/Y OR2X1_LOC

XOR2X1_LOC_524 OR2X1_LOC_524/a_8_216# OR2X1_LOC_524/a_36_216# OR2X1_LOC_524/Y VSS VDD OR2X1_LOC_427/A OR2X1_LOC_47/Y OR2X1_LOC

XOR2X1_LOC_152 OR2X1_LOC_152/a_8_216# OR2X1_LOC_152/a_36_216# OR2X1_LOC_152/Y VSS VDD OR2X1_LOC_152/A OR2X1_LOC_47/Y OR2X1_LOC

XOR2X1_LOC_528 OR2X1_LOC_528/a_8_216# OR2X1_LOC_528/a_36_216# OR2X1_LOC_528/Y VSS VDD OR2X1_LOC_44/Y OR2X1_LOC_7/A OR2X1_LOC

XOR2X1_LOC_122 OR2X1_LOC_122/a_8_216# OR2X1_LOC_122/a_36_216# OR2X1_LOC_122/Y VSS VDD OR2X1_LOC_122/A OR2X1_LOC_44/Y OR2X1_LOC

XOR2X1_LOC_825 OR2X1_LOC_825/a_8_216# OR2X1_LOC_825/a_36_216# OR2X1_LOC_825/Y VSS VDD OR2X1_LOC_96/B OR2X1_LOC_44/Y OR2X1_LOC

XOR2X1_LOC_485 OR2X1_LOC_485/a_8_216# OR2X1_LOC_485/a_36_216# OR2X1_LOC_485/Y VSS VDD OR2X1_LOC_485/A OR2X1_LOC_44/Y OR2X1_LOC

XOR2X1_LOC_297 OR2X1_LOC_297/a_8_216# OR2X1_LOC_297/a_36_216# OR2X1_LOC_297/Y VSS VDD OR2X1_LOC_297/A OR2X1_LOC_44/Y OR2X1_LOC

XOR2X1_LOC_424 OR2X1_LOC_424/a_8_216# OR2X1_LOC_424/a_36_216# OR2X1_LOC_424/Y VSS VDD OR2X1_LOC_89/A OR2X1_LOC_44/Y OR2X1_LOC

XOR2X1_LOC_279 OR2X1_LOC_279/a_8_216# OR2X1_LOC_279/a_36_216# OR2X1_LOC_279/Y VSS VDD OR2X1_LOC_427/A OR2X1_LOC_44/Y OR2X1_LOC

XOR2X1_LOC_45 OR2X1_LOC_45/a_8_216# OR2X1_LOC_45/a_36_216# OR2X1_LOC_45/Y VSS VDD OR2X1_LOC_44/Y OR2X1_LOC_45/B OR2X1_LOC

XOR2X1_LOC_744 OR2X1_LOC_744/a_8_216# OR2X1_LOC_744/a_36_216# OR2X1_LOC_744/Y VSS VDD OR2X1_LOC_744/A OR2X1_LOC_44/Y OR2X1_LOC

XOR2X1_LOC_701 OR2X1_LOC_701/a_8_216# OR2X1_LOC_701/a_36_216# OR2X1_LOC_701/Y VSS VDD OR2X1_LOC_428/A OR2X1_LOC_44/Y OR2X1_LOC

XOR2X1_LOC_757 OR2X1_LOC_757/a_8_216# OR2X1_LOC_757/a_36_216# OR2X1_LOC_757/Y VSS VDD OR2X1_LOC_757/A OR2X1_LOC_44/Y OR2X1_LOC

XOR2X1_LOC_399 OR2X1_LOC_399/a_8_216# OR2X1_LOC_399/a_36_216# OR2X1_LOC_399/Y VSS VDD OR2X1_LOC_399/A OR2X1_LOC_44/Y OR2X1_LOC

XOR2X1_LOC_517 OR2X1_LOC_517/a_8_216# OR2X1_LOC_517/a_36_216# OR2X1_LOC_517/Y VSS VDD OR2X1_LOC_517/A OR2X1_LOC_31/Y OR2X1_LOC

XOR2X1_LOC_315 OR2X1_LOC_315/a_8_216# OR2X1_LOC_315/a_36_216# OR2X1_LOC_315/Y VSS VDD OR2X1_LOC_427/A OR2X1_LOC_31/Y OR2X1_LOC

XOR2X1_LOC_491 OR2X1_LOC_491/a_8_216# OR2X1_LOC_491/a_36_216# OR2X1_LOC_491/Y VSS VDD OR2X1_LOC_485/A OR2X1_LOC_31/Y OR2X1_LOC

XOR2X1_LOC_109 OR2X1_LOC_109/a_8_216# OR2X1_LOC_109/a_36_216# OR2X1_LOC_109/Y VSS VDD OR2X1_LOC_89/A OR2X1_LOC_31/Y OR2X1_LOC

XOR2X1_LOC_600 OR2X1_LOC_600/a_8_216# OR2X1_LOC_600/a_36_216# OR2X1_LOC_600/Y VSS VDD OR2X1_LOC_600/A OR2X1_LOC_31/Y OR2X1_LOC

XOR2X1_LOC_230 OR2X1_LOC_230/a_8_216# OR2X1_LOC_230/a_36_216# OR2X1_LOC_230/Y VSS VDD OR2X1_LOC_31/Y OR2X1_LOC_7/A OR2X1_LOC

XOR2X1_LOC_298 OR2X1_LOC_298/a_8_216# OR2X1_LOC_298/a_36_216# OR2X1_LOC_298/Y VSS VDD OR2X1_LOC_56/A OR2X1_LOC_31/Y OR2X1_LOC

XOR2X1_LOC_224 OR2X1_LOC_224/a_8_216# OR2X1_LOC_224/a_36_216# OR2X1_LOC_224/Y VSS VDD OR2X1_LOC_744/A OR2X1_LOC_31/Y OR2X1_LOC

XOR2X1_LOC_428 OR2X1_LOC_428/a_8_216# OR2X1_LOC_428/a_36_216# OR2X1_LOC_428/Y VSS VDD OR2X1_LOC_428/A OR2X1_LOC_31/Y OR2X1_LOC

XOR2X1_LOC_74 OR2X1_LOC_74/a_8_216# OR2X1_LOC_74/a_36_216# OR2X1_LOC_74/Y VSS VDD OR2X1_LOC_74/A OR2X1_LOC_31/Y OR2X1_LOC

XOR2X1_LOC_32 OR2X1_LOC_32/a_8_216# OR2X1_LOC_32/a_36_216# OR2X1_LOC_32/Y VSS VDD OR2X1_LOC_31/Y OR2X1_LOC_32/B OR2X1_LOC

XOR2X1_LOC_583 OR2X1_LOC_583/a_8_216# OR2X1_LOC_583/a_36_216# OR2X1_LOC_583/Y VSS VDD OR2X1_LOC_52/B OR2X1_LOC_31/Y OR2X1_LOC

XOR2X1_LOC_526 OR2X1_LOC_526/a_8_216# OR2X1_LOC_526/a_36_216# OR2X1_LOC_526/Y VSS VDD OR2X1_LOC_604/A OR2X1_LOC_31/Y OR2X1_LOC

XOR2X1_LOC_505 OR2X1_LOC_505/a_8_216# OR2X1_LOC_505/a_36_216# OR2X1_LOC_505/Y VSS VDD OR2X1_LOC_45/B OR2X1_LOC_18/Y OR2X1_LOC

XOR2X1_LOC_666 OR2X1_LOC_666/a_8_216# OR2X1_LOC_666/a_36_216# OR2X1_LOC_666/Y VSS VDD OR2X1_LOC_666/A OR2X1_LOC_18/Y OR2X1_LOC

XOR2X1_LOC_496 OR2X1_LOC_496/a_8_216# OR2X1_LOC_496/a_36_216# OR2X1_LOC_496/Y VSS VDD OR2X1_LOC_56/A OR2X1_LOC_18/Y OR2X1_LOC

XOR2X1_LOC_432 OR2X1_LOC_432/a_8_216# OR2X1_LOC_432/a_36_216# OR2X1_LOC_432/Y VSS VDD OR2X1_LOC_589/A OR2X1_LOC_18/Y OR2X1_LOC

XOR2X1_LOC_616 OR2X1_LOC_616/a_8_216# OR2X1_LOC_616/a_36_216# OR2X1_LOC_616/Y VSS VDD OR2X1_LOC_600/A OR2X1_LOC_18/Y OR2X1_LOC

XOR2X1_LOC_607 OR2X1_LOC_607/a_8_216# OR2X1_LOC_607/a_36_216# OR2X1_LOC_607/Y VSS VDD OR2X1_LOC_607/A OR2X1_LOC_18/Y OR2X1_LOC

XOR2X1_LOC_257 OR2X1_LOC_257/a_8_216# OR2X1_LOC_257/a_36_216# OR2X1_LOC_257/Y VSS VDD OR2X1_LOC_427/A OR2X1_LOC_18/Y OR2X1_LOC

XOR2X1_LOC_20 OR2X1_LOC_20/a_8_216# OR2X1_LOC_20/a_36_216# OR2X1_LOC_20/Y VSS VDD OR2X1_LOC_20/A OR2X1_LOC_18/Y OR2X1_LOC

XOR2X1_LOC_79 OR2X1_LOC_79/a_8_216# OR2X1_LOC_79/a_36_216# OR2X1_LOC_79/Y VSS VDD OR2X1_LOC_79/A OR2X1_LOC_18/Y OR2X1_LOC

XOR2X1_LOC_521 OR2X1_LOC_521/a_8_216# OR2X1_LOC_521/a_36_216# OR2X1_LOC_521/Y VSS VDD OR2X1_LOC_52/B OR2X1_LOC_18/Y OR2X1_LOC

XOR2X1_LOC_135 OR2X1_LOC_135/a_8_216# OR2X1_LOC_135/a_36_216# OR2X1_LOC_135/Y VSS VDD OR2X1_LOC_427/A OR2X1_LOC_59/Y OR2X1_LOC

XOR2X1_LOC_492 OR2X1_LOC_492/a_8_216# OR2X1_LOC_492/a_36_216# OR2X1_LOC_492/Y VSS VDD OR2X1_LOC_744/A OR2X1_LOC_59/Y OR2X1_LOC

XOR2X1_LOC_482 OR2X1_LOC_482/a_8_216# OR2X1_LOC_482/a_36_216# OR2X1_LOC_482/Y VSS VDD OR2X1_LOC_59/Y OR2X1_LOC_7/A OR2X1_LOC

XOR2X1_LOC_108 OR2X1_LOC_108/a_8_216# OR2X1_LOC_108/a_36_216# OR2X1_LOC_108/Y VSS VDD OR2X1_LOC_485/A OR2X1_LOC_59/Y OR2X1_LOC

XOR2X1_LOC_295 OR2X1_LOC_295/a_8_216# OR2X1_LOC_295/a_36_216# OR2X1_LOC_295/Y VSS VDD OR2X1_LOC_481/A OR2X1_LOC_59/Y OR2X1_LOC

XOR2X1_LOC_252 OR2X1_LOC_252/a_8_216# OR2X1_LOC_252/a_36_216# OR2X1_LOC_252/Y VSS VDD OR2X1_LOC_59/Y OR2X1_LOC_56/A OR2X1_LOC

XOR2X1_LOC_81 OR2X1_LOC_81/a_8_216# OR2X1_LOC_81/a_36_216# OR2X1_LOC_81/Y VSS VDD OR2X1_LOC_80/Y OR2X1_LOC_59/Y OR2X1_LOC

XOR2X1_LOC_60 OR2X1_LOC_60/a_8_216# OR2X1_LOC_60/a_36_216# OR2X1_LOC_60/Y VSS VDD OR2X1_LOC_59/Y OR2X1_LOC_39/A OR2X1_LOC

XOR2X1_LOC_437 OR2X1_LOC_437/a_8_216# OR2X1_LOC_437/a_36_216# OR2X1_LOC_437/Y VSS VDD OR2X1_LOC_437/A OR2X1_LOC_59/Y OR2X1_LOC

XOR2X1_LOC_609 OR2X1_LOC_609/a_8_216# OR2X1_LOC_609/a_36_216# OR2X1_LOC_609/Y VSS VDD OR2X1_LOC_609/A OR2X1_LOC_59/Y OR2X1_LOC

XOR2X1_LOC_75 OR2X1_LOC_75/a_8_216# OR2X1_LOC_75/a_36_216# OR2X1_LOC_75/Y VSS VDD OR2X1_LOC_59/Y OR2X1_LOC_45/B OR2X1_LOC

XOR2X1_LOC_89 OR2X1_LOC_89/a_8_216# OR2X1_LOC_89/a_36_216# OR2X1_LOC_89/Y VSS VDD OR2X1_LOC_89/A OR2X1_LOC_59/Y OR2X1_LOC

XOR2X1_LOC_700 OR2X1_LOC_700/a_8_216# OR2X1_LOC_700/a_36_216# OR2X1_LOC_700/Y VSS VDD OR2X1_LOC_91/A OR2X1_LOC_59/Y OR2X1_LOC

XOR2X1_LOC_755 OR2X1_LOC_755/a_8_216# OR2X1_LOC_755/a_36_216# OR2X1_LOC_755/Y VSS VDD OR2X1_LOC_755/A OR2X1_LOC_59/Y OR2X1_LOC

XOR2X1_LOC_395 OR2X1_LOC_395/a_8_216# OR2X1_LOC_395/a_36_216# OR2X1_LOC_395/Y VSS VDD OR2X1_LOC_600/A OR2X1_LOC_59/Y OR2X1_LOC

XOR2X1_LOC_316 OR2X1_LOC_316/a_8_216# OR2X1_LOC_316/a_36_216# OR2X1_LOC_316/Y VSS VDD OR2X1_LOC_80/Y OR2X1_LOC_12/Y OR2X1_LOC

XOR2X1_LOC_494 OR2X1_LOC_494/a_8_216# OR2X1_LOC_494/a_36_216# OR2X1_LOC_494/Y VSS VDD OR2X1_LOC_494/A OR2X1_LOC_12/Y OR2X1_LOC

XAND2X1_LOC_379 AND2X1_LOC_379/a_36_24# OR2X1_LOC_380/A AND2X1_LOC_379/a_8_24# VSS VDD OR2X1_LOC_12/Y OR2X1_LOC_26/Y AND2X1_LOC

XOR2X1_LOC_603 OR2X1_LOC_603/a_8_216# OR2X1_LOC_603/a_36_216# OR2X1_LOC_603/Y VSS VDD OR2X1_LOC_52/B OR2X1_LOC_12/Y OR2X1_LOC

XAND2X1_LOC_260 AND2X1_LOC_260/a_36_24# OR2X1_LOC_261/A AND2X1_LOC_260/a_8_24# VSS VDD OR2X1_LOC_12/Y OR2X1_LOC_158/A AND2X1_LOC

XAND2X1_LOC_678 AND2X1_LOC_678/a_36_24# OR2X1_LOC_679/A AND2X1_LOC_678/a_8_24# VSS VDD OR2X1_LOC_12/Y OR2X1_LOC_677/Y AND2X1_LOC

XOR2X1_LOC_229 OR2X1_LOC_229/a_8_216# OR2X1_LOC_229/a_36_216# OR2X1_LOC_229/Y VSS VDD OR2X1_LOC_45/B OR2X1_LOC_12/Y OR2X1_LOC

XOR2X1_LOC_13 OR2X1_LOC_13/a_8_216# OR2X1_LOC_13/a_36_216# OR2X1_LOC_13/Y VSS VDD OR2X1_LOC_12/Y OR2X1_LOC_13/B OR2X1_LOC

XOR2X1_LOC_765 OR2X1_LOC_765/a_8_216# OR2X1_LOC_765/a_36_216# OR2X1_LOC_765/Y VSS VDD OR2X1_LOC_16/A OR2X1_LOC_12/Y OR2X1_LOC

XOR2X1_LOC_536 OR2X1_LOC_536/a_8_216# OR2X1_LOC_536/a_36_216# OR2X1_LOC_536/Y VSS VDD OR2X1_LOC_485/A OR2X1_LOC_12/Y OR2X1_LOC

XOR2X1_LOC_131 OR2X1_LOC_131/a_8_216# OR2X1_LOC_131/a_36_216# OR2X1_LOC_131/Y VSS VDD OR2X1_LOC_131/A OR2X1_LOC_12/Y OR2X1_LOC

XAND2X1_LOC_790 AND2X1_LOC_790/a_36_24# AND2X1_LOC_793/B AND2X1_LOC_790/a_8_24# VSS VDD OR2X1_LOC_753/Y OR2X1_LOC_754/Y AND2X1_LOC

XOR2X1_LOC_707 OR2X1_LOC_707/a_8_216# OR2X1_LOC_707/a_36_216# OR2X1_LOC_712/B VSS VDD OR2X1_LOC_707/A OR2X1_LOC_707/B OR2X1_LOC

XAND2X1_LOC_755 AND2X1_LOC_755/a_36_24# OR2X1_LOC_791/B AND2X1_LOC_755/a_8_24# VSS VDD AND2X1_LOC_59/Y OR2X1_LOC_664/Y AND2X1_LOC

XAND2X1_LOC_700 AND2X1_LOC_700/a_36_24# OR2X1_LOC_710/B AND2X1_LOC_700/a_8_24# VSS VDD AND2X1_LOC_59/Y AND2X1_LOC_91/B AND2X1_LOC

XAND2X1_LOC_395 AND2X1_LOC_395/a_36_24# OR2X1_LOC_401/B AND2X1_LOC_395/a_8_24# VSS VDD AND2X1_LOC_59/Y OR2X1_LOC_756/B AND2X1_LOC

XAND2X1_LOC_81 AND2X1_LOC_81/a_36_24# OR2X1_LOC_84/B AND2X1_LOC_81/a_8_24# VSS VDD AND2X1_LOC_59/Y AND2X1_LOC_81/B AND2X1_LOC

XAND2X1_LOC_60 AND2X1_LOC_60/a_36_24# OR2X1_LOC_61/A AND2X1_LOC_60/a_8_24# VSS VDD OR2X1_LOC_154/A AND2X1_LOC_59/Y AND2X1_LOC

XAND2X1_LOC_75 AND2X1_LOC_75/a_36_24# OR2X1_LOC_76/A AND2X1_LOC_75/a_8_24# VSS VDD OR2X1_LOC_160/B AND2X1_LOC_59/Y AND2X1_LOC

XAND2X1_LOC_89 AND2X1_LOC_89/a_36_24# OR2X1_LOC_97/B AND2X1_LOC_89/a_8_24# VSS VDD AND2X1_LOC_59/Y OR2X1_LOC_78/A AND2X1_LOC

XAND2X1_LOC_135 AND2X1_LOC_135/a_36_24# OR2X1_LOC_702/A AND2X1_LOC_135/a_8_24# VSS VDD AND2X1_LOC_59/Y OR2X1_LOC_161/B AND2X1_LOC

XAND2X1_LOC_492 AND2X1_LOC_492/a_36_24# OR2X1_LOC_493/A AND2X1_LOC_492/a_8_24# VSS VDD AND2X1_LOC_59/Y OR2X1_LOC_160/A AND2X1_LOC

XAND2X1_LOC_482 AND2X1_LOC_482/a_36_24# OR2X1_LOC_833/B AND2X1_LOC_482/a_8_24# VSS VDD AND2X1_LOC_7/B AND2X1_LOC_59/Y AND2X1_LOC

XAND2X1_LOC_108 AND2X1_LOC_108/a_36_24# OR2X1_LOC_114/B AND2X1_LOC_108/a_8_24# VSS VDD AND2X1_LOC_59/Y OR2X1_LOC_532/B AND2X1_LOC

XAND2X1_LOC_295 AND2X1_LOC_295/a_36_24# OR2X1_LOC_346/A AND2X1_LOC_295/a_8_24# VSS VDD AND2X1_LOC_59/Y OR2X1_LOC_294/Y AND2X1_LOC

XAND2X1_LOC_252 AND2X1_LOC_252/a_36_24# OR2X1_LOC_254/B AND2X1_LOC_252/a_8_24# VSS VDD AND2X1_LOC_56/B AND2X1_LOC_59/Y AND2X1_LOC

XAND2X1_LOC_437 AND2X1_LOC_437/a_36_24# OR2X1_LOC_440/B AND2X1_LOC_437/a_8_24# VSS VDD AND2X1_LOC_59/Y OR2X1_LOC_151/A AND2X1_LOC

XAND2X1_LOC_609 AND2X1_LOC_609/a_36_24# OR2X1_LOC_646/A AND2X1_LOC_609/a_8_24# VSS VDD AND2X1_LOC_59/Y OR2X1_LOC_608/Y AND2X1_LOC

XAND2X1_LOC_229 AND2X1_LOC_229/a_36_24# OR2X1_LOC_231/B AND2X1_LOC_229/a_8_24# VSS VDD AND2X1_LOC_12/Y OR2X1_LOC_160/B AND2X1_LOC

XAND2X1_LOC_765 AND2X1_LOC_765/a_36_24# OR2X1_LOC_770/B AND2X1_LOC_765/a_8_24# VSS VDD AND2X1_LOC_12/Y OR2X1_LOC_78/B AND2X1_LOC

XAND2X1_LOC_536 AND2X1_LOC_536/a_36_24# OR2X1_LOC_537/A AND2X1_LOC_536/a_8_24# VSS VDD AND2X1_LOC_12/Y OR2X1_LOC_532/B AND2X1_LOC

XAND2X1_LOC_131 AND2X1_LOC_131/a_36_24# OR2X1_LOC_140/A AND2X1_LOC_131/a_8_24# VSS VDD AND2X1_LOC_12/Y OR2X1_LOC_130/Y AND2X1_LOC

XOR2X1_LOC_260 OR2X1_LOC_260/a_8_216# OR2X1_LOC_260/a_36_216# OR2X1_LOC_260/Y VSS VDD OR2X1_LOC_375/A AND2X1_LOC_12/Y OR2X1_LOC

XOR2X1_LOC_678 OR2X1_LOC_678/a_8_216# OR2X1_LOC_678/a_36_216# OR2X1_LOC_678/Y VSS VDD OR2X1_LOC_834/A AND2X1_LOC_12/Y OR2X1_LOC

XAND2X1_LOC_316 AND2X1_LOC_316/a_36_24# OR2X1_LOC_318/A AND2X1_LOC_316/a_8_24# VSS VDD AND2X1_LOC_12/Y AND2X1_LOC_81/B AND2X1_LOC

XAND2X1_LOC_13 AND2X1_LOC_13/a_36_24# OR2X1_LOC_193/A AND2X1_LOC_13/a_8_24# VSS VDD AND2X1_LOC_41/A AND2X1_LOC_12/Y AND2X1_LOC

XAND2X1_LOC_494 AND2X1_LOC_494/a_36_24# OR2X1_LOC_558/A AND2X1_LOC_494/a_8_24# VSS VDD AND2X1_LOC_12/Y OR2X1_LOC_383/Y AND2X1_LOC

XAND2X1_LOC_603 AND2X1_LOC_603/a_36_24# OR2X1_LOC_605/B AND2X1_LOC_603/a_8_24# VSS VDD AND2X1_LOC_12/Y OR2X1_LOC_87/A AND2X1_LOC

XAND2X1_LOC_594 AND2X1_LOC_594/a_36_24# OR2X1_LOC_653/B AND2X1_LOC_594/a_8_24# VSS VDD AND2X1_LOC_95/Y OR2X1_LOC_186/Y AND2X1_LOC

XAND2X1_LOC_533 AND2X1_LOC_533/a_36_24# OR2X1_LOC_788/B AND2X1_LOC_533/a_8_24# VSS VDD AND2X1_LOC_95/Y OR2X1_LOC_532/Y AND2X1_LOC

XAND2X1_LOC_184 AND2X1_LOC_184/a_36_24# OR2X1_LOC_190/A AND2X1_LOC_184/a_8_24# VSS VDD AND2X1_LOC_72/B AND2X1_LOC_95/Y AND2X1_LOC

XAND2X1_LOC_96 AND2X1_LOC_96/a_36_24# OR2X1_LOC_98/A AND2X1_LOC_96/a_8_24# VSS VDD AND2X1_LOC_94/Y AND2X1_LOC_95/Y AND2X1_LOC

XAND2X1_LOC_132 AND2X1_LOC_132/a_36_24# OR2X1_LOC_137/B AND2X1_LOC_132/a_8_24# VSS VDD AND2X1_LOC_91/B AND2X1_LOC_95/Y AND2X1_LOC

XAND2X1_LOC_189 AND2X1_LOC_189/a_36_24# OR2X1_LOC_192/B AND2X1_LOC_189/a_8_24# VSS VDD AND2X1_LOC_95/Y OR2X1_LOC_188/Y AND2X1_LOC

XAND2X1_LOC_134 AND2X1_LOC_134/a_36_24# OR2X1_LOC_768/A AND2X1_LOC_134/a_8_24# VSS VDD AND2X1_LOC_95/Y OR2X1_LOC_161/B AND2X1_LOC

XAND2X1_LOC_125 AND2X1_LOC_125/a_36_24# OR2X1_LOC_128/B AND2X1_LOC_125/a_8_24# VSS VDD AND2X1_LOC_95/Y OR2X1_LOC_756/B AND2X1_LOC

XAND2X1_LOC_826 AND2X1_LOC_826/a_36_24# OR2X1_LOC_837/A AND2X1_LOC_826/a_8_24# VSS VDD AND2X1_LOC_56/B AND2X1_LOC_95/Y AND2X1_LOC

XAND2X1_LOC_420 AND2X1_LOC_420/a_36_24# OR2X1_LOC_447/A AND2X1_LOC_420/a_8_24# VSS VDD AND2X1_LOC_95/Y OR2X1_LOC_532/B AND2X1_LOC

XAND2X1_LOC_487 AND2X1_LOC_487/a_36_24# OR2X1_LOC_489/B AND2X1_LOC_487/a_8_24# VSS VDD OR2X1_LOC_160/B AND2X1_LOC_95/Y AND2X1_LOC

XAND2X1_LOC_626 AND2X1_LOC_626/a_36_24# OR2X1_LOC_629/B AND2X1_LOC_626/a_8_24# VSS VDD AND2X1_LOC_95/Y OR2X1_LOC_161/A AND2X1_LOC

XAND2X1_LOC_406 AND2X1_LOC_406/a_36_24# OR2X1_LOC_475/B AND2X1_LOC_406/a_8_24# VSS VDD AND2X1_LOC_95/Y OR2X1_LOC_405/Y AND2X1_LOC

XAND2X1_LOC_597 AND2X1_LOC_597/a_36_24# OR2X1_LOC_644/B AND2X1_LOC_597/a_8_24# VSS VDD AND2X1_LOC_41/A OR2X1_LOC_596/Y AND2X1_LOC

XOR2X1_LOC_448 OR2X1_LOC_448/a_8_216# OR2X1_LOC_448/a_36_216# OR2X1_LOC_448/Y VSS VDD OR2X1_LOC_448/A OR2X1_LOC_448/B OR2X1_LOC

XOR2X1_LOC_355 OR2X1_LOC_355/a_8_216# OR2X1_LOC_355/a_36_216# OR2X1_LOC_356/A VSS VDD OR2X1_LOC_355/A OR2X1_LOC_355/B OR2X1_LOC

XOR2X1_LOC_176 OR2X1_LOC_176/a_8_216# OR2X1_LOC_176/a_36_216# OR2X1_LOC_176/Y VSS VDD OR2X1_LOC_91/A OR2X1_LOC_26/Y OR2X1_LOC

XOR2X1_LOC_290 OR2X1_LOC_290/a_8_216# OR2X1_LOC_290/a_36_216# OR2X1_LOC_290/Y VSS VDD OR2X1_LOC_26/Y OR2X1_LOC_16/A OR2X1_LOC

XOR2X1_LOC_677 OR2X1_LOC_677/a_8_216# OR2X1_LOC_677/a_36_216# OR2X1_LOC_677/Y VSS VDD OR2X1_LOC_427/A OR2X1_LOC_26/Y OR2X1_LOC

XOR2X1_LOC_83 OR2X1_LOC_83/a_8_216# OR2X1_LOC_83/a_36_216# OR2X1_LOC_83/Y VSS VDD OR2X1_LOC_83/A OR2X1_LOC_26/Y OR2X1_LOC

XOR2X1_LOC_237 OR2X1_LOC_237/a_8_216# OR2X1_LOC_237/a_36_216# OR2X1_LOC_237/Y VSS VDD OR2X1_LOC_428/A OR2X1_LOC_26/Y OR2X1_LOC

XAND2X1_LOC_668 AND2X1_LOC_668/a_36_24# OR2X1_LOC_669/A AND2X1_LOC_668/a_8_24# VSS VDD OR2X1_LOC_26/Y OR2X1_LOC_158/A AND2X1_LOC

XOR2X1_LOC_595 OR2X1_LOC_595/a_8_216# OR2X1_LOC_595/a_36_216# OR2X1_LOC_595/Y VSS VDD OR2X1_LOC_595/A OR2X1_LOC_26/Y OR2X1_LOC

XOR2X1_LOC_27 OR2X1_LOC_27/a_8_216# OR2X1_LOC_27/a_36_216# OR2X1_LOC_27/Y VSS VDD OR2X1_LOC_26/Y OR2X1_LOC_7/A OR2X1_LOC

XOR2X1_LOC_385 OR2X1_LOC_385/a_8_216# OR2X1_LOC_385/a_36_216# OR2X1_LOC_385/Y VSS VDD OR2X1_LOC_600/A OR2X1_LOC_26/Y OR2X1_LOC

XOR2X1_LOC_311 OR2X1_LOC_311/a_8_216# OR2X1_LOC_311/a_36_216# OR2X1_LOC_311/Y VSS VDD OR2X1_LOC_485/A OR2X1_LOC_26/Y OR2X1_LOC

XOR2X1_LOC_146 OR2X1_LOC_146/a_8_216# OR2X1_LOC_146/a_36_216# OR2X1_LOC_146/Y VSS VDD OR2X1_LOC_744/A OR2X1_LOC_36/Y OR2X1_LOC

XOR2X1_LOC_179 OR2X1_LOC_179/a_8_216# OR2X1_LOC_179/a_36_216# OR2X1_LOC_179/Y VSS VDD OR2X1_LOC_600/A OR2X1_LOC_36/Y OR2X1_LOC

XOR2X1_LOC_484 OR2X1_LOC_484/a_8_216# OR2X1_LOC_484/a_36_216# OR2X1_LOC_484/Y VSS VDD OR2X1_LOC_36/Y OR2X1_LOC_13/B OR2X1_LOC

XOR2X1_LOC_495 OR2X1_LOC_495/a_8_216# OR2X1_LOC_495/a_36_216# OR2X1_LOC_495/Y VSS VDD OR2X1_LOC_56/A OR2X1_LOC_36/Y OR2X1_LOC

XOR2X1_LOC_627 OR2X1_LOC_627/a_8_216# OR2X1_LOC_627/a_36_216# OR2X1_LOC_627/Y VSS VDD OR2X1_LOC_36/Y OR2X1_LOC_7/A OR2X1_LOC

XOR2X1_LOC_754 OR2X1_LOC_754/a_8_216# OR2X1_LOC_754/a_36_216# OR2X1_LOC_754/Y VSS VDD OR2X1_LOC_754/A OR2X1_LOC_36/Y OR2X1_LOC

XOR2X1_LOC_69 OR2X1_LOC_69/a_8_216# OR2X1_LOC_69/a_36_216# OR2X1_LOC_69/Y VSS VDD OR2X1_LOC_69/A OR2X1_LOC_36/Y OR2X1_LOC

XOR2X1_LOC_39 OR2X1_LOC_39/a_8_216# OR2X1_LOC_39/a_36_216# OR2X1_LOC_39/Y VSS VDD OR2X1_LOC_39/A OR2X1_LOC_36/Y OR2X1_LOC

XOR2X1_LOC_396 OR2X1_LOC_396/a_8_216# OR2X1_LOC_396/a_36_216# OR2X1_LOC_396/Y VSS VDD OR2X1_LOC_36/Y OR2X1_LOC_45/B OR2X1_LOC

XOR2X1_LOC_320 OR2X1_LOC_320/a_8_216# OR2X1_LOC_320/a_36_216# OR2X1_LOC_320/Y VSS VDD OR2X1_LOC_91/A OR2X1_LOC_36/Y OR2X1_LOC

XOR2X1_LOC_497 OR2X1_LOC_497/a_8_216# OR2X1_LOC_497/a_36_216# OR2X1_LOC_497/Y VSS VDD OR2X1_LOC_71/Y OR2X1_LOC_22/Y OR2X1_LOC

XOR2X1_LOC_615 OR2X1_LOC_615/a_8_216# OR2X1_LOC_615/a_36_216# OR2X1_LOC_615/Y VSS VDD OR2X1_LOC_754/A OR2X1_LOC_22/Y OR2X1_LOC

XOR2X1_LOC_24 OR2X1_LOC_24/a_8_216# OR2X1_LOC_24/a_36_216# OR2X1_LOC_24/Y VSS VDD OR2X1_LOC_45/B OR2X1_LOC_22/Y OR2X1_LOC

XOR2X1_LOC_58 OR2X1_LOC_58/a_8_216# OR2X1_LOC_58/a_36_216# OR2X1_LOC_58/Y VSS VDD OR2X1_LOC_52/B OR2X1_LOC_22/Y OR2X1_LOC

XOR2X1_LOC_522 OR2X1_LOC_522/a_8_216# OR2X1_LOC_522/a_36_216# OR2X1_LOC_522/Y VSS VDD OR2X1_LOC_485/A OR2X1_LOC_22/Y OR2X1_LOC

XOR2X1_LOC_589 OR2X1_LOC_589/a_8_216# OR2X1_LOC_589/a_36_216# OR2X1_LOC_589/Y VSS VDD OR2X1_LOC_589/A OR2X1_LOC_22/Y OR2X1_LOC

XAND2X1_LOC_549 AND2X1_LOC_549/a_36_24# AND2X1_LOC_549/Y AND2X1_LOC_549/a_8_24# VSS VDD OR2X1_LOC_531/Y AND2X1_LOC_548/Y AND2X1_LOC

XOR2X1_LOC_709 OR2X1_LOC_709/a_8_216# OR2X1_LOC_709/a_36_216# OR2X1_LOC_711/B VSS VDD OR2X1_LOC_709/A OR2X1_LOC_709/B OR2X1_LOC

XOR2X1_LOC_706 OR2X1_LOC_706/a_8_216# OR2X1_LOC_706/a_36_216# OR2X1_LOC_713/A VSS VDD OR2X1_LOC_706/A OR2X1_LOC_706/B OR2X1_LOC

XAND2X1_LOC_335 AND2X1_LOC_335/a_36_24# AND2X1_LOC_335/Y AND2X1_LOC_335/a_8_24# VSS VDD OR2X1_LOC_309/Y OR2X1_LOC_310/Y AND2X1_LOC

XAND2X1_LOC_778 AND2X1_LOC_778/a_36_24# AND2X1_LOC_778/Y AND2X1_LOC_778/a_8_24# VSS VDD OR2X1_LOC_371/Y OR2X1_LOC_496/Y AND2X1_LOC

XAND2X1_LOC_198 AND2X1_LOC_198/a_36_24# AND2X1_LOC_208/B AND2X1_LOC_198/a_8_24# VSS VDD OR2X1_LOC_57/Y AND2X1_LOC_197/Y AND2X1_LOC

XOR2X1_LOC_72 OR2X1_LOC_72/a_8_216# OR2X1_LOC_72/a_36_216# OR2X1_LOC_72/Y VSS VDD OR2X1_LOC_71/Y OR2X1_LOC_70/Y OR2X1_LOC

XOR2X1_LOC_184 OR2X1_LOC_184/a_8_216# OR2X1_LOC_184/a_36_216# OR2X1_LOC_184/Y VSS VDD OR2X1_LOC_95/Y OR2X1_LOC_71/Y OR2X1_LOC

XAND2X1_LOC_151 AND2X1_LOC_151/a_36_24# OR2X1_LOC_152/A AND2X1_LOC_151/a_8_24# VSS VDD OR2X1_LOC_56/A OR2X1_LOC_437/A AND2X1_LOC

XAND2X1_LOC_186 AND2X1_LOC_186/a_36_24# OR2X1_LOC_680/A AND2X1_LOC_186/a_8_24# VSS VDD OR2X1_LOC_437/A OR2X1_LOC_816/A AND2X1_LOC

XOR2X1_LOC_292 OR2X1_LOC_292/a_8_216# OR2X1_LOC_292/a_36_216# OR2X1_LOC_292/Y VSS VDD OR2X1_LOC_437/A OR2X1_LOC_40/Y OR2X1_LOC

XOR2X1_LOC_173 OR2X1_LOC_173/a_8_216# OR2X1_LOC_173/a_36_216# OR2X1_LOC_173/Y VSS VDD OR2X1_LOC_437/A OR2X1_LOC_70/Y OR2X1_LOC

XOR2X1_LOC_235 OR2X1_LOC_235/a_8_216# OR2X1_LOC_235/a_36_216# OR2X1_LOC_235/Y VSS VDD OR2X1_LOC_86/A OR2X1_LOC_235/B OR2X1_LOC

XAND2X1_LOC_777 AND2X1_LOC_777/a_36_24# AND2X1_LOC_784/A AND2X1_LOC_777/a_8_24# VSS VDD OR2X1_LOC_246/A OR2X1_LOC_305/Y AND2X1_LOC

XAND2X1_LOC_633 AND2X1_LOC_633/a_36_24# AND2X1_LOC_633/Y AND2X1_LOC_633/a_8_24# VSS VDD OR2X1_LOC_118/Y OR2X1_LOC_278/A AND2X1_LOC

XAND2X1_LOC_541 AND2X1_LOC_541/a_36_24# AND2X1_LOC_541/Y AND2X1_LOC_541/a_8_24# VSS VDD OR2X1_LOC_256/A OR2X1_LOC_272/Y AND2X1_LOC

XAND2X1_LOC_634 AND2X1_LOC_634/a_36_24# AND2X1_LOC_634/Y AND2X1_LOC_634/a_8_24# VSS VDD OR2X1_LOC_290/Y OR2X1_LOC_690/A AND2X1_LOC

XOR2X1_LOC_813 OR2X1_LOC_813/a_8_216# OR2X1_LOC_813/a_36_216# OR2X1_LOC_813/Y VSS VDD OR2X1_LOC_813/A OR2X1_LOC_235/B OR2X1_LOC

XAND2X1_LOC_266 AND2X1_LOC_266/a_36_24# AND2X1_LOC_266/Y AND2X1_LOC_266/a_8_24# VSS VDD OR2X1_LOC_262/Y OR2X1_LOC_813/A AND2X1_LOC

XOR2X1_LOC_622 OR2X1_LOC_622/a_8_216# OR2X1_LOC_622/a_36_216# OR2X1_LOC_624/B VSS VDD OR2X1_LOC_622/A OR2X1_LOC_622/B OR2X1_LOC

XAND2X1_LOC_673 AND2X1_LOC_673/a_36_24# AND2X1_LOC_721/A AND2X1_LOC_673/a_8_24# VSS VDD OR2X1_LOC_670/Y OR2X1_LOC_672/Y AND2X1_LOC

XAND2X1_LOC_69 AND2X1_LOC_69/a_36_24# AND2X1_LOC_69/Y AND2X1_LOC_69/a_8_24# VSS VDD AND2X1_LOC_36/Y OR2X1_LOC_68/Y AND2X1_LOC

XOR2X1_LOC_198 OR2X1_LOC_198/a_8_216# OR2X1_LOC_198/a_36_216# OR2X1_LOC_208/A VSS VDD OR2X1_LOC_198/A AND2X1_LOC_57/Y OR2X1_LOC

XOR2X1_LOC_335 OR2X1_LOC_335/a_8_216# OR2X1_LOC_335/a_36_216# OR2X1_LOC_335/Y VSS VDD OR2X1_LOC_335/A OR2X1_LOC_335/B OR2X1_LOC

XOR2X1_LOC_778 OR2X1_LOC_778/a_8_216# OR2X1_LOC_778/a_36_216# OR2X1_LOC_778/Y VSS VDD OR2X1_LOC_778/A OR2X1_LOC_778/B OR2X1_LOC

XOR2X1_LOC_117 OR2X1_LOC_117/a_8_216# OR2X1_LOC_117/a_36_216# OR2X1_LOC_117/Y VSS VDD OR2X1_LOC_70/Y OR2X1_LOC_65/B OR2X1_LOC

XOR2X1_LOC_262 OR2X1_LOC_262/a_8_216# OR2X1_LOC_262/a_36_216# OR2X1_LOC_262/Y VSS VDD OR2X1_LOC_65/B OR2X1_LOC_40/Y OR2X1_LOC

XOR2X1_LOC_65 OR2X1_LOC_65/a_8_216# OR2X1_LOC_65/a_36_216# OR2X1_LOC_65/Y VSS VDD OR2X1_LOC_64/Y OR2X1_LOC_65/B OR2X1_LOC

XOR2X1_LOC_464 OR2X1_LOC_464/a_8_216# OR2X1_LOC_464/a_36_216# OR2X1_LOC_471/B VSS VDD OR2X1_LOC_464/A OR2X1_LOC_464/B OR2X1_LOC

XAND2X1_LOC_301 AND2X1_LOC_301/a_36_24# AND2X1_LOC_303/A AND2X1_LOC_301/a_8_24# VSS VDD OR2X1_LOC_75/Y OR2X1_LOC_300/Y AND2X1_LOC

XAND2X1_LOC_831 AND2X1_LOC_831/a_36_24# AND2X1_LOC_831/Y AND2X1_LOC_831/a_8_24# VSS VDD OR2X1_LOC_273/Y OR2X1_LOC_300/Y AND2X1_LOC

XAND2X1_LOC_302 AND2X1_LOC_302/a_36_24# AND2X1_LOC_303/B AND2X1_LOC_302/a_8_24# VSS VDD OR2X1_LOC_298/Y OR2X1_LOC_299/Y AND2X1_LOC

XAND2X1_LOC_370 AND2X1_LOC_370/a_36_24# AND2X1_LOC_787/A AND2X1_LOC_370/a_8_24# VSS VDD OR2X1_LOC_309/Y OR2X1_LOC_369/Y AND2X1_LOC

XAND2X1_LOC_543 AND2X1_LOC_543/a_36_24# AND2X1_LOC_543/Y AND2X1_LOC_543/a_8_24# VSS VDD OR2X1_LOC_315/Y OR2X1_LOC_369/Y AND2X1_LOC

XOR2X1_LOC_832 OR2X1_LOC_832/a_8_216# OR2X1_LOC_832/a_36_216# OR2X1_LOC_841/A VSS VDD OR2X1_LOC_435/A OR2X1_LOC_449/B OR2X1_LOC

XOR2X1_LOC_435 OR2X1_LOC_435/a_8_216# OR2X1_LOC_435/a_36_216# OR2X1_LOC_435/Y VSS VDD OR2X1_LOC_435/A OR2X1_LOC_435/B OR2X1_LOC

XOR2X1_LOC_831 OR2X1_LOC_831/a_8_216# OR2X1_LOC_831/a_36_216# OR2X1_LOC_841/B VSS VDD OR2X1_LOC_831/A OR2X1_LOC_831/B OR2X1_LOC

XOR2X1_LOC_828 OR2X1_LOC_828/a_8_216# OR2X1_LOC_828/a_36_216# OR2X1_LOC_828/Y VSS VDD OR2X1_LOC_598/Y OR2X1_LOC_828/B OR2X1_LOC

XOR2X1_LOC_780 OR2X1_LOC_780/a_8_216# OR2X1_LOC_780/a_36_216# OR2X1_LOC_783/A VSS VDD OR2X1_LOC_780/A OR2X1_LOC_780/B OR2X1_LOC

XOR2X1_LOC_156 OR2X1_LOC_156/a_8_216# OR2X1_LOC_156/a_36_216# OR2X1_LOC_156/Y VSS VDD OR2X1_LOC_156/A OR2X1_LOC_156/B OR2X1_LOC

XOR2X1_LOC_708 OR2X1_LOC_708/a_8_216# OR2X1_LOC_708/a_36_216# OR2X1_LOC_708/Y VSS VDD OR2X1_LOC_779/A OR2X1_LOC_708/B OR2X1_LOC

XOR2X1_LOC_308 OR2X1_LOC_308/a_8_216# OR2X1_LOC_308/a_36_216# OR2X1_LOC_308/Y VSS VDD OR2X1_LOC_308/A OR2X1_LOC_512/A OR2X1_LOC

XOR2X1_LOC_147 OR2X1_LOC_147/a_8_216# OR2X1_LOC_147/a_36_216# OR2X1_LOC_149/B VSS VDD OR2X1_LOC_147/A OR2X1_LOC_147/B OR2X1_LOC

XOR2X1_LOC_168 OR2X1_LOC_168/a_8_216# OR2X1_LOC_168/a_36_216# OR2X1_LOC_168/Y VSS VDD OR2X1_LOC_168/A OR2X1_LOC_168/B OR2X1_LOC

XOR2X1_LOC_776 OR2X1_LOC_776/a_8_216# OR2X1_LOC_776/a_36_216# OR2X1_LOC_776/Y VSS VDD OR2X1_LOC_776/A OR2X1_LOC_168/B OR2X1_LOC

XOR2X1_LOC_325 OR2X1_LOC_325/a_8_216# OR2X1_LOC_325/a_36_216# OR2X1_LOC_325/Y VSS VDD OR2X1_LOC_325/A OR2X1_LOC_325/B OR2X1_LOC

XOR2X1_LOC_459 OR2X1_LOC_459/a_8_216# OR2X1_LOC_459/a_36_216# OR2X1_LOC_463/B VSS VDD OR2X1_LOC_459/A OR2X1_LOC_459/B OR2X1_LOC

XOR2X1_LOC_638 OR2X1_LOC_638/a_8_216# OR2X1_LOC_638/a_36_216# OR2X1_LOC_651/B VSS VDD OR2X1_LOC_637/Y OR2X1_LOC_638/B OR2X1_LOC

XOR2X1_LOC_416 OR2X1_LOC_416/a_8_216# OR2X1_LOC_416/a_36_216# OR2X1_LOC_416/Y VSS VDD OR2X1_LOC_416/A OR2X1_LOC_158/A OR2X1_LOC

XAND2X1_LOC_637 AND2X1_LOC_637/a_36_24# AND2X1_LOC_637/Y AND2X1_LOC_637/a_8_24# VSS VDD OR2X1_LOC_585/Y OR2X1_LOC_586/Y AND2X1_LOC

XOR2X1_LOC_481 OR2X1_LOC_481/a_8_216# OR2X1_LOC_481/a_36_216# OR2X1_LOC_481/Y VSS VDD OR2X1_LOC_481/A OR2X1_LOC_3/Y OR2X1_LOC

XAND2X1_LOC_631 AND2X1_LOC_631/a_36_24# AND2X1_LOC_631/Y AND2X1_LOC_631/a_8_24# VSS VDD AND2X1_LOC_483/Y OR2X1_LOC_625/Y AND2X1_LOC

XOR2X1_LOC_196 OR2X1_LOC_196/a_8_216# OR2X1_LOC_196/a_36_216# OR2X1_LOC_196/Y VSS VDD AND2X1_LOC_48/Y OR2X1_LOC_196/B OR2X1_LOC

XOR2X1_LOC_520 OR2X1_LOC_520/a_8_216# OR2X1_LOC_520/a_36_216# OR2X1_LOC_520/Y VSS VDD OR2X1_LOC_520/A OR2X1_LOC_520/B OR2X1_LOC

XOR2X1_LOC_834 OR2X1_LOC_834/a_8_216# OR2X1_LOC_834/a_36_216# OR2X1_LOC_840/A VSS VDD OR2X1_LOC_834/A OR2X1_LOC_779/B OR2X1_LOC

XOR2X1_LOC_779 OR2X1_LOC_779/a_8_216# OR2X1_LOC_779/a_36_216# OR2X1_LOC_779/Y VSS VDD OR2X1_LOC_779/A OR2X1_LOC_779/B OR2X1_LOC

XAND2X1_LOC_98 AND2X1_LOC_98/a_36_24# AND2X1_LOC_98/Y AND2X1_LOC_98/a_8_24# VSS VDD OR2X1_LOC_93/Y OR2X1_LOC_96/Y AND2X1_LOC

XAND2X1_LOC_630 AND2X1_LOC_630/a_36_24# AND2X1_LOC_632/A AND2X1_LOC_630/a_8_24# VSS VDD OR2X1_LOC_628/Y AND2X1_LOC_629/Y AND2X1_LOC

XAND2X1_LOC_448 AND2X1_LOC_448/a_36_24# AND2X1_LOC_448/Y AND2X1_LOC_448/a_8_24# VSS VDD OR2X1_LOC_421/Y OR2X1_LOC_422/Y AND2X1_LOC

XOR2X1_LOC_154 OR2X1_LOC_154/a_8_216# OR2X1_LOC_154/a_36_216# OR2X1_LOC_156/B VSS VDD OR2X1_LOC_154/A AND2X1_LOC_7/B OR2X1_LOC

XAND2X1_LOC_584 AND2X1_LOC_584/a_36_24# OR2X1_LOC_636/A AND2X1_LOC_584/a_8_24# VSS VDD AND2X1_LOC_7/B AND2X1_LOC_51/Y AND2X1_LOC

XAND2X1_LOC_368 AND2X1_LOC_368/a_36_24# OR2X1_LOC_457/B AND2X1_LOC_368/a_8_24# VSS VDD AND2X1_LOC_7/B OR2X1_LOC_270/Y AND2X1_LOC

XAND2X1_LOC_528 AND2X1_LOC_528/a_36_24# OR2X1_LOC_620/B AND2X1_LOC_528/a_8_24# VSS VDD AND2X1_LOC_7/B AND2X1_LOC_44/Y AND2X1_LOC

XOR2X1_LOC_247 OR2X1_LOC_247/a_8_216# OR2X1_LOC_247/a_36_216# OR2X1_LOC_247/Y VSS VDD AND2X1_LOC_41/A AND2X1_LOC_7/B OR2X1_LOC

XAND2X1_LOC_230 AND2X1_LOC_230/a_36_24# OR2X1_LOC_231/A AND2X1_LOC_230/a_8_24# VSS VDD AND2X1_LOC_7/B AND2X1_LOC_31/Y AND2X1_LOC

XAND2X1_LOC_627 AND2X1_LOC_627/a_36_24# OR2X1_LOC_629/A AND2X1_LOC_627/a_8_24# VSS VDD AND2X1_LOC_7/B AND2X1_LOC_36/Y AND2X1_LOC

XOR2X1_LOC_130 OR2X1_LOC_130/a_8_216# OR2X1_LOC_130/a_36_216# OR2X1_LOC_130/Y VSS VDD OR2X1_LOC_130/A AND2X1_LOC_7/B OR2X1_LOC

XAND2X1_LOC_344 AND2X1_LOC_344/a_36_24# AND2X1_LOC_348/A AND2X1_LOC_344/a_8_24# VSS VDD AND2X1_LOC_456/B OR2X1_LOC_256/Y AND2X1_LOC

XOR2X1_LOC_105 OR2X1_LOC_105/a_8_216# OR2X1_LOC_105/a_36_216# OR2X1_LOC_105/Y VSS VDD OR2X1_LOC_756/B OR2X1_LOC_78/A OR2X1_LOC

XAND2X1_LOC_179 AND2X1_LOC_179/a_36_24# OR2X1_LOC_181/A AND2X1_LOC_179/a_8_24# VSS VDD AND2X1_LOC_36/Y OR2X1_LOC_756/B AND2X1_LOC

XAND2X1_LOC_600 AND2X1_LOC_600/a_36_24# OR2X1_LOC_602/B AND2X1_LOC_600/a_8_24# VSS VDD AND2X1_LOC_31/Y OR2X1_LOC_756/B AND2X1_LOC

XAND2X1_LOC_261 AND2X1_LOC_261/a_36_24# OR2X1_LOC_345/A AND2X1_LOC_261/a_8_24# VSS VDD OR2X1_LOC_756/B OR2X1_LOC_260/Y AND2X1_LOC

XAND2X1_LOC_616 AND2X1_LOC_616/a_36_24# OR2X1_LOC_621/B AND2X1_LOC_616/a_8_24# VSS VDD AND2X1_LOC_18/Y OR2X1_LOC_756/B AND2X1_LOC

XOR2X1_LOC_756 OR2X1_LOC_756/a_8_216# OR2X1_LOC_756/a_36_216# OR2X1_LOC_756/Y VSS VDD OR2X1_LOC_161/A OR2X1_LOC_756/B OR2X1_LOC

XAND2X1_LOC_396 AND2X1_LOC_396/a_36_24# OR2X1_LOC_401/A AND2X1_LOC_396/a_8_24# VSS VDD OR2X1_LOC_160/B AND2X1_LOC_36/Y AND2X1_LOC

XAND2X1_LOC_505 AND2X1_LOC_505/a_36_24# OR2X1_LOC_507/A AND2X1_LOC_505/a_8_24# VSS VDD AND2X1_LOC_18/Y OR2X1_LOC_160/B AND2X1_LOC

XAND2X1_LOC_45 AND2X1_LOC_45/a_36_24# OR2X1_LOC_196/B AND2X1_LOC_45/a_8_24# VSS VDD OR2X1_LOC_160/B AND2X1_LOC_44/Y AND2X1_LOC

XAND2X1_LOC_695 AND2X1_LOC_695/a_36_24# OR2X1_LOC_707/A AND2X1_LOC_695/a_8_24# VSS VDD OR2X1_LOC_160/B AND2X1_LOC_47/Y AND2X1_LOC

XOR2X1_LOC_249 OR2X1_LOC_249/a_8_216# OR2X1_LOC_249/a_36_216# OR2X1_LOC_249/Y VSS VDD OR2X1_LOC_154/A OR2X1_LOC_160/B OR2X1_LOC

XOR2X1_LOC_160 OR2X1_LOC_160/a_8_216# OR2X1_LOC_160/a_36_216# OR2X1_LOC_160/Y VSS VDD OR2X1_LOC_160/A OR2X1_LOC_160/B OR2X1_LOC

XAND2X1_LOC_238 AND2X1_LOC_238/a_36_24# OR2X1_LOC_776/A AND2X1_LOC_238/a_8_24# VSS VDD OR2X1_LOC_160/B AND2X1_LOC_51/Y AND2X1_LOC

XOR2X1_LOC_789 OR2X1_LOC_789/a_8_216# OR2X1_LOC_789/a_36_216# OR2X1_LOC_793/B VSS VDD OR2X1_LOC_789/A OR2X1_LOC_789/B OR2X1_LOC

XAND2X1_LOC_557 AND2X1_LOC_557/a_36_24# AND2X1_LOC_557/Y AND2X1_LOC_557/a_8_24# VSS VDD AND2X1_LOC_489/Y OR2X1_LOC_490/Y AND2X1_LOC

XAND2X1_LOC_535 AND2X1_LOC_535/a_36_24# AND2X1_LOC_535/Y AND2X1_LOC_535/a_8_24# VSS VDD OR2X1_LOC_533/Y OR2X1_LOC_534/Y AND2X1_LOC

XAND2X1_LOC_195 AND2X1_LOC_195/a_36_24# AND2X1_LOC_199/A AND2X1_LOC_195/a_8_24# VSS VDD OR2X1_LOC_41/Y OR2X1_LOC_43/Y AND2X1_LOC

XAND2X1_LOC_506 AND2X1_LOC_506/a_36_24# AND2X1_LOC_508/A AND2X1_LOC_506/a_8_24# VSS VDD OR2X1_LOC_239/Y OR2X1_LOC_419/Y AND2X1_LOC

XAND2X1_LOC_447 AND2X1_LOC_447/a_36_24# AND2X1_LOC_447/Y AND2X1_LOC_447/a_8_24# VSS VDD OR2X1_LOC_419/Y OR2X1_LOC_420/Y AND2X1_LOC

XAND2X1_LOC_838 AND2X1_LOC_838/a_36_24# AND2X1_LOC_838/Y AND2X1_LOC_838/a_8_24# VSS VDD OR2X1_LOC_827/Y AND2X1_LOC_838/B AND2X1_LOC

XAND2X1_LOC_138 AND2X1_LOC_138/a_36_24# AND2X1_LOC_139/B AND2X1_LOC_138/a_8_24# VSS VDD OR2X1_LOC_135/Y OR2X1_LOC_136/Y AND2X1_LOC

XOR2X1_LOC_178 OR2X1_LOC_178/a_8_216# OR2X1_LOC_178/a_36_216# OR2X1_LOC_178/Y VSS VDD OR2X1_LOC_158/A OR2X1_LOC_56/A OR2X1_LOC

XOR2X1_LOC_826 OR2X1_LOC_826/a_8_216# OR2X1_LOC_826/a_36_216# OR2X1_LOC_826/Y VSS VDD OR2X1_LOC_95/Y OR2X1_LOC_56/A OR2X1_LOC

XOR2X1_LOC_613 OR2X1_LOC_613/a_8_216# OR2X1_LOC_613/a_36_216# OR2X1_LOC_613/Y VSS VDD OR2X1_LOC_56/A OR2X1_LOC_40/Y OR2X1_LOC

XOR2X1_LOC_67 OR2X1_LOC_67/a_8_216# OR2X1_LOC_67/a_36_216# OR2X1_LOC_67/Y VSS VDD OR2X1_LOC_67/A OR2X1_LOC_56/A OR2X1_LOC

XOR2X1_LOC_312 OR2X1_LOC_312/a_8_216# OR2X1_LOC_312/a_36_216# OR2X1_LOC_312/Y VSS VDD OR2X1_LOC_64/Y OR2X1_LOC_56/A OR2X1_LOC

XAND2X1_LOC_612 AND2X1_LOC_612/a_36_24# OR2X1_LOC_647/B AND2X1_LOC_612/a_8_24# VSS VDD OR2X1_LOC_610/Y AND2X1_LOC_612/B AND2X1_LOC

XOR2X1_LOC_313 OR2X1_LOC_313/a_8_216# OR2X1_LOC_313/a_36_216# OR2X1_LOC_313/Y VSS VDD OR2X1_LOC_91/A OR2X1_LOC_70/Y OR2X1_LOC

XOR2X1_LOC_132 OR2X1_LOC_132/a_8_216# OR2X1_LOC_132/a_36_216# OR2X1_LOC_132/Y VSS VDD OR2X1_LOC_95/Y OR2X1_LOC_91/A OR2X1_LOC

XOR2X1_LOC_305 OR2X1_LOC_305/a_8_216# OR2X1_LOC_305/a_36_216# OR2X1_LOC_305/Y VSS VDD OR2X1_LOC_91/A OR2X1_LOC_3/Y OR2X1_LOC

XAND2X1_LOC_383 AND2X1_LOC_383/a_36_24# OR2X1_LOC_494/A AND2X1_LOC_383/a_8_24# VSS VDD OR2X1_LOC_91/A OR2X1_LOC_428/A AND2X1_LOC

XOR2X1_LOC_91 OR2X1_LOC_91/a_8_216# OR2X1_LOC_91/a_36_216# OR2X1_LOC_91/Y VSS VDD OR2X1_LOC_91/A OR2X1_LOC_51/Y OR2X1_LOC

XOR2X1_LOC_766 OR2X1_LOC_766/a_8_216# OR2X1_LOC_766/a_36_216# OR2X1_LOC_766/Y VSS VDD OR2X1_LOC_91/A OR2X1_LOC_64/Y OR2X1_LOC

XAND2X1_LOC_825 AND2X1_LOC_825/a_36_24# OR2X1_LOC_837/B AND2X1_LOC_825/a_8_24# VSS VDD AND2X1_LOC_44/Y AND2X1_LOC_94/Y AND2X1_LOC

XOR2X1_LOC_670 OR2X1_LOC_670/a_8_216# OR2X1_LOC_670/a_36_216# OR2X1_LOC_670/Y VSS VDD OR2X1_LOC_485/A OR2X1_LOC_40/Y OR2X1_LOC

XAND2X1_LOC_532 AND2X1_LOC_532/a_36_24# OR2X1_LOC_533/A AND2X1_LOC_532/a_8_24# VSS VDD OR2X1_LOC_485/A OR2X1_LOC_744/A AND2X1_LOC

XOR2X1_LOC_822 OR2X1_LOC_822/a_8_216# OR2X1_LOC_822/a_36_216# OR2X1_LOC_822/Y VSS VDD OR2X1_LOC_485/A OR2X1_LOC_64/Y OR2X1_LOC

XOR2X1_LOC_282 OR2X1_LOC_282/a_8_216# OR2X1_LOC_282/a_36_216# OR2X1_LOC_282/Y VSS VDD OR2X1_LOC_158/A OR2X1_LOC_485/A OR2X1_LOC

XOR2X1_LOC_420 OR2X1_LOC_420/a_8_216# OR2X1_LOC_420/a_36_216# OR2X1_LOC_420/Y VSS VDD OR2X1_LOC_485/A OR2X1_LOC_95/Y OR2X1_LOC

XOR2X1_LOC_239 OR2X1_LOC_239/a_8_216# OR2X1_LOC_239/a_36_216# OR2X1_LOC_239/Y VSS VDD OR2X1_LOC_485/A OR2X1_LOC_51/Y OR2X1_LOC

XOR2X1_LOC_172 OR2X1_LOC_172/a_8_216# OR2X1_LOC_172/a_36_216# OR2X1_LOC_172/Y VSS VDD OR2X1_LOC_485/A OR2X1_LOC_70/Y OR2X1_LOC

XAND2X1_LOC_590 AND2X1_LOC_590/a_36_24# OR2X1_LOC_591/A AND2X1_LOC_590/a_8_24# VSS VDD OR2X1_LOC_39/A OR2X1_LOC_485/A AND2X1_LOC

XOR2X1_LOC_342 OR2X1_LOC_342/a_8_216# OR2X1_LOC_342/a_36_216# OR2X1_LOC_349/B VSS VDD OR2X1_LOC_342/A OR2X1_LOC_342/B OR2X1_LOC

XAND2X1_LOC_843 AND2X1_LOC_843/a_36_24# AND2X1_LOC_843/Y AND2X1_LOC_843/a_8_24# VSS VDD OR2X1_LOC_251/Y OR2X1_LOC_278/Y AND2X1_LOC

XAND2X1_LOC_287 AND2X1_LOC_287/a_36_24# AND2X1_LOC_287/Y AND2X1_LOC_287/a_8_24# VSS VDD OR2X1_LOC_278/Y AND2X1_LOC_287/B AND2X1_LOC

XOR2X1_LOC_608 OR2X1_LOC_608/a_8_216# OR2X1_LOC_608/a_36_216# OR2X1_LOC_608/Y VSS VDD OR2X1_LOC_185/A OR2X1_LOC_78/B OR2X1_LOC

XAND2X1_LOC_601 AND2X1_LOC_601/a_36_24# OR2X1_LOC_602/A AND2X1_LOC_601/a_8_24# VSS VDD OR2X1_LOC_78/B AND2X1_LOC_47/Y AND2X1_LOC

XOR2X1_LOC_78 OR2X1_LOC_78/a_8_216# OR2X1_LOC_78/a_36_216# OR2X1_LOC_78/Y VSS VDD OR2X1_LOC_78/A OR2X1_LOC_78/B OR2X1_LOC

XAND2X1_LOC_232 AND2X1_LOC_232/a_36_24# OR2X1_LOC_240/B AND2X1_LOC_232/a_8_24# VSS VDD OR2X1_LOC_78/B OR2X1_LOC_375/A AND2X1_LOC

XAND2X1_LOC_418 AND2X1_LOC_418/a_36_24# OR2X1_LOC_446/A AND2X1_LOC_418/a_8_24# VSS VDD OR2X1_LOC_78/B AND2X1_LOC_51/Y AND2X1_LOC

XAND2X1_LOC_526 AND2X1_LOC_526/a_36_24# OR2X1_LOC_546/A AND2X1_LOC_526/a_8_24# VSS VDD AND2X1_LOC_31/Y OR2X1_LOC_161/A AND2X1_LOC

XAND2X1_LOC_669 AND2X1_LOC_669/a_36_24# OR2X1_LOC_720/A AND2X1_LOC_669/a_8_24# VSS VDD OR2X1_LOC_161/A OR2X1_LOC_668/Y AND2X1_LOC

XOR2X1_LOC_161 OR2X1_LOC_161/a_8_216# OR2X1_LOC_161/a_36_216# OR2X1_LOC_162/A VSS VDD OR2X1_LOC_161/A OR2X1_LOC_161/B OR2X1_LOC

XAND2X1_LOC_525 AND2X1_LOC_525/a_36_24# OR2X1_LOC_546/B AND2X1_LOC_525/a_8_24# VSS VDD AND2X1_LOC_41/A AND2X1_LOC_51/Y AND2X1_LOC

XAND2X1_LOC_504 AND2X1_LOC_504/a_36_24# OR2X1_LOC_507/B AND2X1_LOC_504/a_8_24# VSS VDD AND2X1_LOC_41/A OR2X1_LOC_375/A AND2X1_LOC

XAND2X1_LOC_484 AND2X1_LOC_484/a_36_24# OR2X1_LOC_486/B AND2X1_LOC_484/a_8_24# VSS VDD AND2X1_LOC_41/A AND2X1_LOC_36/Y AND2X1_LOC

XOR2X1_LOC_848 OR2X1_LOC_848/a_8_216# OR2X1_LOC_848/a_36_216# OR2X1_LOC_859/B VSS VDD OR2X1_LOC_848/A OR2X1_LOC_848/B OR2X1_LOC

XAND2X1_LOC_154 AND2X1_LOC_154/a_36_24# AND2X1_LOC_154/Y AND2X1_LOC_154/a_8_24# VSS VDD OR2X1_LOC_7/A OR2X1_LOC_39/A AND2X1_LOC

XAND2X1_LOC_188 AND2X1_LOC_188/a_36_24# OR2X1_LOC_189/A AND2X1_LOC_188/a_8_24# VSS VDD OR2X1_LOC_39/A OR2X1_LOC_816/A AND2X1_LOC

XOR2X1_LOC_617 OR2X1_LOC_617/a_8_216# OR2X1_LOC_617/a_36_216# OR2X1_LOC_617/Y VSS VDD OR2X1_LOC_51/Y OR2X1_LOC_39/A OR2X1_LOC

XOR2X1_LOC_393 OR2X1_LOC_393/a_8_216# OR2X1_LOC_393/a_36_216# OR2X1_LOC_393/Y VSS VDD OR2X1_LOC_40/Y OR2X1_LOC_39/A OR2X1_LOC

XAND2X1_LOC_249 AND2X1_LOC_249/a_36_24# OR2X1_LOC_595/A AND2X1_LOC_249/a_8_24# VSS VDD OR2X1_LOC_45/B OR2X1_LOC_39/A AND2X1_LOC

XAND2X1_LOC_391 AND2X1_LOC_391/a_36_24# AND2X1_LOC_391/Y AND2X1_LOC_391/a_8_24# VSS VDD OR2X1_LOC_382/Y OR2X1_LOC_384/Y AND2X1_LOC

XOR2X1_LOC_823 OR2X1_LOC_823/a_8_216# OR2X1_LOC_823/a_36_216# OR2X1_LOC_823/Y VSS VDD OR2X1_LOC_428/A OR2X1_LOC_51/Y OR2X1_LOC

XOR2X1_LOC_697 OR2X1_LOC_697/a_8_216# OR2X1_LOC_697/a_36_216# OR2X1_LOC_697/Y VSS VDD OR2X1_LOC_428/A OR2X1_LOC_158/A OR2X1_LOC

XOR2X1_LOC_281 OR2X1_LOC_281/a_8_216# OR2X1_LOC_281/a_36_216# OR2X1_LOC_281/Y VSS VDD OR2X1_LOC_428/A OR2X1_LOC_3/Y OR2X1_LOC

XOR2X1_LOC_431 OR2X1_LOC_431/a_8_216# OR2X1_LOC_431/a_36_216# OR2X1_LOC_431/Y VSS VDD OR2X1_LOC_428/A OR2X1_LOC_70/Y OR2X1_LOC

XOR2X1_LOC_759 OR2X1_LOC_759/a_8_216# OR2X1_LOC_759/a_36_216# OR2X1_LOC_759/Y VSS VDD OR2X1_LOC_759/A OR2X1_LOC_428/A OR2X1_LOC

XAND2X1_LOC_32 AND2X1_LOC_32/a_36_24# OR2X1_LOC_34/A AND2X1_LOC_32/a_8_24# VSS VDD OR2X1_LOC_87/B AND2X1_LOC_31/Y AND2X1_LOC

XOR2X1_LOC_134 OR2X1_LOC_134/a_8_216# OR2X1_LOC_134/a_36_216# OR2X1_LOC_134/Y VSS VDD OR2X1_LOC_427/A OR2X1_LOC_95/Y OR2X1_LOC

XAND2X1_LOC_161 AND2X1_LOC_161/a_36_24# AND2X1_LOC_161/Y AND2X1_LOC_161/a_8_24# VSS VDD OR2X1_LOC_427/A OR2X1_LOC_604/A AND2X1_LOC

XOR2X1_LOC_253 OR2X1_LOC_253/a_8_216# OR2X1_LOC_253/a_36_216# OR2X1_LOC_253/Y VSS VDD OR2X1_LOC_427/A OR2X1_LOC_64/Y OR2X1_LOC

XOR2X1_LOC_427 OR2X1_LOC_427/a_8_216# OR2X1_LOC_427/a_36_216# OR2X1_LOC_427/Y VSS VDD OR2X1_LOC_427/A OR2X1_LOC_70/Y OR2X1_LOC

XAND2X1_LOC_676 AND2X1_LOC_676/a_36_24# OR2X1_LOC_679/B AND2X1_LOC_676/a_8_24# VSS VDD OR2X1_LOC_427/A OR2X1_LOC_599/A AND2X1_LOC

XAND2X1_LOC_614 AND2X1_LOC_614/a_36_24# OR2X1_LOC_754/A AND2X1_LOC_614/a_8_24# VSS VDD OR2X1_LOC_89/A OR2X1_LOC_427/A AND2X1_LOC

XOR2X1_LOC_227 OR2X1_LOC_227/a_8_216# OR2X1_LOC_227/a_36_216# OR2X1_LOC_227/Y VSS VDD OR2X1_LOC_227/A OR2X1_LOC_227/B OR2X1_LOC

XOR2X1_LOC_446 OR2X1_LOC_446/a_8_216# OR2X1_LOC_446/a_36_216# OR2X1_LOC_446/Y VSS VDD OR2X1_LOC_446/A OR2X1_LOC_446/B OR2X1_LOC

XOR2X1_LOC_704 OR2X1_LOC_704/a_8_216# OR2X1_LOC_704/a_36_216# OR2X1_LOC_714/A VSS VDD OR2X1_LOC_446/B OR2X1_LOC_317/B OR2X1_LOC

XOR2X1_LOC_333 OR2X1_LOC_333/a_8_216# OR2X1_LOC_333/a_36_216# OR2X1_LOC_338/B VSS VDD OR2X1_LOC_333/A OR2X1_LOC_333/B OR2X1_LOC

XOR2X1_LOC_489 OR2X1_LOC_489/a_8_216# OR2X1_LOC_489/a_36_216# OR2X1_LOC_772/B VSS VDD OR2X1_LOC_489/A OR2X1_LOC_489/B OR2X1_LOC

XOR2X1_LOC_286 OR2X1_LOC_286/a_8_216# OR2X1_LOC_286/a_36_216# OR2X1_LOC_286/Y VSS VDD OR2X1_LOC_285/Y OR2X1_LOC_286/B OR2X1_LOC

XOR2X1_LOC_370 OR2X1_LOC_370/a_8_216# OR2X1_LOC_370/a_36_216# OR2X1_LOC_787/B VSS VDD OR2X1_LOC_543/A OR2X1_LOC_335/B OR2X1_LOC

XOR2X1_LOC_516 OR2X1_LOC_516/a_8_216# OR2X1_LOC_516/a_36_216# OR2X1_LOC_516/Y VSS VDD OR2X1_LOC_516/A OR2X1_LOC_516/B OR2X1_LOC

XOR2X1_LOC_112 OR2X1_LOC_112/a_8_216# OR2X1_LOC_112/a_36_216# OR2X1_LOC_715/B VSS VDD OR2X1_LOC_112/A OR2X1_LOC_112/B OR2X1_LOC

XOR2X1_LOC_332 OR2X1_LOC_332/a_8_216# OR2X1_LOC_332/a_36_216# OR2X1_LOC_339/A VSS VDD OR2X1_LOC_702/A OR2X1_LOC_112/A OR2X1_LOC

XOR2X1_LOC_547 OR2X1_LOC_547/a_8_216# OR2X1_LOC_547/a_36_216# OR2X1_LOC_550/A VSS VDD OR2X1_LOC_620/B OR2X1_LOC_547/B OR2X1_LOC

XOR2X1_LOC_855 OR2X1_LOC_855/a_8_216# OR2X1_LOC_855/a_36_216# OR2X1_LOC_856/A VSS VDD OR2X1_LOC_855/A OR2X1_LOC_691/Y OR2X1_LOC

XOR2X1_LOC_729 OR2X1_LOC_729/a_8_216# OR2X1_LOC_729/a_36_216# OR2X1_LOC_730/A VSS VDD OR2X1_LOC_691/Y OR2X1_LOC_687/Y OR2X1_LOC

XAND2X1_LOC_462 AND2X1_LOC_462/a_36_24# AND2X1_LOC_462/Y AND2X1_LOC_462/a_8_24# VSS VDD OR2X1_LOC_416/Y AND2X1_LOC_462/B AND2X1_LOC

XAND2X1_LOC_240 AND2X1_LOC_240/a_36_24# AND2X1_LOC_240/Y AND2X1_LOC_240/a_8_24# VSS VDD OR2X1_LOC_232/Y OR2X1_LOC_234/Y AND2X1_LOC

XAND2X1_LOC_836 AND2X1_LOC_836/a_36_24# AND2X1_LOC_839/B AND2X1_LOC_836/a_8_24# VSS VDD OR2X1_LOC_823/Y OR2X1_LOC_824/Y AND2X1_LOC

XAND2X1_LOC_334 AND2X1_LOC_334/a_36_24# AND2X1_LOC_334/Y AND2X1_LOC_334/a_8_24# VSS VDD OR2X1_LOC_290/Y OR2X1_LOC_291/Y AND2X1_LOC

XAND2X1_LOC_701 AND2X1_LOC_701/a_36_24# OR2X1_LOC_710/A AND2X1_LOC_701/a_8_24# VSS VDD AND2X1_LOC_44/Y OR2X1_LOC_269/B AND2X1_LOC

XAND2X1_LOC_759 AND2X1_LOC_759/a_36_24# OR2X1_LOC_792/B AND2X1_LOC_759/a_8_24# VSS VDD OR2X1_LOC_269/B OR2X1_LOC_758/Y AND2X1_LOC

XAND2X1_LOC_823 AND2X1_LOC_823/a_36_24# OR2X1_LOC_836/B AND2X1_LOC_823/a_8_24# VSS VDD AND2X1_LOC_51/Y OR2X1_LOC_269/B AND2X1_LOC

XAND2X1_LOC_697 AND2X1_LOC_697/a_36_24# OR2X1_LOC_779/A AND2X1_LOC_697/a_8_24# VSS VDD OR2X1_LOC_375/A OR2X1_LOC_269/B AND2X1_LOC

XAND2X1_LOC_280 AND2X1_LOC_280/a_36_24# OR2X1_LOC_542/B AND2X1_LOC_280/a_8_24# VSS VDD AND2X1_LOC_47/Y OR2X1_LOC_269/B AND2X1_LOC

XOR2X1_LOC_383 OR2X1_LOC_383/a_8_216# OR2X1_LOC_383/a_36_216# OR2X1_LOC_383/Y VSS VDD OR2X1_LOC_269/B AND2X1_LOC_91/B OR2X1_LOC

XAND2X1_LOC_428 AND2X1_LOC_428/a_36_24# OR2X1_LOC_451/B AND2X1_LOC_428/a_8_24# VSS VDD AND2X1_LOC_31/Y OR2X1_LOC_269/B AND2X1_LOC

XAND2X1_LOC_583 AND2X1_LOC_583/a_36_24# OR2X1_LOC_636/B AND2X1_LOC_583/a_8_24# VSS VDD AND2X1_LOC_31/Y OR2X1_LOC_87/A AND2X1_LOC

XAND2X1_LOC_521 AND2X1_LOC_521/a_36_24# OR2X1_LOC_523/B AND2X1_LOC_521/a_8_24# VSS VDD AND2X1_LOC_18/Y OR2X1_LOC_87/A AND2X1_LOC

XAND2X1_LOC_747 AND2X1_LOC_747/a_36_24# OR2X1_LOC_782/B AND2X1_LOC_747/a_8_24# VSS VDD AND2X1_LOC_47/Y OR2X1_LOC_87/A AND2X1_LOC

XAND2X1_LOC_52 AND2X1_LOC_52/a_36_24# AND2X1_LOC_52/Y AND2X1_LOC_52/a_8_24# VSS VDD OR2X1_LOC_87/A AND2X1_LOC_51/Y AND2X1_LOC

XAND2X1_LOC_524 AND2X1_LOC_524/a_36_24# OR2X1_LOC_545/A AND2X1_LOC_524/a_8_24# VSS VDD AND2X1_LOC_47/Y OR2X1_LOC_161/B AND2X1_LOC

XOR2X1_LOC_676 OR2X1_LOC_676/a_8_216# OR2X1_LOC_676/a_36_216# OR2X1_LOC_676/Y VSS VDD OR2X1_LOC_598/Y OR2X1_LOC_161/B OR2X1_LOC

XAND2X1_LOC_315 AND2X1_LOC_315/a_36_24# OR2X1_LOC_318/B AND2X1_LOC_315/a_8_24# VSS VDD AND2X1_LOC_31/Y OR2X1_LOC_161/B AND2X1_LOC

XOR2X1_LOC_614 OR2X1_LOC_614/a_8_216# OR2X1_LOC_614/a_36_216# OR2X1_LOC_614/Y VSS VDD OR2X1_LOC_161/B OR2X1_LOC_78/A OR2X1_LOC

XAND2X1_LOC_279 AND2X1_LOC_279/a_36_24# OR2X1_LOC_284/B AND2X1_LOC_279/a_8_24# VSS VDD AND2X1_LOC_44/Y OR2X1_LOC_161/B AND2X1_LOC

XAND2X1_LOC_257 AND2X1_LOC_257/a_36_24# OR2X1_LOC_259/B AND2X1_LOC_257/a_8_24# VSS VDD AND2X1_LOC_18/Y OR2X1_LOC_161/B AND2X1_LOC

XAND2X1_LOC_130 AND2X1_LOC_130/a_36_24# OR2X1_LOC_131/A AND2X1_LOC_130/a_8_24# VSS VDD OR2X1_LOC_7/A OR2X1_LOC_589/A AND2X1_LOC

XOR2X1_LOC_586 OR2X1_LOC_586/a_8_216# OR2X1_LOC_586/a_36_216# OR2X1_LOC_586/Y VSS VDD OR2X1_LOC_589/A OR2X1_LOC_70/Y OR2X1_LOC

XAND2X1_LOC_789 AND2X1_LOC_789/a_36_24# AND2X1_LOC_789/Y AND2X1_LOC_789/a_8_24# VSS VDD OR2X1_LOC_748/Y OR2X1_LOC_751/Y AND2X1_LOC

XOR2X1_LOC_344 OR2X1_LOC_344/a_8_216# OR2X1_LOC_344/a_36_216# OR2X1_LOC_348/B VSS VDD OR2X1_LOC_344/A OR2X1_LOC_456/A OR2X1_LOC

XOR2X1_LOC_368 OR2X1_LOC_368/a_8_216# OR2X1_LOC_368/a_36_216# OR2X1_LOC_368/Y VSS VDD OR2X1_LOC_368/A OR2X1_LOC_7/A OR2X1_LOC

XOR2X1_LOC_423 OR2X1_LOC_423/a_8_216# OR2X1_LOC_423/a_36_216# OR2X1_LOC_423/Y VSS VDD OR2X1_LOC_64/Y OR2X1_LOC_7/A OR2X1_LOC

XOR2X1_LOC_7 OR2X1_LOC_7/a_8_216# OR2X1_LOC_7/a_36_216# OR2X1_LOC_7/Y VSS VDD OR2X1_LOC_7/A OR2X1_LOC_3/Y OR2X1_LOC

XOR2X1_LOC_584 OR2X1_LOC_584/a_8_216# OR2X1_LOC_584/a_36_216# OR2X1_LOC_584/Y VSS VDD OR2X1_LOC_51/Y OR2X1_LOC_7/A OR2X1_LOC

XAND2X1_LOC_247 AND2X1_LOC_247/a_36_24# OR2X1_LOC_248/A AND2X1_LOC_247/a_8_24# VSS VDD OR2X1_LOC_7/A OR2X1_LOC_13/B AND2X1_LOC

XOR2X1_LOC_183 OR2X1_LOC_183/a_8_216# OR2X1_LOC_183/a_36_216# OR2X1_LOC_183/Y VSS VDD OR2X1_LOC_40/Y OR2X1_LOC_7/A OR2X1_LOC

XAND2X1_LOC_20 AND2X1_LOC_20/a_36_24# OR2X1_LOC_33/B AND2X1_LOC_20/a_8_24# VSS VDD AND2X1_LOC_18/Y AND2X1_LOC_19/Y AND2X1_LOC

XOR2X1_LOC_557 OR2X1_LOC_557/a_8_216# OR2X1_LOC_557/a_36_216# OR2X1_LOC_561/B VSS VDD OR2X1_LOC_557/A OR2X1_LOC_772/B OR2X1_LOC

XOR2X1_LOC_127 OR2X1_LOC_127/a_8_216# OR2X1_LOC_127/a_36_216# OR2X1_LOC_127/Y VSS VDD OR2X1_LOC_744/A OR2X1_LOC_3/Y OR2X1_LOC

XAND2X1_LOC_160 AND2X1_LOC_160/a_36_24# AND2X1_LOC_160/Y AND2X1_LOC_160/a_8_24# VSS VDD OR2X1_LOC_45/B OR2X1_LOC_744/A AND2X1_LOC

XOR2X1_LOC_698 OR2X1_LOC_698/a_8_216# OR2X1_LOC_698/a_36_216# OR2X1_LOC_698/Y VSS VDD OR2X1_LOC_744/A OR2X1_LOC_64/Y OR2X1_LOC

XOR2X1_LOC_764 OR2X1_LOC_764/a_8_216# OR2X1_LOC_764/a_36_216# OR2X1_LOC_764/Y VSS VDD OR2X1_LOC_744/A OR2X1_LOC_40/Y OR2X1_LOC

XOR2X1_LOC_380 OR2X1_LOC_380/a_8_216# OR2X1_LOC_380/a_36_216# OR2X1_LOC_380/Y VSS VDD OR2X1_LOC_380/A OR2X1_LOC_744/A OR2X1_LOC

XAND2X1_LOC_756 AND2X1_LOC_756/a_36_24# OR2X1_LOC_757/A AND2X1_LOC_756/a_8_24# VSS VDD OR2X1_LOC_600/A OR2X1_LOC_604/A AND2X1_LOC

XOR2X1_LOC_125 OR2X1_LOC_125/a_8_216# OR2X1_LOC_125/a_36_216# OR2X1_LOC_125/Y VSS VDD OR2X1_LOC_600/A OR2X1_LOC_95/Y OR2X1_LOC

XOR2X1_LOC_442 OR2X1_LOC_442/a_8_216# OR2X1_LOC_442/a_36_216# OR2X1_LOC_442/Y VSS VDD OR2X1_LOC_600/A OR2X1_LOC_40/Y OR2X1_LOC

XOR2X1_LOC_261 OR2X1_LOC_261/a_8_216# OR2X1_LOC_261/a_36_216# OR2X1_LOC_261/Y VSS VDD OR2X1_LOC_261/A OR2X1_LOC_600/A OR2X1_LOC

XAND2X1_LOC_105 AND2X1_LOC_105/a_36_24# OR2X1_LOC_106/A AND2X1_LOC_105/a_8_24# VSS VDD OR2X1_LOC_89/A OR2X1_LOC_600/A AND2X1_LOC

XAND2X1_LOC_101 AND2X1_LOC_101/a_36_24# AND2X1_LOC_216/A AND2X1_LOC_101/a_8_24# VSS VDD AND2X1_LOC_99/Y AND2X1_LOC_101/B AND2X1_LOC

XOR2X1_LOC_473 OR2X1_LOC_473/a_8_216# OR2X1_LOC_473/a_36_216# OR2X1_LOC_473/Y VSS VDD OR2X1_LOC_473/A OR2X1_LOC_216/A OR2X1_LOC

XOR2X1_LOC_361 OR2X1_LOC_361/a_8_216# OR2X1_LOC_361/a_36_216# OR2X1_LOC_362/A VSS VDD OR2X1_LOC_473/A OR2X1_LOC_267/Y OR2X1_LOC

XAND2X1_LOC_516 AND2X1_LOC_516/a_36_24# OR2X1_LOC_574/A AND2X1_LOC_516/a_8_24# VSS VDD OR2X1_LOC_513/Y OR2X1_LOC_515/Y AND2X1_LOC

XOR2X1_LOC_809 OR2X1_LOC_809/a_8_216# OR2X1_LOC_809/a_36_216# OR2X1_LOC_810/A VSS VDD OR2X1_LOC_802/Y OR2X1_LOC_809/B OR2X1_LOC

XAND2X1_LOC_79 AND2X1_LOC_79/a_36_24# AND2X1_LOC_79/Y AND2X1_LOC_79/a_8_24# VSS VDD AND2X1_LOC_18/Y OR2X1_LOC_78/Y AND2X1_LOC

XAND2X1_LOC_666 AND2X1_LOC_666/a_36_24# OR2X1_LOC_719/A AND2X1_LOC_666/a_8_24# VSS VDD AND2X1_LOC_18/Y OR2X1_LOC_121/A AND2X1_LOC

XAND2X1_LOC_496 AND2X1_LOC_496/a_36_24# OR2X1_LOC_778/A AND2X1_LOC_496/a_8_24# VSS VDD AND2X1_LOC_18/Y AND2X1_LOC_56/B AND2X1_LOC

XAND2X1_LOC_432 AND2X1_LOC_432/a_36_24# OR2X1_LOC_435/B AND2X1_LOC_432/a_8_24# VSS VDD AND2X1_LOC_18/Y OR2X1_LOC_130/A AND2X1_LOC

XAND2X1_LOC_607 AND2X1_LOC_607/a_36_24# OR2X1_LOC_646/B AND2X1_LOC_607/a_8_24# VSS VDD AND2X1_LOC_18/Y OR2X1_LOC_606/Y AND2X1_LOC

XAND2X1_LOC_754 AND2X1_LOC_754/a_36_24# OR2X1_LOC_790/A AND2X1_LOC_754/a_8_24# VSS VDD AND2X1_LOC_36/Y OR2X1_LOC_614/Y AND2X1_LOC

XAND2X1_LOC_320 AND2X1_LOC_320/a_36_24# OR2X1_LOC_324/B AND2X1_LOC_320/a_8_24# VSS VDD AND2X1_LOC_36/Y AND2X1_LOC_91/B AND2X1_LOC

XAND2X1_LOC_146 AND2X1_LOC_146/a_36_24# OR2X1_LOC_148/A AND2X1_LOC_146/a_8_24# VSS VDD AND2X1_LOC_36/Y OR2X1_LOC_160/A AND2X1_LOC

XAND2X1_LOC_39 AND2X1_LOC_39/a_36_24# AND2X1_LOC_39/Y AND2X1_LOC_39/a_8_24# VSS VDD AND2X1_LOC_36/Y OR2X1_LOC_154/A AND2X1_LOC

XAND2X1_LOC_495 AND2X1_LOC_495/a_36_24# OR2X1_LOC_499/B AND2X1_LOC_495/a_8_24# VSS VDD AND2X1_LOC_36/Y AND2X1_LOC_56/B AND2X1_LOC

XAND2X1_LOC_746 AND2X1_LOC_746/a_36_24# OR2X1_LOC_781/A AND2X1_LOC_746/a_8_24# VSS VDD OR2X1_LOC_185/A OR2X1_LOC_375/A AND2X1_LOC

XAND2X1_LOC_178 AND2X1_LOC_178/a_36_24# OR2X1_LOC_181/B AND2X1_LOC_178/a_8_24# VSS VDD AND2X1_LOC_56/B OR2X1_LOC_375/A AND2X1_LOC

XAND2X1_LOC_158 AND2X1_LOC_158/a_36_24# OR2X1_LOC_210/B AND2X1_LOC_158/a_8_24# VSS VDD OR2X1_LOC_156/Y OR2X1_LOC_375/A AND2X1_LOC

XAND2X1_LOC_282 AND2X1_LOC_282/a_36_24# OR2X1_LOC_285/A AND2X1_LOC_282/a_8_24# VSS VDD OR2X1_LOC_532/B OR2X1_LOC_375/A AND2X1_LOC

XAND2X1_LOC_416 AND2X1_LOC_416/a_36_24# OR2X1_LOC_462/B AND2X1_LOC_416/a_8_24# VSS VDD OR2X1_LOC_375/A OR2X1_LOC_415/Y AND2X1_LOC

XAND2X1_LOC_258 AND2X1_LOC_258/a_36_24# OR2X1_LOC_259/A AND2X1_LOC_258/a_8_24# VSS VDD OR2X1_LOC_78/A OR2X1_LOC_375/A AND2X1_LOC

XOR2X1_LOC_314 OR2X1_LOC_314/a_8_216# OR2X1_LOC_314/a_36_216# OR2X1_LOC_314/Y VSS VDD OR2X1_LOC_64/Y OR2X1_LOC_16/A OR2X1_LOC

XOR2X1_LOC_518 OR2X1_LOC_518/a_8_216# OR2X1_LOC_518/a_36_216# OR2X1_LOC_518/Y VSS VDD OR2X1_LOC_74/A OR2X1_LOC_64/Y OR2X1_LOC

XOR2X1_LOC_167 OR2X1_LOC_167/a_8_216# OR2X1_LOC_167/a_36_216# OR2X1_LOC_167/Y VSS VDD OR2X1_LOC_604/A OR2X1_LOC_64/Y OR2X1_LOC

XOR2X1_LOC_107 OR2X1_LOC_107/a_8_216# OR2X1_LOC_107/a_36_216# OR2X1_LOC_107/Y VSS VDD OR2X1_LOC_89/A OR2X1_LOC_64/Y OR2X1_LOC

XOR2X1_LOC_667 OR2X1_LOC_667/a_8_216# OR2X1_LOC_667/a_36_216# OR2X1_LOC_667/Y VSS VDD OR2X1_LOC_517/A OR2X1_LOC_64/Y OR2X1_LOC

XOR2X1_LOC_250 OR2X1_LOC_250/a_8_216# OR2X1_LOC_250/a_36_216# OR2X1_LOC_250/Y VSS VDD OR2X1_LOC_595/A OR2X1_LOC_64/Y OR2X1_LOC

XOR2X1_LOC_829 OR2X1_LOC_829/a_8_216# OR2X1_LOC_829/a_36_216# OR2X1_LOC_829/Y VSS VDD OR2X1_LOC_829/A OR2X1_LOC_64/Y OR2X1_LOC

XOR2X1_LOC_591 OR2X1_LOC_591/a_8_216# OR2X1_LOC_591/a_36_216# OR2X1_LOC_591/Y VSS VDD OR2X1_LOC_591/A OR2X1_LOC_64/Y OR2X1_LOC

XOR2X1_LOC_321 OR2X1_LOC_321/a_8_216# OR2X1_LOC_321/a_36_216# OR2X1_LOC_321/Y VSS VDD OR2X1_LOC_64/Y OR2X1_LOC_13/B OR2X1_LOC

XOR2X1_LOC_503 OR2X1_LOC_503/a_8_216# OR2X1_LOC_503/a_36_216# OR2X1_LOC_503/Y VSS VDD OR2X1_LOC_503/A OR2X1_LOC_64/Y OR2X1_LOC

XOR2X1_LOC_142 OR2X1_LOC_142/a_8_216# OR2X1_LOC_142/a_36_216# OR2X1_LOC_142/Y VSS VDD OR2X1_LOC_64/Y OR2X1_LOC_52/B OR2X1_LOC

XOR2X1_LOC_189 OR2X1_LOC_189/a_8_216# OR2X1_LOC_189/a_36_216# OR2X1_LOC_189/Y VSS VDD OR2X1_LOC_189/A OR2X1_LOC_95/Y OR2X1_LOC

XAND2X1_LOC_758 AND2X1_LOC_758/a_36_24# OR2X1_LOC_759/A AND2X1_LOC_758/a_8_24# VSS VDD OR2X1_LOC_40/Y OR2X1_LOC_95/Y AND2X1_LOC

XOR2X1_LOC_487 OR2X1_LOC_487/a_8_216# OR2X1_LOC_487/a_36_216# OR2X1_LOC_487/Y VSS VDD OR2X1_LOC_95/Y OR2X1_LOC_45/B OR2X1_LOC

XOR2X1_LOC_626 OR2X1_LOC_626/a_8_216# OR2X1_LOC_626/a_36_216# OR2X1_LOC_626/Y VSS VDD OR2X1_LOC_604/A OR2X1_LOC_95/Y OR2X1_LOC

XOR2X1_LOC_406 OR2X1_LOC_406/a_8_216# OR2X1_LOC_406/a_36_216# OR2X1_LOC_406/Y VSS VDD OR2X1_LOC_406/A OR2X1_LOC_95/Y OR2X1_LOC

XOR2X1_LOC_96 OR2X1_LOC_96/a_8_216# OR2X1_LOC_96/a_36_216# OR2X1_LOC_96/Y VSS VDD OR2X1_LOC_95/Y OR2X1_LOC_96/B OR2X1_LOC

XOR2X1_LOC_594 OR2X1_LOC_594/a_8_216# OR2X1_LOC_594/a_36_216# OR2X1_LOC_594/Y VSS VDD OR2X1_LOC_680/A OR2X1_LOC_95/Y OR2X1_LOC

XOR2X1_LOC_533 OR2X1_LOC_533/a_8_216# OR2X1_LOC_533/a_36_216# OR2X1_LOC_533/Y VSS VDD OR2X1_LOC_533/A OR2X1_LOC_95/Y OR2X1_LOC

XOR2X1_LOC_165 OR2X1_LOC_165/a_8_216# OR2X1_LOC_165/a_36_216# OR2X1_LOC_165/Y VSS VDD OR2X1_LOC_74/A OR2X1_LOC_51/Y OR2X1_LOC

XOR2X1_LOC_145 OR2X1_LOC_145/a_8_216# OR2X1_LOC_145/a_36_216# OR2X1_LOC_145/Y VSS VDD OR2X1_LOC_89/A OR2X1_LOC_51/Y OR2X1_LOC

XOR2X1_LOC_680 OR2X1_LOC_680/a_8_216# OR2X1_LOC_680/a_36_216# OR2X1_LOC_680/Y VSS VDD OR2X1_LOC_680/A OR2X1_LOC_51/Y OR2X1_LOC

XAND2X1_LOC_330 AND2X1_LOC_330/a_36_24# OR2X1_LOC_331/A AND2X1_LOC_330/a_8_24# VSS VDD OR2X1_LOC_51/Y OR2X1_LOC_70/Y AND2X1_LOC

XOR2X1_LOC_816 OR2X1_LOC_816/a_8_216# OR2X1_LOC_816/a_36_216# OR2X1_LOC_816/Y VSS VDD OR2X1_LOC_816/A OR2X1_LOC_51/Y OR2X1_LOC

XOR2X1_LOC_251 OR2X1_LOC_251/a_8_216# OR2X1_LOC_251/a_36_216# OR2X1_LOC_251/Y VSS VDD OR2X1_LOC_106/A OR2X1_LOC_51/Y OR2X1_LOC

XOR2X1_LOC_418 OR2X1_LOC_418/a_8_216# OR2X1_LOC_418/a_36_216# OR2X1_LOC_418/Y VSS VDD OR2X1_LOC_51/Y OR2X1_LOC_16/A OR2X1_LOC

XOR2X1_LOC_52 OR2X1_LOC_52/a_8_216# OR2X1_LOC_52/a_36_216# OR2X1_LOC_52/Y VSS VDD OR2X1_LOC_51/Y OR2X1_LOC_52/B OR2X1_LOC

XOR2X1_LOC_238 OR2X1_LOC_238/a_8_216# OR2X1_LOC_238/a_36_216# OR2X1_LOC_238/Y VSS VDD OR2X1_LOC_51/Y OR2X1_LOC_45/B OR2X1_LOC

XOR2X1_LOC_525 OR2X1_LOC_525/a_8_216# OR2X1_LOC_525/a_36_216# OR2X1_LOC_525/Y VSS VDD OR2X1_LOC_51/Y OR2X1_LOC_13/B OR2X1_LOC

XOR2X1_LOC_163 OR2X1_LOC_163/a_8_216# OR2X1_LOC_163/a_36_216# OR2X1_LOC_163/Y VSS VDD OR2X1_LOC_163/A OR2X1_LOC_51/Y OR2X1_LOC

XAND2X1_LOC_451 AND2X1_LOC_451/a_36_24# AND2X1_LOC_451/Y AND2X1_LOC_451/a_8_24# VSS VDD OR2X1_LOC_428/Y OR2X1_LOC_430/Y AND2X1_LOC

XAND2X1_LOC_460 AND2X1_LOC_460/a_36_24# AND2X1_LOC_463/B AND2X1_LOC_460/a_8_24# VSS VDD OR2X1_LOC_380/Y OR2X1_LOC_409/Y AND2X1_LOC

XOR2X1_LOC_769 OR2X1_LOC_769/a_8_216# OR2X1_LOC_769/a_36_216# OR2X1_LOC_771/B VSS VDD OR2X1_LOC_769/A OR2X1_LOC_769/B OR2X1_LOC

XOR2X1_LOC_635 OR2X1_LOC_635/a_8_216# OR2X1_LOC_635/a_36_216# OR2X1_LOC_639/B VSS VDD OR2X1_LOC_635/A OR2X1_LOC_451/B OR2X1_LOC

XOR2X1_LOC_790 OR2X1_LOC_790/a_8_216# OR2X1_LOC_790/a_36_216# OR2X1_LOC_793/A VSS VDD OR2X1_LOC_790/A OR2X1_LOC_790/B OR2X1_LOC

XAND2X1_LOC_394 AND2X1_LOC_394/a_36_24# OR2X1_LOC_400/A AND2X1_LOC_394/a_8_24# VSS VDD AND2X1_LOC_47/Y OR2X1_LOC_160/A AND2X1_LOC

XAND2X1_LOC_152 AND2X1_LOC_152/a_36_24# OR2X1_LOC_209/A AND2X1_LOC_152/a_8_24# VSS VDD AND2X1_LOC_47/Y OR2X1_LOC_151/Y AND2X1_LOC

XAND2X1_LOC_103 AND2X1_LOC_103/a_36_24# OR2X1_LOC_113/B AND2X1_LOC_103/a_8_24# VSS VDD AND2X1_LOC_47/Y OR2X1_LOC_532/B AND2X1_LOC

XAND2X1_LOC_106 AND2X1_LOC_106/a_36_24# OR2X1_LOC_115/B AND2X1_LOC_106/a_8_24# VSS VDD AND2X1_LOC_47/Y OR2X1_LOC_105/Y AND2X1_LOC

XAND2X1_LOC_248 AND2X1_LOC_248/a_36_24# OR2X1_LOC_342/A AND2X1_LOC_248/a_8_24# VSS VDD AND2X1_LOC_47/Y OR2X1_LOC_247/Y AND2X1_LOC

XAND2X1_LOC_744 AND2X1_LOC_744/a_36_24# OR2X1_LOC_780/A AND2X1_LOC_744/a_8_24# VSS VDD AND2X1_LOC_44/Y OR2X1_LOC_160/A AND2X1_LOC

XAND2X1_LOC_757 AND2X1_LOC_757/a_36_24# OR2X1_LOC_791/A AND2X1_LOC_757/a_8_24# VSS VDD AND2X1_LOC_44/Y OR2X1_LOC_756/Y AND2X1_LOC

XAND2X1_LOC_399 AND2X1_LOC_399/a_36_24# OR2X1_LOC_403/B AND2X1_LOC_399/a_8_24# VSS VDD AND2X1_LOC_44/Y OR2X1_LOC_398/Y AND2X1_LOC

XAND2X1_LOC_122 AND2X1_LOC_122/a_36_24# OR2X1_LOC_124/B AND2X1_LOC_122/a_8_24# VSS VDD AND2X1_LOC_44/Y OR2X1_LOC_121/Y AND2X1_LOC

XAND2X1_LOC_485 AND2X1_LOC_485/a_36_24# OR2X1_LOC_705/B AND2X1_LOC_485/a_8_24# VSS VDD AND2X1_LOC_44/Y OR2X1_LOC_532/B AND2X1_LOC

XAND2X1_LOC_297 AND2X1_LOC_297/a_36_24# OR2X1_LOC_347/B AND2X1_LOC_297/a_8_24# VSS VDD AND2X1_LOC_44/Y OR2X1_LOC_296/Y AND2X1_LOC

XAND2X1_LOC_424 AND2X1_LOC_424/a_36_24# OR2X1_LOC_449/A AND2X1_LOC_424/a_8_24# VSS VDD AND2X1_LOC_44/Y OR2X1_LOC_78/A AND2X1_LOC

XAND2X1_LOC_74 AND2X1_LOC_74/a_36_24# OR2X1_LOC_76/B AND2X1_LOC_74/a_8_24# VSS VDD AND2X1_LOC_31/Y OR2X1_LOC_185/A AND2X1_LOC

XAND2X1_LOC_517 AND2X1_LOC_517/a_36_24# OR2X1_LOC_559/B AND2X1_LOC_517/a_8_24# VSS VDD AND2X1_LOC_31/Y OR2X1_LOC_264/Y AND2X1_LOC

XAND2X1_LOC_491 AND2X1_LOC_491/a_36_24# OR2X1_LOC_493/B AND2X1_LOC_491/a_8_24# VSS VDD AND2X1_LOC_31/Y OR2X1_LOC_532/B AND2X1_LOC

XAND2X1_LOC_109 AND2X1_LOC_109/a_36_24# OR2X1_LOC_112/B AND2X1_LOC_109/a_8_24# VSS VDD AND2X1_LOC_31/Y OR2X1_LOC_78/A AND2X1_LOC

XAND2X1_LOC_298 AND2X1_LOC_298/a_36_24# OR2X1_LOC_302/B AND2X1_LOC_298/a_8_24# VSS VDD AND2X1_LOC_31/Y AND2X1_LOC_56/B AND2X1_LOC

XAND2X1_LOC_224 AND2X1_LOC_224/a_36_24# OR2X1_LOC_227/B AND2X1_LOC_224/a_8_24# VSS VDD AND2X1_LOC_31/Y OR2X1_LOC_160/A AND2X1_LOC

XAND2X1_LOC_91 AND2X1_LOC_91/a_36_24# OR2X1_LOC_97/A AND2X1_LOC_91/a_8_24# VSS VDD AND2X1_LOC_51/Y AND2X1_LOC_91/B AND2X1_LOC

XAND2X1_LOC_163 AND2X1_LOC_163/a_36_24# OR2X1_LOC_467/B AND2X1_LOC_163/a_8_24# VSS VDD AND2X1_LOC_51/Y OR2X1_LOC_162/Y AND2X1_LOC

XAND2X1_LOC_165 AND2X1_LOC_165/a_36_24# OR2X1_LOC_168/A AND2X1_LOC_165/a_8_24# VSS VDD AND2X1_LOC_51/Y OR2X1_LOC_185/A AND2X1_LOC

XAND2X1_LOC_145 AND2X1_LOC_145/a_36_24# OR2X1_LOC_148/B AND2X1_LOC_145/a_8_24# VSS VDD AND2X1_LOC_51/Y OR2X1_LOC_78/A AND2X1_LOC

XAND2X1_LOC_680 AND2X1_LOC_680/a_36_24# OR2X1_LOC_728/A AND2X1_LOC_680/a_8_24# VSS VDD AND2X1_LOC_51/Y OR2X1_LOC_186/Y AND2X1_LOC

XAND2X1_LOC_816 AND2X1_LOC_816/a_36_24# OR2X1_LOC_846/A AND2X1_LOC_816/a_8_24# VSS VDD AND2X1_LOC_51/Y OR2X1_LOC_185/Y AND2X1_LOC

XAND2X1_LOC_251 AND2X1_LOC_251/a_36_24# OR2X1_LOC_843/B AND2X1_LOC_251/a_8_24# VSS VDD AND2X1_LOC_51/Y OR2X1_LOC_105/Y AND2X1_LOC

XAND2X1_LOC_617 AND2X1_LOC_617/a_36_24# OR2X1_LOC_621/A AND2X1_LOC_617/a_8_24# VSS VDD OR2X1_LOC_154/A AND2X1_LOC_51/Y AND2X1_LOC

XAND2X1_LOC_239 AND2X1_LOC_239/a_36_24# OR2X1_LOC_506/B AND2X1_LOC_239/a_8_24# VSS VDD AND2X1_LOC_51/Y OR2X1_LOC_532/B AND2X1_LOC

XAND2X1_LOC_450 AND2X1_LOC_450/a_36_24# AND2X1_LOC_450/Y AND2X1_LOC_450/a_8_24# VSS VDD OR2X1_LOC_426/Y OR2X1_LOC_427/Y AND2X1_LOC

XAND2X1_LOC_707 AND2X1_LOC_707/a_36_24# AND2X1_LOC_707/Y AND2X1_LOC_707/a_8_24# VSS VDD OR2X1_LOC_694/Y OR2X1_LOC_695/Y AND2X1_LOC

XOR2X1_LOC_187 OR2X1_LOC_187/a_8_216# OR2X1_LOC_187/a_36_216# OR2X1_LOC_187/Y VSS VDD OR2X1_LOC_680/A OR2X1_LOC_40/Y OR2X1_LOC

XOR2X1_LOC_166 OR2X1_LOC_166/a_8_216# OR2X1_LOC_166/a_36_216# OR2X1_LOC_166/Y VSS VDD OR2X1_LOC_40/Y OR2X1_LOC_16/A OR2X1_LOC

XOR2X1_LOC_441 OR2X1_LOC_441/a_8_216# OR2X1_LOC_441/a_36_216# OR2X1_LOC_441/Y VSS VDD OR2X1_LOC_52/B OR2X1_LOC_40/Y OR2X1_LOC

XOR2X1_LOC_265 OR2X1_LOC_265/a_8_216# OR2X1_LOC_265/a_36_216# OR2X1_LOC_265/Y VSS VDD OR2X1_LOC_517/A OR2X1_LOC_40/Y OR2X1_LOC

XOR2X1_LOC_41 OR2X1_LOC_41/a_8_216# OR2X1_LOC_41/a_36_216# OR2X1_LOC_41/Y VSS VDD OR2X1_LOC_40/Y OR2X1_LOC_13/B OR2X1_LOC

XOR2X1_LOC_745 OR2X1_LOC_745/a_8_216# OR2X1_LOC_745/a_36_216# OR2X1_LOC_745/Y VSS VDD OR2X1_LOC_604/A OR2X1_LOC_40/Y OR2X1_LOC

XOR2X1_LOC_531 OR2X1_LOC_531/a_8_216# OR2X1_LOC_531/a_36_216# OR2X1_LOC_531/Y VSS VDD OR2X1_LOC_74/A OR2X1_LOC_40/Y OR2X1_LOC

XOR2X1_LOC_384 OR2X1_LOC_384/a_8_216# OR2X1_LOC_384/a_36_216# OR2X1_LOC_384/Y VSS VDD OR2X1_LOC_494/A OR2X1_LOC_40/Y OR2X1_LOC

XOR2X1_LOC_171 OR2X1_LOC_171/a_8_216# OR2X1_LOC_171/a_36_216# OR2X1_LOC_171/Y VSS VDD OR2X1_LOC_40/Y OR2X1_LOC_45/B OR2X1_LOC

XOR2X1_LOC_665 OR2X1_LOC_665/a_8_216# OR2X1_LOC_665/a_36_216# OR2X1_LOC_665/Y VSS VDD OR2X1_LOC_755/A OR2X1_LOC_3/Y OR2X1_LOC

XOR2X1_LOC_815 OR2X1_LOC_815/a_8_216# OR2X1_LOC_815/a_36_216# OR2X1_LOC_815/Y VSS VDD OR2X1_LOC_815/A OR2X1_LOC_3/Y OR2X1_LOC

XOR2X1_LOC_751 OR2X1_LOC_751/a_8_216# OR2X1_LOC_751/a_36_216# OR2X1_LOC_751/Y VSS VDD OR2X1_LOC_751/A OR2X1_LOC_3/Y OR2X1_LOC

XOR2X1_LOC_767 OR2X1_LOC_767/a_8_216# OR2X1_LOC_767/a_36_216# OR2X1_LOC_767/Y VSS VDD OR2X1_LOC_79/A OR2X1_LOC_3/Y OR2X1_LOC

XOR2X1_LOC_16 OR2X1_LOC_16/a_8_216# OR2X1_LOC_16/a_36_216# OR2X1_LOC_16/Y VSS VDD OR2X1_LOC_16/A OR2X1_LOC_3/Y OR2X1_LOC

XOR2X1_LOC_397 OR2X1_LOC_397/a_8_216# OR2X1_LOC_397/a_36_216# OR2X1_LOC_397/Y VSS VDD OR2X1_LOC_83/A OR2X1_LOC_3/Y OR2X1_LOC

XOR2X1_LOC_177 OR2X1_LOC_177/a_8_216# OR2X1_LOC_177/a_36_216# OR2X1_LOC_177/Y VSS VDD OR2X1_LOC_70/Y OR2X1_LOC_52/B OR2X1_LOC

XOR2X1_LOC_821 OR2X1_LOC_821/a_8_216# OR2X1_LOC_821/a_36_216# OR2X1_LOC_821/Y VSS VDD OR2X1_LOC_70/Y OR2X1_LOC_13/B OR2X1_LOC

XOR2X1_LOC_118 OR2X1_LOC_118/a_8_216# OR2X1_LOC_118/a_36_216# OR2X1_LOC_118/Y VSS VDD OR2X1_LOC_89/A OR2X1_LOC_70/Y OR2X1_LOC

XOR2X1_LOC_674 OR2X1_LOC_674/a_8_216# OR2X1_LOC_674/a_36_216# OR2X1_LOC_674/Y VSS VDD OR2X1_LOC_329/B OR2X1_LOC_70/Y OR2X1_LOC

XOR2X1_LOC_498 OR2X1_LOC_498/a_8_216# OR2X1_LOC_498/a_36_216# OR2X1_LOC_498/Y VSS VDD OR2X1_LOC_189/A OR2X1_LOC_70/Y OR2X1_LOC

XOR2X1_LOC_604 OR2X1_LOC_604/a_8_216# OR2X1_LOC_604/a_36_216# OR2X1_LOC_604/Y VSS VDD OR2X1_LOC_604/A OR2X1_LOC_70/Y OR2X1_LOC

XOR2X1_LOC_438 OR2X1_LOC_438/a_8_216# OR2X1_LOC_438/a_36_216# OR2X1_LOC_438/Y VSS VDD OR2X1_LOC_70/Y OR2X1_LOC_45/B OR2X1_LOC

XOR2X1_LOC_158 OR2X1_LOC_158/a_8_216# OR2X1_LOC_158/a_36_216# OR2X1_LOC_158/Y VSS VDD OR2X1_LOC_158/A OR2X1_LOC_158/B OR2X1_LOC

XOR2X1_LOC_232 OR2X1_LOC_232/a_8_216# OR2X1_LOC_232/a_36_216# OR2X1_LOC_232/Y VSS VDD OR2X1_LOC_158/A OR2X1_LOC_16/A OR2X1_LOC

XOR2X1_LOC_258 OR2X1_LOC_258/a_8_216# OR2X1_LOC_258/a_36_216# OR2X1_LOC_258/Y VSS VDD OR2X1_LOC_158/A OR2X1_LOC_89/A OR2X1_LOC

XOR2X1_LOC_746 OR2X1_LOC_746/a_8_216# OR2X1_LOC_746/a_36_216# OR2X1_LOC_746/Y VSS VDD OR2X1_LOC_158/A OR2X1_LOC_74/A OR2X1_LOC

XOR2X1_LOC_504 OR2X1_LOC_504/a_8_216# OR2X1_LOC_504/a_36_216# OR2X1_LOC_504/Y VSS VDD OR2X1_LOC_158/A OR2X1_LOC_13/B OR2X1_LOC

XAND2X1_LOC_197 AND2X1_LOC_197/a_36_24# AND2X1_LOC_197/Y AND2X1_LOC_197/a_8_24# VSS VDD OR2X1_LOC_52/Y OR2X1_LOC_56/Y AND2X1_LOC

XAND2X1_LOC_307 AND2X1_LOC_307/a_36_24# AND2X1_LOC_307/Y AND2X1_LOC_307/a_8_24# VSS VDD OR2X1_LOC_304/Y OR2X1_LOC_305/Y AND2X1_LOC

XAND2X1_LOC_355 AND2X1_LOC_355/a_36_24# AND2X1_LOC_356/B AND2X1_LOC_355/a_8_24# VSS VDD OR2X1_LOC_329/Y OR2X1_LOC_331/Y AND2X1_LOC

XOR2X1_LOC_597 OR2X1_LOC_597/a_8_216# OR2X1_LOC_597/a_36_216# OR2X1_LOC_597/Y VSS VDD OR2X1_LOC_597/A OR2X1_LOC_13/B OR2X1_LOC

XAND2X1_LOC_389 AND2X1_LOC_389/a_36_24# AND2X1_LOC_390/B AND2X1_LOC_389/a_8_24# VSS VDD OR2X1_LOC_385/Y OR2X1_LOC_387/Y AND2X1_LOC

XOR2X1_LOC_391 OR2X1_LOC_391/a_8_216# OR2X1_LOC_391/a_36_216# OR2X1_LOC_392/A VSS VDD OR2X1_LOC_391/A OR2X1_LOC_391/B OR2X1_LOC

XOR2X1_LOC_549 OR2X1_LOC_549/a_8_216# OR2X1_LOC_549/a_36_216# OR2X1_LOC_549/Y VSS VDD OR2X1_LOC_549/A OR2X1_LOC_549/B OR2X1_LOC

XOR2X1_LOC_777 OR2X1_LOC_777/a_8_216# OR2X1_LOC_777/a_36_216# OR2X1_LOC_784/B VSS VDD OR2X1_LOC_307/A OR2X1_LOC_777/B OR2X1_LOC

XOR2X1_LOC_633 OR2X1_LOC_633/a_8_216# OR2X1_LOC_633/a_36_216# OR2X1_LOC_633/Y VSS VDD OR2X1_LOC_633/A OR2X1_LOC_633/B OR2X1_LOC

XOR2X1_LOC_541 OR2X1_LOC_541/a_8_216# OR2X1_LOC_541/a_36_216# OR2X1_LOC_553/A VSS VDD OR2X1_LOC_541/A OR2X1_LOC_541/B OR2X1_LOC

XOR2X1_LOC_634 OR2X1_LOC_634/a_8_216# OR2X1_LOC_634/a_36_216# OR2X1_LOC_640/A VSS VDD OR2X1_LOC_634/A OR2X1_LOC_334/B OR2X1_LOC

XOR2X1_LOC_266 OR2X1_LOC_266/a_8_216# OR2X1_LOC_266/a_36_216# OR2X1_LOC_267/A VSS VDD OR2X1_LOC_266/A OR2X1_LOC_786/A OR2X1_LOC

XAND2X1_LOC_813 AND2X1_LOC_813/a_36_24# OR2X1_LOC_845/A AND2X1_LOC_813/a_8_24# VSS VDD OR2X1_LOC_71/A OR2X1_LOC_266/A AND2X1_LOC

XOR2X1_LOC_188 OR2X1_LOC_188/a_8_216# OR2X1_LOC_188/a_36_216# OR2X1_LOC_188/Y VSS VDD OR2X1_LOC_185/Y OR2X1_LOC_154/A OR2X1_LOC

XOR2X1_LOC_590 OR2X1_LOC_590/a_8_216# OR2X1_LOC_590/a_36_216# OR2X1_LOC_590/Y VSS VDD OR2X1_LOC_532/B OR2X1_LOC_154/A OR2X1_LOC

XAND2X1_LOC_380 AND2X1_LOC_380/a_36_24# OR2X1_LOC_460/B AND2X1_LOC_380/a_8_24# VSS VDD OR2X1_LOC_160/A OR2X1_LOC_379/Y AND2X1_LOC

XOR2X1_LOC_532 OR2X1_LOC_532/a_8_216# OR2X1_LOC_532/a_36_216# OR2X1_LOC_532/Y VSS VDD OR2X1_LOC_160/A OR2X1_LOC_532/B OR2X1_LOC

XAND2X1_LOC_235 AND2X1_LOC_235/a_36_24# OR2X1_LOC_243/B AND2X1_LOC_235/a_8_24# VSS VDD OR2X1_LOC_71/A AND2X1_LOC_86/B AND2X1_LOC

XOR2X1_LOC_664 OR2X1_LOC_664/a_8_216# OR2X1_LOC_664/a_36_216# OR2X1_LOC_664/Y VSS VDD OR2X1_LOC_78/A OR2X1_LOC_185/A OR2X1_LOC

XOR2X1_LOC_151 OR2X1_LOC_151/a_8_216# OR2X1_LOC_151/a_36_216# OR2X1_LOC_151/Y VSS VDD OR2X1_LOC_151/A AND2X1_LOC_56/B OR2X1_LOC

XOR2X1_LOC_186 OR2X1_LOC_186/a_8_216# OR2X1_LOC_186/a_36_216# OR2X1_LOC_186/Y VSS VDD OR2X1_LOC_185/Y OR2X1_LOC_151/A OR2X1_LOC

XAND2X1_LOC_622 AND2X1_LOC_622/a_36_24# AND2X1_LOC_624/A AND2X1_LOC_622/a_8_24# VSS VDD OR2X1_LOC_619/Y AND2X1_LOC_621/Y AND2X1_LOC

XAND2X1_LOC_78 AND2X1_LOC_78/a_36_24# OR2X1_LOC_79/A AND2X1_LOC_78/a_8_24# VSS VDD OR2X1_LOC_16/A OR2X1_LOC_89/A AND2X1_LOC

XAND2X1_LOC_664 AND2X1_LOC_664/a_36_24# OR2X1_LOC_755/A AND2X1_LOC_664/a_8_24# VSS VDD OR2X1_LOC_74/A OR2X1_LOC_89/A AND2X1_LOC

XAND2X1_LOC_709 AND2X1_LOC_709/a_36_24# AND2X1_LOC_711/A AND2X1_LOC_709/a_8_24# VSS VDD OR2X1_LOC_698/Y OR2X1_LOC_748/A AND2X1_LOC

XAND2X1_LOC_706 AND2X1_LOC_706/a_36_24# AND2X1_LOC_706/Y AND2X1_LOC_706/a_8_24# VSS VDD OR2X1_LOC_692/Y OR2X1_LOC_693/Y AND2X1_LOC

XOR2X1_LOC_673 OR2X1_LOC_673/a_8_216# OR2X1_LOC_673/a_36_216# OR2X1_LOC_673/Y VSS VDD OR2X1_LOC_673/A OR2X1_LOC_673/B OR2X1_LOC

XAND2X1_LOC_776 AND2X1_LOC_776/a_36_24# AND2X1_LOC_776/Y AND2X1_LOC_776/a_8_24# VSS VDD OR2X1_LOC_164/Y OR2X1_LOC_238/Y AND2X1_LOC

XAND2X1_LOC_168 AND2X1_LOC_168/a_36_24# AND2X1_LOC_168/Y AND2X1_LOC_168/a_8_24# VSS VDD OR2X1_LOC_164/Y OR2X1_LOC_165/Y AND2X1_LOC

XAND2X1_LOC_325 AND2X1_LOC_325/a_36_24# AND2X1_LOC_326/B AND2X1_LOC_325/a_8_24# VSS VDD OR2X1_LOC_322/Y OR2X1_LOC_323/Y AND2X1_LOC

XAND2X1_LOC_459 AND2X1_LOC_459/a_36_24# AND2X1_LOC_459/Y AND2X1_LOC_459/a_8_24# VSS VDD OR2X1_LOC_376/Y OR2X1_LOC_378/Y AND2X1_LOC

XAND2X1_LOC_638 AND2X1_LOC_638/a_36_24# AND2X1_LOC_638/Y AND2X1_LOC_638/a_8_24# VSS VDD OR2X1_LOC_588/Y AND2X1_LOC_637/Y AND2X1_LOC

XAND2X1_LOC_708 AND2X1_LOC_708/a_36_24# AND2X1_LOC_712/B AND2X1_LOC_708/a_8_24# VSS VDD OR2X1_LOC_696/Y OR2X1_LOC_697/Y AND2X1_LOC

XAND2X1_LOC_308 AND2X1_LOC_308/a_36_24# AND2X1_LOC_727/A AND2X1_LOC_308/a_8_24# VSS VDD OR2X1_LOC_306/Y AND2X1_LOC_307/Y AND2X1_LOC

XAND2X1_LOC_147 AND2X1_LOC_147/a_36_24# AND2X1_LOC_147/Y AND2X1_LOC_147/a_8_24# VSS VDD OR2X1_LOC_142/Y OR2X1_LOC_144/Y AND2X1_LOC

XOR2X1_LOC_630 OR2X1_LOC_630/a_8_216# OR2X1_LOC_630/a_36_216# OR2X1_LOC_630/Y VSS VDD OR2X1_LOC_629/Y OR2X1_LOC_630/B OR2X1_LOC

XOR2X1_LOC_389 OR2X1_LOC_389/a_8_216# OR2X1_LOC_389/a_36_216# OR2X1_LOC_390/A VSS VDD OR2X1_LOC_389/A OR2X1_LOC_389/B OR2X1_LOC

XOR2X1_LOC_98 OR2X1_LOC_98/a_8_216# OR2X1_LOC_98/a_36_216# OR2X1_LOC_99/A VSS VDD OR2X1_LOC_98/A OR2X1_LOC_98/B OR2X1_LOC

XOR2X1_LOC_506 OR2X1_LOC_506/a_8_216# OR2X1_LOC_506/a_36_216# OR2X1_LOC_506/Y VSS VDD OR2X1_LOC_506/A OR2X1_LOC_506/B OR2X1_LOC

XOR2X1_LOC_447 OR2X1_LOC_447/a_8_216# OR2X1_LOC_447/a_36_216# OR2X1_LOC_447/Y VSS VDD OR2X1_LOC_447/A OR2X1_LOC_506/A OR2X1_LOC

XOR2X1_LOC_838 OR2X1_LOC_838/a_8_216# OR2X1_LOC_838/a_36_216# OR2X1_LOC_852/B VSS VDD OR2X1_LOC_837/Y OR2X1_LOC_838/B OR2X1_LOC

XOR2X1_LOC_138 OR2X1_LOC_138/a_8_216# OR2X1_LOC_138/a_36_216# OR2X1_LOC_139/A VSS VDD OR2X1_LOC_138/A OR2X1_LOC_702/A OR2X1_LOC

XOR2X1_LOC_195 OR2X1_LOC_195/a_8_216# OR2X1_LOC_195/a_36_216# OR2X1_LOC_199/B VSS VDD OR2X1_LOC_195/A AND2X1_LOC_41/Y OR2X1_LOC

XOR2X1_LOC_535 OR2X1_LOC_535/a_8_216# OR2X1_LOC_535/a_36_216# OR2X1_LOC_854/A VSS VDD OR2X1_LOC_535/A OR2X1_LOC_788/B OR2X1_LOC

XAND2X1_LOC_67 AND2X1_LOC_67/a_36_24# AND2X1_LOC_67/Y AND2X1_LOC_67/a_8_24# VSS VDD AND2X1_LOC_56/B OR2X1_LOC_66/Y AND2X1_LOC

XOR2X1_LOC_612 OR2X1_LOC_612/a_8_216# OR2X1_LOC_612/a_36_216# OR2X1_LOC_612/Y VSS VDD OR2X1_LOC_611/Y OR2X1_LOC_612/B OR2X1_LOC

XAND2X1_LOC_848 AND2X1_LOC_848/a_36_24# AND2X1_LOC_848/Y AND2X1_LOC_848/a_8_24# VSS VDD AND2X1_LOC_848/A AND2X1_LOC_847/Y AND2X1_LOC

XOR2X1_LOC_450 OR2X1_LOC_450/a_8_216# OR2X1_LOC_450/a_36_216# OR2X1_LOC_450/Y VSS VDD OR2X1_LOC_450/A OR2X1_LOC_450/B OR2X1_LOC

XOR2X1_LOC_302 OR2X1_LOC_302/a_8_216# OR2X1_LOC_302/a_36_216# OR2X1_LOC_303/A VSS VDD OR2X1_LOC_302/A OR2X1_LOC_302/B OR2X1_LOC

XOR2X1_LOC_543 OR2X1_LOC_543/a_8_216# OR2X1_LOC_543/a_36_216# OR2X1_LOC_552/A VSS VDD OR2X1_LOC_543/A OR2X1_LOC_318/B OR2X1_LOC

XOR2X1_LOC_301 OR2X1_LOC_301/a_8_216# OR2X1_LOC_301/a_36_216# OR2X1_LOC_303/B VSS VDD OR2X1_LOC_831/A OR2X1_LOC_76/A OR2X1_LOC

XAND2X1_LOC_227 AND2X1_LOC_227/a_36_24# AND2X1_LOC_227/Y AND2X1_LOC_227/a_8_24# VSS VDD OR2X1_LOC_224/Y OR2X1_LOC_226/Y AND2X1_LOC

XAND2X1_LOC_704 AND2X1_LOC_704/a_36_24# AND2X1_LOC_714/B AND2X1_LOC_704/a_8_24# VSS VDD OR2X1_LOC_313/Y OR2X1_LOC_417/Y AND2X1_LOC

XAND2X1_LOC_446 AND2X1_LOC_446/a_36_24# AND2X1_LOC_454/A AND2X1_LOC_446/a_8_24# VSS VDD OR2X1_LOC_417/Y OR2X1_LOC_418/Y AND2X1_LOC

XAND2X1_LOC_333 AND2X1_LOC_333/a_36_24# AND2X1_LOC_338/A AND2X1_LOC_333/a_8_24# VSS VDD OR2X1_LOC_171/Y OR2X1_LOC_289/Y AND2X1_LOC

XAND2X1_LOC_489 AND2X1_LOC_489/a_36_24# AND2X1_LOC_489/Y AND2X1_LOC_489/a_8_24# VSS VDD OR2X1_LOC_487/Y OR2X1_LOC_488/Y AND2X1_LOC

XAND2X1_LOC_286 AND2X1_LOC_286/a_36_24# AND2X1_LOC_286/Y AND2X1_LOC_286/a_8_24# VSS VDD OR2X1_LOC_283/Y AND2X1_LOC_285/Y AND2X1_LOC

XOR2X1_LOC_631 OR2X1_LOC_631/a_8_216# OR2X1_LOC_631/a_36_216# OR2X1_LOC_632/A VSS VDD OR2X1_LOC_631/A OR2X1_LOC_631/B OR2X1_LOC

XOR2X1_LOC_637 OR2X1_LOC_637/a_8_216# OR2X1_LOC_637/a_36_216# OR2X1_LOC_637/Y VSS VDD OR2X1_LOC_637/A OR2X1_LOC_637/B OR2X1_LOC

XOR2X1_LOC_843 OR2X1_LOC_843/a_8_216# OR2X1_LOC_843/a_36_216# OR2X1_LOC_850/A VSS VDD OR2X1_LOC_287/B OR2X1_LOC_843/B OR2X1_LOC

XOR2X1_LOC_287 OR2X1_LOC_287/a_8_216# OR2X1_LOC_287/a_36_216# OR2X1_LOC_288/A VSS VDD OR2X1_LOC_287/A OR2X1_LOC_287/B OR2X1_LOC

XAND2X1_LOC_608 AND2X1_LOC_608/a_36_24# OR2X1_LOC_609/A AND2X1_LOC_608/a_8_24# VSS VDD OR2X1_LOC_16/A OR2X1_LOC_74/A AND2X1_LOC

XAND2X1_LOC_342 AND2X1_LOC_342/a_36_24# AND2X1_LOC_342/Y AND2X1_LOC_342/a_8_24# VSS VDD OR2X1_LOC_246/Y OR2X1_LOC_248/Y AND2X1_LOC

XOR2X1_LOC_669 OR2X1_LOC_669/a_8_216# OR2X1_LOC_669/a_36_216# OR2X1_LOC_669/Y VSS VDD OR2X1_LOC_669/A OR2X1_LOC_604/A OR2X1_LOC

XAND2X1_LOC_779 AND2X1_LOC_779/a_36_24# AND2X1_LOC_779/Y AND2X1_LOC_779/a_8_24# VSS VDD OR2X1_LOC_511/Y OR2X1_LOC_697/Y AND2X1_LOC

XAND2X1_LOC_834 AND2X1_LOC_834/a_36_24# AND2X1_LOC_840/B AND2X1_LOC_834/a_8_24# VSS VDD OR2X1_LOC_511/Y OR2X1_LOC_677/Y AND2X1_LOC

XAND2X1_LOC_196 AND2X1_LOC_196/a_36_24# AND2X1_LOC_196/Y AND2X1_LOC_196/a_8_24# VSS VDD OR2X1_LOC_45/Y OR2X1_LOC_48/Y AND2X1_LOC

XAND2X1_LOC_769 AND2X1_LOC_769/a_36_24# AND2X1_LOC_769/Y AND2X1_LOC_769/a_8_24# VSS VDD OR2X1_LOC_763/Y OR2X1_LOC_764/Y AND2X1_LOC

XAND2X1_LOC_828 AND2X1_LOC_828/a_36_24# OR2X1_LOC_829/A AND2X1_LOC_828/a_8_24# VSS VDD OR2X1_LOC_409/B OR2X1_LOC_599/A AND2X1_LOC

XAND2X1_LOC_520 AND2X1_LOC_520/a_36_24# AND2X1_LOC_520/Y AND2X1_LOC_520/a_8_24# VSS VDD OR2X1_LOC_518/Y OR2X1_LOC_519/Y AND2X1_LOC

XAND2X1_LOC_464 AND2X1_LOC_464/a_36_24# AND2X1_LOC_464/Y AND2X1_LOC_464/a_8_24# VSS VDD AND2X1_LOC_464/A AND2X1_LOC_458/Y AND2X1_LOC

XAND2X1_LOC_780 AND2X1_LOC_780/a_36_24# AND2X1_LOC_783/B AND2X1_LOC_780/a_8_24# VSS VDD OR2X1_LOC_743/Y OR2X1_LOC_744/Y AND2X1_LOC

XAND2X1_LOC_832 AND2X1_LOC_832/a_36_24# AND2X1_LOC_841/B AND2X1_LOC_832/a_8_24# VSS VDD OR2X1_LOC_423/Y OR2X1_LOC_433/Y AND2X1_LOC

XAND2X1_LOC_435 AND2X1_LOC_435/a_36_24# AND2X1_LOC_436/B AND2X1_LOC_435/a_8_24# VSS VDD OR2X1_LOC_432/Y OR2X1_LOC_433/Y AND2X1_LOC

XAND2X1_LOC_156 AND2X1_LOC_156/a_36_24# OR2X1_LOC_158/B AND2X1_LOC_156/a_8_24# VSS VDD AND2X1_LOC_154/Y AND2X1_LOC_155/Y AND2X1_LOC

XAND2X1_LOC_332 AND2X1_LOC_332/a_36_24# AND2X1_LOC_339/B AND2X1_LOC_332/a_8_24# VSS VDD OR2X1_LOC_111/Y OR2X1_LOC_135/Y AND2X1_LOC

XAND2X1_LOC_112 AND2X1_LOC_112/a_36_24# AND2X1_LOC_715/A AND2X1_LOC_112/a_8_24# VSS VDD OR2X1_LOC_109/Y OR2X1_LOC_111/Y AND2X1_LOC

XAND2X1_LOC_547 AND2X1_LOC_547/a_36_24# AND2X1_LOC_547/Y AND2X1_LOC_547/a_8_24# VSS VDD OR2X1_LOC_527/Y OR2X1_LOC_528/Y AND2X1_LOC

XAND2X1_LOC_729 AND2X1_LOC_729/a_36_24# AND2X1_LOC_729/Y AND2X1_LOC_729/a_8_24# VSS VDD AND2X1_LOC_687/Y AND2X1_LOC_729/B AND2X1_LOC

XAND2X1_LOC_855 AND2X1_LOC_855/a_36_24# AND2X1_LOC_856/B AND2X1_LOC_855/a_8_24# VSS VDD AND2X1_LOC_729/B OR2X1_LOC_829/Y AND2X1_LOC

XOR2X1_LOC_101 OR2X1_LOC_101/a_8_216# OR2X1_LOC_101/a_36_216# OR2X1_LOC_656/B VSS VDD OR2X1_LOC_100/Y OR2X1_LOC_99/Y OR2X1_LOC

XAND2X1_LOC_361 AND2X1_LOC_361/a_36_24# AND2X1_LOC_362/B AND2X1_LOC_361/a_8_24# VSS VDD AND2X1_LOC_361/A AND2X1_LOC_276/Y AND2X1_LOC

XAND2X1_LOC_473 AND2X1_LOC_473/a_36_24# AND2X1_LOC_473/Y AND2X1_LOC_473/a_8_24# VSS VDD AND2X1_LOC_116/Y AND2X1_LOC_276/Y AND2X1_LOC

XAND2X1_LOC_809 AND2X1_LOC_809/a_36_24# AND2X1_LOC_810/B AND2X1_LOC_809/a_8_24# VSS VDD AND2X1_LOC_809/A AND2X1_LOC_802/Y AND2X1_LOC

XOR2X1_LOC_462 OR2X1_LOC_462/a_8_216# OR2X1_LOC_462/a_36_216# OR2X1_LOC_472/B VSS VDD OR2X1_LOC_461/Y OR2X1_LOC_462/B OR2X1_LOC

XOR2X1_LOC_240 OR2X1_LOC_240/a_8_216# OR2X1_LOC_240/a_36_216# OR2X1_LOC_243/A VSS VDD OR2X1_LOC_240/A OR2X1_LOC_240/B OR2X1_LOC

XOR2X1_LOC_836 OR2X1_LOC_836/a_8_216# OR2X1_LOC_836/a_36_216# OR2X1_LOC_836/Y VSS VDD OR2X1_LOC_836/A OR2X1_LOC_836/B OR2X1_LOC

XOR2X1_LOC_334 OR2X1_LOC_334/a_8_216# OR2X1_LOC_334/a_36_216# OR2X1_LOC_338/A VSS VDD OR2X1_LOC_334/A OR2X1_LOC_334/B OR2X1_LOC

XAND2X1_LOC_331 AND2X1_LOC_331/a_36_24# OR2X1_LOC_355/A AND2X1_LOC_331/a_8_24# VSS VDD OR2X1_LOC_186/Y OR2X1_LOC_330/Y AND2X1_LOC

XOR2X1_LOC_621 OR2X1_LOC_621/a_8_216# OR2X1_LOC_621/a_36_216# OR2X1_LOC_622/A VSS VDD OR2X1_LOC_621/A OR2X1_LOC_621/B OR2X1_LOC

XOR2X1_LOC_457 OR2X1_LOC_457/a_8_216# OR2X1_LOC_457/a_36_216# OR2X1_LOC_464/B VSS VDD OR2X1_LOC_787/B OR2X1_LOC_457/B OR2X1_LOC

XAND2X1_LOC_483 AND2X1_LOC_483/a_36_24# AND2X1_LOC_483/Y AND2X1_LOC_483/a_8_24# VSS VDD OR2X1_LOC_252/Y OR2X1_LOC_482/Y AND2X1_LOC

XAND2X1_LOC_629 AND2X1_LOC_629/a_36_24# AND2X1_LOC_629/Y AND2X1_LOC_629/a_8_24# VSS VDD OR2X1_LOC_626/Y OR2X1_LOC_627/Y AND2X1_LOC

XAND2X1_LOC_254 AND2X1_LOC_254/a_36_24# AND2X1_LOC_456/B AND2X1_LOC_254/a_8_24# VSS VDD OR2X1_LOC_252/Y OR2X1_LOC_253/Y AND2X1_LOC

XAND2X1_LOC_837 AND2X1_LOC_837/a_36_24# AND2X1_LOC_838/B AND2X1_LOC_837/a_8_24# VSS VDD OR2X1_LOC_825/Y OR2X1_LOC_826/Y AND2X1_LOC

XAND2X1_LOC_284 AND2X1_LOC_284/a_36_24# AND2X1_LOC_287/B AND2X1_LOC_284/a_8_24# VSS VDD OR2X1_LOC_279/Y OR2X1_LOC_280/Y AND2X1_LOC

XOR2X1_LOC_846 OR2X1_LOC_846/a_8_216# OR2X1_LOC_846/a_36_216# OR2X1_LOC_848/B VSS VDD OR2X1_LOC_846/A OR2X1_LOC_846/B OR2X1_LOC

XOR2X1_LOC_285 OR2X1_LOC_285/a_8_216# OR2X1_LOC_285/a_36_216# OR2X1_LOC_285/Y VSS VDD OR2X1_LOC_285/A OR2X1_LOC_285/B OR2X1_LOC

XOR2X1_LOC_254 OR2X1_LOC_254/a_8_216# OR2X1_LOC_254/a_36_216# OR2X1_LOC_456/A VSS VDD OR2X1_LOC_254/A OR2X1_LOC_254/B OR2X1_LOC

XAND2X1_LOC_99 AND2X1_LOC_99/a_36_24# AND2X1_LOC_99/Y AND2X1_LOC_99/a_8_24# VSS VDD AND2X1_LOC_99/A AND2X1_LOC_98/Y AND2X1_LOC

XOR2X1_LOC_116 OR2X1_LOC_116/a_8_216# OR2X1_LOC_116/a_36_216# OR2X1_LOC_216/A VSS VDD OR2X1_LOC_116/A OR2X1_LOC_114/Y OR2X1_LOC

XOR2X1_LOC_267 OR2X1_LOC_267/a_8_216# OR2X1_LOC_267/a_36_216# OR2X1_LOC_267/Y VSS VDD OR2X1_LOC_267/A OR2X1_LOC_641/A OR2X1_LOC

XOR2X1_LOC_802 OR2X1_LOC_802/a_8_216# OR2X1_LOC_802/a_36_216# OR2X1_LOC_802/Y VSS VDD OR2X1_LOC_802/A OR2X1_LOC_798/Y OR2X1_LOC

XAND2X1_LOC_162 AND2X1_LOC_162/a_36_24# OR2X1_LOC_163/A AND2X1_LOC_162/a_8_24# VSS VDD AND2X1_LOC_160/Y AND2X1_LOC_161/Y AND2X1_LOC

XOR2X1_LOC_162 OR2X1_LOC_162/a_8_216# OR2X1_LOC_162/a_36_216# OR2X1_LOC_162/Y VSS VDD OR2X1_LOC_162/A OR2X1_LOC_160/Y OR2X1_LOC

XOR2X1_LOC_331 OR2X1_LOC_331/a_8_216# OR2X1_LOC_331/a_36_216# OR2X1_LOC_331/Y VSS VDD OR2X1_LOC_331/A OR2X1_LOC_680/A OR2X1_LOC

XAND2X1_LOC_621 AND2X1_LOC_621/a_36_24# AND2X1_LOC_621/Y AND2X1_LOC_621/a_8_24# VSS VDD OR2X1_LOC_616/Y OR2X1_LOC_617/Y AND2X1_LOC

XOR2X1_LOC_629 OR2X1_LOC_629/a_8_216# OR2X1_LOC_629/a_36_216# OR2X1_LOC_629/Y VSS VDD OR2X1_LOC_629/A OR2X1_LOC_629/B OR2X1_LOC

XOR2X1_LOC_837 OR2X1_LOC_837/a_8_216# OR2X1_LOC_837/a_36_216# OR2X1_LOC_837/Y VSS VDD OR2X1_LOC_837/A OR2X1_LOC_837/B OR2X1_LOC

XAND2X1_LOC_846 AND2X1_LOC_846/a_36_24# AND2X1_LOC_848/A AND2X1_LOC_846/a_8_24# VSS VDD OR2X1_LOC_815/Y OR2X1_LOC_816/Y AND2X1_LOC

XAND2X1_LOC_285 AND2X1_LOC_285/a_36_24# AND2X1_LOC_285/Y AND2X1_LOC_285/a_8_24# VSS VDD OR2X1_LOC_281/Y OR2X1_LOC_282/Y AND2X1_LOC

XOR2X1_LOC_483 OR2X1_LOC_483/a_8_216# OR2X1_LOC_483/a_36_216# OR2X1_LOC_631/B VSS VDD OR2X1_LOC_833/B OR2X1_LOC_254/B OR2X1_LOC

XOR2X1_LOC_284 OR2X1_LOC_284/a_8_216# OR2X1_LOC_284/a_36_216# OR2X1_LOC_287/A VSS VDD OR2X1_LOC_542/B OR2X1_LOC_284/B OR2X1_LOC

XAND2X1_LOC_457 AND2X1_LOC_457/a_36_24# AND2X1_LOC_464/A AND2X1_LOC_457/a_8_24# VSS VDD OR2X1_LOC_368/Y AND2X1_LOC_787/A AND2X1_LOC

XOR2X1_LOC_99 OR2X1_LOC_99/a_8_216# OR2X1_LOC_99/a_36_216# OR2X1_LOC_99/Y VSS VDD OR2X1_LOC_99/A OR2X1_LOC_99/B OR2X1_LOC

XAND2X1_LOC_267 AND2X1_LOC_267/a_36_24# AND2X1_LOC_361/A AND2X1_LOC_267/a_8_24# VSS VDD OR2X1_LOC_265/Y AND2X1_LOC_266/Y AND2X1_LOC

XAND2X1_LOC_116 AND2X1_LOC_116/a_36_24# AND2X1_LOC_116/Y AND2X1_LOC_116/a_8_24# VSS VDD AND2X1_LOC_114/Y AND2X1_LOC_116/B AND2X1_LOC

XAND2X1_LOC_802 AND2X1_LOC_802/a_36_24# AND2X1_LOC_802/Y AND2X1_LOC_802/a_8_24# VSS VDD AND2X1_LOC_798/Y AND2X1_LOC_802/B AND2X1_LOC

XAND2X1_LOC_97 AND2X1_LOC_97/a_36_24# AND2X1_LOC_99/A AND2X1_LOC_97/a_8_24# VSS VDD OR2X1_LOC_89/Y OR2X1_LOC_91/Y AND2X1_LOC

XOR2X1_LOC_115 OR2X1_LOC_115/a_8_216# OR2X1_LOC_115/a_36_216# OR2X1_LOC_116/A VSS VDD OR2X1_LOC_715/B OR2X1_LOC_115/B OR2X1_LOC

XOR2X1_LOC_114 OR2X1_LOC_114/a_8_216# OR2X1_LOC_114/a_36_216# OR2X1_LOC_114/Y VSS VDD OR2X1_LOC_113/Y OR2X1_LOC_114/B OR2X1_LOC

XOR2X1_LOC_799 OR2X1_LOC_799/a_8_216# OR2X1_LOC_799/a_36_216# OR2X1_LOC_802/A VSS VDD OR2X1_LOC_799/A OR2X1_LOC_539/Y OR2X1_LOC

XOR2X1_LOC_798 OR2X1_LOC_798/a_8_216# OR2X1_LOC_798/a_36_216# OR2X1_LOC_798/Y VSS VDD OR2X1_LOC_436/Y OR2X1_LOC_319/Y OR2X1_LOC

XOR2X1_LOC_97 OR2X1_LOC_97/a_8_216# OR2X1_LOC_97/a_36_216# OR2X1_LOC_99/B VSS VDD OR2X1_LOC_97/A OR2X1_LOC_97/B OR2X1_LOC

XAND2X1_LOC_114 AND2X1_LOC_114/a_36_24# AND2X1_LOC_114/Y AND2X1_LOC_114/a_8_24# VSS VDD OR2X1_LOC_108/Y AND2X1_LOC_113/Y AND2X1_LOC

XAND2X1_LOC_115 AND2X1_LOC_115/a_36_24# AND2X1_LOC_116/B AND2X1_LOC_115/a_8_24# VSS VDD OR2X1_LOC_106/Y AND2X1_LOC_715/A AND2X1_LOC

XAND2X1_LOC_798 AND2X1_LOC_798/a_36_24# AND2X1_LOC_798/Y AND2X1_LOC_798/a_8_24# VSS VDD AND2X1_LOC_798/A AND2X1_LOC_436/Y AND2X1_LOC

XAND2X1_LOC_799 AND2X1_LOC_799/a_36_24# AND2X1_LOC_802/B AND2X1_LOC_799/a_8_24# VSS VDD AND2X1_LOC_539/Y AND2X1_LOC_593/Y AND2X1_LOC

XOR2X1_LOC_113 OR2X1_LOC_113/a_8_216# OR2X1_LOC_113/a_36_216# OR2X1_LOC_113/Y VSS VDD OR2X1_LOC_113/A OR2X1_LOC_113/B OR2X1_LOC

XOR2X1_LOC_593 OR2X1_LOC_593/a_8_216# OR2X1_LOC_593/a_36_216# OR2X1_LOC_799/A VSS VDD OR2X1_LOC_593/A OR2X1_LOC_593/B OR2X1_LOC

XOR2X1_LOC_539 OR2X1_LOC_539/a_8_216# OR2X1_LOC_539/a_36_216# OR2X1_LOC_539/Y VSS VDD OR2X1_LOC_539/A OR2X1_LOC_539/B OR2X1_LOC

XOR2X1_LOC_436 OR2X1_LOC_436/a_8_216# OR2X1_LOC_436/a_36_216# OR2X1_LOC_436/Y VSS VDD OR2X1_LOC_435/Y OR2X1_LOC_436/B OR2X1_LOC

XOR2X1_LOC_319 OR2X1_LOC_319/a_8_216# OR2X1_LOC_319/a_36_216# OR2X1_LOC_319/Y VSS VDD OR2X1_LOC_318/Y OR2X1_LOC_319/B OR2X1_LOC

XAND2X1_LOC_113 AND2X1_LOC_113/a_36_24# AND2X1_LOC_113/Y AND2X1_LOC_113/a_8_24# VSS VDD OR2X1_LOC_103/Y OR2X1_LOC_107/Y AND2X1_LOC

XAND2X1_LOC_319 AND2X1_LOC_319/a_36_24# AND2X1_LOC_798/A AND2X1_LOC_319/a_8_24# VSS VDD AND2X1_LOC_319/A AND2X1_LOC_318/Y AND2X1_LOC

XAND2X1_LOC_436 AND2X1_LOC_436/a_36_24# AND2X1_LOC_436/Y AND2X1_LOC_436/a_8_24# VSS VDD AND2X1_LOC_434/Y AND2X1_LOC_436/B AND2X1_LOC

XAND2X1_LOC_539 AND2X1_LOC_539/a_36_24# AND2X1_LOC_539/Y AND2X1_LOC_539/a_8_24# VSS VDD AND2X1_LOC_537/Y AND2X1_LOC_538/Y AND2X1_LOC

XAND2X1_LOC_593 AND2X1_LOC_593/a_36_24# AND2X1_LOC_593/Y AND2X1_LOC_593/a_8_24# VSS VDD OR2X1_LOC_591/Y AND2X1_LOC_592/Y AND2X1_LOC

XOR2X1_LOC_592 OR2X1_LOC_592/a_8_216# OR2X1_LOC_592/a_36_216# OR2X1_LOC_593/A VSS VDD OR2X1_LOC_592/A OR2X1_LOC_449/B OR2X1_LOC

XOR2X1_LOC_538 OR2X1_LOC_538/a_8_216# OR2X1_LOC_538/a_36_216# OR2X1_LOC_539/A VSS VDD OR2X1_LOC_538/A OR2X1_LOC_193/A OR2X1_LOC

XOR2X1_LOC_537 OR2X1_LOC_537/a_8_216# OR2X1_LOC_537/a_36_216# OR2X1_LOC_539/B VSS VDD OR2X1_LOC_537/A OR2X1_LOC_389/B OR2X1_LOC

XOR2X1_LOC_434 OR2X1_LOC_434/a_8_216# OR2X1_LOC_434/a_36_216# OR2X1_LOC_436/B VSS VDD OR2X1_LOC_434/A OR2X1_LOC_174/A OR2X1_LOC

XOR2X1_LOC_318 OR2X1_LOC_318/a_8_216# OR2X1_LOC_318/a_36_216# OR2X1_LOC_318/Y VSS VDD OR2X1_LOC_318/A OR2X1_LOC_318/B OR2X1_LOC

XOR2X1_LOC_317 OR2X1_LOC_317/a_8_216# OR2X1_LOC_317/a_36_216# OR2X1_LOC_319/B VSS VDD OR2X1_LOC_317/A OR2X1_LOC_317/B OR2X1_LOC

XAND2X1_LOC_317 AND2X1_LOC_317/a_36_24# AND2X1_LOC_319/A AND2X1_LOC_317/a_8_24# VSS VDD OR2X1_LOC_313/Y OR2X1_LOC_314/Y AND2X1_LOC

XAND2X1_LOC_318 AND2X1_LOC_318/a_36_24# AND2X1_LOC_318/Y AND2X1_LOC_318/a_8_24# VSS VDD OR2X1_LOC_315/Y OR2X1_LOC_316/Y AND2X1_LOC

XAND2X1_LOC_434 AND2X1_LOC_434/a_36_24# AND2X1_LOC_434/Y AND2X1_LOC_434/a_8_24# VSS VDD OR2X1_LOC_172/Y OR2X1_LOC_431/Y AND2X1_LOC

XAND2X1_LOC_537 AND2X1_LOC_537/a_36_24# AND2X1_LOC_537/Y AND2X1_LOC_537/a_8_24# VSS VDD OR2X1_LOC_385/Y OR2X1_LOC_536/Y AND2X1_LOC

XAND2X1_LOC_538 AND2X1_LOC_538/a_36_24# AND2X1_LOC_538/Y AND2X1_LOC_538/a_8_24# VSS VDD OR2X1_LOC_13/Y OR2X1_LOC_311/Y AND2X1_LOC

XAND2X1_LOC_592 AND2X1_LOC_592/a_36_24# AND2X1_LOC_592/Y AND2X1_LOC_592/a_8_24# VSS VDD OR2X1_LOC_423/Y OR2X1_LOC_589/Y AND2X1_LOC

C20418 VDD OR2X1_LOC_451/A -0.00fF
C30118 OR2X1_LOC_451/a_8_216# OR2X1_LOC_451/A 0.47fF
C40025 OR2X1_LOC_451/A OR2X1_LOC_451/B 0.05fF
C56903 OR2X1_LOC_451/A VSS 0.15fF
C6044 OR2X1_LOC_582/Y AND2X1_LOC_639/A 0.87fF
C20848 VDD OR2X1_LOC_582/Y 0.04fF
C22216 OR2X1_LOC_427/A OR2X1_LOC_582/Y 0.01fF
C39574 OR2X1_LOC_70/Y OR2X1_LOC_582/Y 0.01fF
C51231 OR2X1_LOC_582/Y AND2X1_LOC_635/a_8_24# 0.01fF
C56805 OR2X1_LOC_582/Y VSS 0.08fF
C7394 OR2X1_LOC_459/B OR2X1_LOC_460/A 0.88fF
C43050 OR2X1_LOC_460/B OR2X1_LOC_460/A 0.28fF
C56283 OR2X1_LOC_460/A VSS 0.15fF
C9632 OR2X1_LOC_197/A OR2X1_LOC_197/a_8_216# 0.47fF
C24775 OR2X1_LOC_197/A OR2X1_LOC_375/A 0.04fF
C57339 OR2X1_LOC_197/A VSS 0.05fF
C4203 OR2X1_LOC_307/a_8_216# OR2X1_LOC_307/B 0.06fF
C6185 OR2X1_LOC_307/B OR2X1_LOC_78/A 0.01fF
C24501 VDD OR2X1_LOC_307/B -0.00fF
C33148 OR2X1_LOC_307/B AND2X1_LOC_47/Y 0.01fF
C34144 AND2X1_LOC_22/Y OR2X1_LOC_307/B 0.04fF
C41056 OR2X1_LOC_307/B OR2X1_LOC_161/A 0.03fF
C43426 OR2X1_LOC_307/B AND2X1_LOC_31/Y 0.05fF
C45684 OR2X1_LOC_308/A OR2X1_LOC_307/B 0.88fF
C48391 OR2X1_LOC_307/B OR2X1_LOC_161/B 0.03fF
C57409 OR2X1_LOC_307/B VSS 0.12fF
C839 AND2X1_LOC_165/a_8_24# OR2X1_LOC_66/A 0.01fF
C1235 OR2X1_LOC_287/B OR2X1_LOC_66/A 0.03fF
C1271 OR2X1_LOC_76/A OR2X1_LOC_66/A 0.14fF
C1328 OR2X1_LOC_436/Y OR2X1_LOC_66/A 0.03fF
C1517 OR2X1_LOC_160/B OR2X1_LOC_66/A 0.42fF
C1612 OR2X1_LOC_553/A OR2X1_LOC_66/A 0.25fF
C2367 OR2X1_LOC_151/A OR2X1_LOC_66/A 0.19fF
C3330 OR2X1_LOC_137/B OR2X1_LOC_66/A 0.03fF
C3610 OR2X1_LOC_66/A OR2X1_LOC_415/Y 0.05fF
C4009 OR2X1_LOC_66/A OR2X1_LOC_168/Y 1.10fF
C4215 OR2X1_LOC_520/B OR2X1_LOC_66/A 0.17fF
C4803 OR2X1_LOC_66/A OR2X1_LOC_308/Y 0.07fF
C4907 AND2X1_LOC_125/a_8_24# OR2X1_LOC_66/A 0.02fF
C4979 OR2X1_LOC_593/A OR2X1_LOC_66/A 0.01fF
C5359 OR2X1_LOC_664/Y OR2X1_LOC_66/A 0.05fF
C5606 OR2X1_LOC_66/A OR2X1_LOC_342/a_8_216# 0.02fF
C5745 OR2X1_LOC_448/A OR2X1_LOC_66/A 0.03fF
C6113 OR2X1_LOC_66/A OR2X1_LOC_390/A 0.09fF
C6315 OR2X1_LOC_168/A OR2X1_LOC_66/A 0.01fF
C6621 AND2X1_LOC_314/a_8_24# OR2X1_LOC_66/A 0.03fF
C6655 OR2X1_LOC_668/Y OR2X1_LOC_66/A 0.01fF
C7026 AND2X1_LOC_311/a_8_24# OR2X1_LOC_66/A 0.09fF
C7256 OR2X1_LOC_84/A OR2X1_LOC_66/A 0.02fF
C7289 OR2X1_LOC_98/B OR2X1_LOC_66/A 0.23fF
C7482 AND2X1_LOC_94/Y OR2X1_LOC_66/A 0.03fF
C7718 OR2X1_LOC_66/A OR2X1_LOC_241/B 0.54fF
C8259 OR2X1_LOC_66/A OR2X1_LOC_339/A 0.01fF
C8297 OR2X1_LOC_208/A OR2X1_LOC_66/A 0.04fF
C8346 OR2X1_LOC_598/Y OR2X1_LOC_66/A 0.23fF
C8413 AND2X1_LOC_40/Y OR2X1_LOC_66/A 1.06fF
C8449 OR2X1_LOC_537/A OR2X1_LOC_66/A 0.03fF
C8753 OR2X1_LOC_66/A OR2X1_LOC_356/A 0.06fF
C9337 OR2X1_LOC_810/A OR2X1_LOC_66/A 0.18fF
C9355 AND2X1_LOC_589/a_8_24# OR2X1_LOC_66/A 0.01fF
C9607 OR2X1_LOC_715/B OR2X1_LOC_66/A 0.08fF
C9616 OR2X1_LOC_784/B OR2X1_LOC_66/A 0.01fF
C10569 AND2X1_LOC_399/a_8_24# OR2X1_LOC_66/A 0.01fF
C10652 OR2X1_LOC_606/Y OR2X1_LOC_66/A 0.07fF
C10942 OR2X1_LOC_828/B OR2X1_LOC_66/A 0.14fF
C11298 OR2X1_LOC_78/A OR2X1_LOC_66/A 0.55fF
C11331 OR2X1_LOC_448/B OR2X1_LOC_66/A 0.02fF
C12240 AND2X1_LOC_669/a_8_24# OR2X1_LOC_66/A 0.01fF
C12541 OR2X1_LOC_121/Y OR2X1_LOC_66/A 0.01fF
C12559 OR2X1_LOC_114/B OR2X1_LOC_66/A 0.03fF
C12586 OR2X1_LOC_538/A OR2X1_LOC_66/A 0.05fF
C12659 AND2X1_LOC_12/Y OR2X1_LOC_66/A 0.27fF
C12720 AND2X1_LOC_79/Y OR2X1_LOC_66/A 0.03fF
C12841 OR2X1_LOC_98/a_8_216# OR2X1_LOC_66/A -0.00fF
C13046 OR2X1_LOC_168/B OR2X1_LOC_66/A 0.03fF
C13121 AND2X1_LOC_59/Y OR2X1_LOC_66/A 1.00fF
C13369 OR2X1_LOC_66/A OR2X1_LOC_342/B 0.01fF
C13944 OR2X1_LOC_833/B OR2X1_LOC_66/A 0.03fF
C14779 OR2X1_LOC_448/Y OR2X1_LOC_66/A 0.01fF
C14841 OR2X1_LOC_592/A OR2X1_LOC_66/A 0.01fF
C15457 OR2X1_LOC_66/A OR2X1_LOC_338/A 0.01fF
C15476 OR2X1_LOC_186/Y OR2X1_LOC_66/A 0.44fF
C15738 OR2X1_LOC_112/B OR2X1_LOC_66/A 0.20fF
C16082 OR2X1_LOC_574/A OR2X1_LOC_66/A 0.03fF
C16705 OR2X1_LOC_66/A OR2X1_LOC_539/B 0.01fF
C16819 OR2X1_LOC_78/B OR2X1_LOC_66/A 10.24fF
C16861 OR2X1_LOC_448/a_8_216# OR2X1_LOC_66/A 0.01fF
C16904 OR2X1_LOC_375/A OR2X1_LOC_66/A 0.36fF
C17212 OR2X1_LOC_66/A OR2X1_LOC_549/A 0.12fF
C17261 OR2X1_LOC_113/Y OR2X1_LOC_66/A 0.01fF
C18796 OR2X1_LOC_779/Y OR2X1_LOC_66/A 0.01fF
C19055 OR2X1_LOC_673/Y OR2X1_LOC_66/A 1.16fF
C19561 AND2X1_LOC_27/a_8_24# OR2X1_LOC_66/A 0.11fF
C19762 OR2X1_LOC_139/A OR2X1_LOC_66/A 0.05fF
C20659 AND2X1_LOC_595/a_8_24# OR2X1_LOC_66/A 0.05fF
C21014 OR2X1_LOC_66/A AND2X1_LOC_235/a_8_24# 0.01fF
C21160 OR2X1_LOC_668/a_8_216# OR2X1_LOC_66/A 0.10fF
C21196 OR2X1_LOC_703/B OR2X1_LOC_66/A 0.29fF
C21209 OR2X1_LOC_87/A OR2X1_LOC_66/A 0.11fF
C21459 OR2X1_LOC_66/A OR2X1_LOC_844/B 0.02fF
C21537 OR2X1_LOC_389/A OR2X1_LOC_66/A 0.03fF
C21569 AND2X1_LOC_177/a_8_24# OR2X1_LOC_66/A 0.01fF
C21656 OR2X1_LOC_403/B OR2X1_LOC_66/A 0.01fF
C22293 OR2X1_LOC_66/A OR2X1_LOC_349/B 0.01fF
C22351 OR2X1_LOC_97/A OR2X1_LOC_66/A 0.02fF
C22463 AND2X1_LOC_290/a_8_24# OR2X1_LOC_66/A 0.14fF
C22815 OR2X1_LOC_691/Y OR2X1_LOC_66/A 0.03fF
C22824 OR2X1_LOC_66/A OR2X1_LOC_713/A 0.07fF
C22917 OR2X1_LOC_249/a_8_216# OR2X1_LOC_66/A 0.02fF
C23339 OR2X1_LOC_720/A OR2X1_LOC_66/A 0.01fF
C23412 OR2X1_LOC_99/B OR2X1_LOC_66/A 0.14fF
C23754 OR2X1_LOC_154/A OR2X1_LOC_66/A 1.06fF
C23922 OR2X1_LOC_99/A OR2X1_LOC_66/A 0.03fF
C23947 OR2X1_LOC_66/A OR2X1_LOC_198/A 0.08fF
C24109 AND2X1_LOC_96/a_8_24# OR2X1_LOC_66/A 0.01fF
C24306 AND2X1_LOC_813/a_8_24# OR2X1_LOC_66/A 0.01fF
C24493 OR2X1_LOC_634/A OR2X1_LOC_66/A 0.90fF
C24846 OR2X1_LOC_267/Y OR2X1_LOC_66/A 0.02fF
C24864 OR2X1_LOC_633/A OR2X1_LOC_66/A 0.03fF
C24984 OR2X1_LOC_520/Y OR2X1_LOC_66/A 0.14fF
C25254 AND2X1_LOC_64/Y OR2X1_LOC_66/A 0.22fF
C25691 OR2X1_LOC_66/A OR2X1_LOC_342/A 0.03fF
C25751 OR2X1_LOC_756/B OR2X1_LOC_66/A 0.75fF
C25898 AND2X1_LOC_677/a_8_24# OR2X1_LOC_66/A 0.07fF
C26225 OR2X1_LOC_379/a_8_216# OR2X1_LOC_66/A 0.01fF
C26296 OR2X1_LOC_719/A OR2X1_LOC_66/A 0.09fF
C26521 OR2X1_LOC_66/A OR2X1_LOC_779/A 0.74fF
C26626 OR2X1_LOC_668/a_36_216# OR2X1_LOC_66/A 0.03fF
C26688 OR2X1_LOC_708/B OR2X1_LOC_66/A 0.01fF
C27120 OR2X1_LOC_87/B OR2X1_LOC_66/A 0.02fF
C27617 OR2X1_LOC_532/B OR2X1_LOC_66/A 0.20fF
C27627 AND2X1_LOC_665/a_8_24# OR2X1_LOC_66/A 0.02fF
C27829 OR2X1_LOC_440/B OR2X1_LOC_66/A 0.03fF
C27945 OR2X1_LOC_99/a_8_216# OR2X1_LOC_66/A 0.01fF
C29145 AND2X1_LOC_52/a_8_24# OR2X1_LOC_66/A 0.02fF
C29529 VDD OR2X1_LOC_66/A 1.81fF
C29553 OR2X1_LOC_98/A OR2X1_LOC_66/A 0.01fF
C29768 OR2X1_LOC_845/A OR2X1_LOC_66/A 0.03fF
C30462 OR2X1_LOC_462/B OR2X1_LOC_66/A 0.02fF
C30754 AND2X1_LOC_83/a_8_24# OR2X1_LOC_66/A 0.08fF
C31583 OR2X1_LOC_66/A OR2X1_LOC_115/B 0.01fF
C31673 OR2X1_LOC_840/A OR2X1_LOC_66/A 0.03fF
C32125 OR2X1_LOC_802/Y OR2X1_LOC_66/A 0.14fF
C32147 AND2X1_LOC_385/a_8_24# OR2X1_LOC_66/A 0.05fF
C32195 AND2X1_LOC_134/a_8_24# OR2X1_LOC_66/A 0.01fF
C32451 OR2X1_LOC_809/B OR2X1_LOC_66/A 0.59fF
C32546 OR2X1_LOC_160/A OR2X1_LOC_66/A 0.19fF
C32610 AND2X1_LOC_86/B OR2X1_LOC_66/A 0.06fF
C32621 OR2X1_LOC_624/B OR2X1_LOC_66/A 0.03fF
C32846 OR2X1_LOC_266/A OR2X1_LOC_66/A 0.01fF
C32868 AND2X1_LOC_607/a_8_24# OR2X1_LOC_66/A 0.14fF
C32965 OR2X1_LOC_447/A OR2X1_LOC_66/A 0.02fF
C33270 OR2X1_LOC_113/a_8_216# OR2X1_LOC_66/A 0.02fF
C33396 AND2X1_LOC_290/a_36_24# OR2X1_LOC_66/A 0.01fF
C33794 OR2X1_LOC_708/Y OR2X1_LOC_66/A 0.01fF
C33829 OR2X1_LOC_185/A OR2X1_LOC_66/A 0.64fF
C33840 OR2X1_LOC_249/Y OR2X1_LOC_66/A 0.11fF
C34285 OR2X1_LOC_702/A OR2X1_LOC_66/A 0.04fF
C34575 AND2X1_LOC_437/a_8_24# OR2X1_LOC_66/A 0.01fF
C34998 OR2X1_LOC_294/Y OR2X1_LOC_66/A 0.03fF
C35071 OR2X1_LOC_379/Y OR2X1_LOC_66/A 0.14fF
C35485 OR2X1_LOC_168/a_8_216# OR2X1_LOC_66/A 0.01fF
C35958 OR2X1_LOC_643/A OR2X1_LOC_66/A 0.04fF
C35960 OR2X1_LOC_778/Y OR2X1_LOC_66/A 0.14fF
C36042 OR2X1_LOC_113/A OR2X1_LOC_66/A 0.03fF
C36206 AND2X1_LOC_91/B OR2X1_LOC_66/A 13.85fF
C36342 OR2X1_LOC_799/A OR2X1_LOC_66/A 0.12fF
C36561 OR2X1_LOC_66/A OR2X1_LOC_446/B 0.03fF
C36567 OR2X1_LOC_66/A OR2X1_LOC_303/B 0.03fF
C36644 OR2X1_LOC_66/A OR2X1_LOC_719/B 0.03fF
C36757 AND2X1_LOC_56/B OR2X1_LOC_66/A 0.19fF
C37173 AND2X1_LOC_166/a_8_24# OR2X1_LOC_66/A 0.03fF
C37634 OR2X1_LOC_83/A OR2X1_LOC_66/A 0.03fF
C37636 OR2X1_LOC_389/B OR2X1_LOC_66/A 0.41fF
C38153 AND2X1_LOC_47/Y OR2X1_LOC_66/A 6.92fF
C38341 OR2X1_LOC_646/B OR2X1_LOC_66/A 0.01fF
C38447 OR2X1_LOC_506/A OR2X1_LOC_66/A 0.09fF
C38735 OR2X1_LOC_66/A OR2X1_LOC_180/B 0.01fF
C38896 AND2X1_LOC_95/Y OR2X1_LOC_66/A 13.47fF
C38901 OR2X1_LOC_633/Y OR2X1_LOC_66/A 0.03fF
C38942 OR2X1_LOC_99/Y OR2X1_LOC_66/A 0.39fF
C39155 OR2X1_LOC_66/A OR2X1_LOC_788/B 0.06fF
C39203 AND2X1_LOC_22/Y OR2X1_LOC_66/A 0.70fF
C40079 OR2X1_LOC_235/B OR2X1_LOC_66/A 0.09fF
C40357 OR2X1_LOC_66/A OR2X1_LOC_779/B 0.14fF
C40477 OR2X1_LOC_709/A OR2X1_LOC_66/A 0.07fF
C40517 AND2X1_LOC_70/Y OR2X1_LOC_66/A 6.41fF
C40895 OR2X1_LOC_362/A OR2X1_LOC_66/A 0.03fF
C40962 OR2X1_LOC_539/A OR2X1_LOC_66/A 0.03fF
C41138 OR2X1_LOC_243/B OR2X1_LOC_66/A 0.05fF
C41270 OR2X1_LOC_66/A OR2X1_LOC_771/B 0.06fF
C41732 OR2X1_LOC_66/A OR2X1_LOC_593/B 0.04fF
C42193 OR2X1_LOC_66/A AND2X1_LOC_44/Y 0.60fF
C42475 OR2X1_LOC_720/B OR2X1_LOC_66/A 0.03fF
C43086 OR2X1_LOC_66/A OR2X1_LOC_708/a_8_216# 0.02fF
C43124 AND2X1_LOC_18/Y OR2X1_LOC_66/A 1.37fF
C43526 OR2X1_LOC_112/a_8_216# OR2X1_LOC_66/A 0.01fF
C43535 OR2X1_LOC_307/A OR2X1_LOC_66/A 0.22fF
C43659 AND2X1_LOC_394/a_8_24# OR2X1_LOC_66/A 0.01fF
C44069 OR2X1_LOC_447/a_8_216# OR2X1_LOC_66/A 0.05fF
C44083 OR2X1_LOC_130/A OR2X1_LOC_66/A 0.04fF
C44537 OR2X1_LOC_449/B OR2X1_LOC_66/A 0.87fF
C45341 OR2X1_LOC_175/B OR2X1_LOC_66/A 0.02fF
C45678 OR2X1_LOC_66/A OR2X1_LOC_389/a_8_216# 0.01fF
C45934 OR2X1_LOC_447/Y OR2X1_LOC_66/A 0.03fF
C46245 OR2X1_LOC_161/A OR2X1_LOC_66/A 1.21fF
C46347 AND2X1_LOC_51/Y OR2X1_LOC_66/A 0.23fF
C46916 OR2X1_LOC_66/A AND2X1_LOC_52/Y 0.03fF
C47060 OR2X1_LOC_439/B OR2X1_LOC_66/A 0.09fF
C47116 AND2X1_LOC_41/A OR2X1_LOC_66/A 0.17fF
C47210 OR2X1_LOC_631/B OR2X1_LOC_66/A 0.07fF
C47859 OR2X1_LOC_66/A OR2X1_LOC_112/A 0.39fF
C47885 AND2X1_LOC_57/Y OR2X1_LOC_66/A 0.05fF
C48301 OR2X1_LOC_66/A OR2X1_LOC_71/A 0.08fF
C48514 OR2X1_LOC_593/a_8_216# OR2X1_LOC_66/A 0.01fF
C48673 AND2X1_LOC_31/Y OR2X1_LOC_66/A 1.84fF
C48913 OR2X1_LOC_809/a_8_216# OR2X1_LOC_66/A 0.01fF
C48927 OR2X1_LOC_66/A OR2X1_LOC_240/A 2.75fF
C49149 OR2X1_LOC_66/A OR2X1_LOC_397/a_8_216# 0.03fF
C49502 AND2X1_LOC_72/B OR2X1_LOC_66/A 0.03fF
C49584 OR2X1_LOC_66/A AND2X1_LOC_36/Y 0.47fF
C50155 OR2X1_LOC_128/B OR2X1_LOC_66/A 0.01fF
C50194 OR2X1_LOC_592/a_8_216# OR2X1_LOC_66/A 0.01fF
C50835 OR2X1_LOC_66/A OR2X1_LOC_537/a_8_216# 0.02fF
C51348 OR2X1_LOC_768/A OR2X1_LOC_66/A 0.01fF
C51871 OR2X1_LOC_269/B OR2X1_LOC_66/A 0.24fF
C52236 OR2X1_LOC_347/B OR2X1_LOC_66/A 0.03fF
C52246 OR2X1_LOC_539/Y OR2X1_LOC_66/A 0.08fF
C52266 OR2X1_LOC_779/a_8_216# OR2X1_LOC_66/A 0.01fF
C52324 AND2X1_LOC_176/a_8_24# OR2X1_LOC_66/A 0.01fF
C52860 OR2X1_LOC_66/A AND2X1_LOC_237/a_8_24# 0.01fF
C52935 OR2X1_LOC_66/A OR2X1_LOC_777/B 0.06fF
C52990 OR2X1_LOC_344/A OR2X1_LOC_66/A 0.03fF
C53332 OR2X1_LOC_66/A OR2X1_LOC_332/a_8_216# 0.01fF
C53371 OR2X1_LOC_198/a_8_216# OR2X1_LOC_66/A 0.04fF
C53405 OR2X1_LOC_66/A OR2X1_LOC_161/B 0.32fF
C53486 OR2X1_LOC_435/B OR2X1_LOC_66/A 0.34fF
C53933 AND2X1_LOC_132/a_8_24# OR2X1_LOC_66/A 0.01fF
C54268 OR2X1_LOC_520/a_8_216# OR2X1_LOC_66/A 0.14fF
C54349 OR2X1_LOC_539/a_8_216# OR2X1_LOC_66/A 0.02fF
C54419 OR2X1_LOC_3/Y OR2X1_LOC_66/A 0.03fF
C54676 OR2X1_LOC_777/a_8_216# OR2X1_LOC_66/A 0.01fF
C54778 OR2X1_LOC_400/A OR2X1_LOC_66/A 0.01fF
C54900 AND2X1_LOC_106/a_8_24# OR2X1_LOC_66/A 0.02fF
C55267 AND2X1_LOC_3/Y OR2X1_LOC_66/A 0.34fF
C55947 AND2X1_LOC_7/B OR2X1_LOC_66/A 0.15fF
C56027 OR2X1_LOC_319/B OR2X1_LOC_66/A 0.17fF
C56039 OR2X1_LOC_318/Y OR2X1_LOC_66/A 0.03fF
C56505 OR2X1_LOC_66/A VSS -4.58fF
C19 AND2X1_LOC_22/Y OR2X1_LOC_198/A 0.12fF
C126 AND2X1_LOC_22/Y OR2X1_LOC_435/A 0.08fF
C603 AND2X1_LOC_22/Y AND2X1_LOC_20/a_8_24# 0.03fF
C768 AND2X1_LOC_22/Y OR2X1_LOC_335/B 0.05fF
C1121 AND2X1_LOC_22/Y OR2X1_LOC_520/Y 0.07fF
C1226 AND2X1_LOC_22/Y AND2X1_LOC_107/a_8_24# 0.06fF
C1418 AND2X1_LOC_64/Y AND2X1_LOC_22/Y 0.43fF
C1512 OR2X1_LOC_512/A AND2X1_LOC_22/Y 0.01fF
C1885 AND2X1_LOC_22/Y OR2X1_LOC_776/Y 0.20fF
C1921 AND2X1_LOC_22/Y OR2X1_LOC_756/B 0.08fF
C2753 OR2X1_LOC_653/B AND2X1_LOC_22/Y 0.01fF
C2757 OR2X1_LOC_614/Y AND2X1_LOC_22/Y 0.27fF
C3324 AND2X1_LOC_22/Y OR2X1_LOC_33/B 0.09fF
C3549 AND2X1_LOC_22/Y OR2X1_LOC_333/A 0.20fF
C3650 OR2X1_LOC_100/Y AND2X1_LOC_22/Y 1.97fF
C3658 AND2X1_LOC_22/Y AND2X1_LOC_58/a_36_24# 0.01fF
C3803 AND2X1_LOC_22/Y OR2X1_LOC_532/B 0.11fF
C4374 AND2X1_LOC_22/Y OR2X1_LOC_855/a_8_216# 0.03fF
C4426 OR2X1_LOC_114/a_8_216# AND2X1_LOC_22/Y 0.07fF
C5659 AND2X1_LOC_22/Y VDD 0.73fF
C5912 AND2X1_LOC_22/Y OR2X1_LOC_845/A 0.05fF
C6426 AND2X1_LOC_22/Y OR2X1_LOC_523/A 0.33fF
C6453 OR2X1_LOC_335/a_8_216# AND2X1_LOC_22/Y 0.01fF
C6515 AND2X1_LOC_22/Y OR2X1_LOC_834/A 0.08fF
C7785 AND2X1_LOC_22/Y OR2X1_LOC_115/B 0.02fF
C7878 AND2X1_LOC_22/Y OR2X1_LOC_840/A 0.03fF
C8299 AND2X1_LOC_754/a_8_24# AND2X1_LOC_22/Y 0.17fF
C8488 AND2X1_LOC_22/Y AND2X1_LOC_134/a_8_24# 0.03fF
C8786 OR2X1_LOC_160/A AND2X1_LOC_22/Y 0.12fF
C9104 OR2X1_LOC_196/Y AND2X1_LOC_22/Y 0.35fF
C10024 AND2X1_LOC_22/Y OR2X1_LOC_608/a_8_216# 0.03fF
C10044 AND2X1_LOC_22/Y OR2X1_LOC_185/A 0.16fF
C10122 AND2X1_LOC_22/Y OR2X1_LOC_435/Y 0.34fF
C10186 AND2X1_LOC_22/Y AND2X1_LOC_431/a_8_24# -0.00fF
C10493 AND2X1_LOC_22/Y AND2X1_LOC_669/a_36_24# 0.01fF
C10814 AND2X1_LOC_22/Y AND2X1_LOC_262/a_8_24# 0.04fF
C11291 OR2X1_LOC_379/Y AND2X1_LOC_22/Y 0.03fF
C11324 AND2X1_LOC_22/Y OR2X1_LOC_114/Y 0.03fF
C11697 AND2X1_LOC_22/Y AND2X1_LOC_20/a_36_24# 0.01fF
C12123 AND2X1_LOC_22/Y OR2X1_LOC_637/A 0.01fF
C12126 AND2X1_LOC_22/Y OR2X1_LOC_436/B 0.01fF
C12186 AND2X1_LOC_22/Y OR2X1_LOC_643/A 0.07fF
C12193 AND2X1_LOC_22/Y OR2X1_LOC_778/Y 0.05fF
C12285 AND2X1_LOC_22/Y OR2X1_LOC_113/A 0.03fF
C12470 AND2X1_LOC_91/B AND2X1_LOC_22/Y 0.25fF
C12575 AND2X1_LOC_22/Y OR2X1_LOC_799/A 0.17fF
C12842 AND2X1_LOC_22/Y OR2X1_LOC_446/B 0.03fF
C12849 AND2X1_LOC_22/Y OR2X1_LOC_303/B 0.57fF
C13066 AND2X1_LOC_22/Y AND2X1_LOC_56/B 0.10fF
C13797 OR2X1_LOC_790/A AND2X1_LOC_22/Y 0.01fF
C14440 AND2X1_LOC_22/Y AND2X1_LOC_47/Y 0.45fF
C14644 AND2X1_LOC_521/a_8_24# AND2X1_LOC_22/Y 0.03fF
C14692 AND2X1_LOC_22/Y OR2X1_LOC_828/a_8_216# 0.03fF
C14715 AND2X1_LOC_22/Y OR2X1_LOC_506/A 0.02fF
C14908 AND2X1_LOC_22/Y AND2X1_LOC_48/Y 0.04fF
C15125 AND2X1_LOC_22/Y AND2X1_LOC_95/Y 0.26fF
C15156 AND2X1_LOC_22/Y OR2X1_LOC_99/Y 0.05fF
C15371 AND2X1_LOC_22/Y AND2X1_LOC_41/Y 0.02fF
C15507 AND2X1_LOC_22/Y OR2X1_LOC_608/a_36_216# 0.02fF
C15652 AND2X1_LOC_22/Y OR2X1_LOC_434/A 0.31fF
C16328 AND2X1_LOC_22/Y OR2X1_LOC_235/B 0.16fF
C16605 AND2X1_LOC_22/Y OR2X1_LOC_779/B 0.01fF
C16758 AND2X1_LOC_22/Y AND2X1_LOC_70/Y 8.99fF
C17170 AND2X1_LOC_22/Y OR2X1_LOC_362/A 0.07fF
C17510 AND2X1_LOC_22/Y OR2X1_LOC_771/B 0.01fF
C17944 AND2X1_LOC_22/Y OR2X1_LOC_593/B 0.03fF
C18440 AND2X1_LOC_22/Y AND2X1_LOC_44/Y 0.21fF
C18663 AND2X1_LOC_22/Y OR2X1_LOC_720/B 0.01fF
C19322 AND2X1_LOC_22/Y AND2X1_LOC_18/Y 13.06fF
C19750 AND2X1_LOC_22/Y OR2X1_LOC_307/A 0.28fF
C20174 OR2X1_LOC_523/B AND2X1_LOC_22/Y 0.01fF
C20242 OR2X1_LOC_101/a_8_216# AND2X1_LOC_22/Y 0.03fF
C20265 AND2X1_LOC_22/Y OR2X1_LOC_130/A 0.42fF
C20275 AND2X1_LOC_22/Y AND2X1_LOC_7/a_8_24# 0.02fF
C20716 AND2X1_LOC_22/Y OR2X1_LOC_449/B 0.03fF
C20973 AND2X1_LOC_22/Y OR2X1_LOC_195/a_8_216# 0.01fF
C22400 AND2X1_LOC_22/Y OR2X1_LOC_161/A 0.94fF
C22500 AND2X1_LOC_22/Y AND2X1_LOC_51/Y 0.81fF
C22880 AND2X1_LOC_22/Y OR2X1_LOC_831/a_8_216# 0.01fF
C23055 AND2X1_LOC_22/Y AND2X1_LOC_52/Y 0.03fF
C23222 AND2X1_LOC_22/Y AND2X1_LOC_41/A 0.10fF
C24728 AND2X1_LOC_22/Y AND2X1_LOC_31/Y 1.36fF
C24959 AND2X1_LOC_22/Y OR2X1_LOC_633/B 0.03fF
C25020 AND2X1_LOC_22/Y AND2X1_LOC_134/a_36_24# 0.01fF
C25510 AND2X1_LOC_22/Y AND2X1_LOC_72/B 0.02fF
C25608 AND2X1_LOC_22/Y AND2X1_LOC_36/Y 2.94fF
C25627 AND2X1_LOC_22/Y OR2X1_LOC_333/a_8_216# 0.02fF
C25717 OR2X1_LOC_635/A AND2X1_LOC_22/Y 0.01fF
C25736 AND2X1_LOC_586/a_8_24# AND2X1_LOC_22/Y 0.01fF
C25920 AND2X1_LOC_22/Y OR2X1_LOC_196/a_8_216# 0.01fF
C26480 AND2X1_LOC_22/Y AND2X1_LOC_522/a_8_24# 0.06fF
C27358 AND2X1_LOC_22/Y AND2X1_LOC_262/a_36_24# 0.01fF
C27378 OR2X1_LOC_768/A AND2X1_LOC_22/Y 0.02fF
C27881 AND2X1_LOC_22/Y OR2X1_LOC_269/B 0.18fF
C28960 AND2X1_LOC_22/Y OR2X1_LOC_777/B 0.03fF
C28996 AND2X1_LOC_22/Y OR2X1_LOC_831/B 0.03fF
C29438 AND2X1_LOC_22/Y OR2X1_LOC_161/B 0.05fF
C29508 AND2X1_LOC_22/Y OR2X1_LOC_435/B 0.21fF
C29962 AND2X1_LOC_22/Y AND2X1_LOC_132/a_8_24# 0.02fF
C31226 OR2X1_LOC_101/a_36_216# AND2X1_LOC_22/Y 0.02fF
C31286 AND2X1_LOC_22/Y AND2X1_LOC_3/Y 0.35fF
C31936 AND2X1_LOC_22/Y AND2X1_LOC_7/B 0.10fF
C32012 AND2X1_LOC_22/Y OR2X1_LOC_318/Y 0.01fF
C33426 AND2X1_LOC_22/Y OR2X1_LOC_76/A 0.50fF
C33495 AND2X1_LOC_22/Y OR2X1_LOC_436/Y 0.01fF
C33713 AND2X1_LOC_22/Y OR2X1_LOC_160/B 0.80fF
C33789 AND2X1_LOC_22/Y OR2X1_LOC_266/a_8_216# 0.03fF
C33979 AND2X1_LOC_22/Y OR2X1_LOC_197/a_8_216# 0.05fF
C34498 AND2X1_LOC_22/Y OR2X1_LOC_151/A 0.03fF
C34990 OR2X1_LOC_769/A AND2X1_LOC_22/Y 0.07fF
C35005 AND2X1_LOC_22/Y OR2X1_LOC_174/A 0.28fF
C35009 AND2X1_LOC_22/Y OR2X1_LOC_435/a_8_216# 0.01fF
C35425 AND2X1_LOC_22/Y OR2X1_LOC_137/B 0.02fF
C36470 AND2X1_LOC_22/Y AND2X1_LOC_497/a_8_24# 0.05fF
C37007 AND2X1_LOC_22/Y AND2X1_LOC_604/a_8_24# 0.01fF
C37414 AND2X1_LOC_22/Y OR2X1_LOC_301/a_8_216# 0.01fF
C37442 AND2X1_LOC_22/Y OR2X1_LOC_828/Y 0.03fF
C37457 AND2X1_LOC_22/Y AND2X1_LOC_522/a_36_24# 0.01fF
C37904 AND2X1_LOC_22/Y AND2X1_LOC_24/a_8_24# 0.03fF
C38070 AND2X1_LOC_22/Y AND2X1_LOC_7/Y 0.01fF
C38298 AND2X1_LOC_22/Y OR2X1_LOC_390/A 0.03fF
C38847 AND2X1_LOC_22/Y OR2X1_LOC_668/Y 0.05fF
C39207 AND2X1_LOC_22/Y OR2X1_LOC_841/A 0.03fF
C40045 AND2X1_LOC_22/Y AND2X1_LOC_615/a_8_24# 0.04fF
C40356 AND2X1_LOC_22/Y OR2X1_LOC_339/A 0.12fF
C40438 AND2X1_LOC_22/Y OR2X1_LOC_831/A 0.38fF
C40446 AND2X1_LOC_22/Y OR2X1_LOC_598/Y 0.06fF
C40483 OR2X1_LOC_335/Y AND2X1_LOC_22/Y 0.09fF
C40502 AND2X1_LOC_40/Y AND2X1_LOC_22/Y 0.15fF
C40939 AND2X1_LOC_22/Y AND2X1_LOC_132/a_36_24# 0.01fF
C41429 AND2X1_LOC_22/Y OR2X1_LOC_810/A 0.16fF
C41430 OR2X1_LOC_307/a_8_216# AND2X1_LOC_22/Y 0.01fF
C41455 AND2X1_LOC_22/Y AND2X1_LOC_589/a_8_24# 0.03fF
C41755 OR2X1_LOC_715/B AND2X1_LOC_22/Y 0.03fF
C42140 AND2X1_LOC_22/Y OR2X1_LOC_338/B 0.06fF
C42252 OR2X1_LOC_656/B AND2X1_LOC_22/Y 0.03fF
C42733 AND2X1_LOC_22/Y OR2X1_LOC_687/Y 0.03fF
C42993 AND2X1_LOC_22/Y OR2X1_LOC_199/B 0.01fF
C43152 AND2X1_LOC_22/Y OR2X1_LOC_828/B 0.03fF
C43519 AND2X1_LOC_22/Y OR2X1_LOC_78/A 0.14fF
C43646 AND2X1_LOC_22/Y OR2X1_LOC_605/A 0.04fF
C44436 AND2X1_LOC_22/Y AND2X1_LOC_669/a_8_24# 0.08fF
C44474 AND2X1_LOC_22/Y AND2X1_LOC_171/a_8_24# 0.02fF
C44642 AND2X1_LOC_22/Y OR2X1_LOC_318/B 0.05fF
C44788 OR2X1_LOC_114/B AND2X1_LOC_22/Y 0.05fF
C44860 AND2X1_LOC_12/Y AND2X1_LOC_22/Y 0.34fF
C44885 AND2X1_LOC_22/Y OR2X1_LOC_841/B 0.05fF
C45255 AND2X1_LOC_22/Y OR2X1_LOC_168/B 0.15fF
C45309 AND2X1_LOC_59/Y AND2X1_LOC_22/Y 1.70fF
C45647 OR2X1_LOC_318/a_8_216# AND2X1_LOC_22/Y 0.01fF
C45706 AND2X1_LOC_22/Y OR2X1_LOC_623/B 0.01fF
C46149 AND2X1_LOC_22/Y OR2X1_LOC_434/a_8_216# 0.02fF
C46151 AND2X1_LOC_22/Y OR2X1_LOC_776/a_8_216# 0.01fF
C47862 AND2X1_LOC_22/Y OR2X1_LOC_338/A 0.83fF
C47999 AND2X1_LOC_81/B AND2X1_LOC_22/Y 0.03fF
C48089 AND2X1_LOC_22/Y OR2X1_LOC_196/B 0.02fF
C48161 AND2X1_LOC_22/Y OR2X1_LOC_112/B 0.31fF
C48477 AND2X1_LOC_22/Y OR2X1_LOC_574/A 0.03fF
C48716 AND2X1_LOC_22/Y OR2X1_LOC_855/A 0.01fF
C48787 AND2X1_LOC_22/Y AND2X1_LOC_58/a_8_24# 0.03fF
C49079 AND2X1_LOC_22/Y OR2X1_LOC_539/B 0.02fF
C49181 AND2X1_LOC_22/Y OR2X1_LOC_78/B 0.34fF
C49231 AND2X1_LOC_22/Y OR2X1_LOC_375/A 0.32fF
C49309 AND2X1_LOC_22/Y OR2X1_LOC_605/B 0.03fF
C49601 AND2X1_LOC_22/Y OR2X1_LOC_549/A 0.07fF
C49640 OR2X1_LOC_113/Y AND2X1_LOC_22/Y 0.06fF
C50448 AND2X1_LOC_22/Y AND2X1_LOC_65/A 0.03fF
C51281 AND2X1_LOC_22/Y AND2X1_LOC_19/Y 2.57fF
C51375 AND2X1_LOC_22/Y OR2X1_LOC_673/Y 0.10fF
C51400 AND2X1_LOC_22/Y OR2X1_LOC_195/A 0.08fF
C51592 AND2X1_LOC_22/Y OR2X1_LOC_769/a_8_216# 0.03fF
C51729 OR2X1_LOC_769/B AND2X1_LOC_22/Y 0.17fF
C52068 AND2X1_LOC_22/Y OR2X1_LOC_139/A 0.03fF
C53236 AND2X1_LOC_22/Y AND2X1_LOC_497/a_36_24# 0.01fF
C53363 AND2X1_LOC_594/a_8_24# AND2X1_LOC_22/Y 0.02fF
C53450 AND2X1_LOC_22/Y OR2X1_LOC_668/a_8_216# 0.07fF
C53492 AND2X1_LOC_22/Y OR2X1_LOC_87/A 0.13fF
C54249 AND2X1_LOC_22/Y OR2X1_LOC_61/B 0.02fF
C54609 OR2X1_LOC_97/A AND2X1_LOC_22/Y 0.07fF
C55023 AND2X1_LOC_22/Y OR2X1_LOC_691/Y 0.06fF
C55573 AND2X1_LOC_22/Y OR2X1_LOC_720/A 0.08fF
C55612 AND2X1_LOC_22/Y OR2X1_LOC_333/B 0.01fF
C56017 OR2X1_LOC_154/A AND2X1_LOC_22/Y 0.25fF
C57870 AND2X1_LOC_22/Y VSS 0.72fF
C315 AND2X1_LOC_64/Y OR2X1_LOC_68/Y 0.03fF
C341 AND2X1_LOC_64/Y AND2X1_LOC_47/Y 0.57fF
C626 AND2X1_LOC_64/Y OR2X1_LOC_506/A 0.09fF
C795 AND2X1_LOC_64/Y OR2X1_LOC_227/Y 0.08fF
C1089 AND2X1_LOC_64/Y AND2X1_LOC_95/Y 0.73fF
C1114 AND2X1_LOC_64/Y OR2X1_LOC_99/Y 0.03fF
C1513 AND2X1_LOC_64/Y OR2X1_LOC_630/a_8_216# 0.01fF
C1518 AND2X1_LOC_64/Y OR2X1_LOC_664/a_8_216# 0.01fF
C1922 AND2X1_LOC_64/Y OR2X1_LOC_509/A 0.01fF
C2342 AND2X1_LOC_64/Y OR2X1_LOC_235/B 0.11fF
C2728 OR2X1_LOC_709/A AND2X1_LOC_64/Y 0.06fF
C2765 AND2X1_LOC_64/Y AND2X1_LOC_70/Y 0.70fF
C3172 AND2X1_LOC_64/Y OR2X1_LOC_362/A 0.22fF
C3501 AND2X1_LOC_64/Y OR2X1_LOC_771/B 0.03fF
C3524 AND2X1_LOC_64/Y OR2X1_LOC_776/A 0.03fF
C3935 AND2X1_LOC_64/Y OR2X1_LOC_593/B 0.01fF
C3959 OR2X1_LOC_506/a_8_216# AND2X1_LOC_64/Y 0.06fF
C4276 AND2X1_LOC_64/Y OR2X1_LOC_317/B 0.03fF
C4355 AND2X1_LOC_64/Y AND2X1_LOC_44/Y 0.98fF
C4916 AND2X1_LOC_64/Y AND2X1_LOC_69/Y 0.01fF
C4998 AND2X1_LOC_64/Y OR2X1_LOC_506/B 0.15fF
C5042 AND2X1_LOC_64/Y OR2X1_LOC_247/Y 0.01fF
C5204 AND2X1_LOC_64/Y AND2X1_LOC_18/Y 0.48fF
C5828 AND2X1_LOC_64/Y AND2X1_LOC_69/a_8_24# 0.02fF
C6098 AND2X1_LOC_64/Y AND2X1_LOC_65/a_8_24# 0.11fF
C6136 AND2X1_LOC_64/Y OR2X1_LOC_447/a_8_216# 0.09fF
C6145 AND2X1_LOC_64/Y OR2X1_LOC_130/A 0.03fF
C6593 AND2X1_LOC_64/Y OR2X1_LOC_449/B 0.06fF
C7817 AND2X1_LOC_64/Y OR2X1_LOC_786/A 0.03fF
C8021 AND2X1_LOC_64/Y OR2X1_LOC_447/Y 0.01fF
C8360 AND2X1_LOC_64/Y OR2X1_LOC_161/A 0.60fF
C8441 AND2X1_LOC_64/Y AND2X1_LOC_51/Y 10.19fF
C9151 AND2X1_LOC_64/Y AND2X1_LOC_41/A 1.61fF
C9219 AND2X1_LOC_64/Y OR2X1_LOC_631/B 0.06fF
C9876 AND2X1_LOC_64/Y OR2X1_LOC_704/a_8_216# 0.01fF
C10283 AND2X1_LOC_64/Y OR2X1_LOC_71/A 0.08fF
C10681 AND2X1_LOC_64/Y AND2X1_LOC_31/Y 1.54fF
C10910 AND2X1_LOC_64/Y OR2X1_LOC_633/B 0.03fF
C11063 AND2X1_LOC_64/Y OR2X1_LOC_608/Y 0.04fF
C11480 AND2X1_LOC_64/Y AND2X1_LOC_72/B 0.04fF
C11575 AND2X1_LOC_64/Y AND2X1_LOC_36/Y 2.36fF
C11626 OR2X1_LOC_506/Y AND2X1_LOC_64/Y 0.05fF
C11671 AND2X1_LOC_64/Y OR2X1_LOC_630/Y 0.16fF
C11717 AND2X1_LOC_64/Y AND2X1_LOC_586/a_8_24# 0.02fF
C12085 AND2X1_LOC_64/Y AND2X1_LOC_167/a_8_24# 0.04fF
C12175 AND2X1_LOC_64/Y OR2X1_LOC_592/a_8_216# 0.05fF
C12499 AND2X1_LOC_64/Y AND2X1_LOC_313/a_8_24# 0.01fF
C13015 AND2X1_LOC_64/Y AND2X1_LOC_504/a_8_24# 0.01fF
C13080 AND2X1_LOC_64/Y OR2X1_LOC_557/A 0.03fF
C13777 OR2X1_LOC_709/a_8_216# AND2X1_LOC_64/Y 0.02fF
C13833 AND2X1_LOC_64/Y AND2X1_LOC_312/a_36_24# 0.01fF
C13895 AND2X1_LOC_64/Y OR2X1_LOC_269/B 0.15fF
C14285 AND2X1_LOC_64/Y OR2X1_LOC_539/Y 0.09fF
C14575 AND2X1_LOC_64/Y OR2X1_LOC_319/Y 0.58fF
C14966 AND2X1_LOC_64/Y OR2X1_LOC_777/B 1.88fF
C15024 AND2X1_LOC_64/Y OR2X1_LOC_831/B 0.03fF
C15418 AND2X1_LOC_64/Y OR2X1_LOC_161/B 2.43fF
C16003 AND2X1_LOC_64/Y AND2X1_LOC_67/Y 0.02fF
C16563 AND2X1_LOC_64/Y OR2X1_LOC_705/B 0.01fF
C16844 AND2X1_LOC_64/Y AND2X1_LOC_72/a_8_24# 0.01fF
C16938 AND2X1_LOC_64/Y AND2X1_LOC_69/a_36_24# 0.01fF
C17201 AND2X1_LOC_64/Y OR2X1_LOC_201/A 0.01fF
C17273 AND2X1_LOC_64/Y AND2X1_LOC_3/Y 0.26fF
C17967 AND2X1_LOC_64/Y AND2X1_LOC_7/B 0.32fF
C18043 AND2X1_LOC_64/Y OR2X1_LOC_319/B 0.18fF
C18058 AND2X1_LOC_64/Y OR2X1_LOC_318/Y 7.13fF
C18135 AND2X1_LOC_64/Y OR2X1_LOC_296/Y 0.01fF
C18519 AND2X1_LOC_64/Y OR2X1_LOC_507/B 0.40fF
C18983 AND2X1_LOC_64/Y OR2X1_LOC_629/A 0.18fF
C19104 AND2X1_LOC_64/Y OR2X1_LOC_473/A 0.07fF
C19416 AND2X1_LOC_64/Y OR2X1_LOC_287/B 0.07fF
C19509 AND2X1_LOC_64/Y OR2X1_LOC_436/Y 0.03fF
C19738 AND2X1_LOC_64/Y OR2X1_LOC_160/B 0.18fF
C19823 AND2X1_LOC_64/Y OR2X1_LOC_799/a_8_216# 0.02fF
C20577 AND2X1_LOC_64/Y OR2X1_LOC_318/A 0.01fF
C20589 AND2X1_LOC_64/Y OR2X1_LOC_151/A 0.43fF
C20934 AND2X1_LOC_64/Y OR2X1_LOC_714/A 0.02fF
C23105 AND2X1_LOC_64/Y OR2X1_LOC_308/Y 1.80fF
C23545 AND2X1_LOC_64/Y OR2X1_LOC_828/Y 0.05fF
C23661 AND2X1_LOC_64/Y OR2X1_LOC_664/Y 0.01fF
C24827 OR2X1_LOC_711/B AND2X1_LOC_64/Y 0.01fF
C24850 AND2X1_LOC_64/Y OR2X1_LOC_324/B 0.03fF
C24880 AND2X1_LOC_64/Y AND2X1_LOC_142/a_8_24# 0.11fF
C24889 AND2X1_LOC_64/Y AND2X1_LOC_314/a_8_24# 0.14fF
C25326 AND2X1_LOC_64/Y OR2X1_LOC_799/a_36_216# 0.02fF
C25785 AND2X1_LOC_64/Y OR2X1_LOC_473/Y 0.45fF
C26126 AND2X1_LOC_64/Y AND2X1_LOC_423/a_8_24# 0.05fF
C26492 AND2X1_LOC_64/Y OR2X1_LOC_598/Y 0.03fF
C26499 AND2X1_LOC_64/Y AND2X1_LOC_131/a_8_24# 0.02fF
C26506 AND2X1_LOC_64/Y AND2X1_LOC_505/a_8_24# 0.01fF
C26541 AND2X1_LOC_64/Y AND2X1_LOC_40/Y 2.15fF
C26907 AND2X1_LOC_64/Y OR2X1_LOC_356/A 0.27fF
C27096 AND2X1_LOC_64/Y AND2X1_LOC_698/a_8_24# 0.04fF
C27443 AND2X1_LOC_64/Y OR2X1_LOC_810/A 0.06fF
C27757 OR2X1_LOC_715/B AND2X1_LOC_64/Y 0.07fF
C27863 AND2X1_LOC_64/Y AND2X1_LOC_81/a_8_24# 0.02fF
C28256 OR2X1_LOC_656/B AND2X1_LOC_64/Y 0.03fF
C28683 AND2X1_LOC_64/Y OR2X1_LOC_687/Y 0.23fF
C28750 AND2X1_LOC_64/Y OR2X1_LOC_401/B 0.29fF
C28990 AND2X1_LOC_64/Y AND2X1_LOC_829/a_8_24# 0.01fF
C29009 AND2X1_LOC_64/Y OR2X1_LOC_535/A 0.01fF
C29095 AND2X1_LOC_64/Y OR2X1_LOC_828/B 0.23fF
C29108 AND2X1_LOC_64/Y OR2X1_LOC_835/B 0.92fF
C29475 AND2X1_LOC_64/Y OR2X1_LOC_78/A 1.25fF
C30332 AND2X1_LOC_64/Y OR2X1_LOC_501/B 0.03fF
C30351 AND2X1_LOC_64/Y OR2X1_LOC_147/B 0.04fF
C30547 AND2X1_LOC_64/Y OR2X1_LOC_318/B 0.03fF
C30563 AND2X1_LOC_64/Y OR2X1_LOC_854/A 0.03fF
C30679 OR2X1_LOC_121/Y AND2X1_LOC_64/Y 0.07fF
C30697 AND2X1_LOC_64/Y OR2X1_LOC_114/B 0.06fF
C30732 AND2X1_LOC_64/Y OR2X1_LOC_538/A 0.03fF
C30791 AND2X1_LOC_12/Y AND2X1_LOC_64/Y 6.59fF
C30846 AND2X1_LOC_64/Y AND2X1_LOC_79/Y 4.54fF
C31176 AND2X1_LOC_64/Y OR2X1_LOC_168/B 0.20fF
C31223 AND2X1_LOC_64/Y AND2X1_LOC_59/Y 6.91fF
C31612 AND2X1_LOC_64/Y OR2X1_LOC_623/B 0.03fF
C31949 AND2X1_LOC_64/Y OR2X1_LOC_507/A 0.03fF
C31974 AND2X1_LOC_64/Y OR2X1_LOC_776/a_8_216# 0.03fF
C32019 AND2X1_LOC_64/Y OR2X1_LOC_254/B 0.15fF
C32421 AND2X1_LOC_64/Y AND2X1_LOC_321/a_8_24# 0.01fF
C33346 AND2X1_LOC_64/Y OR2X1_LOC_84/B 0.07fF
C33663 AND2X1_LOC_64/Y OR2X1_LOC_338/A 0.07fF
C33684 OR2X1_LOC_186/Y AND2X1_LOC_64/Y 0.34fF
C33759 AND2X1_LOC_64/Y AND2X1_LOC_81/B 0.09fF
C34194 AND2X1_LOC_64/Y OR2X1_LOC_574/A 8.03fF
C34201 AND2X1_LOC_64/Y OR2X1_LOC_33/A 0.10fF
C34457 AND2X1_LOC_64/Y OR2X1_LOC_855/A 0.15fF
C34465 AND2X1_LOC_64/Y AND2X1_LOC_627/a_8_24# 0.01fF
C34553 AND2X1_LOC_64/Y OR2X1_LOC_319/a_8_216# 0.06fF
C34980 AND2X1_LOC_64/Y OR2X1_LOC_78/B 0.77fF
C35026 AND2X1_LOC_64/Y OR2X1_LOC_375/A 0.13fF
C35305 AND2X1_LOC_64/Y OR2X1_LOC_843/B 0.16fF
C35315 AND2X1_LOC_64/Y OR2X1_LOC_549/A 0.18fF
C35470 AND2X1_LOC_64/Y OR2X1_LOC_629/a_8_216# 0.01fF
C36182 AND2X1_LOC_64/Y AND2X1_LOC_65/A 0.97fF
C37045 AND2X1_LOC_64/Y AND2X1_LOC_19/Y 0.07fF
C37063 AND2X1_LOC_64/Y AND2X1_LOC_316/a_8_24# 0.01fF
C37112 AND2X1_LOC_64/Y OR2X1_LOC_673/Y 0.07fF
C37420 OR2X1_LOC_335/A AND2X1_LOC_64/Y 0.01fF
C37837 AND2X1_LOC_64/Y OR2X1_LOC_139/A 0.98fF
C37919 AND2X1_LOC_64/Y OR2X1_LOC_324/A 0.01fF
C39002 AND2X1_LOC_64/Y OR2X1_LOC_247/a_8_216# 0.01fF
C39244 AND2X1_LOC_64/Y OR2X1_LOC_703/B 0.01fF
C39259 AND2X1_LOC_64/Y OR2X1_LOC_87/A 0.46fF
C39536 AND2X1_LOC_64/Y OR2X1_LOC_844/B 0.13fF
C39703 AND2X1_LOC_64/Y OR2X1_LOC_403/B 0.03fF
C40347 AND2X1_LOC_64/Y AND2X1_LOC_239/a_8_24# 0.01fF
C40399 AND2X1_LOC_64/Y OR2X1_LOC_97/A 0.06fF
C40453 OR2X1_LOC_302/B AND2X1_LOC_64/Y 0.08fF
C40484 AND2X1_LOC_64/Y OR2X1_LOC_475/B 0.57fF
C40821 AND2X1_LOC_64/Y OR2X1_LOC_691/Y 0.06fF
C40887 AND2X1_LOC_64/Y OR2X1_LOC_629/Y 0.19fF
C41359 AND2X1_LOC_64/Y AND2X1_LOC_314/a_36_24# 0.01fF
C41832 AND2X1_LOC_64/Y OR2X1_LOC_154/A 0.50fF
C42158 AND2X1_LOC_64/Y OR2X1_LOC_435/A 0.03fF
C42419 AND2X1_LOC_64/Y AND2X1_LOC_813/a_8_24# 0.03fF
C43092 AND2X1_LOC_64/Y OR2X1_LOC_776/a_36_216# 0.02fF
C43141 AND2X1_LOC_64/Y OR2X1_LOC_520/Y 0.05fF
C43214 AND2X1_LOC_64/Y AND2X1_LOC_107/a_8_24# 0.01fF
C43393 AND2X1_LOC_64/Y OR2X1_LOC_590/Y 0.10fF
C43954 AND2X1_LOC_64/Y OR2X1_LOC_756/B 0.26fF
C45340 AND2X1_LOC_64/Y OR2X1_LOC_33/B 0.03fF
C45686 OR2X1_LOC_100/Y AND2X1_LOC_64/Y 0.17fF
C45837 AND2X1_LOC_64/Y OR2X1_LOC_532/B 1.11fF
C45843 AND2X1_LOC_64/Y AND2X1_LOC_665/a_8_24# 0.01fF
C46539 AND2X1_LOC_64/Y OR2X1_LOC_729/a_8_216# 0.05fF
C46579 AND2X1_LOC_64/Y OR2X1_LOC_114/a_8_216# 0.01fF
C47050 AND2X1_LOC_64/Y AND2X1_LOC_503/a_8_24# 0.01fF
C47071 AND2X1_LOC_64/Y OR2X1_LOC_547/B 0.04fF
C47504 AND2X1_LOC_64/Y OR2X1_LOC_798/Y 0.01fF
C47837 AND2X1_LOC_64/Y OR2X1_LOC_502/Y 0.02fF
C47896 AND2X1_LOC_64/Y VDD 1.51fF
C48813 AND2X1_LOC_64/Y OR2X1_LOC_462/B 0.14fF
C48815 AND2X1_LOC_64/Y OR2X1_LOC_483/a_8_216# 0.01fF
C49059 AND2X1_LOC_64/Y AND2X1_LOC_591/a_8_24# 0.01fF
C49769 AND2X1_LOC_64/Y AND2X1_LOC_667/a_8_24# 0.11fF
C49963 AND2X1_LOC_64/Y OR2X1_LOC_115/B 1.34fF
C50056 AND2X1_LOC_64/Y OR2X1_LOC_840/A 0.29fF
C50472 AND2X1_LOC_64/Y OR2X1_LOC_216/A 0.74fF
C50918 AND2X1_LOC_64/Y OR2X1_LOC_160/A 0.49fF
C50964 AND2X1_LOC_64/Y OR2X1_LOC_624/B 0.07fF
C51317 AND2X1_LOC_64/Y OR2X1_LOC_447/A 0.09fF
C51714 AND2X1_LOC_64/Y OR2X1_LOC_78/Y 0.03fF
C52131 AND2X1_LOC_64/Y OR2X1_LOC_608/a_8_216# 0.01fF
C52148 AND2X1_LOC_64/Y OR2X1_LOC_185/A 0.59fF
C53366 AND2X1_LOC_64/Y OR2X1_LOC_641/A 0.03fF
C53397 AND2X1_LOC_64/Y AND2X1_LOC_312/a_8_24# 0.03fF
C53442 OR2X1_LOC_379/Y AND2X1_LOC_64/Y 0.03fF
C53472 AND2X1_LOC_64/Y OR2X1_LOC_114/Y 0.04fF
C54129 AND2X1_LOC_64/Y AND2X1_LOC_238/a_8_24# 0.01fF
C54225 AND2X1_LOC_64/Y OR2X1_LOC_637/A 0.03fF
C54281 AND2X1_LOC_64/Y OR2X1_LOC_643/A 0.18fF
C54284 AND2X1_LOC_64/Y OR2X1_LOC_778/Y 0.07fF
C54375 AND2X1_LOC_64/Y OR2X1_LOC_113/A 0.01fF
C54577 AND2X1_LOC_64/Y AND2X1_LOC_91/B 2.78fF
C54680 AND2X1_LOC_64/Y AND2X1_LOC_72/Y 0.01fF
C54681 AND2X1_LOC_64/Y OR2X1_LOC_799/A 4.36fF
C54926 AND2X1_LOC_64/Y OR2X1_LOC_446/B 0.70fF
C55029 AND2X1_LOC_64/Y OR2X1_LOC_719/B 0.22fF
C55123 AND2X1_LOC_64/Y AND2X1_LOC_56/B 11.23fF
C58014 AND2X1_LOC_64/Y VSS 0.61fF
C62 OR2X1_LOC_193/A AND2X1_LOC_3/Y 0.23fF
C207 AND2X1_LOC_3/Y OR2X1_LOC_339/A 1.32fF
C331 OR2X1_LOC_598/Y AND2X1_LOC_3/Y 0.04fF
C404 AND2X1_LOC_40/Y AND2X1_LOC_3/Y 0.20fF
C828 AND2X1_LOC_39/a_8_24# AND2X1_LOC_3/Y 0.01fF
C1355 OR2X1_LOC_810/A AND2X1_LOC_3/Y 0.03fF
C1633 OR2X1_LOC_715/B AND2X1_LOC_3/Y 0.47fF
C2167 OR2X1_LOC_656/B AND2X1_LOC_3/Y 1.15fF
C2180 AND2X1_LOC_767/a_8_24# AND2X1_LOC_3/Y 0.04fF
C2205 OR2X1_LOC_793/A AND2X1_LOC_3/Y 1.81fF
C2647 OR2X1_LOC_687/Y AND2X1_LOC_3/Y 0.03fF
C2700 OR2X1_LOC_401/B AND2X1_LOC_3/Y 0.01fF
C3402 AND2X1_LOC_3/Y OR2X1_LOC_78/A 5.41fF
C4195 OR2X1_LOC_501/B AND2X1_LOC_3/Y 0.03fF
C4224 OR2X1_LOC_147/B AND2X1_LOC_3/Y 0.02fF
C4238 AND2X1_LOC_517/a_8_24# AND2X1_LOC_3/Y 0.01fF
C4536 OR2X1_LOC_121/Y AND2X1_LOC_3/Y 0.08fF
C4573 OR2X1_LOC_114/B AND2X1_LOC_3/Y 0.06fF
C4586 AND2X1_LOC_396/a_8_24# AND2X1_LOC_3/Y 0.02fF
C4610 OR2X1_LOC_538/A AND2X1_LOC_3/Y 0.03fF
C4671 AND2X1_LOC_12/Y AND2X1_LOC_3/Y 1.25fF
C5082 AND2X1_LOC_59/Y AND2X1_LOC_3/Y 0.09fF
C5848 OR2X1_LOC_140/A AND2X1_LOC_3/Y 0.03fF
C5907 OR2X1_LOC_434/a_8_216# AND2X1_LOC_3/Y 0.04fF
C6630 AND2X1_LOC_3/Y AND2X1_LOC_248/a_8_24# 0.01fF
C7136 AND2X1_LOC_3/Y OR2X1_LOC_629/B 0.02fF
C7677 OR2X1_LOC_773/B AND2X1_LOC_3/Y 0.01fF
C7691 AND2X1_LOC_81/B AND2X1_LOC_3/Y 0.03fF
C7985 AND2X1_LOC_765/a_8_24# AND2X1_LOC_3/Y 0.02fF
C8179 OR2X1_LOC_574/A AND2X1_LOC_3/Y 0.03fF
C8442 AND2X1_LOC_3/Y AND2X1_LOC_627/a_8_24# 0.01fF
C8577 AND2X1_LOC_16/a_8_24# AND2X1_LOC_3/Y 0.10fF
C8925 AND2X1_LOC_3/Y OR2X1_LOC_78/B 1.04fF
C8989 OR2X1_LOC_375/A AND2X1_LOC_3/Y 0.31fF
C9301 AND2X1_LOC_3/Y OR2X1_LOC_549/A 0.12fF
C9484 OR2X1_LOC_629/a_8_216# AND2X1_LOC_3/Y 0.02fF
C9797 OR2X1_LOC_499/B AND2X1_LOC_3/Y 0.02fF
C10133 AND2X1_LOC_3/Y AND2X1_LOC_65/A 0.35fF
C11075 OR2X1_LOC_115/a_8_216# AND2X1_LOC_3/Y 0.01fF
C11107 OR2X1_LOC_673/Y AND2X1_LOC_3/Y 0.03fF
C11131 OR2X1_LOC_195/A AND2X1_LOC_3/Y 0.01fF
C11272 AND2X1_LOC_3/Y OR2X1_LOC_769/a_8_216# 0.01fF
C11722 AND2X1_LOC_3/Y OR2X1_LOC_712/B 0.09fF
C11791 OR2X1_LOC_139/A AND2X1_LOC_3/Y 0.10fF
C12944 OR2X1_LOC_247/a_8_216# AND2X1_LOC_3/Y 0.01fF
C13277 OR2X1_LOC_87/A AND2X1_LOC_3/Y 0.26fF
C13313 AND2X1_LOC_3/Y AND2X1_LOC_815/a_8_24# 0.07fF
C14096 OR2X1_LOC_194/B AND2X1_LOC_3/Y 0.01fF
C14355 OR2X1_LOC_97/A AND2X1_LOC_3/Y 0.03fF
C14451 AND2X1_LOC_3/Y OR2X1_LOC_78/a_8_216# 0.02fF
C14471 AND2X1_LOC_3/Y OR2X1_LOC_475/B 0.03fF
C14767 OR2X1_LOC_691/Y AND2X1_LOC_3/Y 0.05fF
C14784 AND2X1_LOC_3/Y OR2X1_LOC_713/A 0.01fF
C14901 OR2X1_LOC_629/Y AND2X1_LOC_3/Y 0.16fF
C15301 OR2X1_LOC_559/B AND2X1_LOC_3/Y 0.03fF
C15316 OR2X1_LOC_639/B AND2X1_LOC_3/Y 0.16fF
C15730 OR2X1_LOC_154/A AND2X1_LOC_3/Y 0.26fF
C15779 OR2X1_LOC_778/A AND2X1_LOC_3/Y 0.03fF
C15895 AND2X1_LOC_3/Y OR2X1_LOC_198/A 0.02fF
C16177 AND2X1_LOC_395/a_8_24# AND2X1_LOC_3/Y 0.02fF
C16463 AND2X1_LOC_3/Y OR2X1_LOC_361/a_8_216# 0.01fF
C16872 AND2X1_LOC_3/Y OR2X1_LOC_267/Y 0.03fF
C17043 OR2X1_LOC_520/Y AND2X1_LOC_3/Y 0.09fF
C17704 AND2X1_LOC_3/Y OR2X1_LOC_342/A 0.09fF
C17797 OR2X1_LOC_756/B AND2X1_LOC_3/Y 0.06fF
C18226 OR2X1_LOC_124/B AND2X1_LOC_3/Y 0.03fF
C18324 OR2X1_LOC_379/a_8_216# AND2X1_LOC_3/Y 0.01fF
C18626 OR2X1_LOC_614/Y AND2X1_LOC_3/Y 0.01fF
C19022 OR2X1_LOC_770/B AND2X1_LOC_3/Y 0.01fF
C19470 AND2X1_LOC_3/Y OR2X1_LOC_113/B 0.03fF
C19507 OR2X1_LOC_450/A AND2X1_LOC_3/Y 0.01fF
C19708 OR2X1_LOC_532/B AND2X1_LOC_3/Y 0.17fF
C19714 AND2X1_LOC_665/a_8_24# AND2X1_LOC_3/Y 0.04fF
C20302 OR2X1_LOC_855/a_8_216# AND2X1_LOC_3/Y 0.01fF
C21650 AND2X1_LOC_3/Y AND2X1_LOC_265/a_8_24# 0.01fF
C21665 VDD AND2X1_LOC_3/Y 1.04fF
C22317 AND2X1_LOC_3/Y AND2X1_LOC_418/a_8_24# 0.02fF
C22534 OR2X1_LOC_676/Y AND2X1_LOC_3/Y 0.09fF
C22563 OR2X1_LOC_834/A AND2X1_LOC_3/Y 0.42fF
C23703 AND2X1_LOC_3/Y OR2X1_LOC_115/B 0.51fF
C24235 AND2X1_LOC_397/a_8_24# AND2X1_LOC_3/Y 0.03fF
C24267 OR2X1_LOC_216/A AND2X1_LOC_3/Y 0.01fF
C24437 AND2X1_LOC_3/Y OR2X1_LOC_750/Y 0.05fF
C24701 OR2X1_LOC_160/A AND2X1_LOC_3/Y 0.27fF
C24764 OR2X1_LOC_624/B AND2X1_LOC_3/Y 0.03fF
C25195 AND2X1_LOC_127/a_8_24# AND2X1_LOC_3/Y 0.11fF
C25476 AND2X1_LOC_3/Y OR2X1_LOC_78/Y 0.02fF
C25923 OR2X1_LOC_185/A AND2X1_LOC_3/Y 0.06fF
C26406 OR2X1_LOC_702/A AND2X1_LOC_3/Y 0.03fF
C27104 AND2X1_LOC_3/Y OR2X1_LOC_294/Y 0.35fF
C27133 AND2X1_LOC_3/Y OR2X1_LOC_641/A 0.04fF
C27220 OR2X1_LOC_379/Y AND2X1_LOC_3/Y 0.59fF
C27255 OR2X1_LOC_114/Y AND2X1_LOC_3/Y 0.03fF
C27719 OR2X1_LOC_707/B AND2X1_LOC_3/Y 0.06fF
C27760 AND2X1_LOC_3/Y OR2X1_LOC_446/A 0.04fF
C28031 OR2X1_LOC_637/A AND2X1_LOC_3/Y 0.01fF
C28098 OR2X1_LOC_643/A AND2X1_LOC_3/Y 0.06fF
C28328 AND2X1_LOC_91/B AND2X1_LOC_3/Y 0.08fF
C28481 AND2X1_LOC_72/Y AND2X1_LOC_3/Y 0.01fF
C28776 AND2X1_LOC_3/Y OR2X1_LOC_719/B 0.22fF
C28807 OR2X1_LOC_542/B AND2X1_LOC_3/Y 0.03fF
C28876 OR2X1_LOC_631/a_8_216# AND2X1_LOC_3/Y 0.02fF
C28911 AND2X1_LOC_56/B AND2X1_LOC_3/Y 0.13fF
C29046 AND2X1_LOC_3/Y AND2X1_LOC_427/a_8_24# 0.02fF
C29672 OR2X1_LOC_402/B AND2X1_LOC_3/Y 0.01fF
C29903 AND2X1_LOC_3/Y AND2X1_LOC_751/a_8_24# 0.04fF
C30268 AND2X1_LOC_47/Y AND2X1_LOC_3/Y 2.45fF
C30579 AND2X1_LOC_695/a_8_24# AND2X1_LOC_3/Y 0.02fF
C30680 AND2X1_LOC_3/Y OR2X1_LOC_227/Y 0.02fF
C30683 AND2X1_LOC_3/Y OR2X1_LOC_284/B 0.01fF
C31016 AND2X1_LOC_95/Y AND2X1_LOC_3/Y 0.20fF
C31054 AND2X1_LOC_3/Y OR2X1_LOC_99/Y 0.25fF
C31214 AND2X1_LOC_3/Y AND2X1_LOC_41/Y 0.03fF
C31417 OR2X1_LOC_630/a_8_216# AND2X1_LOC_3/Y 0.01fF
C31533 AND2X1_LOC_3/Y OR2X1_LOC_434/A 0.44fF
C32180 OR2X1_LOC_235/B AND2X1_LOC_3/Y 0.03fF
C32395 AND2X1_LOC_3/Y OR2X1_LOC_779/B 0.45fF
C32562 OR2X1_LOC_709/A AND2X1_LOC_3/Y 0.35fF
C32566 AND2X1_LOC_3/Y AND2X1_LOC_295/a_8_24# 0.01fF
C32615 AND2X1_LOC_70/Y AND2X1_LOC_3/Y 2.36fF
C32688 AND2X1_LOC_380/a_8_24# AND2X1_LOC_3/Y 0.01fF
C32697 OR2X1_LOC_791/B AND2X1_LOC_3/Y 0.06fF
C32725 OR2X1_LOC_116/a_8_216# AND2X1_LOC_3/Y -0.00fF
C33007 AND2X1_LOC_3/Y OR2X1_LOC_362/A 0.01fF
C33100 OR2X1_LOC_116/A AND2X1_LOC_3/Y 0.01fF
C33308 AND2X1_LOC_3/Y OR2X1_LOC_771/B 0.04fF
C33524 OR2X1_LOC_637/B AND2X1_LOC_3/Y 0.01fF
C33806 AND2X1_LOC_766/a_8_24# AND2X1_LOC_3/Y 0.02fF
C34221 AND2X1_LOC_3/Y AND2X1_LOC_44/Y 2.83fF
C34446 AND2X1_LOC_3/Y OR2X1_LOC_720/B 0.03fF
C34870 AND2X1_LOC_3/Y OR2X1_LOC_793/B 0.03fF
C34938 OR2X1_LOC_506/B AND2X1_LOC_3/Y 0.14fF
C34970 OR2X1_LOC_247/Y AND2X1_LOC_3/Y 0.01fF
C35124 AND2X1_LOC_3/Y AND2X1_LOC_18/Y 0.38fF
C35353 AND2X1_LOC_3/Y OR2X1_LOC_789/A 0.03fF
C35534 AND2X1_LOC_3/Y OR2X1_LOC_307/A 0.74fF
C35773 AND2X1_LOC_3/Y AND2X1_LOC_428/a_8_24# 0.10fF
C36041 OR2X1_LOC_101/a_8_216# AND2X1_LOC_3/Y 0.01fF
C36047 OR2X1_LOC_231/A AND2X1_LOC_3/Y 0.03fF
C36071 OR2X1_LOC_707/A AND2X1_LOC_3/Y 0.04fF
C36073 OR2X1_LOC_130/A AND2X1_LOC_3/Y 1.33fF
C36092 AND2X1_LOC_292/a_8_24# AND2X1_LOC_3/Y 0.01fF
C36186 AND2X1_LOC_3/Y AND2X1_LOC_39/Y 0.06fF
C36475 AND2X1_LOC_487/a_8_24# AND2X1_LOC_3/Y 0.02fF
C36509 AND2X1_LOC_3/Y OR2X1_LOC_449/B 0.03fF
C38035 AND2X1_LOC_3/Y OR2X1_LOC_346/A 0.01fF
C38156 OR2X1_LOC_460/B AND2X1_LOC_3/Y 0.03fF
C38157 AND2X1_LOC_3/Y OR2X1_LOC_161/A 0.23fF
C38237 AND2X1_LOC_3/Y AND2X1_LOC_51/Y 0.12fF
C38598 AND2X1_LOC_3/Y AND2X1_LOC_297/a_8_24# 0.01fF
C38997 AND2X1_LOC_41/A AND2X1_LOC_3/Y 2.06fF
C39079 OR2X1_LOC_631/B AND2X1_LOC_3/Y 0.06fF
C39883 OR2X1_LOC_632/A AND2X1_LOC_3/Y 0.02fF
C40405 OR2X1_LOC_614/a_8_216# AND2X1_LOC_3/Y 0.02fF
C40459 AND2X1_LOC_3/Y AND2X1_LOC_31/Y 1.40fF
C41148 AND2X1_LOC_305/a_8_24# AND2X1_LOC_3/Y 0.10fF
C41250 OR2X1_LOC_288/A AND2X1_LOC_3/Y 0.08fF
C41291 AND2X1_LOC_3/Y AND2X1_LOC_72/B 0.03fF
C41296 AND2X1_LOC_3/Y OR2X1_LOC_451/B 0.24fF
C41375 AND2X1_LOC_3/Y AND2X1_LOC_36/Y 1.03fF
C41535 OR2X1_LOC_630/Y AND2X1_LOC_3/Y 0.01fF
C41572 OR2X1_LOC_635/A AND2X1_LOC_3/Y 0.06fF
C41599 AND2X1_LOC_586/a_8_24# AND2X1_LOC_3/Y 0.01fF
C41649 OR2X1_LOC_346/B AND2X1_LOC_3/Y 0.01fF
C41671 AND2X1_LOC_122/a_8_24# AND2X1_LOC_3/Y 0.01fF
C42347 OR2X1_LOC_856/A AND2X1_LOC_3/Y 0.01fF
C42959 OR2X1_LOC_557/A AND2X1_LOC_3/Y 0.94fF
C43326 OR2X1_LOC_814/Y AND2X1_LOC_3/Y 0.12fF
C43817 AND2X1_LOC_3/Y OR2X1_LOC_269/B 3.84fF
C43837 OR2X1_LOC_460/a_8_216# AND2X1_LOC_3/Y 0.01fF
C44212 AND2X1_LOC_3/Y OR2X1_LOC_347/B 0.01fF
C44216 AND2X1_LOC_3/Y OR2X1_LOC_539/Y 0.03fF
C44549 AND2X1_LOC_184/a_8_24# AND2X1_LOC_3/Y 0.01fF
C44841 AND2X1_LOC_3/Y OR2X1_LOC_777/B 0.03fF
C44903 OR2X1_LOC_770/A AND2X1_LOC_3/Y 0.01fF
C45368 AND2X1_LOC_3/Y OR2X1_LOC_161/B 2.57fF
C45534 OR2X1_LOC_460/Y AND2X1_LOC_3/Y 0.01fF
C45702 AND2X1_LOC_3/Y OR2X1_LOC_707/a_8_216# 0.06fF
C45880 AND2X1_LOC_3/Y OR2X1_LOC_630/B 0.02fF
C46861 AND2X1_LOC_3/Y AND2X1_LOC_230/a_8_24# 0.02fF
C46895 AND2X1_LOC_72/a_8_24# AND2X1_LOC_3/Y 0.02fF
C47172 AND2X1_LOC_3/Y OR2X1_LOC_489/A 0.01fF
C47820 OR2X1_LOC_401/A AND2X1_LOC_3/Y 0.56fF
C48037 AND2X1_LOC_3/Y AND2X1_LOC_7/B 5.25fF
C48249 OR2X1_LOC_296/Y AND2X1_LOC_3/Y 0.03fF
C49054 OR2X1_LOC_629/A AND2X1_LOC_3/Y 0.18fF
C49099 OR2X1_LOC_446/Y AND2X1_LOC_3/Y 0.04fF
C49120 OR2X1_LOC_473/A AND2X1_LOC_3/Y 0.78fF
C49443 OR2X1_LOC_635/a_8_216# AND2X1_LOC_3/Y 0.01fF
C49503 OR2X1_LOC_287/B AND2X1_LOC_3/Y 0.04fF
C49797 OR2X1_LOC_160/B AND2X1_LOC_3/Y 1.18fF
C50601 OR2X1_LOC_151/A AND2X1_LOC_3/Y 0.07fF
C51000 AND2X1_LOC_3/Y AND2X1_LOC_279/a_8_24# 0.01fF
C51059 OR2X1_LOC_287/A AND2X1_LOC_3/Y 0.80fF
C51079 OR2X1_LOC_174/A AND2X1_LOC_3/Y 0.05fF
C51874 AND2X1_LOC_3/Y OR2X1_LOC_631/A 0.03fF
C53694 OR2X1_LOC_664/Y AND2X1_LOC_3/Y 0.05fF
C54103 OR2X1_LOC_446/a_8_216# AND2X1_LOC_3/Y 0.01fF
C54158 AND2X1_LOC_3/Y AND2X1_LOC_7/Y 0.03fF
C54355 AND2X1_LOC_3/Y OR2X1_LOC_390/A 0.03fF
C55690 OR2X1_LOC_190/A AND2X1_LOC_3/Y 0.01fF
C56880 AND2X1_LOC_3/Y VSS 0.68fF
C405 AND2X1_LOC_40/Y OR2X1_LOC_647/B 0.78fF
C1082 AND2X1_LOC_40/Y AND2X1_LOC_7/B 0.20fF
C1214 AND2X1_LOC_40/Y OR2X1_LOC_318/Y 0.03fF
C1325 AND2X1_LOC_40/Y OR2X1_LOC_436/a_8_216# 0.01fF
C1357 AND2X1_LOC_40/Y AND2X1_LOC_441/a_8_24# 0.04fF
C2678 AND2X1_LOC_40/Y OR2X1_LOC_436/Y 0.10fF
C2869 AND2X1_LOC_40/Y OR2X1_LOC_160/B 0.38fF
C2976 AND2X1_LOC_40/Y OR2X1_LOC_553/A 0.09fF
C3683 AND2X1_LOC_40/Y OR2X1_LOC_151/A 0.32fF
C3707 AND2X1_LOC_40/Y AND2X1_LOC_41/a_36_24# 0.01fF
C4123 AND2X1_LOC_40/Y OR2X1_LOC_174/A 0.01fF
C4127 AND2X1_LOC_40/Y OR2X1_LOC_435/a_8_216# 0.01fF
C4906 AND2X1_LOC_40/Y AND2X1_LOC_616/a_8_24# 0.01fF
C5071 AND2X1_LOC_40/Y OR2X1_LOC_285/B 0.17fF
C5232 AND2X1_LOC_40/Y OR2X1_LOC_168/Y 0.07fF
C5422 AND2X1_LOC_394/a_36_24# AND2X1_LOC_40/Y 0.01fF
C6295 AND2X1_LOC_40/Y OR2X1_LOC_593/A 0.01fF
C6489 AND2X1_LOC_40/Y OR2X1_LOC_535/a_36_216# -0.00fF
C6537 AND2X1_LOC_40/Y OR2X1_LOC_828/Y 0.01fF
C7009 AND2X1_LOC_40/Y OR2X1_LOC_61/A 0.13fF
C7274 AND2X1_LOC_40/Y AND2X1_LOC_7/Y 0.03fF
C7480 AND2X1_LOC_40/Y OR2X1_LOC_390/A 0.07fF
C8256 AND2X1_LOC_40/Y OR2X1_LOC_344/a_8_216# 0.01fF
C8646 AND2X1_LOC_40/Y OR2X1_LOC_84/A 0.23fF
C8816 AND2X1_LOC_40/Y OR2X1_LOC_190/A 1.00fF
C9235 AND2X1_LOC_40/Y OR2X1_LOC_325/B 0.03fF
C9280 AND2X1_LOC_40/Y AND2X1_LOC_189/a_8_24# 0.17fF
C9293 AND2X1_LOC_40/Y OR2X1_LOC_285/a_8_216# 0.01fF
C9564 AND2X1_LOC_40/Y OR2X1_LOC_339/A 0.12fF
C9629 AND2X1_LOC_40/Y OR2X1_LOC_673/B 0.03fF
C9643 AND2X1_LOC_40/Y OR2X1_LOC_831/A 0.03fF
C9657 AND2X1_LOC_40/Y OR2X1_LOC_598/Y 0.01fF
C9659 AND2X1_LOC_40/Y AND2X1_LOC_505/a_8_24# 0.10fF
C9695 OR2X1_LOC_335/Y AND2X1_LOC_40/Y 0.03fF
C10460 AND2X1_LOC_40/Y AND2X1_LOC_258/a_36_24# 0.01fF
C10638 AND2X1_LOC_40/Y OR2X1_LOC_810/A 0.03fF
C10662 AND2X1_LOC_40/Y AND2X1_LOC_589/a_8_24# 0.01fF
C10894 OR2X1_LOC_715/B AND2X1_LOC_40/Y 0.01fF
C11180 AND2X1_LOC_40/Y OR2X1_LOC_398/Y 0.03fF
C11413 OR2X1_LOC_656/B AND2X1_LOC_40/Y 0.08fF
C12117 AND2X1_LOC_40/Y AND2X1_LOC_829/a_8_24# 0.01fF
C12297 AND2X1_LOC_40/Y OR2X1_LOC_828/B 0.04fF
C12628 AND2X1_LOC_40/Y OR2X1_LOC_78/A 0.20fF
C13547 AND2X1_LOC_40/Y OR2X1_LOC_147/B 0.06fF
C13623 AND2X1_LOC_40/Y OR2X1_LOC_383/a_8_216# 0.01fF
C13628 AND2X1_LOC_40/Y AND2X1_LOC_171/a_8_24# 0.14fF
C13697 AND2X1_LOC_40/Y OR2X1_LOC_545/B 0.31fF
C13745 AND2X1_LOC_40/Y OR2X1_LOC_318/B 0.03fF
C13755 AND2X1_LOC_40/Y OR2X1_LOC_854/A 0.01fF
C13767 AND2X1_LOC_40/Y OR2X1_LOC_344/a_36_216# 0.02fF
C14012 AND2X1_LOC_12/Y AND2X1_LOC_40/Y 1.34fF
C14427 AND2X1_LOC_40/Y AND2X1_LOC_59/Y 1.88fF
C15186 AND2X1_LOC_40/Y OR2X1_LOC_434/a_8_216# 0.01fF
C15238 AND2X1_LOC_40/Y OR2X1_LOC_254/B 0.55fF
C15268 AND2X1_LOC_40/Y OR2X1_LOC_646/A 0.01fF
C16142 AND2X1_LOC_40/Y OR2X1_LOC_592/A 0.01fF
C16544 AND2X1_LOC_40/Y OR2X1_LOC_84/B 0.47fF
C16808 OR2X1_LOC_186/Y AND2X1_LOC_40/Y 0.49fF
C16974 AND2X1_LOC_40/Y AND2X1_LOC_81/B 0.05fF
C17092 AND2X1_LOC_40/Y OR2X1_LOC_112/B 0.02fF
C17404 AND2X1_LOC_40/Y OR2X1_LOC_574/A 0.03fF
C17610 AND2X1_LOC_40/Y OR2X1_LOC_855/A 0.01fF
C17849 AND2X1_LOC_40/Y AND2X1_LOC_670/a_8_24# 0.04fF
C18017 AND2X1_LOC_40/Y OR2X1_LOC_539/B 0.02fF
C18150 AND2X1_LOC_40/Y OR2X1_LOC_78/B 0.91fF
C18239 AND2X1_LOC_40/Y OR2X1_LOC_375/A 6.37fF
C18539 AND2X1_LOC_40/Y OR2X1_LOC_549/A 0.08fF
C19281 AND2X1_LOC_40/Y OR2X1_LOC_348/B 0.09fF
C19397 AND2X1_LOC_40/Y AND2X1_LOC_65/A 0.55fF
C19491 AND2X1_LOC_40/Y OR2X1_LOC_181/B 0.02fF
C20047 AND2X1_LOC_40/Y OR2X1_LOC_285/Y 0.01fF
C20398 AND2X1_LOC_40/Y OR2X1_LOC_673/Y 0.07fF
C20700 AND2X1_LOC_40/Y OR2X1_LOC_676/a_8_216# 0.01fF
C20729 OR2X1_LOC_769/B AND2X1_LOC_40/Y 0.01fF
C21078 AND2X1_LOC_40/Y OR2X1_LOC_139/A 0.03fF
C21082 AND2X1_LOC_40/Y OR2X1_LOC_758/a_8_216# 0.04fF
C21177 AND2X1_LOC_40/Y OR2X1_LOC_637/Y 0.09fF
C22395 AND2X1_LOC_594/a_8_24# AND2X1_LOC_40/Y 0.01fF
C22558 OR2X1_LOC_703/B AND2X1_LOC_40/Y 0.02fF
C22569 AND2X1_LOC_40/Y OR2X1_LOC_87/A 0.59fF
C22890 AND2X1_LOC_40/Y OR2X1_LOC_389/A 0.25fF
C22930 AND2X1_LOC_40/Y AND2X1_LOC_177/a_8_24# 0.01fF
C23347 AND2X1_LOC_40/Y OR2X1_LOC_61/B 0.02fF
C23509 AND2X1_LOC_40/Y AND2X1_LOC_441/a_36_24# 0.01fF
C23648 AND2X1_LOC_40/Y OR2X1_LOC_97/A 0.05fF
C23919 AND2X1_LOC_40/Y AND2X1_LOC_613/a_8_24# 0.04fF
C24081 AND2X1_LOC_40/Y OR2X1_LOC_691/Y 0.02fF
C24673 AND2X1_LOC_40/Y OR2X1_LOC_333/B 0.04fF
C25038 OR2X1_LOC_154/A AND2X1_LOC_40/Y 0.40fF
C25225 AND2X1_LOC_40/Y OR2X1_LOC_198/A 0.02fF
C26812 AND2X1_LOC_40/Y AND2X1_LOC_600/a_8_24# 0.04fF
C27086 AND2X1_LOC_40/Y OR2X1_LOC_756/B 0.76fF
C27842 OR2X1_LOC_653/B AND2X1_LOC_40/Y 0.01fF
C28762 OR2X1_LOC_100/Y AND2X1_LOC_40/Y 0.04fF
C28796 AND2X1_LOC_40/Y OR2X1_LOC_286/Y 0.02fF
C28928 AND2X1_LOC_40/Y OR2X1_LOC_532/B 0.26fF
C29139 AND2X1_LOC_40/Y OR2X1_LOC_440/B 0.05fF
C29189 AND2X1_LOC_531/a_8_24# AND2X1_LOC_40/Y 0.04fF
C29786 AND2X1_LOC_40/Y OR2X1_LOC_286/B 0.03fF
C30055 AND2X1_LOC_40/Y AND2X1_LOC_503/a_8_24# 0.01fF
C30146 AND2X1_LOC_40/Y AND2X1_LOC_171/a_36_24# 0.01fF
C30659 AND2X1_LOC_40/Y OR2X1_LOC_192/B 0.04fF
C30751 AND2X1_LOC_40/Y OR2X1_LOC_502/Y 0.31fF
C30828 AND2X1_LOC_40/Y AND2X1_LOC_265/a_8_24# 0.03fF
C30843 AND2X1_LOC_40/Y VDD 2.84fF
C31044 AND2X1_LOC_40/Y OR2X1_LOC_444/B 0.05fF
C31675 AND2X1_LOC_40/Y OR2X1_LOC_676/Y 0.08fF
C32027 AND2X1_LOC_40/Y AND2X1_LOC_83/a_8_24# 0.02fF
C32985 AND2X1_LOC_40/Y OR2X1_LOC_840/A 0.03fF
C33671 AND2X1_LOC_40/Y OR2X1_LOC_750/Y 0.01fF
C33897 OR2X1_LOC_160/A AND2X1_LOC_40/Y 7.90fF
C33946 AND2X1_LOC_40/Y AND2X1_LOC_86/B 0.03fF
C33953 AND2X1_LOC_40/Y OR2X1_LOC_624/B 0.09fF
C34666 AND2X1_LOC_40/Y OR2X1_LOC_190/B 0.29fF
C35103 AND2X1_LOC_40/Y OR2X1_LOC_608/a_8_216# 0.19fF
C35127 AND2X1_LOC_40/Y OR2X1_LOC_185/A 0.51fF
C35195 AND2X1_LOC_40/Y OR2X1_LOC_435/Y 0.01fF
C35239 AND2X1_LOC_40/Y AND2X1_LOC_431/a_8_24# 0.01fF
C35402 AND2X1_LOC_40/Y OR2X1_LOC_550/A 0.11fF
C35909 AND2X1_LOC_40/Y AND2X1_LOC_437/a_8_24# 0.01fF
C36031 AND2X1_LOC_40/Y AND2X1_LOC_481/a_8_24# 0.05fF
C36066 AND2X1_LOC_40/Y AND2X1_LOC_442/a_8_24# 0.01fF
C36268 AND2X1_LOC_40/Y OR2X1_LOC_294/Y 0.06fF
C36298 AND2X1_LOC_40/Y OR2X1_LOC_641/A 0.03fF
C36507 AND2X1_LOC_40/Y OR2X1_LOC_286/a_8_216# 0.01fF
C36798 AND2X1_LOC_40/Y AND2X1_LOC_617/a_8_24# 0.01fF
C37191 AND2X1_LOC_40/Y OR2X1_LOC_436/B 0.01fF
C37269 AND2X1_LOC_40/Y OR2X1_LOC_778/Y 0.07fF
C37510 AND2X1_LOC_91/B AND2X1_LOC_40/Y 5.95fF
C37645 AND2X1_LOC_40/Y OR2X1_LOC_799/A 0.08fF
C37771 AND2X1_LOC_40/Y AND2X1_LOC_600/a_36_24# 0.01fF
C37861 AND2X1_LOC_40/Y OR2X1_LOC_303/B 0.03fF
C37980 AND2X1_LOC_40/Y OR2X1_LOC_542/B 0.03fF
C38088 AND2X1_LOC_40/Y AND2X1_LOC_56/B 1.10fF
C38507 AND2X1_LOC_40/Y AND2X1_LOC_166/a_8_24# 0.03fF
C38575 AND2X1_LOC_40/Y AND2X1_LOC_183/a_8_24# 0.23fF
C39004 AND2X1_LOC_40/Y OR2X1_LOC_389/B 0.06fF
C39010 AND2X1_LOC_40/Y AND2X1_LOC_118/a_8_24# 0.07fF
C39264 AND2X1_LOC_745/a_8_24# AND2X1_LOC_40/Y 0.09fF
C39518 AND2X1_LOC_40/Y AND2X1_LOC_47/Y 0.26fF
C39697 AND2X1_LOC_40/Y OR2X1_LOC_646/B 0.35fF
C39761 AND2X1_LOC_40/Y OR2X1_LOC_828/a_8_216# 0.01fF
C39800 AND2X1_LOC_40/Y OR2X1_LOC_506/A 0.03fF
C40011 AND2X1_LOC_40/Y OR2X1_LOC_180/B 0.07fF
C40169 AND2X1_LOC_40/Y AND2X1_LOC_95/Y 2.37fF
C40175 AND2X1_LOC_40/Y OR2X1_LOC_633/Y 0.10fF
C40436 AND2X1_LOC_40/Y OR2X1_LOC_788/B 0.04fF
C40529 AND2X1_LOC_40/Y OR2X1_LOC_621/A 0.22fF
C40757 AND2X1_LOC_40/Y OR2X1_LOC_434/A 0.01fF
C41039 AND2X1_LOC_40/Y OR2X1_LOC_509/A 0.01fF
C41453 AND2X1_LOC_40/Y OR2X1_LOC_235/B 0.07fF
C41545 AND2X1_LOC_393/a_8_24# AND2X1_LOC_40/Y 0.05fF
C41870 AND2X1_LOC_40/Y AND2X1_LOC_70/Y 0.20fF
C41899 AND2X1_LOC_40/Y OR2X1_LOC_703/A 0.03fF
C41949 OR2X1_LOC_791/B AND2X1_LOC_40/Y 0.03fF
C42641 AND2X1_LOC_40/Y OR2X1_LOC_771/B 0.05fF
C42649 AND2X1_LOC_40/Y OR2X1_LOC_209/A 0.03fF
C42800 AND2X1_LOC_40/Y OR2X1_LOC_637/B 0.03fF
C43073 AND2X1_LOC_40/Y OR2X1_LOC_593/B 0.03fF
C43158 AND2X1_LOC_40/Y AND2X1_LOC_41/a_8_24# 0.12fF
C43335 AND2X1_LOC_40/Y OR2X1_LOC_254/a_8_216# 0.01fF
C43551 AND2X1_LOC_40/Y AND2X1_LOC_44/Y 2.93fF
C44393 AND2X1_LOC_40/Y AND2X1_LOC_258/a_8_24# 0.05fF
C44456 AND2X1_LOC_40/Y AND2X1_LOC_18/Y 1.06fF
C44579 OR2X1_LOC_596/Y AND2X1_LOC_40/Y 0.01fF
C44716 AND2X1_LOC_40/Y AND2X1_LOC_485/a_8_24# 0.03fF
C45001 AND2X1_LOC_394/a_8_24# AND2X1_LOC_40/Y 0.03fF
C45436 AND2X1_LOC_40/Y OR2X1_LOC_130/A 0.07fF
C45894 AND2X1_LOC_40/Y OR2X1_LOC_449/B 0.03fF
C46199 AND2X1_LOC_40/Y OR2X1_LOC_621/B 0.23fF
C46431 AND2X1_LOC_40/Y OR2X1_LOC_383/Y 0.10fF
C47091 AND2X1_LOC_40/Y OR2X1_LOC_389/a_8_216# 0.14fF
C47581 AND2X1_LOC_40/Y AND2X1_LOC_265/a_36_24# 0.01fF
C47671 AND2X1_LOC_40/Y OR2X1_LOC_161/A 0.11fF
C47755 AND2X1_LOC_40/Y AND2X1_LOC_51/Y 0.18fF
C48427 AND2X1_LOC_40/Y OR2X1_LOC_439/B 0.03fF
C48487 AND2X1_LOC_40/Y AND2X1_LOC_41/A 0.87fF
C48560 AND2X1_LOC_40/Y OR2X1_LOC_631/B 0.42fF
C48888 AND2X1_LOC_40/Y AND2X1_LOC_253/a_8_24# 0.01fF
C49593 AND2X1_LOC_40/Y OR2X1_LOC_71/A 0.03fF
C49827 AND2X1_LOC_40/Y OR2X1_LOC_593/a_8_216# 0.01fF
C49987 AND2X1_LOC_40/Y AND2X1_LOC_31/Y 0.17fF
C50236 AND2X1_LOC_597/a_8_24# AND2X1_LOC_40/Y 0.18fF
C50263 AND2X1_LOC_40/Y OR2X1_LOC_633/B 0.05fF
C50413 AND2X1_LOC_40/Y OR2X1_LOC_608/Y 0.37fF
C50810 AND2X1_LOC_40/Y AND2X1_LOC_72/B 0.31fF
C50883 AND2X1_LOC_40/Y AND2X1_LOC_36/Y 1.80fF
C51491 AND2X1_LOC_40/Y OR2X1_LOC_592/a_8_216# 0.01fF
C51695 AND2X1_LOC_40/Y OR2X1_LOC_535/a_8_216# 0.01fF
C52149 AND2X1_LOC_40/Y AND2X1_LOC_60/a_8_24# 0.17fF
C52766 AND2X1_LOC_393/a_36_24# AND2X1_LOC_40/Y 0.01fF
C52793 AND2X1_LOC_40/Y AND2X1_LOC_481/a_36_24# 0.01fF
C53168 AND2X1_LOC_40/Y OR2X1_LOC_798/a_8_216# 0.04fF
C53186 AND2X1_LOC_40/Y OR2X1_LOC_269/B 2.37fF
C53674 AND2X1_LOC_40/Y AND2X1_LOC_176/a_8_24# 0.04fF
C53958 AND2X1_LOC_40/Y OR2X1_LOC_637/a_8_216# 0.01fF
C54191 AND2X1_LOC_40/Y OR2X1_LOC_777/B 10.58fF
C54262 AND2X1_LOC_40/Y OR2X1_LOC_344/A 0.09fF
C54358 AND2X1_LOC_40/Y OR2X1_LOC_254/A 0.01fF
C54479 AND2X1_LOC_40/Y OR2X1_LOC_456/A 0.14fF
C54686 AND2X1_LOC_40/Y OR2X1_LOC_161/B 0.35fF
C55727 OR2X1_LOC_644/B AND2X1_LOC_40/Y 0.01fF
C55891 AND2X1_LOC_40/Y AND2X1_LOC_609/a_8_24# 0.01fF
C57900 AND2X1_LOC_40/Y VSS 1.37fF
C166 AND2X1_LOC_70/Y OR2X1_LOC_691/Y 0.05fF
C724 AND2X1_LOC_70/Y OR2X1_LOC_639/B 0.01fF
C790 OR2X1_LOC_333/B AND2X1_LOC_70/Y 0.06fF
C1198 OR2X1_LOC_154/A AND2X1_LOC_70/Y 0.26fF
C1265 AND2X1_LOC_70/Y OR2X1_LOC_778/A 0.01fF
C1399 AND2X1_LOC_70/Y OR2X1_LOC_198/A 0.17fF
C1498 AND2X1_LOC_70/Y OR2X1_LOC_435/A 0.26fF
C1743 AND2X1_LOC_70/Y AND2X1_LOC_821/a_8_24# 0.11fF
C1988 OR2X1_LOC_538/a_8_216# AND2X1_LOC_70/Y 0.01fF
C3034 AND2X1_LOC_70/Y AND2X1_LOC_600/a_8_24# 0.01fF
C3286 OR2X1_LOC_756/B AND2X1_LOC_70/Y 1.42fF
C3633 AND2X1_LOC_70/Y OR2X1_LOC_355/A 0.01fF
C3665 OR2X1_LOC_124/B AND2X1_LOC_70/Y 0.05fF
C4058 OR2X1_LOC_614/Y AND2X1_LOC_70/Y 0.01fF
C5068 AND2X1_LOC_70/Y OR2X1_LOC_532/B 2.58fF
C5677 AND2X1_LOC_70/Y OR2X1_LOC_855/a_8_216# 0.01fF
C6430 AND2X1_LOC_70/Y AND2X1_LOC_432/a_8_24# 0.02fF
C7014 VDD AND2X1_LOC_70/Y 1.07fF
C7720 AND2X1_LOC_70/Y AND2X1_LOC_418/a_8_24# 0.01fF
C8583 AND2X1_LOC_70/Y OR2X1_LOC_602/B 0.01fF
C8974 AND2X1_LOC_70/Y AND2X1_LOC_667/a_8_24# 0.01fF
C9243 AND2X1_LOC_70/Y OR2X1_LOC_840/A 0.03fF
C9672 AND2X1_LOC_70/Y OR2X1_LOC_216/A 0.01fF
C9922 AND2X1_LOC_70/Y OR2X1_LOC_750/Y 0.15fF
C10045 AND2X1_LOC_70/Y OR2X1_LOC_809/B 0.24fF
C10081 AND2X1_LOC_70/Y AND2X1_LOC_177/a_36_24# 0.01fF
C10125 OR2X1_LOC_160/A AND2X1_LOC_70/Y 0.22fF
C10364 AND2X1_LOC_70/Y OR2X1_LOC_532/Y 0.09fF
C10841 AND2X1_LOC_91/a_36_24# AND2X1_LOC_70/Y 0.01fF
C11367 AND2X1_LOC_70/Y OR2X1_LOC_185/A 0.10fF
C11511 AND2X1_LOC_70/Y AND2X1_LOC_431/a_8_24# 0.09fF
C11872 OR2X1_LOC_702/A AND2X1_LOC_70/Y 0.03fF
C12120 AND2X1_LOC_70/Y AND2X1_LOC_262/a_8_24# 0.01fF
C12544 AND2X1_LOC_70/Y OR2X1_LOC_294/Y 0.01fF
C12560 AND2X1_LOC_70/Y OR2X1_LOC_641/A 0.03fF
C12655 OR2X1_LOC_379/Y AND2X1_LOC_70/Y 0.02fF
C13119 AND2X1_LOC_70/Y OR2X1_LOC_541/B 0.08fF
C13304 AND2X1_LOC_70/Y OR2X1_LOC_446/A 0.01fF
C13488 AND2X1_LOC_70/Y OR2X1_LOC_637/A 0.01fF
C13563 AND2X1_LOC_70/Y OR2X1_LOC_643/A 0.03fF
C13572 AND2X1_LOC_70/Y OR2X1_LOC_778/Y 0.03fF
C13807 AND2X1_LOC_91/B AND2X1_LOC_70/Y 0.35fF
C14191 AND2X1_LOC_70/Y OR2X1_LOC_446/B 0.02fF
C14197 AND2X1_LOC_70/Y OR2X1_LOC_303/B 0.06fF
C14267 AND2X1_LOC_70/Y OR2X1_LOC_719/B 0.10fF
C14399 AND2X1_LOC_70/Y AND2X1_LOC_56/B 1.47fF
C15217 OR2X1_LOC_389/B AND2X1_LOC_70/Y 0.02fF
C15722 AND2X1_LOC_70/Y AND2X1_LOC_47/Y 3.37fF
C16025 AND2X1_LOC_70/Y OR2X1_LOC_506/A 0.02fF
C16298 AND2X1_LOC_70/Y OR2X1_LOC_180/B 0.03fF
C16434 AND2X1_LOC_70/Y AND2X1_LOC_95/Y 1.30fF
C18052 OR2X1_LOC_709/A AND2X1_LOC_70/Y 0.04fF
C18122 AND2X1_LOC_70/Y OR2X1_LOC_703/A 0.03fF
C18209 OR2X1_LOC_116/a_8_216# AND2X1_LOC_70/Y 0.01fF
C18526 AND2X1_LOC_70/Y OR2X1_LOC_832/a_8_216# 0.01fF
C18568 OR2X1_LOC_539/A AND2X1_LOC_70/Y 0.01fF
C18613 OR2X1_LOC_116/A AND2X1_LOC_70/Y 0.01fF
C18874 AND2X1_LOC_70/Y OR2X1_LOC_771/B 0.03fF
C19289 AND2X1_LOC_70/Y OR2X1_LOC_593/B 2.91fF
C19779 AND2X1_LOC_70/Y AND2X1_LOC_44/Y 1.74fF
C20023 AND2X1_LOC_70/Y OR2X1_LOC_720/B -0.00fF
C20506 AND2X1_LOC_70/Y OR2X1_LOC_247/Y 0.09fF
C20668 AND2X1_LOC_70/Y AND2X1_LOC_18/Y 3.98fF
C21390 AND2X1_LOC_70/Y AND2X1_LOC_428/a_8_24# 0.01fF
C21639 AND2X1_LOC_70/Y OR2X1_LOC_130/A 0.98fF
C22120 AND2X1_LOC_70/Y OR2X1_LOC_636/A 0.01fF
C22973 AND2X1_LOC_70/Y OR2X1_LOC_355/B 0.03fF
C23003 AND2X1_LOC_70/Y AND2X1_LOC_674/a_8_24# 0.03fF
C23236 AND2X1_LOC_70/Y OR2X1_LOC_786/A 0.01fF
C23746 AND2X1_LOC_70/Y OR2X1_LOC_161/A 0.86fF
C23837 AND2X1_LOC_70/Y AND2X1_LOC_51/Y 12.67fF
C24350 AND2X1_LOC_70/Y AND2X1_LOC_52/Y 0.03fF
C24502 AND2X1_LOC_70/Y AND2X1_LOC_41/A 0.17fF
C24596 AND2X1_LOC_70/Y OR2X1_LOC_631/B 0.02fF
C24647 AND2X1_LOC_70/Y AND2X1_LOC_135/a_8_24# 0.03fF
C25224 AND2X1_LOC_70/Y OR2X1_LOC_112/A 0.08fF
C25704 AND2X1_LOC_70/Y OR2X1_LOC_355/a_8_216# 0.04fF
C25941 AND2X1_LOC_70/Y OR2X1_LOC_614/a_8_216# 0.01fF
C26013 AND2X1_LOC_70/Y AND2X1_LOC_31/Y 3.79fF
C26278 AND2X1_LOC_70/Y OR2X1_LOC_633/B 0.03fF
C26833 AND2X1_LOC_70/Y OR2X1_LOC_451/B 0.01fF
C26912 AND2X1_LOC_70/Y AND2X1_LOC_36/Y 2.05fF
C27081 AND2X1_LOC_586/a_8_24# AND2X1_LOC_70/Y 0.14fF
C27182 AND2X1_LOC_70/Y AND2X1_LOC_122/a_8_24# 0.01fF
C27563 AND2X1_LOC_70/Y OR2X1_LOC_636/B 0.01fF
C27809 AND2X1_LOC_70/Y OR2X1_LOC_856/A 0.06fF
C27838 AND2X1_LOC_70/Y AND2X1_LOC_313/a_8_24# 0.09fF
C28185 AND2X1_LOC_70/Y OR2X1_LOC_537/a_8_216# 0.06fF
C28332 AND2X1_LOC_70/Y OR2X1_LOC_330/Y 0.02fF
C28431 AND2X1_LOC_70/Y AND2X1_LOC_117/a_8_24# 0.01fF
C28783 AND2X1_LOC_584/a_8_24# AND2X1_LOC_70/Y 0.01fF
C29216 AND2X1_LOC_70/Y OR2X1_LOC_269/B 6.86fF
C29536 AND2X1_LOC_70/Y AND2X1_LOC_172/a_8_24# 0.10fF
C30277 AND2X1_LOC_70/Y OR2X1_LOC_777/B 0.06fF
C30700 OR2X1_LOC_198/a_8_216# AND2X1_LOC_70/Y 0.01fF
C30749 AND2X1_LOC_70/Y OR2X1_LOC_161/B 1.51fF
C30833 AND2X1_LOC_70/Y OR2X1_LOC_435/B 0.01fF
C30879 AND2X1_LOC_70/Y AND2X1_LOC_536/a_8_24# 0.01fF
C31254 AND2X1_LOC_70/Y OR2X1_LOC_630/B 0.01fF
C33274 AND2X1_LOC_70/Y AND2X1_LOC_7/B 0.15fF
C33379 OR2X1_LOC_318/Y AND2X1_LOC_70/Y 0.03fF
C33809 AND2X1_LOC_70/Y AND2X1_LOC_331/a_8_24# 0.06fF
C33924 AND2X1_LOC_70/Y OR2X1_LOC_123/B 0.01fF
C34355 AND2X1_LOC_70/Y OR2X1_LOC_446/Y 0.16fF
C34385 AND2X1_LOC_70/Y OR2X1_LOC_473/A 0.15fF
C34590 AND2X1_LOC_70/Y AND2X1_LOC_498/a_8_24# 0.01fF
C34651 AND2X1_LOC_70/Y OR2X1_LOC_635/a_8_216# 0.01fF
C35023 OR2X1_LOC_160/B AND2X1_LOC_70/Y 0.20fF
C35098 AND2X1_LOC_70/Y OR2X1_LOC_553/A 0.03fF
C35842 AND2X1_LOC_70/Y OR2X1_LOC_151/A 0.45fF
C36301 AND2X1_LOC_70/Y OR2X1_LOC_174/A 0.01fF
C37092 AND2X1_LOC_70/Y OR2X1_LOC_631/A 0.01fF
C38189 AND2X1_LOC_70/Y AND2X1_LOC_109/a_8_24# 0.01fF
C38292 AND2X1_LOC_70/Y OR2X1_LOC_308/Y 0.03fF
C38772 AND2X1_LOC_70/Y OR2X1_LOC_828/Y 0.13fF
C39341 AND2X1_LOC_70/Y AND2X1_LOC_601/a_8_24# 0.01fF
C39411 AND2X1_LOC_70/Y OR2X1_LOC_446/a_8_216# 0.01fF
C39645 AND2X1_LOC_70/Y OR2X1_LOC_390/A 0.03fF
C40521 AND2X1_LOC_70/Y OR2X1_LOC_841/A 0.01fF
C41197 AND2X1_LOC_70/Y OR2X1_LOC_241/B 0.07fF
C41313 OR2X1_LOC_188/Y AND2X1_LOC_70/Y 0.08fF
C41467 AND2X1_LOC_70/Y OR2X1_LOC_405/Y 0.01fF
C41555 AND2X1_LOC_70/Y OR2X1_LOC_193/A 0.02fF
C41730 AND2X1_LOC_70/Y OR2X1_LOC_339/A 0.21fF
C41751 OR2X1_LOC_208/A AND2X1_LOC_70/Y 0.01fF
C41783 AND2X1_LOC_70/Y AND2X1_LOC_438/a_8_24# 0.01fF
C41800 AND2X1_LOC_70/Y OR2X1_LOC_831/A 0.03fF
C41811 AND2X1_LOC_70/Y OR2X1_LOC_598/Y 0.12fF
C41816 AND2X1_LOC_70/Y AND2X1_LOC_131/a_8_24# 0.01fF
C41852 OR2X1_LOC_335/Y AND2X1_LOC_70/Y 0.10fF
C41903 AND2X1_LOC_70/Y OR2X1_LOC_537/A 0.06fF
C42835 AND2X1_LOC_70/Y OR2X1_LOC_810/A 0.08fF
C43120 OR2X1_LOC_715/B AND2X1_LOC_70/Y 0.06fF
C43123 AND2X1_LOC_70/Y AND2X1_LOC_626/a_8_24# 0.01fF
C43248 AND2X1_LOC_81/a_8_24# AND2X1_LOC_70/Y 0.01fF
C44094 AND2X1_LOC_70/Y OR2X1_LOC_687/Y 0.03fF
C44509 AND2X1_LOC_70/Y OR2X1_LOC_828/B 0.03fF
C44803 AND2X1_LOC_91/a_8_24# AND2X1_LOC_70/Y 0.02fF
C44862 AND2X1_LOC_70/Y OR2X1_LOC_78/A 1.29fF
C44941 AND2X1_LOC_70/Y OR2X1_LOC_602/A 0.01fF
C45017 AND2X1_LOC_70/Y OR2X1_LOC_605/A 0.07fF
C45747 AND2X1_LOC_70/Y OR2X1_LOC_501/B 0.01fF
C46020 AND2X1_LOC_70/Y OR2X1_LOC_318/B 0.03fF
C46142 OR2X1_LOC_121/Y AND2X1_LOC_70/Y 0.09fF
C46201 AND2X1_LOC_70/Y OR2X1_LOC_538/A 0.04fF
C46261 AND2X1_LOC_12/Y AND2X1_LOC_70/Y 0.35fF
C46333 AND2X1_LOC_70/Y AND2X1_LOC_496/a_8_24# 0.01fF
C46639 AND2X1_LOC_70/Y OR2X1_LOC_168/B 0.01fF
C46724 AND2X1_LOC_59/Y AND2X1_LOC_70/Y 0.31fF
C46772 AND2X1_LOC_70/Y AND2X1_LOC_495/a_8_24# 0.01fF
C47330 AND2X1_LOC_70/Y OR2X1_LOC_544/A 0.01fF
C47536 AND2X1_LOC_70/Y OR2X1_LOC_140/A 0.01fF
C47619 AND2X1_LOC_70/Y OR2X1_LOC_833/B 0.07fF
C48790 AND2X1_LOC_70/Y OR2X1_LOC_629/B 0.01fF
C49185 OR2X1_LOC_186/Y AND2X1_LOC_70/Y 0.42fF
C49489 AND2X1_LOC_70/Y OR2X1_LOC_112/B 0.04fF
C49808 AND2X1_LOC_70/Y OR2X1_LOC_574/A 0.04fF
C50038 AND2X1_LOC_70/Y OR2X1_LOC_855/A 0.01fF
C50436 AND2X1_LOC_70/Y OR2X1_LOC_539/B 0.02fF
C50516 AND2X1_LOC_70/Y OR2X1_LOC_78/B 5.18fF
C50594 AND2X1_LOC_70/Y OR2X1_LOC_375/A 0.17fF
C50666 AND2X1_LOC_70/Y OR2X1_LOC_605/B 0.09fF
C50903 AND2X1_LOC_70/Y OR2X1_LOC_549/A 0.16fF
C51374 AND2X1_LOC_70/Y OR2X1_LOC_499/B 0.01fF
C51748 AND2X1_LOC_70/Y AND2X1_LOC_65/A 0.25fF
C52435 AND2X1_LOC_70/Y OR2X1_LOC_330/a_8_216# 0.02fF
C52667 OR2X1_LOC_115/a_8_216# AND2X1_LOC_70/Y 0.01fF
C52966 OR2X1_LOC_335/A AND2X1_LOC_70/Y 0.03fF
C53062 AND2X1_LOC_583/a_8_24# AND2X1_LOC_70/Y 0.01fF
C53396 OR2X1_LOC_139/A AND2X1_LOC_70/Y 0.08fF
C54441 AND2X1_LOC_70/Y AND2X1_LOC_666/a_8_24# 0.03fF
C54520 AND2X1_LOC_70/Y OR2X1_LOC_247/a_8_216# 0.01fF
C54796 AND2X1_LOC_70/Y OR2X1_LOC_87/A 0.65fF
C55107 AND2X1_LOC_70/Y OR2X1_LOC_389/A 0.01fF
C55156 AND2X1_LOC_70/Y AND2X1_LOC_177/a_8_24# 0.07fF
C55959 OR2X1_LOC_97/A AND2X1_LOC_70/Y 0.05fF
C56797 AND2X1_LOC_70/Y VSS 0.37fF
C110 OR2X1_LOC_47/Y OR2X1_LOC_754/a_8_216# 0.01fF
C443 AND2X1_LOC_547/Y OR2X1_LOC_47/Y 0.02fF
C525 AND2X1_LOC_729/Y OR2X1_LOC_47/Y 0.13fF
C539 AND2X1_LOC_784/A OR2X1_LOC_47/Y 0.09fF
C582 OR2X1_LOC_47/Y AND2X1_LOC_639/A 0.08fF
C1007 OR2X1_LOC_47/Y OR2X1_LOC_52/B 0.22fF
C1014 AND2X1_LOC_489/Y OR2X1_LOC_47/Y 0.02fF
C1322 OR2X1_LOC_47/Y OR2X1_LOC_584/Y 0.01fF
C1400 OR2X1_LOC_47/Y OR2X1_LOC_394/Y 0.37fF
C1441 OR2X1_LOC_280/Y OR2X1_LOC_47/Y 0.02fF
C1477 OR2X1_LOC_22/Y OR2X1_LOC_47/Y 0.14fF
C1819 OR2X1_LOC_47/Y OR2X1_LOC_39/A 0.19fF
C2230 OR2X1_LOC_47/Y AND2X1_LOC_240/a_8_24# 0.04fF
C2657 OR2X1_LOC_51/Y OR2X1_LOC_47/Y 0.17fF
C2712 OR2X1_LOC_680/A OR2X1_LOC_47/Y 0.03fF
C3289 OR2X1_LOC_47/Y AND2X1_LOC_790/a_8_24# 0.02fF
C3478 OR2X1_LOC_47/Y AND2X1_LOC_436/Y 0.03fF
C3513 AND2X1_LOC_344/a_8_24# OR2X1_LOC_47/Y 0.02fF
C3568 OR2X1_LOC_47/Y OR2X1_LOC_588/Y 0.02fF
C3714 OR2X1_LOC_47/Y OR2X1_LOC_152/a_8_216# 0.05fF
C3993 OR2X1_LOC_47/Y OR2X1_LOC_609/A 0.03fF
C4570 OR2X1_LOC_47/Y OR2X1_LOC_183/Y 0.23fF
C4777 OR2X1_LOC_47/Y OR2X1_LOC_248/a_8_216# 0.08fF
C5169 OR2X1_LOC_47/Y OR2X1_LOC_237/Y 0.02fF
C5545 AND2X1_LOC_391/Y OR2X1_LOC_47/Y 0.03fF
C5549 OR2X1_LOC_91/A OR2X1_LOC_47/Y 0.83fF
C6026 OR2X1_LOC_32/B OR2X1_LOC_47/Y 0.10fF
C6053 OR2X1_LOC_47/Y OR2X1_LOC_371/Y 0.04fF
C6467 OR2X1_LOC_490/Y OR2X1_LOC_47/Y 0.05fF
C6468 OR2X1_LOC_47/Y OR2X1_LOC_74/A 0.12fF
C7822 OR2X1_LOC_615/a_8_216# OR2X1_LOC_47/Y 0.01fF
C8238 OR2X1_LOC_47/Y AND2X1_LOC_633/a_8_24# 0.16fF
C8996 OR2X1_LOC_47/Y AND2X1_LOC_614/a_8_24# 0.02fF
C9060 AND2X1_LOC_99/A OR2X1_LOC_47/Y 0.02fF
C9252 OR2X1_LOC_47/Y OR2X1_LOC_152/a_36_216# 0.03fF
C9584 OR2X1_LOC_167/Y OR2X1_LOC_47/Y 0.01fF
C9841 AND2X1_LOC_362/B OR2X1_LOC_47/Y 0.24fF
C10375 OR2X1_LOC_485/A OR2X1_LOC_47/Y 5.49fF
C10464 OR2X1_LOC_47/Y OR2X1_LOC_609/Y 0.06fF
C10633 AND2X1_LOC_802/B OR2X1_LOC_47/Y 0.03fF
C11154 OR2X1_LOC_695/a_8_216# OR2X1_LOC_47/Y 0.06fF
C12363 OR2X1_LOC_47/Y OR2X1_LOC_13/Y 0.02fF
C12850 OR2X1_LOC_441/a_8_216# OR2X1_LOC_47/Y 0.14fF
C13253 OR2X1_LOC_106/a_8_216# OR2X1_LOC_47/Y 0.07fF
C14004 OR2X1_LOC_516/Y OR2X1_LOC_47/Y 0.03fF
C14331 OR2X1_LOC_47/Y AND2X1_LOC_793/B 0.01fF
C14570 AND2X1_LOC_348/A OR2X1_LOC_47/Y 0.01fF
C14923 OR2X1_LOC_47/Y OR2X1_LOC_583/a_8_216# 0.01fF
C15334 VDD OR2X1_LOC_47/Y 2.54fF
C15477 OR2X1_LOC_256/A OR2X1_LOC_47/Y 0.04fF
C15519 OR2X1_LOC_47/Y OR2X1_LOC_67/Y 0.03fF
C15826 OR2X1_LOC_47/Y OR2X1_LOC_248/Y 0.70fF
C16123 OR2X1_LOC_47/Y AND2X1_LOC_457/a_8_24# 0.10fF
C16539 OR2X1_LOC_494/A OR2X1_LOC_47/Y 0.03fF
C16666 OR2X1_LOC_47/Y OR2X1_LOC_427/A 1.44fF
C17971 OR2X1_LOC_47/Y OR2X1_LOC_44/Y 9.11fF
C18279 OR2X1_LOC_45/B OR2X1_LOC_47/Y 5.07fF
C18759 OR2X1_LOC_158/A OR2X1_LOC_47/Y 0.14fF
C18769 OR2X1_LOC_106/a_36_216# OR2X1_LOC_47/Y 0.03fF
C18817 AND2X1_LOC_98/Y OR2X1_LOC_47/Y 0.02fF
C18824 OR2X1_LOC_103/Y OR2X1_LOC_47/Y 0.03fF
C18838 OR2X1_LOC_103/a_8_216# OR2X1_LOC_47/Y 0.01fF
C20587 OR2X1_LOC_47/Y OR2X1_LOC_438/a_8_216# 0.03fF
C20932 OR2X1_LOC_107/a_8_216# OR2X1_LOC_47/Y 0.01fF
C21010 AND2X1_LOC_390/B OR2X1_LOC_47/Y 0.07fF
C21380 OR2X1_LOC_744/A OR2X1_LOC_47/Y 0.29fF
C21436 OR2X1_LOC_47/Y AND2X1_LOC_840/B 0.05fF
C21520 OR2X1_LOC_47/Y OR2X1_LOC_31/Y 3.32fF
C21723 OR2X1_LOC_47/Y AND2X1_LOC_464/A 0.42fF
C21781 OR2X1_LOC_694/Y OR2X1_LOC_47/Y 0.13fF
C22664 OR2X1_LOC_47/Y OR2X1_LOC_56/A 0.22fF
C23068 OR2X1_LOC_47/Y AND2X1_LOC_285/Y 0.02fF
C23126 OR2X1_LOC_91/Y OR2X1_LOC_47/Y 0.15fF
C23153 OR2X1_LOC_189/Y OR2X1_LOC_47/Y 7.71fF
C23159 OR2X1_LOC_152/Y OR2X1_LOC_47/Y 0.24fF
C23177 OR2X1_LOC_291/Y OR2X1_LOC_47/Y 1.99fF
C23256 OR2X1_LOC_47/Y AND2X1_LOC_483/Y 0.17fF
C23518 OR2X1_LOC_494/a_8_216# OR2X1_LOC_47/Y 0.01fF
C23557 OR2X1_LOC_83/A OR2X1_LOC_47/Y 0.07fF
C23927 OR2X1_LOC_441/Y OR2X1_LOC_47/Y 0.06fF
C23961 OR2X1_LOC_47/Y AND2X1_LOC_436/B 0.02fF
C24419 OR2X1_LOC_481/A OR2X1_LOC_47/Y 0.01fF
C24446 OR2X1_LOC_47/Y OR2X1_LOC_71/Y 0.02fF
C24845 OR2X1_LOC_47/Y OR2X1_LOC_246/A 0.05fF
C24876 OR2X1_LOC_47/Y OR2X1_LOC_409/B 0.02fF
C25611 OR2X1_LOC_109/a_8_216# OR2X1_LOC_47/Y 0.01fF
C26037 AND2X1_LOC_319/A OR2X1_LOC_47/Y 0.16fF
C26151 OR2X1_LOC_47/Y AND2X1_LOC_721/A 0.05fF
C26183 OR2X1_LOC_47/Y OR2X1_LOC_331/Y 0.07fF
C26462 OR2X1_LOC_47/Y AND2X1_LOC_361/A 0.85fF
C26878 OR2X1_LOC_47/Y OR2X1_LOC_96/B 0.03fF
C26896 OR2X1_LOC_83/Y OR2X1_LOC_47/Y 0.01fF
C27192 AND2X1_LOC_787/A OR2X1_LOC_47/Y 0.03fF
C28046 OR2X1_LOC_692/Y OR2X1_LOC_47/Y 0.01fF
C28057 AND2X1_LOC_729/a_8_24# OR2X1_LOC_47/Y 0.01fF
C28089 OR2X1_LOC_600/A OR2X1_LOC_47/Y 0.22fF
C28101 OR2X1_LOC_166/a_8_216# OR2X1_LOC_47/Y 0.03fF
C28145 OR2X1_LOC_47/Y OR2X1_LOC_619/Y 0.22fF
C28592 OR2X1_LOC_232/a_8_216# OR2X1_LOC_47/Y 0.01fF
C28624 OR2X1_LOC_601/a_36_216# OR2X1_LOC_47/Y 0.01fF
C29113 OR2X1_LOC_47/Y OR2X1_LOC_406/A 0.01fF
C29320 OR2X1_LOC_329/Y OR2X1_LOC_47/Y 0.01fF
C29809 AND2X1_LOC_113/a_8_24# OR2X1_LOC_47/Y 0.02fF
C30235 OR2X1_LOC_47/Y OR2X1_LOC_393/a_8_216# 0.01fF
C30284 OR2X1_LOC_312/Y OR2X1_LOC_47/Y 0.04fF
C30450 OR2X1_LOC_47/Y OR2X1_LOC_13/B 1.41fF
C30988 OR2X1_LOC_47/Y OR2X1_LOC_428/A 0.74fF
C31007 OR2X1_LOC_47/Y OR2X1_LOC_595/A 0.03fF
C31439 OR2X1_LOC_47/Y OR2X1_LOC_583/Y 0.02fF
C31530 AND2X1_LOC_342/Y OR2X1_LOC_47/Y 0.04fF
C31557 OR2X1_LOC_47/Y OR2X1_LOC_438/a_36_216# 0.03fF
C31833 OR2X1_LOC_47/Y OR2X1_LOC_765/Y 0.03fF
C31933 OR2X1_LOC_26/Y OR2X1_LOC_47/Y 3.84fF
C31940 OR2X1_LOC_47/Y OR2X1_LOC_89/A 0.17fF
C32210 OR2X1_LOC_167/a_8_216# OR2X1_LOC_47/Y 0.01fF
C32790 OR2X1_LOC_47/Y OR2X1_LOC_824/Y 0.07fF
C32837 AND2X1_LOC_727/A OR2X1_LOC_47/Y 0.03fF
C32857 OR2X1_LOC_47/Y OR2X1_LOC_95/Y 0.86fF
C33084 OR2X1_LOC_821/Y OR2X1_LOC_47/Y 0.03fF
C33162 OR2X1_LOC_122/Y OR2X1_LOC_47/Y 0.02fF
C33601 OR2X1_LOC_166/a_36_216# OR2X1_LOC_47/Y 0.01fF
C33621 OR2X1_LOC_438/Y OR2X1_LOC_47/Y 0.43fF
C33651 OR2X1_LOC_47/Y AND2X1_LOC_621/Y 0.03fF
C33821 OR2X1_LOC_47/Y OR2X1_LOC_71/A 0.03fF
C34000 OR2X1_LOC_47/Y OR2X1_LOC_59/Y 0.34fF
C34091 OR2X1_LOC_70/Y OR2X1_LOC_47/Y 0.12fF
C34914 OR2X1_LOC_625/Y OR2X1_LOC_47/Y 0.11fF
C35193 OR2X1_LOC_47/Y OR2X1_LOC_584/a_8_216# 0.01fF
C35215 AND2X1_LOC_535/Y OR2X1_LOC_47/Y 0.03fF
C35293 OR2X1_LOC_246/Y OR2X1_LOC_47/Y 0.18fF
C35626 OR2X1_LOC_47/Y OR2X1_LOC_16/A 0.28fF
C35657 OR2X1_LOC_108/Y OR2X1_LOC_47/Y 0.02fF
C35721 AND2X1_LOC_168/Y OR2X1_LOC_47/Y 0.03fF
C35803 OR2X1_LOC_47/Y AND2X1_LOC_687/Y 0.02fF
C36501 OR2X1_LOC_47/Y AND2X1_LOC_447/Y 0.10fF
C36554 OR2X1_LOC_109/Y OR2X1_LOC_47/Y 0.08fF
C36596 OR2X1_LOC_47/Y AND2X1_LOC_729/B 0.02fF
C37065 AND2X1_LOC_227/Y OR2X1_LOC_47/Y 0.02fF
C37119 OR2X1_LOC_47/Y OR2X1_LOC_753/Y 0.04fF
C37359 OR2X1_LOC_107/Y OR2X1_LOC_47/Y 0.01fF
C37437 OR2X1_LOC_599/A OR2X1_LOC_47/Y 0.83fF
C37724 OR2X1_LOC_177/a_8_216# OR2X1_LOC_47/Y 0.01fF
C37750 OR2X1_LOC_40/Y OR2X1_LOC_47/Y 7.47fF
C37847 OR2X1_LOC_47/Y OR2X1_LOC_7/A 0.73fF
C38104 OR2X1_LOC_176/a_8_216# OR2X1_LOC_47/Y 0.01fF
C38177 OR2X1_LOC_822/a_8_216# OR2X1_LOC_47/Y 0.01fF
C38348 OR2X1_LOC_47/Y OR2X1_LOC_615/Y 0.22fF
C38686 AND2X1_LOC_841/B OR2X1_LOC_47/Y 0.03fF
C38989 AND2X1_LOC_543/Y OR2X1_LOC_47/Y 0.15fF
C39047 OR2X1_LOC_589/A OR2X1_LOC_47/Y 0.32fF
C39055 OR2X1_LOC_47/Y OR2X1_LOC_322/Y 0.15fF
C39084 OR2X1_LOC_166/Y OR2X1_LOC_47/Y 0.03fF
C39600 OR2X1_LOC_47/Y AND2X1_LOC_240/Y 0.01fF
C39984 OR2X1_LOC_3/Y OR2X1_LOC_47/Y 0.62fF
C40380 AND2X1_LOC_113/Y OR2X1_LOC_47/Y 0.01fF
C40823 OR2X1_LOC_47/Y AND2X1_LOC_610/a_8_24# 0.04fF
C40830 OR2X1_LOC_280/a_8_216# OR2X1_LOC_47/Y 0.08fF
C41136 OR2X1_LOC_47/Y OR2X1_LOC_766/a_8_216# 0.01fF
C41299 OR2X1_LOC_64/Y OR2X1_LOC_47/Y 1.11fF
C41477 OR2X1_LOC_47/Y AND2X1_LOC_247/a_8_24# 0.02fF
C41653 OR2X1_LOC_47/Y OR2X1_LOC_232/Y 0.03fF
C42016 OR2X1_LOC_47/Y OR2X1_LOC_524/a_8_216# 0.01fF
C42661 AND2X1_LOC_196/Y OR2X1_LOC_47/Y 0.08fF
C43808 OR2X1_LOC_494/Y OR2X1_LOC_47/Y 0.01fF
C44650 OR2X1_LOC_47/Y AND2X1_LOC_778/Y 0.03fF
C44720 OR2X1_LOC_47/Y AND2X1_LOC_624/A 0.03fF
C44731 OR2X1_LOC_380/A OR2X1_LOC_47/Y 0.02fF
C45561 OR2X1_LOC_524/Y OR2X1_LOC_47/Y 0.65fF
C45902 OR2X1_LOC_47/Y OR2X1_LOC_312/a_8_216# 0.01fF
C46527 OR2X1_LOC_47/Y OR2X1_LOC_612/B 0.03fF
C46934 OR2X1_LOC_47/Y OR2X1_LOC_278/Y 0.02fF
C47180 OR2X1_LOC_47/Y AND2X1_LOC_608/a_8_24# 0.04fF
C47458 OR2X1_LOC_754/A OR2X1_LOC_47/Y 0.06fF
C47649 OR2X1_LOC_47/Y OR2X1_LOC_142/Y 0.03fF
C48334 OR2X1_LOC_47/Y OR2X1_LOC_83/a_8_216# 0.01fF
C48443 OR2X1_LOC_47/Y OR2X1_LOC_754/Y 0.01fF
C48702 OR2X1_LOC_36/Y OR2X1_LOC_47/Y 0.22fF
C48810 OR2X1_LOC_47/Y OR2X1_LOC_419/Y 0.03fF
C48838 OR2X1_LOC_47/Y OR2X1_LOC_152/A 0.05fF
C49002 OR2X1_LOC_177/Y OR2X1_LOC_47/Y 0.06fF
C49024 OR2X1_LOC_604/A OR2X1_LOC_47/Y 0.39fF
C49100 OR2X1_LOC_80/Y OR2X1_LOC_47/Y 0.01fF
C49216 OR2X1_LOC_47/Y OR2X1_LOC_747/a_8_216# 0.18fF
C49408 OR2X1_LOC_176/Y OR2X1_LOC_47/Y 0.28fF
C49932 OR2X1_LOC_164/Y OR2X1_LOC_47/Y 0.06fF
C50033 AND2X1_LOC_633/Y OR2X1_LOC_47/Y 0.18fF
C50241 AND2X1_LOC_539/Y OR2X1_LOC_47/Y 0.03fF
C52052 AND2X1_LOC_342/a_8_24# OR2X1_LOC_47/Y 0.01fF
C52065 OR2X1_LOC_47/Y AND2X1_LOC_610/a_36_24# 0.01fF
C52070 OR2X1_LOC_280/a_36_216# OR2X1_LOC_47/Y 0.03fF
C52374 OR2X1_LOC_47/Y OR2X1_LOC_12/Y 0.20fF
C52378 OR2X1_LOC_47/Y OR2X1_LOC_766/Y 0.01fF
C52472 OR2X1_LOC_47/Y OR2X1_LOC_393/Y 0.34fF
C52695 OR2X1_LOC_47/Y OR2X1_LOC_248/A 0.09fF
C52869 OR2X1_LOC_47/Y OR2X1_LOC_234/Y 0.01fF
C52969 OR2X1_LOC_278/A OR2X1_LOC_47/Y 0.29fF
C53319 OR2X1_LOC_47/Y AND2X1_LOC_848/Y 0.03fF
C54091 OR2X1_LOC_178/Y OR2X1_LOC_47/Y 0.02fF
C54115 OR2X1_LOC_256/Y OR2X1_LOC_47/Y 0.06fF
C54884 AND2X1_LOC_361/a_8_24# OR2X1_LOC_47/Y 0.03fF
C54923 OR2X1_LOC_822/Y OR2X1_LOC_47/Y 0.01fF
C54984 OR2X1_LOC_18/Y OR2X1_LOC_47/Y 0.23fF
C55340 OR2X1_LOC_47/Y AND2X1_LOC_810/B 0.07fF
C56061 OR2X1_LOC_47/Y OR2X1_LOC_437/A 0.41fF
C57101 OR2X1_LOC_47/Y VSS 1.86fF
C482 OR2X1_LOC_416/Y OR2X1_LOC_44/Y 0.03fF
C595 OR2X1_LOC_44/Y AND2X1_LOC_592/a_8_24# 0.02fF
C1269 OR2X1_LOC_485/a_8_216# OR2X1_LOC_44/Y 0.07fF
C1296 OR2X1_LOC_45/a_8_216# OR2X1_LOC_44/Y 0.05fF
C1298 OR2X1_LOC_701/Y OR2X1_LOC_44/Y 0.10fF
C1565 OR2X1_LOC_45/B OR2X1_LOC_44/Y 0.19fF
C1726 AND2X1_LOC_435/a_8_24# OR2X1_LOC_44/Y 0.01fF
C1765 OR2X1_LOC_261/Y OR2X1_LOC_44/Y 0.26fF
C2025 OR2X1_LOC_158/A OR2X1_LOC_44/Y 1.17fF
C2101 OR2X1_LOC_103/Y OR2X1_LOC_44/Y 0.03fF
C2484 OR2X1_LOC_482/Y OR2X1_LOC_44/Y 0.03fF
C2576 OR2X1_LOC_44/Y OR2X1_LOC_586/Y 0.03fF
C2635 OR2X1_LOC_748/A OR2X1_LOC_44/Y 0.04fF
C3028 AND2X1_LOC_848/a_8_24# OR2X1_LOC_44/Y 0.01fF
C3340 OR2X1_LOC_368/a_36_216# OR2X1_LOC_44/Y 0.02fF
C3432 AND2X1_LOC_97/a_36_24# OR2X1_LOC_44/Y 0.01fF
C3590 AND2X1_LOC_848/A OR2X1_LOC_44/Y 0.09fF
C3730 OR2X1_LOC_591/Y OR2X1_LOC_44/Y 0.04fF
C4166 OR2X1_LOC_107/a_8_216# OR2X1_LOC_44/Y 0.02fF
C4230 OR2X1_LOC_316/Y OR2X1_LOC_44/Y 0.11fF
C4287 AND2X1_LOC_390/B OR2X1_LOC_44/Y 0.07fF
C4580 OR2X1_LOC_744/A OR2X1_LOC_44/Y 0.89fF
C4752 OR2X1_LOC_31/Y OR2X1_LOC_44/Y 2.63fF
C4908 AND2X1_LOC_464/A OR2X1_LOC_44/Y 0.05fF
C5419 OR2X1_LOC_179/a_8_216# OR2X1_LOC_44/Y 0.02fF
C5594 OR2X1_LOC_751/A OR2X1_LOC_44/Y 0.28fF
C5845 OR2X1_LOC_56/A OR2X1_LOC_44/Y 0.26fF
C5888 AND2X1_LOC_638/Y OR2X1_LOC_44/Y 0.04fF
C6326 OR2X1_LOC_91/Y OR2X1_LOC_44/Y 11.98fF
C6374 OR2X1_LOC_44/Y OR2X1_LOC_757/Y 0.37fF
C6406 OR2X1_LOC_417/Y OR2X1_LOC_44/Y 0.07fF
C6423 OR2X1_LOC_601/a_8_216# OR2X1_LOC_44/Y 0.05fF
C6806 OR2X1_LOC_44/Y OR2X1_LOC_701/a_8_216# 0.01fF
C7725 OR2X1_LOC_481/A OR2X1_LOC_44/Y 0.03fF
C7760 OR2X1_LOC_71/Y OR2X1_LOC_44/Y 0.03fF
C7875 OR2X1_LOC_44/Y AND2X1_LOC_789/Y 0.09fF
C8236 OR2X1_LOC_409/B OR2X1_LOC_44/Y 0.03fF
C8621 OR2X1_LOC_229/Y OR2X1_LOC_44/Y 0.02fF
C8882 OR2X1_LOC_380/a_8_216# OR2X1_LOC_44/Y 0.01fF
C8947 AND2X1_LOC_344/a_36_24# OR2X1_LOC_44/Y 0.01fF
C8995 OR2X1_LOC_24/a_8_216# OR2X1_LOC_44/Y 0.06fF
C9427 AND2X1_LOC_319/A OR2X1_LOC_44/Y 0.07fF
C9474 OR2X1_LOC_52/a_8_216# OR2X1_LOC_44/Y 0.01fF
C9542 AND2X1_LOC_721/A OR2X1_LOC_44/Y 0.03fF
C9560 OR2X1_LOC_44/Y OR2X1_LOC_331/Y 0.07fF
C9758 OR2X1_LOC_107/a_36_216# OR2X1_LOC_44/Y 0.02fF
C10253 OR2X1_LOC_96/B OR2X1_LOC_44/Y 0.04fF
C10273 OR2X1_LOC_83/Y OR2X1_LOC_44/Y 0.02fF
C10487 AND2X1_LOC_284/a_8_24# OR2X1_LOC_44/Y 0.01fF
C10496 AND2X1_LOC_787/A OR2X1_LOC_44/Y 0.03fF
C11006 OR2X1_LOC_179/a_36_216# OR2X1_LOC_44/Y 0.02fF
C11348 OR2X1_LOC_692/Y OR2X1_LOC_44/Y 0.14fF
C11387 OR2X1_LOC_600/A OR2X1_LOC_44/Y 2.13fF
C11403 OR2X1_LOC_166/a_8_216# OR2X1_LOC_44/Y 0.05fF
C11491 OR2X1_LOC_619/Y OR2X1_LOC_44/Y 0.14fF
C11776 OR2X1_LOC_44/Y AND2X1_LOC_769/Y 0.03fF
C12159 OR2X1_LOC_44/Y AND2X1_LOC_783/B 0.04fF
C12786 OR2X1_LOC_69/A OR2X1_LOC_44/Y 0.02fF
C13223 AND2X1_LOC_779/a_36_24# OR2X1_LOC_44/Y 0.02fF
C13683 OR2X1_LOC_312/Y OR2X1_LOC_44/Y 0.03fF
C13838 OR2X1_LOC_44/Y OR2X1_LOC_13/B 0.15fF
C13947 AND2X1_LOC_199/A OR2X1_LOC_44/Y 0.10fF
C14337 OR2X1_LOC_44/Y OR2X1_LOC_428/A 0.23fF
C14347 OR2X1_LOC_44/Y OR2X1_LOC_595/A 0.03fF
C14778 AND2X1_LOC_592/Y OR2X1_LOC_44/Y 0.05fF
C14958 OR2X1_LOC_279/a_8_216# OR2X1_LOC_44/Y 0.03fF
C15326 OR2X1_LOC_26/Y OR2X1_LOC_44/Y 0.60fF
C15338 OR2X1_LOC_89/A OR2X1_LOC_44/Y 0.47fF
C16118 OR2X1_LOC_45/Y OR2X1_LOC_44/Y 0.08fF
C16176 OR2X1_LOC_591/a_8_216# OR2X1_LOC_44/Y 0.02fF
C16230 AND2X1_LOC_727/A OR2X1_LOC_44/Y 0.03fF
C16259 OR2X1_LOC_95/Y OR2X1_LOC_44/Y 2.17fF
C16515 OR2X1_LOC_297/a_8_216# OR2X1_LOC_44/Y 0.03fF
C16541 AND2X1_LOC_832/a_8_24# OR2X1_LOC_44/Y 0.02fF
C16878 OR2X1_LOC_693/Y OR2X1_LOC_44/Y 0.01fF
C17011 AND2X1_LOC_621/Y OR2X1_LOC_44/Y 0.03fF
C17348 OR2X1_LOC_59/Y OR2X1_LOC_44/Y 2.89fF
C17476 OR2X1_LOC_70/Y OR2X1_LOC_44/Y 0.13fF
C17537 OR2X1_LOC_184/Y OR2X1_LOC_44/Y 0.03fF
C18281 OR2X1_LOC_625/Y OR2X1_LOC_44/Y 0.07fF
C18528 OR2X1_LOC_44/Y OR2X1_LOC_759/Y 0.22fF
C18621 AND2X1_LOC_535/Y OR2X1_LOC_44/Y 0.03fF
C19003 OR2X1_LOC_16/A OR2X1_LOC_44/Y 0.06fF
C19046 OR2X1_LOC_108/Y OR2X1_LOC_44/Y 0.07fF
C19239 AND2X1_LOC_687/Y OR2X1_LOC_44/Y 0.02fF
C19872 OR2X1_LOC_44/Y OR2X1_LOC_759/a_8_216# 0.01fF
C19930 AND2X1_LOC_447/Y OR2X1_LOC_44/Y 0.71fF
C19946 OR2X1_LOC_380/Y OR2X1_LOC_44/Y 0.30fF
C20005 OR2X1_LOC_109/Y OR2X1_LOC_44/Y 0.08fF
C20078 AND2X1_LOC_729/B OR2X1_LOC_44/Y 0.03fF
C20312 AND2X1_LOC_593/a_8_24# OR2X1_LOC_44/Y 0.02fF
C20493 OR2X1_LOC_279/a_36_216# OR2X1_LOC_44/Y 0.03fF
C20560 AND2X1_LOC_227/Y OR2X1_LOC_44/Y 0.06fF
C20896 OR2X1_LOC_599/A OR2X1_LOC_44/Y 0.09fF
C21195 OR2X1_LOC_40/Y OR2X1_LOC_44/Y 0.10fF
C21306 OR2X1_LOC_424/a_8_216# OR2X1_LOC_44/Y 0.05fF
C21358 OR2X1_LOC_7/A OR2X1_LOC_44/Y 9.23fF
C21933 OR2X1_LOC_44/Y OR2X1_LOC_424/Y 0.02fF
C22154 AND2X1_LOC_841/B OR2X1_LOC_44/Y 0.01fF
C22412 AND2X1_LOC_543/Y OR2X1_LOC_44/Y 0.04fF
C22465 AND2X1_LOC_706/a_8_24# OR2X1_LOC_44/Y 0.01fF
C22475 OR2X1_LOC_589/A OR2X1_LOC_44/Y 0.01fF
C22479 OR2X1_LOC_44/Y OR2X1_LOC_322/Y 0.08fF
C22513 OR2X1_LOC_261/a_8_216# OR2X1_LOC_44/Y 0.01fF
C22528 OR2X1_LOC_166/Y OR2X1_LOC_44/Y 0.03fF
C22618 AND2X1_LOC_379/a_8_24# OR2X1_LOC_44/Y 0.01fF
C23488 OR2X1_LOC_3/Y OR2X1_LOC_44/Y 2.83fF
C23562 AND2X1_LOC_462/B OR2X1_LOC_44/Y 0.80fF
C24602 OR2X1_LOC_122/A OR2X1_LOC_44/Y 0.01fF
C24720 OR2X1_LOC_690/A OR2X1_LOC_44/Y 0.08fF
C24761 OR2X1_LOC_64/Y OR2X1_LOC_44/Y 2.70fF
C25601 OR2X1_LOC_7/Y OR2X1_LOC_44/Y 0.43fF
C25969 OR2X1_LOC_279/Y OR2X1_LOC_44/Y 0.31fF
C26621 AND2X1_LOC_828/a_8_24# OR2X1_LOC_44/Y 0.01fF
C26769 OR2X1_LOC_424/a_36_216# OR2X1_LOC_44/Y 0.01fF
C27121 OR2X1_LOC_494/Y OR2X1_LOC_44/Y 0.06fF
C27726 OR2X1_LOC_751/a_8_216# OR2X1_LOC_44/Y 0.01fF
C28049 AND2X1_LOC_624/A OR2X1_LOC_44/Y 0.03fF
C28059 OR2X1_LOC_380/A OR2X1_LOC_44/Y 0.03fF
C28401 OR2X1_LOC_755/a_8_216# OR2X1_LOC_44/Y 0.01fF
C28909 OR2X1_LOC_763/Y OR2X1_LOC_44/Y 0.04fF
C28925 OR2X1_LOC_481/a_8_216# OR2X1_LOC_44/Y 0.01fF
C29456 OR2X1_LOC_44/Y AND2X1_LOC_779/Y 0.01fF
C30132 OR2X1_LOC_278/Y OR2X1_LOC_44/Y 0.03fF
C30396 OR2X1_LOC_89/Y OR2X1_LOC_44/Y 0.21fF
C30419 OR2X1_LOC_744/a_8_216# OR2X1_LOC_44/Y 0.02fF
C30510 OR2X1_LOC_751/Y OR2X1_LOC_44/Y 0.01fF
C31472 OR2X1_LOC_52/Y OR2X1_LOC_44/Y 0.02fF
C31528 OR2X1_LOC_503/Y OR2X1_LOC_44/Y 0.01fF
C31664 OR2X1_LOC_44/Y OR2X1_LOC_748/Y 0.02fF
C31829 OR2X1_LOC_36/Y OR2X1_LOC_44/Y 1.12fF
C31830 OR2X1_LOC_91/a_8_216# OR2X1_LOC_44/Y 0.02fF
C32087 OR2X1_LOC_315/a_8_216# OR2X1_LOC_44/Y 0.01fF
C32119 OR2X1_LOC_604/A OR2X1_LOC_44/Y 0.21fF
C32493 OR2X1_LOC_176/Y OR2X1_LOC_44/Y 0.03fF
C33339 AND2X1_LOC_539/Y OR2X1_LOC_44/Y 0.03fF
C33429 AND2X1_LOC_711/A OR2X1_LOC_44/Y 0.15fF
C33764 OR2X1_LOC_316/a_8_216# OR2X1_LOC_44/Y 0.04fF
C34258 OR2X1_LOC_700/a_8_216# OR2X1_LOC_44/Y 0.01fF
C34381 OR2X1_LOC_764/Y OR2X1_LOC_44/Y 0.01fF
C34871 AND2X1_LOC_197/a_8_24# OR2X1_LOC_44/Y 0.01fF
C35475 OR2X1_LOC_12/Y OR2X1_LOC_44/Y 2.86fF
C35894 OR2X1_LOC_744/a_36_216# OR2X1_LOC_44/Y 0.03fF
C36006 AND2X1_LOC_789/a_8_24# OR2X1_LOC_44/Y 0.01fF
C36460 AND2X1_LOC_848/Y OR2X1_LOC_44/Y 0.04fF
C37193 OR2X1_LOC_597/A OR2X1_LOC_44/Y 0.01fF
C37217 OR2X1_LOC_178/Y OR2X1_LOC_44/Y 0.03fF
C37252 OR2X1_LOC_256/Y OR2X1_LOC_44/Y 0.07fF
C37321 OR2X1_LOC_91/a_36_216# OR2X1_LOC_44/Y 0.02fF
C37586 OR2X1_LOC_829/A OR2X1_LOC_44/Y 0.15fF
C37588 OR2X1_LOC_315/a_36_216# OR2X1_LOC_44/Y 0.01fF
C38071 OR2X1_LOC_57/Y OR2X1_LOC_44/Y 0.02fF
C38077 AND2X1_LOC_508/A OR2X1_LOC_44/Y 0.03fF
C38119 OR2X1_LOC_18/Y OR2X1_LOC_44/Y 10.92fF
C38404 OR2X1_LOC_764/a_8_216# OR2X1_LOC_44/Y 0.01fF
C38867 OR2X1_LOC_368/Y OR2X1_LOC_44/Y 0.04fF
C38884 OR2X1_LOC_229/a_8_216# OR2X1_LOC_44/Y -0.00fF
C39214 OR2X1_LOC_44/Y OR2X1_LOC_437/A 0.35fF
C39398 OR2X1_LOC_755/Y OR2X1_LOC_44/Y 0.02fF
C39873 AND2X1_LOC_729/Y OR2X1_LOC_44/Y 0.07fF
C39895 AND2X1_LOC_784/A OR2X1_LOC_44/Y 0.07fF
C39907 AND2X1_LOC_769/a_8_24# OR2X1_LOC_44/Y 0.01fF
C39912 OR2X1_LOC_481/Y OR2X1_LOC_44/Y 0.31fF
C40004 OR2X1_LOC_44/Y OR2X1_LOC_172/Y 0.33fF
C40292 OR2X1_LOC_44/Y OR2X1_LOC_52/B 0.80fF
C40303 AND2X1_LOC_489/Y OR2X1_LOC_44/Y 0.03fF
C40686 OR2X1_LOC_394/Y OR2X1_LOC_44/Y 0.06fF
C40771 OR2X1_LOC_22/Y OR2X1_LOC_44/Y 0.83fF
C41141 OR2X1_LOC_44/Y OR2X1_LOC_39/A 0.22fF
C41928 OR2X1_LOC_51/Y OR2X1_LOC_44/Y 0.22fF
C42044 OR2X1_LOC_667/a_8_216# OR2X1_LOC_44/Y 0.05fF
C42663 OR2X1_LOC_44/Y OR2X1_LOC_399/a_8_216# 0.06fF
C42815 AND2X1_LOC_436/Y OR2X1_LOC_44/Y 0.03fF
C42857 AND2X1_LOC_344/a_8_24# OR2X1_LOC_44/Y 0.03fF
C42870 AND2X1_LOC_97/a_8_24# OR2X1_LOC_44/Y 0.04fF
C42915 OR2X1_LOC_588/Y OR2X1_LOC_44/Y 0.07fF
C43341 OR2X1_LOC_81/a_8_216# OR2X1_LOC_44/Y 0.14fF
C43718 AND2X1_LOC_197/Y OR2X1_LOC_44/Y 0.01fF
C44195 OR2X1_LOC_511/Y OR2X1_LOC_44/Y 0.13fF
C44246 OR2X1_LOC_297/Y OR2X1_LOC_44/Y 0.02fF
C44800 OR2X1_LOC_44/Y OR2X1_LOC_384/Y 0.03fF
C44989 OR2X1_LOC_91/A OR2X1_LOC_44/Y 1.34fF
C45131 OR2X1_LOC_44/Y OR2X1_LOC_27/Y 0.05fF
C45490 OR2X1_LOC_32/B OR2X1_LOC_44/Y 0.21fF
C45672 OR2X1_LOC_44/Y OR2X1_LOC_423/Y 0.03fF
C45972 OR2X1_LOC_44/Y OR2X1_LOC_757/a_8_216# 0.01fF
C45986 OR2X1_LOC_74/A OR2X1_LOC_44/Y 0.07fF
C46365 OR2X1_LOC_432/a_8_216# OR2X1_LOC_44/Y 0.01fF
C46833 OR2X1_LOC_432/Y OR2X1_LOC_44/Y 0.37fF
C47284 AND2X1_LOC_779/a_8_24# OR2X1_LOC_44/Y 0.02fF
C48176 AND2X1_LOC_847/Y OR2X1_LOC_44/Y 0.06fF
C48574 AND2X1_LOC_99/A OR2X1_LOC_44/Y 0.01fF
C48605 AND2X1_LOC_637/Y OR2X1_LOC_44/Y 0.02fF
C48949 OR2X1_LOC_697/Y OR2X1_LOC_44/Y 0.03fF
C49053 OR2X1_LOC_696/Y OR2X1_LOC_44/Y 0.03fF
C49229 OR2X1_LOC_44/Y OR2X1_LOC_503/a_8_216# 0.01fF
C49308 AND2X1_LOC_362/B OR2X1_LOC_44/Y 0.85fF
C49384 AND2X1_LOC_198/a_8_24# OR2X1_LOC_44/Y 0.01fF
C49722 AND2X1_LOC_706/Y OR2X1_LOC_44/Y 0.03fF
C49768 OR2X1_LOC_58/Y OR2X1_LOC_44/Y 0.03fF
C49888 OR2X1_LOC_81/Y OR2X1_LOC_44/Y 0.06fF
C49910 OR2X1_LOC_485/A OR2X1_LOC_44/Y 0.37fF
C50110 AND2X1_LOC_802/B OR2X1_LOC_44/Y 0.03fF
C50751 OR2X1_LOC_89/a_8_216# OR2X1_LOC_44/Y 0.01fF
C51275 OR2X1_LOC_44/Y OR2X1_LOC_589/Y 0.03fF
C51837 OR2X1_LOC_13/Y OR2X1_LOC_44/Y 0.03fF
C51933 OR2X1_LOC_700/Y OR2X1_LOC_44/Y 0.29fF
C52364 OR2X1_LOC_433/Y OR2X1_LOC_44/Y 0.03fF
C52665 AND2X1_LOC_714/B OR2X1_LOC_44/Y 0.12fF
C53406 OR2X1_LOC_44/Y OR2X1_LOC_589/a_8_216# 0.02fF
C53941 OR2X1_LOC_368/a_8_216# OR2X1_LOC_44/Y 0.02fF
C54788 VDD OR2X1_LOC_44/Y 1.19fF
C54833 AND2X1_LOC_208/B OR2X1_LOC_44/Y 0.01fF
C54870 OR2X1_LOC_315/Y OR2X1_LOC_44/Y 0.11fF
C54917 OR2X1_LOC_251/Y OR2X1_LOC_44/Y 0.15fF
C55593 AND2X1_LOC_457/a_8_24# OR2X1_LOC_44/Y 0.01fF
C55792 OR2X1_LOC_591/A OR2X1_LOC_44/Y 0.01fF
C56018 OR2X1_LOC_494/A OR2X1_LOC_44/Y 0.03fF
C56198 OR2X1_LOC_427/A OR2X1_LOC_44/Y 1.12fF
C56570 OR2X1_LOC_44/Y VSS 0.95fF
C689 OR2X1_LOC_31/Y OR2X1_LOC_589/a_8_216# 0.01fF
C874 OR2X1_LOC_369/Y OR2X1_LOC_31/Y -0.00fF
C1308 OR2X1_LOC_368/a_8_216# OR2X1_LOC_31/Y 0.09fF
C1730 OR2X1_LOC_31/Y OR2X1_LOC_583/a_8_216# 0.01fF
C2172 VDD OR2X1_LOC_31/Y 1.18fF
C2247 OR2X1_LOC_315/Y OR2X1_LOC_31/Y 0.14fF
C2626 OR2X1_LOC_60/Y OR2X1_LOC_31/Y 0.01fF
C2966 OR2X1_LOC_31/Y OR2X1_LOC_56/Y 0.24fF
C2989 OR2X1_LOC_31/Y AND2X1_LOC_457/a_8_24# 0.01fF
C3506 OR2X1_LOC_31/Y OR2X1_LOC_427/A 1.92fF
C4005 OR2X1_LOC_31/Y OR2X1_LOC_416/Y 0.03fF
C4103 OR2X1_LOC_31/Y AND2X1_LOC_592/a_8_24# 0.01fF
C4716 OR2X1_LOC_485/a_8_216# OR2X1_LOC_31/Y 0.01fF
C5012 OR2X1_LOC_45/B OR2X1_LOC_31/Y 0.59fF
C5144 OR2X1_LOC_31/Y AND2X1_LOC_435/a_8_24# 0.01fF
C5465 OR2X1_LOC_158/A OR2X1_LOC_31/Y 4.59fF
C6963 OR2X1_LOC_111/Y OR2X1_LOC_31/Y 0.48fF
C7207 OR2X1_LOC_591/Y OR2X1_LOC_31/Y 0.29fF
C7753 OR2X1_LOC_316/Y OR2X1_LOC_31/Y 0.07fF
C8141 OR2X1_LOC_744/A OR2X1_LOC_31/Y 0.11fF
C8229 OR2X1_LOC_31/Y AND2X1_LOC_840/B 0.20fF
C8237 OR2X1_LOC_31/Y OR2X1_LOC_74/a_8_216# 0.02fF
C8541 OR2X1_LOC_31/Y AND2X1_LOC_464/A 0.01fF
C8588 OR2X1_LOC_694/Y OR2X1_LOC_31/Y 0.09fF
C9442 OR2X1_LOC_31/Y OR2X1_LOC_56/A 0.09fF
C9926 OR2X1_LOC_91/Y OR2X1_LOC_31/Y 0.03fF
C9957 OR2X1_LOC_527/Y OR2X1_LOC_31/Y 0.09fF
C9965 OR2X1_LOC_417/Y OR2X1_LOC_31/Y 0.03fF
C9966 OR2X1_LOC_291/Y OR2X1_LOC_31/Y 0.06fF
C10169 OR2X1_LOC_31/Y OR2X1_LOC_171/Y 0.17fF
C10417 AND2X1_LOC_831/Y OR2X1_LOC_31/Y 0.15fF
C10755 OR2X1_LOC_31/Y AND2X1_LOC_436/B 0.01fF
C10758 AND2X1_LOC_139/B OR2X1_LOC_31/Y 0.13fF
C11651 OR2X1_LOC_246/A OR2X1_LOC_31/Y 0.01fF
C11675 OR2X1_LOC_31/Y OR2X1_LOC_409/B 0.03fF
C11952 OR2X1_LOC_298/a_8_216# OR2X1_LOC_31/Y 0.01fF
C12040 OR2X1_LOC_31/Y OR2X1_LOC_229/Y 0.01fF
C12434 OR2X1_LOC_109/a_8_216# OR2X1_LOC_31/Y 0.09fF
C12893 AND2X1_LOC_319/A OR2X1_LOC_31/Y 0.03fF
C12927 OR2X1_LOC_31/Y OR2X1_LOC_52/a_8_216# 0.01fF
C13749 OR2X1_LOC_31/Y OR2X1_LOC_74/a_36_216# 0.02fF
C14101 OR2X1_LOC_695/Y OR2X1_LOC_31/Y 0.01fF
C14437 AND2X1_LOC_520/a_8_24# OR2X1_LOC_31/Y 0.01fF
C14916 OR2X1_LOC_600/A OR2X1_LOC_31/Y 0.50fF
C14952 AND2X1_LOC_543/a_8_24# OR2X1_LOC_31/Y 0.01fF
C14989 OR2X1_LOC_31/Y OR2X1_LOC_619/Y 0.10fF
C15491 OR2X1_LOC_289/Y OR2X1_LOC_31/Y 0.03fF
C17292 OR2X1_LOC_31/Y OR2X1_LOC_13/B 0.20fF
C17787 OR2X1_LOC_31/Y OR2X1_LOC_428/A 0.66fF
C17800 OR2X1_LOC_31/Y OR2X1_LOC_595/A 0.03fF
C18286 AND2X1_LOC_592/Y OR2X1_LOC_31/Y 0.01fF
C18309 OR2X1_LOC_31/Y OR2X1_LOC_583/Y 0.02fF
C18850 OR2X1_LOC_26/Y OR2X1_LOC_31/Y 8.00fF
C18865 OR2X1_LOC_31/Y OR2X1_LOC_89/A 0.17fF
C19576 OR2X1_LOC_491/a_8_216# OR2X1_LOC_31/Y 0.08fF
C19609 AND2X1_LOC_707/a_8_24# OR2X1_LOC_31/Y 0.01fF
C19704 OR2X1_LOC_31/Y OR2X1_LOC_591/a_8_216# 0.01fF
C19764 OR2X1_LOC_31/Y OR2X1_LOC_95/Y 0.15fF
C20085 AND2X1_LOC_832/a_8_24# OR2X1_LOC_31/Y 0.01fF
C20912 OR2X1_LOC_31/Y OR2X1_LOC_59/Y 2.28fF
C21000 OR2X1_LOC_70/Y OR2X1_LOC_31/Y 0.28fF
C22155 OR2X1_LOC_31/Y OR2X1_LOC_584/a_8_216# 0.01fF
C22579 OR2X1_LOC_31/Y OR2X1_LOC_16/A 0.13fF
C22616 OR2X1_LOC_108/Y OR2X1_LOC_31/Y 0.14fF
C22790 AND2X1_LOC_687/Y OR2X1_LOC_31/Y 0.01fF
C23458 OR2X1_LOC_31/Y AND2X1_LOC_447/Y 0.04fF
C23466 OR2X1_LOC_31/Y OR2X1_LOC_380/Y 0.03fF
C23525 OR2X1_LOC_109/Y OR2X1_LOC_31/Y 0.02fF
C23855 AND2X1_LOC_593/a_8_24# OR2X1_LOC_31/Y 0.01fF
C24360 OR2X1_LOC_599/A OR2X1_LOC_31/Y 0.06fF
C24687 OR2X1_LOC_40/Y OR2X1_LOC_31/Y 1.37fF
C24773 OR2X1_LOC_424/a_8_216# OR2X1_LOC_31/Y 0.01fF
C24802 OR2X1_LOC_31/Y OR2X1_LOC_7/A 0.99fF
C24857 OR2X1_LOC_31/Y OR2X1_LOC_224/a_8_216# 0.02fF
C25374 OR2X1_LOC_31/Y OR2X1_LOC_424/Y 0.01fF
C25458 AND2X1_LOC_707/Y OR2X1_LOC_31/Y 0.05fF
C25580 AND2X1_LOC_841/B OR2X1_LOC_31/Y 0.01fF
C25843 AND2X1_LOC_543/Y OR2X1_LOC_31/Y 0.01fF
C25901 OR2X1_LOC_589/A OR2X1_LOC_31/Y 0.02fF
C25905 OR2X1_LOC_31/Y OR2X1_LOC_322/Y 0.04fF
C25981 OR2X1_LOC_495/Y OR2X1_LOC_31/Y 0.03fF
C26063 OR2X1_LOC_60/a_8_216# OR2X1_LOC_31/Y 0.01fF
C26887 OR2X1_LOC_3/Y OR2X1_LOC_31/Y 0.18fF
C27275 OR2X1_LOC_74/Y OR2X1_LOC_31/Y 0.02fF
C28019 OR2X1_LOC_31/Y OR2X1_LOC_766/a_8_216# 0.01fF
C28161 OR2X1_LOC_31/Y OR2X1_LOC_690/A 0.13fF
C28199 OR2X1_LOC_64/Y OR2X1_LOC_31/Y 1.39fF
C29025 OR2X1_LOC_31/Y OR2X1_LOC_7/Y 0.23fF
C31420 AND2X1_LOC_325/a_8_24# OR2X1_LOC_31/Y 0.02fF
C33686 OR2X1_LOC_273/Y OR2X1_LOC_31/Y 0.31fF
C34460 OR2X1_LOC_31/Y OR2X1_LOC_238/Y 0.02fF
C34949 OR2X1_LOC_31/Y OR2X1_LOC_52/Y 0.01fF
C35276 OR2X1_LOC_36/Y OR2X1_LOC_31/Y 4.18fF
C35381 OR2X1_LOC_31/Y OR2X1_LOC_419/Y 0.56fF
C35613 OR2X1_LOC_315/a_8_216# OR2X1_LOC_31/Y 0.07fF
C35632 OR2X1_LOC_604/A OR2X1_LOC_31/Y 0.08fF
C36139 OR2X1_LOC_31/Y OR2X1_LOC_265/Y 0.10fF
C36349 OR2X1_LOC_31/Y OR2X1_LOC_183/a_8_216# 0.01fF
C36510 OR2X1_LOC_164/Y OR2X1_LOC_31/Y 0.04fF
C36582 OR2X1_LOC_230/a_8_216# OR2X1_LOC_31/Y 0.19fF
C36597 AND2X1_LOC_633/Y OR2X1_LOC_31/Y 0.02fF
C36875 AND2X1_LOC_326/B OR2X1_LOC_31/Y 0.01fF
C37209 OR2X1_LOC_518/a_8_216# OR2X1_LOC_31/Y 0.01fF
C37216 OR2X1_LOC_316/a_8_216# OR2X1_LOC_31/Y 0.01fF
C37311 AND2X1_LOC_112/a_8_24# OR2X1_LOC_31/Y 0.01fF
C37400 OR2X1_LOC_298/Y OR2X1_LOC_31/Y 0.13fF
C37931 OR2X1_LOC_31/Y OR2X1_LOC_595/Y 0.01fF
C38287 AND2X1_LOC_197/a_8_24# OR2X1_LOC_31/Y 0.01fF
C38332 OR2X1_LOC_31/Y OR2X1_LOC_409/Y 0.10fF
C39001 OR2X1_LOC_31/Y OR2X1_LOC_12/Y 1.38fF
C39008 OR2X1_LOC_31/Y OR2X1_LOC_766/Y 0.21fF
C39164 OR2X1_LOC_272/Y OR2X1_LOC_31/Y 0.03fF
C39505 OR2X1_LOC_517/a_8_216# OR2X1_LOC_31/Y 0.05fF
C39929 OR2X1_LOC_31/Y AND2X1_LOC_520/Y 0.04fF
C40872 AND2X1_LOC_318/Y OR2X1_LOC_31/Y 0.16fF
C41325 OR2X1_LOC_31/Y OR2X1_LOC_224/Y 0.01fF
C41676 OR2X1_LOC_18/Y OR2X1_LOC_31/Y 0.22fF
C42415 OR2X1_LOC_31/Y OR2X1_LOC_230/Y 0.01fF
C42421 OR2X1_LOC_31/Y OR2X1_LOC_368/Y 0.01fF
C42750 OR2X1_LOC_31/Y OR2X1_LOC_437/A 0.07fF
C42904 AND2X1_LOC_715/A OR2X1_LOC_31/Y 0.01fF
C43296 OR2X1_LOC_31/Y OR2X1_LOC_323/Y 0.04fF
C43410 AND2X1_LOC_729/Y OR2X1_LOC_31/Y 0.01fF
C43483 OR2X1_LOC_31/Y AND2X1_LOC_639/A 0.02fF
C43578 OR2X1_LOC_31/Y OR2X1_LOC_172/Y 0.43fF
C43883 OR2X1_LOC_31/Y OR2X1_LOC_52/B 0.25fF
C44179 OR2X1_LOC_31/Y OR2X1_LOC_584/Y 0.32fF
C44320 OR2X1_LOC_280/Y OR2X1_LOC_31/Y 0.22fF
C44351 OR2X1_LOC_22/Y OR2X1_LOC_31/Y 0.54fF
C44632 OR2X1_LOC_485/Y OR2X1_LOC_31/Y 0.03fF
C44703 OR2X1_LOC_31/Y OR2X1_LOC_39/A 0.30fF
C44794 OR2X1_LOC_31/Y OR2X1_LOC_428/a_8_216# 0.07fF
C45152 AND2X1_LOC_593/Y OR2X1_LOC_31/Y 0.01fF
C45468 AND2X1_LOC_332/a_8_24# OR2X1_LOC_31/Y 0.03fF
C45519 OR2X1_LOC_51/Y OR2X1_LOC_31/Y 0.21fF
C45562 OR2X1_LOC_31/Y OR2X1_LOC_16/Y 0.02fF
C47360 AND2X1_LOC_197/Y OR2X1_LOC_31/Y 0.01fF
C47638 OR2X1_LOC_31/Y OR2X1_LOC_183/Y 0.01fF
C47834 OR2X1_LOC_31/Y OR2X1_LOC_511/Y 0.03fF
C48202 OR2X1_LOC_600/a_8_216# OR2X1_LOC_31/Y 0.07fF
C48530 OR2X1_LOC_518/Y OR2X1_LOC_31/Y 0.27fF
C48619 OR2X1_LOC_91/A OR2X1_LOC_31/Y 0.60fF
C49075 OR2X1_LOC_32/B OR2X1_LOC_31/Y 0.11fF
C49251 OR2X1_LOC_31/Y OR2X1_LOC_423/Y 0.02fF
C49570 OR2X1_LOC_31/Y OR2X1_LOC_74/A 0.36fF
C50378 OR2X1_LOC_31/Y OR2X1_LOC_432/Y 0.26fF
C51088 AND2X1_LOC_339/B OR2X1_LOC_31/Y 0.08fF
C52167 OR2X1_LOC_31/Y OR2X1_LOC_72/Y 0.03fF
C52507 OR2X1_LOC_696/Y OR2X1_LOC_31/Y 0.03fF
C52859 AND2X1_LOC_198/a_8_24# OR2X1_LOC_31/Y 0.02fF
C52887 OR2X1_LOC_31/Y OR2X1_LOC_595/a_8_216# 0.01fF
C53197 AND2X1_LOC_706/Y OR2X1_LOC_31/Y 0.11fF
C53227 OR2X1_LOC_58/Y OR2X1_LOC_31/Y 0.01fF
C53330 OR2X1_LOC_485/A OR2X1_LOC_31/Y 1.58fF
C54729 OR2X1_LOC_31/Y OR2X1_LOC_589/Y 0.01fF
C55784 OR2X1_LOC_526/Y OR2X1_LOC_31/Y 0.01fF
C55862 OR2X1_LOC_31/Y OR2X1_LOC_433/Y 0.49fF
C56205 AND2X1_LOC_714/B OR2X1_LOC_31/Y 0.09fF
C57053 OR2X1_LOC_31/Y VSS 0.86fF
C44 OR2X1_LOC_18/Y AND2X1_LOC_687/Y 0.06fF
C47 OR2X1_LOC_18/Y AND2X1_LOC_630/a_8_24# 0.03fF
C283 OR2X1_LOC_666/a_8_216# OR2X1_LOC_18/Y 0.07fF
C801 OR2X1_LOC_109/Y OR2X1_LOC_18/Y 0.01fF
C894 OR2X1_LOC_18/Y AND2X1_LOC_729/B 0.03fF
C1388 AND2X1_LOC_227/Y OR2X1_LOC_18/Y 0.05fF
C1412 OR2X1_LOC_18/Y OR2X1_LOC_813/Y 0.01fF
C1716 OR2X1_LOC_599/A OR2X1_LOC_18/Y 0.02fF
C2007 OR2X1_LOC_40/Y OR2X1_LOC_18/Y 1.17fF
C2088 AND2X1_LOC_843/Y OR2X1_LOC_18/Y 0.03fF
C2168 OR2X1_LOC_18/Y OR2X1_LOC_7/A 0.31fF
C3283 AND2X1_LOC_706/a_8_24# OR2X1_LOC_18/Y 0.04fF
C3294 OR2X1_LOC_589/A OR2X1_LOC_18/Y 0.20fF
C3385 OR2X1_LOC_18/Y OR2X1_LOC_495/Y 0.03fF
C3593 OR2X1_LOC_18/Y OR2X1_LOC_384/a_8_216# 0.14fF
C3729 AND2X1_LOC_776/a_8_24# OR2X1_LOC_18/Y 0.01fF
C4257 OR2X1_LOC_3/Y OR2X1_LOC_18/Y 9.00fF
C5473 OR2X1_LOC_173/Y OR2X1_LOC_18/Y 0.02fF
C5475 OR2X1_LOC_18/Y OR2X1_LOC_690/A 0.03fF
C5531 OR2X1_LOC_64/Y OR2X1_LOC_18/Y 0.38fF
C5556 OR2X1_LOC_18/Y AND2X1_LOC_632/A 0.03fF
C5928 AND2X1_LOC_101/B OR2X1_LOC_18/Y 0.71fF
C6819 OR2X1_LOC_18/Y OR2X1_LOC_279/Y 0.19fF
C7130 AND2X1_LOC_456/B OR2X1_LOC_18/Y 0.04fF
C7496 OR2X1_LOC_18/Y AND2X1_LOC_828/a_8_24# 0.01fF
C7982 OR2X1_LOC_494/Y OR2X1_LOC_18/Y 0.05fF
C8175 OR2X1_LOC_18/Y AND2X1_LOC_116/B 0.01fF
C8825 OR2X1_LOC_18/Y AND2X1_LOC_778/Y 0.20fF
C8910 OR2X1_LOC_521/Y OR2X1_LOC_18/Y 0.32fF
C8942 OR2X1_LOC_18/Y AND2X1_LOC_624/A 0.03fF
C11003 OR2X1_LOC_18/Y OR2X1_LOC_278/Y 0.02fF
C11254 OR2X1_LOC_18/Y OR2X1_LOC_504/a_8_216# 0.01fF
C11281 OR2X1_LOC_18/Y OR2X1_LOC_89/Y 0.09fF
C11517 AND2X1_LOC_78/a_8_24# OR2X1_LOC_18/Y 0.03fF
C11683 OR2X1_LOC_18/Y OR2X1_LOC_142/Y 0.03fF
C11880 OR2X1_LOC_18/Y OR2X1_LOC_118/Y 0.03fF
C11927 OR2X1_LOC_18/Y OR2X1_LOC_238/Y 0.03fF
C11929 OR2X1_LOC_18/Y OR2X1_LOC_24/Y 0.65fF
C12767 OR2X1_LOC_18/Y OR2X1_LOC_36/Y 1.09fF
C12912 OR2X1_LOC_18/Y OR2X1_LOC_419/Y 0.05fF
C13067 OR2X1_LOC_315/a_8_216# OR2X1_LOC_18/Y 0.01fF
C13103 OR2X1_LOC_604/A OR2X1_LOC_18/Y 0.06fF
C13986 OR2X1_LOC_164/Y OR2X1_LOC_18/Y 1.16fF
C14759 OR2X1_LOC_20/Y OR2X1_LOC_18/Y 0.02fF
C15298 OR2X1_LOC_764/Y OR2X1_LOC_18/Y 0.01fF
C16376 OR2X1_LOC_18/Y OR2X1_LOC_12/Y 2.67fF
C16477 OR2X1_LOC_837/Y OR2X1_LOC_18/Y 0.09fF
C16594 OR2X1_LOC_272/Y OR2X1_LOC_18/Y 0.08fF
C16792 AND2X1_LOC_776/Y OR2X1_LOC_18/Y 0.09fF
C17030 OR2X1_LOC_79/A OR2X1_LOC_18/Y 0.15fF
C17446 OR2X1_LOC_18/Y OR2X1_LOC_617/Y 0.04fF
C17466 OR2X1_LOC_18/Y AND2X1_LOC_464/Y 0.03fF
C18152 OR2X1_LOC_597/A OR2X1_LOC_18/Y 0.01fF
C18555 OR2X1_LOC_18/Y OR2X1_LOC_829/A 0.01fF
C19392 OR2X1_LOC_18/Y OR2X1_LOC_764/a_8_216# 0.01fF
C19825 OR2X1_LOC_18/Y OR2X1_LOC_230/Y 0.07fF
C20189 OR2X1_LOC_18/Y OR2X1_LOC_437/A 0.08fF
C20296 AND2X1_LOC_715/A OR2X1_LOC_18/Y 0.37fF
C20871 AND2X1_LOC_778/a_8_24# OR2X1_LOC_18/Y 0.02fF
C20887 AND2X1_LOC_769/a_8_24# OR2X1_LOC_18/Y 0.02fF
C20950 OR2X1_LOC_18/Y AND2X1_LOC_639/A 0.01fF
C21009 OR2X1_LOC_18/Y OR2X1_LOC_172/Y 0.07fF
C21315 OR2X1_LOC_18/Y OR2X1_LOC_52/B 0.38fF
C21443 OR2X1_LOC_18/Y AND2X1_LOC_216/A 0.27fF
C21715 OR2X1_LOC_18/Y AND2X1_LOC_286/Y 0.02fF
C21756 OR2X1_LOC_280/Y OR2X1_LOC_18/Y 0.03fF
C21802 OR2X1_LOC_22/Y OR2X1_LOC_18/Y 0.92fF
C22144 OR2X1_LOC_18/Y OR2X1_LOC_39/A 0.31fF
C22638 AND2X1_LOC_78/a_36_24# OR2X1_LOC_18/Y 0.01fF
C22925 OR2X1_LOC_51/Y OR2X1_LOC_18/Y 0.27fF
C23012 OR2X1_LOC_680/A OR2X1_LOC_18/Y 0.06fF
C23976 OR2X1_LOC_18/Y OR2X1_LOC_86/A 0.03fF
C24638 OR2X1_LOC_18/Y OR2X1_LOC_616/a_8_216# 0.18fF
C25666 OR2X1_LOC_18/Y OR2X1_LOC_384/Y 0.04fF
C25810 OR2X1_LOC_91/A OR2X1_LOC_18/Y 0.12fF
C25913 OR2X1_LOC_669/Y OR2X1_LOC_18/Y 0.16fF
C26346 OR2X1_LOC_18/Y OR2X1_LOC_371/Y 0.08fF
C26789 OR2X1_LOC_18/Y OR2X1_LOC_74/A 0.19fF
C27072 OR2X1_LOC_18/Y OR2X1_LOC_626/Y 0.12fF
C27165 OR2X1_LOC_432/a_8_216# OR2X1_LOC_18/Y 0.01fF
C27195 OR2X1_LOC_18/Y AND2X1_LOC_287/Y 0.02fF
C28315 AND2X1_LOC_339/B OR2X1_LOC_18/Y 0.03fF
C28605 OR2X1_LOC_18/Y OR2X1_LOC_521/a_8_216# 0.01fF
C28617 OR2X1_LOC_18/Y OR2X1_LOC_300/Y 0.03fF
C28738 OR2X1_LOC_505/Y OR2X1_LOC_18/Y 0.01fF
C30408 AND2X1_LOC_706/Y OR2X1_LOC_18/Y 0.01fF
C30528 AND2X1_LOC_303/A OR2X1_LOC_18/Y 4.38fF
C30572 OR2X1_LOC_485/A OR2X1_LOC_18/Y 0.82fF
C31391 OR2X1_LOC_18/Y AND2X1_LOC_458/Y 0.01fF
C31418 OR2X1_LOC_18/Y OR2X1_LOC_89/a_8_216# 0.04fF
C32430 OR2X1_LOC_18/Y OR2X1_LOC_171/a_8_216# 0.01fF
C32497 OR2X1_LOC_18/Y OR2X1_LOC_13/Y 0.03fF
C32538 OR2X1_LOC_18/Y OR2X1_LOC_627/Y 0.19fF
C33831 OR2X1_LOC_496/a_8_216# OR2X1_LOC_18/Y 0.01fF
C34132 OR2X1_LOC_516/Y OR2X1_LOC_18/Y 0.03fF
C35209 OR2X1_LOC_131/Y OR2X1_LOC_18/Y 0.03fF
C35489 VDD OR2X1_LOC_18/Y 1.26fF
C35544 AND2X1_LOC_208/B OR2X1_LOC_18/Y 0.02fF
C35588 OR2X1_LOC_315/Y OR2X1_LOC_18/Y 0.53fF
C35630 OR2X1_LOC_251/Y OR2X1_LOC_18/Y 0.02fF
C35738 OR2X1_LOC_18/Y OR2X1_LOC_67/Y 0.05fF
C36667 OR2X1_LOC_494/A OR2X1_LOC_18/Y 0.02fF
C36807 OR2X1_LOC_18/Y OR2X1_LOC_427/A 0.46fF
C36835 OR2X1_LOC_18/Y AND2X1_LOC_464/a_8_24# 0.02fF
C37352 OR2X1_LOC_18/Y OR2X1_LOC_416/Y 0.03fF
C38089 OR2X1_LOC_18/Y OR2X1_LOC_45/a_8_216# 0.02fF
C38166 OR2X1_LOC_18/Y AND2X1_LOC_116/Y 0.01fF
C38171 OR2X1_LOC_18/Y OR2X1_LOC_20/a_8_216# 0.01fF
C38376 OR2X1_LOC_45/B OR2X1_LOC_18/Y 11.02fF
C38545 OR2X1_LOC_18/Y OR2X1_LOC_767/a_8_216# 0.05fF
C38871 OR2X1_LOC_158/A OR2X1_LOC_18/Y 2.18fF
C39298 OR2X1_LOC_482/Y OR2X1_LOC_18/Y 0.03fF
C39395 OR2X1_LOC_18/Y OR2X1_LOC_586/Y 0.42fF
C39517 OR2X1_LOC_18/Y OR2X1_LOC_628/Y 0.06fF
C39708 AND2X1_LOC_195/a_8_24# OR2X1_LOC_18/Y 0.06fF
C41099 OR2X1_LOC_316/Y OR2X1_LOC_18/Y 0.11fF
C41476 OR2X1_LOC_744/A OR2X1_LOC_18/Y 6.11fF
C41575 OR2X1_LOC_18/Y AND2X1_LOC_840/B 0.05fF
C41833 OR2X1_LOC_18/Y OR2X1_LOC_79/a_8_216# 0.05fF
C41843 OR2X1_LOC_18/Y AND2X1_LOC_464/A 0.64fF
C42280 OR2X1_LOC_18/Y OR2X1_LOC_522/Y 0.12fF
C42465 AND2X1_LOC_303/B OR2X1_LOC_18/Y 0.39fF
C42781 OR2X1_LOC_18/Y OR2X1_LOC_56/A 4.63fF
C42821 OR2X1_LOC_18/Y AND2X1_LOC_638/Y 0.05fF
C43297 OR2X1_LOC_91/Y OR2X1_LOC_18/Y 0.03fF
C43362 OR2X1_LOC_527/Y OR2X1_LOC_18/Y 0.06fF
C43545 OR2X1_LOC_18/Y OR2X1_LOC_171/Y 0.52fF
C43652 OR2X1_LOC_18/Y AND2X1_LOC_629/a_8_24# 0.03fF
C43785 OR2X1_LOC_18/Y AND2X1_LOC_276/Y 0.16fF
C44161 OR2X1_LOC_18/Y AND2X1_LOC_139/B 3.31fF
C44661 OR2X1_LOC_481/A OR2X1_LOC_18/Y 0.02fF
C44692 OR2X1_LOC_18/Y OR2X1_LOC_71/Y 1.49fF
C44727 OR2X1_LOC_18/Y OR2X1_LOC_173/a_8_216# 0.01fF
C45124 OR2X1_LOC_18/Y OR2X1_LOC_246/A 0.13fF
C45154 OR2X1_LOC_18/Y OR2X1_LOC_409/B 0.05fF
C45930 OR2X1_LOC_18/Y OR2X1_LOC_24/a_8_216# 0.01fF
C46512 OR2X1_LOC_18/Y AND2X1_LOC_721/A 0.02fF
C46811 AND2X1_LOC_318/a_8_24# OR2X1_LOC_18/Y 0.04fF
C46838 OR2X1_LOC_18/Y AND2X1_LOC_361/A 0.07fF
C47548 OR2X1_LOC_18/Y AND2X1_LOC_284/a_8_24# 0.01fF
C48133 OR2X1_LOC_18/Y OR2X1_LOC_257/a_8_216# 0.02fF
C48145 OR2X1_LOC_18/Y OR2X1_LOC_65/B 0.05fF
C48441 OR2X1_LOC_692/Y OR2X1_LOC_18/Y 0.01fF
C48481 OR2X1_LOC_600/A OR2X1_LOC_18/Y 0.23fF
C48554 OR2X1_LOC_18/Y OR2X1_LOC_619/Y 0.03fF
C48818 OR2X1_LOC_18/Y AND2X1_LOC_769/Y 0.01fF
C49397 OR2X1_LOC_18/Y OR2X1_LOC_45/a_36_216# 0.02fF
C49518 OR2X1_LOC_813/A OR2X1_LOC_18/Y 0.01fF
C49568 OR2X1_LOC_18/Y OR2X1_LOC_406/A 0.02fF
C49685 OR2X1_LOC_505/a_8_216# OR2X1_LOC_18/Y 0.02fF
C50880 OR2X1_LOC_18/Y OR2X1_LOC_13/B 0.35fF
C51350 OR2X1_LOC_18/Y OR2X1_LOC_428/A 0.18fF
C51364 OR2X1_LOC_18/Y OR2X1_LOC_595/A 0.14fF
C51809 OR2X1_LOC_528/Y OR2X1_LOC_18/Y 0.16fF
C51965 OR2X1_LOC_18/Y OR2X1_LOC_279/a_8_216# 0.02fF
C52371 OR2X1_LOC_18/Y OR2X1_LOC_26/Y 0.19fF
C52390 OR2X1_LOC_18/Y OR2X1_LOC_89/A 0.18fF
C53035 OR2X1_LOC_18/Y AND2X1_LOC_473/Y 0.84fF
C53166 OR2X1_LOC_45/Y OR2X1_LOC_18/Y 0.23fF
C53294 OR2X1_LOC_18/Y OR2X1_LOC_95/Y 4.92fF
C53615 OR2X1_LOC_18/Y OR2X1_LOC_257/a_36_216# 0.03fF
C53891 OR2X1_LOC_693/Y OR2X1_LOC_18/Y 0.01fF
C54009 OR2X1_LOC_18/Y AND2X1_LOC_621/Y 0.06fF
C54354 OR2X1_LOC_18/Y OR2X1_LOC_59/Y 0.68fF
C54488 OR2X1_LOC_70/Y OR2X1_LOC_18/Y 0.72fF
C54540 OR2X1_LOC_504/Y OR2X1_LOC_18/Y 0.01fF
C54572 OR2X1_LOC_18/Y OR2X1_LOC_184/Y 0.54fF
C55186 OR2X1_LOC_18/Y OR2X1_LOC_607/A 0.01fF
C55283 OR2X1_LOC_625/Y OR2X1_LOC_18/Y 0.03fF
C55529 OR2X1_LOC_18/Y OR2X1_LOC_767/Y 0.02fF
C56013 OR2X1_LOC_18/Y OR2X1_LOC_16/A 0.12fF
C57234 OR2X1_LOC_18/Y VSS 1.25fF
C82 OR2X1_LOC_59/Y OR2X1_LOC_172/Y 0.01fF
C361 OR2X1_LOC_59/Y OR2X1_LOC_52/B 0.27fF
C397 OR2X1_LOC_755/A OR2X1_LOC_59/Y 0.05fF
C487 AND2X1_LOC_216/A OR2X1_LOC_59/Y 0.16fF
C621 OR2X1_LOC_281/Y OR2X1_LOC_59/Y 0.03fF
C753 OR2X1_LOC_59/Y AND2X1_LOC_286/Y 0.17fF
C802 OR2X1_LOC_280/Y OR2X1_LOC_59/Y 0.03fF
C844 OR2X1_LOC_295/a_36_216# OR2X1_LOC_59/Y 0.03fF
C851 OR2X1_LOC_22/Y OR2X1_LOC_59/Y 0.21fF
C1101 OR2X1_LOC_485/Y OR2X1_LOC_59/Y 0.43fF
C1203 OR2X1_LOC_59/Y OR2X1_LOC_39/A 6.03fF
C1615 AND2X1_LOC_593/Y OR2X1_LOC_59/Y 0.02fF
C1970 OR2X1_LOC_51/Y OR2X1_LOC_59/Y 4.85fF
C2060 OR2X1_LOC_680/A OR2X1_LOC_59/Y 0.11fF
C2837 OR2X1_LOC_178/a_8_216# OR2X1_LOC_59/Y 0.01fF
C3375 OR2X1_LOC_81/a_8_216# OR2X1_LOC_59/Y 0.07fF
C3529 OR2X1_LOC_59/Y OR2X1_LOC_331/a_8_216# 0.01fF
C4010 OR2X1_LOC_59/Y OR2X1_LOC_183/Y 0.04fF
C4151 OR2X1_LOC_511/Y OR2X1_LOC_59/Y 0.03fF
C4193 OR2X1_LOC_297/Y OR2X1_LOC_59/Y 0.01fF
C4894 OR2X1_LOC_91/A OR2X1_LOC_59/Y 0.08fF
C4999 OR2X1_LOC_669/Y OR2X1_LOC_59/Y 0.82fF
C5370 OR2X1_LOC_32/B OR2X1_LOC_59/Y 0.11fF
C5432 OR2X1_LOC_59/Y OR2X1_LOC_371/Y 0.07fF
C5896 OR2X1_LOC_74/A OR2X1_LOC_59/Y 0.31fF
C6150 OR2X1_LOC_59/Y OR2X1_LOC_626/Y 0.08fF
C6248 OR2X1_LOC_59/Y AND2X1_LOC_287/Y 0.03fF
C6665 OR2X1_LOC_59/Y AND2X1_LOC_287/a_8_24# 0.01fF
C7450 AND2X1_LOC_339/B OR2X1_LOC_59/Y 0.07fF
C7456 OR2X1_LOC_482/a_8_216# OR2X1_LOC_59/Y 0.01fF
C7804 OR2X1_LOC_59/Y OR2X1_LOC_300/Y 0.08fF
C7842 OR2X1_LOC_106/Y OR2X1_LOC_59/Y 0.03fF
C8005 AND2X1_LOC_847/Y OR2X1_LOC_59/Y 0.01fF
C8373 AND2X1_LOC_614/a_8_24# OR2X1_LOC_59/Y 0.06fF
C8666 OR2X1_LOC_59/Y OR2X1_LOC_72/Y 0.02fF
C9391 OR2X1_LOC_431/a_8_216# OR2X1_LOC_59/Y 0.01fF
C9630 OR2X1_LOC_58/Y OR2X1_LOC_59/Y 0.01fF
C9747 AND2X1_LOC_303/A OR2X1_LOC_59/Y 4.37fF
C9762 OR2X1_LOC_81/Y OR2X1_LOC_59/Y 0.03fF
C9786 OR2X1_LOC_485/A OR2X1_LOC_59/Y 1.11fF
C10572 AND2X1_LOC_302/a_8_24# OR2X1_LOC_59/Y 0.04fF
C10606 OR2X1_LOC_89/a_8_216# OR2X1_LOC_59/Y 0.07fF
C11423 OR2X1_LOC_69/Y OR2X1_LOC_59/Y 0.02fF
C11554 OR2X1_LOC_437/a_8_216# OR2X1_LOC_59/Y 0.04fF
C11719 OR2X1_LOC_13/Y OR2X1_LOC_59/Y 0.03fF
C11823 OR2X1_LOC_700/Y OR2X1_LOC_59/Y 0.01fF
C12150 OR2X1_LOC_526/Y OR2X1_LOC_59/Y 0.01fF
C13008 OR2X1_LOC_492/a_8_216# OR2X1_LOC_59/Y 0.06fF
C13746 OR2X1_LOC_59/Y OR2X1_LOC_533/A 0.44fF
C14445 OR2X1_LOC_609/a_8_216# OR2X1_LOC_59/Y 0.02fF
C14718 VDD OR2X1_LOC_59/Y 1.25fF
C14827 OR2X1_LOC_491/Y OR2X1_LOC_59/Y 0.03fF
C14833 OR2X1_LOC_251/Y OR2X1_LOC_59/Y 0.03fF
C15131 OR2X1_LOC_60/Y OR2X1_LOC_59/Y 0.01fF
C15242 OR2X1_LOC_666/Y OR2X1_LOC_59/Y 0.09fF
C16024 OR2X1_LOC_427/A OR2X1_LOC_59/Y 0.35fF
C16567 OR2X1_LOC_416/Y OR2X1_LOC_59/Y 0.04fF
C16889 OR2X1_LOC_281/a_8_216# OR2X1_LOC_59/Y 0.03fF
C17297 OR2X1_LOC_485/a_8_216# OR2X1_LOC_59/Y 0.01fF
C17322 OR2X1_LOC_45/a_8_216# OR2X1_LOC_59/Y 0.02fF
C17323 OR2X1_LOC_701/Y OR2X1_LOC_59/Y 0.01fF
C17386 AND2X1_LOC_116/Y OR2X1_LOC_59/Y 1.06fF
C17596 OR2X1_LOC_45/B OR2X1_LOC_59/Y 5.59fF
C17742 OR2X1_LOC_59/Y OR2X1_LOC_767/a_8_216# 0.01fF
C18072 OR2X1_LOC_158/A OR2X1_LOC_59/Y 0.22fF
C18522 OR2X1_LOC_482/Y OR2X1_LOC_59/Y 0.29fF
C18659 OR2X1_LOC_748/A OR2X1_LOC_59/Y 0.02fF
C18711 OR2X1_LOC_304/Y OR2X1_LOC_59/Y 0.21fF
C18747 OR2X1_LOC_628/Y OR2X1_LOC_59/Y 0.07fF
C19052 AND2X1_LOC_848/a_8_24# OR2X1_LOC_59/Y 0.02fF
C19680 AND2X1_LOC_848/A OR2X1_LOC_59/Y 0.05fF
C19983 OR2X1_LOC_609/a_36_216# OR2X1_LOC_59/Y 0.03fF
C20330 OR2X1_LOC_316/Y OR2X1_LOC_59/Y 0.04fF
C20424 OR2X1_LOC_431/Y OR2X1_LOC_59/Y 0.01fF
C20696 OR2X1_LOC_744/A OR2X1_LOC_59/Y 10.06fF
C20780 AND2X1_LOC_840/B OR2X1_LOC_59/Y 0.07fF
C20793 OR2X1_LOC_74/a_8_216# OR2X1_LOC_59/Y 0.02fF
C21047 OR2X1_LOC_79/a_8_216# OR2X1_LOC_59/Y 0.01fF
C21101 AND2X1_LOC_301/a_8_24# OR2X1_LOC_59/Y 0.14fF
C21588 OR2X1_LOC_179/a_8_216# OR2X1_LOC_59/Y 0.01fF
C21983 OR2X1_LOC_56/A OR2X1_LOC_59/Y 8.72fF
C22480 OR2X1_LOC_281/a_36_216# OR2X1_LOC_59/Y 0.02fF
C22516 OR2X1_LOC_91/Y OR2X1_LOC_59/Y 0.16fF
C22568 OR2X1_LOC_59/Y OR2X1_LOC_757/Y 0.01fF
C22588 OR2X1_LOC_527/Y OR2X1_LOC_59/Y 0.07fF
C22600 OR2X1_LOC_291/Y OR2X1_LOC_59/Y 0.26fF
C22869 AND2X1_LOC_330/a_8_24# OR2X1_LOC_59/Y 0.01fF
C22964 OR2X1_LOC_59/Y OR2X1_LOC_701/a_8_216# 0.02fF
C23001 AND2X1_LOC_276/Y OR2X1_LOC_59/Y 0.02fF
C23354 AND2X1_LOC_139/B OR2X1_LOC_59/Y 0.03fF
C23637 OR2X1_LOC_135/a_8_216# OR2X1_LOC_59/Y 0.08fF
C23841 OR2X1_LOC_481/A OR2X1_LOC_59/Y 0.37fF
C24004 OR2X1_LOC_59/Y AND2X1_LOC_789/Y 0.02fF
C24072 OR2X1_LOC_492/Y OR2X1_LOC_59/Y 0.24fF
C24086 OR2X1_LOC_108/a_8_216# OR2X1_LOC_59/Y 0.01fF
C24282 OR2X1_LOC_246/A OR2X1_LOC_59/Y 0.03fF
C24607 OR2X1_LOC_497/Y OR2X1_LOC_59/Y 0.07fF
C25614 OR2X1_LOC_59/Y OR2X1_LOC_331/Y 0.02fF
C26532 AND2X1_LOC_787/A OR2X1_LOC_59/Y 0.25fF
C27113 OR2X1_LOC_65/B OR2X1_LOC_59/Y 0.03fF
C27417 OR2X1_LOC_600/A OR2X1_LOC_59/Y 1.78fF
C27497 OR2X1_LOC_619/Y OR2X1_LOC_59/Y 0.10fF
C27850 AND2X1_LOC_286/a_8_24# OR2X1_LOC_59/Y 0.01fF
C27958 OR2X1_LOC_669/A OR2X1_LOC_59/Y 0.19fF
C28293 OR2X1_LOC_331/A OR2X1_LOC_59/Y 0.01fF
C28439 AND2X1_LOC_473/a_8_24# OR2X1_LOC_59/Y 0.01fF
C28770 OR2X1_LOC_69/A OR2X1_LOC_59/Y 0.02fF
C29856 OR2X1_LOC_59/Y OR2X1_LOC_13/B 0.54fF
C30260 OR2X1_LOC_59/Y OR2X1_LOC_533/a_8_216# -0.00fF
C30348 OR2X1_LOC_59/Y OR2X1_LOC_428/A 1.12fF
C30353 OR2X1_LOC_59/Y OR2X1_LOC_595/A 0.04fF
C30797 OR2X1_LOC_528/Y OR2X1_LOC_59/Y 0.02fF
C30901 OR2X1_LOC_516/A OR2X1_LOC_59/Y 0.03fF
C31353 OR2X1_LOC_26/Y OR2X1_LOC_59/Y 2.11fF
C31368 OR2X1_LOC_89/A OR2X1_LOC_59/Y 7.63fF
C31968 AND2X1_LOC_473/Y OR2X1_LOC_59/Y 0.01fF
C31971 AND2X1_LOC_287/B OR2X1_LOC_59/Y 0.03fF
C32009 OR2X1_LOC_491/a_8_216# OR2X1_LOC_59/Y 0.01fF
C32038 AND2X1_LOC_301/a_36_24# OR2X1_LOC_59/Y 0.01fF
C32102 OR2X1_LOC_45/Y OR2X1_LOC_59/Y 0.05fF
C32117 AND2X1_LOC_843/a_8_24# OR2X1_LOC_59/Y 0.01fF
C32212 AND2X1_LOC_727/A OR2X1_LOC_59/Y 0.03fF
C32246 OR2X1_LOC_95/Y OR2X1_LOC_59/Y 0.09fF
C32516 OR2X1_LOC_297/a_8_216# OR2X1_LOC_59/Y 0.02fF
C32518 OR2X1_LOC_179/Y OR2X1_LOC_59/Y 0.01fF
C32602 AND2X1_LOC_302/a_36_24# OR2X1_LOC_59/Y 0.01fF
C32986 AND2X1_LOC_621/Y OR2X1_LOC_59/Y 0.03fF
C33006 AND2X1_LOC_668/a_8_24# OR2X1_LOC_59/Y 0.01fF
C33509 OR2X1_LOC_70/Y OR2X1_LOC_59/Y 0.12fF
C33611 OR2X1_LOC_184/Y OR2X1_LOC_59/Y 0.01fF
C33616 OR2X1_LOC_437/Y OR2X1_LOC_59/Y 0.90fF
C34234 OR2X1_LOC_625/Y OR2X1_LOC_59/Y 0.07fF
C34495 OR2X1_LOC_59/Y OR2X1_LOC_759/Y 0.01fF
C34510 OR2X1_LOC_59/Y OR2X1_LOC_767/Y 0.02fF
C34603 OR2X1_LOC_484/Y OR2X1_LOC_59/Y 0.51fF
C35007 OR2X1_LOC_59/Y OR2X1_LOC_16/A 0.54fF
C35029 OR2X1_LOC_108/Y OR2X1_LOC_59/Y 0.37fF
C35413 OR2X1_LOC_666/a_8_216# OR2X1_LOC_59/Y 0.01fF
C35833 OR2X1_LOC_59/Y OR2X1_LOC_759/a_8_216# 0.09fF
C35941 OR2X1_LOC_109/Y OR2X1_LOC_59/Y 0.03fF
C36028 AND2X1_LOC_729/B OR2X1_LOC_59/Y 0.03fF
C36492 AND2X1_LOC_227/Y OR2X1_LOC_59/Y 0.10fF
C37103 OR2X1_LOC_40/Y OR2X1_LOC_59/Y 0.21fF
C37174 AND2X1_LOC_843/Y OR2X1_LOC_59/Y 0.02fF
C37249 OR2X1_LOC_7/A OR2X1_LOC_59/Y 0.56fF
C37345 OR2X1_LOC_224/a_8_216# OR2X1_LOC_59/Y 0.01fF
C37773 OR2X1_LOC_615/Y OR2X1_LOC_59/Y 0.03fF
C38349 OR2X1_LOC_589/A OR2X1_LOC_59/Y 0.08fF
C38398 OR2X1_LOC_297/A OR2X1_LOC_59/Y 0.03fF
C38444 OR2X1_LOC_495/Y OR2X1_LOC_59/Y 0.03fF
C38556 OR2X1_LOC_60/a_8_216# OR2X1_LOC_59/Y 0.02fF
C38992 OR2X1_LOC_299/Y OR2X1_LOC_59/Y 0.07fF
C39142 OR2X1_LOC_59/Y OR2X1_LOC_534/Y 0.25fF
C39416 OR2X1_LOC_3/Y OR2X1_LOC_59/Y 0.84fF
C39428 AND2X1_LOC_631/Y OR2X1_LOC_59/Y 0.03fF
C39738 OR2X1_LOC_74/Y OR2X1_LOC_59/Y 0.01fF
C40688 OR2X1_LOC_64/Y OR2X1_LOC_59/Y 5.89fF
C41876 OR2X1_LOC_516/B OR2X1_LOC_59/Y 0.21fF
C42037 AND2X1_LOC_196/Y OR2X1_LOC_59/Y 0.08fF
C42306 AND2X1_LOC_456/B OR2X1_LOC_59/Y 0.05fF
C43145 OR2X1_LOC_494/Y OR2X1_LOC_59/Y 0.03fF
C43323 AND2X1_LOC_116/B OR2X1_LOC_59/Y 0.02fF
C44090 AND2X1_LOC_624/A OR2X1_LOC_59/Y 0.03fF
C44438 AND2X1_LOC_434/a_8_24# OR2X1_LOC_59/Y 0.02fF
C44453 OR2X1_LOC_59/Y OR2X1_LOC_755/a_8_216# 0.03fF
C44552 OR2X1_LOC_669/a_8_216# OR2X1_LOC_59/Y 0.05fF
C45116 AND2X1_LOC_114/Y OR2X1_LOC_59/Y 0.02fF
C45392 AND2X1_LOC_114/a_8_24# OR2X1_LOC_59/Y 0.01fF
C45919 OR2X1_LOC_295/a_8_216# OR2X1_LOC_59/Y 0.09fF
C46254 OR2X1_LOC_59/Y OR2X1_LOC_278/Y 0.04fF
C46441 OR2X1_LOC_75/Y OR2X1_LOC_59/Y 0.07fF
C46574 OR2X1_LOC_89/Y OR2X1_LOC_59/Y 0.12fF
C46804 AND2X1_LOC_78/a_8_24# OR2X1_LOC_59/Y 0.01fF
C47249 OR2X1_LOC_238/Y OR2X1_LOC_59/Y 0.03fF
C47780 OR2X1_LOC_503/Y OR2X1_LOC_59/Y 0.01fF
C48096 OR2X1_LOC_36/Y OR2X1_LOC_59/Y 3.70fF
C48258 OR2X1_LOC_419/Y OR2X1_LOC_59/Y 0.09fF
C48299 OR2X1_LOC_59/Y OR2X1_LOC_526/a_8_216# 0.01fF
C48382 OR2X1_LOC_177/Y OR2X1_LOC_59/Y 0.03fF
C48408 OR2X1_LOC_604/A OR2X1_LOC_59/Y 0.50fF
C48504 OR2X1_LOC_252/a_8_216# OR2X1_LOC_59/Y 0.01fF
C48531 OR2X1_LOC_80/Y OR2X1_LOC_59/Y 0.80fF
C48769 OR2X1_LOC_533/Y OR2X1_LOC_59/Y 0.01fF
C48912 OR2X1_LOC_59/Y OR2X1_LOC_265/Y 0.03fF
C49136 OR2X1_LOC_59/Y OR2X1_LOC_183/a_8_216# 0.01fF
C49268 OR2X1_LOC_164/Y OR2X1_LOC_59/Y 0.03fF
C49434 AND2X1_LOC_633/Y OR2X1_LOC_59/Y 0.02fF
C49677 AND2X1_LOC_711/A OR2X1_LOC_59/Y 0.31fF
C50023 OR2X1_LOC_316/a_8_216# OR2X1_LOC_59/Y 0.08fF
C50520 OR2X1_LOC_700/a_8_216# OR2X1_LOC_59/Y 0.03fF
C50526 OR2X1_LOC_59/Y AND2X1_LOC_434/Y 0.01fF
C51080 AND2X1_LOC_196/a_8_24# OR2X1_LOC_59/Y 0.02fF
C51746 OR2X1_LOC_12/Y OR2X1_LOC_59/Y 0.14fF
C51912 OR2X1_LOC_272/Y OR2X1_LOC_59/Y 0.16fF
C52106 AND2X1_LOC_776/Y OR2X1_LOC_59/Y 0.78fF
C52337 OR2X1_LOC_79/A OR2X1_LOC_59/Y 0.01fF
C52368 OR2X1_LOC_278/A OR2X1_LOC_59/Y 0.14fF
C52580 OR2X1_LOC_135/Y OR2X1_LOC_59/Y 0.52fF
C52701 AND2X1_LOC_848/Y OR2X1_LOC_59/Y 0.09fF
C52733 OR2X1_LOC_283/Y OR2X1_LOC_59/Y 0.27fF
C53478 OR2X1_LOC_178/Y OR2X1_LOC_59/Y 0.04fF
C53627 OR2X1_LOC_258/Y OR2X1_LOC_59/Y 0.05fF
C53876 OR2X1_LOC_759/A OR2X1_LOC_59/Y 0.36fF
C54092 OR2X1_LOC_224/Y OR2X1_LOC_59/Y 0.01fF
C55457 OR2X1_LOC_59/Y OR2X1_LOC_437/A 4.71fF
C55587 OR2X1_LOC_59/Y OR2X1_LOC_755/Y 0.01fF
C56091 AND2X1_LOC_729/Y OR2X1_LOC_59/Y 0.03fF
C56124 AND2X1_LOC_784/A OR2X1_LOC_59/Y 0.07fF
C56613 OR2X1_LOC_59/Y VSS 1.32fF
C124 AND2X1_LOC_707/Y OR2X1_LOC_12/Y 0.13fF
C576 OR2X1_LOC_589/A OR2X1_LOC_12/Y 0.33fF
C750 OR2X1_LOC_60/a_8_216# OR2X1_LOC_12/Y 0.01fF
C1191 OR2X1_LOC_299/Y OR2X1_LOC_12/Y 0.01fF
C1613 OR2X1_LOC_3/Y OR2X1_LOC_12/Y 1.68fF
C2953 OR2X1_LOC_64/Y OR2X1_LOC_12/Y 0.23fF
C3115 OR2X1_LOC_12/Y AND2X1_LOC_247/a_8_24# 0.03fF
C4815 AND2X1_LOC_828/a_8_24# OR2X1_LOC_12/Y 0.01fF
C6082 AND2X1_LOC_130/a_8_24# OR2X1_LOC_12/Y 0.07fF
C7072 AND2X1_LOC_777/a_8_24# OR2X1_LOC_12/Y 0.01fF
C7105 OR2X1_LOC_763/Y OR2X1_LOC_12/Y 0.01fF
C7552 OR2X1_LOC_418/a_8_216# OR2X1_LOC_12/Y 0.01fF
C8386 OR2X1_LOC_12/Y OR2X1_LOC_278/Y 0.03fF
C10095 OR2X1_LOC_36/Y OR2X1_LOC_12/Y 0.30fF
C10298 OR2X1_LOC_12/Y OR2X1_LOC_526/a_8_216# 0.08fF
C10433 OR2X1_LOC_604/A OR2X1_LOC_12/Y 0.21fF
C10494 OR2X1_LOC_306/Y OR2X1_LOC_12/Y 0.05fF
C10903 OR2X1_LOC_12/Y AND2X1_LOC_447/a_8_24# -0.00fF
C11393 OR2X1_LOC_230/a_8_216# OR2X1_LOC_12/Y 0.01fF
C11632 AND2X1_LOC_539/Y OR2X1_LOC_12/Y 0.03fF
C11672 OR2X1_LOC_131/A OR2X1_LOC_12/Y 1.45fF
C12180 OR2X1_LOC_298/Y OR2X1_LOC_12/Y 0.10fF
C12304 AND2X1_LOC_678/a_8_24# OR2X1_LOC_12/Y 0.07fF
C12546 OR2X1_LOC_12/Y AND2X1_LOC_434/Y 0.03fF
C12661 OR2X1_LOC_764/Y OR2X1_LOC_12/Y 0.01fF
C13798 OR2X1_LOC_12/Y OR2X1_LOC_766/Y 0.06fF
C13966 OR2X1_LOC_272/Y OR2X1_LOC_12/Y 0.03fF
C14171 OR2X1_LOC_12/Y OR2X1_LOC_248/A 0.05fF
C14649 OR2X1_LOC_135/Y OR2X1_LOC_12/Y 0.48fF
C14994 OR2X1_LOC_12/Y OR2X1_LOC_536/a_8_216# 0.09fF
C15472 OR2X1_LOC_597/A OR2X1_LOC_12/Y 0.32fF
C15515 OR2X1_LOC_256/Y OR2X1_LOC_12/Y 0.07fF
C15559 OR2X1_LOC_313/a_8_216# OR2X1_LOC_12/Y 0.01fF
C15877 OR2X1_LOC_829/A OR2X1_LOC_12/Y 0.04fF
C16714 OR2X1_LOC_764/a_8_216# OR2X1_LOC_12/Y 0.01fF
C16970 AND2X1_LOC_634/Y OR2X1_LOC_12/Y 0.13fF
C17158 OR2X1_LOC_230/Y OR2X1_LOC_12/Y 0.21fF
C17167 OR2X1_LOC_229/a_8_216# OR2X1_LOC_12/Y 0.01fF
C17505 OR2X1_LOC_12/Y OR2X1_LOC_437/A 0.11fF
C18146 AND2X1_LOC_784/A OR2X1_LOC_12/Y 0.19fF
C18179 AND2X1_LOC_769/a_8_24# OR2X1_LOC_12/Y 0.01fF
C18243 AND2X1_LOC_639/A OR2X1_LOC_12/Y 0.02fF
C18595 OR2X1_LOC_12/Y OR2X1_LOC_52/B 0.58fF
C18780 AND2X1_LOC_216/A OR2X1_LOC_12/Y 0.02fF
C19092 OR2X1_LOC_22/Y OR2X1_LOC_12/Y 0.51fF
C19331 OR2X1_LOC_485/Y OR2X1_LOC_12/Y 0.03fF
C19417 OR2X1_LOC_12/Y OR2X1_LOC_39/A 1.16fF
C20162 OR2X1_LOC_136/Y OR2X1_LOC_12/Y 0.14fF
C20218 OR2X1_LOC_51/Y OR2X1_LOC_12/Y 1.44fF
C20627 AND2X1_LOC_593/a_36_24# OR2X1_LOC_12/Y 0.01fF
C21139 OR2X1_LOC_603/a_8_216# OR2X1_LOC_12/Y 0.08fF
C21170 OR2X1_LOC_12/Y OR2X1_LOC_588/Y 0.12fF
C21571 OR2X1_LOC_313/Y OR2X1_LOC_12/Y 0.51fF
C22441 OR2X1_LOC_511/Y OR2X1_LOC_12/Y 0.07fF
C22458 OR2X1_LOC_248/a_8_216# OR2X1_LOC_12/Y 0.02fF
C23194 OR2X1_LOC_12/Y OR2X1_LOC_131/a_8_216# 0.02fF
C23231 AND2X1_LOC_391/Y OR2X1_LOC_12/Y 0.04fF
C23233 OR2X1_LOC_91/A OR2X1_LOC_12/Y 0.41fF
C23695 OR2X1_LOC_32/B OR2X1_LOC_12/Y 0.01fF
C24180 OR2X1_LOC_490/Y OR2X1_LOC_12/Y 0.07fF
C24182 OR2X1_LOC_74/A OR2X1_LOC_12/Y 0.07fF
C24849 OR2X1_LOC_12/Y AND2X1_LOC_448/a_8_24# 0.01fF
C25262 AND2X1_LOC_704/a_8_24# OR2X1_LOC_12/Y 0.01fF
C25671 AND2X1_LOC_339/B OR2X1_LOC_12/Y 0.03fF
C26008 OR2X1_LOC_12/Y OR2X1_LOC_536/a_36_216# 0.03fF
C26011 OR2X1_LOC_12/Y OR2X1_LOC_300/Y 0.07fF
C26577 AND2X1_LOC_99/A OR2X1_LOC_12/Y 0.03fF
C26636 OR2X1_LOC_12/Y AND2X1_LOC_637/Y 0.02fF
C27770 OR2X1_LOC_12/Y OR2X1_LOC_603/Y 0.02fF
C27793 OR2X1_LOC_58/Y OR2X1_LOC_12/Y 0.40fF
C27924 OR2X1_LOC_485/A OR2X1_LOC_12/Y 1.28fF
C28360 OR2X1_LOC_420/a_8_216# OR2X1_LOC_12/Y 0.03fF
C28719 AND2X1_LOC_302/a_8_24# OR2X1_LOC_12/Y 0.01fF
C29583 OR2X1_LOC_12/Y OR2X1_LOC_418/Y 0.01fF
C29661 AND2X1_LOC_537/Y OR2X1_LOC_12/Y 0.11fF
C29894 OR2X1_LOC_13/Y OR2X1_LOC_12/Y 0.01fF
C30339 OR2X1_LOC_526/Y OR2X1_LOC_12/Y 0.01fF
C30384 OR2X1_LOC_422/Y OR2X1_LOC_12/Y 0.01fF
C30412 AND2X1_LOC_138/a_8_24# OR2X1_LOC_12/Y 0.03fF
C30721 AND2X1_LOC_714/B OR2X1_LOC_12/Y 0.01fF
C32492 OR2X1_LOC_314/Y OR2X1_LOC_12/Y 0.01fF
C32567 OR2X1_LOC_131/Y OR2X1_LOC_12/Y 0.31fF
C32851 VDD OR2X1_LOC_12/Y 0.89fF
C32941 OR2X1_LOC_12/Y AND2X1_LOC_447/a_36_24# -0.02fF
C33055 OR2X1_LOC_256/A OR2X1_LOC_12/Y 0.69fF
C33279 OR2X1_LOC_60/Y OR2X1_LOC_12/Y 0.01fF
C33317 OR2X1_LOC_314/a_8_216# OR2X1_LOC_12/Y 0.01fF
C33387 OR2X1_LOC_248/Y OR2X1_LOC_12/Y 0.10fF
C33815 OR2X1_LOC_591/A OR2X1_LOC_12/Y 0.01fF
C34170 OR2X1_LOC_427/A OR2X1_LOC_12/Y 0.21fF
C34712 OR2X1_LOC_416/Y OR2X1_LOC_12/Y 0.06fF
C35410 OR2X1_LOC_485/a_8_216# OR2X1_LOC_12/Y 0.07fF
C35471 AND2X1_LOC_831/a_8_24# OR2X1_LOC_12/Y 0.04fF
C35766 OR2X1_LOC_45/B OR2X1_LOC_12/Y 0.24fF
C36211 OR2X1_LOC_158/A OR2X1_LOC_12/Y 0.47fF
C36722 OR2X1_LOC_748/A OR2X1_LOC_12/Y 0.09fF
C36764 OR2X1_LOC_304/Y OR2X1_LOC_12/Y 0.03fF
C37981 AND2X1_LOC_317/a_8_24# OR2X1_LOC_12/Y 0.01fF
C38314 OR2X1_LOC_765/a_8_216# OR2X1_LOC_12/Y 0.07fF
C38403 OR2X1_LOC_316/Y OR2X1_LOC_12/Y 0.06fF
C38477 AND2X1_LOC_390/B OR2X1_LOC_12/Y 0.02fF
C38758 OR2X1_LOC_12/Y OR2X1_LOC_604/Y 0.01fF
C38803 OR2X1_LOC_744/A OR2X1_LOC_12/Y 1.51fF
C39138 OR2X1_LOC_12/Y OR2X1_LOC_320/a_8_216# 0.02fF
C39241 OR2X1_LOC_144/Y OR2X1_LOC_12/Y 0.08fF
C39335 OR2X1_LOC_420/Y OR2X1_LOC_12/Y 0.02fF
C40034 OR2X1_LOC_56/A OR2X1_LOC_12/Y 1.13fF
C40050 AND2X1_LOC_638/Y OR2X1_LOC_12/Y 0.03fF
C40515 OR2X1_LOC_290/Y OR2X1_LOC_12/Y 0.03fF
C40573 OR2X1_LOC_12/Y AND2X1_LOC_446/a_8_24# 0.01fF
C40630 OR2X1_LOC_417/Y OR2X1_LOC_12/Y 1.04fF
C40636 OR2X1_LOC_311/Y OR2X1_LOC_12/Y 0.02fF
C40645 AND2X1_LOC_538/Y OR2X1_LOC_12/Y 0.01fF
C40824 OR2X1_LOC_12/Y OR2X1_LOC_171/Y 0.03fF
C41104 AND2X1_LOC_831/Y OR2X1_LOC_12/Y 0.10fF
C41925 OR2X1_LOC_481/A OR2X1_LOC_12/Y 0.04fF
C41975 OR2X1_LOC_71/Y OR2X1_LOC_12/Y 0.03fF
C42410 OR2X1_LOC_246/A OR2X1_LOC_12/Y 0.53fF
C42459 OR2X1_LOC_409/B OR2X1_LOC_12/Y 0.03fF
C42703 OR2X1_LOC_298/a_8_216# OR2X1_LOC_12/Y 0.05fF
C42792 OR2X1_LOC_229/Y OR2X1_LOC_12/Y 0.06fF
C43614 AND2X1_LOC_319/A OR2X1_LOC_12/Y 0.01fF
C43735 OR2X1_LOC_604/a_8_216# OR2X1_LOC_12/Y 0.01fF
C43774 AND2X1_LOC_721/A OR2X1_LOC_12/Y 0.03fF
C44056 OR2X1_LOC_12/Y AND2X1_LOC_361/A 0.07fF
C45328 OR2X1_LOC_65/B OR2X1_LOC_12/Y 0.05fF
C45675 OR2X1_LOC_600/A OR2X1_LOC_12/Y 0.27fF
C45749 OR2X1_LOC_619/Y OR2X1_LOC_12/Y 0.14fF
C46098 OR2X1_LOC_12/Y AND2X1_LOC_769/Y 0.03fF
C46240 OR2X1_LOC_12/Y AND2X1_LOC_454/A 0.01fF
C46325 AND2X1_LOC_539/a_8_24# OR2X1_LOC_12/Y 0.01fF
C46682 AND2X1_LOC_831/a_36_24# OR2X1_LOC_12/Y 0.01fF
C47134 AND2X1_LOC_138/a_36_24# OR2X1_LOC_12/Y 0.01fF
C48272 OR2X1_LOC_12/Y OR2X1_LOC_13/B 17.89fF
C48735 OR2X1_LOC_12/Y OR2X1_LOC_428/A 1.11fF
C48745 OR2X1_LOC_12/Y OR2X1_LOC_595/A 0.07fF
C49163 AND2X1_LOC_592/Y OR2X1_LOC_12/Y 0.06fF
C49252 AND2X1_LOC_342/Y OR2X1_LOC_12/Y 0.30fF
C49372 AND2X1_LOC_712/B OR2X1_LOC_12/Y 0.12fF
C49726 OR2X1_LOC_26/Y OR2X1_LOC_12/Y 0.33fF
C49746 OR2X1_LOC_89/A OR2X1_LOC_12/Y 3.67fF
C49995 OR2X1_LOC_12/Y AND2X1_LOC_590/a_8_24# 0.04fF
C50691 OR2X1_LOC_95/Y OR2X1_LOC_12/Y 0.06fF
C51365 AND2X1_LOC_621/Y OR2X1_LOC_12/Y 0.12fF
C51862 OR2X1_LOC_70/Y OR2X1_LOC_12/Y 0.54fF
C51897 AND2X1_LOC_538/a_8_24# OR2X1_LOC_12/Y 0.09fF
C52618 OR2X1_LOC_625/Y OR2X1_LOC_12/Y 0.10fF
C53374 OR2X1_LOC_12/Y OR2X1_LOC_16/A 0.67fF
C54222 AND2X1_LOC_447/Y OR2X1_LOC_12/Y 0.16fF
C54291 AND2X1_LOC_448/Y OR2X1_LOC_12/Y 0.08fF
C54651 AND2X1_LOC_593/a_8_24# OR2X1_LOC_12/Y 0.04fF
C54846 AND2X1_LOC_227/Y OR2X1_LOC_12/Y 0.03fF
C55183 OR2X1_LOC_599/A OR2X1_LOC_12/Y 0.11fF
C55510 OR2X1_LOC_40/Y OR2X1_LOC_12/Y 0.16fF
C55627 OR2X1_LOC_7/A OR2X1_LOC_12/Y 0.90fF
C56024 OR2X1_LOC_127/Y OR2X1_LOC_12/Y 0.14fF
C56653 OR2X1_LOC_12/Y VSS 0.92fF
C2771 OR2X1_LOC_754/a_8_216# OR2X1_LOC_753/Y 0.01fF
C4056 OR2X1_LOC_22/Y OR2X1_LOC_753/Y 0.02fF
C10435 OR2X1_LOC_615/a_8_216# OR2X1_LOC_753/Y 0.40fF
C12970 OR2X1_LOC_485/A OR2X1_LOC_753/Y 0.02fF
C17929 VDD OR2X1_LOC_753/Y 0.23fF
C19271 OR2X1_LOC_427/A OR2X1_LOC_753/Y 0.33fF
C25586 AND2X1_LOC_285/Y OR2X1_LOC_753/Y 0.02fF
C34507 OR2X1_LOC_89/A OR2X1_LOC_753/Y 0.01fF
C37440 OR2X1_LOC_625/Y OR2X1_LOC_753/Y 0.05fF
C40445 OR2X1_LOC_7/A OR2X1_LOC_753/Y 0.46fF
C50037 OR2X1_LOC_754/A OR2X1_LOC_753/Y 0.27fF
C50989 OR2X1_LOC_753/Y OR2X1_LOC_754/Y 0.20fF
C51247 OR2X1_LOC_36/Y OR2X1_LOC_753/Y 0.07fF
C56495 OR2X1_LOC_753/Y VSS -0.04fF
C5477 OR2X1_LOC_450/B OR2X1_LOC_707/B 0.01fF
C11066 OR2X1_LOC_450/a_8_216# OR2X1_LOC_707/B 0.47fF
C17109 OR2X1_LOC_707/B OR2X1_LOC_449/B 0.01fF
C25865 OR2X1_LOC_707/B OR2X1_LOC_161/B 0.06fF
C26191 OR2X1_LOC_707/B OR2X1_LOC_707/a_8_216# 0.01fF
C29459 OR2X1_LOC_446/Y OR2X1_LOC_707/B 0.20fF
C30144 OR2X1_LOC_160/B OR2X1_LOC_707/B 0.26fF
C48462 OR2X1_LOC_707/B OR2X1_LOC_712/B 0.01fF
C49956 OR2X1_LOC_707/B OR2X1_LOC_87/A 0.15fF
C56210 OR2X1_LOC_450/A OR2X1_LOC_707/B 0.48fF
C57151 OR2X1_LOC_707/B VSS 0.27fF
C164 AND2X1_LOC_59/Y OR2X1_LOC_535/a_8_216# 0.14fF
C290 AND2X1_LOC_59/Y AND2X1_LOC_313/a_8_24# 0.02fF
C882 AND2X1_LOC_59/Y OR2X1_LOC_557/A 0.02fF
C1738 AND2X1_LOC_59/Y OR2X1_LOC_269/B 1.36fF
C1771 AND2X1_LOC_59/Y AND2X1_LOC_75/a_8_24# 0.11fF
C2203 AND2X1_LOC_59/Y AND2X1_LOC_176/a_8_24# 0.02fF
C2578 AND2X1_LOC_59/Y AND2X1_LOC_533/a_8_24# 0.01fF
C2718 AND2X1_LOC_59/Y AND2X1_LOC_237/a_8_24# 0.01fF
C2784 AND2X1_LOC_59/Y OR2X1_LOC_777/B 0.17fF
C2830 AND2X1_LOC_59/Y OR2X1_LOC_831/B 0.10fF
C2838 OR2X1_LOC_188/a_8_216# AND2X1_LOC_59/Y 0.01fF
C2874 AND2X1_LOC_59/Y OR2X1_LOC_344/A 0.04fF
C2987 AND2X1_LOC_59/Y OR2X1_LOC_493/A 0.20fF
C3279 AND2X1_LOC_59/Y OR2X1_LOC_161/B 0.18fF
C3412 AND2X1_LOC_59/Y AND2X1_LOC_536/a_8_24# 0.01fF
C3609 AND2X1_LOC_59/Y AND2X1_LOC_406/a_8_24# 0.01fF
C3906 AND2X1_LOC_59/Y AND2X1_LOC_67/Y 0.05fF
C4137 AND2X1_LOC_59/Y OR2X1_LOC_520/a_8_216# 0.01fF
C4235 OR2X1_LOC_644/B AND2X1_LOC_59/Y 0.14fF
C4370 AND2X1_LOC_59/Y AND2X1_LOC_609/a_8_24# 0.10fF
C4709 AND2X1_LOC_59/Y AND2X1_LOC_518/a_8_24# 0.03fF
C5536 AND2X1_LOC_59/Y OR2X1_LOC_401/A 0.09fF
C5716 AND2X1_LOC_59/Y AND2X1_LOC_7/B 0.38fF
C5860 OR2X1_LOC_319/B AND2X1_LOC_59/Y 0.05fF
C5879 AND2X1_LOC_59/Y OR2X1_LOC_318/Y 0.01fF
C6267 AND2X1_LOC_59/Y AND2X1_LOC_331/a_8_24# 0.02fF
C7238 AND2X1_LOC_59/Y OR2X1_LOC_287/B 0.04fF
C7281 AND2X1_LOC_59/Y OR2X1_LOC_76/A 0.01fF
C7539 AND2X1_LOC_59/Y OR2X1_LOC_160/B 0.48fF
C7644 AND2X1_LOC_59/Y OR2X1_LOC_553/A 0.13fF
C8423 AND2X1_LOC_59/Y OR2X1_LOC_151/A 0.17fF
C8926 AND2X1_LOC_59/Y AND2X1_LOC_482/a_8_24# 0.11fF
C10022 AND2X1_LOC_59/Y OR2X1_LOC_168/Y 0.02fF
C10299 AND2X1_LOC_59/Y OR2X1_LOC_520/B 0.01fF
C10847 AND2X1_LOC_59/Y OR2X1_LOC_308/Y 0.07fF
C11487 AND2X1_LOC_59/Y OR2X1_LOC_664/Y 0.19fF
C11988 AND2X1_LOC_59/Y AND2X1_LOC_7/Y 0.11fF
C13129 AND2X1_LOC_59/Y OR2X1_LOC_841/A 0.06fF
C13698 AND2X1_LOC_59/Y OR2X1_LOC_473/Y 0.01fF
C13761 AND2X1_LOC_59/Y OR2X1_LOC_241/B 0.05fF
C13887 OR2X1_LOC_188/Y AND2X1_LOC_59/Y 0.01fF
C14341 AND2X1_LOC_59/Y OR2X1_LOC_831/A 0.01fF
C14353 AND2X1_LOC_59/Y OR2X1_LOC_598/Y 0.03fF
C14461 AND2X1_LOC_59/Y OR2X1_LOC_537/A 0.01fF
C14751 AND2X1_LOC_59/Y OR2X1_LOC_356/A 0.21fF
C15303 AND2X1_LOC_59/Y OR2X1_LOC_810/A 0.04fF
C15584 OR2X1_LOC_715/B AND2X1_LOC_59/Y 0.08fF
C15712 AND2X1_LOC_59/Y AND2X1_LOC_81/a_8_24# 0.06fF
C16099 OR2X1_LOC_656/B AND2X1_LOC_59/Y 0.03fF
C16855 AND2X1_LOC_59/Y OR2X1_LOC_535/A 0.01fF
C17328 AND2X1_LOC_59/Y OR2X1_LOC_78/A 0.25fF
C17832 AND2X1_LOC_59/Y OR2X1_LOC_97/B 0.05fF
C18434 AND2X1_LOC_59/Y OR2X1_LOC_318/B 0.04fF
C18445 AND2X1_LOC_59/Y OR2X1_LOC_854/A 0.04fF
C18597 OR2X1_LOC_114/B AND2X1_LOC_59/Y 0.02fF
C18642 AND2X1_LOC_59/Y OR2X1_LOC_538/A 0.02fF
C18710 AND2X1_LOC_12/Y AND2X1_LOC_59/Y 0.39fF
C18743 AND2X1_LOC_59/Y OR2X1_LOC_841/B 0.01fF
C18776 AND2X1_LOC_59/Y AND2X1_LOC_79/Y 0.16fF
C19059 AND2X1_LOC_59/Y OR2X1_LOC_168/B 0.22fF
C19422 OR2X1_LOC_318/a_8_216# AND2X1_LOC_59/Y 0.01fF
C19955 AND2X1_LOC_59/Y OR2X1_LOC_776/a_8_216# 0.01fF
C19987 AND2X1_LOC_59/Y OR2X1_LOC_833/B 0.02fF
C21332 AND2X1_LOC_59/Y OR2X1_LOC_84/B 0.28fF
C21398 AND2X1_LOC_59/Y OR2X1_LOC_520/A 0.01fF
C21573 OR2X1_LOC_186/Y AND2X1_LOC_59/Y 0.77fF
C21722 AND2X1_LOC_59/Y AND2X1_LOC_81/B 0.46fF
C22051 AND2X1_LOC_59/Y OR2X1_LOC_493/B 0.23fF
C22192 AND2X1_LOC_59/Y OR2X1_LOC_574/A 0.06fF
C22549 AND2X1_LOC_59/Y AND2X1_LOC_58/a_8_24# 0.01fF
C22826 AND2X1_LOC_59/Y OR2X1_LOC_539/B 0.02fF
C22944 AND2X1_LOC_59/Y OR2X1_LOC_78/B 0.20fF
C23020 AND2X1_LOC_59/Y OR2X1_LOC_375/A 1.23fF
C23291 AND2X1_LOC_59/Y OR2X1_LOC_549/A 0.06fF
C24990 AND2X1_LOC_59/Y AND2X1_LOC_19/Y 0.62fF
C25092 AND2X1_LOC_59/Y OR2X1_LOC_673/Y 0.02fF
C25746 AND2X1_LOC_59/Y OR2X1_LOC_139/A 0.03fF
C26813 AND2X1_LOC_59/Y AND2X1_LOC_666/a_8_24# 0.01fF
C27197 OR2X1_LOC_703/B AND2X1_LOC_59/Y 0.02fF
C27205 AND2X1_LOC_59/Y OR2X1_LOC_87/A 0.38fF
C27489 AND2X1_LOC_59/Y OR2X1_LOC_389/A 0.01fF
C27620 AND2X1_LOC_59/Y OR2X1_LOC_403/B 0.23fF
C27988 AND2X1_LOC_59/Y OR2X1_LOC_61/B 0.14fF
C28296 AND2X1_LOC_59/Y OR2X1_LOC_97/A 0.10fF
C28386 AND2X1_LOC_59/Y OR2X1_LOC_541/A 0.01fF
C28407 AND2X1_LOC_59/Y OR2X1_LOC_475/B 0.04fF
C28706 AND2X1_LOC_59/Y OR2X1_LOC_691/Y 0.03fF
C29181 AND2X1_LOC_700/a_8_24# AND2X1_LOC_59/Y 0.01fF
C29324 AND2X1_LOC_59/Y OR2X1_LOC_333/B 0.03fF
C29707 OR2X1_LOC_154/A AND2X1_LOC_59/Y 0.32fF
C29771 AND2X1_LOC_59/Y OR2X1_LOC_778/A 0.02fF
C30137 AND2X1_LOC_59/Y AND2X1_LOC_395/a_8_24# 0.09fF
C30251 AND2X1_LOC_59/Y AND2X1_LOC_813/a_8_24# 0.17fF
C30989 AND2X1_LOC_59/Y OR2X1_LOC_520/Y 0.04fF
C31713 AND2X1_LOC_59/Y OR2X1_LOC_776/Y 0.04fF
C31756 AND2X1_LOC_59/Y OR2X1_LOC_756/B 0.21fF
C32260 AND2X1_LOC_59/Y OR2X1_LOC_719/A 0.01fF
C33079 AND2X1_LOC_59/Y OR2X1_LOC_87/B 0.03fF
C33290 AND2X1_LOC_59/Y OR2X1_LOC_333/A 0.43fF
C33474 OR2X1_LOC_100/Y AND2X1_LOC_59/Y 0.12fF
C33630 AND2X1_LOC_59/Y OR2X1_LOC_532/B 1.62fF
C33836 AND2X1_LOC_59/Y OR2X1_LOC_440/B 0.01fF
C34426 AND2X1_LOC_59/Y OR2X1_LOC_286/B 0.08fF
C34660 OR2X1_LOC_710/B AND2X1_LOC_59/Y 0.09fF
C35499 AND2X1_LOC_59/Y VDD 2.79fF
C35732 AND2X1_LOC_59/Y OR2X1_LOC_845/A 0.04fF
C36345 AND2X1_LOC_59/Y OR2X1_LOC_676/Y 0.50fF
C36444 AND2X1_LOC_59/Y OR2X1_LOC_462/B 0.02fF
C36935 AND2X1_LOC_59/Y OR2X1_LOC_602/B 0.01fF
C37651 AND2X1_LOC_59/Y OR2X1_LOC_840/A 0.01fF
C38063 AND2X1_LOC_59/Y OR2X1_LOC_216/A 0.13fF
C38294 AND2X1_LOC_59/Y OR2X1_LOC_750/Y 0.09fF
C38548 OR2X1_LOC_160/A AND2X1_LOC_59/Y 0.57fF
C38623 AND2X1_LOC_59/Y OR2X1_LOC_624/B 0.02fF
C38790 AND2X1_LOC_59/Y OR2X1_LOC_532/Y 0.18fF
C38844 AND2X1_LOC_59/Y OR2X1_LOC_266/A 0.16fF
C39109 AND2X1_LOC_59/Y AND2X1_LOC_108/a_8_24# 0.07fF
C39368 AND2X1_LOC_59/Y OR2X1_LOC_78/Y 0.03fF
C39514 AND2X1_LOC_59/Y AND2X1_LOC_491/a_8_24# 0.01fF
C39838 AND2X1_LOC_59/Y OR2X1_LOC_185/A 0.28fF
C40607 AND2X1_LOC_59/Y AND2X1_LOC_437/a_8_24# 0.03fF
C40959 AND2X1_LOC_59/Y OR2X1_LOC_294/Y 0.31fF
C41561 AND2X1_LOC_59/Y OR2X1_LOC_541/B 0.03fF
C42029 AND2X1_LOC_59/Y OR2X1_LOC_778/Y 0.09fF
C42250 AND2X1_LOC_91/B AND2X1_LOC_59/Y 2.41fF
C42753 AND2X1_LOC_59/Y OR2X1_LOC_719/B 0.02fF
C42880 AND2X1_LOC_59/Y AND2X1_LOC_56/B 0.73fF
C44271 AND2X1_LOC_59/Y OR2X1_LOC_68/Y 0.09fF
C44285 AND2X1_LOC_59/Y AND2X1_LOC_47/Y 0.42fF
C44588 AND2X1_LOC_59/Y OR2X1_LOC_506/A 0.04fF
C44822 AND2X1_LOC_59/Y OR2X1_LOC_180/B 0.29fF
C45030 AND2X1_LOC_59/Y AND2X1_LOC_95/Y 0.85fF
C45067 AND2X1_LOC_59/Y OR2X1_LOC_99/Y 0.05fF
C45242 AND2X1_LOC_59/Y OR2X1_LOC_788/B 0.27fF
C45461 AND2X1_LOC_59/Y OR2X1_LOC_664/a_8_216# 0.14fF
C46296 AND2X1_LOC_59/Y OR2X1_LOC_235/B 0.03fF
C46655 OR2X1_LOC_709/A AND2X1_LOC_59/Y 0.07fF
C46660 AND2X1_LOC_59/Y AND2X1_LOC_295/a_8_24# 0.20fF
C47499 AND2X1_LOC_59/Y OR2X1_LOC_771/B 0.05fF
C47521 AND2X1_LOC_59/Y OR2X1_LOC_776/A 0.07fF
C47931 AND2X1_LOC_59/Y OR2X1_LOC_593/B 0.03fF
C48049 AND2X1_LOC_59/Y AND2X1_LOC_41/a_8_24# 0.03fF
C48135 AND2X1_LOC_59/Y AND2X1_LOC_492/a_8_24# 0.01fF
C48440 AND2X1_LOC_59/Y AND2X1_LOC_44/Y 4.63fF
C49302 AND2X1_LOC_59/Y AND2X1_LOC_18/Y 1.23fF
C49376 AND2X1_LOC_59/Y OR2X1_LOC_473/a_8_216# 0.01fF
C50262 AND2X1_LOC_59/Y OR2X1_LOC_130/A 0.09fF
C51821 AND2X1_LOC_59/Y OR2X1_LOC_786/A 0.16fF
C52199 AND2X1_LOC_59/Y OR2X1_LOC_346/A 0.07fF
C52343 AND2X1_LOC_59/Y OR2X1_LOC_161/A 0.34fF
C52426 AND2X1_LOC_59/Y AND2X1_LOC_51/Y 0.21fF
C52736 AND2X1_LOC_59/Y OR2X1_LOC_640/A 0.16fF
C52779 AND2X1_LOC_59/Y OR2X1_LOC_541/a_8_216# 0.01fF
C52787 AND2X1_LOC_59/Y OR2X1_LOC_831/a_8_216# 0.01fF
C53139 AND2X1_LOC_59/Y AND2X1_LOC_41/A 0.54fF
C53224 AND2X1_LOC_59/Y OR2X1_LOC_631/B 0.02fF
C54621 AND2X1_LOC_59/Y AND2X1_LOC_31/Y 5.22fF
C54897 AND2X1_LOC_59/Y OR2X1_LOC_633/B 0.02fF
C55017 AND2X1_LOC_59/Y OR2X1_LOC_608/Y 0.06fF
C55450 AND2X1_LOC_59/Y AND2X1_LOC_72/B 0.02fF
C55520 AND2X1_LOC_59/Y AND2X1_LOC_36/Y 3.20fF
C55706 OR2X1_LOC_325/a_8_216# AND2X1_LOC_59/Y 0.04fF
C55781 AND2X1_LOC_59/Y OR2X1_LOC_346/B 0.37fF
C57899 AND2X1_LOC_59/Y VSS 1.20fF
C48 AND2X1_LOC_12/Y AND2X1_LOC_494/a_8_24# 0.02fF
C210 AND2X1_LOC_12/Y OR2X1_LOC_308/A 0.03fF
C441 AND2X1_LOC_12/Y OR2X1_LOC_557/A 0.11fF
C1309 AND2X1_LOC_12/Y OR2X1_LOC_269/B 0.28fF
C2064 AND2X1_LOC_12/Y OR2X1_LOC_678/Y 0.01fF
C2341 AND2X1_LOC_12/Y OR2X1_LOC_777/B 0.05fF
C2394 AND2X1_LOC_12/Y OR2X1_LOC_831/B 0.03fF
C2397 OR2X1_LOC_506/a_36_216# AND2X1_LOC_12/Y 0.02fF
C2651 AND2X1_LOC_12/Y AND2X1_LOC_13/a_8_24# 0.04fF
C2855 AND2X1_LOC_12/Y OR2X1_LOC_161/B 1.33fF
C2990 AND2X1_LOC_12/Y AND2X1_LOC_536/a_8_24# 0.01fF
C3007 AND2X1_LOC_12/Y OR2X1_LOC_846/a_8_216# 0.01fF
C3355 AND2X1_LOC_12/Y OR2X1_LOC_630/B 0.01fF
C3472 AND2X1_LOC_12/Y AND2X1_LOC_67/Y 0.03fF
C3859 AND2X1_LOC_12/Y OR2X1_LOC_644/B 0.03fF
C4206 AND2X1_LOC_12/Y AND2X1_LOC_230/a_8_24# 0.01fF
C4571 AND2X1_LOC_12/Y OR2X1_LOC_201/A 0.01fF
C4994 AND2X1_LOC_12/Y OR2X1_LOC_772/B 0.60fF
C5283 AND2X1_LOC_12/Y AND2X1_LOC_7/B 0.24fF
C6438 AND2X1_LOC_12/Y OR2X1_LOC_473/A 0.18fF
C6476 AND2X1_LOC_12/Y OR2X1_LOC_513/Y 0.01fF
C6797 AND2X1_LOC_12/Y OR2X1_LOC_287/B 0.05fF
C6834 AND2X1_LOC_12/Y OR2X1_LOC_76/A 0.03fF
C7100 AND2X1_LOC_12/Y OR2X1_LOC_160/B 5.76fF
C7935 AND2X1_LOC_12/Y OR2X1_LOC_318/A 0.01fF
C7967 AND2X1_LOC_12/Y OR2X1_LOC_151/A 0.92fF
C8462 AND2X1_LOC_12/Y OR2X1_LOC_287/A 0.03fF
C9262 AND2X1_LOC_12/Y OR2X1_LOC_631/A 0.01fF
C9454 AND2X1_LOC_12/Y OR2X1_LOC_285/B 0.01fF
C10036 AND2X1_LOC_12/Y OR2X1_LOC_334/a_8_216# 0.01fF
C10452 AND2X1_LOC_12/Y OR2X1_LOC_308/Y 0.01fF
C11040 AND2X1_LOC_12/Y OR2X1_LOC_664/Y 0.09fF
C11137 AND2X1_LOC_12/Y AND2X1_LOC_494/a_36_24# 0.01fF
C11312 AND2X1_LOC_12/Y OR2X1_LOC_61/A 0.02fF
C11384 AND2X1_LOC_12/Y AND2X1_LOC_24/a_8_24# 0.01fF
C11760 AND2X1_LOC_12/Y OR2X1_LOC_706/a_8_216# 0.01fF
C11769 AND2X1_LOC_12/Y OR2X1_LOC_390/A 0.03fF
C12591 AND2X1_LOC_229/a_8_24# AND2X1_LOC_12/Y 0.09fF
C13288 AND2X1_LOC_12/Y OR2X1_LOC_473/Y 0.05fF
C13454 OR2X1_LOC_188/Y AND2X1_LOC_12/Y 0.01fF
C13693 AND2X1_LOC_12/Y OR2X1_LOC_193/A 0.05fF
C13939 AND2X1_LOC_12/Y OR2X1_LOC_598/Y 0.02fF
C13942 AND2X1_LOC_12/Y AND2X1_LOC_131/a_8_24# 0.07fF
C14055 AND2X1_LOC_12/Y OR2X1_LOC_537/A 0.13fF
C14076 AND2X1_LOC_12/Y OR2X1_LOC_848/A 0.46fF
C14081 AND2X1_LOC_12/Y OR2X1_LOC_859/B 0.50fF
C14414 AND2X1_LOC_12/Y AND2X1_LOC_39/a_8_24# 0.01fF
C14654 AND2X1_LOC_12/Y OR2X1_LOC_558/A 0.33fF
C14914 AND2X1_LOC_12/Y OR2X1_LOC_810/A 0.17fF
C15166 OR2X1_LOC_715/B AND2X1_LOC_12/Y 0.03fF
C15514 AND2X1_LOC_12/Y OR2X1_LOC_338/B 0.01fF
C15695 AND2X1_LOC_12/Y OR2X1_LOC_793/A 0.11fF
C16124 AND2X1_LOC_12/Y OR2X1_LOC_687/Y 0.08fF
C16918 AND2X1_LOC_12/Y OR2X1_LOC_78/A 0.10fF
C16962 AND2X1_LOC_12/Y OR2X1_LOC_448/B 0.18fF
C17737 AND2X1_LOC_12/Y OR2X1_LOC_501/B 0.01fF
C17858 AND2X1_LOC_12/Y AND2X1_LOC_171/a_8_24# 0.01fF
C17978 AND2X1_LOC_12/Y OR2X1_LOC_318/B 0.03fF
C18116 OR2X1_LOC_231/B AND2X1_LOC_12/Y 0.05fF
C18126 OR2X1_LOC_121/Y AND2X1_LOC_12/Y 0.08fF
C18159 AND2X1_LOC_12/Y OR2X1_LOC_114/B 0.03fF
C18336 AND2X1_LOC_12/Y AND2X1_LOC_496/a_8_24# 0.01fF
C18753 AND2X1_LOC_12/Y AND2X1_LOC_495/a_8_24# 0.02fF
C19089 AND2X1_LOC_12/Y OR2X1_LOC_623/B 0.03fF
C19194 AND2X1_LOC_12/Y AND2X1_LOC_13/a_36_24# 0.01fF
C19230 AND2X1_LOC_12/Y OR2X1_LOC_544/A 0.05fF
C19566 AND2X1_LOC_12/Y OR2X1_LOC_848/B 0.28fF
C21096 AND2X1_LOC_12/Y OR2X1_LOC_338/A 0.01fF
C21125 OR2X1_LOC_186/Y AND2X1_LOC_12/Y 0.07fF
C21281 AND2X1_LOC_12/Y AND2X1_LOC_81/B 0.03fF
C21385 AND2X1_LOC_12/Y OR2X1_LOC_196/B 0.43fF
C21562 AND2X1_LOC_765/a_8_24# AND2X1_LOC_12/Y 0.02fF
C21757 AND2X1_LOC_12/Y OR2X1_LOC_574/A 0.04fF
C21763 AND2X1_LOC_12/Y OR2X1_LOC_33/A 0.01fF
C22119 AND2X1_LOC_12/Y AND2X1_LOC_16/a_8_24# 0.01fF
C22505 AND2X1_LOC_12/Y OR2X1_LOC_78/B 1.80fF
C22587 AND2X1_LOC_12/Y OR2X1_LOC_375/A 2.53fF
C22649 AND2X1_LOC_12/Y OR2X1_LOC_605/B 0.18fF
C22893 AND2X1_LOC_12/Y OR2X1_LOC_549/A 0.08fF
C23356 AND2X1_LOC_12/Y AND2X1_LOC_498/a_36_24# 0.01fF
C23368 AND2X1_LOC_12/Y OR2X1_LOC_499/B 0.04fF
C23443 AND2X1_LOC_12/Y OR2X1_LOC_391/B 0.76fF
C23496 AND2X1_LOC_12/Y OR2X1_LOC_846/A 0.05fF
C23584 AND2X1_LOC_12/Y OR2X1_LOC_348/B 0.12fF
C23705 AND2X1_LOC_12/Y AND2X1_LOC_65/A 0.03fF
C24116 AND2X1_LOC_12/Y AND2X1_LOC_603/a_8_24# 0.01fF
C24604 AND2X1_LOC_12/Y AND2X1_LOC_316/a_8_24# 0.01fF
C24896 OR2X1_LOC_335/A AND2X1_LOC_12/Y 0.31fF
C25155 AND2X1_LOC_12/Y AND2X1_LOC_27/a_8_24# 0.01fF
C25339 AND2X1_LOC_12/Y OR2X1_LOC_139/A 0.03fF
C25754 AND2X1_LOC_12/Y OR2X1_LOC_138/A 0.04fF
C26262 AND2X1_LOC_12/Y OR2X1_LOC_834/a_8_216# 0.02fF
C26760 AND2X1_LOC_12/Y OR2X1_LOC_87/A 0.39fF
C26838 AND2X1_LOC_12/Y OR2X1_LOC_706/B 0.01fF
C27536 AND2X1_LOC_12/Y OR2X1_LOC_61/B 0.03fF
C27562 AND2X1_LOC_12/Y OR2X1_LOC_194/B 0.01fF
C27788 AND2X1_LOC_12/Y OR2X1_LOC_349/B 0.22fF
C27848 AND2X1_LOC_12/Y OR2X1_LOC_97/A 0.06fF
C27979 AND2X1_LOC_12/Y OR2X1_LOC_475/B 0.03fF
C28030 AND2X1_LOC_12/Y AND2X1_LOC_282/a_8_24# 0.01fF
C28300 AND2X1_LOC_12/Y OR2X1_LOC_691/Y 0.02fF
C28319 AND2X1_LOC_12/Y OR2X1_LOC_713/A 0.03fF
C28413 AND2X1_LOC_12/Y OR2X1_LOC_629/Y 0.05fF
C28901 AND2X1_LOC_12/Y OR2X1_LOC_333/B 0.06fF
C28906 AND2X1_LOC_12/Y OR2X1_LOC_850/A 0.08fF
C29002 AND2X1_LOC_12/Y OR2X1_LOC_590/a_8_216# 0.01fF
C29283 AND2X1_LOC_12/Y OR2X1_LOC_154/A 0.62fF
C29336 AND2X1_LOC_12/Y OR2X1_LOC_778/A 0.01fF
C30070 AND2X1_LOC_12/Y OR2X1_LOC_634/A 0.02fF
C30214 AND2X1_LOC_12/Y OR2X1_LOC_335/B 0.03fF
C30617 AND2X1_LOC_12/Y OR2X1_LOC_34/B 0.03fF
C30741 AND2X1_LOC_12/Y OR2X1_LOC_590/Y 0.01fF
C30938 AND2X1_LOC_12/Y OR2X1_LOC_512/A 0.03fF
C31334 AND2X1_LOC_12/Y OR2X1_LOC_756/B 0.41fF
C31945 AND2X1_LOC_12/Y OR2X1_LOC_557/a_8_216# 0.01fF
C32065 OR2X1_LOC_614/Y AND2X1_LOC_12/Y 0.03fF
C32746 AND2X1_LOC_12/Y OR2X1_LOC_287/a_8_216# 0.01fF
C32871 AND2X1_LOC_12/Y OR2X1_LOC_333/A 0.01fF
C33177 AND2X1_LOC_12/Y OR2X1_LOC_532/B 9.84fF
C33445 AND2X1_LOC_12/Y OR2X1_LOC_391/A 0.19fF
C34022 AND2X1_LOC_12/Y OR2X1_LOC_286/B 0.01fF
C35079 AND2X1_LOC_12/Y VDD 1.32fF
C35164 AND2X1_LOC_12/Y AND2X1_LOC_755/a_8_24# 0.01fF
C35926 AND2X1_LOC_12/Y OR2X1_LOC_676/Y 0.08fF
C35948 AND2X1_LOC_12/Y OR2X1_LOC_834/A 0.63fF
C36226 AND2X1_LOC_12/Y AND2X1_LOC_591/a_8_24# 0.01fF
C37098 AND2X1_LOC_12/Y OR2X1_LOC_115/B 0.37fF
C37227 AND2X1_LOC_12/Y OR2X1_LOC_840/A 0.06fF
C37569 AND2X1_LOC_754/a_8_24# AND2X1_LOC_12/Y 0.02fF
C37647 AND2X1_LOC_12/Y OR2X1_LOC_216/A 0.07fF
C37727 AND2X1_LOC_12/Y AND2X1_LOC_385/a_8_24# 0.02fF
C37761 AND2X1_LOC_12/Y OR2X1_LOC_846/B 0.04fF
C37852 AND2X1_LOC_12/Y OR2X1_LOC_750/Y 0.11fF
C38098 AND2X1_LOC_12/Y OR2X1_LOC_160/A 0.21fF
C38346 AND2X1_LOC_12/Y OR2X1_LOC_130/Y 0.03fF
C38377 OR2X1_LOC_196/Y AND2X1_LOC_12/Y 0.03fF
C39023 AND2X1_LOC_12/Y OR2X1_LOC_285/A 0.01fF
C39420 AND2X1_LOC_12/Y OR2X1_LOC_185/A 0.07fF
C41337 AND2X1_LOC_12/Y AND2X1_LOC_238/a_8_24# 0.01fF
C41589 AND2X1_LOC_12/Y OR2X1_LOC_643/A 0.03fF
C41594 AND2X1_LOC_12/Y OR2X1_LOC_778/Y 0.22fF
C41824 AND2X1_LOC_12/Y AND2X1_LOC_91/B 0.13fF
C41952 AND2X1_LOC_12/Y OR2X1_LOC_308/a_8_216# 0.01fF
C42179 AND2X1_LOC_12/Y OR2X1_LOC_446/B 0.03fF
C42183 AND2X1_LOC_12/Y OR2X1_LOC_303/B 0.03fF
C42470 AND2X1_LOC_12/Y AND2X1_LOC_56/B 0.08fF
C43047 AND2X1_LOC_12/Y OR2X1_LOC_561/B 0.30fF
C43329 AND2X1_LOC_12/Y OR2X1_LOC_389/B 0.03fF
C43463 AND2X1_LOC_12/Y AND2X1_LOC_751/a_8_24# 0.18fF
C43842 AND2X1_LOC_12/Y OR2X1_LOC_68/Y 0.01fF
C43858 AND2X1_LOC_12/Y AND2X1_LOC_47/Y 0.19fF
C44151 AND2X1_LOC_12/Y OR2X1_LOC_506/A 0.02fF
C44547 AND2X1_LOC_12/Y OR2X1_LOC_391/a_8_216# 0.01fF
C44582 AND2X1_LOC_12/Y AND2X1_LOC_95/Y 14.07fF
C44969 AND2X1_LOC_12/Y OR2X1_LOC_706/A 0.06fF
C46089 AND2X1_LOC_12/Y OR2X1_LOC_779/B 0.05fF
C46211 OR2X1_LOC_709/A AND2X1_LOC_12/Y 0.01fF
C46303 AND2X1_LOC_12/Y OR2X1_LOC_703/A 0.06fF
C46358 AND2X1_LOC_12/Y OR2X1_LOC_791/B 0.01fF
C46681 AND2X1_LOC_12/Y OR2X1_LOC_362/A 0.05fF
C47036 AND2X1_LOC_12/Y OR2X1_LOC_771/B 0.03fF
C47063 AND2X1_LOC_12/Y OR2X1_LOC_776/A 0.03fF
C47201 AND2X1_LOC_12/Y OR2X1_LOC_678/a_8_216# 0.03fF
C47503 AND2X1_LOC_12/Y OR2X1_LOC_593/B 0.57fF
C47535 OR2X1_LOC_506/a_8_216# AND2X1_LOC_12/Y 0.03fF
C47688 AND2X1_LOC_12/Y AND2X1_LOC_492/a_8_24# 0.06fF
C47990 AND2X1_LOC_12/Y AND2X1_LOC_44/Y 0.20fF
C48613 AND2X1_LOC_12/Y AND2X1_LOC_69/Y 0.01fF
C48681 AND2X1_LOC_12/Y OR2X1_LOC_506/B 0.05fF
C48869 AND2X1_LOC_12/Y AND2X1_LOC_18/Y 0.81fF
C49138 AND2X1_LOC_12/Y OR2X1_LOC_789/A 0.07fF
C49276 AND2X1_LOC_12/Y OR2X1_LOC_307/A 0.01fF
C49519 AND2X1_LOC_12/Y AND2X1_LOC_69/a_8_24# 0.01fF
C49790 AND2X1_LOC_12/Y AND2X1_LOC_65/a_8_24# 0.01fF
C49847 AND2X1_LOC_12/Y OR2X1_LOC_130/A 0.07fF
C49982 AND2X1_LOC_12/Y AND2X1_LOC_39/Y 0.01fF
C50213 AND2X1_LOC_12/Y OR2X1_LOC_489/a_8_216# 0.01fF
C50288 AND2X1_LOC_12/Y OR2X1_LOC_449/B 0.03fF
C50773 AND2X1_LOC_12/Y OR2X1_LOC_383/Y 0.04fF
C51913 AND2X1_LOC_12/Y OR2X1_LOC_161/A 0.16fF
C51993 AND2X1_LOC_12/Y AND2X1_LOC_51/Y 2.24fF
C52713 AND2X1_LOC_12/Y AND2X1_LOC_41/A 13.38fF
C52804 AND2X1_LOC_12/Y OR2X1_LOC_631/B 0.03fF
C54185 AND2X1_LOC_12/Y AND2X1_LOC_31/Y 0.18fF
C54499 AND2X1_LOC_12/Y AND2X1_LOC_281/a_8_24# 0.01fF
C54835 AND2X1_LOC_12/Y AND2X1_LOC_305/a_8_24# 0.01fF
C54969 AND2X1_LOC_12/Y OR2X1_LOC_288/A 0.01fF
C55001 AND2X1_LOC_12/Y AND2X1_LOC_72/B 0.03fF
C55007 AND2X1_LOC_12/Y OR2X1_LOC_451/B 0.03fF
C55075 AND2X1_LOC_12/Y AND2X1_LOC_36/Y 1.98fF
C55091 AND2X1_LOC_12/Y OR2X1_LOC_333/a_8_216# 0.01fF
C55266 OR2X1_LOC_635/A AND2X1_LOC_12/Y 0.46fF
C55686 AND2X1_LOC_12/Y OR2X1_LOC_392/A 0.01fF
C58020 AND2X1_LOC_12/Y VSS -4.37fF
C318 AND2X1_LOC_95/Y OR2X1_LOC_634/A 0.18fF
C469 AND2X1_LOC_95/Y OR2X1_LOC_335/B 0.36fF
C913 AND2X1_LOC_95/Y OR2X1_LOC_34/B 0.01fF
C924 AND2X1_LOC_95/Y AND2X1_LOC_107/a_8_24# 0.01fF
C1222 AND2X1_LOC_95/Y OR2X1_LOC_464/A 0.03fF
C1627 OR2X1_LOC_756/B AND2X1_LOC_95/Y 2.12fF
C2014 AND2X1_LOC_95/Y OR2X1_LOC_370/a_8_216# 0.02fF
C2112 OR2X1_LOC_379/a_8_216# AND2X1_LOC_95/Y 0.02fF
C2433 OR2X1_LOC_653/B AND2X1_LOC_95/Y 0.01fF
C3089 AND2X1_LOC_95/Y OR2X1_LOC_287/a_8_216# 0.02fF
C3218 AND2X1_LOC_95/Y OR2X1_LOC_333/A 0.01fF
C3290 AND2X1_LOC_95/Y OR2X1_LOC_113/B 0.23fF
C3399 AND2X1_LOC_95/Y OR2X1_LOC_286/Y -0.00fF
C3505 AND2X1_LOC_95/Y OR2X1_LOC_532/B 3.08fF
C4094 AND2X1_LOC_95/Y OR2X1_LOC_729/a_8_216# 0.01fF
C4141 OR2X1_LOC_114/a_8_216# AND2X1_LOC_95/Y 0.01fF
C4310 AND2X1_LOC_95/Y OR2X1_LOC_286/B 0.36fF
C4704 AND2X1_LOC_95/Y OR2X1_LOC_472/B 0.02fF
C4792 AND2X1_LOC_95/Y OR2X1_LOC_552/A 0.03fF
C4973 AND2X1_LOC_95/Y OR2X1_LOC_798/Y 0.09fF
C4975 AND2X1_LOC_95/Y AND2X1_LOC_52/a_8_24# 0.08fF
C5328 VDD AND2X1_LOC_95/Y 2.04fF
C6093 AND2X1_LOC_95/Y OR2X1_LOC_523/A 0.01fF
C6290 AND2X1_LOC_95/Y OR2X1_LOC_462/B 0.72fF
C7460 AND2X1_LOC_95/Y OR2X1_LOC_115/B 0.06fF
C7535 AND2X1_LOC_95/Y OR2X1_LOC_370/a_36_216# 0.02fF
C7583 AND2X1_LOC_95/Y OR2X1_LOC_840/A 0.01fF
C7947 AND2X1_LOC_594/a_36_24# AND2X1_LOC_95/Y 0.01fF
C8172 AND2X1_LOC_95/Y AND2X1_LOC_134/a_8_24# 0.05fF
C8536 OR2X1_LOC_160/A AND2X1_LOC_95/Y 0.22fF
C8600 AND2X1_LOC_95/Y OR2X1_LOC_624/B 0.04fF
C8732 AND2X1_LOC_95/Y OR2X1_LOC_532/Y 0.02fF
C8891 OR2X1_LOC_325/A AND2X1_LOC_95/Y 0.16fF
C9037 AND2X1_LOC_95/Y AND2X1_LOC_108/a_8_24# 0.01fF
C9389 AND2X1_LOC_95/Y OR2X1_LOC_285/A 0.27fF
C9784 AND2X1_LOC_95/Y OR2X1_LOC_185/A 0.12fF
C9856 AND2X1_LOC_95/Y OR2X1_LOC_435/Y 0.13fF
C9903 AND2X1_LOC_95/Y AND2X1_LOC_431/a_8_24# 0.01fF
C10581 AND2X1_LOC_95/Y OR2X1_LOC_802/a_8_216# 0.02fF
C10900 AND2X1_LOC_95/Y OR2X1_LOC_294/Y 0.03fF
C11049 OR2X1_LOC_114/Y AND2X1_LOC_95/Y 0.01fF
C11133 AND2X1_LOC_95/Y OR2X1_LOC_286/a_8_216# 0.01fF
C11848 AND2X1_LOC_95/Y OR2X1_LOC_436/B 0.01fF
C11912 AND2X1_LOC_95/Y OR2X1_LOC_643/A 0.03fF
C11918 AND2X1_LOC_95/Y OR2X1_LOC_778/Y 0.03fF
C11966 AND2X1_LOC_95/Y OR2X1_LOC_113/A 0.01fF
C12138 AND2X1_LOC_91/B AND2X1_LOC_95/Y 0.21fF
C12503 AND2X1_LOC_95/Y OR2X1_LOC_446/B 0.06fF
C12508 AND2X1_LOC_95/Y OR2X1_LOC_303/B 0.03fF
C12760 AND2X1_LOC_95/Y AND2X1_LOC_56/B 9.31fF
C13114 AND2X1_LOC_95/Y OR2X1_LOC_787/B 0.01fF
C14146 AND2X1_LOC_95/Y OR2X1_LOC_287/a_36_216# 0.01fF
C14153 AND2X1_LOC_95/Y AND2X1_LOC_47/Y 0.21fF
C14320 AND2X1_LOC_521/a_8_24# AND2X1_LOC_95/Y 0.01fF
C14442 AND2X1_LOC_95/Y OR2X1_LOC_506/A 0.03fF
C14584 AND2X1_LOC_95/Y AND2X1_LOC_420/a_8_24# 0.03fF
C15072 AND2X1_LOC_95/Y OR2X1_LOC_788/B 0.01fF
C15366 AND2X1_LOC_95/Y OR2X1_LOC_434/A 0.01fF
C16049 AND2X1_LOC_95/Y OR2X1_LOC_235/B 0.03fF
C16474 AND2X1_LOC_95/Y OR2X1_LOC_703/A 1.86fF
C16526 OR2X1_LOC_791/B AND2X1_LOC_95/Y 0.03fF
C16863 AND2X1_LOC_95/Y OR2X1_LOC_362/A 0.49fF
C17058 AND2X1_LOC_95/Y AND2X1_LOC_680/a_8_24# 0.01fF
C17184 AND2X1_LOC_95/Y OR2X1_LOC_771/B 0.03fF
C18100 AND2X1_LOC_95/Y AND2X1_LOC_44/Y 2.93fF
C18374 AND2X1_LOC_95/Y OR2X1_LOC_720/B 0.02fF
C19005 AND2X1_LOC_95/Y AND2X1_LOC_18/Y 0.21fF
C19849 OR2X1_LOC_523/B AND2X1_LOC_95/Y 0.01fF
C19997 AND2X1_LOC_95/Y OR2X1_LOC_130/A 0.15fF
C20390 AND2X1_LOC_95/Y AND2X1_LOC_487/a_8_24# 0.11fF
C20393 AND2X1_LOC_95/Y OR2X1_LOC_128/A 0.02fF
C20431 AND2X1_LOC_95/Y OR2X1_LOC_449/B 0.03fF
C21662 AND2X1_LOC_95/Y OR2X1_LOC_802/a_36_216# 0.02fF
C21669 AND2X1_LOC_95/Y AND2X1_LOC_52/a_36_24# 0.01fF
C22127 AND2X1_LOC_95/Y OR2X1_LOC_161/A 0.72fF
C22209 AND2X1_LOC_95/Y AND2X1_LOC_51/Y 0.82fF
C22752 AND2X1_LOC_95/Y AND2X1_LOC_52/Y 0.03fF
C22941 AND2X1_LOC_95/Y AND2X1_LOC_41/A 0.10fF
C23031 AND2X1_LOC_95/Y OR2X1_LOC_631/B 0.16fF
C23638 AND2X1_LOC_57/Y AND2X1_LOC_95/Y 0.04fF
C24408 AND2X1_LOC_95/Y AND2X1_LOC_31/Y 0.11fF
C25168 AND2X1_LOC_95/Y OR2X1_LOC_288/A 0.02fF
C25209 AND2X1_LOC_95/Y AND2X1_LOC_72/B 1.48fF
C25284 AND2X1_LOC_95/Y AND2X1_LOC_36/Y 0.50fF
C25301 AND2X1_LOC_95/Y OR2X1_LOC_333/a_8_216# 0.03fF
C25435 OR2X1_LOC_325/a_8_216# AND2X1_LOC_95/Y 0.02fF
C25506 AND2X1_LOC_95/Y OR2X1_LOC_346/B 0.15fF
C25876 AND2X1_LOC_95/Y OR2X1_LOC_128/B 0.04fF
C26161 AND2X1_LOC_522/a_8_24# AND2X1_LOC_95/Y 0.01fF
C26201 AND2X1_LOC_95/Y OR2X1_LOC_730/A 0.01fF
C26785 AND2X1_LOC_95/Y OR2X1_LOC_557/A 0.02fF
C27101 OR2X1_LOC_768/A AND2X1_LOC_95/Y 0.10fF
C27604 AND2X1_LOC_95/Y OR2X1_LOC_269/B 0.48fF
C28007 AND2X1_LOC_95/Y OR2X1_LOC_347/B 0.20fF
C28013 AND2X1_LOC_95/Y OR2X1_LOC_539/Y 0.68fF
C28347 AND2X1_LOC_95/Y AND2X1_LOC_184/a_8_24# 0.04fF
C28429 AND2X1_LOC_533/a_8_24# AND2X1_LOC_95/Y 0.04fF
C28618 AND2X1_LOC_95/Y OR2X1_LOC_777/B 0.15fF
C28705 AND2X1_LOC_95/Y OR2X1_LOC_344/A 0.03fF
C29071 OR2X1_LOC_198/a_8_216# AND2X1_LOC_95/Y 0.02fF
C29118 AND2X1_LOC_95/Y OR2X1_LOC_161/B 3.67fF
C29681 AND2X1_LOC_95/Y AND2X1_LOC_132/a_8_24# 0.01fF
C31640 AND2X1_LOC_95/Y AND2X1_LOC_7/B 0.69fF
C31752 OR2X1_LOC_319/B AND2X1_LOC_95/Y 0.13fF
C31828 AND2X1_LOC_95/Y OR2X1_LOC_296/Y 0.03fF
C31850 AND2X1_LOC_95/Y OR2X1_LOC_436/a_8_216# 0.01fF
C32108 AND2X1_LOC_95/Y AND2X1_LOC_103/a_8_24# 0.17fF
C33089 AND2X1_LOC_95/Y OR2X1_LOC_287/B 0.11fF
C33182 AND2X1_LOC_95/Y OR2X1_LOC_436/Y 0.04fF
C33381 OR2X1_LOC_160/B AND2X1_LOC_95/Y 5.91fF
C33508 AND2X1_LOC_95/Y OR2X1_LOC_553/A 0.07fF
C34195 AND2X1_LOC_95/Y OR2X1_LOC_151/A 3.86fF
C34548 OR2X1_LOC_198/a_36_216# AND2X1_LOC_95/Y 0.01fF
C34659 AND2X1_LOC_95/Y OR2X1_LOC_287/A 0.03fF
C34676 AND2X1_LOC_95/Y OR2X1_LOC_174/A 0.01fF
C34688 AND2X1_LOC_95/Y OR2X1_LOC_435/a_8_216# 0.01fF
C35162 AND2X1_LOC_95/Y OR2X1_LOC_137/B 0.26fF
C35189 AND2X1_LOC_95/Y AND2X1_LOC_252/a_8_24# 0.04fF
C35388 AND2X1_LOC_95/Y OR2X1_LOC_415/Y 0.89fF
C35663 AND2X1_LOC_95/Y OR2X1_LOC_285/B 0.26fF
C36162 AND2X1_LOC_95/Y AND2X1_LOC_497/a_8_24# 0.01fF
C36257 AND2X1_LOC_95/Y OR2X1_LOC_334/a_8_216# 0.01fF
C36791 AND2X1_LOC_95/Y AND2X1_LOC_125/a_8_24# 0.01fF
C37268 AND2X1_LOC_95/Y OR2X1_LOC_664/Y 0.03fF
C37479 AND2X1_LOC_95/Y OR2X1_LOC_342/a_8_216# 0.01fF
C37607 AND2X1_LOC_95/Y AND2X1_LOC_24/a_8_24# 0.01fF
C37966 AND2X1_LOC_95/Y OR2X1_LOC_390/A 0.03fF
C38536 AND2X1_LOC_95/Y OR2X1_LOC_668/Y 0.01fF
C39337 AND2X1_LOC_95/Y AND2X1_LOC_94/Y 0.05fF
C39493 AND2X1_LOC_95/Y OR2X1_LOC_473/Y 0.15fF
C39577 AND2X1_LOC_95/Y OR2X1_LOC_241/B 0.09fF
C39680 OR2X1_LOC_188/Y AND2X1_LOC_95/Y 0.05fF
C39730 AND2X1_LOC_95/Y OR2X1_LOC_325/B 0.07fF
C39772 AND2X1_LOC_95/Y AND2X1_LOC_189/a_8_24# 0.02fF
C39788 AND2X1_LOC_95/Y OR2X1_LOC_285/a_8_216# 0.01fF
C39834 AND2X1_LOC_95/Y OR2X1_LOC_405/Y 0.01fF
C40014 AND2X1_LOC_95/Y OR2X1_LOC_339/A 0.03fF
C40084 AND2X1_LOC_95/Y AND2X1_LOC_438/a_8_24# 0.03fF
C40103 AND2X1_LOC_95/Y OR2X1_LOC_598/Y 0.03fF
C40147 OR2X1_LOC_335/Y AND2X1_LOC_95/Y 0.14fF
C40348 AND2X1_LOC_95/Y AND2X1_LOC_826/a_8_24# -0.01fF
C40544 AND2X1_LOC_95/Y OR2X1_LOC_356/A 0.08fF
C40910 AND2X1_LOC_95/Y AND2X1_LOC_416/a_8_24# 0.17fF
C41142 AND2X1_LOC_95/Y OR2X1_LOC_810/A 0.08fF
C41162 AND2X1_LOC_589/a_8_24# AND2X1_LOC_95/Y 0.03fF
C41424 OR2X1_LOC_715/B AND2X1_LOC_95/Y 0.03fF
C41427 AND2X1_LOC_95/Y AND2X1_LOC_626/a_8_24# 0.10fF
C41432 AND2X1_LOC_95/Y OR2X1_LOC_543/A 0.48fF
C41805 AND2X1_LOC_95/Y OR2X1_LOC_338/B 0.01fF
C42370 AND2X1_LOC_95/Y OR2X1_LOC_837/Y 0.01fF
C42734 AND2X1_LOC_95/Y OR2X1_LOC_535/A 0.01fF
C43202 AND2X1_LOC_95/Y OR2X1_LOC_78/A 6.21fF
C44084 OR2X1_LOC_501/B AND2X1_LOC_95/Y 0.03fF
C44119 AND2X1_LOC_95/Y OR2X1_LOC_147/B 0.03fF
C44162 AND2X1_LOC_95/Y AND2X1_LOC_669/a_8_24# 0.01fF
C44197 AND2X1_LOC_171/a_8_24# AND2X1_LOC_95/Y 0.01fF
C44323 AND2X1_LOC_95/Y OR2X1_LOC_318/B 0.08fF
C44470 OR2X1_LOC_114/B AND2X1_LOC_95/Y 0.08fF
C44515 AND2X1_LOC_95/Y OR2X1_LOC_538/A 0.03fF
C44919 AND2X1_LOC_95/Y AND2X1_LOC_184/a_36_24# 0.01fF
C45239 AND2X1_LOC_95/Y OR2X1_LOC_342/B 0.26fF
C45414 AND2X1_LOC_95/Y OR2X1_LOC_623/B 1.38fF
C45570 AND2X1_LOC_95/Y OR2X1_LOC_544/A 0.03fF
C45827 AND2X1_LOC_95/Y OR2X1_LOC_434/a_8_216# 0.01fF
C45868 AND2X1_LOC_95/Y OR2X1_LOC_833/B 0.02fF
C45893 AND2X1_LOC_95/Y OR2X1_LOC_254/B 0.07fF
C46395 AND2X1_LOC_95/Y AND2X1_LOC_252/a_36_24# 0.01fF
C47538 AND2X1_LOC_95/Y OR2X1_LOC_338/A 0.01fF
C47569 OR2X1_LOC_186/Y AND2X1_LOC_95/Y 0.28fF
C47836 AND2X1_LOC_95/Y OR2X1_LOC_112/B 0.02fF
C48144 AND2X1_LOC_95/Y OR2X1_LOC_39/A 0.03fF
C48199 AND2X1_LOC_95/Y OR2X1_LOC_574/A 0.03fF
C48201 AND2X1_LOC_95/Y OR2X1_LOC_33/A 0.01fF
C48422 AND2X1_LOC_95/Y AND2X1_LOC_627/a_8_24# 0.02fF
C48760 AND2X1_LOC_95/Y OR2X1_LOC_539/B 0.02fF
C48889 AND2X1_LOC_95/Y OR2X1_LOC_78/B 0.10fF
C48971 AND2X1_LOC_95/Y OR2X1_LOC_375/A 0.22fF
C49244 AND2X1_LOC_95/Y OR2X1_LOC_549/A 0.08fF
C49301 OR2X1_LOC_325/Y AND2X1_LOC_95/Y 0.04fF
C49998 AND2X1_LOC_95/Y OR2X1_LOC_543/a_8_216# 0.01fF
C50518 AND2X1_LOC_95/Y AND2X1_LOC_603/a_8_24# 0.03fF
C50769 AND2X1_LOC_95/Y OR2X1_LOC_285/Y 0.01fF
C51096 AND2X1_LOC_95/Y OR2X1_LOC_673/Y 0.03fF
C51566 AND2X1_LOC_95/Y AND2X1_LOC_27/a_8_24# 0.01fF
C51768 OR2X1_LOC_139/A AND2X1_LOC_95/Y 0.06fF
C52092 AND2X1_LOC_95/Y OR2X1_LOC_728/A 0.01fF
C53063 AND2X1_LOC_594/a_8_24# AND2X1_LOC_95/Y 0.02fF
C53160 AND2X1_LOC_95/Y OR2X1_LOC_668/a_8_216# 0.01fF
C53188 OR2X1_LOC_703/B AND2X1_LOC_95/Y 0.03fF
C53201 AND2X1_LOC_95/Y OR2X1_LOC_87/A 0.18fF
C53410 AND2X1_LOC_95/Y OR2X1_LOC_844/B 0.01fF
C54209 AND2X1_LOC_95/Y OR2X1_LOC_349/B 0.01fF
C54267 OR2X1_LOC_97/A AND2X1_LOC_95/Y 0.06fF
C54394 AND2X1_LOC_95/Y OR2X1_LOC_475/B 0.03fF
C54704 AND2X1_LOC_95/Y OR2X1_LOC_691/Y 0.09fF
C55271 AND2X1_LOC_95/Y AND2X1_LOC_74/a_8_24# 0.06fF
C55313 AND2X1_LOC_95/Y OR2X1_LOC_720/A 0.01fF
C55352 OR2X1_LOC_333/B AND2X1_LOC_95/Y 0.05fF
C55744 OR2X1_LOC_154/A AND2X1_LOC_95/Y 0.18fF
C56086 AND2X1_LOC_95/Y AND2X1_LOC_96/a_8_24# 0.11fF
C56794 AND2X1_LOC_95/Y VSS -4.24fF
C9729 OR2X1_LOC_596/Y VDD 0.16fF
C10556 OR2X1_LOC_596/Y OR2X1_LOC_676/Y 0.04fF
C17028 OR2X1_LOC_596/Y AND2X1_LOC_56/B 0.01fF
C27158 OR2X1_LOC_596/Y AND2X1_LOC_41/A 0.12fF
C28885 OR2X1_LOC_596/Y AND2X1_LOC_597/a_8_24# 0.23fF
C33369 OR2X1_LOC_596/Y OR2X1_LOC_161/B 0.02fF
C57951 OR2X1_LOC_596/Y VSS 0.07fF
C1037 OR2X1_LOC_448/B OR2X1_LOC_777/B 0.04fF
C10135 OR2X1_LOC_448/A OR2X1_LOC_448/B 0.26fF
C15585 OR2X1_LOC_448/B OR2X1_LOC_78/A 0.11fF
C21210 OR2X1_LOC_448/B OR2X1_LOC_448/a_8_216# 0.07fF
C21240 OR2X1_LOC_448/B OR2X1_LOC_375/A 0.01fF
C25093 OR2X1_LOC_448/B AND2X1_LOC_697/a_8_24# 0.01fF
C27000 OR2X1_LOC_448/B OR2X1_LOC_713/A 0.01fF
C33803 VDD OR2X1_LOC_448/B 0.21fF
C36050 OR2X1_LOC_448/B AND2X1_LOC_697/a_36_24# 0.01fF
C40225 OR2X1_LOC_448/B OR2X1_LOC_778/Y 0.05fF
C44743 OR2X1_LOC_448/B OR2X1_LOC_779/B 0.02fF
C46619 OR2X1_LOC_448/B AND2X1_LOC_44/Y 0.10fF
C50633 OR2X1_LOC_448/B OR2X1_LOC_161/A 0.01fF
C52934 OR2X1_LOC_448/B AND2X1_LOC_31/Y 0.03fF
C56185 OR2X1_LOC_448/B OR2X1_LOC_269/B 0.02fF
C57120 OR2X1_LOC_448/B VSS 0.21fF
C8437 OR2X1_LOC_355/B OR2X1_LOC_355/A 0.04fF
C9938 OR2X1_LOC_355/B OR2X1_LOC_532/B 0.01fF
C11847 VDD OR2X1_LOC_355/B -0.00fF
C14918 OR2X1_LOC_160/A OR2X1_LOC_355/B 0.06fF
C19185 AND2X1_LOC_56/B OR2X1_LOC_355/B 0.03fF
C28551 OR2X1_LOC_355/B AND2X1_LOC_51/Y 0.23fF
C30445 OR2X1_LOC_355/B OR2X1_LOC_355/a_8_216# 0.05fF
C40603 OR2X1_LOC_151/A OR2X1_LOC_355/B 0.08fF
C47184 OR2X1_LOC_355/B OR2X1_LOC_356/A 0.81fF
C53936 OR2X1_LOC_186/Y OR2X1_LOC_355/B 0.01fF
C57251 OR2X1_LOC_355/B VSS 0.11fF
C7 OR2X1_LOC_667/a_8_216# OR2X1_LOC_26/Y 0.01fF
C888 OR2X1_LOC_26/Y OR2X1_LOC_588/Y 0.04fF
C1744 OR2X1_LOC_26/Y AND2X1_LOC_266/Y 0.03fF
C2174 OR2X1_LOC_26/Y OR2X1_LOC_511/Y 0.34fF
C2574 OR2X1_LOC_265/a_8_216# OR2X1_LOC_26/Y 0.01fF
C2623 OR2X1_LOC_26/Y OR2X1_LOC_237/Y 0.04fF
C2965 OR2X1_LOC_26/Y AND2X1_LOC_637/a_36_24# -0.00fF
C2967 OR2X1_LOC_91/A OR2X1_LOC_26/Y 0.32fF
C3024 OR2X1_LOC_823/a_8_216# OR2X1_LOC_26/Y 0.01fF
C3067 OR2X1_LOC_669/Y OR2X1_LOC_26/Y 0.21fF
C3442 OR2X1_LOC_32/B OR2X1_LOC_26/Y 0.34fF
C3490 OR2X1_LOC_26/Y OR2X1_LOC_371/Y 0.07fF
C3905 AND2X1_LOC_673/a_8_24# OR2X1_LOC_26/Y 0.01fF
C3921 OR2X1_LOC_26/Y OR2X1_LOC_74/A 0.27fF
C4260 OR2X1_LOC_26/Y AND2X1_LOC_287/Y 0.01fF
C4655 OR2X1_LOC_26/Y AND2X1_LOC_287/a_8_24# 0.02fF
C5301 OR2X1_LOC_134/Y OR2X1_LOC_26/Y 0.01fF
C5702 OR2X1_LOC_516/a_36_216# OR2X1_LOC_26/Y 0.02fF
C5733 OR2X1_LOC_106/Y OR2X1_LOC_26/Y 0.03fF
C6307 AND2X1_LOC_99/A OR2X1_LOC_26/Y 0.02fF
C6361 OR2X1_LOC_26/Y AND2X1_LOC_637/Y 0.01fF
C6488 OR2X1_LOC_26/Y OR2X1_LOC_72/Y 0.01fF
C6809 OR2X1_LOC_670/a_8_216# OR2X1_LOC_26/Y 0.01fF
C7109 AND2X1_LOC_362/B OR2X1_LOC_26/Y 0.16fF
C7225 OR2X1_LOC_26/Y OR2X1_LOC_595/a_8_216# 0.07fF
C7300 OR2X1_LOC_431/a_8_216# OR2X1_LOC_26/Y 0.14fF
C7576 OR2X1_LOC_58/Y OR2X1_LOC_26/Y 0.03fF
C7689 OR2X1_LOC_81/Y OR2X1_LOC_26/Y 0.05fF
C7710 OR2X1_LOC_485/A OR2X1_LOC_26/Y 0.74fF
C8241 OR2X1_LOC_26/Y OR2X1_LOC_238/a_8_216# 0.01fF
C8332 OR2X1_LOC_26/Y OR2X1_LOC_385/a_8_216# 0.03fF
C9374 OR2X1_LOC_290/a_8_216# OR2X1_LOC_26/Y 0.07fF
C9714 OR2X1_LOC_26/Y OR2X1_LOC_13/Y 0.02fF
C9813 OR2X1_LOC_165/a_36_216# OR2X1_LOC_26/Y 0.02fF
C11287 OR2X1_LOC_516/Y OR2X1_LOC_26/Y 0.03fF
C12407 OR2X1_LOC_131/Y OR2X1_LOC_26/Y 0.03fF
C12691 VDD OR2X1_LOC_26/Y 1.48fF
C12734 OR2X1_LOC_677/Y OR2X1_LOC_26/Y 0.02fF
C12813 OR2X1_LOC_26/Y AND2X1_LOC_267/a_8_24# 0.01fF
C12824 OR2X1_LOC_251/Y OR2X1_LOC_26/Y 0.01fF
C12900 OR2X1_LOC_256/A OR2X1_LOC_26/Y 0.03fF
C12936 OR2X1_LOC_26/Y OR2X1_LOC_67/Y 0.06fF
C13257 OR2X1_LOC_26/Y AND2X1_LOC_834/a_8_24# 0.02fF
C13269 OR2X1_LOC_26/Y OR2X1_LOC_248/Y 0.18fF
C13751 OR2X1_LOC_26/Y OR2X1_LOC_238/a_36_216# 0.02fF
C14072 OR2X1_LOC_26/Y OR2X1_LOC_427/A 0.63fF
C14083 OR2X1_LOC_823/Y OR2X1_LOC_26/Y 0.02fF
C14568 OR2X1_LOC_26/Y OR2X1_LOC_416/Y 0.04fF
C15571 OR2X1_LOC_45/B OR2X1_LOC_26/Y 0.22fF
C15714 OR2X1_LOC_26/Y OR2X1_LOC_767/a_8_216# 0.14fF
C16034 OR2X1_LOC_158/A OR2X1_LOC_26/Y 0.42fF
C16101 OR2X1_LOC_103/Y OR2X1_LOC_26/Y 0.10fF
C16548 OR2X1_LOC_26/Y OR2X1_LOC_586/Y 0.04fF
C16639 OR2X1_LOC_304/Y OR2X1_LOC_26/Y 0.02fF
C16949 OR2X1_LOC_132/a_8_216# OR2X1_LOC_26/Y 0.01fF
C17984 OR2X1_LOC_26/Y OR2X1_LOC_41/a_8_216# 0.01fF
C18183 AND2X1_LOC_541/Y OR2X1_LOC_26/Y 0.01fF
C18306 OR2X1_LOC_316/Y OR2X1_LOC_26/Y 0.04fF
C18385 OR2X1_LOC_431/Y OR2X1_LOC_26/Y 0.18fF
C18392 AND2X1_LOC_101/a_8_24# OR2X1_LOC_26/Y 0.06fF
C18667 OR2X1_LOC_744/A OR2X1_LOC_26/Y 3.43fF
C18772 OR2X1_LOC_26/Y AND2X1_LOC_840/B 0.05fF
C19004 OR2X1_LOC_26/Y AND2X1_LOC_464/A 0.03fF
C19354 OR2X1_LOC_26/Y OR2X1_LOC_385/a_36_216# 0.03fF
C19956 OR2X1_LOC_26/Y OR2X1_LOC_56/A 0.07fF
C20404 OR2X1_LOC_290/Y OR2X1_LOC_26/Y 0.01fF
C20450 OR2X1_LOC_91/Y OR2X1_LOC_26/Y 0.16fF
C20518 OR2X1_LOC_291/Y OR2X1_LOC_26/Y 0.03fF
C20782 AND2X1_LOC_330/a_8_24# OR2X1_LOC_26/Y 0.03fF
C20924 AND2X1_LOC_342/a_36_24# OR2X1_LOC_26/Y 0.01fF
C21274 OR2X1_LOC_667/Y OR2X1_LOC_26/Y 0.01fF
C21841 OR2X1_LOC_26/Y OR2X1_LOC_71/Y 0.05fF
C22252 OR2X1_LOC_26/Y OR2X1_LOC_246/A 0.12fF
C22283 OR2X1_LOC_26/Y OR2X1_LOC_409/B 0.02fF
C22596 OR2X1_LOC_525/Y OR2X1_LOC_26/Y 0.27fF
C23028 OR2X1_LOC_109/a_8_216# OR2X1_LOC_26/Y 0.01fF
C23564 OR2X1_LOC_26/Y AND2X1_LOC_721/A 0.04fF
C23892 OR2X1_LOC_26/Y AND2X1_LOC_361/A 0.21fF
C24298 OR2X1_LOC_26/Y AND2X1_LOC_834/a_36_24# 0.01fF
C24313 OR2X1_LOC_83/Y OR2X1_LOC_26/Y 0.07fF
C24522 AND2X1_LOC_787/A OR2X1_LOC_26/Y 0.03fF
C25099 OR2X1_LOC_26/Y OR2X1_LOC_65/B 0.09fF
C25409 OR2X1_LOC_600/A OR2X1_LOC_26/Y 0.77fF
C25504 OR2X1_LOC_26/Y OR2X1_LOC_619/Y 0.13fF
C25835 OR2X1_LOC_26/Y AND2X1_LOC_286/a_8_24# 0.01fF
C25933 OR2X1_LOC_669/A OR2X1_LOC_26/Y 0.05fF
C25997 AND2X1_LOC_334/a_8_24# OR2X1_LOC_26/Y 0.02fF
C26058 OR2X1_LOC_26/Y OR2X1_LOC_289/Y 0.03fF
C26264 OR2X1_LOC_331/A OR2X1_LOC_26/Y 0.04fF
C26491 OR2X1_LOC_26/Y OR2X1_LOC_406/A 0.01fF
C26779 OR2X1_LOC_26/Y OR2X1_LOC_69/A 0.03fF
C27188 AND2X1_LOC_113/a_8_24# OR2X1_LOC_26/Y 0.03fF
C27657 OR2X1_LOC_312/Y OR2X1_LOC_26/Y 0.03fF
C27807 OR2X1_LOC_26/Y OR2X1_LOC_13/B 1.07fF
C28335 OR2X1_LOC_26/Y OR2X1_LOC_428/A 0.90fF
C28351 OR2X1_LOC_26/Y OR2X1_LOC_595/A 0.47fF
C28877 OR2X1_LOC_516/A OR2X1_LOC_26/Y 0.03fF
C28912 AND2X1_LOC_105/a_8_24# OR2X1_LOC_26/Y 0.03fF
C29349 OR2X1_LOC_26/Y OR2X1_LOC_89/A 1.42fF
C29541 OR2X1_LOC_26/Y AND2X1_LOC_590/a_8_24# 0.03fF
C29995 OR2X1_LOC_26/Y AND2X1_LOC_287/B 0.02fF
C30140 OR2X1_LOC_45/Y OR2X1_LOC_26/Y 0.02fF
C30154 AND2X1_LOC_843/a_8_24# OR2X1_LOC_26/Y 0.02fF
C30176 OR2X1_LOC_26/Y OR2X1_LOC_824/Y 0.44fF
C30232 AND2X1_LOC_727/A OR2X1_LOC_26/Y 0.03fF
C30256 OR2X1_LOC_26/Y OR2X1_LOC_95/Y 2.31fF
C31006 OR2X1_LOC_26/Y AND2X1_LOC_621/Y 0.03fF
C31023 OR2X1_LOC_26/Y AND2X1_LOC_668/a_8_24# 0.04fF
C31463 OR2X1_LOC_70/Y OR2X1_LOC_26/Y 2.69fF
C32962 OR2X1_LOC_26/Y OR2X1_LOC_16/A 1.25fF
C32996 OR2X1_LOC_108/Y OR2X1_LOC_26/Y 0.07fF
C33070 AND2X1_LOC_168/Y OR2X1_LOC_26/Y 0.06fF
C33467 OR2X1_LOC_132/Y OR2X1_LOC_26/Y 0.04fF
C33880 AND2X1_LOC_334/Y OR2X1_LOC_26/Y 0.01fF
C33948 OR2X1_LOC_109/Y OR2X1_LOC_26/Y 0.08fF
C33980 OR2X1_LOC_262/a_8_216# OR2X1_LOC_26/Y 0.01fF
C34013 OR2X1_LOC_26/Y AND2X1_LOC_729/B 0.02fF
C34448 AND2X1_LOC_227/Y OR2X1_LOC_26/Y 0.09fF
C34476 OR2X1_LOC_26/Y OR2X1_LOC_813/Y 0.07fF
C34481 OR2X1_LOC_26/Y OR2X1_LOC_41/Y 0.13fF
C34725 OR2X1_LOC_107/Y OR2X1_LOC_26/Y 0.02fF
C34834 OR2X1_LOC_599/A OR2X1_LOC_26/Y 0.09fF
C35100 OR2X1_LOC_40/Y OR2X1_LOC_26/Y 6.02fF
C35179 AND2X1_LOC_843/Y OR2X1_LOC_26/Y 0.01fF
C35234 OR2X1_LOC_26/Y OR2X1_LOC_7/A 10.81fF
C35456 OR2X1_LOC_176/a_8_216# OR2X1_LOC_26/Y 0.07fF
C35660 OR2X1_LOC_26/Y AND2X1_LOC_836/a_8_24# 0.01fF
C36295 AND2X1_LOC_543/Y OR2X1_LOC_26/Y 0.01fF
C36347 OR2X1_LOC_589/A OR2X1_LOC_26/Y 0.03fF
C36477 AND2X1_LOC_379/a_8_24# OR2X1_LOC_26/Y 0.04fF
C36527 OR2X1_LOC_60/a_8_216# OR2X1_LOC_26/Y 0.06fF
C36782 OR2X1_LOC_26/Y OR2X1_LOC_585/Y 0.01fF
C37356 OR2X1_LOC_3/Y OR2X1_LOC_26/Y 0.29fF
C37730 AND2X1_LOC_113/Y OR2X1_LOC_26/Y 0.01fF
C37951 OR2X1_LOC_26/Y OR2X1_LOC_525/a_8_216# 0.01fF
C38110 AND2X1_LOC_113/a_36_24# OR2X1_LOC_26/Y 0.01fF
C38197 OR2X1_LOC_280/a_8_216# OR2X1_LOC_26/Y 0.01fF
C38260 OR2X1_LOC_26/Y OR2X1_LOC_72/a_8_216# 0.01fF
C38626 OR2X1_LOC_26/Y OR2X1_LOC_690/A 0.04fF
C38664 OR2X1_LOC_64/Y OR2X1_LOC_26/Y 0.36fF
C38866 AND2X1_LOC_541/a_8_24# OR2X1_LOC_26/Y 0.01fF
C39069 AND2X1_LOC_101/B OR2X1_LOC_26/Y 0.03fF
C39832 OR2X1_LOC_516/B OR2X1_LOC_26/Y 0.10fF
C40206 AND2X1_LOC_456/B OR2X1_LOC_26/Y 0.02fF
C41046 OR2X1_LOC_494/Y OR2X1_LOC_26/Y 0.03fF
C41174 OR2X1_LOC_26/Y AND2X1_LOC_839/B 0.01fF
C41283 OR2X1_LOC_26/Y OR2X1_LOC_311/a_8_216# 0.07fF
C41905 AND2X1_LOC_130/a_8_24# OR2X1_LOC_26/Y 0.01fF
C41915 OR2X1_LOC_26/Y AND2X1_LOC_778/Y 0.03fF
C42038 OR2X1_LOC_380/A OR2X1_LOC_26/Y 0.01fF
C42496 OR2X1_LOC_669/a_8_216# OR2X1_LOC_26/Y 0.01fF
C43358 OR2X1_LOC_670/Y OR2X1_LOC_26/Y 0.02fF
C44178 OR2X1_LOC_26/Y OR2X1_LOC_278/Y 0.04fF
C44240 OR2X1_LOC_26/Y AND2X1_LOC_634/a_8_24# 0.02fF
C44265 OR2X1_LOC_273/Y OR2X1_LOC_26/Y 0.09fF
C44834 OR2X1_LOC_26/Y OR2X1_LOC_142/Y 0.18fF
C44864 OR2X1_LOC_134/a_8_216# OR2X1_LOC_26/Y 0.01fF
C45060 OR2X1_LOC_26/Y OR2X1_LOC_118/Y 0.03fF
C45098 OR2X1_LOC_262/Y OR2X1_LOC_26/Y 0.18fF
C45513 OR2X1_LOC_516/a_8_216# OR2X1_LOC_26/Y 0.03fF
C45543 AND2X1_LOC_105/a_36_24# OR2X1_LOC_26/Y 0.02fF
C45560 OR2X1_LOC_26/Y OR2X1_LOC_83/a_8_216# 0.01fF
C45956 OR2X1_LOC_36/Y OR2X1_LOC_26/Y 1.71fF
C46091 OR2X1_LOC_26/Y OR2X1_LOC_419/Y 0.14fF
C46196 OR2X1_LOC_26/Y AND2X1_LOC_590/a_36_24# 0.01fF
C46243 OR2X1_LOC_177/Y OR2X1_LOC_26/Y 0.06fF
C46285 OR2X1_LOC_604/A OR2X1_LOC_26/Y 0.09fF
C46416 OR2X1_LOC_80/Y OR2X1_LOC_26/Y 0.07fF
C46858 OR2X1_LOC_26/Y OR2X1_LOC_265/Y 0.08fF
C47266 OR2X1_LOC_164/Y OR2X1_LOC_26/Y 0.03fF
C47403 AND2X1_LOC_633/Y OR2X1_LOC_26/Y 0.02fF
C47582 OR2X1_LOC_680/a_8_216# OR2X1_LOC_26/Y 0.01fF
C47628 OR2X1_LOC_131/A OR2X1_LOC_26/Y 0.03fF
C47744 OR2X1_LOC_26/Y OR2X1_LOC_237/a_8_216# 0.02fF
C47763 AND2X1_LOC_379/a_36_24# OR2X1_LOC_26/Y 0.01fF
C48108 OR2X1_LOC_26/Y AND2X1_LOC_637/a_8_24# 0.01fF
C48537 OR2X1_LOC_26/Y AND2X1_LOC_434/Y 0.02fF
C49463 AND2X1_LOC_342/a_8_24# OR2X1_LOC_26/Y 0.07fF
C49860 OR2X1_LOC_26/Y OR2X1_LOC_393/Y 0.05fF
C49921 OR2X1_LOC_272/Y OR2X1_LOC_26/Y 0.02fF
C50725 OR2X1_LOC_26/Y AND2X1_LOC_848/Y 0.05fF
C50747 OR2X1_LOC_283/Y OR2X1_LOC_26/Y 0.06fF
C51448 OR2X1_LOC_178/Y OR2X1_LOC_26/Y 0.06fF
C52243 AND2X1_LOC_361/a_8_24# OR2X1_LOC_26/Y 0.01fF
C52898 AND2X1_LOC_634/Y OR2X1_LOC_26/Y 0.01fF
C53416 OR2X1_LOC_26/Y OR2X1_LOC_437/A 0.43fF
C54047 AND2X1_LOC_729/Y OR2X1_LOC_26/Y 0.03fF
C54071 AND2X1_LOC_784/A OR2X1_LOC_26/Y 0.05fF
C54500 OR2X1_LOC_26/Y OR2X1_LOC_52/B 0.19fF
C54513 AND2X1_LOC_489/Y OR2X1_LOC_26/Y 0.02fF
C54622 OR2X1_LOC_26/Y AND2X1_LOC_216/A 0.02fF
C54855 OR2X1_LOC_165/a_8_216# OR2X1_LOC_26/Y 0.07fF
C54866 OR2X1_LOC_26/Y OR2X1_LOC_394/Y 0.01fF
C54893 OR2X1_LOC_26/Y AND2X1_LOC_286/Y 0.01fF
C54938 OR2X1_LOC_280/Y OR2X1_LOC_26/Y 5.67fF
C54975 OR2X1_LOC_22/Y OR2X1_LOC_26/Y 2.56fF
C55235 OR2X1_LOC_485/Y OR2X1_LOC_26/Y 0.02fF
C55346 OR2X1_LOC_26/Y OR2X1_LOC_39/A 2.19fF
C56112 OR2X1_LOC_51/Y OR2X1_LOC_26/Y 7.64fF
C56226 OR2X1_LOC_680/A OR2X1_LOC_26/Y 10.36fF
C57108 OR2X1_LOC_26/Y VSS -4.00fF
C70 OR2X1_LOC_36/Y OR2X1_LOC_7/Y 0.01fF
C500 AND2X1_LOC_196/Y OR2X1_LOC_36/Y 0.01fF
C660 OR2X1_LOC_36/Y OR2X1_LOC_321/a_8_216# 0.02fF
C789 AND2X1_LOC_456/B OR2X1_LOC_36/Y 0.16fF
C1092 OR2X1_LOC_36/Y OR2X1_LOC_395/Y 0.09fF
C2604 OR2X1_LOC_36/Y AND2X1_LOC_624/A 0.03fF
C2954 OR2X1_LOC_36/Y AND2X1_LOC_434/a_8_24# 0.01fF
C3603 OR2X1_LOC_36/Y OR2X1_LOC_172/a_8_216# -0.00fF
C3916 OR2X1_LOC_48/Y OR2X1_LOC_36/Y 0.01fF
C4013 OR2X1_LOC_36/Y AND2X1_LOC_779/Y 0.03fF
C4631 OR2X1_LOC_36/Y OR2X1_LOC_278/Y 0.03fF
C4708 OR2X1_LOC_273/Y OR2X1_LOC_36/Y 0.73fF
C4723 OR2X1_LOC_253/a_8_216# OR2X1_LOC_36/Y 0.01fF
C5109 AND2X1_LOC_78/a_8_24# OR2X1_LOC_36/Y 0.01fF
C5117 OR2X1_LOC_754/A OR2X1_LOC_36/Y 0.14fF
C5250 OR2X1_LOC_36/Y OR2X1_LOC_142/Y 0.02fF
C5425 OR2X1_LOC_36/Y OR2X1_LOC_16/a_8_216# 0.01fF
C5469 OR2X1_LOC_36/Y OR2X1_LOC_118/Y 0.03fF
C5529 OR2X1_LOC_36/Y OR2X1_LOC_238/Y 0.01fF
C5654 OR2X1_LOC_36/Y OR2X1_LOC_39/a_8_216# 0.01fF
C6401 OR2X1_LOC_36/Y OR2X1_LOC_65/a_8_216# 0.02fF
C6463 OR2X1_LOC_36/Y OR2X1_LOC_419/Y 1.82fF
C6666 OR2X1_LOC_604/A OR2X1_LOC_36/Y 0.36fF
C6775 OR2X1_LOC_306/Y OR2X1_LOC_36/Y 0.10fF
C7227 OR2X1_LOC_36/Y OR2X1_LOC_265/Y 0.03fF
C7453 OR2X1_LOC_36/Y OR2X1_LOC_183/a_8_216# 0.06fF
C7750 OR2X1_LOC_36/Y AND2X1_LOC_633/Y 0.02fF
C7929 AND2X1_LOC_539/Y OR2X1_LOC_36/Y 0.03fF
C8015 AND2X1_LOC_326/B OR2X1_LOC_36/Y 0.03fF
C8098 OR2X1_LOC_36/Y OR2X1_LOC_237/a_8_216# 0.01fF
C8897 OR2X1_LOC_36/Y AND2X1_LOC_434/Y 0.08fF
C9009 OR2X1_LOC_36/Y AND2X1_LOC_459/a_8_24# 0.02fF
C9113 OR2X1_LOC_36/Y OR2X1_LOC_595/Y 0.84fF
C9428 OR2X1_LOC_36/Y OR2X1_LOC_69/a_8_216# 0.01fF
C9464 AND2X1_LOC_196/a_8_24# OR2X1_LOC_36/Y 0.01fF
C10293 OR2X1_LOC_272/Y OR2X1_LOC_36/Y 0.02fF
C10599 OR2X1_LOC_36/Y OR2X1_LOC_234/Y 0.02fF
C10708 OR2X1_LOC_79/A OR2X1_LOC_36/Y 0.47fF
C10742 OR2X1_LOC_36/Y OR2X1_LOC_278/A 0.08fF
C10923 OR2X1_LOC_135/Y OR2X1_LOC_36/Y 0.01fF
C11034 OR2X1_LOC_36/Y AND2X1_LOC_520/Y 0.28fF
C11134 OR2X1_LOC_36/Y AND2X1_LOC_856/B 0.26fF
C12026 OR2X1_LOC_36/Y AND2X1_LOC_318/Y 0.01fF
C12303 OR2X1_LOC_698/Y OR2X1_LOC_36/Y 0.01fF
C13827 OR2X1_LOC_36/Y OR2X1_LOC_437/A 0.38fF
C13979 AND2X1_LOC_715/A OR2X1_LOC_36/Y 2.69fF
C14121 OR2X1_LOC_36/Y OR2X1_LOC_754/a_8_216# 0.03fF
C14478 AND2X1_LOC_729/Y OR2X1_LOC_36/Y 0.04fF
C14504 AND2X1_LOC_784/A OR2X1_LOC_36/Y 0.07fF
C14653 OR2X1_LOC_36/Y OR2X1_LOC_172/Y 0.04fF
C14935 OR2X1_LOC_36/Y OR2X1_LOC_52/B 7.04fF
C15187 OR2X1_LOC_36/Y OR2X1_LOC_253/Y 0.01fF
C15297 OR2X1_LOC_36/Y AND2X1_LOC_286/Y 0.03fF
C15339 OR2X1_LOC_280/Y OR2X1_LOC_36/Y 0.51fF
C15373 OR2X1_LOC_22/Y OR2X1_LOC_36/Y 2.68fF
C15609 OR2X1_LOC_485/Y OR2X1_LOC_36/Y 0.06fF
C15699 OR2X1_LOC_36/Y OR2X1_LOC_39/A 0.82fF
C16129 OR2X1_LOC_36/Y AND2X1_LOC_593/Y 0.01fF
C16478 OR2X1_LOC_51/Y OR2X1_LOC_36/Y 0.68fF
C16528 OR2X1_LOC_36/Y OR2X1_LOC_16/Y 0.02fF
C16577 OR2X1_LOC_680/A OR2X1_LOC_36/Y 0.33fF
C16920 AND2X1_LOC_593/a_36_24# OR2X1_LOC_36/Y 0.01fF
C17825 OR2X1_LOC_252/Y OR2X1_LOC_36/Y 0.07fF
C17882 OR2X1_LOC_36/Y OR2X1_LOC_609/A 0.03fF
C18518 OR2X1_LOC_36/Y OR2X1_LOC_183/Y 0.01fF
C18750 OR2X1_LOC_36/Y OR2X1_LOC_511/Y 0.16fF
C19155 OR2X1_LOC_36/Y OR2X1_LOC_237/Y 0.08fF
C19508 OR2X1_LOC_91/A OR2X1_LOC_36/Y 0.73fF
C20012 OR2X1_LOC_32/B OR2X1_LOC_36/Y 0.01fF
C20202 OR2X1_LOC_36/Y OR2X1_LOC_423/Y 0.53fF
C20478 OR2X1_LOC_36/Y OR2X1_LOC_74/A 0.36fF
C20750 OR2X1_LOC_36/Y AND2X1_LOC_254/a_8_24# 0.08fF
C20806 OR2X1_LOC_459/A OR2X1_LOC_36/Y 0.03fF
C20847 OR2X1_LOC_432/a_8_216# OR2X1_LOC_36/Y 0.01fF
C20889 OR2X1_LOC_36/Y AND2X1_LOC_287/Y 0.03fF
C20987 OR2X1_LOC_36/Y OR2X1_LOC_607/Y 0.01fF
C21282 OR2X1_LOC_36/Y OR2X1_LOC_432/Y 0.02fF
C21709 AND2X1_LOC_779/a_8_24# OR2X1_LOC_36/Y 0.01fF
C22082 OR2X1_LOC_816/a_8_216# OR2X1_LOC_36/Y 0.01fF
C22363 OR2X1_LOC_36/Y OR2X1_LOC_300/Y 0.28fF
C23096 OR2X1_LOC_36/Y OR2X1_LOC_65/Y 0.01fF
C23171 OR2X1_LOC_36/Y OR2X1_LOC_72/Y 0.49fF
C23504 OR2X1_LOC_696/Y OR2X1_LOC_36/Y 0.03fF
C23851 OR2X1_LOC_36/Y OR2X1_LOC_595/a_8_216# 0.14fF
C23918 OR2X1_LOC_431/a_8_216# OR2X1_LOC_36/Y 0.01fF
C24149 AND2X1_LOC_706/Y OR2X1_LOC_36/Y 0.02fF
C24305 OR2X1_LOC_665/Y OR2X1_LOC_36/Y 0.03fF
C24317 OR2X1_LOC_485/A OR2X1_LOC_36/Y 0.24fF
C24386 OR2X1_LOC_36/Y OR2X1_LOC_609/Y 0.01fF
C24703 OR2X1_LOC_495/a_8_216# OR2X1_LOC_36/Y 0.07fF
C24787 OR2X1_LOC_36/Y OR2X1_LOC_238/a_8_216# 0.01fF
C24874 OR2X1_LOC_36/Y OR2X1_LOC_376/Y 0.05fF
C25140 OR2X1_LOC_36/Y OR2X1_LOC_754/a_36_216# 0.02fF
C25687 OR2X1_LOC_36/Y OR2X1_LOC_589/Y 0.01fF
C25924 OR2X1_LOC_305/a_8_216# OR2X1_LOC_36/Y 0.01fF
C25994 AND2X1_LOC_537/Y OR2X1_LOC_36/Y 0.03fF
C26672 OR2X1_LOC_526/Y OR2X1_LOC_36/Y 0.03fF
C26758 OR2X1_LOC_36/Y OR2X1_LOC_433/Y 0.03fF
C27473 OR2X1_LOC_492/a_8_216# OR2X1_LOC_36/Y 0.01fF
C27795 OR2X1_LOC_36/Y OR2X1_LOC_589/a_8_216# 0.19fF
C27835 OR2X1_LOC_516/Y OR2X1_LOC_36/Y 0.03fF
C28212 OR2X1_LOC_36/Y AND2X1_LOC_793/B 0.03fF
C28917 OR2X1_LOC_36/Y OR2X1_LOC_609/a_8_216# 0.02fF
C29197 VDD OR2X1_LOC_36/Y 1.17fF
C29292 OR2X1_LOC_315/Y OR2X1_LOC_36/Y 0.30fF
C29321 OR2X1_LOC_36/Y OR2X1_LOC_491/Y 0.01fF
C29326 OR2X1_LOC_251/Y OR2X1_LOC_36/Y 0.03fF
C29426 OR2X1_LOC_36/Y OR2X1_LOC_67/Y 0.07fF
C29977 OR2X1_LOC_36/Y OR2X1_LOC_56/Y 0.01fF
C30215 OR2X1_LOC_36/Y AND2X1_LOC_307/Y 0.15fF
C30524 OR2X1_LOC_36/Y OR2X1_LOC_427/A 0.47fF
C31077 OR2X1_LOC_36/Y OR2X1_LOC_416/Y 0.04fF
C31183 OR2X1_LOC_36/Y AND2X1_LOC_592/a_8_24# 0.01fF
C31546 OR2X1_LOC_36/Y AND2X1_LOC_463/B 0.03fF
C31798 OR2X1_LOC_36/Y OR2X1_LOC_45/a_8_216# 0.01fF
C31827 OR2X1_LOC_36/Y AND2X1_LOC_831/a_8_24# 0.01fF
C32060 OR2X1_LOC_45/B OR2X1_LOC_36/Y 5.76fF
C32204 OR2X1_LOC_36/Y AND2X1_LOC_435/a_8_24# 0.01fF
C32215 OR2X1_LOC_36/Y OR2X1_LOC_767/a_8_216# 0.08fF
C32540 OR2X1_LOC_158/A OR2X1_LOC_36/Y 0.73fF
C32977 OR2X1_LOC_482/Y OR2X1_LOC_36/Y 0.06fF
C33021 OR2X1_LOC_816/Y OR2X1_LOC_36/Y 0.01fF
C33156 OR2X1_LOC_304/Y OR2X1_LOC_36/Y 0.43fF
C34046 OR2X1_LOC_111/Y OR2X1_LOC_36/Y 0.03fF
C34223 OR2X1_LOC_591/Y OR2X1_LOC_36/Y 0.03fF
C34796 OR2X1_LOC_316/Y OR2X1_LOC_36/Y 0.02fF
C34856 AND2X1_LOC_390/B OR2X1_LOC_36/Y 0.07fF
C34879 OR2X1_LOC_431/Y OR2X1_LOC_36/Y 0.01fF
C35125 OR2X1_LOC_744/A OR2X1_LOC_36/Y 0.48fF
C35201 OR2X1_LOC_36/Y AND2X1_LOC_840/B 0.59fF
C35377 OR2X1_LOC_36/Y OR2X1_LOC_320/a_8_216# 0.03fF
C35453 OR2X1_LOC_36/Y OR2X1_LOC_79/a_8_216# 0.01fF
C35701 OR2X1_LOC_36/Y AND2X1_LOC_308/a_8_24# 0.01fF
C35986 OR2X1_LOC_179/a_8_216# OR2X1_LOC_36/Y 0.07fF
C36378 OR2X1_LOC_36/Y OR2X1_LOC_56/A 1.58fF
C36765 OR2X1_LOC_36/Y AND2X1_LOC_285/Y 0.17fF
C36863 OR2X1_LOC_91/Y OR2X1_LOC_36/Y 0.03fF
C36881 OR2X1_LOC_305/Y OR2X1_LOC_36/Y 0.01fF
C36926 OR2X1_LOC_417/Y OR2X1_LOC_36/Y 0.03fF
C36929 OR2X1_LOC_291/Y OR2X1_LOC_36/Y 0.06fF
C36936 OR2X1_LOC_311/Y OR2X1_LOC_36/Y 0.03fF
C37417 AND2X1_LOC_831/Y OR2X1_LOC_36/Y 0.08fF
C37720 OR2X1_LOC_36/Y AND2X1_LOC_436/B 0.01fF
C37726 OR2X1_LOC_36/Y AND2X1_LOC_139/B 0.03fF
C37988 OR2X1_LOC_135/a_8_216# OR2X1_LOC_36/Y 0.01fF
C38251 OR2X1_LOC_36/Y OR2X1_LOC_71/Y 0.03fF
C38448 OR2X1_LOC_492/Y OR2X1_LOC_36/Y 0.01fF
C38673 OR2X1_LOC_36/Y OR2X1_LOC_246/A 0.86fF
C39058 OR2X1_LOC_497/Y OR2X1_LOC_36/Y 0.07fF
C39537 OR2X1_LOC_36/Y OR2X1_LOC_7/a_8_216# 0.01fF
C39813 OR2X1_LOC_235/B OR2X1_LOC_36/Y 0.02fF
C39881 AND2X1_LOC_319/A OR2X1_LOC_36/Y 0.03fF
C40262 AND2X1_LOC_318/a_8_24# OR2X1_LOC_36/Y 0.01fF
C40501 OR2X1_LOC_36/Y OR2X1_LOC_395/a_8_216# 0.02fF
C41586 OR2X1_LOC_36/Y OR2X1_LOC_65/B 0.03fF
C41880 OR2X1_LOC_692/Y OR2X1_LOC_36/Y 0.04fF
C41919 OR2X1_LOC_600/A OR2X1_LOC_36/Y 0.54fF
C42000 OR2X1_LOC_36/Y OR2X1_LOC_619/Y 0.18fF
C42373 OR2X1_LOC_36/Y AND2X1_LOC_286/a_8_24# 0.02fF
C42501 OR2X1_LOC_36/Y OR2X1_LOC_232/a_8_216# 0.14fF
C43319 OR2X1_LOC_36/Y OR2X1_LOC_69/A 0.17fF
C44263 AND2X1_LOC_307/a_8_24# OR2X1_LOC_36/Y 0.01fF
C44387 OR2X1_LOC_36/Y OR2X1_LOC_13/B 1.08fF
C44890 OR2X1_LOC_36/Y OR2X1_LOC_428/A 0.23fF
C45370 AND2X1_LOC_592/Y OR2X1_LOC_36/Y 0.04fF
C45977 OR2X1_LOC_36/Y OR2X1_LOC_89/A 0.12fF
C46662 OR2X1_LOC_36/Y OR2X1_LOC_79/Y 0.01fF
C46706 OR2X1_LOC_491/a_8_216# OR2X1_LOC_36/Y 0.02fF
C46816 OR2X1_LOC_45/Y OR2X1_LOC_36/Y 0.30fF
C46866 OR2X1_LOC_36/Y OR2X1_LOC_824/Y 0.01fF
C46870 OR2X1_LOC_36/Y OR2X1_LOC_591/a_8_216# 0.01fF
C46918 OR2X1_LOC_36/Y AND2X1_LOC_727/A 0.04fF
C46941 OR2X1_LOC_36/Y OR2X1_LOC_95/Y 0.05fF
C47280 OR2X1_LOC_36/Y AND2X1_LOC_832/a_8_24# 0.01fF
C47606 OR2X1_LOC_693/Y OR2X1_LOC_36/Y 0.01fF
C47727 OR2X1_LOC_36/Y AND2X1_LOC_621/Y 0.05fF
C47918 OR2X1_LOC_36/Y OR2X1_LOC_71/A 0.02fF
C48239 OR2X1_LOC_70/Y OR2X1_LOC_36/Y 1.46fF
C48315 OR2X1_LOC_36/Y OR2X1_LOC_184/Y 0.03fF
C48890 OR2X1_LOC_36/Y OR2X1_LOC_607/A 0.04fF
C48981 OR2X1_LOC_625/Y OR2X1_LOC_36/Y 0.08fF
C49712 OR2X1_LOC_36/Y OR2X1_LOC_16/A 1.45fF
C49765 OR2X1_LOC_108/Y OR2X1_LOC_36/Y 0.13fF
C49951 OR2X1_LOC_36/Y AND2X1_LOC_687/Y 0.03fF
C50609 OR2X1_LOC_36/Y AND2X1_LOC_447/Y 0.03fF
C50739 OR2X1_LOC_262/a_8_216# OR2X1_LOC_36/Y 0.05fF
C50770 OR2X1_LOC_36/Y AND2X1_LOC_729/B 0.03fF
C51001 AND2X1_LOC_593/a_8_24# OR2X1_LOC_36/Y 0.04fF
C51056 OR2X1_LOC_39/Y OR2X1_LOC_36/Y 0.01fF
C51216 AND2X1_LOC_227/Y OR2X1_LOC_36/Y 0.03fF
C51540 OR2X1_LOC_599/A OR2X1_LOC_36/Y 0.35fF
C51851 OR2X1_LOC_40/Y OR2X1_LOC_36/Y 0.17fF
C51892 OR2X1_LOC_698/a_8_216# OR2X1_LOC_36/Y 0.01fF
C51940 OR2X1_LOC_36/Y OR2X1_LOC_424/a_8_216# 0.01fF
C51982 OR2X1_LOC_36/Y OR2X1_LOC_7/A 0.63fF
C52003 OR2X1_LOC_320/Y OR2X1_LOC_36/Y 0.01fF
C52242 OR2X1_LOC_491/a_36_216# OR2X1_LOC_36/Y 0.02fF
C52489 OR2X1_LOC_36/Y OR2X1_LOC_615/Y 0.07fF
C52572 OR2X1_LOC_36/Y OR2X1_LOC_424/Y 0.01fF
C52635 AND2X1_LOC_707/Y OR2X1_LOC_36/Y 0.01fF
C52773 OR2X1_LOC_36/Y AND2X1_LOC_841/B 0.01fF
C53097 AND2X1_LOC_706/a_8_24# OR2X1_LOC_36/Y 0.01fF
C53107 OR2X1_LOC_589/A OR2X1_LOC_36/Y 0.52fF
C54087 OR2X1_LOC_3/Y OR2X1_LOC_36/Y 1.40fF
C54921 OR2X1_LOC_280/a_8_216# OR2X1_LOC_36/Y 0.01fF
C54981 OR2X1_LOC_36/Y OR2X1_LOC_607/a_8_216# 0.02fF
C55368 OR2X1_LOC_36/Y OR2X1_LOC_690/A 0.02fF
C55400 OR2X1_LOC_64/Y OR2X1_LOC_36/Y 4.52fF
C57232 OR2X1_LOC_36/Y VSS 0.85fF
C369 OR2X1_LOC_693/Y OR2X1_LOC_22/Y 0.11fF
C990 OR2X1_LOC_70/Y OR2X1_LOC_22/Y 2.22fF
C1011 AND2X1_LOC_538/a_8_24# OR2X1_LOC_22/Y 0.01fF
C1049 OR2X1_LOC_22/Y OR2X1_LOC_184/Y 0.19fF
C1778 OR2X1_LOC_625/Y OR2X1_LOC_22/Y 0.02fF
C2123 AND2X1_LOC_535/Y OR2X1_LOC_22/Y 0.03fF
C2542 OR2X1_LOC_22/Y OR2X1_LOC_16/A 0.30fF
C2587 OR2X1_LOC_108/Y OR2X1_LOC_22/Y 0.94fF
C2738 OR2X1_LOC_22/Y AND2X1_LOC_687/Y 0.02fF
C3564 OR2X1_LOC_22/Y AND2X1_LOC_729/B 0.08fF
C4016 OR2X1_LOC_22/Y AND2X1_LOC_227/Y 0.07fF
C4050 OR2X1_LOC_22/Y OR2X1_LOC_41/Y 0.28fF
C4247 OR2X1_LOC_107/Y OR2X1_LOC_22/Y 0.03fF
C4321 OR2X1_LOC_599/A OR2X1_LOC_22/Y 0.09fF
C4621 OR2X1_LOC_40/Y OR2X1_LOC_22/Y 0.25fF
C4748 OR2X1_LOC_22/Y OR2X1_LOC_7/A 0.62fF
C5157 OR2X1_LOC_22/Y OR2X1_LOC_32/a_8_216# 0.01fF
C5185 OR2X1_LOC_22/Y AND2X1_LOC_115/a_8_24# -0.01fF
C5881 AND2X1_LOC_706/a_8_24# OR2X1_LOC_22/Y 0.02fF
C5891 OR2X1_LOC_589/A OR2X1_LOC_22/Y 0.49fF
C6037 OR2X1_LOC_22/Y OR2X1_LOC_60/a_8_216# 0.01fF
C6317 OR2X1_LOC_22/Y OR2X1_LOC_585/Y 0.08fF
C6908 OR2X1_LOC_3/Y OR2X1_LOC_22/Y 2.56fF
C6975 OR2X1_LOC_22/Y AND2X1_LOC_462/B 0.72fF
C7266 OR2X1_LOC_74/Y OR2X1_LOC_22/Y 0.06fF
C7297 OR2X1_LOC_22/Y AND2X1_LOC_113/Y 0.06fF
C8192 OR2X1_LOC_503/A OR2X1_LOC_22/Y 0.01fF
C8216 OR2X1_LOC_22/Y OR2X1_LOC_690/A 0.40fF
C8252 OR2X1_LOC_22/Y OR2X1_LOC_64/Y 1.30fF
C9090 OR2X1_LOC_22/Y OR2X1_LOC_829/Y 0.01fF
C9528 OR2X1_LOC_22/Y OR2X1_LOC_279/Y 0.16fF
C9849 AND2X1_LOC_456/B OR2X1_LOC_22/Y 0.06fF
C10799 OR2X1_LOC_22/Y AND2X1_LOC_116/B 0.01fF
C10843 OR2X1_LOC_22/Y OR2X1_LOC_311/a_8_216# 0.03fF
C10990 OR2X1_LOC_22/Y AND2X1_LOC_802/Y 0.15fF
C11546 OR2X1_LOC_521/Y OR2X1_LOC_22/Y 0.03fF
C11577 OR2X1_LOC_380/A OR2X1_LOC_22/Y 0.05fF
C11922 OR2X1_LOC_22/Y AND2X1_LOC_434/a_8_24# 0.02fF
C13702 OR2X1_LOC_22/Y OR2X1_LOC_278/Y 0.03fF
C13753 OR2X1_LOC_273/Y OR2X1_LOC_22/Y 0.14fF
C13800 OR2X1_LOC_22/Y OR2X1_LOC_75/Y 0.02fF
C14190 OR2X1_LOC_22/Y OR2X1_LOC_754/A 0.44fF
C14539 OR2X1_LOC_22/Y OR2X1_LOC_118/Y 0.03fF
C14615 OR2X1_LOC_22/Y AND2X1_LOC_855/a_8_24# 0.01fF
C15478 OR2X1_LOC_22/Y OR2X1_LOC_419/Y 0.03fF
C15680 OR2X1_LOC_604/A OR2X1_LOC_22/Y 0.10fF
C15769 OR2X1_LOC_306/Y OR2X1_LOC_22/Y 0.03fF
C15782 OR2X1_LOC_22/Y OR2X1_LOC_80/Y 0.01fF
C16222 OR2X1_LOC_22/Y OR2X1_LOC_265/Y 0.07fF
C16686 OR2X1_LOC_22/Y OR2X1_LOC_230/a_8_216# 0.04fF
C16708 OR2X1_LOC_22/Y AND2X1_LOC_633/Y 0.03fF
C16923 AND2X1_LOC_539/Y OR2X1_LOC_22/Y 0.07fF
C17313 OR2X1_LOC_316/a_8_216# OR2X1_LOC_22/Y 0.05fF
C17843 OR2X1_LOC_22/Y AND2X1_LOC_434/Y 0.44fF
C18048 OR2X1_LOC_22/Y OR2X1_LOC_595/Y 0.02fF
C18351 OR2X1_LOC_837/B OR2X1_LOC_22/Y 0.03fF
C19259 OR2X1_LOC_272/Y OR2X1_LOC_22/Y 0.05fF
C19608 OR2X1_LOC_517/a_8_216# OR2X1_LOC_22/Y 0.01fF
C20064 OR2X1_LOC_22/Y AND2X1_LOC_520/Y 0.01fF
C20141 OR2X1_LOC_22/Y AND2X1_LOC_856/B 0.01fF
C21249 OR2X1_LOC_22/Y OR2X1_LOC_829/A 0.17fF
C21493 OR2X1_LOC_22/Y OR2X1_LOC_224/Y 0.03fF
C21837 OR2X1_LOC_385/Y OR2X1_LOC_22/Y 0.04fF
C22108 OR2X1_LOC_22/Y AND2X1_LOC_810/B 0.07fF
C22874 OR2X1_LOC_22/Y OR2X1_LOC_437/A 0.10fF
C23029 AND2X1_LOC_715/A OR2X1_LOC_22/Y 0.01fF
C23512 AND2X1_LOC_729/Y OR2X1_LOC_22/Y 0.07fF
C23532 AND2X1_LOC_784/A OR2X1_LOC_22/Y 0.03fF
C23653 OR2X1_LOC_22/Y OR2X1_LOC_172/Y 0.15fF
C23948 OR2X1_LOC_22/Y OR2X1_LOC_52/B 0.40fF
C24242 OR2X1_LOC_22/Y OR2X1_LOC_13/a_8_216# 0.03fF
C24358 AND2X1_LOC_356/B OR2X1_LOC_22/Y 0.03fF
C24359 OR2X1_LOC_280/Y OR2X1_LOC_22/Y 0.07fF
C24758 OR2X1_LOC_22/Y OR2X1_LOC_39/A 0.12fF
C25245 OR2X1_LOC_22/Y OR2X1_LOC_226/Y 0.01fF
C25501 OR2X1_LOC_51/Y OR2X1_LOC_22/Y 0.14fF
C25531 OR2X1_LOC_22/Y OR2X1_LOC_58/a_8_216# 0.01fF
C26324 OR2X1_LOC_22/Y AND2X1_LOC_436/Y 0.08fF
C26426 OR2X1_LOC_22/Y OR2X1_LOC_588/Y 0.03fF
C28403 OR2X1_LOC_22/Y OR2X1_LOC_522/a_8_216# 0.08fF
C28480 OR2X1_LOC_22/Y OR2X1_LOC_91/A 0.94fF
C28580 OR2X1_LOC_22/Y OR2X1_LOC_27/Y 0.03fF
C28941 OR2X1_LOC_32/B OR2X1_LOC_22/Y 0.09fF
C29408 OR2X1_LOC_22/Y OR2X1_LOC_74/A 0.16fF
C29785 OR2X1_LOC_432/a_8_216# OR2X1_LOC_22/Y 0.01fF
C30201 OR2X1_LOC_22/Y OR2X1_LOC_432/Y 0.04fF
C30205 OR2X1_LOC_22/Y AND2X1_LOC_287/a_8_24# 0.06fF
C30670 OR2X1_LOC_22/Y OR2X1_LOC_615/a_8_216# 0.02fF
C31232 OR2X1_LOC_22/Y OR2X1_LOC_521/a_8_216# 0.01fF
C31324 OR2X1_LOC_106/Y OR2X1_LOC_22/Y 0.01fF
C31482 OR2X1_LOC_497/a_8_216# OR2X1_LOC_22/Y 0.01fF
C32002 OR2X1_LOC_22/Y OR2X1_LOC_72/Y 0.02fF
C32742 OR2X1_LOC_22/Y OR2X1_LOC_595/a_8_216# 0.02fF
C33038 AND2X1_LOC_706/Y OR2X1_LOC_22/Y 0.03fF
C33066 OR2X1_LOC_58/Y OR2X1_LOC_22/Y 0.43fF
C33206 OR2X1_LOC_485/A OR2X1_LOC_22/Y 9.27fF
C33777 OR2X1_LOC_22/Y OR2X1_LOC_385/a_8_216# 0.10fF
C34039 OR2X1_LOC_32/Y OR2X1_LOC_22/Y 0.04fF
C34942 AND2X1_LOC_537/Y OR2X1_LOC_22/Y 0.02fF
C35087 OR2X1_LOC_22/Y OR2X1_LOC_171/a_8_216# 0.03fF
C35156 OR2X1_LOC_22/Y OR2X1_LOC_13/Y 0.19fF
C35688 OR2X1_LOC_22/Y OR2X1_LOC_433/Y 0.02fF
C36167 OR2X1_LOC_22/Y OR2X1_LOC_615/a_36_216# 0.03fF
C36678 OR2X1_LOC_22/Y OR2X1_LOC_589/a_8_216# 0.03fF
C36736 AND2X1_LOC_798/a_8_24# OR2X1_LOC_22/Y 0.03fF
C38116 VDD OR2X1_LOC_22/Y 0.95fF
C38208 OR2X1_LOC_22/Y OR2X1_LOC_829/a_8_216# 0.01fF
C38248 OR2X1_LOC_251/Y OR2X1_LOC_22/Y 0.03fF
C38325 OR2X1_LOC_22/Y OR2X1_LOC_67/Y 0.08fF
C38558 OR2X1_LOC_60/Y OR2X1_LOC_22/Y 0.01fF
C39508 OR2X1_LOC_22/Y OR2X1_LOC_427/A 0.64fF
C39970 OR2X1_LOC_22/Y OR2X1_LOC_416/Y 0.03fF
C40613 OR2X1_LOC_22/Y OR2X1_LOC_184/a_8_216# 0.03fF
C41063 OR2X1_LOC_45/B OR2X1_LOC_22/Y 0.40fF
C41198 OR2X1_LOC_22/Y AND2X1_LOC_435/a_8_24# 0.01fF
C41214 OR2X1_LOC_22/Y OR2X1_LOC_767/a_8_216# 0.02fF
C41543 OR2X1_LOC_158/A OR2X1_LOC_22/Y 2.94fF
C41628 OR2X1_LOC_103/Y OR2X1_LOC_22/Y 0.08fF
C41648 OR2X1_LOC_103/a_8_216# OR2X1_LOC_22/Y 0.01fF
C42071 OR2X1_LOC_22/Y OR2X1_LOC_586/Y 0.03fF
C43517 OR2X1_LOC_22/Y OR2X1_LOC_41/a_8_216# 0.02fF
C43678 OR2X1_LOC_22/Y AND2X1_LOC_227/a_8_24# 0.01fF
C43732 AND2X1_LOC_541/Y OR2X1_LOC_22/Y 0.02fF
C43768 OR2X1_LOC_107/a_8_216# OR2X1_LOC_22/Y 0.05fF
C43839 OR2X1_LOC_22/Y OR2X1_LOC_316/Y 0.03fF
C43880 AND2X1_LOC_390/B OR2X1_LOC_22/Y 0.15fF
C43895 OR2X1_LOC_431/Y OR2X1_LOC_22/Y 0.42fF
C44163 OR2X1_LOC_309/Y OR2X1_LOC_22/Y 0.01fF
C44194 OR2X1_LOC_744/A OR2X1_LOC_22/Y 0.74fF
C44286 OR2X1_LOC_22/Y OR2X1_LOC_74/a_8_216# 0.05fF
C44610 OR2X1_LOC_694/Y OR2X1_LOC_22/Y 0.01fF
C45003 OR2X1_LOC_22/Y OR2X1_LOC_522/Y 0.03fF
C45421 OR2X1_LOC_118/a_8_216# OR2X1_LOC_22/Y 0.02fF
C45494 OR2X1_LOC_22/Y OR2X1_LOC_56/A 0.21fF
C46016 OR2X1_LOC_91/Y OR2X1_LOC_22/Y 0.07fF
C46073 OR2X1_LOC_291/Y OR2X1_LOC_22/Y 0.12fF
C46075 OR2X1_LOC_311/Y OR2X1_LOC_22/Y 1.36fF
C46081 AND2X1_LOC_538/Y OR2X1_LOC_22/Y 0.01fF
C46267 OR2X1_LOC_22/Y OR2X1_LOC_171/Y 0.39fF
C46513 OR2X1_LOC_22/Y AND2X1_LOC_276/Y 0.01fF
C46897 OR2X1_LOC_22/Y AND2X1_LOC_436/B 0.07fF
C46903 OR2X1_LOC_22/Y AND2X1_LOC_287/a_36_24# 0.01fF
C46908 OR2X1_LOC_22/Y AND2X1_LOC_139/B 0.07fF
C46914 OR2X1_LOC_22/Y OR2X1_LOC_767/a_36_216# 0.02fF
C47457 OR2X1_LOC_22/Y OR2X1_LOC_71/Y 2.30fF
C47706 OR2X1_LOC_108/a_8_216# OR2X1_LOC_22/Y 0.05fF
C47813 OR2X1_LOC_517/Y OR2X1_LOC_22/Y 0.03fF
C47871 OR2X1_LOC_22/Y OR2X1_LOC_246/A 1.33fF
C47895 OR2X1_LOC_22/Y OR2X1_LOC_409/B 0.03fF
C48065 AND2X1_LOC_798/a_36_24# OR2X1_LOC_22/Y 0.01fF
C48270 OR2X1_LOC_497/Y OR2X1_LOC_22/Y 0.03fF
C48677 OR2X1_LOC_22/Y OR2X1_LOC_24/a_8_216# 0.05fF
C49066 OR2X1_LOC_22/Y AND2X1_LOC_319/A 0.07fF
C49534 OR2X1_LOC_22/Y AND2X1_LOC_361/A 0.07fF
C50266 OR2X1_LOC_695/Y OR2X1_LOC_22/Y 0.09fF
C50774 OR2X1_LOC_22/Y OR2X1_LOC_65/B 0.03fF
C51053 OR2X1_LOC_692/Y OR2X1_LOC_22/Y 0.03fF
C51093 OR2X1_LOC_600/A OR2X1_LOC_22/Y 0.20fF
C51157 OR2X1_LOC_22/Y OR2X1_LOC_619/Y 0.14fF
C51671 AND2X1_LOC_539/a_8_24# OR2X1_LOC_22/Y 0.01fF
C52844 AND2X1_LOC_113/a_8_24# OR2X1_LOC_22/Y 0.03fF
C53308 OR2X1_LOC_312/Y OR2X1_LOC_22/Y 0.06fF
C53483 OR2X1_LOC_22/Y OR2X1_LOC_13/B 0.77fF
C53982 OR2X1_LOC_22/Y OR2X1_LOC_428/A 12.95fF
C53995 OR2X1_LOC_22/Y OR2X1_LOC_595/A 2.95fF
C54578 OR2X1_LOC_22/Y OR2X1_LOC_279/a_8_216# 0.04fF
C54985 OR2X1_LOC_22/Y OR2X1_LOC_89/A 0.18fF
C55663 OR2X1_LOC_22/Y AND2X1_LOC_473/Y 0.10fF
C55672 OR2X1_LOC_22/Y AND2X1_LOC_287/B 0.04fF
C55833 OR2X1_LOC_45/Y OR2X1_LOC_22/Y 0.41fF
C55909 OR2X1_LOC_22/Y AND2X1_LOC_727/A 0.03fF
C55932 OR2X1_LOC_22/Y OR2X1_LOC_95/Y 0.23fF
C57307 OR2X1_LOC_22/Y VSS 0.85fF
C2437 AND2X1_LOC_548/Y AND2X1_LOC_549/a_8_24# 0.03fF
C9099 AND2X1_LOC_548/Y OR2X1_LOC_437/A 0.01fF
C10956 AND2X1_LOC_548/Y OR2X1_LOC_39/A 0.01fF
C11836 OR2X1_LOC_680/A AND2X1_LOC_548/Y 0.89fF
C13485 AND2X1_LOC_548/Y AND2X1_LOC_549/a_36_24# 0.01fF
C15665 AND2X1_LOC_548/Y OR2X1_LOC_74/A 0.11fF
C24484 VDD AND2X1_LOC_548/Y 0.01fF
C27385 OR2X1_LOC_45/B AND2X1_LOC_548/Y 0.03fF
C40512 OR2X1_LOC_528/Y AND2X1_LOC_548/Y 0.06fF
C42060 AND2X1_LOC_548/Y OR2X1_LOC_95/Y 0.26fF
C47092 OR2X1_LOC_40/Y AND2X1_LOC_548/Y 0.14fF
C53956 AND2X1_LOC_548/Y AND2X1_LOC_624/A 0.05fF
C57558 AND2X1_LOC_548/Y VSS 0.11fF
C1146 OR2X1_LOC_709/A OR2X1_LOC_154/A 0.09fF
C6981 OR2X1_LOC_709/A VDD 0.21fF
C7853 OR2X1_LOC_709/A OR2X1_LOC_676/Y 0.01fF
C9198 OR2X1_LOC_709/A OR2X1_LOC_840/A 0.10fF
C9286 OR2X1_LOC_709/A OR2X1_LOC_789/a_8_216# 0.01fF
C10486 OR2X1_LOC_709/A OR2X1_LOC_447/A 0.02fF
C11828 OR2X1_LOC_709/A OR2X1_LOC_702/A 1.01fF
C13518 OR2X1_LOC_709/A OR2X1_LOC_778/Y 0.10fF
C13778 OR2X1_LOC_709/A AND2X1_LOC_91/B 0.16fF
C14156 OR2X1_LOC_709/A OR2X1_LOC_446/B 0.40fF
C14344 OR2X1_LOC_709/A AND2X1_LOC_56/B 0.06fF
C15677 OR2X1_LOC_709/A AND2X1_LOC_47/Y 0.03fF
C15964 OR2X1_LOC_709/A OR2X1_LOC_506/A 0.03fF
C19681 OR2X1_LOC_709/A OR2X1_LOC_317/B 0.08fF
C19734 OR2X1_LOC_709/A AND2X1_LOC_44/Y 0.46fF
C20315 OR2X1_LOC_709/A OR2X1_LOC_793/B 0.01fF
C20631 OR2X1_LOC_709/A AND2X1_LOC_18/Y 0.03fF
C20951 OR2X1_LOC_709/A OR2X1_LOC_789/A 0.22fF
C21570 OR2X1_LOC_709/A OR2X1_LOC_447/a_8_216# 0.02fF
C22042 OR2X1_LOC_709/A OR2X1_LOC_449/B 0.09fF
C23409 OR2X1_LOC_709/A OR2X1_LOC_447/Y 0.02fF
C23697 OR2X1_LOC_709/A OR2X1_LOC_161/A 0.03fF
C23783 OR2X1_LOC_709/A AND2X1_LOC_51/Y 0.05fF
C25181 OR2X1_LOC_709/A OR2X1_LOC_704/a_8_216# 0.04fF
C25968 OR2X1_LOC_709/A AND2X1_LOC_31/Y 0.03fF
C26874 OR2X1_LOC_709/A AND2X1_LOC_36/Y 0.07fF
C27797 OR2X1_LOC_709/A AND2X1_LOC_313/a_8_24# 0.04fF
C29171 OR2X1_LOC_709/A OR2X1_LOC_269/B 0.10fF
C30241 OR2X1_LOC_709/A OR2X1_LOC_777/B 0.02fF
C30707 OR2X1_LOC_709/A OR2X1_LOC_161/B 0.07fF
C32932 OR2X1_LOC_709/A OR2X1_LOC_789/B 0.01fF
C33249 OR2X1_LOC_709/A AND2X1_LOC_7/B 0.01fF
C34993 OR2X1_LOC_709/A OR2X1_LOC_160/B 0.13fF
C36132 OR2X1_LOC_709/A OR2X1_LOC_714/A 0.04fF
C38261 OR2X1_LOC_709/A OR2X1_LOC_308/Y 1.17fF
C38463 OR2X1_LOC_709/A AND2X1_LOC_516/a_8_24# 0.01fF
C38796 OR2X1_LOC_709/A AND2X1_LOC_313/a_36_24# 0.01fF
C41378 OR2X1_LOC_709/A AND2X1_LOC_423/a_8_24# 0.02fF
C41497 OR2X1_LOC_709/A OR2X1_LOC_193/A 0.54fF
C43081 OR2X1_LOC_709/A OR2X1_LOC_715/B 0.11fF
C43628 OR2X1_LOC_709/A OR2X1_LOC_793/A 0.18fF
C44042 OR2X1_LOC_709/A OR2X1_LOC_687/Y 0.03fF
C44830 OR2X1_LOC_709/A OR2X1_LOC_78/A 0.07fF
C47099 OR2X1_LOC_709/A OR2X1_LOC_623/B 0.03fF
C49752 OR2X1_LOC_709/A OR2X1_LOC_574/A 0.05fF
C50483 OR2X1_LOC_709/A OR2X1_LOC_78/B 0.09fF
C50808 OR2X1_LOC_709/A OR2X1_LOC_515/Y 0.01fF
C52612 OR2X1_LOC_709/A AND2X1_LOC_423/a_36_24# 0.01fF
C53819 OR2X1_LOC_709/A OR2X1_LOC_138/A 0.31fF
C58094 OR2X1_LOC_709/A VSS -0.65fF
C5730 VDD OR2X1_LOC_706/A 0.21fF
C13880 OR2X1_LOC_790/A OR2X1_LOC_706/A 0.28fF
C18507 OR2X1_LOC_706/A AND2X1_LOC_44/Y 0.01fF
C19404 OR2X1_LOC_706/A AND2X1_LOC_18/Y 0.01fF
C23302 AND2X1_LOC_41/A OR2X1_LOC_706/A 0.01fF
C33781 OR2X1_LOC_160/B OR2X1_LOC_706/A 0.23fF
C42489 AND2X1_LOC_45/a_8_24# OR2X1_LOC_706/A 0.20fF
C48204 OR2X1_LOC_196/B OR2X1_LOC_706/A 0.28fF
C49264 OR2X1_LOC_706/A OR2X1_LOC_78/B 0.03fF
C49371 OR2X1_LOC_706/A OR2X1_LOC_375/A 0.01fF
C53696 OR2X1_LOC_706/B OR2X1_LOC_706/A 0.16fF
C57214 OR2X1_LOC_706/A VSS -0.32fF
C666 OR2X1_LOC_310/Y OR2X1_LOC_56/A 0.03fF
C2008 OR2X1_LOC_310/Y AND2X1_LOC_335/a_8_24# 0.01fF
C6159 OR2X1_LOC_310/Y AND2X1_LOC_335/Y 0.79fF
C15943 OR2X1_LOC_40/Y OR2X1_LOC_310/Y 0.01fF
C32267 OR2X1_LOC_310/Y AND2X1_LOC_318/Y 0.06fF
C34722 AND2X1_LOC_784/A OR2X1_LOC_310/Y 0.03fF
C49684 VDD OR2X1_LOC_310/Y 0.04fF
C53025 OR2X1_LOC_158/A OR2X1_LOC_310/Y 0.08fF
C57546 OR2X1_LOC_310/Y VSS 0.08fF
C575 OR2X1_LOC_371/Y OR2X1_LOC_406/A 0.01fF
C3502 OR2X1_LOC_89/A OR2X1_LOC_371/Y 0.07fF
C4361 OR2X1_LOC_95/Y OR2X1_LOC_371/Y 0.10fF
C5567 OR2X1_LOC_70/Y OR2X1_LOC_371/Y 0.03fF
C10997 AND2X1_LOC_776/a_8_24# OR2X1_LOC_371/Y 0.01fF
C12885 OR2X1_LOC_64/Y OR2X1_LOC_371/Y 0.15fF
C18944 OR2X1_LOC_371/Y OR2X1_LOC_142/Y 0.06fF
C19216 OR2X1_LOC_238/Y OR2X1_LOC_371/Y 0.02fF
C20186 OR2X1_LOC_419/Y OR2X1_LOC_371/Y 0.10fF
C20361 OR2X1_LOC_604/A OR2X1_LOC_371/Y 0.10fF
C21279 OR2X1_LOC_164/Y OR2X1_LOC_371/Y 0.05fF
C24127 AND2X1_LOC_776/Y OR2X1_LOC_371/Y 0.27fF
C24781 AND2X1_LOC_464/Y OR2X1_LOC_371/Y 0.04fF
C27398 OR2X1_LOC_371/Y OR2X1_LOC_437/A 0.10fF
C28109 AND2X1_LOC_778/a_8_24# OR2X1_LOC_371/Y -0.00fF
C28949 OR2X1_LOC_280/Y OR2X1_LOC_371/Y 0.07fF
C29325 OR2X1_LOC_371/Y OR2X1_LOC_39/A 0.10fF
C30102 OR2X1_LOC_51/Y OR2X1_LOC_371/Y 0.07fF
C37792 OR2X1_LOC_485/A OR2X1_LOC_371/Y 0.07fF
C38624 AND2X1_LOC_458/Y OR2X1_LOC_371/Y 0.03fF
C41394 OR2X1_LOC_516/Y OR2X1_LOC_371/Y 0.03fF
C44198 OR2X1_LOC_427/A OR2X1_LOC_371/Y 0.07fF
C44238 AND2X1_LOC_464/a_8_24# OR2X1_LOC_371/Y 0.02fF
C45799 OR2X1_LOC_45/B OR2X1_LOC_371/Y 0.01fF
C49041 AND2X1_LOC_840/B OR2X1_LOC_371/Y 0.19fF
C49314 AND2X1_LOC_464/A OR2X1_LOC_371/Y 0.13fF
C50233 OR2X1_LOC_56/A OR2X1_LOC_371/Y 0.07fF
C50798 OR2X1_LOC_527/Y OR2X1_LOC_371/Y 0.28fF
C55694 OR2X1_LOC_600/A OR2X1_LOC_371/Y 0.07fF
C56538 OR2X1_LOC_371/Y VSS 0.51fF
C30018 OR2X1_LOC_57/Y AND2X1_LOC_198/a_8_24# 0.23fF
C35431 VDD OR2X1_LOC_57/Y 0.12fF
C57510 OR2X1_LOC_57/Y VSS 0.06fF
C95 OR2X1_LOC_485/A OR2X1_LOC_71/Y 0.09fF
C4775 OR2X1_LOC_131/Y OR2X1_LOC_71/Y 0.43fF
C5061 VDD OR2X1_LOC_71/Y 0.53fF
C5207 OR2X1_LOC_256/A OR2X1_LOC_71/Y 0.03fF
C5242 OR2X1_LOC_71/Y OR2X1_LOC_67/Y 0.01fF
C6036 OR2X1_LOC_487/Y OR2X1_LOC_71/Y 0.01fF
C6398 OR2X1_LOC_71/Y OR2X1_LOC_427/A 0.06fF
C7350 AND2X1_LOC_557/a_8_24# OR2X1_LOC_71/Y 0.01fF
C7595 OR2X1_LOC_71/Y OR2X1_LOC_184/a_8_216# 0.08fF
C8054 OR2X1_LOC_45/B OR2X1_LOC_71/Y 0.04fF
C8551 OR2X1_LOC_158/A OR2X1_LOC_71/Y 0.05fF
C11092 OR2X1_LOC_744/A OR2X1_LOC_71/Y 0.12fF
C12311 OR2X1_LOC_118/a_8_216# OR2X1_LOC_71/Y 0.01fF
C12367 OR2X1_LOC_71/Y OR2X1_LOC_56/A 0.02fF
C12875 OR2X1_LOC_91/Y OR2X1_LOC_71/Y 0.03fF
C14634 OR2X1_LOC_246/A OR2X1_LOC_71/Y 0.02fF
C15015 OR2X1_LOC_497/Y OR2X1_LOC_71/Y 0.03fF
C15249 OR2X1_LOC_71/Y AND2X1_LOC_249/a_8_24# 0.01fF
C16250 OR2X1_LOC_71/Y AND2X1_LOC_361/A 0.28fF
C17502 OR2X1_LOC_71/Y OR2X1_LOC_65/B 0.08fF
C17835 OR2X1_LOC_600/A OR2X1_LOC_71/Y 0.03fF
C18893 OR2X1_LOC_813/A OR2X1_LOC_71/Y 0.35fF
C20278 OR2X1_LOC_71/Y OR2X1_LOC_13/B 0.03fF
C20490 OR2X1_LOC_71/Y AND2X1_LOC_266/a_8_24# 0.01fF
C20810 OR2X1_LOC_71/Y OR2X1_LOC_428/A 0.02fF
C20833 OR2X1_LOC_71/Y OR2X1_LOC_595/A 0.04fF
C21852 OR2X1_LOC_71/Y OR2X1_LOC_89/A 0.04fF
C22759 OR2X1_LOC_488/Y OR2X1_LOC_71/Y 0.01fF
C22796 OR2X1_LOC_71/Y OR2X1_LOC_95/Y 0.31fF
C23691 OR2X1_LOC_71/Y OR2X1_LOC_71/A 0.01fF
C23982 OR2X1_LOC_70/Y OR2X1_LOC_71/Y 0.02fF
C24046 OR2X1_LOC_184/Y OR2X1_LOC_71/Y 0.09fF
C26935 AND2X1_LOC_227/Y OR2X1_LOC_71/Y 0.89fF
C27603 OR2X1_LOC_40/Y OR2X1_LOC_71/Y 0.03fF
C27722 OR2X1_LOC_71/Y OR2X1_LOC_7/A 0.06fF
C29719 OR2X1_LOC_71/Y AND2X1_LOC_489/a_8_24# 0.01fF
C29846 OR2X1_LOC_3/Y OR2X1_LOC_71/Y 0.06fF
C31083 OR2X1_LOC_503/A OR2X1_LOC_71/Y 0.02fF
C31135 OR2X1_LOC_64/Y OR2X1_LOC_71/Y 0.11fF
C32301 AND2X1_LOC_557/Y OR2X1_LOC_71/Y 0.01fF
C33546 OR2X1_LOC_494/Y OR2X1_LOC_71/Y 0.02fF
C37387 OR2X1_LOC_71/Y OR2X1_LOC_118/Y 1.95fF
C37422 OR2X1_LOC_262/Y OR2X1_LOC_71/Y 0.03fF
C38570 OR2X1_LOC_604/A OR2X1_LOC_71/Y 0.05fF
C39111 OR2X1_LOC_71/Y OR2X1_LOC_265/Y 0.01fF
C45761 OR2X1_LOC_71/Y OR2X1_LOC_437/A 0.03fF
C46954 AND2X1_LOC_489/Y OR2X1_LOC_71/Y 0.01fF
C47070 OR2X1_LOC_71/Y AND2X1_LOC_216/A 0.02fF
C47423 OR2X1_LOC_280/Y OR2X1_LOC_71/Y 0.02fF
C47815 OR2X1_LOC_71/Y OR2X1_LOC_39/A 0.23fF
C50389 OR2X1_LOC_71/Y AND2X1_LOC_266/Y 0.01fF
C51224 OR2X1_LOC_487/a_8_216# OR2X1_LOC_71/Y 0.01fF
C51511 OR2X1_LOC_71/Y OR2X1_LOC_131/a_8_216# 0.01fF
C51550 OR2X1_LOC_91/A OR2X1_LOC_71/Y 0.03fF
C52488 OR2X1_LOC_490/Y OR2X1_LOC_71/Y 0.15fF
C54392 OR2X1_LOC_106/Y OR2X1_LOC_71/Y 0.02fF
C54561 OR2X1_LOC_497/a_8_216# OR2X1_LOC_71/Y 0.01fF
C55753 AND2X1_LOC_362/B OR2X1_LOC_71/Y 0.03fF
C57076 OR2X1_LOC_71/Y VSS 0.50fF
C822 OR2X1_LOC_32/B OR2X1_LOC_69/A 0.03fF
C5059 OR2X1_LOC_81/Y OR2X1_LOC_69/A 0.01fF
C6778 OR2X1_LOC_69/A OR2X1_LOC_69/Y 0.01fF
C22923 OR2X1_LOC_600/A OR2X1_LOC_69/A 0.03fF
C30413 OR2X1_LOC_69/A OR2X1_LOC_16/A 0.03fF
C43752 OR2X1_LOC_80/Y OR2X1_LOC_69/A 0.02fF
C51957 OR2X1_LOC_69/A OR2X1_LOC_52/B 0.87fF
C52778 OR2X1_LOC_69/A OR2X1_LOC_39/A 0.03fF
C54871 OR2X1_LOC_81/a_8_216# OR2X1_LOC_69/A 0.01fF
C56645 OR2X1_LOC_69/A VSS 0.01fF
C1948 AND2X1_LOC_41/A AND2X1_LOC_65/A 0.07fF
C3493 AND2X1_LOC_31/Y AND2X1_LOC_65/A 0.02fF
C3749 OR2X1_LOC_633/B AND2X1_LOC_65/A 0.03fF
C5838 AND2X1_LOC_117/a_8_24# AND2X1_LOC_65/A 0.10fF
C8304 AND2X1_LOC_65/A OR2X1_LOC_161/B 0.03fF
C10806 AND2X1_LOC_65/A AND2X1_LOC_7/B 0.04fF
C11406 OR2X1_LOC_123/B AND2X1_LOC_65/A 0.04fF
C12539 OR2X1_LOC_160/B AND2X1_LOC_65/A 3.31fF
C21123 OR2X1_LOC_656/B AND2X1_LOC_65/A 0.53fF
C22376 AND2X1_LOC_65/A OR2X1_LOC_78/A 0.63fF
C26617 AND2X1_LOC_81/B AND2X1_LOC_65/A 0.03fF
C27826 AND2X1_LOC_65/A OR2X1_LOC_78/B 0.17fF
C27884 OR2X1_LOC_375/A AND2X1_LOC_65/A 0.07fF
C28225 AND2X1_LOC_65/A OR2X1_LOC_549/A 0.10fF
C30693 OR2X1_LOC_139/A AND2X1_LOC_65/A 0.28fF
C32082 OR2X1_LOC_87/A AND2X1_LOC_65/A 0.02fF
C33325 AND2X1_LOC_65/A OR2X1_LOC_475/B 0.40fF
C34648 OR2X1_LOC_267/A AND2X1_LOC_65/A 0.79fF
C40466 AND2X1_LOC_65/A AND2X1_LOC_265/a_8_24# 0.03fF
C40480 VDD AND2X1_LOC_65/A 0.27fF
C42431 AND2X1_LOC_667/a_8_24# AND2X1_LOC_65/A 0.03fF
C43608 OR2X1_LOC_160/A AND2X1_LOC_65/A 0.02fF
C44878 OR2X1_LOC_185/A AND2X1_LOC_65/A 0.09fF
C46131 AND2X1_LOC_65/A OR2X1_LOC_641/A 0.08fF
C47165 OR2X1_LOC_643/A AND2X1_LOC_65/A 0.07fF
C53375 AND2X1_LOC_65/A AND2X1_LOC_44/Y 0.65fF
C54224 AND2X1_LOC_65/A AND2X1_LOC_18/Y 0.05fF
C55140 OR2X1_LOC_231/A AND2X1_LOC_65/A 0.08fF
C56775 AND2X1_LOC_65/A VSS -0.95fF
C142 OR2X1_LOC_625/Y OR2X1_LOC_437/A 0.24fF
C545 OR2X1_LOC_484/Y OR2X1_LOC_437/A 0.01fF
C590 OR2X1_LOC_246/Y OR2X1_LOC_437/A 0.02fF
C947 OR2X1_LOC_16/A OR2X1_LOC_437/A 0.07fF
C987 OR2X1_LOC_108/Y OR2X1_LOC_437/A 1.05fF
C1041 AND2X1_LOC_168/Y OR2X1_LOC_437/A 0.08fF
C1876 OR2X1_LOC_109/Y OR2X1_LOC_437/A 0.10fF
C2460 AND2X1_LOC_227/Y OR2X1_LOC_437/A 0.03fF
C3134 OR2X1_LOC_40/Y OR2X1_LOC_437/A 0.60fF
C3232 OR2X1_LOC_7/A OR2X1_LOC_437/A 2.05fF
C3313 OR2X1_LOC_224/a_8_216# OR2X1_LOC_437/A 0.01fF
C4020 AND2X1_LOC_841/B OR2X1_LOC_437/A 0.07fF
C4290 AND2X1_LOC_543/Y OR2X1_LOC_437/A 0.02fF
C4331 OR2X1_LOC_437/A OR2X1_LOC_322/Y 0.19fF
C5172 AND2X1_LOC_489/a_8_24# OR2X1_LOC_437/A 0.02fF
C5263 OR2X1_LOC_3/Y OR2X1_LOC_437/A 0.09fF
C6568 OR2X1_LOC_64/Y OR2X1_LOC_437/A 0.25fF
C6774 AND2X1_LOC_247/a_8_24# OR2X1_LOC_437/A 0.01fF
C7814 OR2X1_LOC_516/B OR2X1_LOC_437/A 0.03fF
C7892 OR2X1_LOC_279/Y OR2X1_LOC_437/A 0.19fF
C8270 AND2X1_LOC_456/B OR2X1_LOC_437/A 0.04fF
C9080 OR2X1_LOC_494/Y OR2X1_LOC_437/A 0.01fF
C9988 AND2X1_LOC_624/A OR2X1_LOC_437/A 0.09fF
C12066 OR2X1_LOC_278/Y OR2X1_LOC_437/A 0.03fF
C12800 OR2X1_LOC_437/A OR2X1_LOC_142/Y 0.06fF
C13831 OR2X1_LOC_91/a_8_216# OR2X1_LOC_437/A 0.03fF
C13982 OR2X1_LOC_419/Y OR2X1_LOC_437/A 0.19fF
C14165 OR2X1_LOC_177/Y OR2X1_LOC_437/A 0.05fF
C14185 OR2X1_LOC_604/A OR2X1_LOC_437/A 0.19fF
C14550 OR2X1_LOC_176/Y OR2X1_LOC_437/A 0.02fF
C14919 OR2X1_LOC_437/A OR2X1_LOC_183/a_8_216# 0.03fF
C15399 AND2X1_LOC_326/B OR2X1_LOC_437/A 0.01fF
C15460 OR2X1_LOC_237/a_8_216# OR2X1_LOC_437/A 0.15fF
C17205 AND2X1_LOC_342/a_8_24# OR2X1_LOC_437/A 0.02fF
C17845 OR2X1_LOC_248/A OR2X1_LOC_437/A 0.01fF
C18393 OR2X1_LOC_135/Y OR2X1_LOC_437/A 0.10fF
C18474 AND2X1_LOC_848/Y OR2X1_LOC_437/A 5.95fF
C18477 AND2X1_LOC_186/a_8_24# OR2X1_LOC_437/A 0.04fF
C19295 OR2X1_LOC_256/Y OR2X1_LOC_437/A 0.03fF
C19896 OR2X1_LOC_224/Y OR2X1_LOC_437/A 0.08fF
C20591 OR2X1_LOC_165/Y OR2X1_LOC_437/A 0.02fF
C21032 OR2X1_LOC_237/a_36_216# OR2X1_LOC_437/A 0.15fF
C21434 AND2X1_LOC_715/A OR2X1_LOC_437/A 0.07fF
C21923 AND2X1_LOC_784/A OR2X1_LOC_437/A 0.16fF
C22369 OR2X1_LOC_52/B OR2X1_LOC_437/A 0.03fF
C22710 OR2X1_LOC_281/Y OR2X1_LOC_437/A 0.08fF
C22788 OR2X1_LOC_165/a_8_216# OR2X1_LOC_437/A 0.03fF
C22842 OR2X1_LOC_280/Y OR2X1_LOC_437/A 0.12fF
C23193 OR2X1_LOC_39/A OR2X1_LOC_437/A 1.74fF
C23917 OR2X1_LOC_136/Y OR2X1_LOC_437/A 0.01fF
C23978 OR2X1_LOC_51/Y OR2X1_LOC_437/A 0.17fF
C24041 OR2X1_LOC_680/A OR2X1_LOC_437/A 0.12fF
C24796 OR2X1_LOC_178/a_8_216# OR2X1_LOC_437/A 0.04fF
C24832 AND2X1_LOC_344/a_8_24# OR2X1_LOC_437/A 0.02fF
C25936 OR2X1_LOC_437/A OR2X1_LOC_183/Y 0.04fF
C26119 OR2X1_LOC_248/a_8_216# OR2X1_LOC_437/A 0.03fF
C26524 OR2X1_LOC_237/Y OR2X1_LOC_437/A 0.05fF
C26893 AND2X1_LOC_391/Y OR2X1_LOC_437/A 0.07fF
C26895 OR2X1_LOC_91/A OR2X1_LOC_437/A 0.43fF
C26963 OR2X1_LOC_669/Y OR2X1_LOC_437/A 0.07fF
C27824 OR2X1_LOC_74/A OR2X1_LOC_437/A 1.35fF
C31562 AND2X1_LOC_168/a_8_24# OR2X1_LOC_437/A 0.04fF
C31600 AND2X1_LOC_303/A OR2X1_LOC_437/A 0.01fF
C31629 OR2X1_LOC_485/A OR2X1_LOC_437/A 0.27fF
C32272 AND2X1_LOC_383/a_8_24# OR2X1_LOC_437/A 0.02fF
C34907 OR2X1_LOC_492/a_8_216# OR2X1_LOC_437/A 0.01fF
C35216 OR2X1_LOC_516/Y OR2X1_LOC_437/A 0.07fF
C35298 OR2X1_LOC_369/Y OR2X1_LOC_437/A -0.03fF
C35770 AND2X1_LOC_348/A OR2X1_LOC_437/A 0.01fF
C36568 VDD OR2X1_LOC_437/A 1.99fF
C36632 OR2X1_LOC_491/Y OR2X1_LOC_437/A 0.01fF
C36637 OR2X1_LOC_251/Y OR2X1_LOC_437/A 0.03fF
C36712 OR2X1_LOC_256/A OR2X1_LOC_437/A 0.09fF
C37064 OR2X1_LOC_248/Y OR2X1_LOC_437/A 0.36fF
C37371 AND2X1_LOC_370/a_8_24# OR2X1_LOC_437/A 0.05fF
C37520 OR2X1_LOC_487/Y OR2X1_LOC_437/A 0.01fF
C37785 OR2X1_LOC_494/A OR2X1_LOC_437/A 0.14fF
C37871 OR2X1_LOC_427/A OR2X1_LOC_437/A 0.28fF
C39531 OR2X1_LOC_45/B OR2X1_LOC_437/A 0.13fF
C39595 OR2X1_LOC_292/a_8_216# OR2X1_LOC_437/A 0.03fF
C39951 OR2X1_LOC_158/A OR2X1_LOC_437/A 0.40fF
C39979 AND2X1_LOC_98/Y OR2X1_LOC_437/A 0.02fF
C40372 OR2X1_LOC_482/Y OR2X1_LOC_437/A 0.17fF
C42584 OR2X1_LOC_309/Y OR2X1_LOC_437/A 0.01fF
C42605 OR2X1_LOC_744/A OR2X1_LOC_437/A 1.02fF
C42629 AND2X1_LOC_168/a_36_24# OR2X1_LOC_437/A 0.01fF
C42670 AND2X1_LOC_840/B OR2X1_LOC_437/A 0.05fF
C42978 AND2X1_LOC_464/A OR2X1_LOC_437/A 0.02fF
C43510 AND2X1_LOC_303/B OR2X1_LOC_437/A 0.08fF
C43890 OR2X1_LOC_56/A OR2X1_LOC_437/A 0.48fF
C44373 OR2X1_LOC_91/Y OR2X1_LOC_437/A 0.12fF
C44765 OR2X1_LOC_494/a_8_216# OR2X1_LOC_437/A 0.03fF
C45203 AND2X1_LOC_335/a_8_24# OR2X1_LOC_437/A 0.04fF
C45627 OR2X1_LOC_484/a_8_216# OR2X1_LOC_437/A 0.01fF
C45719 OR2X1_LOC_481/A OR2X1_LOC_437/A 0.03fF
C46038 OR2X1_LOC_492/Y OR2X1_LOC_437/A 0.02fF
C46195 OR2X1_LOC_246/A OR2X1_LOC_437/A 0.10fF
C46587 OR2X1_LOC_497/Y OR2X1_LOC_437/A 0.19fF
C47640 AND2X1_LOC_721/A OR2X1_LOC_437/A 0.24fF
C48654 AND2X1_LOC_787/A OR2X1_LOC_437/A 0.58fF
C49554 OR2X1_LOC_600/A OR2X1_LOC_437/A 0.62fF
C50048 OR2X1_LOC_669/A OR2X1_LOC_437/A 0.11fF
C50849 OR2X1_LOC_292/Y OR2X1_LOC_437/A 0.02fF
C51744 OR2X1_LOC_312/Y OR2X1_LOC_437/A 0.10fF
C51938 OR2X1_LOC_13/B OR2X1_LOC_437/A 0.49fF
C52376 OR2X1_LOC_437/A OR2X1_LOC_142/a_8_216# 0.01fF
C52449 OR2X1_LOC_428/A OR2X1_LOC_437/A 0.38fF
C52911 OR2X1_LOC_528/Y OR2X1_LOC_437/A 0.06fF
C52979 OR2X1_LOC_516/A OR2X1_LOC_437/A 0.12fF
C52983 AND2X1_LOC_342/Y OR2X1_LOC_437/A 0.08fF
C53430 OR2X1_LOC_89/A OR2X1_LOC_437/A 0.22fF
C54099 AND2X1_LOC_287/B OR2X1_LOC_437/A 0.09fF
C54142 OR2X1_LOC_491/a_8_216# OR2X1_LOC_437/A 0.02fF
C54257 OR2X1_LOC_488/Y OR2X1_LOC_437/A 0.05fF
C54280 AND2X1_LOC_727/A OR2X1_LOC_437/A 0.03fF
C54314 OR2X1_LOC_95/Y OR2X1_LOC_437/A 0.34fF
C55050 AND2X1_LOC_621/Y OR2X1_LOC_437/A 0.07fF
C55541 OR2X1_LOC_70/Y OR2X1_LOC_437/A 0.07fF
C55643 OR2X1_LOC_437/Y OR2X1_LOC_437/A 0.12fF
C56379 OR2X1_LOC_437/A VSS -8.26fF
C2193 OR2X1_LOC_821/Y OR2X1_LOC_86/A 0.01fF
C3186 OR2X1_LOC_70/Y OR2X1_LOC_86/A 0.50fF
C6164 OR2X1_LOC_813/Y OR2X1_LOC_86/A 0.02fF
C6944 OR2X1_LOC_86/A OR2X1_LOC_7/A 0.05fF
C10428 OR2X1_LOC_64/Y OR2X1_LOC_86/A 0.10fF
C10804 AND2X1_LOC_101/B OR2X1_LOC_86/A 0.16fF
C15818 OR2X1_LOC_86/A OR2X1_LOC_278/Y 0.01fF
C26189 OR2X1_LOC_86/A AND2X1_LOC_216/A 0.20fF
C40536 OR2X1_LOC_86/A OR2X1_LOC_67/Y 0.01fF
C47332 OR2X1_LOC_821/a_8_216# OR2X1_LOC_86/A 0.39fF
C50052 OR2X1_LOC_246/A OR2X1_LOC_86/A 0.03fF
C51192 OR2X1_LOC_235/B OR2X1_LOC_86/A 0.04fF
C54238 OR2X1_LOC_813/A OR2X1_LOC_86/A 0.37fF
C55667 OR2X1_LOC_86/A OR2X1_LOC_13/B 0.08fF
C56971 OR2X1_LOC_86/A VSS 0.42fF
C42 OR2X1_LOC_246/A OR2X1_LOC_595/a_8_216# 0.11fF
C517 OR2X1_LOC_485/A OR2X1_LOC_246/A 0.03fF
C5461 VDD OR2X1_LOC_246/A 1.15fF
C5670 OR2X1_LOC_246/A OR2X1_LOC_67/Y 0.07fF
C7358 OR2X1_LOC_246/A OR2X1_LOC_416/Y 0.01fF
C8493 OR2X1_LOC_45/B OR2X1_LOC_246/A 0.01fF
C8638 OR2X1_LOC_246/A OR2X1_LOC_767/a_8_216# 0.16fF
C8932 OR2X1_LOC_158/A OR2X1_LOC_246/A 0.10fF
C11132 OR2X1_LOC_316/Y OR2X1_LOC_246/A 0.03fF
C11507 OR2X1_LOC_744/A OR2X1_LOC_246/A 0.02fF
C12783 OR2X1_LOC_246/A OR2X1_LOC_56/A 0.01fF
C13319 OR2X1_LOC_305/Y OR2X1_LOC_246/A 0.02fF
C14149 OR2X1_LOC_246/A OR2X1_LOC_767/a_36_216# 0.15fF
C16656 OR2X1_LOC_246/A AND2X1_LOC_361/A 0.03fF
C17914 OR2X1_LOC_246/A OR2X1_LOC_65/B 0.03fF
C18361 OR2X1_LOC_246/A OR2X1_LOC_619/Y 0.01fF
C20692 OR2X1_LOC_246/A OR2X1_LOC_13/B 0.18fF
C21238 OR2X1_LOC_246/A OR2X1_LOC_595/A 0.31fF
C22270 OR2X1_LOC_246/A OR2X1_LOC_89/A 0.55fF
C23395 OR2X1_LOC_821/Y OR2X1_LOC_246/A 0.03fF
C24094 OR2X1_LOC_246/A OR2X1_LOC_71/A 0.47fF
C24371 OR2X1_LOC_70/Y OR2X1_LOC_246/A 0.02fF
C25583 OR2X1_LOC_246/Y OR2X1_LOC_246/A 0.02fF
C27352 AND2X1_LOC_227/Y OR2X1_LOC_246/A 0.10fF
C27374 OR2X1_LOC_246/A OR2X1_LOC_813/Y 0.12fF
C28022 OR2X1_LOC_40/Y OR2X1_LOC_246/A 0.01fF
C29252 OR2X1_LOC_589/A OR2X1_LOC_246/A 0.27fF
C30254 OR2X1_LOC_3/Y OR2X1_LOC_246/A 0.26fF
C31536 OR2X1_LOC_64/Y OR2X1_LOC_246/A 0.03fF
C35710 AND2X1_LOC_777/a_8_24# OR2X1_LOC_246/A 0.10fF
C36904 OR2X1_LOC_246/A OR2X1_LOC_278/Y 0.03fF
C36981 OR2X1_LOC_273/Y OR2X1_LOC_246/A 0.01fF
C37779 OR2X1_LOC_246/A OR2X1_LOC_118/Y 0.02fF
C40212 OR2X1_LOC_131/A OR2X1_LOC_246/A 1.22fF
C41328 OR2X1_LOC_246/A OR2X1_LOC_595/Y 0.51fF
C42587 OR2X1_LOC_272/Y OR2X1_LOC_246/A 0.03fF
C43264 OR2X1_LOC_135/Y OR2X1_LOC_246/A 0.10fF
C46925 AND2X1_LOC_784/A OR2X1_LOC_246/A 0.30fF
C47404 OR2X1_LOC_246/A OR2X1_LOC_52/B 0.10fF
C48248 OR2X1_LOC_246/A OR2X1_LOC_39/A 0.10fF
C48914 OR2X1_LOC_136/Y OR2X1_LOC_246/A 0.10fF
C51911 OR2X1_LOC_246/A OR2X1_LOC_131/a_8_216# 0.18fF
C51954 OR2X1_LOC_91/A OR2X1_LOC_246/A 0.14fF
C52915 OR2X1_LOC_246/A OR2X1_LOC_74/A 0.13fF
C54424 AND2X1_LOC_339/B OR2X1_LOC_246/A 0.03fF
C54716 OR2X1_LOC_246/A OR2X1_LOC_300/Y 0.03fF
C57100 OR2X1_LOC_246/A VSS 0.99fF
C2262 OR2X1_LOC_3/Y OR2X1_LOC_278/A 0.01fF
C8653 OR2X1_LOC_278/A OR2X1_LOC_612/B 0.05fF
C9216 OR2X1_LOC_278/A AND2X1_LOC_608/a_8_24# 0.01fF
C9882 OR2X1_LOC_278/A OR2X1_LOC_118/Y 0.38fF
C12042 OR2X1_LOC_278/A AND2X1_LOC_633/Y 0.02fF
C20073 OR2X1_LOC_278/A OR2X1_LOC_39/A 0.32fF
C22258 OR2X1_LOC_278/A OR2X1_LOC_609/A 0.07fF
C24782 OR2X1_LOC_278/A OR2X1_LOC_74/A 0.04fF
C25243 OR2X1_LOC_278/A OR2X1_LOC_607/Y 0.11fF
C26395 OR2X1_LOC_278/A AND2X1_LOC_633/a_8_24# 0.07fF
C33510 VDD OR2X1_LOC_278/A 0.19fF
C33718 OR2X1_LOC_278/A OR2X1_LOC_67/Y 0.79fF
C36375 OR2X1_LOC_45/B OR2X1_LOC_278/A 0.15fF
C39450 OR2X1_LOC_744/A OR2X1_LOC_278/A 0.15fF
C41255 OR2X1_LOC_291/Y OR2X1_LOC_278/A 0.83fF
C46455 OR2X1_LOC_278/A OR2X1_LOC_619/Y 3.79fF
C52161 OR2X1_LOC_278/A OR2X1_LOC_71/A 0.01fF
C56176 OR2X1_LOC_40/Y OR2X1_LOC_278/A 0.07fF
C57142 OR2X1_LOC_278/A VSS 0.40fF
C523 OR2X1_LOC_117/Y OR2X1_LOC_256/A 0.07fF
C2198 OR2X1_LOC_744/A OR2X1_LOC_256/A 0.03fF
C6990 OR2X1_LOC_256/A AND2X1_LOC_721/A 0.04fF
C7338 OR2X1_LOC_256/A AND2X1_LOC_361/A 0.02fF
C8654 OR2X1_LOC_256/A OR2X1_LOC_65/B 0.02fF
C11343 OR2X1_LOC_256/A OR2X1_LOC_13/B 0.04fF
C11893 OR2X1_LOC_256/A OR2X1_LOC_595/A 0.02fF
C12451 AND2X1_LOC_342/Y OR2X1_LOC_256/A 0.33fF
C12911 OR2X1_LOC_256/A OR2X1_LOC_89/A 0.05fF
C13818 OR2X1_LOC_256/A OR2X1_LOC_95/Y 9.35fF
C17042 OR2X1_LOC_132/Y OR2X1_LOC_256/A 0.08fF
C18062 OR2X1_LOC_256/A OR2X1_LOC_813/Y 0.03fF
C18861 OR2X1_LOC_256/A OR2X1_LOC_7/A 0.32fF
C20995 OR2X1_LOC_3/Y OR2X1_LOC_256/A 0.03fF
C22309 OR2X1_LOC_64/Y OR2X1_LOC_256/A 0.03fF
C22546 AND2X1_LOC_541/a_8_24# OR2X1_LOC_256/A 0.09fF
C27689 OR2X1_LOC_256/A OR2X1_LOC_278/Y 0.03fF
C28550 OR2X1_LOC_256/A OR2X1_LOC_118/Y 0.03fF
C33232 OR2X1_LOC_272/Y OR2X1_LOC_256/A 0.01fF
C34859 OR2X1_LOC_256/Y OR2X1_LOC_256/A 0.07fF
C39478 OR2X1_LOC_51/Y OR2X1_LOC_256/A 0.07fF
C42498 AND2X1_LOC_391/Y OR2X1_LOC_256/A 0.72fF
C43441 OR2X1_LOC_490/Y OR2X1_LOC_256/A 0.07fF
C46019 AND2X1_LOC_99/A OR2X1_LOC_256/A 0.03fF
C47436 OR2X1_LOC_485/A OR2X1_LOC_256/A 0.42fF
C52387 VDD OR2X1_LOC_256/A 0.21fF
C52582 OR2X1_LOC_256/A OR2X1_LOC_67/Y 0.14fF
C52918 OR2X1_LOC_256/A OR2X1_LOC_248/Y 0.09fF
C55763 OR2X1_LOC_158/A OR2X1_LOC_256/A 0.01fF
C57144 OR2X1_LOC_256/A VSS -0.09fF
C1376 OR2X1_LOC_690/A OR2X1_LOC_27/a_8_216# 0.01fF
C7701 OR2X1_LOC_690/A OR2X1_LOC_52/B 0.06fF
C8586 OR2X1_LOC_690/A OR2X1_LOC_39/A 0.11fF
C12426 OR2X1_LOC_690/A OR2X1_LOC_27/Y 0.03fF
C12799 OR2X1_LOC_32/B OR2X1_LOC_690/A 0.01fF
C16932 OR2X1_LOC_58/Y OR2X1_LOC_690/A 0.01fF
C18697 OR2X1_LOC_290/a_8_216# OR2X1_LOC_690/A 0.01fF
C19037 OR2X1_LOC_690/A OR2X1_LOC_13/Y 0.02fF
C22081 VDD OR2X1_LOC_690/A 0.68fF
C23941 OR2X1_LOC_416/Y OR2X1_LOC_690/A 0.02fF
C25395 OR2X1_LOC_158/A OR2X1_LOC_690/A 0.04fF
C29226 OR2X1_LOC_690/A OR2X1_LOC_56/A 0.03fF
C29692 OR2X1_LOC_290/Y OR2X1_LOC_690/A 0.23fF
C32254 OR2X1_LOC_690/A OR2X1_LOC_24/a_8_216# 0.11fF
C32298 OR2X1_LOC_7/a_8_216# OR2X1_LOC_690/A 0.14fF
C34689 OR2X1_LOC_600/A OR2X1_LOC_690/A 0.03fF
C42327 OR2X1_LOC_690/A OR2X1_LOC_16/A 0.06fF
C43373 OR2X1_LOC_690/A OR2X1_LOC_24/a_36_216# 0.03fF
C43398 AND2X1_LOC_729/B OR2X1_LOC_690/A 0.01fF
C44678 OR2X1_LOC_7/A OR2X1_LOC_690/A 0.03fF
C45110 OR2X1_LOC_32/a_8_216# OR2X1_LOC_690/A 0.40fF
C46893 OR2X1_LOC_3/Y OR2X1_LOC_690/A 0.16fF
C46985 AND2X1_LOC_462/B OR2X1_LOC_690/A 0.01fF
C49086 OR2X1_LOC_7/Y OR2X1_LOC_690/A 0.60fF
C54964 OR2X1_LOC_52/Y OR2X1_LOC_690/A 0.02fF
C56862 OR2X1_LOC_690/A VSS 0.76fF
C9824 VDD OR2X1_LOC_813/A 0.12fF
C10003 OR2X1_LOC_813/A OR2X1_LOC_67/Y 0.01fF
C15723 OR2X1_LOC_744/A OR2X1_LOC_813/A 0.03fF
C20465 OR2X1_LOC_235/B OR2X1_LOC_813/A 0.04fF
C25148 OR2X1_LOC_813/A AND2X1_LOC_266/a_8_24# 0.11fF
C28307 OR2X1_LOC_813/A OR2X1_LOC_71/A 0.14fF
C35751 OR2X1_LOC_813/A OR2X1_LOC_64/Y 0.03fF
C42096 OR2X1_LOC_813/A OR2X1_LOC_118/Y 0.02fF
C54976 OR2X1_LOC_813/A AND2X1_LOC_266/Y 0.02fF
C57306 OR2X1_LOC_813/A VSS 0.44fF
C1784 AND2X1_LOC_36/Y OR2X1_LOC_622/B 0.05fF
C19293 OR2X1_LOC_622/A OR2X1_LOC_622/B 0.16fF
C29973 OR2X1_LOC_622/a_8_216# OR2X1_LOC_622/B 0.47fF
C56470 OR2X1_LOC_622/B VSS 0.16fF
C8475 OR2X1_LOC_96/Y OR2X1_LOC_672/Y 0.02fF
C12390 OR2X1_LOC_670/Y OR2X1_LOC_672/Y 0.08fF
C15204 OR2X1_LOC_604/A OR2X1_LOC_672/Y 0.07fF
C37637 VDD OR2X1_LOC_672/Y 0.19fF
C41022 OR2X1_LOC_158/A OR2X1_LOC_672/Y 0.01fF
C44997 OR2X1_LOC_672/Y OR2X1_LOC_56/A 0.01fF
C47084 OR2X1_LOC_672/Y AND2X1_LOC_789/Y 0.02fF
C53522 OR2X1_LOC_672/Y OR2X1_LOC_428/A 0.01fF
C55441 OR2X1_LOC_672/Y OR2X1_LOC_95/Y 0.01fF
C57116 OR2X1_LOC_672/Y VSS 0.26fF
C4648 VDD OR2X1_LOC_68/Y 0.16fF
C9030 OR2X1_LOC_185/A OR2X1_LOC_68/Y 0.01fF
C11397 AND2X1_LOC_91/B OR2X1_LOC_68/Y 0.19fF
C18884 OR2X1_LOC_68/Y AND2X1_LOC_69/a_8_24# 0.23fF
C21447 OR2X1_LOC_68/Y AND2X1_LOC_51/Y 0.01fF
C23655 OR2X1_LOC_68/Y AND2X1_LOC_31/Y 0.02fF
C24538 OR2X1_LOC_68/Y AND2X1_LOC_36/Y 0.11fF
C47415 OR2X1_LOC_574/A OR2X1_LOC_68/Y 0.09fF
C52463 OR2X1_LOC_68/Y OR2X1_LOC_87/A 0.01fF
C57248 OR2X1_LOC_68/Y VSS 0.07fF
C8361 AND2X1_LOC_57/Y OR2X1_LOC_154/A 0.03fF
C8579 AND2X1_LOC_57/Y OR2X1_LOC_198/A 0.17fF
C30858 AND2X1_LOC_57/Y AND2X1_LOC_51/Y 0.09fF
C31592 AND2X1_LOC_57/Y AND2X1_LOC_41/A 0.06fF
C37800 AND2X1_LOC_57/Y OR2X1_LOC_198/a_8_216# 0.05fF
C58097 AND2X1_LOC_57/Y VSS 0.22fF
C2383 OR2X1_LOC_335/A OR2X1_LOC_161/A 0.04fF
C7928 OR2X1_LOC_335/A OR2X1_LOC_269/B 0.14fF
C13515 OR2X1_LOC_335/A OR2X1_LOC_76/A 0.03fF
C23710 OR2X1_LOC_335/A OR2X1_LOC_605/A 0.26fF
C24674 OR2X1_LOC_335/A OR2X1_LOC_318/B 0.02fF
C29092 OR2X1_LOC_335/A OR2X1_LOC_375/A 0.01fF
C29154 OR2X1_LOC_335/A OR2X1_LOC_605/B 0.11fF
C33323 OR2X1_LOC_335/A OR2X1_LOC_87/A 0.01fF
C35619 OR2X1_LOC_335/A OR2X1_LOC_590/a_8_216# 0.01fF
C35862 OR2X1_LOC_335/A OR2X1_LOC_154/A 0.01fF
C36753 OR2X1_LOC_335/A OR2X1_LOC_335/B 0.42fF
C37368 OR2X1_LOC_335/A OR2X1_LOC_590/Y 0.01fF
C42958 OR2X1_LOC_335/A AND2X1_LOC_591/a_8_24# 0.01fF
C46161 OR2X1_LOC_335/A OR2X1_LOC_185/A 0.71fF
C54107 OR2X1_LOC_335/A OR2X1_LOC_593/B 1.48fF
C58110 OR2X1_LOC_335/A VSS 0.05fF
C853 AND2X1_LOC_72/B AND2X1_LOC_248/a_8_24# 0.01fF
C7608 AND2X1_LOC_72/B OR2X1_LOC_844/B 0.84fF
C9950 OR2X1_LOC_154/A AND2X1_LOC_72/B 0.03fF
C11930 AND2X1_LOC_72/B OR2X1_LOC_342/A 0.01fF
C13845 OR2X1_LOC_532/B AND2X1_LOC_72/B 0.02fF
C15760 VDD AND2X1_LOC_72/B 0.48fF
C17804 AND2X1_LOC_72/B OR2X1_LOC_115/B 0.26fF
C18864 OR2X1_LOC_160/A AND2X1_LOC_72/B 0.08fF
C19337 AND2X1_LOC_127/a_8_24# AND2X1_LOC_72/B 0.01fF
C21342 AND2X1_LOC_72/B OR2X1_LOC_294/Y 1.19fF
C22595 AND2X1_LOC_91/B AND2X1_LOC_72/B 0.03fF
C23066 AND2X1_LOC_72/B OR2X1_LOC_719/B 0.03fF
C24458 AND2X1_LOC_47/Y AND2X1_LOC_72/B 0.04fF
C26798 AND2X1_LOC_72/B AND2X1_LOC_295/a_8_24# 0.01fF
C28477 AND2X1_LOC_72/B AND2X1_LOC_44/Y 0.02fF
C29133 OR2X1_LOC_247/Y AND2X1_LOC_72/B 0.02fF
C29353 AND2X1_LOC_72/B AND2X1_LOC_18/Y 0.02fF
C30293 AND2X1_LOC_292/a_8_24# AND2X1_LOC_72/B 0.01fF
C30669 OR2X1_LOC_128/A AND2X1_LOC_72/B 0.01fF
C32242 AND2X1_LOC_72/B OR2X1_LOC_346/A 0.01fF
C32323 AND2X1_LOC_72/B OR2X1_LOC_161/A 1.29fF
C32786 AND2X1_LOC_72/B AND2X1_LOC_297/a_8_24# 0.10fF
C33240 OR2X1_LOC_631/B AND2X1_LOC_72/B 0.05fF
C35759 OR2X1_LOC_346/B AND2X1_LOC_72/B 0.01fF
C38265 AND2X1_LOC_72/B OR2X1_LOC_347/B 0.01fF
C38944 AND2X1_LOC_72/B OR2X1_LOC_777/B 0.03fF
C39470 AND2X1_LOC_72/B OR2X1_LOC_161/B 0.03fF
C40846 AND2X1_LOC_72/a_8_24# AND2X1_LOC_72/B 0.11fF
C42175 OR2X1_LOC_296/Y AND2X1_LOC_72/B 0.35fF
C43825 OR2X1_LOC_160/B AND2X1_LOC_72/B 0.03fF
C44662 OR2X1_LOC_151/A AND2X1_LOC_72/B 1.33fF
C46646 AND2X1_LOC_72/B AND2X1_LOC_497/a_8_24# 0.04fF
C47865 OR2X1_LOC_664/Y AND2X1_LOC_72/B 0.03fF
C53740 AND2X1_LOC_72/B OR2X1_LOC_78/A 0.03fF
C54545 OR2X1_LOC_501/B AND2X1_LOC_72/B 0.03fF
C54940 OR2X1_LOC_114/B AND2X1_LOC_72/B 0.01fF
C56853 AND2X1_LOC_72/B VSS 0.28fF
C8671 AND2X1_LOC_31/Y OR2X1_LOC_778/B 0.42fF
C12980 OR2X1_LOC_831/B OR2X1_LOC_778/B 0.08fF
C17641 OR2X1_LOC_160/B OR2X1_LOC_778/B 0.03fF
C39844 OR2X1_LOC_778/A OR2X1_LOC_778/B 0.01fF
C43788 OR2X1_LOC_532/B OR2X1_LOC_778/B 0.01fF
C44875 OR2X1_LOC_778/B OR2X1_LOC_778/a_8_216# 0.03fF
C45732 VDD OR2X1_LOC_778/B 0.05fF
C50538 OR2X1_LOC_778/B OR2X1_LOC_778/a_36_216# 0.01fF
C52313 OR2X1_LOC_778/Y OR2X1_LOC_778/B 0.86fF
C54490 AND2X1_LOC_47/Y OR2X1_LOC_778/B 0.03fF
C56568 OR2X1_LOC_778/B VSS 0.18fF
C1098 OR2X1_LOC_134/Y OR2X1_LOC_65/B 0.14fF
C2105 AND2X1_LOC_99/A OR2X1_LOC_65/B 0.06fF
C2309 OR2X1_LOC_65/B OR2X1_LOC_72/Y 0.02fF
C3456 OR2X1_LOC_485/A OR2X1_LOC_65/B 0.09fF
C7030 OR2X1_LOC_117/a_8_216# OR2X1_LOC_65/B 0.02fF
C8137 OR2X1_LOC_131/Y OR2X1_LOC_65/B 0.15fF
C8451 VDD OR2X1_LOC_65/B 0.79fF
C8691 OR2X1_LOC_65/B OR2X1_LOC_67/Y 0.05fF
C11097 OR2X1_LOC_65/B AND2X1_LOC_116/Y 0.01fF
C11308 OR2X1_LOC_45/B OR2X1_LOC_65/B 0.13fF
C12592 OR2X1_LOC_117/a_36_216# OR2X1_LOC_65/B 0.03fF
C12668 OR2X1_LOC_132/a_8_216# OR2X1_LOC_65/B 0.02fF
C13935 AND2X1_LOC_541/Y OR2X1_LOC_65/B 0.04fF
C14387 OR2X1_LOC_744/A OR2X1_LOC_65/B 0.04fF
C15610 OR2X1_LOC_65/B OR2X1_LOC_56/A 0.04fF
C18554 OR2X1_LOC_65/B AND2X1_LOC_249/a_8_24# -0.00fF
C19595 OR2X1_LOC_65/B AND2X1_LOC_361/A 0.25fF
C23613 OR2X1_LOC_65/B OR2X1_LOC_13/B 0.03fF
C23801 OR2X1_LOC_65/B AND2X1_LOC_266/a_8_24# 0.01fF
C24122 OR2X1_LOC_65/B OR2X1_LOC_595/A 0.75fF
C25120 OR2X1_LOC_89/A OR2X1_LOC_65/B 0.86fF
C26010 OR2X1_LOC_95/Y OR2X1_LOC_65/B 0.06fF
C27252 OR2X1_LOC_70/Y OR2X1_LOC_65/B 0.03fF
C30236 AND2X1_LOC_227/Y OR2X1_LOC_65/B 0.52fF
C30874 OR2X1_LOC_40/Y OR2X1_LOC_65/B 0.09fF
C31028 OR2X1_LOC_65/B OR2X1_LOC_7/A 0.03fF
C32067 OR2X1_LOC_589/A OR2X1_LOC_65/B 0.02fF
C33113 OR2X1_LOC_3/Y OR2X1_LOC_65/B 0.08fF
C34395 OR2X1_LOC_64/Y OR2X1_LOC_65/B 0.08fF
C34572 AND2X1_LOC_541/a_8_24# OR2X1_LOC_65/B -0.00fF
C40669 OR2X1_LOC_65/B OR2X1_LOC_118/Y 0.04fF
C40711 OR2X1_LOC_262/Y OR2X1_LOC_65/B 0.08fF
C41646 OR2X1_LOC_65/B OR2X1_LOC_65/a_8_216# 0.02fF
C43182 OR2X1_LOC_131/A OR2X1_LOC_65/B 0.01fF
C50298 OR2X1_LOC_65/B OR2X1_LOC_52/B 0.95fF
C50427 OR2X1_LOC_65/B AND2X1_LOC_216/A 0.02fF
C51086 OR2X1_LOC_65/B OR2X1_LOC_39/A 0.02fF
C52862 OR2X1_LOC_65/B OR2X1_LOC_65/a_36_216# 0.03fF
C53657 OR2X1_LOC_65/B AND2X1_LOC_266/Y 0.04fF
C54743 OR2X1_LOC_65/B OR2X1_LOC_131/a_8_216# 0.01fF
C54791 OR2X1_LOC_91/A OR2X1_LOC_65/B 0.03fF
C55805 OR2X1_LOC_490/Y OR2X1_LOC_65/B 0.02fF
C55808 OR2X1_LOC_74/A OR2X1_LOC_65/B 0.06fF
C56970 OR2X1_LOC_65/B VSS -0.60fF
C10779 OR2X1_LOC_464/A AND2X1_LOC_31/Y 0.03fF
C13244 OR2X1_LOC_464/A OR2X1_LOC_675/A 0.01fF
C15508 OR2X1_LOC_464/A OR2X1_LOC_161/B 0.03fF
C16521 OR2X1_LOC_464/B OR2X1_LOC_464/A 0.15fF
C19603 OR2X1_LOC_76/A OR2X1_LOC_464/A 0.03fF
C19842 OR2X1_LOC_160/B OR2X1_LOC_464/A 0.03fF
C30464 OR2X1_LOC_147/B OR2X1_LOC_464/A 0.03fF
C30657 OR2X1_LOC_464/A OR2X1_LOC_318/B 0.03fF
C41488 AND2X1_LOC_74/a_8_24# OR2X1_LOC_464/A 0.01fF
C45985 OR2X1_LOC_464/A OR2X1_LOC_532/B 0.04fF
C47204 OR2X1_LOC_76/B OR2X1_LOC_464/A 0.01fF
C50651 OR2X1_LOC_457/B OR2X1_LOC_464/A 0.03fF
C52291 OR2X1_LOC_185/A OR2X1_LOC_464/A 0.02fF
C55153 OR2X1_LOC_542/B OR2X1_LOC_464/A 0.06fF
C55284 AND2X1_LOC_56/B OR2X1_LOC_464/A 0.03fF
C55588 OR2X1_LOC_464/A OR2X1_LOC_787/B 0.02fF
C56153 OR2X1_LOC_457/a_8_216# OR2X1_LOC_464/A 0.01fF
C57158 OR2X1_LOC_464/A VSS 0.19fF
C9507 OR2X1_LOC_16/A OR2X1_LOC_300/Y 0.10fF
C12895 OR2X1_LOC_589/A OR2X1_LOC_300/Y 0.04fF
C13864 OR2X1_LOC_3/Y OR2X1_LOC_300/Y 0.03fF
C20673 OR2X1_LOC_273/Y OR2X1_LOC_300/Y 0.01fF
C25009 OR2X1_LOC_595/Y OR2X1_LOC_300/Y 0.06fF
C45184 VDD OR2X1_LOC_300/Y 0.08fF
C47109 OR2X1_LOC_416/Y OR2X1_LOC_300/Y 0.01fF
C48263 OR2X1_LOC_45/B OR2X1_LOC_300/Y 0.71fF
C50889 OR2X1_LOC_316/Y OR2X1_LOC_300/Y 0.01fF
C51641 AND2X1_LOC_301/a_8_24# OR2X1_LOC_300/Y 0.01fF
C53516 AND2X1_LOC_831/Y OR2X1_LOC_300/Y 0.02fF
C56303 OR2X1_LOC_300/Y VSS 0.27fF
C6704 OR2X1_LOC_74/A OR2X1_LOC_607/A 0.11fF
C15747 OR2X1_LOC_607/A OR2X1_LOC_67/Y 0.03fF
C41137 OR2X1_LOC_607/a_8_216# OR2X1_LOC_607/A 0.47fF
C56581 OR2X1_LOC_607/A VSS 0.15fF
C5979 OR2X1_LOC_299/Y OR2X1_LOC_52/B 0.13fF
C16186 AND2X1_LOC_302/a_8_24# OR2X1_LOC_299/Y 0.01fF
C20374 VDD OR2X1_LOC_299/Y 0.04fF
C27256 AND2X1_LOC_303/B OR2X1_LOC_299/Y 0.80fF
C27557 OR2X1_LOC_299/Y OR2X1_LOC_56/A 0.04fF
C33099 OR2X1_LOC_299/Y OR2X1_LOC_619/Y 0.03fF
C57138 OR2X1_LOC_299/Y VSS 0.08fF
C15602 AND2X1_LOC_99/A OR2X1_LOC_122/A 0.01fF
C16341 AND2X1_LOC_362/B OR2X1_LOC_122/A 0.05fF
C17663 OR2X1_LOC_122/a_8_216# OR2X1_LOC_122/A 0.47fF
C21961 VDD OR2X1_LOC_122/A -0.00fF
C29124 OR2X1_LOC_122/A OR2X1_LOC_56/A 0.04fF
C46805 OR2X1_LOC_3/Y OR2X1_LOC_122/A 0.01fF
C57517 OR2X1_LOC_122/A VSS 0.15fF
C630 OR2X1_LOC_369/Y OR2X1_LOC_309/Y 0.32fF
C7505 OR2X1_LOC_369/Y AND2X1_LOC_543/a_8_24# 0.09fF
C9767 OR2X1_LOC_369/Y OR2X1_LOC_312/Y 0.05fF
C16029 OR2X1_LOC_369/Y OR2X1_LOC_109/Y 0.01fF
C17365 OR2X1_LOC_369/Y OR2X1_LOC_7/A 0.03fF
C18511 OR2X1_LOC_369/Y OR2X1_LOC_322/Y 0.06fF
C35964 OR2X1_LOC_369/Y AND2X1_LOC_784/A 0.05fF
C41965 OR2X1_LOC_369/Y OR2X1_LOC_74/A -0.03fF
C50928 OR2X1_LOC_369/Y VDD 0.14fF
C51712 OR2X1_LOC_369/Y AND2X1_LOC_370/a_8_24# 0.09fF
C58067 OR2X1_LOC_369/Y VSS 0.14fF
C4046 OR2X1_LOC_435/A AND2X1_LOC_18/Y 0.01fF
C4905 OR2X1_LOC_130/A OR2X1_LOC_435/A 0.02fF
C5335 OR2X1_LOC_449/B OR2X1_LOC_435/A 0.14fF
C9465 AND2X1_LOC_31/Y OR2X1_LOC_435/A 0.01fF
C14277 OR2X1_LOC_435/B OR2X1_LOC_435/A 1.13fF
C16817 OR2X1_LOC_318/Y OR2X1_LOC_435/A 0.04fF
C19816 OR2X1_LOC_435/a_8_216# OR2X1_LOC_435/A 0.08fF
C26221 OR2X1_LOC_810/A OR2X1_LOC_435/A 0.03fF
C26240 AND2X1_LOC_589/a_8_24# OR2X1_LOC_435/A 0.01fF
C28249 OR2X1_LOC_78/A OR2X1_LOC_435/A 0.01fF
C32671 OR2X1_LOC_112/B OR2X1_LOC_435/A 0.43fF
C32982 OR2X1_LOC_574/A OR2X1_LOC_435/A 0.01fF
C39186 OR2X1_LOC_97/A OR2X1_LOC_435/A 0.01fF
C49695 OR2X1_LOC_160/A OR2X1_LOC_435/A 0.03fF
C50948 OR2X1_LOC_185/A OR2X1_LOC_435/A 0.17fF
C53346 AND2X1_LOC_91/B OR2X1_LOC_435/A 0.01fF
C53487 OR2X1_LOC_799/A OR2X1_LOC_435/A 0.31fF
C55304 AND2X1_LOC_47/Y OR2X1_LOC_435/A 0.04fF
C55569 OR2X1_LOC_506/A OR2X1_LOC_435/A 0.36fF
C56740 OR2X1_LOC_435/A VSS 0.21fF
C2158 OR2X1_LOC_831/B OR2X1_LOC_318/B 0.35fF
C10891 OR2X1_LOC_87/A OR2X1_LOC_831/B 0.07fF
C12087 OR2X1_LOC_541/A OR2X1_LOC_831/B 0.50fF
C13455 OR2X1_LOC_154/A OR2X1_LOC_831/B 0.32fF
C17344 OR2X1_LOC_532/B OR2X1_LOC_831/B 0.03fF
C19312 VDD OR2X1_LOC_831/B 0.25fF
C21524 OR2X1_LOC_840/A OR2X1_LOC_831/B 0.08fF
C23651 OR2X1_LOC_185/A OR2X1_LOC_831/B 0.03fF
C25755 OR2X1_LOC_778/Y OR2X1_LOC_831/B 0.07fF
C27971 AND2X1_LOC_47/Y OR2X1_LOC_831/B 5.64fF
C31478 OR2X1_LOC_831/B OR2X1_LOC_593/B 0.01fF
C32823 OR2X1_LOC_831/B AND2X1_LOC_18/Y 0.03fF
C35924 AND2X1_LOC_51/Y OR2X1_LOC_831/B 0.08fF
C36275 OR2X1_LOC_831/a_8_216# OR2X1_LOC_831/B 0.05fF
C36627 AND2X1_LOC_41/A OR2X1_LOC_831/B 0.03fF
C38161 AND2X1_LOC_31/Y OR2X1_LOC_831/B 0.03fF
C39102 OR2X1_LOC_831/B AND2X1_LOC_36/Y 0.16fF
C45621 OR2X1_LOC_831/B AND2X1_LOC_7/B 0.02fF
C47471 OR2X1_LOC_160/B OR2X1_LOC_831/B 0.01fF
C53645 OR2X1_LOC_831/B OR2X1_LOC_241/B 0.01fF
C54187 OR2X1_LOC_831/A OR2X1_LOC_831/B 0.34fF
C56776 OR2X1_LOC_831/B VSS 0.50fF
C374 OR2X1_LOC_637/a_8_216# OR2X1_LOC_828/B 0.01fF
C6677 OR2X1_LOC_769/A OR2X1_LOC_828/B 0.15fF
C9207 OR2X1_LOC_828/B OR2X1_LOC_828/Y 1.00fF
C14721 OR2X1_LOC_828/B AND2X1_LOC_829/a_8_24# 0.01fF
C20259 OR2X1_LOC_828/B OR2X1_LOC_855/A 0.01fF
C23357 OR2X1_LOC_769/B OR2X1_LOC_828/B 0.01fF
C23777 OR2X1_LOC_637/Y OR2X1_LOC_828/B 0.01fF
C27762 OR2X1_LOC_828/B OR2X1_LOC_198/A 0.25fF
C33407 VDD OR2X1_LOC_828/B 0.11fF
C36433 OR2X1_LOC_160/A OR2X1_LOC_828/B 0.03fF
C40703 AND2X1_LOC_56/B OR2X1_LOC_828/B 0.03fF
C42407 OR2X1_LOC_828/a_8_216# OR2X1_LOC_828/B 0.03fF
C50349 OR2X1_LOC_828/B AND2X1_LOC_51/Y 0.04fF
C51857 AND2X1_LOC_764/a_8_24# OR2X1_LOC_828/B 0.01fF
C52525 OR2X1_LOC_828/B AND2X1_LOC_31/Y 0.03fF
C56975 OR2X1_LOC_828/B VSS 0.25fF
C2265 OR2X1_LOC_87/A OR2X1_LOC_780/B 0.01fF
C3479 AND2X1_LOC_744/a_8_24# OR2X1_LOC_780/B 0.27fF
C10679 VDD OR2X1_LOC_780/B 0.21fF
C13729 OR2X1_LOC_160/A OR2X1_LOC_780/B 0.15fF
C14537 OR2X1_LOC_780/B AND2X1_LOC_424/a_8_24# 0.04fF
C19753 OR2X1_LOC_780/A OR2X1_LOC_780/B 0.04fF
C23405 OR2X1_LOC_780/B AND2X1_LOC_44/Y 0.32fF
C25571 OR2X1_LOC_780/B AND2X1_LOC_424/a_36_24# 0.01fF
C25625 OR2X1_LOC_780/B OR2X1_LOC_449/B 0.09fF
C30725 OR2X1_LOC_780/B OR2X1_LOC_780/a_8_216# 0.02fF
C34297 OR2X1_LOC_780/B OR2X1_LOC_161/B 0.23fF
C37883 OR2X1_LOC_446/Y OR2X1_LOC_780/B 0.11fF
C38586 OR2X1_LOC_160/B OR2X1_LOC_780/B 0.11fF
C48606 OR2X1_LOC_780/B OR2X1_LOC_78/A 0.02fF
C57040 OR2X1_LOC_780/B VSS 0.36fF
C12236 OR2X1_LOC_156/A OR2X1_LOC_87/A 0.13fF
C14771 OR2X1_LOC_156/A OR2X1_LOC_154/A 0.14fF
C23720 OR2X1_LOC_156/A OR2X1_LOC_160/A 0.30fF
C40449 OR2X1_LOC_154/a_8_216# OR2X1_LOC_156/A 0.41fF
C47005 OR2X1_LOC_156/A AND2X1_LOC_7/B 0.35fF
C48774 OR2X1_LOC_156/A OR2X1_LOC_160/B 0.22fF
C51706 OR2X1_LOC_156/B OR2X1_LOC_156/A 0.15fF
C58060 OR2X1_LOC_156/A VSS 0.29fF
C179 OR2X1_LOC_608/a_8_216# OR2X1_LOC_502/Y 0.39fF
C200 OR2X1_LOC_185/A OR2X1_LOC_502/Y 0.22fF
C33708 OR2X1_LOC_78/A OR2X1_LOC_502/Y 0.02fF
C37943 AND2X1_LOC_81/B OR2X1_LOC_502/Y 0.01fF
C39199 OR2X1_LOC_78/B OR2X1_LOC_502/Y 0.01fF
C52087 VDD OR2X1_LOC_502/Y 0.08fF
C56349 OR2X1_LOC_502/Y VSS 0.22fF
C5764 OR2X1_LOC_708/B AND2X1_LOC_44/Y 0.03fF
C6618 OR2X1_LOC_708/B OR2X1_LOC_708/a_8_216# 0.03fF
C9826 OR2X1_LOC_708/B OR2X1_LOC_161/A 0.10fF
C12072 OR2X1_LOC_708/B AND2X1_LOC_31/Y 0.03fF
C12205 OR2X1_LOC_708/B OR2X1_LOC_708/a_36_216# 0.01fF
C28302 OR2X1_LOC_710/A OR2X1_LOC_708/B 0.82fF
C30947 OR2X1_LOC_708/B OR2X1_LOC_78/A 0.34fF
C43344 OR2X1_LOC_154/A OR2X1_LOC_708/B 0.14fF
C46218 OR2X1_LOC_708/B OR2X1_LOC_779/A 0.01fF
C49353 VDD OR2X1_LOC_708/B 0.02fF
C57063 OR2X1_LOC_708/B VSS 0.13fF
C465 OR2X1_LOC_512/A AND2X1_LOC_47/Y 0.01fF
C2720 OR2X1_LOC_512/A OR2X1_LOC_779/B 0.01fF
C4441 OR2X1_LOC_512/A AND2X1_LOC_44/Y 0.01fF
C5725 OR2X1_LOC_512/A OR2X1_LOC_307/A 0.25fF
C9276 OR2X1_LOC_512/A AND2X1_LOC_41/A 0.04fF
C10783 OR2X1_LOC_512/A AND2X1_LOC_31/Y 0.01fF
C12997 OR2X1_LOC_308/A OR2X1_LOC_512/A 0.47fF
C14050 OR2X1_LOC_512/A OR2X1_LOC_269/B 0.01fF
C15513 OR2X1_LOC_512/A OR2X1_LOC_161/B 0.01fF
C19848 OR2X1_LOC_512/A OR2X1_LOC_160/B 0.18fF
C27586 OR2X1_LOC_307/a_8_216# OR2X1_LOC_512/A 0.48fF
C29580 OR2X1_LOC_512/A OR2X1_LOC_78/A 0.01fF
C35133 OR2X1_LOC_512/A OR2X1_LOC_375/A 0.04fF
C40920 OR2X1_LOC_512/A OR2X1_LOC_713/A 0.02fF
C48858 OR2X1_LOC_512/A OR2X1_LOC_834/A 0.22fF
C54781 OR2X1_LOC_512/A OR2X1_LOC_308/a_8_216# 0.07fF
C57871 OR2X1_LOC_512/A VSS 0.38fF
C10659 OR2X1_LOC_147/A AND2X1_LOC_51/Y 0.01fF
C11340 OR2X1_LOC_147/A AND2X1_LOC_41/A 0.15fF
C16091 OR2X1_LOC_147/A OR2X1_LOC_269/B 0.24fF
C18832 OR2X1_LOC_147/A OR2X1_LOC_705/B 0.21fF
C20217 OR2X1_LOC_147/A AND2X1_LOC_7/B 0.03fF
C29043 OR2X1_LOC_710/A OR2X1_LOC_147/A 0.09fF
C32548 OR2X1_LOC_147/B OR2X1_LOC_147/A 0.06fF
C37213 OR2X1_LOC_147/A OR2X1_LOC_375/A 0.01fF
C43435 OR2X1_LOC_147/A OR2X1_LOC_546/A 0.21fF
C44111 OR2X1_LOC_154/A OR2X1_LOC_147/A 0.13fF
C49232 OR2X1_LOC_710/B OR2X1_LOC_147/A 0.04fF
C53134 OR2X1_LOC_160/A OR2X1_LOC_147/A 0.05fF
C57443 OR2X1_LOC_147/A VSS 0.04fF
C11835 OR2X1_LOC_168/B AND2X1_LOC_601/a_8_24# 0.20fF
C12371 OR2X1_LOC_168/B OR2X1_LOC_168/A 0.04fF
C13054 OR2X1_LOC_841/A OR2X1_LOC_168/B 0.01fF
C17268 OR2X1_LOC_168/B OR2X1_LOC_78/A 0.02fF
C18666 OR2X1_LOC_841/B OR2X1_LOC_168/B 0.03fF
C19881 OR2X1_LOC_168/B OR2X1_LOC_776/a_8_216# 0.01fF
C22123 OR2X1_LOC_168/B OR2X1_LOC_574/A 0.17fF
C22889 OR2X1_LOC_168/B OR2X1_LOC_78/B 0.19fF
C28241 OR2X1_LOC_97/A OR2X1_LOC_168/B 0.17fF
C35423 VDD OR2X1_LOC_168/B 0.30fF
C37580 OR2X1_LOC_840/A OR2X1_LOC_168/B 0.03fF
C41474 OR2X1_LOC_168/a_8_216# OR2X1_LOC_168/B 0.07fF
C42192 AND2X1_LOC_91/B OR2X1_LOC_168/B 0.13fF
C44234 OR2X1_LOC_168/B AND2X1_LOC_47/Y 0.01fF
C44512 OR2X1_LOC_168/B OR2X1_LOC_506/A 0.19fF
C47469 OR2X1_LOC_168/B OR2X1_LOC_776/A 0.08fF
C47886 OR2X1_LOC_168/B OR2X1_LOC_593/B 0.03fF
C50644 OR2X1_LOC_168/B OR2X1_LOC_449/B 0.02fF
C52359 OR2X1_LOC_168/B AND2X1_LOC_51/Y 2.24fF
C52720 OR2X1_LOC_831/a_8_216# OR2X1_LOC_168/B 0.07fF
C54573 OR2X1_LOC_168/B AND2X1_LOC_31/Y 0.08fF
C55478 OR2X1_LOC_168/B AND2X1_LOC_36/Y 0.10fF
C57577 OR2X1_LOC_168/B VSS 0.25fF
C13456 OR2X1_LOC_325/B OR2X1_LOC_538/A 0.04fF
C16317 OR2X1_LOC_186/Y OR2X1_LOC_325/B 1.76fF
C22057 OR2X1_LOC_325/B OR2X1_LOC_87/A 0.03fF
C23189 OR2X1_LOC_97/A OR2X1_LOC_325/B 0.12fF
C30364 VDD OR2X1_LOC_325/B 0.02fF
C33673 OR2X1_LOC_325/B OR2X1_LOC_532/Y 0.06fF
C33786 OR2X1_LOC_325/A OR2X1_LOC_325/B 0.56fF
C37425 OR2X1_LOC_325/B OR2X1_LOC_303/B 0.03fF
C39040 OR2X1_LOC_325/B AND2X1_LOC_47/Y 0.09fF
C39593 OR2X1_LOC_325/B OR2X1_LOC_180/B 0.03fF
C41390 OR2X1_LOC_325/B OR2X1_LOC_703/A 0.05fF
C47928 OR2X1_LOC_325/B OR2X1_LOC_439/B 0.03fF
C50539 OR2X1_LOC_325/a_8_216# OR2X1_LOC_325/B 0.47fF
C54213 OR2X1_LOC_325/B OR2X1_LOC_161/B 0.01fF
C57662 OR2X1_LOC_325/B VSS 0.49fF
C19562 OR2X1_LOC_459/B OR2X1_LOC_459/a_8_216# 0.02fF
C20414 OR2X1_LOC_459/B OR2X1_LOC_375/A 0.03fF
C24592 OR2X1_LOC_459/A OR2X1_LOC_459/B 0.15fF
C30536 OR2X1_LOC_459/B OR2X1_LOC_463/B 0.01fF
C57119 OR2X1_LOC_459/B VSS 0.14fF
C6571 OR2X1_LOC_638/B VDD 0.21fF
C13487 OR2X1_LOC_638/B OR2X1_LOC_638/a_8_216# 0.05fF
C25618 OR2X1_LOC_638/B AND2X1_LOC_31/Y 0.03fF
C50179 OR2X1_LOC_638/B OR2X1_LOC_375/A 0.02fF
C53071 OR2X1_LOC_638/B OR2X1_LOC_637/Y 0.17fF
C57865 OR2X1_LOC_638/B VSS 0.22fF
C21396 OR2X1_LOC_837/B OR2X1_LOC_416/A 0.43fF
C26877 OR2X1_LOC_416/A OR2X1_LOC_52/B 0.25fF
C44619 OR2X1_LOC_158/A OR2X1_LOC_416/A 0.04fF
C57060 OR2X1_LOC_416/A VSS 0.31fF
C14003 OR2X1_LOC_585/Y AND2X1_LOC_637/Y 0.82fF
C20247 VDD OR2X1_LOC_585/Y -0.00fF
C24151 OR2X1_LOC_585/Y OR2X1_LOC_586/Y 0.02fF
C29754 OR2X1_LOC_409/B OR2X1_LOC_585/Y 0.01fF
C45012 OR2X1_LOC_3/Y OR2X1_LOC_585/Y 0.10fF
C55560 OR2X1_LOC_585/Y AND2X1_LOC_637/a_8_24# 0.02fF
C56690 OR2X1_LOC_585/Y VSS 0.02fF
C64 OR2X1_LOC_485/A OR2X1_LOC_481/A 0.01fF
C2279 OR2X1_LOC_481/A OR2X1_LOC_295/Y 0.01fF
C4243 AND2X1_LOC_348/A OR2X1_LOC_481/A 0.02fF
C5010 VDD OR2X1_LOC_481/A 0.36fF
C5926 OR2X1_LOC_382/Y OR2X1_LOC_481/A 0.41fF
C6214 OR2X1_LOC_494/A OR2X1_LOC_481/A 0.31fF
C6346 OR2X1_LOC_481/A OR2X1_LOC_427/A 0.11fF
C8498 OR2X1_LOC_158/A OR2X1_LOC_481/A 0.06fF
C9028 OR2X1_LOC_748/A OR2X1_LOC_481/A 0.06fF
C9990 OR2X1_LOC_481/A AND2X1_LOC_848/A 0.03fF
C11227 OR2X1_LOC_481/A OR2X1_LOC_257/Y 0.01fF
C12323 OR2X1_LOC_481/A OR2X1_LOC_56/A 0.20fF
C13227 OR2X1_LOC_494/a_8_216# OR2X1_LOC_481/A 0.47fF
C14305 OR2X1_LOC_481/A AND2X1_LOC_789/Y 0.07fF
C17447 OR2X1_LOC_481/A OR2X1_LOC_257/a_8_216# 0.01fF
C17775 OR2X1_LOC_600/A OR2X1_LOC_481/A 0.03fF
C19147 OR2X1_LOC_292/Y OR2X1_LOC_481/A 0.02fF
C20758 OR2X1_LOC_481/A OR2X1_LOC_428/A 0.06fF
C21821 OR2X1_LOC_481/A OR2X1_LOC_89/A 0.06fF
C24721 OR2X1_LOC_481/A OR2X1_LOC_625/Y 0.02fF
C27541 OR2X1_LOC_40/Y OR2X1_LOC_481/A 0.06fF
C29812 OR2X1_LOC_3/Y OR2X1_LOC_481/A 0.16fF
C36150 OR2X1_LOC_481/A OR2X1_LOC_295/a_8_216# 0.19fF
C38515 OR2X1_LOC_604/A OR2X1_LOC_481/A 0.24fF
C39829 AND2X1_LOC_711/A OR2X1_LOC_481/A 0.08fF
C42930 OR2X1_LOC_481/A AND2X1_LOC_848/Y 0.03fF
C43763 OR2X1_LOC_256/Y OR2X1_LOC_481/A 0.01fF
C43860 OR2X1_LOC_481/A OR2X1_LOC_258/Y 0.02fF
C51316 OR2X1_LOC_481/A OR2X1_LOC_384/Y 0.04fF
C51504 OR2X1_LOC_481/A OR2X1_LOC_91/A 2.00fF
C54494 OR2X1_LOC_481/A AND2X1_LOC_847/Y 0.01fF
C57374 OR2X1_LOC_481/A VSS -0.16fF
C424 OR2X1_LOC_625/Y OR2X1_LOC_754/a_8_216# 0.02fF
C2907 OR2X1_LOC_51/Y OR2X1_LOC_625/Y 0.12fF
C3580 OR2X1_LOC_625/Y AND2X1_LOC_790/a_8_24# 0.06fF
C3775 AND2X1_LOC_344/a_8_24# OR2X1_LOC_625/Y 0.02fF
C5039 OR2X1_LOC_625/Y OR2X1_LOC_248/a_8_216# -0.00fF
C8143 OR2X1_LOC_625/Y OR2X1_LOC_615/a_8_216# 0.01fF
C9253 OR2X1_LOC_625/Y AND2X1_LOC_614/a_8_24# 0.06fF
C10649 OR2X1_LOC_625/Y OR2X1_LOC_248/a_36_216# 0.03fF
C10666 OR2X1_LOC_665/Y OR2X1_LOC_625/Y 0.03fF
C10678 OR2X1_LOC_485/A OR2X1_LOC_625/Y 0.11fF
C11513 OR2X1_LOC_625/Y OR2X1_LOC_754/a_36_216# 0.01fF
C13685 OR2X1_LOC_625/Y OR2X1_LOC_615/a_36_216# 0.01fF
C14627 OR2X1_LOC_625/Y AND2X1_LOC_793/B -0.02fF
C14822 AND2X1_LOC_348/A OR2X1_LOC_625/Y 0.02fF
C15587 VDD OR2X1_LOC_625/Y 1.30fF
C16130 OR2X1_LOC_625/Y OR2X1_LOC_248/Y 0.22fF
C16805 OR2X1_LOC_494/A OR2X1_LOC_625/Y 0.01fF
C16967 OR2X1_LOC_625/Y OR2X1_LOC_427/A 0.28fF
C18976 OR2X1_LOC_158/A OR2X1_LOC_625/Y 0.03fF
C19425 OR2X1_LOC_482/Y OR2X1_LOC_625/Y 0.21fF
C19650 OR2X1_LOC_625/Y OR2X1_LOC_628/Y 0.11fF
C21632 OR2X1_LOC_744/A OR2X1_LOC_625/Y 0.99fF
C22927 OR2X1_LOC_625/Y OR2X1_LOC_56/A 0.07fF
C23306 OR2X1_LOC_625/Y AND2X1_LOC_285/Y 0.03fF
C23546 OR2X1_LOC_625/Y AND2X1_LOC_483/Y 0.04fF
C23767 OR2X1_LOC_494/a_8_216# OR2X1_LOC_625/Y 0.01fF
C26448 OR2X1_LOC_625/Y AND2X1_LOC_721/A 0.01fF
C28346 OR2X1_LOC_600/A OR2X1_LOC_625/Y 0.07fF
C30719 OR2X1_LOC_625/Y OR2X1_LOC_13/B 0.13fF
C31241 OR2X1_LOC_625/Y OR2X1_LOC_428/A 0.02fF
C31837 OR2X1_LOC_625/Y AND2X1_LOC_483/a_8_24# 0.01fF
C32224 OR2X1_LOC_625/Y OR2X1_LOC_89/A 0.09fF
C33915 OR2X1_LOC_625/Y AND2X1_LOC_621/Y 0.06fF
C34696 OR2X1_LOC_494/a_36_216# OR2X1_LOC_625/Y 0.01fF
C38145 OR2X1_LOC_625/Y OR2X1_LOC_7/A 0.30fF
C38690 OR2X1_LOC_625/Y OR2X1_LOC_615/Y 0.03fF
C40275 OR2X1_LOC_3/Y OR2X1_LOC_625/Y 0.04fF
C41640 OR2X1_LOC_625/Y OR2X1_LOC_64/Y 0.04fF
C41760 OR2X1_LOC_625/Y AND2X1_LOC_247/a_8_24# 0.02fF
C43230 AND2X1_LOC_456/B OR2X1_LOC_625/Y 0.07fF
C44059 OR2X1_LOC_494/Y OR2X1_LOC_625/Y 0.03fF
C45024 OR2X1_LOC_625/Y AND2X1_LOC_624/A 0.03fF
C47248 OR2X1_LOC_625/Y OR2X1_LOC_278/Y 0.01fF
C47766 OR2X1_LOC_625/Y OR2X1_LOC_754/A 0.19fF
C48714 OR2X1_LOC_625/Y OR2X1_LOC_754/Y 0.07fF
C49274 OR2X1_LOC_604/A OR2X1_LOC_625/Y 0.10fF
C52981 OR2X1_LOC_625/Y OR2X1_LOC_248/A 0.01fF
C53624 OR2X1_LOC_625/Y AND2X1_LOC_848/Y 0.07fF
C54382 OR2X1_LOC_256/Y OR2X1_LOC_625/Y 0.38fF
C57336 OR2X1_LOC_625/Y VSS 0.08fF
C18890 OR2X1_LOC_399/A OR2X1_LOC_399/a_8_216# 0.47fF
C51358 OR2X1_LOC_399/A OR2X1_LOC_16/A 0.11fF
C55791 OR2X1_LOC_3/Y OR2X1_LOC_399/A 0.01fF
C57730 OR2X1_LOC_399/A VSS 0.15fF
C647 OR2X1_LOC_405/Y AND2X1_LOC_7/B 0.06fF
C23272 OR2X1_LOC_97/A OR2X1_LOC_405/Y 0.01fF
C23388 OR2X1_LOC_405/Y OR2X1_LOC_475/B 0.02fF
C24666 OR2X1_LOC_154/A OR2X1_LOC_405/Y 0.01fF
C28546 OR2X1_LOC_405/Y OR2X1_LOC_532/B 0.01fF
C30443 VDD OR2X1_LOC_405/Y 0.19fF
C44064 OR2X1_LOC_405/Y AND2X1_LOC_18/Y 0.02fF
C57059 OR2X1_LOC_405/Y VSS 0.26fF
C2201 OR2X1_LOC_614/Y AND2X1_LOC_48/Y 0.01fF
C13851 AND2X1_LOC_47/Y AND2X1_LOC_48/Y 0.01fF
C25035 AND2X1_LOC_36/Y AND2X1_LOC_48/Y 0.02fF
C25356 AND2X1_LOC_48/Y OR2X1_LOC_196/a_8_216# 0.47fF
C27348 OR2X1_LOC_269/B AND2X1_LOC_48/Y 0.01fF
C42971 OR2X1_LOC_78/A AND2X1_LOC_48/Y 0.01fF
C47498 OR2X1_LOC_196/B AND2X1_LOC_48/Y 0.04fF
C56284 AND2X1_LOC_48/Y VSS 0.03fF
C362 OR2X1_LOC_706/B AND2X1_LOC_44/Y 0.01fF
C5092 AND2X1_LOC_41/A OR2X1_LOC_706/B 0.04fF
C15696 OR2X1_LOC_160/B OR2X1_LOC_706/B 0.01fF
C20379 OR2X1_LOC_706/B OR2X1_LOC_706/a_8_216# 0.47fF
C29866 OR2X1_LOC_196/B OR2X1_LOC_706/B 0.11fF
C31078 OR2X1_LOC_706/B OR2X1_LOC_375/A 0.05fF
C52536 OR2X1_LOC_706/B AND2X1_LOC_47/Y 0.05fF
C57269 OR2X1_LOC_706/B VSS 0.16fF
C6330 OR2X1_LOC_520/A OR2X1_LOC_520/a_8_216# 0.47fF
C12482 OR2X1_LOC_520/B OR2X1_LOC_520/A 0.05fF
C37718 VDD OR2X1_LOC_520/A -0.00fF
C38677 OR2X1_LOC_462/B OR2X1_LOC_520/A 0.01fF
C40768 OR2X1_LOC_160/A OR2X1_LOC_520/A 0.02fF
C57364 OR2X1_LOC_520/A VSS 0.14fF
C34 OR2X1_LOC_779/B OR2X1_LOC_713/A 0.22fF
C3237 AND2X1_LOC_677/a_8_24# OR2X1_LOC_779/B 0.01fF
C3890 OR2X1_LOC_779/B OR2X1_LOC_779/A 0.37fF
C6885 VDD OR2X1_LOC_779/B 0.21fF
C7765 OR2X1_LOC_834/A OR2X1_LOC_779/B 0.17fF
C9085 OR2X1_LOC_840/A OR2X1_LOC_779/B 0.01fF
C13397 OR2X1_LOC_778/Y OR2X1_LOC_779/B 0.17fF
C13763 OR2X1_LOC_308/a_8_216# OR2X1_LOC_779/B 0.01fF
C14010 OR2X1_LOC_446/B OR2X1_LOC_779/B 0.03fF
C15534 AND2X1_LOC_47/Y OR2X1_LOC_779/B 0.01fF
C19636 AND2X1_LOC_44/Y OR2X1_LOC_779/B 0.79fF
C20964 OR2X1_LOC_307/A OR2X1_LOC_779/B 0.35fF
C21898 OR2X1_LOC_449/B OR2X1_LOC_779/B 0.03fF
C23251 OR2X1_LOC_447/Y OR2X1_LOC_779/B 0.09fF
C23570 OR2X1_LOC_161/A OR2X1_LOC_779/B 0.01fF
C23634 AND2X1_LOC_51/Y OR2X1_LOC_779/B 0.08fF
C24365 AND2X1_LOC_41/A OR2X1_LOC_779/B 0.10fF
C25317 AND2X1_LOC_677/a_36_24# OR2X1_LOC_779/B -0.00fF
C25813 AND2X1_LOC_31/Y OR2X1_LOC_779/B 0.03fF
C29033 OR2X1_LOC_269/B OR2X1_LOC_779/B 0.03fF
C29455 OR2X1_LOC_779/a_8_216# OR2X1_LOC_779/B 0.08fF
C29835 OR2X1_LOC_678/Y OR2X1_LOC_779/B 0.01fF
C30110 OR2X1_LOC_777/B OR2X1_LOC_779/B 0.02fF
C30608 OR2X1_LOC_161/B OR2X1_LOC_779/B 0.20fF
C31892 OR2X1_LOC_777/a_8_216# OR2X1_LOC_779/B 0.01fF
C38113 OR2X1_LOC_308/Y OR2X1_LOC_779/B 0.01fF
C39153 OR2X1_LOC_448/A OR2X1_LOC_779/B 0.03fF
C42982 OR2X1_LOC_784/B OR2X1_LOC_779/B 0.01fF
C44712 OR2X1_LOC_78/A OR2X1_LOC_779/B 0.04fF
C48331 OR2X1_LOC_448/Y OR2X1_LOC_779/B -0.00fF
C50445 OR2X1_LOC_375/A OR2X1_LOC_779/B 0.84fF
C52194 OR2X1_LOC_779/Y OR2X1_LOC_779/B 0.02fF
C54160 OR2X1_LOC_834/a_8_216# OR2X1_LOC_779/B 0.01fF
C56361 OR2X1_LOC_779/B VSS 0.51fF
C4444 OR2X1_LOC_93/Y OR2X1_LOC_51/Y 0.01fF
C7475 OR2X1_LOC_93/Y OR2X1_LOC_91/A 0.12fF
C17225 VDD OR2X1_LOC_93/Y 0.12fF
C32840 OR2X1_LOC_93/Y OR2X1_LOC_428/A 0.01fF
C39649 OR2X1_LOC_40/Y OR2X1_LOC_93/Y 0.02fF
C43971 OR2X1_LOC_93/Y OR2X1_LOC_96/Y 0.08fF
C55088 OR2X1_LOC_93/Y AND2X1_LOC_98/a_8_24# 0.23fF
C57470 OR2X1_LOC_93/Y VSS 0.06fF
C3823 OR2X1_LOC_482/Y OR2X1_LOC_628/Y 0.02fF
C7222 OR2X1_LOC_628/Y OR2X1_LOC_56/A 0.09fF
C7848 OR2X1_LOC_628/Y AND2X1_LOC_483/Y 0.86fF
C15044 OR2X1_LOC_628/Y AND2X1_LOC_629/Y 0.04fF
C16105 OR2X1_LOC_528/Y OR2X1_LOC_628/Y 0.07fF
C16269 OR2X1_LOC_628/Y AND2X1_LOC_483/a_8_24# 0.01fF
C17562 OR2X1_LOC_628/Y OR2X1_LOC_95/Y 0.19fF
C18366 OR2X1_LOC_628/Y AND2X1_LOC_621/Y 0.07fF
C22583 OR2X1_LOC_40/Y OR2X1_LOC_628/Y 0.07fF
C22726 OR2X1_LOC_628/Y OR2X1_LOC_7/A 0.24fF
C23185 OR2X1_LOC_628/Y OR2X1_LOC_615/Y 0.01fF
C24800 OR2X1_LOC_628/Y AND2X1_LOC_631/Y 0.02fF
C26072 OR2X1_LOC_628/Y AND2X1_LOC_632/A 0.04fF
C27633 AND2X1_LOC_456/B OR2X1_LOC_628/Y 0.50fF
C29363 OR2X1_LOC_628/Y AND2X1_LOC_624/A 0.07fF
C42541 OR2X1_LOC_628/Y OR2X1_LOC_39/A 0.07fF
C43313 OR2X1_LOC_51/Y OR2X1_LOC_628/Y 0.02fF
C43399 OR2X1_LOC_680/A OR2X1_LOC_628/Y 0.07fF
C44686 OR2X1_LOC_252/Y OR2X1_LOC_628/Y 0.02fF
C47416 OR2X1_LOC_628/Y OR2X1_LOC_74/A 0.22fF
C49480 OR2X1_LOC_628/Y AND2X1_LOC_631/a_8_24# 0.03fF
C51209 OR2X1_LOC_665/Y OR2X1_LOC_628/Y 0.07fF
C56202 VDD OR2X1_LOC_628/Y 0.04fF
C57071 OR2X1_LOC_628/Y VSS 0.19fF
C9195 OR2X1_LOC_422/Y OR2X1_LOC_428/A 0.01fF
C9867 AND2X1_LOC_712/B OR2X1_LOC_422/Y 0.12fF
C14843 OR2X1_LOC_422/Y AND2X1_LOC_448/Y 0.80fF
C16137 OR2X1_LOC_422/Y OR2X1_LOC_7/A 0.01fF
C24929 OR2X1_LOC_422/Y OR2X1_LOC_421/Y 0.10fF
C35181 OR2X1_LOC_422/Y OR2X1_LOC_52/B 0.01fF
C41411 OR2X1_LOC_422/Y AND2X1_LOC_448/a_8_24# 0.01fF
C49708 VDD OR2X1_LOC_422/Y 0.04fF
C52600 OR2X1_LOC_45/B OR2X1_LOC_422/Y 0.01fF
C53061 OR2X1_LOC_158/A OR2X1_LOC_422/Y 0.21fF
C57320 OR2X1_LOC_422/Y VSS 0.08fF
C16097 OR2X1_LOC_838/B OR2X1_LOC_20/A 1.11fF
C21513 OR2X1_LOC_837/Y OR2X1_LOC_20/A 0.18fF
C56377 OR2X1_LOC_20/A VSS 0.18fF
C412 AND2X1_LOC_7/B OR2X1_LOC_241/B 2.12fF
C541 OR2X1_LOC_188/Y AND2X1_LOC_7/B 0.05fF
C602 OR2X1_LOC_471/B AND2X1_LOC_7/B 0.01fF
C622 AND2X1_LOC_423/a_8_24# AND2X1_LOC_7/B 0.01fF
C719 OR2X1_LOC_193/A AND2X1_LOC_7/B 0.03fF
C944 AND2X1_LOC_7/B OR2X1_LOC_339/A 0.12fF
C1107 OR2X1_LOC_537/A AND2X1_LOC_7/B 0.03fF
C1414 OR2X1_LOC_710/A AND2X1_LOC_7/B 0.13fF
C1508 AND2X1_LOC_39/a_8_24# AND2X1_LOC_7/B 0.01fF
C1945 OR2X1_LOC_610/a_8_216# AND2X1_LOC_7/B 0.16fF
C1999 OR2X1_LOC_810/A AND2X1_LOC_7/B 3.52fF
C2316 OR2X1_LOC_715/B AND2X1_LOC_7/B 0.53fF
C2320 AND2X1_LOC_626/a_8_24# AND2X1_LOC_7/B 0.04fF
C2863 OR2X1_LOC_793/A AND2X1_LOC_7/B 0.15fF
C3274 OR2X1_LOC_687/Y AND2X1_LOC_7/B 0.07fF
C4042 OR2X1_LOC_78/A AND2X1_LOC_7/B 0.27fF
C4869 OR2X1_LOC_147/B AND2X1_LOC_7/B 0.03fF
C4980 OR2X1_LOC_545/B AND2X1_LOC_7/B 0.03fF
C5198 OR2X1_LOC_121/Y AND2X1_LOC_7/B 0.01fF
C6129 OR2X1_LOC_623/B AND2X1_LOC_7/B 0.07fF
C6563 OR2X1_LOC_833/B AND2X1_LOC_7/B 1.07fF
C7039 AND2X1_LOC_32/a_8_24# AND2X1_LOC_7/B 0.01fF
C8253 AND2X1_LOC_7/B OR2X1_LOC_338/A 0.34fF
C8280 OR2X1_LOC_186/Y AND2X1_LOC_7/B 0.01fF
C8393 AND2X1_LOC_81/B AND2X1_LOC_7/B 1.22fF
C8477 OR2X1_LOC_196/B AND2X1_LOC_7/B 0.23fF
C8828 OR2X1_LOC_574/A AND2X1_LOC_7/B 0.11fF
C9107 AND2X1_LOC_7/B AND2X1_LOC_627/a_8_24# 0.10fF
C9175 AND2X1_LOC_58/a_8_24# AND2X1_LOC_7/B 0.01fF
C9193 AND2X1_LOC_16/a_8_24# AND2X1_LOC_7/B 0.01fF
C9503 AND2X1_LOC_7/B OR2X1_LOC_539/B 0.02fF
C9585 OR2X1_LOC_78/B AND2X1_LOC_7/B 0.16fF
C9644 OR2X1_LOC_375/A AND2X1_LOC_7/B 0.25fF
C9906 AND2X1_LOC_7/B OR2X1_LOC_515/Y 0.13fF
C9970 AND2X1_LOC_7/B OR2X1_LOC_549/A 0.15fF
C10871 OR2X1_LOC_181/B AND2X1_LOC_7/B 0.03fF
C11687 AND2X1_LOC_19/Y AND2X1_LOC_7/B 0.02fF
C11707 AND2X1_LOC_316/a_8_24# AND2X1_LOC_7/B 0.03fF
C12160 AND2X1_LOC_536/a_36_24# AND2X1_LOC_7/B 0.01fF
C12250 AND2X1_LOC_27/a_8_24# AND2X1_LOC_7/B 0.08fF
C12475 OR2X1_LOC_139/A AND2X1_LOC_7/B 0.07fF
C12938 AND2X1_LOC_7/B OR2X1_LOC_138/A 0.02fF
C13395 AND2X1_LOC_626/a_36_24# AND2X1_LOC_7/B 0.01fF
C13635 OR2X1_LOC_247/a_8_216# AND2X1_LOC_7/B 0.07fF
C13902 OR2X1_LOC_87/A AND2X1_LOC_7/B 0.61fF
C14587 AND2X1_LOC_7/B OR2X1_LOC_130/a_8_216# 0.05fF
C14698 OR2X1_LOC_61/B AND2X1_LOC_7/B 0.01fF
C14711 OR2X1_LOC_194/B AND2X1_LOC_7/B 0.05fF
C15040 OR2X1_LOC_97/A AND2X1_LOC_7/B 2.92fF
C15087 OR2X1_LOC_541/A AND2X1_LOC_7/B 0.08fF
C15105 AND2X1_LOC_7/B OR2X1_LOC_475/B 0.10fF
C15119 AND2X1_LOC_290/a_8_24# AND2X1_LOC_7/B 0.01fF
C15429 OR2X1_LOC_691/Y AND2X1_LOC_7/B 0.03fF
C15950 OR2X1_LOC_639/B AND2X1_LOC_7/B 0.02fF
C16007 OR2X1_LOC_333/B AND2X1_LOC_7/B 0.03fF
C16048 OR2X1_LOC_99/B AND2X1_LOC_7/B 0.02fF
C16374 OR2X1_LOC_154/A AND2X1_LOC_7/B 8.44fF
C16440 OR2X1_LOC_778/A AND2X1_LOC_7/B 0.02fF
C16580 OR2X1_LOC_99/A AND2X1_LOC_7/B 0.05fF
C17200 AND2X1_LOC_20/a_8_24# AND2X1_LOC_7/B 0.01fF
C17211 OR2X1_LOC_634/A AND2X1_LOC_7/B 0.03fF
C17552 AND2X1_LOC_7/B OR2X1_LOC_633/A 0.11fF
C18502 OR2X1_LOC_756/B AND2X1_LOC_7/B 0.28fF
C19846 OR2X1_LOC_87/B AND2X1_LOC_7/B 0.03fF
C19893 OR2X1_LOC_33/B AND2X1_LOC_7/B 0.01fF
C20370 OR2X1_LOC_532/B AND2X1_LOC_7/B 0.25fF
C20701 OR2X1_LOC_99/a_8_216# AND2X1_LOC_7/B 0.06fF
C21497 OR2X1_LOC_710/B AND2X1_LOC_7/B 0.03fF
C21540 OR2X1_LOC_547/B AND2X1_LOC_7/B 0.03fF
C21764 AND2X1_LOC_7/B OR2X1_LOC_552/A 0.06fF
C22342 VDD AND2X1_LOC_7/B 1.25fF
C22518 OR2X1_LOC_444/B AND2X1_LOC_7/B 0.13fF
C22830 OR2X1_LOC_334/B AND2X1_LOC_7/B 0.04fF
C23188 OR2X1_LOC_676/Y AND2X1_LOC_7/B 0.08fF
C23274 OR2X1_LOC_462/B AND2X1_LOC_7/B 0.03fF
C24457 OR2X1_LOC_840/A AND2X1_LOC_7/B 0.10fF
C24887 OR2X1_LOC_216/A AND2X1_LOC_7/B 0.20fF
C24930 OR2X1_LOC_457/B AND2X1_LOC_7/B 0.01fF
C24941 AND2X1_LOC_385/a_8_24# AND2X1_LOC_7/B 0.06fF
C25131 AND2X1_LOC_7/B OR2X1_LOC_750/Y 0.98fF
C25336 OR2X1_LOC_160/A AND2X1_LOC_7/B 5.29fF
C26569 OR2X1_LOC_185/A AND2X1_LOC_7/B 0.08fF
C27074 OR2X1_LOC_702/A AND2X1_LOC_7/B 0.01fF
C28283 AND2X1_LOC_7/B OR2X1_LOC_541/B 0.08fF
C28721 OR2X1_LOC_778/Y AND2X1_LOC_7/B 0.03fF
C28995 AND2X1_LOC_91/B AND2X1_LOC_7/B 0.16fF
C29101 AND2X1_LOC_72/Y AND2X1_LOC_7/B 0.02fF
C29357 AND2X1_LOC_7/B OR2X1_LOC_446/B 0.09fF
C29457 AND2X1_LOC_7/B OR2X1_LOC_719/B 0.02fF
C29480 OR2X1_LOC_542/B AND2X1_LOC_7/B 0.03fF
C29559 AND2X1_LOC_56/B AND2X1_LOC_7/B 12.81fF
C30424 OR2X1_LOC_389/B AND2X1_LOC_7/B 0.03fF
C30593 AND2X1_LOC_7/B AND2X1_LOC_751/a_8_24# 0.04fF
C30954 AND2X1_LOC_47/Y AND2X1_LOC_7/B 8.39fF
C31231 OR2X1_LOC_506/A AND2X1_LOC_7/B 0.15fF
C31650 OR2X1_LOC_633/Y AND2X1_LOC_7/B 0.03fF
C31893 AND2X1_LOC_7/B AND2X1_LOC_41/Y 0.03fF
C34025 AND2X1_LOC_7/B OR2X1_LOC_771/B 0.05fF
C34042 AND2X1_LOC_7/B OR2X1_LOC_776/A 0.01fF
C34865 AND2X1_LOC_7/B OR2X1_LOC_317/B 0.06fF
C34944 AND2X1_LOC_7/B AND2X1_LOC_44/Y 0.70fF
C35792 AND2X1_LOC_7/B AND2X1_LOC_18/Y 0.37fF
C35845 OR2X1_LOC_473/a_8_216# AND2X1_LOC_7/B 0.03fF
C36085 AND2X1_LOC_7/B OR2X1_LOC_789/A 0.03fF
C36635 AND2X1_LOC_65/a_8_24# AND2X1_LOC_7/B 0.01fF
C36656 OR2X1_LOC_231/A AND2X1_LOC_7/B 0.13fF
C36672 OR2X1_LOC_447/a_8_216# AND2X1_LOC_7/B 0.01fF
C36679 OR2X1_LOC_130/A AND2X1_LOC_7/B 0.17fF
C36699 AND2X1_LOC_7/a_8_24# AND2X1_LOC_7/B 0.01fF
C36846 AND2X1_LOC_7/B AND2X1_LOC_39/Y 0.01fF
C37137 OR2X1_LOC_449/B AND2X1_LOC_7/B 0.07fF
C38506 OR2X1_LOC_447/Y AND2X1_LOC_7/B 0.32fF
C38746 OR2X1_LOC_709/B AND2X1_LOC_7/B 0.11fF
C38835 OR2X1_LOC_161/A AND2X1_LOC_7/B 0.29fF
C38919 AND2X1_LOC_51/Y AND2X1_LOC_7/B 0.34fF
C39261 AND2X1_LOC_7/B OR2X1_LOC_541/a_8_216# 0.02fF
C39641 AND2X1_LOC_41/A AND2X1_LOC_7/B 18.11fF
C39718 OR2X1_LOC_631/B AND2X1_LOC_7/B 0.03fF
C39996 AND2X1_LOC_524/a_8_24# AND2X1_LOC_7/B 0.03fF
C41172 AND2X1_LOC_31/Y AND2X1_LOC_7/B 0.18fF
C41354 OR2X1_LOC_473/a_36_216# AND2X1_LOC_7/B 0.02fF
C41641 AND2X1_LOC_7/B AND2X1_LOC_751/a_36_24# 0.01fF
C42022 AND2X1_LOC_7/B OR2X1_LOC_451/B 0.08fF
C42112 AND2X1_LOC_7/B AND2X1_LOC_36/Y 11.29fF
C42135 AND2X1_LOC_7/B OR2X1_LOC_334/A 0.21fF
C42157 OR2X1_LOC_154/a_8_216# AND2X1_LOC_7/B 0.06fF
C42208 AND2X1_LOC_368/a_8_24# AND2X1_LOC_7/B 0.01fF
C42211 OR2X1_LOC_633/a_8_216# AND2X1_LOC_7/B 0.47fF
C43072 AND2X1_LOC_313/a_8_24# AND2X1_LOC_7/B 0.01fF
C43452 AND2X1_LOC_60/a_8_24# AND2X1_LOC_7/B 0.01fF
C44012 AND2X1_LOC_584/a_8_24# AND2X1_LOC_7/B -0.00fF
C44460 AND2X1_LOC_7/B OR2X1_LOC_269/B 0.99fF
C44796 AND2X1_LOC_172/a_8_24# AND2X1_LOC_7/B 0.01fF
C45257 OR2X1_LOC_678/Y AND2X1_LOC_7/B 0.01fF
C45572 AND2X1_LOC_7/B OR2X1_LOC_777/B 0.09fF
C45625 OR2X1_LOC_188/a_8_216# AND2X1_LOC_7/B -0.04fF
C45644 AND2X1_LOC_7/B OR2X1_LOC_344/A 0.04fF
C45722 OR2X1_LOC_493/A AND2X1_LOC_7/B 0.98fF
C45800 AND2X1_LOC_13/a_8_24# AND2X1_LOC_7/B 0.08fF
C46087 AND2X1_LOC_7/B OR2X1_LOC_161/B 0.64fF
C46174 AND2X1_LOC_536/a_8_24# AND2X1_LOC_7/B 0.04fF
C46459 AND2X1_LOC_7/B AND2X1_LOC_406/a_8_24# 0.02fF
C46716 AND2X1_LOC_67/Y AND2X1_LOC_7/B 0.18fF
C47556 AND2X1_LOC_230/a_8_24# AND2X1_LOC_7/B 0.09fF
C47938 OR2X1_LOC_201/A AND2X1_LOC_7/B 0.01fF
C48024 AND2X1_LOC_7/a_36_24# AND2X1_LOC_7/B 0.01fF
C48041 OR2X1_LOC_647/B AND2X1_LOC_7/B 0.07fF
C48862 OR2X1_LOC_296/Y AND2X1_LOC_7/B 0.01fF
C49836 OR2X1_LOC_473/A AND2X1_LOC_7/B 0.05fF
C49904 AND2X1_LOC_7/B OR2X1_LOC_513/Y 0.01fF
C50455 OR2X1_LOC_160/B AND2X1_LOC_7/B 0.96fF
C50519 AND2X1_LOC_7/B OR2X1_LOC_553/A 0.11fF
C51255 OR2X1_LOC_151/A AND2X1_LOC_7/B 0.07fF
C51297 AND2X1_LOC_67/a_8_24# AND2X1_LOC_7/B 0.04fF
C51586 AND2X1_LOC_7/B OR2X1_LOC_714/A 0.01fF
C51739 OR2X1_LOC_174/A AND2X1_LOC_7/B 0.01fF
C51759 AND2X1_LOC_482/a_8_24# AND2X1_LOC_7/B 0.04fF
C53760 AND2X1_LOC_7/B OR2X1_LOC_308/Y 0.09fF
C53909 AND2X1_LOC_516/a_8_24# AND2X1_LOC_7/B 0.01fF
C54518 AND2X1_LOC_7/B OR2X1_LOC_181/A 0.11fF
C54610 OR2X1_LOC_61/A AND2X1_LOC_7/B 0.01fF
C54821 AND2X1_LOC_7/Y AND2X1_LOC_7/B 0.03fF
C55031 AND2X1_LOC_7/B OR2X1_LOC_390/A 0.03fF
C55481 OR2X1_LOC_711/B AND2X1_LOC_7/B 0.12fF
C56643 AND2X1_LOC_7/B VSS -5.59fF
C1280 OR2X1_LOC_256/Y OR2X1_LOC_7/A 0.04fF
C3430 OR2X1_LOC_3/Y OR2X1_LOC_256/Y 0.03fF
C4813 OR2X1_LOC_256/Y AND2X1_LOC_247/a_8_24# 0.01fF
C6208 AND2X1_LOC_456/B OR2X1_LOC_256/Y 0.23fF
C7050 OR2X1_LOC_494/Y OR2X1_LOC_256/Y 0.01fF
C15867 OR2X1_LOC_256/Y OR2X1_LOC_248/A 0.01fF
C22009 OR2X1_LOC_256/Y OR2X1_LOC_51/Y 0.12fF
C22932 OR2X1_LOC_256/Y AND2X1_LOC_344/a_8_24# 0.05fF
C24241 OR2X1_LOC_256/Y OR2X1_LOC_248/a_8_216# 0.02fF
C24956 AND2X1_LOC_391/Y OR2X1_LOC_256/Y 0.07fF
C29703 OR2X1_LOC_256/Y OR2X1_LOC_485/A 0.01fF
C33849 OR2X1_LOC_256/Y AND2X1_LOC_348/A 0.01fF
C34607 VDD OR2X1_LOC_256/Y 0.35fF
C35155 OR2X1_LOC_256/Y OR2X1_LOC_248/Y 0.52fF
C37947 OR2X1_LOC_158/A OR2X1_LOC_256/Y 0.10fF
C40556 OR2X1_LOC_256/Y OR2X1_LOC_744/A 0.07fF
C41869 OR2X1_LOC_256/Y OR2X1_LOC_56/A 0.03fF
C42773 OR2X1_LOC_256/Y OR2X1_LOC_494/a_8_216# 0.01fF
C45587 OR2X1_LOC_256/Y AND2X1_LOC_721/A 0.01fF
C47575 OR2X1_LOC_256/Y OR2X1_LOC_600/A 0.03fF
C50016 OR2X1_LOC_256/Y OR2X1_LOC_13/B 0.04fF
C51046 OR2X1_LOC_256/Y AND2X1_LOC_342/Y 0.05fF
C57666 OR2X1_LOC_256/Y VSS -0.17fF
C908 OR2X1_LOC_756/B AND2X1_LOC_47/Y 0.17fF
C1075 OR2X1_LOC_756/B OR2X1_LOC_34/A 0.01fF
C1215 OR2X1_LOC_756/B OR2X1_LOC_506/A 0.03fF
C1468 OR2X1_LOC_756/B OR2X1_LOC_180/B 0.06fF
C1957 OR2X1_LOC_756/B OR2X1_LOC_621/A 0.07fF
C2206 OR2X1_LOC_756/B OR2X1_LOC_434/A 0.01fF
C2972 AND2X1_LOC_393/a_8_24# OR2X1_LOC_756/B 0.02fF
C3315 OR2X1_LOC_756/B OR2X1_LOC_703/A 0.03fF
C3368 OR2X1_LOC_791/B OR2X1_LOC_756/B 0.03fF
C3673 OR2X1_LOC_756/B OR2X1_LOC_362/A 0.04fF
C4008 OR2X1_LOC_756/B OR2X1_LOC_771/B 0.14fF
C4859 OR2X1_LOC_756/B AND2X1_LOC_44/Y 0.07fF
C5377 OR2X1_LOC_756/B OR2X1_LOC_260/Y 0.07fF
C5727 OR2X1_LOC_756/B AND2X1_LOC_18/Y 0.59fF
C6703 OR2X1_LOC_756/B OR2X1_LOC_130/A 0.04fF
C6973 OR2X1_LOC_549/a_8_216# OR2X1_LOC_756/B 0.01fF
C7129 OR2X1_LOC_756/B AND2X1_LOC_487/a_8_24# 0.01fF
C7171 OR2X1_LOC_756/B OR2X1_LOC_449/B 0.03fF
C8519 OR2X1_LOC_400/B OR2X1_LOC_756/B 0.03fF
C8589 OR2X1_LOC_756/B AND2X1_LOC_442/a_36_24# 0.01fF
C8885 OR2X1_LOC_756/B OR2X1_LOC_161/A 0.18fF
C8973 OR2X1_LOC_756/B AND2X1_LOC_51/Y 0.87fF
C9681 OR2X1_LOC_756/B AND2X1_LOC_41/A 0.18fF
C10037 OR2X1_LOC_756/B AND2X1_LOC_524/a_8_24# 0.18fF
C10523 OR2X1_LOC_756/Y OR2X1_LOC_756/B 0.02fF
C10993 OR2X1_LOC_756/B OR2X1_LOC_593/a_8_216# 0.01fF
C11173 OR2X1_LOC_756/B AND2X1_LOC_31/Y 0.16fF
C11946 OR2X1_LOC_756/B OR2X1_LOC_288/A 0.01fF
C12062 OR2X1_LOC_756/B AND2X1_LOC_36/Y 0.26fF
C12080 OR2X1_LOC_756/B OR2X1_LOC_333/a_8_216# 0.02fF
C12086 OR2X1_LOC_756/B OR2X1_LOC_334/A 0.01fF
C12732 OR2X1_LOC_756/B OR2X1_LOC_592/a_8_216# 0.01fF
C13621 OR2X1_LOC_756/B OR2X1_LOC_557/A 0.06fF
C13967 OR2X1_LOC_756/B OR2X1_LOC_814/Y 0.02fF
C14441 OR2X1_LOC_756/B OR2X1_LOC_269/B 0.05fF
C14890 OR2X1_LOC_756/B AND2X1_LOC_176/a_8_24# 0.13fF
C15438 OR2X1_LOC_756/B OR2X1_LOC_777/B 0.05fF
C15520 OR2X1_LOC_756/B OR2X1_LOC_545/A 0.13fF
C15922 OR2X1_LOC_756/B OR2X1_LOC_161/B 0.55fF
C16002 OR2X1_LOC_756/B OR2X1_LOC_435/B 0.09fF
C17356 OR2X1_LOC_400/A OR2X1_LOC_756/B 0.01fF
C17614 OR2X1_LOC_756/B OR2X1_LOC_489/A 0.01fF
C18298 OR2X1_LOC_756/B OR2X1_LOC_401/A 0.01fF
C18614 OR2X1_LOC_318/Y OR2X1_LOC_756/B 0.03fF
C18745 OR2X1_LOC_756/B OR2X1_LOC_436/a_8_216# 0.01fF
C19618 OR2X1_LOC_756/B AND2X1_LOC_165/a_8_24# 0.01fF
C19992 OR2X1_LOC_756/B OR2X1_LOC_287/B 0.09fF
C20063 OR2X1_LOC_756/B OR2X1_LOC_436/Y 0.01fF
C20263 OR2X1_LOC_756/B OR2X1_LOC_160/B 0.24fF
C20359 OR2X1_LOC_756/B OR2X1_LOC_553/A 0.03fF
C21093 OR2X1_LOC_756/B OR2X1_LOC_151/A 0.29fF
C21582 OR2X1_LOC_756/B OR2X1_LOC_287/A 0.26fF
C21602 OR2X1_LOC_756/B OR2X1_LOC_174/A 0.26fF
C21609 OR2X1_LOC_756/B OR2X1_LOC_435/a_8_216# 0.01fF
C22422 OR2X1_LOC_756/B AND2X1_LOC_616/a_8_24# 0.03fF
C22532 OR2X1_LOC_756/B AND2X1_LOC_251/a_8_24# 0.02fF
C22609 OR2X1_LOC_756/B OR2X1_LOC_285/B 0.01fF
C22806 OR2X1_LOC_756/B OR2X1_LOC_168/Y 0.34fF
C23211 OR2X1_LOC_756/B OR2X1_LOC_334/a_8_216# 0.02fF
C23748 OR2X1_LOC_756/B AND2X1_LOC_125/a_8_24# 0.11fF
C23830 OR2X1_LOC_756/B OR2X1_LOC_593/A 0.01fF
C24521 OR2X1_LOC_756/B AND2X1_LOC_24/a_8_24# 0.01fF
C24898 OR2X1_LOC_756/B OR2X1_LOC_390/A 0.05fF
C25126 OR2X1_LOC_756/B OR2X1_LOC_168/A 0.01fF
C25517 OR2X1_LOC_756/B AND2X1_LOC_816/a_8_24# 0.01fF
C25979 OR2X1_LOC_756/B OR2X1_LOC_84/A -0.00fF
C26177 OR2X1_LOC_756/B OR2X1_LOC_190/A 0.03fF
C26540 OR2X1_LOC_188/Y OR2X1_LOC_756/B 0.02fF
C26924 OR2X1_LOC_756/B OR2X1_LOC_339/A 0.24fF
C26977 OR2X1_LOC_756/B AND2X1_LOC_438/a_8_24# 0.01fF
C27058 OR2X1_LOC_335/Y OR2X1_LOC_756/B 0.02fF
C27079 OR2X1_LOC_791/A OR2X1_LOC_756/B 0.12fF
C28008 OR2X1_LOC_756/B OR2X1_LOC_810/A 0.08fF
C28026 OR2X1_LOC_756/B AND2X1_LOC_589/a_8_24# 0.01fF
C28280 OR2X1_LOC_715/B OR2X1_LOC_756/B 0.01fF
C28631 OR2X1_LOC_756/B OR2X1_LOC_338/B 0.01fF
C28788 AND2X1_LOC_767/a_8_24# OR2X1_LOC_756/B 0.01fF
C29922 AND2X1_LOC_91/a_8_24# OR2X1_LOC_756/B 0.01fF
C29996 OR2X1_LOC_756/B OR2X1_LOC_78/A 0.33fF
C30891 OR2X1_LOC_756/B OR2X1_LOC_147/B 0.03fF
C30971 OR2X1_LOC_756/B AND2X1_LOC_171/a_8_24# 0.01fF
C30977 OR2X1_LOC_756/B OR2X1_LOC_843/a_8_216# 0.02fF
C31042 OR2X1_LOC_756/B OR2X1_LOC_545/B 0.02fF
C31257 OR2X1_LOC_756/B AND2X1_LOC_396/a_8_24# 0.01fF
C31886 OR2X1_LOC_756/B OR2X1_LOC_549/Y 0.01fF
C32256 OR2X1_LOC_756/B OR2X1_LOC_544/A 0.01fF
C32532 OR2X1_LOC_756/B OR2X1_LOC_434/a_8_216# 0.01fF
C33515 OR2X1_LOC_756/B OR2X1_LOC_592/A 0.02fF
C34127 OR2X1_LOC_756/B OR2X1_LOC_338/A 0.70fF
C34259 OR2X1_LOC_773/B OR2X1_LOC_756/B 0.01fF
C34411 OR2X1_LOC_756/B OR2X1_LOC_112/B 0.02fF
C34751 OR2X1_LOC_756/B OR2X1_LOC_574/A 0.03fF
C34760 OR2X1_LOC_756/B OR2X1_LOC_33/A 0.01fF
C35335 OR2X1_LOC_756/B OR2X1_LOC_539/B 0.02fF
C35460 OR2X1_LOC_756/B OR2X1_LOC_78/B 0.81fF
C35553 OR2X1_LOC_756/B OR2X1_LOC_375/A 0.28fF
C35850 OR2X1_LOC_756/B OR2X1_LOC_843/B 0.04fF
C36479 OR2X1_LOC_756/B OR2X1_LOC_846/A 0.01fF
C36572 OR2X1_LOC_756/B OR2X1_LOC_348/B 0.09fF
C36758 OR2X1_LOC_756/B OR2X1_LOC_181/B 0.02fF
C36854 OR2X1_LOC_756/B AND2X1_LOC_261/a_8_24# 0.19fF
C37665 OR2X1_LOC_756/B OR2X1_LOC_673/Y 0.01fF
C38150 OR2X1_LOC_756/B AND2X1_LOC_27/a_8_24# 0.01fF
C38339 OR2X1_LOC_756/B OR2X1_LOC_139/A 0.03fF
C38409 OR2X1_LOC_756/B AND2X1_LOC_179/a_8_24# 0.14fF
C39667 AND2X1_LOC_594/a_8_24# OR2X1_LOC_756/B 0.01fF
C39805 OR2X1_LOC_703/B OR2X1_LOC_756/B 0.02fF
C39820 OR2X1_LOC_756/B OR2X1_LOC_87/A 0.03fF
C39856 OR2X1_LOC_756/B AND2X1_LOC_815/a_8_24# 0.01fF
C40201 OR2X1_LOC_756/B OR2X1_LOC_403/B 0.01fF
C40762 OR2X1_LOC_756/B AND2X1_LOC_250/a_8_24# 0.02fF
C40843 OR2X1_LOC_756/B OR2X1_LOC_349/B 0.20fF
C40886 OR2X1_LOC_97/A OR2X1_LOC_756/B 0.01fF
C41066 OR2X1_LOC_756/B AND2X1_LOC_282/a_8_24# 0.02fF
C41988 OR2X1_LOC_756/B OR2X1_LOC_333/B 0.04fF
C41995 OR2X1_LOC_756/B OR2X1_LOC_850/A 0.03fF
C42403 OR2X1_LOC_154/A OR2X1_LOC_756/B 0.05fF
C42478 OR2X1_LOC_756/B OR2X1_LOC_345/A 0.08fF
C42833 AND2X1_LOC_395/a_8_24# OR2X1_LOC_756/B 0.05fF
C43185 OR2X1_LOC_756/B OR2X1_LOC_634/A 0.02fF
C43542 OR2X1_LOC_756/B OR2X1_LOC_756/a_8_216# 0.09fF
C43776 OR2X1_LOC_756/B OR2X1_LOC_34/B 0.01fF
C43983 OR2X1_LOC_756/B AND2X1_LOC_82/Y 0.01fF
C44222 OR2X1_LOC_756/B AND2X1_LOC_600/a_8_24# 0.07fF
C44465 OR2X1_LOC_756/B AND2X1_LOC_616/a_36_24# 0.01fF
C45288 OR2X1_LOC_653/B OR2X1_LOC_756/B 0.01fF
C45912 OR2X1_LOC_756/B OR2X1_LOC_33/B 0.01fF
C45960 OR2X1_LOC_756/B OR2X1_LOC_287/a_8_216# 0.02fF
C46110 OR2X1_LOC_756/B OR2X1_LOC_333/A 0.01fF
C46434 OR2X1_LOC_756/B OR2X1_LOC_532/B 0.64fF
C46478 OR2X1_LOC_756/B OR2X1_LOC_343/B 0.15fF
C47349 OR2X1_LOC_756/B OR2X1_LOC_286/B 0.01fF
C48439 OR2X1_LOC_756/B VDD 2.38fF
C48523 AND2X1_LOC_755/a_8_24# OR2X1_LOC_756/B 0.02fF
C48860 OR2X1_LOC_756/B OR2X1_LOC_334/B 0.01fF
C49204 OR2X1_LOC_756/B OR2X1_LOC_756/a_36_216# 0.03fF
C49661 OR2X1_LOC_756/B AND2X1_LOC_83/a_8_24# 0.02fF
C49705 OR2X1_LOC_756/B AND2X1_LOC_179/a_36_24# 0.01fF
C50572 OR2X1_LOC_756/B OR2X1_LOC_840/A 0.03fF
C50603 OR2X1_LOC_756/B OR2X1_LOC_260/a_8_216# 0.02fF
C51066 OR2X1_LOC_756/B AND2X1_LOC_385/a_8_24# 0.11fF
C51437 OR2X1_LOC_160/A OR2X1_LOC_756/B 0.10fF
C51490 OR2X1_LOC_756/B AND2X1_LOC_86/B 0.07fF
C51505 OR2X1_LOC_756/B OR2X1_LOC_624/B 0.02fF
C52216 OR2X1_LOC_756/B OR2X1_LOC_78/Y 0.08fF
C52307 OR2X1_LOC_756/B OR2X1_LOC_285/A 0.01fF
C52709 OR2X1_LOC_756/B OR2X1_LOC_185/A 0.65fF
C52788 OR2X1_LOC_756/B OR2X1_LOC_435/Y 0.01fF
C52842 OR2X1_LOC_756/B AND2X1_LOC_431/a_8_24# 0.01fF
C53677 OR2X1_LOC_756/B AND2X1_LOC_442/a_8_24# 0.03fF
C54373 OR2X1_LOC_168/a_8_216# OR2X1_LOC_756/B 0.01fF
C54385 OR2X1_LOC_756/B AND2X1_LOC_617/a_8_24# 0.03fF
C54769 OR2X1_LOC_756/B OR2X1_LOC_436/B 0.01fF
C54834 OR2X1_LOC_756/B OR2X1_LOC_778/Y 0.03fF
C55070 AND2X1_LOC_91/B OR2X1_LOC_756/B 0.65fF
C55245 OR2X1_LOC_756/B OR2X1_LOC_799/A 0.04fF
C55373 OR2X1_LOC_756/B AND2X1_LOC_600/a_36_24# 0.01fF
C55467 OR2X1_LOC_756/B OR2X1_LOC_303/B 0.03fF
C55614 OR2X1_LOC_756/B OR2X1_LOC_105/a_8_216# 0.05fF
C55697 OR2X1_LOC_756/B AND2X1_LOC_56/B 0.15fF
C57854 OR2X1_LOC_756/B VSS 0.79fF
C152 OR2X1_LOC_160/B OR2X1_LOC_61/A 0.10fF
C589 OR2X1_LOC_160/B OR2X1_LOC_706/a_8_216# -0.02fF
C1484 AND2X1_LOC_229/a_8_24# OR2X1_LOC_160/B 0.03fF
C2217 OR2X1_LOC_160/B OR2X1_LOC_241/B 0.92fF
C2327 OR2X1_LOC_188/Y OR2X1_LOC_160/B 0.05fF
C2557 OR2X1_LOC_160/B OR2X1_LOC_193/A 0.02fF
C2752 OR2X1_LOC_208/A OR2X1_LOC_160/B 1.16fF
C2788 OR2X1_LOC_160/B AND2X1_LOC_438/a_8_24# 0.04fF
C2814 OR2X1_LOC_160/B AND2X1_LOC_505/a_8_24# 0.03fF
C2847 OR2X1_LOC_335/Y OR2X1_LOC_160/B 0.10fF
C2898 OR2X1_LOC_160/B OR2X1_LOC_537/A 0.01fF
C3185 OR2X1_LOC_138/a_8_216# OR2X1_LOC_160/B 0.06fF
C3771 OR2X1_LOC_160/B OR2X1_LOC_810/A 0.10fF
C4389 OR2X1_LOC_160/B OR2X1_LOC_338/B 0.01fF
C4502 OR2X1_LOC_656/B OR2X1_LOC_160/B 0.07fF
C4515 AND2X1_LOC_767/a_8_24# OR2X1_LOC_160/B 0.04fF
C4622 OR2X1_LOC_160/B AND2X1_LOC_45/a_8_24# 0.09fF
C4942 OR2X1_LOC_160/B OR2X1_LOC_687/Y 0.07fF
C5708 OR2X1_LOC_160/B OR2X1_LOC_78/A 0.12fF
C6697 OR2X1_LOC_160/B AND2X1_LOC_171/a_8_24# 0.03fF
C6740 OR2X1_LOC_160/B AND2X1_LOC_75/a_36_24# 0.01fF
C6860 OR2X1_LOC_160/B OR2X1_LOC_318/B 0.03fF
C7002 OR2X1_LOC_114/B OR2X1_LOC_160/B 0.03fF
C7158 OR2X1_LOC_160/B AND2X1_LOC_496/a_8_24# 0.06fF
C7951 OR2X1_LOC_160/B OR2X1_LOC_623/B 0.07fF
C8348 OR2X1_LOC_160/B OR2X1_LOC_507/A 0.10fF
C9279 OR2X1_LOC_160/B OR2X1_LOC_448/Y 0.11fF
C9982 OR2X1_LOC_160/B OR2X1_LOC_338/A 0.01fF
C10115 OR2X1_LOC_773/B OR2X1_LOC_160/B 0.03fF
C10128 AND2X1_LOC_81/B OR2X1_LOC_160/B 0.03fF
C10220 OR2X1_LOC_160/B OR2X1_LOC_196/B 0.07fF
C11296 OR2X1_LOC_160/B OR2X1_LOC_78/B 0.38fF
C11371 OR2X1_LOC_160/B OR2X1_LOC_375/A 3.67fF
C11695 OR2X1_LOC_160/B OR2X1_LOC_549/A 0.14fF
C12169 OR2X1_LOC_160/B OR2X1_LOC_499/B 0.09fF
C12532 AND2X1_LOC_229/a_36_24# OR2X1_LOC_160/B 0.01fF
C12983 OR2X1_LOC_160/B AND2X1_LOC_603/a_8_24# 0.05fF
C13278 OR2X1_LOC_160/B OR2X1_LOC_779/Y 0.03fF
C13538 OR2X1_LOC_160/B OR2X1_LOC_673/Y 0.03fF
C13858 OR2X1_LOC_160/B AND2X1_LOC_505/a_36_24# 0.01fF
C14202 OR2X1_LOC_160/B OR2X1_LOC_712/B 0.01fF
C14242 OR2X1_LOC_139/A OR2X1_LOC_160/B 0.74fF
C14670 OR2X1_LOC_160/B OR2X1_LOC_138/A 0.06fF
C15098 AND2X1_LOC_595/a_8_24# OR2X1_LOC_160/B 0.04fF
C15247 OR2X1_LOC_160/B AND2X1_LOC_666/a_8_24# 0.01fF
C15614 OR2X1_LOC_160/B OR2X1_LOC_87/A 6.33fF
C15842 OR2X1_LOC_160/B OR2X1_LOC_844/B 0.06fF
C15927 OR2X1_LOC_160/B OR2X1_LOC_389/A 0.01fF
C16388 OR2X1_LOC_160/B OR2X1_LOC_61/B 0.03fF
C16750 OR2X1_LOC_97/A OR2X1_LOC_160/B 0.12fF
C16821 OR2X1_LOC_160/B OR2X1_LOC_541/A 0.02fF
C16826 AND2X1_LOC_744/a_8_24# OR2X1_LOC_160/B 0.01fF
C17186 OR2X1_LOC_160/B OR2X1_LOC_691/Y 0.03fF
C17203 OR2X1_LOC_160/B OR2X1_LOC_713/A 0.01fF
C17296 OR2X1_LOC_160/B OR2X1_LOC_249/a_8_216# 0.07fF
C17759 OR2X1_LOC_160/B OR2X1_LOC_333/B 0.26fF
C18181 OR2X1_LOC_154/A OR2X1_LOC_160/B 2.91fF
C18197 OR2X1_LOC_160/B OR2X1_LOC_267/A 0.01fF
C18245 OR2X1_LOC_160/B OR2X1_LOC_778/A 0.10fF
C18964 OR2X1_LOC_538/a_8_216# OR2X1_LOC_160/B 0.01fF
C19145 OR2X1_LOC_160/B OR2X1_LOC_335/B 0.03fF
C20823 OR2X1_LOC_160/B OR2X1_LOC_719/A 0.02fF
C21878 OR2X1_LOC_160/B OR2X1_LOC_333/A 0.01fF
C21935 OR2X1_LOC_160/B OR2X1_LOC_113/B 0.20fF
C21950 OR2X1_LOC_160/B OR2X1_LOC_450/A 0.11fF
C22174 OR2X1_LOC_160/B OR2X1_LOC_532/B 0.11fF
C23264 OR2X1_LOC_160/B OR2X1_LOC_778/a_8_216# 0.05fF
C24048 OR2X1_LOC_160/B AND2X1_LOC_603/a_36_24# 0.01fF
C24063 OR2X1_LOC_160/B AND2X1_LOC_265/a_8_24# 0.04fF
C24077 OR2X1_LOC_160/B VDD 1.42fF
C24840 OR2X1_LOC_335/a_8_216# OR2X1_LOC_160/B 0.06fF
C24893 OR2X1_LOC_160/B OR2X1_LOC_676/Y 0.07fF
C24910 OR2X1_LOC_160/B OR2X1_LOC_834/A 0.06fF
C25902 OR2X1_LOC_160/B AND2X1_LOC_667/a_8_24# 0.03fF
C26087 OR2X1_LOC_160/B OR2X1_LOC_115/B 0.03fF
C26185 OR2X1_LOC_160/B OR2X1_LOC_840/A 0.05fF
C26852 OR2X1_LOC_160/B OR2X1_LOC_750/Y 0.07fF
C27075 OR2X1_LOC_160/A OR2X1_LOC_160/B 1.83fF
C27162 OR2X1_LOC_160/B OR2X1_LOC_624/B 0.49fF
C27780 OR2X1_LOC_113/a_8_216# OR2X1_LOC_160/B 0.02fF
C27851 OR2X1_LOC_160/B OR2X1_LOC_78/Y 0.05fF
C27869 OR2X1_LOC_160/B AND2X1_LOC_424/a_8_24# 0.01fF
C28349 OR2X1_LOC_160/B OR2X1_LOC_185/A 0.05fF
C28354 OR2X1_LOC_160/B OR2X1_LOC_249/Y 0.01fF
C28812 OR2X1_LOC_702/A OR2X1_LOC_160/B 0.72fF
C29513 OR2X1_LOC_160/B OR2X1_LOC_641/A 6.23fF
C29637 OR2X1_LOC_160/B OR2X1_LOC_449/A 0.01fF
C30022 OR2X1_LOC_160/B OR2X1_LOC_541/B 0.01fF
C30289 OR2X1_LOC_160/B AND2X1_LOC_238/a_8_24# 0.01fF
C30467 OR2X1_LOC_160/B OR2X1_LOC_643/A 0.08fF
C30471 OR2X1_LOC_160/B OR2X1_LOC_778/Y 0.15fF
C30542 OR2X1_LOC_160/B OR2X1_LOC_113/A 0.01fF
C30709 AND2X1_LOC_91/B OR2X1_LOC_160/B 0.64fF
C30842 OR2X1_LOC_308/a_8_216# OR2X1_LOC_160/B 0.03fF
C31106 OR2X1_LOC_160/B OR2X1_LOC_446/B 0.07fF
C31198 OR2X1_LOC_160/B OR2X1_LOC_719/B 0.02fF
C31320 OR2X1_LOC_160/B AND2X1_LOC_56/B 0.06fF
C32681 OR2X1_LOC_160/B AND2X1_LOC_47/Y 0.59fF
C32973 OR2X1_LOC_160/B AND2X1_LOC_695/a_8_24# 0.01fF
C33087 OR2X1_LOC_160/B OR2X1_LOC_780/A 0.01fF
C34197 OR2X1_LOC_160/B AND2X1_LOC_173/a_8_24# 0.01fF
C34585 OR2X1_LOC_160/B OR2X1_LOC_235/B 0.03fF
C35374 OR2X1_LOC_160/B OR2X1_LOC_362/A 0.07fF
C35452 OR2X1_LOC_539/A OR2X1_LOC_160/B 0.01fF
C35865 OR2X1_LOC_160/B OR2X1_LOC_678/a_8_216# 0.03fF
C36202 OR2X1_LOC_156/a_8_216# OR2X1_LOC_160/B 0.01fF
C36617 OR2X1_LOC_160/B AND2X1_LOC_44/Y 3.99fF
C36848 OR2X1_LOC_160/B OR2X1_LOC_720/B 0.03fF
C37522 OR2X1_LOC_160/B AND2X1_LOC_18/Y 5.33fF
C37916 OR2X1_LOC_160/B OR2X1_LOC_307/A 0.03fF
C38461 OR2X1_LOC_160/B OR2X1_LOC_707/A 0.01fF
C38466 OR2X1_LOC_160/B OR2X1_LOC_130/A 0.21fF
C38892 OR2X1_LOC_160/B AND2X1_LOC_487/a_8_24# 0.04fF
C38934 OR2X1_LOC_160/B OR2X1_LOC_449/B 5.09fF
C40257 OR2X1_LOC_160/B OR2X1_LOC_447/Y 0.03fF
C40574 OR2X1_LOC_160/B OR2X1_LOC_161/A 0.18fF
C40658 OR2X1_LOC_160/B AND2X1_LOC_51/Y 4.48fF
C41009 OR2X1_LOC_160/B OR2X1_LOC_541/a_8_216# 0.01fF
C41389 OR2X1_LOC_160/B AND2X1_LOC_41/A 1.31fF
C41489 OR2X1_LOC_160/B OR2X1_LOC_631/B 0.03fF
C41536 OR2X1_LOC_160/B AND2X1_LOC_135/a_8_24# 0.01fF
C42289 OR2X1_LOC_105/Y OR2X1_LOC_160/B 0.02fF
C42983 OR2X1_LOC_160/B AND2X1_LOC_31/Y 0.45fF
C43906 OR2X1_LOC_160/B AND2X1_LOC_36/Y 0.06fF
C43926 OR2X1_LOC_160/B OR2X1_LOC_333/a_8_216# 0.01fF
C43944 OR2X1_LOC_154/a_8_216# OR2X1_LOC_160/B 0.01fF
C43995 OR2X1_LOC_160/B OR2X1_LOC_630/Y 0.07fF
C45219 OR2X1_LOC_308/A OR2X1_LOC_160/B 0.03fF
C45419 OR2X1_LOC_160/B OR2X1_LOC_557/A 0.03fF
C45453 OR2X1_LOC_160/B OR2X1_LOC_675/A 0.01fF
C45729 OR2X1_LOC_768/A OR2X1_LOC_160/B 0.02fF
C46290 OR2X1_LOC_160/B OR2X1_LOC_269/B 0.12fF
C46343 OR2X1_LOC_160/B AND2X1_LOC_75/a_8_24# 0.04fF
C47355 OR2X1_LOC_160/B AND2X1_LOC_237/a_8_24# 0.01fF
C47429 OR2X1_LOC_160/B OR2X1_LOC_777/B 0.07fF
C47475 OR2X1_LOC_188/a_8_216# OR2X1_LOC_160/B 0.01fF
C47481 OR2X1_LOC_156/Y OR2X1_LOC_160/B 0.15fF
C47921 OR2X1_LOC_160/B OR2X1_LOC_161/B 0.26fF
C48042 OR2X1_LOC_160/B AND2X1_LOC_536/a_8_24# 0.01fF
C48308 OR2X1_LOC_160/B OR2X1_LOC_707/a_8_216# -0.00fF
C49453 OR2X1_LOC_160/B AND2X1_LOC_106/a_8_24# 0.04fF
C49635 OR2X1_LOC_160/B OR2X1_LOC_489/A 0.03fF
C50153 OR2X1_LOC_160/B OR2X1_LOC_489/B -0.01fF
C51522 OR2X1_LOC_160/B OR2X1_LOC_446/Y 0.15fF
C51881 OR2X1_LOC_160/B OR2X1_LOC_287/B 0.04fF
C51908 OR2X1_LOC_160/B OR2X1_LOC_76/A 0.13fF
C52247 OR2X1_LOC_160/B OR2X1_LOC_553/A 0.50fF
C53000 OR2X1_LOC_160/B OR2X1_LOC_151/A 0.07fF
C55062 OR2X1_LOC_156/B OR2X1_LOC_160/B 0.01fF
C55466 OR2X1_LOC_160/B OR2X1_LOC_308/Y 0.01fF
C57848 OR2X1_LOC_160/B VSS 0.98fF
C449 OR2X1_LOC_789/B OR2X1_LOC_193/A 0.13fF
C15137 OR2X1_LOC_789/B OR2X1_LOC_691/Y 0.01fF
C24289 OR2X1_LOC_789/B OR2X1_LOC_789/a_8_216# 0.47fF
C35490 OR2X1_LOC_789/B AND2X1_LOC_18/Y 0.11fF
C35762 OR2X1_LOC_789/B OR2X1_LOC_789/A 0.17fF
C41778 OR2X1_LOC_789/B AND2X1_LOC_36/Y 0.01fF
C57823 OR2X1_LOC_789/B VSS 0.16fF
C2926 OR2X1_LOC_490/Y OR2X1_LOC_595/A 0.01fF
C4784 OR2X1_LOC_490/Y OR2X1_LOC_95/Y 0.07fF
C6002 OR2X1_LOC_70/Y OR2X1_LOC_490/Y 0.09fF
C11979 OR2X1_LOC_3/Y OR2X1_LOC_490/Y 0.01fF
C19614 OR2X1_LOC_490/Y OR2X1_LOC_118/Y 0.03fF
C28946 AND2X1_LOC_489/Y OR2X1_LOC_490/Y 0.02fF
C33500 OR2X1_LOC_490/Y OR2X1_LOC_91/A 0.14fF
C36322 OR2X1_LOC_106/Y OR2X1_LOC_490/Y 0.01fF
C36870 OR2X1_LOC_490/Y AND2X1_LOC_99/A 0.09fF
C37630 AND2X1_LOC_362/B OR2X1_LOC_490/Y 0.68fF
C41897 OR2X1_LOC_117/a_8_216# OR2X1_LOC_490/Y 0.42fF
C42970 OR2X1_LOC_490/Y OR2X1_LOC_131/Y 0.01fF
C43261 VDD OR2X1_LOC_490/Y 0.24fF
C43479 OR2X1_LOC_490/Y OR2X1_LOC_67/Y 0.01fF
C49391 OR2X1_LOC_490/Y OR2X1_LOC_744/A 0.20fF
C50658 OR2X1_LOC_490/Y OR2X1_LOC_56/A 0.02fF
C54515 OR2X1_LOC_490/Y AND2X1_LOC_361/A 0.01fF
C56133 OR2X1_LOC_490/Y OR2X1_LOC_600/A 0.03fF
C57753 OR2X1_LOC_490/Y VSS 0.10fF
C7390 AND2X1_LOC_593/Y OR2X1_LOC_534/Y 0.21fF
C19496 OR2X1_LOC_533/A OR2X1_LOC_534/Y 0.19fF
C20544 VDD OR2X1_LOC_534/Y 0.12fF
C26120 AND2X1_LOC_390/B OR2X1_LOC_534/Y 0.01fF
C28254 OR2X1_LOC_417/Y OR2X1_LOC_534/Y 0.09fF
C31327 OR2X1_LOC_534/Y OR2X1_LOC_331/Y 0.07fF
C33245 OR2X1_LOC_619/Y OR2X1_LOC_534/Y 0.03fF
C35587 OR2X1_LOC_13/B OR2X1_LOC_534/Y 0.03fF
C39218 OR2X1_LOC_70/Y OR2X1_LOC_534/Y 0.01fF
C42997 AND2X1_LOC_535/a_8_24# OR2X1_LOC_534/Y 0.09fF
C54521 OR2X1_LOC_533/Y OR2X1_LOC_534/Y 0.18fF
C56404 OR2X1_LOC_534/Y VSS 0.18fF
C13140 AND2X1_LOC_847/Y OR2X1_LOC_297/A 0.01fF
C21190 OR2X1_LOC_427/A OR2X1_LOC_297/A 0.01fF
C23239 OR2X1_LOC_158/A OR2X1_LOC_297/A 0.01fF
C23799 OR2X1_LOC_748/A OR2X1_LOC_297/A 0.02fF
C27031 OR2X1_LOC_56/A OR2X1_LOC_297/A 0.01fF
C29017 OR2X1_LOC_297/A AND2X1_LOC_789/Y 0.02fF
C32460 OR2X1_LOC_600/A OR2X1_LOC_297/A 0.03fF
C35367 OR2X1_LOC_297/A OR2X1_LOC_428/A 0.81fF
C36411 OR2X1_LOC_89/A OR2X1_LOC_297/A 0.01fF
C53463 OR2X1_LOC_604/A OR2X1_LOC_297/A 0.04fF
C56714 OR2X1_LOC_297/A VSS 0.18fF
C1899 OR2X1_LOC_43/Y OR2X1_LOC_600/A 0.08fF
C10567 OR2X1_LOC_43/Y AND2X1_LOC_729/B 0.02fF
C11089 OR2X1_LOC_43/Y OR2X1_LOC_41/Y 0.23fF
C24879 OR2X1_LOC_43/Y AND2X1_LOC_434/Y 0.08fF
C42180 OR2X1_LOC_43/Y OR2X1_LOC_13/Y 0.01fF
C45247 VDD OR2X1_LOC_43/Y 0.16fF
C49604 OR2X1_LOC_43/Y AND2X1_LOC_195/a_8_24# 0.23fF
C57701 OR2X1_LOC_43/Y VSS 0.07fF
C2726 OR2X1_LOC_419/Y AND2X1_LOC_624/A 0.03fF
C5638 OR2X1_LOC_419/Y OR2X1_LOC_238/Y 0.05fF
C6820 OR2X1_LOC_177/Y OR2X1_LOC_419/Y 0.03fF
C6842 OR2X1_LOC_604/A OR2X1_LOC_419/Y 0.17fF
C7353 OR2X1_LOC_419/Y AND2X1_LOC_447/a_8_24# 0.01fF
C7758 OR2X1_LOC_164/Y OR2X1_LOC_419/Y 0.05fF
C10400 OR2X1_LOC_419/Y OR2X1_LOC_239/a_8_216# 0.01fF
C14617 AND2X1_LOC_729/Y OR2X1_LOC_419/Y 0.48fF
C14632 AND2X1_LOC_784/A OR2X1_LOC_419/Y 0.10fF
C15757 OR2X1_LOC_485/Y OR2X1_LOC_419/Y 0.14fF
C15831 OR2X1_LOC_419/Y OR2X1_LOC_39/A 0.11fF
C16279 AND2X1_LOC_593/Y OR2X1_LOC_419/Y 0.01fF
C16644 OR2X1_LOC_51/Y OR2X1_LOC_419/Y 0.06fF
C16701 OR2X1_LOC_680/A OR2X1_LOC_419/Y 0.10fF
C19213 OR2X1_LOC_600/a_8_216# OR2X1_LOC_419/Y 0.39fF
C20600 OR2X1_LOC_74/A OR2X1_LOC_419/Y 0.17fF
C21477 OR2X1_LOC_419/Y OR2X1_LOC_239/Y 0.49fF
C24423 OR2X1_LOC_485/A OR2X1_LOC_419/Y 0.09fF
C24836 OR2X1_LOC_420/a_8_216# OR2X1_LOC_419/Y 0.01fF
C28009 OR2X1_LOC_516/Y OR2X1_LOC_419/Y 0.06fF
C29359 VDD OR2X1_LOC_419/Y 2.74fF
C30290 OR2X1_LOC_419/Y OR2X1_LOC_591/A 0.02fF
C30666 OR2X1_LOC_427/A OR2X1_LOC_419/Y 0.10fF
C32227 OR2X1_LOC_45/B OR2X1_LOC_419/Y 0.06fF
C33140 OR2X1_LOC_482/Y OR2X1_LOC_419/Y 0.03fF
C35260 OR2X1_LOC_744/A OR2X1_LOC_419/Y 0.16fF
C35312 AND2X1_LOC_840/B OR2X1_LOC_419/Y 0.10fF
C35778 OR2X1_LOC_420/Y OR2X1_LOC_419/Y 0.22fF
C36528 OR2X1_LOC_419/Y OR2X1_LOC_56/A 0.05fF
C37001 OR2X1_LOC_91/Y OR2X1_LOC_419/Y 0.10fF
C37375 AND2X1_LOC_330/a_8_24# OR2X1_LOC_419/Y 0.32fF
C39181 OR2X1_LOC_497/Y OR2X1_LOC_419/Y 0.49fF
C39579 OR2X1_LOC_109/a_8_216# OR2X1_LOC_419/Y 0.10fF
C41152 AND2X1_LOC_787/A OR2X1_LOC_419/Y 0.03fF
C42084 OR2X1_LOC_600/A OR2X1_LOC_419/Y 0.22fF
C42965 OR2X1_LOC_331/A OR2X1_LOC_419/Y 0.01fF
C44536 OR2X1_LOC_419/Y OR2X1_LOC_13/B 0.10fF
C45546 OR2X1_LOC_528/Y OR2X1_LOC_419/Y 0.07fF
C45629 OR2X1_LOC_516/A OR2X1_LOC_419/Y 0.01fF
C46101 OR2X1_LOC_89/A OR2X1_LOC_419/Y 1.28fF
C46362 OR2X1_LOC_419/Y AND2X1_LOC_590/a_8_24# 0.11fF
C46879 OR2X1_LOC_491/a_8_216# OR2X1_LOC_419/Y 0.12fF
C47038 AND2X1_LOC_727/A OR2X1_LOC_419/Y 0.03fF
C47078 OR2X1_LOC_95/Y OR2X1_LOC_419/Y 0.69fF
C47857 OR2X1_LOC_419/Y AND2X1_LOC_621/Y 0.03fF
C48353 OR2X1_LOC_70/Y OR2X1_LOC_419/Y 3.36fF
C48421 OR2X1_LOC_184/Y OR2X1_LOC_419/Y 0.05fF
C48659 AND2X1_LOC_330/a_36_24# OR2X1_LOC_419/Y 0.06fF
C49522 OR2X1_LOC_484/Y OR2X1_LOC_419/Y 0.10fF
C49916 OR2X1_LOC_108/Y OR2X1_LOC_419/Y 0.10fF
C50772 OR2X1_LOC_419/Y AND2X1_LOC_447/Y 0.01fF
C50829 OR2X1_LOC_109/Y OR2X1_LOC_419/Y 0.09fF
C51320 AND2X1_LOC_227/Y OR2X1_LOC_419/Y 0.05fF
C52004 OR2X1_LOC_40/Y OR2X1_LOC_419/Y 0.08fF
C52421 OR2X1_LOC_491/a_36_216# OR2X1_LOC_419/Y 0.17fF
C53315 OR2X1_LOC_495/Y OR2X1_LOC_419/Y 0.05fF
C55509 OR2X1_LOC_64/Y OR2X1_LOC_419/Y 0.76fF
C56925 OR2X1_LOC_419/Y VSS 0.53fF
C30581 OR2X1_LOC_827/Y AND2X1_LOC_838/Y 0.23fF
C42932 OR2X1_LOC_827/Y AND2X1_LOC_838/a_8_24# 0.08fF
C50852 OR2X1_LOC_827/Y AND2X1_LOC_838/B 0.10fF
C57422 OR2X1_LOC_827/Y VSS -0.06fF
C752 OR2X1_LOC_589/A OR2X1_LOC_272/Y 0.02fF
C1799 OR2X1_LOC_3/Y OR2X1_LOC_272/Y 0.11fF
C3122 OR2X1_LOC_272/Y OR2X1_LOC_64/Y 0.05fF
C9043 OR2X1_LOC_272/Y AND2X1_LOC_78/a_8_24# 0.16fF
C14567 OR2X1_LOC_272/Y OR2X1_LOC_79/A 0.19fF
C18810 OR2X1_LOC_272/Y OR2X1_LOC_52/B 0.05fF
C18897 OR2X1_LOC_272/Y AND2X1_LOC_216/A 0.30fF
C19628 OR2X1_LOC_272/Y OR2X1_LOC_39/A 0.02fF
C23413 OR2X1_LOC_272/Y OR2X1_LOC_91/A 0.05fF
C24348 OR2X1_LOC_272/Y OR2X1_LOC_74/A 0.05fF
C25776 OR2X1_LOC_134/Y OR2X1_LOC_272/Y 0.04fF
C33033 VDD OR2X1_LOC_272/Y 0.53fF
C36087 OR2X1_LOC_272/Y OR2X1_LOC_767/a_8_216# 0.01fF
C36379 OR2X1_LOC_158/A OR2X1_LOC_272/Y 0.03fF
C41639 OR2X1_LOC_272/Y AND2X1_LOC_139/B 0.03fF
C48398 OR2X1_LOC_272/Y OR2X1_LOC_13/B 0.03fF
C48900 OR2X1_LOC_272/Y OR2X1_LOC_595/A 0.03fF
C49933 OR2X1_LOC_272/Y OR2X1_LOC_89/A 0.35fF
C50843 OR2X1_LOC_272/Y OR2X1_LOC_95/Y 0.02fF
C53082 OR2X1_LOC_272/Y OR2X1_LOC_767/Y 0.01fF
C54015 OR2X1_LOC_132/Y OR2X1_LOC_272/Y 0.09fF
C55010 OR2X1_LOC_272/Y AND2X1_LOC_227/Y 0.02fF
C57432 OR2X1_LOC_272/Y VSS -0.25fF
C12331 OR2X1_LOC_3/Y OR2X1_LOC_459/A 0.04fF
C30077 OR2X1_LOC_459/A OR2X1_LOC_39/A 0.09fF
C43586 VDD OR2X1_LOC_459/A 0.21fF
C57603 OR2X1_LOC_459/A VSS 0.12fF
C5646 OR2X1_LOC_136/Y OR2X1_LOC_40/Y 0.01fF
C6939 OR2X1_LOC_136/Y OR2X1_LOC_589/A 0.84fF
C7978 OR2X1_LOC_136/Y OR2X1_LOC_3/Y 0.05fF
C24511 AND2X1_LOC_784/A OR2X1_LOC_136/Y 0.42fF
C31946 OR2X1_LOC_136/Y AND2X1_LOC_339/B 0.02fF
C34177 OR2X1_LOC_136/Y AND2X1_LOC_303/A 0.08fF
C36674 OR2X1_LOC_136/Y AND2X1_LOC_138/a_8_24# 0.11fF
C39197 OR2X1_LOC_136/Y VDD 0.27fF
C47678 OR2X1_LOC_136/Y AND2X1_LOC_831/Y 0.03fF
C54530 OR2X1_LOC_136/Y OR2X1_LOC_13/B 0.06fF
C57934 OR2X1_LOC_136/Y VSS 0.06fF
C218 OR2X1_LOC_56/A OR2X1_LOC_627/Y 0.01fF
C1824 OR2X1_LOC_56/A OR2X1_LOC_521/a_36_216# 0.01fF
C1864 OR2X1_LOC_516/Y OR2X1_LOC_56/A 0.03fF
C2263 OR2X1_LOC_56/A AND2X1_LOC_793/B 0.07fF
C2464 AND2X1_LOC_348/A OR2X1_LOC_56/A 0.03fF
C2628 OR2X1_LOC_442/a_8_216# OR2X1_LOC_56/A 0.20fF
C2661 AND2X1_LOC_798/A OR2X1_LOC_56/A 0.03fF
C3254 VDD OR2X1_LOC_56/A 1.17fF
C3384 OR2X1_LOC_251/Y OR2X1_LOC_56/A 0.07fF
C3416 OR2X1_LOC_826/a_8_216# OR2X1_LOC_56/A 0.04fF
C4098 OR2X1_LOC_382/Y OR2X1_LOC_56/A 0.01fF
C4165 OR2X1_LOC_495/a_36_216# OR2X1_LOC_56/A 0.02fF
C4413 OR2X1_LOC_494/A OR2X1_LOC_56/A 0.08fF
C4517 OR2X1_LOC_427/A OR2X1_LOC_56/A 5.92fF
C4555 AND2X1_LOC_464/a_8_24# OR2X1_LOC_56/A 0.01fF
C5333 OR2X1_LOC_281/a_8_216# OR2X1_LOC_56/A 0.01fF
C5375 OR2X1_LOC_67/a_36_216# OR2X1_LOC_56/A 0.03fF
C5804 OR2X1_LOC_45/a_8_216# OR2X1_LOC_56/A 0.03fF
C5889 AND2X1_LOC_116/Y OR2X1_LOC_56/A 0.04fF
C6106 OR2X1_LOC_45/B OR2X1_LOC_56/A 0.82fF
C6170 OR2X1_LOC_292/a_8_216# OR2X1_LOC_56/A 0.02fF
C6547 OR2X1_LOC_158/A OR2X1_LOC_56/A 19.94fF
C7032 OR2X1_LOC_816/Y OR2X1_LOC_56/A 0.02fF
C7187 OR2X1_LOC_304/Y OR2X1_LOC_56/A 0.13fF
C7596 OR2X1_LOC_117/Y OR2X1_LOC_56/A 0.02fF
C8769 AND2X1_LOC_541/Y OR2X1_LOC_56/A 0.04fF
C8862 OR2X1_LOC_316/Y OR2X1_LOC_56/A 0.03fF
C8933 AND2X1_LOC_390/B OR2X1_LOC_56/A 0.14fF
C8958 OR2X1_LOC_431/Y OR2X1_LOC_56/A 0.02fF
C9224 OR2X1_LOC_744/A OR2X1_LOC_56/A 0.17fF
C9330 AND2X1_LOC_840/B OR2X1_LOC_56/A 0.05fF
C9373 OR2X1_LOC_282/a_8_216# OR2X1_LOC_56/A 0.05fF
C9552 OR2X1_LOC_56/A OR2X1_LOC_320/a_8_216# 0.01fF
C9590 OR2X1_LOC_56/A AND2X1_LOC_464/A 0.03fF
C10078 OR2X1_LOC_179/a_8_216# OR2X1_LOC_56/A 0.01fF
C10150 AND2X1_LOC_303/B OR2X1_LOC_56/A 0.21fF
C10885 OR2X1_LOC_56/A AND2X1_LOC_285/Y 0.03fF
C10960 OR2X1_LOC_91/Y OR2X1_LOC_56/A 0.03fF
C11031 OR2X1_LOC_527/Y OR2X1_LOC_56/A 0.03fF
C11057 OR2X1_LOC_311/Y OR2X1_LOC_56/A 0.06fF
C11064 AND2X1_LOC_538/Y OR2X1_LOC_56/A 0.09fF
C11329 OR2X1_LOC_494/a_8_216# OR2X1_LOC_56/A 0.05fF
C11460 AND2X1_LOC_276/Y OR2X1_LOC_56/A 0.06fF
C11526 AND2X1_LOC_831/Y OR2X1_LOC_56/A 0.07fF
C11771 AND2X1_LOC_335/a_8_24# OR2X1_LOC_56/A 0.03fF
C11780 OR2X1_LOC_441/Y OR2X1_LOC_56/A 0.06fF
C12102 OR2X1_LOC_135/a_8_216# OR2X1_LOC_56/A 0.08fF
C12561 OR2X1_LOC_108/a_8_216# OR2X1_LOC_56/A 0.01fF
C13640 OR2X1_LOC_7/a_8_216# OR2X1_LOC_56/A 0.02fF
C13981 AND2X1_LOC_319/A OR2X1_LOC_56/A 0.42fF
C14139 AND2X1_LOC_721/A OR2X1_LOC_56/A 0.03fF
C14411 OR2X1_LOC_56/A AND2X1_LOC_361/A 0.02fF
C14803 OR2X1_LOC_96/B OR2X1_LOC_56/A 0.04fF
C15940 OR2X1_LOC_600/A OR2X1_LOC_56/A 6.28fF
C15941 AND2X1_LOC_335/Y OR2X1_LOC_56/A 0.02fF
C16033 OR2X1_LOC_619/Y OR2X1_LOC_56/A 0.16fF
C16989 AND2X1_LOC_473/a_8_24# OR2X1_LOC_56/A 0.05fF
C17087 OR2X1_LOC_56/A OR2X1_LOC_406/A 0.29fF
C18425 OR2X1_LOC_56/A OR2X1_LOC_13/B 0.33fF
C18913 OR2X1_LOC_56/A OR2X1_LOC_428/A 1.21fF
C18920 OR2X1_LOC_56/A OR2X1_LOC_595/A 1.51fF
C19376 OR2X1_LOC_528/Y OR2X1_LOC_56/A 0.32fF
C19467 OR2X1_LOC_516/A OR2X1_LOC_56/A 0.10fF
C19971 OR2X1_LOC_89/A OR2X1_LOC_56/A 0.67fF
C20403 OR2X1_LOC_282/Y OR2X1_LOC_56/A 0.05fF
C20619 AND2X1_LOC_473/Y OR2X1_LOC_56/A 1.10fF
C20735 OR2X1_LOC_45/Y OR2X1_LOC_56/A 0.52fF
C20863 AND2X1_LOC_727/A OR2X1_LOC_56/A 0.06fF
C20908 OR2X1_LOC_95/Y OR2X1_LOC_56/A 0.45fF
C21129 OR2X1_LOC_122/Y OR2X1_LOC_56/A 0.01fF
C21149 OR2X1_LOC_179/Y OR2X1_LOC_56/A 0.02fF
C21590 OR2X1_LOC_438/Y OR2X1_LOC_56/A 0.07fF
C21631 AND2X1_LOC_621/Y OR2X1_LOC_56/A 0.12fF
C22140 OR2X1_LOC_70/Y OR2X1_LOC_56/A 0.11fF
C23244 AND2X1_LOC_535/Y OR2X1_LOC_56/A 0.03fF
C23635 OR2X1_LOC_56/A OR2X1_LOC_16/A 0.17fF
C23658 OR2X1_LOC_108/Y OR2X1_LOC_56/A 0.29fF
C24557 OR2X1_LOC_109/Y OR2X1_LOC_56/A 0.03fF
C24652 AND2X1_LOC_729/B OR2X1_LOC_56/A 0.03fF
C25029 OR2X1_LOC_106/A OR2X1_LOC_56/A 0.16fF
C25130 AND2X1_LOC_227/Y OR2X1_LOC_56/A 0.02fF
C25730 OR2X1_LOC_40/Y OR2X1_LOC_56/A 0.45fF
C25756 OR2X1_LOC_698/a_8_216# OR2X1_LOC_56/A 0.05fF
C25859 OR2X1_LOC_7/A OR2X1_LOC_56/A 0.53fF
C25875 OR2X1_LOC_320/Y OR2X1_LOC_56/A 0.01fF
C25949 OR2X1_LOC_224/a_8_216# OR2X1_LOC_56/A 0.01fF
C26376 OR2X1_LOC_615/Y OR2X1_LOC_56/A 0.12fF
C26972 OR2X1_LOC_589/A OR2X1_LOC_56/A 0.12fF
C27311 OR2X1_LOC_56/A OR2X1_LOC_384/a_8_216# 0.01fF
C27420 AND2X1_LOC_776/a_8_24# OR2X1_LOC_56/A 0.01fF
C28004 OR2X1_LOC_3/Y OR2X1_LOC_56/A 1.64fF
C28016 AND2X1_LOC_631/Y OR2X1_LOC_56/A 0.03fF
C28367 AND2X1_LOC_113/Y OR2X1_LOC_56/A 0.03fF
C29275 OR2X1_LOC_64/Y OR2X1_LOC_56/A 0.34fF
C29484 AND2X1_LOC_541/a_8_24# OR2X1_LOC_56/A 0.17fF
C29944 OR2X1_LOC_96/Y OR2X1_LOC_56/A 0.01fF
C30163 OR2X1_LOC_7/Y OR2X1_LOC_56/A 0.03fF
C30567 AND2X1_LOC_196/Y OR2X1_LOC_56/A 0.01fF
C30731 OR2X1_LOC_56/A OR2X1_LOC_321/a_8_216# 0.01fF
C30844 AND2X1_LOC_456/B OR2X1_LOC_56/A 0.03fF
C31374 OR2X1_LOC_321/Y OR2X1_LOC_56/A 0.01fF
C31804 AND2X1_LOC_116/B OR2X1_LOC_56/A 0.19fF
C31848 OR2X1_LOC_96/a_8_216# OR2X1_LOC_56/A 0.02fF
C31983 OR2X1_LOC_56/A AND2X1_LOC_802/Y 0.03fF
C32443 OR2X1_LOC_56/A AND2X1_LOC_778/Y 0.04fF
C32569 AND2X1_LOC_624/A OR2X1_LOC_56/A 0.07fF
C32911 OR2X1_LOC_56/A AND2X1_LOC_434/a_8_24# 0.04fF
C33443 AND2X1_LOC_777/a_8_24# OR2X1_LOC_56/A 0.01fF
C33594 AND2X1_LOC_114/Y OR2X1_LOC_56/A 0.01fF
C33646 OR2X1_LOC_56/A OR2X1_LOC_172/a_8_216# -0.03fF
C33721 OR2X1_LOC_56/A OR2X1_LOC_312/a_8_216# 0.02fF
C33854 AND2X1_LOC_114/a_8_24# OR2X1_LOC_56/A 0.01fF
C33918 OR2X1_LOC_48/Y OR2X1_LOC_56/A 0.01fF
C34649 OR2X1_LOC_56/A OR2X1_LOC_278/Y 0.03fF
C34782 OR2X1_LOC_253/a_8_216# OR2X1_LOC_56/A 0.03fF
C35313 OR2X1_LOC_56/A OR2X1_LOC_142/Y 0.04fF
C35467 OR2X1_LOC_56/A OR2X1_LOC_16/a_8_216# 0.08fF
C35505 OR2X1_LOC_118/Y OR2X1_LOC_56/A 0.02fF
C35572 OR2X1_LOC_56/A OR2X1_LOC_238/Y 0.12fF
C36645 OR2X1_LOC_177/Y OR2X1_LOC_56/A 0.03fF
C36662 OR2X1_LOC_604/A OR2X1_LOC_56/A 1.48fF
C36743 OR2X1_LOC_252/a_8_216# OR2X1_LOC_56/A 0.08fF
C37459 OR2X1_LOC_56/A OR2X1_LOC_183/a_8_216# 0.03fF
C37567 OR2X1_LOC_164/Y OR2X1_LOC_56/A 0.02fF
C37887 AND2X1_LOC_539/Y OR2X1_LOC_56/A 0.03fF
C37946 AND2X1_LOC_326/B OR2X1_LOC_56/A 0.03fF
C38400 AND2X1_LOC_319/a_36_24# OR2X1_LOC_56/A 0.01fF
C38472 OR2X1_LOC_298/Y OR2X1_LOC_56/A 0.07fF
C38845 OR2X1_LOC_56/A AND2X1_LOC_434/Y 0.14fF
C39421 AND2X1_LOC_196/a_8_24# OR2X1_LOC_56/A 0.03fF
C39424 AND2X1_LOC_260/a_8_24# OR2X1_LOC_56/A 0.01fF
C40450 AND2X1_LOC_776/Y OR2X1_LOC_56/A 0.15fF
C40883 OR2X1_LOC_135/Y OR2X1_LOC_56/A 0.10fF
C41030 AND2X1_LOC_848/Y OR2X1_LOC_56/A 0.07fF
C41127 AND2X1_LOC_464/Y OR2X1_LOC_56/A 0.01fF
C41842 OR2X1_LOC_178/Y OR2X1_LOC_56/A 0.56fF
C42062 AND2X1_LOC_318/Y OR2X1_LOC_56/A 0.20fF
C42304 OR2X1_LOC_698/Y OR2X1_LOC_56/A 0.03fF
C42512 OR2X1_LOC_224/Y OR2X1_LOC_56/A 0.01fF
C42850 OR2X1_LOC_385/Y OR2X1_LOC_56/A 0.08fF
C43097 OR2X1_LOC_56/A AND2X1_LOC_810/B 0.07fF
C43996 AND2X1_LOC_715/A OR2X1_LOC_56/A 0.06fF
C44010 OR2X1_LOC_56/A AND2X1_LOC_434/a_36_24# 0.01fF
C44513 AND2X1_LOC_729/Y OR2X1_LOC_56/A 0.04fF
C44544 AND2X1_LOC_784/A OR2X1_LOC_56/A 0.10fF
C44553 AND2X1_LOC_778/a_8_24# OR2X1_LOC_56/A 0.01fF
C44714 OR2X1_LOC_56/A OR2X1_LOC_172/Y 0.02fF
C44808 OR2X1_LOC_56/A OR2X1_LOC_312/a_36_216# 0.03fF
C44993 OR2X1_LOC_56/A OR2X1_LOC_52/B 9.09fF
C45268 OR2X1_LOC_281/Y OR2X1_LOC_56/A 0.16fF
C45282 OR2X1_LOC_56/A OR2X1_LOC_253/Y 0.03fF
C45434 AND2X1_LOC_356/B OR2X1_LOC_56/A 0.09fF
C45441 OR2X1_LOC_280/Y OR2X1_LOC_56/A 0.03fF
C45815 OR2X1_LOC_56/A OR2X1_LOC_39/A 0.22fF
C46634 OR2X1_LOC_51/Y OR2X1_LOC_56/A 0.29fF
C46678 OR2X1_LOC_56/A OR2X1_LOC_16/Y 0.13fF
C46741 OR2X1_LOC_680/A OR2X1_LOC_56/A 0.06fF
C47545 OR2X1_LOC_178/a_8_216# OR2X1_LOC_56/A 0.03fF
C48070 OR2X1_LOC_252/Y OR2X1_LOC_56/A 0.02fF
C48733 OR2X1_LOC_56/A OR2X1_LOC_183/Y 0.13fF
C49330 OR2X1_LOC_237/Y OR2X1_LOC_56/A 0.03fF
C49558 OR2X1_LOC_56/A OR2X1_LOC_384/Y 0.03fF
C49690 OR2X1_LOC_91/A OR2X1_LOC_56/A 0.85fF
C50663 OR2X1_LOC_74/A OR2X1_LOC_56/A 4.86fF
C50684 AND2X1_LOC_196/a_36_24# OR2X1_LOC_56/A 0.01fF
C50921 OR2X1_LOC_56/A AND2X1_LOC_254/a_8_24# 0.03fF
C51442 AND2X1_LOC_151/a_8_24# OR2X1_LOC_56/A -0.00fF
C52105 OR2X1_LOC_134/Y OR2X1_LOC_56/A 0.02fF
C52172 OR2X1_LOC_816/a_8_216# OR2X1_LOC_56/A 0.02fF
C52482 OR2X1_LOC_56/A OR2X1_LOC_521/a_8_216# 0.03fF
C52553 OR2X1_LOC_106/Y OR2X1_LOC_56/A 0.04fF
C52601 OR2X1_LOC_505/Y OR2X1_LOC_56/A 0.01fF
C53113 AND2X1_LOC_99/A OR2X1_LOC_56/A 0.02fF
C53147 OR2X1_LOC_627/a_8_216# OR2X1_LOC_56/A 0.03fF
C53257 AND2X1_LOC_319/a_8_24# OR2X1_LOC_56/A 0.04fF
C54023 OR2X1_LOC_431/a_8_216# OR2X1_LOC_56/A 0.03fF
C54411 OR2X1_LOC_665/Y OR2X1_LOC_56/A 0.07fF
C54427 OR2X1_LOC_485/A OR2X1_LOC_56/A 0.22fF
C54806 OR2X1_LOC_495/a_8_216# OR2X1_LOC_56/A 0.02fF
C55058 AND2X1_LOC_383/a_8_24# OR2X1_LOC_56/A 0.01fF
C55135 OR2X1_LOC_122/a_8_216# OR2X1_LOC_56/A 0.02fF
C55236 AND2X1_LOC_458/Y OR2X1_LOC_56/A 0.01fF
C55239 AND2X1_LOC_302/a_8_24# OR2X1_LOC_56/A 0.09fF
C56093 OR2X1_LOC_67/a_8_216# OR2X1_LOC_56/A 0.03fF
C56208 AND2X1_LOC_537/Y OR2X1_LOC_56/A 0.10fF
C56716 OR2X1_LOC_56/A VSS -7.20fF
C1766 OR2X1_LOC_83/A AND2X1_LOC_612/B 0.23fF
C8168 AND2X1_LOC_612/B AND2X1_LOC_612/a_8_24# 0.03fF
C13064 AND2X1_LOC_612/B OR2X1_LOC_397/a_8_216# 0.47fF
C19209 AND2X1_LOC_612/B OR2X1_LOC_647/B 0.03fF
C23701 AND2X1_LOC_612/B OR2X1_LOC_415/Y 0.02fF
C36879 AND2X1_LOC_612/B OR2X1_LOC_375/A 0.03fF
C49795 VDD AND2X1_LOC_612/B 0.01fF
C56922 AND2X1_LOC_612/B VSS -0.12fF
C270 OR2X1_LOC_292/Y OR2X1_LOC_91/A 0.08fF
C1257 OR2X1_LOC_312/Y OR2X1_LOC_91/A 0.07fF
C1433 OR2X1_LOC_91/A OR2X1_LOC_13/B 3.20fF
C1918 OR2X1_LOC_91/A OR2X1_LOC_428/A 2.36fF
C1930 OR2X1_LOC_91/A OR2X1_LOC_595/A 0.07fF
C2519 AND2X1_LOC_342/Y OR2X1_LOC_91/A 0.12fF
C2985 OR2X1_LOC_91/A OR2X1_LOC_89/A 0.13fF
C3688 AND2X1_LOC_707/a_8_24# OR2X1_LOC_91/A 0.03fF
C3867 OR2X1_LOC_91/A AND2X1_LOC_727/A 0.01fF
C3901 OR2X1_LOC_91/A OR2X1_LOC_95/Y 0.08fF
C5034 OR2X1_LOC_70/Y OR2X1_LOC_91/A 0.69fF
C6539 OR2X1_LOC_91/A OR2X1_LOC_16/A 0.05fF
C6658 AND2X1_LOC_168/Y OR2X1_LOC_91/A 0.02fF
C6799 OR2X1_LOC_91/A AND2X1_LOC_687/Y 0.11fF
C7045 OR2X1_LOC_132/Y OR2X1_LOC_91/A 0.26fF
C7643 OR2X1_LOC_91/A AND2X1_LOC_729/B 0.07fF
C8152 AND2X1_LOC_227/Y OR2X1_LOC_91/A 0.03fF
C8196 OR2X1_LOC_91/A OR2X1_LOC_813/Y 0.19fF
C8504 OR2X1_LOC_599/A OR2X1_LOC_91/A 0.03fF
C8780 OR2X1_LOC_40/Y OR2X1_LOC_91/A 0.27fF
C8929 OR2X1_LOC_91/A OR2X1_LOC_7/A 0.28fF
C8948 OR2X1_LOC_320/Y OR2X1_LOC_91/A 0.01fF
C9156 OR2X1_LOC_176/a_8_216# OR2X1_LOC_91/A 0.01fF
C9311 OR2X1_LOC_127/Y OR2X1_LOC_91/A 0.10fF
C9594 AND2X1_LOC_707/Y OR2X1_LOC_91/A 0.03fF
C9713 OR2X1_LOC_91/A AND2X1_LOC_841/B 0.07fF
C10025 OR2X1_LOC_589/A OR2X1_LOC_91/A 4.15fF
C10344 OR2X1_LOC_91/A OR2X1_LOC_384/a_8_216# 0.06fF
C11024 OR2X1_LOC_3/Y OR2X1_LOC_91/A 4.30fF
C11798 AND2X1_LOC_99/Y OR2X1_LOC_91/A 0.06fF
C12114 OR2X1_LOC_91/A OR2X1_LOC_766/a_8_216# 0.10fF
C12345 OR2X1_LOC_91/A OR2X1_LOC_64/Y 1.71fF
C13035 OR2X1_LOC_96/Y OR2X1_LOC_91/A 0.05fF
C13222 OR2X1_LOC_91/A OR2X1_LOC_829/Y 0.10fF
C13828 OR2X1_LOC_91/A OR2X1_LOC_321/a_8_216# 0.03fF
C16491 AND2X1_LOC_777/a_8_24# OR2X1_LOC_91/A 0.12fF
C17719 OR2X1_LOC_91/A OR2X1_LOC_278/Y 0.03fF
C18629 OR2X1_LOC_91/A OR2X1_LOC_118/Y 0.03fF
C19828 OR2X1_LOC_604/A OR2X1_LOC_91/A 0.23fF
C19935 OR2X1_LOC_306/Y OR2X1_LOC_91/A 0.03fF
C20219 OR2X1_LOC_176/Y OR2X1_LOC_91/A 0.04fF
C21037 AND2X1_LOC_539/Y OR2X1_LOC_91/A 0.03fF
C21105 AND2X1_LOC_326/B OR2X1_LOC_91/A 0.03fF
C21993 OR2X1_LOC_91/A AND2X1_LOC_434/Y 0.07fF
C24100 AND2X1_LOC_98/a_8_24# OR2X1_LOC_91/A 0.03fF
C24173 OR2X1_LOC_91/A AND2X1_LOC_520/Y 0.10fF
C25144 OR2X1_LOC_91/A AND2X1_LOC_318/Y 0.02fF
C25579 OR2X1_LOC_91/A OR2X1_LOC_597/Y 0.09fF
C27020 AND2X1_LOC_715/A OR2X1_LOC_91/A 0.07fF
C27533 AND2X1_LOC_784/A OR2X1_LOC_91/A 0.10fF
C27992 OR2X1_LOC_91/A OR2X1_LOC_52/B 0.10fF
C28781 OR2X1_LOC_91/A OR2X1_LOC_39/A 0.07fF
C29552 OR2X1_LOC_51/Y OR2X1_LOC_91/A 0.08fF
C32327 OR2X1_LOC_91/A OR2X1_LOC_384/Y 0.02fF
C32383 OR2X1_LOC_518/Y OR2X1_LOC_91/A 0.03fF
C32488 AND2X1_LOC_391/Y OR2X1_LOC_91/A 0.09fF
C33502 OR2X1_LOC_91/A OR2X1_LOC_74/A 0.21fF
C34986 OR2X1_LOC_134/Y OR2X1_LOC_91/A 0.24fF
C35520 OR2X1_LOC_91/A AND2X1_LOC_847/Y 0.01fF
C37259 OR2X1_LOC_485/A OR2X1_LOC_91/A 0.06fF
C37901 AND2X1_LOC_383/a_8_24# OR2X1_LOC_91/A 0.09fF
C38013 OR2X1_LOC_695/a_8_216# OR2X1_LOC_91/A 0.02fF
C38957 OR2X1_LOC_305/a_8_216# OR2X1_LOC_91/A 0.06fF
C40048 AND2X1_LOC_714/B OR2X1_LOC_91/A 0.03fF
C41452 AND2X1_LOC_348/A OR2X1_LOC_91/A 0.05fF
C41838 OR2X1_LOC_125/a_8_216# OR2X1_LOC_91/A 0.03fF
C41929 OR2X1_LOC_314/Y OR2X1_LOC_91/A 0.09fF
C41981 OR2X1_LOC_131/Y OR2X1_LOC_91/A 0.03fF
C42264 VDD OR2X1_LOC_91/A 0.55fF
C42551 OR2X1_LOC_91/A OR2X1_LOC_67/Y 0.03fF
C42844 OR2X1_LOC_91/A OR2X1_LOC_248/Y 0.03fF
C43181 OR2X1_LOC_382/Y OR2X1_LOC_91/A 0.05fF
C43317 OR2X1_LOC_91/A AND2X1_LOC_307/Y 0.03fF
C43518 OR2X1_LOC_494/A OR2X1_LOC_91/A 0.08fF
C43658 OR2X1_LOC_91/A OR2X1_LOC_427/A 0.17fF
C45035 OR2X1_LOC_91/A AND2X1_LOC_116/Y 0.03fF
C45258 OR2X1_LOC_45/B OR2X1_LOC_91/A 0.91fF
C45713 OR2X1_LOC_158/A OR2X1_LOC_91/A 0.68fF
C45773 AND2X1_LOC_98/Y OR2X1_LOC_91/A 0.01fF
C46314 OR2X1_LOC_748/A OR2X1_LOC_91/A 0.02fF
C46640 OR2X1_LOC_132/a_8_216# OR2X1_LOC_91/A 0.03fF
C47345 OR2X1_LOC_111/Y OR2X1_LOC_91/A 0.04fF
C48080 OR2X1_LOC_91/A OR2X1_LOC_316/Y 0.03fF
C48153 AND2X1_LOC_390/B OR2X1_LOC_91/A 0.07fF
C48193 AND2X1_LOC_101/a_8_24# OR2X1_LOC_91/A 0.02fF
C48452 OR2X1_LOC_744/A OR2X1_LOC_91/A 0.14fF
C48734 OR2X1_LOC_91/A OR2X1_LOC_320/a_8_216# 0.02fF
C48819 OR2X1_LOC_694/Y OR2X1_LOC_91/A 0.04fF
C49180 AND2X1_LOC_383/a_36_24# OR2X1_LOC_91/A 0.01fF
C50192 OR2X1_LOC_91/Y OR2X1_LOC_91/A 0.01fF
C50287 OR2X1_LOC_311/Y OR2X1_LOC_91/A 0.03fF
C50750 OR2X1_LOC_91/A AND2X1_LOC_831/Y 0.07fF
C51012 OR2X1_LOC_519/Y OR2X1_LOC_91/A 0.16fF
C51678 OR2X1_LOC_91/A AND2X1_LOC_789/Y 0.02fF
C51949 OR2X1_LOC_91/A OR2X1_LOC_125/Y 0.06fF
C53142 AND2X1_LOC_319/A OR2X1_LOC_91/A 0.03fF
C53287 OR2X1_LOC_91/A AND2X1_LOC_721/A 0.03fF
C53594 OR2X1_LOC_91/A AND2X1_LOC_361/A 0.07fF
C54279 OR2X1_LOC_695/Y OR2X1_LOC_91/A 0.01fF
C54322 AND2X1_LOC_391/a_8_24# OR2X1_LOC_91/A 0.07fF
C54362 OR2X1_LOC_127/a_8_216# OR2X1_LOC_91/A 0.05fF
C54666 AND2X1_LOC_520/a_8_24# OR2X1_LOC_91/A 0.01fF
C55084 OR2X1_LOC_692/Y OR2X1_LOC_91/A 0.10fF
C55122 OR2X1_LOC_600/A OR2X1_LOC_91/A 3.98fF
C55125 AND2X1_LOC_335/Y OR2X1_LOC_91/A 0.03fF
C55230 OR2X1_LOC_91/A OR2X1_LOC_619/Y 0.08fF
C57274 OR2X1_LOC_91/A VSS -4.30fF
C852 AND2X1_LOC_94/Y AND2X1_LOC_825/a_8_24# 0.09fF
C15467 AND2X1_LOC_94/Y OR2X1_LOC_397/Y 0.09fF
C29956 VDD AND2X1_LOC_94/Y 0.40fF
C37222 AND2X1_LOC_94/Y AND2X1_LOC_56/B 0.07fF
C38067 AND2X1_LOC_94/Y OR2X1_LOC_83/A 0.10fF
C49381 AND2X1_LOC_94/Y OR2X1_LOC_240/A 0.07fF
C54838 OR2X1_LOC_3/Y AND2X1_LOC_94/Y 0.01fF
C57593 AND2X1_LOC_94/Y VSS 0.39fF
C314 OR2X1_LOC_492/Y OR2X1_LOC_485/A 0.01fF
C335 OR2X1_LOC_108/a_8_216# OR2X1_LOC_485/A 0.01fF
C910 OR2X1_LOC_485/A OR2X1_LOC_497/Y 0.03fF
C1686 OR2X1_LOC_235/B OR2X1_LOC_485/A 0.09fF
C1760 OR2X1_LOC_485/A AND2X1_LOC_319/A 0.02fF
C1861 OR2X1_LOC_485/A AND2X1_LOC_721/A 0.02fF
C2897 AND2X1_LOC_787/A OR2X1_LOC_485/A 0.03fF
C3036 AND2X1_LOC_532/a_8_24# OR2X1_LOC_485/A 0.03fF
C3753 AND2X1_LOC_729/a_8_24# OR2X1_LOC_485/A 0.02fF
C3788 OR2X1_LOC_485/A OR2X1_LOC_600/A 0.25fF
C3872 OR2X1_LOC_485/A OR2X1_LOC_619/Y 0.03fF
C4338 OR2X1_LOC_485/A AND2X1_LOC_539/a_8_24# 0.01fF
C4597 OR2X1_LOC_331/A OR2X1_LOC_485/A 0.06fF
C4972 OR2X1_LOC_329/Y OR2X1_LOC_485/A 0.01fF
C6130 OR2X1_LOC_485/A OR2X1_LOC_13/B 0.28fF
C6636 OR2X1_LOC_485/A OR2X1_LOC_428/A 0.42fF
C7245 OR2X1_LOC_516/A OR2X1_LOC_485/A 0.03fF
C7253 OR2X1_LOC_485/A AND2X1_LOC_342/Y 0.23fF
C7304 OR2X1_LOC_485/A OR2X1_LOC_279/a_8_216# 0.03fF
C7730 OR2X1_LOC_485/A OR2X1_LOC_89/A 1.49fF
C7943 OR2X1_LOC_485/A AND2X1_LOC_590/a_8_24# 0.16fF
C8003 OR2X1_LOC_167/a_8_216# OR2X1_LOC_485/A 0.01fF
C8473 OR2X1_LOC_491/a_8_216# OR2X1_LOC_485/A 0.01fF
C8584 OR2X1_LOC_45/Y OR2X1_LOC_485/A 0.23fF
C8670 OR2X1_LOC_485/A AND2X1_LOC_727/A 0.03fF
C8696 OR2X1_LOC_485/A OR2X1_LOC_95/Y 0.94fF
C8858 OR2X1_LOC_821/Y OR2X1_LOC_485/A 0.40fF
C8959 OR2X1_LOC_179/Y OR2X1_LOC_485/A 0.01fF
C9435 OR2X1_LOC_485/A AND2X1_LOC_621/Y 0.05fF
C9601 OR2X1_LOC_485/A OR2X1_LOC_71/A 0.54fF
C9915 OR2X1_LOC_70/Y OR2X1_LOC_485/A 9.68fF
C9934 AND2X1_LOC_538/a_8_24# OR2X1_LOC_485/A 0.02fF
C9960 OR2X1_LOC_485/A OR2X1_LOC_184/Y 0.01fF
C11014 OR2X1_LOC_484/Y OR2X1_LOC_485/A 0.56fF
C11102 OR2X1_LOC_246/Y OR2X1_LOC_485/A 0.26fF
C11377 OR2X1_LOC_485/A OR2X1_LOC_16/A 0.07fF
C11420 OR2X1_LOC_108/Y OR2X1_LOC_485/A 0.19fF
C11611 OR2X1_LOC_485/A AND2X1_LOC_687/Y 0.02fF
C12296 OR2X1_LOC_485/A AND2X1_LOC_447/Y 0.12fF
C12364 OR2X1_LOC_109/Y OR2X1_LOC_485/A 0.24fF
C12447 OR2X1_LOC_485/A AND2X1_LOC_729/B 0.08fF
C12861 OR2X1_LOC_485/A OR2X1_LOC_279/a_36_216# 0.01fF
C12918 OR2X1_LOC_485/A AND2X1_LOC_227/Y 0.03fF
C13286 OR2X1_LOC_599/A OR2X1_LOC_485/A 0.04fF
C13567 OR2X1_LOC_40/Y OR2X1_LOC_485/A 0.88fF
C13711 OR2X1_LOC_485/A OR2X1_LOC_7/A 0.34fF
C13771 OR2X1_LOC_485/A OR2X1_LOC_224/a_8_216# 0.01fF
C14001 OR2X1_LOC_822/a_8_216# OR2X1_LOC_485/A 0.01fF
C14213 OR2X1_LOC_485/A OR2X1_LOC_615/Y 0.20fF
C14484 OR2X1_LOC_485/A AND2X1_LOC_841/B 0.03fF
C14793 OR2X1_LOC_589/A OR2X1_LOC_485/A 0.18fF
C14899 OR2X1_LOC_485/A OR2X1_LOC_495/Y 0.03fF
C15772 OR2X1_LOC_3/Y OR2X1_LOC_485/A 0.04fF
C17041 OR2X1_LOC_503/A OR2X1_LOC_485/A 0.01fF
C17103 OR2X1_LOC_485/A OR2X1_LOC_64/Y 5.80fF
C17227 OR2X1_LOC_485/A AND2X1_LOC_247/a_8_24# 0.01fF
C18275 OR2X1_LOC_516/B OR2X1_LOC_485/A 0.23fF
C18414 OR2X1_LOC_485/A AND2X1_LOC_196/Y 0.15fF
C18713 AND2X1_LOC_456/B OR2X1_LOC_485/A 0.06fF
C19506 OR2X1_LOC_822/a_36_216# OR2X1_LOC_485/A 0.02fF
C19516 OR2X1_LOC_494/Y OR2X1_LOC_485/A 0.01fF
C19741 OR2X1_LOC_485/A OR2X1_LOC_311/a_8_216# 0.01fF
C20460 OR2X1_LOC_485/A AND2X1_LOC_624/A 0.03fF
C20814 OR2X1_LOC_485/A AND2X1_LOC_434/a_8_24# 0.01fF
C21501 OR2X1_LOC_485/A OR2X1_LOC_172/a_8_216# 0.01fF
C21607 OR2X1_LOC_485/A OR2X1_LOC_312/a_8_216# 0.02fF
C21772 OR2X1_LOC_485/A AND2X1_LOC_114/a_8_24# 0.08fF
C22617 OR2X1_LOC_485/A OR2X1_LOC_278/Y 0.06fF
C23077 OR2X1_LOC_485/A OR2X1_LOC_601/Y 0.01fF
C23101 OR2X1_LOC_485/A OR2X1_LOC_754/A 0.08fF
C23252 OR2X1_LOC_485/A OR2X1_LOC_142/Y 0.02fF
C23503 OR2X1_LOC_485/A OR2X1_LOC_238/Y 0.03fF
C24575 OR2X1_LOC_177/Y OR2X1_LOC_485/A 0.03fF
C24603 OR2X1_LOC_604/A OR2X1_LOC_485/A 1.10fF
C25121 OR2X1_LOC_485/A AND2X1_LOC_447/a_8_24# 0.01fF
C25333 OR2X1_LOC_485/A OR2X1_LOC_183/a_8_216# 0.01fF
C25484 OR2X1_LOC_485/A OR2X1_LOC_164/Y 0.03fF
C25766 AND2X1_LOC_539/Y OR2X1_LOC_485/A 0.04fF
C26720 OR2X1_LOC_485/A AND2X1_LOC_434/Y 0.24fF
C27285 AND2X1_LOC_196/a_8_24# OR2X1_LOC_485/A 0.08fF
C27660 AND2X1_LOC_342/a_8_24# OR2X1_LOC_485/A 0.02fF
C28267 OR2X1_LOC_485/A OR2X1_LOC_248/A 0.01fF
C28448 OR2X1_LOC_485/A OR2X1_LOC_594/a_8_216# 0.01fF
C28904 OR2X1_LOC_485/A AND2X1_LOC_848/Y 0.03fF
C29657 OR2X1_LOC_597/A OR2X1_LOC_485/A 0.21fF
C29670 OR2X1_LOC_178/Y OR2X1_LOC_485/A 0.01fF
C30056 OR2X1_LOC_485/A OR2X1_LOC_829/A 0.19fF
C30287 OR2X1_LOC_485/A OR2X1_LOC_224/Y 0.01fF
C30300 OR2X1_LOC_485/A OR2X1_LOC_597/Y 0.01fF
C30522 OR2X1_LOC_485/A AND2X1_LOC_508/A 0.09fF
C32238 AND2X1_LOC_729/Y OR2X1_LOC_485/A 0.04fF
C32262 AND2X1_LOC_784/A OR2X1_LOC_485/A 0.07fF
C32403 OR2X1_LOC_485/A OR2X1_LOC_172/Y 0.01fF
C32733 OR2X1_LOC_485/A OR2X1_LOC_52/B 0.08fF
C32994 OR2X1_LOC_485/A OR2X1_LOC_13/a_8_216# 0.02fF
C33165 OR2X1_LOC_280/Y OR2X1_LOC_485/A 0.06fF
C33449 OR2X1_LOC_485/Y OR2X1_LOC_485/A 0.01fF
C33568 OR2X1_LOC_485/A OR2X1_LOC_39/A 0.37fF
C33967 OR2X1_LOC_485/A AND2X1_LOC_593/Y 0.03fF
C34061 OR2X1_LOC_485/A OR2X1_LOC_226/Y 0.01fF
C34287 OR2X1_LOC_485/A OR2X1_LOC_51/Y 0.41fF
C34370 OR2X1_LOC_680/A OR2X1_LOC_485/A 0.48fF
C35129 OR2X1_LOC_178/a_8_216# OR2X1_LOC_485/A 0.01fF
C35141 OR2X1_LOC_485/A AND2X1_LOC_436/Y 0.02fF
C35183 AND2X1_LOC_344/a_8_24# OR2X1_LOC_485/A 0.01fF
C36280 OR2X1_LOC_485/A OR2X1_LOC_183/Y 0.01fF
C36503 OR2X1_LOC_485/A OR2X1_LOC_248/a_8_216# -0.00fF
C36801 OR2X1_LOC_600/a_8_216# OR2X1_LOC_485/A 0.01fF
C37178 OR2X1_LOC_485/A OR2X1_LOC_522/a_8_216# 0.07fF
C37253 AND2X1_LOC_391/Y OR2X1_LOC_485/A 0.03fF
C38222 OR2X1_LOC_485/A OR2X1_LOC_74/A 0.12fF
C39056 OR2X1_LOC_485/A AND2X1_LOC_287/a_8_24# 0.06fF
C39071 OR2X1_LOC_485/A OR2X1_LOC_235/a_8_216# 0.03fF
C39089 OR2X1_LOC_485/A OR2X1_LOC_239/Y 0.04fF
C39544 OR2X1_LOC_485/A OR2X1_LOC_615/a_8_216# 0.14fF
C40046 OR2X1_LOC_485/A OR2X1_LOC_536/a_36_216# 0.01fF
C40298 OR2X1_LOC_485/A OR2X1_LOC_497/a_8_216# 0.02fF
C40632 OR2X1_LOC_485/A AND2X1_LOC_614/a_8_24# 0.01fF
C40659 OR2X1_LOC_485/A OR2X1_LOC_597/a_8_216# 0.01fF
C41251 OR2X1_LOC_485/A OR2X1_LOC_167/Y 0.01fF
C42535 OR2X1_LOC_485/A OR2X1_LOC_420/a_8_216# 0.02fF
C43870 OR2X1_LOC_485/A AND2X1_LOC_537/Y 0.02fF
C44095 OR2X1_LOC_485/A OR2X1_LOC_13/Y 0.01fF
C44555 OR2X1_LOC_526/Y OR2X1_LOC_485/A 0.01fF
C45382 OR2X1_LOC_492/a_8_216# OR2X1_LOC_485/A 0.01fF
C45741 OR2X1_LOC_516/Y OR2X1_LOC_485/A 0.11fF
C46382 AND2X1_LOC_348/A OR2X1_LOC_485/A 0.01fF
C47238 VDD OR2X1_LOC_485/A 0.61fF
C47347 OR2X1_LOC_485/A AND2X1_LOC_447/a_36_24# -0.00fF
C47361 OR2X1_LOC_485/A OR2X1_LOC_491/Y 0.01fF
C47368 OR2X1_LOC_251/Y OR2X1_LOC_485/A 0.03fF
C47464 OR2X1_LOC_485/A OR2X1_LOC_67/Y 0.01fF
C47788 OR2X1_LOC_485/A OR2X1_LOC_248/Y 0.41fF
C48127 OR2X1_LOC_600/Y OR2X1_LOC_485/A 0.01fF
C48226 OR2X1_LOC_485/A OR2X1_LOC_591/A 0.09fF
C48585 OR2X1_LOC_485/A OR2X1_LOC_427/A 14.75fF
C49709 OR2X1_LOC_485/A OR2X1_LOC_184/a_8_216# 0.02fF
C49886 OR2X1_LOC_485/A OR2X1_LOC_45/a_8_216# 0.01fF
C50149 OR2X1_LOC_45/B OR2X1_LOC_485/A 0.10fF
C50339 OR2X1_LOC_485/A OR2X1_LOC_235/a_36_216# 0.01fF
C50606 OR2X1_LOC_158/A OR2X1_LOC_485/A 1.55fF
C50688 OR2X1_LOC_485/A AND2X1_LOC_98/Y 0.16fF
C50707 OR2X1_LOC_485/A OR2X1_LOC_594/Y 0.13fF
C51024 OR2X1_LOC_482/Y OR2X1_LOC_485/A 0.09fF
C52644 OR2X1_LOC_485/A AND2X1_LOC_227/a_8_24# 0.02fF
C52880 AND2X1_LOC_390/B OR2X1_LOC_485/A 0.07fF
C52896 OR2X1_LOC_485/A OR2X1_LOC_431/Y 0.05fF
C53175 OR2X1_LOC_744/A OR2X1_LOC_485/A 0.56fF
C53254 OR2X1_LOC_485/A AND2X1_LOC_840/B 0.12fF
C53288 OR2X1_LOC_485/A OR2X1_LOC_282/a_8_216# 0.07fF
C53730 OR2X1_LOC_485/A OR2X1_LOC_420/Y 0.01fF
C54024 OR2X1_LOC_179/a_8_216# OR2X1_LOC_485/A 0.01fF
C54825 OR2X1_LOC_485/A AND2X1_LOC_285/Y 0.02fF
C54920 OR2X1_LOC_91/Y OR2X1_LOC_485/A 0.10fF
C54977 OR2X1_LOC_417/Y OR2X1_LOC_485/A 0.03fF
C54983 OR2X1_LOC_311/Y OR2X1_LOC_485/A 0.04fF
C54987 OR2X1_LOC_485/A AND2X1_LOC_538/Y 0.01fF
C54990 OR2X1_LOC_485/A OR2X1_LOC_601/a_8_216# 0.02fF
C55276 AND2X1_LOC_330/a_8_24# OR2X1_LOC_485/A 0.17fF
C55311 OR2X1_LOC_494/a_8_216# OR2X1_LOC_485/A 0.01fF
C55801 OR2X1_LOC_485/A AND2X1_LOC_436/B 0.02fF
C57496 OR2X1_LOC_485/A VSS -2.58fF
C11928 OR2X1_LOC_342/B OR2X1_LOC_342/a_8_216# 0.01fF
C28487 OR2X1_LOC_342/B OR2X1_LOC_349/B 0.80fF
C52564 OR2X1_LOC_161/A OR2X1_LOC_342/B 0.01fF
C56451 OR2X1_LOC_342/B VSS -0.07fF
C1290 OR2X1_LOC_669/a_8_216# OR2X1_LOC_278/Y 0.01fF
C4595 OR2X1_LOC_250/Y OR2X1_LOC_278/Y 0.18fF
C4912 OR2X1_LOC_604/A OR2X1_LOC_278/Y 0.05fF
C9376 AND2X1_LOC_848/Y OR2X1_LOC_278/Y 0.03fF
C9394 OR2X1_LOC_283/Y OR2X1_LOC_278/Y 0.05fF
C13348 AND2X1_LOC_216/A OR2X1_LOC_278/Y 0.02fF
C13616 OR2X1_LOC_278/Y AND2X1_LOC_286/Y 0.01fF
C14762 OR2X1_LOC_51/Y OR2X1_LOC_278/Y 2.61fF
C14885 OR2X1_LOC_667/a_8_216# OR2X1_LOC_278/Y 0.01fF
C17713 AND2X1_LOC_391/Y OR2X1_LOC_278/Y 0.12fF
C17828 OR2X1_LOC_669/Y OR2X1_LOC_278/Y 0.02fF
C18757 OR2X1_LOC_74/A OR2X1_LOC_278/Y 0.89fF
C19127 OR2X1_LOC_278/Y AND2X1_LOC_287/Y 0.01fF
C19521 OR2X1_LOC_278/Y AND2X1_LOC_287/a_8_24# 0.01fF
C19558 OR2X1_LOC_235/a_8_216# OR2X1_LOC_278/Y 0.01fF
C27468 VDD OR2X1_LOC_278/Y 0.31fF
C27605 OR2X1_LOC_251/Y OR2X1_LOC_278/Y 1.95fF
C28811 OR2X1_LOC_427/A OR2X1_LOC_278/Y 0.06fF
C30831 OR2X1_LOC_158/A OR2X1_LOC_278/Y 0.03fF
C30900 AND2X1_LOC_98/Y OR2X1_LOC_278/Y 0.04fF
C33142 AND2X1_LOC_101/a_8_24# OR2X1_LOC_278/Y 0.01fF
C33406 OR2X1_LOC_744/A OR2X1_LOC_278/Y 0.03fF
C34173 OR2X1_LOC_821/a_8_216# OR2X1_LOC_278/Y 0.01fF
C35068 AND2X1_LOC_285/Y OR2X1_LOC_278/Y 0.03fF
C35974 OR2X1_LOC_667/Y OR2X1_LOC_278/Y 0.01fF
C36033 OR2X1_LOC_235/Y OR2X1_LOC_278/Y 0.01fF
C38030 OR2X1_LOC_235/B OR2X1_LOC_278/Y 0.03fF
C38258 AND2X1_LOC_721/A OR2X1_LOC_278/Y 0.04fF
C40109 OR2X1_LOC_600/A OR2X1_LOC_278/Y 0.59fF
C40576 AND2X1_LOC_286/a_8_24# OR2X1_LOC_278/Y 0.01fF
C40674 OR2X1_LOC_669/A OR2X1_LOC_278/Y 0.01fF
C41924 AND2X1_LOC_99/a_8_24# OR2X1_LOC_278/Y 0.01fF
C42645 OR2X1_LOC_278/Y OR2X1_LOC_13/B 0.05fF
C43143 OR2X1_LOC_278/Y OR2X1_LOC_428/A 0.02fF
C43758 AND2X1_LOC_105/a_8_24# OR2X1_LOC_278/Y 0.01fF
C44192 OR2X1_LOC_89/A OR2X1_LOC_278/Y 0.03fF
C44847 AND2X1_LOC_287/B OR2X1_LOC_278/Y 0.15fF
C44957 OR2X1_LOC_251/a_8_216# OR2X1_LOC_278/Y 0.01fF
C45144 OR2X1_LOC_95/Y OR2X1_LOC_278/Y 0.03fF
C45317 OR2X1_LOC_821/Y OR2X1_LOC_278/Y 0.26fF
C45890 AND2X1_LOC_668/a_8_24# OR2X1_LOC_278/Y 0.01fF
C46099 OR2X1_LOC_278/Y OR2X1_LOC_71/A 0.17fF
C49426 OR2X1_LOC_106/A OR2X1_LOC_278/Y 0.01fF
C49551 OR2X1_LOC_813/Y OR2X1_LOC_278/Y 0.38fF
C49809 OR2X1_LOC_250/a_8_216# OR2X1_LOC_278/Y 0.01fF
C50128 OR2X1_LOC_40/Y OR2X1_LOC_278/Y 0.03fF
C50284 OR2X1_LOC_7/A OR2X1_LOC_278/Y 0.05fF
C50967 OR2X1_LOC_813/a_8_216# OR2X1_LOC_278/Y 0.01fF
C51951 OR2X1_LOC_278/Y AND2X1_LOC_240/Y 0.02fF
C52389 OR2X1_LOC_3/Y OR2X1_LOC_278/Y 0.02fF
C53138 AND2X1_LOC_99/Y OR2X1_LOC_278/Y 0.01fF
C53704 OR2X1_LOC_64/Y OR2X1_LOC_278/Y 0.10fF
C54035 AND2X1_LOC_101/B OR2X1_LOC_278/Y 0.17fF
C55234 AND2X1_LOC_456/B OR2X1_LOC_278/Y 0.02fF
C56052 OR2X1_LOC_494/Y OR2X1_LOC_278/Y 0.03fF
C56602 OR2X1_LOC_278/Y VSS 0.08fF
C684 AND2X1_LOC_41/A OR2X1_LOC_78/B 0.14fF
C830 AND2X1_LOC_135/a_8_24# OR2X1_LOC_78/B 0.04fF
C1090 AND2X1_LOC_83/a_36_24# OR2X1_LOC_78/B 0.01fF
C1435 OR2X1_LOC_78/B OR2X1_LOC_112/A 0.37fF
C1828 OR2X1_LOC_78/B OR2X1_LOC_71/A 0.03fF
C2266 AND2X1_LOC_31/Y OR2X1_LOC_78/B 0.35fF
C2559 OR2X1_LOC_633/B OR2X1_LOC_78/B 0.03fF
C2699 OR2X1_LOC_78/B OR2X1_LOC_608/Y 0.01fF
C3174 OR2X1_LOC_78/B AND2X1_LOC_36/Y 0.44fF
C3297 OR2X1_LOC_633/a_8_216# OR2X1_LOC_78/B 0.01fF
C3312 OR2X1_LOC_635/A OR2X1_LOC_78/B 0.01fF
C3997 OR2X1_LOC_78/B OR2X1_LOC_535/a_8_216# 0.01fF
C4369 OR2X1_LOC_78/B OR2X1_LOC_537/a_8_216# 0.04fF
C4422 AND2X1_LOC_60/a_8_24# OR2X1_LOC_78/B 0.03fF
C4537 AND2X1_LOC_504/a_8_24# OR2X1_LOC_78/B 0.18fF
C4609 OR2X1_LOC_557/A OR2X1_LOC_78/B 0.06fF
C5389 OR2X1_LOC_78/B OR2X1_LOC_798/a_8_216# 0.01fF
C5409 OR2X1_LOC_78/B OR2X1_LOC_269/B 5.09fF
C5718 AND2X1_LOC_172/a_8_24# OR2X1_LOC_78/B 0.01fF
C5824 OR2X1_LOC_78/B OR2X1_LOC_539/Y 1.55fF
C6511 OR2X1_LOC_770/A OR2X1_LOC_78/B 0.01fF
C6927 OR2X1_LOC_78/B OR2X1_LOC_332/a_8_216# 0.01fF
C6988 OR2X1_LOC_78/B OR2X1_LOC_161/B 4.66fF
C8018 OR2X1_LOC_539/a_8_216# OR2X1_LOC_78/B 0.01fF
C8220 OR2X1_LOC_78/B AND2X1_LOC_609/a_8_24# 0.02fF
C8931 OR2X1_LOC_647/B OR2X1_LOC_78/B 0.07fF
C9398 OR2X1_LOC_401/A OR2X1_LOC_78/B 0.01fF
C9679 OR2X1_LOC_319/B OR2X1_LOC_78/B 0.04fF
C9697 OR2X1_LOC_318/Y OR2X1_LOC_78/B 0.03fF
C11007 OR2X1_LOC_287/B OR2X1_LOC_78/B 0.06fF
C11105 OR2X1_LOC_436/Y OR2X1_LOC_78/B 0.04fF
C11394 OR2X1_LOC_78/B OR2X1_LOC_799/a_8_216# 0.01fF
C12134 OR2X1_LOC_151/A OR2X1_LOC_78/B 5.67fF
C15435 OR2X1_LOC_78/B OR2X1_LOC_537/a_36_216# 0.02fF
C15484 OR2X1_LOC_61/A OR2X1_LOC_78/B 0.03fF
C15620 AND2X1_LOC_601/a_8_24# OR2X1_LOC_78/B 0.08fF
C15918 OR2X1_LOC_78/B OR2X1_LOC_390/A 0.03fF
C16161 OR2X1_LOC_168/A OR2X1_LOC_78/B 0.02fF
C16465 OR2X1_LOC_243/A OR2X1_LOC_78/B 0.08fF
C16775 AND2X1_LOC_229/a_8_24# OR2X1_LOC_78/B 0.13fF
C17409 AND2X1_LOC_135/a_36_24# OR2X1_LOC_78/B 0.01fF
C17806 OR2X1_LOC_193/A OR2X1_LOC_78/B 0.44fF
C17987 OR2X1_LOC_78/B OR2X1_LOC_339/A 0.19fF
C18091 AND2X1_LOC_505/a_8_24# OR2X1_LOC_78/B 0.03fF
C18578 AND2X1_LOC_39/a_8_24# OR2X1_LOC_78/B 0.02fF
C19379 OR2X1_LOC_715/B OR2X1_LOC_78/B 0.10fF
C19914 OR2X1_LOC_656/B OR2X1_LOC_78/B 0.10fF
C19921 AND2X1_LOC_767/a_8_24# OR2X1_LOC_78/B 0.01fF
C19952 OR2X1_LOC_793/A OR2X1_LOC_78/B 0.02fF
C20015 AND2X1_LOC_45/a_8_24# OR2X1_LOC_78/B 0.05fF
C20347 OR2X1_LOC_687/Y OR2X1_LOC_78/B 0.19fF
C20429 OR2X1_LOC_401/B OR2X1_LOC_78/B 0.01fF
C20656 OR2X1_LOC_535/A OR2X1_LOC_78/B 0.12fF
C21120 OR2X1_LOC_78/A OR2X1_LOC_78/B 1.11fF
C22266 OR2X1_LOC_78/B OR2X1_LOC_854/A 0.21fF
C22407 AND2X1_LOC_396/a_8_24# OR2X1_LOC_78/B 0.01fF
C22417 AND2X1_LOC_172/a_36_24# OR2X1_LOC_78/B 0.01fF
C22436 OR2X1_LOC_538/A OR2X1_LOC_78/B 0.03fF
C22520 OR2X1_LOC_78/B OR2X1_LOC_802/A 0.01fF
C23664 OR2X1_LOC_507/A OR2X1_LOC_78/B 0.01fF
C23815 OR2X1_LOC_646/A OR2X1_LOC_78/B 0.01fF
C25299 OR2X1_LOC_186/Y OR2X1_LOC_78/B 0.12fF
C25404 OR2X1_LOC_773/B OR2X1_LOC_78/B 0.01fF
C25419 AND2X1_LOC_81/B OR2X1_LOC_78/B 0.01fF
C25565 OR2X1_LOC_112/B OR2X1_LOC_78/B 0.23fF
C25705 AND2X1_LOC_765/a_8_24# OR2X1_LOC_78/B 0.03fF
C25866 OR2X1_LOC_574/A OR2X1_LOC_78/B 0.03fF
C26214 AND2X1_LOC_58/a_8_24# OR2X1_LOC_78/B 0.01fF
C26227 AND2X1_LOC_16/a_8_24# OR2X1_LOC_78/B 0.05fF
C26489 OR2X1_LOC_78/B OR2X1_LOC_539/B 0.01fF
C26679 OR2X1_LOC_375/A OR2X1_LOC_78/B 0.81fF
C26975 OR2X1_LOC_78/B OR2X1_LOC_549/A 0.37fF
C28800 OR2X1_LOC_673/Y OR2X1_LOC_78/B 0.07fF
C29495 OR2X1_LOC_139/A OR2X1_LOC_78/B 0.03fF
C30915 OR2X1_LOC_703/B OR2X1_LOC_78/B 0.37fF
C30932 OR2X1_LOC_87/A OR2X1_LOC_78/B 0.70fF
C31013 AND2X1_LOC_45/a_36_24# OR2X1_LOC_78/B 0.01fF
C31701 OR2X1_LOC_61/B OR2X1_LOC_78/B -0.01fF
C31724 OR2X1_LOC_194/B OR2X1_LOC_78/B 0.01fF
C31982 OR2X1_LOC_97/A OR2X1_LOC_78/B 0.03fF
C32055 OR2X1_LOC_78/B OR2X1_LOC_78/a_8_216# 0.02fF
C32418 OR2X1_LOC_691/Y OR2X1_LOC_78/B 0.03fF
C33047 OR2X1_LOC_333/B OR2X1_LOC_78/B 0.03fF
C33441 OR2X1_LOC_154/A OR2X1_LOC_78/B 0.38fF
C33873 AND2X1_LOC_395/a_8_24# OR2X1_LOC_78/B 0.01fF
C34191 AND2X1_LOC_20/a_8_24# OR2X1_LOC_78/B 0.01fF
C34542 OR2X1_LOC_78/B OR2X1_LOC_633/A 0.02fF
C35011 AND2X1_LOC_82/Y OR2X1_LOC_78/B 0.10fF
C36253 OR2X1_LOC_614/Y OR2X1_LOC_78/B 0.11fF
C36824 OR2X1_LOC_33/B OR2X1_LOC_78/B 0.01fF
C37159 OR2X1_LOC_100/Y OR2X1_LOC_78/B 0.04fF
C37187 AND2X1_LOC_16/a_36_24# OR2X1_LOC_78/B 0.02fF
C37322 OR2X1_LOC_532/B OR2X1_LOC_78/B 0.36fF
C37565 OR2X1_LOC_78/B OR2X1_LOC_78/a_36_216# 0.01fF
C38441 AND2X1_LOC_503/a_8_24# OR2X1_LOC_78/B 0.05fF
C38885 OR2X1_LOC_798/Y OR2X1_LOC_78/B 0.05fF
C39255 VDD OR2X1_LOC_78/B 2.12fF
C40070 OR2X1_LOC_676/Y OR2X1_LOC_78/B 0.57fF
C40498 AND2X1_LOC_83/a_8_24# OR2X1_LOC_78/B 0.03fF
C41436 OR2X1_LOC_840/A OR2X1_LOC_78/B 1.52fF
C41813 AND2X1_LOC_754/a_8_24# OR2X1_LOC_78/B 0.03fF
C41933 OR2X1_LOC_802/Y OR2X1_LOC_78/B 0.06fF
C42272 OR2X1_LOC_809/B OR2X1_LOC_78/B 0.14fF
C42359 OR2X1_LOC_160/A OR2X1_LOC_78/B 0.34fF
C42434 AND2X1_LOC_86/B OR2X1_LOC_78/B 0.12fF
C42446 OR2X1_LOC_624/B OR2X1_LOC_78/B 0.08fF
C42673 OR2X1_LOC_196/Y OR2X1_LOC_78/B 0.03fF
C42785 OR2X1_LOC_447/A OR2X1_LOC_78/B 0.16fF
C43172 OR2X1_LOC_78/B OR2X1_LOC_78/Y 1.43fF
C43637 OR2X1_LOC_608/a_8_216# OR2X1_LOC_78/B 0.03fF
C43668 OR2X1_LOC_185/A OR2X1_LOC_78/B 0.36fF
C43787 AND2X1_LOC_431/a_8_24# OR2X1_LOC_78/B 0.03fF
C44473 OR2X1_LOC_802/a_8_216# OR2X1_LOC_78/B 0.01fF
C44848 OR2X1_LOC_78/B OR2X1_LOC_641/A 0.07fF
C45374 OR2X1_LOC_168/a_8_216# OR2X1_LOC_78/B 0.06fF
C46118 AND2X1_LOC_91/B OR2X1_LOC_78/B 0.17fF
C46271 OR2X1_LOC_799/A OR2X1_LOC_78/B 0.03fF
C46522 OR2X1_LOC_78/B OR2X1_LOC_446/B 0.01fF
C46770 AND2X1_LOC_56/B OR2X1_LOC_78/B 0.09fF
C47677 OR2X1_LOC_389/B OR2X1_LOC_78/B 0.05fF
C48219 AND2X1_LOC_47/Y OR2X1_LOC_78/B 0.26fF
C48393 OR2X1_LOC_78/B OR2X1_LOC_646/B 0.05fF
C48506 OR2X1_LOC_506/A OR2X1_LOC_78/B 0.03fF
C49118 OR2X1_LOC_78/B OR2X1_LOC_788/B 0.04fF
C49696 OR2X1_LOC_78/B AND2X1_LOC_232/a_8_24# -0.00fF
C49733 OR2X1_LOC_509/A OR2X1_LOC_78/B 0.02fF
C50118 OR2X1_LOC_235/B OR2X1_LOC_78/B 0.07fF
C51241 OR2X1_LOC_78/B OR2X1_LOC_771/B 0.11fF
C51715 AND2X1_LOC_766/a_8_24# OR2X1_LOC_78/B 0.01fF
C52127 OR2X1_LOC_78/B AND2X1_LOC_44/Y 2.48fF
C53045 OR2X1_LOC_78/B AND2X1_LOC_18/Y 0.65fF
C53317 OR2X1_LOC_78/B OR2X1_LOC_789/A 0.03fF
C53439 OR2X1_LOC_112/a_8_216# OR2X1_LOC_78/B 0.01fF
C53966 OR2X1_LOC_130/A OR2X1_LOC_78/B 0.11fF
C54101 OR2X1_LOC_78/B AND2X1_LOC_39/Y 0.01fF
C54407 OR2X1_LOC_449/B OR2X1_LOC_78/B 0.06fF
C54915 AND2X1_LOC_431/a_36_24# OR2X1_LOC_78/B 0.01fF
C55210 AND2X1_LOC_503/a_36_24# OR2X1_LOC_78/B 0.01fF
C56078 OR2X1_LOC_240/B OR2X1_LOC_78/B 0.05fF
C56085 OR2X1_LOC_78/B OR2X1_LOC_161/A 0.11fF
C56203 AND2X1_LOC_51/Y OR2X1_LOC_78/B 0.31fF
C56757 OR2X1_LOC_78/B VSS 0.54fF
C8 OR2X1_LOC_605/B OR2X1_LOC_161/A 0.01fF
C148 OR2X1_LOC_161/A OR2X1_LOC_515/Y 0.16fF
C260 OR2X1_LOC_161/A OR2X1_LOC_549/A 0.03fF
C645 OR2X1_LOC_161/A OR2X1_LOC_161/a_8_216# 0.01fF
C1026 OR2X1_LOC_161/A OR2X1_LOC_348/B 0.03fF
C1217 AND2X1_LOC_311/a_36_24# OR2X1_LOC_161/A 0.01fF
C1818 OR2X1_LOC_779/Y OR2X1_LOC_161/A 0.01fF
C2785 OR2X1_LOC_161/A OR2X1_LOC_712/B 0.04fF
C2841 OR2X1_LOC_139/A OR2X1_LOC_161/A 0.07fF
C3447 OR2X1_LOC_307/a_36_216# OR2X1_LOC_161/A 0.01fF
C3587 OR2X1_LOC_161/A OR2X1_LOC_259/B 0.02fF
C4149 AND2X1_LOC_526/a_8_24# OR2X1_LOC_161/A 0.01fF
C4189 OR2X1_LOC_668/a_8_216# OR2X1_LOC_161/A 0.01fF
C4214 OR2X1_LOC_703/B OR2X1_LOC_161/A 0.03fF
C4219 OR2X1_LOC_87/A OR2X1_LOC_161/A 0.28fF
C4423 OR2X1_LOC_161/A OR2X1_LOC_844/B 0.02fF
C4519 OR2X1_LOC_389/A OR2X1_LOC_161/A 0.01fF
C5222 OR2X1_LOC_161/A OR2X1_LOC_349/B 0.01fF
C5284 OR2X1_LOC_97/A OR2X1_LOC_161/A 0.03fF
C5728 OR2X1_LOC_691/Y OR2X1_LOC_161/A 0.03fF
C6063 OR2X1_LOC_161/A OR2X1_LOC_546/A 0.01fF
C6756 OR2X1_LOC_154/A OR2X1_LOC_161/A 0.27fF
C7588 OR2X1_LOC_538/a_8_216# OR2X1_LOC_161/A 0.04fF
C8188 AND2X1_LOC_107/a_8_24# OR2X1_LOC_161/A 0.01fF
C8795 OR2X1_LOC_161/A OR2X1_LOC_342/A 0.02fF
C9025 AND2X1_LOC_677/a_8_24# OR2X1_LOC_161/A 0.02fF
C9636 OR2X1_LOC_161/A OR2X1_LOC_779/A 0.03fF
C9670 OR2X1_LOC_614/Y OR2X1_LOC_161/A 0.03fF
C10744 OR2X1_LOC_532/B OR2X1_LOC_161/A 0.24fF
C10928 OR2X1_LOC_440/B OR2X1_LOC_161/A 0.04fF
C11395 OR2X1_LOC_114/a_8_216# OR2X1_LOC_161/A 0.01fF
C12652 VDD OR2X1_LOC_161/A 2.66fF
C13343 OR2X1_LOC_161/A AND2X1_LOC_418/a_8_24# 0.01fF
C13421 OR2X1_LOC_161/A OR2X1_LOC_523/A 0.01fF
C13514 OR2X1_LOC_676/Y OR2X1_LOC_161/A 0.07fF
C14705 OR2X1_LOC_161/A OR2X1_LOC_115/B 0.12fF
C14823 OR2X1_LOC_840/A OR2X1_LOC_161/A 0.10fF
C14870 AND2X1_LOC_145/a_8_24# OR2X1_LOC_161/A 0.01fF
C15605 OR2X1_LOC_809/B OR2X1_LOC_161/A 0.07fF
C15669 OR2X1_LOC_160/A OR2X1_LOC_161/A 3.92fF
C16229 AND2X1_LOC_108/a_8_24# OR2X1_LOC_161/A 0.01fF
C16945 OR2X1_LOC_161/A OR2X1_LOC_708/Y 0.03fF
C16986 OR2X1_LOC_185/A OR2X1_LOC_161/A 0.09fF
C17441 OR2X1_LOC_702/A OR2X1_LOC_161/A 0.03fF
C18285 OR2X1_LOC_114/Y OR2X1_LOC_161/A 0.03fF
C18700 OR2X1_LOC_161/A OR2X1_LOC_541/B 0.02fF
C18859 OR2X1_LOC_161/A OR2X1_LOC_446/A 0.02fF
C19156 OR2X1_LOC_778/Y OR2X1_LOC_161/A 0.04fF
C19218 OR2X1_LOC_113/A OR2X1_LOC_161/A 0.01fF
C19383 AND2X1_LOC_91/B OR2X1_LOC_161/A 0.11fF
C19749 OR2X1_LOC_161/A OR2X1_LOC_446/B 1.34fF
C19752 OR2X1_LOC_161/A OR2X1_LOC_303/B 0.06fF
C19904 OR2X1_LOC_542/B OR2X1_LOC_161/A 0.03fF
C20007 AND2X1_LOC_56/B OR2X1_LOC_161/A 0.07fF
C21143 AND2X1_LOC_745/a_8_24# OR2X1_LOC_161/A 0.11fF
C21405 AND2X1_LOC_47/Y OR2X1_LOC_161/A 11.54fF
C21535 OR2X1_LOC_161/A OR2X1_LOC_186/a_8_216# 0.01fF
C21575 AND2X1_LOC_521/a_8_24# OR2X1_LOC_161/A 0.01fF
C21698 OR2X1_LOC_506/A OR2X1_LOC_161/A 0.07fF
C21842 OR2X1_LOC_161/A OR2X1_LOC_284/B 0.03fF
C21932 OR2X1_LOC_161/A OR2X1_LOC_180/B 0.03fF
C22349 OR2X1_LOC_161/A OR2X1_LOC_788/B 0.05fF
C22871 OR2X1_LOC_161/A OR2X1_LOC_162/A 0.01fF
C23353 OR2X1_LOC_235/B OR2X1_LOC_161/A 1.50fF
C23774 OR2X1_LOC_703/A OR2X1_LOC_161/A 0.20fF
C24143 OR2X1_LOC_161/A OR2X1_LOC_362/A 0.02fF
C24219 OR2X1_LOC_539/A OR2X1_LOC_161/A 0.01fF
C24867 OR2X1_LOC_161/A OR2X1_LOC_593/B 0.06fF
C25342 OR2X1_LOC_161/A AND2X1_LOC_44/Y 0.30fF
C25896 OR2X1_LOC_148/B OR2X1_LOC_161/A 0.01fF
C26153 OR2X1_LOC_161/A AND2X1_LOC_258/a_8_24# 0.01fF
C26167 OR2X1_LOC_161/A OR2X1_LOC_708/a_8_216# 0.04fF
C26217 OR2X1_LOC_161/A AND2X1_LOC_18/Y 0.15fF
C26610 OR2X1_LOC_161/A OR2X1_LOC_307/A 0.02fF
C26979 OR2X1_LOC_161/A OR2X1_LOC_186/a_36_216# 0.02fF
C27043 OR2X1_LOC_523/B OR2X1_LOC_161/A 0.01fF
C27611 OR2X1_LOC_449/B OR2X1_LOC_161/A 0.10fF
C28956 OR2X1_LOC_447/Y OR2X1_LOC_161/A 0.07fF
C29149 OR2X1_LOC_346/A OR2X1_LOC_161/A 0.02fF
C29347 AND2X1_LOC_51/Y OR2X1_LOC_161/A 0.68fF
C29694 OR2X1_LOC_161/A OR2X1_LOC_541/a_8_216# 0.14fF
C30069 AND2X1_LOC_41/A OR2X1_LOC_161/A 0.46fF
C30149 OR2X1_LOC_631/B OR2X1_LOC_161/A 0.03fF
C30188 AND2X1_LOC_135/a_8_24# OR2X1_LOC_161/A -0.06fF
C30729 OR2X1_LOC_161/A OR2X1_LOC_112/A 0.01fF
C30887 OR2X1_LOC_284/a_8_216# OR2X1_LOC_161/A 0.01fF
C30920 OR2X1_LOC_756/Y OR2X1_LOC_161/A 0.01fF
C31416 AND2X1_LOC_701/a_8_24# OR2X1_LOC_161/A 0.04fF
C31556 AND2X1_LOC_31/Y OR2X1_LOC_161/A 0.18fF
C32328 OR2X1_LOC_161/A OR2X1_LOC_451/B 0.03fF
C32413 OR2X1_LOC_161/A AND2X1_LOC_36/Y 1.02fF
C32675 OR2X1_LOC_346/B OR2X1_LOC_161/A 0.12fF
C33004 AND2X1_LOC_167/a_8_24# OR2X1_LOC_161/A 0.06fF
C33054 OR2X1_LOC_128/B OR2X1_LOC_161/A 0.36fF
C33333 AND2X1_LOC_522/a_8_24# OR2X1_LOC_161/A 0.01fF
C33755 OR2X1_LOC_308/A OR2X1_LOC_161/A 0.01fF
C33795 OR2X1_LOC_161/A OR2X1_LOC_160/Y 0.56fF
C34801 OR2X1_LOC_161/A OR2X1_LOC_269/B 0.29fF
C34881 AND2X1_LOC_146/a_8_24# OR2X1_LOC_161/A 0.01fF
C35163 OR2X1_LOC_161/A OR2X1_LOC_347/B 0.12fF
C35184 OR2X1_LOC_161/A OR2X1_LOC_779/a_8_216# 0.03fF
C35372 OR2X1_LOC_161/A OR2X1_LOC_319/Y 0.01fF
C35806 OR2X1_LOC_161/A OR2X1_LOC_777/B 0.09fF
C36294 OR2X1_LOC_161/A OR2X1_LOC_161/B 0.58fF
C36412 AND2X1_LOC_536/a_8_24# OR2X1_LOC_161/A 0.03fF
C37105 OR2X1_LOC_161/A OR2X1_LOC_259/A 0.03fF
C37581 OR2X1_LOC_161/A OR2X1_LOC_777/a_8_216# 0.03fF
C38956 OR2X1_LOC_319/B OR2X1_LOC_161/A 0.12fF
C38974 OR2X1_LOC_318/Y OR2X1_LOC_161/A 0.01fF
C39062 OR2X1_LOC_296/Y OR2X1_LOC_161/A 0.02fF
C39406 AND2X1_LOC_173/a_36_24# OR2X1_LOC_161/A 0.01fF
C39892 OR2X1_LOC_629/A OR2X1_LOC_161/A 0.04fF
C40309 OR2X1_LOC_76/A OR2X1_LOC_161/A 0.02fF
C40346 OR2X1_LOC_148/A OR2X1_LOC_161/A 0.01fF
C40680 OR2X1_LOC_161/A OR2X1_LOC_553/A 0.14fF
C40693 OR2X1_LOC_161/A OR2X1_LOC_779/a_36_216# 0.01fF
C41423 OR2X1_LOC_151/A OR2X1_LOC_161/A 1.02fF
C41913 OR2X1_LOC_287/A OR2X1_LOC_161/A -0.01fF
C41934 AND2X1_LOC_757/a_8_24# OR2X1_LOC_161/A 0.01fF
C43111 OR2X1_LOC_161/A OR2X1_LOC_168/Y 0.03fF
C43188 OR2X1_LOC_161/A OR2X1_LOC_777/a_36_216# 0.01fF
C43440 AND2X1_LOC_497/a_8_24# OR2X1_LOC_161/A 0.01fF
C44126 AND2X1_LOC_125/a_8_24# OR2X1_LOC_161/A 0.01fF
C44392 OR2X1_LOC_161/A OR2X1_LOC_301/a_8_216# 0.01fF
C44604 OR2X1_LOC_664/Y OR2X1_LOC_161/A 0.03fF
C44790 OR2X1_LOC_161/A OR2X1_LOC_342/a_8_216# 0.01fF
C44979 OR2X1_LOC_448/A OR2X1_LOC_161/A 0.01fF
C45091 OR2X1_LOC_446/a_8_216# OR2X1_LOC_161/A 0.07fF
C45322 OR2X1_LOC_161/A OR2X1_LOC_706/a_8_216# 0.05fF
C45630 AND2X1_LOC_280/a_8_24# OR2X1_LOC_161/A 0.01fF
C45905 OR2X1_LOC_161/A OR2X1_LOC_668/Y 0.12fF
C46283 AND2X1_LOC_311/a_8_24# OR2X1_LOC_161/A 0.02fF
C46709 OR2X1_LOC_190/A OR2X1_LOC_161/A 0.03fF
C46955 OR2X1_LOC_161/A OR2X1_LOC_241/B 0.01fF
C47097 OR2X1_LOC_188/Y OR2X1_LOC_161/A 0.02fF
C47591 OR2X1_LOC_831/A OR2X1_LOC_161/A 0.02fF
C47667 OR2X1_LOC_791/A OR2X1_LOC_161/A 0.09fF
C47956 OR2X1_LOC_710/A OR2X1_LOC_161/A 0.02fF
C48017 OR2X1_LOC_161/A OR2X1_LOC_356/A 0.11fF
C48587 OR2X1_LOC_810/A OR2X1_LOC_161/A 0.03fF
C48588 OR2X1_LOC_307/a_8_216# OR2X1_LOC_161/A 0.03fF
C48850 OR2X1_LOC_715/B OR2X1_LOC_161/A 0.10fF
C48856 OR2X1_LOC_161/A AND2X1_LOC_626/a_8_24# 0.23fF
C48865 OR2X1_LOC_161/A OR2X1_LOC_784/B 0.01fF
C49794 AND2X1_LOC_167/a_36_24# OR2X1_LOC_161/A 0.01fF
C49850 OR2X1_LOC_687/Y OR2X1_LOC_161/A 0.15fF
C50115 OR2X1_LOC_535/A OR2X1_LOC_161/A 0.01fF
C50592 OR2X1_LOC_78/A OR2X1_LOC_161/A 2.17fF
C50743 OR2X1_LOC_605/A OR2X1_LOC_161/A 0.01fF
C51425 OR2X1_LOC_501/B OR2X1_LOC_161/A 0.03fF
C51655 OR2X1_LOC_161/A OR2X1_LOC_318/B 0.02fF
C51669 OR2X1_LOC_161/A OR2X1_LOC_854/A 0.03fF
C51824 OR2X1_LOC_114/B OR2X1_LOC_161/A 0.06fF
C51865 OR2X1_LOC_538/A OR2X1_LOC_161/A 0.07fF
C53173 OR2X1_LOC_833/B OR2X1_LOC_161/A 0.04fF
C54019 OR2X1_LOC_448/Y OR2X1_LOC_161/A 0.48fF
C54320 OR2X1_LOC_161/A OR2X1_LOC_629/B 0.51fF
C54718 OR2X1_LOC_186/Y OR2X1_LOC_161/A 0.36fF
C54947 OR2X1_LOC_196/B OR2X1_LOC_161/A 0.07fF
C55353 OR2X1_LOC_574/A OR2X1_LOC_161/A 0.07fF
C55561 OR2X1_LOC_161/A AND2X1_LOC_627/a_8_24# 0.17fF
C55712 OR2X1_LOC_319/a_8_216# OR2X1_LOC_161/A 0.03fF
C56136 OR2X1_LOC_448/a_8_216# OR2X1_LOC_161/A 0.04fF
C56194 OR2X1_LOC_375/A OR2X1_LOC_161/A 0.15fF
C56749 OR2X1_LOC_161/A VSS 1.43fF
C757 AND2X1_LOC_41/A OR2X1_LOC_375/A 1.98fF
C1094 AND2X1_LOC_41/A OR2X1_LOC_549/A 0.14fF
C1935 AND2X1_LOC_229/a_36_24# AND2X1_LOC_41/A 0.01fF
C3641 OR2X1_LOC_139/A AND2X1_LOC_41/A 0.29fF
C4508 OR2X1_LOC_834/a_8_216# AND2X1_LOC_41/A 0.01fF
C4629 AND2X1_LOC_41/A AND2X1_LOC_697/a_8_24# 0.04fF
C4647 AND2X1_LOC_41/A AND2X1_LOC_666/a_8_24# 0.10fF
C4991 AND2X1_LOC_41/A OR2X1_LOC_87/A 0.23fF
C5294 OR2X1_LOC_389/A AND2X1_LOC_41/A 0.01fF
C5651 AND2X1_LOC_41/A OR2X1_LOC_130/a_8_216# 0.01fF
C5799 AND2X1_LOC_41/A OR2X1_LOC_61/B 0.09fF
C6062 AND2X1_LOC_41/A AND2X1_LOC_239/a_8_24# 0.01fF
C6120 OR2X1_LOC_97/A AND2X1_LOC_41/A 0.03fF
C6189 AND2X1_LOC_41/A OR2X1_LOC_541/A 0.09fF
C6538 OR2X1_LOC_691/Y AND2X1_LOC_41/A 0.03fF
C6553 AND2X1_LOC_41/A OR2X1_LOC_713/A 1.05fF
C6914 AND2X1_LOC_41/A OR2X1_LOC_546/A 0.26fF
C7035 AND2X1_LOC_700/a_8_24# AND2X1_LOC_41/A 0.02fF
C7190 OR2X1_LOC_333/B AND2X1_LOC_41/A 0.03fF
C7597 OR2X1_LOC_154/A AND2X1_LOC_41/A 0.46fF
C7612 AND2X1_LOC_41/A OR2X1_LOC_267/A 0.05fF
C7649 AND2X1_LOC_41/A OR2X1_LOC_778/A 0.02fF
C7778 AND2X1_LOC_41/A OR2X1_LOC_198/A 0.04fF
C8045 AND2X1_LOC_41/A OR2X1_LOC_267/a_8_216# 0.01fF
C8153 AND2X1_LOC_41/A AND2X1_LOC_821/a_8_24# 0.03fF
C8747 AND2X1_LOC_41/A OR2X1_LOC_267/Y 0.01fF
C10059 OR2X1_LOC_124/B AND2X1_LOC_41/A 0.01fF
C10451 AND2X1_LOC_41/A OR2X1_LOC_779/A 0.03fF
C11539 AND2X1_LOC_41/A OR2X1_LOC_532/B 0.07fF
C12596 OR2X1_LOC_710/B AND2X1_LOC_41/A 0.03fF
C13470 VDD AND2X1_LOC_41/A 1.00fF
C14306 OR2X1_LOC_676/Y AND2X1_LOC_41/A 0.12fF
C14330 OR2X1_LOC_834/A AND2X1_LOC_41/A 0.02fF
C15592 OR2X1_LOC_840/A AND2X1_LOC_41/A 0.01fF
C16011 OR2X1_LOC_216/A AND2X1_LOC_41/A 0.03fF
C16093 AND2X1_LOC_385/a_8_24# AND2X1_LOC_41/A 0.03fF
C16264 AND2X1_LOC_41/A OR2X1_LOC_750/Y 0.04fF
C16479 OR2X1_LOC_160/A AND2X1_LOC_41/A 0.93fF
C16749 AND2X1_LOC_41/A OR2X1_LOC_130/Y 0.01fF
C17738 OR2X1_LOC_185/A AND2X1_LOC_41/A 0.03fF
C18935 AND2X1_LOC_41/A OR2X1_LOC_294/Y 0.09fF
C18950 AND2X1_LOC_41/A OR2X1_LOC_641/A 0.02fF
C19478 AND2X1_LOC_41/A OR2X1_LOC_541/B 0.02fF
C19967 OR2X1_LOC_643/A AND2X1_LOC_41/A 0.03fF
C19976 AND2X1_LOC_41/A OR2X1_LOC_778/Y 0.10fF
C20213 AND2X1_LOC_91/B AND2X1_LOC_41/A 0.06fF
C20308 OR2X1_LOC_308/a_8_216# AND2X1_LOC_41/A 0.02fF
C20579 AND2X1_LOC_41/A OR2X1_LOC_446/B 0.07fF
C20802 AND2X1_LOC_41/A AND2X1_LOC_56/B 1.56fF
C21317 AND2X1_LOC_41/A AND2X1_LOC_666/a_36_24# 0.01fF
C21543 OR2X1_LOC_790/A AND2X1_LOC_41/A 0.02fF
C21686 OR2X1_LOC_389/B AND2X1_LOC_41/A 0.03fF
C21849 AND2X1_LOC_41/A AND2X1_LOC_751/a_8_24# 0.03fF
C22214 AND2X1_LOC_41/A AND2X1_LOC_47/Y 0.22fF
C22512 AND2X1_LOC_41/A OR2X1_LOC_506/A 0.31fF
C25260 AND2X1_LOC_41/A OR2X1_LOC_776/A 0.17fF
C25364 OR2X1_LOC_678/a_8_216# AND2X1_LOC_41/A 0.02fF
C25686 OR2X1_LOC_506/a_8_216# AND2X1_LOC_41/A 0.01fF
C26139 AND2X1_LOC_41/A AND2X1_LOC_44/Y 0.40fF
C26353 AND2X1_LOC_41/A OR2X1_LOC_720/B 0.03fF
C26825 AND2X1_LOC_41/A OR2X1_LOC_506/B 0.01fF
C27021 AND2X1_LOC_41/A AND2X1_LOC_18/Y 3.61fF
C27314 AND2X1_LOC_41/A OR2X1_LOC_789/A 0.03fF
C27416 AND2X1_LOC_41/A OR2X1_LOC_307/A 0.01fF
C27964 AND2X1_LOC_41/A OR2X1_LOC_130/A 0.21fF
C28422 AND2X1_LOC_41/A OR2X1_LOC_449/B 0.07fF
C29759 AND2X1_LOC_41/A OR2X1_LOC_447/Y 0.07fF
C30063 OR2X1_LOC_790/B AND2X1_LOC_41/A 0.12fF
C30148 AND2X1_LOC_41/A AND2X1_LOC_51/Y 0.61fF
C30477 AND2X1_LOC_41/A OR2X1_LOC_541/a_8_216# 0.06fF
C30956 OR2X1_LOC_631/B AND2X1_LOC_41/A 0.04fF
C31603 OR2X1_LOC_149/B AND2X1_LOC_41/A 0.18fF
C32315 AND2X1_LOC_41/A AND2X1_LOC_31/Y 0.10fF
C32616 AND2X1_LOC_597/a_8_24# AND2X1_LOC_41/A 0.01fF
C32630 AND2X1_LOC_385/a_36_24# AND2X1_LOC_41/A 0.01fF
C32992 AND2X1_LOC_41/A AND2X1_LOC_305/a_8_24# -0.01fF
C33256 AND2X1_LOC_41/A AND2X1_LOC_36/Y 0.62fF
C33299 OR2X1_LOC_506/Y AND2X1_LOC_41/A 0.07fF
C34154 OR2X1_LOC_856/A AND2X1_LOC_41/A 0.05fF
C34523 OR2X1_LOC_308/A AND2X1_LOC_41/A 0.01fF
C34677 AND2X1_LOC_504/a_8_24# AND2X1_LOC_41/A 0.04fF
C35580 AND2X1_LOC_41/A OR2X1_LOC_269/B 0.28fF
C36591 AND2X1_LOC_41/A OR2X1_LOC_777/B 0.09fF
C36628 OR2X1_LOC_188/a_8_216# AND2X1_LOC_41/A -0.02fF
C36839 AND2X1_LOC_41/A AND2X1_LOC_13/a_8_24# 0.04fF
C37048 OR2X1_LOC_198/a_8_216# AND2X1_LOC_41/A 0.05fF
C37084 AND2X1_LOC_41/A OR2X1_LOC_161/B 0.81fF
C37199 AND2X1_LOC_536/a_8_24# AND2X1_LOC_41/A 0.08fF
C37711 AND2X1_LOC_41/A AND2X1_LOC_67/Y 0.45fF
C38073 OR2X1_LOC_644/B AND2X1_LOC_41/A 0.01fF
C38246 AND2X1_LOC_41/A OR2X1_LOC_705/B 0.31fF
C38961 AND2X1_LOC_41/A OR2X1_LOC_790/a_8_216# 0.02fF
C39847 AND2X1_LOC_41/A OR2X1_LOC_296/Y 0.01fF
C40156 OR2X1_LOC_507/B AND2X1_LOC_41/A 0.01fF
C40656 OR2X1_LOC_147/a_8_216# AND2X1_LOC_41/A 0.01fF
C40764 AND2X1_LOC_41/A OR2X1_LOC_473/A 0.05fF
C41505 AND2X1_LOC_41/A OR2X1_LOC_553/A 0.08fF
C42246 OR2X1_LOC_151/A AND2X1_LOC_41/A 0.07fF
C42322 AND2X1_LOC_41/A AND2X1_LOC_67/a_8_24# 0.02fF
C44779 AND2X1_LOC_41/A OR2X1_LOC_308/Y 0.13fF
C45829 AND2X1_LOC_504/a_36_24# AND2X1_LOC_41/A 0.01fF
C45967 AND2X1_LOC_41/A AND2X1_LOC_7/Y 0.03fF
C46156 AND2X1_LOC_41/A OR2X1_LOC_706/a_8_216# 0.01fF
C46165 AND2X1_LOC_41/A OR2X1_LOC_390/A 0.03fF
C47066 AND2X1_LOC_229/a_8_24# AND2X1_LOC_41/A 0.08fF
C47816 AND2X1_LOC_41/A OR2X1_LOC_241/B 0.41fF
C47932 OR2X1_LOC_188/Y AND2X1_LOC_41/A 0.01fF
C48183 AND2X1_LOC_41/A OR2X1_LOC_193/A 0.01fF
C48362 OR2X1_LOC_208/A AND2X1_LOC_41/A 0.03fF
C48524 OR2X1_LOC_537/A AND2X1_LOC_41/A 0.03fF
C48755 OR2X1_LOC_710/A AND2X1_LOC_41/A 0.01fF
C49388 AND2X1_LOC_41/A OR2X1_LOC_810/A 0.03fF
C49673 OR2X1_LOC_715/B AND2X1_LOC_41/A 0.03fF
C50177 OR2X1_LOC_656/B AND2X1_LOC_41/A 0.02fF
C50222 AND2X1_LOC_41/A OR2X1_LOC_793/A 0.01fF
C50301 AND2X1_LOC_41/A AND2X1_LOC_45/a_8_24# 0.02fF
C50631 OR2X1_LOC_687/Y AND2X1_LOC_41/A 0.07fF
C51378 AND2X1_LOC_41/A OR2X1_LOC_78/A 0.92fF
C52248 OR2X1_LOC_147/B AND2X1_LOC_41/A 0.75fF
C52592 OR2X1_LOC_121/Y AND2X1_LOC_41/A 0.01fF
C53539 AND2X1_LOC_41/A OR2X1_LOC_623/B 0.07fF
C53665 AND2X1_LOC_41/A AND2X1_LOC_13/a_36_24# 0.01fF
C53882 OR2X1_LOC_507/A AND2X1_LOC_41/A 0.64fF
C53953 AND2X1_LOC_41/A OR2X1_LOC_833/B 0.19fF
C54353 AND2X1_LOC_321/a_8_24# AND2X1_LOC_41/A 0.10fF
C55683 AND2X1_LOC_81/B AND2X1_LOC_41/A 0.05fF
C55787 AND2X1_LOC_41/A OR2X1_LOC_196/B 0.07fF
C56179 OR2X1_LOC_574/A AND2X1_LOC_41/A 0.05fF
C57435 AND2X1_LOC_41/A VSS 0.69fF
C265 OR2X1_LOC_848/A OR2X1_LOC_489/A 0.01fF
C805 OR2X1_LOC_848/A OR2X1_LOC_772/B 0.03fF
C836 OR2X1_LOC_489/B OR2X1_LOC_848/A 0.01fF
C15288 OR2X1_LOC_848/B OR2X1_LOC_848/A 0.47fF
C17008 OR2X1_LOC_773/B OR2X1_LOC_848/A 0.01fF
C19164 OR2X1_LOC_391/B OR2X1_LOC_848/A 0.40fF
C19223 OR2X1_LOC_848/A OR2X1_LOC_846/A 0.09fF
C27764 OR2X1_LOC_848/A OR2X1_LOC_557/a_8_216# 0.02fF
C28327 OR2X1_LOC_770/B OR2X1_LOC_848/A 0.17fF
C29233 OR2X1_LOC_848/A OR2X1_LOC_391/A 0.19fF
C30899 VDD OR2X1_LOC_848/A 0.27fF
C33605 OR2X1_LOC_848/A OR2X1_LOC_846/B 0.04fF
C38754 OR2X1_LOC_848/A OR2X1_LOC_561/B 0.40fF
C40190 OR2X1_LOC_848/A OR2X1_LOC_391/a_8_216# 0.02fF
C42681 OR2X1_LOC_848/A OR2X1_LOC_771/B 0.01fF
C43764 OR2X1_LOC_848/A OR2X1_LOC_848/a_8_216# 0.06fF
C45867 OR2X1_LOC_848/A OR2X1_LOC_391/a_36_216# 0.01fF
C45871 OR2X1_LOC_848/A OR2X1_LOC_489/a_8_216# 0.02fF
C51470 OR2X1_LOC_848/A OR2X1_LOC_392/A 0.01fF
C52418 OR2X1_LOC_848/A OR2X1_LOC_557/A 0.01fF
C53237 OR2X1_LOC_848/A OR2X1_LOC_269/B 0.01fF
C54283 OR2X1_LOC_770/A OR2X1_LOC_848/A 0.09fF
C54863 OR2X1_LOC_846/a_8_216# OR2X1_LOC_848/A 0.03fF
C57552 OR2X1_LOC_848/A VSS -4.79fF
C43 AND2X1_LOC_727/A OR2X1_LOC_39/A 0.03fF
C74 OR2X1_LOC_95/Y OR2X1_LOC_39/A 0.14fF
C815 AND2X1_LOC_621/Y OR2X1_LOC_39/A 0.15fF
C1043 OR2X1_LOC_39/A OR2X1_LOC_71/A 0.86fF
C1340 OR2X1_LOC_70/Y OR2X1_LOC_39/A 1.89fF
C1385 OR2X1_LOC_504/Y OR2X1_LOC_39/A 0.43fF
C1417 OR2X1_LOC_437/Y OR2X1_LOC_39/A 0.38fF
C2505 OR2X1_LOC_484/Y OR2X1_LOC_39/A 0.23fF
C2866 OR2X1_LOC_16/A OR2X1_LOC_39/A 0.10fF
C2905 OR2X1_LOC_108/Y OR2X1_LOC_39/A 0.19fF
C3824 OR2X1_LOC_109/Y OR2X1_LOC_39/A 0.05fF
C4163 OR2X1_LOC_39/Y OR2X1_LOC_39/A 0.06fF
C4656 OR2X1_LOC_599/A OR2X1_LOC_39/A 0.07fF
C4925 OR2X1_LOC_40/Y OR2X1_LOC_39/A 0.18fF
C5078 OR2X1_LOC_7/A OR2X1_LOC_39/A 0.13fF
C5497 OR2X1_LOC_32/a_8_216# OR2X1_LOC_39/A 0.01fF
C5552 AND2X1_LOC_115/a_8_24# OR2X1_LOC_39/A 0.02fF
C5595 OR2X1_LOC_615/Y OR2X1_LOC_39/A 0.03fF
C6186 OR2X1_LOC_589/A OR2X1_LOC_39/A 0.02fF
C6272 OR2X1_LOC_495/Y OR2X1_LOC_39/A 0.07fF
C6378 OR2X1_LOC_60/a_8_216# OR2X1_LOC_39/A 0.03fF
C7250 OR2X1_LOC_3/Y OR2X1_LOC_39/A 0.18fF
C7265 AND2X1_LOC_631/Y OR2X1_LOC_39/A 0.03fF
C7610 OR2X1_LOC_74/Y OR2X1_LOC_39/A 0.04fF
C8123 OR2X1_LOC_280/a_8_216# OR2X1_LOC_39/A 0.04fF
C8533 OR2X1_LOC_393/a_36_216# OR2X1_LOC_39/A 0.03fF
C8624 OR2X1_LOC_64/Y OR2X1_LOC_39/A 0.10fF
C9761 OR2X1_LOC_516/B OR2X1_LOC_39/A 0.28fF
C11130 AND2X1_LOC_116/B OR2X1_LOC_39/A 0.01fF
C11533 AND2X1_LOC_154/Y OR2X1_LOC_39/A 0.04fF
C11866 OR2X1_LOC_521/Y OR2X1_LOC_39/A 0.02fF
C11898 AND2X1_LOC_624/A OR2X1_LOC_39/A 0.06fF
C13645 OR2X1_LOC_612/B OR2X1_LOC_39/A 0.03fF
C14120 OR2X1_LOC_273/Y OR2X1_LOC_39/A 0.03fF
C14170 OR2X1_LOC_75/Y OR2X1_LOC_39/A 0.03fF
C14260 OR2X1_LOC_39/A OR2X1_LOC_504/a_8_216# 0.01fF
C14302 OR2X1_LOC_744/a_8_216# OR2X1_LOC_39/A 0.01fF
C14675 OR2X1_LOC_39/A OR2X1_LOC_142/Y 0.02fF
C14867 OR2X1_LOC_118/Y OR2X1_LOC_39/A 0.02fF
C14921 OR2X1_LOC_238/Y OR2X1_LOC_39/A 0.06fF
C15056 OR2X1_LOC_39/A OR2X1_LOC_39/a_8_216# 0.09fF
C15385 OR2X1_LOC_503/Y OR2X1_LOC_39/A 0.01fF
C15983 OR2X1_LOC_177/Y OR2X1_LOC_39/A 0.05fF
C16015 OR2X1_LOC_604/A OR2X1_LOC_39/A 0.42fF
C16554 OR2X1_LOC_39/A OR2X1_LOC_265/Y 0.07fF
C16957 OR2X1_LOC_164/Y OR2X1_LOC_39/A 0.01fF
C17044 AND2X1_LOC_155/Y OR2X1_LOC_39/A 0.01fF
C17076 AND2X1_LOC_633/Y OR2X1_LOC_39/A 0.03fF
C17334 OR2X1_LOC_612/Y OR2X1_LOC_39/A 0.01fF
C17397 OR2X1_LOC_237/a_8_216# OR2X1_LOC_39/A 0.04fF
C17473 OR2X1_LOC_60/a_36_216# OR2X1_LOC_39/A 0.02fF
C17623 OR2X1_LOC_316/a_8_216# OR2X1_LOC_39/A 0.01fF
C17706 OR2X1_LOC_20/Y OR2X1_LOC_39/A 0.10fF
C18428 OR2X1_LOC_595/Y OR2X1_LOC_39/A 0.05fF
C18643 OR2X1_LOC_674/a_8_216# OR2X1_LOC_39/A 0.06fF
C18682 OR2X1_LOC_837/B OR2X1_LOC_39/A 0.03fF
C18736 OR2X1_LOC_69/a_8_216# OR2X1_LOC_39/A 0.03fF
C19494 OR2X1_LOC_837/Y OR2X1_LOC_39/A 0.07fF
C19941 OR2X1_LOC_517/a_8_216# OR2X1_LOC_39/A 0.02fF
C20395 AND2X1_LOC_520/Y OR2X1_LOC_39/A 0.05fF
C20419 AND2X1_LOC_186/a_8_24# OR2X1_LOC_39/A 0.01fF
C23017 OR2X1_LOC_237/a_36_216# OR2X1_LOC_39/A 0.01fF
C23320 AND2X1_LOC_715/A OR2X1_LOC_39/A 0.02fF
C23845 AND2X1_LOC_729/Y OR2X1_LOC_39/A 0.05fF
C23864 AND2X1_LOC_784/A OR2X1_LOC_39/A 0.10fF
C24288 OR2X1_LOC_39/A OR2X1_LOC_52/B 0.11fF
C24716 OR2X1_LOC_280/Y OR2X1_LOC_39/A 0.09fF
C24963 OR2X1_LOC_485/Y OR2X1_LOC_39/A 0.05fF
C25347 OR2X1_LOC_744/Y OR2X1_LOC_39/A 0.23fF
C25800 OR2X1_LOC_51/Y OR2X1_LOC_39/A 0.22fF
C25836 OR2X1_LOC_58/a_8_216# OR2X1_LOC_39/A 0.01fF
C25899 OR2X1_LOC_680/A OR2X1_LOC_39/A 7.79fF
C26342 OR2X1_LOC_626/a_8_216# OR2X1_LOC_39/A 0.01fF
C28456 OR2X1_LOC_237/Y OR2X1_LOC_39/A 0.06fF
C28708 OR2X1_LOC_39/A OR2X1_LOC_522/a_8_216# 0.03fF
C29268 OR2X1_LOC_32/B OR2X1_LOC_39/A 0.09fF
C29715 OR2X1_LOC_69/a_36_216# OR2X1_LOC_39/A 0.02fF
C29755 OR2X1_LOC_74/A OR2X1_LOC_39/A 0.28fF
C30036 OR2X1_LOC_39/A OR2X1_LOC_626/Y 0.34fF
C30930 OR2X1_LOC_517/a_36_216# OR2X1_LOC_39/A 0.01fF
C31394 AND2X1_LOC_633/a_8_24# OR2X1_LOC_39/A 0.01fF
C31709 OR2X1_LOC_505/Y OR2X1_LOC_39/A 0.09fF
C32600 OR2X1_LOC_697/Y OR2X1_LOC_39/A 0.03fF
C33060 OR2X1_LOC_595/a_8_216# OR2X1_LOC_39/A 0.02fF
C33398 OR2X1_LOC_58/Y OR2X1_LOC_39/A 0.04fF
C33952 OR2X1_LOC_495/a_8_216# OR2X1_LOC_39/A 0.02fF
C34035 OR2X1_LOC_238/a_8_216# OR2X1_LOC_39/A 0.02fF
C34190 OR2X1_LOC_39/A OR2X1_LOC_522/a_36_216# 0.01fF
C34354 OR2X1_LOC_32/Y OR2X1_LOC_39/A 0.23fF
C35192 OR2X1_LOC_69/Y OR2X1_LOC_39/A 0.06fF
C35385 OR2X1_LOC_39/A OR2X1_LOC_743/Y 0.01fF
C36704 OR2X1_LOC_492/a_8_216# OR2X1_LOC_39/A 0.09fF
C37077 OR2X1_LOC_516/Y OR2X1_LOC_39/A 1.95fF
C37784 OR2X1_LOC_472/B OR2X1_LOC_39/A 0.15fF
C38464 VDD OR2X1_LOC_39/A 6.30fF
C38550 OR2X1_LOC_315/Y OR2X1_LOC_39/A 0.03fF
C38717 OR2X1_LOC_39/A OR2X1_LOC_67/Y 0.03fF
C38904 OR2X1_LOC_60/Y OR2X1_LOC_39/A 0.02fF
C39447 OR2X1_LOC_462/B OR2X1_LOC_39/A 0.17fF
C39831 OR2X1_LOC_427/A OR2X1_LOC_39/A 0.24fF
C40329 OR2X1_LOC_416/Y OR2X1_LOC_39/A 0.01fF
C41392 OR2X1_LOC_45/B OR2X1_LOC_39/A 0.29fF
C41877 OR2X1_LOC_158/A OR2X1_LOC_39/A 0.20fF
C42317 OR2X1_LOC_482/Y OR2X1_LOC_39/A 0.15fF
C44170 OR2X1_LOC_316/Y OR2X1_LOC_39/A 0.01fF
C44290 OR2X1_LOC_416/a_8_216# OR2X1_LOC_39/A 0.01fF
C44521 OR2X1_LOC_744/A OR2X1_LOC_39/A 1.56fF
C44621 AND2X1_LOC_840/B OR2X1_LOC_39/A 0.11fF
C44634 OR2X1_LOC_74/a_8_216# OR2X1_LOC_39/A 0.04fF
C45331 OR2X1_LOC_39/A OR2X1_LOC_522/Y 0.02fF
C45926 AND2X1_LOC_56/B OR2X1_LOC_39/A 3.56fF
C46369 OR2X1_LOC_91/Y OR2X1_LOC_39/A 0.17fF
C46446 OR2X1_LOC_527/Y OR2X1_LOC_39/A 0.35fF
C46464 OR2X1_LOC_291/Y OR2X1_LOC_39/A 0.05fF
C46621 OR2X1_LOC_39/A AND2X1_LOC_780/a_8_24# 0.01fF
C46875 AND2X1_LOC_276/Y OR2X1_LOC_39/A 0.02fF
C47293 AND2X1_LOC_139/B OR2X1_LOC_39/A 0.07fF
C48028 OR2X1_LOC_492/Y OR2X1_LOC_39/A 0.16fF
C48180 OR2X1_LOC_517/Y OR2X1_LOC_39/A 0.04fF
C48583 OR2X1_LOC_497/Y OR2X1_LOC_39/A 0.04fF
C48836 OR2X1_LOC_39/A AND2X1_LOC_249/a_8_24# 0.01fF
C48964 OR2X1_LOC_109/a_8_216# OR2X1_LOC_39/A 0.30fF
C49348 OR2X1_LOC_235/B OR2X1_LOC_39/A 0.01fF
C50514 AND2X1_LOC_787/A OR2X1_LOC_39/A 0.05fF
C51403 OR2X1_LOC_612/a_8_216# OR2X1_LOC_39/A 0.06fF
C51408 OR2X1_LOC_600/A OR2X1_LOC_39/A 0.13fF
C51482 OR2X1_LOC_619/Y OR2X1_LOC_39/A 0.71fF
C52157 OR2X1_LOC_39/A AND2X1_LOC_783/B 0.01fF
C52259 OR2X1_LOC_331/A OR2X1_LOC_39/A 0.43fF
C52628 OR2X1_LOC_505/a_8_216# OR2X1_LOC_39/A 0.01fF
C53605 OR2X1_LOC_393/a_8_216# OR2X1_LOC_39/A 0.05fF
C53832 OR2X1_LOC_39/A OR2X1_LOC_13/B 0.84fF
C54282 OR2X1_LOC_39/A OR2X1_LOC_428/A 0.05fF
C54295 OR2X1_LOC_39/A OR2X1_LOC_595/A 0.03fF
C54446 AND2X1_LOC_154/a_8_24# OR2X1_LOC_39/A 0.01fF
C54748 OR2X1_LOC_528/Y OR2X1_LOC_39/A 0.04fF
C54850 OR2X1_LOC_516/A OR2X1_LOC_39/A 0.01fF
C55363 OR2X1_LOC_89/A OR2X1_LOC_39/A 1.14fF
C55379 OR2X1_LOC_461/Y OR2X1_LOC_39/A 0.09fF
C55536 OR2X1_LOC_39/A AND2X1_LOC_590/a_8_24# 0.02fF
C55997 AND2X1_LOC_473/Y OR2X1_LOC_39/A 0.05fF
C56532 OR2X1_LOC_39/A VSS 1.02fF
C216 OR2X1_LOC_382/Y OR2X1_LOC_158/A 0.01fF
C9653 OR2X1_LOC_382/Y OR2X1_LOC_600/A 0.03fF
C12555 OR2X1_LOC_382/Y OR2X1_LOC_428/A 0.02fF
C13617 OR2X1_LOC_382/Y OR2X1_LOC_89/A 0.01fF
C19400 OR2X1_LOC_382/Y OR2X1_LOC_40/Y 0.01fF
C21718 OR2X1_LOC_382/Y OR2X1_LOC_3/Y 0.03fF
C30397 OR2X1_LOC_382/Y OR2X1_LOC_604/A 0.11fF
C43034 OR2X1_LOC_382/Y OR2X1_LOC_384/Y 0.08fF
C52254 OR2X1_LOC_382/Y AND2X1_LOC_348/A 0.11fF
C53064 OR2X1_LOC_382/Y VDD 0.23fF
C58058 OR2X1_LOC_382/Y VSS 0.18fF
C973 OR2X1_LOC_428/A OR2X1_LOC_183/Y 0.02fF
C1551 OR2X1_LOC_237/Y OR2X1_LOC_428/A 0.01fF
C1789 OR2X1_LOC_384/Y OR2X1_LOC_428/A 0.68fF
C1857 OR2X1_LOC_522/a_8_216# OR2X1_LOC_428/A 0.01fF
C1916 AND2X1_LOC_391/Y OR2X1_LOC_428/A 0.01fF
C2681 OR2X1_LOC_428/A OR2X1_LOC_423/Y 0.01fF
C2894 AND2X1_LOC_673/a_8_24# OR2X1_LOC_428/A 0.01fF
C2914 OR2X1_LOC_74/A OR2X1_LOC_428/A 0.07fF
C3618 AND2X1_LOC_448/a_8_24# OR2X1_LOC_428/A 0.01fF
C4787 OR2X1_LOC_106/Y OR2X1_LOC_428/A 0.02fF
C4882 AND2X1_LOC_847/Y OR2X1_LOC_428/A 0.01fF
C5459 AND2X1_LOC_319/a_8_24# OR2X1_LOC_428/A 0.03fF
C5747 OR2X1_LOC_670/a_8_216# OR2X1_LOC_428/A 0.01fF
C6070 AND2X1_LOC_362/B OR2X1_LOC_428/A 0.06fF
C6229 OR2X1_LOC_431/a_8_216# OR2X1_LOC_428/A 0.04fF
C6480 AND2X1_LOC_706/Y OR2X1_LOC_428/A 0.07fF
C7364 AND2X1_LOC_383/a_8_24# OR2X1_LOC_428/A 0.04fF
C8410 OR2X1_LOC_305/a_8_216# OR2X1_LOC_428/A 0.06fF
C8492 AND2X1_LOC_537/Y OR2X1_LOC_428/A 0.07fF
C8722 AND2X1_LOC_285/a_8_24# OR2X1_LOC_428/A 0.08fF
C8724 OR2X1_LOC_13/Y OR2X1_LOC_428/A 0.03fF
C8788 OR2X1_LOC_700/Y OR2X1_LOC_428/A 0.02fF
C8902 OR2X1_LOC_295/Y OR2X1_LOC_428/A 0.04fF
C9213 OR2X1_LOC_433/Y OR2X1_LOC_428/A 0.03fF
C9563 AND2X1_LOC_714/B OR2X1_LOC_428/A 0.12fF
C10310 OR2X1_LOC_428/A OR2X1_LOC_589/a_8_216# 0.04fF
C10347 AND2X1_LOC_798/a_8_24# OR2X1_LOC_428/A 0.05fF
C11044 AND2X1_LOC_798/A OR2X1_LOC_428/A 0.07fF
C11239 OR2X1_LOC_125/a_8_216# OR2X1_LOC_428/A 0.01fF
C11679 VDD OR2X1_LOC_428/A 1.89fF
C11789 OR2X1_LOC_251/Y OR2X1_LOC_428/A 0.02fF
C12690 AND2X1_LOC_307/Y OR2X1_LOC_428/A 0.05fF
C12930 OR2X1_LOC_494/A OR2X1_LOC_428/A 0.01fF
C13033 OR2X1_LOC_427/A OR2X1_LOC_428/A 0.28fF
C13873 OR2X1_LOC_281/a_8_216# OR2X1_LOC_428/A 0.15fF
C14631 OR2X1_LOC_45/B OR2X1_LOC_428/A 0.20fF
C14684 OR2X1_LOC_292/a_8_216# OR2X1_LOC_428/A 0.02fF
C15063 OR2X1_LOC_158/A OR2X1_LOC_428/A 1.02fF
C15108 OR2X1_LOC_103/Y OR2X1_LOC_428/A 0.04fF
C15126 OR2X1_LOC_103/a_8_216# OR2X1_LOC_428/A 0.14fF
C15521 OR2X1_LOC_586/Y OR2X1_LOC_428/A 0.07fF
C15569 OR2X1_LOC_748/A OR2X1_LOC_428/A 0.04fF
C15613 OR2X1_LOC_304/Y OR2X1_LOC_428/A 0.53fF
C16586 AND2X1_LOC_848/A OR2X1_LOC_428/A 0.02fF
C17263 OR2X1_LOC_316/Y OR2X1_LOC_428/A 0.02fF
C17311 AND2X1_LOC_390/B OR2X1_LOC_428/A 0.07fF
C17336 OR2X1_LOC_431/Y OR2X1_LOC_428/A 0.02fF
C17578 OR2X1_LOC_309/Y OR2X1_LOC_428/A 0.12fF
C17599 OR2X1_LOC_744/A OR2X1_LOC_428/A 0.12fF
C18206 AND2X1_LOC_308/a_8_24# OR2X1_LOC_428/A 0.04fF
C18438 AND2X1_LOC_383/a_36_24# OR2X1_LOC_428/A 0.02fF
C18453 OR2X1_LOC_522/Y OR2X1_LOC_428/A 0.01fF
C19414 OR2X1_LOC_91/Y OR2X1_LOC_428/A 0.03fF
C19427 OR2X1_LOC_305/Y OR2X1_LOC_428/A 0.04fF
C19476 OR2X1_LOC_417/Y OR2X1_LOC_428/A 0.03fF
C19489 OR2X1_LOC_311/Y OR2X1_LOC_428/A 0.06fF
C19980 AND2X1_LOC_831/Y OR2X1_LOC_428/A 0.12fF
C20266 AND2X1_LOC_436/B OR2X1_LOC_428/A 0.72fF
C20595 OR2X1_LOC_135/a_8_216# OR2X1_LOC_428/A 0.03fF
C20979 OR2X1_LOC_428/A AND2X1_LOC_789/Y 0.04fF
C21222 OR2X1_LOC_125/Y OR2X1_LOC_428/A 0.04fF
C21259 OR2X1_LOC_409/B OR2X1_LOC_428/A 0.03fF
C22431 AND2X1_LOC_319/A OR2X1_LOC_428/A 0.04fF
C22611 AND2X1_LOC_721/A OR2X1_LOC_428/A 0.04fF
C23646 AND2X1_LOC_391/a_8_24# OR2X1_LOC_428/A 0.01fF
C23677 OR2X1_LOC_127/a_8_216# OR2X1_LOC_428/A 0.02fF
C24440 OR2X1_LOC_600/A OR2X1_LOC_428/A 0.18fF
C24486 OR2X1_LOC_619/Y OR2X1_LOC_428/A 0.10fF
C24957 AND2X1_LOC_454/A OR2X1_LOC_428/A 0.39fF
C25709 OR2X1_LOC_292/Y OR2X1_LOC_428/A 0.01fF
C26631 OR2X1_LOC_312/Y OR2X1_LOC_428/A 0.09fF
C26675 AND2X1_LOC_307/a_8_24# OR2X1_LOC_428/A 0.03fF
C26847 OR2X1_LOC_428/A OR2X1_LOC_13/B 0.53fF
C27953 AND2X1_LOC_712/B OR2X1_LOC_428/A 0.01fF
C28355 OR2X1_LOC_89/A OR2X1_LOC_428/A 0.09fF
C29105 OR2X1_LOC_45/Y OR2X1_LOC_428/A 0.09fF
C29217 AND2X1_LOC_727/A OR2X1_LOC_428/A 0.06fF
C29258 OR2X1_LOC_95/Y OR2X1_LOC_428/A 0.11fF
C30455 OR2X1_LOC_70/Y OR2X1_LOC_428/A 0.26fF
C31525 OR2X1_LOC_428/A OR2X1_LOC_759/Y 0.03fF
C31594 AND2X1_LOC_535/Y OR2X1_LOC_428/A 0.07fF
C31947 OR2X1_LOC_16/A OR2X1_LOC_428/A 0.10fF
C31962 OR2X1_LOC_108/Y OR2X1_LOC_428/A 0.02fF
C32811 OR2X1_LOC_428/A OR2X1_LOC_759/a_8_216# 0.06fF
C32905 OR2X1_LOC_109/Y OR2X1_LOC_428/A 0.03fF
C32913 AND2X1_LOC_448/Y OR2X1_LOC_428/A 0.07fF
C32991 AND2X1_LOC_729/B OR2X1_LOC_428/A 0.03fF
C33498 AND2X1_LOC_227/Y OR2X1_LOC_428/A 0.02fF
C33557 OR2X1_LOC_41/Y OR2X1_LOC_428/A 0.30fF
C33805 OR2X1_LOC_599/A OR2X1_LOC_428/A 0.03fF
C34113 OR2X1_LOC_40/Y OR2X1_LOC_428/A 0.69fF
C34218 OR2X1_LOC_7/A OR2X1_LOC_428/A 0.27fF
C34591 OR2X1_LOC_127/Y OR2X1_LOC_428/A 0.01fF
C34701 AND2X1_LOC_115/a_8_24# OR2X1_LOC_428/A 0.16fF
C34710 AND2X1_LOC_308/a_36_24# OR2X1_LOC_428/A 0.01fF
C34946 AND2X1_LOC_707/Y OR2X1_LOC_428/A 0.10fF
C35339 OR2X1_LOC_589/A OR2X1_LOC_428/A 0.12fF
C35686 OR2X1_LOC_384/a_8_216# OR2X1_LOC_428/A 0.01fF
C36346 OR2X1_LOC_3/Y OR2X1_LOC_428/A 0.43fF
C37160 OR2X1_LOC_280/a_8_216# OR2X1_LOC_428/A 0.01fF
C37623 OR2X1_LOC_64/Y OR2X1_LOC_428/A 0.67fF
C37627 AND2X1_LOC_307/a_36_24# OR2X1_LOC_428/A 0.01fF
C38316 OR2X1_LOC_96/Y OR2X1_LOC_428/A 0.01fF
C39228 AND2X1_LOC_456/B OR2X1_LOC_428/A 0.02fF
C40017 OR2X1_LOC_494/Y OR2X1_LOC_428/A 0.75fF
C40171 AND2X1_LOC_116/B OR2X1_LOC_428/A 0.06fF
C40426 AND2X1_LOC_802/Y OR2X1_LOC_428/A 0.05fF
C40916 OR2X1_LOC_521/Y OR2X1_LOC_428/A 0.02fF
C41327 AND2X1_LOC_434/a_8_24# OR2X1_LOC_428/A 0.08fF
C41937 AND2X1_LOC_635/a_8_24# OR2X1_LOC_428/A 0.08fF
C42311 OR2X1_LOC_670/Y OR2X1_LOC_428/A 0.03fF
C42812 OR2X1_LOC_295/a_8_216# OR2X1_LOC_428/A 0.14fF
C43065 OR2X1_LOC_421/Y OR2X1_LOC_428/A 0.01fF
C45234 OR2X1_LOC_604/A OR2X1_LOC_428/A 0.31fF
C45325 OR2X1_LOC_306/Y OR2X1_LOC_428/A 0.05fF
C46525 AND2X1_LOC_539/Y OR2X1_LOC_428/A 0.03fF
C46578 AND2X1_LOC_711/A OR2X1_LOC_428/A 0.02fF
C46580 AND2X1_LOC_326/B OR2X1_LOC_428/A 0.03fF
C46638 OR2X1_LOC_237/a_8_216# OR2X1_LOC_428/A 0.05fF
C47064 AND2X1_LOC_319/a_36_24# OR2X1_LOC_428/A 0.01fF
C47505 AND2X1_LOC_434/Y OR2X1_LOC_428/A 0.14fF
C49599 OR2X1_LOC_135/Y OR2X1_LOC_428/A 0.03fF
C49630 AND2X1_LOC_98/a_8_24# OR2X1_LOC_428/A 0.01fF
C49689 AND2X1_LOC_848/Y OR2X1_LOC_428/A 0.03fF
C49783 AND2X1_LOC_856/B OR2X1_LOC_428/A 0.08fF
C50471 OR2X1_LOC_178/Y OR2X1_LOC_428/A 0.04fF
C50585 OR2X1_LOC_258/Y OR2X1_LOC_428/A 0.02fF
C50689 AND2X1_LOC_318/Y OR2X1_LOC_428/A 0.03fF
C51401 OR2X1_LOC_385/Y OR2X1_LOC_428/A 0.03fF
C51684 AND2X1_LOC_810/B OR2X1_LOC_428/A 0.14fF
C52558 AND2X1_LOC_715/A OR2X1_LOC_428/A 0.08fF
C53060 AND2X1_LOC_729/Y OR2X1_LOC_428/A 0.07fF
C53083 AND2X1_LOC_784/A OR2X1_LOC_428/A 0.07fF
C53153 AND2X1_LOC_639/A OR2X1_LOC_428/A 0.19fF
C53263 OR2X1_LOC_428/A OR2X1_LOC_172/Y 0.06fF
C53520 OR2X1_LOC_52/B OR2X1_LOC_428/A 0.37fF
C53533 AND2X1_LOC_489/Y OR2X1_LOC_428/A 0.02fF
C53815 OR2X1_LOC_281/Y OR2X1_LOC_428/A 0.33fF
C53923 AND2X1_LOC_356/B OR2X1_LOC_428/A 0.03fF
C53929 OR2X1_LOC_280/Y OR2X1_LOC_428/A 0.01fF
C55068 OR2X1_LOC_51/Y OR2X1_LOC_428/A 0.78fF
C55603 OR2X1_LOC_423/a_8_216# OR2X1_LOC_428/A 0.01fF
C55952 OR2X1_LOC_178/a_8_216# OR2X1_LOC_428/A 0.14fF
C56418 OR2X1_LOC_428/A VSS 1.83fF
C5247 OR2X1_LOC_87/B OR2X1_LOC_771/B 0.07fF
C6179 OR2X1_LOC_87/B AND2X1_LOC_44/Y 0.18fF
C13443 OR2X1_LOC_87/B AND2X1_LOC_36/Y 5.54fF
C36858 OR2X1_LOC_87/B OR2X1_LOC_375/A 0.06fF
C38949 AND2X1_LOC_19/Y OR2X1_LOC_87/B 0.05fF
C41160 OR2X1_LOC_87/A OR2X1_LOC_87/B 0.39fF
C42299 OR2X1_LOC_97/A OR2X1_LOC_87/B 0.03fF
C49773 VDD OR2X1_LOC_87/B 0.31fF
C50726 OR2X1_LOC_462/B OR2X1_LOC_87/B 0.03fF
C52798 OR2X1_LOC_160/A OR2X1_LOC_87/B 0.03fF
C57036 OR2X1_LOC_87/B VSS 0.30fF
C8490 AND2X1_LOC_82/Y AND2X1_LOC_51/Y 0.02fF
C13137 AND2X1_LOC_82/Y OR2X1_LOC_557/A 0.05fF
C19461 OR2X1_LOC_287/B AND2X1_LOC_82/Y 1.06fF
C29509 AND2X1_LOC_82/Y OR2X1_LOC_78/A 0.65fF
C34094 AND2X1_LOC_765/a_8_24# AND2X1_LOC_82/Y 0.05fF
C40497 AND2X1_LOC_82/Y OR2X1_LOC_78/a_8_216# 0.01fF
C47927 VDD AND2X1_LOC_82/Y 0.16fF
C49157 AND2X1_LOC_82/Y AND2X1_LOC_83/a_8_24# 0.11fF
C50476 AND2X1_LOC_397/a_8_24# AND2X1_LOC_82/Y 0.09fF
C51009 AND2X1_LOC_82/Y AND2X1_LOC_86/B 0.03fF
C51756 AND2X1_LOC_82/Y OR2X1_LOC_78/Y 0.37fF
C55971 OR2X1_LOC_402/B AND2X1_LOC_82/Y 0.84fF
C57719 AND2X1_LOC_82/Y VSS 0.16fF
C1032 AND2X1_LOC_81/B AND2X1_LOC_31/Y 0.03fF
C1335 AND2X1_LOC_81/B OR2X1_LOC_633/B 0.02fF
C1451 AND2X1_LOC_81/B OR2X1_LOC_608/Y 0.01fF
C1995 OR2X1_LOC_506/Y AND2X1_LOC_81/B 0.01fF
C3420 AND2X1_LOC_81/B AND2X1_LOC_504/a_8_24# 0.01fF
C5445 AND2X1_LOC_81/B OR2X1_LOC_493/A 0.05fF
C6936 AND2X1_LOC_81/B AND2X1_LOC_609/a_8_24# 0.01fF
C7696 AND2X1_LOC_81/B OR2X1_LOC_647/B 0.01fF
C8951 AND2X1_LOC_81/B OR2X1_LOC_507/B 0.01fF
C10925 AND2X1_LOC_81/B OR2X1_LOC_151/A 0.03fF
C16203 AND2X1_LOC_81/B OR2X1_LOC_473/Y 0.33fF
C16899 AND2X1_LOC_81/B AND2X1_LOC_505/a_8_24# 0.01fF
C17867 AND2X1_LOC_81/B OR2X1_LOC_810/A 0.06fF
C18167 OR2X1_LOC_715/B AND2X1_LOC_81/B 0.03fF
C18323 AND2X1_LOC_81/B AND2X1_LOC_81/a_8_24# 0.11fF
C19938 AND2X1_LOC_81/B OR2X1_LOC_78/A 0.08fF
C22486 AND2X1_LOC_81/B OR2X1_LOC_507/A 0.01fF
C22644 AND2X1_LOC_81/B OR2X1_LOC_646/A 0.01fF
C25500 AND2X1_LOC_81/B OR2X1_LOC_375/A 0.11fF
C25777 AND2X1_LOC_81/B OR2X1_LOC_549/A 0.03fF
C27540 AND2X1_LOC_81/B AND2X1_LOC_316/a_8_24# 0.09fF
C28308 AND2X1_LOC_81/B OR2X1_LOC_139/A 0.05fF
C29724 AND2X1_LOC_81/B OR2X1_LOC_87/A 0.08fF
C30365 AND2X1_LOC_81/B OR2X1_LOC_130/a_8_216# 0.05fF
C30762 AND2X1_LOC_81/B AND2X1_LOC_239/a_8_24# 0.01fF
C32209 OR2X1_LOC_154/A AND2X1_LOC_81/B 0.01fF
C35992 OR2X1_LOC_100/Y AND2X1_LOC_81/B 0.01fF
C36130 AND2X1_LOC_81/B OR2X1_LOC_532/B 0.10fF
C37250 AND2X1_LOC_81/B AND2X1_LOC_503/a_8_24# 0.01fF
C38029 AND2X1_LOC_81/B VDD 0.57fF
C40644 AND2X1_LOC_81/B OR2X1_LOC_216/A 0.20fF
C41125 OR2X1_LOC_160/A AND2X1_LOC_81/B 0.05fF
C41360 AND2X1_LOC_81/B OR2X1_LOC_130/Y 0.03fF
C42427 AND2X1_LOC_81/B OR2X1_LOC_608/a_8_216# 0.01fF
C42463 AND2X1_LOC_81/B OR2X1_LOC_185/A 0.03fF
C43647 AND2X1_LOC_81/B OR2X1_LOC_641/A 0.03fF
C44641 AND2X1_LOC_81/B OR2X1_LOC_643/A 0.03fF
C47150 AND2X1_LOC_81/B OR2X1_LOC_646/B 0.16fF
C47288 AND2X1_LOC_81/B OR2X1_LOC_506/A 0.03fF
C48557 AND2X1_LOC_81/B OR2X1_LOC_509/A 0.01fF
C50059 AND2X1_LOC_81/B OR2X1_LOC_771/B 0.05fF
C50498 OR2X1_LOC_506/a_8_216# AND2X1_LOC_81/B 0.01fF
C50958 AND2X1_LOC_81/B AND2X1_LOC_44/Y 0.03fF
C51630 AND2X1_LOC_81/B OR2X1_LOC_506/B 0.01fF
C51849 AND2X1_LOC_81/B AND2X1_LOC_18/Y 0.03fF
C51900 AND2X1_LOC_81/B OR2X1_LOC_473/a_8_216# 0.14fF
C54946 AND2X1_LOC_81/B AND2X1_LOC_51/Y 2.53fF
C57892 AND2X1_LOC_81/B VSS -0.49fF
C214 OR2X1_LOC_45/B OR2X1_LOC_427/A 0.15fF
C489 OR2X1_LOC_427/A OR2X1_LOC_428/Y 0.01fF
C664 OR2X1_LOC_158/A OR2X1_LOC_427/A 0.37fF
C745 OR2X1_LOC_103/Y OR2X1_LOC_427/A 0.01fF
C1286 OR2X1_LOC_748/A OR2X1_LOC_427/A 0.01fF
C2249 OR2X1_LOC_146/Y OR2X1_LOC_427/A 0.01fF
C2430 OR2X1_LOC_591/Y OR2X1_LOC_427/A 0.08fF
C2456 OR2X1_LOC_427/A OR2X1_LOC_583/a_36_216# 0.02fF
C2570 AND2X1_LOC_317/a_8_24# OR2X1_LOC_427/A 0.01fF
C2615 OR2X1_LOC_438/a_8_216# OR2X1_LOC_427/A 0.01fF
C2865 OR2X1_LOC_427/A OR2X1_LOC_765/a_8_216# 0.01fF
C2873 AND2X1_LOC_541/Y OR2X1_LOC_427/A 0.01fF
C2909 OR2X1_LOC_107/a_8_216# OR2X1_LOC_427/A 0.03fF
C3042 AND2X1_LOC_390/B OR2X1_LOC_427/A 0.07fF
C3272 OR2X1_LOC_427/A OR2X1_LOC_604/Y 0.01fF
C3329 OR2X1_LOC_744/A OR2X1_LOC_427/A 0.23fF
C3419 OR2X1_LOC_427/A AND2X1_LOC_840/B 0.10fF
C3672 OR2X1_LOC_427/A AND2X1_LOC_464/A 0.03fF
C3770 OR2X1_LOC_144/Y OR2X1_LOC_427/A 0.03fF
C4575 OR2X1_LOC_427/A OR2X1_LOC_426/Y 0.01fF
C4921 OR2X1_LOC_427/A AND2X1_LOC_285/Y 0.02fF
C5023 OR2X1_LOC_91/Y OR2X1_LOC_427/A 0.10fF
C5048 OR2X1_LOC_427/A AND2X1_LOC_446/a_8_24# 0.01fF
C5054 OR2X1_LOC_189/Y OR2X1_LOC_427/A 0.03fF
C5101 OR2X1_LOC_417/Y OR2X1_LOC_427/A 0.04fF
C5105 OR2X1_LOC_311/Y OR2X1_LOC_427/A 0.03fF
C5166 OR2X1_LOC_427/A AND2X1_LOC_483/Y 0.03fF
C5496 OR2X1_LOC_427/A AND2X1_LOC_276/Y 0.01fF
C5822 OR2X1_LOC_441/Y OR2X1_LOC_427/A 0.06fF
C6152 OR2X1_LOC_135/a_8_216# OR2X1_LOC_427/A 0.02fF
C6500 OR2X1_LOC_427/A AND2X1_LOC_789/Y 0.09fF
C6876 OR2X1_LOC_427/A OR2X1_LOC_409/B 0.03fF
C7001 OR2X1_LOC_146/a_8_216# OR2X1_LOC_427/A 0.01fF
C7201 OR2X1_LOC_497/Y OR2X1_LOC_427/A 0.07fF
C7601 OR2X1_LOC_109/a_8_216# OR2X1_LOC_427/A 0.03fF
C8073 AND2X1_LOC_319/A OR2X1_LOC_427/A 0.03fF
C8194 OR2X1_LOC_604/a_8_216# OR2X1_LOC_427/A 0.02fF
C8227 OR2X1_LOC_427/A AND2X1_LOC_721/A 0.03fF
C8554 OR2X1_LOC_427/A AND2X1_LOC_361/A 0.33fF
C8668 OR2X1_LOC_427/A OR2X1_LOC_430/Y 0.01fF
C9332 AND2X1_LOC_147/a_8_24# OR2X1_LOC_427/A 0.03fF
C10093 OR2X1_LOC_600/A OR2X1_LOC_427/A 0.36fF
C10190 OR2X1_LOC_427/A OR2X1_LOC_619/Y 0.03fF
C10660 OR2X1_LOC_427/A AND2X1_LOC_454/A 0.03fF
C10855 OR2X1_LOC_427/A AND2X1_LOC_783/B 0.01fF
C11178 OR2X1_LOC_427/A OR2X1_LOC_406/A -0.04fF
C11843 AND2X1_LOC_113/a_8_24# OR2X1_LOC_427/A 0.02fF
C12380 AND2X1_LOC_307/a_8_24# OR2X1_LOC_427/A 0.08fF
C12506 OR2X1_LOC_427/A OR2X1_LOC_13/B 0.93fF
C13647 OR2X1_LOC_427/A OR2X1_LOC_279/a_8_216# 0.05fF
C13689 AND2X1_LOC_712/B OR2X1_LOC_427/A 0.94fF
C13921 OR2X1_LOC_427/A OR2X1_LOC_765/Y 0.03fF
C14085 OR2X1_LOC_427/A OR2X1_LOC_89/A 15.38fF
C14176 OR2X1_LOC_427/A AND2X1_LOC_451/a_8_24# 0.01fF
C14856 OR2X1_LOC_427/a_8_216# OR2X1_LOC_427/A 0.01fF
C14889 OR2X1_LOC_427/A OR2X1_LOC_591/a_8_216# 0.02fF
C14983 OR2X1_LOC_427/A OR2X1_LOC_95/Y 0.96fF
C15239 OR2X1_LOC_427/A OR2X1_LOC_257/a_36_216# 0.02fF
C15622 OR2X1_LOC_438/Y OR2X1_LOC_427/A 0.04fF
C15642 OR2X1_LOC_427/A OR2X1_LOC_427/Y 0.01fF
C15656 OR2X1_LOC_427/A AND2X1_LOC_621/Y 0.09fF
C16168 OR2X1_LOC_70/Y OR2X1_LOC_427/A 4.74fF
C16196 AND2X1_LOC_538/a_8_24# OR2X1_LOC_427/A 0.06fF
C16242 OR2X1_LOC_184/Y OR2X1_LOC_427/A 0.18fF
C17650 OR2X1_LOC_427/A OR2X1_LOC_16/A 0.12fF
C17680 OR2X1_LOC_108/Y OR2X1_LOC_427/A 0.07fF
C18671 OR2X1_LOC_109/Y OR2X1_LOC_427/A 0.02fF
C18685 OR2X1_LOC_427/A AND2X1_LOC_448/Y 0.03fF
C18773 AND2X1_LOC_729/B OR2X1_LOC_427/A 0.03fF
C19212 OR2X1_LOC_679/A OR2X1_LOC_427/A 0.03fF
C19227 AND2X1_LOC_227/Y OR2X1_LOC_427/A 0.03fF
C19464 OR2X1_LOC_107/Y OR2X1_LOC_427/A 0.01fF
C19564 OR2X1_LOC_599/A OR2X1_LOC_427/A 0.08fF
C19834 OR2X1_LOC_177/a_8_216# OR2X1_LOC_427/A 0.01fF
C19864 OR2X1_LOC_40/Y OR2X1_LOC_427/A 0.11fF
C20018 OR2X1_LOC_427/A OR2X1_LOC_7/A 0.36fF
C20538 OR2X1_LOC_427/A OR2X1_LOC_615/Y 0.24fF
C21117 OR2X1_LOC_589/A OR2X1_LOC_427/A 0.03fF
C21128 OR2X1_LOC_427/A OR2X1_LOC_322/Y 0.01fF
C21223 OR2X1_LOC_495/Y OR2X1_LOC_427/A 0.03fF
C21233 OR2X1_LOC_427/A AND2X1_LOC_450/a_8_24# 0.02fF
C21462 OR2X1_LOC_427/A OR2X1_LOC_384/a_8_216# 0.02fF
C22182 OR2X1_LOC_3/Y OR2X1_LOC_427/A 0.16fF
C22565 AND2X1_LOC_113/Y OR2X1_LOC_427/A 0.01fF
C22962 AND2X1_LOC_113/a_36_24# OR2X1_LOC_427/A 0.01fF
C23473 OR2X1_LOC_64/Y OR2X1_LOC_427/A 0.16fF
C23640 OR2X1_LOC_427/A OR2X1_LOC_89/a_36_216# 0.02fF
C23806 AND2X1_LOC_161/a_8_24# OR2X1_LOC_427/A 0.06fF
C24108 OR2X1_LOC_427/A OR2X1_LOC_524/a_8_216# 0.01fF
C24989 AND2X1_LOC_456/B OR2X1_LOC_427/A 0.06fF
C25778 OR2X1_LOC_494/Y OR2X1_LOC_427/A 0.03fF
C26602 OR2X1_LOC_427/A AND2X1_LOC_778/Y 0.07fF
C26718 OR2X1_LOC_427/A AND2X1_LOC_624/A 0.06fF
C27496 OR2X1_LOC_524/Y OR2X1_LOC_427/A 0.01fF
C27663 OR2X1_LOC_427/A AND2X1_LOC_635/a_8_24# 0.01fF
C28055 OR2X1_LOC_427/A OR2X1_LOC_418/a_8_216# 0.01fF
C28182 OR2X1_LOC_427/A AND2X1_LOC_779/Y 0.04fF
C29079 OR2X1_LOC_427/A OR2X1_LOC_89/Y 0.03fF
C29312 OR2X1_LOC_754/A OR2X1_LOC_427/A 0.08fF
C29481 OR2X1_LOC_427/A OR2X1_LOC_142/Y 2.39fF
C29717 OR2X1_LOC_427/A OR2X1_LOC_238/Y 0.03fF
C30276 OR2X1_LOC_427/A OR2X1_LOC_754/Y 0.02fF
C30682 OR2X1_LOC_427/A OR2X1_LOC_152/A 0.03fF
C30827 OR2X1_LOC_177/Y OR2X1_LOC_427/A 0.14fF
C30854 OR2X1_LOC_604/A OR2X1_LOC_427/A 0.78fF
C31738 OR2X1_LOC_164/Y OR2X1_LOC_427/A 0.11fF
C31894 OR2X1_LOC_427/A AND2X1_LOC_450/Y 0.01fF
C32976 OR2X1_LOC_427/A AND2X1_LOC_434/Y 0.07fF
C33565 OR2X1_LOC_427/A AND2X1_LOC_260/a_8_24# 0.03fF
C35037 OR2X1_LOC_135/Y OR2X1_LOC_427/A 0.01fF
C35153 OR2X1_LOC_427/A AND2X1_LOC_848/Y 0.03fF
C36001 OR2X1_LOC_313/a_8_216# OR2X1_LOC_427/A 0.01fF
C36357 OR2X1_LOC_697/a_8_216# OR2X1_LOC_427/A 0.06fF
C36687 AND2X1_LOC_361/a_8_24# OR2X1_LOC_427/A -0.02fF
C36855 OR2X1_LOC_385/Y OR2X1_LOC_427/A 0.07fF
C38139 OR2X1_LOC_427/A OR2X1_LOC_754/a_8_216# 0.01fF
C38415 AND2X1_LOC_547/Y OR2X1_LOC_427/A 0.02fF
C38525 AND2X1_LOC_729/Y OR2X1_LOC_427/A 0.03fF
C38641 OR2X1_LOC_427/A AND2X1_LOC_639/A 0.04fF
C39028 OR2X1_LOC_427/A OR2X1_LOC_52/B 0.27fF
C39039 AND2X1_LOC_489/Y OR2X1_LOC_427/A 0.03fF
C39283 OR2X1_LOC_427/A OR2X1_LOC_584/Y 0.03fF
C39459 OR2X1_LOC_280/Y OR2X1_LOC_427/A 0.23fF
C39928 OR2X1_LOC_427/A OR2X1_LOC_428/a_8_216# 0.01fF
C40571 OR2X1_LOC_51/Y OR2X1_LOC_427/A 2.02fF
C40664 OR2X1_LOC_680/A OR2X1_LOC_427/A 0.07fF
C41271 OR2X1_LOC_427/A AND2X1_LOC_790/a_8_24# 0.01fF
C41549 OR2X1_LOC_603/a_8_216# OR2X1_LOC_427/A 0.01fF
C41562 OR2X1_LOC_145/a_8_216# OR2X1_LOC_427/A 0.01fF
C41678 OR2X1_LOC_145/Y OR2X1_LOC_427/A 0.02fF
C41969 OR2X1_LOC_313/Y OR2X1_LOC_427/A 0.01fF
C42356 OR2X1_LOC_677/a_8_216# OR2X1_LOC_427/A 0.06fF
C42862 OR2X1_LOC_427/A OR2X1_LOC_511/Y 0.01fF
C42984 OR2X1_LOC_427/A AND2X1_LOC_451/Y 0.08fF
C43754 OR2X1_LOC_669/Y OR2X1_LOC_427/A 0.07fF
C44637 OR2X1_LOC_427/A OR2X1_LOC_74/A 16.42fF
C44656 OR2X1_LOC_427/A OR2X1_LOC_261/A 0.01fF
C45039 OR2X1_LOC_427/A AND2X1_LOC_287/Y 0.36fF
C45752 AND2X1_LOC_704/a_8_24# OR2X1_LOC_427/A 0.01fF
C45845 AND2X1_LOC_779/a_8_24# OR2X1_LOC_427/A 0.02fF
C45959 OR2X1_LOC_615/a_8_216# OR2X1_LOC_427/A 0.01fF
C46158 OR2X1_LOC_134/Y OR2X1_LOC_427/A 0.01fF
C46610 OR2X1_LOC_106/Y OR2X1_LOC_427/A 0.07fF
C47141 OR2X1_LOC_427/A AND2X1_LOC_614/a_8_24# 0.01fF
C47751 OR2X1_LOC_680/Y OR2X1_LOC_427/A 0.03fF
C47771 OR2X1_LOC_696/Y OR2X1_LOC_427/A 0.03fF
C48006 AND2X1_LOC_362/B OR2X1_LOC_427/A 0.04fF
C48430 OR2X1_LOC_427/A OR2X1_LOC_603/Y 0.01fF
C49425 OR2X1_LOC_427/A OR2X1_LOC_89/a_8_216# 0.02fF
C50260 OR2X1_LOC_427/A OR2X1_LOC_418/Y 0.01fF
C51368 AND2X1_LOC_714/B OR2X1_LOC_427/A 0.03fF
C52123 OR2X1_LOC_516/Y OR2X1_LOC_427/A 0.07fF
C52505 OR2X1_LOC_427/A AND2X1_LOC_793/B 0.01fF
C53076 OR2X1_LOC_427/A OR2X1_LOC_583/a_8_216# 0.03fF
C53178 OR2X1_LOC_314/Y OR2X1_LOC_427/A 0.01fF
C53495 AND2X1_LOC_361/a_36_24# OR2X1_LOC_427/A -0.02fF
C53515 VDD OR2X1_LOC_427/A 0.75fF
C53563 OR2X1_LOC_677/Y OR2X1_LOC_427/A 0.03fF
C53659 OR2X1_LOC_251/Y OR2X1_LOC_427/A 0.06fF
C53787 OR2X1_LOC_427/A OR2X1_LOC_163/Y 0.16fF
C53973 OR2X1_LOC_314/a_8_216# OR2X1_LOC_427/A 0.01fF
C54264 OR2X1_LOC_427/A AND2X1_LOC_457/a_8_24# 0.01fF
C54445 OR2X1_LOC_427/A OR2X1_LOC_591/A 0.01fF
C54684 OR2X1_LOC_494/A OR2X1_LOC_427/A 0.03fF
C57043 OR2X1_LOC_427/A VSS 1.39fF
C9648 OR2X1_LOC_87/A OR2X1_LOC_227/A 0.03fF
C14385 OR2X1_LOC_227/a_8_216# OR2X1_LOC_227/A 0.47fF
C21092 OR2X1_LOC_160/A OR2X1_LOC_227/A 0.03fF
C23588 OR2X1_LOC_641/A OR2X1_LOC_227/A 0.02fF
C32455 OR2X1_LOC_130/A OR2X1_LOC_227/A 0.05fF
C36885 AND2X1_LOC_31/Y OR2X1_LOC_227/A 0.01fF
C56367 OR2X1_LOC_227/A VSS 0.13fF
C1128 OR2X1_LOC_532/B OR2X1_LOC_446/B 0.03fF
C2737 OR2X1_LOC_798/Y OR2X1_LOC_446/B 0.22fF
C3137 VDD OR2X1_LOC_446/B 0.13fF
C3968 OR2X1_LOC_676/Y OR2X1_LOC_446/B 0.05fF
C3980 OR2X1_LOC_834/A OR2X1_LOC_446/B 0.03fF
C5194 OR2X1_LOC_840/A OR2X1_LOC_446/B 0.01fF
C5662 OR2X1_LOC_802/Y OR2X1_LOC_446/B 0.90fF
C6071 OR2X1_LOC_160/A OR2X1_LOC_446/B 0.21fF
C6482 OR2X1_LOC_447/A OR2X1_LOC_446/B 0.02fF
C7400 OR2X1_LOC_185/A OR2X1_LOC_446/B 0.03fF
C7873 OR2X1_LOC_702/A OR2X1_LOC_446/B 0.01fF
C8272 OR2X1_LOC_802/a_8_216# OR2X1_LOC_446/B 0.01fF
C9587 OR2X1_LOC_778/Y OR2X1_LOC_446/B 0.14fF
C9877 AND2X1_LOC_91/B OR2X1_LOC_446/B 0.03fF
C9977 OR2X1_LOC_799/A OR2X1_LOC_446/B 0.09fF
C10430 AND2X1_LOC_56/B OR2X1_LOC_446/B 0.07fF
C11772 AND2X1_LOC_47/Y OR2X1_LOC_446/B 0.12fF
C12064 OR2X1_LOC_506/A OR2X1_LOC_446/B 0.03fF
C15675 OR2X1_LOC_446/B OR2X1_LOC_317/B 0.14fF
C15768 AND2X1_LOC_44/Y OR2X1_LOC_446/B 0.03fF
C17570 OR2X1_LOC_447/a_8_216# OR2X1_LOC_446/B 0.01fF
C18041 OR2X1_LOC_449/B OR2X1_LOC_446/B 0.06fF
C19413 OR2X1_LOC_447/Y OR2X1_LOC_446/B 0.09fF
C19817 AND2X1_LOC_51/Y OR2X1_LOC_446/B 0.06fF
C22101 AND2X1_LOC_31/Y OR2X1_LOC_446/B 0.06fF
C23043 AND2X1_LOC_36/Y OR2X1_LOC_446/B 0.76fF
C23953 OR2X1_LOC_446/B OR2X1_LOC_730/A 0.02fF
C25283 OR2X1_LOC_269/B OR2X1_LOC_446/B 0.14fF
C25674 OR2X1_LOC_539/Y OR2X1_LOC_446/B 0.01fF
C25939 OR2X1_LOC_446/B OR2X1_LOC_319/Y 0.06fF
C26050 OR2X1_LOC_678/Y OR2X1_LOC_446/B 0.08fF
C26320 OR2X1_LOC_777/B OR2X1_LOC_446/B 0.02fF
C26840 OR2X1_LOC_161/B OR2X1_LOC_446/B 0.07fF
C29431 OR2X1_LOC_319/B OR2X1_LOC_446/B 0.15fF
C29450 OR2X1_LOC_318/Y OR2X1_LOC_446/B 0.03fF
C30504 OR2X1_LOC_446/B OR2X1_LOC_513/Y 0.03fF
C30850 OR2X1_LOC_436/Y OR2X1_LOC_446/B 0.01fF
C31172 OR2X1_LOC_799/a_8_216# OR2X1_LOC_446/B 0.01fF
C31904 OR2X1_LOC_151/A OR2X1_LOC_446/B 0.07fF
C34353 OR2X1_LOC_446/B OR2X1_LOC_308/Y 0.05fF
C34529 AND2X1_LOC_516/a_8_24# OR2X1_LOC_446/B 0.01fF
C35375 OR2X1_LOC_446/a_8_216# OR2X1_LOC_446/B 0.02fF
C37458 AND2X1_LOC_423/a_8_24# OR2X1_LOC_446/B 0.01fF
C39122 OR2X1_LOC_715/B OR2X1_LOC_446/B 0.20fF
C40013 OR2X1_LOC_687/Y OR2X1_LOC_446/B 0.03fF
C40813 OR2X1_LOC_78/A OR2X1_LOC_446/B 0.03fF
C40897 OR2X1_LOC_446/a_36_216# OR2X1_LOC_446/B 0.03fF
C42151 OR2X1_LOC_538/A OR2X1_LOC_446/B 0.03fF
C42189 OR2X1_LOC_802/A OR2X1_LOC_446/B 0.03fF
C43043 OR2X1_LOC_623/B OR2X1_LOC_446/B 0.03fF
C45145 OR2X1_LOC_186/Y OR2X1_LOC_446/B 0.57fF
C45301 OR2X1_LOC_196/B OR2X1_LOC_446/B 0.10fF
C45691 OR2X1_LOC_574/A OR2X1_LOC_446/B 5.68fF
C46568 OR2X1_LOC_375/A OR2X1_LOC_446/B 0.03fF
C46832 OR2X1_LOC_446/B OR2X1_LOC_515/Y 0.14fF
C50888 OR2X1_LOC_87/A OR2X1_LOC_446/B 0.02fF
C52454 OR2X1_LOC_446/B OR2X1_LOC_713/A 0.07fF
C53384 OR2X1_LOC_154/A OR2X1_LOC_446/B 0.08fF
C56424 OR2X1_LOC_446/B VSS 0.49fF
C10502 AND2X1_LOC_51/Y OR2X1_LOC_333/A 0.05fF
C43583 OR2X1_LOC_333/B OR2X1_LOC_333/A 0.01fF
C56302 OR2X1_LOC_333/A VSS -0.11fF
C28190 AND2X1_LOC_91/B OR2X1_LOC_489/A 0.01fF
C43631 OR2X1_LOC_489/A OR2X1_LOC_269/B 0.02fF
C47572 OR2X1_LOC_489/B OR2X1_LOC_489/A 1.23fF
C56732 OR2X1_LOC_489/A VSS -0.15fF
C564 OR2X1_LOC_286/a_8_216# OR2X1_LOC_286/B 0.08fF
C14651 OR2X1_LOC_288/A OR2X1_LOC_286/B 0.02fF
C17112 OR2X1_LOC_286/B OR2X1_LOC_269/B 0.35fF
C25227 OR2X1_LOC_285/B OR2X1_LOC_286/B 0.10fF
C39993 OR2X1_LOC_285/Y OR2X1_LOC_286/B 0.06fF
C51110 VDD OR2X1_LOC_286/B 0.21fF
C51174 AND2X1_LOC_755/a_8_24# OR2X1_LOC_286/B 0.20fF
C56833 OR2X1_LOC_286/B VSS 0.28fF
C27194 OR2X1_LOC_335/B OR2X1_LOC_543/A 0.38fF
C29927 OR2X1_LOC_335/B OR2X1_LOC_318/B 0.16fF
C34420 OR2X1_LOC_335/B OR2X1_LOC_375/A 0.01fF
C35987 OR2X1_LOC_335/B AND2X1_LOC_603/a_8_24# 0.02fF
C38678 OR2X1_LOC_335/B OR2X1_LOC_87/A 0.11fF
C43756 OR2X1_LOC_335/B OR2X1_LOC_370/a_8_216# 0.47fF
C48079 OR2X1_LOC_335/a_8_216# OR2X1_LOC_335/B 0.07fF
C51583 OR2X1_LOC_185/A OR2X1_LOC_335/B 0.39fF
C54557 AND2X1_LOC_56/B OR2X1_LOC_335/B 0.03fF
C57137 OR2X1_LOC_335/B VSS 0.41fF
C9433 OR2X1_LOC_814/Y AND2X1_LOC_815/a_8_24# 0.23fF
C17689 VDD OR2X1_LOC_814/Y 0.16fF
C24463 AND2X1_LOC_91/B OR2X1_LOC_814/Y 0.01fF
C45493 OR2X1_LOC_287/B OR2X1_LOC_814/Y 0.01fF
C57549 OR2X1_LOC_814/Y VSS 0.07fF
C11545 AND2X1_LOC_44/Y OR2X1_LOC_750/Y 0.68fF
C21027 OR2X1_LOC_269/B OR2X1_LOC_750/Y 0.29fF
C22662 OR2X1_LOC_161/B OR2X1_LOC_750/Y 0.65fF
C22768 AND2X1_LOC_536/a_8_24# OR2X1_LOC_750/Y 0.07fF
C33690 OR2X1_LOC_537/A OR2X1_LOC_750/Y 0.01fF
C46927 OR2X1_LOC_389/A OR2X1_LOC_750/Y 0.02fF
C48223 OR2X1_LOC_691/Y OR2X1_LOC_750/Y 0.02fF
C53036 OR2X1_LOC_532/B OR2X1_LOC_750/Y 0.26fF
C54970 VDD OR2X1_LOC_750/Y 0.74fF
C56268 OR2X1_LOC_750/Y VSS -0.81fF
C10853 OR2X1_LOC_516/A OR2X1_LOC_516/Y 0.01fF
C18291 OR2X1_LOC_516/A AND2X1_LOC_840/B 0.03fF
C24107 OR2X1_LOC_516/A AND2X1_LOC_787/A 0.04fF
C24973 OR2X1_LOC_516/A OR2X1_LOC_600/A 0.17fF
C31049 OR2X1_LOC_516/A OR2X1_LOC_70/Y 0.03fF
C39384 OR2X1_LOC_516/A OR2X1_LOC_516/B 0.66fF
C44386 OR2X1_LOC_516/A OR2X1_LOC_142/Y 0.03fF
C45050 OR2X1_LOC_516/A OR2X1_LOC_516/a_8_216# 0.01fF
C53672 OR2X1_LOC_516/A AND2X1_LOC_784/A 0.02fF
C54051 OR2X1_LOC_516/A OR2X1_LOC_52/B 0.03fF
C55758 OR2X1_LOC_516/A OR2X1_LOC_680/A 0.03fF
C58127 OR2X1_LOC_516/A VSS 0.17fF
C300 OR2X1_LOC_112/B OR2X1_LOC_112/A 0.10fF
C4314 OR2X1_LOC_139/A OR2X1_LOC_112/A 0.03fF
C8326 OR2X1_LOC_154/A OR2X1_LOC_112/A 0.11fF
C14198 VDD OR2X1_LOC_112/A 0.21fF
C17143 OR2X1_LOC_809/B OR2X1_LOC_112/A 0.23fF
C18941 OR2X1_LOC_702/A OR2X1_LOC_112/A 0.03fF
C24424 AND2X1_LOC_173/a_8_24# OR2X1_LOC_112/A 0.20fF
C29886 OR2X1_LOC_175/B OR2X1_LOC_112/A 0.04fF
C36622 OR2X1_LOC_539/Y OR2X1_LOC_112/A 0.01fF
C43005 OR2X1_LOC_151/A OR2X1_LOC_112/A 0.03fF
C53351 OR2X1_LOC_538/A OR2X1_LOC_112/A 0.03fF
C56338 OR2X1_LOC_112/A VSS 0.21fF
C2586 OR2X1_LOC_547/B AND2X1_LOC_56/B 1.61fF
C7909 OR2X1_LOC_547/B AND2X1_LOC_44/Y 0.02fF
C15079 OR2X1_LOC_547/B AND2X1_LOC_36/Y 1.46fF
C21318 OR2X1_LOC_547/B AND2X1_LOC_528/a_8_24# 0.04fF
C32225 OR2X1_LOC_547/B OR2X1_LOC_620/B 0.01fF
C37118 OR2X1_LOC_186/Y OR2X1_LOC_547/B 0.09fF
C57557 OR2X1_LOC_547/B VSS -0.03fF
C2760 OR2X1_LOC_325/A OR2X1_LOC_532/Y 0.23fF
C10534 OR2X1_LOC_325/A OR2X1_LOC_703/A 0.01fF
C12128 OR2X1_LOC_325/A AND2X1_LOC_44/Y 0.94fF
C19471 OR2X1_LOC_325/A OR2X1_LOC_325/a_8_216# 0.02fF
C38443 OR2X1_LOC_325/A OR2X1_LOC_538/A 0.01fF
C41367 OR2X1_LOC_186/Y OR2X1_LOC_325/A 0.07fF
C55579 OR2X1_LOC_325/A VDD 0.21fF
C58066 OR2X1_LOC_325/A VSS 0.16fF
C1854 OR2X1_LOC_691/Y AND2X1_LOC_44/Y 0.03fF
C2481 OR2X1_LOC_691/Y OR2X1_LOC_793/B 0.01fF
C2781 OR2X1_LOC_691/Y AND2X1_LOC_18/Y 0.03fF
C3075 OR2X1_LOC_691/Y OR2X1_LOC_789/A 0.01fF
C3700 OR2X1_LOC_691/Y OR2X1_LOC_130/A 0.02fF
C5823 OR2X1_LOC_691/Y AND2X1_LOC_51/Y 0.03fF
C8157 OR2X1_LOC_691/Y AND2X1_LOC_31/Y 0.03fF
C9064 OR2X1_LOC_691/Y AND2X1_LOC_36/Y 0.01fF
C9211 AND2X1_LOC_586/a_8_24# OR2X1_LOC_691/Y 0.01fF
C9975 OR2X1_LOC_691/Y OR2X1_LOC_856/A 0.01fF
C11344 OR2X1_LOC_691/Y OR2X1_LOC_269/B 0.03fF
C12949 OR2X1_LOC_691/Y OR2X1_LOC_161/B 0.03fF
C23760 OR2X1_LOC_691/Y OR2X1_LOC_193/A 0.02fF
C24035 OR2X1_LOC_691/Y OR2X1_LOC_598/Y 0.11fF
C24403 OR2X1_LOC_138/a_8_216# OR2X1_LOC_691/Y 0.01fF
C25265 OR2X1_LOC_715/B OR2X1_LOC_691/Y 0.03fF
C26192 OR2X1_LOC_687/Y OR2X1_LOC_691/Y 0.15fF
C26599 OR2X1_LOC_691/Y OR2X1_LOC_835/B 0.83fF
C29087 OR2X1_LOC_691/Y OR2X1_LOC_623/B 0.03fF
C35317 OR2X1_LOC_139/A OR2X1_LOC_691/Y 0.01fF
C39286 OR2X1_LOC_154/A OR2X1_LOC_691/Y 0.03fF
C39509 OR2X1_LOC_691/Y OR2X1_LOC_198/A 0.45fF
C41849 OR2X1_LOC_379/a_8_216# OR2X1_LOC_691/Y 0.01fF
C43277 OR2X1_LOC_691/Y OR2X1_LOC_532/B 0.01fF
C43924 OR2X1_LOC_691/Y OR2X1_LOC_855/a_8_216# 0.03fF
C43936 OR2X1_LOC_691/Y OR2X1_LOC_729/a_8_216# 0.12fF
C45241 VDD OR2X1_LOC_691/Y 0.31fF
C47616 OR2X1_LOC_691/Y OR2X1_LOC_789/a_8_216# 0.01fF
C48372 OR2X1_LOC_691/Y OR2X1_LOC_809/B 0.01fF
C48436 OR2X1_LOC_160/A OR2X1_LOC_691/Y 0.04fF
C49682 OR2X1_LOC_691/Y OR2X1_LOC_185/A 0.23fF
C50158 OR2X1_LOC_702/A OR2X1_LOC_691/Y 0.02fF
C50939 OR2X1_LOC_379/Y OR2X1_LOC_691/Y 0.43fF
C51757 OR2X1_LOC_691/Y OR2X1_LOC_637/A 0.01fF
C52641 OR2X1_LOC_691/Y AND2X1_LOC_56/B 0.07fF
C53716 OR2X1_LOC_691/Y AND2X1_LOC_751/a_8_24# 0.01fF
C54010 OR2X1_LOC_691/Y AND2X1_LOC_47/Y 0.03fF
C55034 OR2X1_LOC_691/Y OR2X1_LOC_855/a_36_216# 0.02fF
C57732 OR2X1_LOC_691/Y VSS -0.34fF
C974 OR2X1_LOC_837/B AND2X1_LOC_462/B 0.65fF
C11230 AND2X1_LOC_462/B OR2X1_LOC_27/Y 0.21fF
C20939 VDD AND2X1_LOC_462/B 0.02fF
C22811 AND2X1_LOC_462/B OR2X1_LOC_416/Y 0.17fF
C33722 AND2X1_LOC_462/B AND2X1_LOC_462/a_8_24# 0.01fF
C56988 AND2X1_LOC_462/B VSS 0.28fF
C3712 OR2X1_LOC_232/Y OR2X1_LOC_234/Y 0.09fF
C33336 VDD OR2X1_LOC_234/Y 0.10fF
C36663 OR2X1_LOC_158/A OR2X1_LOC_234/Y 0.09fF
C46286 OR2X1_LOC_619/Y OR2X1_LOC_234/Y 0.01fF
C46802 OR2X1_LOC_232/a_8_216# OR2X1_LOC_234/Y 0.40fF
C53858 OR2X1_LOC_234/Y OR2X1_LOC_16/A 0.02fF
C56772 OR2X1_LOC_234/Y VSS 0.11fF
C14898 OR2X1_LOC_823/Y OR2X1_LOC_824/Y 0.04fF
C16893 OR2X1_LOC_158/A OR2X1_LOC_824/Y 0.07fF
C26323 OR2X1_LOC_824/Y OR2X1_LOC_619/Y 0.72fF
C36488 OR2X1_LOC_824/Y AND2X1_LOC_836/a_8_24# 0.06fF
C42053 OR2X1_LOC_824/Y AND2X1_LOC_839/B 0.02fF
C56933 OR2X1_LOC_824/Y VSS -0.16fF
C481 OR2X1_LOC_291/Y OR2X1_LOC_69/Y 0.03fF
C3539 OR2X1_LOC_291/Y OR2X1_LOC_609/a_8_216# 0.02fF
C3828 VDD OR2X1_LOC_291/Y 0.38fF
C5611 OR2X1_LOC_291/Y OR2X1_LOC_416/Y 0.02fF
C6684 OR2X1_LOC_45/B OR2X1_LOC_291/Y 0.03fF
C7165 OR2X1_LOC_158/A OR2X1_LOC_291/Y 0.07fF
C9061 OR2X1_LOC_291/Y OR2X1_LOC_609/a_36_216# 0.02fF
C9469 OR2X1_LOC_291/Y OR2X1_LOC_316/Y 0.02fF
C9815 OR2X1_LOC_291/Y OR2X1_LOC_744/A 0.03fF
C11518 OR2X1_LOC_290/Y OR2X1_LOC_291/Y 0.05fF
C16619 OR2X1_LOC_291/Y OR2X1_LOC_619/Y 0.07fF
C17138 OR2X1_LOC_291/Y AND2X1_LOC_334/a_8_24# 0.11fF
C22387 OR2X1_LOC_291/Y OR2X1_LOC_71/A 0.02fF
C24210 OR2X1_LOC_291/Y OR2X1_LOC_16/A 0.32fF
C26293 OR2X1_LOC_40/Y OR2X1_LOC_291/Y 0.05fF
C27538 OR2X1_LOC_589/A OR2X1_LOC_291/Y 0.03fF
C28568 OR2X1_LOC_3/Y OR2X1_LOC_291/Y 0.03fF
C29381 OR2X1_LOC_291/Y AND2X1_LOC_610/a_8_24# 0.02fF
C34899 OR2X1_LOC_291/Y OR2X1_LOC_612/B 0.03fF
C35424 OR2X1_LOC_291/Y AND2X1_LOC_608/a_8_24# 0.26fF
C43903 OR2X1_LOC_291/Y AND2X1_LOC_634/Y 0.02fF
C45581 OR2X1_LOC_291/Y OR2X1_LOC_52/B 0.03fF
C48675 OR2X1_LOC_291/Y OR2X1_LOC_609/A 0.04fF
C50765 OR2X1_LOC_291/Y OR2X1_LOC_32/B 0.07fF
C51208 OR2X1_LOC_291/Y OR2X1_LOC_74/A 0.49fF
C57607 OR2X1_LOC_291/Y VSS 0.23fF
C905 OR2X1_LOC_269/B OR2X1_LOC_383/a_8_216# 0.01fF
C1027 OR2X1_LOC_269/B OR2X1_LOC_318/B 0.03fF
C1207 OR2X1_LOC_114/B OR2X1_LOC_269/B 0.03fF
C1251 OR2X1_LOC_538/A OR2X1_LOC_269/B 0.03fF
C2118 OR2X1_LOC_623/B OR2X1_LOC_269/B 0.01fF
C2597 OR2X1_LOC_833/B OR2X1_LOC_269/B 0.02fF
C2624 OR2X1_LOC_254/B OR2X1_LOC_269/B 0.03fF
C2629 OR2X1_LOC_848/B OR2X1_LOC_269/B 0.01fF
C4114 OR2X1_LOC_186/Y OR2X1_LOC_269/B 0.03fF
C4239 OR2X1_LOC_773/B OR2X1_LOC_269/B 0.02fF
C5268 OR2X1_LOC_269/B OR2X1_LOC_539/B 0.27fF
C5491 OR2X1_LOC_375/A OR2X1_LOC_269/B 1.86fF
C5795 OR2X1_LOC_269/B OR2X1_LOC_549/A 0.07fF
C6351 OR2X1_LOC_391/B OR2X1_LOC_269/B 0.06fF
C6419 OR2X1_LOC_846/A OR2X1_LOC_269/B 0.03fF
C7249 AND2X1_LOC_823/a_8_24# OR2X1_LOC_269/B 0.05fF
C7324 OR2X1_LOC_285/Y OR2X1_LOC_269/B 0.01fF
C7713 OR2X1_LOC_195/A OR2X1_LOC_269/B 0.03fF
C8082 AND2X1_LOC_384/a_8_24# OR2X1_LOC_269/B 0.01fF
C8397 AND2X1_LOC_701/a_36_24# OR2X1_LOC_269/B 0.01fF
C8429 OR2X1_LOC_269/B OR2X1_LOC_758/a_8_216# 0.01fF
C9371 OR2X1_LOC_834/a_8_216# OR2X1_LOC_269/B 0.01fF
C9471 AND2X1_LOC_697/a_8_24# OR2X1_LOC_269/B 0.11fF
C9481 AND2X1_LOC_666/a_8_24# OR2X1_LOC_269/B 0.01fF
C9850 OR2X1_LOC_87/A OR2X1_LOC_269/B 0.08fF
C10152 OR2X1_LOC_389/A OR2X1_LOC_269/B 0.01fF
C10654 OR2X1_LOC_194/B OR2X1_LOC_269/B 0.05fF
C10917 OR2X1_LOC_97/A OR2X1_LOC_269/B 0.03fF
C11358 OR2X1_LOC_269/B OR2X1_LOC_713/A 0.09fF
C11837 AND2X1_LOC_700/a_8_24# OR2X1_LOC_269/B 0.01fF
C11925 OR2X1_LOC_639/B OR2X1_LOC_269/B 0.05fF
C11955 OR2X1_LOC_333/B OR2X1_LOC_269/B 0.12fF
C12366 OR2X1_LOC_154/A OR2X1_LOC_269/B 0.29fF
C12513 OR2X1_LOC_269/B OR2X1_LOC_198/A 0.01fF
C12898 AND2X1_LOC_821/a_8_24# OR2X1_LOC_269/B 0.03fF
C13196 OR2X1_LOC_538/a_8_216# OR2X1_LOC_269/B 0.01fF
C13850 OR2X1_LOC_269/B OR2X1_LOC_590/Y 0.02fF
C14974 OR2X1_LOC_719/A OR2X1_LOC_269/B 0.01fF
C15068 OR2X1_LOC_269/B OR2X1_LOC_557/a_8_216# 0.01fF
C15153 OR2X1_LOC_269/B OR2X1_LOC_779/A 0.01fF
C15183 OR2X1_LOC_614/Y OR2X1_LOC_269/B 0.01fF
C16135 OR2X1_LOC_286/Y OR2X1_LOC_269/B 0.01fF
C16254 OR2X1_LOC_532/B OR2X1_LOC_269/B 0.26fF
C16513 OR2X1_LOC_391/A OR2X1_LOC_269/B 0.44fF
C17341 OR2X1_LOC_710/B OR2X1_LOC_269/B 0.24fF
C18203 VDD OR2X1_LOC_269/B 2.36fF
C19063 OR2X1_LOC_676/Y OR2X1_LOC_269/B 0.07fF
C19084 OR2X1_LOC_834/A OR2X1_LOC_269/B 0.02fF
C19368 OR2X1_LOC_269/B AND2X1_LOC_591/a_8_24# -0.01fF
C20402 OR2X1_LOC_840/A OR2X1_LOC_269/B 0.01fF
C20475 OR2X1_LOC_789/a_8_216# OR2X1_LOC_269/B 0.05fF
C20743 AND2X1_LOC_754/a_8_24# OR2X1_LOC_269/B 0.01fF
C20955 OR2X1_LOC_846/B OR2X1_LOC_269/B 0.02fF
C21316 OR2X1_LOC_160/A OR2X1_LOC_269/B 0.14fF
C21532 OR2X1_LOC_269/B OR2X1_LOC_532/Y 0.02fF
C21584 OR2X1_LOC_196/Y OR2X1_LOC_269/B 0.01fF
C22605 OR2X1_LOC_185/A OR2X1_LOC_269/B 0.08fF
C22730 AND2X1_LOC_431/a_8_24# OR2X1_LOC_269/B 0.04fF
C23081 OR2X1_LOC_702/A OR2X1_LOC_269/B 0.03fF
C23382 OR2X1_LOC_269/B AND2X1_LOC_437/a_8_24# 0.04fF
C23731 OR2X1_LOC_294/Y OR2X1_LOC_269/B 0.03fF
C23952 OR2X1_LOC_286/a_8_216# OR2X1_LOC_269/B 0.10fF
C24255 OR2X1_LOC_538/a_36_216# OR2X1_LOC_269/B 0.02fF
C24276 OR2X1_LOC_541/B OR2X1_LOC_269/B 0.09fF
C24727 OR2X1_LOC_778/Y OR2X1_LOC_269/B 0.05fF
C24933 AND2X1_LOC_91/B OR2X1_LOC_269/B 0.70fF
C25068 OR2X1_LOC_308/a_8_216# OR2X1_LOC_269/B 0.01fF
C25289 OR2X1_LOC_269/B OR2X1_LOC_303/B 0.03fF
C25393 OR2X1_LOC_269/B OR2X1_LOC_719/B 0.02fF
C25417 OR2X1_LOC_542/B OR2X1_LOC_269/B 0.01fF
C25532 AND2X1_LOC_56/B OR2X1_LOC_269/B 0.28fF
C26104 OR2X1_LOC_269/B OR2X1_LOC_561/B 0.01fF
C26231 OR2X1_LOC_790/A OR2X1_LOC_269/B 0.01fF
C26873 AND2X1_LOC_47/Y OR2X1_LOC_269/B 1.91fF
C27408 OR2X1_LOC_269/B OR2X1_LOC_180/B 0.03fF
C27568 OR2X1_LOC_391/a_8_216# OR2X1_LOC_269/B 0.01fF
C27813 OR2X1_LOC_269/B AND2X1_LOC_41/Y 0.03fF
C29212 OR2X1_LOC_758/Y OR2X1_LOC_269/B 0.10fF
C29250 OR2X1_LOC_703/A OR2X1_LOC_269/B 0.03fF
C29301 OR2X1_LOC_791/B OR2X1_LOC_269/B 0.02fF
C29691 OR2X1_LOC_539/A OR2X1_LOC_269/B 0.01fF
C29931 OR2X1_LOC_269/B OR2X1_LOC_771/B 0.07fF
C30368 OR2X1_LOC_269/B OR2X1_LOC_593/B 2.90fF
C30746 OR2X1_LOC_269/B OR2X1_LOC_317/B 0.35fF
C30863 OR2X1_LOC_269/B AND2X1_LOC_44/Y 1.41fF
C31024 OR2X1_LOC_848/a_8_216# OR2X1_LOC_269/B -0.00fF
C31742 AND2X1_LOC_18/Y OR2X1_LOC_269/B 5.02fF
C32115 OR2X1_LOC_307/A OR2X1_LOC_269/B 0.01fF
C32686 OR2X1_LOC_130/A OR2X1_LOC_269/B 0.02fF
C33051 OR2X1_LOC_489/a_8_216# OR2X1_LOC_269/B 0.01fF
C33128 OR2X1_LOC_449/B OR2X1_LOC_269/B 0.03fF
C33291 OR2X1_LOC_269/B OR2X1_LOC_195/a_8_216# 0.09fF
C33641 OR2X1_LOC_383/Y OR2X1_LOC_269/B 0.01fF
C34440 OR2X1_LOC_447/Y OR2X1_LOC_269/B 0.10fF
C34882 AND2X1_LOC_51/Y OR2X1_LOC_269/B 0.20fF
C35698 AND2X1_LOC_135/a_8_24# OR2X1_LOC_269/B 0.05fF
C36008 AND2X1_LOC_253/a_8_24# OR2X1_LOC_269/B 0.04fF
C36384 OR2X1_LOC_284/a_8_216# OR2X1_LOC_269/B 0.07fF
C36894 AND2X1_LOC_701/a_8_24# OR2X1_LOC_269/B 0.03fF
C37040 AND2X1_LOC_31/Y OR2X1_LOC_269/B 0.73fF
C37370 AND2X1_LOC_281/a_8_24# OR2X1_LOC_269/B 0.14fF
C37819 OR2X1_LOC_288/A OR2X1_LOC_269/B 0.03fF
C37932 OR2X1_LOC_269/B AND2X1_LOC_36/Y 1.00fF
C38296 OR2X1_LOC_269/B OR2X1_LOC_196/a_8_216# 0.01fF
C38534 OR2X1_LOC_392/A OR2X1_LOC_269/B 0.03fF
C38900 OR2X1_LOC_856/A OR2X1_LOC_269/B 0.02fF
C39121 AND2X1_LOC_494/a_8_24# OR2X1_LOC_269/B 0.01fF
C39224 OR2X1_LOC_269/B OR2X1_LOC_537/a_8_216# 0.05fF
C39512 OR2X1_LOC_557/A OR2X1_LOC_269/B 0.16fF
C39821 OR2X1_LOC_269/B AND2X1_LOC_437/a_36_24# 0.01fF
C41143 AND2X1_LOC_533/a_8_24# OR2X1_LOC_269/B 0.03fF
C41274 OR2X1_LOC_269/B AND2X1_LOC_237/a_8_24# 0.01fF
C41340 OR2X1_LOC_269/B OR2X1_LOC_777/B 0.02fF
C41362 OR2X1_LOC_269/B AND2X1_LOC_591/a_36_24# 0.01fF
C41450 OR2X1_LOC_269/B OR2X1_LOC_344/A 0.03fF
C41834 OR2X1_LOC_198/a_8_216# OR2X1_LOC_269/B 0.01fF
C41885 OR2X1_LOC_269/B OR2X1_LOC_161/B 2.69fF
C42007 AND2X1_LOC_536/a_8_24# OR2X1_LOC_269/B 0.01fF
C42020 OR2X1_LOC_846/a_8_216# OR2X1_LOC_269/B 0.01fF
C44165 OR2X1_LOC_772/B OR2X1_LOC_269/B 0.01fF
C44190 OR2X1_LOC_489/B OR2X1_LOC_269/B 0.03fF
C46407 OR2X1_LOC_553/A OR2X1_LOC_269/B 0.27fF
C47177 OR2X1_LOC_151/A OR2X1_LOC_269/B 0.15fF
C47276 AND2X1_LOC_253/a_36_24# OR2X1_LOC_269/B 0.01fF
C47669 OR2X1_LOC_287/A OR2X1_LOC_269/B 0.42fF
C47724 AND2X1_LOC_482/a_8_24# OR2X1_LOC_269/B 0.01fF
C48222 AND2X1_LOC_252/a_8_24# OR2X1_LOC_269/B 0.01fF
C49662 OR2X1_LOC_269/B OR2X1_LOC_308/Y 0.08fF
C50307 OR2X1_LOC_835/A OR2X1_LOC_269/B 0.05fF
C50678 OR2X1_LOC_448/A OR2X1_LOC_269/B 0.01fF
C50990 OR2X1_LOC_269/B OR2X1_LOC_390/A 0.03fF
C51248 AND2X1_LOC_280/a_8_24# OR2X1_LOC_269/B 0.01fF
C51565 AND2X1_LOC_822/a_8_24# OR2X1_LOC_269/B 0.04fF
C52284 OR2X1_LOC_190/A OR2X1_LOC_269/B 0.03fF
C52385 AND2X1_LOC_533/a_36_24# OR2X1_LOC_269/B 0.01fF
C52508 OR2X1_LOC_269/B OR2X1_LOC_241/B 0.13fF
C52639 OR2X1_LOC_188/Y OR2X1_LOC_269/B 0.03fF
C52760 OR2X1_LOC_285/a_8_216# OR2X1_LOC_269/B 0.01fF
C52765 AND2X1_LOC_615/a_8_24# OR2X1_LOC_269/B 0.01fF
C52875 OR2X1_LOC_193/A OR2X1_LOC_269/B 0.09fF
C53011 OR2X1_LOC_269/B OR2X1_LOC_339/A 0.01fF
C53055 OR2X1_LOC_208/A OR2X1_LOC_269/B 0.01fF
C53117 OR2X1_LOC_831/A OR2X1_LOC_269/B 0.03fF
C53242 OR2X1_LOC_859/B OR2X1_LOC_269/B 0.01fF
C53537 OR2X1_LOC_269/B OR2X1_LOC_356/A 0.88fF
C53839 OR2X1_LOC_269/B OR2X1_LOC_558/A 0.01fF
C54079 OR2X1_LOC_810/A OR2X1_LOC_269/B 0.05fF
C54111 AND2X1_LOC_281/a_36_24# OR2X1_LOC_269/B 0.01fF
C55358 OR2X1_LOC_687/Y OR2X1_LOC_269/B 0.03fF
C55535 OR2X1_LOC_269/B OR2X1_LOC_199/B 0.06fF
C55796 OR2X1_LOC_835/B OR2X1_LOC_269/B 0.15fF
C56130 OR2X1_LOC_78/A OR2X1_LOC_269/B 11.08fF
C56543 OR2X1_LOC_269/B VSS -5.04fF
C1666 OR2X1_LOC_32/B OR2X1_LOC_393/a_8_216# 0.05fF
C7046 OR2X1_LOC_32/B OR2X1_LOC_16/A 5.66fF
C9264 OR2X1_LOC_40/Y OR2X1_LOC_32/B 0.20fF
C9837 OR2X1_LOC_32/B OR2X1_LOC_32/a_8_216# 0.03fF
C10508 OR2X1_LOC_589/A OR2X1_LOC_32/B 0.21fF
C10706 OR2X1_LOC_32/B OR2X1_LOC_60/a_8_216# 0.03fF
C11535 OR2X1_LOC_3/Y OR2X1_LOC_32/B 0.03fF
C20425 OR2X1_LOC_32/B OR2X1_LOC_80/Y 0.03fF
C21391 OR2X1_LOC_32/B AND2X1_LOC_633/Y 0.02fF
C21951 OR2X1_LOC_316/a_8_216# OR2X1_LOC_32/B 0.03fF
C22986 OR2X1_LOC_837/B OR2X1_LOC_32/B 0.43fF
C23829 OR2X1_LOC_32/B OR2X1_LOC_393/Y 0.13fF
C28479 OR2X1_LOC_32/B OR2X1_LOC_52/B 0.11fF
C36590 OR2X1_LOC_32/B OR2X1_LOC_72/Y 0.09fF
C39454 OR2X1_LOC_32/B OR2X1_LOC_69/Y 0.13fF
C42776 VDD OR2X1_LOC_32/B 0.11fF
C43022 OR2X1_LOC_32/B OR2X1_LOC_67/Y 0.02fF
C45745 OR2X1_LOC_45/B OR2X1_LOC_32/B 0.01fF
C46221 OR2X1_LOC_158/A OR2X1_LOC_32/B 0.58fF
C48903 OR2X1_LOC_744/A OR2X1_LOC_32/B 0.20fF
C55621 OR2X1_LOC_32/B OR2X1_LOC_600/A 0.07fF
C57472 OR2X1_LOC_32/B VSS 0.52fF
C261 OR2X1_LOC_87/A AND2X1_LOC_44/Y 0.48fF
C917 OR2X1_LOC_87/A AND2X1_LOC_69/Y 0.03fF
C988 OR2X1_LOC_506/B OR2X1_LOC_87/A 0.03fF
C1193 OR2X1_LOC_87/A AND2X1_LOC_18/Y 0.16fF
C1809 AND2X1_LOC_69/a_8_24# OR2X1_LOC_87/A 0.01fF
C1845 OR2X1_LOC_87/A AND2X1_LOC_428/a_8_24# 0.02fF
C2081 AND2X1_LOC_65/a_8_24# OR2X1_LOC_87/A 0.05fF
C2122 OR2X1_LOC_231/A OR2X1_LOC_87/A 0.14fF
C2157 OR2X1_LOC_87/A OR2X1_LOC_707/A 0.05fF
C2164 OR2X1_LOC_87/A OR2X1_LOC_130/A 1.12fF
C2184 OR2X1_LOC_87/A AND2X1_LOC_7/a_8_24# 0.17fF
C2638 OR2X1_LOC_87/A OR2X1_LOC_449/B 0.07fF
C2662 OR2X1_LOC_636/A OR2X1_LOC_87/A 0.02fF
C3953 OR2X1_LOC_447/Y OR2X1_LOC_87/A 0.07fF
C4259 OR2X1_LOC_116/a_36_216# OR2X1_LOC_87/A 0.02fF
C4275 AND2X1_LOC_525/a_8_24# OR2X1_LOC_87/A 0.05fF
C4302 OR2X1_LOC_87/A AND2X1_LOC_51/Y 0.55fF
C4810 OR2X1_LOC_87/A AND2X1_LOC_52/Y 0.22fF
C4927 OR2X1_LOC_87/A OR2X1_LOC_439/B 0.03fF
C5721 OR2X1_LOC_149/B OR2X1_LOC_87/A 0.07fF
C6439 OR2X1_LOC_614/a_8_216# OR2X1_LOC_87/A 0.01fF
C6484 OR2X1_LOC_87/A AND2X1_LOC_31/Y 0.21fF
C6827 OR2X1_LOC_87/A OR2X1_LOC_633/B 0.82fF
C7380 OR2X1_LOC_87/A OR2X1_LOC_451/B 0.02fF
C7452 OR2X1_LOC_87/A AND2X1_LOC_36/Y 0.13fF
C7508 OR2X1_LOC_154/a_8_216# OR2X1_LOC_87/A 0.02fF
C7520 OR2X1_LOC_506/Y OR2X1_LOC_87/A 0.04fF
C7615 OR2X1_LOC_635/A OR2X1_LOC_87/A 0.01fF
C8167 OR2X1_LOC_636/B OR2X1_LOC_87/A 0.02fF
C8831 OR2X1_LOC_87/A OR2X1_LOC_160/Y 0.03fF
C9430 AND2X1_LOC_584/a_8_24# OR2X1_LOC_87/A 0.01fF
C9781 AND2X1_LOC_312/a_36_24# OR2X1_LOC_87/A 0.01fF
C10844 OR2X1_LOC_87/A OR2X1_LOC_777/B 0.07fF
C10898 OR2X1_LOC_156/Y OR2X1_LOC_87/A 0.09fF
C11335 OR2X1_LOC_87/A OR2X1_LOC_161/B 0.16fF
C11691 OR2X1_LOC_87/A OR2X1_LOC_707/a_8_216# 0.02fF
C12485 OR2X1_LOC_87/A OR2X1_LOC_705/B 0.15fF
C12775 OR2X1_LOC_87/A AND2X1_LOC_230/a_8_24# 0.02fF
C13182 OR2X1_LOC_201/A OR2X1_LOC_87/A 0.09fF
C13280 OR2X1_LOC_87/A OR2X1_LOC_647/B 0.39fF
C14169 OR2X1_LOC_87/A AND2X1_LOC_441/a_8_24# 0.01fF
C15011 OR2X1_LOC_446/Y OR2X1_LOC_87/A 0.29fF
C15270 OR2X1_LOC_635/a_8_216# OR2X1_LOC_87/A 0.01fF
C15360 OR2X1_LOC_76/A OR2X1_LOC_87/A 0.03fF
C15380 OR2X1_LOC_148/A OR2X1_LOC_87/A 0.03fF
C16401 OR2X1_LOC_318/A OR2X1_LOC_87/A 0.05fF
C16429 OR2X1_LOC_151/A OR2X1_LOC_87/A 11.18fF
C18561 OR2X1_LOC_156/B OR2X1_LOC_87/A 0.02fF
C18848 OR2X1_LOC_87/A OR2X1_LOC_783/A 0.02fF
C18932 OR2X1_LOC_87/A OR2X1_LOC_308/Y 0.65fF
C20059 OR2X1_LOC_446/a_8_216# OR2X1_LOC_87/A 0.02fF
C20110 OR2X1_LOC_87/A AND2X1_LOC_7/Y 0.19fF
C20829 AND2X1_LOC_142/a_8_24# OR2X1_LOC_87/A 0.04fF
C21141 AND2X1_LOC_229/a_8_24# OR2X1_LOC_87/A 0.04fF
C21808 OR2X1_LOC_473/Y OR2X1_LOC_87/A 0.08fF
C22453 OR2X1_LOC_87/A AND2X1_LOC_438/a_8_24# 0.06fF
C23467 OR2X1_LOC_810/A OR2X1_LOC_87/A 0.07fF
C23744 OR2X1_LOC_715/B OR2X1_LOC_87/A 0.10fF
C23856 OR2X1_LOC_87/A AND2X1_LOC_230/a_36_24# 0.01fF
C24240 AND2X1_LOC_65/a_36_24# OR2X1_LOC_87/A 0.01fF
C24694 OR2X1_LOC_687/Y OR2X1_LOC_87/A 0.07fF
C25422 OR2X1_LOC_87/A OR2X1_LOC_78/A 0.25fF
C25556 OR2X1_LOC_605/A OR2X1_LOC_87/A 0.12fF
C26297 OR2X1_LOC_147/B OR2X1_LOC_87/A 0.03fF
C26428 OR2X1_LOC_545/B OR2X1_LOC_87/A 0.01fF
C26484 OR2X1_LOC_87/A OR2X1_LOC_318/B 0.03fF
C26606 OR2X1_LOC_231/B OR2X1_LOC_87/A 0.06fF
C26619 OR2X1_LOC_121/Y OR2X1_LOC_87/A 0.07fF
C27711 OR2X1_LOC_87/A OR2X1_LOC_544/A 0.03fF
C28088 OR2X1_LOC_646/A OR2X1_LOC_87/A 0.03fF
C28865 OR2X1_LOC_448/Y OR2X1_LOC_87/A 0.14fF
C29577 OR2X1_LOC_186/Y OR2X1_LOC_87/A 0.07fF
C29727 AND2X1_LOC_747/a_8_24# OR2X1_LOC_87/A 0.01fF
C30186 OR2X1_LOC_574/A OR2X1_LOC_87/A 0.03fF
C30513 AND2X1_LOC_58/a_8_24# OR2X1_LOC_87/A 0.11fF
C31005 OR2X1_LOC_87/A OR2X1_LOC_375/A 7.45fF
C31059 OR2X1_LOC_605/B OR2X1_LOC_87/A 0.15fF
C31290 OR2X1_LOC_87/A OR2X1_LOC_549/A 0.08fF
C31787 AND2X1_LOC_142/a_36_24# OR2X1_LOC_87/A 0.01fF
C32074 AND2X1_LOC_229/a_36_24# OR2X1_LOC_87/A 0.01fF
C32512 OR2X1_LOC_87/A AND2X1_LOC_603/a_8_24# 0.05fF
C32791 OR2X1_LOC_87/A OR2X1_LOC_779/Y 0.02fF
C33014 AND2X1_LOC_19/Y OR2X1_LOC_87/A 0.23fF
C33042 AND2X1_LOC_316/a_8_24# OR2X1_LOC_87/A 0.04fF
C33465 AND2X1_LOC_583/a_8_24# OR2X1_LOC_87/A 0.15fF
C33736 OR2X1_LOC_87/A OR2X1_LOC_712/B 0.02fF
C33796 OR2X1_LOC_139/A OR2X1_LOC_87/A 0.07fF
C35198 OR2X1_LOC_782/B OR2X1_LOC_87/A 0.01fF
C35575 AND2X1_LOC_177/a_8_24# OR2X1_LOC_87/A 0.01fF
C36306 OR2X1_LOC_97/A OR2X1_LOC_87/A 0.05fF
C36396 AND2X1_LOC_744/a_8_24# OR2X1_LOC_87/A 0.01fF
C36413 OR2X1_LOC_87/A OR2X1_LOC_475/B 0.10fF
C37047 OR2X1_LOC_87/A OR2X1_LOC_546/A 0.03fF
C37293 OR2X1_LOC_639/B OR2X1_LOC_87/A 0.03fF
C37456 OR2X1_LOC_87/A OR2X1_LOC_590/a_8_216# 0.01fF
C37470 OR2X1_LOC_87/A OR2X1_LOC_160/a_8_216# 0.05fF
C37732 OR2X1_LOC_154/A OR2X1_LOC_87/A 1.47fF
C37875 OR2X1_LOC_87/A OR2X1_LOC_198/A 0.08fF
C38856 OR2X1_LOC_87/A OR2X1_LOC_267/Y 0.03fF
C39041 OR2X1_LOC_520/Y OR2X1_LOC_87/A 0.03fF
C39220 OR2X1_LOC_87/A OR2X1_LOC_590/Y 0.07fF
C39935 OR2X1_LOC_87/A OR2X1_LOC_227/a_8_216# 0.06fF
C40572 OR2X1_LOC_614/Y OR2X1_LOC_87/A 0.02fF
C41483 OR2X1_LOC_450/A OR2X1_LOC_87/A 0.03fF
C41685 OR2X1_LOC_87/A OR2X1_LOC_532/B 0.42fF
C42728 OR2X1_LOC_87/A AND2X1_LOC_224/a_8_24# 0.01fF
C43278 AND2X1_LOC_52/a_8_24# OR2X1_LOC_87/A 0.01fF
C43677 VDD OR2X1_LOC_87/A 1.71fF
C43848 OR2X1_LOC_444/B OR2X1_LOC_87/A 0.03fF
C44331 OR2X1_LOC_87/A AND2X1_LOC_418/a_8_24# 0.02fF
C44427 OR2X1_LOC_335/a_8_216# OR2X1_LOC_87/A 0.02fF
C44826 OR2X1_LOC_87/A AND2X1_LOC_591/a_8_24# 0.04fF
C45875 OR2X1_LOC_840/A OR2X1_LOC_87/A 0.14fF
C45927 AND2X1_LOC_145/a_8_24# OR2X1_LOC_87/A 0.05fF
C46331 OR2X1_LOC_216/A OR2X1_LOC_87/A 0.07fF
C46835 OR2X1_LOC_160/A OR2X1_LOC_87/A 0.22fF
C47157 OR2X1_LOC_87/A AND2X1_LOC_607/a_8_24# 0.02fF
C47693 OR2X1_LOC_87/A AND2X1_LOC_424/a_8_24# 0.04fF
C48172 OR2X1_LOC_185/A OR2X1_LOC_87/A 0.56fF
C48603 AND2X1_LOC_158/a_8_24# OR2X1_LOC_87/A 0.03fF
C49058 OR2X1_LOC_87/A AND2X1_LOC_442/a_8_24# 0.01fF
C49315 OR2X1_LOC_87/A OR2X1_LOC_641/A 0.08fF
C49375 AND2X1_LOC_312/a_8_24# OR2X1_LOC_87/A 0.04fF
C49450 OR2X1_LOC_114/Y OR2X1_LOC_87/A 0.12fF
C49459 OR2X1_LOC_87/A OR2X1_LOC_449/A 0.03fF
C50004 OR2X1_LOC_87/A OR2X1_LOC_446/A 0.02fF
C50073 OR2X1_LOC_87/A AND2X1_LOC_238/a_8_24# 0.03fF
C50098 OR2X1_LOC_335/a_36_216# OR2X1_LOC_87/A 0.02fF
C50317 OR2X1_LOC_643/A OR2X1_LOC_87/A 0.07fF
C50323 OR2X1_LOC_87/A OR2X1_LOC_778/Y 0.10fF
C50512 AND2X1_LOC_91/B OR2X1_LOC_87/A 0.03fF
C50892 OR2X1_LOC_87/A OR2X1_LOC_303/B 0.03fF
C51120 AND2X1_LOC_56/B OR2X1_LOC_87/A 5.13fF
C51259 OR2X1_LOC_87/A AND2X1_LOC_427/a_8_24# 0.04fF
C51977 OR2X1_LOC_87/A AND2X1_LOC_118/a_8_24# 0.01fF
C52473 OR2X1_LOC_87/A AND2X1_LOC_47/Y 0.14fF
C52657 AND2X1_LOC_521/a_8_24# OR2X1_LOC_87/A 0.04fF
C52784 OR2X1_LOC_506/A OR2X1_LOC_87/A 0.02fF
C52800 OR2X1_LOC_87/A AND2X1_LOC_695/a_8_24# 0.04fF
C52930 OR2X1_LOC_87/A OR2X1_LOC_227/Y -0.01fF
C53016 OR2X1_LOC_87/A OR2X1_LOC_180/B 0.55fF
C53241 OR2X1_LOC_87/A OR2X1_LOC_99/Y 0.03fF
C53418 OR2X1_LOC_87/A AND2X1_LOC_41/Y 0.03fF
C53894 OR2X1_LOC_87/A OR2X1_LOC_227/B 0.01fF
C54067 OR2X1_LOC_210/B OR2X1_LOC_87/A 0.01fF
C54403 OR2X1_LOC_235/B OR2X1_LOC_87/A 0.03fF
C54826 OR2X1_LOC_703/A OR2X1_LOC_87/A 0.03fF
C54894 OR2X1_LOC_116/a_8_216# OR2X1_LOC_87/A 0.02fF
C55297 AND2X1_LOC_316/a_36_24# OR2X1_LOC_87/A 0.01fF
C55524 OR2X1_LOC_87/A OR2X1_LOC_771/B 0.18fF
C55538 OR2X1_LOC_87/A OR2X1_LOC_776/A 0.16fF
C55972 OR2X1_LOC_87/A OR2X1_LOC_593/B 0.01fF
C56002 OR2X1_LOC_156/a_8_216# OR2X1_LOC_87/A 0.01fF
C56073 AND2X1_LOC_41/a_8_24# OR2X1_LOC_87/A 0.01fF
C57135 OR2X1_LOC_87/A VSS 0.90fF
C10640 OR2X1_LOC_80/Y OR2X1_LOC_393/Y 0.18fF
C15319 OR2X1_LOC_80/Y OR2X1_LOC_52/B 0.02fF
C18313 OR2X1_LOC_80/Y OR2X1_LOC_81/a_8_216# 0.18fF
C24697 OR2X1_LOC_81/Y OR2X1_LOC_80/Y 0.06fF
C29623 VDD OR2X1_LOC_80/Y 0.33fF
C32966 OR2X1_LOC_158/A OR2X1_LOC_80/Y 0.01fF
C35545 OR2X1_LOC_744/A OR2X1_LOC_80/Y 0.01fF
C41165 OR2X1_LOC_83/Y OR2X1_LOC_80/Y 0.54fF
C50129 OR2X1_LOC_80/Y OR2X1_LOC_16/A 0.02fF
C57157 OR2X1_LOC_80/Y VSS 0.26fF
C683 OR2X1_LOC_687/Y OR2X1_LOC_161/B 0.03fF
C1442 AND2X1_LOC_91/a_8_24# OR2X1_LOC_161/B 0.01fF
C1501 OR2X1_LOC_78/A OR2X1_LOC_161/B 0.54fF
C1557 OR2X1_LOC_602/A OR2X1_LOC_161/B 0.02fF
C2370 OR2X1_LOC_501/B OR2X1_LOC_161/B 0.07fF
C2403 OR2X1_LOC_147/B OR2X1_LOC_161/B 15.77fF
C2553 OR2X1_LOC_545/B OR2X1_LOC_161/B 0.01fF
C2643 OR2X1_LOC_318/B OR2X1_LOC_161/B 0.10fF
C2655 OR2X1_LOC_161/B OR2X1_LOC_854/A 0.14fF
C2811 OR2X1_LOC_538/A OR2X1_LOC_161/B 0.04fF
C3663 OR2X1_LOC_623/B OR2X1_LOC_161/B 0.03fF
C3822 OR2X1_LOC_544/A OR2X1_LOC_161/B 0.04fF
C4035 OR2X1_LOC_140/A OR2X1_LOC_161/B 0.01fF
C4093 OR2X1_LOC_254/B OR2X1_LOC_161/B 0.04fF
C4889 OR2X1_LOC_448/Y OR2X1_LOC_161/B 0.02fF
C5332 OR2X1_LOC_84/B OR2X1_LOC_161/B 0.13fF
C5641 OR2X1_LOC_186/Y OR2X1_LOC_161/B 0.06fF
C6212 OR2X1_LOC_574/A OR2X1_LOC_161/B 0.30fF
C6473 AND2X1_LOC_627/a_8_24# OR2X1_LOC_161/B 0.01fF
C6579 AND2X1_LOC_16/a_8_24# OR2X1_LOC_161/B 0.02fF
C6581 OR2X1_LOC_319/a_8_216# OR2X1_LOC_161/B 0.01fF
C7047 OR2X1_LOC_375/A OR2X1_LOC_161/B 0.41fF
C7402 OR2X1_LOC_161/B OR2X1_LOC_549/A 0.07fF
C7559 OR2X1_LOC_629/a_8_216# OR2X1_LOC_161/B 0.01fF
C7811 OR2X1_LOC_161/B OR2X1_LOC_161/a_8_216# 0.03fF
C7883 OR2X1_LOC_499/B OR2X1_LOC_161/B 0.01fF
C8142 OR2X1_LOC_543/a_8_216# OR2X1_LOC_161/B 0.02fF
C8177 OR2X1_LOC_161/B OR2X1_LOC_348/B 0.09fF
C9578 OR2X1_LOC_676/a_8_216# OR2X1_LOC_161/B 0.03fF
C9925 OR2X1_LOC_161/B OR2X1_LOC_712/B 0.01fF
C9962 OR2X1_LOC_139/A OR2X1_LOC_161/B 0.22fF
C10893 AND2X1_LOC_315/a_8_24# OR2X1_LOC_161/B 0.05fF
C11076 OR2X1_LOC_247/a_8_216# OR2X1_LOC_161/B 0.01fF
C11323 OR2X1_LOC_703/B OR2X1_LOC_161/B 0.04fF
C12489 OR2X1_LOC_97/A OR2X1_LOC_161/B 0.01fF
C12962 OR2X1_LOC_161/B OR2X1_LOC_713/A 0.15fF
C13034 OR2X1_LOC_629/Y OR2X1_LOC_161/B 0.02fF
C13684 OR2X1_LOC_543/a_36_216# OR2X1_LOC_161/B 0.02fF
C13926 OR2X1_LOC_154/A OR2X1_LOC_161/B 0.20fF
C13936 OR2X1_LOC_267/A OR2X1_LOC_161/B 0.01fF
C13971 OR2X1_LOC_778/A OR2X1_LOC_161/B 0.01fF
C14339 OR2X1_LOC_267/a_8_216# OR2X1_LOC_161/B 0.15fF
C14656 OR2X1_LOC_361/a_8_216# OR2X1_LOC_161/B 0.02fF
C14702 OR2X1_LOC_538/a_8_216# OR2X1_LOC_161/B 0.01fF
C15042 OR2X1_LOC_267/Y OR2X1_LOC_161/B 0.06fF
C15654 AND2X1_LOC_600/a_8_24# OR2X1_LOC_161/B 0.01fF
C16080 AND2X1_LOC_677/a_8_24# OR2X1_LOC_161/B 0.04fF
C16742 OR2X1_LOC_614/Y OR2X1_LOC_161/B 0.01fF
C17589 OR2X1_LOC_450/A OR2X1_LOC_161/B 0.24fF
C17784 OR2X1_LOC_532/B OR2X1_LOC_161/B 1.81fF
C17795 AND2X1_LOC_665/a_8_24# OR2X1_LOC_161/B 0.01fF
C18458 OR2X1_LOC_162/Y OR2X1_LOC_161/B 0.01fF
C19191 OR2X1_LOC_552/A OR2X1_LOC_161/B 0.03fF
C19775 VDD OR2X1_LOC_161/B 2.21fF
C20442 OR2X1_LOC_161/B AND2X1_LOC_418/a_8_24# 0.01fF
C20624 OR2X1_LOC_676/Y OR2X1_LOC_161/B 0.01fF
C20644 OR2X1_LOC_834/A OR2X1_LOC_161/B 0.01fF
C20714 OR2X1_LOC_483/a_8_216# OR2X1_LOC_161/B 0.01fF
C21247 OR2X1_LOC_602/B OR2X1_LOC_161/B 0.02fF
C21870 OR2X1_LOC_115/B OR2X1_LOC_161/B 0.08fF
C21954 OR2X1_LOC_840/A OR2X1_LOC_161/B 0.05fF
C22440 OR2X1_LOC_457/B OR2X1_LOC_161/B 0.03fF
C22543 AND2X1_LOC_134/a_8_24# OR2X1_LOC_161/B 0.11fF
C22828 OR2X1_LOC_809/B OR2X1_LOC_161/B 0.02fF
C22878 OR2X1_LOC_160/A OR2X1_LOC_161/B 0.17fF
C23210 OR2X1_LOC_450/B OR2X1_LOC_161/B 0.25fF
C24029 AND2X1_LOC_163/a_8_24# OR2X1_LOC_161/B 0.02fF
C24110 OR2X1_LOC_185/A OR2X1_LOC_161/B 0.73fF
C24565 OR2X1_LOC_702/A OR2X1_LOC_161/B 0.03fF
C24968 AND2X1_LOC_481/a_8_24# OR2X1_LOC_161/B 0.01fF
C25250 OR2X1_LOC_294/Y OR2X1_LOC_161/B 0.07fF
C25270 OR2X1_LOC_641/A OR2X1_LOC_161/B 0.29fF
C25369 OR2X1_LOC_114/Y OR2X1_LOC_161/B 0.02fF
C25375 OR2X1_LOC_449/A OR2X1_LOC_161/B 0.06fF
C25921 OR2X1_LOC_161/B OR2X1_LOC_446/A 0.03fF
C26206 OR2X1_LOC_643/A OR2X1_LOC_161/B 0.03fF
C26212 OR2X1_LOC_778/Y OR2X1_LOC_161/B 0.10fF
C26470 AND2X1_LOC_91/B OR2X1_LOC_161/B 0.71fF
C26579 AND2X1_LOC_72/Y OR2X1_LOC_161/B 0.01fF
C26848 OR2X1_LOC_161/B OR2X1_LOC_303/B 0.07fF
C26934 OR2X1_LOC_161/B OR2X1_LOC_719/B 0.01fF
C26955 OR2X1_LOC_542/B OR2X1_LOC_161/B 0.03fF
C27015 OR2X1_LOC_631/a_8_216# OR2X1_LOC_161/B 0.02fF
C27052 AND2X1_LOC_56/B OR2X1_LOC_161/B 0.27fF
C27261 AND2X1_LOC_427/a_8_24# OR2X1_LOC_161/B 0.15fF
C27446 AND2X1_LOC_315/a_36_24# OR2X1_LOC_161/B 0.01fF
C27882 OR2X1_LOC_457/a_8_216# OR2X1_LOC_161/B 0.05fF
C28435 AND2X1_LOC_47/Y OR2X1_LOC_161/B 0.84fF
C28586 OR2X1_LOC_161/B OR2X1_LOC_186/a_8_216# 0.01fF
C28700 OR2X1_LOC_506/A OR2X1_LOC_161/B 0.21fF
C28710 AND2X1_LOC_695/a_8_24# OR2X1_LOC_161/B 0.01fF
C28828 OR2X1_LOC_780/A OR2X1_LOC_161/B 0.04fF
C28861 AND2X1_LOC_420/a_8_24# OR2X1_LOC_161/B 0.02fF
C29392 OR2X1_LOC_161/B OR2X1_LOC_788/B 0.01fF
C29465 OR2X1_LOC_467/B OR2X1_LOC_161/B 0.04fF
C29545 OR2X1_LOC_630/a_8_216# OR2X1_LOC_161/B 0.02fF
C29554 OR2X1_LOC_664/a_8_216# OR2X1_LOC_161/B 0.01fF
C29878 OR2X1_LOC_161/B OR2X1_LOC_162/A 0.02fF
C30357 OR2X1_LOC_235/B OR2X1_LOC_161/B 0.03fF
C30777 OR2X1_LOC_703/A OR2X1_LOC_161/B 0.03fF
C31173 OR2X1_LOC_362/A OR2X1_LOC_161/B 0.01fF
C31222 OR2X1_LOC_539/A OR2X1_LOC_161/B 0.01fF
C32142 OR2X1_LOC_254/a_8_216# OR2X1_LOC_161/B 0.04fF
C32359 AND2X1_LOC_44/Y OR2X1_LOC_161/B 0.70fF
C32622 OR2X1_LOC_720/B OR2X1_LOC_161/B 0.14fF
C33101 OR2X1_LOC_247/Y OR2X1_LOC_161/B 0.01fF
C33276 AND2X1_LOC_18/Y OR2X1_LOC_161/B 0.21fF
C33606 OR2X1_LOC_161/B OR2X1_LOC_789/A 0.03fF
C33712 OR2X1_LOC_307/A OR2X1_LOC_161/B 0.25fF
C34192 OR2X1_LOC_707/A OR2X1_LOC_161/B 0.03fF
C34638 OR2X1_LOC_449/B OR2X1_LOC_161/B 9.84fF
C35799 OR2X1_LOC_786/A OR2X1_LOC_161/B 0.03fF
C35931 OR2X1_LOC_555/A OR2X1_LOC_161/B 0.05fF
C36002 OR2X1_LOC_447/Y OR2X1_LOC_161/B 0.12fF
C36368 AND2X1_LOC_51/Y OR2X1_LOC_161/B 0.70fF
C37039 OR2X1_LOC_439/B OR2X1_LOC_161/B 0.01fF
C37156 OR2X1_LOC_631/B OR2X1_LOC_161/B 0.43fF
C37204 AND2X1_LOC_135/a_8_24# OR2X1_LOC_161/B 0.01fF
C37530 AND2X1_LOC_253/a_8_24# OR2X1_LOC_161/B 0.06fF
C37957 OR2X1_LOC_632/A OR2X1_LOC_161/B 0.03fF
C38072 AND2X1_LOC_677/a_36_24# OR2X1_LOC_161/B 0.01fF
C38211 AND2X1_LOC_427/a_36_24# OR2X1_LOC_161/B 0.01fF
C38224 OR2X1_LOC_161/B OR2X1_LOC_71/A 0.01fF
C38639 AND2X1_LOC_31/Y OR2X1_LOC_161/B 0.77fF
C38881 AND2X1_LOC_597/a_8_24# OR2X1_LOC_161/B 0.01fF
C39262 AND2X1_LOC_305/a_8_24# OR2X1_LOC_161/B 0.09fF
C39480 OR2X1_LOC_161/B OR2X1_LOC_451/B 0.02fF
C39568 AND2X1_LOC_36/Y OR2X1_LOC_161/B 0.20fF
C39646 OR2X1_LOC_630/Y OR2X1_LOC_161/B 0.01fF
C39672 OR2X1_LOC_635/A OR2X1_LOC_161/B 0.46fF
C39839 OR2X1_LOC_780/a_8_216# OR2X1_LOC_161/B 0.02fF
C40044 AND2X1_LOC_167/a_8_24# OR2X1_LOC_161/B 0.01fF
C40851 OR2X1_LOC_161/B OR2X1_LOC_160/Y 0.02fF
C42590 OR2X1_LOC_161/B OR2X1_LOC_319/Y 0.01fF
C42991 OR2X1_LOC_161/B OR2X1_LOC_777/B 0.10fF
C43061 OR2X1_LOC_344/A OR2X1_LOC_161/B 0.03fF
C43129 OR2X1_LOC_254/A OR2X1_LOC_161/B 0.01fF
C43215 AND2X1_LOC_13/a_8_24# OR2X1_LOC_161/B 0.01fF
C43854 OR2X1_LOC_161/B OR2X1_LOC_707/a_8_216# 0.01fF
C43972 OR2X1_LOC_630/B OR2X1_LOC_161/B 0.02fF
C44469 OR2X1_LOC_644/B OR2X1_LOC_161/B -0.02fF
C44923 AND2X1_LOC_72/a_8_24# OR2X1_LOC_161/B 0.01fF
C46166 OR2X1_LOC_319/B OR2X1_LOC_161/B 0.61fF
C46263 OR2X1_LOC_296/Y OR2X1_LOC_161/B 0.01fF
C47176 OR2X1_LOC_629/A OR2X1_LOC_161/B 0.13fF
C47268 OR2X1_LOC_446/Y OR2X1_LOC_161/B 0.25fF
C47303 OR2X1_LOC_473/A OR2X1_LOC_161/B 0.31fF
C48014 OR2X1_LOC_553/A OR2X1_LOC_161/B 0.07fF
C48021 OR2X1_LOC_266/a_8_216# OR2X1_LOC_161/B 0.01fF
C48747 OR2X1_LOC_151/A OR2X1_LOC_161/B 0.24fF
C49146 OR2X1_LOC_161/B AND2X1_LOC_279/a_8_24# 0.11fF
C50036 OR2X1_LOC_631/A OR2X1_LOC_161/B 0.02fF
C50419 OR2X1_LOC_168/Y OR2X1_LOC_161/B 0.03fF
C51085 OR2X1_LOC_783/A OR2X1_LOC_161/B 0.01fF
C51219 OR2X1_LOC_161/B OR2X1_LOC_308/Y 0.07fF
C51795 OR2X1_LOC_664/Y OR2X1_LOC_161/B 0.35fF
C52094 OR2X1_LOC_161/B OR2X1_LOC_162/a_8_216# 0.01fF
C52257 OR2X1_LOC_446/a_8_216# OR2X1_LOC_161/B 0.01fF
C53427 AND2X1_LOC_311/a_8_24# OR2X1_LOC_161/B 0.01fF
C53838 OR2X1_LOC_190/A OR2X1_LOC_161/B 0.03fF
C54182 OR2X1_LOC_188/Y OR2X1_LOC_161/B 0.03fF
C54376 OR2X1_LOC_193/A OR2X1_LOC_161/B 0.18fF
C54630 AND2X1_LOC_438/a_8_24# OR2X1_LOC_161/B 0.01fF
C54648 OR2X1_LOC_598/Y OR2X1_LOC_161/B 0.05fF
C54672 OR2X1_LOC_335/Y OR2X1_LOC_161/B 0.02fF
C55608 OR2X1_LOC_810/A OR2X1_LOC_161/B 0.10fF
C55611 OR2X1_LOC_307/a_8_216# OR2X1_LOC_161/B 0.06fF
C55941 OR2X1_LOC_715/B OR2X1_LOC_161/B 0.03fF
C55953 OR2X1_LOC_543/A OR2X1_LOC_161/B 0.03fF
C56455 OR2X1_LOC_161/B VSS 1.07fF
C1473 OR2X1_LOC_135/Y OR2X1_LOC_589/A 0.02fF
C1814 OR2X1_LOC_589/A OR2X1_LOC_536/a_8_216# 0.01fF
C2364 OR2X1_LOC_597/A OR2X1_LOC_589/A 0.07fF
C2778 OR2X1_LOC_589/A OR2X1_LOC_829/A 0.80fF
C3053 OR2X1_LOC_589/A OR2X1_LOC_597/Y 0.04fF
C3342 OR2X1_LOC_589/A OR2X1_LOC_385/Y 0.01fF
C4909 AND2X1_LOC_729/Y OR2X1_LOC_589/A 0.03fF
C5357 OR2X1_LOC_589/A OR2X1_LOC_52/B 0.08fF
C6528 OR2X1_LOC_589/A OR2X1_LOC_536/Y 0.01fF
C8835 OR2X1_LOC_589/A AND2X1_LOC_266/Y 0.15fF
C9640 OR2X1_LOC_589/A OR2X1_LOC_265/a_8_216# 0.01fF
C10962 OR2X1_LOC_589/A OR2X1_LOC_74/A 0.03fF
C11314 OR2X1_LOC_589/A OR2X1_LOC_432/a_8_216# 0.03fF
C11770 OR2X1_LOC_589/A OR2X1_LOC_432/Y 0.02fF
C12105 OR2X1_LOC_589/A AND2X1_LOC_537/a_8_24# 0.01fF
C12520 AND2X1_LOC_339/B OR2X1_LOC_589/A 0.02fF
C13447 OR2X1_LOC_589/A OR2X1_LOC_597/a_8_216# 0.11fF
C13710 OR2X1_LOC_589/A OR2X1_LOC_72/Y 0.22fF
C14660 AND2X1_LOC_706/Y OR2X1_LOC_589/A 0.11fF
C16436 OR2X1_LOC_589/A OR2X1_LOC_69/Y 0.30fF
C16514 OR2X1_LOC_589/A AND2X1_LOC_537/Y 0.01fF
C17277 OR2X1_LOC_589/A OR2X1_LOC_433/Y 0.03fF
C17284 OR2X1_LOC_589/A AND2X1_LOC_138/a_8_24# 0.17fF
C19794 VDD OR2X1_LOC_589/A 0.85fF
C19851 OR2X1_LOC_589/A OR2X1_LOC_829/a_8_216# 0.05fF
C19894 OR2X1_LOC_589/A AND2X1_LOC_267/a_8_24# 0.01fF
C20805 OR2X1_LOC_589/A AND2X1_LOC_307/Y 0.03fF
C21679 OR2X1_LOC_589/A OR2X1_LOC_416/Y 0.02fF
C22470 OR2X1_LOC_589/A AND2X1_LOC_831/a_8_24# 0.17fF
C22789 OR2X1_LOC_45/B OR2X1_LOC_589/A 0.19fF
C22894 OR2X1_LOC_589/A AND2X1_LOC_435/a_8_24# 0.02fF
C23201 OR2X1_LOC_158/A OR2X1_LOC_589/A 0.03fF
C25366 OR2X1_LOC_589/A OR2X1_LOC_316/Y 0.02fF
C25412 OR2X1_LOC_589/A AND2X1_LOC_390/B 0.07fF
C25718 OR2X1_LOC_589/A OR2X1_LOC_744/A 0.40fF
C26035 OR2X1_LOC_589/A OR2X1_LOC_320/a_8_216# 0.07fF
C27552 OR2X1_LOC_589/A OR2X1_LOC_311/Y 0.03fF
C28032 OR2X1_LOC_589/A AND2X1_LOC_831/Y 0.50fF
C28333 OR2X1_LOC_589/A AND2X1_LOC_436/B 0.09fF
C28339 OR2X1_LOC_589/A AND2X1_LOC_139/B 0.23fF
C29290 OR2X1_LOC_589/A OR2X1_LOC_409/B 0.16fF
C30436 OR2X1_LOC_589/A AND2X1_LOC_319/A 0.19fF
C30882 OR2X1_LOC_589/A AND2X1_LOC_361/A 0.01fF
C32391 OR2X1_LOC_589/A AND2X1_LOC_729/a_8_24# 0.02fF
C32491 OR2X1_LOC_589/A OR2X1_LOC_619/Y 0.10fF
C34592 OR2X1_LOC_589/A OR2X1_LOC_393/a_8_216# 0.39fF
C34915 OR2X1_LOC_589/A OR2X1_LOC_13/B 1.41fF
C35344 OR2X1_LOC_589/A OR2X1_LOC_595/A 0.16fF
C36364 OR2X1_LOC_589/A OR2X1_LOC_89/A 0.07fF
C37284 OR2X1_LOC_589/A OR2X1_LOC_95/Y 0.03fF
C38496 OR2X1_LOC_70/Y OR2X1_LOC_589/A 0.97fF
C40008 OR2X1_LOC_589/A OR2X1_LOC_16/A 0.06fF
C40214 OR2X1_LOC_589/A AND2X1_LOC_687/Y 0.28fF
C41012 OR2X1_LOC_589/A OR2X1_LOC_262/a_8_216# 0.01fF
C41065 OR2X1_LOC_589/A AND2X1_LOC_729/B 0.08fF
C41578 OR2X1_LOC_589/A AND2X1_LOC_227/Y 0.05fF
C41896 OR2X1_LOC_599/A OR2X1_LOC_589/A 0.49fF
C42206 OR2X1_LOC_40/Y OR2X1_LOC_589/A 0.11fF
C42355 OR2X1_LOC_589/A OR2X1_LOC_7/A 0.03fF
C42376 OR2X1_LOC_589/A OR2X1_LOC_320/Y 0.14fF
C44528 OR2X1_LOC_3/Y OR2X1_LOC_589/A 0.02fF
C45475 OR2X1_LOC_589/A OR2X1_LOC_72/a_8_216# 0.01fF
C45855 OR2X1_LOC_589/A OR2X1_LOC_64/Y 0.14fF
C49170 OR2X1_LOC_589/A AND2X1_LOC_130/a_8_24# 0.11fF
C49175 OR2X1_LOC_589/A AND2X1_LOC_729/a_36_24# 0.01fF
C52251 OR2X1_LOC_589/A OR2X1_LOC_262/Y 0.17fF
C53512 OR2X1_LOC_306/Y OR2X1_LOC_589/A 0.03fF
C53912 OR2X1_LOC_589/A OR2X1_LOC_265/Y 0.22fF
C54437 OR2X1_LOC_589/A AND2X1_LOC_633/Y 0.02fF
C54619 AND2X1_LOC_539/Y OR2X1_LOC_589/A 0.03fF
C54658 OR2X1_LOC_589/A OR2X1_LOC_131/A 0.03fF
C55531 OR2X1_LOC_589/A AND2X1_LOC_434/Y 0.07fF
C57645 OR2X1_LOC_589/A VSS 0.93fF
C10454 AND2X1_LOC_789/a_8_24# OR2X1_LOC_748/Y 0.23fF
C29029 VDD OR2X1_LOC_748/Y 0.12fF
C41753 OR2X1_LOC_600/A OR2X1_LOC_748/Y 0.01fF
C53911 OR2X1_LOC_3/Y OR2X1_LOC_748/Y 0.02fF
C56419 OR2X1_LOC_748/Y VSS 0.06fF
C1964 OR2X1_LOC_147/B OR2X1_LOC_344/A 0.03fF
C3689 OR2X1_LOC_833/B OR2X1_LOC_344/A 0.02fF
C3711 OR2X1_LOC_254/B OR2X1_LOC_344/A 0.01fF
C6962 OR2X1_LOC_344/A OR2X1_LOC_549/A 0.08fF
C17389 OR2X1_LOC_532/B OR2X1_LOC_344/A 0.03fF
C19344 VDD OR2X1_LOC_344/A 0.35fF
C23693 OR2X1_LOC_185/A OR2X1_LOC_344/A 0.02fF
C26522 OR2X1_LOC_344/A OR2X1_LOC_719/B 0.02fF
C26534 OR2X1_LOC_542/B OR2X1_LOC_344/A 0.03fF
C26620 AND2X1_LOC_56/B OR2X1_LOC_344/A 0.04fF
C32852 AND2X1_LOC_18/Y OR2X1_LOC_344/A 0.04fF
C39145 OR2X1_LOC_344/A AND2X1_LOC_36/Y 0.12fF
C42829 OR2X1_LOC_456/A OR2X1_LOC_344/A 0.20fF
C48825 AND2X1_LOC_482/a_8_24# OR2X1_LOC_344/A 0.01fF
C49297 AND2X1_LOC_252/a_8_24# OR2X1_LOC_344/A 0.01fF
C53414 OR2X1_LOC_190/A OR2X1_LOC_344/A 0.07fF
C56506 OR2X1_LOC_344/A VSS -0.05fF
C297 OR2X1_LOC_135/Y OR2X1_LOC_7/A 0.07fF
C438 OR2X1_LOC_7/A AND2X1_LOC_848/Y 0.07fF
C445 AND2X1_LOC_154/a_36_24# OR2X1_LOC_7/A 0.01fF
C814 AND2X1_LOC_160/a_8_24# OR2X1_LOC_7/A 0.05fF
C1249 OR2X1_LOC_178/Y OR2X1_LOC_7/A 0.04fF
C1681 OR2X1_LOC_697/a_8_216# OR2X1_LOC_7/A -0.04fF
C2222 OR2X1_LOC_385/Y OR2X1_LOC_7/A 0.68fF
C2489 OR2X1_LOC_7/A AND2X1_LOC_810/B 0.07fF
C2884 OR2X1_LOC_7/A OR2X1_LOC_230/Y 0.02fF
C2888 OR2X1_LOC_7/A OR2X1_LOC_368/Y 0.18fF
C2916 OR2X1_LOC_229/a_8_216# OR2X1_LOC_7/A -0.03fF
C3494 OR2X1_LOC_7/A OR2X1_LOC_754/a_8_216# 0.03fF
C3737 OR2X1_LOC_7/A OR2X1_LOC_323/Y 0.08fF
C3877 AND2X1_LOC_729/Y OR2X1_LOC_7/A 0.07fF
C3907 AND2X1_LOC_784/A OR2X1_LOC_7/A 0.07fF
C4286 OR2X1_LOC_7/A OR2X1_LOC_52/B 4.28fF
C4391 OR2X1_LOC_7/A AND2X1_LOC_216/A 0.15fF
C4715 OR2X1_LOC_280/Y OR2X1_LOC_7/A 0.07fF
C5334 OR2X1_LOC_7/A OR2X1_LOC_744/Y 0.01fF
C5393 OR2X1_LOC_536/Y OR2X1_LOC_7/A 0.03fF
C5605 OR2X1_LOC_226/Y OR2X1_LOC_7/A 0.03fF
C5864 OR2X1_LOC_51/Y OR2X1_LOC_7/A 2.92fF
C6385 OR2X1_LOC_423/a_8_216# OR2X1_LOC_7/A 0.10fF
C6427 AND2X1_LOC_802/a_8_24# OR2X1_LOC_7/A 0.02fF
C6496 OR2X1_LOC_7/A AND2X1_LOC_790/a_8_24# 0.03fF
C6696 OR2X1_LOC_178/a_8_216# OR2X1_LOC_7/A 0.01fF
C6710 OR2X1_LOC_7/A AND2X1_LOC_436/Y 0.03fF
C6751 AND2X1_LOC_344/a_8_24# OR2X1_LOC_7/A 0.04fF
C7236 OR2X1_LOC_252/Y OR2X1_LOC_7/A 0.17fF
C7906 OR2X1_LOC_7/A OR2X1_LOC_183/Y 0.35fF
C8150 OR2X1_LOC_248/a_8_216# OR2X1_LOC_7/A 0.01fF
C8919 AND2X1_LOC_391/Y OR2X1_LOC_7/A 0.07fF
C9045 OR2X1_LOC_7/A OR2X1_LOC_27/Y 0.15fF
C9599 OR2X1_LOC_7/A OR2X1_LOC_423/Y 0.05fF
C9900 OR2X1_LOC_74/A OR2X1_LOC_7/A 0.25fF
C10156 OR2X1_LOC_7/A AND2X1_LOC_254/a_8_24# 0.07fF
C10570 OR2X1_LOC_7/A AND2X1_LOC_448/a_8_24# 0.05fF
C10982 AND2X1_LOC_537/a_8_24# OR2X1_LOC_7/A 0.05fF
C11146 OR2X1_LOC_615/a_8_216# OR2X1_LOC_7/A 0.03fF
C11381 OR2X1_LOC_482/a_8_216# OR2X1_LOC_7/A 0.09fF
C12276 OR2X1_LOC_7/A AND2X1_LOC_614/a_8_24# 0.01fF
C12743 OR2X1_LOC_697/Y OR2X1_LOC_7/A 0.03fF
C12869 OR2X1_LOC_696/Y OR2X1_LOC_7/A 0.01fF
C13070 OR2X1_LOC_7/A OR2X1_LOC_503/a_8_216# 0.01fF
C13531 AND2X1_LOC_706/Y OR2X1_LOC_7/A 0.07fF
C13705 OR2X1_LOC_665/Y OR2X1_LOC_7/A 0.03fF
C14476 OR2X1_LOC_695/a_8_216# OR2X1_LOC_7/A 0.04fF
C14509 AND2X1_LOC_302/a_8_24# OR2X1_LOC_7/A 0.02fF
C15091 OR2X1_LOC_7/A OR2X1_LOC_589/Y 0.03fF
C15387 AND2X1_LOC_537/Y OR2X1_LOC_7/A 4.03fF
C15548 OR2X1_LOC_7/A OR2X1_LOC_743/Y 0.02fF
C16459 AND2X1_LOC_714/B OR2X1_LOC_7/A 0.23fF
C16922 OR2X1_LOC_482/a_36_216# OR2X1_LOC_7/A 0.03fF
C17587 OR2X1_LOC_7/A AND2X1_LOC_793/B 0.01fF
C17747 OR2X1_LOC_368/a_8_216# OR2X1_LOC_7/A 0.03fF
C17810 AND2X1_LOC_348/A OR2X1_LOC_7/A 0.03fF
C18378 OR2X1_LOC_131/Y OR2X1_LOC_7/A 0.03fF
C18657 VDD OR2X1_LOC_7/A 0.91fF
C18763 OR2X1_LOC_315/Y OR2X1_LOC_7/A 0.49fF
C18885 OR2X1_LOC_7/A OR2X1_LOC_67/Y 0.03fF
C19195 OR2X1_LOC_248/Y OR2X1_LOC_7/A 0.78fF
C19208 OR2X1_LOC_666/Y OR2X1_LOC_7/A 0.02fF
C19877 OR2X1_LOC_494/A OR2X1_LOC_7/A 0.01fF
C21608 OR2X1_LOC_45/B OR2X1_LOC_7/A 0.96fF
C22064 OR2X1_LOC_158/A OR2X1_LOC_7/A 0.28fF
C22100 AND2X1_LOC_537/a_36_24# OR2X1_LOC_7/A 0.01fF
C22146 AND2X1_LOC_98/Y OR2X1_LOC_7/A 0.02fF
C22508 OR2X1_LOC_482/Y OR2X1_LOC_7/A 0.06fF
C24342 AND2X1_LOC_390/B OR2X1_LOC_7/A 0.14fF
C24585 OR2X1_LOC_309/Y OR2X1_LOC_7/A 0.03fF
C24631 OR2X1_LOC_744/A OR2X1_LOC_7/A 0.52fF
C25014 OR2X1_LOC_694/Y OR2X1_LOC_7/A 0.02fF
C25392 OR2X1_LOC_7/A OR2X1_LOC_522/Y 0.14fF
C25478 OR2X1_LOC_179/a_8_216# OR2X1_LOC_7/A 0.02fF
C25542 AND2X1_LOC_303/B OR2X1_LOC_7/A -0.02fF
C26273 OR2X1_LOC_7/A AND2X1_LOC_285/Y 0.03fF
C26351 OR2X1_LOC_91/Y OR2X1_LOC_7/A 0.10fF
C26368 OR2X1_LOC_305/Y OR2X1_LOC_7/A 0.03fF
C26424 OR2X1_LOC_417/Y OR2X1_LOC_7/A 0.07fF
C26432 OR2X1_LOC_311/Y OR2X1_LOC_7/A 0.03fF
C26500 AND2X1_LOC_483/Y OR2X1_LOC_7/A 0.56fF
C26587 OR2X1_LOC_7/A AND2X1_LOC_780/a_8_24# 0.04fF
C26592 OR2X1_LOC_7/A OR2X1_LOC_171/Y 0.03fF
C26736 OR2X1_LOC_494/a_8_216# OR2X1_LOC_7/A 0.03fF
C27139 OR2X1_LOC_7/A AND2X1_LOC_448/a_36_24# 0.01fF
C27229 OR2X1_LOC_7/A AND2X1_LOC_436/B 0.07fF
C27950 OR2X1_LOC_108/a_8_216# OR2X1_LOC_7/A 0.01fF
C28444 OR2X1_LOC_298/a_8_216# OR2X1_LOC_7/A 0.01fF
C28505 OR2X1_LOC_497/Y OR2X1_LOC_7/A 0.07fF
C28529 OR2X1_LOC_7/A OR2X1_LOC_229/Y 0.03fF
C29327 AND2X1_LOC_319/A OR2X1_LOC_7/A 0.07fF
C29374 OR2X1_LOC_52/a_8_216# OR2X1_LOC_7/A 0.02fF
C29395 AND2X1_LOC_708/a_8_24# OR2X1_LOC_7/A 0.09fF
C29443 AND2X1_LOC_721/A OR2X1_LOC_7/A 0.03fF
C29474 OR2X1_LOC_7/A OR2X1_LOC_331/Y 0.03fF
C29778 OR2X1_LOC_7/A AND2X1_LOC_361/A 0.09fF
C30491 OR2X1_LOC_695/Y OR2X1_LOC_7/A 0.01fF
C31346 OR2X1_LOC_600/A OR2X1_LOC_7/A 0.41fF
C31383 AND2X1_LOC_543/a_8_24# OR2X1_LOC_7/A 0.01fF
C31419 OR2X1_LOC_7/A OR2X1_LOC_619/Y 0.28fF
C31862 OR2X1_LOC_7/A AND2X1_LOC_454/A 0.29fF
C31912 AND2X1_LOC_539/a_8_24# OR2X1_LOC_7/A 0.06fF
C32053 OR2X1_LOC_7/A AND2X1_LOC_783/B 0.01fF
C33607 OR2X1_LOC_312/Y OR2X1_LOC_7/A 0.03fF
C33632 AND2X1_LOC_307/a_8_24# OR2X1_LOC_7/A 0.06fF
C33745 OR2X1_LOC_7/A OR2X1_LOC_13/B 0.84fF
C34233 OR2X1_LOC_7/A OR2X1_LOC_595/A 0.07fF
C34358 AND2X1_LOC_154/a_8_24# OR2X1_LOC_7/A 0.07fF
C34686 OR2X1_LOC_528/Y OR2X1_LOC_7/A 0.14fF
C34831 AND2X1_LOC_342/Y OR2X1_LOC_7/A 0.08fF
C34886 AND2X1_LOC_483/a_8_24# OR2X1_LOC_7/A 0.18fF
C34909 AND2X1_LOC_712/B OR2X1_LOC_7/A 0.17fF
C35114 OR2X1_LOC_7/A OR2X1_LOC_765/Y 0.02fF
C35250 OR2X1_LOC_89/A OR2X1_LOC_7/A 0.35fF
C35978 AND2X1_LOC_707/a_8_24# OR2X1_LOC_7/A 0.03fF
C36119 OR2X1_LOC_488/Y OR2X1_LOC_7/A 0.10fF
C36143 AND2X1_LOC_727/A OR2X1_LOC_7/A 0.03fF
C36165 OR2X1_LOC_95/Y OR2X1_LOC_7/A 0.71fF
C36435 OR2X1_LOC_179/Y OR2X1_LOC_7/A 0.01fF
C36873 OR2X1_LOC_7/A AND2X1_LOC_621/Y 0.11fF
C37385 OR2X1_LOC_70/Y OR2X1_LOC_7/A 0.15fF
C38468 OR2X1_LOC_7/A OR2X1_LOC_584/a_8_216# 0.02fF
C38493 AND2X1_LOC_535/Y OR2X1_LOC_7/A 0.03fF
C38618 OR2X1_LOC_246/Y OR2X1_LOC_7/A 0.03fF
C38905 OR2X1_LOC_7/A OR2X1_LOC_16/A 14.31fF
C38948 OR2X1_LOC_108/Y OR2X1_LOC_7/A 0.50fF
C39811 OR2X1_LOC_7/A AND2X1_LOC_447/Y 0.01fF
C39882 OR2X1_LOC_109/Y OR2X1_LOC_7/A 0.03fF
C39888 OR2X1_LOC_7/A AND2X1_LOC_448/Y 0.02fF
C39937 AND2X1_LOC_729/B OR2X1_LOC_7/A 0.19fF
C40352 AND2X1_LOC_798/Y OR2X1_LOC_7/A 0.05fF
C40368 AND2X1_LOC_708/a_36_24# OR2X1_LOC_7/A 0.01fF
C40398 AND2X1_LOC_227/Y OR2X1_LOC_7/A 0.13fF
C40428 OR2X1_LOC_813/Y OR2X1_LOC_7/A 0.07fF
C40737 OR2X1_LOC_599/A OR2X1_LOC_7/A 0.06fF
C41048 OR2X1_LOC_40/Y OR2X1_LOC_7/A 0.21fF
C41264 OR2X1_LOC_224/a_8_216# OR2X1_LOC_7/A 0.01fF
C41731 OR2X1_LOC_7/A OR2X1_LOC_615/Y 0.15fF
C41802 OR2X1_LOC_7/A OR2X1_LOC_424/Y -0.03fF
C41886 AND2X1_LOC_707/Y OR2X1_LOC_7/A 0.19fF
C42012 AND2X1_LOC_841/B OR2X1_LOC_7/A 9.11fF
C42298 AND2X1_LOC_543/Y OR2X1_LOC_7/A 0.01fF
C42363 OR2X1_LOC_7/A OR2X1_LOC_322/Y 0.51fF
C43171 OR2X1_LOC_7/A AND2X1_LOC_780/a_36_24# 0.01fF
C43391 OR2X1_LOC_3/Y OR2X1_LOC_7/A 6.85fF
C44492 OR2X1_LOC_7/A OR2X1_LOC_766/a_8_216# 0.05fF
C44700 OR2X1_LOC_64/Y OR2X1_LOC_7/A 0.53fF
C44838 OR2X1_LOC_7/A AND2X1_LOC_247/a_8_24# 0.03fF
C45113 AND2X1_LOC_101/B OR2X1_LOC_7/A 0.73fF
C45606 OR2X1_LOC_7/A OR2X1_LOC_7/Y 1.75fF
C46352 AND2X1_LOC_456/B OR2X1_LOC_7/A 0.31fF
C46715 OR2X1_LOC_7/A AND2X1_LOC_828/a_8_24# 0.06fF
C47231 OR2X1_LOC_494/Y OR2X1_LOC_7/A 0.03fF
C47245 AND2X1_LOC_707/a_36_24# OR2X1_LOC_7/A 0.01fF
C47620 OR2X1_LOC_7/A AND2X1_LOC_802/Y 0.07fF
C47807 AND2X1_LOC_154/Y OR2X1_LOC_7/A 0.22fF
C48075 AND2X1_LOC_130/a_8_24# OR2X1_LOC_7/A 0.03fF
C48206 OR2X1_LOC_7/A AND2X1_LOC_624/A 0.06fF
C49515 OR2X1_LOC_48/Y OR2X1_LOC_7/A 0.21fF
C49764 OR2X1_LOC_7/A OR2X1_LOC_584/a_36_216# 0.02fF
C49810 AND2X1_LOC_160/Y OR2X1_LOC_7/A 0.03fF
C50171 OR2X1_LOC_7/A OR2X1_LOC_421/Y 0.26fF
C50500 OR2X1_LOC_7/A OR2X1_LOC_504/a_8_216# 0.07fF
C50563 OR2X1_LOC_7/A OR2X1_LOC_744/a_8_216# 0.04fF
C50782 OR2X1_LOC_754/A OR2X1_LOC_7/A 0.09fF
C51118 OR2X1_LOC_7/A OR2X1_LOC_118/Y 0.03fF
C51605 OR2X1_LOC_52/Y OR2X1_LOC_7/A 0.11fF
C51650 OR2X1_LOC_503/Y OR2X1_LOC_7/A 0.01fF
C51703 OR2X1_LOC_7/A OR2X1_LOC_754/Y 0.05fF
C52290 OR2X1_LOC_604/A OR2X1_LOC_7/A 1.96fF
C53034 OR2X1_LOC_7/A OR2X1_LOC_183/a_8_216# 0.21fF
C53284 AND2X1_LOC_155/Y OR2X1_LOC_7/A 0.01fF
C53290 OR2X1_LOC_230/a_8_216# OR2X1_LOC_7/A 0.05fF
C53504 AND2X1_LOC_539/Y OR2X1_LOC_7/A 0.03fF
C54054 OR2X1_LOC_298/Y OR2X1_LOC_7/A 0.05fF
C54114 OR2X1_LOC_7/A OR2X1_LOC_27/a_8_216# 0.01fF
C54426 OR2X1_LOC_7/A AND2X1_LOC_434/Y 0.79fF
C55377 AND2X1_LOC_342/a_8_24# OR2X1_LOC_7/A 0.04fF
C55630 OR2X1_LOC_7/A OR2X1_LOC_766/Y 0.01fF
C55982 OR2X1_LOC_7/A OR2X1_LOC_248/A 0.03fF
C55995 OR2X1_LOC_7/A OR2X1_LOC_504/a_36_216# 0.02fF
C56939 OR2X1_LOC_7/A VSS -29.87fF
C34125 OR2X1_LOC_97/A AND2X1_LOC_19/Y 0.02fF
C36299 AND2X1_LOC_19/Y AND2X1_LOC_20/a_8_24# 0.11fF
C36770 OR2X1_LOC_520/Y AND2X1_LOC_19/Y 1.24fF
C41380 VDD AND2X1_LOC_19/Y 0.31fF
C44511 OR2X1_LOC_160/A AND2X1_LOC_19/Y 0.01fF
C45807 OR2X1_LOC_185/A AND2X1_LOC_19/Y 0.03fF
C54226 AND2X1_LOC_19/Y AND2X1_LOC_44/Y 0.01fF
C56101 AND2X1_LOC_19/Y OR2X1_LOC_130/A 0.04fF
C57532 AND2X1_LOC_19/Y VSS 0.25fF
C3734 AND2X1_LOC_765/a_8_24# OR2X1_LOC_557/A 0.19fF
C4682 OR2X1_LOC_557/A OR2X1_LOC_375/A 0.03fF
C5535 OR2X1_LOC_391/B OR2X1_LOC_557/A 0.01fF
C9042 OR2X1_LOC_557/A AND2X1_LOC_815/a_8_24# 0.06fF
C15017 AND2X1_LOC_79/a_8_24# OR2X1_LOC_557/A 0.01fF
C15200 OR2X1_LOC_557/A OR2X1_LOC_113/B 0.01fF
C17361 VDD OR2X1_LOC_557/A 0.53fF
C20098 OR2X1_LOC_557/A OR2X1_LOC_846/B 0.09fF
C21267 OR2X1_LOC_557/A OR2X1_LOC_78/Y 0.03fF
C24133 AND2X1_LOC_91/B OR2X1_LOC_557/A 0.10fF
C28099 AND2X1_LOC_393/a_8_24# OR2X1_LOC_557/A 0.01fF
C29096 OR2X1_LOC_557/A OR2X1_LOC_771/B 0.03fF
C33599 OR2X1_LOC_400/B OR2X1_LOC_557/A 0.01fF
C34033 OR2X1_LOC_557/A AND2X1_LOC_51/Y 1.94fF
C37109 OR2X1_LOC_557/A AND2X1_LOC_36/Y 0.02fF
C44148 AND2X1_LOC_103/a_8_24# OR2X1_LOC_557/A 0.01fF
C45130 OR2X1_LOC_287/B OR2X1_LOC_557/A 2.24fF
C51239 OR2X1_LOC_557/A OR2X1_LOC_84/A -0.00fF
C57198 OR2X1_LOC_557/A VSS -1.01fF
C540 OR2X1_LOC_744/A OR2X1_LOC_589/a_8_216# 0.01fF
C979 OR2X1_LOC_744/A AND2X1_LOC_793/B 0.60fF
C986 OR2X1_LOC_744/A OR2X1_LOC_533/A 0.01fF
C1683 OR2X1_LOC_131/Y OR2X1_LOC_744/A 0.49fF
C1960 VDD OR2X1_LOC_744/A 1.19fF
C2004 OR2X1_LOC_744/A OR2X1_LOC_677/Y 0.03fF
C2078 OR2X1_LOC_744/A OR2X1_LOC_491/Y 0.01fF
C2232 OR2X1_LOC_744/A OR2X1_LOC_67/Y 0.03fF
C2522 OR2X1_LOC_744/A AND2X1_LOC_834/a_8_24# 0.02fF
C2536 OR2X1_LOC_744/A OR2X1_LOC_248/Y 0.19fF
C4204 AND2X1_LOC_557/a_8_24# OR2X1_LOC_744/A 0.02fF
C4846 OR2X1_LOC_45/B OR2X1_LOC_744/A 1.58fF
C4953 OR2X1_LOC_744/A AND2X1_LOC_435/a_8_24# 0.01fF
C5269 OR2X1_LOC_158/A OR2X1_LOC_744/A 1.01fF
C5321 OR2X1_LOC_744/A OR2X1_LOC_103/Y 0.03fF
C5327 OR2X1_LOC_744/A OR2X1_LOC_594/Y 0.10fF
C5700 OR2X1_LOC_482/Y OR2X1_LOC_744/A 0.10fF
C5736 OR2X1_LOC_744/A OR2X1_LOC_816/Y 0.14fF
C7469 AND2X1_LOC_541/Y OR2X1_LOC_744/A 0.15fF
C7571 OR2X1_LOC_744/A OR2X1_LOC_316/Y 0.03fF
C7621 AND2X1_LOC_390/B OR2X1_LOC_744/A 0.07fF
C7897 OR2X1_LOC_309/Y OR2X1_LOC_744/A 0.03fF
C8032 OR2X1_LOC_744/A AND2X1_LOC_840/B 0.05fF
C8759 OR2X1_LOC_744/A OR2X1_LOC_522/Y 0.07fF
C8822 OR2X1_LOC_179/a_8_216# OR2X1_LOC_744/A 0.02fF
C9163 OR2X1_LOC_118/a_8_216# OR2X1_LOC_744/A 0.01fF
C9250 OR2X1_LOC_744/A AND2X1_LOC_638/Y 0.36fF
C9746 OR2X1_LOC_91/Y OR2X1_LOC_744/A 0.07fF
C9812 OR2X1_LOC_417/Y OR2X1_LOC_744/A 0.03fF
C9985 OR2X1_LOC_744/A AND2X1_LOC_780/a_8_24# 0.02fF
C10184 OR2X1_LOC_744/A OR2X1_LOC_83/A 0.27fF
C10562 OR2X1_LOC_744/A AND2X1_LOC_436/B 0.10fF
C10897 OR2X1_LOC_744/A OR2X1_LOC_484/a_8_216# 0.01fF
C11277 OR2X1_LOC_492/Y OR2X1_LOC_744/A 0.04fF
C11285 OR2X1_LOC_108/a_8_216# OR2X1_LOC_744/A 0.03fF
C11543 OR2X1_LOC_744/A OR2X1_LOC_409/B 0.83fF
C11673 OR2X1_LOC_146/a_8_216# OR2X1_LOC_744/A 0.18fF
C11811 OR2X1_LOC_525/Y OR2X1_LOC_744/A 0.19fF
C11853 OR2X1_LOC_744/A OR2X1_LOC_497/Y 0.07fF
C12110 OR2X1_LOC_744/A AND2X1_LOC_249/a_8_24# 0.01fF
C12163 OR2X1_LOC_744/A OR2X1_LOC_380/a_8_216# 0.05fF
C12696 OR2X1_LOC_744/A AND2X1_LOC_319/A 0.03fF
C12847 OR2X1_LOC_744/A AND2X1_LOC_721/A 0.03fF
C12892 OR2X1_LOC_744/A OR2X1_LOC_331/Y 0.03fF
C13149 OR2X1_LOC_744/A AND2X1_LOC_318/a_8_24# 0.06fF
C13174 OR2X1_LOC_744/A AND2X1_LOC_361/A 0.07fF
C13583 OR2X1_LOC_83/Y OR2X1_LOC_744/A 0.01fF
C13960 AND2X1_LOC_532/a_8_24# OR2X1_LOC_744/A 0.01fF
C14686 OR2X1_LOC_692/Y OR2X1_LOC_744/A 0.01fF
C14716 OR2X1_LOC_744/A OR2X1_LOC_600/A 6.00fF
C14786 OR2X1_LOC_744/A OR2X1_LOC_619/Y 0.13fF
C15088 OR2X1_LOC_744/A AND2X1_LOC_769/Y 0.01fF
C15461 OR2X1_LOC_744/A AND2X1_LOC_783/B 0.01fF
C16969 OR2X1_LOC_744/A OR2X1_LOC_312/Y 0.06fF
C17148 OR2X1_LOC_744/A OR2X1_LOC_13/B 0.17fF
C17294 OR2X1_LOC_744/A AND2X1_LOC_266/a_8_24# 0.01fF
C17549 OR2X1_LOC_744/A OR2X1_LOC_142/a_8_216# 0.01fF
C17608 OR2X1_LOC_744/A OR2X1_LOC_595/A 0.08fF
C18201 OR2X1_LOC_744/A AND2X1_LOC_342/Y 0.39fF
C18690 OR2X1_LOC_744/A OR2X1_LOC_89/A 0.13fF
C19375 OR2X1_LOC_491/a_8_216# OR2X1_LOC_744/A 0.02fF
C19593 OR2X1_LOC_744/A AND2X1_LOC_727/A 0.03fF
C19630 OR2X1_LOC_744/A OR2X1_LOC_95/Y 0.40fF
C19859 OR2X1_LOC_122/Y OR2X1_LOC_744/A 0.06fF
C19880 OR2X1_LOC_179/Y OR2X1_LOC_744/A 0.01fF
C19900 OR2X1_LOC_744/A AND2X1_LOC_832/a_8_24# 0.02fF
C20229 OR2X1_LOC_693/Y OR2X1_LOC_744/A 0.01fF
C20843 OR2X1_LOC_70/Y OR2X1_LOC_744/A 0.34fF
C20947 OR2X1_LOC_744/A OR2X1_LOC_184/Y 0.07fF
C21959 AND2X1_LOC_535/Y OR2X1_LOC_744/A 0.03fF
C21992 OR2X1_LOC_744/A OR2X1_LOC_484/Y 0.10fF
C22373 OR2X1_LOC_744/A OR2X1_LOC_16/A 0.89fF
C22392 OR2X1_LOC_108/Y OR2X1_LOC_744/A 1.15fF
C22622 OR2X1_LOC_744/A AND2X1_LOC_687/Y 0.02fF
C23329 OR2X1_LOC_109/Y OR2X1_LOC_744/A 0.03fF
C23844 OR2X1_LOC_744/A AND2X1_LOC_798/Y 0.23fF
C23898 OR2X1_LOC_744/A AND2X1_LOC_227/Y 0.09fF
C24214 OR2X1_LOC_599/A OR2X1_LOC_744/A 0.82fF
C24478 OR2X1_LOC_40/Y OR2X1_LOC_744/A 0.28fF
C24551 OR2X1_LOC_744/A AND2X1_LOC_843/Y 0.11fF
C24737 OR2X1_LOC_744/A OR2X1_LOC_224/a_8_216# 0.02fF
C25151 OR2X1_LOC_744/A OR2X1_LOC_615/Y 0.07fF
C25385 OR2X1_LOC_744/A AND2X1_LOC_841/B 8.65fF
C25712 AND2X1_LOC_706/a_8_24# OR2X1_LOC_744/A 0.01fF
C25824 OR2X1_LOC_744/A AND2X1_LOC_379/a_8_24# 0.01fF
C26725 OR2X1_LOC_3/Y OR2X1_LOC_744/A 0.67fF
C27115 OR2X1_LOC_744/A AND2X1_LOC_113/Y 0.01fF
C28039 OR2X1_LOC_744/A OR2X1_LOC_64/Y 0.37fF
C29155 OR2X1_LOC_516/B OR2X1_LOC_744/A 0.02fF
C29574 AND2X1_LOC_456/B OR2X1_LOC_744/A 0.03fF
C29929 OR2X1_LOC_744/A AND2X1_LOC_828/a_8_24# 0.01fF
C30761 OR2X1_LOC_744/A AND2X1_LOC_802/Y 0.16fF
C31240 OR2X1_LOC_744/A AND2X1_LOC_325/a_8_24# 0.06fF
C31339 OR2X1_LOC_744/A OR2X1_LOC_380/A 0.15fF
C32170 OR2X1_LOC_763/Y OR2X1_LOC_744/A 0.09fF
C32266 OR2X1_LOC_744/A AND2X1_LOC_114/Y 0.12fF
C32583 OR2X1_LOC_744/A AND2X1_LOC_114/a_8_24# 0.02fF
C33729 OR2X1_LOC_744/A OR2X1_LOC_744/a_8_216# 0.20fF
C34080 OR2X1_LOC_744/A OR2X1_LOC_142/Y 0.07fF
C34245 OR2X1_LOC_744/A OR2X1_LOC_118/Y 0.03fF
C34756 OR2X1_LOC_744/A OR2X1_LOC_83/a_8_216# 0.01fF
C34848 OR2X1_LOC_744/A OR2X1_LOC_503/Y 0.10fF
C35409 OR2X1_LOC_604/A OR2X1_LOC_744/A 0.18fF
C35828 OR2X1_LOC_176/Y OR2X1_LOC_744/A 0.50fF
C36187 OR2X1_LOC_744/A OR2X1_LOC_183/a_8_216# 0.02fF
C36418 OR2X1_LOC_744/A AND2X1_LOC_155/Y 0.09fF
C36468 OR2X1_LOC_744/A AND2X1_LOC_633/Y 0.01fF
C36619 AND2X1_LOC_539/Y OR2X1_LOC_744/A 0.16fF
C36654 OR2X1_LOC_131/A OR2X1_LOC_744/A 0.03fF
C37551 OR2X1_LOC_744/A AND2X1_LOC_434/Y 0.07fF
C37672 OR2X1_LOC_764/Y OR2X1_LOC_744/A 0.01fF
C38517 AND2X1_LOC_355/a_8_24# OR2X1_LOC_744/A 0.03fF
C38916 OR2X1_LOC_744/A OR2X1_LOC_393/Y 0.09fF
C39307 OR2X1_LOC_744/A OR2X1_LOC_594/a_8_216# 0.01fF
C39810 OR2X1_LOC_744/A OR2X1_LOC_283/Y 1.46fF
C40101 AND2X1_LOC_160/a_8_24# OR2X1_LOC_744/A 0.09fF
C40523 OR2X1_LOC_597/A OR2X1_LOC_744/A 0.03fF
C40533 OR2X1_LOC_178/Y OR2X1_LOC_744/A 0.03fF
C40898 OR2X1_LOC_744/A OR2X1_LOC_829/A 0.03fF
C41188 OR2X1_LOC_744/A OR2X1_LOC_224/Y 0.02fF
C41773 OR2X1_LOC_744/A OR2X1_LOC_764/a_8_216# 0.01fF
C41797 OR2X1_LOC_744/A AND2X1_LOC_810/B 0.24fF
C43107 OR2X1_LOC_744/A OR2X1_LOC_323/Y 0.43fF
C43227 AND2X1_LOC_729/Y OR2X1_LOC_744/A 0.10fF
C43254 AND2X1_LOC_784/A OR2X1_LOC_744/A 0.07fF
C43279 AND2X1_LOC_769/a_8_24# OR2X1_LOC_744/A 0.01fF
C43711 OR2X1_LOC_744/A OR2X1_LOC_52/B 0.13fF
C43728 AND2X1_LOC_489/Y OR2X1_LOC_744/A 0.09fF
C43851 OR2X1_LOC_744/A AND2X1_LOC_216/A 0.02fF
C44081 OR2X1_LOC_744/A OR2X1_LOC_394/Y 0.01fF
C44139 AND2X1_LOC_356/B OR2X1_LOC_744/A 0.03fF
C44144 OR2X1_LOC_280/Y OR2X1_LOC_744/A 0.46fF
C44412 OR2X1_LOC_485/Y OR2X1_LOC_744/A 0.27fF
C44817 OR2X1_LOC_744/A OR2X1_LOC_744/Y 0.01fF
C44940 OR2X1_LOC_744/A AND2X1_LOC_593/Y 0.53fF
C45310 OR2X1_LOC_744/A OR2X1_LOC_51/Y 0.41fF
C45403 OR2X1_LOC_744/A OR2X1_LOC_680/A 0.07fF
C45921 OR2X1_LOC_744/A AND2X1_LOC_802/a_8_24# 0.01fF
C46181 OR2X1_LOC_178/a_8_216# OR2X1_LOC_744/A -0.01fF
C46191 OR2X1_LOC_744/A AND2X1_LOC_436/Y 0.04fF
C46312 OR2X1_LOC_744/A OR2X1_LOC_588/Y 0.68fF
C47216 OR2X1_LOC_744/A AND2X1_LOC_266/Y 0.01fF
C47463 OR2X1_LOC_744/A OR2X1_LOC_183/Y 0.02fF
C47654 OR2X1_LOC_744/A OR2X1_LOC_511/Y 0.05fF
C47923 AND2X1_LOC_799/a_8_24# OR2X1_LOC_744/A 0.01fF
C48400 OR2X1_LOC_744/A OR2X1_LOC_131/a_8_216# 0.01fF
C48447 AND2X1_LOC_391/Y OR2X1_LOC_744/A 0.04fF
C49108 OR2X1_LOC_744/A OR2X1_LOC_423/Y 0.15fF
C49355 OR2X1_LOC_744/A AND2X1_LOC_114/a_36_24# 0.01fF
C49392 OR2X1_LOC_744/A OR2X1_LOC_74/A 0.10fF
C49741 OR2X1_LOC_744/A OR2X1_LOC_432/a_8_216# 0.01fF
C50166 OR2X1_LOC_744/A OR2X1_LOC_432/Y 0.01fF
C50558 OR2X1_LOC_744/A OR2X1_LOC_594/a_36_216# -0.00fF
C51022 OR2X1_LOC_744/A AND2X1_LOC_633/a_8_24# 0.01fF
C51271 OR2X1_LOC_106/Y OR2X1_LOC_744/A 0.08fF
C51439 OR2X1_LOC_744/A OR2X1_LOC_497/a_8_216# 0.04fF
C51846 OR2X1_LOC_744/A AND2X1_LOC_99/A 0.03fF
C51893 OR2X1_LOC_744/A AND2X1_LOC_637/Y 0.02fF
C52594 AND2X1_LOC_362/B OR2X1_LOC_744/A 1.49fF
C53010 AND2X1_LOC_706/Y OR2X1_LOC_744/A 0.01fF
C53404 AND2X1_LOC_802/B OR2X1_LOC_744/A 0.05fF
C54594 OR2X1_LOC_744/A OR2X1_LOC_589/Y 0.01fF
C55047 OR2X1_LOC_744/A OR2X1_LOC_743/Y 0.01fF
C55552 OR2X1_LOC_526/Y OR2X1_LOC_744/A 0.14fF
C55641 OR2X1_LOC_744/A OR2X1_LOC_433/Y 0.01fF
C57580 OR2X1_LOC_744/A VSS 1.31fF
C896 OR2X1_LOC_600/A AND2X1_LOC_837/a_8_24# 0.01fF
C2015 OR2X1_LOC_600/A AND2X1_LOC_847/Y 0.01fF
C2465 AND2X1_LOC_99/A OR2X1_LOC_600/A 0.03fF
C3223 AND2X1_LOC_362/B OR2X1_LOC_600/A 0.07fF
C3651 OR2X1_LOC_58/Y OR2X1_LOC_600/A 0.03fF
C3778 OR2X1_LOC_665/Y OR2X1_LOC_600/A 0.09fF
C4139 OR2X1_LOC_495/a_8_216# OR2X1_LOC_600/A 0.06fF
C4147 OR2X1_LOC_600/A AND2X1_LOC_838/a_8_24# 0.01fF
C4341 OR2X1_LOC_600/A OR2X1_LOC_385/a_8_216# 0.14fF
C4460 OR2X1_LOC_122/a_8_216# OR2X1_LOC_600/A 0.05fF
C5300 OR2X1_LOC_290/a_8_216# OR2X1_LOC_600/A 0.05fF
C5441 OR2X1_LOC_665/a_8_216# OR2X1_LOC_600/A 0.01fF
C5684 OR2X1_LOC_600/A OR2X1_LOC_13/Y 0.03fF
C5917 OR2X1_LOC_600/A OR2X1_LOC_295/Y 0.01fF
C7383 OR2X1_LOC_516/Y OR2X1_LOC_600/A 0.11fF
C7756 OR2X1_LOC_600/A OR2X1_LOC_533/A 0.16fF
C8186 OR2X1_LOC_600/A AND2X1_LOC_846/a_8_24# 0.01fF
C8354 OR2X1_LOC_125/a_8_216# OR2X1_LOC_600/A 0.07fF
C8770 VDD OR2X1_LOC_600/A 1.35fF
C8845 OR2X1_LOC_600/A OR2X1_LOC_616/Y 0.83fF
C8886 OR2X1_LOC_251/Y OR2X1_LOC_600/A 0.30fF
C8928 OR2X1_LOC_826/a_8_216# OR2X1_LOC_600/A 0.01fF
C10632 OR2X1_LOC_600/A OR2X1_LOC_416/Y 0.03fF
C10995 AND2X1_LOC_557/a_8_24# OR2X1_LOC_600/A 0.04fF
C11674 OR2X1_LOC_45/B OR2X1_LOC_600/A 0.20fF
C11948 OR2X1_LOC_600/A AND2X1_LOC_838/B 0.02fF
C12106 OR2X1_LOC_158/A OR2X1_LOC_600/A 3.65fF
C12167 OR2X1_LOC_600/A AND2X1_LOC_98/Y 0.22fF
C12181 OR2X1_LOC_600/A OR2X1_LOC_103/Y 0.03fF
C12184 OR2X1_LOC_600/A OR2X1_LOC_594/Y 0.07fF
C12618 OR2X1_LOC_600/A OR2X1_LOC_586/Y 0.05fF
C12683 OR2X1_LOC_748/A OR2X1_LOC_600/A 0.06fF
C13218 OR2X1_LOC_600/A OR2X1_LOC_815/A 0.03fF
C13714 OR2X1_LOC_600/A AND2X1_LOC_848/A 0.18fF
C14261 AND2X1_LOC_541/Y OR2X1_LOC_600/A 0.04fF
C14371 OR2X1_LOC_600/A OR2X1_LOC_316/Y 0.03fF
C14438 OR2X1_LOC_825/a_8_216# OR2X1_LOC_600/A 0.01fF
C14787 OR2X1_LOC_600/A AND2X1_LOC_840/B 0.05fF
C14960 OR2X1_LOC_600/A OR2X1_LOC_257/Y 0.01fF
C15077 OR2X1_LOC_600/A AND2X1_LOC_464/A 0.03fF
C15546 OR2X1_LOC_179/a_8_216# OR2X1_LOC_600/A 0.01fF
C15713 OR2X1_LOC_600/A OR2X1_LOC_751/A 0.01fF
C16447 OR2X1_LOC_91/Y OR2X1_LOC_600/A 0.12fF
C16530 OR2X1_LOC_417/Y OR2X1_LOC_600/A 0.04fF
C16730 OR2X1_LOC_600/A OR2X1_LOC_171/Y 2.75fF
C17977 OR2X1_LOC_600/A AND2X1_LOC_789/Y 0.15fF
C18065 OR2X1_LOC_108/a_8_216# OR2X1_LOC_600/A 0.01fF
C18270 OR2X1_LOC_600/A OR2X1_LOC_125/Y 0.03fF
C19398 OR2X1_LOC_235/B OR2X1_LOC_600/A 0.07fF
C19640 OR2X1_LOC_600/A AND2X1_LOC_721/A 0.03fF
C19671 OR2X1_LOC_600/A OR2X1_LOC_331/Y 0.07fF
C20613 AND2X1_LOC_787/A OR2X1_LOC_600/A 0.05fF
C20697 AND2X1_LOC_391/a_8_24# OR2X1_LOC_600/A 0.03fF
C20731 OR2X1_LOC_127/a_8_216# OR2X1_LOC_600/A 0.02fF
C21165 OR2X1_LOC_600/A OR2X1_LOC_257/a_8_216# 0.01fF
C23780 OR2X1_LOC_312/Y OR2X1_LOC_600/A 0.03fF
C23971 OR2X1_LOC_600/A OR2X1_LOC_13/B 0.13fF
C24447 OR2X1_LOC_600/A OR2X1_LOC_595/A 0.07fF
C24886 OR2X1_LOC_528/Y OR2X1_LOC_600/A 0.03fF
C25001 OR2X1_LOC_600/A AND2X1_LOC_105/a_8_24# 0.01fF
C25431 OR2X1_LOC_600/A OR2X1_LOC_89/A 0.10fF
C26181 OR2X1_LOC_600/A OR2X1_LOC_251/a_8_216# 0.02fF
C26207 OR2X1_LOC_45/Y OR2X1_LOC_600/A 0.43fF
C26308 OR2X1_LOC_600/A AND2X1_LOC_727/A 0.03fF
C26343 OR2X1_LOC_600/A OR2X1_LOC_95/Y 0.88fF
C26586 OR2X1_LOC_179/Y OR2X1_LOC_600/A 0.01fF
C27073 OR2X1_LOC_600/A AND2X1_LOC_621/Y 0.03fF
C27307 OR2X1_LOC_600/A OR2X1_LOC_71/A 0.07fF
C27548 OR2X1_LOC_70/Y OR2X1_LOC_600/A 0.10fF
C27555 AND2X1_LOC_557/a_36_24# OR2X1_LOC_600/A 0.01fF
C29051 OR2X1_LOC_600/A OR2X1_LOC_16/A 11.19fF
C29082 OR2X1_LOC_108/Y OR2X1_LOC_600/A 0.24fF
C29159 AND2X1_LOC_168/Y OR2X1_LOC_600/A 0.50fF
C29940 OR2X1_LOC_600/A AND2X1_LOC_447/Y 0.01fF
C30017 OR2X1_LOC_109/Y OR2X1_LOC_600/A 0.07fF
C30106 OR2X1_LOC_600/A AND2X1_LOC_729/B 0.03fF
C30479 OR2X1_LOC_600/A OR2X1_LOC_106/A 0.04fF
C30569 OR2X1_LOC_600/A AND2X1_LOC_227/Y 0.03fF
C30620 OR2X1_LOC_600/A OR2X1_LOC_41/Y 0.46fF
C30867 OR2X1_LOC_600/A OR2X1_LOC_250/a_8_216# 0.01fF
C30939 OR2X1_LOC_600/A OR2X1_LOC_258/a_8_216# 0.01fF
C31205 OR2X1_LOC_40/Y OR2X1_LOC_600/A 0.32fF
C31428 OR2X1_LOC_600/A OR2X1_LOC_224/a_8_216# 0.01fF
C31672 OR2X1_LOC_600/A OR2X1_LOC_251/a_36_216# 0.02fF
C31710 OR2X1_LOC_127/Y OR2X1_LOC_600/A 0.01fF
C32372 AND2X1_LOC_543/Y OR2X1_LOC_600/A 0.01fF
C32444 OR2X1_LOC_600/A OR2X1_LOC_261/a_8_216# 0.03fF
C32628 OR2X1_LOC_600/A OR2X1_LOC_60/a_8_216# 0.05fF
C32646 OR2X1_LOC_600/A AND2X1_LOC_664/a_8_24# 0.01fF
C33470 OR2X1_LOC_3/Y OR2X1_LOC_600/A 0.35fF
C34747 OR2X1_LOC_600/A OR2X1_LOC_64/Y 0.07fF
C34930 OR2X1_LOC_600/A AND2X1_LOC_247/a_8_24# 0.03fF
C36416 OR2X1_LOC_825/Y OR2X1_LOC_600/A 0.21fF
C37745 OR2X1_LOC_600/A OR2X1_LOC_751/a_8_216# 0.01fF
C37930 AND2X1_LOC_709/a_8_24# OR2X1_LOC_600/A 0.01fF
C38006 OR2X1_LOC_600/A AND2X1_LOC_624/A 0.32fF
C39327 OR2X1_LOC_600/A AND2X1_LOC_114/a_8_24# 0.05fF
C39837 OR2X1_LOC_600/A OR2X1_LOC_295/a_8_216# 0.01fF
C40545 OR2X1_LOC_751/Y OR2X1_LOC_600/A 0.23fF
C40822 OR2X1_LOC_600/A OR2X1_LOC_142/Y 0.03fF
C41059 OR2X1_LOC_600/A OR2X1_LOC_238/Y 0.03fF
C41470 OR2X1_LOC_516/a_8_216# OR2X1_LOC_600/A 0.01fF
C41889 OR2X1_LOC_600/A OR2X1_LOC_250/Y 0.14fF
C42209 OR2X1_LOC_177/Y OR2X1_LOC_600/A 0.03fF
C42226 OR2X1_LOC_604/A OR2X1_LOC_600/A 0.23fF
C42228 AND2X1_LOC_758/a_8_24# OR2X1_LOC_600/A 0.01fF
C42668 OR2X1_LOC_533/Y OR2X1_LOC_600/A 0.06fF
C42780 OR2X1_LOC_600/A OR2X1_LOC_265/Y 0.39fF
C43548 AND2X1_LOC_711/A OR2X1_LOC_600/A 0.03fF
C43956 AND2X1_LOC_338/A OR2X1_LOC_600/A 0.08fF
C44416 OR2X1_LOC_600/A AND2X1_LOC_434/Y 0.15fF
C45786 OR2X1_LOC_600/A OR2X1_LOC_393/Y 0.03fF
C46210 AND2X1_LOC_789/a_8_24# OR2X1_LOC_600/A 0.01fF
C46612 OR2X1_LOC_815/a_8_216# OR2X1_LOC_600/A 0.01fF
C46710 OR2X1_LOC_600/A AND2X1_LOC_848/Y 0.03fF
C46792 OR2X1_LOC_600/A OR2X1_LOC_617/Y 0.03fF
C47096 AND2X1_LOC_756/a_8_24# OR2X1_LOC_600/A 0.15fF
C47547 OR2X1_LOC_178/Y OR2X1_LOC_600/A 0.03fF
C47680 OR2X1_LOC_600/A OR2X1_LOC_258/Y 0.01fF
C47798 OR2X1_LOC_600/A OR2X1_LOC_815/Y 0.01fF
C47955 OR2X1_LOC_759/A OR2X1_LOC_600/A 0.18fF
C48058 OR2X1_LOC_600/A AND2X1_LOC_838/Y 0.79fF
C48214 OR2X1_LOC_600/A OR2X1_LOC_224/Y 0.01fF
C48834 OR2X1_LOC_600/A OR2X1_LOC_165/Y 0.03fF
C49159 OR2X1_LOC_600/A OR2X1_LOC_230/Y 0.14fF
C49207 AND2X1_LOC_709/a_36_24# OR2X1_LOC_600/A -0.00fF
C50154 AND2X1_LOC_729/Y OR2X1_LOC_600/A 0.09fF
C50181 AND2X1_LOC_784/A OR2X1_LOC_600/A 0.07fF
C50386 OR2X1_LOC_600/A OR2X1_LOC_172/Y 0.07fF
C50612 OR2X1_LOC_600/A OR2X1_LOC_52/B 0.13fF
C50628 AND2X1_LOC_489/Y OR2X1_LOC_600/A 0.03fF
C50668 OR2X1_LOC_755/A OR2X1_LOC_600/A 0.99fF
C51036 OR2X1_LOC_280/Y OR2X1_LOC_600/A 0.10fF
C51554 OR2X1_LOC_600/A OR2X1_LOC_826/Y 0.02fF
C51826 OR2X1_LOC_600/A AND2X1_LOC_593/Y 3.04fF
C52159 OR2X1_LOC_600/A OR2X1_LOC_51/Y 0.41fF
C52253 OR2X1_LOC_680/A OR2X1_LOC_600/A 0.06fF
C52606 OR2X1_LOC_757/A OR2X1_LOC_600/A 0.05fF
C53017 OR2X1_LOC_178/a_8_216# OR2X1_LOC_600/A 0.01fF
C53026 OR2X1_LOC_600/A AND2X1_LOC_436/Y 0.03fF
C54178 OR2X1_LOC_600/A OR2X1_LOC_183/Y 0.04fF
C54772 OR2X1_LOC_600/A OR2X1_LOC_237/Y 0.03fF
C55117 AND2X1_LOC_391/Y OR2X1_LOC_600/A 1.32fF
C56134 OR2X1_LOC_600/A OR2X1_LOC_74/A 0.19fF
C56167 OR2X1_LOC_600/A OR2X1_LOC_261/A 0.18fF
C57436 OR2X1_LOC_600/A VSS 1.12fF
C8291 AND2X1_LOC_101/B AND2X1_LOC_216/A 0.46fF
C22519 VDD AND2X1_LOC_101/B 0.01fF
C22772 AND2X1_LOC_101/B OR2X1_LOC_67/Y 0.01fF
C28132 AND2X1_LOC_101/B AND2X1_LOC_101/a_8_24# 0.01fF
C37507 AND2X1_LOC_101/B OR2X1_LOC_13/B 0.10fF
C41200 OR2X1_LOC_70/Y AND2X1_LOC_101/B 0.01fF
C44340 AND2X1_LOC_101/B OR2X1_LOC_813/Y 0.09fF
C47370 OR2X1_LOC_3/Y AND2X1_LOC_101/B 0.08fF
C48663 AND2X1_LOC_101/B OR2X1_LOC_64/Y 0.25fF
C57449 AND2X1_LOC_101/B VSS 0.30fF
C3155 OR2X1_LOC_473/A OR2X1_LOC_810/A 0.29fF
C5113 OR2X1_LOC_473/A OR2X1_LOC_78/A 0.10fF
C6320 OR2X1_LOC_121/Y OR2X1_LOC_473/A 0.03fF
C7685 OR2X1_LOC_140/A OR2X1_LOC_473/A 0.37fF
C9955 OR2X1_LOC_574/A OR2X1_LOC_473/A 0.15fF
C10775 OR2X1_LOC_473/A OR2X1_LOC_375/A 0.02fF
C11072 OR2X1_LOC_473/A OR2X1_LOC_549/A 0.03fF
C15636 OR2X1_LOC_473/A OR2X1_LOC_130/a_8_216# 0.18fF
C18312 OR2X1_LOC_473/A OR2X1_LOC_361/a_8_216# 0.03fF
C18703 OR2X1_LOC_473/A OR2X1_LOC_267/Y 0.04fF
C21505 OR2X1_LOC_473/A OR2X1_LOC_532/B 0.72fF
C23475 VDD OR2X1_LOC_473/A 0.07fF
C25459 OR2X1_LOC_473/A OR2X1_LOC_115/B 0.09fF
C25988 OR2X1_LOC_216/A OR2X1_LOC_473/A 0.05fF
C26441 OR2X1_LOC_160/A OR2X1_LOC_473/A 0.74fF
C32307 OR2X1_LOC_473/A OR2X1_LOC_506/A 0.02fF
C37825 OR2X1_LOC_473/A OR2X1_LOC_130/A 0.29fF
C39999 OR2X1_LOC_473/A AND2X1_LOC_51/Y 0.43fF
C46932 OR2X1_LOC_473/A OR2X1_LOC_493/A 0.19fF
C47887 OR2X1_LOC_473/A AND2X1_LOC_67/Y 0.31fF
C52388 OR2X1_LOC_151/A OR2X1_LOC_473/A 0.15fF
C53693 OR2X1_LOC_473/A OR2X1_LOC_631/A 0.83fF
C57202 OR2X1_LOC_473/A VSS 0.45fF
C7362 OR2X1_LOC_623/B OR2X1_LOC_513/Y 0.13fF
C10810 OR2X1_LOC_375/A OR2X1_LOC_513/Y 0.01fF
C11022 OR2X1_LOC_513/Y OR2X1_LOC_515/Y 0.15fF
C16636 OR2X1_LOC_513/Y OR2X1_LOC_713/A 0.01fF
C17567 OR2X1_LOC_154/A OR2X1_LOC_513/Y 0.01fF
C23539 VDD OR2X1_LOC_513/Y 0.18fF
C24354 OR2X1_LOC_676/Y OR2X1_LOC_513/Y 0.01fF
C24363 OR2X1_LOC_834/A OR2X1_LOC_513/Y 0.09fF
C35284 OR2X1_LOC_678/a_8_216# OR2X1_LOC_513/Y 0.40fF
C36094 AND2X1_LOC_44/Y OR2X1_LOC_513/Y 0.01fF
C43311 AND2X1_LOC_36/Y OR2X1_LOC_513/Y 0.01fF
C46519 OR2X1_LOC_678/Y OR2X1_LOC_513/Y 0.01fF
C56360 OR2X1_LOC_513/Y VSS 0.25fF
C1635 OR2X1_LOC_809/B OR2X1_LOC_802/Y 0.10fF
C7681 OR2X1_LOC_809/B AND2X1_LOC_47/Y 0.05fF
C13003 OR2X1_LOC_112/a_8_216# OR2X1_LOC_809/B 0.03fF
C17947 OR2X1_LOC_809/B AND2X1_LOC_31/Y 0.07fF
C18221 OR2X1_LOC_809/B OR2X1_LOC_809/a_8_216# 0.02fF
C21638 OR2X1_LOC_809/B OR2X1_LOC_539/Y 0.01fF
C27823 OR2X1_LOC_151/A OR2X1_LOC_809/B 0.06fF
C34119 OR2X1_LOC_138/a_8_216# OR2X1_LOC_809/B 0.40fF
C34716 OR2X1_LOC_809/B OR2X1_LOC_810/A 0.03fF
C35017 OR2X1_LOC_715/B OR2X1_LOC_809/B 0.15fF
C37970 OR2X1_LOC_809/B OR2X1_LOC_538/A 0.03fF
C40882 OR2X1_LOC_186/Y OR2X1_LOC_809/B 0.11fF
C41186 OR2X1_LOC_809/B OR2X1_LOC_112/B 0.19fF
C45688 OR2X1_LOC_809/B OR2X1_LOC_138/A 0.09fF
C53235 OR2X1_LOC_809/B OR2X1_LOC_532/B 0.24fF
C55113 VDD OR2X1_LOC_809/B 0.07fF
C57676 OR2X1_LOC_809/B VSS 0.41fF
C796 AND2X1_LOC_666/a_8_24# AND2X1_LOC_18/Y 0.03fF
C1145 OR2X1_LOC_668/a_8_216# AND2X1_LOC_18/Y 0.02fF
C1631 OR2X1_LOC_403/B AND2X1_LOC_18/Y 0.01fF
C1991 OR2X1_LOC_61/B AND2X1_LOC_18/Y 0.03fF
C2011 OR2X1_LOC_194/B AND2X1_LOC_18/Y 0.10fF
C2338 OR2X1_LOC_97/A AND2X1_LOC_18/Y 0.04fF
C2417 OR2X1_LOC_541/A AND2X1_LOC_18/Y 0.05fF
C3317 OR2X1_LOC_559/B AND2X1_LOC_18/Y 0.01fF
C3337 OR2X1_LOC_720/A AND2X1_LOC_18/Y 0.02fF
C3382 OR2X1_LOC_333/B AND2X1_LOC_18/Y 0.03fF
C3741 OR2X1_LOC_154/A AND2X1_LOC_18/Y 3.07fF
C3759 OR2X1_LOC_267/A AND2X1_LOC_18/Y 0.13fF
C4264 AND2X1_LOC_813/a_8_24# AND2X1_LOC_18/Y 0.01fF
C4463 AND2X1_LOC_20/a_8_24# AND2X1_LOC_18/Y -0.00fF
C4937 OR2X1_LOC_520/Y AND2X1_LOC_18/Y 0.03fF
C5037 AND2X1_LOC_107/a_8_24# AND2X1_LOC_18/Y 0.02fF
C6520 OR2X1_LOC_653/B AND2X1_LOC_18/Y 0.01fF
C7196 AND2X1_LOC_79/a_8_24# AND2X1_LOC_18/Y 0.06fF
C7506 OR2X1_LOC_100/Y AND2X1_LOC_18/Y 0.08fF
C7658 OR2X1_LOC_532/B AND2X1_LOC_18/Y 0.24fF
C8387 OR2X1_LOC_114/a_8_216# AND2X1_LOC_18/Y 0.02fF
C9049 AND2X1_LOC_432/a_8_24# AND2X1_LOC_18/Y 0.02fF
C9368 AND2X1_LOC_496/a_36_24# AND2X1_LOC_18/Y 0.01fF
C9604 AND2X1_LOC_18/Y AND2X1_LOC_265/a_8_24# 0.13fF
C9614 VDD AND2X1_LOC_18/Y 1.16fF
C9866 OR2X1_LOC_845/A AND2X1_LOC_18/Y 0.07fF
C10359 AND2X1_LOC_18/Y OR2X1_LOC_523/A 0.04fF
C10465 OR2X1_LOC_676/Y AND2X1_LOC_18/Y 0.07fF
C11655 AND2X1_LOC_18/Y OR2X1_LOC_115/B 0.02fF
C12334 AND2X1_LOC_134/a_8_24# AND2X1_LOC_18/Y 0.02fF
C12648 OR2X1_LOC_160/A AND2X1_LOC_18/Y 0.54fF
C12711 AND2X1_LOC_86/B AND2X1_LOC_18/Y 0.01fF
C12721 OR2X1_LOC_624/B AND2X1_LOC_18/Y 0.18fF
C12978 OR2X1_LOC_266/A AND2X1_LOC_18/Y 0.01fF
C12995 AND2X1_LOC_18/Y AND2X1_LOC_607/a_8_24# 0.03fF
C13461 OR2X1_LOC_78/Y AND2X1_LOC_18/Y 0.01fF
C13922 OR2X1_LOC_608/a_8_216# AND2X1_LOC_18/Y 0.04fF
C13941 OR2X1_LOC_185/A AND2X1_LOC_18/Y 6.66fF
C14425 OR2X1_LOC_702/A AND2X1_LOC_18/Y 0.13fF
C14680 AND2X1_LOC_262/a_8_24# AND2X1_LOC_18/Y 0.03fF
C14813 AND2X1_LOC_481/a_8_24# AND2X1_LOC_18/Y 0.14fF
C15099 AND2X1_LOC_18/Y OR2X1_LOC_641/A 0.05fF
C15196 OR2X1_LOC_114/Y AND2X1_LOC_18/Y 0.01fF
C15589 AND2X1_LOC_18/Y OR2X1_LOC_541/B 0.06fF
C16056 OR2X1_LOC_643/A AND2X1_LOC_18/Y 0.15fF
C16128 OR2X1_LOC_113/A AND2X1_LOC_18/Y 0.01fF
C16307 AND2X1_LOC_91/B AND2X1_LOC_18/Y 0.32fF
C16776 AND2X1_LOC_18/Y OR2X1_LOC_719/B 0.02fF
C16800 OR2X1_LOC_542/B AND2X1_LOC_18/Y 0.03fF
C16916 AND2X1_LOC_56/B AND2X1_LOC_18/Y 1.46fF
C18308 AND2X1_LOC_47/Y AND2X1_LOC_18/Y 1.11fF
C18495 AND2X1_LOC_521/a_8_24# AND2X1_LOC_18/Y 0.05fF
C18779 AND2X1_LOC_18/Y OR2X1_LOC_227/Y 0.03fF
C19057 OR2X1_LOC_99/Y AND2X1_LOC_18/Y 0.20fF
C19267 AND2X1_LOC_18/Y AND2X1_LOC_41/Y 0.06fF
C19361 OR2X1_LOC_621/A AND2X1_LOC_18/Y 0.17fF
C19594 OR2X1_LOC_434/A AND2X1_LOC_18/Y 0.52fF
C20257 OR2X1_LOC_235/B AND2X1_LOC_18/Y 0.05fF
C21063 AND2X1_LOC_18/Y OR2X1_LOC_362/A 0.07fF
C21075 OR2X1_LOC_832/a_8_216# AND2X1_LOC_18/Y 0.01fF
C21446 AND2X1_LOC_18/Y OR2X1_LOC_771/B 0.06fF
C22347 AND2X1_LOC_18/Y AND2X1_LOC_44/Y 0.51fF
C22601 OR2X1_LOC_720/B AND2X1_LOC_18/Y 0.03fF
C23531 AND2X1_LOC_18/Y OR2X1_LOC_789/A 0.03fF
C23743 AND2X1_LOC_394/a_8_24# AND2X1_LOC_18/Y 0.01fF
C24051 OR2X1_LOC_523/B AND2X1_LOC_18/Y 0.09fF
C24128 OR2X1_LOC_101/a_8_216# AND2X1_LOC_18/Y 0.02fF
C24134 OR2X1_LOC_231/A AND2X1_LOC_18/Y 0.03fF
C24168 OR2X1_LOC_130/A AND2X1_LOC_18/Y 0.62fF
C25839 OR2X1_LOC_555/A AND2X1_LOC_18/Y 0.18fF
C26213 OR2X1_LOC_790/B AND2X1_LOC_18/Y 0.23fF
C26291 AND2X1_LOC_51/Y AND2X1_LOC_18/Y 0.11fF
C26647 AND2X1_LOC_18/Y OR2X1_LOC_541/a_8_216# 0.01fF
C27116 OR2X1_LOC_631/B AND2X1_LOC_18/Y 0.03fF
C28149 AND2X1_LOC_18/Y OR2X1_LOC_71/A 0.02fF
C28552 AND2X1_LOC_31/Y AND2X1_LOC_18/Y 0.63fF
C28798 OR2X1_LOC_633/B AND2X1_LOC_18/Y 0.03fF
C29424 AND2X1_LOC_18/Y AND2X1_LOC_36/Y 2.38fF
C29538 OR2X1_LOC_630/Y AND2X1_LOC_18/Y 0.07fF
C30331 AND2X1_LOC_522/a_8_24# AND2X1_LOC_18/Y 0.03fF
C30727 AND2X1_LOC_60/a_8_24# AND2X1_LOC_18/Y 0.01fF
C31237 OR2X1_LOC_768/A AND2X1_LOC_18/Y 0.01fF
C32013 AND2X1_LOC_172/a_8_24# AND2X1_LOC_18/Y 0.01fF
C32788 AND2X1_LOC_18/Y OR2X1_LOC_777/B 0.03fF
C32830 OR2X1_LOC_188/a_8_216# AND2X1_LOC_18/Y -0.00fF
C33049 OR2X1_LOC_456/A AND2X1_LOC_18/Y 0.44fF
C33337 OR2X1_LOC_435/B AND2X1_LOC_18/Y 0.01fF
C33830 AND2X1_LOC_132/a_8_24# AND2X1_LOC_18/Y 0.01fF
C34662 OR2X1_LOC_400/A AND2X1_LOC_18/Y 0.01fF
C35090 OR2X1_LOC_790/a_8_216# AND2X1_LOC_18/Y 0.01fF
C35897 OR2X1_LOC_318/Y AND2X1_LOC_18/Y 0.07fF
C37600 AND2X1_LOC_18/Y OR2X1_LOC_553/A 0.24fF
C38335 OR2X1_LOC_151/A AND2X1_LOC_18/Y 0.14fF
C38840 OR2X1_LOC_174/A AND2X1_LOC_18/Y 0.11fF
C38879 AND2X1_LOC_482/a_8_24# AND2X1_LOC_18/Y 0.01fF
C39322 OR2X1_LOC_137/B AND2X1_LOC_18/Y 0.03fF
C39364 AND2X1_LOC_252/a_8_24# AND2X1_LOC_18/Y 0.01fF
C39671 AND2X1_LOC_18/Y AND2X1_LOC_616/a_8_24# 0.10fF
C40330 AND2X1_LOC_497/a_8_24# AND2X1_LOC_18/Y 0.04fF
C40726 AND2X1_LOC_109/a_8_24# AND2X1_LOC_18/Y 0.01fF
C41764 OR2X1_LOC_61/A AND2X1_LOC_18/Y 0.01fF
C42205 AND2X1_LOC_18/Y OR2X1_LOC_390/A 0.04fF
C42777 OR2X1_LOC_668/Y AND2X1_LOC_18/Y 0.02fF
C42985 AND2X1_LOC_18/Y OR2X1_LOC_344/a_8_216# 0.14fF
C43082 AND2X1_LOC_229/a_8_24# AND2X1_LOC_18/Y 0.01fF
C43128 OR2X1_LOC_841/A AND2X1_LOC_18/Y 0.10fF
C43355 OR2X1_LOC_84/A AND2X1_LOC_18/Y 0.03fF
C43553 OR2X1_LOC_190/A AND2X1_LOC_18/Y 0.03fF
C43823 AND2X1_LOC_18/Y OR2X1_LOC_241/B 0.70fF
C43942 OR2X1_LOC_188/Y AND2X1_LOC_18/Y 0.01fF
C44138 OR2X1_LOC_193/A AND2X1_LOC_18/Y 0.03fF
C44322 AND2X1_LOC_18/Y OR2X1_LOC_339/A 0.07fF
C44401 AND2X1_LOC_505/a_8_24# AND2X1_LOC_18/Y 0.03fF
C45405 OR2X1_LOC_810/A AND2X1_LOC_18/Y 0.17fF
C45695 OR2X1_LOC_715/B AND2X1_LOC_18/Y 0.10fF
C46228 OR2X1_LOC_656/B AND2X1_LOC_18/Y 0.01fF
C46273 OR2X1_LOC_793/A AND2X1_LOC_18/Y 0.01fF
C46360 AND2X1_LOC_45/a_8_24# AND2X1_LOC_18/Y 0.01fF
C46740 AND2X1_LOC_399/a_8_24# AND2X1_LOC_18/Y 0.01fF
C47550 OR2X1_LOC_78/A AND2X1_LOC_18/Y 0.18fF
C48456 OR2X1_LOC_147/B AND2X1_LOC_18/Y 0.03fF
C48468 AND2X1_LOC_517/a_8_24# AND2X1_LOC_18/Y 0.02fF
C48494 AND2X1_LOC_669/a_8_24# AND2X1_LOC_18/Y 0.02fF
C48757 OR2X1_LOC_231/B AND2X1_LOC_18/Y 0.03fF
C48782 OR2X1_LOC_114/B AND2X1_LOC_18/Y 0.03fF
C48934 AND2X1_LOC_79/Y AND2X1_LOC_18/Y 0.03fF
C48944 AND2X1_LOC_496/a_8_24# AND2X1_LOC_18/Y 0.07fF
C50138 OR2X1_LOC_833/B AND2X1_LOC_18/Y 0.01fF
C50157 OR2X1_LOC_254/B AND2X1_LOC_18/Y 0.01fF
C51921 OR2X1_LOC_196/B AND2X1_LOC_18/Y 0.09fF
C51978 OR2X1_LOC_112/B AND2X1_LOC_18/Y 0.02fF
C52294 OR2X1_LOC_574/A AND2X1_LOC_18/Y 0.10fF
C52636 AND2X1_LOC_58/a_8_24# AND2X1_LOC_18/Y 0.01fF
C52941 AND2X1_LOC_18/Y OR2X1_LOC_539/B 0.13fF
C53114 OR2X1_LOC_375/A AND2X1_LOC_18/Y 1.64fF
C53415 AND2X1_LOC_18/Y OR2X1_LOC_549/A 0.15fF
C53465 OR2X1_LOC_113/Y AND2X1_LOC_18/Y 0.01fF
C53885 OR2X1_LOC_499/B AND2X1_LOC_18/Y 0.12fF
C54135 AND2X1_LOC_18/Y OR2X1_LOC_348/B 0.77fF
C55232 OR2X1_LOC_673/Y AND2X1_LOC_18/Y 0.51fF
C55263 OR2X1_LOC_195/A AND2X1_LOC_18/Y 0.98fF
C55534 AND2X1_LOC_505/a_36_24# AND2X1_LOC_18/Y 0.01fF
C55942 OR2X1_LOC_139/A AND2X1_LOC_18/Y 0.07fF
C56641 AND2X1_LOC_18/Y VSS -5.89fF
C162 OR2X1_LOC_833/B AND2X1_LOC_36/Y 0.08fF
C186 OR2X1_LOC_254/B AND2X1_LOC_36/Y 0.01fF
C213 OR2X1_LOC_646/A AND2X1_LOC_36/Y 0.06fF
C617 AND2X1_LOC_32/a_8_24# AND2X1_LOC_36/Y 0.01fF
C1426 OR2X1_LOC_629/B AND2X1_LOC_36/Y 0.01fF
C1803 AND2X1_LOC_36/Y OR2X1_LOC_338/A 0.07fF
C1822 OR2X1_LOC_186/Y AND2X1_LOC_36/Y 0.07fF
C2000 OR2X1_LOC_196/B AND2X1_LOC_36/Y 0.03fF
C2404 OR2X1_LOC_574/A AND2X1_LOC_36/Y 0.01fF
C2698 OR2X1_LOC_855/A AND2X1_LOC_36/Y 0.28fF
C2701 AND2X1_LOC_627/a_8_24# AND2X1_LOC_36/Y 0.03fF
C3222 OR2X1_LOC_375/A AND2X1_LOC_36/Y 8.48fF
C3458 AND2X1_LOC_36/Y OR2X1_LOC_515/Y 0.01fF
C3559 AND2X1_LOC_36/Y OR2X1_LOC_549/A 0.29fF
C4022 OR2X1_LOC_499/B AND2X1_LOC_36/Y 0.01fF
C4416 OR2X1_LOC_181/B AND2X1_LOC_36/Y 0.18fF
C5280 OR2X1_LOC_195/A AND2X1_LOC_36/Y 0.01fF
C5632 OR2X1_LOC_769/B AND2X1_LOC_36/Y 0.07fF
C6014 OR2X1_LOC_139/A AND2X1_LOC_36/Y 0.04fF
C6054 AND2X1_LOC_179/a_8_24# AND2X1_LOC_36/Y 0.08fF
C6442 AND2X1_LOC_36/Y OR2X1_LOC_138/A 0.01fF
C6921 AND2X1_LOC_626/a_36_24# AND2X1_LOC_36/Y 0.01fF
C7891 OR2X1_LOC_403/B AND2X1_LOC_36/Y 0.03fF
C7914 OR2X1_LOC_622/a_8_216# AND2X1_LOC_36/Y 0.01fF
C7921 AND2X1_LOC_528/a_36_24# AND2X1_LOC_36/Y 0.01fF
C8663 OR2X1_LOC_97/A AND2X1_LOC_36/Y 0.03fF
C8736 AND2X1_LOC_290/a_8_24# AND2X1_LOC_36/Y 0.01fF
C9411 AND2X1_LOC_36/Y OR2X1_LOC_546/A 0.53fF
C9660 AND2X1_LOC_484/a_36_24# AND2X1_LOC_36/Y 0.01fF
C10011 OR2X1_LOC_154/A AND2X1_LOC_36/Y 2.56fF
C10063 OR2X1_LOC_778/A AND2X1_LOC_36/Y 0.01fF
C10226 AND2X1_LOC_36/Y OR2X1_LOC_198/A 0.02fF
C11163 OR2X1_LOC_633/A AND2X1_LOC_36/Y 0.03fF
C12543 OR2X1_LOC_379/a_8_216# AND2X1_LOC_36/Y 0.01fF
C12908 OR2X1_LOC_614/Y AND2X1_LOC_36/Y 0.26fF
C13494 AND2X1_LOC_79/a_8_24# AND2X1_LOC_36/Y 0.14fF
C13954 OR2X1_LOC_532/B AND2X1_LOC_36/Y 3.45fF
C14590 OR2X1_LOC_855/a_8_216# AND2X1_LOC_36/Y 0.01fF
C15841 VDD AND2X1_LOC_36/Y 1.73fF
C16306 OR2X1_LOC_334/B AND2X1_LOC_36/Y 0.01fF
C16706 OR2X1_LOC_676/Y AND2X1_LOC_36/Y 0.09fF
C16782 OR2X1_LOC_462/B AND2X1_LOC_36/Y 0.03fF
C17132 AND2X1_LOC_83/a_8_24# AND2X1_LOC_36/Y 0.01fF
C18016 OR2X1_LOC_840/A AND2X1_LOC_36/Y 0.14fF
C18083 OR2X1_LOC_789/a_8_216# AND2X1_LOC_36/Y 0.02fF
C18418 AND2X1_LOC_754/a_8_24# AND2X1_LOC_36/Y 0.01fF
C18916 OR2X1_LOC_160/A AND2X1_LOC_36/Y 0.27fF
C18947 AND2X1_LOC_86/B AND2X1_LOC_36/Y 0.03fF
C18956 OR2X1_LOC_624/B AND2X1_LOC_36/Y 0.45fF
C19243 OR2X1_LOC_196/Y AND2X1_LOC_36/Y 0.09fF
C19336 OR2X1_LOC_447/A AND2X1_LOC_36/Y 0.03fF
C19740 OR2X1_LOC_78/Y AND2X1_LOC_36/Y 0.11fF
C19856 AND2X1_LOC_491/a_8_24# AND2X1_LOC_36/Y 0.03fF
C20215 OR2X1_LOC_185/A AND2X1_LOC_36/Y 0.67fF
C21133 AND2X1_LOC_442/a_8_24# AND2X1_LOC_36/Y 0.07fF
C21508 OR2X1_LOC_379/Y AND2X1_LOC_36/Y 0.04fF
C21930 AND2X1_LOC_617/a_8_24# AND2X1_LOC_36/Y 0.01fF
C22336 OR2X1_LOC_637/A AND2X1_LOC_36/Y 0.01fF
C22384 OR2X1_LOC_778/Y AND2X1_LOC_36/Y 0.05fF
C22700 AND2X1_LOC_91/B AND2X1_LOC_36/Y 0.29fF
C22821 AND2X1_LOC_72/Y AND2X1_LOC_36/Y 0.03fF
C23099 OR2X1_LOC_147/a_36_216# AND2X1_LOC_36/Y 0.02fF
C23135 AND2X1_LOC_36/Y OR2X1_LOC_719/B 0.02fF
C23154 OR2X1_LOC_542/B AND2X1_LOC_36/Y 0.03fF
C23234 AND2X1_LOC_56/B AND2X1_LOC_36/Y 1.46fF
C23980 OR2X1_LOC_790/A AND2X1_LOC_36/Y 0.03fF
C24268 AND2X1_LOC_36/Y AND2X1_LOC_751/a_8_24# 0.01fF
C24558 AND2X1_LOC_47/Y AND2X1_LOC_36/Y 0.26fF
C24779 OR2X1_LOC_34/A AND2X1_LOC_36/Y 0.01fF
C24790 AND2X1_LOC_627/a_36_24# AND2X1_LOC_36/Y 0.01fF
C24803 OR2X1_LOC_646/B AND2X1_LOC_36/Y 0.03fF
C24865 OR2X1_LOC_506/A AND2X1_LOC_36/Y 0.13fF
C25286 OR2X1_LOC_633/Y AND2X1_LOC_36/Y 0.10fF
C25315 OR2X1_LOC_99/Y AND2X1_LOC_36/Y 0.15fF
C25536 AND2X1_LOC_36/Y AND2X1_LOC_41/Y 0.03fF
C25640 OR2X1_LOC_621/A AND2X1_LOC_36/Y 0.01fF
C26507 OR2X1_LOC_235/B AND2X1_LOC_36/Y 0.07fF
C26552 AND2X1_LOC_393/a_8_24# AND2X1_LOC_36/Y 0.01fF
C27651 AND2X1_LOC_36/Y OR2X1_LOC_771/B 9.25fF
C27673 AND2X1_LOC_36/Y OR2X1_LOC_776/A 0.06fF
C28482 AND2X1_LOC_36/Y OR2X1_LOC_317/B 0.03fF
C28572 AND2X1_LOC_36/Y AND2X1_LOC_44/Y 0.43fF
C29102 OR2X1_LOC_793/B AND2X1_LOC_36/Y 0.21fF
C29705 AND2X1_LOC_36/Y OR2X1_LOC_789/A 0.51fF
C30019 AND2X1_LOC_69/a_8_24# AND2X1_LOC_36/Y 0.10fF
C30344 OR2X1_LOC_447/a_8_216# AND2X1_LOC_36/Y 0.01fF
C30369 AND2X1_LOC_7/a_8_24# AND2X1_LOC_36/Y 0.01fF
C30786 OR2X1_LOC_449/B AND2X1_LOC_36/Y 0.04fF
C31041 AND2X1_LOC_36/Y OR2X1_LOC_195/a_8_216# 0.01fF
C31124 OR2X1_LOC_621/B AND2X1_LOC_36/Y 0.12fF
C32004 OR2X1_LOC_400/B AND2X1_LOC_36/Y 0.05fF
C32091 OR2X1_LOC_447/Y AND2X1_LOC_36/Y 0.01fF
C32319 OR2X1_LOC_709/B AND2X1_LOC_36/Y 0.18fF
C32408 OR2X1_LOC_240/B AND2X1_LOC_36/Y 0.05fF
C32479 AND2X1_LOC_51/Y AND2X1_LOC_36/Y 0.28fF
C32872 OR2X1_LOC_831/a_8_216# AND2X1_LOC_36/Y 0.01fF
C33304 OR2X1_LOC_631/B AND2X1_LOC_36/Y 0.02fF
C33668 AND2X1_LOC_524/a_8_24# AND2X1_LOC_36/Y 0.05fF
C33965 AND2X1_LOC_36/Y OR2X1_LOC_704/a_8_216# 0.01fF
C34345 AND2X1_LOC_36/Y OR2X1_LOC_71/A 0.07fF
C34766 AND2X1_LOC_31/Y AND2X1_LOC_36/Y 5.99fF
C35028 OR2X1_LOC_240/A AND2X1_LOC_36/Y 0.02fF
C35032 OR2X1_LOC_633/B AND2X1_LOC_36/Y 0.06fF
C35774 OR2X1_LOC_633/a_8_216# AND2X1_LOC_36/Y 0.01fF
C35817 AND2X1_LOC_586/a_8_24# AND2X1_LOC_36/Y 0.02fF
C35995 AND2X1_LOC_36/Y OR2X1_LOC_196/a_8_216# 0.01fF
C36563 OR2X1_LOC_856/A AND2X1_LOC_36/Y 0.01fF
C36578 AND2X1_LOC_313/a_8_24# AND2X1_LOC_36/Y 0.01fF
C37834 OR2X1_LOC_709/a_8_216# AND2X1_LOC_36/Y 0.01fF
C37905 OR2X1_LOC_240/a_8_216# AND2X1_LOC_36/Y 0.01fF
C37999 AND2X1_LOC_146/a_8_24# AND2X1_LOC_36/Y 0.09fF
C39064 AND2X1_LOC_36/Y OR2X1_LOC_777/B 0.05fF
C39285 OR2X1_LOC_456/A AND2X1_LOC_36/Y 0.15fF
C39997 OR2X1_LOC_630/B AND2X1_LOC_36/Y 0.01fF
C40504 OR2X1_LOC_644/B AND2X1_LOC_36/Y 0.02fF
C40617 OR2X1_LOC_673/A AND2X1_LOC_36/Y 0.03fF
C40653 OR2X1_LOC_705/B AND2X1_LOC_36/Y 0.08fF
C41377 OR2X1_LOC_647/B AND2X1_LOC_36/Y 0.07fF
C41828 AND2X1_LOC_528/a_8_24# AND2X1_LOC_36/Y 0.04fF
C42152 OR2X1_LOC_621/a_8_216# AND2X1_LOC_36/Y 0.01fF
C43130 OR2X1_LOC_147/a_8_216# AND2X1_LOC_36/Y 0.03fF
C43469 AND2X1_LOC_498/a_8_24# AND2X1_LOC_36/Y 0.01fF
C43470 AND2X1_LOC_320/a_8_24# AND2X1_LOC_36/Y 0.10fF
C43562 OR2X1_LOC_287/B AND2X1_LOC_36/Y 0.02fF
C43969 OR2X1_LOC_553/A AND2X1_LOC_36/Y 0.07fF
C44736 OR2X1_LOC_151/A AND2X1_LOC_36/Y 0.12fF
C44737 AND2X1_LOC_524/a_36_24# AND2X1_LOC_36/Y 0.01fF
C45086 AND2X1_LOC_36/Y OR2X1_LOC_714/A 0.01fF
C45240 AND2X1_LOC_482/a_8_24# AND2X1_LOC_36/Y 0.01fF
C45714 AND2X1_LOC_252/a_8_24# AND2X1_LOC_36/Y 0.01fF
C46084 AND2X1_LOC_616/a_8_24# AND2X1_LOC_36/Y 0.01fF
C47364 AND2X1_LOC_36/Y OR2X1_LOC_308/Y 0.09fF
C47540 AND2X1_LOC_516/a_8_24# AND2X1_LOC_36/Y 0.01fF
C48486 AND2X1_LOC_7/Y AND2X1_LOC_36/Y 0.01fF
C49104 OR2X1_LOC_711/B AND2X1_LOC_36/Y 0.08fF
C49184 OR2X1_LOC_243/A AND2X1_LOC_36/Y 0.01fF
C49785 OR2X1_LOC_84/A AND2X1_LOC_36/Y 0.01fF
C50008 OR2X1_LOC_190/A AND2X1_LOC_36/Y 0.15fF
C50388 OR2X1_LOC_188/Y AND2X1_LOC_36/Y 1.20fF
C50458 AND2X1_LOC_423/a_8_24# AND2X1_LOC_36/Y 0.01fF
C50527 OR2X1_LOC_193/A AND2X1_LOC_36/Y 0.02fF
C50821 OR2X1_LOC_673/B AND2X1_LOC_36/Y 0.02fF
C50827 OR2X1_LOC_831/A AND2X1_LOC_36/Y 0.20fF
C50837 OR2X1_LOC_598/Y AND2X1_LOC_36/Y 0.17fF
C51383 AND2X1_LOC_698/a_8_24# AND2X1_LOC_36/Y 0.01fF
C52054 OR2X1_LOC_715/B AND2X1_LOC_36/Y 0.12fF
C52057 AND2X1_LOC_626/a_8_24# AND2X1_LOC_36/Y 0.04fF
C52587 OR2X1_LOC_793/A AND2X1_LOC_36/Y 0.17fF
C53008 OR2X1_LOC_687/Y AND2X1_LOC_36/Y 0.03fF
C53258 AND2X1_LOC_36/Y OR2X1_LOC_199/B 0.11fF
C53338 OR2X1_LOC_622/A AND2X1_LOC_36/Y 0.28fF
C53433 OR2X1_LOC_835/B AND2X1_LOC_36/Y 0.07fF
C53804 OR2X1_LOC_78/A AND2X1_LOC_36/Y 0.17fF
C54627 OR2X1_LOC_501/B AND2X1_LOC_36/Y 0.01fF
C54649 OR2X1_LOC_147/B AND2X1_LOC_36/Y 0.10fF
C54714 AND2X1_LOC_484/a_8_24# AND2X1_LOC_36/Y 0.01fF
C54755 OR2X1_LOC_545/B AND2X1_LOC_36/Y 0.03fF
C54836 OR2X1_LOC_318/B AND2X1_LOC_36/Y 0.16fF
C55018 AND2X1_LOC_396/a_8_24# AND2X1_LOC_36/Y 0.06fF
C55092 OR2X1_LOC_841/B AND2X1_LOC_36/Y 0.04fF
C55119 AND2X1_LOC_79/Y AND2X1_LOC_36/Y 0.01fF
C55129 AND2X1_LOC_496/a_8_24# AND2X1_LOC_36/Y 0.01fF
C55545 AND2X1_LOC_495/a_8_24# AND2X1_LOC_36/Y 0.01fF
C55940 OR2X1_LOC_623/B AND2X1_LOC_36/Y 0.03fF
C56471 AND2X1_LOC_36/Y VSS -4.77fF
C9 AND2X1_LOC_525/a_8_24# OR2X1_LOC_375/A 0.01fF
C31 OR2X1_LOC_375/A AND2X1_LOC_51/Y 1.52fF
C54 OR2X1_LOC_836/Y OR2X1_LOC_375/A 0.02fF
C553 OR2X1_LOC_375/A AND2X1_LOC_52/Y 0.05fF
C1531 OR2X1_LOC_149/B OR2X1_LOC_375/A 0.72fF
C1877 OR2X1_LOC_375/A OR2X1_LOC_71/A 0.03fF
C2145 AND2X1_LOC_145/a_36_24# OR2X1_LOC_375/A 0.01fF
C2253 OR2X1_LOC_614/a_8_216# OR2X1_LOC_375/A 0.05fF
C2311 OR2X1_LOC_375/A AND2X1_LOC_31/Y 0.97fF
C2640 OR2X1_LOC_633/B OR2X1_LOC_375/A 1.75fF
C3156 OR2X1_LOC_375/A OR2X1_LOC_451/B 0.11fF
C3292 OR2X1_LOC_506/Y OR2X1_LOC_375/A 0.01fF
C3367 OR2X1_LOC_633/a_8_216# OR2X1_LOC_375/A 0.01fF
C3390 OR2X1_LOC_635/A OR2X1_LOC_375/A 0.07fF
C3474 AND2X1_LOC_122/a_8_24# OR2X1_LOC_375/A 0.01fF
C4617 AND2X1_LOC_504/a_8_24# OR2X1_LOC_375/A 0.11fF
C4695 AND2X1_LOC_117/a_8_24# OR2X1_LOC_375/A 0.01fF
C5523 OR2X1_LOC_546/B OR2X1_LOC_375/A 0.01fF
C6247 OR2X1_LOC_678/Y OR2X1_LOC_375/A 0.01fF
C6507 OR2X1_LOC_375/A OR2X1_LOC_777/B 5.11fF
C6574 OR2X1_LOC_188/a_8_216# OR2X1_LOC_375/A 0.01fF
C6580 OR2X1_LOC_156/Y OR2X1_LOC_375/A 0.10fF
C6840 OR2X1_LOC_456/A OR2X1_LOC_375/A 0.03fF
C7216 OR2X1_LOC_460/Y OR2X1_LOC_375/A 0.02fF
C7633 AND2X1_LOC_132/a_8_24# OR2X1_LOC_375/A 0.03fF
C7706 AND2X1_LOC_67/Y OR2X1_LOC_375/A 0.12fF
C7911 OR2X1_LOC_375/A OR2X1_LOC_259/A 0.01fF
C8234 OR2X1_LOC_673/A OR2X1_LOC_375/A 0.02fF
C8261 OR2X1_LOC_705/B OR2X1_LOC_375/A 0.53fF
C8965 OR2X1_LOC_790/a_8_216# OR2X1_LOC_375/A 0.02fF
C8992 OR2X1_LOC_375/A OR2X1_LOC_647/B 0.03fF
C10167 OR2X1_LOC_375/A AND2X1_LOC_232/a_36_24# 0.01fF
C10289 OR2X1_LOC_123/B OR2X1_LOC_375/A 0.02fF
C11090 OR2X1_LOC_287/B OR2X1_LOC_375/A 0.03fF
C11111 OR2X1_LOC_97/a_8_216# OR2X1_LOC_375/A 0.01fF
C11123 OR2X1_LOC_76/A OR2X1_LOC_375/A 0.03fF
C11147 OR2X1_LOC_148/A OR2X1_LOC_375/A 0.03fF
C11492 OR2X1_LOC_375/A OR2X1_LOC_553/A 0.07fF
C11646 OR2X1_LOC_375/A OR2X1_LOC_197/a_8_216# 0.02fF
C12199 OR2X1_LOC_151/A OR2X1_LOC_375/A 0.03fF
C12282 AND2X1_LOC_67/a_8_24# OR2X1_LOC_375/A 0.01fF
C12299 OR2X1_LOC_651/B OR2X1_LOC_375/A 0.04fF
C13666 OR2X1_LOC_375/A OR2X1_LOC_378/Y 0.21fF
C14685 OR2X1_LOC_375/A OR2X1_LOC_308/Y 0.01fF
C15647 OR2X1_LOC_448/A OR2X1_LOC_375/A 0.09fF
C15786 OR2X1_LOC_375/A AND2X1_LOC_7/Y 0.04fF
C15967 OR2X1_LOC_375/A OR2X1_LOC_706/a_8_216# 0.01fF
C16145 AND2X1_LOC_89/a_8_24# OR2X1_LOC_375/A 0.04fF
C16287 AND2X1_LOC_280/a_8_24# OR2X1_LOC_375/A 0.07fF
C16611 AND2X1_LOC_525/a_36_24# OR2X1_LOC_375/A 0.01fF
C16721 OR2X1_LOC_375/A OR2X1_LOC_344/a_8_216# 0.02fF
C17140 OR2X1_LOC_375/A OR2X1_LOC_98/B 0.09fF
C17317 OR2X1_LOC_190/A OR2X1_LOC_375/A 0.07fF
C17536 OR2X1_LOC_375/A OR2X1_LOC_241/B 0.06fF
C17652 OR2X1_LOC_188/Y OR2X1_LOC_375/A 0.09fF
C17752 AND2X1_LOC_189/a_8_24# OR2X1_LOC_375/A 0.01fF
C17893 OR2X1_LOC_193/A OR2X1_LOC_375/A 0.03fF
C18130 OR2X1_LOC_673/B OR2X1_LOC_375/A 0.06fF
C18946 OR2X1_LOC_375/A AND2X1_LOC_416/a_8_24# 0.10fF
C19165 OR2X1_LOC_810/A OR2X1_LOC_375/A 0.05fF
C19443 OR2X1_LOC_715/B OR2X1_LOC_375/A 0.03fF
C19448 OR2X1_LOC_375/A OR2X1_LOC_543/A 0.01fF
C19604 AND2X1_LOC_81/a_8_24# OR2X1_LOC_375/A 0.01fF
C20017 OR2X1_LOC_793/A OR2X1_LOC_375/A 0.01fF
C20082 AND2X1_LOC_45/a_8_24# OR2X1_LOC_375/A 0.01fF
C20432 OR2X1_LOC_687/Y OR2X1_LOC_375/A 0.03fF
C20641 OR2X1_LOC_375/A OR2X1_LOC_199/B 0.05fF
C21211 OR2X1_LOC_375/A OR2X1_LOC_78/A 1.89fF
C21739 OR2X1_LOC_97/B OR2X1_LOC_375/A 1.60fF
C22116 OR2X1_LOC_147/B OR2X1_LOC_375/A 0.05fF
C22303 OR2X1_LOC_375/A OR2X1_LOC_318/B 0.03fF
C22443 OR2X1_LOC_121/Y OR2X1_LOC_375/A 0.27fF
C22750 OR2X1_LOC_375/A OR2X1_LOC_98/a_8_216# 0.03fF
C23394 OR2X1_LOC_375/A OR2X1_LOC_623/B 0.03fF
C23741 OR2X1_LOC_507/A OR2X1_LOC_375/A 0.03fF
C25485 OR2X1_LOC_773/B OR2X1_LOC_375/A 0.08fF
C25574 OR2X1_LOC_196/B OR2X1_LOC_375/A 0.04fF
C25938 OR2X1_LOC_574/A OR2X1_LOC_375/A 0.05fF
C26807 OR2X1_LOC_605/B OR2X1_LOC_375/A 0.01fF
C27054 OR2X1_LOC_375/A OR2X1_LOC_549/A 0.25fF
C27749 OR2X1_LOC_375/A OR2X1_LOC_543/a_8_216# 0.01fF
C27766 OR2X1_LOC_375/A OR2X1_LOC_348/B 2.75fF
C28014 OR2X1_LOC_181/B OR2X1_LOC_375/A 0.03fF
C28186 OR2X1_LOC_375/A OR2X1_LOC_98/a_36_216# 0.02fF
C28318 OR2X1_LOC_375/A AND2X1_LOC_603/a_8_24# 0.01fF
C28870 OR2X1_LOC_673/Y OR2X1_LOC_375/A 0.03fF
C29550 OR2X1_LOC_139/A OR2X1_LOC_375/A 0.12fF
C29647 OR2X1_LOC_637/Y OR2X1_LOC_375/A 0.03fF
C30490 OR2X1_LOC_834/a_8_216# OR2X1_LOC_375/A 0.01fF
C30592 AND2X1_LOC_697/a_8_24# OR2X1_LOC_375/A 0.01fF
C30966 OR2X1_LOC_668/a_8_216# OR2X1_LOC_375/A 0.04fF
C31628 OR2X1_LOC_375/A OR2X1_LOC_130/a_8_216# 0.01fF
C32045 OR2X1_LOC_97/A OR2X1_LOC_375/A 3.27fF
C32148 OR2X1_LOC_541/A OR2X1_LOC_375/A 0.03fF
C32197 OR2X1_LOC_375/A AND2X1_LOC_282/a_8_24# 0.11fF
C32498 OR2X1_LOC_375/A OR2X1_LOC_713/A 0.43fF
C32828 OR2X1_LOC_375/A OR2X1_LOC_546/A 0.04fF
C32983 AND2X1_LOC_700/a_8_24# OR2X1_LOC_375/A 0.01fF
C33153 OR2X1_LOC_99/B OR2X1_LOC_375/A 0.01fF
C33237 OR2X1_LOC_590/a_8_216# OR2X1_LOC_375/A 0.01fF
C33527 OR2X1_LOC_154/A OR2X1_LOC_375/A 0.42fF
C33547 OR2X1_LOC_267/A OR2X1_LOC_375/A 0.03fF
C33588 OR2X1_LOC_778/A OR2X1_LOC_375/A 0.02fF
C33699 OR2X1_LOC_375/A OR2X1_LOC_198/A 0.01fF
C34264 OR2X1_LOC_634/A OR2X1_LOC_375/A 0.22fF
C34582 OR2X1_LOC_375/A OR2X1_LOC_267/Y 0.03fF
C34616 OR2X1_LOC_375/A OR2X1_LOC_633/A 0.11fF
C34629 OR2X1_LOC_673/a_8_216# OR2X1_LOC_375/A 0.01fF
C34995 OR2X1_LOC_375/A OR2X1_LOC_590/Y 0.01fF
C35932 OR2X1_LOC_124/B OR2X1_LOC_375/A 0.01fF
C35938 OR2X1_LOC_375/A OR2X1_LOC_370/a_8_216# 0.01fF
C36285 OR2X1_LOC_375/A OR2X1_LOC_779/A 0.01fF
C36324 OR2X1_LOC_614/Y OR2X1_LOC_375/A 0.01fF
C36845 OR2X1_LOC_463/B OR2X1_LOC_375/A 0.13fF
C37395 OR2X1_LOC_532/B OR2X1_LOC_375/A 2.03fF
C38470 OR2X1_LOC_710/B OR2X1_LOC_375/A 0.01fF
C38655 OR2X1_LOC_472/B OR2X1_LOC_375/A 0.39fF
C38739 OR2X1_LOC_375/A OR2X1_LOC_552/A 0.48fF
C38972 AND2X1_LOC_52/a_8_24# OR2X1_LOC_375/A 0.02fF
C39169 OR2X1_LOC_375/A OR2X1_LOC_192/B 0.01fF
C39333 VDD OR2X1_LOC_375/A 2.44fF
C40133 OR2X1_LOC_676/Y OR2X1_LOC_375/A 0.08fF
C40154 OR2X1_LOC_834/A OR2X1_LOC_375/A 0.01fF
C40256 OR2X1_LOC_462/B OR2X1_LOC_375/A 0.03fF
C40474 OR2X1_LOC_375/A AND2X1_LOC_591/a_8_24# 0.01fF
C41215 OR2X1_LOC_375/A AND2X1_LOC_667/a_8_24# 0.01fF
C41519 OR2X1_LOC_840/A OR2X1_LOC_375/A 0.01fF
C41554 OR2X1_LOC_260/a_8_216# OR2X1_LOC_375/A 0.18fF
C41571 AND2X1_LOC_145/a_8_24# OR2X1_LOC_375/A 0.04fF
C41950 OR2X1_LOC_216/A OR2X1_LOC_375/A 0.04fF
C42461 OR2X1_LOC_160/A OR2X1_LOC_375/A 0.10fF
C42505 OR2X1_LOC_624/B OR2X1_LOC_375/A 0.07fF
C42698 OR2X1_LOC_375/A OR2X1_LOC_130/Y 0.01fF
C43737 OR2X1_LOC_185/A OR2X1_LOC_375/A 0.28fF
C44202 AND2X1_LOC_158/a_8_24# OR2X1_LOC_375/A 0.04fF
C44472 OR2X1_LOC_375/A AND2X1_LOC_262/a_8_24# 0.01fF
C44648 AND2X1_LOC_481/a_8_24# OR2X1_LOC_375/A 0.04fF
C44912 OR2X1_LOC_375/A OR2X1_LOC_641/A 0.03fF
C45784 OR2X1_LOC_673/a_36_216# OR2X1_LOC_375/A 0.02fF
C45937 OR2X1_LOC_643/A OR2X1_LOC_375/A 0.03fF
C45942 OR2X1_LOC_375/A OR2X1_LOC_778/Y 0.13fF
C46180 AND2X1_LOC_91/B OR2X1_LOC_375/A 0.43fF
C46309 OR2X1_LOC_638/a_8_216# OR2X1_LOC_375/A 0.01fF
C46323 OR2X1_LOC_308/a_8_216# OR2X1_LOC_375/A 0.01fF
C46721 OR2X1_LOC_542/B OR2X1_LOC_375/A 0.03fF
C46845 AND2X1_LOC_56/B OR2X1_LOC_375/A 0.11fF
C47190 OR2X1_LOC_375/A OR2X1_LOC_787/B 0.01fF
C47605 OR2X1_LOC_790/A OR2X1_LOC_375/A 0.26fF
C47757 AND2X1_LOC_118/a_8_24# OR2X1_LOC_375/A 0.01fF
C48276 AND2X1_LOC_47/Y OR2X1_LOC_375/A 1.06fF
C48459 AND2X1_LOC_521/a_8_24# OR2X1_LOC_375/A 0.08fF
C48974 OR2X1_LOC_633/Y OR2X1_LOC_375/A 0.05fF
C49177 OR2X1_LOC_375/A AND2X1_LOC_41/Y 1.03fF
C49784 OR2X1_LOC_375/A AND2X1_LOC_232/a_8_24# 0.14fF
C50190 OR2X1_LOC_235/B OR2X1_LOC_375/A 0.14fF
C50696 OR2X1_LOC_791/B OR2X1_LOC_375/A 0.04fF
C51179 OR2X1_LOC_243/B OR2X1_LOC_375/A 0.03fF
C51286 OR2X1_LOC_375/A OR2X1_LOC_771/B 0.08fF
C51291 OR2X1_LOC_375/A OR2X1_LOC_209/A 0.02fF
C51435 OR2X1_LOC_678/a_8_216# OR2X1_LOC_375/A 0.01fF
C51741 OR2X1_LOC_375/A OR2X1_LOC_593/B 0.01fF
C51762 OR2X1_LOC_506/a_8_216# OR2X1_LOC_375/A 0.01fF
C51831 AND2X1_LOC_41/a_8_24# OR2X1_LOC_375/A 0.01fF
C52180 OR2X1_LOC_375/A AND2X1_LOC_44/Y 1.12fF
C52908 OR2X1_LOC_506/B OR2X1_LOC_375/A 0.01fF
C53037 OR2X1_LOC_375/A AND2X1_LOC_258/a_8_24# 0.06fF
C53525 OR2X1_LOC_375/A OR2X1_LOC_307/A 0.01fF
C54060 OR2X1_LOC_375/A AND2X1_LOC_612/a_8_24# 0.10fF
C54475 OR2X1_LOC_375/A OR2X1_LOC_449/B 0.03fF
C55609 OR2X1_LOC_375/A OR2X1_LOC_786/A 0.01fF
C55861 OR2X1_LOC_447/Y OR2X1_LOC_375/A 0.03fF
C56183 OR2X1_LOC_240/B OR2X1_LOC_375/A 0.02fF
C56186 OR2X1_LOC_790/B OR2X1_LOC_375/A 0.21fF
C56890 OR2X1_LOC_375/A VSS 0.75fF
C36 OR2X1_LOC_64/Y OR2X1_LOC_265/Y 0.03fF
C426 OR2X1_LOC_164/Y OR2X1_LOC_64/Y 0.40fF
C717 AND2X1_LOC_539/Y OR2X1_LOC_64/Y 0.02fF
C816 AND2X1_LOC_326/B OR2X1_LOC_64/Y 0.03fF
C1270 AND2X1_LOC_112/a_8_24# OR2X1_LOC_64/Y 0.01fF
C1709 OR2X1_LOC_64/Y AND2X1_LOC_434/Y 0.01fF
C1806 OR2X1_LOC_764/Y OR2X1_LOC_64/Y 0.02fF
C3322 AND2X1_LOC_776/Y OR2X1_LOC_64/Y 0.20fF
C3542 OR2X1_LOC_79/A OR2X1_LOC_64/Y 0.01fF
C3933 OR2X1_LOC_283/Y OR2X1_LOC_64/Y 0.05fF
C4612 OR2X1_LOC_597/A OR2X1_LOC_64/Y 0.01fF
C4814 OR2X1_LOC_64/Y AND2X1_LOC_318/Y 0.05fF
C4981 OR2X1_LOC_64/Y OR2X1_LOC_829/A 0.01fF
C5203 OR2X1_LOC_64/Y OR2X1_LOC_224/Y 0.01fF
C5212 OR2X1_LOC_64/Y OR2X1_LOC_597/Y 0.01fF
C5812 OR2X1_LOC_64/Y OR2X1_LOC_764/a_8_216# 0.01fF
C6736 AND2X1_LOC_715/A OR2X1_LOC_64/Y 0.04fF
C7279 AND2X1_LOC_729/Y OR2X1_LOC_64/Y 0.51fF
C7303 AND2X1_LOC_784/A OR2X1_LOC_64/Y 0.14fF
C7320 AND2X1_LOC_769/a_8_24# OR2X1_LOC_64/Y 0.01fF
C7745 OR2X1_LOC_64/Y OR2X1_LOC_52/B 0.32fF
C7754 AND2X1_LOC_489/Y OR2X1_LOC_64/Y 0.02fF
C8215 OR2X1_LOC_280/Y OR2X1_LOC_64/Y 0.03fF
C8534 OR2X1_LOC_485/Y OR2X1_LOC_64/Y 0.28fF
C9012 OR2X1_LOC_64/Y AND2X1_LOC_593/Y 0.01fF
C9111 OR2X1_LOC_64/Y OR2X1_LOC_226/Y 0.01fF
C9386 OR2X1_LOC_51/Y OR2X1_LOC_64/Y 2.25fF
C9473 OR2X1_LOC_680/A OR2X1_LOC_64/Y 1.55fF
C9483 OR2X1_LOC_667/a_8_216# OR2X1_LOC_64/Y 0.07fF
C10007 OR2X1_LOC_64/Y AND2X1_LOC_790/a_8_24# 0.17fF
C10218 OR2X1_LOC_64/Y AND2X1_LOC_436/Y 0.06fF
C10277 AND2X1_LOC_97/a_8_24# OR2X1_LOC_64/Y 0.26fF
C10311 OR2X1_LOC_64/Y OR2X1_LOC_588/Y 0.26fF
C10839 OR2X1_LOC_64/Y OR2X1_LOC_331/a_8_216# 0.04fF
C11129 OR2X1_LOC_64/Y AND2X1_LOC_266/Y 0.13fF
C11936 OR2X1_LOC_64/Y OR2X1_LOC_265/a_8_216# 0.06fF
C13321 OR2X1_LOC_64/Y OR2X1_LOC_74/A 0.12fF
C14141 OR2X1_LOC_64/Y OR2X1_LOC_235/a_8_216# 0.18fF
C14880 OR2X1_LOC_816/a_8_216# OR2X1_LOC_64/Y 0.01fF
C15355 OR2X1_LOC_497/a_8_216# OR2X1_LOC_64/Y 0.06fF
C15690 OR2X1_LOC_64/Y OR2X1_LOC_597/a_8_216# 0.15fF
C15739 AND2X1_LOC_99/A OR2X1_LOC_64/Y 0.12fF
C15778 OR2X1_LOC_64/Y AND2X1_LOC_637/Y 0.03fF
C16262 OR2X1_LOC_696/Y OR2X1_LOC_64/Y 0.09fF
C16291 OR2X1_LOC_167/Y OR2X1_LOC_64/Y 0.02fF
C16433 OR2X1_LOC_64/Y OR2X1_LOC_503/a_8_216# 0.06fF
C16500 AND2X1_LOC_362/B OR2X1_LOC_64/Y 0.02fF
C17507 OR2X1_LOC_420/a_8_216# OR2X1_LOC_64/Y 0.02fF
C17875 OR2X1_LOC_695/a_8_216# OR2X1_LOC_64/Y 0.02fF
C19963 AND2X1_LOC_714/B OR2X1_LOC_64/Y 0.03fF
C21067 OR2X1_LOC_64/Y AND2X1_LOC_793/B 0.35fF
C22048 OR2X1_LOC_64/Y OR2X1_LOC_503/a_36_216# 0.03fF
C22142 VDD OR2X1_LOC_64/Y 1.98fF
C22212 OR2X1_LOC_829/a_8_216# OR2X1_LOC_64/Y 0.14fF
C22245 OR2X1_LOC_251/Y OR2X1_LOC_64/Y 0.07fF
C22345 OR2X1_LOC_64/Y OR2X1_LOC_67/Y 0.07fF
C23091 OR2X1_LOC_64/Y OR2X1_LOC_591/A 0.05fF
C23107 OR2X1_LOC_420/a_36_216# OR2X1_LOC_64/Y 0.02fF
C23129 OR2X1_LOC_64/Y AND2X1_LOC_307/Y 0.02fF
C24088 OR2X1_LOC_64/Y AND2X1_LOC_592/a_8_24# 0.03fF
C24560 OR2X1_LOC_64/Y OR2X1_LOC_184/a_8_216# 0.01fF
C24994 OR2X1_LOC_45/B OR2X1_LOC_64/Y 0.38fF
C25443 OR2X1_LOC_158/A OR2X1_LOC_64/Y 0.15fF
C25525 OR2X1_LOC_103/Y OR2X1_LOC_64/Y 0.01fF
C25543 OR2X1_LOC_103/a_8_216# OR2X1_LOC_64/Y 0.01fF
C25858 OR2X1_LOC_482/Y OR2X1_LOC_64/Y 0.83fF
C25903 OR2X1_LOC_816/Y OR2X1_LOC_64/Y 0.12fF
C26909 OR2X1_LOC_111/Y OR2X1_LOC_64/Y 0.15fF
C27159 OR2X1_LOC_591/Y OR2X1_LOC_64/Y 0.01fF
C27488 OR2X1_LOC_64/Y AND2X1_LOC_227/a_8_24# 0.01fF
C27599 OR2X1_LOC_107/a_8_216# OR2X1_LOC_64/Y 0.07fF
C27709 AND2X1_LOC_390/B OR2X1_LOC_64/Y 0.04fF
C27733 AND2X1_LOC_101/a_8_24# OR2X1_LOC_64/Y 0.01fF
C28000 OR2X1_LOC_309/Y OR2X1_LOC_64/Y 0.03fF
C28119 OR2X1_LOC_64/Y AND2X1_LOC_840/B 0.12fF
C28316 OR2X1_LOC_64/Y OR2X1_LOC_320/a_8_216# 0.11fF
C28378 OR2X1_LOC_64/Y OR2X1_LOC_79/a_8_216# 0.01fF
C28434 OR2X1_LOC_694/Y OR2X1_LOC_64/Y 0.01fF
C28792 OR2X1_LOC_821/a_8_216# OR2X1_LOC_64/Y 0.01fF
C29309 OR2X1_LOC_64/Y AND2X1_LOC_638/Y 0.01fF
C29796 OR2X1_LOC_91/Y OR2X1_LOC_64/Y 0.52fF
C29831 OR2X1_LOC_527/Y OR2X1_LOC_64/Y 0.13fF
C29839 OR2X1_LOC_417/Y OR2X1_LOC_64/Y 0.03fF
C29847 OR2X1_LOC_311/Y OR2X1_LOC_64/Y 0.02fF
C30291 OR2X1_LOC_64/Y AND2X1_LOC_831/Y 0.41fF
C30610 OR2X1_LOC_64/Y AND2X1_LOC_436/B 0.02fF
C30985 OR2X1_LOC_484/a_8_216# OR2X1_LOC_64/Y 0.01fF
C31355 OR2X1_LOC_492/Y OR2X1_LOC_64/Y 0.07fF
C31889 OR2X1_LOC_497/Y OR2X1_LOC_64/Y 0.53fF
C32249 OR2X1_LOC_109/a_8_216# OR2X1_LOC_64/Y 0.13fF
C32666 OR2X1_LOC_235/B OR2X1_LOC_64/Y 0.66fF
C32740 AND2X1_LOC_319/A OR2X1_LOC_64/Y 0.10fF
C32836 OR2X1_LOC_64/Y AND2X1_LOC_721/A 0.03fF
C32866 OR2X1_LOC_64/Y OR2X1_LOC_331/Y 0.19fF
C33170 OR2X1_LOC_64/Y AND2X1_LOC_361/A 0.07fF
C33858 AND2X1_LOC_787/A OR2X1_LOC_64/Y 0.03fF
C33931 OR2X1_LOC_695/Y OR2X1_LOC_64/Y 0.01fF
C34702 OR2X1_LOC_692/Y OR2X1_LOC_64/Y 0.04fF
C34715 AND2X1_LOC_729/a_8_24# OR2X1_LOC_64/Y 0.01fF
C34748 AND2X1_LOC_335/Y OR2X1_LOC_64/Y 0.03fF
C34850 OR2X1_LOC_64/Y OR2X1_LOC_619/Y 0.04fF
C35110 OR2X1_LOC_64/Y AND2X1_LOC_769/Y 0.03fF
C35261 OR2X1_LOC_64/Y AND2X1_LOC_454/A 0.09fF
C35606 OR2X1_LOC_331/A OR2X1_LOC_64/Y 0.03fF
C35994 OR2X1_LOC_329/Y OR2X1_LOC_64/Y 0.01fF
C36471 AND2X1_LOC_99/a_8_24# OR2X1_LOC_64/Y 0.01fF
C36940 OR2X1_LOC_312/Y OR2X1_LOC_64/Y 0.03fF
C37110 OR2X1_LOC_64/Y OR2X1_LOC_13/B 1.86fF
C37640 OR2X1_LOC_64/Y OR2X1_LOC_595/A 0.51fF
C38074 AND2X1_LOC_592/Y OR2X1_LOC_64/Y 0.01fF
C38232 OR2X1_LOC_64/Y AND2X1_LOC_105/a_8_24# 0.01fF
C38681 OR2X1_LOC_64/Y OR2X1_LOC_89/A 3.67fF
C38953 OR2X1_LOC_167/a_8_216# OR2X1_LOC_64/Y 0.08fF
C39363 OR2X1_LOC_64/Y OR2X1_LOC_79/Y 0.02fF
C39429 AND2X1_LOC_707/a_8_24# OR2X1_LOC_64/Y 0.11fF
C39467 OR2X1_LOC_251/a_8_216# OR2X1_LOC_64/Y 0.01fF
C39507 OR2X1_LOC_64/Y AND2X1_LOC_843/a_8_24# 0.16fF
C39534 OR2X1_LOC_64/Y OR2X1_LOC_591/a_8_216# 0.05fF
C39582 OR2X1_LOC_64/Y AND2X1_LOC_727/A 0.04fF
C39606 OR2X1_LOC_64/Y OR2X1_LOC_95/Y 9.17fF
C39802 OR2X1_LOC_821/Y OR2X1_LOC_64/Y 0.04fF
C40511 OR2X1_LOC_64/Y OR2X1_LOC_71/A 0.08fF
C40789 OR2X1_LOC_70/Y OR2X1_LOC_64/Y 0.34fF
C40856 OR2X1_LOC_64/Y OR2X1_LOC_184/Y 0.04fF
C42001 OR2X1_LOC_484/Y OR2X1_LOC_64/Y 0.70fF
C42087 OR2X1_LOC_246/Y OR2X1_LOC_64/Y 0.18fF
C42382 OR2X1_LOC_64/Y OR2X1_LOC_16/A 0.14fF
C42437 OR2X1_LOC_108/Y OR2X1_LOC_64/Y 0.07fF
C42606 OR2X1_LOC_64/Y AND2X1_LOC_687/Y 0.04fF
C43291 OR2X1_LOC_64/Y AND2X1_LOC_447/Y 0.02fF
C43370 OR2X1_LOC_109/Y OR2X1_LOC_64/Y 0.13fF
C43419 OR2X1_LOC_64/Y AND2X1_LOC_729/B 0.01fF
C43720 AND2X1_LOC_593/a_8_24# OR2X1_LOC_64/Y 0.02fF
C43852 OR2X1_LOC_64/Y OR2X1_LOC_106/A 0.01fF
C43920 AND2X1_LOC_227/Y OR2X1_LOC_64/Y 0.07fF
C43945 OR2X1_LOC_64/Y OR2X1_LOC_813/Y 0.52fF
C44235 OR2X1_LOC_250/a_8_216# OR2X1_LOC_64/Y 0.01fF
C44268 OR2X1_LOC_599/A OR2X1_LOC_64/Y 0.17fF
C44575 OR2X1_LOC_40/Y OR2X1_LOC_64/Y 0.28fF
C44626 OR2X1_LOC_698/a_8_216# OR2X1_LOC_64/Y 0.07fF
C44659 AND2X1_LOC_843/Y OR2X1_LOC_64/Y 0.32fF
C44680 OR2X1_LOC_64/Y OR2X1_LOC_424/a_8_216# 0.01fF
C44711 OR2X1_LOC_320/Y OR2X1_LOC_64/Y 0.29fF
C45021 OR2X1_LOC_822/a_8_216# OR2X1_LOC_64/Y 0.18fF
C45218 OR2X1_LOC_64/Y OR2X1_LOC_615/Y 0.02fF
C45305 OR2X1_LOC_64/Y OR2X1_LOC_424/Y 0.01fF
C45390 AND2X1_LOC_707/Y OR2X1_LOC_64/Y 0.02fF
C45455 OR2X1_LOC_813/a_8_216# OR2X1_LOC_64/Y 0.01fF
C45531 OR2X1_LOC_64/Y AND2X1_LOC_841/B 0.07fF
C45957 OR2X1_LOC_64/Y OR2X1_LOC_495/Y 0.11fF
C45999 AND2X1_LOC_379/a_8_24# OR2X1_LOC_64/Y 0.01fF
C46356 AND2X1_LOC_776/a_8_24# OR2X1_LOC_64/Y 0.03fF
C46933 OR2X1_LOC_3/Y OR2X1_LOC_64/Y 0.38fF
C47756 AND2X1_LOC_99/Y OR2X1_LOC_64/Y 0.03fF
C48093 OR2X1_LOC_64/Y OR2X1_LOC_766/a_8_216# 0.03fF
C48240 OR2X1_LOC_503/A OR2X1_LOC_64/Y 0.05fF
C49444 OR2X1_LOC_516/B OR2X1_LOC_64/Y 0.02fF
C49760 OR2X1_LOC_64/Y OR2X1_LOC_321/a_8_216# 0.01fF
C49872 AND2X1_LOC_456/B OR2X1_LOC_64/Y 0.02fF
C50197 OR2X1_LOC_64/Y AND2X1_LOC_828/a_8_24# 0.01fF
C50400 OR2X1_LOC_321/Y OR2X1_LOC_64/Y 0.01fF
C50759 OR2X1_LOC_64/Y AND2X1_LOC_843/a_36_24# 0.01fF
C51582 OR2X1_LOC_380/A OR2X1_LOC_64/Y 0.88fF
C52457 OR2X1_LOC_763/Y OR2X1_LOC_64/Y 0.33fF
C52690 OR2X1_LOC_64/Y OR2X1_LOC_312/a_8_216# 0.01fF
C53576 OR2X1_LOC_64/Y OR2X1_LOC_766/a_36_216# 0.03fF
C53592 OR2X1_LOC_64/Y OR2X1_LOC_421/Y 0.10fF
C54136 AND2X1_LOC_78/a_8_24# OR2X1_LOC_64/Y 0.01fF
C54510 OR2X1_LOC_64/Y OR2X1_LOC_118/Y 0.03fF
C54556 OR2X1_LOC_64/Y OR2X1_LOC_238/Y 0.03fF
C55378 OR2X1_LOC_250/Y OR2X1_LOC_64/Y 0.16fF
C55684 OR2X1_LOC_177/Y OR2X1_LOC_64/Y 0.22fF
C55717 OR2X1_LOC_604/A OR2X1_LOC_64/Y 0.24fF
C55834 OR2X1_LOC_306/Y OR2X1_LOC_64/Y 0.02fF
C57264 OR2X1_LOC_64/Y VSS 1.27fF
C427 OR2X1_LOC_536/Y OR2X1_LOC_95/Y 0.02fF
C492 AND2X1_LOC_593/Y OR2X1_LOC_95/Y 0.03fF
C581 OR2X1_LOC_95/Y OR2X1_LOC_226/Y 0.01fF
C877 OR2X1_LOC_51/Y OR2X1_LOC_95/Y 3.67fF
C964 OR2X1_LOC_680/A OR2X1_LOC_95/Y 0.37fF
C1337 OR2X1_LOC_757/A OR2X1_LOC_95/Y 0.02fF
C1416 OR2X1_LOC_626/a_8_216# OR2X1_LOC_95/Y 0.17fF
C1751 OR2X1_LOC_95/Y AND2X1_LOC_436/Y 0.02fF
C2395 OR2X1_LOC_95/Y OR2X1_LOC_331/a_8_216# 0.06fF
C2723 OR2X1_LOC_387/Y OR2X1_LOC_95/Y 0.02fF
C3452 OR2X1_LOC_600/a_8_216# OR2X1_LOC_95/Y 0.01fF
C4785 OR2X1_LOC_74/A OR2X1_LOC_95/Y 0.16fF
C4804 OR2X1_LOC_95/Y OR2X1_LOC_261/A 0.01fF
C5074 OR2X1_LOC_95/Y OR2X1_LOC_626/Y 0.06fF
C5940 AND2X1_LOC_537/a_8_24# OR2X1_LOC_95/Y 0.01fF
C6262 OR2X1_LOC_134/Y OR2X1_LOC_95/Y 0.21fF
C6399 OR2X1_LOC_95/Y OR2X1_LOC_586/a_8_216# 0.01fF
C6711 OR2X1_LOC_106/Y OR2X1_LOC_95/Y 0.03fF
C6791 OR2X1_LOC_505/Y OR2X1_LOC_95/Y 0.03fF
C7261 OR2X1_LOC_95/Y OR2X1_LOC_597/a_8_216# 0.01fF
C7311 AND2X1_LOC_99/A OR2X1_LOC_95/Y 0.03fF
C7829 OR2X1_LOC_167/Y OR2X1_LOC_95/Y 0.01fF
C8096 AND2X1_LOC_362/B OR2X1_LOC_95/Y 0.01fF
C9086 OR2X1_LOC_420/a_8_216# OR2X1_LOC_95/Y 0.03fF
C9249 OR2X1_LOC_95/Y OR2X1_LOC_385/a_8_216# 0.39fF
C10329 OR2X1_LOC_95/Y OR2X1_LOC_67/a_8_216# 0.04fF
C10403 AND2X1_LOC_537/Y OR2X1_LOC_95/Y 0.01fF
C10675 AND2X1_LOC_549/Y OR2X1_LOC_95/Y 0.03fF
C10683 OR2X1_LOC_95/Y OR2X1_LOC_627/Y 0.02fF
C11869 OR2X1_LOC_406/Y OR2X1_LOC_95/Y 0.03fF
C12251 OR2X1_LOC_516/Y OR2X1_LOC_95/Y 0.03fF
C12594 OR2X1_LOC_95/Y OR2X1_LOC_533/A 0.07fF
C13251 OR2X1_LOC_125/a_8_216# OR2X1_LOC_95/Y 0.10fF
C13366 OR2X1_LOC_131/Y OR2X1_LOC_95/Y 0.03fF
C13652 VDD OR2X1_LOC_95/Y 1.41fF
C13766 AND2X1_LOC_389/a_8_24# OR2X1_LOC_95/Y 0.01fF
C13835 OR2X1_LOC_674/Y OR2X1_LOC_95/Y 0.01fF
C14187 OR2X1_LOC_95/Y OR2X1_LOC_248/Y 0.04fF
C14507 OR2X1_LOC_600/Y OR2X1_LOC_95/Y 0.02fF
C14557 OR2X1_LOC_95/Y OR2X1_LOC_531/a_8_216# 0.01fF
C14611 OR2X1_LOC_420/a_36_216# OR2X1_LOC_95/Y 0.03fF
C15012 OR2X1_LOC_95/Y AND2X1_LOC_464/a_8_24# 0.03fF
C16087 OR2X1_LOC_95/Y OR2X1_LOC_184/a_8_216# 0.18fF
C16525 OR2X1_LOC_45/B OR2X1_LOC_95/Y 0.56fF
C17010 OR2X1_LOC_158/A OR2X1_LOC_95/Y 3.15fF
C17066 OR2X1_LOC_103/Y OR2X1_LOC_95/Y 1.03fF
C17084 OR2X1_LOC_103/a_8_216# OR2X1_LOC_95/Y 0.01fF
C17490 OR2X1_LOC_95/Y OR2X1_LOC_586/Y 0.09fF
C17871 OR2X1_LOC_132/a_8_216# OR2X1_LOC_95/Y 0.02fF
C17963 OR2X1_LOC_117/Y OR2X1_LOC_95/Y 0.07fF
C18765 OR2X1_LOC_125/a_36_216# OR2X1_LOC_95/Y 0.03fF
C19086 OR2X1_LOC_95/Y AND2X1_LOC_227/a_8_24# 0.01fF
C19152 AND2X1_LOC_541/Y OR2X1_LOC_95/Y 0.01fF
C19181 OR2X1_LOC_107/a_8_216# OR2X1_LOC_95/Y 0.01fF
C19280 AND2X1_LOC_390/B OR2X1_LOC_95/Y 0.01fF
C19285 OR2X1_LOC_825/a_8_216# OR2X1_LOC_95/Y 0.01fF
C19694 AND2X1_LOC_840/B OR2X1_LOC_95/Y 0.12fF
C19994 OR2X1_LOC_95/Y AND2X1_LOC_464/A 0.02fF
C20137 OR2X1_LOC_420/Y OR2X1_LOC_95/Y 0.01fF
C20615 OR2X1_LOC_95/Y OR2X1_LOC_751/A 0.04fF
C21417 OR2X1_LOC_91/Y OR2X1_LOC_95/Y 0.13fF
C21458 OR2X1_LOC_527/Y OR2X1_LOC_95/Y 0.03fF
C21464 OR2X1_LOC_417/Y OR2X1_LOC_95/Y 0.03fF
C21483 OR2X1_LOC_601/a_8_216# OR2X1_LOC_95/Y 0.01fF
C22253 OR2X1_LOC_95/Y AND2X1_LOC_436/B 0.02fF
C23200 OR2X1_LOC_95/Y OR2X1_LOC_409/B 0.01fF
C23542 OR2X1_LOC_497/Y OR2X1_LOC_95/Y 0.06fF
C24357 AND2X1_LOC_319/A OR2X1_LOC_95/Y 0.02fF
C24455 AND2X1_LOC_721/A OR2X1_LOC_95/Y 0.03fF
C24483 OR2X1_LOC_95/Y OR2X1_LOC_331/Y 0.18fF
C24793 OR2X1_LOC_95/Y AND2X1_LOC_361/A 0.11fF
C25196 OR2X1_LOC_96/B OR2X1_LOC_95/Y 0.41fF
C25465 AND2X1_LOC_787/A OR2X1_LOC_95/Y 0.03fF
C25613 OR2X1_LOC_406/a_8_216# OR2X1_LOC_95/Y 0.02fF
C26314 AND2X1_LOC_729/a_8_24# OR2X1_LOC_95/Y 0.01fF
C26379 AND2X1_LOC_543/a_8_24# OR2X1_LOC_95/Y 0.01fF
C26418 OR2X1_LOC_95/Y OR2X1_LOC_619/Y 0.03fF
C27242 OR2X1_LOC_331/A OR2X1_LOC_95/Y 0.18fF
C27612 OR2X1_LOC_329/Y OR2X1_LOC_95/Y 0.01fF
C28116 AND2X1_LOC_113/a_8_24# OR2X1_LOC_95/Y 0.01fF
C28576 OR2X1_LOC_312/Y OR2X1_LOC_95/Y 0.03fF
C28735 OR2X1_LOC_95/Y OR2X1_LOC_13/B 0.12fF
C29141 OR2X1_LOC_95/Y OR2X1_LOC_533/a_8_216# 0.07fF
C29269 OR2X1_LOC_95/Y OR2X1_LOC_595/A 0.07fF
C29720 OR2X1_LOC_528/Y OR2X1_LOC_95/Y 0.16fF
C29824 AND2X1_LOC_342/Y OR2X1_LOC_95/Y 0.07fF
C30273 OR2X1_LOC_89/A OR2X1_LOC_95/Y 0.13fF
C30527 OR2X1_LOC_167/a_8_216# OR2X1_LOC_95/Y 0.01fF
C31139 OR2X1_LOC_488/Y OR2X1_LOC_95/Y 0.09fF
C31152 AND2X1_LOC_727/A OR2X1_LOC_95/Y 0.03fF
C31902 OR2X1_LOC_95/Y AND2X1_LOC_621/Y 0.03fF
C32338 OR2X1_LOC_70/Y OR2X1_LOC_95/Y 0.44fF
C32382 OR2X1_LOC_504/Y OR2X1_LOC_95/Y 0.03fF
C32415 OR2X1_LOC_184/Y OR2X1_LOC_95/Y 0.02fF
C33936 OR2X1_LOC_95/Y OR2X1_LOC_16/A 0.05fF
C33955 OR2X1_LOC_108/Y OR2X1_LOC_95/Y 0.07fF
C34098 AND2X1_LOC_687/Y OR2X1_LOC_95/Y 0.01fF
C34374 OR2X1_LOC_132/Y OR2X1_LOC_95/Y 0.07fF
C34820 OR2X1_LOC_95/Y AND2X1_LOC_447/Y 0.01fF
C34898 OR2X1_LOC_109/Y OR2X1_LOC_95/Y 0.07fF
C35350 AND2X1_LOC_227/Y OR2X1_LOC_95/Y 0.08fF
C35379 OR2X1_LOC_813/Y OR2X1_LOC_95/Y 0.03fF
C35669 OR2X1_LOC_107/Y OR2X1_LOC_95/Y 0.05fF
C35733 OR2X1_LOC_599/A OR2X1_LOC_95/Y 0.01fF
C36051 OR2X1_LOC_40/Y OR2X1_LOC_95/Y 5.63fF
C36491 OR2X1_LOC_531/Y OR2X1_LOC_95/Y 0.02fF
C36556 OR2X1_LOC_406/a_36_216# OR2X1_LOC_95/Y 0.03fF
C36629 OR2X1_LOC_95/Y OR2X1_LOC_615/Y 0.11fF
C36933 AND2X1_LOC_841/B OR2X1_LOC_95/Y 0.03fF
C37231 AND2X1_LOC_543/Y OR2X1_LOC_95/Y 0.26fF
C37291 OR2X1_LOC_95/Y OR2X1_LOC_322/Y 0.01fF
C37373 OR2X1_LOC_495/Y OR2X1_LOC_95/Y 0.48fF
C38276 OR2X1_LOC_3/Y OR2X1_LOC_95/Y 0.03fF
C38285 AND2X1_LOC_631/Y OR2X1_LOC_95/Y 0.03fF
C38684 AND2X1_LOC_113/Y OR2X1_LOC_95/Y 0.01fF
C39618 AND2X1_LOC_632/A OR2X1_LOC_95/Y 0.12fF
C39822 AND2X1_LOC_541/a_8_24# OR2X1_LOC_95/Y -0.01fF
C40270 OR2X1_LOC_96/Y OR2X1_LOC_95/Y 0.01fF
C40787 OR2X1_LOC_189/A OR2X1_LOC_95/Y 0.11fF
C41282 OR2X1_LOC_825/Y OR2X1_LOC_95/Y 0.09fF
C42195 OR2X1_LOC_95/Y OR2X1_LOC_96/a_8_216# 0.01fF
C42992 OR2X1_LOC_95/Y AND2X1_LOC_624/A 0.03fF
C44136 OR2X1_LOC_95/Y OR2X1_LOC_312/a_8_216# 0.01fF
C45610 OR2X1_LOC_95/Y OR2X1_LOC_601/Y 0.43fF
C45801 OR2X1_LOC_95/Y OR2X1_LOC_142/Y 0.12fF
C45840 OR2X1_LOC_134/a_8_216# OR2X1_LOC_95/Y 0.03fF
C46030 OR2X1_LOC_95/Y OR2X1_LOC_118/Y 0.03fF
C46064 OR2X1_LOC_95/Y OR2X1_LOC_238/Y 0.03fF
C47294 OR2X1_LOC_177/Y OR2X1_LOC_95/Y 0.03fF
C47322 OR2X1_LOC_604/A OR2X1_LOC_95/Y 1.07fF
C47325 AND2X1_LOC_758/a_8_24# OR2X1_LOC_95/Y 0.11fF
C47777 AND2X1_LOC_549/a_8_24# OR2X1_LOC_95/Y 0.15fF
C47822 OR2X1_LOC_95/Y AND2X1_LOC_447/a_8_24# 0.01fF
C48238 OR2X1_LOC_164/Y OR2X1_LOC_95/Y 0.03fF
C49908 OR2X1_LOC_674/a_8_216# OR2X1_LOC_95/Y 0.01fF
C50009 OR2X1_LOC_95/Y AND2X1_LOC_260/a_8_24# 0.14fF
C51062 AND2X1_LOC_541/a_36_24# OR2X1_LOC_95/Y 0.01fF
C51151 OR2X1_LOC_95/Y OR2X1_LOC_594/a_8_216# 0.07fF
C51663 OR2X1_LOC_617/Y OR2X1_LOC_95/Y 0.02fF
C51680 AND2X1_LOC_464/Y OR2X1_LOC_95/Y 0.01fF
C51811 OR2X1_LOC_95/Y OR2X1_LOC_536/a_8_216# 0.01fF
C52783 OR2X1_LOC_95/Y OR2X1_LOC_829/A 0.05fF
C52817 OR2X1_LOC_759/A OR2X1_LOC_95/Y 0.02fF
C53009 OR2X1_LOC_95/Y OR2X1_LOC_597/Y 0.01fF
C53208 AND2X1_LOC_361/a_8_24# OR2X1_LOC_95/Y 0.01fF
C53328 OR2X1_LOC_385/Y OR2X1_LOC_95/Y 0.51fF
C54003 OR2X1_LOC_95/Y OR2X1_LOC_368/Y 0.08fF
C54851 OR2X1_LOC_95/Y OR2X1_LOC_323/Y 0.10fF
C54978 AND2X1_LOC_729/Y OR2X1_LOC_95/Y 0.58fF
C54992 AND2X1_LOC_784/A OR2X1_LOC_95/Y 0.07fF
C55439 OR2X1_LOC_95/Y OR2X1_LOC_52/B 0.03fF
C55902 OR2X1_LOC_280/Y OR2X1_LOC_95/Y 0.13fF
C56972 OR2X1_LOC_95/Y VSS 0.79fF
C586 OR2X1_LOC_51/Y AND2X1_LOC_287/B 0.04fF
C642 AND2X1_LOC_707/a_8_24# OR2X1_LOC_51/Y 0.01fF
C680 OR2X1_LOC_51/Y OR2X1_LOC_251/a_8_216# 0.04fF
C716 OR2X1_LOC_51/Y AND2X1_LOC_843/a_8_24# 0.01fF
C837 OR2X1_LOC_51/Y AND2X1_LOC_727/A 0.02fF
C1607 OR2X1_LOC_51/Y AND2X1_LOC_621/Y 0.23fF
C2106 OR2X1_LOC_70/Y OR2X1_LOC_51/Y 0.93fF
C2128 AND2X1_LOC_333/a_8_24# OR2X1_LOC_51/Y 0.01fF
C2171 OR2X1_LOC_504/Y OR2X1_LOC_51/Y 0.04fF
C3221 OR2X1_LOC_51/Y OR2X1_LOC_584/a_8_216# 0.01fF
C3638 OR2X1_LOC_51/Y OR2X1_LOC_16/A 0.61fF
C3726 AND2X1_LOC_168/Y OR2X1_LOC_51/Y 0.01fF
C3862 OR2X1_LOC_51/Y AND2X1_LOC_687/Y -0.01fF
C4069 OR2X1_LOC_666/a_8_216# OR2X1_LOC_51/Y 0.01fF
C4457 OR2X1_LOC_51/Y AND2X1_LOC_334/Y 0.03fF
C4525 OR2X1_LOC_109/Y OR2X1_LOC_51/Y 0.07fF
C4534 OR2X1_LOC_51/Y AND2X1_LOC_448/Y 0.03fF
C4618 OR2X1_LOC_51/Y AND2X1_LOC_729/B 0.03fF
C4986 OR2X1_LOC_51/Y OR2X1_LOC_106/A 0.01fF
C5337 OR2X1_LOC_250/a_8_216# OR2X1_LOC_51/Y 0.01fF
C5382 OR2X1_LOC_599/A OR2X1_LOC_51/Y 0.02fF
C5698 OR2X1_LOC_40/Y OR2X1_LOC_51/Y 3.05fF
C5782 OR2X1_LOC_51/Y AND2X1_LOC_843/Y 0.01fF
C6090 OR2X1_LOC_176/a_8_216# OR2X1_LOC_51/Y 0.14fF
C6178 OR2X1_LOC_51/Y OR2X1_LOC_251/a_36_216# 0.02fF
C6369 OR2X1_LOC_51/Y OR2X1_LOC_615/Y 0.02fF
C6502 AND2X1_LOC_707/Y OR2X1_LOC_51/Y 0.01fF
C6958 AND2X1_LOC_543/Y OR2X1_LOC_51/Y 0.01fF
C6999 OR2X1_LOC_51/Y OR2X1_LOC_322/Y 0.01fF
C7077 OR2X1_LOC_51/Y OR2X1_LOC_495/Y 0.01fF
C8058 OR2X1_LOC_3/Y OR2X1_LOC_51/Y 0.21fF
C8721 OR2X1_LOC_51/Y OR2X1_LOC_525/a_8_216# 0.01fF
C9159 OR2X1_LOC_51/Y OR2X1_LOC_766/a_8_216# 0.01fF
C10248 OR2X1_LOC_51/Y OR2X1_LOC_7/Y 0.16fF
C10498 OR2X1_LOC_516/B OR2X1_LOC_51/Y 0.01fF
C10626 OR2X1_LOC_51/Y AND2X1_LOC_483/a_36_24# 0.01fF
C10906 AND2X1_LOC_456/B OR2X1_LOC_51/Y 0.05fF
C11733 OR2X1_LOC_494/Y OR2X1_LOC_51/Y 0.03fF
C12669 OR2X1_LOC_51/Y AND2X1_LOC_624/A 0.13fF
C12684 OR2X1_LOC_380/A OR2X1_LOC_51/Y 0.03fF
C13163 OR2X1_LOC_51/Y OR2X1_LOC_669/a_8_216# 0.01fF
C13993 OR2X1_LOC_51/Y OR2X1_LOC_670/Y 0.01fF
C14023 OR2X1_LOC_51/Y OR2X1_LOC_418/a_8_216# 0.01fF
C14037 OR2X1_LOC_48/Y OR2X1_LOC_51/Y 0.03fF
C14296 AND2X1_LOC_160/Y OR2X1_LOC_51/Y 0.07fF
C14879 OR2X1_LOC_51/Y OR2X1_LOC_253/a_8_216# 0.01fF
C15049 OR2X1_LOC_51/Y OR2X1_LOC_504/a_8_216# 0.14fF
C15078 OR2X1_LOC_51/Y OR2X1_LOC_744/a_8_216# 0.01fF
C15426 OR2X1_LOC_51/Y OR2X1_LOC_142/Y 0.02fF
C15645 OR2X1_LOC_51/Y OR2X1_LOC_238/Y 0.01fF
C16112 OR2X1_LOC_51/Y OR2X1_LOC_52/Y 0.02fF
C16438 OR2X1_LOC_250/Y OR2X1_LOC_51/Y 0.19fF
C16780 OR2X1_LOC_177/Y OR2X1_LOC_51/Y 0.03fF
C16801 OR2X1_LOC_604/A OR2X1_LOC_51/Y 1.48fF
C16894 OR2X1_LOC_51/Y OR2X1_LOC_252/a_8_216# 0.01fF
C17194 OR2X1_LOC_176/Y OR2X1_LOC_51/Y 0.04fF
C17209 OR2X1_LOC_533/Y OR2X1_LOC_51/Y 0.01fF
C17324 OR2X1_LOC_51/Y OR2X1_LOC_265/Y 0.03fF
C17491 OR2X1_LOC_51/Y OR2X1_LOC_163/A 0.05fF
C17773 OR2X1_LOC_51/Y AND2X1_LOC_155/Y 0.01fF
C18022 OR2X1_LOC_680/a_8_216# OR2X1_LOC_51/Y 0.16fF
C18499 AND2X1_LOC_338/A OR2X1_LOC_51/Y 0.01fF
C19408 OR2X1_LOC_674/a_8_216# OR2X1_LOC_51/Y 0.01fF
C20222 OR2X1_LOC_51/Y OR2X1_LOC_766/Y 0.01fF
C20368 OR2X1_LOC_51/Y OR2X1_LOC_239/a_8_216# 0.11fF
C21089 AND2X1_LOC_98/a_8_24# OR2X1_LOC_51/Y 0.02fF
C21202 OR2X1_LOC_51/Y AND2X1_LOC_848/Y 0.03fF
C21219 OR2X1_LOC_283/Y OR2X1_LOC_51/Y 0.54fF
C21572 AND2X1_LOC_160/a_8_24# OR2X1_LOC_51/Y 0.18fF
C22888 AND2X1_LOC_508/A OR2X1_LOC_51/Y 0.52fF
C24568 AND2X1_LOC_729/Y OR2X1_LOC_51/Y 0.02fF
C24594 AND2X1_LOC_784/A OR2X1_LOC_51/Y 0.07fF
C24682 OR2X1_LOC_51/Y AND2X1_LOC_639/A 0.17fF
C25016 OR2X1_LOC_51/Y OR2X1_LOC_52/B 0.70fF
C25305 OR2X1_LOC_51/Y OR2X1_LOC_584/Y 0.01fF
C25311 OR2X1_LOC_51/Y OR2X1_LOC_253/Y 0.02fF
C25340 AND2X1_LOC_161/Y OR2X1_LOC_51/Y 0.01fF
C25377 OR2X1_LOC_165/a_8_216# OR2X1_LOC_51/Y 0.13fF
C25407 OR2X1_LOC_51/Y AND2X1_LOC_286/Y 0.01fF
C25449 OR2X1_LOC_280/Y OR2X1_LOC_51/Y 0.12fF
C25728 OR2X1_LOC_485/Y OR2X1_LOC_51/Y 0.02fF
C26116 OR2X1_LOC_51/Y OR2X1_LOC_744/Y 0.01fF
C26224 OR2X1_LOC_51/Y AND2X1_LOC_593/Y 0.65fF
C26668 OR2X1_LOC_680/A OR2X1_LOC_51/Y 0.54fF
C26687 OR2X1_LOC_667/a_8_216# OR2X1_LOC_51/Y 0.01fF
C27418 OR2X1_LOC_51/Y AND2X1_LOC_436/Y 0.83fF
C27501 OR2X1_LOC_51/Y OR2X1_LOC_603/a_8_216# 0.01fF
C27506 OR2X1_LOC_145/a_8_216# OR2X1_LOC_51/Y 0.01fF
C27518 OR2X1_LOC_51/Y OR2X1_LOC_588/Y 0.03fF
C27923 OR2X1_LOC_51/Y OR2X1_LOC_252/Y 0.55fF
C27928 OR2X1_LOC_51/Y OR2X1_LOC_313/Y 0.03fF
C28128 OR2X1_LOC_51/Y OR2X1_LOC_331/a_8_216# 0.01fF
C28542 OR2X1_LOC_51/Y OR2X1_LOC_163/a_8_216# 0.07fF
C28767 OR2X1_LOC_51/Y OR2X1_LOC_511/Y 0.01fF
C29192 OR2X1_LOC_51/Y OR2X1_LOC_237/Y 0.15fF
C29549 AND2X1_LOC_391/Y OR2X1_LOC_51/Y 0.12fF
C29596 OR2X1_LOC_823/a_8_216# OR2X1_LOC_51/Y 0.01fF
C29656 OR2X1_LOC_51/Y OR2X1_LOC_669/Y 0.18fF
C30493 OR2X1_LOC_51/Y AND2X1_LOC_673/a_8_24# 0.02fF
C30507 OR2X1_LOC_51/Y OR2X1_LOC_74/A 0.37fF
C30821 AND2X1_LOC_162/a_8_24# OR2X1_LOC_51/Y 0.01fF
C30907 OR2X1_LOC_51/Y AND2X1_LOC_287/Y 0.01fF
C31308 OR2X1_LOC_51/Y AND2X1_LOC_287/a_8_24# 0.01fF
C31362 OR2X1_LOC_51/Y OR2X1_LOC_239/Y 0.16fF
C31620 AND2X1_LOC_704/a_8_24# OR2X1_LOC_51/Y 0.01fF
C31989 AND2X1_LOC_339/B OR2X1_LOC_51/Y 0.03fF
C31993 OR2X1_LOC_482/a_8_216# OR2X1_LOC_51/Y 0.15fF
C32032 OR2X1_LOC_51/Y OR2X1_LOC_816/a_8_216# 0.05fF
C33020 OR2X1_LOC_51/Y OR2X1_LOC_627/a_8_216# 0.01fF
C33352 OR2X1_LOC_697/Y OR2X1_LOC_51/Y 0.42fF
C33435 OR2X1_LOC_670/a_8_216# OR2X1_LOC_51/Y 0.01fF
C33489 OR2X1_LOC_680/Y OR2X1_LOC_51/Y 0.23fF
C34130 OR2X1_LOC_51/Y OR2X1_LOC_603/Y 0.02fF
C34249 AND2X1_LOC_303/A OR2X1_LOC_51/Y 0.09fF
C34275 OR2X1_LOC_665/Y OR2X1_LOC_51/Y 0.15fF
C34692 OR2X1_LOC_495/a_8_216# OR2X1_LOC_51/Y 0.01fF
C34827 OR2X1_LOC_51/Y OR2X1_LOC_238/a_8_216# 0.19fF
C35064 OR2X1_LOC_695/a_8_216# OR2X1_LOC_51/Y 0.01fF
C35962 OR2X1_LOC_51/Y OR2X1_LOC_418/Y 0.01fF
C36200 OR2X1_LOC_51/Y OR2X1_LOC_171/a_8_216# 0.13fF
C36246 OR2X1_LOC_51/Y OR2X1_LOC_13/Y 0.03fF
C36264 OR2X1_LOC_51/Y OR2X1_LOC_627/Y 0.01fF
C36664 OR2X1_LOC_526/Y OR2X1_LOC_51/Y 0.02fF
C37078 AND2X1_LOC_714/B OR2X1_LOC_51/Y 0.01fF
C37865 OR2X1_LOC_516/Y OR2X1_LOC_51/Y 0.03fF
C38257 OR2X1_LOC_51/Y OR2X1_LOC_533/A 0.02fF
C38814 OR2X1_LOC_51/Y OR2X1_LOC_583/a_8_216# 0.01fF
C38825 OR2X1_LOC_125/a_8_216# OR2X1_LOC_51/Y 0.01fF
C39242 VDD OR2X1_LOC_51/Y 1.94fF
C39292 OR2X1_LOC_677/Y OR2X1_LOC_51/Y 0.02fF
C39381 OR2X1_LOC_251/Y OR2X1_LOC_51/Y 0.26fF
C39498 OR2X1_LOC_51/Y OR2X1_LOC_674/Y 0.01fF
C39540 OR2X1_LOC_51/Y OR2X1_LOC_163/Y 0.03fF
C39778 OR2X1_LOC_51/Y AND2X1_LOC_834/a_8_24# 0.02fF
C39792 OR2X1_LOC_51/Y OR2X1_LOC_248/Y 0.04fF
C39817 OR2X1_LOC_666/Y OR2X1_LOC_51/Y 0.22fF
C42199 OR2X1_LOC_45/B OR2X1_LOC_51/Y 1.14fF
C42690 OR2X1_LOC_158/A OR2X1_LOC_51/Y 0.59fF
C42737 OR2X1_LOC_51/Y AND2X1_LOC_98/Y 0.01fF
C42751 OR2X1_LOC_51/Y OR2X1_LOC_594/Y 0.04fF
C43115 OR2X1_LOC_482/Y OR2X1_LOC_51/Y 1.26fF
C44244 OR2X1_LOC_51/Y OR2X1_LOC_146/Y 0.05fF
C45264 OR2X1_LOC_51/Y OR2X1_LOC_604/Y 0.01fF
C45402 OR2X1_LOC_51/Y AND2X1_LOC_840/B 0.12fF
C45680 OR2X1_LOC_51/Y AND2X1_LOC_464/A 0.03fF
C45723 OR2X1_LOC_694/Y OR2X1_LOC_51/Y 0.01fF
C47196 OR2X1_LOC_91/Y OR2X1_LOC_51/Y 0.18fF
C47223 OR2X1_LOC_51/Y AND2X1_LOC_446/a_8_24# 0.01fF
C47286 OR2X1_LOC_417/Y OR2X1_LOC_51/Y 0.06fF
C47376 OR2X1_LOC_51/Y AND2X1_LOC_483/Y 0.02fF
C47473 OR2X1_LOC_51/Y AND2X1_LOC_780/a_8_24# 0.01fF
C47477 OR2X1_LOC_51/Y OR2X1_LOC_171/Y 0.53fF
C47541 OR2X1_LOC_51/Y AND2X1_LOC_254/a_36_24# 0.01fF
C47553 AND2X1_LOC_330/a_8_24# OR2X1_LOC_51/Y 0.10fF
C48043 OR2X1_LOC_667/Y OR2X1_LOC_51/Y 0.02fF
C49018 OR2X1_LOC_51/Y OR2X1_LOC_409/B 0.03fF
C49158 OR2X1_LOC_146/a_8_216# OR2X1_LOC_51/Y 0.15fF
C49288 OR2X1_LOC_525/Y OR2X1_LOC_51/Y 0.03fF
C50180 OR2X1_LOC_51/Y AND2X1_LOC_319/A 0.44fF
C50238 OR2X1_LOC_51/Y OR2X1_LOC_52/a_8_216# 0.17fF
C50314 OR2X1_LOC_51/Y OR2X1_LOC_604/a_8_216# 0.01fF
C50357 OR2X1_LOC_51/Y AND2X1_LOC_721/A 0.08fF
C50382 OR2X1_LOC_51/Y OR2X1_LOC_331/Y 0.13fF
C51277 AND2X1_LOC_787/A OR2X1_LOC_51/Y 0.04fF
C51336 OR2X1_LOC_695/Y OR2X1_LOC_51/Y 0.01fF
C52238 OR2X1_LOC_51/Y OR2X1_LOC_619/Y 0.05fF
C52605 OR2X1_LOC_51/Y AND2X1_LOC_286/a_8_24# 0.01fF
C52707 OR2X1_LOC_51/Y OR2X1_LOC_669/A 0.04fF
C52730 OR2X1_LOC_51/Y AND2X1_LOC_454/A 0.01fF
C52865 OR2X1_LOC_51/Y OR2X1_LOC_289/Y 0.02fF
C52968 OR2X1_LOC_51/Y AND2X1_LOC_783/B 0.03fF
C53052 OR2X1_LOC_331/A OR2X1_LOC_51/Y 0.01fF
C54401 OR2X1_LOC_312/Y OR2X1_LOC_51/Y 0.03fF
C54593 OR2X1_LOC_51/Y OR2X1_LOC_13/B 0.34fF
C54989 OR2X1_LOC_51/Y OR2X1_LOC_533/a_8_216# -0.00fF
C55533 OR2X1_LOC_528/Y OR2X1_LOC_51/Y 0.03fF
C55544 OR2X1_LOC_51/Y OR2X1_LOC_583/Y 0.01fF
C55644 OR2X1_LOC_51/Y AND2X1_LOC_342/Y 0.07fF
C55679 OR2X1_LOC_51/Y AND2X1_LOC_105/a_8_24# 0.01fF
C55723 OR2X1_LOC_51/Y AND2X1_LOC_483/a_8_24# 0.14fF
C55979 OR2X1_LOC_51/Y OR2X1_LOC_765/Y 0.16fF
C56143 OR2X1_LOC_51/Y OR2X1_LOC_89/A 0.30fF
C57419 OR2X1_LOC_51/Y VSS 1.81fF
C7271 VDD OR2X1_LOC_430/Y 0.16fF
C10458 OR2X1_LOC_428/Y OR2X1_LOC_430/Y 0.19fF
C24089 OR2X1_LOC_430/Y AND2X1_LOC_451/a_8_24# 0.23fF
C26086 OR2X1_LOC_70/Y OR2X1_LOC_430/Y 0.01fF
C40738 OR2X1_LOC_604/A OR2X1_LOC_430/Y 0.02fF
C56956 OR2X1_LOC_430/Y VSS 0.07fF
C23650 OR2X1_LOC_409/Y AND2X1_LOC_460/a_8_24# 0.01fF
C32253 VDD OR2X1_LOC_409/Y 0.04fF
C34565 OR2X1_LOC_409/Y AND2X1_LOC_463/B 0.78fF
C57046 OR2X1_LOC_409/Y VSS 0.02fF
C4750 OR2X1_LOC_769/B AND2X1_LOC_31/Y 0.05fF
C8842 OR2X1_LOC_769/B OR2X1_LOC_637/a_8_216# 0.47fF
C15143 OR2X1_LOC_769/B OR2X1_LOC_769/A 0.05fF
C31548 OR2X1_LOC_769/B OR2X1_LOC_769/a_8_216# 0.03fF
C48479 OR2X1_LOC_769/B OR2X1_LOC_637/A 0.16fF
C53800 OR2X1_LOC_769/B OR2X1_LOC_771/B 0.02fF
C53917 OR2X1_LOC_769/B OR2X1_LOC_637/B 0.13fF
C58120 OR2X1_LOC_769/B VSS 0.30fF
C13040 OR2X1_LOC_635/A OR2X1_LOC_614/Y 0.02fF
C34866 OR2X1_LOC_635/A OR2X1_LOC_614/a_8_216# -0.05fF
C35727 OR2X1_LOC_635/A OR2X1_LOC_451/B 0.28fF
C53913 OR2X1_LOC_635/A OR2X1_LOC_78/A 0.01fF
C58112 OR2X1_LOC_635/A VSS 0.34fF
C22346 OR2X1_LOC_790/B AND2X1_LOC_41/Y 0.01fF
C38107 OR2X1_LOC_790/B OR2X1_LOC_790/a_8_216# 0.01fF
C49412 OR2X1_LOC_790/B OR2X1_LOC_793/A 0.80fF
C58082 OR2X1_LOC_790/B VSS 0.10fF
C569 AND2X1_LOC_47/Y AND2X1_LOC_600/a_8_24# 0.01fF
C809 AND2X1_LOC_47/Y OR2X1_LOC_342/A 0.01fF
C1705 OR2X1_LOC_614/Y AND2X1_LOC_47/Y 0.16fF
C2593 AND2X1_LOC_47/Y OR2X1_LOC_113/B 0.08fF
C2770 AND2X1_LOC_47/Y OR2X1_LOC_532/B 0.88fF
C4083 AND2X1_LOC_47/Y AND2X1_LOC_432/a_8_24# 0.01fF
C4665 VDD AND2X1_LOC_47/Y 1.73fF
C4844 AND2X1_LOC_47/Y OR2X1_LOC_845/A 0.21fF
C5494 OR2X1_LOC_676/Y AND2X1_LOC_47/Y 0.07fF
C5583 OR2X1_LOC_462/B AND2X1_LOC_47/Y 0.02fF
C6068 AND2X1_LOC_47/Y OR2X1_LOC_602/B 0.05fF
C6472 AND2X1_LOC_47/Y OR2X1_LOC_416/Y 0.08fF
C6699 AND2X1_LOC_47/Y OR2X1_LOC_115/B 0.02fF
C6843 OR2X1_LOC_840/A AND2X1_LOC_47/Y 1.25fF
C7206 AND2X1_LOC_754/a_8_24# AND2X1_LOC_47/Y 0.01fF
C7328 OR2X1_LOC_802/Y AND2X1_LOC_47/Y 0.18fF
C7751 OR2X1_LOC_160/A AND2X1_LOC_47/Y 0.14fF
C7788 AND2X1_LOC_86/B AND2X1_LOC_47/Y 0.01fF
C7795 OR2X1_LOC_624/B AND2X1_LOC_47/Y 1.06fF
C8057 OR2X1_LOC_196/Y AND2X1_LOC_47/Y 0.01fF
C8063 AND2X1_LOC_47/Y OR2X1_LOC_266/A 0.01fF
C8293 AND2X1_LOC_127/a_8_24# AND2X1_LOC_47/Y -0.00fF
C8517 OR2X1_LOC_113/a_8_216# AND2X1_LOC_47/Y 0.01fF
C9047 OR2X1_LOC_185/A AND2X1_LOC_47/Y 0.17fF
C9538 OR2X1_LOC_702/A AND2X1_LOC_47/Y 0.03fF
C10219 AND2X1_LOC_47/Y OR2X1_LOC_294/Y 0.01fF
C11166 OR2X1_LOC_643/A AND2X1_LOC_47/Y 0.03fF
C11170 AND2X1_LOC_47/Y OR2X1_LOC_778/Y 0.12fF
C11430 AND2X1_LOC_91/B AND2X1_LOC_47/Y 0.21fF
C11784 AND2X1_LOC_47/Y OR2X1_LOC_303/B 0.03fF
C11931 OR2X1_LOC_542/B AND2X1_LOC_47/Y 0.03fF
C12017 AND2X1_LOC_56/B AND2X1_LOC_47/Y 0.12fF
C12774 OR2X1_LOC_790/A AND2X1_LOC_47/Y 0.01fF
C13562 AND2X1_LOC_47/Y OR2X1_LOC_186/a_8_216# 0.05fF
C13727 OR2X1_LOC_506/A AND2X1_LOC_47/Y 0.02fF
C13730 AND2X1_LOC_47/Y AND2X1_LOC_695/a_8_24# 0.11fF
C13836 AND2X1_LOC_47/Y OR2X1_LOC_284/B 0.09fF
C14157 OR2X1_LOC_633/Y AND2X1_LOC_47/Y 7.73fF
C15336 OR2X1_LOC_235/B AND2X1_LOC_47/Y 0.10fF
C15681 AND2X1_LOC_47/Y AND2X1_LOC_295/a_8_24# 0.01fF
C15745 OR2X1_LOC_703/A AND2X1_LOC_47/Y 0.03fF
C16138 AND2X1_LOC_47/Y OR2X1_LOC_362/A 0.03fF
C16155 OR2X1_LOC_832/a_8_216# AND2X1_LOC_47/Y 0.01fF
C16430 AND2X1_LOC_47/Y OR2X1_LOC_771/B 0.03fF
C16896 AND2X1_LOC_47/Y OR2X1_LOC_593/B 0.05fF
C17384 AND2X1_LOC_47/Y AND2X1_LOC_44/Y 0.31fF
C18069 AND2X1_LOC_47/Y OR2X1_LOC_247/Y 0.02fF
C18833 AND2X1_LOC_394/a_8_24# AND2X1_LOC_47/Y 0.04fF
C19244 AND2X1_LOC_47/Y OR2X1_LOC_130/A 0.05fF
C19253 AND2X1_LOC_47/Y AND2X1_LOC_7/a_8_24# 0.01fF
C19257 AND2X1_LOC_47/Y AND2X1_LOC_292/a_8_24# 0.02fF
C19679 OR2X1_LOC_128/A AND2X1_LOC_47/Y 0.04fF
C19703 AND2X1_LOC_47/Y OR2X1_LOC_449/B 0.11fF
C19889 AND2X1_LOC_47/Y OR2X1_LOC_195/a_8_216# 0.01fF
C21276 AND2X1_LOC_47/Y OR2X1_LOC_346/A 0.01fF
C21457 AND2X1_LOC_47/Y AND2X1_LOC_51/Y 0.19fF
C21801 OR2X1_LOC_640/A AND2X1_LOC_47/Y 0.02fF
C21823 AND2X1_LOC_47/Y AND2X1_LOC_297/a_8_24# 0.02fF
C22274 OR2X1_LOC_631/B AND2X1_LOC_47/Y 0.03fF
C22592 AND2X1_LOC_524/a_8_24# AND2X1_LOC_47/Y 0.01fF
C23286 AND2X1_LOC_47/Y OR2X1_LOC_71/A 0.08fF
C23669 AND2X1_LOC_47/Y AND2X1_LOC_31/Y 1.90fF
C23974 AND2X1_LOC_47/Y OR2X1_LOC_240/A 0.01fF
C24723 OR2X1_LOC_630/Y AND2X1_LOC_47/Y 0.80fF
C24795 AND2X1_LOC_47/Y OR2X1_LOC_346/B 0.01fF
C24892 AND2X1_LOC_47/Y OR2X1_LOC_196/a_8_216# 0.01fF
C25180 OR2X1_LOC_128/B AND2X1_LOC_47/Y 0.02fF
C25841 OR2X1_LOC_308/A AND2X1_LOC_47/Y 0.01fF
C27289 AND2X1_LOC_47/Y OR2X1_LOC_347/B 0.01fF
C27294 AND2X1_LOC_47/Y OR2X1_LOC_539/Y 0.08fF
C27622 AND2X1_LOC_184/a_8_24# AND2X1_LOC_47/Y 0.02fF
C27895 AND2X1_LOC_47/Y OR2X1_LOC_777/B 0.06fF
C28035 OR2X1_LOC_545/A AND2X1_LOC_47/Y 0.01fF
C28510 OR2X1_LOC_435/B AND2X1_LOC_47/Y 0.08fF
C28965 AND2X1_LOC_132/a_8_24# AND2X1_LOC_47/Y 0.02fF
C29492 OR2X1_LOC_673/A AND2X1_LOC_47/Y 0.04fF
C29823 OR2X1_LOC_400/A AND2X1_LOC_47/Y 0.01fF
C29904 AND2X1_LOC_47/Y AND2X1_LOC_106/a_8_24# 0.09fF
C30270 AND2X1_LOC_47/Y OR2X1_LOC_647/B 0.08fF
C31073 OR2X1_LOC_318/Y AND2X1_LOC_47/Y 0.17fF
C31438 AND2X1_LOC_103/a_8_24# AND2X1_LOC_47/Y 0.10fF
C31960 OR2X1_LOC_446/Y AND2X1_LOC_47/Y 0.03fF
C32393 OR2X1_LOC_436/Y AND2X1_LOC_47/Y 0.03fF
C33525 OR2X1_LOC_151/A AND2X1_LOC_47/Y 0.57fF
C33665 OR2X1_LOC_191/B AND2X1_LOC_47/Y 0.02fF
C33932 AND2X1_LOC_47/Y AND2X1_LOC_279/a_8_24# 0.10fF
C34430 OR2X1_LOC_137/B AND2X1_LOC_47/Y 0.01fF
C35382 AND2X1_LOC_47/Y AND2X1_LOC_497/a_8_24# 0.02fF
C36148 OR2X1_LOC_151/Y AND2X1_LOC_47/Y 0.10fF
C36547 OR2X1_LOC_664/Y AND2X1_LOC_47/Y 0.03fF
C36947 AND2X1_LOC_47/Y AND2X1_LOC_601/a_8_24# 0.01fF
C37036 AND2X1_LOC_47/Y AND2X1_LOC_7/Y 0.01fF
C37264 AND2X1_LOC_47/Y OR2X1_LOC_706/a_8_216# 0.03fF
C37418 AND2X1_LOC_89/a_8_24# AND2X1_LOC_47/Y 0.01fF
C37525 AND2X1_LOC_47/Y AND2X1_LOC_280/a_8_24# 0.10fF
C38163 OR2X1_LOC_841/A AND2X1_LOC_47/Y 0.01fF
C38328 AND2X1_LOC_47/Y OR2X1_LOC_84/A 0.19fF
C38601 OR2X1_LOC_190/A AND2X1_LOC_47/Y 0.01fF
C38807 AND2X1_LOC_47/Y OR2X1_LOC_241/B 0.17fF
C39086 AND2X1_LOC_47/Y AND2X1_LOC_615/a_8_24# 0.01fF
C39423 AND2X1_LOC_47/Y AND2X1_LOC_438/a_8_24# 0.01fF
C39431 OR2X1_LOC_673/B AND2X1_LOC_47/Y 0.02fF
C39443 OR2X1_LOC_831/A AND2X1_LOC_47/Y 0.01fF
C39501 OR2X1_LOC_335/Y AND2X1_LOC_47/Y 0.03fF
C40342 OR2X1_LOC_610/a_8_216# AND2X1_LOC_47/Y 0.05fF
C40387 OR2X1_LOC_810/A AND2X1_LOC_47/Y 4.20fF
C40390 OR2X1_LOC_307/a_8_216# AND2X1_LOC_47/Y 0.01fF
C40697 OR2X1_LOC_715/B AND2X1_LOC_47/Y 0.14fF
C40926 AND2X1_LOC_47/Y OR2X1_LOC_398/Y 0.01fF
C41693 OR2X1_LOC_687/Y AND2X1_LOC_47/Y 0.06fF
C41695 AND2X1_LOC_47/Y OR2X1_LOC_781/A 0.15fF
C41699 AND2X1_LOC_399/a_8_24# AND2X1_LOC_47/Y 0.02fF
C41702 AND2X1_LOC_152/a_8_24# AND2X1_LOC_47/Y 0.02fF
C41901 AND2X1_LOC_47/Y OR2X1_LOC_199/B 0.01fF
C42418 AND2X1_LOC_91/a_8_24# AND2X1_LOC_47/Y 0.01fF
C42495 AND2X1_LOC_47/Y OR2X1_LOC_78/A 2.34fF
C42572 AND2X1_LOC_47/Y OR2X1_LOC_602/A 0.01fF
C42864 AND2X1_LOC_47/Y OR2X1_LOC_706/a_36_216# 0.02fF
C43006 OR2X1_LOC_97/B AND2X1_LOC_47/Y 0.18fF
C43363 OR2X1_LOC_501/B AND2X1_LOC_47/Y 0.14fF
C43389 OR2X1_LOC_147/B AND2X1_LOC_47/Y 0.06fF
C43487 OR2X1_LOC_545/B AND2X1_LOC_47/Y 0.01fF
C43554 AND2X1_LOC_47/Y OR2X1_LOC_318/B 0.03fF
C43769 OR2X1_LOC_114/B AND2X1_LOC_47/Y 3.29fF
C43810 OR2X1_LOC_538/A AND2X1_LOC_47/Y 0.03fF
C43893 AND2X1_LOC_47/Y AND2X1_LOC_79/Y 0.03fF
C44683 AND2X1_LOC_47/Y OR2X1_LOC_623/B 0.01fF
C44787 AND2X1_LOC_47/Y OR2X1_LOC_544/A 0.01fF
C45877 AND2X1_LOC_47/Y AND2X1_LOC_248/a_8_24# 0.04fF
C46812 OR2X1_LOC_186/Y AND2X1_LOC_47/Y 0.03fF
C46997 OR2X1_LOC_196/B AND2X1_LOC_47/Y 0.07fF
C47427 OR2X1_LOC_574/A AND2X1_LOC_47/Y 0.01fF
C48572 AND2X1_LOC_47/Y OR2X1_LOC_549/A 1.31fF
C48616 OR2X1_LOC_113/Y AND2X1_LOC_47/Y 0.52fF
C49042 OR2X1_LOC_499/B AND2X1_LOC_47/Y 0.03fF
C50402 OR2X1_LOC_673/Y AND2X1_LOC_47/Y 0.20fF
C50422 OR2X1_LOC_195/A AND2X1_LOC_47/Y 0.01fF
C52273 AND2X1_LOC_47/Y AND2X1_LOC_235/a_8_24# 0.03fF
C52679 AND2X1_LOC_47/Y OR2X1_LOC_844/B 0.07fF
C52921 OR2X1_LOC_403/B AND2X1_LOC_47/Y 0.01fF
C53612 OR2X1_LOC_97/A AND2X1_LOC_47/Y 0.12fF
C53708 OR2X1_LOC_541/A AND2X1_LOC_47/Y 0.03fF
C54614 AND2X1_LOC_47/Y OR2X1_LOC_99/B 0.14fF
C54980 OR2X1_LOC_154/A AND2X1_LOC_47/Y 0.48fF
C55093 AND2X1_LOC_47/Y OR2X1_LOC_99/A 0.03fF
C55517 AND2X1_LOC_47/Y AND2X1_LOC_813/a_8_24# 0.02fF
C55819 OR2X1_LOC_634/A AND2X1_LOC_47/Y 0.02fF
C56180 AND2X1_LOC_47/Y OR2X1_LOC_633/A 0.54fF
C57124 AND2X1_LOC_47/Y VSS 0.78fF
C215 OR2X1_LOC_668/a_8_216# AND2X1_LOC_44/Y 0.01fF
C518 AND2X1_LOC_44/Y OR2X1_LOC_844/B 0.01fF
C587 OR2X1_LOC_389/A AND2X1_LOC_44/Y 0.03fF
C718 AND2X1_LOC_528/a_36_24# AND2X1_LOC_44/Y 0.01fF
C951 OR2X1_LOC_532/a_8_216# AND2X1_LOC_44/Y 0.02fF
C1108 OR2X1_LOC_194/B AND2X1_LOC_44/Y 0.01fF
C1443 OR2X1_LOC_97/A AND2X1_LOC_44/Y 0.03fF
C1506 AND2X1_LOC_744/a_8_24# AND2X1_LOC_44/Y 0.01fF
C1866 AND2X1_LOC_44/Y OR2X1_LOC_713/A 0.44fF
C2426 OR2X1_LOC_639/B AND2X1_LOC_44/Y 0.11fF
C2446 OR2X1_LOC_720/A AND2X1_LOC_44/Y 0.06fF
C2483 OR2X1_LOC_333/B AND2X1_LOC_44/Y 0.09fF
C2509 OR2X1_LOC_99/B AND2X1_LOC_44/Y 0.01fF
C2867 OR2X1_LOC_154/A AND2X1_LOC_44/Y 0.37fF
C3643 OR2X1_LOC_634/A AND2X1_LOC_44/Y 0.09fF
C3992 OR2X1_LOC_267/Y AND2X1_LOC_44/Y 0.03fF
C4091 OR2X1_LOC_520/Y AND2X1_LOC_44/Y 0.03fF
C4176 AND2X1_LOC_107/a_8_24# AND2X1_LOC_44/Y 0.01fF
C4808 AND2X1_LOC_44/Y OR2X1_LOC_342/A 0.01fF
C5224 OR2X1_LOC_124/B AND2X1_LOC_44/Y 0.28fF
C5626 AND2X1_LOC_44/Y OR2X1_LOC_779/A 0.06fF
C6721 OR2X1_LOC_532/B AND2X1_LOC_44/Y 1.17fF
C7444 OR2X1_LOC_114/a_8_216# AND2X1_LOC_44/Y 0.01fF
C7845 OR2X1_LOC_710/B AND2X1_LOC_44/Y 0.13fF
C8733 VDD AND2X1_LOC_44/Y 1.80fF
C9511 AND2X1_LOC_44/Y OR2X1_LOC_523/A 0.01fF
C9579 OR2X1_LOC_676/Y AND2X1_LOC_44/Y 0.09fF
C9592 OR2X1_LOC_834/A AND2X1_LOC_44/Y 0.01fF
C9665 OR2X1_LOC_462/B AND2X1_LOC_44/Y 0.01fF
C10788 OR2X1_LOC_115/B AND2X1_LOC_44/Y 0.05fF
C10861 OR2X1_LOC_840/A AND2X1_LOC_44/Y 0.01fF
C11752 OR2X1_LOC_160/A AND2X1_LOC_44/Y 0.69fF
C12006 OR2X1_LOC_532/Y AND2X1_LOC_44/Y 0.07fF
C12283 AND2X1_LOC_127/a_8_24# AND2X1_LOC_44/Y 0.01fF
C13012 OR2X1_LOC_708/Y AND2X1_LOC_44/Y 0.01fF
C13042 OR2X1_LOC_185/A AND2X1_LOC_44/Y 0.17fF
C13803 AND2X1_LOC_262/a_8_24# AND2X1_LOC_44/Y 0.01fF
C13946 AND2X1_LOC_481/a_8_24# AND2X1_LOC_44/Y 0.03fF
C14229 OR2X1_LOC_294/Y AND2X1_LOC_44/Y 0.01fF
C14241 OR2X1_LOC_641/A AND2X1_LOC_44/Y 0.03fF
C14336 OR2X1_LOC_114/Y AND2X1_LOC_44/Y 0.01fF
C15159 OR2X1_LOC_643/A AND2X1_LOC_44/Y 0.03fF
C15168 OR2X1_LOC_778/Y AND2X1_LOC_44/Y 0.36fF
C15230 OR2X1_LOC_113/A AND2X1_LOC_44/Y 0.01fF
C15417 AND2X1_LOC_91/B AND2X1_LOC_44/Y 0.22fF
C15512 OR2X1_LOC_308/a_8_216# AND2X1_LOC_44/Y 0.01fF
C15896 OR2X1_LOC_542/B AND2X1_LOC_44/Y 0.03fF
C15981 AND2X1_LOC_56/B AND2X1_LOC_44/Y 0.47fF
C16873 OR2X1_LOC_389/B AND2X1_LOC_44/Y 0.09fF
C17564 AND2X1_LOC_521/a_8_24# AND2X1_LOC_44/Y 0.01fF
C17776 OR2X1_LOC_780/A AND2X1_LOC_44/Y 0.09fF
C17811 AND2X1_LOC_44/Y OR2X1_LOC_284/B 0.01fF
C18107 OR2X1_LOC_633/Y AND2X1_LOC_44/Y 0.03fF
C18137 OR2X1_LOC_99/Y AND2X1_LOC_44/Y 0.03fF
C18394 AND2X1_LOC_44/Y AND2X1_LOC_41/Y 0.02fF
C19360 OR2X1_LOC_235/B AND2X1_LOC_44/Y 0.09fF
C19739 AND2X1_LOC_295/a_8_24# AND2X1_LOC_44/Y 0.01fF
C20192 OR2X1_LOC_362/A AND2X1_LOC_44/Y 0.51fF
C20539 OR2X1_LOC_771/B AND2X1_LOC_44/Y 0.03fF
C20551 AND2X1_LOC_44/Y OR2X1_LOC_209/A 0.28fF
C20643 OR2X1_LOC_678/a_8_216# AND2X1_LOC_44/Y 0.01fF
C21677 OR2X1_LOC_720/B AND2X1_LOC_44/Y -0.00fF
C22297 AND2X1_LOC_44/Y AND2X1_LOC_258/a_8_24# 0.03fF
C22313 AND2X1_LOC_44/Y OR2X1_LOC_708/a_8_216# 0.01fF
C22623 AND2X1_LOC_485/a_8_24# AND2X1_LOC_44/Y 0.04fF
C22795 OR2X1_LOC_307/A AND2X1_LOC_44/Y 0.01fF
C23174 OR2X1_LOC_523/B AND2X1_LOC_44/Y 0.03fF
C23281 OR2X1_LOC_130/A AND2X1_LOC_44/Y 0.56fF
C23297 AND2X1_LOC_292/a_8_24# AND2X1_LOC_44/Y 0.01fF
C23449 AND2X1_LOC_44/Y AND2X1_LOC_39/Y 0.03fF
C23682 OR2X1_LOC_128/A AND2X1_LOC_44/Y 0.01fF
C23717 OR2X1_LOC_449/B AND2X1_LOC_44/Y 0.03fF
C24835 AND2X1_LOC_44/Y OR2X1_LOC_389/a_8_216# 0.02fF
C24844 OR2X1_LOC_786/A AND2X1_LOC_44/Y 0.04fF
C25036 OR2X1_LOC_447/Y AND2X1_LOC_44/Y 0.03fF
C25251 OR2X1_LOC_346/A AND2X1_LOC_44/Y 0.01fF
C25403 AND2X1_LOC_51/Y AND2X1_LOC_44/Y 0.23fF
C25739 AND2X1_LOC_297/a_8_24# AND2X1_LOC_44/Y 0.01fF
C27277 AND2X1_LOC_44/Y OR2X1_LOC_71/A 0.85fF
C27467 AND2X1_LOC_701/a_8_24# AND2X1_LOC_44/Y 0.01fF
C27656 AND2X1_LOC_31/Y AND2X1_LOC_44/Y 4.26fF
C27898 OR2X1_LOC_240/A AND2X1_LOC_44/Y 0.08fF
C27903 OR2X1_LOC_633/B AND2X1_LOC_44/Y 0.05fF
C28079 AND2X1_LOC_44/Y OR2X1_LOC_608/Y 0.07fF
C28578 AND2X1_LOC_44/Y OR2X1_LOC_333/a_8_216# 0.03fF
C28732 OR2X1_LOC_346/B AND2X1_LOC_44/Y 0.01fF
C28758 AND2X1_LOC_122/a_8_24# AND2X1_LOC_44/Y 0.04fF
C29187 OR2X1_LOC_636/B AND2X1_LOC_44/Y 0.19fF
C29440 AND2X1_LOC_522/a_8_24# AND2X1_LOC_44/Y 0.01fF
C30048 AND2X1_LOC_117/a_8_24# AND2X1_LOC_44/Y 0.01fF
C31245 OR2X1_LOC_347/B AND2X1_LOC_44/Y 0.01fF
C31266 OR2X1_LOC_779/a_8_216# AND2X1_LOC_44/Y 0.01fF
C31599 AND2X1_LOC_184/a_8_24# AND2X1_LOC_44/Y 0.01fF
C31619 OR2X1_LOC_678/Y AND2X1_LOC_44/Y 0.01fF
C31899 AND2X1_LOC_44/Y OR2X1_LOC_777/B 0.05fF
C32111 AND2X1_LOC_13/a_8_24# AND2X1_LOC_44/Y 0.02fF
C33236 AND2X1_LOC_44/Y OR2X1_LOC_259/A 0.01fF
C33562 OR2X1_LOC_705/B AND2X1_LOC_44/Y 0.41fF
C33577 AND2X1_LOC_44/Y AND2X1_LOC_609/a_8_24# 0.04fF
C34644 AND2X1_LOC_528/a_8_24# AND2X1_LOC_44/Y 0.03fF
C35085 OR2X1_LOC_296/Y AND2X1_LOC_44/Y 0.05fF
C35514 OR2X1_LOC_123/B AND2X1_LOC_44/Y 0.05fF
C35559 AND2X1_LOC_825/a_8_24# AND2X1_LOC_44/Y -0.00fF
C36000 OR2X1_LOC_446/Y AND2X1_LOC_44/Y 0.28fF
C36235 AND2X1_LOC_320/a_8_24# AND2X1_LOC_44/Y 0.01fF
C36359 OR2X1_LOC_97/a_8_216# AND2X1_LOC_44/Y 0.01fF
C37475 OR2X1_LOC_151/A AND2X1_LOC_44/Y 0.14fF
C37867 AND2X1_LOC_44/Y AND2X1_LOC_279/a_8_24# 0.01fF
C39471 AND2X1_LOC_497/a_8_24# AND2X1_LOC_44/Y 0.01fF
C39584 AND2X1_LOC_44/Y OR2X1_LOC_333/a_36_216# 0.02fF
C39957 AND2X1_LOC_44/Y OR2X1_LOC_308/Y 0.11fF
C40541 OR2X1_LOC_664/Y AND2X1_LOC_44/Y 0.03fF
C41083 AND2X1_LOC_7/Y AND2X1_LOC_44/Y 0.02fF
C41286 AND2X1_LOC_44/Y OR2X1_LOC_706/a_8_216# 0.01fF
C41789 OR2X1_LOC_324/B AND2X1_LOC_44/Y 0.21fF
C41819 AND2X1_LOC_142/a_8_24# AND2X1_LOC_44/Y 0.02fF
C41855 OR2X1_LOC_668/Y AND2X1_LOC_44/Y 0.01fF
C42664 OR2X1_LOC_190/A AND2X1_LOC_44/Y 0.01fF
C43216 OR2X1_LOC_193/A AND2X1_LOC_44/Y 0.03fF
C43888 OR2X1_LOC_710/A AND2X1_LOC_44/Y 0.01fF
C43982 AND2X1_LOC_39/a_8_24# AND2X1_LOC_44/Y 0.03fF
C44330 AND2X1_LOC_416/a_8_24# AND2X1_LOC_44/Y 0.01fF
C44471 OR2X1_LOC_810/A AND2X1_LOC_44/Y 0.05fF
C44666 AND2X1_LOC_44/Y AND2X1_LOC_609/a_36_24# 0.01fF
C44798 OR2X1_LOC_784/B AND2X1_LOC_44/Y 0.11fF
C44904 AND2X1_LOC_81/a_8_24# AND2X1_LOC_44/Y 0.01fF
C45096 AND2X1_LOC_44/Y OR2X1_LOC_398/Y 0.33fF
C45302 OR2X1_LOC_656/B AND2X1_LOC_44/Y 0.03fF
C45337 OR2X1_LOC_793/A AND2X1_LOC_44/Y 0.07fF
C45412 AND2X1_LOC_45/a_8_24# AND2X1_LOC_44/Y 0.01fF
C45758 OR2X1_LOC_687/Y AND2X1_LOC_44/Y 0.03fF
C45798 OR2X1_LOC_620/B AND2X1_LOC_44/Y 0.23fF
C46590 OR2X1_LOC_78/A AND2X1_LOC_44/Y 1.53fF
C47137 OR2X1_LOC_97/B AND2X1_LOC_44/Y 0.21fF
C47515 OR2X1_LOC_501/B AND2X1_LOC_44/Y 0.18fF
C47539 OR2X1_LOC_147/B AND2X1_LOC_44/Y 0.09fF
C47576 AND2X1_LOC_669/a_8_24# AND2X1_LOC_44/Y 0.01fF
C47892 OR2X1_LOC_121/Y AND2X1_LOC_44/Y 0.01fF
C47914 OR2X1_LOC_114/B AND2X1_LOC_44/Y 0.01fF
C48794 OR2X1_LOC_623/B AND2X1_LOC_44/Y 0.03fF
C49670 AND2X1_LOC_321/a_8_24# AND2X1_LOC_44/Y 0.02fF
C50012 AND2X1_LOC_44/Y AND2X1_LOC_248/a_8_24# 0.01fF
C50562 OR2X1_LOC_84/B AND2X1_LOC_44/Y 0.07fF
C50864 OR2X1_LOC_186/Y AND2X1_LOC_44/Y 0.02fF
C51033 OR2X1_LOC_196/B AND2X1_LOC_44/Y 0.04fF
C51770 AND2X1_LOC_16/a_8_24# AND2X1_LOC_44/Y -0.06fF
C52154 OR2X1_LOC_448/a_8_216# AND2X1_LOC_44/Y 0.01fF
C52533 AND2X1_LOC_44/Y OR2X1_LOC_549/A 0.18fF
C53130 OR2X1_LOC_486/B AND2X1_LOC_44/Y 0.16fF
C53264 AND2X1_LOC_44/Y OR2X1_LOC_348/B 0.03fF
C54036 OR2X1_LOC_779/Y AND2X1_LOC_44/Y 0.01fF
C54042 AND2X1_LOC_44/Y OR2X1_LOC_330/a_8_216# 0.05fF
C54301 OR2X1_LOC_673/Y AND2X1_LOC_44/Y 0.02fF
C54974 AND2X1_LOC_44/Y OR2X1_LOC_712/B 0.06fF
C55022 OR2X1_LOC_139/A AND2X1_LOC_44/Y 0.07fF
C55111 OR2X1_LOC_324/A AND2X1_LOC_44/Y 0.04fF
C55817 AND2X1_LOC_44/Y OR2X1_LOC_259/B 0.04fF
C55976 OR2X1_LOC_834/a_8_216# AND2X1_LOC_44/Y 0.01fF
C56456 AND2X1_LOC_44/Y VSS 0.85fF
C122 OR2X1_LOC_448/Y AND2X1_LOC_31/Y 0.01fF
C876 AND2X1_LOC_31/Y OR2X1_LOC_338/A 0.02fF
C918 OR2X1_LOC_186/Y AND2X1_LOC_31/Y 0.11fF
C1084 OR2X1_LOC_196/B AND2X1_LOC_31/Y 0.72fF
C1131 OR2X1_LOC_112/B AND2X1_LOC_31/Y 0.06fF
C1481 OR2X1_LOC_574/A AND2X1_LOC_31/Y 0.06fF
C2294 OR2X1_LOC_448/a_8_216# AND2X1_LOC_31/Y 0.01fF
C2563 AND2X1_LOC_31/Y OR2X1_LOC_515/Y 0.34fF
C4099 OR2X1_LOC_779/Y AND2X1_LOC_31/Y 0.01fF
C4348 AND2X1_LOC_316/a_8_24# AND2X1_LOC_31/Y 0.01fF
C4755 AND2X1_LOC_583/a_8_24# AND2X1_LOC_31/Y 0.01fF
C5022 AND2X1_LOC_31/Y OR2X1_LOC_712/B 0.03fF
C5098 OR2X1_LOC_139/A AND2X1_LOC_31/Y 0.03fF
C5165 OR2X1_LOC_637/Y AND2X1_LOC_31/Y 0.02fF
C6051 AND2X1_LOC_315/a_8_24# AND2X1_LOC_31/Y 0.01fF
C7698 OR2X1_LOC_97/A AND2X1_LOC_31/Y 0.10fF
C7769 OR2X1_LOC_541/A AND2X1_LOC_31/Y 0.01fF
C7789 AND2X1_LOC_31/Y OR2X1_LOC_475/B 0.03fF
C8173 AND2X1_LOC_31/Y OR2X1_LOC_713/A 0.03fF
C8702 AND2X1_LOC_74/a_8_24# AND2X1_LOC_31/Y 0.01fF
C8711 OR2X1_LOC_639/B AND2X1_LOC_31/Y 0.13fF
C9124 OR2X1_LOC_154/A AND2X1_LOC_31/Y 0.58fF
C10398 OR2X1_LOC_520/Y AND2X1_LOC_31/Y 0.01fF
C10869 AND2X1_LOC_600/a_8_24# AND2X1_LOC_31/Y 0.01fF
C11270 AND2X1_LOC_677/a_8_24# AND2X1_LOC_31/Y 0.01fF
C11273 OR2X1_LOC_227/a_8_216# AND2X1_LOC_31/Y 0.01fF
C11944 AND2X1_LOC_31/Y OR2X1_LOC_779/A 0.01fF
C11965 OR2X1_LOC_614/Y AND2X1_LOC_31/Y 0.01fF
C13029 OR2X1_LOC_532/B AND2X1_LOC_31/Y 7.61fF
C14112 AND2X1_LOC_31/Y AND2X1_LOC_224/a_8_24# 0.01fF
C14177 AND2X1_LOC_31/Y OR2X1_LOC_778/a_8_216# 0.01fF
C14209 OR2X1_LOC_76/B AND2X1_LOC_31/Y 0.01fF
C14374 AND2X1_LOC_31/Y OR2X1_LOC_552/A 0.13fF
C14393 AND2X1_LOC_31/Y AND2X1_LOC_432/a_8_24# 0.01fF
C14988 AND2X1_LOC_31/Y OR2X1_LOC_302/A 0.14fF
C14999 VDD AND2X1_LOC_31/Y 1.48fF
C15395 OR2X1_LOC_334/B AND2X1_LOC_31/Y 0.02fF
C15791 OR2X1_LOC_676/Y AND2X1_LOC_31/Y 0.07fF
C15802 OR2X1_LOC_834/A AND2X1_LOC_31/Y 0.01fF
C16347 OR2X1_LOC_602/B AND2X1_LOC_31/Y 0.05fF
C17135 OR2X1_LOC_840/A AND2X1_LOC_31/Y 0.03fF
C17563 OR2X1_LOC_802/Y AND2X1_LOC_31/Y 0.02fF
C17993 OR2X1_LOC_160/A AND2X1_LOC_31/Y 5.25fF
C19265 AND2X1_LOC_31/Y OR2X1_LOC_708/Y 0.01fF
C19290 OR2X1_LOC_185/A AND2X1_LOC_31/Y 0.39fF
C19343 OR2X1_LOC_435/Y AND2X1_LOC_31/Y 0.14fF
C19774 OR2X1_LOC_702/A AND2X1_LOC_31/Y 0.05fF
C20514 AND2X1_LOC_31/Y OR2X1_LOC_641/A 0.03fF
C20586 OR2X1_LOC_379/Y AND2X1_LOC_31/Y 0.03fF
C21437 OR2X1_LOC_637/A AND2X1_LOC_31/Y 0.06fF
C21488 OR2X1_LOC_643/A AND2X1_LOC_31/Y 0.03fF
C21492 OR2X1_LOC_778/Y AND2X1_LOC_31/Y 0.09fF
C21760 AND2X1_LOC_91/B AND2X1_LOC_31/Y 0.16fF
C21851 OR2X1_LOC_638/a_8_216# AND2X1_LOC_31/Y 0.01fF
C22326 AND2X1_LOC_56/B AND2X1_LOC_31/Y 0.11fF
C22712 AND2X1_LOC_31/Y OR2X1_LOC_787/B 0.29fF
C23169 OR2X1_LOC_457/a_8_216# AND2X1_LOC_31/Y 0.05fF
C23871 AND2X1_LOC_31/Y OR2X1_LOC_186/a_8_216# 0.01fF
C23899 AND2X1_LOC_31/Y OR2X1_LOC_34/A 0.06fF
C23997 OR2X1_LOC_506/A AND2X1_LOC_31/Y 0.04fF
C24117 AND2X1_LOC_31/Y OR2X1_LOC_227/Y 0.09fF
C25133 AND2X1_LOC_31/Y OR2X1_LOC_227/B 0.04fF
C26034 OR2X1_LOC_703/A AND2X1_LOC_31/Y 0.03fF
C26415 OR2X1_LOC_832/a_8_216# AND2X1_LOC_31/Y 0.01fF
C26730 AND2X1_LOC_31/Y OR2X1_LOC_771/B 0.13fF
C26757 AND2X1_LOC_31/Y OR2X1_LOC_776/A 1.82fF
C27190 AND2X1_LOC_31/Y OR2X1_LOC_593/B 0.02fF
C28233 AND2X1_LOC_69/Y AND2X1_LOC_31/Y 0.01fF
C28506 AND2X1_LOC_31/Y OR2X1_LOC_708/a_8_216# 0.01fF
C28952 AND2X1_LOC_31/Y OR2X1_LOC_307/A 0.01fF
C29090 AND2X1_LOC_69/a_8_24# AND2X1_LOC_31/Y 0.01fF
C29165 AND2X1_LOC_31/Y AND2X1_LOC_428/a_8_24# 0.01fF
C29412 AND2X1_LOC_65/a_8_24# AND2X1_LOC_31/Y 0.01fF
C29422 OR2X1_LOC_231/A AND2X1_LOC_31/Y 0.01fF
C29453 OR2X1_LOC_130/A AND2X1_LOC_31/Y 0.06fF
C29892 AND2X1_LOC_31/Y OR2X1_LOC_449/B 0.09fF
C29908 OR2X1_LOC_636/A AND2X1_LOC_31/Y 0.01fF
C30753 AND2X1_LOC_674/a_8_24# AND2X1_LOC_31/Y 0.01fF
C31230 OR2X1_LOC_447/Y AND2X1_LOC_31/Y 0.03fF
C31614 AND2X1_LOC_31/Y AND2X1_LOC_51/Y 1.85fF
C33709 AND2X1_LOC_701/a_8_24# AND2X1_LOC_31/Y 0.01fF
C33770 OR2X1_LOC_614/a_8_216# AND2X1_LOC_31/Y 0.01fF
C34103 OR2X1_LOC_809/a_8_216# AND2X1_LOC_31/Y 0.06fF
C34642 AND2X1_LOC_31/Y OR2X1_LOC_451/B 0.04fF
C35358 OR2X1_LOC_636/B AND2X1_LOC_31/Y 0.35fF
C36063 OR2X1_LOC_308/A AND2X1_LOC_31/Y 0.01fF
C36237 OR2X1_LOC_675/A AND2X1_LOC_31/Y 0.01fF
C36599 AND2X1_LOC_584/a_8_24# AND2X1_LOC_31/Y 0.01fF
C37028 AND2X1_LOC_31/Y AND2X1_LOC_298/a_8_24# 0.10fF
C37398 OR2X1_LOC_832/a_36_216# AND2X1_LOC_31/Y 0.02fF
C37461 AND2X1_LOC_31/Y OR2X1_LOC_539/Y 0.07fF
C37472 AND2X1_LOC_31/Y OR2X1_LOC_779/a_8_216# 0.01fF
C37824 OR2X1_LOC_678/Y AND2X1_LOC_31/Y 0.13fF
C37842 OR2X1_LOC_637/a_8_216# AND2X1_LOC_31/Y 0.06fF
C38086 AND2X1_LOC_31/Y OR2X1_LOC_777/B 0.12fF
C38705 OR2X1_LOC_435/B AND2X1_LOC_31/Y 0.01fF
C39217 AND2X1_LOC_67/Y AND2X1_LOC_31/Y 0.02fF
C39934 AND2X1_LOC_31/Y OR2X1_LOC_777/a_8_216# 0.01fF
C39985 AND2X1_LOC_31/Y AND2X1_LOC_230/a_8_24# 0.01fF
C40391 OR2X1_LOC_201/A AND2X1_LOC_31/Y 0.01fF
C41268 OR2X1_LOC_318/Y AND2X1_LOC_31/Y 0.03fF
C42616 OR2X1_LOC_635/a_8_216# AND2X1_LOC_31/Y 0.01fF
C42684 OR2X1_LOC_76/A AND2X1_LOC_31/Y 0.03fF
C42721 OR2X1_LOC_436/Y AND2X1_LOC_31/Y 0.03fF
C43818 OR2X1_LOC_318/A AND2X1_LOC_31/Y 0.01fF
C43834 OR2X1_LOC_151/A AND2X1_LOC_31/Y 0.36fF
C43891 OR2X1_LOC_651/B AND2X1_LOC_31/Y 0.06fF
C46203 AND2X1_LOC_109/a_8_24# AND2X1_LOC_31/Y 0.06fF
C47456 AND2X1_LOC_601/a_8_24# AND2X1_LOC_31/Y 0.01fF
C48359 AND2X1_LOC_822/a_8_24# AND2X1_LOC_31/Y 0.03fF
C48632 AND2X1_LOC_229/a_8_24# AND2X1_LOC_31/Y 0.01fF
C48676 OR2X1_LOC_841/A AND2X1_LOC_31/Y 0.07fF
C48686 AND2X1_LOC_311/a_8_24# AND2X1_LOC_31/Y 0.01fF
C49188 OR2X1_LOC_473/Y AND2X1_LOC_31/Y 0.02fF
C49565 AND2X1_LOC_31/Y AND2X1_LOC_615/a_8_24# 0.03fF
C50302 OR2X1_LOC_710/A AND2X1_LOC_31/Y 0.01fF
C50884 OR2X1_LOC_810/A AND2X1_LOC_31/Y 0.06fF
C50885 OR2X1_LOC_307/a_8_216# AND2X1_LOC_31/Y 0.01fF
C51169 OR2X1_LOC_715/B AND2X1_LOC_31/Y 3.89fF
C51184 AND2X1_LOC_31/Y OR2X1_LOC_543/A 0.03fF
C51187 AND2X1_LOC_31/Y OR2X1_LOC_784/B 0.02fF
C51668 OR2X1_LOC_656/B AND2X1_LOC_31/Y 0.02fF
C52085 OR2X1_LOC_687/Y AND2X1_LOC_31/Y 0.06fF
C52529 OR2X1_LOC_835/B AND2X1_LOC_31/Y 0.07fF
C52907 AND2X1_LOC_31/Y OR2X1_LOC_78/A 2.41fF
C52955 OR2X1_LOC_602/A AND2X1_LOC_31/Y 0.01fF
C53788 OR2X1_LOC_147/B AND2X1_LOC_31/Y 0.05fF
C53795 AND2X1_LOC_517/a_8_24# AND2X1_LOC_31/Y 0.11fF
C53931 AND2X1_LOC_31/Y OR2X1_LOC_318/B 0.22fF
C54089 OR2X1_LOC_231/B AND2X1_LOC_31/Y 0.01fF
C54150 OR2X1_LOC_538/A AND2X1_LOC_31/Y 0.20fF
C54197 OR2X1_LOC_841/B AND2X1_LOC_31/Y 0.03fF
C55006 AND2X1_LOC_31/Y OR2X1_LOC_623/B 0.54fF
C55931 AND2X1_LOC_32/a_8_24# AND2X1_LOC_31/Y 0.12fF
C56838 AND2X1_LOC_31/Y VSS 0.61fF
C225 AND2X1_LOC_51/Y OR2X1_LOC_515/Y 0.65fF
C347 AND2X1_LOC_51/Y OR2X1_LOC_549/A 0.07fF
C996 AND2X1_LOC_51/Y OR2X1_LOC_846/A 0.01fF
C1790 AND2X1_LOC_823/a_8_24# AND2X1_LOC_51/Y 0.01fF
C1879 AND2X1_LOC_51/Y OR2X1_LOC_330/a_8_216# 0.09fF
C2166 AND2X1_LOC_316/a_8_24# AND2X1_LOC_51/Y 0.01fF
C2600 AND2X1_LOC_583/a_8_24# AND2X1_LOC_51/Y 0.01fF
C2715 AND2X1_LOC_27/a_8_24# AND2X1_LOC_51/Y 0.01fF
C2927 OR2X1_LOC_139/A AND2X1_LOC_51/Y 0.01fF
C3248 AND2X1_LOC_51/Y OR2X1_LOC_728/A 0.04fF
C4659 AND2X1_LOC_177/a_8_24# AND2X1_LOC_51/Y 0.03fF
C5302 AND2X1_LOC_51/Y AND2X1_LOC_239/a_8_24# 0.03fF
C5369 OR2X1_LOC_97/A AND2X1_LOC_51/Y 0.03fF
C5846 AND2X1_LOC_51/Y OR2X1_LOC_713/A 0.19fF
C6132 AND2X1_LOC_51/Y OR2X1_LOC_546/A 0.02fF
C6282 AND2X1_LOC_700/a_8_24# AND2X1_LOC_51/Y 0.04fF
C6379 OR2X1_LOC_639/B AND2X1_LOC_51/Y 0.03fF
C6425 OR2X1_LOC_333/B AND2X1_LOC_51/Y 0.11fF
C6844 OR2X1_LOC_154/A AND2X1_LOC_51/Y 0.34fF
C6991 AND2X1_LOC_51/Y OR2X1_LOC_198/A 0.35fF
C7377 AND2X1_LOC_821/a_8_24# AND2X1_LOC_51/Y 0.01fF
C7653 OR2X1_LOC_634/A AND2X1_LOC_51/Y 0.02fF
C8244 OR2X1_LOC_34/B AND2X1_LOC_51/Y 0.05fF
C8250 AND2X1_LOC_107/a_8_24# AND2X1_LOC_51/Y 0.03fF
C8698 AND2X1_LOC_600/a_8_24# AND2X1_LOC_51/Y 0.02fF
C9303 AND2X1_LOC_51/Y OR2X1_LOC_355/A 0.04fF
C9458 OR2X1_LOC_379/a_8_216# AND2X1_LOC_51/Y 0.14fF
C9763 OR2X1_LOC_614/Y AND2X1_LOC_51/Y 0.01fF
C10326 AND2X1_LOC_51/Y OR2X1_LOC_33/B 0.03fF
C10348 AND2X1_LOC_79/a_8_24# AND2X1_LOC_51/Y 0.01fF
C10589 AND2X1_LOC_51/Y OR2X1_LOC_113/B 0.52fF
C10798 OR2X1_LOC_532/B AND2X1_LOC_51/Y 0.13fF
C11418 OR2X1_LOC_162/Y AND2X1_LOC_51/Y 0.10fF
C11431 AND2X1_LOC_51/Y OR2X1_LOC_729/a_8_216# 0.02fF
C11885 OR2X1_LOC_710/B AND2X1_LOC_51/Y 0.01fF
C12358 AND2X1_LOC_52/a_8_24# AND2X1_LOC_51/Y 0.14fF
C12736 VDD AND2X1_LOC_51/Y 2.52fF
C12856 OR2X1_LOC_836/B AND2X1_LOC_51/Y 0.34fF
C13233 OR2X1_LOC_334/B AND2X1_LOC_51/Y 0.03fF
C13398 AND2X1_LOC_51/Y AND2X1_LOC_418/a_8_24# 0.02fF
C13608 OR2X1_LOC_676/Y AND2X1_LOC_51/Y 0.46fF
C13626 OR2X1_LOC_834/A AND2X1_LOC_51/Y 0.03fF
C13996 AND2X1_LOC_83/a_8_24# AND2X1_LOC_51/Y 0.01fF
C14205 OR2X1_LOC_602/B AND2X1_LOC_51/Y 0.01fF
C14763 AND2X1_LOC_51/Y OR2X1_LOC_115/B 0.03fF
C14915 OR2X1_LOC_840/A AND2X1_LOC_51/Y 0.06fF
C14955 AND2X1_LOC_145/a_8_24# AND2X1_LOC_51/Y 0.16fF
C15296 OR2X1_LOC_216/A AND2X1_LOC_51/Y 0.36fF
C15389 OR2X1_LOC_846/B AND2X1_LOC_51/Y 0.13fF
C15744 OR2X1_LOC_160/A AND2X1_LOC_51/Y 0.30fF
C15796 OR2X1_LOC_624/B AND2X1_LOC_51/Y 0.01fF
C15954 AND2X1_LOC_51/Y OR2X1_LOC_532/Y 0.01fF
C15990 AND2X1_LOC_51/Y OR2X1_LOC_130/Y 0.13fF
C16184 OR2X1_LOC_447/A AND2X1_LOC_51/Y 0.01fF
C16568 AND2X1_LOC_51/Y OR2X1_LOC_78/Y 0.02fF
C16960 AND2X1_LOC_163/a_8_24# AND2X1_LOC_51/Y 0.01fF
C17054 OR2X1_LOC_185/A AND2X1_LOC_51/Y 0.04fF
C17493 AND2X1_LOC_158/a_8_24# AND2X1_LOC_51/Y 0.17fF
C18344 OR2X1_LOC_379/Y AND2X1_LOC_51/Y 0.04fF
C18373 OR2X1_LOC_114/Y AND2X1_LOC_51/Y 0.03fF
C18978 AND2X1_LOC_51/Y AND2X1_LOC_238/a_8_24# 0.07fF
C19220 OR2X1_LOC_643/A AND2X1_LOC_51/Y 0.03fF
C19224 OR2X1_LOC_778/Y AND2X1_LOC_51/Y 0.04fF
C19449 AND2X1_LOC_91/B AND2X1_LOC_51/Y 1.08fF
C19634 OR2X1_LOC_799/A AND2X1_LOC_51/Y 0.22fF
C20024 OR2X1_LOC_105/a_8_216# AND2X1_LOC_51/Y 0.06fF
C20081 AND2X1_LOC_56/B AND2X1_LOC_51/Y 1.94fF
C21784 OR2X1_LOC_506/A AND2X1_LOC_51/Y 0.59fF
C21888 AND2X1_LOC_420/a_8_24# AND2X1_LOC_51/Y 0.02fF
C22001 AND2X1_LOC_51/Y OR2X1_LOC_180/B 0.03fF
C22401 AND2X1_LOC_51/Y OR2X1_LOC_788/B 0.02fF
C22539 OR2X1_LOC_467/B AND2X1_LOC_51/Y 0.18fF
C23097 OR2X1_LOC_210/B AND2X1_LOC_51/Y 0.13fF
C23438 OR2X1_LOC_235/B AND2X1_LOC_51/Y 0.03fF
C23510 AND2X1_LOC_393/a_8_24# AND2X1_LOC_51/Y 0.01fF
C23859 OR2X1_LOC_703/A AND2X1_LOC_51/Y 0.03fF
C24231 AND2X1_LOC_51/Y OR2X1_LOC_362/A 0.03fF
C24372 AND2X1_LOC_680/a_8_24# AND2X1_LOC_51/Y 0.05fF
C24491 AND2X1_LOC_51/Y OR2X1_LOC_771/B 0.10fF
C24516 AND2X1_LOC_51/Y OR2X1_LOC_776/A 0.03fF
C24934 AND2X1_LOC_51/Y OR2X1_LOC_593/B 0.03fF
C24961 OR2X1_LOC_506/a_8_216# AND2X1_LOC_51/Y 0.02fF
C25320 AND2X1_LOC_51/Y OR2X1_LOC_317/B 0.02fF
C25967 OR2X1_LOC_148/B AND2X1_LOC_51/Y 0.13fF
C26017 AND2X1_LOC_69/Y AND2X1_LOC_51/Y 0.01fF
C26078 OR2X1_LOC_506/B AND2X1_LOC_51/Y 0.39fF
C26892 AND2X1_LOC_69/a_8_24# AND2X1_LOC_51/Y 0.01fF
C26944 AND2X1_LOC_51/Y AND2X1_LOC_428/a_8_24# 0.01fF
C27266 OR2X1_LOC_130/A AND2X1_LOC_51/Y 0.08fF
C27688 OR2X1_LOC_449/B AND2X1_LOC_51/Y 0.09fF
C27705 OR2X1_LOC_636/A AND2X1_LOC_51/Y 0.01fF
C28052 OR2X1_LOC_317/a_8_216# AND2X1_LOC_51/Y 0.01fF
C28895 AND2X1_LOC_52/a_36_24# AND2X1_LOC_51/Y 0.01fF
C28945 OR2X1_LOC_400/B AND2X1_LOC_51/Y 0.01fF
C29394 AND2X1_LOC_525/a_8_24# AND2X1_LOC_51/Y 0.03fF
C29792 OR2X1_LOC_831/a_8_216# AND2X1_LOC_51/Y 0.02fF
C29911 AND2X1_LOC_51/Y AND2X1_LOC_52/Y 0.02fF
C29999 AND2X1_LOC_51/Y AND2X1_LOC_238/a_36_24# 0.01fF
C30881 OR2X1_LOC_149/B AND2X1_LOC_51/Y 0.03fF
C31019 OR2X1_LOC_105/Y AND2X1_LOC_51/Y 0.01fF
C31333 AND2X1_LOC_51/Y OR2X1_LOC_355/a_8_216# 0.01fF
C31458 AND2X1_LOC_145/a_36_24# AND2X1_LOC_51/Y 0.01fF
C31554 OR2X1_LOC_614/a_8_216# AND2X1_LOC_51/Y 0.01fF
C32396 AND2X1_LOC_51/Y OR2X1_LOC_451/B 0.01fF
C32523 AND2X1_LOC_51/Y OR2X1_LOC_333/a_8_216# 0.01fF
C32534 AND2X1_LOC_51/Y OR2X1_LOC_334/A 0.16fF
C32590 OR2X1_LOC_506/Y AND2X1_LOC_51/Y 0.01fF
C33194 OR2X1_LOC_636/B AND2X1_LOC_51/Y 0.01fF
C33447 OR2X1_LOC_856/A AND2X1_LOC_51/Y 0.02fF
C33488 AND2X1_LOC_51/Y OR2X1_LOC_730/A 0.04fF
C33886 AND2X1_LOC_51/Y OR2X1_LOC_160/Y 0.02fF
C33962 OR2X1_LOC_330/Y AND2X1_LOC_51/Y 0.01fF
C34403 AND2X1_LOC_584/a_8_24# AND2X1_LOC_51/Y 0.01fF
C35624 OR2X1_LOC_678/Y AND2X1_LOC_51/Y 0.05fF
C35866 AND2X1_LOC_51/Y OR2X1_LOC_777/B 0.05fF
C36079 OR2X1_LOC_493/A AND2X1_LOC_51/Y 0.94fF
C36329 OR2X1_LOC_198/a_8_216# AND2X1_LOC_51/Y 0.03fF
C36967 AND2X1_LOC_67/Y AND2X1_LOC_51/Y 0.02fF
C37487 OR2X1_LOC_705/B AND2X1_LOC_51/Y 0.26fF
C39043 OR2X1_LOC_319/B AND2X1_LOC_51/Y 0.01fF
C39441 AND2X1_LOC_103/a_8_24# AND2X1_LOC_51/Y 0.01fF
C39474 AND2X1_LOC_331/a_8_24# AND2X1_LOC_51/Y 0.02fF
C39933 OR2X1_LOC_147/a_8_216# AND2X1_LOC_51/Y 0.01fF
C39965 AND2X1_LOC_165/a_8_24# AND2X1_LOC_51/Y 0.09fF
C40295 OR2X1_LOC_635/a_8_216# AND2X1_LOC_51/Y 0.01fF
C40354 OR2X1_LOC_287/B AND2X1_LOC_51/Y 0.07fF
C40410 OR2X1_LOC_148/A AND2X1_LOC_51/Y 0.10fF
C40761 OR2X1_LOC_831/a_36_216# AND2X1_LOC_51/Y 0.02fF
C41496 OR2X1_LOC_318/A AND2X1_LOC_51/Y 0.01fF
C41514 OR2X1_LOC_151/A AND2X1_LOC_51/Y 0.14fF
C41883 OR2X1_LOC_198/a_36_216# AND2X1_LOC_51/Y 0.03fF
C43645 AND2X1_LOC_51/Y OR2X1_LOC_334/a_8_216# 0.01fF
C44022 AND2X1_LOC_51/Y OR2X1_LOC_308/Y 0.02fF
C44274 AND2X1_LOC_516/a_8_24# AND2X1_LOC_51/Y 0.06fF
C44682 OR2X1_LOC_835/A AND2X1_LOC_51/Y 0.01fF
C45049 AND2X1_LOC_24/a_8_24# AND2X1_LOC_51/Y 0.01fF
C45115 AND2X1_LOC_601/a_8_24# AND2X1_LOC_51/Y 0.02fF
C45964 AND2X1_LOC_314/a_8_24# AND2X1_LOC_51/Y 0.02fF
C46028 AND2X1_LOC_822/a_8_24# AND2X1_LOC_51/Y 0.01fF
C46042 AND2X1_LOC_525/a_36_24# AND2X1_LOC_51/Y 0.01fF
C46056 AND2X1_LOC_51/Y AND2X1_LOC_816/a_8_24# 0.01fF
C46943 OR2X1_LOC_473/Y AND2X1_LOC_51/Y 0.15fF
C47611 OR2X1_LOC_208/A AND2X1_LOC_51/Y 0.02fF
C47685 OR2X1_LOC_598/Y AND2X1_LOC_51/Y 0.02fF
C48100 AND2X1_LOC_51/Y OR2X1_LOC_356/A 0.25fF
C48151 OR2X1_LOC_614/a_36_216# AND2X1_LOC_51/Y -0.00fF
C48662 OR2X1_LOC_810/A AND2X1_LOC_51/Y 1.76fF
C48947 OR2X1_LOC_715/B AND2X1_LOC_51/Y 0.10fF
C49291 AND2X1_LOC_51/Y OR2X1_LOC_338/B 0.05fF
C49920 OR2X1_LOC_687/Y AND2X1_LOC_51/Y 0.03fF
C50362 OR2X1_LOC_835/B AND2X1_LOC_51/Y 0.22fF
C50590 AND2X1_LOC_91/a_8_24# AND2X1_LOC_51/Y 0.06fF
C50698 AND2X1_LOC_51/Y OR2X1_LOC_78/A 0.42fF
C50762 OR2X1_LOC_602/A AND2X1_LOC_51/Y 0.04fF
C51541 OR2X1_LOC_147/B AND2X1_LOC_51/Y 0.02fF
C51556 OR2X1_LOC_317/A AND2X1_LOC_51/Y 0.04fF
C51717 AND2X1_LOC_51/Y OR2X1_LOC_318/B 0.03fF
C51880 OR2X1_LOC_121/Y AND2X1_LOC_51/Y 0.07fF
C51937 OR2X1_LOC_538/A AND2X1_LOC_51/Y 0.03fF
C52033 AND2X1_LOC_79/Y AND2X1_LOC_51/Y 0.01fF
C54773 AND2X1_LOC_51/Y OR2X1_LOC_338/A 0.17fF
C54803 OR2X1_LOC_186/Y AND2X1_LOC_51/Y 0.04fF
C55409 OR2X1_LOC_574/A AND2X1_LOC_51/Y 0.76fF
C55411 AND2X1_LOC_51/Y OR2X1_LOC_33/A 0.01fF
C56824 AND2X1_LOC_51/Y VSS 1.00fF
C3304 VDD OR2X1_LOC_426/Y 0.12fF
C21658 OR2X1_LOC_426/Y OR2X1_LOC_427/Y 0.05fF
C22183 OR2X1_LOC_70/Y OR2X1_LOC_426/Y 0.01fF
C27145 OR2X1_LOC_426/Y AND2X1_LOC_450/a_8_24# 0.23fF
C36700 OR2X1_LOC_604/A OR2X1_LOC_426/Y 0.02fF
C49067 OR2X1_LOC_426/Y AND2X1_LOC_451/Y 0.01fF
C57000 OR2X1_LOC_426/Y VSS 0.06fF
C5221 OR2X1_LOC_45/B OR2X1_LOC_694/Y 0.05fF
C14279 OR2X1_LOC_694/Y OR2X1_LOC_695/Y 0.21fF
C27160 OR2X1_LOC_3/Y OR2X1_LOC_694/Y 0.03fF
C44104 OR2X1_LOC_694/Y OR2X1_LOC_52/B 0.03fF
C54308 OR2X1_LOC_695/a_8_216# OR2X1_LOC_694/Y 0.41fF
C57630 OR2X1_LOC_694/Y VSS 0.21fF
C155 OR2X1_LOC_40/Y OR2X1_LOC_135/Y 0.01fF
C190 OR2X1_LOC_40/Y OR2X1_LOC_815/a_8_216# 0.01fF
C194 OR2X1_LOC_40/Y AND2X1_LOC_98/a_8_24# 0.01fF
C287 OR2X1_LOC_40/Y AND2X1_LOC_848/Y 0.15fF
C357 OR2X1_LOC_40/Y OR2X1_LOC_617/Y 0.06fF
C1241 OR2X1_LOC_40/Y OR2X1_LOC_258/Y 0.61fF
C1320 OR2X1_LOC_40/Y AND2X1_LOC_318/Y 0.02fF
C1349 OR2X1_LOC_40/Y OR2X1_LOC_815/Y 0.02fF
C1511 OR2X1_LOC_40/Y OR2X1_LOC_759/A 0.05fF
C1545 OR2X1_LOC_40/Y OR2X1_LOC_698/Y 0.01fF
C1967 OR2X1_LOC_40/Y AND2X1_LOC_508/A 0.02fF
C2067 OR2X1_LOC_40/Y OR2X1_LOC_385/Y 0.03fF
C2323 OR2X1_LOC_40/Y OR2X1_LOC_764/a_8_216# 0.09fF
C2344 OR2X1_LOC_40/Y AND2X1_LOC_810/B 0.42fF
C2424 OR2X1_LOC_40/Y OR2X1_LOC_165/Y 0.01fF
C3238 OR2X1_LOC_40/Y AND2X1_LOC_715/A 0.03fF
C3724 AND2X1_LOC_729/Y OR2X1_LOC_40/Y 0.03fF
C3751 AND2X1_LOC_784/A OR2X1_LOC_40/Y 0.10fF
C4143 OR2X1_LOC_40/Y OR2X1_LOC_52/B 0.96fF
C4190 OR2X1_LOC_40/Y OR2X1_LOC_755/A 0.93fF
C4493 OR2X1_LOC_165/a_8_216# OR2X1_LOC_40/Y 0.01fF
C5791 OR2X1_LOC_40/Y OR2X1_LOC_680/A 10.75fF
C6143 OR2X1_LOC_757/A OR2X1_LOC_40/Y 0.07fF
C6232 OR2X1_LOC_40/Y OR2X1_LOC_626/a_8_216# 0.02fF
C6552 OR2X1_LOC_40/Y AND2X1_LOC_436/Y 0.16fF
C6888 OR2X1_LOC_40/Y OR2X1_LOC_152/a_8_216# 0.02fF
C7000 OR2X1_LOC_40/Y OR2X1_LOC_745/a_36_216# 0.02fF
C7132 OR2X1_LOC_40/Y OR2X1_LOC_609/A 0.03fF
C7545 OR2X1_LOC_40/Y AND2X1_LOC_266/Y 0.03fF
C7584 OR2X1_LOC_40/Y OR2X1_LOC_387/Y 0.11fF
C8401 OR2X1_LOC_40/Y OR2X1_LOC_265/a_8_216# 0.03fF
C8664 OR2X1_LOC_40/Y OR2X1_LOC_384/Y 0.01fF
C8777 AND2X1_LOC_391/Y OR2X1_LOC_40/Y 0.01fF
C9737 OR2X1_LOC_40/Y AND2X1_LOC_673/a_8_24# 0.01fF
C9757 OR2X1_LOC_40/Y OR2X1_LOC_74/A 1.74fF
C10020 OR2X1_LOC_40/Y OR2X1_LOC_626/Y 0.03fF
C10542 OR2X1_LOC_40/Y OR2X1_LOC_235/a_8_216# 0.01fF
C10578 OR2X1_LOC_40/Y OR2X1_LOC_239/Y 0.06fF
C11708 OR2X1_LOC_40/Y OR2X1_LOC_505/Y 0.01fF
C11834 OR2X1_LOC_40/Y OR2X1_LOC_626/a_36_216# 0.02fF
C12433 OR2X1_LOC_40/Y OR2X1_LOC_72/Y 0.01fF
C12450 OR2X1_LOC_40/Y OR2X1_LOC_152/a_36_216# 0.02fF
C12558 OR2X1_LOC_40/Y AND2X1_LOC_758/a_36_24# 0.01fF
C12665 OR2X1_LOC_670/a_8_216# OR2X1_LOC_40/Y 0.08fF
C12706 OR2X1_LOC_40/Y OR2X1_LOC_680/Y 0.03fF
C13401 OR2X1_LOC_40/Y OR2X1_LOC_764/a_36_216# 0.03fF
C13475 OR2X1_LOC_40/Y AND2X1_LOC_168/a_8_24# 0.02fF
C13522 OR2X1_LOC_40/Y AND2X1_LOC_303/A 0.31fF
C13554 OR2X1_LOC_40/Y OR2X1_LOC_665/Y 0.01fF
C13678 OR2X1_LOC_40/Y OR2X1_LOC_609/Y 0.15fF
C13802 AND2X1_LOC_802/B OR2X1_LOC_40/Y 0.03fF
C14235 AND2X1_LOC_383/a_8_24# OR2X1_LOC_40/Y 0.01fF
C15194 OR2X1_LOC_40/Y OR2X1_LOC_69/Y 0.01fF
C15248 OR2X1_LOC_40/Y OR2X1_LOC_665/a_8_216# 0.01fF
C15256 OR2X1_LOC_40/Y AND2X1_LOC_537/Y 0.02fF
C15328 OR2X1_LOC_40/Y OR2X1_LOC_437/a_8_216# 0.01fF
C15439 OR2X1_LOC_40/Y OR2X1_LOC_171/a_8_216# 0.01fF
C15479 OR2X1_LOC_40/Y OR2X1_LOC_13/Y 0.03fF
C15498 OR2X1_LOC_40/Y OR2X1_LOC_627/Y 0.03fF
C15674 OR2X1_LOC_40/Y OR2X1_LOC_295/Y 0.07fF
C15951 OR2X1_LOC_40/Y OR2X1_LOC_441/a_8_216# 0.03fF
C16788 OR2X1_LOC_40/Y OR2X1_LOC_496/a_8_216# 0.14fF
C17150 OR2X1_LOC_516/Y OR2X1_LOC_40/Y 0.07fF
C17670 OR2X1_LOC_40/Y AND2X1_LOC_348/A 0.03fF
C17812 OR2X1_LOC_40/Y OR2X1_LOC_442/a_8_216# 0.07fF
C17902 OR2X1_LOC_40/Y AND2X1_LOC_846/a_8_24# 0.01fF
C18067 OR2X1_LOC_125/a_8_216# OR2X1_LOC_40/Y 0.01fF
C18509 OR2X1_LOC_40/Y VDD 2.02fF
C18592 OR2X1_LOC_40/Y OR2X1_LOC_616/Y 0.44fF
C18655 OR2X1_LOC_40/Y AND2X1_LOC_389/a_8_24# 0.03fF
C18767 OR2X1_LOC_40/Y OR2X1_LOC_674/Y 0.01fF
C18798 OR2X1_LOC_40/Y OR2X1_LOC_67/Y 3.78fF
C19313 AND2X1_LOC_370/a_8_24# OR2X1_LOC_40/Y 0.02fF
C19429 OR2X1_LOC_40/Y OR2X1_LOC_531/a_8_216# 0.15fF
C19747 OR2X1_LOC_494/A OR2X1_LOC_40/Y 0.01fF
C21494 OR2X1_LOC_45/B OR2X1_LOC_40/Y 1.46fF
C21552 OR2X1_LOC_40/Y OR2X1_LOC_292/a_8_216# 0.03fF
C21926 OR2X1_LOC_40/Y OR2X1_LOC_158/A 1.67fF
C21971 OR2X1_LOC_40/Y AND2X1_LOC_98/Y 0.01fF
C22364 OR2X1_LOC_40/Y OR2X1_LOC_482/Y 0.12fF
C22438 OR2X1_LOC_40/Y OR2X1_LOC_586/Y 0.07fF
C22499 OR2X1_LOC_40/Y OR2X1_LOC_748/A 0.02fF
C22554 OR2X1_LOC_40/Y OR2X1_LOC_304/Y 0.13fF
C23015 OR2X1_LOC_40/Y OR2X1_LOC_815/A 0.01fF
C23493 OR2X1_LOC_40/Y AND2X1_LOC_848/A 0.01fF
C23906 OR2X1_LOC_40/Y OR2X1_LOC_41/a_8_216# 0.07fF
C24217 OR2X1_LOC_40/Y AND2X1_LOC_390/B 0.01fF
C24247 OR2X1_LOC_40/Y OR2X1_LOC_431/Y 0.46fF
C24453 OR2X1_LOC_40/Y OR2X1_LOC_309/Y 0.01fF
C24563 OR2X1_LOC_40/Y AND2X1_LOC_840/B 0.02fF
C25390 OR2X1_LOC_40/Y AND2X1_LOC_303/B 0.03fF
C26222 OR2X1_LOC_91/Y OR2X1_LOC_40/Y 0.40fF
C26282 OR2X1_LOC_40/Y OR2X1_LOC_527/Y 0.03fF
C26493 OR2X1_LOC_40/Y OR2X1_LOC_171/Y 0.07fF
C27009 OR2X1_LOC_40/Y OR2X1_LOC_292/a_36_216# 0.03fF
C27014 OR2X1_LOC_40/Y AND2X1_LOC_335/a_8_24# 0.02fF
C27024 OR2X1_LOC_40/Y OR2X1_LOC_441/Y 0.50fF
C27059 OR2X1_LOC_519/Y OR2X1_LOC_40/Y 0.01fF
C27111 OR2X1_LOC_40/Y OR2X1_LOC_235/Y 0.02fF
C27658 OR2X1_LOC_40/Y OR2X1_LOC_173/a_8_216# 0.02fF
C27739 OR2X1_LOC_40/Y AND2X1_LOC_789/Y 0.06fF
C28017 OR2X1_LOC_40/Y OR2X1_LOC_125/Y 0.02fF
C28056 OR2X1_LOC_40/Y OR2X1_LOC_409/B 0.02fF
C28341 OR2X1_LOC_40/Y AND2X1_LOC_676/a_8_24# 0.04fF
C29106 OR2X1_LOC_40/Y OR2X1_LOC_235/B 0.07fF
C29345 OR2X1_LOC_40/Y AND2X1_LOC_721/A 0.01fF
C29370 OR2X1_LOC_40/Y OR2X1_LOC_331/Y 0.01fF
C29624 OR2X1_LOC_40/Y AND2X1_LOC_361/A 0.02fF
C30317 AND2X1_LOC_787/A OR2X1_LOC_40/Y 0.03fF
C30398 AND2X1_LOC_391/a_8_24# OR2X1_LOC_40/Y 0.01fF
C30432 OR2X1_LOC_40/Y OR2X1_LOC_127/a_8_216# 0.01fF
C31206 OR2X1_LOC_40/Y AND2X1_LOC_335/Y 0.01fF
C31281 OR2X1_LOC_40/Y OR2X1_LOC_619/Y 0.24fF
C32269 OR2X1_LOC_40/Y OR2X1_LOC_406/A 0.04fF
C32390 OR2X1_LOC_505/a_8_216# OR2X1_LOC_40/Y 0.01fF
C32463 OR2X1_LOC_40/Y OR2X1_LOC_292/Y 0.01fF
C33434 OR2X1_LOC_40/Y OR2X1_LOC_312/Y 0.03fF
C33661 OR2X1_LOC_40/Y OR2X1_LOC_13/B 0.25fF
C34536 OR2X1_LOC_528/Y OR2X1_LOC_40/Y 0.05fF
C35123 OR2X1_LOC_40/Y OR2X1_LOC_89/A 0.16fF
C35902 OR2X1_LOC_45/Y OR2X1_LOC_40/Y 0.07fF
C36018 OR2X1_LOC_40/Y AND2X1_LOC_727/A 0.03fF
C36222 OR2X1_LOC_40/Y OR2X1_LOC_821/Y 0.02fF
C36683 OR2X1_LOC_40/Y OR2X1_LOC_438/Y 0.16fF
C36719 OR2X1_LOC_40/Y AND2X1_LOC_621/Y 0.10fF
C36959 OR2X1_LOC_40/Y OR2X1_LOC_71/A 0.06fF
C37238 OR2X1_LOC_40/Y OR2X1_LOC_70/Y 0.30fF
C37289 OR2X1_LOC_40/Y OR2X1_LOC_504/Y 0.65fF
C37344 OR2X1_LOC_40/Y OR2X1_LOC_437/Y 0.17fF
C38340 OR2X1_LOC_40/Y AND2X1_LOC_535/Y 0.06fF
C38462 OR2X1_LOC_40/Y OR2X1_LOC_246/Y 0.16fF
C38779 OR2X1_LOC_40/Y OR2X1_LOC_16/A 0.65fF
C38804 OR2X1_LOC_40/Y OR2X1_LOC_108/Y 0.03fF
C38875 AND2X1_LOC_168/Y OR2X1_LOC_40/Y 0.14fF
C39314 OR2X1_LOC_40/Y AND2X1_LOC_676/a_36_24# 0.01fF
C39763 OR2X1_LOC_40/Y OR2X1_LOC_262/a_8_216# 0.03fF
C39825 OR2X1_LOC_40/Y AND2X1_LOC_729/B 0.03fF
C40253 OR2X1_LOC_40/Y OR2X1_LOC_679/A 0.03fF
C40266 OR2X1_LOC_40/Y AND2X1_LOC_227/Y 0.03fF
C40596 OR2X1_LOC_599/A OR2X1_LOC_40/Y 0.08fF
C40629 OR2X1_LOC_40/Y OR2X1_LOC_258/a_8_216# 0.01fF
C40641 OR2X1_LOC_40/Y AND2X1_LOC_389/a_36_24# 0.02fF
C41393 OR2X1_LOC_187/a_8_216# OR2X1_LOC_40/Y 0.07fF
C41443 OR2X1_LOC_40/Y OR2X1_LOC_127/Y 0.21fF
C41617 OR2X1_LOC_40/Y OR2X1_LOC_615/Y 0.03fF
C41798 OR2X1_LOC_40/Y OR2X1_LOC_813/a_8_216# 0.02fF
C41866 OR2X1_LOC_40/Y AND2X1_LOC_841/B 0.03fF
C42291 OR2X1_LOC_40/Y OR2X1_LOC_495/Y 0.09fF
C42444 OR2X1_LOC_40/Y AND2X1_LOC_664/a_8_24# 0.01fF
C42563 OR2X1_LOC_40/Y OR2X1_LOC_384/a_8_216# 0.01fF
C42826 OR2X1_LOC_40/Y AND2X1_LOC_147/Y 0.03fF
C43247 OR2X1_LOC_40/Y OR2X1_LOC_3/Y 2.56fF
C43263 OR2X1_LOC_40/Y AND2X1_LOC_631/Y 0.07fF
C44091 OR2X1_LOC_40/Y AND2X1_LOC_610/a_8_24# 0.10fF
C44186 OR2X1_LOC_40/Y OR2X1_LOC_72/a_8_216# 0.02fF
C44518 OR2X1_LOC_40/Y OR2X1_LOC_173/Y 0.01fF
C45267 OR2X1_LOC_40/Y OR2X1_LOC_96/Y 0.01fF
C47945 OR2X1_LOC_40/Y AND2X1_LOC_709/a_8_24# 0.01fF
C48046 OR2X1_LOC_40/Y AND2X1_LOC_624/A 0.08fF
C48812 OR2X1_LOC_40/Y OR2X1_LOC_524/Y 5.32fF
C48916 OR2X1_LOC_40/Y OR2X1_LOC_763/Y 0.02fF
C49064 OR2X1_LOC_40/Y OR2X1_LOC_746/Y 0.06fF
C49327 OR2X1_LOC_40/Y OR2X1_LOC_670/Y 0.02fF
C49775 OR2X1_LOC_40/Y OR2X1_LOC_612/B 0.03fF
C49826 OR2X1_LOC_40/Y OR2X1_LOC_295/a_8_216# 0.01fF
C50411 OR2X1_LOC_40/Y AND2X1_LOC_608/a_8_24# 0.01fF
C50830 OR2X1_LOC_40/Y OR2X1_LOC_142/Y 0.14fF
C51017 OR2X1_LOC_40/Y OR2X1_LOC_262/Y 0.04fF
C51852 OR2X1_LOC_40/Y OR2X1_LOC_91/a_8_216# 0.02fF
C52117 OR2X1_LOC_177/Y OR2X1_LOC_40/Y 0.02fF
C52137 OR2X1_LOC_604/A OR2X1_LOC_40/Y 0.68fF
C52138 OR2X1_LOC_40/Y OR2X1_LOC_745/a_8_216# 0.01fF
C52140 OR2X1_LOC_40/Y AND2X1_LOC_758/a_8_24# 0.06fF
C52550 OR2X1_LOC_176/Y OR2X1_LOC_40/Y 0.05fF
C52666 OR2X1_LOC_40/Y OR2X1_LOC_265/Y 0.01fF
C53012 OR2X1_LOC_40/Y OR2X1_LOC_813/a_36_216# 0.03fF
C53193 OR2X1_LOC_40/Y AND2X1_LOC_633/Y 0.02fF
C53373 AND2X1_LOC_539/Y OR2X1_LOC_40/Y 0.03fF
C53438 OR2X1_LOC_40/Y AND2X1_LOC_711/A 0.01fF
C54255 OR2X1_LOC_40/Y AND2X1_LOC_434/Y 0.14fF
C54366 OR2X1_LOC_496/Y OR2X1_LOC_40/Y 0.06fF
C54699 OR2X1_LOC_40/Y OR2X1_LOC_674/a_8_216# 0.02fF
C55662 OR2X1_LOC_40/Y OR2X1_LOC_239/a_8_216# 0.14fF
C57883 OR2X1_LOC_40/Y VSS 1.36fF
C945 OR2X1_LOC_3/Y AND2X1_LOC_196/a_8_24# 0.06fF
C1618 OR2X1_LOC_3/Y OR2X1_LOC_766/Y 0.02fF
C2148 AND2X1_LOC_789/a_8_24# OR2X1_LOC_3/Y 0.01fF
C2499 OR2X1_LOC_3/Y OR2X1_LOC_135/Y 0.75fF
C2538 OR2X1_LOC_3/Y OR2X1_LOC_815/a_8_216# 0.02fF
C2645 OR2X1_LOC_3/Y AND2X1_LOC_848/Y 0.03fF
C3018 AND2X1_LOC_160/a_8_24# OR2X1_LOC_3/Y 0.01fF
C3800 OR2X1_LOC_759/A OR2X1_LOC_3/Y 0.02fF
C3831 OR2X1_LOC_3/Y OR2X1_LOC_697/a_8_216# -0.00fF
C3843 OR2X1_LOC_3/Y OR2X1_LOC_698/Y 0.01fF
C5974 AND2X1_LOC_784/A OR2X1_LOC_3/Y 0.41fF
C6005 OR2X1_LOC_3/Y OR2X1_LOC_481/Y 0.01fF
C6028 OR2X1_LOC_3/Y AND2X1_LOC_639/A 0.02fF
C6103 OR2X1_LOC_3/Y OR2X1_LOC_172/Y 0.27fF
C6192 OR2X1_LOC_3/Y OR2X1_LOC_397/Y 0.34fF
C6387 OR2X1_LOC_3/Y OR2X1_LOC_52/B 0.23fF
C6490 OR2X1_LOC_3/Y AND2X1_LOC_216/A 0.22fF
C6675 OR2X1_LOC_3/Y OR2X1_LOC_281/Y 0.33fF
C8048 OR2X1_LOC_3/Y OR2X1_LOC_815/a_36_216# 0.03fF
C8100 OR2X1_LOC_3/Y OR2X1_LOC_16/Y 0.34fF
C8540 OR2X1_LOC_757/A OR2X1_LOC_3/Y 0.09fF
C8629 OR2X1_LOC_3/Y OR2X1_LOC_423/a_8_216# 0.01fF
C8756 OR2X1_LOC_3/Y OR2X1_LOC_399/a_8_216# 0.01fF
C9022 OR2X1_LOC_3/Y OR2X1_LOC_588/Y 0.03fF
C9870 OR2X1_LOC_3/Y AND2X1_LOC_266/Y 0.15fF
C10849 OR2X1_LOC_3/Y OR2X1_LOC_384/Y 0.79fF
C10973 OR2X1_LOC_3/Y OR2X1_LOC_131/a_8_216# 0.01fF
C11018 AND2X1_LOC_391/Y OR2X1_LOC_3/Y 0.04fF
C11552 AND2X1_LOC_777/a_36_24# OR2X1_LOC_3/Y 0.01fF
C11706 OR2X1_LOC_3/Y OR2X1_LOC_423/Y 0.01fF
C11980 OR2X1_LOC_3/Y OR2X1_LOC_74/A 0.10fF
C13545 OR2X1_LOC_3/Y AND2X1_LOC_339/B 0.03fF
C13593 OR2X1_LOC_3/Y OR2X1_LOC_816/a_8_216# 0.03fF
C13679 OR2X1_LOC_3/Y AND2X1_LOC_633/a_8_24# 0.01fF
C13931 OR2X1_LOC_106/Y OR2X1_LOC_3/Y 0.01fF
C14107 OR2X1_LOC_3/Y AND2X1_LOC_847/Y 0.01fF
C14495 OR2X1_LOC_3/Y AND2X1_LOC_99/A 0.12fF
C14882 OR2X1_LOC_3/Y OR2X1_LOC_697/Y 0.01fF
C15006 OR2X1_LOC_3/Y OR2X1_LOC_696/Y 0.01fF
C15325 OR2X1_LOC_3/Y OR2X1_LOC_595/a_8_216# 0.02fF
C15379 OR2X1_LOC_3/Y OR2X1_LOC_431/a_8_216# 0.01fF
C15763 OR2X1_LOC_3/Y OR2X1_LOC_665/Y 0.02fF
C16345 OR2X1_LOC_3/Y OR2X1_LOC_376/Y 0.02fF
C16413 AND2X1_LOC_383/a_8_24# OR2X1_LOC_3/Y 0.01fF
C16522 OR2X1_LOC_122/a_8_216# OR2X1_LOC_3/Y 0.01fF
C16579 OR2X1_LOC_695/a_8_216# OR2X1_LOC_3/Y 0.02fF
C17453 OR2X1_LOC_3/Y OR2X1_LOC_67/a_8_216# 0.01fF
C17463 OR2X1_LOC_305/a_8_216# OR2X1_LOC_3/Y 0.02fF
C17517 OR2X1_LOC_3/Y OR2X1_LOC_665/a_8_216# 0.01fF
C17522 OR2X1_LOC_3/Y AND2X1_LOC_537/Y 0.07fF
C17745 OR2X1_LOC_3/Y OR2X1_LOC_13/Y 0.03fF
C18638 AND2X1_LOC_714/B OR2X1_LOC_3/Y 0.07fF
C18645 OR2X1_LOC_106/a_8_216# OR2X1_LOC_3/Y -0.00fF
C19112 OR2X1_LOC_3/Y OR2X1_LOC_816/a_36_216# 0.03fF
C19452 OR2X1_LOC_117/a_8_216# OR2X1_LOC_3/Y 0.01fF
C19778 OR2X1_LOC_3/Y AND2X1_LOC_793/B 0.03fF
C20352 OR2X1_LOC_3/Y OR2X1_LOC_583/a_8_216# 0.02fF
C20515 OR2X1_LOC_3/Y OR2X1_LOC_131/Y 0.04fF
C20803 VDD OR2X1_LOC_3/Y 1.01fF
C21019 OR2X1_LOC_3/Y OR2X1_LOC_67/Y 0.07fF
C21377 OR2X1_LOC_3/Y OR2X1_LOC_248/Y 0.02fF
C21604 OR2X1_LOC_3/Y OR2X1_LOC_56/Y 0.01fF
C21832 OR2X1_LOC_3/Y AND2X1_LOC_307/Y 0.15fF
C22034 OR2X1_LOC_494/A OR2X1_LOC_3/Y 0.01fF
C22729 OR2X1_LOC_3/Y OR2X1_LOC_416/Y 0.03fF
C23041 OR2X1_LOC_3/Y OR2X1_LOC_281/a_8_216# 0.01fF
C23073 OR2X1_LOC_305/a_36_216# OR2X1_LOC_3/Y 0.02fF
C23462 OR2X1_LOC_3/Y OR2X1_LOC_45/a_8_216# 0.01fF
C23740 OR2X1_LOC_45/B OR2X1_LOC_3/Y 3.80fF
C23838 OR2X1_LOC_3/Y OR2X1_LOC_292/a_8_216# 0.01fF
C23895 OR2X1_LOC_3/Y OR2X1_LOC_767/a_8_216# 0.02fF
C23924 OR2X1_LOC_3/Y OR2X1_LOC_261/Y 0.01fF
C24201 OR2X1_LOC_158/A OR2X1_LOC_3/Y 1.93fF
C24640 OR2X1_LOC_3/Y OR2X1_LOC_816/Y 0.03fF
C24744 OR2X1_LOC_3/Y OR2X1_LOC_748/A 0.02fF
C24771 OR2X1_LOC_3/Y OR2X1_LOC_304/Y 0.17fF
C25156 OR2X1_LOC_3/Y OR2X1_LOC_117/Y 0.22fF
C25202 OR2X1_LOC_3/Y OR2X1_LOC_815/A 0.01fF
C25309 OR2X1_LOC_3/Y OR2X1_LOC_399/Y 0.02fF
C26355 OR2X1_LOC_3/Y OR2X1_LOC_316/Y 0.03fF
C26360 OR2X1_LOC_3/Y OR2X1_LOC_595/a_36_216# 0.01fF
C26434 OR2X1_LOC_3/Y OR2X1_LOC_431/Y 0.03fF
C26841 OR2X1_LOC_3/Y OR2X1_LOC_282/a_8_216# 0.01fF
C27741 OR2X1_LOC_3/Y OR2X1_LOC_751/A 0.10fF
C27920 OR2X1_LOC_3/Y OR2X1_LOC_118/a_8_216# 0.01fF
C28100 OR2X1_LOC_3/Y AND2X1_LOC_56/B 0.03fF
C28417 OR2X1_LOC_3/Y AND2X1_LOC_285/Y 0.01fF
C28514 OR2X1_LOC_305/Y OR2X1_LOC_3/Y 0.14fF
C28566 OR2X1_LOC_3/Y OR2X1_LOC_417/Y 0.03fF
C29333 OR2X1_LOC_3/Y AND2X1_LOC_139/B 0.03fF
C29616 OR2X1_LOC_135/a_8_216# OR2X1_LOC_3/Y 0.01fF
C29954 OR2X1_LOC_3/Y AND2X1_LOC_789/Y 0.03fF
C30280 OR2X1_LOC_3/Y OR2X1_LOC_409/B 0.03fF
C30897 OR2X1_LOC_3/Y AND2X1_LOC_249/a_8_24# 0.01fF
C31107 OR2X1_LOC_3/Y OR2X1_LOC_7/a_8_216# 0.01fF
C31445 OR2X1_LOC_3/Y AND2X1_LOC_319/A 0.07fF
C31515 OR2X1_LOC_3/Y AND2X1_LOC_708/a_8_24# 0.01fF
C31567 OR2X1_LOC_3/Y AND2X1_LOC_721/A 0.02fF
C31863 OR2X1_LOC_3/Y AND2X1_LOC_361/A 0.07fF
C32617 OR2X1_LOC_3/Y OR2X1_LOC_695/Y 0.01fF
C32659 AND2X1_LOC_391/a_8_24# OR2X1_LOC_3/Y 0.01fF
C32699 OR2X1_LOC_127/a_8_216# OR2X1_LOC_3/Y 0.09fF
C33561 OR2X1_LOC_3/Y OR2X1_LOC_619/Y 0.13fF
C34008 OR2X1_LOC_3/Y AND2X1_LOC_454/A 0.46fF
C34769 OR2X1_LOC_3/Y OR2X1_LOC_292/Y 0.01fF
C35719 OR2X1_LOC_3/Y AND2X1_LOC_307/a_8_24# 0.03fF
C35851 OR2X1_LOC_3/Y OR2X1_LOC_13/B 0.10fF
C36039 OR2X1_LOC_3/Y AND2X1_LOC_266/a_8_24# 0.01fF
C36361 OR2X1_LOC_3/Y OR2X1_LOC_595/A 1.89fF
C36796 OR2X1_LOC_3/Y OR2X1_LOC_583/Y 0.04fF
C36891 OR2X1_LOC_3/Y AND2X1_LOC_342/Y 0.04fF
C36965 OR2X1_LOC_3/Y AND2X1_LOC_712/B 0.39fF
C37220 OR2X1_LOC_3/Y OR2X1_LOC_765/Y 0.03fF
C37376 OR2X1_LOC_3/Y OR2X1_LOC_89/A 0.71fF
C37801 OR2X1_LOC_3/Y OR2X1_LOC_282/Y 0.21fF
C38076 OR2X1_LOC_3/Y AND2X1_LOC_707/a_8_24# 0.01fF
C38152 OR2X1_LOC_45/Y OR2X1_LOC_3/Y 1.18fF
C38173 OR2X1_LOC_127/a_36_216# OR2X1_LOC_3/Y 0.03fF
C38549 OR2X1_LOC_122/Y OR2X1_LOC_3/Y 0.33fF
C39541 OR2X1_LOC_70/Y OR2X1_LOC_3/Y 0.91fF
C39915 OR2X1_LOC_3/Y OR2X1_LOC_240/A 0.07fF
C40098 OR2X1_LOC_3/Y OR2X1_LOC_397/a_8_216# 0.01fF
C40549 OR2X1_LOC_3/Y OR2X1_LOC_767/Y 0.02fF
C40606 OR2X1_LOC_3/Y OR2X1_LOC_584/a_8_216# 0.02fF
C41023 OR2X1_LOC_3/Y OR2X1_LOC_16/A 0.36fF
C42106 OR2X1_LOC_3/Y AND2X1_LOC_729/B 0.03fF
C42604 OR2X1_LOC_3/Y AND2X1_LOC_227/Y 0.05fF
C43295 OR2X1_LOC_3/Y OR2X1_LOC_698/a_8_216# 0.01fF
C44068 AND2X1_LOC_707/Y OR2X1_LOC_3/Y 0.14fF
C44567 OR2X1_LOC_3/Y OR2X1_LOC_261/a_8_216# 0.01fF
C44664 OR2X1_LOC_3/Y AND2X1_LOC_379/a_8_24# 0.03fF
C44813 OR2X1_LOC_3/Y OR2X1_LOC_384/a_8_216# 0.01fF
C46725 OR2X1_LOC_3/Y OR2X1_LOC_766/a_8_216# 0.02fF
C47851 OR2X1_LOC_3/Y OR2X1_LOC_7/Y 0.01fF
C48309 OR2X1_LOC_3/Y AND2X1_LOC_196/Y 0.06fF
C50006 OR2X1_LOC_3/Y OR2X1_LOC_751/a_8_216# 0.01fF
C50669 OR2X1_LOC_3/Y AND2X1_LOC_434/a_8_24# 0.02fF
C51145 AND2X1_LOC_777/a_8_24# OR2X1_LOC_3/Y 0.03fF
C51183 OR2X1_LOC_3/Y OR2X1_LOC_481/a_8_216# 0.07fF
C51597 OR2X1_LOC_3/Y OR2X1_LOC_48/Y 0.04fF
C51899 OR2X1_LOC_3/Y AND2X1_LOC_160/Y 0.01fF
C52276 OR2X1_LOC_3/Y OR2X1_LOC_421/Y 0.01fF
C52456 OR2X1_LOC_3/Y OR2X1_LOC_273/Y 0.07fF
C52791 OR2X1_LOC_751/Y OR2X1_LOC_3/Y 0.01fF
C53211 OR2X1_LOC_3/Y OR2X1_LOC_16/a_8_216# 0.01fF
C53240 OR2X1_LOC_3/Y OR2X1_LOC_118/Y 0.07fF
C53271 OR2X1_LOC_3/Y OR2X1_LOC_262/Y 0.45fF
C53411 OR2X1_LOC_3/Y OR2X1_LOC_39/a_8_216# 0.09fF
C54399 OR2X1_LOC_604/A OR2X1_LOC_3/Y 0.09fF
C55434 OR2X1_LOC_3/Y AND2X1_LOC_633/Y 0.01fF
C55671 OR2X1_LOC_3/Y OR2X1_LOC_131/A 0.09fF
C57765 OR2X1_LOC_3/Y VSS 0.84fF
C18 AND2X1_LOC_729/Y OR2X1_LOC_70/Y 0.04fF
C41 AND2X1_LOC_784/A OR2X1_LOC_70/Y 0.07fF
C57 AND2X1_LOC_769/a_8_24# OR2X1_LOC_70/Y 0.06fF
C94 OR2X1_LOC_70/Y AND2X1_LOC_639/A 0.04fF
C178 OR2X1_LOC_70/Y OR2X1_LOC_172/Y 0.31fF
C403 OR2X1_LOC_70/Y OR2X1_LOC_674/a_36_216# 0.02fF
C473 OR2X1_LOC_70/Y OR2X1_LOC_52/B 0.16fF
C579 OR2X1_LOC_70/Y AND2X1_LOC_216/A 0.02fF
C764 OR2X1_LOC_70/Y OR2X1_LOC_584/Y 0.03fF
C938 OR2X1_LOC_70/Y AND2X1_LOC_356/B 0.03fF
C1247 OR2X1_LOC_70/Y OR2X1_LOC_485/Y 0.07fF
C1432 OR2X1_LOC_70/Y OR2X1_LOC_428/a_8_216# 0.01fF
C1757 OR2X1_LOC_70/Y AND2X1_LOC_593/Y 0.12fF
C2210 OR2X1_LOC_70/Y OR2X1_LOC_680/A 0.11fF
C2671 OR2X1_LOC_70/Y OR2X1_LOC_498/a_8_216# 0.07fF
C2986 OR2X1_LOC_70/Y AND2X1_LOC_436/Y 0.01fF
C3470 OR2X1_LOC_70/Y OR2X1_LOC_313/Y 0.01fF
C3625 OR2X1_LOC_70/Y OR2X1_LOC_331/a_8_216# 0.01fF
C3914 OR2X1_LOC_70/Y AND2X1_LOC_266/Y 0.03fF
C4372 OR2X1_LOC_70/Y AND2X1_LOC_451/Y 0.01fF
C4661 OR2X1_LOC_70/Y OR2X1_LOC_265/a_8_216# 0.01fF
C4983 OR2X1_LOC_70/Y OR2X1_LOC_131/a_8_216# 0.15fF
C6003 OR2X1_LOC_70/Y OR2X1_LOC_74/A 0.17fF
C6344 OR2X1_LOC_70/Y OR2X1_LOC_432/a_8_216# 0.14fF
C6817 OR2X1_LOC_70/Y OR2X1_LOC_432/Y 0.18fF
C7139 AND2X1_LOC_704/a_8_24# OR2X1_LOC_70/Y 0.01fF
C7581 OR2X1_LOC_70/Y AND2X1_LOC_339/B 0.03fF
C7664 OR2X1_LOC_70/Y OR2X1_LOC_586/a_8_216# 0.09fF
C9096 OR2X1_LOC_70/Y OR2X1_LOC_167/Y 0.16fF
C9517 OR2X1_LOC_70/Y OR2X1_LOC_431/a_8_216# 0.08fF
C9739 AND2X1_LOC_706/Y OR2X1_LOC_70/Y 0.05fF
C11038 OR2X1_LOC_70/Y AND2X1_LOC_436/a_8_24# 0.01fF
C11185 OR2X1_LOC_70/Y AND2X1_LOC_635/a_36_24# -0.00fF
C11560 OR2X1_LOC_70/Y OR2X1_LOC_418/Y 0.01fF
C11846 OR2X1_LOC_70/Y OR2X1_LOC_13/Y 0.02fF
C12702 AND2X1_LOC_714/B OR2X1_LOC_70/Y 0.01fF
C13477 OR2X1_LOC_516/Y OR2X1_LOC_70/Y 0.03fF
C14521 OR2X1_LOC_70/Y OR2X1_LOC_314/Y 0.01fF
C14572 OR2X1_LOC_70/Y OR2X1_LOC_131/Y 0.04fF
C14848 VDD OR2X1_LOC_70/Y 2.03fF
C14962 OR2X1_LOC_70/Y AND2X1_LOC_267/a_8_24# 0.01fF
C14992 OR2X1_LOC_70/Y AND2X1_LOC_389/a_8_24# 0.11fF
C15292 OR2X1_LOC_314/a_8_216# OR2X1_LOC_70/Y 0.02fF
C16677 OR2X1_LOC_70/Y OR2X1_LOC_416/Y 0.03fF
C17449 OR2X1_LOC_70/Y OR2X1_LOC_45/a_8_216# 0.01fF
C17720 OR2X1_LOC_45/B OR2X1_LOC_70/Y 0.29fF
C17986 OR2X1_LOC_70/Y OR2X1_LOC_428/Y 0.01fF
C18219 OR2X1_LOC_158/A OR2X1_LOC_70/Y 0.10fF
C18222 AND2X1_LOC_704/a_36_24# OR2X1_LOC_70/Y -0.00fF
C18760 OR2X1_LOC_70/Y OR2X1_LOC_586/Y 0.09fF
C18837 OR2X1_LOC_70/Y OR2X1_LOC_304/Y 0.32fF
C20055 OR2X1_LOC_70/Y AND2X1_LOC_317/a_8_24# 0.02fF
C20091 OR2X1_LOC_70/Y OR2X1_LOC_438/a_8_216# 0.01fF
C20356 OR2X1_LOC_70/Y OR2X1_LOC_765/a_8_216# 0.01fF
C20469 OR2X1_LOC_70/Y OR2X1_LOC_316/Y 0.03fF
C20531 OR2X1_LOC_70/Y AND2X1_LOC_390/B 0.58fF
C20558 OR2X1_LOC_70/Y OR2X1_LOC_431/Y 0.01fF
C20937 OR2X1_LOC_70/Y AND2X1_LOC_840/B 0.03fF
C21641 OR2X1_LOC_821/a_8_216# OR2X1_LOC_70/Y 0.07fF
C22063 OR2X1_LOC_70/Y OR2X1_LOC_118/a_8_216# 0.03fF
C22661 OR2X1_LOC_91/Y OR2X1_LOC_70/Y 0.07fF
C22681 OR2X1_LOC_70/Y AND2X1_LOC_446/a_8_24# 0.02fF
C22694 OR2X1_LOC_189/Y OR2X1_LOC_70/Y 0.03fF
C22717 OR2X1_LOC_70/Y OR2X1_LOC_527/Y 0.11fF
C22731 OR2X1_LOC_70/Y OR2X1_LOC_417/Y 0.04fF
C22734 OR2X1_LOC_70/Y OR2X1_LOC_311/Y 0.04fF
C22997 AND2X1_LOC_330/a_8_24# OR2X1_LOC_70/Y 0.01fF
C23479 OR2X1_LOC_70/Y AND2X1_LOC_436/B 0.11fF
C24028 OR2X1_LOC_70/Y OR2X1_LOC_173/a_8_216# 0.06fF
C24405 OR2X1_LOC_70/Y OR2X1_LOC_409/B 0.06fF
C24675 OR2X1_LOC_70/Y OR2X1_LOC_298/a_8_216# 0.05fF
C25122 OR2X1_LOC_70/Y OR2X1_LOC_109/a_8_216# 0.03fF
C25557 OR2X1_LOC_70/Y AND2X1_LOC_319/A 0.17fF
C25648 OR2X1_LOC_70/Y OR2X1_LOC_604/a_8_216# 0.01fF
C25694 OR2X1_LOC_70/Y OR2X1_LOC_331/Y 0.12fF
C25975 OR2X1_LOC_70/Y AND2X1_LOC_361/A 0.08fF
C26658 AND2X1_LOC_787/A OR2X1_LOC_70/Y 0.03fF
C27572 OR2X1_LOC_166/a_8_216# OR2X1_LOC_70/Y 0.01fF
C27644 OR2X1_LOC_70/Y OR2X1_LOC_619/Y 0.10fF
C28121 OR2X1_LOC_70/Y AND2X1_LOC_454/A 0.01fF
C28209 OR2X1_LOC_70/Y OR2X1_LOC_289/Y 0.03fF
C28433 OR2X1_LOC_331/A OR2X1_LOC_70/Y 0.37fF
C28620 OR2X1_LOC_70/Y OR2X1_LOC_406/A 0.48fF
C28808 OR2X1_LOC_329/Y OR2X1_LOC_70/Y 0.02fF
C29800 OR2X1_LOC_70/Y OR2X1_LOC_312/Y 0.68fF
C29858 OR2X1_LOC_70/Y OR2X1_LOC_75/a_8_216# 0.05fF
C29943 OR2X1_LOC_70/Y OR2X1_LOC_13/B 0.33fF
C30355 OR2X1_LOC_70/Y OR2X1_LOC_533/a_8_216# 0.01fF
C30469 OR2X1_LOC_70/Y OR2X1_LOC_595/A 0.24fF
C30942 OR2X1_LOC_528/Y OR2X1_LOC_70/Y 0.02fF
C31351 OR2X1_LOC_70/Y OR2X1_LOC_765/Y 0.01fF
C31477 OR2X1_LOC_70/Y OR2X1_LOC_89/A 2.92fF
C31575 OR2X1_LOC_70/Y AND2X1_LOC_451/a_8_24# 0.02fF
C32114 OR2X1_LOC_70/Y OR2X1_LOC_79/Y 0.02fF
C32232 OR2X1_LOC_45/Y OR2X1_LOC_70/Y 0.32fF
C32255 OR2X1_LOC_70/Y OR2X1_LOC_427/a_8_216# 0.03fF
C32316 OR2X1_LOC_70/Y AND2X1_LOC_727/A 0.03fF
C33080 OR2X1_LOC_438/Y OR2X1_LOC_70/Y 0.10fF
C33098 OR2X1_LOC_70/Y OR2X1_LOC_427/Y 0.01fF
C33124 OR2X1_LOC_70/Y AND2X1_LOC_621/Y 0.03fF
C33928 AND2X1_LOC_330/a_36_24# OR2X1_LOC_70/Y 0.01fF
C34719 AND2X1_LOC_535/Y OR2X1_LOC_70/Y 0.01fF
C34763 OR2X1_LOC_70/Y OR2X1_LOC_484/Y 0.07fF
C35105 OR2X1_LOC_70/Y OR2X1_LOC_16/A 0.34fF
C36074 OR2X1_LOC_70/Y OR2X1_LOC_109/Y 0.04fF
C36142 OR2X1_LOC_70/Y AND2X1_LOC_729/B 0.02fF
C36580 OR2X1_LOC_70/Y AND2X1_LOC_227/Y 0.10fF
C36603 OR2X1_LOC_70/Y OR2X1_LOC_813/Y 0.01fF
C36911 OR2X1_LOC_599/A OR2X1_LOC_70/Y 0.04fF
C37203 OR2X1_LOC_177/a_8_216# OR2X1_LOC_70/Y 0.01fF
C37254 OR2X1_LOC_70/Y AND2X1_LOC_535/a_8_24# 0.01fF
C38016 AND2X1_LOC_707/Y OR2X1_LOC_70/Y 0.02fF
C38162 OR2X1_LOC_70/Y AND2X1_LOC_841/B 0.17fF
C38542 OR2X1_LOC_166/Y OR2X1_LOC_70/Y 0.01fF
C38592 OR2X1_LOC_70/Y OR2X1_LOC_495/Y 0.03fF
C38608 OR2X1_LOC_70/Y AND2X1_LOC_450/a_8_24# 0.02fF
C40412 OR2X1_LOC_70/Y OR2X1_LOC_72/a_8_216# 0.02fF
C42074 OR2X1_LOC_70/Y OR2X1_LOC_189/A 0.06fF
C43491 OR2X1_LOC_70/Y OR2X1_LOC_311/a_8_216# 0.14fF
C43671 OR2X1_LOC_70/Y AND2X1_LOC_802/Y 0.03fF
C44124 OR2X1_LOC_70/Y AND2X1_LOC_778/Y 1.20fF
C44237 OR2X1_LOC_70/Y AND2X1_LOC_624/A 0.05fF
C44590 OR2X1_LOC_70/Y AND2X1_LOC_434/a_8_24# 0.01fF
C45047 OR2X1_LOC_524/Y OR2X1_LOC_70/Y 0.02fF
C45179 OR2X1_LOC_70/Y AND2X1_LOC_635/a_8_24# 0.01fF
C45253 OR2X1_LOC_70/Y OR2X1_LOC_172/a_8_216# 0.01fF
C45579 OR2X1_LOC_70/Y OR2X1_LOC_418/a_8_216# 0.01fF
C46538 OR2X1_LOC_70/Y OR2X1_LOC_75/Y 0.06fF
C47105 OR2X1_LOC_70/Y OR2X1_LOC_142/Y 0.03fF
C47342 OR2X1_LOC_70/Y OR2X1_LOC_118/Y 0.02fF
C47379 OR2X1_LOC_70/Y OR2X1_LOC_262/Y 1.04fF
C48526 OR2X1_LOC_177/Y OR2X1_LOC_70/Y 0.04fF
C48545 OR2X1_LOC_604/A OR2X1_LOC_70/Y 0.22fF
C48906 OR2X1_LOC_533/Y OR2X1_LOC_70/Y 0.01fF
C49039 OR2X1_LOC_70/Y OR2X1_LOC_265/Y 8.97fF
C49333 OR2X1_LOC_70/Y AND2X1_LOC_809/a_8_24# 0.11fF
C49585 OR2X1_LOC_70/Y AND2X1_LOC_450/Y 0.01fF
C49727 AND2X1_LOC_539/Y OR2X1_LOC_70/Y 0.79fF
C49801 OR2X1_LOC_70/Y OR2X1_LOC_131/A 0.31fF
C50332 OR2X1_LOC_70/Y OR2X1_LOC_298/Y 0.01fF
C50685 OR2X1_LOC_70/Y AND2X1_LOC_434/Y 0.03fF
C51091 OR2X1_LOC_70/Y OR2X1_LOC_674/a_8_216# 0.03fF
C51590 OR2X1_LOC_70/Y AND2X1_LOC_355/a_8_24# 0.01fF
C51667 OR2X1_LOC_70/Y OR2X1_LOC_72/a_36_216# 0.03fF
C52215 AND2X1_LOC_776/Y OR2X1_LOC_70/Y 0.26fF
C52703 OR2X1_LOC_70/Y OR2X1_LOC_135/Y 0.08fF
C53705 OR2X1_LOC_313/a_8_216# OR2X1_LOC_70/Y 0.09fF
C54542 OR2X1_LOC_70/Y OR2X1_LOC_385/Y 0.06fF
C54790 OR2X1_LOC_70/Y AND2X1_LOC_810/B 0.01fF
C56148 AND2X1_LOC_547/Y OR2X1_LOC_70/Y 0.04fF
C57784 OR2X1_LOC_70/Y VSS 1.33fF
C128 OR2X1_LOC_158/A OR2X1_LOC_56/Y 0.03fF
C1255 OR2X1_LOC_158/A OR2X1_LOC_416/Y 0.03fF
C1548 OR2X1_LOC_158/A OR2X1_LOC_281/a_8_216# 0.01fF
C2062 OR2X1_LOC_158/A AND2X1_LOC_116/Y 0.09fF
C2318 OR2X1_LOC_45/B OR2X1_LOC_158/A 0.35fF
C2393 OR2X1_LOC_158/A OR2X1_LOC_292/a_8_216# 0.01fF
C2458 OR2X1_LOC_158/A AND2X1_LOC_435/a_8_24# 0.06fF
C3206 OR2X1_LOC_158/A OR2X1_LOC_482/Y 0.03fF
C3328 OR2X1_LOC_158/A OR2X1_LOC_748/A 0.03fF
C4278 OR2X1_LOC_158/A AND2X1_LOC_848/A 0.16fF
C4913 OR2X1_LOC_158/A OR2X1_LOC_316/Y 0.04fF
C4966 OR2X1_LOC_158/A AND2X1_LOC_390/B 0.07fF
C5351 OR2X1_LOC_158/A OR2X1_LOC_74/a_8_216# 0.02fF
C5385 OR2X1_LOC_158/A OR2X1_LOC_282/a_8_216# 0.19fF
C5522 OR2X1_LOC_158/A OR2X1_LOC_257/Y 0.01fF
C6147 OR2X1_LOC_179/a_8_216# OR2X1_LOC_158/A 0.01fF
C6995 OR2X1_LOC_158/A AND2X1_LOC_285/Y 0.29fF
C7087 OR2X1_LOC_91/Y OR2X1_LOC_158/A 0.03fF
C7160 OR2X1_LOC_158/A OR2X1_LOC_417/Y 0.03fF
C7170 OR2X1_LOC_158/A OR2X1_LOC_311/Y 0.03fF
C7381 OR2X1_LOC_158/A AND2X1_LOC_780/a_8_24# 0.01fF
C7582 OR2X1_LOC_158/A AND2X1_LOC_276/Y 0.14fF
C7645 OR2X1_LOC_158/A AND2X1_LOC_831/Y 0.07fF
C7899 OR2X1_LOC_158/A AND2X1_LOC_335/a_8_24# 0.05fF
C7958 OR2X1_LOC_519/Y OR2X1_LOC_158/A 0.01fF
C7970 OR2X1_LOC_158/A AND2X1_LOC_436/B 0.65fF
C7976 OR2X1_LOC_158/A AND2X1_LOC_139/B 0.07fF
C8561 OR2X1_LOC_158/A AND2X1_LOC_462/Y 0.03fF
C8686 OR2X1_LOC_158/A AND2X1_LOC_789/Y 0.29fF
C8742 OR2X1_LOC_158/A OR2X1_LOC_108/a_8_216# 0.02fF
C8837 OR2X1_LOC_158/A OR2X1_LOC_517/Y 0.08fF
C8967 OR2X1_LOC_158/A OR2X1_LOC_409/B 0.03fF
C9282 OR2X1_LOC_158/A OR2X1_LOC_497/Y 0.06fF
C10483 OR2X1_LOC_158/A AND2X1_LOC_198/a_36_24# 0.01fF
C10932 OR2X1_LOC_158/A OR2X1_LOC_96/B 0.03fF
C11212 OR2X1_LOC_158/A AND2X1_LOC_284/a_8_24# 0.04fF
C11768 OR2X1_LOC_158/A OR2X1_LOC_257/a_8_216# 0.02fF
C12107 OR2X1_LOC_158/A AND2X1_LOC_335/Y 0.01fF
C12185 OR2X1_LOC_158/A OR2X1_LOC_619/Y 0.21fF
C12644 OR2X1_LOC_158/A OR2X1_LOC_669/A 0.41fF
C12671 OR2X1_LOC_158/A AND2X1_LOC_454/A 0.04fF
C12673 OR2X1_LOC_158/A OR2X1_LOC_232/a_8_216# 0.07fF
C12940 OR2X1_LOC_158/A AND2X1_LOC_783/B 0.01fF
C13162 OR2X1_LOC_158/A AND2X1_LOC_473/a_8_24# 0.02fF
C14585 OR2X1_LOC_158/A OR2X1_LOC_13/B 1.19fF
C15073 OR2X1_LOC_158/A OR2X1_LOC_595/A 0.01fF
C15161 OR2X1_LOC_158/A AND2X1_LOC_154/a_8_24# 0.09fF
C15580 OR2X1_LOC_158/A AND2X1_LOC_342/Y 0.05fF
C15626 OR2X1_LOC_158/A OR2X1_LOC_279/a_8_216# 0.01fF
C15655 OR2X1_LOC_158/A AND2X1_LOC_712/B 0.29fF
C16052 OR2X1_LOC_158/A OR2X1_LOC_89/A 0.36fF
C16485 OR2X1_LOC_158/A OR2X1_LOC_282/Y 0.01fF
C16722 OR2X1_LOC_158/A AND2X1_LOC_473/Y 0.10fF
C16978 OR2X1_LOC_158/A AND2X1_LOC_727/A 0.03fF
C17253 OR2X1_LOC_179/Y OR2X1_LOC_158/A 0.01fF
C17679 OR2X1_LOC_158/A AND2X1_LOC_621/Y 0.02fF
C17692 OR2X1_LOC_158/A AND2X1_LOC_668/a_8_24# 0.14fF
C19345 OR2X1_LOC_158/A AND2X1_LOC_535/Y 0.03fF
C19758 OR2X1_LOC_158/A OR2X1_LOC_16/A 0.14fF
C19789 OR2X1_LOC_158/A OR2X1_LOC_108/Y 0.17fF
C20660 OR2X1_LOC_158/A OR2X1_LOC_380/Y 0.03fF
C20704 OR2X1_LOC_158/A OR2X1_LOC_109/Y 0.03fF
C20717 OR2X1_LOC_158/A AND2X1_LOC_448/Y 0.01fF
C21293 OR2X1_LOC_158/A AND2X1_LOC_227/Y 0.03fF
C21619 OR2X1_LOC_599/A OR2X1_LOC_158/A 0.03fF
C21645 OR2X1_LOC_158/A OR2X1_LOC_258/a_8_216# 0.20fF
C21989 OR2X1_LOC_158/A AND2X1_LOC_843/Y 0.02fF
C22171 OR2X1_LOC_158/A OR2X1_LOC_224/a_8_216# 0.05fF
C22324 OR2X1_LOC_158/A AND2X1_LOC_284/a_36_24# 0.01fF
C22496 OR2X1_LOC_158/A OR2X1_LOC_32/a_8_216# 0.03fF
C22787 AND2X1_LOC_707/Y OR2X1_LOC_158/A 0.11fF
C23385 OR2X1_LOC_158/A OR2X1_LOC_60/a_8_216# 0.01fF
C24213 OR2X1_LOC_158/A AND2X1_LOC_473/a_36_24# 0.01fF
C24492 OR2X1_LOC_158/A OR2X1_LOC_74/Y 0.03fF
C25760 OR2X1_LOC_158/A AND2X1_LOC_161/a_8_24# 0.01fF
C26124 OR2X1_LOC_158/A OR2X1_LOC_96/Y 0.01fF
C26691 OR2X1_LOC_158/A OR2X1_LOC_279/Y 0.09fF
C26999 OR2X1_LOC_158/A AND2X1_LOC_456/B 0.04fF
C28005 OR2X1_LOC_158/A AND2X1_LOC_116/B 0.02fF
C28048 OR2X1_LOC_158/A OR2X1_LOC_96/a_8_216# 0.01fF
C28216 OR2X1_LOC_158/A AND2X1_LOC_802/Y 0.03fF
C28382 OR2X1_LOC_158/A AND2X1_LOC_154/Y 0.04fF
C28643 OR2X1_LOC_158/A AND2X1_LOC_709/a_8_24# 0.01fF
C28729 OR2X1_LOC_158/A AND2X1_LOC_624/A 0.09fF
C29729 OR2X1_LOC_158/A AND2X1_LOC_114/Y 0.01fF
C29884 OR2X1_LOC_158/A OR2X1_LOC_312/a_8_216# 0.05fF
C29961 OR2X1_LOC_158/A AND2X1_LOC_335/a_36_24# 0.01fF
C29972 OR2X1_LOC_158/A OR2X1_LOC_837/A 0.03fF
C30008 OR2X1_LOC_158/A AND2X1_LOC_114/a_8_24# 0.02fF
C30360 OR2X1_LOC_158/A AND2X1_LOC_160/Y 0.02fF
C30503 OR2X1_LOC_158/A OR2X1_LOC_295/a_8_216# 0.01fF
C30735 OR2X1_LOC_158/A OR2X1_LOC_421/Y 1.04fF
C30933 OR2X1_LOC_158/A OR2X1_LOC_273/Y 0.01fF
C31157 OR2X1_LOC_158/A OR2X1_LOC_744/a_8_216# 0.01fF
C31737 OR2X1_LOC_158/A OR2X1_LOC_24/Y 0.03fF
C32858 OR2X1_LOC_604/A OR2X1_LOC_158/A 0.95fF
C33378 OR2X1_LOC_158/A OR2X1_LOC_265/Y 0.07fF
C33589 OR2X1_LOC_158/A OR2X1_LOC_163/A 0.04fF
C33874 OR2X1_LOC_158/A AND2X1_LOC_155/Y 0.17fF
C33923 OR2X1_LOC_158/A AND2X1_LOC_633/Y 0.02fF
C34085 AND2X1_LOC_539/Y OR2X1_LOC_158/A 0.03fF
C34136 OR2X1_LOC_158/A AND2X1_LOC_711/A 0.01fF
C34138 OR2X1_LOC_158/A AND2X1_LOC_326/B 0.03fF
C34224 OR2X1_LOC_158/A AND2X1_LOC_668/a_36_24# 0.01fF
C34472 OR2X1_LOC_316/a_8_216# OR2X1_LOC_158/A 0.02fF
C35016 OR2X1_LOC_158/A AND2X1_LOC_434/Y 0.07fF
C35232 OR2X1_LOC_158/A OR2X1_LOC_595/Y 0.01fF
C35438 OR2X1_LOC_158/A OR2X1_LOC_837/B 0.07fF
C35554 OR2X1_LOC_158/A AND2X1_LOC_260/a_8_24# 0.27fF
C36265 OR2X1_LOC_158/A OR2X1_LOC_837/Y 0.07fF
C36661 OR2X1_LOC_517/a_8_216# OR2X1_LOC_158/A 0.03fF
C36708 OR2X1_LOC_158/A AND2X1_LOC_161/a_36_24# 0.02fF
C37131 OR2X1_LOC_158/A AND2X1_LOC_520/Y 0.02fF
C37150 OR2X1_LOC_158/A AND2X1_LOC_848/Y 0.06fF
C37923 OR2X1_LOC_178/Y OR2X1_LOC_158/A 0.01fF
C38050 OR2X1_LOC_158/A OR2X1_LOC_258/Y 0.01fF
C38136 OR2X1_LOC_158/A AND2X1_LOC_318/Y 0.10fF
C38338 OR2X1_LOC_759/A OR2X1_LOC_158/A 0.04fF
C38356 OR2X1_LOC_158/A OR2X1_LOC_697/a_8_216# 0.07fF
C38368 OR2X1_LOC_158/A OR2X1_LOC_698/Y 0.02fF
C39198 OR2X1_LOC_158/A AND2X1_LOC_810/B 0.07fF
C39653 OR2X1_LOC_158/A AND2X1_LOC_709/a_36_24# -0.00fF
C40038 OR2X1_LOC_158/A AND2X1_LOC_715/A 0.06fF
C40555 AND2X1_LOC_729/Y OR2X1_LOC_158/A 0.07fF
C40587 AND2X1_LOC_784/A OR2X1_LOC_158/A 0.09fF
C41021 OR2X1_LOC_158/A OR2X1_LOC_52/B 0.74fF
C41038 OR2X1_LOC_158/A AND2X1_LOC_489/Y 0.14fF
C41314 OR2X1_LOC_158/A OR2X1_LOC_281/Y 0.01fF
C41353 OR2X1_LOC_158/A AND2X1_LOC_161/Y 0.01fF
C41446 OR2X1_LOC_158/A AND2X1_LOC_286/Y 0.04fF
C41484 OR2X1_LOC_158/A AND2X1_LOC_356/B 0.03fF
C41490 OR2X1_LOC_158/A OR2X1_LOC_280/Y 4.57fF
C42178 OR2X1_LOC_158/A OR2X1_LOC_744/Y 0.01fF
C42715 OR2X1_LOC_158/A OR2X1_LOC_58/a_8_216# 0.05fF
C42724 OR2X1_LOC_158/A OR2X1_LOC_16/Y 0.03fF
C43209 OR2X1_LOC_158/A OR2X1_LOC_423/a_8_216# 0.01fF
C44414 OR2X1_LOC_158/A AND2X1_LOC_197/Y 0.07fF
C44677 OR2X1_LOC_158/A OR2X1_LOC_163/a_8_216# 0.01fF
C44740 OR2X1_LOC_158/A OR2X1_LOC_183/Y 0.04fF
C45809 OR2X1_LOC_158/A OR2X1_LOC_669/Y 0.02fF
C45848 OR2X1_LOC_158/A OR2X1_LOC_27/Y 0.03fF
C46414 OR2X1_LOC_158/A AND2X1_LOC_116/a_8_24# 0.02fF
C46493 OR2X1_LOC_158/A OR2X1_LOC_423/Y 0.01fF
C46753 OR2X1_LOC_158/A OR2X1_LOC_74/A 1.31fF
C46777 OR2X1_LOC_158/A OR2X1_LOC_261/A 0.01fF
C47079 OR2X1_LOC_158/A AND2X1_LOC_162/a_8_24# 0.01fF
C47161 OR2X1_LOC_158/A AND2X1_LOC_287/Y 0.02fF
C47500 OR2X1_LOC_158/A AND2X1_LOC_448/a_8_24# 0.01fF
C48669 OR2X1_LOC_158/A OR2X1_LOC_521/a_8_216# 0.04fF
C48729 OR2X1_LOC_106/Y OR2X1_LOC_158/A 0.03fF
C49438 OR2X1_LOC_158/A AND2X1_LOC_319/a_8_24# 0.06fF
C49510 OR2X1_LOC_158/A OR2X1_LOC_72/Y 0.03fF
C50085 OR2X1_LOC_158/A AND2X1_LOC_198/a_8_24# 0.04fF
C50127 OR2X1_LOC_158/A OR2X1_LOC_595/a_8_216# 0.01fF
C50462 AND2X1_LOC_706/Y OR2X1_LOC_158/A 0.07fF
C50473 OR2X1_LOC_158/A OR2X1_LOC_58/Y 0.05fF
C51416 OR2X1_LOC_158/A OR2X1_LOC_32/Y 0.13fF
C52503 OR2X1_LOC_158/A OR2X1_LOC_743/Y 0.01fF
C52557 OR2X1_LOC_158/A AND2X1_LOC_285/a_8_24# 0.01fF
C52756 OR2X1_LOC_158/A OR2X1_LOC_295/Y 0.01fF
C53079 OR2X1_LOC_158/A OR2X1_LOC_433/Y 0.03fF
C53394 OR2X1_LOC_158/A AND2X1_LOC_714/B 0.03fF
C53877 OR2X1_LOC_158/A OR2X1_LOC_58/a_36_216# 0.01fF
C54885 OR2X1_LOC_158/A AND2X1_LOC_798/A 0.03fF
C55081 OR2X1_LOC_125/a_8_216# OR2X1_LOC_158/A 0.14fF
C55521 OR2X1_LOC_158/A VDD 1.56fF
C55634 OR2X1_LOC_158/A OR2X1_LOC_251/Y 0.02fF
C55835 OR2X1_LOC_158/A OR2X1_LOC_163/Y 0.09fF
C55965 OR2X1_LOC_158/A OR2X1_LOC_60/Y 0.01fF
C56066 OR2X1_LOC_158/A OR2X1_LOC_248/Y 0.01fF
C57839 OR2X1_LOC_158/A VSS 1.15fF
C29614 OR2X1_LOC_52/Y OR2X1_LOC_56/Y 0.05fF
C32978 AND2X1_LOC_197/a_8_24# OR2X1_LOC_56/Y 0.01fF
C40042 OR2X1_LOC_56/Y OR2X1_LOC_16/Y 0.15fF
C41782 AND2X1_LOC_197/Y OR2X1_LOC_56/Y 0.21fF
C47513 AND2X1_LOC_198/a_8_24# OR2X1_LOC_56/Y 0.01fF
C52972 VDD OR2X1_LOC_56/Y 0.33fF
C53001 AND2X1_LOC_208/B OR2X1_LOC_56/Y 0.01fF
C56759 OR2X1_LOC_56/Y VSS 0.04fF
C2923 OR2X1_LOC_45/B OR2X1_LOC_304/Y 0.09fF
C5596 OR2X1_LOC_431/Y OR2X1_LOC_304/Y 0.73fF
C8870 OR2X1_LOC_135/a_8_216# OR2X1_LOC_304/Y 0.01fF
C17443 OR2X1_LOC_45/Y OR2X1_LOC_304/Y 0.31fF
C37626 OR2X1_LOC_135/Y OR2X1_LOC_304/Y 0.23fF
C41665 OR2X1_LOC_304/Y OR2X1_LOC_52/B 0.06fF
C50811 OR2X1_LOC_431/a_8_216# OR2X1_LOC_304/Y 0.01fF
C56162 VDD OR2X1_LOC_304/Y 0.04fF
C57250 OR2X1_LOC_304/Y VSS -0.06fF
C13128 OR2X1_LOC_52/B OR2X1_LOC_421/Y 0.01fF
C15193 OR2X1_LOC_423/a_8_216# OR2X1_LOC_421/Y 0.44fF
C18396 OR2X1_LOC_421/Y OR2X1_LOC_423/Y 0.05fF
C19338 OR2X1_LOC_421/Y AND2X1_LOC_448/a_8_24# -0.00fF
C20757 OR2X1_LOC_423/a_36_216# OR2X1_LOC_421/Y 0.01fF
C27390 VDD OR2X1_LOC_421/Y 0.26fF
C30310 OR2X1_LOC_45/B OR2X1_LOC_421/Y 0.24fF
C35137 OR2X1_LOC_417/Y OR2X1_LOC_421/Y 0.03fF
C40097 OR2X1_LOC_619/Y OR2X1_LOC_421/Y 0.03fF
C40597 AND2X1_LOC_454/A OR2X1_LOC_421/Y 0.15fF
C43717 AND2X1_LOC_712/B OR2X1_LOC_421/Y 0.10fF
C48770 AND2X1_LOC_447/Y OR2X1_LOC_421/Y 0.03fF
C50814 OR2X1_LOC_421/Y OR2X1_LOC_424/Y 0.05fF
C50868 AND2X1_LOC_707/Y OR2X1_LOC_421/Y 1.30fF
C56520 OR2X1_LOC_421/Y VSS 0.18fF
C10018 OR2X1_LOC_329/Y VDD 0.17fF
C15638 OR2X1_LOC_329/Y AND2X1_LOC_390/B 0.02fF
C18584 OR2X1_LOC_329/Y AND2X1_LOC_436/B 0.02fF
C20962 OR2X1_LOC_329/Y OR2X1_LOC_331/Y 0.09fF
C24993 OR2X1_LOC_329/Y OR2X1_LOC_312/Y 0.02fF
C25198 OR2X1_LOC_329/Y OR2X1_LOC_13/B 0.03fF
C30330 OR2X1_LOC_329/Y OR2X1_LOC_16/A 0.04fF
C32106 OR2X1_LOC_329/Y OR2X1_LOC_599/A 0.85fF
C44775 AND2X1_LOC_539/Y OR2X1_LOC_329/Y 0.02fF
C45717 OR2X1_LOC_329/Y AND2X1_LOC_434/Y 0.07fF
C51396 AND2X1_LOC_729/Y OR2X1_LOC_329/Y 0.03fF
C52279 OR2X1_LOC_329/Y AND2X1_LOC_356/B 0.02fF
C57920 OR2X1_LOC_329/Y VSS 0.08fF
C733 OR2X1_LOC_597/A OR2X1_LOC_599/A 0.02fF
C57989 OR2X1_LOC_597/A VSS 0.29fF
C24751 OR2X1_LOC_385/Y OR2X1_LOC_387/Y 0.22fF
C41068 VDD OR2X1_LOC_387/Y 0.16fF
C41209 OR2X1_LOC_387/Y AND2X1_LOC_389/a_8_24# 0.23fF
C45061 OR2X1_LOC_387/Y OR2X1_LOC_586/Y 0.02fF
C57599 OR2X1_LOC_387/Y VSS -0.00fF
C4607 OR2X1_LOC_391/B OR2X1_LOC_392/A 0.05fF
C8101 OR2X1_LOC_391/B OR2X1_LOC_846/a_8_216# 0.09fF
C10212 OR2X1_LOC_391/B OR2X1_LOC_772/B 0.29fF
C10243 OR2X1_LOC_391/B OR2X1_LOC_489/B 0.03fF
C24693 OR2X1_LOC_391/B OR2X1_LOC_848/B 0.11fF
C26331 OR2X1_LOC_391/B OR2X1_LOC_773/B 0.04fF
C28549 OR2X1_LOC_391/B OR2X1_LOC_846/A 0.22fF
C37033 OR2X1_LOC_391/B OR2X1_LOC_557/a_8_216# 0.02fF
C42951 OR2X1_LOC_391/B OR2X1_LOC_846/B 0.28fF
C48352 OR2X1_LOC_391/B OR2X1_LOC_561/B 0.21fF
C49820 OR2X1_LOC_391/B OR2X1_LOC_391/a_8_216# 0.06fF
C55294 OR2X1_LOC_391/B OR2X1_LOC_489/a_8_216# 0.05fF
C57983 OR2X1_LOC_391/B VSS 0.33fF
C253 OR2X1_LOC_240/B OR2X1_LOC_549/A 0.03fF
C2922 OR2X1_LOC_240/A OR2X1_LOC_549/A 0.09fF
C2930 OR2X1_LOC_633/B OR2X1_LOC_549/A 0.01fF
C3659 OR2X1_LOC_633/a_8_216# OR2X1_LOC_549/A 0.03fF
C3772 AND2X1_LOC_122/a_8_24# OR2X1_LOC_549/A 0.01fF
C4971 AND2X1_LOC_117/a_8_24# OR2X1_LOC_549/A 0.03fF
C5744 OR2X1_LOC_240/a_8_216# OR2X1_LOC_549/A 0.40fF
C6897 OR2X1_LOC_777/B OR2X1_LOC_549/A 0.07fF
C7152 OR2X1_LOC_456/A OR2X1_LOC_549/A 0.01fF
C7888 OR2X1_LOC_630/B OR2X1_LOC_549/A 0.01fF
C10579 OR2X1_LOC_123/B OR2X1_LOC_549/A 0.04fF
C11271 AND2X1_LOC_498/a_8_24# OR2X1_LOC_549/A 0.01fF
C12523 OR2X1_LOC_151/A OR2X1_LOC_549/A 0.12fF
C13058 AND2X1_LOC_482/a_8_24# OR2X1_LOC_549/A 0.01fF
C13526 AND2X1_LOC_252/a_8_24# OR2X1_LOC_549/A 0.01fF
C13783 OR2X1_LOC_415/Y OR2X1_LOC_549/A 0.01fF
C13830 OR2X1_LOC_631/A OR2X1_LOC_549/A 0.01fF
C14817 AND2X1_LOC_122/a_36_24# OR2X1_LOC_549/A 0.01fF
C16857 OR2X1_LOC_243/A OR2X1_LOC_549/A 0.03fF
C17603 OR2X1_LOC_190/A OR2X1_LOC_549/A 0.07fF
C18000 OR2X1_LOC_188/Y OR2X1_LOC_549/A 0.03fF
C18492 AND2X1_LOC_131/a_8_24# OR2X1_LOC_549/A 0.03fF
C19462 OR2X1_LOC_810/A OR2X1_LOC_549/A 0.10fF
C19773 OR2X1_LOC_715/B OR2X1_LOC_549/A 0.31fF
C19776 AND2X1_LOC_626/a_8_24# OR2X1_LOC_549/A 0.02fF
C19910 AND2X1_LOC_81/a_8_24# OR2X1_LOC_549/A 0.02fF
C21534 OR2X1_LOC_78/A OR2X1_LOC_549/A 1.50fF
C22408 OR2X1_LOC_147/B OR2X1_LOC_549/A 0.07fF
C22798 OR2X1_LOC_121/Y OR2X1_LOC_549/A 0.39fF
C22948 AND2X1_LOC_496/a_8_24# OR2X1_LOC_549/A 0.01fF
C23324 AND2X1_LOC_495/a_8_24# OR2X1_LOC_549/A 0.02fF
C24049 OR2X1_LOC_140/A OR2X1_LOC_549/A 0.14fF
C24118 OR2X1_LOC_833/B OR2X1_LOC_549/A 0.02fF
C25285 OR2X1_LOC_629/B OR2X1_LOC_549/A 0.01fF
C26238 OR2X1_LOC_574/A OR2X1_LOC_549/A 0.10fF
C27840 OR2X1_LOC_499/B OR2X1_LOC_549/A 0.02fF
C29136 OR2X1_LOC_115/a_8_216# OR2X1_LOC_549/A 0.03fF
C29883 OR2X1_LOC_139/A OR2X1_LOC_549/A 0.10fF
C33817 OR2X1_LOC_154/A OR2X1_LOC_549/A 0.10fF
C34975 OR2X1_LOC_633/A OR2X1_LOC_549/A 0.17fF
C36236 OR2X1_LOC_124/B OR2X1_LOC_549/A -0.02fF
C37688 OR2X1_LOC_532/B OR2X1_LOC_549/A 0.20fF
C39643 VDD OR2X1_LOC_549/A 1.95fF
C41541 AND2X1_LOC_667/a_8_24# OR2X1_LOC_549/A 0.03fF
C41738 OR2X1_LOC_115/B OR2X1_LOC_549/A 0.11fF
C42255 OR2X1_LOC_216/A OR2X1_LOC_549/A 0.03fF
C42742 OR2X1_LOC_160/A OR2X1_LOC_549/A 0.14fF
C43029 OR2X1_LOC_130/Y OR2X1_LOC_549/A 0.03fF
C44020 OR2X1_LOC_185/A OR2X1_LOC_549/A 0.07fF
C44807 AND2X1_LOC_262/a_8_24# OR2X1_LOC_549/A 0.02fF
C45250 OR2X1_LOC_641/A OR2X1_LOC_549/A 0.07fF
C45356 OR2X1_LOC_114/Y OR2X1_LOC_549/A 0.04fF
C45760 OR2X1_LOC_541/B OR2X1_LOC_549/A 0.02fF
C46244 OR2X1_LOC_643/A OR2X1_LOC_549/A 0.07fF
C46541 AND2X1_LOC_91/B OR2X1_LOC_549/A 0.10fF
C46652 AND2X1_LOC_72/Y OR2X1_LOC_549/A 0.01fF
C47026 OR2X1_LOC_549/A OR2X1_LOC_719/B 0.02fF
C47058 OR2X1_LOC_542/B OR2X1_LOC_549/A 0.07fF
C47154 AND2X1_LOC_56/B OR2X1_LOC_549/A 0.44fF
C48063 AND2X1_LOC_118/a_8_24# OR2X1_LOC_549/A 0.01fF
C49121 OR2X1_LOC_549/B OR2X1_LOC_549/A 0.04fF
C50072 AND2X1_LOC_232/a_8_24# OR2X1_LOC_549/A 0.01fF
C50988 OR2X1_LOC_116/a_8_216# OR2X1_LOC_549/A 0.04fF
C51382 OR2X1_LOC_116/A OR2X1_LOC_549/A 0.04fF
C51631 OR2X1_LOC_771/B OR2X1_LOC_549/A 0.09fF
C52763 OR2X1_LOC_720/B OR2X1_LOC_549/A -0.02fF
C54611 OR2X1_LOC_549/a_8_216# OR2X1_LOC_549/A 0.02fF
C55960 OR2X1_LOC_786/A OR2X1_LOC_549/A 0.02fF
C56261 OR2X1_LOC_549/A VSS 0.61fF
C1009 OR2X1_LOC_78/A OR2X1_LOC_777/B 0.11fF
C1881 OR2X1_LOC_317/A OR2X1_LOC_777/B 0.13fF
C2076 OR2X1_LOC_318/B OR2X1_LOC_777/B 0.03fF
C2284 OR2X1_LOC_114/B OR2X1_LOC_777/B 0.06fF
C2306 OR2X1_LOC_538/A OR2X1_LOC_777/B 0.03fF
C3619 OR2X1_LOC_833/B OR2X1_LOC_777/B 0.07fF
C4763 OR2X1_LOC_629/B OR2X1_LOC_777/B 0.01fF
C5154 OR2X1_LOC_186/Y OR2X1_LOC_777/B 0.02fF
C7013 OR2X1_LOC_629/a_8_216# OR2X1_LOC_777/B 0.04fF
C10837 OR2X1_LOC_703/B OR2X1_LOC_777/B 0.06fF
C11989 OR2X1_LOC_97/A OR2X1_LOC_777/B 0.03fF
C12050 OR2X1_LOC_541/A OR2X1_LOC_777/B 0.03fF
C12455 OR2X1_LOC_777/B OR2X1_LOC_713/A 0.03fF
C13423 OR2X1_LOC_154/A OR2X1_LOC_777/B 0.10fF
C15154 AND2X1_LOC_600/a_8_24# OR2X1_LOC_777/B 0.03fF
C17287 OR2X1_LOC_532/B OR2X1_LOC_777/B 0.05fF
C19270 VDD OR2X1_LOC_777/B 0.99fF
C22350 OR2X1_LOC_160/A OR2X1_LOC_777/B 0.07fF
C23612 OR2X1_LOC_185/A OR2X1_LOC_777/B 0.03fF
C25273 OR2X1_LOC_541/B OR2X1_LOC_777/B 0.13fF
C25708 OR2X1_LOC_778/Y OR2X1_LOC_777/B 0.07fF
C25980 AND2X1_LOC_91/B OR2X1_LOC_777/B 0.09fF
C26328 OR2X1_LOC_777/B OR2X1_LOC_303/B 0.05fF
C26538 AND2X1_LOC_56/B OR2X1_LOC_777/B 0.05fF
C28496 OR2X1_LOC_777/B OR2X1_LOC_180/B 0.17fF
C28879 OR2X1_LOC_777/B OR2X1_LOC_788/B 0.03fF
C31434 OR2X1_LOC_777/B OR2X1_LOC_593/B 0.03fF
C33716 OR2X1_LOC_447/a_8_216# OR2X1_LOC_777/B 0.14fF
C35464 OR2X1_LOC_447/Y OR2X1_LOC_777/B 0.04fF
C36640 OR2X1_LOC_631/B OR2X1_LOC_777/B 0.07fF
C37898 OR2X1_LOC_169/B OR2X1_LOC_777/B 0.14fF
C44307 OR2X1_LOC_777/a_8_216# OR2X1_LOC_777/B 0.06fF
C45650 OR2X1_LOC_319/B OR2X1_LOC_777/B 0.07fF
C45715 OR2X1_LOC_296/Y OR2X1_LOC_777/B 0.03fF
C46617 OR2X1_LOC_629/A OR2X1_LOC_777/B 0.99fF
C48295 OR2X1_LOC_151/A OR2X1_LOC_777/B 0.14fF
C49912 OR2X1_LOC_168/Y OR2X1_LOC_777/B 0.19fF
C50749 OR2X1_LOC_777/B OR2X1_LOC_308/Y 0.03fF
C52548 AND2X1_LOC_314/a_8_24# OR2X1_LOC_777/B 0.17fF
C53569 OR2X1_LOC_777/B OR2X1_LOC_241/B 0.04fF
C53742 OR2X1_LOC_188/Y OR2X1_LOC_777/B 0.03fF
C54147 OR2X1_LOC_831/A OR2X1_LOC_777/B 0.03fF
C54565 OR2X1_LOC_777/B OR2X1_LOC_356/A 0.21fF
C56452 OR2X1_LOC_777/B VSS -0.62fF
C1505 AND2X1_LOC_232/a_8_24# OR2X1_LOC_633/A 0.03fF
C1929 OR2X1_LOC_235/B OR2X1_LOC_633/A 0.08fF
C7930 OR2X1_LOC_240/B OR2X1_LOC_633/A 0.01fF
C9905 OR2X1_LOC_633/A OR2X1_LOC_71/A 0.09fF
C10537 OR2X1_LOC_633/A OR2X1_LOC_240/A 0.01fF
C13472 OR2X1_LOC_240/a_8_216# OR2X1_LOC_633/A 0.03fF
C16127 OR2X1_LOC_673/A OR2X1_LOC_633/A 0.04fF
C18068 AND2X1_LOC_232/a_36_24# OR2X1_LOC_633/A 0.01fF
C19018 OR2X1_LOC_287/B OR2X1_LOC_633/A 0.05fF
C24503 OR2X1_LOC_243/A OR2X1_LOC_633/A 0.02fF
C28630 OR2X1_LOC_622/A OR2X1_LOC_633/A 0.03fF
C29065 OR2X1_LOC_78/A OR2X1_LOC_633/A 0.14fF
C39338 OR2X1_LOC_622/a_8_216# OR2X1_LOC_633/A 0.05fF
C45454 OR2X1_LOC_532/B OR2X1_LOC_633/A 0.87fF
C47496 VDD OR2X1_LOC_633/A 0.51fF
C51785 OR2X1_LOC_185/A OR2X1_LOC_633/A 0.10fF
C56551 OR2X1_LOC_633/A VSS 0.65fF
C2023 VDD OR2X1_LOC_541/B 0.30fF
C9403 AND2X1_LOC_56/B OR2X1_LOC_541/B 0.04fF
C19123 OR2X1_LOC_541/B OR2X1_LOC_541/a_8_216# 0.49fF
C30131 OR2X1_LOC_541/B OR2X1_LOC_553/A 0.01fF
C36156 OR2X1_LOC_541/B OR2X1_LOC_241/B 0.14fF
C36267 OR2X1_LOC_188/Y OR2X1_LOC_541/B 0.01fF
C42428 OR2X1_LOC_833/B OR2X1_LOC_541/B 0.02fF
C51020 OR2X1_LOC_541/A OR2X1_LOC_541/B 0.16fF
C56592 OR2X1_LOC_541/B VSS 0.25fF
C7983 OR2X1_LOC_634/A OR2X1_LOC_640/A 0.01fF
C10204 OR2X1_LOC_634/A OR2X1_LOC_240/A 0.12fF
C10827 OR2X1_LOC_634/A OR2X1_LOC_334/A 0.09fF
C17861 OR2X1_LOC_634/A AND2X1_LOC_825/a_8_24# 0.20fF
C23805 OR2X1_LOC_634/A AND2X1_LOC_89/a_8_24# 0.17fF
C26529 OR2X1_LOC_634/A AND2X1_LOC_416/a_8_24# 0.01fF
C28717 OR2X1_LOC_634/A OR2X1_LOC_78/A 0.70fF
C29238 OR2X1_LOC_634/A OR2X1_LOC_97/B 0.06fF
C32853 OR2X1_LOC_634/A OR2X1_LOC_338/A 0.02fF
C36865 OR2X1_LOC_634/A AND2X1_LOC_27/a_8_24# 0.17fF
C42486 OR2X1_LOC_634/A OR2X1_LOC_34/B 0.13fF
C46408 OR2X1_LOC_472/B OR2X1_LOC_634/A 0.33fF
C47113 VDD OR2X1_LOC_634/A 0.64fF
C47607 OR2X1_LOC_634/A OR2X1_LOC_334/B 0.08fF
C48109 OR2X1_LOC_462/B OR2X1_LOC_634/A 0.05fF
C53098 OR2X1_LOC_634/A OR2X1_LOC_634/a_8_216# 0.01fF
C54408 OR2X1_LOC_634/A AND2X1_LOC_56/B 0.02fF
C57455 OR2X1_LOC_634/A VSS 0.38fF
C3678 OR2X1_LOC_185/A OR2X1_LOC_266/A 0.01fF
C6039 AND2X1_LOC_91/B OR2X1_LOC_266/A 0.22fF
C10006 OR2X1_LOC_235/B OR2X1_LOC_266/A 0.06fF
C15456 OR2X1_LOC_786/A OR2X1_LOC_266/A 0.17fF
C17912 OR2X1_LOC_266/A OR2X1_LOC_71/A 0.14fF
C27448 OR2X1_LOC_266/a_8_216# OR2X1_LOC_266/A 0.18fF
C38451 AND2X1_LOC_79/Y OR2X1_LOC_266/A 0.07fF
C44886 OR2X1_LOC_673/Y OR2X1_LOC_266/A 0.02fF
C50256 AND2X1_LOC_813/a_8_24# OR2X1_LOC_266/A 0.01fF
C55507 VDD OR2X1_LOC_266/A 0.08fF
C55755 OR2X1_LOC_845/A OR2X1_LOC_266/A 1.12fF
C56719 OR2X1_LOC_266/A VSS -0.20fF
C655 OR2X1_LOC_139/A OR2X1_LOC_130/A 0.07fF
C1342 AND2X1_LOC_589/a_36_24# OR2X1_LOC_130/A 0.01fF
C3276 OR2X1_LOC_97/A OR2X1_LOC_130/A 0.12fF
C3396 OR2X1_LOC_130/A OR2X1_LOC_475/B 0.03fF
C4653 OR2X1_LOC_154/A OR2X1_LOC_130/A 0.17fF
C5151 AND2X1_LOC_821/a_8_24# OR2X1_LOC_130/A 0.13fF
C5923 OR2X1_LOC_520/Y OR2X1_LOC_130/A 0.05fF
C6652 OR2X1_LOC_130/A OR2X1_LOC_776/Y 0.19fF
C6868 OR2X1_LOC_130/A OR2X1_LOC_227/a_8_216# 0.03fF
C7519 OR2X1_LOC_653/B OR2X1_LOC_130/A 0.01fF
C8149 OR2X1_LOC_130/A OR2X1_LOC_33/B 0.02fF
C8658 OR2X1_LOC_130/A OR2X1_LOC_532/B 0.21fF
C9639 OR2X1_LOC_130/A AND2X1_LOC_224/a_8_24# 0.03fF
C9972 OR2X1_LOC_130/A AND2X1_LOC_432/a_8_24# 0.03fF
C10545 VDD OR2X1_LOC_130/A 1.43fF
C11501 OR2X1_LOC_462/B OR2X1_LOC_130/A 0.52fF
C13625 OR2X1_LOC_160/A OR2X1_LOC_130/A 9.11fF
C14871 OR2X1_LOC_185/A OR2X1_LOC_130/A 0.23fF
C16017 OR2X1_LOC_130/A OR2X1_LOC_641/A 0.07fF
C16108 OR2X1_LOC_379/Y OR2X1_LOC_130/A 0.03fF
C16244 AND2X1_LOC_821/a_36_24# OR2X1_LOC_130/A 0.01fF
C17021 OR2X1_LOC_643/A OR2X1_LOC_130/A 0.07fF
C17396 OR2X1_LOC_799/A OR2X1_LOC_130/A 0.02fF
C17838 AND2X1_LOC_56/B OR2X1_LOC_130/A 0.07fF
C19560 OR2X1_LOC_506/A OR2X1_LOC_130/A 0.11fF
C19701 OR2X1_LOC_130/A OR2X1_LOC_227/Y -0.00fF
C20687 OR2X1_LOC_130/A OR2X1_LOC_227/B 0.02fF
C25053 OR2X1_LOC_231/A OR2X1_LOC_130/A 0.06fF
C30520 AND2X1_LOC_586/a_8_24# OR2X1_LOC_130/A 0.11fF
C31667 OR2X1_LOC_130/A AND2X1_LOC_224/a_36_24# 0.01fF
C33929 OR2X1_LOC_493/A OR2X1_LOC_130/A 0.51fF
C34271 OR2X1_LOC_435/B OR2X1_LOC_130/A 0.02fF
C34855 OR2X1_LOC_130/A AND2X1_LOC_67/Y 0.08fF
C35608 OR2X1_LOC_130/A AND2X1_LOC_230/a_8_24# 0.14fF
C39289 OR2X1_LOC_318/A OR2X1_LOC_130/A 0.03fF
C39312 OR2X1_LOC_151/A OR2X1_LOC_130/A 0.07fF
C41701 OR2X1_LOC_130/A AND2X1_LOC_109/a_8_24# 0.03fF
C42814 AND2X1_LOC_24/a_8_24# OR2X1_LOC_130/A 0.14fF
C43178 OR2X1_LOC_130/A OR2X1_LOC_390/A 0.01fF
C44017 AND2X1_LOC_229/a_8_24# OR2X1_LOC_130/A 0.04fF
C46417 OR2X1_LOC_810/A OR2X1_LOC_130/A 0.07fF
C46429 AND2X1_LOC_589/a_8_24# OR2X1_LOC_130/A 0.03fF
C46692 OR2X1_LOC_715/B OR2X1_LOC_130/A 0.10fF
C48190 OR2X1_LOC_835/B OR2X1_LOC_130/A 0.04fF
C48450 AND2X1_LOC_432/a_36_24# OR2X1_LOC_130/A 0.01fF
C48521 OR2X1_LOC_130/A OR2X1_LOC_78/A 0.12fF
C49699 OR2X1_LOC_231/B OR2X1_LOC_130/A 0.02fF
C50549 OR2X1_LOC_318/a_8_216# OR2X1_LOC_130/A 0.05fF
C52611 OR2X1_LOC_130/A OR2X1_LOC_338/A 0.02fF
C52922 OR2X1_LOC_130/A OR2X1_LOC_112/B 0.04fF
C53976 AND2X1_LOC_24/a_36_24# OR2X1_LOC_130/A 0.01fF
C57081 OR2X1_LOC_130/A VSS 0.75fF
C380 OR2X1_LOC_154/A AND2X1_LOC_173/a_8_24# 0.06fF
C763 OR2X1_LOC_154/A OR2X1_LOC_235/B -0.03fF
C855 OR2X1_LOC_154/A AND2X1_LOC_393/a_8_24# 0.14fF
C1601 OR2X1_LOC_154/A OR2X1_LOC_362/A 0.07fF
C1667 OR2X1_LOC_539/A OR2X1_LOC_154/A 0.01fF
C1915 OR2X1_LOC_154/A OR2X1_LOC_771/B 0.14fF
C2779 OR2X1_LOC_154/A OR2X1_LOC_317/B 0.03fF
C3338 AND2X1_LOC_595/a_36_24# OR2X1_LOC_154/A 0.01fF
C3481 OR2X1_LOC_154/A AND2X1_LOC_69/Y 0.02fF
C4221 OR2X1_LOC_154/A AND2X1_LOC_394/a_8_24# 0.20fF
C4317 OR2X1_LOC_154/A AND2X1_LOC_79/a_36_24# 0.01fF
C4322 OR2X1_LOC_154/A AND2X1_LOC_69/a_8_24# 0.01fF
C4582 OR2X1_LOC_154/A AND2X1_LOC_65/a_8_24# 0.03fF
C4634 OR2X1_LOC_154/A OR2X1_LOC_447/a_8_216# 0.04fF
C5076 OR2X1_LOC_154/A OR2X1_LOC_449/B 0.07fF
C5893 OR2X1_LOC_154/A OR2X1_LOC_175/B 0.02fF
C6177 OR2X1_LOC_154/A OR2X1_LOC_389/a_8_216# 0.01fF
C6332 OR2X1_LOC_154/A OR2X1_LOC_400/B 0.02fF
C6422 OR2X1_LOC_154/A OR2X1_LOC_447/Y 0.45fF
C6617 OR2X1_LOC_709/B OR2X1_LOC_154/A 0.01fF
C7666 OR2X1_LOC_154/A OR2X1_LOC_631/B 0.03fF
C8318 OR2X1_LOC_154/A OR2X1_LOC_704/a_8_216# 0.04fF
C8518 OR2X1_LOC_154/A OR2X1_LOC_105/Y 0.01fF
C10071 OR2X1_LOC_154/a_8_216# OR2X1_LOC_154/A 0.04fF
C10157 OR2X1_LOC_154/A OR2X1_LOC_630/Y 0.10fF
C10941 OR2X1_LOC_154/A AND2X1_LOC_313/a_8_24# 0.02fF
C11253 OR2X1_LOC_154/A OR2X1_LOC_537/a_8_216# 0.03fF
C11316 OR2X1_LOC_154/A AND2X1_LOC_60/a_8_24# 0.04fF
C11838 OR2X1_LOC_154/A OR2X1_LOC_768/A 0.01fF
C12200 OR2X1_LOC_709/a_8_216# OR2X1_LOC_154/A 0.04fF
C12769 OR2X1_LOC_154/A OR2X1_LOC_539/Y 0.06fF
C13168 OR2X1_LOC_154/A OR2X1_LOC_678/Y 0.02fF
C13459 OR2X1_LOC_188/a_8_216# OR2X1_LOC_154/A 0.05fF
C13834 OR2X1_LOC_154/A OR2X1_LOC_332/a_8_216# 0.05fF
C14532 OR2X1_LOC_154/A AND2X1_LOC_67/Y 0.03fF
C14894 OR2X1_LOC_539/a_8_216# OR2X1_LOC_154/A 0.05fF
C15284 OR2X1_LOC_154/A OR2X1_LOC_400/A 0.06fF
C15392 OR2X1_LOC_154/A AND2X1_LOC_106/a_8_24# 0.04fF
C15646 OR2X1_LOC_154/A OR2X1_LOC_201/A 0.01fF
C16634 OR2X1_LOC_154/A OR2X1_LOC_436/a_8_216# 0.05fF
C16939 OR2X1_LOC_154/A AND2X1_LOC_103/a_8_24# -0.04fF
C17691 OR2X1_LOC_709/a_36_216# OR2X1_LOC_154/A 0.01fF
C17952 OR2X1_LOC_154/A OR2X1_LOC_436/Y 0.03fF
C19007 OR2X1_LOC_154/A OR2X1_LOC_151/A 0.17fF
C19332 OR2X1_LOC_154/A OR2X1_LOC_714/A 0.03fF
C19504 OR2X1_LOC_154/A OR2X1_LOC_174/A 0.01fF
C21531 OR2X1_LOC_154/A OR2X1_LOC_308/Y 0.07fF
C21767 OR2X1_LOC_154/A AND2X1_LOC_516/a_8_24# 0.01fF
C22433 OR2X1_LOC_154/A OR2X1_LOC_61/A 0.04fF
C22906 OR2X1_LOC_154/A OR2X1_LOC_390/A 0.04fF
C23303 OR2X1_LOC_711/B OR2X1_LOC_154/A 0.12fF
C23969 OR2X1_LOC_154/A OR2X1_LOC_84/A 0.43fF
C24328 OR2X1_LOC_154/A OR2X1_LOC_473/Y 0.03fF
C24390 OR2X1_LOC_154/A OR2X1_LOC_241/B 0.13fF
C24630 OR2X1_LOC_154/A AND2X1_LOC_423/a_8_24# 0.01fF
C24873 OR2X1_LOC_154/A OR2X1_LOC_339/A 0.01fF
C24904 OR2X1_LOC_208/A OR2X1_LOC_154/A 0.02fF
C25076 OR2X1_LOC_154/A OR2X1_LOC_537/A 0.01fF
C25343 OR2X1_LOC_154/A OR2X1_LOC_138/a_8_216# 0.06fF
C25447 OR2X1_LOC_154/A AND2X1_LOC_39/a_8_24# 0.04fF
C25935 OR2X1_LOC_154/A OR2X1_LOC_810/A 0.18fF
C26219 OR2X1_LOC_715/B OR2X1_LOC_154/A 0.10fF
C26449 OR2X1_LOC_154/A AND2X1_LOC_106/a_36_24# 0.01fF
C26490 OR2X1_LOC_154/A OR2X1_LOC_398/Y 0.05fF
C26710 OR2X1_LOC_154/A AND2X1_LOC_65/a_36_24# 0.01fF
C27212 OR2X1_LOC_154/A OR2X1_LOC_687/Y 0.07fF
C27949 OR2X1_LOC_154/A OR2X1_LOC_78/A 0.20fF
C29184 OR2X1_LOC_154/A OR2X1_LOC_114/B 0.05fF
C29219 OR2X1_LOC_154/A OR2X1_LOC_538/A 0.03fF
C29337 OR2X1_LOC_154/A AND2X1_LOC_79/Y 0.03fF
C29348 OR2X1_LOC_154/A AND2X1_LOC_496/a_8_24# 0.34fF
C30103 OR2X1_LOC_154/A OR2X1_LOC_623/B 0.07fF
C32280 OR2X1_LOC_154/A OR2X1_LOC_196/B 0.34fF
C32710 OR2X1_LOC_154/A OR2X1_LOC_574/A 0.11fF
C33287 OR2X1_LOC_154/A OR2X1_LOC_539/B 0.07fF
C33726 OR2X1_LOC_154/A OR2X1_LOC_515/Y 0.36fF
C34277 OR2X1_LOC_154/A OR2X1_LOC_499/B 0.04fF
C35570 OR2X1_LOC_154/A AND2X1_LOC_316/a_8_24# 0.02fF
C35633 OR2X1_LOC_154/A OR2X1_LOC_673/Y 0.01fF
C36297 OR2X1_LOC_154/A OR2X1_LOC_139/A 12.45fF
C36702 OR2X1_LOC_154/A OR2X1_LOC_138/A 0.02fF
C37172 AND2X1_LOC_595/a_8_24# OR2X1_LOC_154/A 0.04fF
C37920 OR2X1_LOC_154/A OR2X1_LOC_844/B 0.05fF
C38028 OR2X1_LOC_154/A OR2X1_LOC_389/A 0.02fF
C38160 OR2X1_LOC_154/A OR2X1_LOC_403/B 0.05fF
C38522 OR2X1_LOC_154/A OR2X1_LOC_61/B 0.33fF
C38859 OR2X1_LOC_154/A OR2X1_LOC_97/A 0.03fF
C38954 OR2X1_LOC_154/A OR2X1_LOC_541/A 0.05fF
C39436 OR2X1_LOC_154/A OR2X1_LOC_249/a_8_216# 0.17fF
C39978 OR2X1_LOC_154/A OR2X1_LOC_590/a_8_216# 0.01fF
C41784 OR2X1_LOC_154/A OR2X1_LOC_590/Y 0.04fF
C43843 OR2X1_LOC_154/A AND2X1_LOC_79/a_8_24# 0.07fF
C44050 OR2X1_LOC_154/A OR2X1_LOC_113/B 0.01fF
C44288 OR2X1_LOC_154/A OR2X1_LOC_532/B 0.33fF
C45386 OR2X1_LOC_710/B OR2X1_LOC_154/A 0.03fF
C45991 OR2X1_LOC_154/A AND2X1_LOC_496/a_36_24# 0.06fF
C46265 OR2X1_LOC_154/A VDD 2.40fF
C47187 OR2X1_LOC_154/A OR2X1_LOC_676/Y 0.03fF
C47514 OR2X1_LOC_154/A AND2X1_LOC_591/a_8_24# 0.02fF
C47599 OR2X1_LOC_154/A AND2X1_LOC_83/a_8_24# 0.04fF
C48414 OR2X1_LOC_154/A OR2X1_LOC_115/B 0.01fF
C48549 OR2X1_LOC_154/A OR2X1_LOC_840/A 0.17fF
C49012 OR2X1_LOC_154/A AND2X1_LOC_385/a_8_24# 0.01fF
C49410 OR2X1_LOC_154/A OR2X1_LOC_160/A 0.27fF
C49486 OR2X1_LOC_154/A OR2X1_LOC_624/B 1.02fF
C49839 OR2X1_LOC_154/A OR2X1_LOC_447/A 0.02fF
C50100 OR2X1_LOC_113/a_8_216# OR2X1_LOC_154/A 0.04fF
C50207 OR2X1_LOC_154/A OR2X1_LOC_78/Y 0.02fF
C50694 OR2X1_LOC_154/A OR2X1_LOC_185/A 0.03fF
C50703 OR2X1_LOC_154/A OR2X1_LOC_249/Y -0.02fF
C51142 OR2X1_LOC_154/A OR2X1_LOC_702/A 0.10fF
C52355 OR2X1_LOC_154/A AND2X1_LOC_617/a_8_24# 0.10fF
C52586 OR2X1_LOC_154/A AND2X1_LOC_238/a_8_24# 0.02fF
C52751 OR2X1_LOC_154/A OR2X1_LOC_436/B 0.01fF
C52816 OR2X1_LOC_154/A OR2X1_LOC_643/A 0.07fF
C52824 OR2X1_LOC_154/A OR2X1_LOC_778/Y 0.26fF
C52886 OR2X1_LOC_154/A OR2X1_LOC_113/A 0.03fF
C53053 AND2X1_LOC_91/B OR2X1_LOC_154/A 0.43fF
C53180 OR2X1_LOC_154/A AND2X1_LOC_39/a_36_24# 0.01fF
C53679 OR2X1_LOC_154/A AND2X1_LOC_56/B 0.49fF
C54480 OR2X1_LOC_154/A OR2X1_LOC_389/B 0.14fF
C55309 OR2X1_LOC_154/A OR2X1_LOC_506/A 0.03fF
C57980 OR2X1_LOC_154/A VSS -10.29fF
C1093 OR2X1_LOC_160/A OR2X1_LOC_115/B 0.15fF
C1234 OR2X1_LOC_160/A OR2X1_LOC_840/A 0.10fF
C1645 OR2X1_LOC_160/A OR2X1_LOC_216/A 0.01fF
C1714 OR2X1_LOC_160/A OR2X1_LOC_802/Y 0.03fF
C2185 OR2X1_LOC_160/A AND2X1_LOC_86/B 0.01fF
C2349 OR2X1_LOC_160/A OR2X1_LOC_532/Y 0.03fF
C2676 OR2X1_LOC_160/A AND2X1_LOC_127/a_8_24# 0.05fF
C2961 OR2X1_LOC_160/A AND2X1_LOC_424/a_8_24# 0.02fF
C3364 OR2X1_LOC_160/A OR2X1_LOC_114/a_36_216# 0.01fF
C3410 OR2X1_LOC_160/A OR2X1_LOC_185/A 0.31fF
C4503 OR2X1_LOC_160/A OR2X1_LOC_641/A 0.03fF
C4605 OR2X1_LOC_379/Y OR2X1_LOC_160/A 0.16fF
C4650 OR2X1_LOC_160/A OR2X1_LOC_114/Y 0.04fF
C4658 OR2X1_LOC_160/A OR2X1_LOC_449/A 0.01fF
C5474 OR2X1_LOC_160/A OR2X1_LOC_643/A 0.07fF
C5483 OR2X1_LOC_160/A OR2X1_LOC_778/Y 0.10fF
C5557 OR2X1_LOC_160/A OR2X1_LOC_113/A 0.05fF
C5703 AND2X1_LOC_91/B OR2X1_LOC_160/A 0.37fF
C5898 OR2X1_LOC_160/A OR2X1_LOC_799/A 0.05fF
C5995 OR2X1_LOC_160/A AND2X1_LOC_698/a_36_24# 0.01fF
C6312 OR2X1_LOC_160/A AND2X1_LOC_56/B 1.56fF
C7885 OR2X1_LOC_160/A OR2X1_LOC_186/a_8_216# 0.04fF
C7968 OR2X1_LOC_160/A OR2X1_LOC_646/B 0.11fF
C8068 OR2X1_LOC_160/A OR2X1_LOC_506/A 0.10fF
C8205 OR2X1_LOC_160/A OR2X1_LOC_780/A 0.01fF
C8575 OR2X1_LOC_160/A OR2X1_LOC_99/Y 0.03fF
C9206 OR2X1_LOC_160/A OR2X1_LOC_227/B 0.01fF
C9735 OR2X1_LOC_160/A OR2X1_LOC_235/B 0.19fF
C10207 AND2X1_LOC_380/a_8_24# OR2X1_LOC_160/A 0.03fF
C10517 OR2X1_LOC_160/A OR2X1_LOC_362/A 0.15fF
C10712 OR2X1_LOC_160/A AND2X1_LOC_680/a_8_24# 0.04fF
C10735 OR2X1_LOC_160/A OR2X1_LOC_243/B 0.95fF
C10833 OR2X1_LOC_160/A OR2X1_LOC_771/B 0.05fF
C10986 OR2X1_LOC_160/A OR2X1_LOC_637/B 0.25fF
C11286 OR2X1_LOC_156/a_8_216# OR2X1_LOC_160/A 0.02fF
C11447 OR2X1_LOC_160/A AND2X1_LOC_492/a_8_24# 0.11fF
C11666 OR2X1_LOC_160/A OR2X1_LOC_317/B 0.01fF
C12715 OR2X1_LOC_160/A OR2X1_LOC_473/a_8_216# 0.06fF
C13558 OR2X1_LOC_160/A AND2X1_LOC_65/a_8_24# 0.01fF
C13590 OR2X1_LOC_160/A OR2X1_LOC_231/A 0.03fF
C14052 OR2X1_LOC_160/A OR2X1_LOC_128/A 0.05fF
C14088 OR2X1_LOC_160/A OR2X1_LOC_449/B 0.07fF
C14408 OR2X1_LOC_317/a_8_216# OR2X1_LOC_160/A 0.02fF
C15369 OR2X1_LOC_160/A OR2X1_LOC_447/Y 0.03fF
C17314 AND2X1_LOC_764/a_8_24# OR2X1_LOC_160/A 0.02fF
C17568 OR2X1_LOC_160/A OR2X1_LOC_71/A 0.04fF
C17669 OR2X1_LOC_160/A OR2X1_LOC_355/a_8_216# 0.03fF
C18318 OR2X1_LOC_160/A OR2X1_LOC_633/B 0.14fF
C18955 OR2X1_LOC_154/a_8_216# OR2X1_LOC_160/A 0.02fF
C19551 OR2X1_LOC_160/A OR2X1_LOC_128/B 0.02fF
C19885 OR2X1_LOC_160/A OR2X1_LOC_730/A 0.02fF
C20365 OR2X1_LOC_160/A OR2X1_LOC_330/Y 0.02fF
C21710 OR2X1_LOC_160/A OR2X1_LOC_539/Y 0.07fF
C22394 OR2X1_LOC_156/Y OR2X1_LOC_160/A 0.15fF
C22566 OR2X1_LOC_160/A OR2X1_LOC_493/A 0.11fF
C22954 OR2X1_LOC_160/A OR2X1_LOC_435/B 0.07fF
C23480 OR2X1_LOC_160/A AND2X1_LOC_67/Y 0.39fF
C23755 OR2X1_LOC_160/A OR2X1_LOC_520/a_8_216# 0.05fF
C23983 OR2X1_LOC_160/A OR2X1_LOC_705/B 0.03fF
C24257 OR2X1_LOC_160/A AND2X1_LOC_230/a_8_24# 0.01fF
C24600 OR2X1_LOC_160/A OR2X1_LOC_201/A 0.01fF
C24705 OR2X1_LOC_160/A OR2X1_LOC_647/B 0.07fF
C25853 OR2X1_LOC_160/A AND2X1_LOC_331/a_8_24# 0.02fF
C26417 OR2X1_LOC_160/A OR2X1_LOC_446/Y 0.06fF
C26669 OR2X1_LOC_160/A AND2X1_LOC_320/a_8_24# 0.15fF
C26860 OR2X1_LOC_160/A OR2X1_LOC_436/Y 0.03fF
C27862 OR2X1_LOC_160/A OR2X1_LOC_318/A 0.11fF
C27883 OR2X1_LOC_160/A OR2X1_LOC_151/A 0.70fF
C28369 OR2X1_LOC_769/A OR2X1_LOC_160/A 0.02fF
C29166 OR2X1_LOC_160/A OR2X1_LOC_631/A 0.11fF
C29793 OR2X1_LOC_160/A OR2X1_LOC_520/B 0.12fF
C29851 OR2X1_LOC_160/A AND2X1_LOC_497/a_8_24# 0.04fF
C29971 OR2X1_LOC_156/B OR2X1_LOC_160/A 0.01fF
C30238 OR2X1_LOC_160/A OR2X1_LOC_783/A 0.03fF
C30349 OR2X1_LOC_160/A OR2X1_LOC_308/Y 0.04fF
C30987 OR2X1_LOC_160/A OR2X1_LOC_835/A 0.02fF
C32072 OR2X1_LOC_711/B OR2X1_LOC_160/A 0.34fF
C32131 OR2X1_LOC_160/A OR2X1_LOC_324/B 0.10fF
C32177 OR2X1_LOC_160/A AND2X1_LOC_314/a_8_24# 0.01fF
C32471 AND2X1_LOC_229/a_8_24# OR2X1_LOC_160/A 0.04fF
C32771 OR2X1_LOC_160/A OR2X1_LOC_84/A 0.27fF
C33141 OR2X1_LOC_160/A OR2X1_LOC_473/Y 0.05fF
C34198 OR2X1_LOC_160/A OR2X1_LOC_356/A 0.01fF
C34397 OR2X1_LOC_160/A AND2X1_LOC_698/a_8_24# 0.03fF
C34806 OR2X1_LOC_160/A OR2X1_LOC_810/A 8.93fF
C35061 OR2X1_LOC_715/B OR2X1_LOC_160/A 0.21fF
C35314 OR2X1_LOC_160/A OR2X1_LOC_398/Y 0.04fF
C36035 OR2X1_LOC_160/A OR2X1_LOC_687/Y 0.03fF
C36105 OR2X1_LOC_160/A OR2X1_LOC_606/Y 0.03fF
C36440 OR2X1_LOC_160/A OR2X1_LOC_835/B 0.16fF
C36750 OR2X1_LOC_160/A OR2X1_LOC_78/A 0.40fF
C37619 OR2X1_LOC_160/A OR2X1_LOC_501/B 0.09fF
C37678 OR2X1_LOC_160/A OR2X1_LOC_317/A 0.02fF
C37961 OR2X1_LOC_231/B OR2X1_LOC_160/A 0.04fF
C37972 OR2X1_LOC_121/Y OR2X1_LOC_160/A 0.07fF
C38001 OR2X1_LOC_160/A OR2X1_LOC_114/B 0.01fF
C38040 OR2X1_LOC_160/A OR2X1_LOC_538/A 0.03fF
C38970 OR2X1_LOC_160/A OR2X1_LOC_623/B 0.10fF
C39346 AND2X1_LOC_764/a_36_24# OR2X1_LOC_160/A 0.01fF
C39469 OR2X1_LOC_160/A OR2X1_LOC_646/A 0.03fF
C40226 OR2X1_LOC_160/A OR2X1_LOC_448/Y 0.02fF
C40922 OR2X1_LOC_160/A OR2X1_LOC_338/A 0.07fF
C40948 OR2X1_LOC_186/Y OR2X1_LOC_160/A 0.05fF
C41611 OR2X1_LOC_160/A OR2X1_LOC_574/A 0.26fF
C42806 OR2X1_LOC_160/A OR2X1_LOC_113/Y 0.01fF
C44312 OR2X1_LOC_160/A OR2X1_LOC_330/a_8_216# 0.01fF
C44618 OR2X1_LOC_160/A OR2X1_LOC_673/Y 0.01fF
C45303 OR2X1_LOC_160/A OR2X1_LOC_139/A 0.03fF
C45664 OR2X1_LOC_160/A OR2X1_LOC_728/A 0.05fF
C46606 OR2X1_LOC_160/A AND2X1_LOC_235/a_8_24# 0.01fF
C47053 OR2X1_LOC_160/A OR2X1_LOC_844/B 0.02fF
C47492 OR2X1_LOC_160/A OR2X1_LOC_532/a_8_216# 0.05fF
C47519 OR2X1_LOC_160/A OR2X1_LOC_130/a_8_216# 0.04fF
C47986 OR2X1_LOC_160/A OR2X1_LOC_97/A 0.06fF
C48087 AND2X1_LOC_744/a_8_24# OR2X1_LOC_160/A 0.04fF
C48118 OR2X1_LOC_160/A OR2X1_LOC_475/B 0.03fF
C48739 OR2X1_LOC_160/A OR2X1_LOC_546/A 0.16fF
C49123 OR2X1_LOC_160/A OR2X1_LOC_160/a_8_216# 0.18fF
C50701 OR2X1_LOC_160/A OR2X1_LOC_520/Y 0.03fF
C51405 OR2X1_LOC_160/A OR2X1_LOC_776/Y 0.07fF
C51580 OR2X1_LOC_160/A OR2X1_LOC_227/a_8_216# 0.01fF
C51781 OR2X1_LOC_160/A OR2X1_LOC_355/A 0.02fF
C53292 OR2X1_LOC_160/A OR2X1_LOC_532/B 0.98fF
C53908 OR2X1_LOC_160/A OR2X1_LOC_729/a_8_216# 0.03fF
C53965 OR2X1_LOC_160/A OR2X1_LOC_114/a_8_216# 0.02fF
C54261 OR2X1_LOC_160/A AND2X1_LOC_224/a_8_24# 0.01fF
C55209 OR2X1_LOC_160/A VDD 1.90fF
C55345 OR2X1_LOC_160/A OR2X1_LOC_836/B 0.01fF
C55670 OR2X1_LOC_160/A OR2X1_LOC_334/B 0.14fF
C56204 OR2X1_LOC_160/A OR2X1_LOC_462/B 0.03fF
C57941 OR2X1_LOC_160/A VSS 0.58fF
C2237 AND2X1_LOC_86/B OR2X1_LOC_624/B 0.07fF
C3003 AND2X1_LOC_86/B OR2X1_LOC_78/Y 0.03fF
C3451 OR2X1_LOC_185/A AND2X1_LOC_86/B 0.01fF
C5080 AND2X1_LOC_86/B AND2X1_LOC_617/a_8_24# 0.03fF
C5756 AND2X1_LOC_91/B AND2X1_LOC_86/B 0.01fF
C9793 OR2X1_LOC_235/B AND2X1_LOC_86/B 0.02fF
C17604 AND2X1_LOC_86/B OR2X1_LOC_71/A 0.08fF
C26827 OR2X1_LOC_287/B AND2X1_LOC_86/B 0.03fF
C53324 AND2X1_LOC_86/B OR2X1_LOC_532/B 0.03fF
C55270 VDD AND2X1_LOC_86/B 0.48fF
C57589 AND2X1_LOC_86/B VSS 0.43fF
C101 OR2X1_LOC_185/A OR2X1_LOC_192/B 0.31fF
C285 VDD OR2X1_LOC_185/A 1.01fF
C1284 OR2X1_LOC_462/B OR2X1_LOC_185/A 0.01fF
C1287 OR2X1_LOC_185/A OR2X1_LOC_483/a_8_216# 0.02fF
C2527 OR2X1_LOC_840/A OR2X1_LOC_185/A 0.11fF
C5004 OR2X1_LOC_185/A AND2X1_LOC_74/a_36_24# 0.01fF
C5761 OR2X1_LOC_185/A OR2X1_LOC_641/A 0.23fF
C6524 OR2X1_LOC_185/A AND2X1_LOC_238/a_8_24# 0.01fF
C6766 OR2X1_LOC_185/A OR2X1_LOC_643/A 0.18fF
C6772 OR2X1_LOC_185/A OR2X1_LOC_778/Y 0.05fF
C7008 AND2X1_LOC_91/B OR2X1_LOC_185/A 0.03fF
C7176 OR2X1_LOC_799/A OR2X1_LOC_185/A 0.07fF
C7536 OR2X1_LOC_185/A OR2X1_LOC_542/B 0.03fF
C7646 OR2X1_LOC_185/A AND2X1_LOC_56/B 1.45fF
C7993 OR2X1_LOC_185/A OR2X1_LOC_787/B 0.67fF
C8347 OR2X1_LOC_185/A AND2X1_LOC_235/a_36_24# 0.01fF
C9370 OR2X1_LOC_185/A OR2X1_LOC_506/A 0.02fF
C10202 OR2X1_LOC_185/A OR2X1_LOC_664/a_8_216# 0.02fF
C11398 OR2X1_LOC_185/A OR2X1_LOC_703/A 0.06fF
C11969 OR2X1_LOC_185/A OR2X1_LOC_243/B 0.15fF
C12083 OR2X1_LOC_185/A OR2X1_LOC_771/B 0.07fF
C12088 OR2X1_LOC_185/A OR2X1_LOC_209/A 0.15fF
C12103 OR2X1_LOC_185/A OR2X1_LOC_776/A 0.02fF
C12534 OR2X1_LOC_185/A OR2X1_LOC_593/B 0.04fF
C12823 OR2X1_LOC_185/A OR2X1_LOC_254/a_8_216# 0.01fF
C13672 OR2X1_LOC_185/A AND2X1_LOC_69/Y 0.01fF
C15283 OR2X1_LOC_185/A OR2X1_LOC_449/B 0.01fF
C16405 OR2X1_LOC_185/A OR2X1_LOC_786/A 0.02fF
C17821 OR2X1_LOC_185/A OR2X1_LOC_631/B 0.39fF
C18216 OR2X1_LOC_185/A AND2X1_LOC_253/a_8_24# 0.01fF
C18891 OR2X1_LOC_185/A OR2X1_LOC_71/A 0.02fF
C19139 OR2X1_LOC_185/A OR2X1_LOC_593/a_8_216# 0.01fF
C19602 OR2X1_LOC_185/A OR2X1_LOC_633/B 0.03fF
C20873 OR2X1_LOC_185/A OR2X1_LOC_592/a_8_216# 0.06fF
C21775 OR2X1_LOC_185/A AND2X1_LOC_117/a_8_24# 0.02fF
C23005 OR2X1_LOC_185/A OR2X1_LOC_539/Y 0.03fF
C23785 OR2X1_LOC_185/A OR2X1_LOC_254/A 0.01fF
C23903 OR2X1_LOC_185/A OR2X1_LOC_456/A 0.01fF
C24420 OR2X1_LOC_185/A AND2X1_LOC_406/a_8_24# 0.01fF
C25558 OR2X1_LOC_185/A AND2X1_LOC_518/a_8_24# 0.04fF
C26701 OR2X1_LOC_318/Y OR2X1_LOC_185/A 7.27fF
C28097 OR2X1_LOC_185/A OR2X1_LOC_76/A 0.03fF
C28131 OR2X1_LOC_185/A OR2X1_LOC_436/Y 0.03fF
C28445 OR2X1_LOC_185/A OR2X1_LOC_553/A 0.02fF
C28453 OR2X1_LOC_185/A OR2X1_LOC_266/a_8_216# 0.02fF
C29123 OR2X1_LOC_318/A OR2X1_LOC_185/A 0.02fF
C29148 OR2X1_LOC_151/A OR2X1_LOC_185/A 0.10fF
C30155 OR2X1_LOC_185/A AND2X1_LOC_252/a_8_24# 0.17fF
C31060 OR2X1_LOC_185/A OR2X1_LOC_520/B 0.10fF
C31800 OR2X1_LOC_185/A OR2X1_LOC_151/Y 0.03fF
C31816 OR2X1_LOC_185/A OR2X1_LOC_593/A 0.01fF
C32190 OR2X1_LOC_185/A OR2X1_LOC_664/Y 0.01fF
C33501 OR2X1_LOC_185/A OR2X1_LOC_243/A 0.02fF
C33691 OR2X1_LOC_185/A OR2X1_LOC_344/a_8_216# 0.01fF
C34041 OR2X1_LOC_185/A OR2X1_LOC_84/A 0.02fF
C34222 OR2X1_LOC_190/A OR2X1_LOC_185/A 0.03fF
C34379 OR2X1_LOC_185/A OR2X1_LOC_473/Y 0.16fF
C34454 OR2X1_LOC_185/A OR2X1_LOC_241/B 0.04fF
C34569 OR2X1_LOC_188/Y OR2X1_LOC_185/A 0.02fF
C36049 OR2X1_LOC_185/A OR2X1_LOC_810/A 0.03fF
C36317 OR2X1_LOC_715/B OR2X1_LOC_185/A 0.05fF
C36334 OR2X1_LOC_185/A OR2X1_LOC_543/A 0.48fF
C36581 OR2X1_LOC_185/A OR2X1_LOC_398/Y -0.06fF
C36813 OR2X1_LOC_656/B OR2X1_LOC_185/A 0.03fF
C37274 OR2X1_LOC_687/Y OR2X1_LOC_185/A 0.14fF
C38025 OR2X1_LOC_185/A OR2X1_LOC_78/A 0.47fF
C38965 OR2X1_LOC_185/A OR2X1_LOC_147/B 0.06fF
C38980 OR2X1_LOC_185/A AND2X1_LOC_517/a_8_24# 0.02fF
C39160 OR2X1_LOC_185/A OR2X1_LOC_318/B 3.55fF
C39345 OR2X1_LOC_538/A OR2X1_LOC_185/A 0.03fF
C39437 OR2X1_LOC_185/A OR2X1_LOC_802/A 0.10fF
C39475 OR2X1_LOC_185/A AND2X1_LOC_79/Y 0.01fF
C40087 OR2X1_LOC_318/a_8_216# OR2X1_LOC_185/A 0.01fF
C40173 OR2X1_LOC_185/A OR2X1_LOC_623/B 0.09fF
C40651 OR2X1_LOC_185/A OR2X1_LOC_833/B 0.03fF
C40672 OR2X1_LOC_185/A OR2X1_LOC_254/B 0.64fF
C41616 OR2X1_LOC_592/A OR2X1_LOC_185/A 0.03fF
C42019 OR2X1_LOC_84/B OR2X1_LOC_185/A 0.35fF
C42081 OR2X1_LOC_185/A AND2X1_LOC_518/a_36_24# 0.01fF
C42277 OR2X1_LOC_186/Y OR2X1_LOC_185/A 0.03fF
C42894 OR2X1_LOC_185/A OR2X1_LOC_574/A 0.04fF
C43273 OR2X1_LOC_319/a_8_216# OR2X1_LOC_185/A 0.05fF
C43792 OR2X1_LOC_185/A OR2X1_LOC_605/B 0.04fF
C44769 OR2X1_LOC_185/A OR2X1_LOC_348/B 0.01fF
C45009 OR2X1_LOC_185/A OR2X1_LOC_181/B 0.04fF
C45316 OR2X1_LOC_185/A AND2X1_LOC_603/a_8_24# 0.01fF
C46630 OR2X1_LOC_139/A OR2X1_LOC_185/A 0.03fF
C47941 OR2X1_LOC_185/A AND2X1_LOC_235/a_8_24# 0.01fF
C49225 OR2X1_LOC_97/A OR2X1_LOC_185/A 0.03fF
C49373 OR2X1_LOC_185/A OR2X1_LOC_475/B 0.04fF
C50224 OR2X1_LOC_185/A AND2X1_LOC_74/a_8_24# 0.14fF
C50424 OR2X1_LOC_185/A OR2X1_LOC_590/a_8_216# 0.01fF
C50710 OR2X1_LOC_185/A OR2X1_LOC_267/A 0.01fF
C51922 OR2X1_LOC_520/Y OR2X1_LOC_185/A 0.49fF
C52110 OR2X1_LOC_185/A OR2X1_LOC_590/Y 0.01fF
C52659 OR2X1_LOC_185/A OR2X1_LOC_776/Y 0.43fF
C53106 OR2X1_LOC_185/A OR2X1_LOC_370/a_8_216# 0.15fF
C54393 OR2X1_LOC_100/Y OR2X1_LOC_185/A 0.06fF
C54539 OR2X1_LOC_185/A OR2X1_LOC_532/B 0.17fF
C55161 OR2X1_LOC_185/A OR2X1_LOC_729/a_8_216# 0.05fF
C56111 OR2X1_LOC_185/A OR2X1_LOC_798/Y 0.03fF
C57647 OR2X1_LOC_185/A VSS 1.40fF
C100 OR2X1_LOC_151/A OR2X1_LOC_308/Y 0.07fF
C529 OR2X1_LOC_151/A OR2X1_LOC_535/a_36_216# 0.02fF
C699 OR2X1_LOC_151/A OR2X1_LOC_664/Y 0.03fF
C1942 OR2X1_LOC_324/B OR2X1_LOC_151/A 0.05fF
C1974 OR2X1_LOC_151/A AND2X1_LOC_142/a_8_24# 0.04fF
C1984 OR2X1_LOC_151/A AND2X1_LOC_314/a_8_24# 0.03fF
C2384 OR2X1_LOC_151/A AND2X1_LOC_311/a_8_24# 0.01fF
C2962 OR2X1_LOC_151/A OR2X1_LOC_473/Y 0.03fF
C4030 OR2X1_LOC_151/A OR2X1_LOC_356/A 0.02fF
C4540 OR2X1_LOC_151/A OR2X1_LOC_810/A 0.10fF
C4840 OR2X1_LOC_715/B OR2X1_LOC_151/A 0.10fF
C6551 OR2X1_LOC_151/A OR2X1_LOC_78/A 0.31fF
C6594 AND2X1_LOC_331/a_36_24# OR2X1_LOC_151/A 0.01fF
C7461 OR2X1_LOC_501/B OR2X1_LOC_151/A 0.07fF
C7466 AND2X1_LOC_320/a_36_24# OR2X1_LOC_151/A 0.01fF
C7488 OR2X1_LOC_151/A OR2X1_LOC_147/B 0.14fF
C7507 OR2X1_LOC_151/A OR2X1_LOC_317/A 0.09fF
C7724 OR2X1_LOC_151/A OR2X1_LOC_854/A 0.01fF
C7834 OR2X1_LOC_121/Y OR2X1_LOC_151/A 0.07fF
C7894 OR2X1_LOC_151/A OR2X1_LOC_538/A 0.08fF
C8790 OR2X1_LOC_151/A OR2X1_LOC_623/B 0.20fF
C9160 OR2X1_LOC_151/A OR2X1_LOC_140/A 0.01fF
C9656 OR2X1_LOC_151/A AND2X1_LOC_321/a_8_24# 0.04fF
C9978 OR2X1_LOC_151/A AND2X1_LOC_248/a_8_24# 0.01fF
C10817 OR2X1_LOC_186/Y OR2X1_LOC_151/A 0.13fF
C11386 OR2X1_LOC_151/A OR2X1_LOC_574/A 0.09fF
C11764 OR2X1_LOC_319/a_8_216# OR2X1_LOC_151/A 0.03fF
C13030 OR2X1_LOC_151/A OR2X1_LOC_499/B 0.01fF
C13172 OR2X1_LOC_151/A OR2X1_LOC_486/B 0.02fF
C14114 OR2X1_LOC_151/A OR2X1_LOC_330/a_8_216# 0.02fF
C15144 OR2X1_LOC_151/A OR2X1_LOC_324/A 0.07fF
C16412 OR2X1_LOC_703/B OR2X1_LOC_151/A 0.08fF
C17121 OR2X1_LOC_151/A OR2X1_LOC_532/a_8_216# 0.06fF
C17566 OR2X1_LOC_97/A OR2X1_LOC_151/A 0.03fF
C17657 OR2X1_LOC_151/A OR2X1_LOC_475/B 0.03fF
C18115 OR2X1_LOC_151/A OR2X1_LOC_629/Y 0.14fF
C18560 OR2X1_LOC_151/A AND2X1_LOC_314/a_36_24# 0.01fF
C19078 OR2X1_LOC_151/A OR2X1_LOC_778/A 0.01fF
C19770 OR2X1_LOC_151/A OR2X1_LOC_361/a_8_216# 0.02fF
C20172 OR2X1_LOC_151/A OR2X1_LOC_267/Y 0.04fF
C20699 OR2X1_LOC_151/A AND2X1_LOC_321/a_36_24# 0.01fF
C21028 OR2X1_LOC_151/A OR2X1_LOC_342/A 0.01fF
C21487 OR2X1_LOC_151/A OR2X1_LOC_355/A 0.09fF
C23016 OR2X1_LOC_151/A OR2X1_LOC_532/B 0.79fF
C23217 OR2X1_LOC_151/A OR2X1_LOC_440/B 0.01fF
C24347 OR2X1_LOC_151/A OR2X1_LOC_151/a_8_216# 0.01fF
C24882 VDD OR2X1_LOC_151/A 0.43fF
C26914 OR2X1_LOC_151/A OR2X1_LOC_115/B 0.20fF
C27007 OR2X1_LOC_151/A OR2X1_LOC_840/A 0.10fF
C27422 OR2X1_LOC_151/A OR2X1_LOC_216/A 0.07fF
C28158 OR2X1_LOC_151/A OR2X1_LOC_532/Y 0.03fF
C28322 OR2X1_LOC_151/A OR2X1_LOC_447/A 0.07fF
C28428 OR2X1_LOC_151/A AND2X1_LOC_127/a_8_24# 0.01fF
C29218 OR2X1_LOC_151/A OR2X1_LOC_435/Y 0.05fF
C29935 OR2X1_LOC_151/A AND2X1_LOC_437/a_8_24# 0.01fF
C30325 OR2X1_LOC_151/A OR2X1_LOC_294/Y 0.02fF
C30441 OR2X1_LOC_114/Y OR2X1_LOC_151/A 0.34fF
C31313 OR2X1_LOC_151/A OR2X1_LOC_778/Y 0.14fF
C31560 AND2X1_LOC_91/B OR2X1_LOC_151/A 0.29fF
C32050 OR2X1_LOC_151/A OR2X1_LOC_631/a_8_216# 0.02fF
C32092 OR2X1_LOC_151/A AND2X1_LOC_56/B 1.23fF
C33688 OR2X1_LOC_151/A OR2X1_LOC_186/a_8_216# 0.02fF
C33802 OR2X1_LOC_151/A OR2X1_LOC_506/A 0.07fF
C33963 OR2X1_LOC_151/A AND2X1_LOC_420/a_8_24# 0.03fF
C34062 OR2X1_LOC_151/A OR2X1_LOC_180/B 0.43fF
C34442 OR2X1_LOC_151/A OR2X1_LOC_788/B 0.12fF
C34614 OR2X1_LOC_151/A OR2X1_LOC_630/a_8_216# 0.02fF
C35040 OR2X1_LOC_151/A AND2X1_LOC_173/a_8_24# 0.04fF
C35801 OR2X1_LOC_151/A AND2X1_LOC_295/a_8_24# 0.01fF
C35928 OR2X1_LOC_116/a_8_216# OR2X1_LOC_151/A 0.05fF
C36323 OR2X1_LOC_116/A OR2X1_LOC_151/A 0.02fF
C36569 OR2X1_LOC_151/A OR2X1_LOC_209/A 0.04fF
C37405 OR2X1_LOC_151/A OR2X1_LOC_317/B 0.04fF
C38137 OR2X1_LOC_151/A OR2X1_LOC_506/B 0.03fF
C38194 OR2X1_LOC_151/A OR2X1_LOC_247/Y 0.02fF
C38632 OR2X1_LOC_151/A AND2X1_LOC_485/a_8_24# 0.12fF
C39334 OR2X1_LOC_151/A AND2X1_LOC_292/a_8_24# 0.01fF
C39721 OR2X1_LOC_128/A OR2X1_LOC_151/A 0.04fF
C39755 OR2X1_LOC_151/A OR2X1_LOC_449/B 0.07fF
C40063 OR2X1_LOC_317/a_8_216# OR2X1_LOC_151/A 0.04fF
C41315 OR2X1_LOC_151/A OR2X1_LOC_346/A 0.01fF
C41865 OR2X1_LOC_151/A AND2X1_LOC_297/a_8_24# 0.01fF
C42335 OR2X1_LOC_151/A OR2X1_LOC_631/B 0.05fF
C43170 OR2X1_LOC_151/A OR2X1_LOC_632/A 0.03fF
C43496 OR2X1_LOC_151/A OR2X1_LOC_355/a_8_216# 0.02fF
C44786 OR2X1_LOC_506/Y OR2X1_LOC_151/A 0.01fF
C44843 OR2X1_LOC_151/A OR2X1_LOC_630/Y 0.38fF
C44935 OR2X1_LOC_151/A OR2X1_LOC_346/B 0.01fF
C45292 OR2X1_LOC_151/A AND2X1_LOC_167/a_8_24# 0.03fF
C45338 OR2X1_LOC_128/B OR2X1_LOC_151/A 0.01fF
C45608 OR2X1_LOC_151/A OR2X1_LOC_535/a_8_216# 0.03fF
C46190 OR2X1_LOC_330/Y OR2X1_LOC_151/A 0.04fF
C47592 OR2X1_LOC_151/A OR2X1_LOC_347/B 0.01fF
C47597 OR2X1_LOC_151/A OR2X1_LOC_539/Y 0.03fF
C47664 OR2X1_LOC_151/A AND2X1_LOC_176/a_8_24# 0.01fF
C47866 OR2X1_LOC_151/A OR2X1_LOC_319/Y 0.10fF
C49210 OR2X1_LOC_151/A OR2X1_LOC_630/B 0.02fF
C49911 OR2X1_LOC_151/A OR2X1_LOC_705/B 0.03fF
C50499 OR2X1_LOC_151/A OR2X1_LOC_201/A 0.13fF
C51346 OR2X1_LOC_319/B OR2X1_LOC_151/A 0.11fF
C51360 OR2X1_LOC_318/Y OR2X1_LOC_151/A 0.02fF
C51434 OR2X1_LOC_151/A OR2X1_LOC_296/Y 0.08fF
C51459 OR2X1_LOC_151/A OR2X1_LOC_436/a_8_216# 0.04fF
C51779 AND2X1_LOC_331/a_8_24# OR2X1_LOC_151/A 0.03fF
C52590 AND2X1_LOC_320/a_8_24# OR2X1_LOC_151/A 0.03fF
C52795 OR2X1_LOC_151/A OR2X1_LOC_436/Y 0.03fF
C55072 OR2X1_LOC_151/A OR2X1_LOC_631/A 0.02fF
C55383 OR2X1_LOC_151/A AND2X1_LOC_485/a_36_24# 0.01fF
C55463 OR2X1_LOC_151/A OR2X1_LOC_168/Y 0.47fF
C57768 OR2X1_LOC_151/A VSS -4.85fF
C2735 OR2X1_LOC_619/Y OR2X1_LOC_72/Y 0.07fF
C3694 AND2X1_LOC_706/Y OR2X1_LOC_619/Y 0.01fF
C3887 OR2X1_LOC_158/B OR2X1_LOC_619/Y 0.01fF
C4624 AND2X1_LOC_302/a_8_24# OR2X1_LOC_619/Y 0.02fF
C5541 AND2X1_LOC_537/Y OR2X1_LOC_619/Y 0.07fF
C8838 VDD OR2X1_LOC_619/Y 1.53fF
C9076 OR2X1_LOC_619/Y OR2X1_LOC_67/Y 0.07fF
C9101 OR2X1_LOC_619/Y OR2X1_LOC_163/Y 0.01fF
C10709 OR2X1_LOC_416/Y OR2X1_LOC_619/Y 0.03fF
C11745 OR2X1_LOC_45/B OR2X1_LOC_619/Y 0.13fF
C14454 OR2X1_LOC_316/Y OR2X1_LOC_619/Y 0.03fF
C14505 AND2X1_LOC_390/B OR2X1_LOC_619/Y 0.07fF
C15082 OR2X1_LOC_619/Y OR2X1_LOC_320/a_8_216# 0.01fF
C15683 AND2X1_LOC_303/B OR2X1_LOC_619/Y -0.03fF
C16562 OR2X1_LOC_305/Y OR2X1_LOC_619/Y 0.01fF
C16617 OR2X1_LOC_417/Y OR2X1_LOC_619/Y 13.69fF
C16790 OR2X1_LOC_619/Y OR2X1_LOC_171/Y 1.75fF
C18641 OR2X1_LOC_298/a_8_216# OR2X1_LOC_619/Y 0.02fF
C19472 OR2X1_LOC_235/B OR2X1_LOC_619/Y 0.07fF
C19723 OR2X1_LOC_619/Y OR2X1_LOC_331/Y 0.07fF
C20632 OR2X1_LOC_619/Y OR2X1_LOC_320/a_36_216# 0.01fF
C21613 AND2X1_LOC_335/Y OR2X1_LOC_619/Y 0.02fF
C23866 OR2X1_LOC_312/Y OR2X1_LOC_619/Y 0.07fF
C24034 OR2X1_LOC_619/Y OR2X1_LOC_13/B 0.15fF
C24946 AND2X1_LOC_592/Y OR2X1_LOC_619/Y 0.03fF
C25143 AND2X1_LOC_712/B OR2X1_LOC_619/Y 0.01fF
C25520 OR2X1_LOC_89/A OR2X1_LOC_619/Y 0.03fF
C26383 AND2X1_LOC_727/A OR2X1_LOC_619/Y 0.06fF
C27179 OR2X1_LOC_619/Y AND2X1_LOC_621/Y 0.33fF
C27353 OR2X1_LOC_619/Y OR2X1_LOC_71/A 0.07fF
C27659 AND2X1_LOC_333/a_8_24# OR2X1_LOC_619/Y 0.06fF
C29126 OR2X1_LOC_619/Y OR2X1_LOC_16/A 0.13fF
C29650 OR2X1_LOC_298/a_36_216# OR2X1_LOC_619/Y 0.01fF
C30027 OR2X1_LOC_619/Y AND2X1_LOC_447/Y 0.07fF
C30120 OR2X1_LOC_619/Y AND2X1_LOC_448/Y 0.02fF
C30990 OR2X1_LOC_599/A OR2X1_LOC_619/Y 0.03fF
C31299 AND2X1_LOC_535/a_8_24# OR2X1_LOC_619/Y 0.03fF
C31432 OR2X1_LOC_320/Y OR2X1_LOC_619/Y 0.03fF
C32164 AND2X1_LOC_841/B OR2X1_LOC_619/Y 0.07fF
C32636 OR2X1_LOC_619/Y AND2X1_LOC_622/a_8_24# 0.10fF
C34419 OR2X1_LOC_607/a_8_216# OR2X1_LOC_619/Y 0.04fF
C36262 OR2X1_LOC_619/Y OR2X1_LOC_321/a_8_216# 0.02fF
C36887 OR2X1_LOC_321/Y OR2X1_LOC_619/Y 0.03fF
C37742 AND2X1_LOC_154/Y OR2X1_LOC_619/Y 0.03fF
C39020 AND2X1_LOC_777/a_8_24# OR2X1_LOC_619/Y 0.02fF
C39750 AND2X1_LOC_160/Y OR2X1_LOC_619/Y 0.02fF
C40451 OR2X1_LOC_619/Y AND2X1_LOC_608/a_8_24# 0.06fF
C40696 OR2X1_LOC_619/Y OR2X1_LOC_601/Y 0.03fF
C41091 OR2X1_LOC_118/Y OR2X1_LOC_619/Y 0.03fF
C41831 OR2X1_LOC_619/Y OR2X1_LOC_321/a_36_216# 0.01fF
C42065 OR2X1_LOC_619/Y OR2X1_LOC_65/a_8_216# 0.04fF
C42321 OR2X1_LOC_604/A OR2X1_LOC_619/Y 0.05fF
C42718 OR2X1_LOC_176/Y OR2X1_LOC_619/Y 0.02fF
C42727 OR2X1_LOC_533/Y OR2X1_LOC_619/Y 0.06fF
C42867 OR2X1_LOC_619/Y OR2X1_LOC_265/Y 0.07fF
C43023 OR2X1_LOC_619/Y OR2X1_LOC_163/A 0.01fF
C43348 AND2X1_LOC_155/Y OR2X1_LOC_619/Y 0.16fF
C43556 AND2X1_LOC_539/Y OR2X1_LOC_619/Y 0.05fF
C44153 OR2X1_LOC_298/Y OR2X1_LOC_619/Y 0.04fF
C46643 OR2X1_LOC_135/Y OR2X1_LOC_619/Y 0.10fF
C47825 AND2X1_LOC_318/Y OR2X1_LOC_619/Y 0.02fF
C48943 OR2X1_LOC_158/a_8_216# OR2X1_LOC_619/Y 0.01fF
C49731 AND2X1_LOC_715/A OR2X1_LOC_619/Y 0.07fF
C50245 AND2X1_LOC_729/Y OR2X1_LOC_619/Y 0.07fF
C50273 AND2X1_LOC_784/A OR2X1_LOC_619/Y 0.02fF
C50438 OR2X1_LOC_619/Y OR2X1_LOC_172/Y 0.05fF
C50718 OR2X1_LOC_619/Y OR2X1_LOC_52/B 2.26fF
C51004 AND2X1_LOC_161/Y OR2X1_LOC_619/Y 0.01fF
C51906 AND2X1_LOC_593/Y OR2X1_LOC_619/Y 0.03fF
C53111 OR2X1_LOC_619/Y AND2X1_LOC_436/Y 0.03fF
C54487 AND2X1_LOC_156/a_8_24# OR2X1_LOC_619/Y 0.01fF
C54692 AND2X1_LOC_799/a_8_24# OR2X1_LOC_619/Y 0.03fF
C54702 OR2X1_LOC_619/Y OR2X1_LOC_158/Y 0.01fF
C56915 OR2X1_LOC_619/Y VSS -3.41fF
C1603 OR2X1_LOC_584/a_8_216# OR2X1_LOC_52/B 0.03fF
C2018 OR2X1_LOC_16/A OR2X1_LOC_52/B 0.21fF
C2260 AND2X1_LOC_687/Y OR2X1_LOC_52/B -0.11fF
C2955 AND2X1_LOC_447/Y OR2X1_LOC_52/B 0.01fF
C3037 AND2X1_LOC_448/Y OR2X1_LOC_52/B 0.05fF
C3098 AND2X1_LOC_729/B OR2X1_LOC_52/B 0.15fF
C3530 AND2X1_LOC_708/a_36_24# OR2X1_LOC_52/B 0.01fF
C3886 OR2X1_LOC_599/A OR2X1_LOC_52/B 0.07fF
C4120 OR2X1_LOC_177/a_8_216# OR2X1_LOC_52/B 0.02fF
C4697 OR2X1_LOC_32/a_8_216# OR2X1_LOC_52/B 0.01fF
C4856 OR2X1_LOC_52/B OR2X1_LOC_424/Y -0.01fF
C4911 AND2X1_LOC_707/Y OR2X1_LOC_52/B 0.03fF
C6169 OR2X1_LOC_52/B AND2X1_LOC_780/a_36_24# 0.01fF
C6752 OR2X1_LOC_74/Y OR2X1_LOC_52/B 0.03fF
C7029 OR2X1_LOC_52/B OR2X1_LOC_525/a_8_216# 0.06fF
C7532 OR2X1_LOC_766/a_8_216# OR2X1_LOC_52/B 0.03fF
C8665 OR2X1_LOC_7/Y OR2X1_LOC_52/B 0.01fF
C8943 OR2X1_LOC_516/B OR2X1_LOC_52/B 0.03fF
C9693 AND2X1_LOC_828/a_8_24# OR2X1_LOC_52/B 0.02fF
C9701 OR2X1_LOC_177/a_36_216# OR2X1_LOC_52/B 0.03fF
C10175 AND2X1_LOC_707/a_36_24# OR2X1_LOC_52/B 0.01fF
C10718 AND2X1_LOC_154/Y OR2X1_LOC_52/B 0.58fF
C11077 AND2X1_LOC_624/A OR2X1_LOC_52/B 0.06fF
C11871 OR2X1_LOC_524/Y OR2X1_LOC_52/B 0.11fF
C12070 OR2X1_LOC_52/B OR2X1_LOC_746/Y 0.01fF
C12707 AND2X1_LOC_160/Y OR2X1_LOC_52/B 0.13fF
C13309 OR2X1_LOC_273/Y OR2X1_LOC_52/B 0.02fF
C13498 OR2X1_LOC_744/a_8_216# OR2X1_LOC_52/B 0.03fF
C13856 OR2X1_LOC_52/B OR2X1_LOC_142/Y 0.03fF
C14561 OR2X1_LOC_52/Y OR2X1_LOC_52/B 0.01fF
C14985 OR2X1_LOC_65/a_8_216# OR2X1_LOC_52/B 0.06fF
C15202 OR2X1_LOC_604/A OR2X1_LOC_52/B 0.14fF
C15203 OR2X1_LOC_745/a_8_216# OR2X1_LOC_52/B 0.02fF
C15717 OR2X1_LOC_52/B OR2X1_LOC_265/Y 0.07fF
C16209 AND2X1_LOC_155/Y OR2X1_LOC_52/B 0.02fF
C16219 OR2X1_LOC_230/a_8_216# OR2X1_LOC_52/B 0.04fF
C16241 AND2X1_LOC_633/Y OR2X1_LOC_52/B 0.02fF
C16828 OR2X1_LOC_316/a_8_216# OR2X1_LOC_52/B 0.02fF
C16993 OR2X1_LOC_52/B OR2X1_LOC_746/a_8_216# 0.02fF
C17020 OR2X1_LOC_298/Y OR2X1_LOC_52/B 0.02fF
C17074 OR2X1_LOC_52/B OR2X1_LOC_27/a_8_216# 0.03fF
C17362 AND2X1_LOC_434/Y OR2X1_LOC_52/B 0.07fF
C17560 OR2X1_LOC_595/Y OR2X1_LOC_52/B 0.02fF
C17809 OR2X1_LOC_837/B OR2X1_LOC_52/B 0.03fF
C17870 OR2X1_LOC_69/a_8_216# OR2X1_LOC_52/B 0.01fF
C18600 OR2X1_LOC_766/Y OR2X1_LOC_52/B 0.03fF
C19106 OR2X1_LOC_517/a_8_216# OR2X1_LOC_52/B 0.03fF
C19447 OR2X1_LOC_135/Y OR2X1_LOC_52/B 0.07fF
C19581 AND2X1_LOC_520/Y OR2X1_LOC_52/B 0.01fF
C19986 AND2X1_LOC_160/a_8_24# OR2X1_LOC_52/B 0.04fF
C20815 OR2X1_LOC_697/a_8_216# OR2X1_LOC_52/B 0.04fF
C21374 OR2X1_LOC_385/Y OR2X1_LOC_52/B 0.72fF
C22041 OR2X1_LOC_229/a_8_216# OR2X1_LOC_52/B -0.03fF
C22688 OR2X1_LOC_52/B OR2X1_LOC_27/a_36_216# 0.02fF
C23046 AND2X1_LOC_729/Y OR2X1_LOC_52/B 0.03fF
C23064 AND2X1_LOC_784/A OR2X1_LOC_52/B 0.75fF
C23752 OR2X1_LOC_584/Y OR2X1_LOC_52/B 0.23fF
C24198 OR2X1_LOC_485/Y OR2X1_LOC_52/B 0.03fF
C24537 OR2X1_LOC_744/Y OR2X1_LOC_52/B 0.01fF
C25048 OR2X1_LOC_58/a_8_216# OR2X1_LOC_52/B 0.01fF
C25117 OR2X1_LOC_680/A OR2X1_LOC_52/B 0.10fF
C25551 OR2X1_LOC_423/a_8_216# OR2X1_LOC_52/B 0.03fF
C26356 OR2X1_LOC_81/a_8_216# OR2X1_LOC_52/B 0.03fF
C27231 OR2X1_LOC_511/Y OR2X1_LOC_52/B 3.83fF
C27861 OR2X1_LOC_316/a_36_216# OR2X1_LOC_52/B 0.02fF
C28632 OR2X1_LOC_52/B OR2X1_LOC_423/Y 0.03fF
C28907 OR2X1_LOC_69/a_36_216# OR2X1_LOC_52/B -0.00fF
C28933 OR2X1_LOC_74/A OR2X1_LOC_52/B 1.42fF
C29626 OR2X1_LOC_52/B AND2X1_LOC_448/a_8_24# 0.03fF
C30139 AND2X1_LOC_779/a_8_24# OR2X1_LOC_52/B 0.03fF
C31496 OR2X1_LOC_65/Y OR2X1_LOC_52/B 0.28fF
C31589 OR2X1_LOC_52/B OR2X1_LOC_72/Y 0.05fF
C31780 OR2X1_LOC_697/Y OR2X1_LOC_52/B 0.12fF
C31891 OR2X1_LOC_696/Y OR2X1_LOC_52/B 0.01fF
C32221 OR2X1_LOC_595/a_8_216# OR2X1_LOC_52/B 0.02fF
C32587 OR2X1_LOC_58/Y OR2X1_LOC_52/B 0.04fF
C32713 OR2X1_LOC_81/Y OR2X1_LOC_52/B 0.04fF
C33523 OR2X1_LOC_695/a_8_216# OR2X1_LOC_52/B 0.03fF
C33560 AND2X1_LOC_302/a_8_24# OR2X1_LOC_52/B 0.04fF
C33593 OR2X1_LOC_32/Y OR2X1_LOC_52/B 0.01fF
C34373 OR2X1_LOC_69/Y OR2X1_LOC_52/B 0.01fF
C34433 AND2X1_LOC_537/Y OR2X1_LOC_52/B 4.21fF
C35120 OR2X1_LOC_526/Y OR2X1_LOC_52/B 0.03fF
C35507 AND2X1_LOC_714/B OR2X1_LOC_52/B 0.07fF
C36266 OR2X1_LOC_516/Y OR2X1_LOC_52/B 0.03fF
C36426 AND2X1_LOC_160/a_36_24# OR2X1_LOC_52/B 0.01fF
C37635 VDD OR2X1_LOC_52/B 0.92fF
C39543 OR2X1_LOC_416/Y OR2X1_LOC_52/B 0.03fF
C40231 OR2X1_LOC_485/a_8_216# OR2X1_LOC_52/B 0.05fF
C40559 OR2X1_LOC_45/B OR2X1_LOC_52/B 0.29fF
C43333 OR2X1_LOC_316/Y OR2X1_LOC_52/B 0.03fF
C43386 AND2X1_LOC_390/B OR2X1_LOC_52/B 0.07fF
C43796 AND2X1_LOC_840/B OR2X1_LOC_52/B 0.07fF
C43805 OR2X1_LOC_74/a_8_216# OR2X1_LOC_52/B 0.03fF
C44653 AND2X1_LOC_303/B OR2X1_LOC_52/B -0.02fF
C45548 OR2X1_LOC_189/Y OR2X1_LOC_52/B 0.15fF
C45580 OR2X1_LOC_417/Y OR2X1_LOC_52/B 0.07fF
C45592 OR2X1_LOC_311/Y OR2X1_LOC_52/B 0.03fF
C45748 OR2X1_LOC_52/B AND2X1_LOC_780/a_8_24# 0.04fF
C45750 OR2X1_LOC_52/B OR2X1_LOC_171/Y 0.02fF
C46004 AND2X1_LOC_276/Y OR2X1_LOC_52/B 0.05fF
C46293 OR2X1_LOC_52/B AND2X1_LOC_448/a_36_24# 0.01fF
C46350 OR2X1_LOC_441/Y OR2X1_LOC_52/B 0.11fF
C46410 AND2X1_LOC_139/B OR2X1_LOC_52/B 0.07fF
C47334 OR2X1_LOC_517/Y OR2X1_LOC_52/B 0.03fF
C47424 OR2X1_LOC_409/B OR2X1_LOC_52/B 0.06fF
C47698 OR2X1_LOC_298/a_8_216# OR2X1_LOC_52/B 0.03fF
C47803 OR2X1_LOC_229/Y OR2X1_LOC_52/B 0.01fF
C48602 AND2X1_LOC_319/A OR2X1_LOC_52/B 0.07fF
C48649 OR2X1_LOC_52/a_8_216# OR2X1_LOC_52/B 0.07fF
C48670 AND2X1_LOC_708/a_8_24# OR2X1_LOC_52/B 0.03fF
C49485 OR2X1_LOC_83/Y OR2X1_LOC_52/B 0.04fF
C49792 OR2X1_LOC_695/Y OR2X1_LOC_52/B 0.01fF
C51143 AND2X1_LOC_454/A OR2X1_LOC_52/B 0.02fF
C51210 AND2X1_LOC_539/a_8_24# OR2X1_LOC_52/B 0.02fF
C51363 OR2X1_LOC_52/B AND2X1_LOC_783/B 0.03fF
C51696 OR2X1_LOC_52/B OR2X1_LOC_745/Y 0.01fF
C52884 AND2X1_LOC_307/a_8_24# OR2X1_LOC_52/B 0.03fF
C53002 OR2X1_LOC_52/B OR2X1_LOC_13/B 0.23fF
C53432 OR2X1_LOC_52/B OR2X1_LOC_142/a_8_216# 0.06fF
C53534 OR2X1_LOC_52/B OR2X1_LOC_595/A 0.14fF
C53684 AND2X1_LOC_154/a_8_24# OR2X1_LOC_52/B 0.02fF
C54130 AND2X1_LOC_712/B OR2X1_LOC_52/B 0.02fF
C54364 OR2X1_LOC_765/Y OR2X1_LOC_52/B 0.02fF
C54517 OR2X1_LOC_89/A OR2X1_LOC_52/B 0.14fF
C55170 AND2X1_LOC_473/Y OR2X1_LOC_52/B 0.01fF
C55259 AND2X1_LOC_707/a_8_24# OR2X1_LOC_52/B 0.02fF
C55412 AND2X1_LOC_727/A OR2X1_LOC_52/B 0.03fF
C56182 OR2X1_LOC_438/Y OR2X1_LOC_52/B 0.02fF
C56217 AND2X1_LOC_621/Y OR2X1_LOC_52/B 0.05fF
C56531 OR2X1_LOC_52/B VSS 1.59fF
C749 OR2X1_LOC_45/B OR2X1_LOC_416/Y 0.06fF
C1540 OR2X1_LOC_45/B OR2X1_LOC_45/a_8_216# 0.08fF
C1561 OR2X1_LOC_45/B AND2X1_LOC_831/a_8_24# 0.01fF
C4118 OR2X1_LOC_45/B OR2X1_LOC_438/a_8_216# 0.06fF
C4359 OR2X1_LOC_45/B AND2X1_LOC_227/a_8_24# 0.17fF
C4473 OR2X1_LOC_45/B OR2X1_LOC_316/Y 0.06fF
C4531 OR2X1_LOC_45/B AND2X1_LOC_390/B 0.07fF
C4557 OR2X1_LOC_45/B OR2X1_LOC_431/Y 0.02fF
C4902 OR2X1_LOC_45/B AND2X1_LOC_840/B 0.03fF
C5193 OR2X1_LOC_45/B OR2X1_LOC_79/a_8_216# 0.02fF
C5223 OR2X1_LOC_45/B AND2X1_LOC_301/a_8_24# 0.02fF
C5381 OR2X1_LOC_45/B AND2X1_LOC_308/a_8_24# 0.02fF
C5709 OR2X1_LOC_45/B OR2X1_LOC_695/a_36_216# 0.02fF
C6601 OR2X1_LOC_45/B OR2X1_LOC_91/Y 0.03fF
C6608 OR2X1_LOC_45/B OR2X1_LOC_305/Y 0.02fF
C6671 OR2X1_LOC_45/B OR2X1_LOC_527/Y 0.11fF
C6679 OR2X1_LOC_45/B OR2X1_LOC_417/Y 0.07fF
C6689 OR2X1_LOC_45/B OR2X1_LOC_311/Y 0.03fF
C6911 OR2X1_LOC_45/B OR2X1_LOC_171/Y 2.76fF
C7173 OR2X1_LOC_45/B AND2X1_LOC_831/Y 0.01fF
C7495 OR2X1_LOC_45/B AND2X1_LOC_139/B 0.03fF
C7816 OR2X1_LOC_45/B OR2X1_LOC_135/a_8_216# 0.01fF
C8819 OR2X1_LOC_45/B OR2X1_LOC_497/Y 0.02fF
C9121 OR2X1_LOC_45/B AND2X1_LOC_249/a_8_24# 0.11fF
C9662 OR2X1_LOC_45/B AND2X1_LOC_319/A 0.07fF
C9740 OR2X1_LOC_45/B AND2X1_LOC_708/a_8_24# 0.01fF
C10067 OR2X1_LOC_45/B AND2X1_LOC_318/a_8_24# 0.01fF
C10085 OR2X1_LOC_45/B AND2X1_LOC_361/A 0.30fF
C10333 OR2X1_LOC_45/B OR2X1_LOC_395/a_8_216# 0.01fF
C10803 OR2X1_LOC_45/B OR2X1_LOC_79/a_36_216# 0.02fF
C10825 OR2X1_LOC_45/B OR2X1_LOC_695/Y 0.02fF
C10901 OR2X1_LOC_45/B OR2X1_LOC_406/a_8_216# 0.01fF
C11650 OR2X1_LOC_45/B OR2X1_LOC_692/Y 0.01fF
C12202 OR2X1_LOC_45/B AND2X1_LOC_454/A 0.02fF
C12266 OR2X1_LOC_45/B AND2X1_LOC_334/a_8_24# 0.03fF
C12943 OR2X1_LOC_45/B OR2X1_LOC_505/a_8_216# 0.05fF
C13972 OR2X1_LOC_45/B AND2X1_LOC_307/a_8_24# 0.01fF
C14042 OR2X1_LOC_45/B OR2X1_LOC_75/a_8_216# 0.03fF
C14152 OR2X1_LOC_45/B OR2X1_LOC_13/B 0.17fF
C14643 OR2X1_LOC_45/B OR2X1_LOC_595/A 0.03fF
C15069 OR2X1_LOC_45/B OR2X1_LOC_528/Y 0.25fF
C15209 OR2X1_LOC_45/B AND2X1_LOC_712/B 0.15fF
C15590 OR2X1_LOC_45/B OR2X1_LOC_89/A 0.05fF
C16289 OR2X1_LOC_45/B AND2X1_LOC_473/Y 0.02fF
C16315 OR2X1_LOC_45/B AND2X1_LOC_707/a_8_24# 0.03fF
C16354 OR2X1_LOC_45/B OR2X1_LOC_45/Y 0.47fF
C17258 OR2X1_LOC_45/B AND2X1_LOC_621/Y 0.03fF
C17769 OR2X1_LOC_45/B OR2X1_LOC_504/Y 0.32fF
C19303 OR2X1_LOC_45/B OR2X1_LOC_16/A 0.24fF
C19325 OR2X1_LOC_45/B OR2X1_LOC_108/Y 0.02fF
C19514 OR2X1_LOC_45/B AND2X1_LOC_687/Y 0.01fF
C20205 OR2X1_LOC_45/B AND2X1_LOC_447/Y 0.01fF
C20207 OR2X1_LOC_45/B AND2X1_LOC_334/Y 0.01fF
C20262 OR2X1_LOC_45/B AND2X1_LOC_448/Y 0.01fF
C20323 OR2X1_LOC_45/B AND2X1_LOC_729/B 0.03fF
C20828 OR2X1_LOC_45/B AND2X1_LOC_227/Y 0.11fF
C21140 OR2X1_LOC_45/B OR2X1_LOC_599/A 0.03fF
C21158 OR2X1_LOC_45/B AND2X1_LOC_267/a_36_24# 0.01fF
C21927 OR2X1_LOC_45/B OR2X1_LOC_531/Y 0.02fF
C22247 OR2X1_LOC_45/B OR2X1_LOC_424/Y 0.01fF
C22307 OR2X1_LOC_45/B AND2X1_LOC_707/Y 0.79fF
C23203 OR2X1_LOC_45/B AND2X1_LOC_776/a_8_24# 0.01fF
C25056 OR2X1_LOC_45/B OR2X1_LOC_75/a_36_216# 0.01fF
C26870 OR2X1_LOC_45/B OR2X1_LOC_395/Y 0.14fF
C28217 OR2X1_LOC_45/B AND2X1_LOC_778/Y 0.01fF
C28297 OR2X1_LOC_45/B AND2X1_LOC_624/A 0.10fF
C28633 OR2X1_LOC_45/B AND2X1_LOC_434/a_8_24# 0.02fF
C29061 OR2X1_LOC_45/B OR2X1_LOC_524/Y 0.01fF
C29909 OR2X1_LOC_45/B AND2X1_LOC_160/Y 0.01fF
C30456 OR2X1_LOC_45/B OR2X1_LOC_273/Y 0.01fF
C30519 OR2X1_LOC_45/B OR2X1_LOC_75/Y 0.50fF
C31098 OR2X1_LOC_45/B OR2X1_LOC_142/Y 0.03fF
C31243 OR2X1_LOC_45/B OR2X1_LOC_118/Y 0.02fF
C31279 OR2X1_LOC_45/B OR2X1_LOC_262/Y 0.27fF
C31289 OR2X1_LOC_45/B OR2X1_LOC_238/Y 0.03fF
C32370 OR2X1_LOC_45/B OR2X1_LOC_315/a_8_216# 0.01fF
C32385 OR2X1_LOC_45/B OR2X1_LOC_604/A 0.06fF
C32472 OR2X1_LOC_45/B OR2X1_LOC_306/Y 0.06fF
C32864 OR2X1_LOC_45/B AND2X1_LOC_549/a_8_24# 0.03fF
C32870 OR2X1_LOC_45/B AND2X1_LOC_506/a_8_24# 0.03fF
C32926 OR2X1_LOC_45/B OR2X1_LOC_265/Y 0.11fF
C33195 OR2X1_LOC_45/B OR2X1_LOC_183/a_8_216# 0.09fF
C33454 OR2X1_LOC_45/B AND2X1_LOC_633/Y 0.03fF
C33679 OR2X1_LOC_45/B AND2X1_LOC_539/Y 0.03fF
C34526 OR2X1_LOC_45/B AND2X1_LOC_434/Y 0.07fF
C34627 OR2X1_LOC_45/B OR2X1_LOC_496/Y 0.61fF
C34809 OR2X1_LOC_45/B OR2X1_LOC_595/Y 0.02fF
C36166 OR2X1_LOC_45/B AND2X1_LOC_776/Y 0.10fF
C36594 OR2X1_LOC_45/B OR2X1_LOC_135/Y 0.02fF
C36670 OR2X1_LOC_45/B AND2X1_LOC_520/Y 0.28fF
C36768 OR2X1_LOC_45/B AND2X1_LOC_856/B 1.24fF
C36773 OR2X1_LOC_45/B AND2X1_LOC_464/Y 0.01fF
C37080 OR2X1_LOC_45/B AND2X1_LOC_160/a_8_24# 0.01fF
C37686 OR2X1_LOC_45/B AND2X1_LOC_318/Y 0.01fF
C37911 OR2X1_LOC_45/B OR2X1_LOC_697/a_8_216# 0.01fF
C38344 OR2X1_LOC_45/B AND2X1_LOC_508/A 0.03fF
C38691 OR2X1_LOC_45/B OR2X1_LOC_183/a_36_216# 0.03fF
C38962 OR2X1_LOC_45/B AND2X1_LOC_634/Y 0.04fF
C39172 OR2X1_LOC_45/B OR2X1_LOC_230/Y 0.03fF
C39630 OR2X1_LOC_45/B AND2X1_LOC_715/A 0.02fF
C40106 OR2X1_LOC_45/B AND2X1_LOC_778/a_8_24# 0.01fF
C40306 OR2X1_LOC_45/B OR2X1_LOC_172/Y 0.25fF
C41003 OR2X1_LOC_45/B OR2X1_LOC_280/Y 0.08fF
C41967 OR2X1_LOC_45/B OR2X1_LOC_226/Y 0.06fF
C42282 OR2X1_LOC_45/B OR2X1_LOC_680/A 0.18fF
C42761 OR2X1_LOC_45/B OR2X1_LOC_423/a_8_216# 0.02fF
C43633 OR2X1_LOC_45/B OR2X1_LOC_609/A 0.08fF
C44019 OR2X1_LOC_45/B AND2X1_LOC_266/Y 1.81fF
C44292 OR2X1_LOC_45/B OR2X1_LOC_183/Y 0.02fF
C44869 OR2X1_LOC_45/B OR2X1_LOC_237/Y 0.33fF
C44914 OR2X1_LOC_45/B OR2X1_LOC_487/a_8_216# 0.07fF
C46006 OR2X1_LOC_45/B OR2X1_LOC_423/Y 0.03fF
C46248 OR2X1_LOC_45/B OR2X1_LOC_74/A 13.05fF
C47009 OR2X1_LOC_45/B AND2X1_LOC_448/a_8_24# 0.02fF
C47162 OR2X1_LOC_45/B OR2X1_LOC_239/Y 0.01fF
C47893 OR2X1_LOC_45/B AND2X1_LOC_339/B 0.03fF
C47996 OR2X1_LOC_45/B AND2X1_LOC_633/a_8_24# 0.01fF
C49195 OR2X1_LOC_45/B OR2X1_LOC_697/Y 0.18fF
C49328 OR2X1_LOC_45/B OR2X1_LOC_696/Y 0.03fF
C49770 OR2X1_LOC_45/B OR2X1_LOC_431/a_8_216# 0.01fF
C50109 OR2X1_LOC_45/B AND2X1_LOC_303/A 0.01fF
C50544 OR2X1_LOC_45/B OR2X1_LOC_495/a_8_216# 0.09fF
C50672 OR2X1_LOC_45/B OR2X1_LOC_238/a_8_216# 0.02fF
C50925 OR2X1_LOC_45/B OR2X1_LOC_695/a_8_216# 0.02fF
C50951 OR2X1_LOC_45/B AND2X1_LOC_458/Y 0.01fF
C51797 OR2X1_LOC_45/B OR2X1_LOC_305/a_8_216# 0.01fF
C51882 OR2X1_LOC_45/B AND2X1_LOC_537/Y 0.07fF
C52048 OR2X1_LOC_45/B OR2X1_LOC_171/a_8_216# 0.06fF
C52964 OR2X1_LOC_45/B AND2X1_LOC_714/B 0.07fF
C53339 OR2X1_LOC_45/B OR2X1_LOC_406/Y 0.06fF
C53395 OR2X1_LOC_45/B OR2X1_LOC_496/a_8_216# 0.01fF
C53770 OR2X1_LOC_45/B OR2X1_LOC_516/Y 0.10fF
C54638 OR2X1_LOC_45/B OR2X1_LOC_528/a_8_216# 0.06fF
C54760 OR2X1_LOC_45/B OR2X1_LOC_609/a_8_216# 0.40fF
C55063 OR2X1_LOC_45/B VDD 1.30fF
C55132 OR2X1_LOC_45/B OR2X1_LOC_315/Y 0.06fF
C55165 OR2X1_LOC_45/B AND2X1_LOC_267/a_8_24# 0.06fF
C55343 OR2X1_LOC_45/B OR2X1_LOC_67/Y 0.03fF
C56102 OR2X1_LOC_45/B AND2X1_LOC_307/Y 0.01fF
C56174 OR2X1_LOC_45/B OR2X1_LOC_238/a_36_216# 0.03fF
C58129 OR2X1_LOC_45/B VSS -5.64fF
C6 OR2X1_LOC_680/A OR2X1_LOC_89/A 0.03fF
C378 OR2X1_LOC_757/A OR2X1_LOC_89/A 0.73fF
C850 AND2X1_LOC_97/a_8_24# OR2X1_LOC_89/A 0.12fF
C2194 OR2X1_LOC_511/Y OR2X1_LOC_89/A 0.02fF
C2801 OR2X1_LOC_89/A OR2X1_LOC_384/Y 0.13fF
C2944 OR2X1_LOC_89/A OR2X1_LOC_131/a_8_216# 0.01fF
C3931 OR2X1_LOC_74/A OR2X1_LOC_89/A 0.14fF
C3946 OR2X1_LOC_89/A OR2X1_LOC_261/A 0.79fF
C5055 AND2X1_LOC_779/a_8_24# OR2X1_LOC_89/A 0.01fF
C5143 OR2X1_LOC_615/a_8_216# OR2X1_LOC_89/A 0.01fF
C5752 OR2X1_LOC_106/Y OR2X1_LOC_89/A 0.18fF
C6250 OR2X1_LOC_89/A AND2X1_LOC_614/a_8_24# 0.01fF
C6327 AND2X1_LOC_99/A OR2X1_LOC_89/A 0.01fF
C6864 OR2X1_LOC_680/Y OR2X1_LOC_89/A 0.15fF
C6884 OR2X1_LOC_696/Y OR2X1_LOC_89/A 0.01fF
C7122 AND2X1_LOC_362/B OR2X1_LOC_89/A 0.10fF
C7555 AND2X1_LOC_706/Y OR2X1_LOC_89/A 0.01fF
C7719 OR2X1_LOC_665/Y OR2X1_LOC_89/A 0.01fF
C8627 OR2X1_LOC_89/A OR2X1_LOC_89/a_8_216# 0.05fF
C10173 OR2X1_LOC_526/Y OR2X1_LOC_89/A 0.03fF
C11302 OR2X1_LOC_516/Y OR2X1_LOC_89/A 0.03fF
C11681 OR2X1_LOC_89/A AND2X1_LOC_793/B 0.34fF
C12063 OR2X1_LOC_89/A AND2X1_LOC_846/a_8_24# 0.01fF
C12424 OR2X1_LOC_131/Y OR2X1_LOC_89/A 0.01fF
C12713 VDD OR2X1_LOC_89/A 0.78fF
C12753 OR2X1_LOC_677/Y OR2X1_LOC_89/A 0.03fF
C12830 OR2X1_LOC_491/Y OR2X1_LOC_89/A 0.07fF
C12836 OR2X1_LOC_251/Y OR2X1_LOC_89/A 0.05fF
C13694 OR2X1_LOC_89/A OR2X1_LOC_591/A 0.02fF
C13933 OR2X1_LOC_494/A OR2X1_LOC_89/A 0.03fF
C14979 AND2X1_LOC_557/a_8_24# OR2X1_LOC_89/A 0.01fF
C15158 OR2X1_LOC_89/A OR2X1_LOC_184/a_8_216# 0.01fF
C15726 OR2X1_LOC_89/A OR2X1_LOC_767/a_8_216# 0.05fF
C16119 OR2X1_LOC_103/Y OR2X1_LOC_89/A 0.32fF
C16150 OR2X1_LOC_103/a_8_216# OR2X1_LOC_89/A 0.01fF
C16472 OR2X1_LOC_482/Y OR2X1_LOC_89/A 0.17fF
C16512 OR2X1_LOC_816/Y OR2X1_LOC_89/A 0.04fF
C16616 OR2X1_LOC_748/A OR2X1_LOC_89/A 0.01fF
C17117 OR2X1_LOC_89/A OR2X1_LOC_815/A 0.01fF
C17544 OR2X1_LOC_146/Y OR2X1_LOC_89/A 0.08fF
C17569 OR2X1_LOC_89/A AND2X1_LOC_848/A 0.01fF
C17733 OR2X1_LOC_591/Y OR2X1_LOC_89/A 0.01fF
C18131 OR2X1_LOC_89/A AND2X1_LOC_227/a_8_24# 0.01fF
C18791 AND2X1_LOC_840/B OR2X1_LOC_89/A 0.23fF
C18821 OR2X1_LOC_282/a_8_216# OR2X1_LOC_89/A 0.02fF
C19138 OR2X1_LOC_144/Y OR2X1_LOC_89/A 0.10fF
C20369 OR2X1_LOC_89/A AND2X1_LOC_285/Y 0.03fF
C20464 OR2X1_LOC_91/Y OR2X1_LOC_89/A 2.32fF
C20527 OR2X1_LOC_527/Y OR2X1_LOC_89/A 0.84fF
C20536 OR2X1_LOC_417/Y OR2X1_LOC_89/A 0.03fF
C21270 OR2X1_LOC_441/Y OR2X1_LOC_89/A 0.03fF
C21310 OR2X1_LOC_667/Y OR2X1_LOC_89/A 0.02fF
C22442 OR2X1_LOC_146/a_8_216# OR2X1_LOC_89/A 0.01fF
C22612 OR2X1_LOC_525/Y OR2X1_LOC_89/A 0.03fF
C22659 OR2X1_LOC_497/Y OR2X1_LOC_89/A 0.63fF
C23578 AND2X1_LOC_721/A OR2X1_LOC_89/A 0.03fF
C23908 OR2X1_LOC_89/A AND2X1_LOC_361/A 0.09fF
C24346 OR2X1_LOC_282/a_36_216# OR2X1_LOC_89/A 0.02fF
C25102 OR2X1_LOC_257/a_8_216# OR2X1_LOC_89/A 0.06fF
C26511 OR2X1_LOC_89/A OR2X1_LOC_406/A 0.01fF
C27821 OR2X1_LOC_89/A OR2X1_LOC_13/B 0.31fF
C28363 OR2X1_LOC_89/A OR2X1_LOC_595/A 4.49fF
C28929 AND2X1_LOC_105/a_8_24# OR2X1_LOC_89/A 0.09fF
C30195 OR2X1_LOC_89/A OR2X1_LOC_591/a_8_216# 0.01fF
C30243 AND2X1_LOC_727/A OR2X1_LOC_89/A 0.03fF
C30983 OR2X1_LOC_438/Y OR2X1_LOC_89/A 0.03fF
C31020 OR2X1_LOC_89/A AND2X1_LOC_621/Y 13.91fF
C31550 OR2X1_LOC_184/Y OR2X1_LOC_89/A 0.13fF
C32487 OR2X1_LOC_89/A OR2X1_LOC_767/Y 0.06fF
C32981 OR2X1_LOC_89/A OR2X1_LOC_16/A 0.01fF
C33019 OR2X1_LOC_108/Y OR2X1_LOC_89/A 0.07fF
C33960 OR2X1_LOC_109/Y OR2X1_LOC_89/A 0.01fF
C34255 AND2X1_LOC_593/a_8_24# OR2X1_LOC_89/A 0.01fF
C34464 AND2X1_LOC_227/Y OR2X1_LOC_89/A 0.08fF
C34847 OR2X1_LOC_599/A OR2X1_LOC_89/A 1.08fF
C34875 OR2X1_LOC_89/A OR2X1_LOC_258/a_8_216# 0.01fF
C35752 OR2X1_LOC_89/A OR2X1_LOC_615/Y 0.71fF
C36449 OR2X1_LOC_495/Y OR2X1_LOC_89/A 0.03fF
C36550 AND2X1_LOC_664/a_8_24# OR2X1_LOC_89/A 0.01fF
C38612 OR2X1_LOC_503/A OR2X1_LOC_89/A 0.03fF
C39903 AND2X1_LOC_557/Y OR2X1_LOC_89/A 0.01fF
C40223 AND2X1_LOC_456/B OR2X1_LOC_89/A 0.03fF
C40339 OR2X1_LOC_89/A OR2X1_LOC_258/a_36_216# 0.02fF
C41072 OR2X1_LOC_494/Y OR2X1_LOC_89/A 0.03fF
C41930 OR2X1_LOC_89/A AND2X1_LOC_778/Y 0.03fF
C42041 OR2X1_LOC_89/A AND2X1_LOC_624/A 0.03fF
C43500 OR2X1_LOC_89/A AND2X1_LOC_779/Y 0.01fF
C44466 OR2X1_LOC_89/A OR2X1_LOC_89/Y 0.14fF
C44694 OR2X1_LOC_754/A OR2X1_LOC_89/A 0.03fF
C44846 OR2X1_LOC_89/A OR2X1_LOC_142/Y 0.08fF
C45011 OR2X1_LOC_89/A OR2X1_LOC_442/Y 0.11fF
C45125 OR2X1_LOC_89/A OR2X1_LOC_238/Y 0.03fF
C46125 OR2X1_LOC_89/A OR2X1_LOC_152/A 0.14fF
C46268 OR2X1_LOC_177/Y OR2X1_LOC_89/A 0.04fF
C46305 OR2X1_LOC_604/A OR2X1_LOC_89/A 0.23fF
C47285 OR2X1_LOC_164/Y OR2X1_LOC_89/A 0.03fF
C47652 OR2X1_LOC_131/A OR2X1_LOC_89/A 0.69fF
C48304 OR2X1_LOC_89/A AND2X1_LOC_678/a_8_24# 0.05fF
C49069 OR2X1_LOC_89/A AND2X1_LOC_260/a_8_24# 0.01fF
C50371 OR2X1_LOC_79/A OR2X1_LOC_89/A 0.01fF
C50624 OR2X1_LOC_815/a_8_216# OR2X1_LOC_89/A 0.01fF
C50742 OR2X1_LOC_89/A AND2X1_LOC_848/Y 0.03fF
C51682 OR2X1_LOC_89/A OR2X1_LOC_815/Y 0.01fF
C51886 OR2X1_LOC_759/A OR2X1_LOC_89/A 0.04fF
C51920 OR2X1_LOC_698/Y OR2X1_LOC_89/A 0.03fF
C52066 OR2X1_LOC_224/Y OR2X1_LOC_89/A 0.03fF
C54063 AND2X1_LOC_729/Y OR2X1_LOC_89/A 0.03fF
C54527 AND2X1_LOC_489/Y OR2X1_LOC_89/A 1.15fF
C54554 OR2X1_LOC_755/A OR2X1_LOC_89/A 0.01fF
C54636 OR2X1_LOC_89/A AND2X1_LOC_216/A 0.16fF
C54952 OR2X1_LOC_280/Y OR2X1_LOC_89/A 0.03fF
C55789 AND2X1_LOC_593/Y OR2X1_LOC_89/A 0.03fF
C55896 OR2X1_LOC_89/A OR2X1_LOC_226/Y 0.21fF
C56998 OR2X1_LOC_89/A VSS 0.77fF
C11528 AND2X1_LOC_56/B OR2X1_LOC_83/A 0.03fF
C23487 OR2X1_LOC_83/A OR2X1_LOC_240/A 0.03fF
C42424 OR2X1_LOC_83/A OR2X1_LOC_394/a_8_216# 0.01fF
C46381 OR2X1_LOC_83/A OR2X1_LOC_394/Y 0.01fF
C57122 OR2X1_LOC_83/A VSS 0.20fF
C3071 OR2X1_LOC_261/Y OR2X1_LOC_748/A 0.01fF
C4233 OR2X1_LOC_748/A AND2X1_LOC_848/a_8_24# 0.01fF
C4809 OR2X1_LOC_748/A AND2X1_LOC_848/A 0.04fF
C8132 OR2X1_LOC_748/A OR2X1_LOC_701/a_8_216# 0.01fF
C9176 OR2X1_LOC_748/A AND2X1_LOC_789/Y 0.28fF
C17783 OR2X1_LOC_748/A OR2X1_LOC_297/a_8_216# 0.01fF
C19819 OR2X1_LOC_748/A OR2X1_LOC_759/Y 0.01fF
C23769 OR2X1_LOC_748/A OR2X1_LOC_261/a_8_216# 0.01fF
C29200 OR2X1_LOC_748/A AND2X1_LOC_709/a_8_24# 0.07fF
C33420 OR2X1_LOC_604/A OR2X1_LOC_748/A 0.04fF
C34683 OR2X1_LOC_748/A AND2X1_LOC_711/A 0.27fF
C35548 OR2X1_LOC_748/A OR2X1_LOC_700/a_8_216# 0.01fF
C37731 OR2X1_LOC_748/A AND2X1_LOC_848/Y 0.04fF
C38644 OR2X1_LOC_748/A OR2X1_LOC_258/Y 0.03fF
C38932 OR2X1_LOC_759/A OR2X1_LOC_748/A 0.59fF
C38986 OR2X1_LOC_698/Y OR2X1_LOC_748/A 0.09fF
C40161 OR2X1_LOC_748/A AND2X1_LOC_709/a_36_24# 0.01fF
C41195 OR2X1_LOC_481/Y OR2X1_LOC_748/A 0.01fF
C45541 OR2X1_LOC_748/A OR2X1_LOC_297/Y 0.01fF
C47383 OR2X1_LOC_748/A OR2X1_LOC_261/A 0.02fF
C49420 OR2X1_LOC_748/A AND2X1_LOC_847/Y 0.01fF
C53215 OR2X1_LOC_700/Y OR2X1_LOC_748/A 0.01fF
C57524 OR2X1_LOC_748/A VSS -1.10fF
C14254 VDD OR2X1_LOC_693/Y 0.16fF
C26930 OR2X1_LOC_692/Y OR2X1_LOC_693/Y 0.21fF
C37879 OR2X1_LOC_693/Y AND2X1_LOC_706/a_8_24# 0.23fF
C57688 OR2X1_LOC_693/Y VSS 0.07fF
C16153 OR2X1_LOC_673/a_8_216# OR2X1_LOC_673/A 0.08fF
C18905 OR2X1_LOC_673/A OR2X1_LOC_532/B 0.61fF
C20914 VDD OR2X1_LOC_673/A 0.26fF
C27558 AND2X1_LOC_91/B OR2X1_LOC_673/A 0.09fF
C31456 OR2X1_LOC_235/B OR2X1_LOC_673/A 0.01fF
C55767 OR2X1_LOC_673/B OR2X1_LOC_673/A 0.04fF
C57155 OR2X1_LOC_673/A VSS 0.21fF
C7898 OR2X1_LOC_177/Y OR2X1_LOC_164/Y 0.03fF
C7932 OR2X1_LOC_604/A OR2X1_LOC_164/Y 0.07fF
C11688 AND2X1_LOC_776/Y OR2X1_LOC_164/Y 0.04fF
C21720 OR2X1_LOC_164/Y OR2X1_LOC_74/A 0.02fF
C30409 VDD OR2X1_LOC_164/Y 0.29fF
C36402 OR2X1_LOC_164/Y AND2X1_LOC_840/B 0.11fF
C38068 OR2X1_LOC_91/Y OR2X1_LOC_164/Y 0.10fF
C38138 OR2X1_LOC_527/Y OR2X1_LOC_164/Y 0.13fF
C42225 AND2X1_LOC_787/A OR2X1_LOC_164/Y 0.02fF
C51872 OR2X1_LOC_109/Y OR2X1_LOC_164/Y 0.78fF
C54719 AND2X1_LOC_776/a_8_24# OR2X1_LOC_164/Y 0.01fF
C57325 OR2X1_LOC_164/Y VSS 0.40fF
C4019 OR2X1_LOC_368/Y OR2X1_LOC_322/Y 0.01fF
C4829 OR2X1_LOC_322/Y OR2X1_LOC_323/Y 0.78fF
C10970 OR2X1_LOC_74/A OR2X1_LOC_322/Y 0.10fF
C18917 OR2X1_LOC_368/a_8_216# OR2X1_LOC_322/Y 0.03fF
C19799 VDD OR2X1_LOC_322/Y 0.49fF
C19875 OR2X1_LOC_315/Y OR2X1_LOC_322/Y 0.02fF
C20605 AND2X1_LOC_457/a_8_24# OR2X1_LOC_322/Y 0.02fF
C26098 AND2X1_LOC_464/A OR2X1_LOC_322/Y 0.01fF
C27475 OR2X1_LOC_91/Y OR2X1_LOC_322/Y 0.07fF
C31581 AND2X1_LOC_787/A OR2X1_LOC_322/Y 0.03fF
C32450 AND2X1_LOC_543/a_8_24# OR2X1_LOC_322/Y 0.04fF
C34669 OR2X1_LOC_312/Y OR2X1_LOC_322/Y 0.15fF
C40965 OR2X1_LOC_109/Y OR2X1_LOC_322/Y 0.48fF
C43464 AND2X1_LOC_543/Y OR2X1_LOC_322/Y 0.23fF
C53387 OR2X1_LOC_177/Y OR2X1_LOC_322/Y 0.02fF
C56300 OR2X1_LOC_322/Y VSS 0.33fF
C47858 VDD OR2X1_LOC_376/Y -0.00fF
C56345 OR2X1_LOC_376/Y VSS 0.10fF
C5398 OR2X1_LOC_380/Y OR2X1_LOC_588/Y 0.73fF
C8118 AND2X1_LOC_379/a_8_24# OR2X1_LOC_588/Y 0.06fF
C13655 OR2X1_LOC_380/A OR2X1_LOC_588/Y 0.06fF
C33983 OR2X1_LOC_588/Y AND2X1_LOC_637/Y 0.14fF
C40159 VDD OR2X1_LOC_588/Y 0.05fF
C49977 OR2X1_LOC_409/B OR2X1_LOC_588/Y 0.81fF
C50618 OR2X1_LOC_380/a_8_216# OR2X1_LOC_588/Y 0.01fF
C56639 OR2X1_LOC_588/Y VSS 0.24fF
C7734 OR2X1_LOC_696/Y OR2X1_LOC_591/a_8_216# 0.57fF
C12415 OR2X1_LOC_599/A OR2X1_LOC_696/Y 0.01fF
C21266 AND2X1_LOC_160/Y OR2X1_LOC_696/Y 0.15fF
C23820 OR2X1_LOC_604/A OR2X1_LOC_696/Y 0.02fF
C40260 OR2X1_LOC_697/Y OR2X1_LOC_696/Y 0.44fF
C46341 VDD OR2X1_LOC_696/Y 0.15fF
C47377 OR2X1_LOC_696/Y OR2X1_LOC_591/A 0.15fF
C57562 OR2X1_LOC_696/Y VSS 0.28fF
C31814 OR2X1_LOC_503/A OR2X1_LOC_497/Y 0.79fF
C57755 OR2X1_LOC_503/A VSS 0.21fF
C8379 AND2X1_LOC_539/Y OR2X1_LOC_306/Y 0.02fF
C9308 OR2X1_LOC_306/Y AND2X1_LOC_434/Y 0.03fF
C11553 OR2X1_LOC_306/Y AND2X1_LOC_856/B 0.16fF
C12617 OR2X1_LOC_306/Y OR2X1_LOC_829/A 0.15fF
C29609 OR2X1_LOC_306/Y VDD 0.01fF
C29689 OR2X1_LOC_306/Y OR2X1_LOC_829/a_8_216# 0.39fF
C35221 OR2X1_LOC_306/Y AND2X1_LOC_390/B 0.04fF
C36100 OR2X1_LOC_306/Y AND2X1_LOC_308/a_8_24# 0.10fF
C37365 OR2X1_LOC_306/Y OR2X1_LOC_311/Y 0.04fF
C44801 OR2X1_LOC_306/Y OR2X1_LOC_13/B 0.05fF
C47378 OR2X1_LOC_306/Y AND2X1_LOC_727/A 0.01fF
C51146 OR2X1_LOC_306/Y AND2X1_LOC_729/B 0.03fF
C57960 OR2X1_LOC_306/Y VSS 0.37fF
C2444 VDD OR2X1_LOC_144/Y 0.19fF
C2492 OR2X1_LOC_677/Y OR2X1_LOC_144/Y 0.12fF
C20788 OR2X1_LOC_144/Y AND2X1_LOC_621/Y 0.19fF
C24323 OR2X1_LOC_679/A OR2X1_LOC_144/Y 0.01fF
C34505 OR2X1_LOC_144/Y OR2X1_LOC_142/Y 0.06fF
C37764 OR2X1_LOC_144/Y AND2X1_LOC_678/a_8_24# 0.24fF
C43709 AND2X1_LOC_729/Y OR2X1_LOC_144/Y 0.31fF
C49858 OR2X1_LOC_144/Y OR2X1_LOC_74/A 0.07fF
C52796 OR2X1_LOC_680/Y OR2X1_LOC_144/Y 0.01fF
C56030 OR2X1_LOC_526/Y OR2X1_LOC_144/Y 0.01fF
C57278 OR2X1_LOC_144/Y VSS 0.07fF
C1986 OR2X1_LOC_78/A OR2X1_LOC_630/B 0.03fF
C2876 OR2X1_LOC_501/B OR2X1_LOC_630/B 1.11fF
C8427 OR2X1_LOC_499/B OR2X1_LOC_630/B 0.02fF
C13525 OR2X1_LOC_629/Y OR2X1_LOC_630/B 0.07fF
C27528 AND2X1_LOC_56/B OR2X1_LOC_630/B 0.01fF
C30050 OR2X1_LOC_630/a_8_216# OR2X1_LOC_630/B 0.05fF
C56579 OR2X1_LOC_630/B VSS 0.22fF
C19582 OR2X1_LOC_448/A AND2X1_LOC_697/a_8_24# 0.20fF
C21544 OR2X1_LOC_448/A OR2X1_LOC_713/A 0.01fF
C28323 VDD OR2X1_LOC_448/A 0.21fF
C57121 OR2X1_LOC_448/A VSS 0.21fF
C4044 OR2X1_LOC_389/A OR2X1_LOC_389/a_8_216# 0.01fF
C20638 OR2X1_LOC_389/A OR2X1_LOC_390/A 0.01fF
C22920 OR2X1_LOC_389/A OR2X1_LOC_537/A 1.13fF
C42023 OR2X1_LOC_389/A OR2X1_LOC_532/B 0.01fF
C57724 OR2X1_LOC_389/A VSS 0.23fF
C13057 OR2X1_LOC_98/B OR2X1_LOC_98/a_8_216# 0.01fF
C24119 OR2X1_LOC_98/B OR2X1_LOC_99/A 0.88fF
C56860 OR2X1_LOC_98/B VSS 0.10fF
C5987 OR2X1_LOC_378/Y AND2X1_LOC_459/a_8_24# 0.01fF
C26270 VDD OR2X1_LOC_378/Y 0.06fF
C30179 AND2X1_LOC_459/Y OR2X1_LOC_378/Y 0.01fF
C56522 OR2X1_LOC_378/Y VSS 0.14fF
C1156 OR2X1_LOC_506/A OR2X1_LOC_776/Y 0.14fF
C3101 OR2X1_LOC_506/A OR2X1_LOC_532/B 0.47fF
C4926 VDD OR2X1_LOC_506/A 0.85fF
C7142 OR2X1_LOC_840/A OR2X1_LOC_506/A 0.05fF
C8342 OR2X1_LOC_506/A OR2X1_LOC_130/Y 0.09fF
C8526 OR2X1_LOC_447/A OR2X1_LOC_506/A 0.07fF
C9013 OR2X1_LOC_506/A AND2X1_LOC_491/a_8_24# 0.17fF
C11725 AND2X1_LOC_91/B OR2X1_LOC_506/A 0.09fF
C11878 OR2X1_LOC_799/A OR2X1_LOC_506/A 0.03fF
C12337 AND2X1_LOC_56/B OR2X1_LOC_506/A 0.07fF
C14173 OR2X1_LOC_506/A AND2X1_LOC_420/a_8_24# 0.05fF
C16620 AND2X1_LOC_680/a_8_24# OR2X1_LOC_506/A 0.01fF
C17199 OR2X1_LOC_506/A OR2X1_LOC_593/B 0.02fF
C18334 OR2X1_LOC_506/A AND2X1_LOC_69/Y 0.13fF
C19217 AND2X1_LOC_69/a_8_24# OR2X1_LOC_506/A 0.17fF
C19534 OR2X1_LOC_506/A OR2X1_LOC_447/a_8_216# 0.08fF
C20013 OR2X1_LOC_506/A OR2X1_LOC_449/B 0.29fF
C27580 OR2X1_LOC_506/A OR2X1_LOC_539/Y 0.03fF
C29332 OR2X1_LOC_506/A AND2X1_LOC_67/Y 0.04fF
C31343 OR2X1_LOC_319/B OR2X1_LOC_506/A 0.07fF
C31356 OR2X1_LOC_318/Y OR2X1_LOC_506/A 0.08fF
C32274 AND2X1_LOC_165/a_8_24# OR2X1_LOC_506/A 0.07fF
C32757 OR2X1_LOC_436/Y OR2X1_LOC_506/A 0.09fF
C33868 AND2X1_LOC_67/a_8_24# OR2X1_LOC_506/A 0.01fF
C36232 OR2X1_LOC_506/A OR2X1_LOC_308/Y 0.05fF
C39379 OR2X1_LOC_506/A AND2X1_LOC_423/a_8_24# 0.20fF
C40706 OR2X1_LOC_810/A OR2X1_LOC_506/A 0.01fF
C42788 OR2X1_LOC_506/A OR2X1_LOC_78/A 0.07fF
C43896 OR2X1_LOC_506/A OR2X1_LOC_318/B 0.02fF
C43910 OR2X1_LOC_506/A OR2X1_LOC_854/A 0.03fF
C44011 OR2X1_LOC_121/Y OR2X1_LOC_506/A 0.01fF
C44089 OR2X1_LOC_538/A OR2X1_LOC_506/A 0.03fF
C45407 OR2X1_LOC_506/A OR2X1_LOC_776/a_8_216# 0.14fF
C47118 OR2X1_LOC_186/Y OR2X1_LOC_506/A 0.03fF
C47617 OR2X1_LOC_493/B OR2X1_LOC_506/A 0.04fF
C47750 OR2X1_LOC_574/A OR2X1_LOC_506/A 0.03fF
C51698 OR2X1_LOC_506/A OR2X1_LOC_728/A 0.03fF
C53419 OR2X1_LOC_506/A OR2X1_LOC_130/a_8_216# 0.01fF
C53880 OR2X1_LOC_97/A OR2X1_LOC_506/A 0.02fF
C57163 OR2X1_LOC_506/A VSS 0.85fF
C8640 OR2X1_LOC_837/Y OR2X1_LOC_838/B 0.07fF
C19663 OR2X1_LOC_838/a_8_216# OR2X1_LOC_838/B 0.05fF
C56822 OR2X1_LOC_838/B VSS 0.22fF
C23103 OR2X1_LOC_541/A OR2X1_LOC_241/B 0.03fF
C23212 OR2X1_LOC_188/Y OR2X1_LOC_541/A 0.02fF
C39014 OR2X1_LOC_541/A OR2X1_LOC_778/A 0.61fF
C44026 OR2X1_LOC_541/A OR2X1_LOC_778/a_8_216# 0.05fF
C51465 OR2X1_LOC_541/A OR2X1_LOC_778/Y 0.01fF
C57305 OR2X1_LOC_541/A VSS 0.37fF
C42667 VDD OR2X1_LOC_138/A -0.00fF
C43513 OR2X1_LOC_676/Y OR2X1_LOC_138/A 0.01fF
C47632 OR2X1_LOC_702/A OR2X1_LOC_138/A 0.27fF
C50132 AND2X1_LOC_56/B OR2X1_LOC_138/A 0.04fF
C56317 OR2X1_LOC_138/A VSS 0.37fF
C4199 OR2X1_LOC_296/Y OR2X1_LOC_78/A 0.01fF
C9284 OR2X1_LOC_296/Y AND2X1_LOC_627/a_8_24# 0.01fF
C10316 OR2X1_LOC_296/Y OR2X1_LOC_629/a_8_216# 0.01fF
C13792 OR2X1_LOC_296/Y OR2X1_LOC_247/a_8_216# 0.01fF
C15705 OR2X1_LOC_629/Y OR2X1_LOC_296/Y 0.75fF
C22550 VDD OR2X1_LOC_296/Y 0.31fF
C27936 OR2X1_LOC_296/Y OR2X1_LOC_294/Y 0.04fF
C35784 OR2X1_LOC_296/Y OR2X1_LOC_247/Y 0.59fF
C39910 OR2X1_LOC_631/B OR2X1_LOC_296/Y 0.01fF
C57308 OR2X1_LOC_296/Y VSS 0.19fF
C41517 VDD OR2X1_LOC_195/A -0.00fF
C51328 OR2X1_LOC_195/A AND2X1_LOC_41/Y 0.23fF
C57464 OR2X1_LOC_195/A VSS 0.21fF
C3669 OR2X1_LOC_319/B OR2X1_LOC_535/A 0.01fF
C12515 OR2X1_LOC_535/A OR2X1_LOC_356/A 0.08fF
C16340 OR2X1_LOC_535/A OR2X1_LOC_538/A 0.02fF
C24951 OR2X1_LOC_703/B OR2X1_LOC_535/A 0.05fF
C40954 OR2X1_LOC_535/A AND2X1_LOC_166/a_8_24# 0.08fF
C42998 OR2X1_LOC_535/A OR2X1_LOC_788/B 0.08fF
C57808 OR2X1_LOC_535/A VSS -0.16fF
C3215 OR2X1_LOC_609/A OR2X1_LOC_71/A 0.02fF
C4031 OR2X1_LOC_673/Y OR2X1_LOC_71/A 0.01fF
C5688 OR2X1_LOC_74/A OR2X1_LOC_71/A 0.04fF
C5955 AND2X1_LOC_235/a_8_24# OR2X1_LOC_71/A 0.01fF
C6495 OR2X1_LOC_235/a_8_216# OR2X1_LOC_71/A 0.01fF
C12598 OR2X1_LOC_532/B OR2X1_LOC_71/A 0.02fF
C14594 VDD OR2X1_LOC_71/A 1.12fF
C14782 OR2X1_LOC_67/Y OR2X1_LOC_71/A 0.03fF
C21369 AND2X1_LOC_91/B OR2X1_LOC_71/A 0.02fF
C21909 AND2X1_LOC_56/B OR2X1_LOC_71/A 0.01fF
C23204 OR2X1_LOC_235/Y OR2X1_LOC_71/A 0.01fF
C25221 OR2X1_LOC_235/B OR2X1_LOC_71/A 0.56fF
C26166 OR2X1_LOC_243/B OR2X1_LOC_71/A 0.01fF
C26327 OR2X1_LOC_771/B OR2X1_LOC_71/A 0.03fF
C27303 OR2X1_LOC_612/a_8_216# OR2X1_LOC_71/A 0.01fF
C32286 OR2X1_LOC_821/Y OR2X1_LOC_71/A 0.35fF
C34513 OR2X1_LOC_246/Y OR2X1_LOC_71/A 0.01fF
C34884 OR2X1_LOC_16/A OR2X1_LOC_71/A 0.10fF
C36351 OR2X1_LOC_813/Y OR2X1_LOC_71/A 0.01fF
C37815 OR2X1_LOC_813/a_8_216# OR2X1_LOC_71/A 0.01fF
C38800 AND2X1_LOC_240/Y OR2X1_LOC_71/A 0.02fF
C40022 AND2X1_LOC_610/a_8_24# OR2X1_LOC_71/A 0.03fF
C45679 OR2X1_LOC_612/B OR2X1_LOC_71/A 0.01fF
C46366 AND2X1_LOC_608/a_8_24# OR2X1_LOC_71/A 0.03fF
C47568 OR2X1_LOC_611/Y OR2X1_LOC_71/A 0.03fF
C48475 OR2X1_LOC_84/A OR2X1_LOC_71/A 0.02fF
C49566 OR2X1_LOC_612/Y OR2X1_LOC_71/A 0.05fF
C51031 OR2X1_LOC_71/A OR2X1_LOC_398/Y -0.01fF
C52486 OR2X1_LOC_78/A OR2X1_LOC_71/A 0.03fF
C56380 OR2X1_LOC_71/A VSS 0.34fF
C7563 VDD OR2X1_LOC_96/B -0.00fF
C36151 OR2X1_LOC_96/B OR2X1_LOC_96/a_8_216# 0.08fF
C41018 OR2X1_LOC_604/A OR2X1_LOC_96/B 0.04fF
C57077 OR2X1_LOC_96/B VSS -0.20fF
C59 OR2X1_LOC_532/B AND2X1_LOC_617/a_8_24# 0.01fF
C513 OR2X1_LOC_643/A OR2X1_LOC_532/B 0.03fF
C521 OR2X1_LOC_532/B OR2X1_LOC_778/Y 0.10fF
C760 AND2X1_LOC_91/B OR2X1_LOC_532/B 0.53fF
C1397 AND2X1_LOC_56/B OR2X1_LOC_532/B 0.27fF
C2942 OR2X1_LOC_532/B OR2X1_LOC_186/a_8_216# 0.01fF
C3005 AND2X1_LOC_521/a_8_24# OR2X1_LOC_532/B 0.01fF
C3017 OR2X1_LOC_532/B OR2X1_LOC_646/B 0.43fF
C3510 OR2X1_LOC_633/Y OR2X1_LOC_532/B 0.01fF
C3846 OR2X1_LOC_621/A OR2X1_LOC_532/B 0.21fF
C4686 OR2X1_LOC_235/B OR2X1_LOC_532/B 0.06fF
C4746 AND2X1_LOC_393/a_8_24# OR2X1_LOC_532/B 0.01fF
C5140 OR2X1_LOC_791/B OR2X1_LOC_532/B 0.04fF
C5468 OR2X1_LOC_532/B OR2X1_LOC_362/A 0.10fF
C5538 OR2X1_LOC_539/A OR2X1_LOC_532/B 0.01fF
C5775 OR2X1_LOC_532/B OR2X1_LOC_771/B 0.06fF
C5786 OR2X1_LOC_532/B OR2X1_LOC_209/A 0.09fF
C5806 OR2X1_LOC_532/B OR2X1_LOC_776/A 0.03fF
C6018 OR2X1_LOC_483/a_36_216# OR2X1_LOC_532/B 0.03fF
C6206 OR2X1_LOC_532/B OR2X1_LOC_593/B 0.03fF
C6239 OR2X1_LOC_506/a_8_216# OR2X1_LOC_532/B 0.05fF
C6395 AND2X1_LOC_492/a_8_24# OR2X1_LOC_532/B 0.04fF
C6949 OR2X1_LOC_532/B OR2X1_LOC_720/B 0.02fF
C7422 OR2X1_LOC_506/B OR2X1_LOC_532/B 0.01fF
C7715 OR2X1_LOC_473/a_8_216# OR2X1_LOC_532/B 0.01fF
C7872 OR2X1_LOC_532/B AND2X1_LOC_485/a_8_24# 0.01fF
C8548 OR2X1_LOC_523/B OR2X1_LOC_532/B 0.01fF
C8675 OR2X1_LOC_532/B AND2X1_LOC_292/a_8_24# 0.17fF
C8726 OR2X1_LOC_532/B AND2X1_LOC_108/a_36_24# 0.01fF
C9066 OR2X1_LOC_532/B OR2X1_LOC_449/B 0.03fF
C9401 OR2X1_LOC_621/B OR2X1_LOC_532/B 0.20fF
C9452 OR2X1_LOC_317/a_8_216# OR2X1_LOC_532/B 0.01fF
C9951 AND2X1_LOC_674/a_8_24# OR2X1_LOC_532/B 0.01fF
C10334 OR2X1_LOC_400/B OR2X1_LOC_532/B 0.03fF
C10738 OR2X1_LOC_240/B OR2X1_LOC_532/B 0.01fF
C11599 OR2X1_LOC_631/B OR2X1_LOC_532/B 0.07fF
C11627 AND2X1_LOC_135/a_8_24# OR2X1_LOC_532/B 0.01fF
C12737 OR2X1_LOC_532/B OR2X1_LOC_355/a_8_216# 0.01fF
C13325 OR2X1_LOC_809/a_8_216# OR2X1_LOC_532/B 0.02fF
C13335 OR2X1_LOC_532/B OR2X1_LOC_240/A 0.02fF
C13341 OR2X1_LOC_633/B OR2X1_LOC_532/B 0.04fF
C13365 OR2X1_LOC_532/B AND2X1_LOC_281/a_8_24# 0.01fF
C13801 OR2X1_LOC_288/A OR2X1_LOC_532/B 0.01fF
C14043 OR2X1_LOC_506/Y OR2X1_LOC_532/B 0.01fF
C14115 OR2X1_LOC_633/a_8_216# OR2X1_LOC_532/B 0.01fF
C14181 OR2X1_LOC_532/B OR2X1_LOC_346/B 0.23fF
C14515 AND2X1_LOC_167/a_8_24# OR2X1_LOC_532/B 0.01fF
C14847 AND2X1_LOC_522/a_8_24# OR2X1_LOC_532/B 0.01fF
C14866 OR2X1_LOC_856/A OR2X1_LOC_532/B 0.02fF
C15347 OR2X1_LOC_330/Y OR2X1_LOC_532/B 0.02fF
C15423 OR2X1_LOC_675/A OR2X1_LOC_532/B -0.00fF
C15725 OR2X1_LOC_768/A OR2X1_LOC_532/B 0.01fF
C16224 OR2X1_LOC_240/a_8_216# OR2X1_LOC_532/B 0.01fF
C16581 AND2X1_LOC_172/a_8_24# OR2X1_LOC_532/B 0.01fF
C16653 OR2X1_LOC_532/B OR2X1_LOC_539/Y 0.07fF
C16910 OR2X1_LOC_532/B OR2X1_LOC_319/Y 0.01fF
C17487 OR2X1_LOC_493/A OR2X1_LOC_532/B 0.18fF
C17734 OR2X1_LOC_198/a_8_216# OR2X1_LOC_532/B 0.01fF
C17927 AND2X1_LOC_536/a_8_24# OR2X1_LOC_532/B 0.01fF
C18430 AND2X1_LOC_67/Y OR2X1_LOC_532/B 0.02fF
C18842 OR2X1_LOC_809/a_36_216# OR2X1_LOC_532/B 0.01fF
C18929 OR2X1_LOC_532/B OR2X1_LOC_705/B 0.01fF
C19709 OR2X1_LOC_532/B OR2X1_LOC_647/B 0.02fF
C20479 OR2X1_LOC_319/B OR2X1_LOC_532/B 0.13fF
C20903 AND2X1_LOC_103/a_8_24# OR2X1_LOC_532/B 0.03fF
C20938 AND2X1_LOC_331/a_8_24# OR2X1_LOC_532/B 0.01fF
C21768 AND2X1_LOC_320/a_8_24# OR2X1_LOC_532/B 0.01fF
C21848 OR2X1_LOC_287/B OR2X1_LOC_532/B 0.05fF
C21877 OR2X1_LOC_76/A OR2X1_LOC_532/B 0.03fF
C21902 OR2X1_LOC_436/Y OR2X1_LOC_532/B 0.03fF
C22251 OR2X1_LOC_532/B OR2X1_LOC_553/A 0.07fF
C23461 OR2X1_LOC_287/A OR2X1_LOC_532/B 0.03fF
C23476 OR2X1_LOC_174/A OR2X1_LOC_532/B 0.01fF
C23484 OR2X1_LOC_435/a_8_216# OR2X1_LOC_532/B 0.02fF
C23507 AND2X1_LOC_482/a_8_24# OR2X1_LOC_532/B 0.06fF
C23938 OR2X1_LOC_137/B OR2X1_LOC_532/B 0.25fF
C24205 OR2X1_LOC_532/B OR2X1_LOC_415/Y 0.51fF
C24286 OR2X1_LOC_532/B AND2X1_LOC_616/a_8_24# 0.01fF
C24397 OR2X1_LOC_532/B OR2X1_LOC_285/B 0.09fF
C25278 OR2X1_LOC_532/B AND2X1_LOC_109/a_8_24# 0.05fF
C25389 OR2X1_LOC_532/B OR2X1_LOC_308/Y 0.03fF
C26007 OR2X1_LOC_664/Y OR2X1_LOC_532/B 0.72fF
C27243 OR2X1_LOC_324/B OR2X1_LOC_532/B 0.23fF
C27267 AND2X1_LOC_142/a_8_24# OR2X1_LOC_532/B 0.01fF
C27278 AND2X1_LOC_314/a_8_24# OR2X1_LOC_532/B 0.01fF
C27288 OR2X1_LOC_243/A OR2X1_LOC_532/B 0.01fF
C27291 OR2X1_LOC_532/B OR2X1_LOC_668/Y 0.02fF
C27643 AND2X1_LOC_311/a_8_24# OR2X1_LOC_532/B 0.06fF
C27792 OR2X1_LOC_532/B OR2X1_LOC_84/A 0.01fF
C28189 OR2X1_LOC_473/Y OR2X1_LOC_532/B 0.04fF
C28245 OR2X1_LOC_532/B OR2X1_LOC_241/B 0.07fF
C28402 OR2X1_LOC_188/Y OR2X1_LOC_532/B 0.03fF
C28537 AND2X1_LOC_492/a_36_24# OR2X1_LOC_532/B 0.01fF
C28590 OR2X1_LOC_193/A OR2X1_LOC_532/B 0.28fF
C28780 OR2X1_LOC_208/A OR2X1_LOC_532/B 0.01fF
C28830 OR2X1_LOC_673/B OR2X1_LOC_532/B 0.03fF
C28863 AND2X1_LOC_131/a_8_24# OR2X1_LOC_532/B 0.03fF
C28957 OR2X1_LOC_537/A OR2X1_LOC_532/B 0.01fF
C29264 OR2X1_LOC_532/B OR2X1_LOC_356/A 0.01fF
C29832 OR2X1_LOC_810/A OR2X1_LOC_532/B 0.01fF
C30138 OR2X1_LOC_715/B OR2X1_LOC_532/B 8.09fF
C31507 OR2X1_LOC_835/B OR2X1_LOC_532/B 0.10fF
C31834 OR2X1_LOC_532/B OR2X1_LOC_78/A 1.08fF
C32738 OR2X1_LOC_147/B OR2X1_LOC_532/B 0.04fF
C32745 OR2X1_LOC_317/A OR2X1_LOC_532/B 0.01fF
C32760 OR2X1_LOC_532/B AND2X1_LOC_669/a_8_24# 0.01fF
C33052 OR2X1_LOC_121/Y OR2X1_LOC_532/B 0.07fF
C33078 OR2X1_LOC_114/B OR2X1_LOC_532/B 0.02fF
C33123 OR2X1_LOC_538/A OR2X1_LOC_532/B 0.04fF
C33218 OR2X1_LOC_532/B AND2X1_LOC_79/Y 0.01fF
C33999 OR2X1_LOC_532/B OR2X1_LOC_623/B 0.06fF
C34429 OR2X1_LOC_254/B OR2X1_LOC_532/B 0.09fF
C34447 OR2X1_LOC_646/A OR2X1_LOC_532/B 0.02fF
C34869 AND2X1_LOC_321/a_8_24# OR2X1_LOC_532/B 0.01fF
C36009 OR2X1_LOC_186/Y OR2X1_LOC_532/B 1.45fF
C36224 OR2X1_LOC_532/B OR2X1_LOC_112/B 0.10fF
C36466 OR2X1_LOC_493/B OR2X1_LOC_532/B 0.21fF
C36566 OR2X1_LOC_574/A OR2X1_LOC_532/B 0.41fF
C36922 OR2X1_LOC_319/a_8_216# OR2X1_LOC_532/B 0.01fF
C36999 AND2X1_LOC_670/a_8_24# OR2X1_LOC_532/B 0.03fF
C37168 OR2X1_LOC_532/B OR2X1_LOC_539/B 0.16fF
C37334 AND2X1_LOC_103/a_36_24# OR2X1_LOC_532/B 0.01fF
C39219 OR2X1_LOC_532/B OR2X1_LOC_330/a_8_216# 0.01fF
C39558 OR2X1_LOC_673/Y OR2X1_LOC_532/B 0.55fF
C40186 OR2X1_LOC_139/A OR2X1_LOC_532/B 0.13fF
C40337 OR2X1_LOC_324/A OR2X1_LOC_532/B 0.01fF
C41662 OR2X1_LOC_668/a_8_216# OR2X1_LOC_532/B 0.01fF
C41681 OR2X1_LOC_703/B OR2X1_LOC_532/B 0.01fF
C41771 OR2X1_LOC_532/B AND2X1_LOC_109/a_36_24# 0.01fF
C42313 OR2X1_LOC_532/B OR2X1_LOC_532/a_8_216# 0.02fF
C42852 OR2X1_LOC_97/A OR2X1_LOC_532/B 1.17fF
C43864 OR2X1_LOC_532/B OR2X1_LOC_720/A 0.01fF
C43977 OR2X1_LOC_532/B OR2X1_LOC_590/a_8_216# 0.18fF
C44424 OR2X1_LOC_532/B OR2X1_LOC_198/A 0.16fF
C44782 AND2X1_LOC_821/a_8_24# OR2X1_LOC_532/B 0.01fF
C45044 OR2X1_LOC_532/B OR2X1_LOC_361/a_8_216# 0.01fF
C45109 OR2X1_LOC_538/a_8_216# OR2X1_LOC_532/B 0.01fF
C45422 OR2X1_LOC_532/B OR2X1_LOC_267/Y 0.02fF
C45466 OR2X1_LOC_673/a_8_216# OR2X1_LOC_532/B 0.04fF
C46391 OR2X1_LOC_532/B OR2X1_LOC_776/Y 0.46fF
C46793 OR2X1_LOC_532/B OR2X1_LOC_355/A 0.01fF
C47876 AND2X1_LOC_79/a_8_24# OR2X1_LOC_532/B 0.01fF
C47891 OR2X1_LOC_287/a_8_216# OR2X1_LOC_532/B 0.01fF
C49462 OR2X1_LOC_532/B OR2X1_LOC_778/a_8_216# 0.01fF
C49511 OR2X1_LOC_76/B OR2X1_LOC_532/B 0.06fF
C50289 VDD OR2X1_LOC_532/B 2.30fF
C50375 AND2X1_LOC_755/a_8_24# OR2X1_LOC_532/B 0.23fF
C50700 OR2X1_LOC_532/B OR2X1_LOC_361/a_36_216# 0.01fF
C50983 OR2X1_LOC_532/B OR2X1_LOC_523/A 0.01fF
C51202 OR2X1_LOC_483/a_8_216# OR2X1_LOC_532/B 0.03fF
C51486 AND2X1_LOC_83/a_8_24# OR2X1_LOC_532/B 0.01fF
C52287 OR2X1_LOC_532/B OR2X1_LOC_115/B 0.03fF
C52425 OR2X1_LOC_840/A OR2X1_LOC_532/B 0.03fF
C52856 OR2X1_LOC_216/A OR2X1_LOC_532/B 0.29fF
C52897 OR2X1_LOC_802/Y OR2X1_LOC_532/B 0.01fF
C52953 AND2X1_LOC_134/a_8_24# OR2X1_LOC_532/B 0.01fF
C53331 OR2X1_LOC_624/B OR2X1_LOC_532/B 0.59fF
C53524 OR2X1_LOC_532/B OR2X1_LOC_532/Y 0.01fF
C53738 OR2X1_LOC_447/A OR2X1_LOC_532/B 0.01fF
C53823 OR2X1_LOC_532/B AND2X1_LOC_108/a_8_24# 0.14fF
C54181 AND2X1_LOC_491/a_8_24# OR2X1_LOC_532/B 0.11fF
C55002 OR2X1_LOC_702/A OR2X1_LOC_532/B 0.03fF
C55731 OR2X1_LOC_532/B OR2X1_LOC_294/Y 0.02fF
C55873 OR2X1_LOC_114/Y OR2X1_LOC_532/B 0.03fF
C57019 OR2X1_LOC_532/B VSS 0.64fF
C333 OR2X1_LOC_78/A OR2X1_LOC_779/a_8_216# 0.01fF
C390 AND2X1_LOC_176/a_8_24# OR2X1_LOC_78/A 0.01fF
C728 AND2X1_LOC_533/a_8_24# OR2X1_LOC_78/A 0.06fF
C1568 OR2X1_LOC_435/B OR2X1_LOC_78/A 0.23fF
C2828 OR2X1_LOC_78/A OR2X1_LOC_777/a_8_216# 0.01fF
C2978 AND2X1_LOC_72/a_8_24# OR2X1_LOC_78/A 0.01fF
C3303 OR2X1_LOC_201/A OR2X1_LOC_78/A 0.04fF
C3404 OR2X1_LOC_647/B OR2X1_LOC_78/A 0.19fF
C4115 OR2X1_LOC_318/Y OR2X1_LOC_78/A 0.07fF
C5009 OR2X1_LOC_629/A OR2X1_LOC_78/A 0.01fF
C5064 AND2X1_LOC_165/a_8_24# OR2X1_LOC_78/A 0.03fF
C5084 OR2X1_LOC_446/Y OR2X1_LOC_78/A 0.01fF
C5420 OR2X1_LOC_287/B OR2X1_LOC_78/A 0.86fF
C5449 OR2X1_LOC_97/a_8_216# OR2X1_LOC_78/A 0.01fF
C5502 OR2X1_LOC_148/A OR2X1_LOC_78/A 0.01fF
C7037 OR2X1_LOC_287/A OR2X1_LOC_78/A -0.00fF
C7063 OR2X1_LOC_435/a_8_216# OR2X1_LOC_78/A 0.01fF
C7896 OR2X1_LOC_78/A OR2X1_LOC_631/A 0.02fF
C7919 OR2X1_LOC_78/A AND2X1_LOC_616/a_8_24# 0.07fF
C8303 OR2X1_LOC_78/A OR2X1_LOC_168/Y 0.42fF
C9122 OR2X1_LOC_78/A OR2X1_LOC_308/Y 0.07fF
C9359 OR2X1_LOC_593/A OR2X1_LOC_78/A 0.01fF
C9734 OR2X1_LOC_664/Y OR2X1_LOC_78/A 0.07fF
C10582 AND2X1_LOC_89/a_8_24# OR2X1_LOC_78/A 0.03fF
C10677 OR2X1_LOC_168/A OR2X1_LOC_78/A 0.05fF
C10751 AND2X1_LOC_280/a_8_24# OR2X1_LOC_78/A 0.02fF
C11742 OR2X1_LOC_190/A OR2X1_LOC_78/A 0.02fF
C11900 OR2X1_LOC_473/Y OR2X1_LOC_78/A 0.03fF
C12201 OR2X1_LOC_78/A AND2X1_LOC_615/a_8_24# 0.01fF
C12569 AND2X1_LOC_505/a_8_24# OR2X1_LOC_78/A 0.02fF
C12971 OR2X1_LOC_710/A OR2X1_LOC_78/A 0.01fF
C13010 OR2X1_LOC_78/A OR2X1_LOC_356/A 0.07fF
C13041 OR2X1_LOC_614/a_36_216# OR2X1_LOC_78/A 0.03fF
C13517 OR2X1_LOC_610/a_8_216# OR2X1_LOC_78/A 0.03fF
C13580 OR2X1_LOC_810/A OR2X1_LOC_78/A 0.12fF
C13581 OR2X1_LOC_307/a_8_216# OR2X1_LOC_78/A 0.01fF
C13600 AND2X1_LOC_589/a_8_24# OR2X1_LOC_78/A 0.02fF
C13866 OR2X1_LOC_715/B OR2X1_LOC_78/A 2.84fF
C13878 OR2X1_LOC_78/A OR2X1_LOC_784/B 0.01fF
C14015 AND2X1_LOC_81/a_8_24# OR2X1_LOC_78/A 0.01fF
C14373 OR2X1_LOC_656/B OR2X1_LOC_78/A 0.01fF
C14809 OR2X1_LOC_687/Y OR2X1_LOC_78/A 0.03fF
C16076 OR2X1_LOC_97/B OR2X1_LOC_78/A 0.08fF
C16382 OR2X1_LOC_501/B OR2X1_LOC_78/A 0.12fF
C16549 OR2X1_LOC_97/a_36_216# OR2X1_LOC_78/A 0.01fF
C16781 OR2X1_LOC_121/Y OR2X1_LOC_78/A 0.07fF
C16809 OR2X1_LOC_114/B OR2X1_LOC_78/A 0.04fF
C16843 OR2X1_LOC_538/A OR2X1_LOC_78/A 0.03fF
C17693 OR2X1_LOC_78/A OR2X1_LOC_623/B 0.01fF
C18086 OR2X1_LOC_140/A OR2X1_LOC_78/A 0.02fF
C18092 OR2X1_LOC_507/A OR2X1_LOC_78/A 0.01fF
C19053 OR2X1_LOC_448/Y OR2X1_LOC_78/A 0.21fF
C19117 OR2X1_LOC_592/A OR2X1_LOC_78/A 0.02fF
C19385 OR2X1_LOC_78/A OR2X1_LOC_629/B 0.02fF
C19802 OR2X1_LOC_186/Y OR2X1_LOC_78/A 0.03fF
C20381 OR2X1_LOC_574/A OR2X1_LOC_78/A 0.29fF
C20637 OR2X1_LOC_78/A AND2X1_LOC_627/a_8_24# 0.01fF
C21172 OR2X1_LOC_448/a_8_216# OR2X1_LOC_78/A 0.03fF
C21663 AND2X1_LOC_89/a_36_24# OR2X1_LOC_78/A 0.01fF
C21700 OR2X1_LOC_629/a_8_216# OR2X1_LOC_78/A 0.01fF
C22015 OR2X1_LOC_499/B OR2X1_LOC_78/A 0.02fF
C23084 OR2X1_LOC_779/Y OR2X1_LOC_78/A 0.01fF
C23323 OR2X1_LOC_115/a_8_216# OR2X1_LOC_78/A 0.02fF
C23371 OR2X1_LOC_673/Y OR2X1_LOC_78/A 0.15fF
C23994 OR2X1_LOC_78/A OR2X1_LOC_712/B 0.05fF
C24047 OR2X1_LOC_139/A OR2X1_LOC_78/A 0.01fF
C25049 AND2X1_LOC_697/a_8_24# OR2X1_LOC_78/A 0.04fF
C25164 OR2X1_LOC_247/a_8_216# OR2X1_LOC_78/A 0.01fF
C25253 OR2X1_LOC_78/A AND2X1_LOC_235/a_8_24# 0.05fF
C25300 AND2X1_LOC_594/a_8_24# OR2X1_LOC_78/A 0.02fF
C25357 AND2X1_LOC_526/a_8_24# OR2X1_LOC_78/A 0.01fF
C25410 OR2X1_LOC_703/B OR2X1_LOC_78/A 0.01fF
C25660 OR2X1_LOC_78/A OR2X1_LOC_844/B 0.42fF
C25765 AND2X1_LOC_177/a_8_24# OR2X1_LOC_78/A 0.02fF
C26533 OR2X1_LOC_97/A OR2X1_LOC_78/A 0.04fF
C26588 OR2X1_LOC_78/A OR2X1_LOC_78/a_8_216# 0.13fF
C26630 OR2X1_LOC_78/A OR2X1_LOC_475/B 0.26fF
C26640 OR2X1_LOC_448/a_36_216# OR2X1_LOC_78/A 0.03fF
C26970 OR2X1_LOC_78/A OR2X1_LOC_713/A 0.07fF
C27076 OR2X1_LOC_629/Y OR2X1_LOC_78/A 0.01fF
C27313 OR2X1_LOC_78/A OR2X1_LOC_546/A 0.01fF
C28021 OR2X1_LOC_778/A OR2X1_LOC_78/A 0.02fF
C28129 OR2X1_LOC_99/A OR2X1_LOC_78/A 0.03fF
C28655 OR2X1_LOC_78/A OR2X1_LOC_361/a_8_216# 0.02fF
C29048 OR2X1_LOC_78/A OR2X1_LOC_267/Y 0.13fF
C29303 AND2X1_LOC_107/a_8_24# OR2X1_LOC_78/A 0.07fF
C29953 OR2X1_LOC_776/Y OR2X1_LOC_78/A 0.43fF
C30150 AND2X1_LOC_677/a_8_24# OR2X1_LOC_78/A 0.01fF
C30742 OR2X1_LOC_78/A OR2X1_LOC_779/A 0.01fF
C30776 OR2X1_LOC_614/Y OR2X1_LOC_78/A 0.74fF
C31630 OR2X1_LOC_78/A OR2X1_LOC_113/B 0.02fF
C31843 AND2X1_LOC_665/a_8_24# OR2X1_LOC_78/A 0.09fF
C32020 OR2X1_LOC_440/B OR2X1_LOC_78/A 0.01fF
C32054 OR2X1_LOC_78/A OR2X1_LOC_78/a_36_216# 0.01fF
C32961 AND2X1_LOC_503/a_8_24# OR2X1_LOC_78/A 0.02fF
C33753 OR2X1_LOC_78/A AND2X1_LOC_265/a_8_24# 0.08fF
C33763 VDD OR2X1_LOC_78/A 1.75fF
C34243 OR2X1_LOC_115/a_36_216# OR2X1_LOC_78/A 0.02fF
C34595 OR2X1_LOC_834/A OR2X1_LOC_78/A 0.01fF
C35796 OR2X1_LOC_78/A OR2X1_LOC_115/B 0.12fF
C35905 OR2X1_LOC_840/A OR2X1_LOC_78/A 0.10fF
C36019 AND2X1_LOC_697/a_36_24# OR2X1_LOC_78/A 0.01fF
C36252 AND2X1_LOC_754/a_8_24# OR2X1_LOC_78/A 0.01fF
C36290 AND2X1_LOC_397/a_8_24# OR2X1_LOC_78/A 0.01fF
C36327 OR2X1_LOC_216/A OR2X1_LOC_78/A 0.29fF
C36822 OR2X1_LOC_624/B OR2X1_LOC_78/A 0.07fF
C37060 OR2X1_LOC_196/Y OR2X1_LOC_78/A 0.01fF
C37325 AND2X1_LOC_108/a_8_24# OR2X1_LOC_78/A 0.01fF
C37579 OR2X1_LOC_78/A AND2X1_LOC_424/a_8_24# 0.03fF
C37986 OR2X1_LOC_78/A OR2X1_LOC_708/Y 0.01fF
C38100 OR2X1_LOC_435/Y OR2X1_LOC_78/A 0.04fF
C38820 AND2X1_LOC_262/a_8_24# OR2X1_LOC_78/A 0.01fF
C38853 OR2X1_LOC_78/A AND2X1_LOC_437/a_8_24# 0.04fF
C39225 OR2X1_LOC_294/Y OR2X1_LOC_78/A 0.05fF
C39235 OR2X1_LOC_78/A OR2X1_LOC_641/A 0.03fF
C39374 OR2X1_LOC_114/Y OR2X1_LOC_78/A 0.02fF
C39753 OR2X1_LOC_168/a_8_216# OR2X1_LOC_78/A 0.05fF
C40176 OR2X1_LOC_643/A OR2X1_LOC_78/A 0.05fF
C40182 OR2X1_LOC_778/Y OR2X1_LOC_78/A 0.10fF
C40457 AND2X1_LOC_91/B OR2X1_LOC_78/A 0.19fF
C40594 AND2X1_LOC_72/Y OR2X1_LOC_78/A 0.03fF
C40598 OR2X1_LOC_799/A OR2X1_LOC_78/A 0.23fF
C40820 OR2X1_LOC_78/A OR2X1_LOC_303/B 0.07fF
C40904 OR2X1_LOC_78/A OR2X1_LOC_719/B 0.03fF
C40931 OR2X1_LOC_542/B OR2X1_LOC_78/A 0.04fF
C40975 OR2X1_LOC_105/a_8_216# OR2X1_LOC_78/A 0.02fF
C41016 OR2X1_LOC_631/a_8_216# OR2X1_LOC_78/A 0.01fF
C41057 AND2X1_LOC_56/B OR2X1_LOC_78/A 0.09fF
C41814 OR2X1_LOC_790/A OR2X1_LOC_78/A 0.01fF
C41850 OR2X1_LOC_402/B OR2X1_LOC_78/A 0.38fF
C41954 AND2X1_LOC_118/a_8_24# OR2X1_LOC_78/A 0.01fF
C42938 OR2X1_LOC_78/A OR2X1_LOC_227/Y 0.02fF
C42942 OR2X1_LOC_78/A OR2X1_LOC_284/B 0.12fF
C43049 OR2X1_LOC_78/A OR2X1_LOC_180/B 0.05fF
C43207 OR2X1_LOC_633/Y OR2X1_LOC_78/A 6.10fF
C43453 OR2X1_LOC_78/A OR2X1_LOC_788/B 3.83fF
C43549 OR2X1_LOC_621/A OR2X1_LOC_78/A 0.19fF
C43657 OR2X1_LOC_630/a_8_216# OR2X1_LOC_78/A 0.01fF
C43669 OR2X1_LOC_664/a_8_216# OR2X1_LOC_78/A 0.03fF
C44061 OR2X1_LOC_509/A OR2X1_LOC_78/A 0.04fF
C44457 OR2X1_LOC_235/B OR2X1_LOC_78/A 0.09fF
C44832 AND2X1_LOC_295/a_8_24# OR2X1_LOC_78/A 0.05fF
C44891 OR2X1_LOC_703/A OR2X1_LOC_78/A 0.03fF
C45289 OR2X1_LOC_78/A OR2X1_LOC_362/A 0.66fF
C45637 OR2X1_LOC_78/A OR2X1_LOC_771/B 0.03fF
C45944 AND2X1_LOC_107/a_36_24# OR2X1_LOC_78/A 0.01fF
C46094 OR2X1_LOC_78/A OR2X1_LOC_593/B 0.01fF
C46521 OR2X1_LOC_78/A OR2X1_LOC_317/B 0.03fF
C46677 OR2X1_LOC_105/a_36_216# OR2X1_LOC_78/A 0.03fF
C47353 OR2X1_LOC_506/B OR2X1_LOC_78/A 0.05fF
C47392 OR2X1_LOC_247/Y OR2X1_LOC_78/A 0.01fF
C47490 OR2X1_LOC_78/A AND2X1_LOC_258/a_8_24# 0.03fF
C47506 OR2X1_LOC_78/A OR2X1_LOC_708/a_8_216# 0.01fF
C47959 OR2X1_LOC_78/A OR2X1_LOC_307/A 0.01fF
C48938 OR2X1_LOC_449/B OR2X1_LOC_78/A 0.10fF
C49209 OR2X1_LOC_621/B OR2X1_LOC_78/A 0.39fF
C50079 OR2X1_LOC_786/A OR2X1_LOC_78/A 0.01fF
C50311 OR2X1_LOC_447/Y OR2X1_LOC_78/A 0.10fF
C50484 OR2X1_LOC_346/A OR2X1_LOC_78/A 0.07fF
C51315 OR2X1_LOC_78/A OR2X1_LOC_439/B 0.01fF
C51449 OR2X1_LOC_631/B OR2X1_LOC_78/A 0.08fF
C52174 OR2X1_LOC_284/a_8_216# OR2X1_LOC_78/A 0.02fF
C52256 OR2X1_LOC_632/A OR2X1_LOC_78/A 0.01fF
C52721 OR2X1_LOC_593/a_8_216# OR2X1_LOC_78/A 0.01fF
C52741 AND2X1_LOC_701/a_8_24# OR2X1_LOC_78/A 0.01fF
C52840 OR2X1_LOC_614/a_8_216# OR2X1_LOC_78/A 0.02fF
C53170 OR2X1_LOC_633/B OR2X1_LOC_78/A 0.05fF
C53848 OR2X1_LOC_506/Y OR2X1_LOC_78/A 0.01fF
C53890 OR2X1_LOC_630/Y OR2X1_LOC_78/A 0.01fF
C53901 OR2X1_LOC_633/a_8_216# OR2X1_LOC_78/A 0.01fF
C53988 OR2X1_LOC_346/B OR2X1_LOC_78/A 0.03fF
C54125 OR2X1_LOC_78/A OR2X1_LOC_196/a_8_216# 0.01fF
C54410 OR2X1_LOC_592/a_8_216# OR2X1_LOC_78/A 0.01fF
C54786 OR2X1_LOC_664/a_36_216# OR2X1_LOC_78/A 0.02fF
C55056 OR2X1_LOC_308/A OR2X1_LOC_78/A 0.01fF
C55221 AND2X1_LOC_504/a_8_24# OR2X1_LOC_78/A 0.09fF
C55303 AND2X1_LOC_117/a_8_24# OR2X1_LOC_78/A 0.07fF
C56229 AND2X1_LOC_146/a_8_24# OR2X1_LOC_78/A 0.01fF
C56758 OR2X1_LOC_78/A VSS 0.95fF
C912 AND2X1_LOC_56/B OR2X1_LOC_33/B 0.22fF
C2020 AND2X1_LOC_56/B OR2X1_LOC_729/a_8_216# 0.03fF
C2580 OR2X1_LOC_76/B AND2X1_LOC_56/B 0.12fF
C2687 OR2X1_LOC_472/B AND2X1_LOC_56/B 0.03fF
C2749 AND2X1_LOC_56/B OR2X1_LOC_552/A 0.02fF
C2773 AND2X1_LOC_56/B OR2X1_LOC_151/a_8_216# 0.02fF
C3166 AND2X1_LOC_56/B OR2X1_LOC_192/B 0.09fF
C3347 VDD AND2X1_LOC_56/B 1.30fF
C3515 AND2X1_LOC_56/B OR2X1_LOC_444/B 0.01fF
C3802 OR2X1_LOC_334/B AND2X1_LOC_56/B 0.02fF
C4138 OR2X1_LOC_676/Y AND2X1_LOC_56/B 0.01fF
C4241 OR2X1_LOC_462/B AND2X1_LOC_56/B 0.03fF
C5135 AND2X1_LOC_56/B OR2X1_LOC_416/Y 0.16fF
C5423 OR2X1_LOC_840/A AND2X1_LOC_56/B 0.10fF
C6535 AND2X1_LOC_56/B OR2X1_LOC_532/Y 0.01fF
C6754 AND2X1_LOC_56/B OR2X1_LOC_447/A 0.01fF
C7340 AND2X1_LOC_56/B OR2X1_LOC_620/A 0.01fF
C8163 OR2X1_LOC_702/A AND2X1_LOC_56/B 0.84fF
C8311 AND2X1_LOC_56/B OR2X1_LOC_151/a_36_216# 0.03fF
C8913 AND2X1_LOC_312/a_8_24# AND2X1_LOC_56/B 0.12fF
C8956 OR2X1_LOC_379/Y AND2X1_LOC_56/B 0.03fF
C9785 AND2X1_LOC_56/B OR2X1_LOC_637/A 0.17fF
C9854 AND2X1_LOC_56/B OR2X1_LOC_778/Y 0.10fF
C10056 AND2X1_LOC_91/B AND2X1_LOC_56/B 0.16fF
C10533 AND2X1_LOC_56/B OR2X1_LOC_719/B 0.02fF
C10563 AND2X1_LOC_56/B OR2X1_LOC_542/B 0.12fF
C10963 AND2X1_LOC_56/B OR2X1_LOC_787/B 0.01fF
C12182 AND2X1_LOC_56/B OR2X1_LOC_34/A 0.03fF
C12309 AND2X1_LOC_56/B OR2X1_LOC_828/a_8_216# 0.01fF
C12467 AND2X1_LOC_56/B AND2X1_LOC_420/a_8_24# 0.03fF
C14977 AND2X1_LOC_56/B AND2X1_LOC_680/a_8_24# 0.03fF
C15094 AND2X1_LOC_56/B OR2X1_LOC_771/B 0.03fF
C15100 AND2X1_LOC_56/B OR2X1_LOC_209/A 0.03fF
C17976 AND2X1_LOC_56/B AND2X1_LOC_39/Y 0.04fF
C18331 AND2X1_LOC_56/B OR2X1_LOC_449/B 0.07fF
C18672 OR2X1_LOC_317/a_8_216# AND2X1_LOC_56/B 0.03fF
C20071 OR2X1_LOC_461/Y AND2X1_LOC_56/B 0.01fF
C22025 AND2X1_LOC_56/B OR2X1_LOC_355/a_8_216# 0.03fF
C22626 AND2X1_LOC_597/a_8_24# AND2X1_LOC_56/B 0.01fF
C23265 AND2X1_LOC_56/B OR2X1_LOC_334/A 0.03fF
C23422 AND2X1_LOC_586/a_8_24# AND2X1_LOC_56/B 0.04fF
C23555 AND2X1_LOC_56/B AND2X1_LOC_420/a_36_24# 0.01fF
C24171 AND2X1_LOC_56/B OR2X1_LOC_730/A 0.02fF
C24637 OR2X1_LOC_330/Y AND2X1_LOC_56/B 0.02fF
C25523 AND2X1_LOC_56/B AND2X1_LOC_298/a_8_24# 0.11fF
C26821 AND2X1_LOC_56/B AND2X1_LOC_13/a_8_24# 0.02fF
C30113 AND2X1_LOC_331/a_8_24# AND2X1_LOC_56/B 0.04fF
C30226 AND2X1_LOC_56/B AND2X1_LOC_825/a_8_24# 0.03fF
C30929 AND2X1_LOC_498/a_8_24# AND2X1_LOC_56/B 0.13fF
C30931 AND2X1_LOC_320/a_8_24# AND2X1_LOC_56/B 0.03fF
C31413 AND2X1_LOC_56/B OR2X1_LOC_553/A 0.07fF
C32645 AND2X1_LOC_56/B AND2X1_LOC_482/a_8_24# 0.01fF
C33331 AND2X1_LOC_56/B OR2X1_LOC_415/Y 0.02fF
C34174 AND2X1_LOC_56/B OR2X1_LOC_334/a_8_216# 0.01fF
C34324 AND2X1_LOC_586/a_36_24# AND2X1_LOC_56/B 0.01fF
C34556 AND2X1_LOC_56/B OR2X1_LOC_308/Y 0.07fF
C35044 AND2X1_LOC_56/B OR2X1_LOC_828/Y 0.01fF
C35349 AND2X1_LOC_56/B OR2X1_LOC_181/A 0.02fF
C35552 AND2X1_LOC_56/B AND2X1_LOC_24/a_8_24# 0.05fF
C36390 OR2X1_LOC_324/B AND2X1_LOC_56/B 0.01fF
C36432 AND2X1_LOC_314/a_8_24# AND2X1_LOC_56/B 0.03fF
C36522 OR2X1_LOC_462/a_8_216# AND2X1_LOC_56/B 0.05fF
C37448 AND2X1_LOC_56/B OR2X1_LOC_241/B 0.38fF
C37550 OR2X1_LOC_188/Y AND2X1_LOC_56/B 0.06fF
C37660 AND2X1_LOC_56/B AND2X1_LOC_189/a_8_24# 0.01fF
C37780 AND2X1_LOC_56/B OR2X1_LOC_193/A 0.03fF
C38017 OR2X1_LOC_598/Y AND2X1_LOC_56/B 0.06fF
C38254 AND2X1_LOC_56/B AND2X1_LOC_826/a_8_24# 0.10fF
C38520 AND2X1_LOC_56/B AND2X1_LOC_39/a_8_24# 0.02fF
C39328 OR2X1_LOC_715/B AND2X1_LOC_56/B 0.14fF
C39332 AND2X1_LOC_56/B AND2X1_LOC_626/a_8_24# 0.01fF
C39885 AND2X1_LOC_56/B OR2X1_LOC_793/A 0.03fF
C40191 OR2X1_LOC_837/Y AND2X1_LOC_56/B 0.01fF
C40271 OR2X1_LOC_687/Y AND2X1_LOC_56/B 1.64fF
C40539 AND2X1_LOC_56/B AND2X1_LOC_829/a_8_24# 0.18fF
C41101 AND2X1_LOC_331/a_36_24# AND2X1_LOC_56/B 0.01fF
C41941 OR2X1_LOC_501/B AND2X1_LOC_56/B 0.24fF
C41943 AND2X1_LOC_320/a_36_24# AND2X1_LOC_56/B 0.01fF
C41977 OR2X1_LOC_147/B AND2X1_LOC_56/B 0.06fF
C41996 OR2X1_LOC_317/A AND2X1_LOC_56/B 0.05fF
C42116 AND2X1_LOC_56/B OR2X1_LOC_545/B 0.03fF
C42167 AND2X1_LOC_56/B OR2X1_LOC_318/B 5.14fF
C42319 OR2X1_LOC_121/Y AND2X1_LOC_56/B 0.09fF
C42521 AND2X1_LOC_56/B AND2X1_LOC_496/a_8_24# 0.01fF
C42921 AND2X1_LOC_56/B AND2X1_LOC_495/a_8_24# 0.04fF
C43286 AND2X1_LOC_56/B OR2X1_LOC_623/B 1.47fF
C43746 AND2X1_LOC_56/B OR2X1_LOC_833/B 0.01fF
C44159 AND2X1_LOC_321/a_8_24# AND2X1_LOC_56/B 0.04fF
C44865 AND2X1_LOC_56/B OR2X1_LOC_397/Y 0.03fF
C44934 AND2X1_LOC_56/B OR2X1_LOC_629/B 0.01fF
C45319 AND2X1_LOC_56/B OR2X1_LOC_338/A 0.20fF
C45346 OR2X1_LOC_186/Y AND2X1_LOC_56/B 0.11fF
C45973 OR2X1_LOC_574/A AND2X1_LOC_56/B 0.10fF
C45980 AND2X1_LOC_56/B OR2X1_LOC_33/A 0.04fF
C46207 AND2X1_LOC_56/B OR2X1_LOC_855/A 0.03fF
C46364 AND2X1_LOC_56/B AND2X1_LOC_16/a_8_24# -0.00fF
C47044 AND2X1_LOC_56/B OR2X1_LOC_515/Y 0.01fF
C47681 OR2X1_LOC_499/B AND2X1_LOC_56/B 0.03fF
C47879 AND2X1_LOC_56/B OR2X1_LOC_543/a_8_216# 0.01fF
C48166 AND2X1_LOC_56/B OR2X1_LOC_181/B 0.07fF
C48713 AND2X1_LOC_56/B OR2X1_LOC_330/a_8_216# 0.02fF
C49320 OR2X1_LOC_676/a_8_216# AND2X1_LOC_56/B 0.01fF
C49517 AND2X1_LOC_56/B AND2X1_LOC_27/a_8_24# 0.01fF
C49838 OR2X1_LOC_324/A AND2X1_LOC_56/B 0.10fF
C50046 AND2X1_LOC_56/B OR2X1_LOC_728/A 0.05fF
C51738 AND2X1_LOC_56/B OR2X1_LOC_532/a_8_216# 0.04fF
C51926 AND2X1_LOC_56/B OR2X1_LOC_194/B 0.04fF
C52293 OR2X1_LOC_302/B AND2X1_LOC_56/B 0.15fF
C52479 AND2X1_LOC_56/B AND2X1_LOC_613/a_8_24# 0.01fF
C52768 OR2X1_LOC_629/Y AND2X1_LOC_56/B 0.17fF
C53727 AND2X1_LOC_56/B OR2X1_LOC_778/A 0.01fF
C53822 AND2X1_LOC_56/B OR2X1_LOC_198/A 0.02fF
C54144 AND2X1_LOC_56/B AND2X1_LOC_821/a_8_24# 0.05fF
C54960 AND2X1_LOC_56/B OR2X1_LOC_34/B 0.01fF
C56034 AND2X1_LOC_56/B OR2X1_LOC_355/A 0.05fF
C56089 AND2X1_LOC_56/B OR2X1_LOC_370/a_8_216# 0.07fF
C57405 AND2X1_LOC_56/B VSS 0.91fF
C3962 OR2X1_LOC_611/Y OR2X1_LOC_612/B 0.06fF
C41582 OR2X1_LOC_611/Y OR2X1_LOC_612/a_8_216# 0.39fF
C49386 OR2X1_LOC_611/Y OR2X1_LOC_16/A 0.01fF
C57462 OR2X1_LOC_611/Y VSS 0.18fF
C251 AND2X1_LOC_91/B AND2X1_LOC_399/a_36_24# 0.01fF
C1063 AND2X1_LOC_91/B OR2X1_LOC_391/A 0.62fF
C2763 AND2X1_LOC_91/B VDD 4.07fF
C2988 AND2X1_LOC_91/B OR2X1_LOC_845/A 0.17fF
C4159 AND2X1_LOC_91/B OR2X1_LOC_602/B 0.04fF
C4759 AND2X1_LOC_91/B OR2X1_LOC_115/B 0.34fF
C4851 AND2X1_LOC_91/B OR2X1_LOC_840/A 0.10fF
C5767 AND2X1_LOC_91/B OR2X1_LOC_624/B 0.07fF
C5997 AND2X1_LOC_91/B OR2X1_LOC_532/Y 0.01fF
C6510 AND2X1_LOC_91/B OR2X1_LOC_78/Y 0.06fF
C9179 AND2X1_LOC_91/B AND2X1_LOC_384/a_36_24# 0.01fF
C9227 AND2X1_LOC_91/B OR2X1_LOC_643/A 0.34fF
C9233 AND2X1_LOC_91/B OR2X1_LOC_778/Y 0.14fF
C10000 AND2X1_LOC_91/B OR2X1_LOC_105/a_8_216# 0.01fF
C10472 AND2X1_LOC_91/B AND2X1_LOC_166/a_8_24# 0.05fF
C11996 AND2X1_LOC_91/B OR2X1_LOC_180/B 0.03fF
C12416 AND2X1_LOC_91/B OR2X1_LOC_788/B 0.04fF
C13416 AND2X1_LOC_91/B OR2X1_LOC_235/B 0.01fF
C14227 AND2X1_LOC_91/B OR2X1_LOC_362/A 0.03fF
C14234 AND2X1_LOC_91/B OR2X1_LOC_832/a_8_216# 0.28fF
C14554 AND2X1_LOC_91/B OR2X1_LOC_771/B 0.03fF
C14577 AND2X1_LOC_91/B OR2X1_LOC_776/A 0.10fF
C15030 AND2X1_LOC_91/B AND2X1_LOC_766/a_8_24# 0.05fF
C15346 AND2X1_LOC_91/B OR2X1_LOC_317/B 0.03fF
C16719 AND2X1_LOC_91/B OR2X1_LOC_307/A 0.09fF
C16813 AND2X1_LOC_91/B AND2X1_LOC_394/a_8_24# 0.01fF
C17236 AND2X1_LOC_91/B OR2X1_LOC_447/a_8_216# 0.02fF
C17629 AND2X1_LOC_91/B AND2X1_LOC_487/a_8_24# 0.02fF
C18195 AND2X1_LOC_91/B OR2X1_LOC_383/Y 0.05fF
C19071 AND2X1_LOC_91/B OR2X1_LOC_447/Y 0.24fF
C20268 AND2X1_LOC_91/B OR2X1_LOC_631/B 0.03fF
C20935 AND2X1_LOC_91/B OR2X1_LOC_704/a_8_216# 0.01fF
C21058 AND2X1_LOC_91/B OR2X1_LOC_105/Y 0.03fF
C22378 AND2X1_LOC_91/B AND2X1_LOC_305/a_8_24# 0.05fF
C22809 AND2X1_LOC_91/B OR2X1_LOC_630/Y 0.10fF
C22852 AND2X1_LOC_91/B OR2X1_LOC_447/a_36_216# 0.02fF
C23221 AND2X1_LOC_91/B OR2X1_LOC_392/A 0.01fF
C23597 AND2X1_LOC_91/B AND2X1_LOC_313/a_8_24# 0.01fF
C23763 AND2X1_LOC_91/B AND2X1_LOC_494/a_8_24# 0.05fF
C25259 AND2X1_LOC_91/B OR2X1_LOC_832/a_36_216# 0.01fF
C25378 AND2X1_LOC_91/B AND2X1_LOC_176/a_8_24# 0.06fF
C27845 AND2X1_LOC_91/B OR2X1_LOC_400/A 0.01fF
C28674 AND2X1_LOC_91/B OR2X1_LOC_489/B -0.02fF
C28751 AND2X1_LOC_91/B OR2X1_LOC_401/A 0.03fF
C29058 AND2X1_LOC_91/B OR2X1_LOC_319/B 0.07fF
C30422 AND2X1_LOC_91/B OR2X1_LOC_287/B 0.06fF
C31869 AND2X1_LOC_91/B OR2X1_LOC_714/A 0.01fF
C32458 AND2X1_LOC_91/B AND2X1_LOC_166/a_36_24# 0.01fF
C32899 AND2X1_LOC_91/B AND2X1_LOC_251/a_8_24# 0.02fF
C33201 AND2X1_LOC_91/B OR2X1_LOC_168/Y 0.09fF
C34031 AND2X1_LOC_91/B OR2X1_LOC_308/Y 0.16fF
C34694 AND2X1_LOC_91/B AND2X1_LOC_494/a_36_24# -0.02fF
C35031 AND2X1_LOC_91/B AND2X1_LOC_601/a_8_24# 0.04fF
C35849 AND2X1_LOC_91/B AND2X1_LOC_314/a_8_24# 0.03fF
C35940 AND2X1_LOC_91/B AND2X1_LOC_816/a_8_24# 0.02fF
C36210 AND2X1_LOC_91/B OR2X1_LOC_841/A 0.14fF
C36341 AND2X1_LOC_91/B AND2X1_LOC_176/a_36_24# 0.01fF
C36407 AND2X1_LOC_91/B OR2X1_LOC_84/A 0.02fF
C37849 AND2X1_LOC_91/B OR2X1_LOC_356/A 0.42fF
C38201 AND2X1_LOC_91/B OR2X1_LOC_558/A 0.01fF
C38401 AND2X1_LOC_91/B OR2X1_LOC_810/A 0.10fF
C39049 AND2X1_LOC_91/B OR2X1_LOC_398/Y 0.49fF
C39240 AND2X1_LOC_91/B AND2X1_LOC_767/a_8_24# 0.04fF
C39705 AND2X1_LOC_91/B AND2X1_LOC_399/a_8_24# 0.02fF
C39758 AND2X1_LOC_91/B OR2X1_LOC_401/B 0.18fF
C40400 AND2X1_LOC_91/B AND2X1_LOC_91/a_8_24# 0.05fF
C40522 AND2X1_LOC_91/B OR2X1_LOC_602/A 0.05fF
C41413 AND2X1_LOC_91/B OR2X1_LOC_383/a_8_216# 0.08fF
C41591 AND2X1_LOC_91/B OR2X1_LOC_318/B 0.03fF
C41749 AND2X1_LOC_91/B OR2X1_LOC_114/B 0.03fF
C41758 AND2X1_LOC_91/B AND2X1_LOC_396/a_8_24# 0.04fF
C41768 AND2X1_LOC_91/B OR2X1_LOC_538/A 0.03fF
C41874 AND2X1_LOC_91/B AND2X1_LOC_79/Y 0.03fF
C42292 AND2X1_LOC_91/B AND2X1_LOC_495/a_8_24# 0.16fF
C44759 OR2X1_LOC_186/Y AND2X1_LOC_91/B 0.03fF
C44853 AND2X1_LOC_91/B OR2X1_LOC_773/B 0.03fF
C46534 AND2X1_LOC_91/B OR2X1_LOC_843/B 0.08fF
C47194 AND2X1_LOC_91/B OR2X1_LOC_846/A 0.01fF
C48163 AND2X1_LOC_91/B OR2X1_LOC_330/a_8_216# 0.04fF
C48435 AND2X1_LOC_91/B OR2X1_LOC_673/Y 0.12fF
C48775 AND2X1_LOC_91/B AND2X1_LOC_384/a_8_24# 0.09fF
C50501 AND2X1_LOC_91/B OR2X1_LOC_703/B 0.06fF
C50560 AND2X1_LOC_91/B AND2X1_LOC_815/a_8_24# 0.01fF
C50795 AND2X1_LOC_91/B OR2X1_LOC_844/B 0.29fF
C50955 AND2X1_LOC_91/B OR2X1_LOC_403/B 0.04fF
C51165 AND2X1_LOC_91/B OR2X1_LOC_532/a_8_216# 0.05fF
C51474 AND2X1_LOC_91/B AND2X1_LOC_250/a_8_24# 0.15fF
C51649 AND2X1_LOC_91/B OR2X1_LOC_97/A 0.08fF
C52071 AND2X1_LOC_91/B OR2X1_LOC_713/A 0.14fF
C52542 AND2X1_LOC_91/B AND2X1_LOC_700/a_8_24# 0.11fF
C52598 AND2X1_LOC_91/B AND2X1_LOC_314/a_36_24# 0.01fF
C53464 AND2X1_LOC_91/B AND2X1_LOC_395/a_8_24# 0.04fF
C53617 AND2X1_LOC_91/B AND2X1_LOC_813/a_8_24# 0.01fF
C54184 AND2X1_LOC_91/B OR2X1_LOC_673/a_8_216# 0.49fF
C54799 AND2X1_LOC_91/B AND2X1_LOC_600/a_8_24# 0.09fF
C58013 AND2X1_LOC_91/B VSS 0.75fF
C7141 OR2X1_LOC_297/a_8_216# AND2X1_LOC_847/Y 0.03fF
C8572 AND2X1_LOC_847/Y OR2X1_LOC_701/a_36_216# 0.01fF
C13115 OR2X1_LOC_261/a_8_216# AND2X1_LOC_847/Y 0.01fF
C18225 OR2X1_LOC_297/a_36_216# AND2X1_LOC_847/Y 0.01fF
C19621 OR2X1_LOC_481/a_8_216# AND2X1_LOC_847/Y 0.03fF
C24976 AND2X1_LOC_847/Y OR2X1_LOC_700/a_8_216# 0.03fF
C25129 OR2X1_LOC_481/a_36_216# AND2X1_LOC_847/Y 0.01fF
C27187 AND2X1_LOC_847/Y AND2X1_LOC_848/Y 0.02fF
C30453 AND2X1_LOC_847/Y OR2X1_LOC_700/a_36_216# 0.01fF
C30588 OR2X1_LOC_481/Y AND2X1_LOC_847/Y 0.02fF
C34817 OR2X1_LOC_297/Y AND2X1_LOC_847/Y 0.02fF
C36500 OR2X1_LOC_261/A AND2X1_LOC_847/Y 0.02fF
C42436 OR2X1_LOC_700/Y AND2X1_LOC_847/Y 0.02fF
C45357 VDD AND2X1_LOC_847/Y 0.88fF
C48143 OR2X1_LOC_701/Y AND2X1_LOC_847/Y 0.02fF
C48594 OR2X1_LOC_261/Y AND2X1_LOC_847/Y 0.02fF
C49831 AND2X1_LOC_847/Y AND2X1_LOC_848/a_8_24# 0.01fF
C50425 AND2X1_LOC_848/A AND2X1_LOC_847/Y 0.23fF
C53664 AND2X1_LOC_847/Y OR2X1_LOC_701/a_8_216# 0.03fF
C54661 AND2X1_LOC_847/Y AND2X1_LOC_789/Y 0.02fF
C56881 AND2X1_LOC_847/Y VSS 0.05fF
C14404 OR2X1_LOC_450/B OR2X1_LOC_449/B 0.39fF
C53449 OR2X1_LOC_450/A OR2X1_LOC_450/B 0.12fF
C55543 VDD OR2X1_LOC_450/B 0.21fF
C57635 OR2X1_LOC_450/B VSS 0.01fF
C5282 OR2X1_LOC_303/A OR2X1_LOC_302/A 0.86fF
C18185 AND2X1_LOC_298/a_8_24# OR2X1_LOC_302/A 0.08fF
C27337 OR2X1_LOC_302/A OR2X1_LOC_308/Y 0.14fF
C44851 OR2X1_LOC_302/B OR2X1_LOC_302/A 0.01fF
C50497 OR2X1_LOC_302/a_8_216# OR2X1_LOC_302/A 0.01fF
C52147 VDD OR2X1_LOC_302/A -0.00fF
C56550 OR2X1_LOC_302/A VSS -0.05fF
C33069 VDD OR2X1_LOC_606/Y 0.05fF
C36410 OR2X1_LOC_606/Y AND2X1_LOC_607/a_8_24# 0.01fF
C41974 OR2X1_LOC_606/Y OR2X1_LOC_646/B 0.01fF
C42570 OR2X1_LOC_606/Y OR2X1_LOC_99/Y 1.08fF
C57183 OR2X1_LOC_606/Y VSS 0.10fF
C14740 OR2X1_LOC_147/B OR2X1_LOC_543/A 0.05fF
C14970 OR2X1_LOC_543/A OR2X1_LOC_318/B 0.20fF
C20503 OR2X1_LOC_543/A OR2X1_LOC_543/a_8_216# 0.01fF
C28654 OR2X1_LOC_543/A OR2X1_LOC_370/a_8_216# 0.01fF
C31474 OR2X1_LOC_543/A OR2X1_LOC_552/A -0.00fF
C39668 OR2X1_LOC_543/A OR2X1_LOC_787/B 0.03fF
C43148 OR2X1_LOC_703/A OR2X1_LOC_543/A 0.30fF
C56651 OR2X1_LOC_543/A VSS 0.19fF
C2543 OR2X1_LOC_831/A OR2X1_LOC_76/A 0.05fF
C13700 OR2X1_LOC_831/A OR2X1_LOC_318/B 0.76fF
C32901 OR2X1_LOC_840/A OR2X1_LOC_831/A 0.01fF
C37185 OR2X1_LOC_831/A OR2X1_LOC_778/Y 0.05fF
C37812 OR2X1_LOC_831/A OR2X1_LOC_303/B 0.61fF
C43019 OR2X1_LOC_831/A OR2X1_LOC_593/B 0.04fF
C57670 OR2X1_LOC_831/A VSS 0.39fF
C7890 OR2X1_LOC_121/Y AND2X1_LOC_67/a_8_24# 0.23fF
C9153 OR2X1_LOC_121/Y OR2X1_LOC_631/A 0.02fF
C13824 OR2X1_LOC_121/Y AND2X1_LOC_131/a_8_24# 0.01fF
C14775 OR2X1_LOC_121/Y OR2X1_LOC_810/A 0.10fF
C15075 OR2X1_LOC_121/Y OR2X1_LOC_715/B 0.08fF
C24495 OR2X1_LOC_121/Y OR2X1_LOC_115/a_8_216# 0.03fF
C25242 OR2X1_LOC_121/Y OR2X1_LOC_139/A 0.10fF
C34996 OR2X1_LOC_121/Y VDD 0.81fF
C35446 OR2X1_LOC_121/Y OR2X1_LOC_115/a_36_216# 0.01fF
C37536 OR2X1_LOC_121/Y OR2X1_LOC_216/A 0.01fF
C38267 OR2X1_LOC_121/Y OR2X1_LOC_130/Y 0.01fF
C41445 OR2X1_LOC_121/Y OR2X1_LOC_643/A 0.43fF
C46232 OR2X1_LOC_121/Y OR2X1_LOC_116/a_8_216# 0.02fF
C46653 OR2X1_LOC_121/Y OR2X1_LOC_116/A 0.01fF
C51828 OR2X1_LOC_121/Y OR2X1_LOC_116/a_36_216# 0.01fF
C55242 OR2X1_LOC_121/Y AND2X1_LOC_122/a_8_24# 0.02fF
C58099 OR2X1_LOC_121/Y VSS 0.03fF
C406 VDD OR2X1_LOC_815/A -0.00fF
C38115 OR2X1_LOC_815/a_8_216# OR2X1_LOC_815/A 0.47fF
C39445 OR2X1_LOC_759/A OR2X1_LOC_815/A 0.01fF
C42144 OR2X1_LOC_755/A OR2X1_LOC_815/A 0.04fF
C44201 OR2X1_LOC_757/A OR2X1_LOC_815/A 0.01fF
C56938 OR2X1_LOC_815/A VSS 0.15fF
C4827 AND2X1_LOC_227/Y OR2X1_LOC_226/Y 0.80fF
C16574 OR2X1_LOC_604/A OR2X1_LOC_226/Y 0.01fF
C22357 OR2X1_LOC_224/Y OR2X1_LOC_226/Y 0.04fF
C39044 VDD OR2X1_LOC_226/Y 0.04fF
C44548 OR2X1_LOC_226/Y AND2X1_LOC_227/a_8_24# 0.01fF
C49094 OR2X1_LOC_497/Y OR2X1_LOC_226/Y 0.11fF
C56952 OR2X1_LOC_226/Y VSS 0.08fF
C479 OR2X1_LOC_417/Y OR2X1_LOC_418/Y 0.34fF
C1657 AND2X1_LOC_714/B OR2X1_LOC_417/Y 0.15fF
C3827 VDD OR2X1_LOC_417/Y 0.46fF
C4549 AND2X1_LOC_799/a_36_24# OR2X1_LOC_417/Y 0.01fF
C9516 OR2X1_LOC_417/Y AND2X1_LOC_390/B 0.07fF
C9764 OR2X1_LOC_417/Y OR2X1_LOC_604/Y 0.23fF
C11579 OR2X1_LOC_417/Y AND2X1_LOC_446/a_8_24# 0.01fF
C14630 OR2X1_LOC_417/Y OR2X1_LOC_604/a_8_216# 0.01fF
C14679 OR2X1_LOC_417/Y OR2X1_LOC_331/Y 0.07fF
C17094 OR2X1_LOC_417/Y AND2X1_LOC_454/A 0.01fF
C18951 OR2X1_LOC_417/Y OR2X1_LOC_13/B 0.07fF
C19972 AND2X1_LOC_592/Y OR2X1_LOC_417/Y 0.03fF
C20134 OR2X1_LOC_417/Y AND2X1_LOC_712/B 0.01fF
C21439 OR2X1_LOC_417/Y AND2X1_LOC_727/A 0.03fF
C25067 OR2X1_LOC_417/Y AND2X1_LOC_447/Y 0.07fF
C25986 OR2X1_LOC_599/A OR2X1_LOC_417/Y 0.03fF
C26307 AND2X1_LOC_535/a_8_24# OR2X1_LOC_417/Y 0.04fF
C26670 OR2X1_LOC_176/a_8_216# OR2X1_LOC_417/Y 0.01fF
C35703 OR2X1_LOC_417/Y OR2X1_LOC_601/Y 0.03fF
C37257 OR2X1_LOC_604/A OR2X1_LOC_417/Y 0.09fF
C37275 AND2X1_LOC_535/a_36_24# OR2X1_LOC_417/Y 0.01fF
C37621 OR2X1_LOC_176/Y OR2X1_LOC_417/Y 0.30fF
C38467 AND2X1_LOC_539/Y OR2X1_LOC_417/Y 0.03fF
C45122 AND2X1_LOC_729/Y OR2X1_LOC_417/Y 0.07fF
C45138 AND2X1_LOC_784/A OR2X1_LOC_417/Y 0.03fF
C46883 OR2X1_LOC_417/Y AND2X1_LOC_593/Y 0.07fF
C48159 OR2X1_LOC_417/Y AND2X1_LOC_436/Y 0.03fF
C48243 OR2X1_LOC_417/Y OR2X1_LOC_603/a_8_216# 0.01fF
C48637 OR2X1_LOC_417/Y OR2X1_LOC_313/Y 0.10fF
C49763 AND2X1_LOC_799/a_8_24# OR2X1_LOC_417/Y 0.03fF
C52309 AND2X1_LOC_704/a_8_24# OR2X1_LOC_417/Y 0.01fF
C54811 OR2X1_LOC_417/Y OR2X1_LOC_603/Y 0.01fF
C54817 AND2X1_LOC_706/Y OR2X1_LOC_417/Y 0.39fF
C57621 OR2X1_LOC_417/Y VSS -0.57fF
C2182 AND2X1_LOC_339/B OR2X1_LOC_289/Y 0.04fF
C9462 VDD OR2X1_LOC_289/Y 0.12fF
C17391 OR2X1_LOC_289/Y OR2X1_LOC_171/Y 0.29fF
C28219 AND2X1_LOC_333/a_8_24# OR2X1_LOC_289/Y 0.05fF
C43437 OR2X1_LOC_289/Y OR2X1_LOC_265/Y 0.03fF
C57098 OR2X1_LOC_289/Y VSS 0.09fF
C3525 OR2X1_LOC_487/a_8_216# OR2X1_LOC_488/Y 0.40fF
C13604 VDD OR2X1_LOC_488/Y 0.08fF
C14580 OR2X1_LOC_487/Y OR2X1_LOC_488/Y 0.08fF
C47258 OR2X1_LOC_604/A OR2X1_LOC_488/Y 0.05fF
C57313 OR2X1_LOC_488/Y VSS 0.22fF
C398 OR2X1_LOC_283/Y AND2X1_LOC_843/Y 0.80fF
C5421 AND2X1_LOC_456/B OR2X1_LOC_283/Y 0.01fF
C20029 OR2X1_LOC_283/Y AND2X1_LOC_286/Y 0.10fF
C33865 VDD OR2X1_LOC_283/Y 0.04fF
C33984 OR2X1_LOC_251/Y OR2X1_LOC_283/Y 0.16fF
C47217 OR2X1_LOC_283/Y AND2X1_LOC_286/a_8_24# 0.10fF
C51519 OR2X1_LOC_283/Y AND2X1_LOC_843/a_8_24# 0.04fF
C57433 OR2X1_LOC_283/Y VSS 0.22fF
C1933 VDD OR2X1_LOC_309/Y 0.12fF
C10481 OR2X1_LOC_309/Y AND2X1_LOC_335/a_8_24# 0.23fF
C16927 OR2X1_LOC_309/Y OR2X1_LOC_312/Y 0.03fF
C25361 OR2X1_LOC_309/Y AND2X1_LOC_841/B 0.03fF
C43212 AND2X1_LOC_784/A OR2X1_LOC_309/Y 0.05fF
C57815 OR2X1_LOC_309/Y VSS 0.19fF
C1455 OR2X1_LOC_400/A OR2X1_LOC_398/Y 0.01fF
C10066 OR2X1_LOC_84/A OR2X1_LOC_398/Y 0.43fF
C13386 AND2X1_LOC_399/a_8_24# OR2X1_LOC_398/Y 0.09fF
C21887 OR2X1_LOC_673/Y OR2X1_LOC_398/Y 0.01fF
C24427 OR2X1_LOC_403/B OR2X1_LOC_398/Y 0.01fF
C32288 VDD OR2X1_LOC_398/Y 0.09fF
C43002 OR2X1_LOC_235/B OR2X1_LOC_398/Y 0.05fF
C44146 OR2X1_LOC_771/B OR2X1_LOC_398/Y 0.03fF
C46540 AND2X1_LOC_394/a_8_24# OR2X1_LOC_398/Y 0.01fF
C56341 OR2X1_LOC_398/Y VSS 0.29fF
C12065 OR2X1_LOC_598/Y AND2X1_LOC_829/a_8_24# 0.08fF
C17571 OR2X1_LOC_598/Y OR2X1_LOC_855/A 0.45fF
C25171 OR2X1_LOC_598/Y OR2X1_LOC_198/A 0.02fF
C27474 OR2X1_LOC_379/a_8_216# OR2X1_LOC_598/Y 0.01fF
C29478 OR2X1_LOC_855/a_8_216# OR2X1_LOC_598/Y 0.01fF
C30769 VDD OR2X1_LOC_598/Y 0.12fF
C36321 OR2X1_LOC_379/Y OR2X1_LOC_598/Y 0.01fF
C37120 OR2X1_LOC_598/Y OR2X1_LOC_637/A 0.26fF
C50965 AND2X1_LOC_586/a_8_24# OR2X1_LOC_598/Y 0.24fF
C55637 OR2X1_LOC_644/B OR2X1_LOC_598/Y 0.02fF
C57595 OR2X1_LOC_598/Y VSS 0.45fF
C5831 OR2X1_LOC_810/A OR2X1_LOC_631/A 0.03fF
C12694 OR2X1_LOC_574/A OR2X1_LOC_631/A 0.04fF
C28203 OR2X1_LOC_631/A OR2X1_LOC_115/B 0.03fF
C56751 OR2X1_LOC_631/A VSS 0.19fF
C5603 OR2X1_LOC_415/Y AND2X1_LOC_416/a_8_24# 0.11fF
C20622 AND2X1_LOC_96/a_8_24# OR2X1_LOC_415/Y 0.17fF
C26093 VDD OR2X1_LOC_415/Y 0.50fF
C26114 OR2X1_LOC_98/A OR2X1_LOC_415/Y 0.13fF
C42704 OR2X1_LOC_240/B OR2X1_LOC_415/Y 0.05fF
C43299 OR2X1_LOC_415/Y OR2X1_LOC_396/Y 0.02fF
C45332 OR2X1_LOC_240/A OR2X1_LOC_415/Y 0.44fF
C53864 OR2X1_LOC_240/a_36_216# OR2X1_LOC_415/Y 0.03fF
C54134 OR2X1_LOC_395/Y OR2X1_LOC_415/Y 0.28fF
C56469 OR2X1_LOC_415/Y VSS 0.26fF
C1496 VDD OR2X1_LOC_294/Y 0.41fF
C8748 OR2X1_LOC_542/B OR2X1_LOC_294/Y 0.03fF
C10669 OR2X1_LOC_294/Y OR2X1_LOC_284/B 0.01fF
C12510 OR2X1_LOC_294/Y AND2X1_LOC_295/a_8_24# 0.07fF
C14936 OR2X1_LOC_247/Y OR2X1_LOC_294/Y 0.02fF
C16014 AND2X1_LOC_292/a_8_24# OR2X1_LOC_294/Y 0.01fF
C18020 OR2X1_LOC_294/Y OR2X1_LOC_346/A 0.01fF
C18553 OR2X1_LOC_294/Y AND2X1_LOC_297/a_8_24# 0.01fF
C19008 OR2X1_LOC_631/B OR2X1_LOC_294/Y 0.03fF
C21618 OR2X1_LOC_346/B OR2X1_LOC_294/Y 0.01fF
C24121 OR2X1_LOC_294/Y OR2X1_LOC_347/B 0.01fF
C24448 AND2X1_LOC_184/a_8_24# OR2X1_LOC_294/Y 0.01fF
C30710 OR2X1_LOC_294/Y AND2X1_LOC_279/a_8_24# 0.01fF
C33364 OR2X1_LOC_664/Y OR2X1_LOC_294/Y 0.03fF
C35364 OR2X1_LOC_190/A OR2X1_LOC_294/Y 0.39fF
C40071 OR2X1_LOC_147/B OR2X1_LOC_294/Y 0.03fF
C40468 OR2X1_LOC_114/B OR2X1_LOC_294/Y 0.01fF
C42628 OR2X1_LOC_294/Y AND2X1_LOC_248/a_8_24# 0.01fF
C49013 OR2X1_LOC_247/a_8_216# OR2X1_LOC_294/Y 0.40fF
C53814 OR2X1_LOC_294/Y OR2X1_LOC_342/A 0.01fF
C56770 OR2X1_LOC_294/Y VSS 0.29fF
C7954 VDD OR2X1_LOC_637/B 0.21fF
C13571 OR2X1_LOC_379/Y OR2X1_LOC_637/B 0.01fF
C14381 OR2X1_LOC_637/A OR2X1_LOC_637/B 0.14fF
C19081 AND2X1_LOC_380/a_8_24# OR2X1_LOC_637/B 0.20fF
C30903 OR2X1_LOC_637/B OR2X1_LOC_637/a_8_216# 0.07fF
C37158 OR2X1_LOC_769/A OR2X1_LOC_637/B 0.32fF
C53810 OR2X1_LOC_637/B OR2X1_LOC_769/a_8_216# 0.01fF
C57289 OR2X1_LOC_637/B VSS 0.26fF
C954 OR2X1_LOC_287/B AND2X1_LOC_816/a_8_24# 0.01fF
C3485 OR2X1_LOC_287/B OR2X1_LOC_810/A 0.05fF
C4248 AND2X1_LOC_767/a_8_24# OR2X1_LOC_287/B 0.01fF
C4736 OR2X1_LOC_287/B OR2X1_LOC_401/B 0.01fF
C6390 OR2X1_LOC_287/B OR2X1_LOC_843/a_8_216# 0.19fF
C6706 AND2X1_LOC_396/a_8_24# OR2X1_LOC_287/B 0.01fF
C11369 OR2X1_LOC_287/B OR2X1_LOC_843/B 0.27fF
C15363 OR2X1_LOC_287/B AND2X1_LOC_815/a_8_24# 0.01fF
C16285 OR2X1_LOC_287/B AND2X1_LOC_250/a_8_24# 0.01fF
C16337 OR2X1_LOC_287/B OR2X1_LOC_349/B 0.02fF
C16517 OR2X1_LOC_287/B OR2X1_LOC_78/a_8_216# 0.01fF
C17484 OR2X1_LOC_287/B OR2X1_LOC_850/A 0.01fF
C21180 OR2X1_LOC_770/B OR2X1_LOC_287/B -0.00fF
C21423 OR2X1_LOC_287/B OR2X1_LOC_287/a_8_216# 0.02fF
C21874 OR2X1_LOC_287/B OR2X1_LOC_343/B 0.01fF
C23789 VDD OR2X1_LOC_287/B 0.91fF
C26280 OR2X1_LOC_287/B AND2X1_LOC_397/a_8_24# 0.01fF
C27569 OR2X1_LOC_287/B OR2X1_LOC_78/Y 0.03fF
C28062 OR2X1_LOC_287/B OR2X1_LOC_249/Y 0.02fF
C30976 OR2X1_LOC_105/a_8_216# OR2X1_LOC_287/B 0.01fF
C31775 OR2X1_LOC_287/B OR2X1_LOC_402/B 0.01fF
C32314 OR2X1_LOC_287/B OR2X1_LOC_287/a_36_216# 0.03fF
C34816 OR2X1_LOC_791/B OR2X1_LOC_287/B 0.02fF
C35113 OR2X1_LOC_287/B OR2X1_LOC_362/A 0.06fF
C35391 OR2X1_LOC_287/B OR2X1_LOC_771/B 0.03fF
C35899 AND2X1_LOC_766/a_8_24# OR2X1_LOC_287/B 0.01fF
C41994 OR2X1_LOC_105/Y OR2X1_LOC_287/B 0.03fF
C49884 OR2X1_LOC_489/B OR2X1_LOC_287/B -0.00fF
C49943 OR2X1_LOC_287/B OR2X1_LOC_401/A 0.01fF
C53165 OR2X1_LOC_287/B OR2X1_LOC_287/A 0.01fF
C55802 OR2X1_LOC_287/B OR2X1_LOC_664/Y 0.03fF
C57802 OR2X1_LOC_287/B VSS 0.33fF
C370 AND2X1_LOC_634/Y OR2X1_LOC_16/A 0.01fF
C1556 AND2X1_LOC_729/Y OR2X1_LOC_16/A 0.03fF
C3207 OR2X1_LOC_536/Y OR2X1_LOC_16/A 0.01fF
C4893 OR2X1_LOC_313/Y OR2X1_LOC_16/A 0.08fF
C4933 OR2X1_LOC_609/A OR2X1_LOC_16/A 0.48fF
C7557 OR2X1_LOC_74/A OR2X1_LOC_16/A 0.09fF
C8738 AND2X1_LOC_537/a_8_24# OR2X1_LOC_16/A 0.02fF
C9132 AND2X1_LOC_339/B OR2X1_LOC_16/A 0.05fF
C10013 OR2X1_LOC_16/A OR2X1_LOC_597/a_8_216# 0.01fF
C10621 OR2X1_LOC_167/Y OR2X1_LOC_16/A 0.03fF
C11245 OR2X1_LOC_58/Y OR2X1_LOC_16/A 0.03fF
C11332 AND2X1_LOC_303/A OR2X1_LOC_16/A 0.06fF
C13020 OR2X1_LOC_290/a_8_216# OR2X1_LOC_16/A 0.01fF
C13175 AND2X1_LOC_537/Y OR2X1_LOC_16/A 0.03fF
C15977 OR2X1_LOC_314/Y OR2X1_LOC_16/A 0.05fF
C16320 VDD OR2X1_LOC_16/A 1.24fF
C16766 OR2X1_LOC_60/Y OR2X1_LOC_16/A 0.09fF
C16807 OR2X1_LOC_314/a_8_216# OR2X1_LOC_16/A 0.05fF
C17346 AND2X1_LOC_307/Y OR2X1_LOC_16/A 0.14fF
C18228 OR2X1_LOC_416/Y OR2X1_LOC_16/A 0.05fF
C21583 AND2X1_LOC_317/a_8_24# OR2X1_LOC_16/A 0.04fF
C21903 OR2X1_LOC_765/a_8_216# OR2X1_LOC_16/A 0.06fF
C21999 OR2X1_LOC_316/Y OR2X1_LOC_16/A 0.05fF
C22062 AND2X1_LOC_390/B OR2X1_LOC_16/A 0.07fF
C22819 AND2X1_LOC_301/a_8_24# OR2X1_LOC_16/A 0.01fF
C24085 OR2X1_LOC_290/Y OR2X1_LOC_16/A 0.15fF
C24146 OR2X1_LOC_305/Y OR2X1_LOC_16/A 0.03fF
C24220 OR2X1_LOC_311/Y OR2X1_LOC_16/A 0.03fF
C24233 OR2X1_LOC_601/a_8_216# OR2X1_LOC_16/A 0.03fF
C24391 OR2X1_LOC_16/A OR2X1_LOC_171/Y 0.13fF
C24938 AND2X1_LOC_436/B OR2X1_LOC_16/A 0.02fF
C26973 OR2X1_LOC_235/B OR2X1_LOC_16/A 0.65fF
C27048 AND2X1_LOC_319/A OR2X1_LOC_16/A 0.05fF
C27118 OR2X1_LOC_52/a_8_216# OR2X1_LOC_16/A 0.01fF
C29032 AND2X1_LOC_729/a_8_24# OR2X1_LOC_16/A 0.01fF
C29047 OR2X1_LOC_612/a_8_216# OR2X1_LOC_16/A -0.00fF
C29059 OR2X1_LOC_166/a_8_216# OR2X1_LOC_16/A 0.02fF
C29597 OR2X1_LOC_232/a_8_216# OR2X1_LOC_16/A 0.02fF
C29654 AND2X1_LOC_334/a_8_24# OR2X1_LOC_16/A 0.01fF
C29671 OR2X1_LOC_601/a_36_216# OR2X1_LOC_16/A 0.03fF
C31297 OR2X1_LOC_312/Y OR2X1_LOC_16/A 0.05fF
C31389 OR2X1_LOC_75/a_8_216# OR2X1_LOC_16/A 0.01fF
C31498 OR2X1_LOC_16/A OR2X1_LOC_13/B 0.10fF
C32844 OR2X1_LOC_765/Y OR2X1_LOC_16/A 0.04fF
C33259 OR2X1_LOC_167/a_8_216# OR2X1_LOC_16/A 0.01fF
C34537 OR2X1_LOC_166/a_36_216# OR2X1_LOC_16/A 0.03fF
C35082 OR2X1_LOC_232/a_36_216# OR2X1_LOC_16/A 0.03fF
C36203 OR2X1_LOC_584/a_8_216# OR2X1_LOC_16/A 0.06fF
C36811 AND2X1_LOC_687/Y OR2X1_LOC_16/A 0.01fF
C37495 AND2X1_LOC_447/Y OR2X1_LOC_16/A 0.02fF
C37498 AND2X1_LOC_334/Y OR2X1_LOC_16/A 0.01fF
C37628 AND2X1_LOC_729/B OR2X1_LOC_16/A 0.09fF
C38428 OR2X1_LOC_599/A OR2X1_LOC_16/A 0.04fF
C39693 AND2X1_LOC_841/B OR2X1_LOC_16/A 0.03fF
C40037 OR2X1_LOC_166/Y OR2X1_LOC_16/A 0.02fF
C41893 AND2X1_LOC_610/a_8_24# OR2X1_LOC_16/A 0.01fF
C43275 OR2X1_LOC_7/Y OR2X1_LOC_16/A 0.26fF
C46987 OR2X1_LOC_16/A OR2X1_LOC_312/a_8_216# 0.01fF
C47182 OR2X1_LOC_418/a_8_216# OR2X1_LOC_16/A 0.09fF
C47618 OR2X1_LOC_612/B OR2X1_LOC_16/A 0.03fF
C48077 OR2X1_LOC_273/Y OR2X1_LOC_16/A 0.06fF
C48167 OR2X1_LOC_75/Y OR2X1_LOC_16/A 0.04fF
C48274 OR2X1_LOC_16/A AND2X1_LOC_608/a_8_24# 0.01fF
C48503 AND2X1_LOC_78/a_8_24# OR2X1_LOC_16/A 0.10fF
C48799 OR2X1_LOC_16/A OR2X1_LOC_16/a_8_216# 0.18fF
C49364 OR2X1_LOC_52/Y OR2X1_LOC_16/A 0.02fF
C50044 OR2X1_LOC_604/A OR2X1_LOC_16/A 0.18fF
C50542 OR2X1_LOC_16/A OR2X1_LOC_265/Y 0.03fF
C51054 AND2X1_LOC_633/Y OR2X1_LOC_16/A 0.03fF
C51236 AND2X1_LOC_539/Y OR2X1_LOC_16/A 0.13fF
C51310 OR2X1_LOC_612/Y OR2X1_LOC_16/A 0.02fF
C52134 OR2X1_LOC_16/A AND2X1_LOC_434/Y 0.30fF
C52407 OR2X1_LOC_595/Y OR2X1_LOC_16/A 0.05fF
C53477 OR2X1_LOC_393/Y OR2X1_LOC_16/A 0.03fF
C53945 OR2X1_LOC_79/A OR2X1_LOC_16/A 0.16fF
C54194 OR2X1_LOC_135/Y OR2X1_LOC_16/A 2.07fF
C54553 OR2X1_LOC_16/A OR2X1_LOC_536/a_8_216# 0.01fF
C55148 OR2X1_LOC_313/a_8_216# OR2X1_LOC_16/A 0.05fF
C55489 OR2X1_LOC_829/A OR2X1_LOC_16/A 0.30fF
C55783 OR2X1_LOC_597/Y OR2X1_LOC_16/A 0.01fF
C56064 OR2X1_LOC_385/Y OR2X1_LOC_16/A 0.05fF
C56582 OR2X1_LOC_16/A VSS -3.88fF
C591 OR2X1_LOC_511/Y OR2X1_LOC_13/B 0.25fF
C604 OR2X1_LOC_248/a_8_216# OR2X1_LOC_13/B 0.01fF
C1407 OR2X1_LOC_13/B OR2X1_LOC_131/a_8_216# 0.02fF
C1429 AND2X1_LOC_391/Y OR2X1_LOC_13/B 0.03fF
C2381 OR2X1_LOC_74/A OR2X1_LOC_13/B 0.21fF
C2792 AND2X1_LOC_287/Y OR2X1_LOC_13/B 0.19fF
C3954 AND2X1_LOC_339/B OR2X1_LOC_13/B 0.03fF
C4793 OR2X1_LOC_597/a_8_216# OR2X1_LOC_13/B 0.02fF
C4818 AND2X1_LOC_99/A OR2X1_LOC_13/B 0.01fF
C5314 OR2X1_LOC_167/Y OR2X1_LOC_13/B 0.02fF
C6996 OR2X1_LOC_89/a_8_216# OR2X1_LOC_13/B 0.03fF
C7372 AND2X1_LOC_436/a_8_24# OR2X1_LOC_13/B 0.01fF
C7931 AND2X1_LOC_537/Y OR2X1_LOC_13/B 0.01fF
C8225 OR2X1_LOC_13/Y OR2X1_LOC_13/B 0.05fF
C8731 AND2X1_LOC_138/a_8_24# OR2X1_LOC_13/B 0.03fF
C10208 OR2X1_LOC_533/A OR2X1_LOC_13/B 0.02fF
C10367 OR2X1_LOC_597/a_36_216# OR2X1_LOC_13/B 0.03fF
C11179 VDD OR2X1_LOC_13/B 0.79fF
C11229 OR2X1_LOC_829/a_8_216# OR2X1_LOC_13/B 0.04fF
C11262 OR2X1_LOC_251/Y OR2X1_LOC_13/B 0.07fF
C11390 OR2X1_LOC_67/Y OR2X1_LOC_13/B 0.07fF
C11700 OR2X1_LOC_248/Y OR2X1_LOC_13/B 0.13fF
C12156 AND2X1_LOC_307/Y OR2X1_LOC_13/B 0.03fF
C13047 OR2X1_LOC_416/Y OR2X1_LOC_13/B 0.03fF
C13832 AND2X1_LOC_831/a_8_24# OR2X1_LOC_13/B 0.03fF
C14629 AND2X1_LOC_98/Y OR2X1_LOC_13/B 0.02fF
C15018 OR2X1_LOC_482/Y OR2X1_LOC_13/B 0.03fF
C16470 OR2X1_LOC_41/a_8_216# OR2X1_LOC_13/B 0.08fF
C16754 OR2X1_LOC_316/Y OR2X1_LOC_13/B 0.03fF
C16798 AND2X1_LOC_390/B OR2X1_LOC_13/B 0.09fF
C17206 AND2X1_LOC_840/B OR2X1_LOC_13/B 0.08fF
C17432 OR2X1_LOC_13/B OR2X1_LOC_320/a_8_216# 0.03fF
C17939 OR2X1_LOC_821/a_8_216# OR2X1_LOC_13/B 0.01fF
C18013 AND2X1_LOC_809/A OR2X1_LOC_13/B 0.10fF
C18961 OR2X1_LOC_311/Y OR2X1_LOC_13/B 0.10fF
C18968 AND2X1_LOC_538/Y OR2X1_LOC_13/B -0.01fF
C19272 AND2X1_LOC_330/a_8_24# OR2X1_LOC_13/B 0.01fF
C19436 AND2X1_LOC_831/Y OR2X1_LOC_13/B 0.06fF
C19763 AND2X1_LOC_436/B OR2X1_LOC_13/B -0.01fF
C20145 OR2X1_LOC_484/a_8_216# OR2X1_LOC_13/B 0.08fF
C21917 AND2X1_LOC_319/A OR2X1_LOC_13/B 0.02fF
C22065 AND2X1_LOC_721/A OR2X1_LOC_13/B 0.06fF
C22111 OR2X1_LOC_13/B OR2X1_LOC_331/Y 1.09fF
C22343 OR2X1_LOC_829/a_36_216# OR2X1_LOC_13/B 0.01fF
C22368 AND2X1_LOC_361/A OR2X1_LOC_13/B 0.07fF
C23090 AND2X1_LOC_284/a_8_24# OR2X1_LOC_13/B 0.03fF
C23981 OR2X1_LOC_166/a_8_216# OR2X1_LOC_13/B 0.01fF
C24506 AND2X1_LOC_539/a_8_24# OR2X1_LOC_13/B 0.01fF
C24813 OR2X1_LOC_331/A OR2X1_LOC_13/B 0.11fF
C26138 OR2X1_LOC_312/Y OR2X1_LOC_13/B 0.07fF
C26739 OR2X1_LOC_533/a_8_216# OR2X1_LOC_13/B 0.05fF
C26775 OR2X1_LOC_13/B OR2X1_LOC_142/a_8_216# 0.02fF
C26861 OR2X1_LOC_13/B OR2X1_LOC_595/A 0.24fF
C27369 AND2X1_LOC_342/Y OR2X1_LOC_13/B 0.04fF
C27404 OR2X1_LOC_279/a_8_216# OR2X1_LOC_13/B 0.03fF
C29979 AND2X1_LOC_538/a_8_24# OR2X1_LOC_13/B 0.01fF
C31109 AND2X1_LOC_535/Y OR2X1_LOC_13/B 0.01fF
C31185 OR2X1_LOC_246/Y OR2X1_LOC_13/B 0.20fF
C32448 AND2X1_LOC_729/B OR2X1_LOC_13/B 0.09fF
C32873 OR2X1_LOC_106/A OR2X1_LOC_13/B 0.03fF
C32960 AND2X1_LOC_227/Y OR2X1_LOC_13/B 0.03fF
C33001 OR2X1_LOC_813/Y OR2X1_LOC_13/B 0.35fF
C33266 OR2X1_LOC_250/a_8_216# OR2X1_LOC_13/B 0.02fF
C33672 AND2X1_LOC_535/a_8_24# OR2X1_LOC_13/B 0.02fF
C33704 AND2X1_LOC_843/Y OR2X1_LOC_13/B 0.02fF
C33751 OR2X1_LOC_320/Y OR2X1_LOC_13/B 0.58fF
C34504 AND2X1_LOC_841/B OR2X1_LOC_13/B 0.07fF
C34940 OR2X1_LOC_166/Y OR2X1_LOC_13/B 0.03fF
C36506 OR2X1_LOC_13/B OR2X1_LOC_525/a_8_216# 0.07fF
C37302 OR2X1_LOC_13/B AND2X1_LOC_247/a_8_24# 0.01fF
C37944 OR2X1_LOC_829/Y OR2X1_LOC_13/B 0.01fF
C38293 OR2X1_LOC_516/B OR2X1_LOC_13/B 0.01fF
C38355 OR2X1_LOC_279/Y OR2X1_LOC_13/B 0.02fF
C38740 AND2X1_LOC_456/B OR2X1_LOC_13/B 0.02fF
C39581 OR2X1_LOC_494/Y OR2X1_LOC_13/B 0.07fF
C39785 OR2X1_LOC_13/B OR2X1_LOC_311/a_8_216# 0.01fF
C39940 AND2X1_LOC_802/Y OR2X1_LOC_13/B 0.04fF
C40375 AND2X1_LOC_130/a_8_24# OR2X1_LOC_13/B 0.03fF
C42950 OR2X1_LOC_89/Y OR2X1_LOC_13/B 0.02fF
C43498 OR2X1_LOC_118/Y OR2X1_LOC_13/B 0.03fF
C43569 AND2X1_LOC_855/a_8_24# OR2X1_LOC_13/B 0.02fF
C44365 OR2X1_LOC_250/Y OR2X1_LOC_13/B 0.91fF
C44726 OR2X1_LOC_604/A OR2X1_LOC_13/B 0.17fF
C45155 OR2X1_LOC_533/Y OR2X1_LOC_13/B 0.09fF
C45590 AND2X1_LOC_809/a_8_24# OR2X1_LOC_13/B 0.03fF
C46003 AND2X1_LOC_539/Y OR2X1_LOC_13/B 0.12fF
C46970 AND2X1_LOC_434/Y OR2X1_LOC_13/B 2.24fF
C47929 AND2X1_LOC_342/a_8_24# OR2X1_LOC_13/B 0.24fF
C47942 AND2X1_LOC_355/a_8_24# OR2X1_LOC_13/B 0.01fF
C48590 OR2X1_LOC_13/B OR2X1_LOC_248/A 0.01fF
C49076 OR2X1_LOC_135/Y OR2X1_LOC_13/B 0.03fF
C49227 AND2X1_LOC_856/B OR2X1_LOC_13/B 0.01fF
C50394 OR2X1_LOC_829/A OR2X1_LOC_13/B 0.10fF
C51197 AND2X1_LOC_810/B OR2X1_LOC_13/B 0.01fF
C51629 AND2X1_LOC_130/a_36_24# OR2X1_LOC_13/B 0.01fF
C52573 AND2X1_LOC_784/A OR2X1_LOC_13/B 0.07fF
C53303 OR2X1_LOC_13/a_8_216# OR2X1_LOC_13/B 0.01fF
C53435 AND2X1_LOC_356/B OR2X1_LOC_13/B 0.01fF
C53775 OR2X1_LOC_485/Y OR2X1_LOC_13/B 0.35fF
C54206 AND2X1_LOC_593/Y OR2X1_LOC_13/B 0.02fF
C54655 OR2X1_LOC_680/A OR2X1_LOC_13/B 0.36fF
C55487 AND2X1_LOC_97/a_8_24# OR2X1_LOC_13/B 0.01fF
C56122 OR2X1_LOC_13/B OR2X1_LOC_331/a_8_216# 0.03fF
C56414 OR2X1_LOC_13/B VSS -5.53fF
C1044 OR2X1_LOC_74/A OR2X1_LOC_406/A 0.03fF
C1182 OR2X1_LOC_505/a_8_216# OR2X1_LOC_74/A 0.03fF
C2225 OR2X1_LOC_312/Y OR2X1_LOC_74/A 0.03fF
C2929 OR2X1_LOC_74/A OR2X1_LOC_595/A 0.15fF
C3372 OR2X1_LOC_528/Y OR2X1_LOC_74/A 10.35fF
C4949 OR2X1_LOC_821/Y OR2X1_LOC_74/A 0.01fF
C5464 OR2X1_LOC_438/Y OR2X1_LOC_74/A 0.03fF
C5511 OR2X1_LOC_74/A AND2X1_LOC_621/Y 0.12fF
C6035 OR2X1_LOC_504/Y OR2X1_LOC_74/A 0.19fF
C6059 OR2X1_LOC_437/Y OR2X1_LOC_74/A -0.02fF
C6659 OR2X1_LOC_505/a_36_216# OR2X1_LOC_74/A 0.02fF
C7264 OR2X1_LOC_246/Y OR2X1_LOC_74/A 0.03fF
C7665 AND2X1_LOC_168/Y OR2X1_LOC_74/A 0.39fF
C8596 OR2X1_LOC_109/Y OR2X1_LOC_74/A 0.11fF
C8623 OR2X1_LOC_262/a_8_216# OR2X1_LOC_74/A 0.06fF
C9084 OR2X1_LOC_679/A OR2X1_LOC_74/A 0.03fF
C9126 OR2X1_LOC_813/Y OR2X1_LOC_74/A 0.15fF
C9460 OR2X1_LOC_599/A OR2X1_LOC_74/A 0.03fF
C9724 OR2X1_LOC_177/a_8_216# OR2X1_LOC_74/A 0.02fF
C10200 OR2X1_LOC_531/Y OR2X1_LOC_74/A 0.01fF
C10376 OR2X1_LOC_74/A OR2X1_LOC_615/Y 0.03fF
C10588 OR2X1_LOC_813/a_8_216# OR2X1_LOC_74/A 0.01fF
C10918 AND2X1_LOC_543/Y OR2X1_LOC_74/A 0.04fF
C11569 OR2X1_LOC_74/A AND2X1_LOC_240/Y 0.03fF
C11992 OR2X1_LOC_74/A AND2X1_LOC_631/Y 0.08fF
C12352 OR2X1_LOC_74/Y OR2X1_LOC_74/A 0.02fF
C14007 OR2X1_LOC_96/Y OR2X1_LOC_74/A 0.02fF
C15709 AND2X1_LOC_147/a_36_24# OR2X1_LOC_74/A 0.01fF
C16496 AND2X1_LOC_325/a_8_24# OR2X1_LOC_74/A 0.03fF
C16597 OR2X1_LOC_74/A AND2X1_LOC_624/A 0.07fF
C18829 OR2X1_LOC_273/Y OR2X1_LOC_74/A 0.02fF
C19388 OR2X1_LOC_74/A OR2X1_LOC_142/Y 0.07fF
C19615 OR2X1_LOC_74/A OR2X1_LOC_118/Y 0.03fF
C20481 OR2X1_LOC_91/a_8_216# OR2X1_LOC_74/A 0.16fF
C20629 OR2X1_LOC_74/A OR2X1_LOC_152/A 0.03fF
C20763 OR2X1_LOC_177/Y OR2X1_LOC_74/A 0.02fF
C20789 OR2X1_LOC_604/A OR2X1_LOC_74/A 0.23fF
C21181 OR2X1_LOC_176/Y OR2X1_LOC_74/A 0.05fF
C21261 AND2X1_LOC_549/a_8_24# OR2X1_LOC_74/A 0.04fF
C21269 AND2X1_LOC_506/a_8_24# OR2X1_LOC_74/A 0.04fF
C21355 OR2X1_LOC_74/A OR2X1_LOC_265/Y 0.07fF
C22423 OR2X1_LOC_518/a_8_216# OR2X1_LOC_74/A 0.03fF
C22548 AND2X1_LOC_112/a_8_24# OR2X1_LOC_74/A 0.05fF
C22599 OR2X1_LOC_74/A OR2X1_LOC_746/a_8_216# 0.02fF
C23178 OR2X1_LOC_74/A OR2X1_LOC_595/Y 0.03fF
C24653 OR2X1_LOC_517/a_8_216# OR2X1_LOC_74/A 0.08fF
C25106 OR2X1_LOC_74/A AND2X1_LOC_520/Y 0.02fF
C25132 AND2X1_LOC_186/a_8_24# OR2X1_LOC_74/A 0.03fF
C26057 AND2X1_LOC_318/Y OR2X1_LOC_74/A 0.02fF
C26275 OR2X1_LOC_759/A OR2X1_LOC_74/A 0.03fF
C26745 AND2X1_LOC_508/A OR2X1_LOC_74/A 0.03fF
C27200 OR2X1_LOC_165/Y OR2X1_LOC_74/A 0.06fF
C27479 OR2X1_LOC_74/A OR2X1_LOC_368/Y 0.11fF
C27546 AND2X1_LOC_325/a_36_24# OR2X1_LOC_74/A 0.01fF
C27987 AND2X1_LOC_715/A OR2X1_LOC_74/A 0.14fF
C28371 OR2X1_LOC_74/A OR2X1_LOC_323/Y 0.02fF
C28492 AND2X1_LOC_729/Y OR2X1_LOC_74/A 0.03fF
C28517 AND2X1_LOC_784/A OR2X1_LOC_74/A 0.24fF
C29305 OR2X1_LOC_165/a_8_216# OR2X1_LOC_74/A 0.02fF
C30597 OR2X1_LOC_680/A OR2X1_LOC_74/A 0.10fF
C30967 OR2X1_LOC_757/A OR2X1_LOC_74/A 0.03fF
C31836 OR2X1_LOC_252/Y OR2X1_LOC_74/A 0.03fF
C32188 AND2X1_LOC_549/a_36_24# OR2X1_LOC_74/A 0.01fF
C32192 OR2X1_LOC_677/a_8_216# OR2X1_LOC_74/A 0.03fF
C32193 AND2X1_LOC_506/a_36_24# OR2X1_LOC_74/A 0.01fF
C33529 OR2X1_LOC_74/A OR2X1_LOC_746/a_36_216# 0.03fF
C34402 AND2X1_LOC_673/a_8_24# OR2X1_LOC_74/A 0.17fF
C35229 OR2X1_LOC_235/a_8_216# OR2X1_LOC_74/A 0.01fF
C37052 OR2X1_LOC_74/A OR2X1_LOC_72/Y 0.07fF
C37384 OR2X1_LOC_680/Y OR2X1_LOC_74/A 0.03fF
C37697 OR2X1_LOC_677/a_36_216# OR2X1_LOC_74/A 0.02fF
C37747 OR2X1_LOC_74/A OR2X1_LOC_595/a_8_216# 0.05fF
C38127 AND2X1_LOC_168/a_8_24# OR2X1_LOC_74/A 0.04fF
C39987 OR2X1_LOC_437/a_8_216# OR2X1_LOC_74/A 0.02fF
C40189 OR2X1_LOC_74/A OR2X1_LOC_627/Y 0.14fF
C41444 OR2X1_LOC_406/Y OR2X1_LOC_74/A 0.03fF
C41846 OR2X1_LOC_516/Y OR2X1_LOC_74/A 0.53fF
C42391 OR2X1_LOC_368/a_8_216# OR2X1_LOC_74/A 0.24fF
C42810 OR2X1_LOC_528/a_8_216# OR2X1_LOC_74/A 0.03fF
C43262 VDD OR2X1_LOC_74/A 1.53fF
C43306 OR2X1_LOC_677/Y OR2X1_LOC_74/A 0.03fF
C43353 OR2X1_LOC_315/Y OR2X1_LOC_74/A 0.02fF
C43480 OR2X1_LOC_74/A OR2X1_LOC_67/Y 0.07fF
C44204 OR2X1_LOC_74/A OR2X1_LOC_531/a_8_216# 0.01fF
C48314 OR2X1_LOC_111/Y OR2X1_LOC_74/A 0.09fF
C48328 OR2X1_LOC_146/Y OR2X1_LOC_74/A 0.03fF
C49021 OR2X1_LOC_316/Y OR2X1_LOC_74/A 0.03fF
C49431 AND2X1_LOC_168/a_36_24# OR2X1_LOC_74/A 0.01fF
C49491 AND2X1_LOC_840/B OR2X1_LOC_74/A 0.10fF
C49496 OR2X1_LOC_74/A OR2X1_LOC_74/a_8_216# 0.04fF
C51138 OR2X1_LOC_91/Y OR2X1_LOC_74/A 0.26fF
C51195 OR2X1_LOC_527/Y OR2X1_LOC_74/A 0.07fF
C51645 AND2X1_LOC_831/Y OR2X1_LOC_74/A 0.01fF
C51930 OR2X1_LOC_441/Y OR2X1_LOC_74/A 14.70fF
C51979 AND2X1_LOC_139/B OR2X1_LOC_74/A 0.07fF
C52001 OR2X1_LOC_235/Y OR2X1_LOC_74/A 0.01fF
C52603 OR2X1_LOC_74/A AND2X1_LOC_789/Y 0.02fF
C52852 OR2X1_LOC_517/Y OR2X1_LOC_74/A 0.04fF
C53975 OR2X1_LOC_528/a_36_216# OR2X1_LOC_74/A 0.02fF
C54018 OR2X1_LOC_235/B OR2X1_LOC_74/A 0.02fF
C54190 AND2X1_LOC_721/A OR2X1_LOC_74/A 0.60fF
C55208 AND2X1_LOC_787/A OR2X1_LOC_74/A 0.03fF
C55334 AND2X1_LOC_147/a_8_24# OR2X1_LOC_74/A 0.05fF
C55371 OR2X1_LOC_74/A OR2X1_LOC_406/a_8_216# 0.02fF
C55638 OR2X1_LOC_821/a_36_216# OR2X1_LOC_74/A 0.03fF
C56197 AND2X1_LOC_543/a_8_24# OR2X1_LOC_74/A 0.02fF
C57015 OR2X1_LOC_74/A VSS -6.14fF
C16045 VDD OR2X1_LOC_246/Y 0.03fF
C16584 OR2X1_LOC_246/Y OR2X1_LOC_248/Y 0.09fF
C26883 OR2X1_LOC_246/Y AND2X1_LOC_721/A 0.02fF
C33811 OR2X1_LOC_821/Y OR2X1_LOC_246/Y 0.30fF
C38909 OR2X1_LOC_246/Y OR2X1_LOC_822/a_8_216# 0.40fF
C57796 OR2X1_LOC_246/Y VSS -0.18fF
C348 OR2X1_LOC_235/B OR2X1_LOC_720/A 0.01fF
C784 OR2X1_LOC_235/B OR2X1_LOC_267/A 0.03fF
C1367 OR2X1_LOC_235/B AND2X1_LOC_813/a_8_24# 0.03fF
C1946 OR2X1_LOC_235/B OR2X1_LOC_673/a_8_216# 0.02fF
C2176 OR2X1_LOC_235/B AND2X1_LOC_107/a_8_24# 0.01fF
C5315 OR2X1_LOC_114/a_8_216# OR2X1_LOC_235/B 0.01fF
C6587 VDD OR2X1_LOC_235/B 2.18fF
C6852 OR2X1_LOC_235/B OR2X1_LOC_845/A 0.06fF
C7391 OR2X1_LOC_235/B OR2X1_LOC_523/A 0.01fF
C9769 OR2X1_LOC_235/B OR2X1_LOC_235/a_36_216# 0.03fF
C12292 OR2X1_LOC_114/Y OR2X1_LOC_235/B 0.16fF
C13176 OR2X1_LOC_235/B OR2X1_LOC_643/A 0.03fF
C15234 OR2X1_LOC_235/B OR2X1_LOC_235/Y 0.01fF
C15506 AND2X1_LOC_521/a_8_24# OR2X1_LOC_235/B 0.02fF
C18088 OR2X1_LOC_235/B OR2X1_LOC_362/A 0.02fF
C18450 OR2X1_LOC_235/B OR2X1_LOC_771/B 0.07fF
C19620 OR2X1_LOC_235/B OR2X1_LOC_720/B 0.79fF
C20774 AND2X1_LOC_394/a_8_24# OR2X1_LOC_235/B 0.03fF
C21081 OR2X1_LOC_523/B OR2X1_LOC_235/B 0.01fF
C27393 AND2X1_LOC_522/a_8_24# OR2X1_LOC_235/B 0.01fF
C28321 OR2X1_LOC_768/A OR2X1_LOC_235/B 0.01fF
C30908 OR2X1_LOC_235/B AND2X1_LOC_132/a_8_24# 0.01fF
C30969 OR2X1_LOC_235/B AND2X1_LOC_240/Y 0.02fF
C31757 OR2X1_LOC_400/A OR2X1_LOC_235/B 0.02fF
C36372 OR2X1_LOC_235/B OR2X1_LOC_137/B 0.01fF
C39790 OR2X1_LOC_235/B OR2X1_LOC_668/Y 0.01fF
C40328 OR2X1_LOC_235/B OR2X1_LOC_84/A 0.02fF
C42422 OR2X1_LOC_235/B OR2X1_LOC_810/A 0.05fF
C43710 OR2X1_LOC_235/B AND2X1_LOC_399/a_8_24# 0.04fF
C45413 OR2X1_LOC_235/B AND2X1_LOC_669/a_8_24# 0.01fF
C45735 OR2X1_LOC_114/B OR2X1_LOC_235/B 0.01fF
C45891 OR2X1_LOC_235/B AND2X1_LOC_79/Y 0.07fF
C52306 OR2X1_LOC_235/B OR2X1_LOC_673/Y -0.00fF
C54816 OR2X1_LOC_235/B OR2X1_LOC_235/a_8_216# 0.02fF
C54829 OR2X1_LOC_235/B OR2X1_LOC_403/B 0.01fF
C57778 OR2X1_LOC_235/B VSS 0.22fF
C189 OR2X1_LOC_604/A OR2X1_LOC_96/Y 0.07fF
C353 OR2X1_LOC_604/A OR2X1_LOC_617/a_8_216# 0.15fF
C785 OR2X1_LOC_604/A OR2X1_LOC_279/Y 0.10fF
C1112 OR2X1_LOC_604/A AND2X1_LOC_456/B 0.06fF
C2177 OR2X1_LOC_604/A OR2X1_LOC_96/a_8_216# 0.47fF
C2533 OR2X1_LOC_604/A AND2X1_LOC_154/Y 0.01fF
C2903 OR2X1_LOC_604/A AND2X1_LOC_624/A 0.10fF
C3348 OR2X1_LOC_604/A OR2X1_LOC_669/a_8_216# 0.10fF
C3938 OR2X1_LOC_604/A OR2X1_LOC_746/Y 0.16fF
C4173 OR2X1_LOC_604/A OR2X1_LOC_418/a_8_216# 0.01fF
C4446 OR2X1_LOC_604/A AND2X1_LOC_160/Y 0.01fF
C4608 OR2X1_LOC_604/A OR2X1_LOC_295/a_8_216# 0.11fF
C5019 OR2X1_LOC_604/A OR2X1_LOC_253/a_8_216# 0.03fF
C5213 OR2X1_LOC_604/A OR2X1_LOC_744/a_8_216# 0.01fF
C5371 OR2X1_LOC_604/A OR2X1_LOC_601/Y 0.01fF
C5414 OR2X1_LOC_604/A OR2X1_LOC_754/A 0.40fF
C5844 OR2X1_LOC_604/A OR2X1_LOC_238/Y 0.03fF
C6977 OR2X1_LOC_177/Y OR2X1_LOC_604/A 0.03fF
C6998 OR2X1_LOC_604/A OR2X1_LOC_745/a_8_216# 0.12fF
C7086 OR2X1_LOC_604/A OR2X1_LOC_252/a_8_216# 0.07fF
C7425 OR2X1_LOC_533/Y OR2X1_LOC_604/A 0.03fF
C7531 OR2X1_LOC_604/A AND2X1_LOC_447/a_8_24# 0.08fF
C7675 OR2X1_LOC_604/A OR2X1_LOC_96/a_36_216# 0.01fF
C7798 OR2X1_LOC_604/A OR2X1_LOC_183/a_8_216# 0.30fF
C8039 OR2X1_LOC_604/A AND2X1_LOC_155/Y 0.01fF
C8115 OR2X1_LOC_604/A AND2X1_LOC_450/Y -0.00fF
C8797 OR2X1_LOC_604/A OR2X1_LOC_746/a_8_216# 0.01fF
C9779 OR2X1_LOC_604/A AND2X1_LOC_260/a_8_24# 0.05fF
C11364 OR2X1_LOC_604/A AND2X1_LOC_848/Y 0.20fF
C11441 OR2X1_LOC_604/A OR2X1_LOC_617/Y 0.06fF
C11732 AND2X1_LOC_756/a_8_24# OR2X1_LOC_604/A 0.11fF
C11753 OR2X1_LOC_604/A AND2X1_LOC_160/a_8_24# 0.01fF
C12214 OR2X1_LOC_313/a_8_216# OR2X1_LOC_604/A 0.01fF
C12293 OR2X1_LOC_604/A OR2X1_LOC_258/Y 0.02fF
C12579 OR2X1_LOC_604/A OR2X1_LOC_697/a_8_216# 0.14fF
C12590 OR2X1_LOC_604/A OR2X1_LOC_698/Y 0.01fF
C14766 AND2X1_LOC_729/Y OR2X1_LOC_604/A 0.07fF
C14790 AND2X1_LOC_784/A OR2X1_LOC_604/A 0.10fF
C15474 OR2X1_LOC_604/A OR2X1_LOC_281/Y 0.09fF
C15489 OR2X1_LOC_604/A OR2X1_LOC_253/Y 0.02fF
C15637 OR2X1_LOC_604/A OR2X1_LOC_280/Y 0.10fF
C15671 OR2X1_LOC_604/A OR2X1_LOC_295/a_36_216# 0.01fF
C15917 OR2X1_LOC_604/A OR2X1_LOC_485/Y 0.09fF
C16311 OR2X1_LOC_604/A OR2X1_LOC_744/Y 0.21fF
C16420 OR2X1_LOC_604/A AND2X1_LOC_593/Y 0.03fF
C16895 OR2X1_LOC_604/A OR2X1_LOC_680/A 0.07fF
C17335 OR2X1_LOC_604/A OR2X1_LOC_626/a_8_216# 0.05fF
C17624 OR2X1_LOC_604/A AND2X1_LOC_436/Y 0.08fF
C17710 OR2X1_LOC_604/A OR2X1_LOC_603/a_8_216# 0.01fF
C18158 OR2X1_LOC_604/A OR2X1_LOC_252/Y 0.01fF
C18164 OR2X1_LOC_604/A OR2X1_LOC_313/Y 0.02fF
C18875 OR2X1_LOC_604/A OR2X1_LOC_183/Y 0.03fF
C19024 OR2X1_LOC_604/A OR2X1_LOC_511/Y 0.17fF
C19170 OR2X1_LOC_604/A AND2X1_LOC_451/Y 0.81fF
C19371 OR2X1_LOC_604/A OR2X1_LOC_600/a_8_216# 0.01fF
C19450 OR2X1_LOC_604/A OR2X1_LOC_237/Y 0.03fF
C19495 OR2X1_LOC_604/A OR2X1_LOC_487/a_8_216# 0.30fF
C19936 OR2X1_LOC_604/A OR2X1_LOC_669/Y 1.05fF
C20820 OR2X1_LOC_604/A OR2X1_LOC_261/A -0.01fF
C21065 OR2X1_LOC_604/A AND2X1_LOC_254/a_8_24# -0.04fF
C21077 OR2X1_LOC_604/A OR2X1_LOC_626/Y 0.03fF
C21925 OR2X1_LOC_604/A AND2X1_LOC_704/a_8_24# 0.02fF
C22385 OR2X1_LOC_604/A OR2X1_LOC_816/a_8_216# 0.03fF
C23351 OR2X1_LOC_604/A OR2X1_LOC_627/a_8_216# 0.06fF
C23683 OR2X1_LOC_604/A OR2X1_LOC_697/Y 0.08fF
C24444 OR2X1_LOC_604/A OR2X1_LOC_603/Y 0.02fF
C24507 OR2X1_LOC_604/A AND2X1_LOC_168/a_8_24# 0.13fF
C24590 OR2X1_LOC_604/A OR2X1_LOC_665/Y 0.07fF
C25002 OR2X1_LOC_604/A OR2X1_LOC_420/a_8_216# 0.01fF
C25387 OR2X1_LOC_604/A AND2X1_LOC_458/Y 0.26fF
C26245 OR2X1_LOC_604/A OR2X1_LOC_418/Y 0.38fF
C26486 OR2X1_LOC_604/A OR2X1_LOC_743/Y -0.01fF
C26537 OR2X1_LOC_604/A AND2X1_LOC_285/a_8_24# 0.07fF
C26555 OR2X1_LOC_604/A OR2X1_LOC_627/Y 0.03fF
C26740 OR2X1_LOC_604/A OR2X1_LOC_295/Y 0.06fF
C26974 OR2X1_LOC_604/A OR2X1_LOC_526/Y 0.01fF
C27383 OR2X1_LOC_604/A AND2X1_LOC_714/B 0.12fF
C28554 OR2X1_LOC_604/A AND2X1_LOC_793/B 0.07fF
C28557 OR2X1_LOC_604/A OR2X1_LOC_533/A 0.03fF
C29177 OR2X1_LOC_604/A OR2X1_LOC_314/Y 0.38fF
C29517 OR2X1_LOC_604/A VDD 6.36fF
C29610 OR2X1_LOC_604/A AND2X1_LOC_447/a_36_24# 0.02fF
C29638 OR2X1_LOC_604/A OR2X1_LOC_251/Y 0.03fF
C29799 OR2X1_LOC_604/A OR2X1_LOC_163/Y 0.03fF
C29986 OR2X1_LOC_314/a_8_216# OR2X1_LOC_604/A 0.01fF
C30373 OR2X1_LOC_604/A OR2X1_LOC_600/Y 0.01fF
C30461 OR2X1_LOC_604/A OR2X1_LOC_591/A 0.03fF
C31681 OR2X1_LOC_604/A OR2X1_LOC_281/a_8_216# 0.35fF
C32056 OR2X1_LOC_604/A OR2X1_LOC_485/a_8_216# 0.01fF
C32691 OR2X1_LOC_604/A OR2X1_LOC_428/Y 0.02fF
C32933 OR2X1_LOC_604/A OR2X1_LOC_594/Y 0.14fF
C34532 OR2X1_LOC_591/Y OR2X1_LOC_604/A 0.02fF
C34657 OR2X1_LOC_604/A AND2X1_LOC_317/a_8_24# 0.01fF
C35003 OR2X1_LOC_604/A OR2X1_LOC_765/a_8_216# 0.01fF
C35360 OR2X1_LOC_604/A OR2X1_LOC_604/Y 0.21fF
C35564 OR2X1_LOC_604/A OR2X1_LOC_282/a_8_216# 0.07fF
C35684 OR2X1_LOC_604/A OR2X1_LOC_257/Y 0.06fF
C35805 OR2X1_LOC_604/A AND2X1_LOC_464/A 0.03fF
C35969 OR2X1_LOC_604/A OR2X1_LOC_420/Y 0.08fF
C36467 OR2X1_LOC_604/A OR2X1_LOC_751/A 0.17fF
C37093 OR2X1_LOC_604/A AND2X1_LOC_285/Y 0.03fF
C37182 OR2X1_LOC_91/Y OR2X1_LOC_604/A 0.10fF
C37206 OR2X1_LOC_604/A AND2X1_LOC_446/a_8_24# 0.02fF
C37276 OR2X1_LOC_604/A OR2X1_LOC_601/a_8_216# 0.01fF
C37465 OR2X1_LOC_604/A AND2X1_LOC_780/a_8_24# 0.01fF
C37960 OR2X1_LOC_604/A OR2X1_LOC_441/Y 0.03fF
C39344 OR2X1_LOC_604/A OR2X1_LOC_497/Y 0.10fF
C40136 OR2X1_LOC_604/A AND2X1_LOC_319/A 0.01fF
C40213 OR2X1_LOC_604/A AND2X1_LOC_708/a_8_24# 0.01fF
C40265 OR2X1_LOC_604/A OR2X1_LOC_604/a_8_216# 0.14fF
C40349 OR2X1_LOC_604/A OR2X1_LOC_331/Y 0.07fF
C41305 AND2X1_LOC_787/A OR2X1_LOC_604/A 0.01fF
C41428 AND2X1_LOC_532/a_8_24# OR2X1_LOC_604/A 0.16fF
C41881 OR2X1_LOC_604/A OR2X1_LOC_257/a_8_216# 0.04fF
C42786 OR2X1_LOC_604/A OR2X1_LOC_669/A 0.29fF
C42813 OR2X1_LOC_604/A AND2X1_LOC_454/A 0.25fF
C43051 OR2X1_LOC_604/A AND2X1_LOC_783/B 0.01fF
C43101 OR2X1_LOC_604/A AND2X1_LOC_285/a_36_24# 0.01fF
C43581 OR2X1_LOC_604/A OR2X1_LOC_292/Y 0.04fF
C44534 OR2X1_LOC_604/A OR2X1_LOC_312/Y 0.01fF
C45360 OR2X1_LOC_604/A AND2X1_LOC_154/a_8_24# 0.01fF
C45696 OR2X1_LOC_528/Y OR2X1_LOC_604/A 0.07fF
C45888 OR2X1_LOC_604/A AND2X1_LOC_712/B 0.03fF
C46146 OR2X1_LOC_604/A OR2X1_LOC_765/Y 0.01fF
C46439 OR2X1_LOC_604/A AND2X1_LOC_451/a_8_24# 0.01fF
C46543 OR2X1_LOC_604/A AND2X1_LOC_590/a_8_24# 0.01fF
C46582 OR2X1_LOC_167/a_8_216# OR2X1_LOC_604/A 0.12fF
C46786 OR2X1_LOC_604/A OR2X1_LOC_282/Y 0.05fF
C47011 OR2X1_LOC_604/A AND2X1_LOC_287/B 0.09fF
C47166 OR2X1_LOC_604/A OR2X1_LOC_427/a_8_216# 0.01fF
C47281 OR2X1_LOC_604/A AND2X1_LOC_727/A 0.03fF
C47609 OR2X1_LOC_604/A OR2X1_LOC_257/a_36_216# 0.01fF
C48026 OR2X1_LOC_604/A OR2X1_LOC_427/Y 0.02fF
C48044 OR2X1_LOC_604/A AND2X1_LOC_621/Y 0.09fF
C50069 OR2X1_LOC_604/A OR2X1_LOC_108/Y 0.10fF
C50916 OR2X1_LOC_604/A AND2X1_LOC_447/Y 0.10fF
C50974 OR2X1_LOC_604/A OR2X1_LOC_109/Y 0.10fF
C51531 OR2X1_LOC_604/A AND2X1_LOC_227/Y 0.28fF
C51856 OR2X1_LOC_599/A OR2X1_LOC_604/A 0.03fF
C52168 OR2X1_LOC_604/A OR2X1_LOC_698/a_8_216# 0.03fF
C52975 AND2X1_LOC_707/Y OR2X1_LOC_604/A 0.01fF
C53500 OR2X1_LOC_604/A OR2X1_LOC_495/Y 0.25fF
C53510 OR2X1_LOC_604/A AND2X1_LOC_450/a_8_24# 0.01fF
C56047 OR2X1_LOC_604/A AND2X1_LOC_161/a_8_24# 0.15fF
C57895 OR2X1_LOC_604/A VSS 1.27fF
C7663 OR2X1_LOC_599/A OR2X1_LOC_511/Y 0.02fF
C10870 OR2X1_LOC_511/Y OR2X1_LOC_525/a_8_216# 0.03fF
C16348 OR2X1_LOC_511/Y OR2X1_LOC_525/a_36_216# 0.02fF
C26755 AND2X1_LOC_729/Y OR2X1_LOC_511/Y 0.03fF
C27915 OR2X1_LOC_485/Y OR2X1_LOC_511/Y 0.03fF
C28862 OR2X1_LOC_680/A OR2X1_LOC_511/Y 0.01fF
C33921 AND2X1_LOC_779/a_8_24# OR2X1_LOC_511/Y 0.23fF
C35561 OR2X1_LOC_697/Y OR2X1_LOC_511/Y 0.06fF
C38914 OR2X1_LOC_526/Y OR2X1_LOC_511/Y 0.03fF
C41472 VDD OR2X1_LOC_511/Y 0.17fF
C41520 OR2X1_LOC_677/Y OR2X1_LOC_511/Y 0.01fF
C42014 OR2X1_LOC_511/Y AND2X1_LOC_834/a_8_24# 0.01fF
C44137 OR2X1_LOC_485/a_8_216# OR2X1_LOC_511/Y 0.02fF
C47742 OR2X1_LOC_511/Y AND2X1_LOC_840/B 0.01fF
C51478 OR2X1_LOC_525/Y OR2X1_LOC_511/Y 0.22fF
C55290 OR2X1_LOC_485/a_36_216# OR2X1_LOC_511/Y 0.02fF
C57023 OR2X1_LOC_511/Y VSS 0.17fF
C8109 OR2X1_LOC_406/Y OR2X1_LOC_406/A 0.01fF
C8191 OR2X1_LOC_496/a_8_216# OR2X1_LOC_406/A 0.02fF
C8542 OR2X1_LOC_516/Y OR2X1_LOC_406/A 0.07fF
C9899 VDD OR2X1_LOC_406/A 0.21fF
C15848 AND2X1_LOC_840/B OR2X1_LOC_406/A 0.45fF
C17546 OR2X1_LOC_91/Y OR2X1_LOC_406/A 0.08fF
C17582 OR2X1_LOC_527/Y OR2X1_LOC_406/A 0.01fF
C21875 OR2X1_LOC_406/a_8_216# OR2X1_LOC_406/A 0.01fF
C28178 AND2X1_LOC_621/Y OR2X1_LOC_406/A 0.07fF
C30992 AND2X1_LOC_778/a_36_24# OR2X1_LOC_406/A 0.01fF
C31123 OR2X1_LOC_109/Y OR2X1_LOC_406/A 0.01fF
C34014 AND2X1_LOC_776/a_8_24# OR2X1_LOC_406/A 0.01fF
C39085 OR2X1_LOC_406/A AND2X1_LOC_778/Y 0.23fF
C39165 AND2X1_LOC_624/A OR2X1_LOC_406/A 0.06fF
C41955 OR2X1_LOC_406/A OR2X1_LOC_142/Y 0.07fF
C45648 OR2X1_LOC_496/Y OR2X1_LOC_406/A 0.01fF
C51253 AND2X1_LOC_778/a_8_24# OR2X1_LOC_406/A 0.01fF
C53342 OR2X1_LOC_680/A OR2X1_LOC_406/A 0.07fF
C56466 OR2X1_LOC_406/A VSS -0.19fF
C6886 OR2X1_LOC_48/Y AND2X1_LOC_196/a_8_24# 0.01fF
C26709 VDD OR2X1_LOC_48/Y 0.05fF
C36975 OR2X1_LOC_48/Y OR2X1_LOC_7/a_8_216# 0.39fF
C54165 OR2X1_LOC_48/Y AND2X1_LOC_196/Y 0.01fF
C57640 OR2X1_LOC_48/Y VSS 0.20fF
C5978 OR2X1_LOC_763/Y OR2X1_LOC_764/Y 0.21fF
C10098 OR2X1_LOC_763/Y OR2X1_LOC_764/a_8_216# 0.39fF
C26263 OR2X1_LOC_763/Y VDD 0.08fF
C57878 OR2X1_LOC_763/Y VSS 0.11fF
C1157 OR2X1_LOC_599/A OR2X1_LOC_829/A 0.02fF
C1430 OR2X1_LOC_599/A OR2X1_LOC_597/Y 0.01fF
C3439 AND2X1_LOC_729/Y OR2X1_LOC_599/A 0.11fF
C4952 OR2X1_LOC_599/A OR2X1_LOC_536/Y 0.01fF
C5049 OR2X1_LOC_599/A AND2X1_LOC_593/Y 0.04fF
C6335 OR2X1_LOC_145/a_8_216# OR2X1_LOC_599/A 0.01fF
C6446 OR2X1_LOC_599/A OR2X1_LOC_145/Y 0.01fF
C6632 OR2X1_LOC_599/A AND2X1_LOC_828/a_36_24# 0.01fF
C9148 OR2X1_LOC_599/A OR2X1_LOC_423/Y 0.01fF
C10561 OR2X1_LOC_599/A AND2X1_LOC_537/a_8_24# 0.01fF
C10636 AND2X1_LOC_779/a_8_24# OR2X1_LOC_599/A 0.03fF
C11852 OR2X1_LOC_599/A OR2X1_LOC_597/a_8_216# 0.01fF
C12302 OR2X1_LOC_599/A OR2X1_LOC_697/Y 0.01fF
C15694 OR2X1_LOC_599/A OR2X1_LOC_433/Y 0.01fF
C16764 OR2X1_LOC_599/A OR2X1_LOC_589/a_8_216# 0.01fF
C18196 OR2X1_LOC_599/A VDD 0.02fF
C19169 OR2X1_LOC_599/A OR2X1_LOC_591/A 0.05fF
C20210 OR2X1_LOC_599/A AND2X1_LOC_592/a_8_24# 0.01fF
C21304 OR2X1_LOC_599/A AND2X1_LOC_435/a_8_24# 0.01fF
C23309 OR2X1_LOC_591/Y OR2X1_LOC_599/A 0.06fF
C26716 OR2X1_LOC_599/A OR2X1_LOC_441/Y 0.03fF
C26768 OR2X1_LOC_599/A AND2X1_LOC_436/B 0.02fF
C27717 OR2X1_LOC_599/A OR2X1_LOC_409/B 0.33fF
C27854 OR2X1_LOC_146/a_8_216# OR2X1_LOC_599/A 0.01fF
C28040 OR2X1_LOC_599/A AND2X1_LOC_676/a_8_24# 0.04fF
C28882 OR2X1_LOC_599/A AND2X1_LOC_319/A 0.21fF
C31658 OR2X1_LOC_599/A AND2X1_LOC_783/B 0.01fF
C34227 AND2X1_LOC_592/Y OR2X1_LOC_599/A 0.01fF
C35656 OR2X1_LOC_599/A OR2X1_LOC_591/a_8_216# 0.03fF
C36024 OR2X1_LOC_599/A AND2X1_LOC_832/a_8_24# 0.02fF
C36446 OR2X1_LOC_599/A AND2X1_LOC_621/Y 0.02fF
C38682 OR2X1_LOC_599/A AND2X1_LOC_687/Y 0.02fF
C39032 OR2X1_LOC_599/A AND2X1_LOC_676/a_36_24# 0.01fF
C39359 OR2X1_LOC_599/A AND2X1_LOC_447/Y 0.05fF
C39756 AND2X1_LOC_593/a_8_24# OR2X1_LOC_599/A 0.04fF
C40699 OR2X1_LOC_599/A OR2X1_LOC_424/a_8_216# 0.01fF
C41566 OR2X1_LOC_599/A AND2X1_LOC_841/B 0.18fF
C42510 OR2X1_LOC_599/A AND2X1_LOC_147/Y 0.14fF
C46227 OR2X1_LOC_599/A AND2X1_LOC_828/a_8_24# 0.03fF
C47737 OR2X1_LOC_599/A AND2X1_LOC_624/A 0.03fF
C48541 OR2X1_LOC_599/A OR2X1_LOC_524/Y 0.34fF
C49147 OR2X1_LOC_599/A AND2X1_LOC_779/Y 0.04fF
C57912 OR2X1_LOC_599/A VSS 0.86fF
C57689 OR2X1_LOC_692/Y VSS 0.13fF
C4511 OR2X1_LOC_519/Y VDD 0.09fF
C12865 OR2X1_LOC_519/Y AND2X1_LOC_831/Y 0.01fF
C16811 OR2X1_LOC_519/Y AND2X1_LOC_520/a_8_24# 0.01fF
C39319 OR2X1_LOC_519/Y AND2X1_LOC_326/B 0.02fF
C42417 OR2X1_LOC_519/Y AND2X1_LOC_520/Y 0.12fF
C45923 AND2X1_LOC_784/A OR2X1_LOC_519/Y 0.01fF
C58001 OR2X1_LOC_519/Y VSS 0.16fF
C48062 VDD AND2X1_LOC_458/Y 0.24fF
C49421 AND2X1_LOC_458/Y AND2X1_LOC_464/a_8_24# 0.19fF
C54293 AND2X1_LOC_458/Y AND2X1_LOC_464/A 0.10fF
C56852 AND2X1_LOC_458/Y VSS 0.07fF
C1148 OR2X1_LOC_409/B OR2X1_LOC_385/a_8_216# 0.01fF
C12838 AND2X1_LOC_638/Y OR2X1_LOC_409/B 0.31fF
C18701 OR2X1_LOC_409/B AND2X1_LOC_769/Y 0.01fF
C33513 OR2X1_LOC_409/B AND2X1_LOC_828/a_8_24# 0.10fF
C40734 OR2X1_LOC_409/B AND2X1_LOC_637/a_8_24# 0.01fF
C41261 OR2X1_LOC_764/Y OR2X1_LOC_409/B 0.01fF
C45188 OR2X1_LOC_385/Y OR2X1_LOC_409/B 0.01fF
C46965 AND2X1_LOC_769/a_8_24# OR2X1_LOC_409/B 0.01fF
C51985 OR2X1_LOC_409/B AND2X1_LOC_637/a_36_24# -0.00fF
C54531 OR2X1_LOC_409/B OR2X1_LOC_586/a_8_216# 0.47fF
C55440 OR2X1_LOC_409/B AND2X1_LOC_637/Y 0.02fF
C56873 OR2X1_LOC_409/B VSS 0.69fF
C958 OR2X1_LOC_743/Y AND2X1_LOC_780/a_8_24# 0.23fF
C43080 OR2X1_LOC_697/Y OR2X1_LOC_743/Y -0.00fF
C49144 VDD OR2X1_LOC_743/Y 0.12fF
C56442 OR2X1_LOC_743/Y VSS -0.07fF
C2114 OR2X1_LOC_433/Y AND2X1_LOC_436/B 0.01fF
C3191 OR2X1_LOC_433/Y OR2X1_LOC_589/a_36_216# -0.00fF
C40441 OR2X1_LOC_433/Y OR2X1_LOC_423/Y 0.01fF
C41540 OR2X1_LOC_432/Y OR2X1_LOC_433/Y 0.33fF
C44451 AND2X1_LOC_706/Y OR2X1_LOC_433/Y 0.06fF
C46107 OR2X1_LOC_433/Y OR2X1_LOC_589/Y 0.10fF
C47586 AND2X1_LOC_714/B OR2X1_LOC_433/Y 0.13fF
C48351 OR2X1_LOC_433/Y OR2X1_LOC_589/a_8_216# 0.01fF
C49732 VDD OR2X1_LOC_433/Y 0.20fF
C52764 OR2X1_LOC_433/Y AND2X1_LOC_435/a_8_24# 0.24fF
C56624 OR2X1_LOC_433/Y VSS 0.17fF
C7419 OR2X1_LOC_273/Y OR2X1_LOC_595/Y 0.01fF
C22208 OR2X1_LOC_273/Y OR2X1_LOC_595/a_8_216# 0.02fF
C27554 VDD OR2X1_LOC_273/Y 0.23fF
C29411 OR2X1_LOC_273/Y OR2X1_LOC_416/Y 0.04fF
C30198 OR2X1_LOC_273/Y AND2X1_LOC_831/a_8_24# 0.23fF
C33134 OR2X1_LOC_273/Y OR2X1_LOC_316/Y 0.03fF
C33137 OR2X1_LOC_273/Y OR2X1_LOC_595/a_36_216# 0.03fF
C57366 OR2X1_LOC_273/Y VSS 0.26fF
C3509 AND2X1_LOC_154/Y AND2X1_LOC_155/Y 0.22fF
C6211 AND2X1_LOC_155/Y OR2X1_LOC_744/a_8_216# 0.49fF
C20099 AND2X1_LOC_155/Y AND2X1_LOC_156/a_8_24# 0.03fF
C30501 VDD AND2X1_LOC_155/Y 0.01fF
C42117 AND2X1_LOC_155/Y AND2X1_LOC_156/a_36_24# 0.01fF
C57386 AND2X1_LOC_155/Y VSS 0.30fF
C2429 OR2X1_LOC_109/Y OR2X1_LOC_323/Y 0.27fF
C10443 AND2X1_LOC_325/a_8_24# OR2X1_LOC_323/Y 0.07fF
C37062 VDD OR2X1_LOC_323/Y 0.44fF
C37133 OR2X1_LOC_315/Y OR2X1_LOC_323/Y 0.08fF
C50077 AND2X1_LOC_543/a_8_24# OR2X1_LOC_323/Y 0.23fF
C52240 OR2X1_LOC_312/Y OR2X1_LOC_323/Y 0.42fF
C56254 OR2X1_LOC_323/Y VSS 0.43fF
C859 VDD OR2X1_LOC_111/Y 0.25fF
C9139 OR2X1_LOC_111/Y AND2X1_LOC_831/Y 0.09fF
C13180 AND2X1_LOC_520/a_8_24# OR2X1_LOC_111/Y 0.02fF
C22243 OR2X1_LOC_109/Y OR2X1_LOC_111/Y 0.40fF
C35641 AND2X1_LOC_326/B OR2X1_LOC_111/Y 0.01fF
C35955 OR2X1_LOC_518/a_8_216# OR2X1_LOC_111/Y 0.13fF
C36055 OR2X1_LOC_111/Y AND2X1_LOC_112/a_8_24# 0.24fF
C38538 OR2X1_LOC_135/Y OR2X1_LOC_111/Y 0.01fF
C38659 OR2X1_LOC_111/Y AND2X1_LOC_520/Y 0.01fF
C41603 OR2X1_LOC_111/Y AND2X1_LOC_715/A 0.01fF
C44164 AND2X1_LOC_332/a_8_24# OR2X1_LOC_111/Y 0.04fF
C47214 OR2X1_LOC_518/Y OR2X1_LOC_111/Y 0.05fF
C49840 AND2X1_LOC_339/B OR2X1_LOC_111/Y 0.01fF
C57393 OR2X1_LOC_111/Y VSS 0.26fF
C2036 OR2X1_LOC_406/Y OR2X1_LOC_527/Y 0.18fF
C2110 OR2X1_LOC_527/Y OR2X1_LOC_496/a_8_216# 0.03fF
C2448 OR2X1_LOC_516/Y OR2X1_LOC_527/Y 0.07fF
C2516 OR2X1_LOC_527/Y AND2X1_LOC_547/a_8_24# -0.00fF
C3819 VDD OR2X1_LOC_527/Y 0.04fF
C9894 OR2X1_LOC_527/Y AND2X1_LOC_840/B 0.10fF
C11578 OR2X1_LOC_189/Y OR2X1_LOC_527/Y 0.07fF
C15752 OR2X1_LOC_527/Y OR2X1_LOC_406/a_8_216# 0.01fF
C19965 OR2X1_LOC_528/Y OR2X1_LOC_527/Y 0.01fF
C22211 OR2X1_LOC_527/Y AND2X1_LOC_621/Y 0.07fF
C28011 AND2X1_LOC_776/a_8_24# OR2X1_LOC_527/Y 0.01fF
C33030 OR2X1_LOC_527/Y AND2X1_LOC_778/Y 0.29fF
C33143 OR2X1_LOC_527/Y AND2X1_LOC_624/A 0.07fF
C35871 OR2X1_LOC_527/Y OR2X1_LOC_142/Y 0.07fF
C39526 OR2X1_LOC_496/Y OR2X1_LOC_527/Y 0.04fF
C40992 AND2X1_LOC_776/Y OR2X1_LOC_527/Y 0.91fF
C45136 AND2X1_LOC_778/a_8_24# OR2X1_LOC_527/Y 0.01fF
C47363 OR2X1_LOC_527/Y OR2X1_LOC_680/A 0.07fF
C57681 OR2X1_LOC_527/Y VSS 0.15fF
C339 AND2X1_LOC_729/B OR2X1_LOC_829/A 0.10fF
C2660 AND2X1_LOC_729/Y AND2X1_LOC_729/B 0.03fF
C3374 AND2X1_LOC_729/B OR2X1_LOC_13/a_8_216# 0.01fF
C14194 AND2X1_LOC_537/Y AND2X1_LOC_729/B 0.02fF
C14419 AND2X1_LOC_729/B OR2X1_LOC_13/Y 1.99fF
C17383 VDD AND2X1_LOC_729/B 0.76fF
C17451 OR2X1_LOC_829/a_8_216# AND2X1_LOC_729/B 0.01fF
C21653 AND2X1_LOC_195/a_8_24# AND2X1_LOC_729/B 0.01fF
C22794 AND2X1_LOC_729/B OR2X1_LOC_41/a_8_216# 0.01fF
C23111 AND2X1_LOC_390/B AND2X1_LOC_729/B 0.62fF
C25208 OR2X1_LOC_311/Y AND2X1_LOC_729/B 0.12fF
C25218 AND2X1_LOC_538/Y AND2X1_LOC_729/B 0.01fF
C28498 OR2X1_LOC_829/a_36_216# AND2X1_LOC_729/B 0.01fF
C30083 AND2X1_LOC_729/a_8_24# AND2X1_LOC_729/B 0.11fF
C30673 AND2X1_LOC_539/a_8_24# AND2X1_LOC_729/B 0.07fF
C32597 AND2X1_LOC_199/A AND2X1_LOC_729/B 0.01fF
C36161 AND2X1_LOC_538/a_8_24# AND2X1_LOC_729/B 0.01fF
C39202 AND2X1_LOC_729/B OR2X1_LOC_41/Y 0.02fF
C44294 AND2X1_LOC_729/B OR2X1_LOC_829/Y 0.14fF
C44321 AND2X1_LOC_729/B OR2X1_LOC_7/Y 0.09fF
C46112 AND2X1_LOC_729/B OR2X1_LOC_311/a_8_216# 0.01fF
C49964 AND2X1_LOC_729/B AND2X1_LOC_855/a_8_24# 0.05fF
C52234 AND2X1_LOC_539/Y AND2X1_LOC_729/B 0.73fF
C53196 AND2X1_LOC_729/B AND2X1_LOC_434/Y 0.01fF
C55433 AND2X1_LOC_729/B AND2X1_LOC_856/B 0.01fF
C57087 AND2X1_LOC_729/B VSS -0.76fF
C9654 OR2X1_LOC_485/Y OR2X1_LOC_516/B 0.24fF
C10596 OR2X1_LOC_516/B OR2X1_LOC_680/A 0.03fF
C21905 OR2X1_LOC_516/Y OR2X1_LOC_516/B 0.01fF
C23282 VDD OR2X1_LOC_516/B 0.18fF
C29244 OR2X1_LOC_516/B AND2X1_LOC_840/B 0.03fF
C35012 AND2X1_LOC_787/A OR2X1_LOC_516/B 0.03fF
C36707 OR2X1_LOC_331/A OR2X1_LOC_516/B 0.82fF
C40723 OR2X1_LOC_516/B AND2X1_LOC_727/A 0.02fF
C43183 OR2X1_LOC_516/B OR2X1_LOC_484/Y 0.28fF
C55482 OR2X1_LOC_516/B OR2X1_LOC_142/Y 0.03fF
C56145 OR2X1_LOC_516/a_8_216# OR2X1_LOC_516/B 0.01fF
C57749 OR2X1_LOC_516/B VSS 0.21fF
C13339 OR2X1_LOC_100/Y OR2X1_LOC_608/Y 0.27fF
C18858 OR2X1_LOC_100/Y AND2X1_LOC_609/a_8_24# 0.23fF
C32592 OR2X1_LOC_100/Y AND2X1_LOC_517/a_8_24# 0.08fF
C45438 OR2X1_LOC_100/Y OR2X1_LOC_520/Y 0.01fF
C50120 OR2X1_LOC_100/Y VDD 0.20fF
C54368 OR2X1_LOC_100/Y OR2X1_LOC_608/a_8_216# 0.03fF
C58026 OR2X1_LOC_100/Y VSS 0.29fF
C4187 VDD AND2X1_LOC_276/Y 0.46fF
C6877 AND2X1_LOC_116/Y AND2X1_LOC_276/Y 0.06fF
C7651 OR2X1_LOC_103/Y AND2X1_LOC_276/Y 0.17fF
C9753 AND2X1_LOC_541/Y AND2X1_LOC_276/Y 0.17fF
C15351 AND2X1_LOC_276/Y AND2X1_LOC_361/A 0.04fF
C17935 AND2X1_LOC_276/Y AND2X1_LOC_473/a_8_24# 0.14fF
C21614 AND2X1_LOC_276/Y AND2X1_LOC_473/Y 0.12fF
C26051 AND2X1_LOC_227/Y AND2X1_LOC_276/Y 0.16fF
C28970 AND2X1_LOC_276/Y AND2X1_LOC_473/a_36_24# 0.01fF
C33545 OR2X1_LOC_521/Y AND2X1_LOC_276/Y 0.04fF
C45004 AND2X1_LOC_715/A AND2X1_LOC_276/Y 0.04fF
C53089 OR2X1_LOC_134/Y AND2X1_LOC_276/Y 0.06fF
C53420 AND2X1_LOC_276/Y OR2X1_LOC_521/a_8_216# 0.13fF
C53518 OR2X1_LOC_106/Y AND2X1_LOC_276/Y 0.02fF
C56960 AND2X1_LOC_276/Y VSS -0.23fF
C2893 VDD AND2X1_LOC_809/A 0.25fF
C8595 AND2X1_LOC_390/B AND2X1_LOC_809/A 0.04fF
C10707 OR2X1_LOC_311/Y AND2X1_LOC_809/A 0.03fF
C22900 AND2X1_LOC_535/Y AND2X1_LOC_809/A 0.01fF
C31659 AND2X1_LOC_809/A AND2X1_LOC_802/Y 0.28fF
C37117 AND2X1_LOC_809/A AND2X1_LOC_809/a_8_24# 0.19fF
C37526 AND2X1_LOC_539/Y AND2X1_LOC_809/A 0.01fF
C38465 AND2X1_LOC_809/A AND2X1_LOC_434/Y 0.04fF
C57024 AND2X1_LOC_809/A VSS 0.10fF
C12027 OR2X1_LOC_461/Y OR2X1_LOC_472/B 0.01fF
C13704 OR2X1_LOC_462/B OR2X1_LOC_461/Y 0.06fF
C46047 OR2X1_LOC_461/Y OR2X1_LOC_462/a_8_216# 0.39fF
C57569 OR2X1_LOC_461/Y VSS 0.18fF
C15218 VDD OR2X1_LOC_240/A 0.11fF
C16179 OR2X1_LOC_462/B OR2X1_LOC_240/A 0.24fF
C31815 OR2X1_LOC_240/B OR2X1_LOC_240/A 0.04fF
C34599 OR2X1_LOC_240/A OR2X1_LOC_397/a_8_216# 0.16fF
C37306 OR2X1_LOC_240/a_8_216# OR2X1_LOC_240/A 0.18fF
C45757 OR2X1_LOC_240/A OR2X1_LOC_397/a_36_216# 0.01fF
C56502 OR2X1_LOC_240/A VSS 0.41fF
C11515 OR2X1_LOC_836/A AND2X1_LOC_823/a_8_24# 0.08fF
C22636 OR2X1_LOC_836/A OR2X1_LOC_836/B 0.07fF
C57548 OR2X1_LOC_836/A VSS 0.25fF
C1823 OR2X1_LOC_334/A OR2X1_LOC_338/A 0.09fF
C5797 AND2X1_LOC_27/a_8_24# OR2X1_LOC_334/A 0.01fF
C8693 OR2X1_LOC_97/A OR2X1_LOC_334/A 0.01fF
C16316 OR2X1_LOC_334/B OR2X1_LOC_334/A 0.48fF
C21918 OR2X1_LOC_634/a_8_216# OR2X1_LOC_334/A 0.47fF
C56256 OR2X1_LOC_334/A VSS 0.22fF
C56845 OR2X1_LOC_751/A VSS 0.11fF
C19697 OR2X1_LOC_715/B OR2X1_LOC_515/Y 0.01fF
C20634 OR2X1_LOC_687/Y OR2X1_LOC_515/Y 0.12fF
C23594 OR2X1_LOC_623/B OR2X1_LOC_515/Y 0.72fF
C25753 OR2X1_LOC_196/B OR2X1_LOC_515/Y 0.33fF
C39583 VDD OR2X1_LOC_515/Y 0.20fF
C40397 OR2X1_LOC_676/Y OR2X1_LOC_515/Y 0.09fF
C44405 OR2X1_LOC_702/A OR2X1_LOC_515/Y 0.10fF
C56274 OR2X1_LOC_515/Y VSS 0.56fF
C34487 OR2X1_LOC_186/Y OR2X1_LOC_355/A 0.01fF
C36398 OR2X1_LOC_622/A OR2X1_LOC_624/B 0.73fF
C3418 OR2X1_LOC_147/B OR2X1_LOC_464/B 0.11fF
C33227 AND2X1_LOC_483/Y AND2X1_LOC_624/A 0.03fF
C55033 OR2X1_LOC_665/Y AND2X1_LOC_483/Y 0.03fF
C21323 AND2X1_LOC_483/Y OR2X1_LOC_816/A 0.11fF
C26996 AND2X1_LOC_483/Y OR2X1_LOC_615/Y 0.38fF
C48704 OR2X1_LOC_252/Y AND2X1_LOC_483/Y 0.18fF
C40772 OR2X1_LOC_613/Y AND2X1_LOC_629/Y 0.14fF
C14046 AND2X1_LOC_456/B OR2X1_LOC_669/Y 0.01fF
C9770 AND2X1_LOC_456/B AND2X1_LOC_286/Y 0.58fF
C5394 AND2X1_LOC_456/B AND2X1_LOC_848/Y 0.03fF
C23825 OR2X1_LOC_251/Y AND2X1_LOC_456/B 0.02fF
C32118 OR2X1_LOC_667/Y AND2X1_LOC_456/B 0.04fF
C9637 AND2X1_LOC_456/B OR2X1_LOC_253/Y 0.79fF
C38406 AND2X1_LOC_456/B OR2X1_LOC_666/A 0.02fF
C15235 AND2X1_LOC_456/B AND2X1_LOC_287/Y 0.48fF
C46277 AND2X1_LOC_456/B AND2X1_LOC_843/Y 0.01fF
C40891 AND2X1_LOC_456/B OR2X1_LOC_816/A 1.23fF
C34425 AND2X1_LOC_456/B AND2X1_LOC_721/A 0.04fF
C46899 AND2X1_LOC_456/B OR2X1_LOC_615/Y 0.03fF
C36805 AND2X1_LOC_456/B OR2X1_LOC_669/A 0.01fF
C52182 OR2X1_LOC_494/Y AND2X1_LOC_456/B 0.47fF
C24261 AND2X1_LOC_456/B OR2X1_LOC_666/Y 0.01fF
C3713 OR2X1_LOC_669/Y AND2X1_LOC_287/B 0.03fF
C51353 AND2X1_LOC_848/Y AND2X1_LOC_287/B 0.03fF
C13491 OR2X1_LOC_251/Y AND2X1_LOC_287/B 0.08fF
C26585 OR2X1_LOC_669/A AND2X1_LOC_287/B 0.77fF
C40585 OR2X1_LOC_279/Y AND2X1_LOC_287/B 0.01fF
C787 OR2X1_LOC_848/B OR2X1_LOC_392/A 0.71fF
C44353 OR2X1_LOC_848/B OR2X1_LOC_561/B 0.04fF
C34711 OR2X1_LOC_848/B OR2X1_LOC_391/A 0.07fF
C15406 OR2X1_LOC_285/Y OR2X1_LOC_285/B 0.03fF
C53632 OR2X1_LOC_190/A OR2X1_LOC_456/A 0.10fF
C51002 AND2X1_LOC_99/Y OR2X1_LOC_517/A 0.08fF
C43412 AND2X1_LOC_99/Y OR2X1_LOC_813/Y 0.03fF
C10959 OR2X1_LOC_216/A AND2X1_LOC_492/a_8_24# 0.05fF
C18901 OR2X1_LOC_216/A AND2X1_LOC_239/a_36_24# 0.01fF
C57570 OR2X1_LOC_216/A VSS -0.21fF
C37445 OR2X1_LOC_139/A OR2X1_LOC_267/Y 0.03fF
C46644 OR2X1_LOC_185/Y OR2X1_LOC_267/Y 0.03fF
C31587 OR2X1_LOC_140/A OR2X1_LOC_267/Y 0.06fF
C53899 OR2X1_LOC_643/A OR2X1_LOC_267/Y 0.03fF
C26443 OR2X1_LOC_436/Y OR2X1_LOC_802/Y 0.01fF
C21301 OR2X1_LOC_802/Y OR2X1_LOC_539/Y 0.05fF
C17857 OR2X1_LOC_802/Y OR2X1_LOC_809/a_8_216# 0.11fF
C57196 OR2X1_LOC_802/Y VSS 0.10fF
C30431 OR2X1_LOC_163/A OR2X1_LOC_163/Y 0.01fF
C15434 AND2X1_LOC_436/B OR2X1_LOC_331/Y 0.02fF
C30278 AND2X1_LOC_841/B OR2X1_LOC_331/Y 0.03fF
C12529 AND2X1_LOC_390/B OR2X1_LOC_331/Y 0.02fF
C49161 AND2X1_LOC_356/B OR2X1_LOC_331/Y 0.01fF
C30650 OR2X1_LOC_166/Y OR2X1_LOC_331/Y 0.18fF
C20540 OR2X1_LOC_331/A OR2X1_LOC_331/Y 0.11fF
C40750 OR2X1_LOC_533/Y OR2X1_LOC_331/Y 0.16fF
C1099 OR2X1_LOC_167/Y OR2X1_LOC_331/Y 0.02fF
C5832 OR2X1_LOC_533/A OR2X1_LOC_331/Y 0.01fF
C21900 OR2X1_LOC_312/Y OR2X1_LOC_331/Y 0.51fF
C26839 AND2X1_LOC_535/Y OR2X1_LOC_331/Y 0.03fF
C50443 OR2X1_LOC_680/A OR2X1_LOC_331/Y 0.13fF
C55737 AND2X1_LOC_729/Y AND2X1_LOC_621/Y 0.03fF
C31866 AND2X1_LOC_727/A AND2X1_LOC_621/Y 0.07fF
C17 OR2X1_LOC_755/A AND2X1_LOC_621/Y 0.10fF
C43736 AND2X1_LOC_621/Y AND2X1_LOC_624/A 20.56fF
C33173 OR2X1_LOC_504/Y AND2X1_LOC_621/Y 0.03fF
C32601 OR2X1_LOC_438/Y AND2X1_LOC_621/Y 0.03fF
C48011 OR2X1_LOC_177/Y AND2X1_LOC_621/Y 0.03fF
C9422 OR2X1_LOC_665/Y AND2X1_LOC_621/Y 0.07fF
C22959 OR2X1_LOC_441/Y AND2X1_LOC_621/Y 0.03fF
C24234 OR2X1_LOC_525/Y AND2X1_LOC_621/Y 0.06fF
C8601 OR2X1_LOC_680/Y AND2X1_LOC_621/Y 0.03fF
C53528 OR2X1_LOC_759/A AND2X1_LOC_621/Y 0.03fF
C46581 AND2X1_LOC_621/Y OR2X1_LOC_142/Y 0.03fF
C46726 AND2X1_LOC_621/Y OR2X1_LOC_442/Y 0.02fF
C2047 OR2X1_LOC_757/A AND2X1_LOC_621/Y 0.03fF
C13001 OR2X1_LOC_516/Y AND2X1_LOC_621/Y 0.07fF
C52412 OR2X1_LOC_617/Y AND2X1_LOC_621/Y 0.15fF
C43346 AND2X1_LOC_154/Y AND2X1_LOC_621/Y 0.14fF
C6340 AND2X1_LOC_621/Y OR2X1_LOC_239/Y 0.03fF
C44176 OR2X1_LOC_613/Y AND2X1_LOC_621/Y 0.01fF
C31655 AND2X1_LOC_621/Y OR2X1_LOC_816/A 0.06fF
C53972 AND2X1_LOC_508/A AND2X1_LOC_621/Y 0.03fF
C1701 OR2X1_LOC_680/A AND2X1_LOC_621/Y 0.03fF
C47877 AND2X1_LOC_621/Y OR2X1_LOC_152/A 0.03fF
C37415 AND2X1_LOC_621/Y OR2X1_LOC_615/Y 0.03fF
C19248 OR2X1_LOC_146/Y AND2X1_LOC_621/Y 0.02fF
C14407 OR2X1_LOC_677/Y AND2X1_LOC_621/Y 0.03fF
C36113 OR2X1_LOC_679/A AND2X1_LOC_621/Y 0.04fF
C2998 OR2X1_LOC_252/Y AND2X1_LOC_621/Y 0.03fF
C14459 OR2X1_LOC_616/Y AND2X1_LOC_621/Y 0.14fF
C50283 OR2X1_LOC_496/Y AND2X1_LOC_621/Y 0.03fF
C14917 OR2X1_LOC_666/Y AND2X1_LOC_621/Y 0.03fF
C11804 OR2X1_LOC_526/Y AND2X1_LOC_621/Y 0.08fF
C30430 OR2X1_LOC_528/Y AND2X1_LOC_621/Y 0.01fF
C27914 OR2X1_LOC_501/B OR2X1_LOC_629/Y 0.01fF
C42076 OR2X1_LOC_837/Y AND2X1_LOC_462/Y 0.01fF
C7556 OR2X1_LOC_837/A OR2X1_LOC_837/Y 0.02fF
C38732 AND2X1_LOC_848/A AND2X1_LOC_848/Y 0.07fF
C35697 AND2X1_LOC_711/A AND2X1_LOC_848/A 0.01fF
C42659 OR2X1_LOC_755/A AND2X1_LOC_848/A 0.23fF
C39620 OR2X1_LOC_258/Y AND2X1_LOC_848/A 0.01fF
C39918 OR2X1_LOC_759/A AND2X1_LOC_848/A 0.02fF
C39954 OR2X1_LOC_698/Y AND2X1_LOC_848/A 0.05fF
C10191 AND2X1_LOC_848/A AND2X1_LOC_789/Y 0.21fF
C56062 AND2X1_LOC_848/A AND2X1_LOC_793/B 0.03fF
C54232 OR2X1_LOC_295/Y AND2X1_LOC_848/A 0.02fF
C3780 OR2X1_LOC_251/Y AND2X1_LOC_285/Y 0.02fF
C20821 OR2X1_LOC_282/Y AND2X1_LOC_285/Y 0.80fF
C21036 OR2X1_LOC_816/A AND2X1_LOC_285/Y 0.03fF
C26809 OR2X1_LOC_615/Y AND2X1_LOC_285/Y 0.02fF
C31802 OR2X1_LOC_632/A OR2X1_LOC_631/B 0.01fF
C33460 OR2X1_LOC_631/B OR2X1_LOC_630/Y 0.04fF
C45502 OR2X1_LOC_664/Y OR2X1_LOC_631/B 0.18fF
C15542 OR2X1_LOC_631/B OR2X1_LOC_115/B 0.05fF
C21 OR2X1_LOC_631/B OR2X1_LOC_574/A 0.02fF
C40751 OR2X1_LOC_631/B OR2X1_LOC_629/A 0.16fF
C26915 OR2X1_LOC_631/B OR2X1_LOC_247/Y 0.03fF
C55228 OR2X1_LOC_631/B OR2X1_LOC_629/B 0.02fF
C54046 OR2X1_LOC_254/B OR2X1_LOC_631/B 0.05fF
C54033 OR2X1_LOC_631/B OR2X1_LOC_833/B 0.02fF
C52308 OR2X1_LOC_501/B OR2X1_LOC_631/B 0.03fF
C20428 OR2X1_LOC_631/B AND2X1_LOC_72/Y 0.03fF
C20741 OR2X1_LOC_631/B OR2X1_LOC_719/B 0.03fF
C45088 OR2X1_LOC_287/A OR2X1_LOC_288/A 0.10fF
C36363 OR2X1_LOC_791/B OR2X1_LOC_287/A 0.20fF
C35779 OR2X1_LOC_177/Y AND2X1_LOC_464/A 0.01fF
C17301 OR2X1_LOC_312/Y AND2X1_LOC_464/A 0.01fF
C26049 AND2X1_LOC_543/Y AND2X1_LOC_464/A 0.01fF
C23680 OR2X1_LOC_109/Y AND2X1_LOC_464/A 0.02fF
C44493 OR2X1_LOC_280/Y AND2X1_LOC_464/A 0.03fF
C42006 OR2X1_LOC_656/B OR2X1_LOC_99/Y 0.24fF
C17223 OR2X1_LOC_99/Y OR2X1_LOC_771/B 0.05fF
C14372 OR2X1_LOC_99/Y OR2X1_LOC_646/B 0.01fF
C867 OR2X1_LOC_520/Y OR2X1_LOC_99/Y 0.02fF
C49043 AND2X1_LOC_489/Y AND2X1_LOC_361/A 0.02fF
C28987 AND2X1_LOC_227/Y AND2X1_LOC_361/A 0.01fF
C36409 OR2X1_LOC_517/A AND2X1_LOC_361/A 0.09fF
C41154 OR2X1_LOC_265/Y AND2X1_LOC_361/A 0.03fF
C49137 AND2X1_LOC_216/A AND2X1_LOC_361/A 0.02fF
C41908 OR2X1_LOC_131/A AND2X1_LOC_361/A 0.11fF
C56016 OR2X1_LOC_134/Y AND2X1_LOC_361/A 0.04fF
C22915 AND2X1_LOC_361/A OR2X1_LOC_595/A 1.01fF
C27973 OR2X1_LOC_132/Y AND2X1_LOC_361/A 0.02fF
C15711 AND2X1_LOC_139/B AND2X1_LOC_361/A 0.02fF
C52398 AND2X1_LOC_266/Y AND2X1_LOC_361/A 0.08fF
C12670 AND2X1_LOC_541/Y AND2X1_LOC_361/A 0.03fF
C237 OR2X1_LOC_106/Y AND2X1_LOC_361/A 0.74fF
C10623 OR2X1_LOC_103/Y AND2X1_LOC_361/A 0.17fF
C27310 AND2X1_LOC_116/B AND2X1_LOC_116/Y 0.26fF
C12441 AND2X1_LOC_116/Y AND2X1_LOC_473/a_8_24# 0.20fF
C45642 AND2X1_LOC_116/a_8_24# AND2X1_LOC_116/Y 0.01fF
C4425 AND2X1_LOC_802/Y AND2X1_LOC_434/Y 0.02fF
C35455 AND2X1_LOC_319/A AND2X1_LOC_802/Y 0.81fF
C12990 AND2X1_LOC_436/Y AND2X1_LOC_802/Y 0.03fF
C46743 AND2X1_LOC_798/Y AND2X1_LOC_802/Y 0.16fF
C20157 AND2X1_LOC_802/B AND2X1_LOC_802/Y 0.11fF
C3576 AND2X1_LOC_539/Y AND2X1_LOC_802/Y 0.10fF
C24273 AND2X1_LOC_798/A AND2X1_LOC_802/Y 0.46fF
C3176 AND2X1_LOC_802/Y AND2X1_LOC_809/a_8_24# 0.03fF
C12697 AND2X1_LOC_802/a_8_24# AND2X1_LOC_802/Y 0.03fF
C18727 AND2X1_LOC_319/a_8_24# AND2X1_LOC_802/Y 0.01fF
C23552 AND2X1_LOC_798/a_8_24# AND2X1_LOC_802/Y 0.04fF
C40095 AND2X1_LOC_362/B AND2X1_LOC_99/A 0.04fF
C19062 AND2X1_LOC_99/A OR2X1_LOC_517/A 0.03fF
C22118 AND2X1_LOC_99/A OR2X1_LOC_118/Y 0.02fF
C5293 AND2X1_LOC_99/A OR2X1_LOC_595/A 0.03fF
C4521 AND2X1_LOC_99/A OR2X1_LOC_666/A 0.37fF
C46052 AND2X1_LOC_99/A OR2X1_LOC_67/Y 0.22fF
C49336 AND2X1_LOC_99/A AND2X1_LOC_98/Y 0.02fF
C50271 AND2X1_LOC_99/A OR2X1_LOC_117/Y 0.66fF
C31372 AND2X1_LOC_99/A OR2X1_LOC_67/A 0.01fF
C7566 OR2X1_LOC_122/Y AND2X1_LOC_99/A 0.02fF
C38818 OR2X1_LOC_106/Y AND2X1_LOC_99/A 0.03fF
C49994 OR2X1_LOC_116/A OR2X1_LOC_66/Y 0.01fF
C865 OR2X1_LOC_185/Y OR2X1_LOC_114/Y 0.05fF
C37332 OR2X1_LOC_114/Y OR2X1_LOC_810/A 0.05fF
C13125 OR2X1_LOC_114/Y OR2X1_LOC_362/A 0.01fF
C8214 OR2X1_LOC_114/Y OR2X1_LOC_113/A 0.81fF
C6899 OR2X1_LOC_436/Y OR2X1_LOC_802/A 0.01fF
C34727 OR2X1_LOC_798/Y OR2X1_LOC_802/A 0.13fF
C1721 OR2X1_LOC_539/Y OR2X1_LOC_802/A 0.01fF
C40195 OR2X1_LOC_802/a_8_216# OR2X1_LOC_802/A 0.39fF
C2525 OR2X1_LOC_799/A OR2X1_LOC_798/Y 0.25fF
C23495 OR2X1_LOC_798/Y OR2X1_LOC_436/Y 0.01fF
C22067 OR2X1_LOC_318/Y OR2X1_LOC_798/Y 0.05fF
C722 OR2X1_LOC_798/Y OR2X1_LOC_802/a_8_216# 0.01fF
C23803 OR2X1_LOC_798/Y OR2X1_LOC_799/a_8_216# 0.48fF
C40019 OR2X1_LOC_99/B OR2X1_LOC_99/A 0.27fF
C51572 OR2X1_LOC_329/B AND2X1_LOC_114/Y 0.01fF
C9396 AND2X1_LOC_715/A AND2X1_LOC_116/B 0.01fF
C49873 OR2X1_LOC_329/B AND2X1_LOC_116/B 0.02fF
C54081 OR2X1_LOC_521/Y AND2X1_LOC_116/B 0.81fF
C17731 OR2X1_LOC_106/Y AND2X1_LOC_116/B 0.03fF
C17780 VDD AND2X1_LOC_798/Y -0.00fF
C52663 AND2X1_LOC_539/Y AND2X1_LOC_798/Y 0.19fF
C35347 AND2X1_LOC_802/B AND2X1_LOC_436/Y 0.01fF
C35101 AND2X1_LOC_802/B AND2X1_LOC_802/a_8_24# 0.10fF
C47488 AND2X1_LOC_802/B VDD 0.01fF
C51335 OR2X1_LOC_113/Y OR2X1_LOC_362/A 0.13fF
C22859 OR2X1_LOC_113/Y OR2X1_LOC_114/B 0.16fF
C31570 OR2X1_LOC_113/Y OR2X1_LOC_844/B 0.02fF
C46317 OR2X1_LOC_113/Y OR2X1_LOC_643/A 0.01fF
C26681 OR2X1_LOC_799/A OR2X1_LOC_435/B 0.04fF
C45506 OR2X1_LOC_799/A OR2X1_LOC_574/A 0.15fF
C48136 OR2X1_LOC_405/A OR2X1_LOC_799/A 0.03fF
C15084 OR2X1_LOC_799/A OR2X1_LOC_593/B 0.17fF
C17831 OR2X1_LOC_799/A OR2X1_LOC_449/B 0.25fF
C44217 OR2X1_LOC_592/A OR2X1_LOC_799/A 0.03fF
C25477 OR2X1_LOC_799/A OR2X1_LOC_539/Y 0.16fF
C46502 OR2X1_LOC_436/Y OR2X1_LOC_539/Y 0.05fF
C45006 OR2X1_LOC_318/Y OR2X1_LOC_539/Y 0.03fF
C18233 OR2X1_LOC_798/Y OR2X1_LOC_539/Y 0.44fF
C37728 OR2X1_LOC_809/a_8_216# OR2X1_LOC_539/Y 0.04fF
C41348 OR2X1_LOC_539/Y OR2X1_LOC_319/Y 0.03fF
C46826 OR2X1_LOC_539/Y OR2X1_LOC_799/a_8_216# 0.01fF
C56610 OR2X1_LOC_539/Y VSS -0.32fF
C6576 OR2X1_LOC_436/Y OR2X1_LOC_854/A 0.03fF
C14039 OR2X1_LOC_139/A OR2X1_LOC_436/Y 0.15fF
C401 OR2X1_LOC_436/Y OR2X1_LOC_390/A 0.01fF
C9802 OR2X1_LOC_186/Y OR2X1_LOC_436/Y 0.02fF
C23122 OR2X1_LOC_185/Y OR2X1_LOC_436/Y 0.03fF
C10001 OR2X1_LOC_436/Y OR2X1_LOC_112/B 0.02fF
C3560 OR2X1_LOC_436/Y OR2X1_LOC_810/A 0.23fF
C10353 OR2X1_LOC_574/A OR2X1_LOC_436/Y 0.03fF
C3860 OR2X1_LOC_715/B OR2X1_LOC_436/Y 0.04fF
C12871 OR2X1_LOC_405/A OR2X1_LOC_436/Y 0.03fF
C45235 OR2X1_LOC_319/B OR2X1_LOC_319/Y 0.03fF
C46748 OR2X1_LOC_436/Y OR2X1_LOC_319/Y 0.14fF
C5679 OR2X1_LOC_319/a_8_216# OR2X1_LOC_319/Y -0.00fF
C40903 OR2X1_LOC_798/a_8_216# OR2X1_LOC_319/Y 0.07fF
C42990 AND2X1_LOC_227/Y AND2X1_LOC_113/Y 0.01fF
C24613 OR2X1_LOC_103/Y AND2X1_LOC_113/Y 0.01fF
C6033 AND2X1_LOC_319/A AND2X1_LOC_798/A 0.17fF
C50223 AND2X1_LOC_798/a_8_24# AND2X1_LOC_798/A 0.18fF
C57191 AND2X1_LOC_798/A VSS 0.15fF
C24052 AND2X1_LOC_436/Y AND2X1_LOC_810/B 0.03fF
C7530 AND2X1_LOC_841/B AND2X1_LOC_436/Y 0.03fF
C1715 AND2X1_LOC_727/A AND2X1_LOC_436/Y 0.01fF
C45872 AND2X1_LOC_390/B AND2X1_LOC_436/Y 0.02fF
C7923 OR2X1_LOC_166/Y AND2X1_LOC_436/Y 0.01fF
C43617 OR2X1_LOC_594/Y AND2X1_LOC_436/Y 0.01fF
C34351 OR2X1_LOC_167/Y AND2X1_LOC_436/Y 0.26fF
C39130 AND2X1_LOC_436/Y OR2X1_LOC_533/A 0.02fF
C55265 OR2X1_LOC_312/Y AND2X1_LOC_436/Y 0.03fF
C4067 AND2X1_LOC_535/Y AND2X1_LOC_436/Y 1.13fF
C27500 OR2X1_LOC_680/A AND2X1_LOC_436/Y 0.18fF
C4087 OR2X1_LOC_484/Y AND2X1_LOC_436/Y 0.13fF
C10423 AND2X1_LOC_539/Y AND2X1_LOC_434/Y 0.04fF
C41385 AND2X1_LOC_539/Y AND2X1_LOC_319/A 0.02fF
C17630 AND2X1_LOC_539/Y AND2X1_LOC_593/Y 0.09fF
C41612 AND2X1_LOC_539/Y OR2X1_LOC_331/Y 0.06fF
C18898 AND2X1_LOC_539/Y AND2X1_LOC_436/Y 0.02fF
C26038 AND2X1_LOC_539/Y AND2X1_LOC_802/B 0.61fF
C9106 AND2X1_LOC_539/Y AND2X1_LOC_809/a_8_24# 0.01fF
C18610 AND2X1_LOC_539/Y AND2X1_LOC_802/a_8_24# 0.01fF
C30788 AND2X1_LOC_539/Y OR2X1_LOC_829/a_8_216# 0.01fF
C24262 AND2X1_LOC_729/Y AND2X1_LOC_593/Y 0.07fF
C466 AND2X1_LOC_727/A AND2X1_LOC_593/Y 0.01fF
C16835 OR2X1_LOC_533/Y AND2X1_LOC_593/Y 0.11fF
C42405 AND2X1_LOC_593/Y OR2X1_LOC_594/Y 0.17fF
C4124 AND2X1_LOC_593/Y AND2X1_LOC_447/Y 0.07fF
C16820 OR2X1_LOC_176/Y AND2X1_LOC_593/Y 0.03fF
C14132 OR2X1_LOC_574/A OR2X1_LOC_593/A 0.08fF
C39676 OR2X1_LOC_593/A OR2X1_LOC_593/B 0.06fF
C42511 OR2X1_LOC_449/B OR2X1_LOC_593/A 0.02fF
C42030 OR2X1_LOC_539/A OR2X1_LOC_193/A 0.01fF
C12347 OR2X1_LOC_539/A OR2X1_LOC_702/A 0.78fF
C15810 OR2X1_LOC_539/B OR2X1_LOC_390/A 0.04fF
C31907 OR2X1_LOC_97/A OR2X1_LOC_539/B 0.02fF
C17876 OR2X1_LOC_339/A OR2X1_LOC_539/B 0.03fF
C49296 OR2X1_LOC_434/A OR2X1_LOC_539/B 0.05fF
C12497 OR2X1_LOC_174/A OR2X1_LOC_539/B 0.23fF
C32893 OR2X1_LOC_333/B OR2X1_LOC_539/B 0.02fF
C48786 OR2X1_LOC_139/A OR2X1_LOC_436/B 0.01fF
C8382 OR2X1_LOC_186/Y OR2X1_LOC_318/Y 0.03fF
C15117 OR2X1_LOC_97/A OR2X1_LOC_318/Y 0.02fF
C46264 OR2X1_LOC_318/Y OR2X1_LOC_435/B 0.16fF
C18566 OR2X1_LOC_318/Y OR2X1_LOC_776/Y 0.73fF
C37273 OR2X1_LOC_318/Y OR2X1_LOC_449/B 0.08fF
C5348 OR2X1_LOC_318/Y OR2X1_LOC_538/A 0.12fF
C5173 OR2X1_LOC_319/B OR2X1_LOC_854/A 0.02fF
C8366 OR2X1_LOC_186/Y OR2X1_LOC_319/B 0.02fF
C8952 OR2X1_LOC_319/B OR2X1_LOC_574/A 0.03fF
C24562 OR2X1_LOC_319/B OR2X1_LOC_840/A 0.10fF
C28836 OR2X1_LOC_319/B OR2X1_LOC_778/Y 0.10fF
C11404 OR2X1_LOC_405/A OR2X1_LOC_319/B 0.09fF
C1528 OR2X1_LOC_319/B OR2X1_LOC_356/A 0.15fF
C37263 OR2X1_LOC_319/B OR2X1_LOC_449/B 0.07fF
C14016 OR2X1_LOC_319/B OR2X1_LOC_703/B 0.03fF
C33397 OR2X1_LOC_319/B OR2X1_LOC_703/A 0.01fF
C46668 AND2X1_LOC_319/A AND2X1_LOC_810/B 0.08fF
C48177 AND2X1_LOC_729/Y AND2X1_LOC_319/A 0.02fF
C1574 AND2X1_LOC_706/Y AND2X1_LOC_319/A 0.07fF
C49028 AND2X1_LOC_356/B AND2X1_LOC_319/A 0.33fF
C29982 AND2X1_LOC_707/Y AND2X1_LOC_319/A 0.07fF
C51513 OR2X1_LOC_313/Y AND2X1_LOC_319/A 0.01fF
C26652 AND2X1_LOC_535/Y AND2X1_LOC_319/A 0.02fF
C31753 OR2X1_LOC_329/B AND2X1_LOC_319/A 0.44fF
C14546 OR2X1_LOC_311/Y AND2X1_LOC_319/A 0.16fF
C54852 AND2X1_LOC_319/A OR2X1_LOC_432/Y 0.19fF
C52331 AND2X1_LOC_318/Y AND2X1_LOC_473/Y 0.02fF
C52535 AND2X1_LOC_727/A AND2X1_LOC_318/Y 0.02fF
C13674 AND2X1_LOC_326/B AND2X1_LOC_318/Y 0.02fF
C20130 AND2X1_LOC_784/A AND2X1_LOC_318/Y 0.02fF
C47770 AND2X1_LOC_335/Y AND2X1_LOC_318/Y 0.51fF
C72 OR2X1_LOC_109/Y AND2X1_LOC_318/Y 0.02fF
C13631 AND2X1_LOC_856/B AND2X1_LOC_434/Y 0.01fF
C40146 AND2X1_LOC_436/B AND2X1_LOC_434/Y 0.01fF
C55212 AND2X1_LOC_841/B AND2X1_LOC_434/Y 0.07fF
C14690 OR2X1_LOC_829/A AND2X1_LOC_434/Y 0.10fF
C37260 AND2X1_LOC_390/B AND2X1_LOC_434/Y 0.01fF
C17771 AND2X1_LOC_356/B AND2X1_LOC_434/Y 0.01fF
C53747 OR2X1_LOC_41/Y AND2X1_LOC_434/Y 0.01fF
C55564 OR2X1_LOC_166/Y AND2X1_LOC_434/Y 0.16fF
C2589 OR2X1_LOC_829/Y AND2X1_LOC_434/Y 0.01fF
C25934 OR2X1_LOC_167/Y AND2X1_LOC_434/Y 0.01fF
C17118 AND2X1_LOC_434/Y OR2X1_LOC_172/Y 0.01fF
C46788 OR2X1_LOC_312/Y AND2X1_LOC_434/Y 0.07fF
C662 OR2X1_LOC_329/B AND2X1_LOC_434/Y 0.07fF
C39453 OR2X1_LOC_311/Y AND2X1_LOC_434/Y 0.15fF
C28657 OR2X1_LOC_13/Y AND2X1_LOC_434/Y 0.02fF
C49310 OR2X1_LOC_45/Y AND2X1_LOC_434/Y 0.95fF
C41530 AND2X1_LOC_339/B AND2X1_LOC_537/Y 0.22fF
C54576 AND2X1_LOC_390/B AND2X1_LOC_537/Y 0.04fF
C488 OR2X1_LOC_305/Y AND2X1_LOC_537/Y 0.07fF
C55854 AND2X1_LOC_303/B AND2X1_LOC_537/Y 0.06fF
C43844 AND2X1_LOC_303/A AND2X1_LOC_537/Y 0.02fF
C544 OR2X1_LOC_311/Y AND2X1_LOC_537/Y 0.02fF
C28636 AND2X1_LOC_537/Y OR2X1_LOC_595/Y 0.14fF
C30497 OR2X1_LOC_135/Y AND2X1_LOC_537/Y 0.15fF
C9527 AND2X1_LOC_390/B AND2X1_LOC_538/Y 0.02fF
C11631 OR2X1_LOC_311/Y AND2X1_LOC_538/Y 0.02fF
C6969 AND2X1_LOC_592/Y AND2X1_LOC_706/Y 0.16fF
C33293 AND2X1_LOC_592/Y AND2X1_LOC_447/Y 0.02fF
C35279 AND2X1_LOC_592/Y OR2X1_LOC_424/Y 0.89fF
C212 OR2X1_LOC_132/a_8_216# VDD 0.21fF
C313 OR2X1_LOC_533/a_8_216# OR2X1_LOC_331/a_8_216# 0.47fF
C430 OR2X1_LOC_280/a_8_216# OR2X1_LOC_237/a_8_216# 0.47fF
C747 VDD AND2X1_LOC_158/a_8_24# -0.00fF
C758 VDD AND2X1_LOC_638/a_8_24# -0.00fF
C1239 VDD OR2X1_LOC_438/a_8_216# 0.21fF
C1697 VDD AND2X1_LOC_101/a_8_24# -0.00fF
C2300 VDD OR2X1_LOC_320/a_8_216# 0.21fF
C3293 AND2X1_LOC_83/a_8_24# AND2X1_LOC_617/a_8_24# 0.23fF
C3731 VDD AND2X1_LOC_166/a_8_24# -0.00fF
C3811 VDD AND2X1_LOC_183/a_8_24# -0.00fF
C4066 AND2X1_LOC_60/a_8_24# AND2X1_LOC_58/a_8_24# 0.23fF
C4135 VDD OR2X1_LOC_457/a_8_216# 0.21fF
C4148 VDD OR2X1_LOC_701/a_8_216# 0.21fF
C4838 OR2X1_LOC_135/a_8_216# VDD 0.21fF
C4897 VDD OR2X1_LOC_828/a_8_216# 0.21fF
C4932 VDD AND2X1_LOC_695/a_8_24# -0.00fF
C5118 VDD OR2X1_LOC_173/a_8_216# 0.21fF
C5257 VDD OR2X1_LOC_108/a_8_216# 0.21fF
C5493 AND2X1_LOC_631/a_8_24# AND2X1_LOC_483/a_8_24# 0.23fF
C5734 VDD OR2X1_LOC_298/a_8_216# 0.21fF
C5788 VDD OR2X1_LOC_664/a_8_216# 0.21fF
C5890 OR2X1_LOC_481/a_8_216# OR2X1_LOC_700/a_8_216# 0.47fF
C6200 VDD OR2X1_LOC_109/a_8_216# 0.21fF
C6242 VDD OR2X1_LOC_24/a_8_216# 0.21fF
C6279 AND2X1_LOC_701/a_8_24# AND2X1_LOC_526/a_8_24# 0.23fF
C6676 AND2X1_LOC_393/a_8_24# VDD -0.00fF
C6723 VDD OR2X1_LOC_52/a_8_216# 0.21fF
C6801 OR2X1_LOC_178/a_8_216# OR2X1_LOC_224/a_8_216# 0.47fF
C7459 VDD OR2X1_LOC_832/a_8_216# 0.21fF
C8438 VDD OR2X1_LOC_257/a_8_216# 0.21fF
C8749 VDD AND2X1_LOC_729/a_8_24# -0.00fF
C9289 VDD OR2X1_LOC_613/a_8_216# 0.21fF
C9566 VDD AND2X1_LOC_258/a_8_24# -0.00fF
C9580 VDD OR2X1_LOC_708/a_8_216# 0.21fF
C10510 OR2X1_LOC_101/a_8_216# VDD 0.21fF
C10530 VDD OR2X1_LOC_447/a_8_216# 0.21fF
C10724 OR2X1_LOC_626/a_8_216# OR2X1_LOC_617/a_8_216# 0.47fF
C11046 OR2X1_LOC_83/a_8_216# OR2X1_LOC_394/a_8_216# 0.47fF
C11082 VDD OR2X1_LOC_75/a_8_216# 0.21fF
C11188 VDD OR2X1_LOC_195/a_8_216# 0.21fF
C11378 OR2X1_LOC_813/a_8_216# OR2X1_LOC_235/a_8_216# 0.47fF
C12275 VDD AND2X1_LOC_105/a_8_24# -0.00fF
C12284 AND2X1_LOC_522/a_8_24# AND2X1_LOC_107/a_8_24# 0.23fF
C12718 VDD AND2X1_LOC_525/a_8_24# -0.00fF
C12956 VDD AND2X1_LOC_590/a_8_24# -0.00fF
C13132 OR2X1_LOC_831/a_8_216# VDD 0.21fF
C13476 VDD OR2X1_LOC_251/a_8_216# 0.21fF
C13841 VDD AND2X1_LOC_524/a_8_24# -0.00fF
C13909 VDD AND2X1_LOC_253/a_8_24# -0.00fF
C15598 AND2X1_LOC_767/a_8_24# AND2X1_LOC_396/a_8_24# 0.23fF
C15858 VDD OR2X1_LOC_333/a_8_216# 0.21fF
C15906 VDD OR2X1_LOC_584/a_8_216# 0.21fF
C16010 AND2X1_LOC_586/a_8_24# VDD -0.00fF
C16164 VDD OR2X1_LOC_780/a_8_216# 0.21fF
C16169 AND2X1_LOC_99/a_8_24# AND2X1_LOC_101/a_8_24# 0.23fF
C16694 VDD OR2X1_LOC_535/a_8_216# 0.21fF
C16741 AND2X1_LOC_680/a_8_24# AND2X1_LOC_420/a_8_24# 0.23fF
C17181 VDD AND2X1_LOC_60/a_8_24# -0.00fF
C17193 VDD OR2X1_LOC_759/a_8_216# 0.21fF
C17298 VDD AND2X1_LOC_504/a_8_24# -0.00fF
C18234 VDD OR2X1_LOC_258/a_8_216# 0.21fF
C18235 OR2X1_LOC_848/a_8_216# OR2X1_LOC_391/a_8_216# 0.47fF
C18529 VDD AND2X1_LOC_172/a_8_24# -0.00fF
C18899 OR2X1_LOC_176/a_8_216# VDD 0.21fF
C19198 VDD AND2X1_LOC_237/a_8_24# -0.00fF
C19316 OR2X1_LOC_188/a_8_216# VDD -0.00fF
C20420 OR2X1_LOC_816/a_8_216# OR2X1_LOC_253/a_8_216# 0.47fF
C20583 OR2X1_LOC_484/a_8_216# OR2X1_LOC_142/a_8_216# 0.47fF
C20662 OR2X1_LOC_285/a_8_216# OR2X1_LOC_758/a_8_216# 0.47fF
C20811 OR2X1_LOC_167/a_8_216# OR2X1_LOC_601/a_8_216# 0.47fF
C21073 VDD OR2X1_LOC_777/a_8_216# 0.21fF
C21470 VDD OR2X1_LOC_525/a_8_216# 0.21fF
C21541 AND2X1_LOC_266/a_8_24# AND2X1_LOC_249/a_8_24# 0.23fF
C21635 VDD OR2X1_LOC_790/a_8_216# 0.21fF
C22095 VDD AND2X1_LOC_528/a_8_24# -0.00fF
C22377 VDD OR2X1_LOC_621/a_8_216# 0.21fF
C22466 VDD AND2X1_LOC_161/a_8_24# -0.00fF
C22529 AND2X1_LOC_117/a_8_24# AND2X1_LOC_262/a_8_24# 0.23fF
C22862 VDD AND2X1_LOC_103/a_8_24# -0.00fF
C24711 AND2X1_LOC_379/a_8_24# AND2X1_LOC_638/a_8_24# 0.23fF
C25125 VDD OR2X1_LOC_751/a_8_216# 0.21fF
C25353 AND2X1_LOC_757/a_8_24# VDD -0.00fF
C26422 VDD OR2X1_LOC_172/a_8_216# 0.21fF
C26654 AND2X1_LOC_843/a_8_24# AND2X1_LOC_286/a_8_24# 0.23fF
C26665 AND2X1_LOC_186/a_8_24# AND2X1_LOC_188/a_8_24# 0.23fF
C27245 VDD AND2X1_LOC_109/a_8_24# -0.00fF
C27574 AND2X1_LOC_312/a_8_24# AND2X1_LOC_528/a_8_24# 0.23fF
C27736 AND2X1_LOC_399/a_8_24# AND2X1_LOC_813/a_8_24# 0.23fF
C27743 OR2X1_LOC_597/a_8_216# OR2X1_LOC_536/a_8_216# 0.47fF
C27984 VDD AND2X1_LOC_78/a_8_24# -0.00fF
C28042 OR2X1_LOC_290/a_8_216# OR2X1_LOC_27/a_8_216# 0.47fF
C28133 OR2X1_LOC_516/a_8_216# OR2X1_LOC_442/a_8_216# 0.47fF
C28361 VDD AND2X1_LOC_601/a_8_24# -0.00fF
C29161 VDD AND2X1_LOC_314/a_8_24# -0.00fF
C29489 AND2X1_LOC_229/a_8_24# VDD -0.00fF
C29974 OR2X1_LOC_41/a_8_216# OR2X1_LOC_311/a_8_216# 0.47fF
C30032 VDD AND2X1_LOC_447/a_8_24# -0.00fF
C30286 VDD OR2X1_LOC_183/a_8_216# 0.21fF
C30444 AND2X1_LOC_481/a_8_24# AND2X1_LOC_279/a_8_24# 0.23fF
C30509 VDD OR2X1_LOC_230/a_8_216# 0.21fF
C30720 OR2X1_LOC_680/a_8_216# VDD 0.21fF
C31260 VDD OR2X1_LOC_746/a_8_216# 0.21fF
C31767 VDD AND2X1_LOC_459/a_8_24# -0.00fF
C32171 VDD AND2X1_LOC_196/a_8_24# -0.00fF
C33433 AND2X1_LOC_184/a_8_24# AND2X1_LOC_292/a_8_24# 0.23fF
C35062 VDD AND2X1_LOC_178/a_8_24# -0.00fF
C36439 OR2X1_LOC_670/a_8_216# OR2X1_LOC_823/a_8_216# 0.47fF
C37336 AND2X1_LOC_536/a_8_24# AND2X1_LOC_135/a_8_24# 0.23fF
C37574 VDD OR2X1_LOC_837/a_8_216# 0.21fF
C37910 VDD OR2X1_LOC_13/a_8_216# 0.21fF
C37992 OR2X1_LOC_165/a_8_216# VDD 0.21fF
C38600 VDD OR2X1_LOC_428/a_8_216# 0.21fF
C39357 VDD OR2X1_LOC_667/a_8_216# 0.21fF
C39773 VDD OR2X1_LOC_498/a_8_216# 0.21fF
C40610 VDD OR2X1_LOC_81/a_8_216# 0.21fF
C41001 VDD OR2X1_LOC_616/a_8_216# 0.21fF
C41714 VDD OR2X1_LOC_769/a_8_216# 0.21fF
C42197 VDD OR2X1_LOC_522/a_8_216# 0.21fF
C42473 AND2X1_LOC_280/a_8_24# AND2X1_LOC_258/a_8_24# 0.23fF
C42557 OR2X1_LOC_635/a_8_216# OR2X1_LOC_614/a_8_216# 0.47fF
C43157 VDD OR2X1_LOC_834/a_8_216# 0.21fF
C43245 VDD OR2X1_LOC_757/a_8_216# 0.21fF
C43265 VDD AND2X1_LOC_697/a_8_24# -0.00fF
C43624 VDD OR2X1_LOC_668/a_8_216# 0.21fF
C44318 VDD OR2X1_LOC_532/a_8_216# 0.21fF
C44531 VDD OR2X1_LOC_836/a_8_216# 0.21fF
C44930 VDD AND2X1_LOC_633/a_8_24# -0.00fF
C45129 OR2X1_LOC_416/a_8_216# OR2X1_LOC_58/a_8_216# 0.47fF
C45167 VDD OR2X1_LOC_521/a_8_216# 0.21fF
C45383 VDD OR2X1_LOC_497/a_8_216# 0.21fF
C45832 VDD OR2X1_LOC_627/a_8_216# 0.21fF
C46049 AND2X1_LOC_187/a_8_24# AND2X1_LOC_441/a_8_24# 0.23fF
C46703 VDD OR2X1_LOC_595/a_8_216# 0.21fF
C46808 VDD OR2X1_LOC_431/a_8_216# 0.21fF
C46836 OR2X1_LOC_838/a_8_216# OR2X1_LOC_20/a_8_216# 0.47fF
C47123 OR2X1_LOC_538/a_8_216# VDD 0.21fF
C47904 AND2X1_LOC_383/a_8_24# VDD -0.00fF
C48097 VDD OR2X1_LOC_89/a_8_216# 0.21fF
C48431 VDD AND2X1_LOC_436/a_8_24# -0.00fF
C48885 VDD OR2X1_LOC_67/a_8_216# 0.21fF
C48897 OR2X1_LOC_305/a_8_216# VDD 0.21fF
C49034 VDD OR2X1_LOC_437/a_8_216# 0.21fF
C49262 AND2X1_LOC_177/a_8_24# AND2X1_LOC_437/a_8_24# 0.23fF
C49620 OR2X1_LOC_118/a_8_216# OR2X1_LOC_131/a_8_216# 0.47fF
C50503 OR2X1_LOC_302/a_8_216# VDD 0.21fF
C50535 AND2X1_LOC_531/a_8_24# VDD -0.00fF
C50605 VDD OR2X1_LOC_99/a_8_216# 0.21fF
C50942 OR2X1_LOC_114/a_8_216# VDD 0.21fF
C51314 OR2X1_LOC_368/a_8_216# VDD 0.21fF
C51349 VDD OR2X1_LOC_778/a_8_216# 0.21fF
C51379 VDD AND2X1_LOC_503/a_8_24# -0.00fF
C51619 VDD OR2X1_LOC_151/a_8_216# 0.21fF
C51793 VDD AND2X1_LOC_52/a_8_24# -0.00fF
C52858 VDD AND2X1_LOC_418/a_8_24# -0.00fF
C53092 VDD OR2X1_LOC_531/a_8_216# 0.21fF
C54274 AND2X1_LOC_297/a_8_24# AND2X1_LOC_248/a_8_24# 0.23fF
C54313 VDD OR2X1_LOC_281/a_8_216# 0.21fF
C54730 VDD OR2X1_LOC_485/a_8_216# 0.21fF
C54798 AND2X1_LOC_385/a_8_24# VDD -0.00fF
C55190 OR2X1_LOC_316/a_8_216# OR2X1_LOC_60/a_8_216# 0.47fF
C55220 VDD OR2X1_LOC_767/a_8_216# 0.21fF
C55324 AND2X1_LOC_482/a_8_24# AND2X1_LOC_252/a_8_24# 0.23fF
C55599 OR2X1_LOC_103/a_8_216# VDD 0.21fF
C56032 VDD AND2X1_LOC_424/a_8_24# -0.00fF
C56427 AND2X1_LOC_406/a_8_24# VSS 0.10fF
C56468 AND2X1_LOC_438/a_8_24# VSS 0.10fF
C56521 AND2X1_LOC_459/a_8_24# VSS 0.10fF
C56529 AND2X1_LOC_607/a_8_24# VSS 0.10fF
C56596 AND2X1_LOC_298/a_8_24# VSS 0.10fF
C56599 AND2X1_LOC_254/a_8_24# VSS 0.10fF
C56604 AND2X1_LOC_265/a_8_24# VSS 0.10fF
C56631 AND2X1_LOC_457/a_8_24# VSS 0.10fF
C56642 AND2X1_LOC_627/a_8_24# VSS 0.10fF
C56675 AND2X1_LOC_434/a_8_24# VSS 0.10fF
C56689 AND2X1_LOC_637/a_8_24# VSS 0.10fF
C56692 AND2X1_LOC_604/a_8_24# VSS 0.10fF
C56698 AND2X1_LOC_829/a_8_24# VSS 0.10fF
C56717 AND2X1_LOC_285/a_8_24# VSS 0.10fF
C56793 AND2X1_LOC_487/a_8_24# VSS 0.10fF
C56796 AND2X1_LOC_498/a_8_24# VSS 0.10fF
C56804 AND2X1_LOC_635/a_8_24# VSS 0.10fF
C56850 AND2X1_LOC_431/a_8_24# VSS 0.10fF
C56868 AND2X1_LOC_667/a_8_24# VSS 0.10fF
C56888 AND2X1_LOC_260/a_8_24# VSS 0.10fF
C56907 AND2X1_LOC_485/a_8_24# VSS 0.10fF
C56910 AND2X1_LOC_677/a_8_24# VSS 0.10fF
C56923 AND2X1_LOC_633/a_8_24# VSS 0.10fF
C56964 AND2X1_LOC_698/a_8_24# VSS 0.10fF
C56968 AND2X1_LOC_665/a_8_24# VSS 0.10fF
C57018 AND2X1_LOC_108/a_8_24# VSS 0.10fF
C57022 AND2X1_LOC_834/a_8_24# VSS 0.10fF
C57031 AND2X1_LOC_823/a_8_24# VSS 0.10fF
C57037 AND2X1_LOC_290/a_8_24# VSS 0.10fF
C57045 AND2X1_LOC_460/a_8_24# VSS 0.10fF
C57080 AND2X1_LOC_118/a_8_24# VSS 0.10fF
C57088 AND2X1_LOC_822/a_8_24# VSS 0.10fF
C57172 AND2X1_LOC_105/a_8_24# VSS 0.10fF
C57249 AND2X1_LOC_307/a_8_24# VSS 0.10fF
C57270 AND2X1_LOC_670/a_8_24# VSS 0.10fF
C57281 AND2X1_LOC_114/a_8_24# VSS 0.10fF
C57287 AND2X1_LOC_79/a_8_24# VSS 0.10fF
C57292 AND2X1_LOC_13/a_8_24# VSS 0.10fF
C57297 AND2X1_LOC_24/a_8_24# VSS 0.10fF
C57326 AND2X1_LOC_179/a_8_24# VSS 0.10fF
C57343 AND2X1_LOC_78/a_8_24# VSS 0.10fF
C57345 AND2X1_LOC_89/a_8_24# VSS 0.10fF
C57352 AND2X1_LOC_305/a_8_24# VSS 0.10fF
C57431 AND2X1_LOC_518/a_8_24# VSS 0.10fF
C57447 AND2X1_LOC_166/a_8_24# VSS 0.10fF
C57448 AND2X1_LOC_122/a_8_24# VSS 0.10fF
C57478 AND2X1_LOC_325/a_8_24# VSS 0.10fF
C57492 AND2X1_LOC_517/a_8_24# VSS 0.10fF
C57507 AND2X1_LOC_154/a_8_24# VSS 0.10fF
C57513 AND2X1_LOC_176/a_8_24# VSS 0.10fF
C57526 AND2X1_LOC_97/a_8_24# VSS 0.10fF
C57534 AND2X1_LOC_75/a_8_24# VSS 0.10fF
C57539 AND2X1_LOC_313/a_8_24# VSS 0.10fF
C57544 AND2X1_LOC_302/a_8_24# VSS 0.10fF
C57554 AND2X1_LOC_538/a_8_24# VSS 0.10fF
C57591 AND2X1_LOC_74/a_8_24# VSS 0.10fF
C57613 AND2X1_LOC_301/a_8_24# VSS 0.10fF
C57639 AND2X1_LOC_196/a_8_24# VSS 0.10fF
C57685 AND2X1_LOC_503/a_8_24# VSS 0.10fF
C57769 AND2X1_LOC_183/a_8_24# VSS 0.10fF
C57791 AND2X1_LOC_320/a_8_24# VSS 0.10fF
C57810 AND2X1_LOC_589/a_8_24# VSS 0.10fF
C57832 AND2X1_LOC_160/a_8_24# VSS 0.10fF
C57915 AND2X1_LOC_521/a_8_24# VSS 0.10fF
C57968 AND2X1_LOC_756/a_8_24# VSS 0.10fF
C58008 AND2X1_LOC_777/a_8_24# VSS 0.10fF
C58071 AND2X1_LOC_583/a_8_24# VSS 0.10fF
C1792 AND2X1_LOC_729/Y AND2X1_LOC_687/Y 0.01fF
C11456 AND2X1_LOC_706/Y AND2X1_LOC_687/Y 0.17fF
C39806 AND2X1_LOC_707/Y AND2X1_LOC_687/Y 0.82fF
C33853 OR2X1_LOC_687/Y OR2X1_LOC_676/Y 0.07fF
C52946 OR2X1_LOC_687/Y OR2X1_LOC_451/B 0.04fF
C13113 OR2X1_LOC_715/B OR2X1_LOC_687/Y 0.10fF
C19226 OR2X1_LOC_687/Y OR2X1_LOC_196/B 0.65fF
C26204 OR2X1_LOC_687/Y OR2X1_LOC_713/A 0.03fF
C56126 OR2X1_LOC_687/Y OR2X1_LOC_678/Y 0.03fF
C16980 OR2X1_LOC_687/Y OR2X1_LOC_623/B 0.33fF
C12905 OR2X1_LOC_334/a_8_216# OR2X1_LOC_338/A 0.01fF
C14248 AND2X1_LOC_24/a_8_24# OR2X1_LOC_338/A 0.10fF
C27933 AND2X1_LOC_27/a_8_24# OR2X1_LOC_338/A 0.25fF
C38331 OR2X1_LOC_334/B OR2X1_LOC_338/A 0.04fF
C39351 OR2X1_LOC_243/A AND2X1_LOC_232/a_8_24# 0.23fF
C45883 OR2X1_LOC_240/B OR2X1_LOC_243/A 0.05fF
C28582 OR2X1_LOC_462/a_8_216# OR2X1_LOC_472/B 0.01fF
C1636 AND2X1_LOC_798/Y AND2X1_LOC_810/B 0.04fF
C4860 OR2X1_LOC_329/B AND2X1_LOC_810/B 1.53fF
C8719 AND2X1_LOC_802/Y AND2X1_LOC_810/B 0.32fF
C23791 AND2X1_LOC_802/a_8_24# AND2X1_LOC_810/B 0.01fF
C25257 AND2X1_LOC_810/B AND2X1_LOC_809/a_36_24# 0.01fF
C29712 AND2X1_LOC_319/a_8_24# AND2X1_LOC_810/B 0.01fF
C31144 AND2X1_LOC_802/B AND2X1_LOC_810/B 0.02fF
C34466 AND2X1_LOC_798/a_8_24# AND2X1_LOC_810/B 0.03fF
C6377 AND2X1_LOC_473/Y OR2X1_LOC_521/a_8_216# 0.18fF
C11953 AND2X1_LOC_473/Y OR2X1_LOC_521/a_36_216# 0.12fF
C18953 OR2X1_LOC_316/Y AND2X1_LOC_473/Y 0.02fF
C27078 AND2X1_LOC_473/a_8_24# AND2X1_LOC_473/Y 0.02fF
C38326 OR2X1_LOC_329/B AND2X1_LOC_473/Y 1.24fF
C5258 AND2X1_LOC_362/B OR2X1_LOC_666/A 0.84fF
C6087 AND2X1_LOC_362/B OR2X1_LOC_595/A 0.31fF
C22318 AND2X1_LOC_362/B OR2X1_LOC_89/Y 0.01fF
C32075 AND2X1_LOC_362/B OR2X1_LOC_67/A 0.03fF
C34613 AND2X1_LOC_362/B AND2X1_LOC_97/a_8_24# 0.01fF
C42231 OR2X1_LOC_122/a_8_216# AND2X1_LOC_362/B 0.05fF
C42360 AND2X1_LOC_362/B OR2X1_LOC_89/a_8_216# 0.01fF
C44381 AND2X1_LOC_362/B OR2X1_LOC_106/a_8_216# 0.07fF
C15237 OR2X1_LOC_656/B AND2X1_LOC_517/a_8_24# 0.01fF
C21681 OR2X1_LOC_656/B OR2X1_LOC_405/A 0.12fF
C32504 OR2X1_LOC_656/B AND2X1_LOC_265/a_8_24# 0.01fF
C38952 OR2X1_LOC_656/B OR2X1_LOC_264/Y 0.08fF
C47236 OR2X1_LOC_101/a_8_216# OR2X1_LOC_656/B 0.01fF
C3708 AND2X1_LOC_729/Y OR2X1_LOC_167/a_36_216# 0.01fF
C6233 AND2X1_LOC_729/Y OR2X1_LOC_329/B 0.43fF
C11749 AND2X1_LOC_729/Y OR2X1_LOC_312/a_8_216# 0.04fF
C14645 AND2X1_LOC_729/Y OR2X1_LOC_526/a_8_216# 0.01fF
C15260 AND2X1_LOC_729/Y AND2X1_LOC_447/a_8_24# 0.02fF
C16650 AND2X1_LOC_729/Y AND2X1_LOC_678/a_8_24# 0.01fF
C27093 AND2X1_LOC_729/Y OR2X1_LOC_600/a_8_216# 0.04fF
C32693 AND2X1_LOC_729/Y OR2X1_LOC_420/a_8_216# 0.05fF
C37226 AND2X1_LOC_729/Y OR2X1_LOC_677/Y 0.02fF
C38134 AND2X1_LOC_729/Y OR2X1_LOC_591/A 0.01fF
C39823 AND2X1_LOC_729/Y OR2X1_LOC_485/a_8_216# 0.01fF
C43789 AND2X1_LOC_729/Y OR2X1_LOC_420/Y 0.02fF
C45135 AND2X1_LOC_729/Y OR2X1_LOC_601/a_8_216# 0.05fF
C45907 AND2X1_LOC_729/Y AND2X1_LOC_436/B 0.03fF
C49378 AND2X1_LOC_729/Y AND2X1_LOC_147/a_8_24# 0.01fF
C50125 AND2X1_LOC_729/Y AND2X1_LOC_729/a_8_24# 0.02fF
C54250 AND2X1_LOC_729/Y AND2X1_LOC_590/a_8_24# 0.01fF
C54297 AND2X1_LOC_729/Y OR2X1_LOC_167/a_8_216# 0.04fF
C35813 AND2X1_LOC_547/Y AND2X1_LOC_547/a_8_24# 0.01fF
C5717 OR2X1_LOC_329/B AND2X1_LOC_715/A 0.09fF
C15857 OR2X1_LOC_518/a_8_216# AND2X1_LOC_715/A 0.47fF
C29828 AND2X1_LOC_715/A OR2X1_LOC_521/a_8_216# 0.01fF
C42339 AND2X1_LOC_715/A OR2X1_LOC_316/Y 0.02fF
C1025 AND2X1_LOC_520/a_8_24# AND2X1_LOC_339/B 0.19fF
C3840 AND2X1_LOC_339/B OR2X1_LOC_75/a_8_216# 0.01fF
C31959 AND2X1_LOC_332/a_8_24# AND2X1_LOC_339/B 0.01fF
C34941 OR2X1_LOC_518/Y AND2X1_LOC_339/B 0.14fF
C42302 AND2X1_LOC_339/B AND2X1_LOC_138/a_8_24# 0.01fF
C31029 OR2X1_LOC_158/a_8_216# OR2X1_LOC_158/B 0.02fF
C36745 OR2X1_LOC_158/B OR2X1_LOC_158/Y 0.01fF
C42046 OR2X1_LOC_158/a_36_216# OR2X1_LOC_158/B 0.01fF
C47256 VDD OR2X1_LOC_158/B 0.04fF
C47493 OR2X1_LOC_158/B OR2X1_LOC_163/Y 0.22fF
C57385 OR2X1_LOC_158/B VSS 0.15fF
C746 AND2X1_LOC_436/B AND2X1_LOC_436/a_8_24# 0.06fF
C3192 AND2X1_LOC_436/B OR2X1_LOC_589/a_8_216# 0.47fF
C4528 VDD AND2X1_LOC_436/B 0.39fF
C10272 AND2X1_LOC_390/B AND2X1_LOC_436/B 0.46fF
C12412 OR2X1_LOC_311/Y AND2X1_LOC_436/B 0.01fF
C19607 OR2X1_LOC_312/Y AND2X1_LOC_436/B 1.06fF
C24540 AND2X1_LOC_535/Y AND2X1_LOC_436/B -0.00fF
C28003 AND2X1_LOC_841/B AND2X1_LOC_436/B 0.19fF
C28375 OR2X1_LOC_166/Y AND2X1_LOC_436/B 0.02fF
C29631 OR2X1_LOC_329/B AND2X1_LOC_436/B 0.02fF
C39247 AND2X1_LOC_539/Y AND2X1_LOC_436/B 0.10fF
C41161 AND2X1_LOC_355/a_8_24# AND2X1_LOC_436/B 0.04fF
C46864 AND2X1_LOC_356/B AND2X1_LOC_436/B 0.07fF
C54967 OR2X1_LOC_167/Y AND2X1_LOC_436/B 0.41fF
C55584 AND2X1_LOC_706/Y AND2X1_LOC_436/B 0.02fF
C56623 AND2X1_LOC_436/B VSS 0.26fF
C15860 AND2X1_LOC_841/B OR2X1_LOC_589/Y 0.01fF
C41164 AND2X1_LOC_841/B AND2X1_LOC_798/Y 0.03fF
C48419 AND2X1_LOC_841/B AND2X1_LOC_802/Y 0.07fF
C48852 AND2X1_LOC_325/a_8_24# AND2X1_LOC_841/B 0.03fF
C52492 OR2X1_LOC_744/Y AND2X1_LOC_783/B 0.78fF
C35253 AND2X1_LOC_464/Y AND2X1_LOC_464/a_8_24# 0.01fF
C24062 OR2X1_LOC_518/Y AND2X1_LOC_520/Y 0.79fF
C39414 OR2X1_LOC_316/Y AND2X1_LOC_520/Y 0.02fF
C13784 AND2X1_LOC_539/Y OR2X1_LOC_829/A 0.01fF
C17102 OR2X1_LOC_829/A OR2X1_LOC_536/a_8_216# 0.28fF
C18620 OR2X1_LOC_385/Y OR2X1_LOC_829/A 0.06fF
C21924 OR2X1_LOC_536/Y OR2X1_LOC_829/A 0.11fF
C27382 AND2X1_LOC_537/a_8_24# OR2X1_LOC_829/A 0.09fF
C35000 VDD OR2X1_LOC_829/A 0.62fF
C40614 AND2X1_LOC_390/B OR2X1_LOC_829/A 0.12fF
C42849 OR2X1_LOC_311/Y OR2X1_LOC_829/A 0.03fF
C56760 OR2X1_LOC_829/A VSS 0.26fF
C3565 AND2X1_LOC_196/a_8_24# AND2X1_LOC_196/Y 0.01fF
C10972 OR2X1_LOC_484/a_8_216# AND2X1_LOC_840/B 0.27fF
C26248 AND2X1_LOC_776/a_8_24# AND2X1_LOC_840/B 0.10fF
C27143 OR2X1_LOC_329/B AND2X1_LOC_840/B 0.04fF
C27415 AND2X1_LOC_840/B OR2X1_LOC_525/a_8_216# 0.04fF
C45496 OR2X1_LOC_680/A AND2X1_LOC_840/B 0.20fF
C4675 OR2X1_LOC_669/Y AND2X1_LOC_668/a_8_24# 0.01fF
C16188 OR2X1_LOC_669/a_8_216# OR2X1_LOC_669/Y 0.01fF
C55809 OR2X1_LOC_669/A OR2X1_LOC_669/Y 0.01fF
C12802 AND2X1_LOC_342/Y OR2X1_LOC_248/Y 0.17fF
C15639 AND2X1_LOC_98/Y AND2X1_LOC_342/Y 0.03fF
C10291 OR2X1_LOC_609/A AND2X1_LOC_610/a_8_24# 0.01fF
C15750 OR2X1_LOC_609/A OR2X1_LOC_612/B 1.33fF
C57020 OR2X1_LOC_609/A VSS 0.29fF
C34939 OR2X1_LOC_288/A AND2X1_LOC_281/a_8_24# 0.23fF
C4479 AND2X1_LOC_764/a_8_24# OR2X1_LOC_637/Y 0.24fF
C15563 OR2X1_LOC_769/A OR2X1_LOC_637/Y 0.05fF
C42270 VDD OR2X1_LOC_637/Y 0.22fF
C49277 OR2X1_LOC_637/Y OR2X1_LOC_638/a_8_216# 0.18fF
C57243 OR2X1_LOC_637/Y VSS -0.01fF
C39930 AND2X1_LOC_489/Y AND2X1_LOC_557/a_8_24# 0.04fF
C53545 AND2X1_LOC_489/Y OR2X1_LOC_595/A 0.07fF
C50198 AND2X1_LOC_333/a_8_24# AND2X1_LOC_338/A 0.01fF
C20128 OR2X1_LOC_604/a_8_216# AND2X1_LOC_454/A 0.47fF
C53260 OR2X1_LOC_423/a_8_216# AND2X1_LOC_454/A 0.10fF
C1610 AND2X1_LOC_714/B AND2X1_LOC_446/a_8_24# 0.20fF
C11759 AND2X1_LOC_714/B AND2X1_LOC_832/a_8_24# 0.04fF
C46498 AND2X1_LOC_714/B OR2X1_LOC_589/Y 0.14fF
C46711 AND2X1_LOC_714/B OR2X1_LOC_418/Y 0.01fF
C1064 AND2X1_LOC_227/Y OR2X1_LOC_224/Y 0.02fF
C1292 AND2X1_LOC_361/a_8_24# AND2X1_LOC_227/Y 0.01fF
C6900 AND2X1_LOC_227/Y AND2X1_LOC_266/Y 0.09fF
C7728 AND2X1_LOC_227/Y OR2X1_LOC_265/a_8_216# 0.01fF
C11160 OR2X1_LOC_497/a_8_216# AND2X1_LOC_227/Y 0.01fF
C17960 AND2X1_LOC_227/Y AND2X1_LOC_267/a_8_24# 0.01fF
C20375 AND2X1_LOC_227/Y OR2X1_LOC_184/a_8_216# 0.01fF
C21400 OR2X1_LOC_103/a_8_216# AND2X1_LOC_227/Y 0.01fF
C22197 OR2X1_LOC_132/a_8_216# AND2X1_LOC_227/Y 0.01fF
C23386 AND2X1_LOC_227/Y AND2X1_LOC_227/a_8_24# 0.01fF
C23472 OR2X1_LOC_107/a_8_216# AND2X1_LOC_227/Y 0.01fF
C32277 AND2X1_LOC_113/a_8_24# AND2X1_LOC_227/Y 0.01fF
C33511 AND2X1_LOC_227/Y OR2X1_LOC_595/A 0.17fF
C39906 OR2X1_LOC_107/Y AND2X1_LOC_227/Y 0.02fF
C43502 AND2X1_LOC_227/Y OR2X1_LOC_72/a_8_216# 0.03fF
C44130 AND2X1_LOC_541/a_8_24# AND2X1_LOC_227/Y 0.01fF
C47305 AND2X1_LOC_130/a_8_24# AND2X1_LOC_227/Y 0.01fF
C47367 AND2X1_LOC_227/Y OR2X1_LOC_517/A 0.03fF
C50199 OR2X1_LOC_134/a_8_216# AND2X1_LOC_227/Y 0.01fF
C52801 OR2X1_LOC_131/A AND2X1_LOC_227/Y 0.04fF
C54654 AND2X1_LOC_227/Y OR2X1_LOC_72/a_36_216# 0.01fF
C34823 OR2X1_LOC_303/B OR2X1_LOC_301/a_8_216# 0.02fF
C45153 OR2X1_LOC_186/Y OR2X1_LOC_303/B 0.01fF
C39739 OR2X1_LOC_543/a_8_216# OR2X1_LOC_552/A 0.01fF
C47526 OR2X1_LOC_303/A OR2X1_LOC_186/Y 0.04fF
C9185 OR2X1_LOC_450/a_8_216# OR2X1_LOC_450/Y -0.00fF
C36777 OR2X1_LOC_292/a_8_216# AND2X1_LOC_848/Y 0.02fF
C38108 AND2X1_LOC_848/a_8_24# AND2X1_LOC_848/Y 0.01fF
C42384 OR2X1_LOC_292/a_36_216# AND2X1_LOC_848/Y 0.01fF
C47308 OR2X1_LOC_669/A AND2X1_LOC_848/Y 0.20fF
C52361 AND2X1_LOC_848/Y AND2X1_LOC_668/a_8_24# 0.04fF
C5877 OR2X1_LOC_612/B OR2X1_LOC_612/Y 0.01fF
C43568 OR2X1_LOC_612/a_8_216# OR2X1_LOC_612/Y -0.00fF
C4232 AND2X1_LOC_67/a_36_24# AND2X1_LOC_67/Y 0.01fF
C6493 AND2X1_LOC_67/Y OR2X1_LOC_66/Y 0.02fF
C9446 OR2X1_LOC_405/A AND2X1_LOC_67/Y 0.02fF
C12605 AND2X1_LOC_67/Y OR2X1_LOC_130/a_8_216# 0.47fF
C19651 OR2X1_LOC_185/Y AND2X1_LOC_67/Y 0.17fF
C49419 AND2X1_LOC_67/a_8_24# AND2X1_LOC_67/Y 0.03fF
C20926 OR2X1_LOC_186/Y OR2X1_LOC_854/A 0.39fF
C608 OR2X1_LOC_139/A AND2X1_LOC_65/a_8_24# 0.02fF
C28471 OR2X1_LOC_139/A OR2X1_LOC_66/Y 0.01fF
C31234 OR2X1_LOC_405/A OR2X1_LOC_139/A 0.13fF
C36311 OR2X1_LOC_139/A OR2X1_LOC_267/A 0.01fF
C36694 OR2X1_LOC_139/A OR2X1_LOC_267/a_8_216# 0.02fF
C41409 OR2X1_LOC_185/Y OR2X1_LOC_139/A 0.01fF
C9348 OR2X1_LOC_447/Y OR2X1_LOC_779/A 0.03fF
C24936 OR2X1_LOC_447/Y OR2X1_LOC_317/B 0.04fF
C30415 OR2X1_LOC_447/Y OR2X1_LOC_704/a_8_216# 0.42fF
C34908 OR2X1_LOC_447/Y OR2X1_LOC_779/a_8_216# 0.02fF
C40365 OR2X1_LOC_447/Y OR2X1_LOC_779/a_36_216# 0.02fF
C44767 OR2X1_LOC_99/A OR2X1_LOC_99/a_8_216# 0.04fF
C46476 VDD OR2X1_LOC_99/A 0.05fF
C55900 OR2X1_LOC_633/Y OR2X1_LOC_99/A 0.03fF
C56859 OR2X1_LOC_99/A VSS 0.14fF
C8422 OR2X1_LOC_539/a_36_216# OR2X1_LOC_390/A 0.01fF
C13024 OR2X1_LOC_434/a_8_216# OR2X1_LOC_390/A 0.01fF
C17667 OR2X1_LOC_405/A OR2X1_LOC_390/A 0.02fF
C31295 AND2X1_LOC_385/a_8_24# OR2X1_LOC_390/A 0.24fF
C36735 OR2X1_LOC_389/B OR2X1_LOC_390/A 0.02fF
C38543 OR2X1_LOC_434/A OR2X1_LOC_390/A 0.55fF
C49961 OR2X1_LOC_537/a_8_216# OR2X1_LOC_390/A 0.01fF
C53505 OR2X1_LOC_539/a_8_216# OR2X1_LOC_390/A 0.01fF
C25797 OR2X1_LOC_630/a_8_216# OR2X1_LOC_630/Y 0.01fF
C931 OR2X1_LOC_680/A AND2X1_LOC_727/A 0.03fF
C1420 AND2X1_LOC_727/A AND2X1_LOC_802/a_8_24# 0.01fF
C3352 AND2X1_LOC_799/a_8_24# AND2X1_LOC_727/A 0.01fF
C5568 AND2X1_LOC_151/a_8_24# AND2X1_LOC_727/A 0.01fF
C7405 AND2X1_LOC_727/A AND2X1_LOC_319/a_8_24# 0.01fF
C8877 AND2X1_LOC_802/B AND2X1_LOC_727/A 0.01fF
C12222 AND2X1_LOC_798/a_8_24# AND2X1_LOC_727/A 0.01fF
C12562 AND2X1_LOC_727/A OR2X1_LOC_533/A 0.01fF
C14614 AND2X1_LOC_307/Y AND2X1_LOC_727/A 0.01fF
C20140 AND2X1_LOC_308/a_8_24# AND2X1_LOC_727/A 0.01fF
C22607 OR2X1_LOC_484/a_8_216# AND2X1_LOC_727/A 0.01fF
C25553 AND2X1_LOC_532/a_8_24# AND2X1_LOC_727/A 0.01fF
C29134 AND2X1_LOC_727/A OR2X1_LOC_142/a_8_216# 0.01fF
C35290 AND2X1_LOC_727/A AND2X1_LOC_798/Y 0.01fF
C38580 OR2X1_LOC_329/B AND2X1_LOC_727/A 0.03fF
C42401 AND2X1_LOC_727/A AND2X1_LOC_802/Y 0.01fF
C47081 AND2X1_LOC_727/A OR2X1_LOC_152/A 0.09fF
C51127 AND2X1_LOC_727/A OR2X1_LOC_594/a_8_216# 0.01fF
C4194 AND2X1_LOC_712/B AND2X1_LOC_448/a_8_24# 0.02fF
C6334 OR2X1_LOC_697/Y AND2X1_LOC_712/B 0.79fF
C23137 AND2X1_LOC_708/a_8_24# AND2X1_LOC_712/B 0.01fF
C43308 AND2X1_LOC_160/Y AND2X1_LOC_712/B 0.11fF
C51526 OR2X1_LOC_697/a_8_216# AND2X1_LOC_712/B 0.02fF
C9969 OR2X1_LOC_518/a_8_216# AND2X1_LOC_326/B 0.01fF
C10032 AND2X1_LOC_326/B AND2X1_LOC_112/a_8_24# 0.01fF
C21018 OR2X1_LOC_518/Y AND2X1_LOC_326/B -0.00fF
C43076 AND2X1_LOC_520/a_8_24# AND2X1_LOC_326/B 0.01fF
C55999 OR2X1_LOC_329/B AND2X1_LOC_326/B 0.03fF
C325 AND2X1_LOC_168/Y OR2X1_LOC_165/Y 0.80fF
C2537 OR2X1_LOC_165/a_8_216# AND2X1_LOC_168/Y 0.01fF
C11405 AND2X1_LOC_168/Y AND2X1_LOC_168/a_8_24# 0.01fF
C1467 AND2X1_LOC_776/Y AND2X1_LOC_776/a_8_24# 0.09fF
C2336 AND2X1_LOC_776/Y OR2X1_LOC_329/B 0.48fF
C9814 OR2X1_LOC_673/Y AND2X1_LOC_132/a_8_24# 0.01fF
C22628 OR2X1_LOC_673/Y AND2X1_LOC_399/a_8_24# 0.02fF
C36157 OR2X1_LOC_673/Y AND2X1_LOC_813/a_8_24# 0.01fF
C44277 OR2X1_LOC_673/Y AND2X1_LOC_134/a_8_24# 0.01fF
C55774 AND2X1_LOC_394/a_8_24# OR2X1_LOC_673/Y 0.02fF
C499 AND2X1_LOC_706/Y OR2X1_LOC_589/a_36_216# -0.00fF
C8789 AND2X1_LOC_706/Y AND2X1_LOC_832/a_8_24# 0.02fF
C13483 AND2X1_LOC_706/Y OR2X1_LOC_424/a_8_216# 0.03fF
C18982 AND2X1_LOC_706/Y OR2X1_LOC_424/a_36_216# 0.01fF
C38384 AND2X1_LOC_706/Y OR2X1_LOC_432/a_8_216# 0.50fF
C38858 AND2X1_LOC_706/Y OR2X1_LOC_432/Y 0.40fF
C43405 AND2X1_LOC_706/Y OR2X1_LOC_589/Y 0.15fF
C45591 AND2X1_LOC_706/Y OR2X1_LOC_589/a_8_216# 0.04fF
C49072 AND2X1_LOC_706/Y AND2X1_LOC_592/a_8_24# 0.04fF
C50114 AND2X1_LOC_706/Y AND2X1_LOC_435/a_8_24# 0.03fF
C5904 AND2X1_LOC_711/A OR2X1_LOC_295/a_8_216# 0.47fF
C13865 OR2X1_LOC_759/A AND2X1_LOC_711/A 0.42fF
C52113 AND2X1_LOC_711/A OR2X1_LOC_759/a_8_216# 0.01fF
C1640 OR2X1_LOC_517/A OR2X1_LOC_118/Y 0.03fF
C2518 OR2X1_LOC_250/Y OR2X1_LOC_517/A 0.01fF
C4082 OR2X1_LOC_131/A OR2X1_LOC_517/A 0.10fF
C6623 OR2X1_LOC_517/a_8_216# OR2X1_LOC_517/A 0.01fF
C18045 OR2X1_LOC_134/Y OR2X1_LOC_517/A 0.05fF
C25078 OR2X1_LOC_131/Y OR2X1_LOC_517/A 0.01fF
C25474 OR2X1_LOC_251/Y OR2X1_LOC_517/A 0.03fF
C25600 OR2X1_LOC_517/A OR2X1_LOC_67/Y 0.03fF
C28033 OR2X1_LOC_517/A AND2X1_LOC_116/Y 0.03fF
C29567 OR2X1_LOC_132/a_8_216# OR2X1_LOC_517/A 0.03fF
C29679 OR2X1_LOC_117/Y OR2X1_LOC_517/A 0.85fF
C33895 OR2X1_LOC_517/A AND2X1_LOC_139/B 0.04fF
C34724 OR2X1_LOC_517/Y OR2X1_LOC_517/A 0.01fF
C40914 OR2X1_LOC_517/A OR2X1_LOC_595/A 0.25fF
C41553 OR2X1_LOC_517/A AND2X1_LOC_105/a_8_24# 0.09fF
C42775 OR2X1_LOC_251/a_8_216# OR2X1_LOC_517/A 0.01fF
C46222 OR2X1_LOC_132/Y OR2X1_LOC_517/A 0.12fF
C47275 OR2X1_LOC_517/A OR2X1_LOC_106/A 0.58fF
C47653 OR2X1_LOC_250/a_8_216# OR2X1_LOC_517/A 0.01fF
C54700 AND2X1_LOC_130/a_8_24# OR2X1_LOC_517/A 0.04fF
C11114 OR2X1_LOC_755/A AND2X1_LOC_624/A 0.05fF
C19530 OR2X1_LOC_755/A OR2X1_LOC_815/a_8_216# 0.02fF
C20611 OR2X1_LOC_755/A OR2X1_LOC_815/Y 0.01fF
C20825 OR2X1_LOC_759/A OR2X1_LOC_755/A 0.01fF
C25486 OR2X1_LOC_757/A OR2X1_LOC_755/A 0.04fF
C32750 OR2X1_LOC_755/A OR2X1_LOC_665/Y 0.01fF
C34444 OR2X1_LOC_755/A OR2X1_LOC_665/a_8_216# 0.49fF
C37050 OR2X1_LOC_755/A AND2X1_LOC_846/a_8_24# 0.01fF
C45588 OR2X1_LOC_755/A OR2X1_LOC_757/Y 0.09fF
C57588 OR2X1_LOC_755/A VSS 0.20fF
C9489 AND2X1_LOC_78/a_8_24# OR2X1_LOC_79/A 0.09fF
C39746 OR2X1_LOC_79/A OR2X1_LOC_79/a_8_216# 0.47fF
C57342 OR2X1_LOC_79/A VSS -0.10fF
C2747 AND2X1_LOC_624/A OR2X1_LOC_152/A 0.03fF
C4581 AND2X1_LOC_624/A OR2X1_LOC_746/a_8_216# 0.01fF
C7203 AND2X1_LOC_186/a_8_24# AND2X1_LOC_624/A 0.05fF
C8452 OR2X1_LOC_759/A AND2X1_LOC_624/A 0.03fF
C12763 OR2X1_LOC_680/A AND2X1_LOC_624/A 0.08fF
C13145 OR2X1_LOC_757/A AND2X1_LOC_624/A 0.03fF
C14059 OR2X1_LOC_252/Y AND2X1_LOC_624/A 0.09fF
C16881 AND2X1_LOC_624/A AND2X1_LOC_254/a_8_24# 0.02fF
C22223 OR2X1_LOC_665/a_8_216# AND2X1_LOC_624/A 0.06fF
C25429 OR2X1_LOC_677/Y AND2X1_LOC_624/A 0.15fF
C25482 OR2X1_LOC_616/Y AND2X1_LOC_624/A 0.03fF
C37278 OR2X1_LOC_406/a_8_216# AND2X1_LOC_624/A 0.05fF
C41117 AND2X1_LOC_154/a_8_24# AND2X1_LOC_624/A 0.01fF
C41636 AND2X1_LOC_483/a_8_24# AND2X1_LOC_624/A 0.02fF
C42726 AND2X1_LOC_624/A OR2X1_LOC_816/A 0.06fF
C48010 OR2X1_LOC_177/a_8_216# AND2X1_LOC_624/A 0.06fF
C568 OR2X1_LOC_186/Y OR2X1_LOC_355/a_8_216# 0.01fF
C1152 OR2X1_LOC_186/Y OR2X1_LOC_809/a_8_216# 0.01fF
C1958 OR2X1_LOC_186/Y OR2X1_LOC_325/a_8_216# 0.10fF
C2378 OR2X1_LOC_186/Y AND2X1_LOC_167/a_8_24# 0.17fF
C3252 OR2X1_LOC_186/Y OR2X1_LOC_330/Y 0.12fF
C4104 OR2X1_LOC_186/Y OR2X1_LOC_798/a_8_216# -0.00fF
C4489 OR2X1_LOC_186/Y OR2X1_LOC_539/Y 0.05fF
C4772 OR2X1_LOC_186/Y OR2X1_LOC_319/Y 0.02fF
C7998 OR2X1_LOC_186/Y AND2X1_LOC_528/a_8_24# 0.07fF
C8781 OR2X1_LOC_186/Y AND2X1_LOC_331/a_8_24# 0.01fF
C10077 OR2X1_LOC_186/Y OR2X1_LOC_799/a_8_216# 0.01fF
C13338 OR2X1_LOC_186/Y OR2X1_LOC_308/Y 0.15fF
C15135 OR2X1_LOC_186/Y AND2X1_LOC_314/a_8_24# 0.01fF
C15496 OR2X1_LOC_186/Y AND2X1_LOC_311/a_8_24# 0.23fF
C17175 OR2X1_LOC_186/Y OR2X1_LOC_356/A 0.01fF
C18027 OR2X1_LOC_186/Y OR2X1_LOC_715/B 0.19fF
C19042 OR2X1_LOC_186/Y OR2X1_LOC_620/B 0.07fF
C20676 OR2X1_LOC_186/Y OR2X1_LOC_147/B 0.07fF
C20688 OR2X1_LOC_186/Y OR2X1_LOC_317/A 0.01fF
C21074 OR2X1_LOC_186/Y OR2X1_LOC_538/A 1.59fF
C21148 OR2X1_LOC_186/Y OR2X1_LOC_802/A 0.01fF
C24275 OR2X1_LOC_186/Y OR2X1_LOC_112/B 0.06fF
C24556 OR2X1_LOC_186/Y OR2X1_LOC_574/A 0.03fF
C27028 OR2X1_LOC_186/Y OR2X1_LOC_405/A 0.49fF
C29463 OR2X1_LOC_186/Y AND2X1_LOC_594/a_8_24# 0.11fF
C29572 OR2X1_LOC_186/Y OR2X1_LOC_703/B 0.23fF
C31569 OR2X1_LOC_186/Y OR2X1_LOC_547/a_8_216# 0.08fF
C37153 OR2X1_LOC_186/Y OR2X1_LOC_185/Y 0.06fF
C37534 OR2X1_LOC_186/Y OR2X1_LOC_798/Y 0.01fF
C37903 OR2X1_LOC_186/Y VDD 0.86fF
C40052 OR2X1_LOC_186/Y OR2X1_LOC_840/A 0.05fF
C40554 OR2X1_LOC_186/Y OR2X1_LOC_802/Y 0.01fF
C41236 OR2X1_LOC_186/Y OR2X1_LOC_532/Y 0.04fF
C41395 OR2X1_LOC_186/Y OR2X1_LOC_447/A 0.01fF
C42636 OR2X1_LOC_186/Y OR2X1_LOC_550/A 0.06fF
C43134 OR2X1_LOC_186/Y OR2X1_LOC_802/a_8_216# 0.01fF
C43546 OR2X1_LOC_186/Y AND2X1_LOC_312/a_8_24# 0.07fF
C44484 OR2X1_LOC_186/Y OR2X1_LOC_778/Y 0.05fF
C49205 OR2X1_LOC_186/Y OR2X1_LOC_703/A 0.17fF
C49804 OR2X1_LOC_186/Y AND2X1_LOC_680/a_8_24# 0.11fF
C52102 OR2X1_LOC_186/Y OR2X1_LOC_112/a_8_216# 0.14fF
C53102 OR2X1_LOC_186/Y OR2X1_LOC_449/B 0.03fF
C53446 OR2X1_LOC_186/Y OR2X1_LOC_317/a_8_216# 0.01fF
C58076 OR2X1_LOC_186/Y VSS 0.57fF
C8604 OR2X1_LOC_151/Y AND2X1_LOC_152/a_8_24# 0.01fF
C27507 VDD OR2X1_LOC_151/Y 0.04fF
C39231 OR2X1_LOC_151/Y OR2X1_LOC_209/A 0.79fF
C57641 OR2X1_LOC_151/Y VSS 0.08fF
C24 OR2X1_LOC_185/Y OR2X1_LOC_702/A 0.02fF
C1745 OR2X1_LOC_185/Y OR2X1_LOC_643/A 0.05fF
C4079 OR2X1_LOC_185/Y OR2X1_LOC_186/a_8_216# 0.19fF
C6646 OR2X1_LOC_185/Y OR2X1_LOC_362/A 0.06fF
C7005 OR2X1_LOC_185/Y OR2X1_LOC_776/A 0.13fF
C7481 OR2X1_LOC_506/a_8_216# OR2X1_LOC_185/Y 0.09fF
C8610 OR2X1_LOC_185/Y OR2X1_LOC_793/B 0.21fF
C8682 OR2X1_LOC_185/Y OR2X1_LOC_506/B 0.11fF
C14500 OR2X1_LOC_185/Y OR2X1_LOC_809/a_8_216# 0.04fF
C15980 OR2X1_LOC_185/Y AND2X1_LOC_522/a_8_24# 0.28fF
C17829 OR2X1_LOC_185/Y OR2X1_LOC_539/Y 0.07fF
C18544 OR2X1_LOC_506/a_36_216# OR2X1_LOC_185/Y 0.15fF
C18717 OR2X1_LOC_185/Y OR2X1_LOC_493/A 0.14fF
C19093 OR2X1_LOC_185/Y OR2X1_LOC_435/B 0.20fF
C24226 OR2X1_LOC_185/Y AND2X1_LOC_67/a_8_24# 0.03fF
C24620 OR2X1_LOC_185/Y OR2X1_LOC_435/a_8_216# 0.02fF
C26455 OR2X1_LOC_185/Y AND2X1_LOC_109/a_8_24# 0.06fF
C27051 OR2X1_LOC_185/Y AND2X1_LOC_522/a_36_24# 0.06fF
C28535 OR2X1_LOC_185/Y AND2X1_LOC_816/a_8_24# 0.01fF
C29360 OR2X1_LOC_185/Y OR2X1_LOC_473/Y 0.03fF
C29425 OR2X1_LOC_185/Y OR2X1_LOC_241/B 0.22fF
C30042 OR2X1_LOC_185/Y AND2X1_LOC_131/a_8_24# 0.26fF
C30100 OR2X1_LOC_185/Y OR2X1_LOC_435/a_36_216# 0.02fF
C30404 OR2X1_LOC_185/Y OR2X1_LOC_138/a_8_216# 0.01fF
C31037 OR2X1_LOC_185/Y OR2X1_LOC_810/A 0.10fF
C31305 OR2X1_LOC_185/Y OR2X1_LOC_715/B 0.35fF
C34274 OR2X1_LOC_185/Y OR2X1_LOC_538/A 0.34fF
C35143 OR2X1_LOC_185/Y AND2X1_LOC_67/a_36_24# 0.01fF
C37435 OR2X1_LOC_185/Y OR2X1_LOC_112/B 0.03fF
C37758 OR2X1_LOC_185/Y OR2X1_LOC_574/A 0.10fF
C39533 OR2X1_LOC_185/Y OR2X1_LOC_846/A 0.01fF
C39816 OR2X1_LOC_185/Y AND2X1_LOC_311/a_36_24# 0.01fF
C41028 OR2X1_LOC_185/Y AND2X1_LOC_131/a_36_24# 0.06fF
C43552 OR2X1_LOC_185/Y OR2X1_LOC_130/a_8_216# 0.02fF
C43744 OR2X1_LOC_185/Y OR2X1_LOC_194/B 0.01fF
C44021 OR2X1_LOC_185/Y OR2X1_LOC_97/A 0.03fF
C45556 OR2X1_LOC_185/Y OR2X1_LOC_778/A 0.02fF
C46239 OR2X1_LOC_185/Y OR2X1_LOC_361/a_8_216# 0.20fF
C47642 OR2X1_LOC_185/Y OR2X1_LOC_776/Y 0.07fF
C49290 OR2X1_LOC_185/Y OR2X1_LOC_113/B 0.05fF
C52264 OR2X1_LOC_185/Y OR2X1_LOC_676/Y 0.07fF
C53469 OR2X1_LOC_185/Y OR2X1_LOC_115/B 0.05fF
C53700 OR2X1_LOC_185/Y OR2X1_LOC_789/a_8_216# 0.03fF
C54002 OR2X1_LOC_185/Y OR2X1_LOC_216/A 0.07fF
C54048 OR2X1_LOC_185/Y OR2X1_LOC_802/Y 0.01fF
C54687 OR2X1_LOC_185/Y OR2X1_LOC_130/Y 0.09fF
C10937 OR2X1_LOC_114/B OR2X1_LOC_664/Y 0.03fF
C12322 OR2X1_LOC_664/Y OR2X1_LOC_833/B 0.08fF
C27925 VDD OR2X1_LOC_664/Y 0.22fF
C28868 OR2X1_LOC_664/Y OR2X1_LOC_483/a_8_216# 0.44fF
C31503 OR2X1_LOC_664/Y AND2X1_LOC_108/a_8_24# 0.02fF
C37693 OR2X1_LOC_664/a_8_216# OR2X1_LOC_664/Y 0.05fF
C48203 OR2X1_LOC_664/Y OR2X1_LOC_346/B 1.29fF
C57646 OR2X1_LOC_664/Y VSS 0.30fF
C55218 OR2X1_LOC_243/B AND2X1_LOC_235/a_8_24# 0.01fF
C19315 OR2X1_LOC_325/a_8_216# OR2X1_LOC_532/Y 0.03fF
C34443 OR2X1_LOC_532/Y OR2X1_LOC_356/A 0.05fF
C43036 OR2X1_LOC_325/Y OR2X1_LOC_532/Y 0.02fF
C44538 OR2X1_LOC_532/Y OR2X1_LOC_330/a_8_216# 0.40fF
C55456 VDD OR2X1_LOC_532/Y 0.20fF
C56483 OR2X1_LOC_532/Y VSS -0.29fF
C23827 AND2X1_LOC_380/a_8_24# OR2X1_LOC_460/B 0.01fF
C34825 OR2X1_LOC_460/B OR2X1_LOC_460/a_8_216# 0.47fF
C58056 OR2X1_LOC_460/B VSS 0.16fF
C3891 OR2X1_LOC_590/Y OR2X1_LOC_593/B 0.01fF
C47863 VDD OR2X1_LOC_590/Y 0.15fF
C49019 OR2X1_LOC_590/Y AND2X1_LOC_591/a_8_24# 0.23fF
C56298 OR2X1_LOC_590/Y VSS 0.04fF
C2045 OR2X1_LOC_188/Y OR2X1_LOC_76/A 0.04fF
C8315 OR2X1_LOC_188/Y OR2X1_LOC_190/A 1.02fF
C8566 OR2X1_LOC_188/Y OR2X1_LOC_241/B 0.03fF
C13014 OR2X1_LOC_188/Y OR2X1_LOC_147/B 0.03fF
C13245 OR2X1_LOC_188/Y OR2X1_LOC_318/B 0.03fF
C21627 OR2X1_LOC_188/Y AND2X1_LOC_666/a_8_24# 0.01fF
C27097 OR2X1_LOC_188/Y OR2X1_LOC_719/A 0.31fF
C29526 OR2X1_LOC_188/Y OR2X1_LOC_76/B 0.02fF
C30320 OR2X1_LOC_188/Y VDD 0.49fF
C32916 OR2X1_LOC_188/Y OR2X1_LOC_457/B 0.22fF
C34140 OR2X1_LOC_188/Y OR2X1_LOC_190/B 0.10fF
C37483 OR2X1_LOC_188/Y OR2X1_LOC_542/B 0.03fF
C38003 OR2X1_LOC_188/Y AND2X1_LOC_183/a_8_24# 0.01fF
C47560 OR2X1_LOC_188/Y OR2X1_LOC_541/a_8_216# 0.01fF
C49996 OR2X1_LOC_188/Y OR2X1_LOC_121/A 0.01fF
C50470 OR2X1_LOC_188/Y AND2X1_LOC_368/a_8_24# 0.01fF
C51848 OR2X1_LOC_188/Y OR2X1_LOC_675/A 0.02fF
C52682 OR2X1_LOC_188/Y AND2X1_LOC_75/a_8_24# 0.01fF
C53652 OR2X1_LOC_188/Y AND2X1_LOC_237/a_8_24# 0.01fF
C58054 OR2X1_LOC_188/Y VSS -0.47fF
C3118 OR2X1_LOC_267/A OR2X1_LOC_720/B 0.03fF
C46291 VDD OR2X1_LOC_267/A 0.08fF
C51855 OR2X1_LOC_267/A OR2X1_LOC_641/A 0.04fF
C57143 OR2X1_LOC_267/A VSS 0.11fF
C45874 OR2X1_LOC_640/A AND2X1_LOC_89/a_8_24# 0.08fF
C15345 AND2X1_LOC_666/a_8_24# OR2X1_LOC_553/A 0.25fF
C26766 OR2X1_LOC_457/B OR2X1_LOC_553/A 0.01fF
C31852 AND2X1_LOC_183/a_8_24# OR2X1_LOC_553/A 0.03fF
C43577 OR2X1_LOC_553/A OR2X1_LOC_121/A 0.01fF
C44106 AND2X1_LOC_368/a_8_24# OR2X1_LOC_553/A 0.04fF
C46466 AND2X1_LOC_75/a_8_24# OR2X1_LOC_553/A 0.04fF
C47434 OR2X1_LOC_553/A AND2X1_LOC_237/a_8_24# 0.07fF
C49980 OR2X1_LOC_270/Y OR2X1_LOC_553/A 0.07fF
C25405 OR2X1_LOC_633/Y OR2X1_LOC_633/a_8_216# 0.01fF
C33125 OR2X1_LOC_633/Y OR2X1_LOC_97/a_8_216# 0.04fF
C41079 OR2X1_LOC_633/Y OR2X1_LOC_610/a_8_216# 0.03fF
C52323 OR2X1_LOC_633/Y OR2X1_LOC_610/a_36_216# 0.02fF
C1080 OR2X1_LOC_777/a_8_216# OR2X1_LOC_784/B -0.00fF
C1748 AND2X1_LOC_390/B OR2X1_LOC_829/a_8_216# 0.04fF
C5489 AND2X1_LOC_390/B OR2X1_LOC_586/Y 0.79fF
C12816 AND2X1_LOC_390/B OR2X1_LOC_829/a_36_216# 0.01fF
C14446 OR2X1_LOC_166/a_8_216# AND2X1_LOC_390/B 0.03fF
C15028 AND2X1_LOC_390/B AND2X1_LOC_539/a_8_24# 0.03fF
C19985 OR2X1_LOC_166/a_36_216# AND2X1_LOC_390/B 0.01fF
C20563 AND2X1_LOC_390/B AND2X1_LOC_538/a_8_24# 0.03fF
C24237 AND2X1_LOC_535/a_8_24# AND2X1_LOC_390/B 0.02fF
C26731 OR2X1_LOC_329/B AND2X1_LOC_390/B 0.07fF
C28563 AND2X1_LOC_390/B OR2X1_LOC_829/Y 0.03fF
C30454 AND2X1_LOC_390/B AND2X1_LOC_802/Y 0.01fF
C34038 AND2X1_LOC_390/B AND2X1_LOC_855/a_8_24# 0.04fF
C35945 AND2X1_LOC_390/B AND2X1_LOC_809/a_8_24# 0.01fF
C38219 AND2X1_LOC_355/a_8_24# AND2X1_LOC_390/B 0.01fF
C41208 OR2X1_LOC_385/Y AND2X1_LOC_390/B 0.01fF
C43685 AND2X1_LOC_390/B OR2X1_LOC_13/a_8_216# 0.03fF
C49347 AND2X1_LOC_390/B OR2X1_LOC_13/a_36_216# 0.01fF
C54020 AND2X1_LOC_390/B AND2X1_LOC_436/a_8_24# 0.02fF
C18806 AND2X1_LOC_355/a_8_24# AND2X1_LOC_356/B 0.01fF
C3563 AND2X1_LOC_307/Y AND2X1_LOC_308/a_8_24# 0.01fF
C4727 OR2X1_LOC_305/Y AND2X1_LOC_307/Y 0.91fF
C12024 AND2X1_LOC_307/a_8_24# AND2X1_LOC_307/Y 0.01fF
C34709 OR2X1_LOC_135/Y AND2X1_LOC_307/Y 0.19fF
C49928 OR2X1_LOC_305/a_8_216# AND2X1_LOC_307/Y 0.03fF
C53187 VDD AND2X1_LOC_307/Y 0.04fF
C57194 AND2X1_LOC_307/Y VSS 0.07fF
C21309 AND2X1_LOC_197/a_8_24# AND2X1_LOC_197/Y 0.01fF
C35491 AND2X1_LOC_197/Y AND2X1_LOC_198/a_8_24# 0.01fF
C40942 VDD AND2X1_LOC_197/Y 0.02fF
C41005 AND2X1_LOC_197/Y AND2X1_LOC_208/B 0.83fF
C57509 AND2X1_LOC_197/Y VSS 0.08fF
C2248 OR2X1_LOC_680/A OR2X1_LOC_504/Y 0.03fF
C28824 OR2X1_LOC_505/a_8_216# OR2X1_LOC_504/Y 0.01fF
C3939 OR2X1_LOC_745/a_8_216# OR2X1_LOC_746/Y 0.39fF
C8049 AND2X1_LOC_709/a_8_24# OR2X1_LOC_258/Y 0.24fF
C9931 OR2X1_LOC_295/a_8_216# OR2X1_LOC_258/Y 0.01fF
C17768 OR2X1_LOC_759/A OR2X1_LOC_258/Y 0.03fF
C17817 OR2X1_LOC_698/Y OR2X1_LOC_258/Y 0.23fF
C9245 OR2X1_LOC_232/Y AND2X1_LOC_240/a_8_24# 0.23fF
C22406 VDD OR2X1_LOC_232/Y 0.12fF
C56773 OR2X1_LOC_232/Y VSS 0.06fF
C36660 OR2X1_LOC_177/a_8_216# OR2X1_LOC_438/Y 0.40fF
C27630 OR2X1_LOC_189/A OR2X1_LOC_498/Y 0.01fF
C39572 OR2X1_LOC_680/A OR2X1_LOC_674/Y 0.03fF
C17403 OR2X1_LOC_118/Y AND2X1_LOC_266/Y 0.81fF
C18572 OR2X1_LOC_118/Y OR2X1_LOC_131/a_8_216# 0.01fF
C35427 OR2X1_LOC_118/a_8_216# OR2X1_LOC_118/Y 0.01fF
C38392 OR2X1_LOC_118/Y AND2X1_LOC_249/a_8_24# 0.01fF
C43700 OR2X1_LOC_118/Y AND2X1_LOC_266/a_8_24# 0.01fF
C44015 OR2X1_LOC_118/Y OR2X1_LOC_595/A 0.03fF
C36626 OR2X1_LOC_821/Y OR2X1_LOC_822/a_8_216# 0.03fF
C37059 OR2X1_LOC_821/Y OR2X1_LOC_813/a_8_216# 0.03fF
C16866 OR2X1_LOC_177/Y OR2X1_LOC_680/A 0.03fF
C39707 OR2X1_LOC_177/Y OR2X1_LOC_109/a_8_216# 0.01fF
C31545 OR2X1_LOC_595/A OR2X1_LOC_767/Y 0.05fF
C9295 OR2X1_LOC_751/Y AND2X1_LOC_789/a_8_24# 0.01fF
C27870 OR2X1_LOC_751/Y VDD 0.06fF
C37035 OR2X1_LOC_751/Y AND2X1_LOC_789/Y 0.81fF
C57966 OR2X1_LOC_751/Y VSS 0.10fF
C16623 OR2X1_LOC_815/a_8_216# OR2X1_LOC_815/Y -0.00fF
C17901 OR2X1_LOC_759/A OR2X1_LOC_815/Y 0.02fF
C34188 OR2X1_LOC_815/Y AND2X1_LOC_846/a_8_24# 0.23fF
C34861 VDD OR2X1_LOC_815/Y 0.12fF
C38660 OR2X1_LOC_816/Y OR2X1_LOC_815/Y 0.08fF
C56982 OR2X1_LOC_815/Y VSS -0.03fF
C7302 OR2X1_LOC_665/Y AND2X1_LOC_483/a_8_24# 0.03fF
C8432 OR2X1_LOC_665/Y OR2X1_LOC_816/A 0.03fF
C18386 OR2X1_LOC_665/Y AND2X1_LOC_483/a_36_24# 0.01fF
C30082 OR2X1_LOC_759/A OR2X1_LOC_665/Y 0.16fF
C32998 OR2X1_LOC_665/Y OR2X1_LOC_253/Y 0.06fF
C34732 OR2X1_LOC_757/A OR2X1_LOC_665/Y 0.01fF
C38486 OR2X1_LOC_665/Y AND2X1_LOC_254/a_8_24# 0.04fF
C49531 OR2X1_LOC_665/a_36_216# OR2X1_LOC_665/Y 0.01fF
C55257 OR2X1_LOC_665/Y AND2X1_LOC_254/a_36_24# 0.01fF
C22921 AND2X1_LOC_333/a_8_24# OR2X1_LOC_171/Y 0.01fF
C41280 AND2X1_LOC_348/A OR2X1_LOC_384/Y 0.01fF
C42127 VDD OR2X1_LOC_384/Y 0.19fF
C56477 OR2X1_LOC_384/Y VSS 0.25fF
C18948 VDD OR2X1_LOC_531/Y 0.12fF
C53067 OR2X1_LOC_531/Y AND2X1_LOC_549/a_8_24# 0.23fF
C57559 OR2X1_LOC_531/Y VSS 0.06fF
C14949 OR2X1_LOC_41/Y OR2X1_LOC_13/Y 0.13fF
C17911 VDD OR2X1_LOC_41/Y 0.21fF
C23276 OR2X1_LOC_41/a_8_216# OR2X1_LOC_41/Y 0.01fF
C56976 OR2X1_LOC_41/Y VSS 0.39fF
C19150 OR2X1_LOC_265/Y AND2X1_LOC_266/Y 0.55fF
C19968 OR2X1_LOC_265/a_8_216# OR2X1_LOC_265/Y 0.01fF
C30161 OR2X1_LOC_265/Y AND2X1_LOC_267/a_8_24# 0.25fF
C35614 OR2X1_LOC_316/Y OR2X1_LOC_265/Y 0.03fF
C55872 OR2X1_LOC_72/a_8_216# OR2X1_LOC_265/Y 0.03fF
C2022 OR2X1_LOC_441/a_8_216# OR2X1_LOC_441/Y 0.01fF
C4526 OR2X1_LOC_677/Y OR2X1_LOC_441/Y 0.03fF
C16452 OR2X1_LOC_441/Y AND2X1_LOC_147/a_8_24# 0.07fF
C37841 OR2X1_LOC_441/Y OR2X1_LOC_152/A 0.03fF
C39748 OR2X1_LOC_441/Y OR2X1_LOC_746/a_8_216# 0.06fF
C49730 OR2X1_LOC_677/a_8_216# OR2X1_LOC_441/Y 0.06fF
C15970 OR2X1_LOC_166/Y AND2X1_LOC_436/a_8_24# 0.01fF
C32468 OR2X1_LOC_166/a_8_216# OR2X1_LOC_166/Y 0.01fF
C7074 AND2X1_LOC_707/Y OR2X1_LOC_423/a_8_216# 0.03fF
C12626 AND2X1_LOC_707/Y OR2X1_LOC_423/a_36_216# 0.01fF
C54550 AND2X1_LOC_450/a_8_24# AND2X1_LOC_450/Y 0.01fF
C2050 OR2X1_LOC_506/B AND2X1_LOC_239/a_8_24# 0.01fF
C21675 OR2X1_LOC_506/a_8_216# OR2X1_LOC_506/B 0.03fF
C1947 OR2X1_LOC_621/A AND2X1_LOC_616/a_36_24# 0.01fF
C3807 OR2X1_LOC_621/A AND2X1_LOC_670/a_36_24# 0.01fF
C5689 VDD OR2X1_LOC_621/A 0.21fF
C8898 OR2X1_LOC_621/A OR2X1_LOC_624/B 0.01fF
C21051 OR2X1_LOC_621/A OR2X1_LOC_621/B 0.62fF
C31985 OR2X1_LOC_621/A OR2X1_LOC_621/a_8_216# 0.01fF
C35844 OR2X1_LOC_621/A AND2X1_LOC_616/a_8_24# 0.21fF
C40456 OR2X1_LOC_673/B OR2X1_LOC_621/A 0.02fF
C48942 OR2X1_LOC_621/A AND2X1_LOC_670/a_8_24# 0.11fF
C57587 OR2X1_LOC_621/A VSS -0.06fF
C22488 OR2X1_LOC_843/a_8_216# OR2X1_LOC_843/B 0.02fF
C32198 AND2X1_LOC_250/a_8_24# OR2X1_LOC_843/B 0.20fF
C44016 OR2X1_LOC_249/Y OR2X1_LOC_843/B 0.35fF
C8180 OR2X1_LOC_846/a_8_216# OR2X1_LOC_846/A 0.14fF
C19215 OR2X1_LOC_846/a_36_216# OR2X1_LOC_846/A 0.01fF
C40234 VDD OR2X1_LOC_846/A 0.01fF
C43014 OR2X1_LOC_846/B OR2X1_LOC_846/A 0.52fF
C48390 OR2X1_LOC_846/A OR2X1_LOC_561/B 0.26fF
C56823 OR2X1_LOC_846/A VSS 0.11fF
C31580 OR2X1_LOC_405/A OR2X1_LOC_728/A 0.03fF
C11493 AND2X1_LOC_145/a_8_24# OR2X1_LOC_148/B 0.01fF
C28858 VDD OR2X1_LOC_168/A -0.00fF
C31047 OR2X1_LOC_840/A OR2X1_LOC_168/A 0.05fF
C34863 OR2X1_LOC_168/a_8_216# OR2X1_LOC_168/A 0.47fF
C43866 OR2X1_LOC_168/A OR2X1_LOC_449/B 0.04fF
C57512 OR2X1_LOC_168/A VSS 0.15fF
C26940 OR2X1_LOC_467/B OR2X1_LOC_160/Y 0.03fF
C147 OR2X1_LOC_97/A OR2X1_LOC_832/a_8_216# 0.01fF
C9958 OR2X1_LOC_97/A AND2X1_LOC_60/a_8_24# 0.01fF
C11241 OR2X1_LOC_97/A AND2X1_LOC_172/a_8_24# 0.01fF
C20000 OR2X1_LOC_97/A AND2X1_LOC_109/a_8_24# 0.01fF
C21110 OR2X1_LOC_97/A AND2X1_LOC_601/a_8_24# 0.01fF
C23582 OR2X1_LOC_97/A AND2X1_LOC_438/a_8_24# 0.02fF
C26473 AND2X1_LOC_91/a_8_24# OR2X1_LOC_97/A 0.01fF
C29563 OR2X1_LOC_97/A AND2X1_LOC_32/a_8_24# 0.01fF
C31633 OR2X1_LOC_97/A AND2X1_LOC_58/a_8_24# 0.01fF
C33761 OR2X1_LOC_405/A OR2X1_LOC_97/A 0.03fF
C37540 OR2X1_LOC_97/A AND2X1_LOC_290/a_8_24# 0.01fF
C39638 OR2X1_LOC_97/A AND2X1_LOC_20/a_8_24# 0.01fF
C40638 OR2X1_LOC_97/A AND2X1_LOC_600/a_8_24# 0.01fF
C44243 OR2X1_LOC_97/A AND2X1_LOC_432/a_8_24# 0.01fF
C45266 OR2X1_LOC_97/A OR2X1_LOC_334/B 0.01fF
C50905 OR2X1_LOC_97/A OR2X1_LOC_634/a_8_216# 0.01fF
C2515 OR2X1_LOC_227/a_8_216# OR2X1_LOC_227/B 0.01fF
C5182 AND2X1_LOC_224/a_8_24# OR2X1_LOC_227/B 0.02fF
C11663 OR2X1_LOC_641/A OR2X1_LOC_227/B 0.08fF
C56460 OR2X1_LOC_227/B VSS 0.17fF
C10976 OR2X1_LOC_302/B AND2X1_LOC_298/a_8_24# 0.02fF
C27477 OR2X1_LOC_302/B OR2X1_LOC_147/B 0.14fF
C44854 OR2X1_LOC_302/B VDD 0.21fF
C58108 OR2X1_LOC_302/B VSS 0.11fF
C1421 OR2X1_LOC_809/a_8_216# OR2X1_LOC_112/B 0.02fF
C5991 OR2X1_LOC_435/B OR2X1_LOC_112/B 0.04fF
C6916 OR2X1_LOC_809/a_36_216# OR2X1_LOC_112/B 0.03fF
C11571 OR2X1_LOC_435/a_8_216# OR2X1_LOC_112/B 0.15fF
C27299 OR2X1_LOC_405/A OR2X1_LOC_112/B 0.03fF
C40804 OR2X1_LOC_802/Y OR2X1_LOC_112/B 0.06fF
C42622 OR2X1_LOC_435/Y OR2X1_LOC_112/B 0.10fF
C52384 OR2X1_LOC_112/a_8_216# OR2X1_LOC_112/B 0.01fF
C27478 OR2X1_LOC_405/A OR2X1_LOC_493/B 0.02fF
C42451 OR2X1_LOC_493/B AND2X1_LOC_491/a_8_24# 0.01fF
C52300 OR2X1_LOC_264/Y OR2X1_LOC_559/B 0.01fF
C9074 AND2X1_LOC_142/a_36_24# OR2X1_LOC_705/B 0.01fF
C37477 AND2X1_LOC_525/a_8_24# OR2X1_LOC_705/B 0.10fF
C48338 OR2X1_LOC_147/a_8_216# OR2X1_LOC_705/B 0.01fF
C54152 AND2X1_LOC_142/a_8_24# OR2X1_LOC_705/B 0.01fF
C26150 OR2X1_LOC_791/A OR2X1_LOC_756/a_8_216# 0.47fF
C44110 OR2X1_LOC_791/A OR2X1_LOC_260/Y 0.02fF
C49304 OR2X1_LOC_756/Y OR2X1_LOC_791/A 0.01fF
C5065 VDD OR2X1_LOC_780/A 0.21fF
C9023 OR2X1_LOC_780/A AND2X1_LOC_424/a_8_24# 0.20fF
C57041 OR2X1_LOC_780/A VSS 0.15fF
C12593 OR2X1_LOC_128/B OR2X1_LOC_342/A 0.37fF
C31178 OR2X1_LOC_114/B OR2X1_LOC_342/A 0.04fF
C48366 VDD OR2X1_LOC_342/A 0.21fF
C51888 AND2X1_LOC_127/a_8_24# OR2X1_LOC_342/A 0.25fF
C56364 OR2X1_LOC_342/A VSS 0.20fF
C5259 OR2X1_LOC_631/a_8_216# OR2X1_LOC_115/B 0.03fF
C32815 AND2X1_LOC_131/a_8_24# OR2X1_LOC_115/B 0.01fF
C40240 OR2X1_LOC_66/Y OR2X1_LOC_115/B 0.01fF
C43544 OR2X1_LOC_115/a_8_216# OR2X1_LOC_115/B 0.05fF
C20661 AND2X1_LOC_103/a_8_24# OR2X1_LOC_113/B 0.01fF
C53809 OR2X1_LOC_113/a_8_216# OR2X1_LOC_113/B 0.03fF
C7208 OR2X1_LOC_209/A OR2X1_LOC_151/a_8_216# 0.01fF
C21676 AND2X1_LOC_485/a_8_24# OR2X1_LOC_209/A 0.04fF
C38080 AND2X1_LOC_485/a_36_24# OR2X1_LOC_209/A 0.01fF
C44840 AND2X1_LOC_152/a_8_24# OR2X1_LOC_209/A 0.01fF
C11874 OR2X1_LOC_793/A AND2X1_LOC_39/a_8_24# 0.05fF
C42214 OR2X1_LOC_793/A AND2X1_LOC_41/Y 0.01fF
C3986 OR2X1_LOC_639/B AND2X1_LOC_428/a_8_24# 0.25fF
C9540 OR2X1_LOC_639/B OR2X1_LOC_451/B 0.19fF
C11500 AND2X1_LOC_584/a_8_24# OR2X1_LOC_639/B 0.04fF
C15039 OR2X1_LOC_639/B AND2X1_LOC_428/a_36_24# 0.01fF
C35540 AND2X1_LOC_583/a_8_24# OR2X1_LOC_639/B 0.03fF
C38815 AND2X1_LOC_584/a_36_24# OR2X1_LOC_639/B 0.01fF
C46764 AND2X1_LOC_583/a_36_24# OR2X1_LOC_639/B 0.01fF
C11649 OR2X1_LOC_78/Y OR2X1_LOC_771/B 0.03fF
C13412 OR2X1_LOC_379/Y OR2X1_LOC_771/B 0.01fF
C38402 OR2X1_LOC_520/B OR2X1_LOC_771/B 0.60fF
C3129 OR2X1_LOC_427/a_8_216# AND2X1_LOC_451/Y 0.49fF
C3942 OR2X1_LOC_427/Y AND2X1_LOC_451/Y 0.01fF
C9500 AND2X1_LOC_450/a_8_24# AND2X1_LOC_451/Y 0.01fF
C36164 OR2X1_LOC_158/a_8_216# OR2X1_LOC_163/Y 0.40fF
C38240 AND2X1_LOC_161/Y OR2X1_LOC_163/Y 0.02fF
C41440 OR2X1_LOC_163/a_8_216# OR2X1_LOC_163/Y 0.01fF
C43863 AND2X1_LOC_162/a_8_24# OR2X1_LOC_163/Y 0.01fF
C5818 OR2X1_LOC_525/Y OR2X1_LOC_677/Y 0.01fF
C6285 OR2X1_LOC_525/Y AND2X1_LOC_834/a_8_24# 0.02fF
C40505 OR2X1_LOC_680/a_8_216# OR2X1_LOC_525/Y 0.01fF
C49396 OR2X1_LOC_525/Y OR2X1_LOC_680/A 0.02fF
C23900 OR2X1_LOC_495/a_8_216# OR2X1_LOC_238/Y 0.41fF
C52735 AND2X1_LOC_776/a_8_24# OR2X1_LOC_238/Y 0.11fF
C53610 OR2X1_LOC_329/B OR2X1_LOC_238/Y 0.10fF
C39565 OR2X1_LOC_52/a_8_216# OR2X1_LOC_52/Y 0.01fF
C37299 OR2X1_LOC_313/Y OR2X1_LOC_418/Y 0.18fF
C41008 AND2X1_LOC_704/a_8_24# OR2X1_LOC_418/Y 0.24fF
C48911 VDD OR2X1_LOC_418/Y 0.19fF
C56622 OR2X1_LOC_418/Y VSS 0.12fF
C9343 OR2X1_LOC_251/Y AND2X1_LOC_286/a_8_24# 0.01fF
C9440 OR2X1_LOC_251/Y OR2X1_LOC_669/A 0.01fF
C11808 OR2X1_LOC_251/Y OR2X1_LOC_595/A 0.01fF
C12394 OR2X1_LOC_251/Y AND2X1_LOC_105/a_8_24# 0.01fF
C13613 OR2X1_LOC_251/Y OR2X1_LOC_251/a_8_216# 0.08fF
C14503 OR2X1_LOC_251/Y AND2X1_LOC_668/a_8_24# 0.01fF
C17892 OR2X1_LOC_251/Y OR2X1_LOC_106/A 0.03fF
C18287 OR2X1_LOC_251/Y OR2X1_LOC_250/a_8_216# 0.03fF
C23857 OR2X1_LOC_251/Y OR2X1_LOC_250/a_36_216# 0.01fF
C25950 OR2X1_LOC_251/Y OR2X1_LOC_669/a_8_216# 0.01fF
C39492 OR2X1_LOC_251/Y OR2X1_LOC_667/a_8_216# 0.04fF
C44188 OR2X1_LOC_251/Y AND2X1_LOC_287/a_8_24# 0.01fF
C50753 OR2X1_LOC_251/Y OR2X1_LOC_667/a_36_216# 0.02fF
C22435 OR2X1_LOC_698/a_8_216# OR2X1_LOC_816/Y 0.57fF
C38834 OR2X1_LOC_759/A OR2X1_LOC_816/Y 0.02fF
C55994 VDD OR2X1_LOC_816/Y 0.17fF
C57418 OR2X1_LOC_816/Y VSS 0.01fF
C8676 OR2X1_LOC_331/A OR2X1_LOC_533/A 0.15fF
C9628 OR2X1_LOC_331/A VDD 0.03fF
C17646 AND2X1_LOC_330/a_8_24# OR2X1_LOC_331/A 0.02fF
C53132 OR2X1_LOC_331/A OR2X1_LOC_680/A 0.06fF
C54549 OR2X1_LOC_331/A OR2X1_LOC_331/a_8_216# 0.04fF
C57855 OR2X1_LOC_331/A VSS 0.14fF
C2156 OR2X1_LOC_680/Y AND2X1_LOC_147/a_8_24# 0.01fF
C46368 OR2X1_LOC_680/Y OR2X1_LOC_677/Y 0.03fF
C30893 OR2X1_LOC_165/Y AND2X1_LOC_168/a_8_24# 0.01fF
C35888 VDD OR2X1_LOC_165/Y 0.04fF
C43712 OR2X1_LOC_91/Y OR2X1_LOC_165/Y 0.05fF
C47946 AND2X1_LOC_787/A OR2X1_LOC_165/Y 0.21fF
C57324 OR2X1_LOC_165/Y VSS 0.08fF
C28936 OR2X1_LOC_533/Y OR2X1_LOC_533/A 0.04fF
C11408 AND2X1_LOC_532/a_8_24# OR2X1_LOC_594/Y 0.25fF
C13096 OR2X1_LOC_823/a_8_216# OR2X1_LOC_96/Y 0.01fF
C16909 OR2X1_LOC_670/a_8_216# OR2X1_LOC_96/Y 0.01fF
C22845 VDD OR2X1_LOC_96/Y 0.30fF
C53560 OR2X1_LOC_96/Y OR2X1_LOC_670/Y 0.01fF
C57469 OR2X1_LOC_96/Y VSS 0.10fF
C6160 OR2X1_LOC_406/Y OR2X1_LOC_406/a_8_216# 0.01fF
C14433 OR2X1_LOC_617/a_8_216# OR2X1_LOC_626/Y 0.01fF
C21174 OR2X1_LOC_252/a_8_216# OR2X1_LOC_626/Y 0.39fF
C25456 OR2X1_LOC_617/Y OR2X1_LOC_626/Y 0.16fF
C30892 OR2X1_LOC_680/A OR2X1_LOC_626/Y 0.03fF
C31341 OR2X1_LOC_626/a_8_216# OR2X1_LOC_626/Y 0.01fF
C40510 OR2X1_LOC_626/Y OR2X1_LOC_627/Y 0.01fF
C56527 OR2X1_LOC_626/Y VSS 0.20fF
C21672 OR2X1_LOC_487/Y AND2X1_LOC_489/a_8_24# 0.23fF
C42961 OR2X1_LOC_487/a_8_216# OR2X1_LOC_487/Y -0.00fF
C53159 VDD OR2X1_LOC_487/Y 0.12fF
C57380 OR2X1_LOC_487/Y VSS 0.06fF
C1240 OR2X1_LOC_759/A OR2X1_LOC_258/a_8_216# 0.01fF
C3014 OR2X1_LOC_759/A AND2X1_LOC_664/a_8_24# 0.01fF
C8355 OR2X1_LOC_759/A AND2X1_LOC_709/a_8_24# 0.18fF
C12557 AND2X1_LOC_758/a_8_24# OR2X1_LOC_759/A 0.01fF
C16795 OR2X1_LOC_759/A OR2X1_LOC_815/a_8_216# 0.01fF
C16972 OR2X1_LOC_759/A OR2X1_LOC_617/Y 0.03fF
C18117 OR2X1_LOC_759/A OR2X1_LOC_698/Y 0.55fF
C22485 OR2X1_LOC_759/A OR2X1_LOC_680/A 0.03fF
C22860 OR2X1_LOC_757/A OR2X1_LOC_759/A 2.01fF
C31785 OR2X1_LOC_759/A OR2X1_LOC_665/a_8_216# 0.01fF
C34032 OR2X1_LOC_759/A AND2X1_LOC_793/B 0.34fF
C34406 OR2X1_LOC_759/A AND2X1_LOC_846/a_8_24# 0.01fF
C35018 OR2X1_LOC_759/A VDD 0.22fF
C35083 OR2X1_LOC_759/A OR2X1_LOC_616/Y 0.01fF
C44334 OR2X1_LOC_759/A AND2X1_LOC_789/Y 0.02fF
C51307 OR2X1_LOC_528/Y OR2X1_LOC_759/A 0.03fF
C57882 OR2X1_LOC_759/A VSS 0.04fF
C5455 OR2X1_LOC_152/A OR2X1_LOC_142/Y 0.03fF
C13446 AND2X1_LOC_778/a_8_24# OR2X1_LOC_142/Y 0.02fF
C15483 OR2X1_LOC_680/A OR2X1_LOC_142/Y 14.00fF
C17163 OR2X1_LOC_677/a_8_216# OR2X1_LOC_142/Y 0.18fF
C20230 AND2X1_LOC_151/a_8_24# OR2X1_LOC_142/Y 0.01fF
C28208 OR2X1_LOC_677/Y OR2X1_LOC_142/Y 0.02fF
C40005 AND2X1_LOC_147/a_8_24# OR2X1_LOC_142/Y -0.00fF
C1605 AND2X1_LOC_539/Y OR2X1_LOC_829/Y 0.02fF
C22998 VDD OR2X1_LOC_829/Y 0.15fF
C30667 OR2X1_LOC_311/Y OR2X1_LOC_829/Y 0.02fF
C55432 OR2X1_LOC_829/Y AND2X1_LOC_855/a_8_24# 0.23fF
C57086 OR2X1_LOC_829/Y VSS 0.07fF
C46758 OR2X1_LOC_250/Y OR2X1_LOC_251/a_8_216# 0.01fF
C51113 OR2X1_LOC_250/Y OR2X1_LOC_106/A 0.02fF
C18106 VDD OR2X1_LOC_107/Y 0.16fF
C21611 OR2X1_LOC_107/Y OR2X1_LOC_103/Y 0.23fF
C32541 OR2X1_LOC_107/Y AND2X1_LOC_113/a_8_24# 0.23fF
C57720 OR2X1_LOC_107/Y VSS -0.09fF
C41516 AND2X1_LOC_802/B OR2X1_LOC_167/Y 0.02fF
C42500 OR2X1_LOC_167/Y AND2X1_LOC_436/a_8_24# 0.13fF
C50613 OR2X1_LOC_518/Y AND2X1_LOC_831/Y 0.13fF
C54579 OR2X1_LOC_518/Y AND2X1_LOC_520/a_8_24# 0.01fF
C58040 OR2X1_LOC_518/Y VSS 0.10fF
C34313 OR2X1_LOC_313/a_8_216# OR2X1_LOC_314/Y 0.40fF
C40238 OR2X1_LOC_313/Y OR2X1_LOC_314/Y 0.22fF
C51847 VDD OR2X1_LOC_314/Y 0.08fF
C57299 OR2X1_LOC_314/Y VSS 0.22fF
C2709 OR2X1_LOC_462/B OR2X1_LOC_416/a_8_216# 0.02fF
C21652 OR2X1_LOC_462/B OR2X1_LOC_520/a_8_216# 0.01fF
C22236 OR2X1_LOC_462/B AND2X1_LOC_518/a_8_24# 0.01fF
C27686 OR2X1_LOC_462/B OR2X1_LOC_520/B 0.01fF
C29728 OR2X1_LOC_462/B AND2X1_LOC_89/a_8_24# 0.01fF
C30207 OR2X1_LOC_462/B OR2X1_LOC_462/a_8_216# 0.02fF
C35199 OR2X1_LOC_462/B OR2X1_LOC_97/B 0.01fF
C41203 OR2X1_LOC_462/B OR2X1_LOC_462/a_36_216# 0.03fF
C11053 OR2X1_LOC_791/B OR2X1_LOC_285/A 0.01fF
C30202 OR2X1_LOC_285/B OR2X1_LOC_285/A 0.05fF
C56889 OR2X1_LOC_285/A VSS 0.18fF
C11104 AND2X1_LOC_158/a_8_24# OR2X1_LOC_210/B 0.01fF
C27485 OR2X1_LOC_210/B OR2X1_LOC_160/Y 0.05fF
C23807 AND2X1_LOC_178/a_8_24# OR2X1_LOC_181/B 0.02fF
C30883 OR2X1_LOC_181/B AND2X1_LOC_179/a_8_24# 0.02fF
C11781 AND2X1_LOC_498/a_8_24# OR2X1_LOC_499/B 0.09fF
C23427 OR2X1_LOC_499/B AND2X1_LOC_496/a_8_24# 0.01fF
C28344 AND2X1_LOC_498/a_36_24# OR2X1_LOC_499/B -0.00fF
C25993 AND2X1_LOC_145/a_8_24# OR2X1_LOC_148/A 0.22fF
C668 AND2X1_LOC_320/a_8_24# OR2X1_LOC_324/B 0.01fF
C1052 OR2X1_LOC_614/Y OR2X1_LOC_790/A 0.01fF
C7397 OR2X1_LOC_196/Y OR2X1_LOC_790/A 0.16fF
C40654 OR2X1_LOC_790/A AND2X1_LOC_45/a_8_24# 0.05fF
C58044 OR2X1_LOC_790/A VSS 0.28fF
C8874 OR2X1_LOC_405/A OR2X1_LOC_435/B 1.33fF
C55721 OR2X1_LOC_435/B OR2X1_LOC_810/A 0.07fF
C55750 AND2X1_LOC_589/a_8_24# OR2X1_LOC_435/B 0.03fF
C57220 OR2X1_LOC_435/B VSS -0.06fF
C9699 OR2X1_LOC_778/A OR2X1_LOC_121/A 0.02fF
C35214 OR2X1_LOC_405/A OR2X1_LOC_778/A 0.01fF
C45470 OR2X1_LOC_778/A OR2X1_LOC_778/a_8_216# 0.04fF
C15878 OR2X1_LOC_719/A AND2X1_LOC_237/a_8_24# 0.21fF
C29863 AND2X1_LOC_813/a_8_24# AND2X1_LOC_79/Y 0.04fF
C40838 AND2X1_LOC_813/a_36_24# AND2X1_LOC_79/Y 0.01fF
C4325 OR2X1_LOC_147/B OR2X1_LOC_270/Y 0.03fF
C6020 OR2X1_LOC_833/B OR2X1_LOC_270/Y 0.01fF
C6032 OR2X1_LOC_254/B OR2X1_LOC_270/Y 0.01fF
C28914 OR2X1_LOC_542/B OR2X1_LOC_270/Y 0.03fF
C41661 AND2X1_LOC_368/a_8_24# OR2X1_LOC_270/Y 0.11fF
C51203 AND2X1_LOC_482/a_8_24# OR2X1_LOC_270/Y 0.01fF
C51660 OR2X1_LOC_270/Y AND2X1_LOC_252/a_8_24# 0.01fF
C55821 OR2X1_LOC_190/A OR2X1_LOC_270/Y 0.03fF
C17995 OR2X1_LOC_810/A OR2X1_LOC_66/Y 0.05fF
C20870 OR2X1_LOC_405/A OR2X1_LOC_810/A 0.13fF
C21264 AND2X1_LOC_316/a_8_24# OR2X1_LOC_810/A 0.05fF
C24093 OR2X1_LOC_810/A OR2X1_LOC_130/a_8_216# 0.14fF
C27296 OR2X1_LOC_810/A AND2X1_LOC_107/a_8_24# 0.22fF
C29539 OR2X1_LOC_810/A OR2X1_LOC_130/a_36_216# 0.17fF
C30111 OR2X1_LOC_810/A OR2X1_LOC_391/A 0.06fF
C34366 OR2X1_LOC_802/Y OR2X1_LOC_810/A 0.02fF
C38256 OR2X1_LOC_810/A OR2X1_LOC_113/A 0.04fF
C38995 OR2X1_LOC_105/a_8_216# OR2X1_LOC_810/A 0.17fF
C45469 OR2X1_LOC_473/a_8_216# OR2X1_LOC_810/A 0.15fF
C50249 OR2X1_LOC_105/Y OR2X1_LOC_810/A 0.08fF
C51089 OR2X1_LOC_473/a_36_216# OR2X1_LOC_810/A 0.12fF
C3078 OR2X1_LOC_574/A OR2X1_LOC_592/a_8_216# 0.11fF
C3120 OR2X1_LOC_574/A AND2X1_LOC_491/a_36_24# 0.08fF
C7775 OR2X1_LOC_574/A AND2X1_LOC_69/a_36_24# 0.06fF
C10688 OR2X1_LOC_574/A OR2X1_LOC_799/a_8_216# 0.06fF
C16174 OR2X1_LOC_574/A OR2X1_LOC_799/a_36_216# 0.16fF
C23011 OR2X1_LOC_574/A OR2X1_LOC_776/a_8_216# 0.16fF
C27619 OR2X1_LOC_405/A OR2X1_LOC_574/A 0.13fF
C33941 OR2X1_LOC_574/A OR2X1_LOC_776/a_36_216# 0.12fF
C38106 OR2X1_LOC_798/Y OR2X1_LOC_574/A 0.01fF
C42567 OR2X1_LOC_574/A AND2X1_LOC_491/a_8_24# 0.30fF
C45933 OR2X1_LOC_631/a_8_216# OR2X1_LOC_574/A 0.03fF
C52919 OR2X1_LOC_574/A AND2X1_LOC_69/a_8_24# 0.32fF
C3006 AND2X1_LOC_107/a_8_24# OR2X1_LOC_362/A 0.01fF
C6149 OR2X1_LOC_114/a_8_216# OR2X1_LOC_362/A 0.02fF
C11788 OR2X1_LOC_249/Y OR2X1_LOC_362/A 0.22fF
C14065 OR2X1_LOC_113/A OR2X1_LOC_362/A 0.01fF
C25748 OR2X1_LOC_105/Y OR2X1_LOC_362/A 0.02fF
C37587 AND2X1_LOC_251/a_8_24# OR2X1_LOC_362/A 0.01fF
C46300 OR2X1_LOC_843/a_8_216# OR2X1_LOC_362/A 0.01fF
C56232 AND2X1_LOC_250/a_8_24# OR2X1_LOC_362/A 0.01fF
C44622 AND2X1_LOC_65/a_8_24# OR2X1_LOC_473/Y 0.18fF
C3450 OR2X1_LOC_106/A OR2X1_LOC_67/A 0.02fF
C33401 OR2X1_LOC_106/A OR2X1_LOC_595/A 0.18fF
C35167 OR2X1_LOC_251/a_8_216# OR2X1_LOC_106/A 0.01fF
C35586 OR2X1_LOC_122/Y OR2X1_LOC_106/A 0.09fF
C39870 OR2X1_LOC_250/a_8_216# OR2X1_LOC_106/A 0.48fF
C57171 OR2X1_LOC_106/A VSS 0.49fF
C7659 OR2X1_LOC_757/A AND2X1_LOC_664/a_8_24# 0.01fF
C17250 OR2X1_LOC_757/A AND2X1_LOC_758/a_8_24# 0.01fF
C21551 OR2X1_LOC_757/A OR2X1_LOC_815/a_8_216# 0.03fF
C21708 OR2X1_LOC_757/A OR2X1_LOC_617/Y 0.03fF
C27006 OR2X1_LOC_757/A OR2X1_LOC_815/a_36_216# 0.01fF
C27125 OR2X1_LOC_757/A OR2X1_LOC_680/A 0.03fF
C36441 OR2X1_LOC_757/A OR2X1_LOC_665/a_8_216# 0.01fF
C39688 OR2X1_LOC_757/A VDD 0.08fF
C39774 OR2X1_LOC_757/A OR2X1_LOC_616/Y 0.01fF
C55988 OR2X1_LOC_528/Y OR2X1_LOC_757/A 0.18fF
C57967 OR2X1_LOC_757/A VSS -0.53fF
C27427 OR2X1_LOC_380/a_8_216# OR2X1_LOC_380/Y -0.00fF
C56706 OR2X1_LOC_380/Y VSS 0.11fF
C17068 OR2X1_LOC_764/Y AND2X1_LOC_769/a_8_24# 0.23fF
C31760 OR2X1_LOC_764/Y VDD 0.16fF
C57877 OR2X1_LOC_764/Y VSS 0.07fF
C1283 OR2X1_LOC_698/Y OR2X1_LOC_258/a_8_216# 0.01fF
C35047 VDD OR2X1_LOC_698/Y 0.33fF
C57579 OR2X1_LOC_698/Y VSS -0.11fF
C13045 AND2X1_LOC_160/Y AND2X1_LOC_161/Y 0.10fF
C18545 AND2X1_LOC_160/Y AND2X1_LOC_162/a_8_24# 0.09fF
C21131 AND2X1_LOC_160/Y OR2X1_LOC_697/Y 0.01fF
C26995 VDD AND2X1_LOC_160/Y 0.21fF
C37699 AND2X1_LOC_160/Y AND2X1_LOC_708/a_8_24# 0.21fF
C57699 AND2X1_LOC_160/Y VSS 0.20fF
C2282 OR2X1_LOC_391/A OR2X1_LOC_561/B 0.02fF
C6531 OR2X1_LOC_846/B OR2X1_LOC_561/B 0.07fF
C13356 OR2X1_LOC_391/a_8_216# OR2X1_LOC_561/B 0.02fF
C16732 OR2X1_LOC_848/a_8_216# OR2X1_LOC_561/B 0.01fF
C27759 OR2X1_LOC_846/a_8_216# OR2X1_LOC_561/B 0.42fF
C25880 AND2X1_LOC_24/a_8_24# OR2X1_LOC_33/B 0.01fF
C8012 OR2X1_LOC_224/a_8_216# OR2X1_LOC_183/Y 0.01fF
C19644 OR2X1_LOC_183/a_8_216# OR2X1_LOC_183/Y 0.01fF
C24587 OR2X1_LOC_224/Y OR2X1_LOC_183/Y 0.79fF
C29428 OR2X1_LOC_178/a_8_216# OR2X1_LOC_183/Y 0.01fF
C22834 OR2X1_LOC_248/a_8_216# OR2X1_LOC_248/A 0.47fF
C33230 VDD OR2X1_LOC_248/A -0.00fF
C44101 AND2X1_LOC_721/A OR2X1_LOC_248/A 0.01fF
C56413 OR2X1_LOC_248/A VSS 0.15fF
C37496 OR2X1_LOC_583/a_8_216# OR2X1_LOC_584/Y 0.39fF
C33241 OR2X1_LOC_7/a_8_216# OR2X1_LOC_7/Y 0.01fF
C33669 OR2X1_LOC_52/a_8_216# OR2X1_LOC_7/Y 0.01fF
C55376 OR2X1_LOC_7/Y OR2X1_LOC_16/a_8_216# 0.40fF
C4811 AND2X1_LOC_832/a_8_24# OR2X1_LOC_423/Y 0.04fF
C39422 OR2X1_LOC_423/Y OR2X1_LOC_589/Y 0.25fF
C45037 OR2X1_LOC_423/Y AND2X1_LOC_592/a_8_24# 0.03fF
C1529 OR2X1_LOC_109/Y OR2X1_LOC_368/Y 0.01fF
C3979 AND2X1_LOC_543/Y OR2X1_LOC_368/Y 0.78fF
C35340 OR2X1_LOC_368/a_8_216# OR2X1_LOC_368/Y 0.02fF
C44007 OR2X1_LOC_91/Y OR2X1_LOC_368/Y 0.11fF
C51387 OR2X1_LOC_312/Y OR2X1_LOC_368/Y 0.01fF
C54008 OR2X1_LOC_368/A OR2X1_LOC_368/Y 0.06fF
C56632 OR2X1_LOC_368/Y VSS 0.12fF
C38723 AND2X1_LOC_531/a_8_24# OR2X1_LOC_348/B 0.23fF
C9589 AND2X1_LOC_848/a_8_24# AND2X1_LOC_789/Y 0.01fF
C13442 OR2X1_LOC_701/a_8_216# AND2X1_LOC_789/Y 0.02fF
C23176 OR2X1_LOC_297/a_8_216# AND2X1_LOC_789/Y 0.02fF
C26130 AND2X1_LOC_848/a_36_24# AND2X1_LOC_789/Y 0.01fF
C26436 OR2X1_LOC_759/a_8_216# AND2X1_LOC_789/Y 0.01fF
C29008 OR2X1_LOC_261/a_8_216# AND2X1_LOC_789/Y 0.01fF
C35419 OR2X1_LOC_481/a_8_216# AND2X1_LOC_789/Y 0.01fF
C40833 OR2X1_LOC_700/a_8_216# AND2X1_LOC_789/Y 0.02fF
C53829 AND2X1_LOC_789/a_36_24# AND2X1_LOC_789/Y 0.01fF
C39449 OR2X1_LOC_385/Y OR2X1_LOC_586/Y 0.30fF
C51685 OR2X1_LOC_586/Y OR2X1_LOC_385/a_8_216# 0.03fF
C56040 VDD OR2X1_LOC_586/Y 0.05fF
C56218 AND2X1_LOC_389/a_8_24# OR2X1_LOC_586/Y 0.01fF
C56549 OR2X1_LOC_586/Y VSS -0.45fF
C4045 AND2X1_LOC_130/a_8_24# OR2X1_LOC_131/A 0.14fF
C21048 OR2X1_LOC_131/A OR2X1_LOC_131/a_8_216# 0.11fF
C30763 VDD OR2X1_LOC_131/A 0.44fF
C46573 OR2X1_LOC_131/A OR2X1_LOC_595/A 0.26fF
C57644 OR2X1_LOC_131/A VSS 0.32fF
C12392 OR2X1_LOC_542/B OR2X1_LOC_284/B 0.61fF
C43859 OR2X1_LOC_147/B OR2X1_LOC_284/B 0.08fF
C44225 OR2X1_LOC_114/B OR2X1_LOC_284/B 0.05fF
C56454 OR2X1_LOC_284/B VSS 0.25fF
C13281 OR2X1_LOC_614/Y OR2X1_LOC_196/a_8_216# 0.01fF
C49189 OR2X1_LOC_614/Y VDD 0.37fF
C51711 OR2X1_LOC_614/Y AND2X1_LOC_754/a_8_24# 0.05fF
C52528 OR2X1_LOC_196/Y OR2X1_LOC_614/Y 0.02fF
C58045 OR2X1_LOC_614/Y VSS 0.19fF
C7686 OR2X1_LOC_318/A OR2X1_LOC_318/B 0.23fF
C10265 AND2X1_LOC_604/a_8_24# OR2X1_LOC_318/B 0.01fF
C10622 OR2X1_LOC_318/B OR2X1_LOC_301/a_8_216# 0.01fF
C18788 OR2X1_LOC_318/a_8_216# OR2X1_LOC_318/B 0.08fF
C19249 OR2X1_LOC_776/a_8_216# OR2X1_LOC_318/B 0.01fF
C23301 OR2X1_LOC_318/B OR2X1_LOC_543/a_8_216# 0.07fF
C52072 OR2X1_LOC_831/a_8_216# OR2X1_LOC_318/B 0.01fF
C16055 AND2X1_LOC_597/a_8_24# OR2X1_LOC_676/Y 0.04fF
C20382 OR2X1_LOC_676/Y AND2X1_LOC_13/a_8_24# 0.02fF
C28392 OR2X1_LOC_676/Y AND2X1_LOC_516/a_8_24# 0.03fF
C32052 OR2X1_LOC_676/Y AND2X1_LOC_39/a_8_24# 0.03fF
C39731 OR2X1_LOC_676/Y AND2X1_LOC_16/a_8_24# 0.03fF
C7554 AND2X1_LOC_52/Y OR2X1_LOC_198/A 0.01fF
C12902 AND2X1_LOC_52/a_8_24# AND2X1_LOC_52/Y 0.01fF
C41456 AND2X1_LOC_52/Y OR2X1_LOC_197/a_8_216# 0.01fF
C8829 OR2X1_LOC_782/B OR2X1_LOC_160/Y 0.08fF
C29725 AND2X1_LOC_747/a_8_24# OR2X1_LOC_782/B 0.01fF
C19324 AND2X1_LOC_521/a_8_24# OR2X1_LOC_523/B 0.01fF
C6293 AND2X1_LOC_583/a_8_24# OR2X1_LOC_636/B 0.02fF
C15762 VDD OR2X1_LOC_451/B 0.21fF
C25555 OR2X1_LOC_451/a_8_216# OR2X1_LOC_451/B 0.08fF
C29985 AND2X1_LOC_428/a_8_24# OR2X1_LOC_451/B 0.01fF
C37453 AND2X1_LOC_584/a_8_24# OR2X1_LOC_451/B 0.20fF
C43430 OR2X1_LOC_635/a_8_216# OR2X1_LOC_451/B 0.08fF
C56426 OR2X1_LOC_451/B VSS 0.50fF
C1343 AND2X1_LOC_384/a_8_24# OR2X1_LOC_383/Y 0.24fF
C9848 OR2X1_LOC_383/Y OR2X1_LOC_391/A 0.05fF
C11488 VDD OR2X1_LOC_383/Y 0.20fF
C56992 OR2X1_LOC_383/Y VSS 0.04fF
C5811 OR2X1_LOC_542/B OR2X1_LOC_457/B 0.14fF
C15666 OR2X1_LOC_542/B OR2X1_LOC_254/a_8_216# 0.05fF
C21548 OR2X1_LOC_542/B OR2X1_LOC_284/a_8_216# 0.47fF
C26573 OR2X1_LOC_464/a_8_216# OR2X1_LOC_542/B 0.06fF
C26601 OR2X1_LOC_542/B OR2X1_LOC_254/A 0.02fF
C43662 OR2X1_LOC_254/B OR2X1_LOC_542/B 0.03fF
C6462 OR2X1_LOC_779/A OR2X1_LOC_708/a_8_216# 0.01fF
C15556 OR2X1_LOC_779/a_8_216# OR2X1_LOC_779/A 0.01fF
C34169 OR2X1_LOC_448/Y OR2X1_LOC_779/A 0.10fF
C38112 OR2X1_LOC_779/Y OR2X1_LOC_779/A 0.01fF
C42171 OR2X1_LOC_713/A OR2X1_LOC_779/A 0.16fF
C53426 OR2X1_LOC_708/Y OR2X1_LOC_779/A 0.01fF
C56240 OR2X1_LOC_779/A VSS 0.02fF
C41170 AND2X1_LOC_823/a_8_24# OR2X1_LOC_836/B 0.02fF
C52281 VDD OR2X1_LOC_836/B -0.00fF
C57030 OR2X1_LOC_836/B VSS 0.13fF
C34580 AND2X1_LOC_759/a_8_24# OR2X1_LOC_792/B 0.01fF
C22934 AND2X1_LOC_334/Y OR2X1_LOC_316/Y 0.01fF
C35696 OR2X1_LOC_837/A AND2X1_LOC_462/Y 0.24fF
C5758 OR2X1_LOC_405/A OR2X1_LOC_730/A 0.01fF
C11128 OR2X1_LOC_856/A OR2X1_LOC_198/A 1.07fF
C22420 OR2X1_LOC_379/Y OR2X1_LOC_856/A 0.73fF
C15055 OR2X1_LOC_434/a_8_216# OR2X1_LOC_339/A 0.10fF
C35063 AND2X1_LOC_431/a_8_24# OR2X1_LOC_339/A 0.11fF
C40569 OR2X1_LOC_434/A OR2X1_LOC_339/A 0.20fF
C7235 OR2X1_LOC_715/B AND2X1_LOC_109/a_8_24# 0.13fF
C7567 OR2X1_LOC_715/B AND2X1_LOC_516/a_8_24# 0.02fF
C18348 OR2X1_LOC_715/B OR2X1_LOC_66/Y 0.03fF
C21142 OR2X1_LOC_715/B OR2X1_LOC_405/A 0.11fF
C24200 OR2X1_LOC_715/B AND2X1_LOC_516/a_36_24# 0.01fF
C34652 OR2X1_LOC_715/B OR2X1_LOC_802/Y 0.35fF
C36392 OR2X1_LOC_715/B OR2X1_LOC_435/Y 0.28fF
C44454 OR2X1_LOC_715/B AND2X1_LOC_492/a_8_24# 0.03fF
C51414 OR2X1_LOC_715/B OR2X1_LOC_809/a_8_216# 0.71fF
C12021 OR2X1_LOC_516/Y OR2X1_LOC_816/A 0.07fF
C28615 OR2X1_LOC_516/Y AND2X1_LOC_506/a_8_24# 0.02fF
C31654 OR2X1_LOC_516/Y OR2X1_LOC_239/a_8_216# 0.02fF
C37114 OR2X1_LOC_516/Y OR2X1_LOC_239/a_36_216# 0.01fF
C37924 OR2X1_LOC_516/Y OR2X1_LOC_680/A 1.44fF
C6228 OR2X1_LOC_457/B OR2X1_LOC_787/B 0.14fF
C11831 OR2X1_LOC_457/a_8_216# OR2X1_LOC_787/B 0.07fF
C53523 AND2X1_LOC_74/a_8_24# OR2X1_LOC_787/B 0.08fF
C55846 OR2X1_LOC_286/a_8_216# OR2X1_LOC_286/Y 0.01fF
C24695 OR2X1_LOC_772/B OR2X1_LOC_846/B 0.04fF
C37703 OR2X1_LOC_317/B OR2X1_LOC_714/A 0.03fF
C43310 OR2X1_LOC_704/a_8_216# OR2X1_LOC_714/A -0.00fF
C16192 AND2X1_LOC_744/a_8_24# OR2X1_LOC_446/Y 0.05fF
C21325 OR2X1_LOC_450/A OR2X1_LOC_446/Y 0.01fF
C27265 OR2X1_LOC_446/Y AND2X1_LOC_424/a_8_24# 0.02fF
C30811 OR2X1_LOC_446/Y AND2X1_LOC_427/a_8_24# 0.24fF
C32291 OR2X1_LOC_446/Y AND2X1_LOC_695/a_8_24# 0.01fF
C37803 OR2X1_LOC_446/Y OR2X1_LOC_707/A 0.01fF
C47595 OR2X1_LOC_446/Y OR2X1_LOC_707/a_8_216# 0.01fF
C4201 OR2X1_LOC_227/Y AND2X1_LOC_224/a_8_24# 0.23fF
C11576 OR2X1_LOC_264/Y OR2X1_LOC_227/Y 0.07fF
C12859 OR2X1_LOC_754/A OR2X1_LOC_754/a_8_216# 0.13fF
C20550 OR2X1_LOC_754/A OR2X1_LOC_615/a_8_216# 0.13fF
C27994 VDD OR2X1_LOC_754/A 0.05fF
C45373 OR2X1_LOC_754/A OR2X1_LOC_816/A 0.11fF
C51245 OR2X1_LOC_754/A OR2X1_LOC_615/Y 0.26fF
C57284 OR2X1_LOC_754/A VSS -0.10fF
C38064 OR2X1_LOC_427/Y AND2X1_LOC_450/a_8_24# 0.04fF
C56999 OR2X1_LOC_427/Y VSS 0.22fF
C29504 OR2X1_LOC_253/Y AND2X1_LOC_254/a_8_24# 0.01fF
C37921 VDD OR2X1_LOC_253/Y 0.04fF
C56600 OR2X1_LOC_253/Y VSS 0.08fF
C8454 AND2X1_LOC_161/a_8_24# AND2X1_LOC_161/Y 0.01fF
C29555 AND2X1_LOC_161/Y AND2X1_LOC_162/a_8_24# 0.19fF
C37945 VDD AND2X1_LOC_161/Y 0.24fF
C57698 AND2X1_LOC_161/Y VSS -0.11fF
C15029 OR2X1_LOC_134/Y AND2X1_LOC_541/a_8_24# 0.01fF
C20984 OR2X1_LOC_134/a_8_216# OR2X1_LOC_134/Y 0.01fF
C49160 OR2X1_LOC_132/a_8_216# OR2X1_LOC_134/Y 0.05fF
C5249 OR2X1_LOC_334/B OR2X1_LOC_34/A 1.10fF
C45755 AND2X1_LOC_32/a_8_24# OR2X1_LOC_34/A 0.05fF
C36977 OR2X1_LOC_759/a_8_216# OR2X1_LOC_759/Y 0.03fF
C1687 VDD OR2X1_LOC_431/Y 0.09fF
C19190 OR2X1_LOC_45/Y OR2X1_LOC_431/Y 0.16fF
C31400 OR2X1_LOC_431/Y AND2X1_LOC_434/a_8_24# 0.04fF
C43110 OR2X1_LOC_431/Y OR2X1_LOC_172/Y 0.11fF
C57440 OR2X1_LOC_431/Y VSS 0.16fF
C37908 VDD OR2X1_LOC_281/Y -0.00fF
C40080 OR2X1_LOC_281/a_8_216# OR2X1_LOC_281/Y 0.01fF
C40908 OR2X1_LOC_292/a_8_216# OR2X1_LOC_281/Y 0.39fF
C56718 OR2X1_LOC_281/Y VSS 0.21fF
C857 OR2X1_LOC_697/Y AND2X1_LOC_708/a_8_24# 0.12fF
C28350 AND2X1_LOC_160/a_8_24# OR2X1_LOC_697/Y 0.01fF
C46200 VDD OR2X1_LOC_697/Y 0.32fF
C57648 OR2X1_LOC_697/Y VSS -0.19fF
C20435 OR2X1_LOC_823/Y AND2X1_LOC_836/a_8_24# 0.23fF
C43723 OR2X1_LOC_823/a_8_216# OR2X1_LOC_823/Y -0.00fF
C53532 VDD OR2X1_LOC_823/Y 0.12fF
C57674 OR2X1_LOC_823/Y VSS -0.14fF
C42838 AND2X1_LOC_391/Y OR2X1_LOC_248/Y 0.07fF
C54359 AND2X1_LOC_391/Y OR2X1_LOC_127/a_8_216# 0.03fF
C691 AND2X1_LOC_266/Y OR2X1_LOC_595/A 0.27fF
C1890 OR2X1_LOC_595/A OR2X1_LOC_131/a_8_216# 0.01fF
C4800 OR2X1_LOC_106/Y OR2X1_LOC_595/A 0.09fF
C11382 OR2X1_LOC_131/Y OR2X1_LOC_595/A 0.01fF
C11693 VDD OR2X1_LOC_595/A 0.34fF
C13974 AND2X1_LOC_557/a_8_24# OR2X1_LOC_595/A 0.02fF
C14747 OR2X1_LOC_767/a_8_216# OR2X1_LOC_595/A 0.01fF
C18889 OR2X1_LOC_118/a_8_216# OR2X1_LOC_595/A 0.07fF
C26547 OR2X1_LOC_666/A OR2X1_LOC_595/A 0.03fF
C26998 AND2X1_LOC_266/a_8_24# OR2X1_LOC_595/A 0.01fF
C38882 AND2X1_LOC_557/Y OR2X1_LOC_595/A 0.05fF
C44066 OR2X1_LOC_262/Y OR2X1_LOC_595/A 0.26fF
C53499 OR2X1_LOC_67/A OR2X1_LOC_595/A 0.03fF
C56321 OR2X1_LOC_595/A VSS -1.29fF
C4735 OR2X1_LOC_617/a_8_216# OR2X1_LOC_617/Y 0.01fF
C7347 OR2X1_LOC_617/Y AND2X1_LOC_621/a_8_24# 0.09fF
C7716 OR2X1_LOC_613/Y OR2X1_LOC_617/Y 0.03fF
C11536 OR2X1_LOC_252/a_8_216# OR2X1_LOC_617/Y 0.01fF
C21368 OR2X1_LOC_680/A OR2X1_LOC_617/Y 0.03fF
C21811 OR2X1_LOC_626/a_8_216# OR2X1_LOC_617/Y 0.01fF
C33911 VDD OR2X1_LOC_617/Y 0.22fF
C33989 OR2X1_LOC_616/Y OR2X1_LOC_617/Y 0.20fF
C41976 OR2X1_LOC_617/Y AND2X1_LOC_629/a_8_24# 0.23fF
C50216 OR2X1_LOC_528/Y OR2X1_LOC_617/Y 0.42fF
C57185 OR2X1_LOC_617/Y VSS 0.25fF
C11074 OR2X1_LOC_189/A OR2X1_LOC_498/a_8_216# 0.01fF
C23330 VDD OR2X1_LOC_189/A 0.21fF
C57376 OR2X1_LOC_189/A VSS -0.47fF
C14565 AND2X1_LOC_154/Y AND2X1_LOC_156/a_8_24# 0.03fF
C25028 VDD AND2X1_LOC_154/Y 0.21fF
C40730 AND2X1_LOC_154/a_8_24# AND2X1_LOC_154/Y 0.01fF
C57387 AND2X1_LOC_154/Y VSS 0.26fF
C2512 OR2X1_LOC_666/A AND2X1_LOC_287/Y 0.15fF
C6713 OR2X1_LOC_666/A OR2X1_LOC_89/a_8_216# 0.01fF
C18632 OR2X1_LOC_91/Y OR2X1_LOC_666/A 0.02fF
C22810 OR2X1_LOC_666/A AND2X1_LOC_284/a_8_24# 0.01fF
C27172 OR2X1_LOC_666/A OR2X1_LOC_279/a_8_216# 0.01fF
C38092 OR2X1_LOC_666/A OR2X1_LOC_279/Y 0.24fF
C39248 OR2X1_LOC_494/Y OR2X1_LOC_666/A 0.06fF
C42652 OR2X1_LOC_666/A OR2X1_LOC_89/Y 0.01fF
C53167 OR2X1_LOC_280/Y OR2X1_LOC_666/A 0.02fF
C55205 AND2X1_LOC_97/a_8_24# OR2X1_LOC_666/A 0.01fF
C29242 OR2X1_LOC_859/B OR2X1_LOC_391/A 0.02fF
C6645 AND2X1_LOC_666/a_8_24# OR2X1_LOC_121/A 0.04fF
C27298 OR2X1_LOC_776/A OR2X1_LOC_121/A 0.16fF
C32459 OR2X1_LOC_541/a_8_216# OR2X1_LOC_121/A 0.01fF
C38719 OR2X1_LOC_188/a_8_216# OR2X1_LOC_121/A 0.41fF
C49857 OR2X1_LOC_241/B OR2X1_LOC_121/A 0.03fF
C2425 OR2X1_LOC_264/Y AND2X1_LOC_265/a_8_24# 0.05fF
C4272 OR2X1_LOC_264/Y AND2X1_LOC_667/a_8_24# 0.03fF
C7153 OR2X1_LOC_264/Y AND2X1_LOC_517/a_36_24# 0.01fF
C7937 OR2X1_LOC_264/Y OR2X1_LOC_641/A 0.04fF
C8941 OR2X1_LOC_264/Y OR2X1_LOC_643/A 0.03fF
C41053 OR2X1_LOC_264/Y AND2X1_LOC_517/a_8_24# 0.03fF
C53999 OR2X1_LOC_264/Y OR2X1_LOC_520/Y 0.02fF
C34885 AND2X1_LOC_525/a_8_24# OR2X1_LOC_546/B 0.01fF
C6092 VDD OR2X1_LOC_162/A -0.00fF
C27351 OR2X1_LOC_162/A OR2X1_LOC_160/Y 0.06fF
C38303 OR2X1_LOC_162/A OR2X1_LOC_162/a_8_216# 0.39fF
C50434 OR2X1_LOC_161/a_8_216# OR2X1_LOC_162/A -0.00fF
C56383 OR2X1_LOC_162/A VSS 0.18fF
C6115 AND2X1_LOC_525/a_8_24# OR2X1_LOC_546/A 0.02fF
C11748 AND2X1_LOC_146/a_8_24# OR2X1_LOC_546/A 0.20fF
C16761 OR2X1_LOC_147/a_8_216# OR2X1_LOC_546/A 0.02fF
C34496 OR2X1_LOC_446/a_8_216# OR2X1_LOC_446/A 0.47fF
C56376 OR2X1_LOC_446/A VSS 0.15fF
C12640 VDD OR2X1_LOC_240/B 0.21fF
C22935 OR2X1_LOC_240/B AND2X1_LOC_232/a_8_24# 0.04fF
C34742 OR2X1_LOC_240/B OR2X1_LOC_240/a_8_216# 0.06fF
C57370 OR2X1_LOC_240/B VSS 0.17fF
C3016 OR2X1_LOC_624/B OR2X1_LOC_78/Y 0.02fF
C12093 AND2X1_LOC_766/a_8_24# OR2X1_LOC_78/Y 0.01fF
C23214 OR2X1_LOC_770/A OR2X1_LOC_78/Y 0.01fF
C25911 OR2X1_LOC_401/A OR2X1_LOC_78/Y 0.01fF
C36861 OR2X1_LOC_401/B OR2X1_LOC_78/Y 0.01fF
C38854 AND2X1_LOC_396/a_8_24# OR2X1_LOC_78/Y 0.01fF
C42219 AND2X1_LOC_765/a_8_24# OR2X1_LOC_78/Y 0.01fF
C50621 AND2X1_LOC_395/a_8_24# OR2X1_LOC_78/Y 0.01fF
C53434 OR2X1_LOC_770/B OR2X1_LOC_78/Y -0.00fF
C56009 VDD OR2X1_LOC_78/Y 0.59fF
C56756 OR2X1_LOC_78/Y VSS 0.19fF
C15368 VDD OR2X1_LOC_608/Y 0.06fF
C56428 OR2X1_LOC_608/Y VSS 0.10fF
C48618 OR2X1_LOC_420/a_8_216# OR2X1_LOC_591/A 0.47fF
C56885 OR2X1_LOC_591/A VSS 0.28fF
C11161 AND2X1_LOC_434/a_8_24# OR2X1_LOC_172/Y 0.04fF
C15910 OR2X1_LOC_230/a_8_216# OR2X1_LOC_172/Y 0.04fF
C39991 OR2X1_LOC_45/a_8_216# OR2X1_LOC_172/Y 0.44fF
C5336 OR2X1_LOC_239/Y OR2X1_LOC_816/A 0.06fF
C22149 AND2X1_LOC_506/a_8_24# OR2X1_LOC_239/Y 0.23fF
C25160 OR2X1_LOC_239/a_8_216# OR2X1_LOC_239/Y 0.01fF
C2534 VDD OR2X1_LOC_420/Y 0.15fF
C36483 OR2X1_LOC_420/Y AND2X1_LOC_447/a_8_24# 0.23fF
C57441 OR2X1_LOC_420/Y VSS -0.12fF
C10165 OR2X1_LOC_282/Y AND2X1_LOC_285/a_8_24# 0.01fF
C13188 VDD OR2X1_LOC_282/Y 0.04fF
C57495 OR2X1_LOC_282/Y VSS 0.08fF
C10600 OR2X1_LOC_533/A OR2X1_LOC_533/a_8_216# 0.01fF
C51206 VDD OR2X1_LOC_533/A 0.21fF
C56448 OR2X1_LOC_533/A VSS -0.05fF
C17890 OR2X1_LOC_670/Y AND2X1_LOC_673/a_8_24# 0.23fF
C26683 VDD OR2X1_LOC_670/Y 0.12fF
C57117 OR2X1_LOC_670/Y VSS 0.06fF
C3073 OR2X1_LOC_837/B AND2X1_LOC_825/a_8_24# 0.01fF
C6688 OR2X1_LOC_837/A OR2X1_LOC_837/B 0.12fF
C17753 OR2X1_LOC_837/B OR2X1_LOC_837/a_8_216# 0.02fF
C22631 OR2X1_LOC_837/B OR2X1_LOC_27/Y 0.03fF
C27049 OR2X1_LOC_58/Y OR2X1_LOC_837/B 0.03fF
C32073 VDD OR2X1_LOC_837/B 0.31fF
C33985 OR2X1_LOC_837/B OR2X1_LOC_416/Y 0.03fF
C45105 OR2X1_LOC_837/B AND2X1_LOC_462/a_8_24# 0.07fF
C55327 OR2X1_LOC_837/B OR2X1_LOC_32/a_8_216# 0.05fF
C57483 OR2X1_LOC_837/B VSS 0.17fF
C532 OR2X1_LOC_91/Y OR2X1_LOC_437/a_8_216# 0.03fF
C9320 OR2X1_LOC_91/Y OR2X1_LOC_107/a_8_216# 0.05fF
C10591 OR2X1_LOC_91/Y OR2X1_LOC_179/a_8_216# 0.05fF
C21420 OR2X1_LOC_91/Y OR2X1_LOC_368/A 0.03fF
C28785 OR2X1_LOC_91/Y OR2X1_LOC_329/B 0.07fF
C35417 OR2X1_LOC_91/Y OR2X1_LOC_89/Y 0.01fF
C36866 OR2X1_LOC_91/Y OR2X1_LOC_91/a_8_216# 0.03fF
C37154 OR2X1_LOC_91/Y OR2X1_LOC_315/a_8_216# 0.08fF
C45882 OR2X1_LOC_165/a_8_216# OR2X1_LOC_91/Y 0.05fF
C47307 OR2X1_LOC_91/Y OR2X1_LOC_680/A 0.03fF
C54830 OR2X1_LOC_91/Y AND2X1_LOC_168/a_8_24# 0.04fF
C55807 OR2X1_LOC_91/Y OR2X1_LOC_89/a_8_216# 0.04fF
C21360 OR2X1_LOC_494/A OR2X1_LOC_384/a_8_216# 0.48fF
C52585 OR2X1_LOC_494/A AND2X1_LOC_348/A 0.27fF
C57939 OR2X1_LOC_494/A VSS 0.43fF
C3761 OR2X1_LOC_305/Y VDD 0.16fF
C18815 OR2X1_LOC_305/Y AND2X1_LOC_307/a_8_24# 0.01fF
C33968 AND2X1_LOC_777/a_8_24# OR2X1_LOC_305/Y 0.11fF
C41438 OR2X1_LOC_305/Y OR2X1_LOC_135/Y 0.01fF
C58000 OR2X1_LOC_305/Y VSS 0.24fF
C21106 OR2X1_LOC_132/a_8_216# OR2X1_LOC_132/Y 0.05fF
C43085 OR2X1_LOC_132/Y AND2X1_LOC_541/a_8_24# 0.23fF
C15324 OR2X1_LOC_313/Y OR2X1_LOC_418/a_8_216# 0.01fF
C40584 VDD OR2X1_LOC_313/Y 0.22fF
C45915 OR2X1_LOC_313/Y AND2X1_LOC_317/a_8_24# 0.24fF
C57300 OR2X1_LOC_313/Y VSS 0.22fF
C1307 OR2X1_LOC_610/a_8_216# OR2X1_LOC_647/B 0.03fF
C19647 OR2X1_LOC_610/Y OR2X1_LOC_647/B 0.04fF
C36101 AND2X1_LOC_612/a_8_24# OR2X1_LOC_647/B 0.02fF
C6187 AND2X1_LOC_802/B OR2X1_LOC_312/Y 0.03fF
C10145 OR2X1_LOC_368/a_8_216# OR2X1_LOC_312/Y 0.01fF
C11796 OR2X1_LOC_312/Y AND2X1_LOC_457/a_8_24# 0.01fF
C23828 AND2X1_LOC_543/a_8_24# OR2X1_LOC_312/Y 0.01fF
C35988 OR2X1_LOC_329/B OR2X1_LOC_312/Y 0.29fF
C39741 OR2X1_LOC_312/Y AND2X1_LOC_802/Y 0.24fF
C47794 AND2X1_LOC_355/a_8_24# OR2X1_LOC_312/Y 0.01fF
C21938 OR2X1_LOC_607/a_8_216# OR2X1_LOC_67/Y 0.02fF
C32874 OR2X1_LOC_607/a_36_216# OR2X1_LOC_67/Y 0.01fF
C51114 OR2X1_LOC_117/a_8_216# OR2X1_LOC_67/Y 0.01fF
C25907 OR2X1_LOC_613/Y OR2X1_LOC_616/Y 0.14fF
C48953 OR2X1_LOC_187/a_8_216# OR2X1_LOC_613/Y 0.01fF
C55410 OR2X1_LOC_613/Y AND2X1_LOC_621/a_8_24# 0.01fF
C10404 OR2X1_LOC_825/Y OR2X1_LOC_826/Y 0.21fF
C30774 OR2X1_LOC_826/Y AND2X1_LOC_837/a_8_24# 0.23fF
C38625 VDD OR2X1_LOC_826/Y 0.16fF
C56883 OR2X1_LOC_826/Y VSS 0.07fF
C658 OR2X1_LOC_680/A OR2X1_LOC_816/A 0.03fF
C1338 OR2X1_LOC_816/A AND2X1_LOC_790/a_8_24# 0.03fF
C5810 OR2X1_LOC_615/a_8_216# OR2X1_LOC_816/A 0.03fF
C6557 AND2X1_LOC_631/a_8_24# OR2X1_LOC_816/A 0.01fF
C12395 OR2X1_LOC_816/A AND2X1_LOC_793/B 0.01fF
C13943 OR2X1_LOC_666/Y OR2X1_LOC_816/A 0.12fF
C17169 OR2X1_LOC_482/Y OR2X1_LOC_816/A 10.04fF
C23290 OR2X1_LOC_497/Y OR2X1_LOC_816/A 0.01fF
C29468 OR2X1_LOC_528/Y OR2X1_LOC_816/A 0.13fF
C29615 AND2X1_LOC_483/a_8_24# OR2X1_LOC_816/A 0.01fF
C36438 OR2X1_LOC_615/Y OR2X1_LOC_816/A 0.58fF
C38022 AND2X1_LOC_631/Y OR2X1_LOC_816/A 0.91fF
C46423 OR2X1_LOC_816/A OR2X1_LOC_754/Y 0.05fF
C51361 AND2X1_LOC_186/a_8_24# OR2X1_LOC_816/A 0.01fF
C54330 OR2X1_LOC_816/A OR2X1_LOC_754/a_8_216# 0.03fF
C41417 OR2X1_LOC_179/a_8_216# OR2X1_LOC_178/Y 0.01fF
C10225 OR2X1_LOC_316/Y AND2X1_LOC_139/B 0.03fF
C7011 OR2X1_LOC_600/a_8_216# AND2X1_LOC_447/Y 0.03fF
C25087 OR2X1_LOC_601/a_8_216# AND2X1_LOC_447/Y 0.12fF
C39752 OR2X1_LOC_424/a_8_216# AND2X1_LOC_447/Y 0.14fF
C51411 AND2X1_LOC_447/Y AND2X1_LOC_447/a_8_24# 0.01fF
C13504 AND2X1_LOC_506/a_8_24# AND2X1_LOC_508/A 0.01fF
C16532 AND2X1_LOC_508/A OR2X1_LOC_239/a_8_216# 0.01fF
C28664 OR2X1_LOC_166/a_8_216# AND2X1_LOC_535/Y 0.01fF
C37667 AND2X1_LOC_535/Y AND2X1_LOC_798/Y 0.16fF
C40919 AND2X1_LOC_535/Y OR2X1_LOC_329/B 0.03fF
C44797 AND2X1_LOC_535/Y AND2X1_LOC_802/Y 0.03fF
C50463 AND2X1_LOC_535/Y AND2X1_LOC_809/a_8_24# 0.01fF
C52712 AND2X1_LOC_535/Y AND2X1_LOC_355/a_8_24# 0.01fF
C25552 AND2X1_LOC_557/Y AND2X1_LOC_557/a_8_24# 0.01fF
C52993 OR2X1_LOC_405/A OR2X1_LOC_776/A 0.07fF
C17207 VDD OR2X1_LOC_160/Y 0.12fF
C22039 AND2X1_LOC_158/a_8_24# OR2X1_LOC_160/Y 0.24fF
C40422 OR2X1_LOC_156/Y OR2X1_LOC_160/Y 0.18fF
C49617 OR2X1_LOC_160/Y OR2X1_LOC_162/a_8_216# 0.07fF
C56334 OR2X1_LOC_160/Y VSS 0.26fF
C291 VDD OR2X1_LOC_249/Y 0.24fF
C47608 AND2X1_LOC_595/a_8_24# OR2X1_LOC_249/Y 0.23fF
C49089 OR2X1_LOC_249/Y AND2X1_LOC_250/a_8_24# 0.01fF
C54570 OR2X1_LOC_249/Y OR2X1_LOC_343/B 0.01fF
C56900 OR2X1_LOC_249/Y VSS 0.21fF
C8453 OR2X1_LOC_450/A OR2X1_LOC_707/A 0.05fF
C34517 OR2X1_LOC_707/A OR2X1_LOC_707/a_8_216# 0.47fF
C57105 OR2X1_LOC_707/A VSS 0.15fF
C2360 OR2X1_LOC_196/B OR2X1_LOC_196/a_8_216# 0.07fF
C1581 AND2X1_LOC_504/a_8_24# OR2X1_LOC_507/A 0.20fF
C15102 AND2X1_LOC_505/a_8_24# OR2X1_LOC_507/A 0.01fF
C16629 AND2X1_LOC_395/a_8_24# OR2X1_LOC_401/A 0.21fF
C34232 AND2X1_LOC_766/a_8_24# OR2X1_LOC_401/A 0.01fF
C9613 OR2X1_LOC_756/Y OR2X1_LOC_756/a_8_216# 0.01fF
C14312 OR2X1_LOC_756/Y VDD 0.05fF
C43642 OR2X1_LOC_756/Y AND2X1_LOC_757/a_8_24# 0.01fF
C57929 OR2X1_LOC_756/Y VSS 0.10fF
C9367 OR2X1_LOC_621/B AND2X1_LOC_670/a_36_24# 0.01fF
C14413 OR2X1_LOC_621/B OR2X1_LOC_624/B 0.27fF
C37508 OR2X1_LOC_621/B OR2X1_LOC_621/a_8_216# 0.01fF
C46116 OR2X1_LOC_673/B OR2X1_LOC_621/B 0.94fF
C54416 OR2X1_LOC_621/B AND2X1_LOC_670/a_8_24# 0.04fF
C57586 OR2X1_LOC_621/B VSS -0.11fF
C3477 OR2X1_LOC_260/Y OR2X1_LOC_345/A 0.01fF
C49597 AND2X1_LOC_600/a_8_24# OR2X1_LOC_602/B 0.01fF
C14325 OR2X1_LOC_105/Y VDD 0.13fF
C20832 OR2X1_LOC_105/Y OR2X1_LOC_643/A 0.02fF
C39524 OR2X1_LOC_105/Y AND2X1_LOC_106/a_8_24# 0.11fF
C44565 OR2X1_LOC_105/Y AND2X1_LOC_251/a_8_24# 0.11fF
C57853 OR2X1_LOC_105/Y VSS 0.34fF
C11590 OR2X1_LOC_506/a_8_216# OR2X1_LOC_130/Y 0.40fF
C41551 OR2X1_LOC_66/Y OR2X1_LOC_130/Y 0.18fF
C55473 VDD OR2X1_LOC_130/Y 0.27fF
C56285 OR2X1_LOC_130/Y VSS 0.07fF
C8893 OR2X1_LOC_629/A OR2X1_LOC_629/B 0.39fF
C11141 OR2X1_LOC_629/A OR2X1_LOC_629/a_8_216# 0.51fF
C23387 VDD OR2X1_LOC_629/A 0.02fF
C57132 OR2X1_LOC_629/A VSS 0.20fF
C24987 AND2X1_LOC_65/a_8_24# OR2X1_LOC_231/A 0.20fF
C35581 OR2X1_LOC_231/A AND2X1_LOC_230/a_8_24# 0.01fF
C55700 OR2X1_LOC_405/A OR2X1_LOC_231/A 0.03fF
C9477 VDD OR2X1_LOC_247/Y 0.33fF
C34493 AND2X1_LOC_72/a_8_24# OR2X1_LOC_247/Y 0.23fF
C56995 OR2X1_LOC_247/Y VSS 0.16fF
C26651 OR2X1_LOC_620/B OR2X1_LOC_547/a_8_216# 0.47fF
C6780 OR2X1_LOC_457/B OR2X1_LOC_457/a_8_216# 0.07fF
C37255 OR2X1_LOC_147/B OR2X1_LOC_457/B 0.03fF
C57213 OR2X1_LOC_457/B VSS 0.09fF
C824 AND2X1_LOC_583/a_8_24# OR2X1_LOC_636/A 0.09fF
C26950 OR2X1_LOC_156/B VDD -0.00fF
C39163 OR2X1_LOC_156/B OR2X1_LOC_156/a_8_216# 0.39fF
C58104 OR2X1_LOC_156/B VSS 0.17fF
C9256 AND2X1_LOC_448/Y AND2X1_LOC_448/a_8_24# 0.05fF
C42624 AND2X1_LOC_630/a_8_24# AND2X1_LOC_632/A 0.01fF
C10317 AND2X1_LOC_98/Y AND2X1_LOC_721/A 0.02fF
C13950 AND2X1_LOC_98/Y AND2X1_LOC_99/a_8_24# 0.06fF
C55142 OR2X1_LOC_125/a_8_216# AND2X1_LOC_98/Y 0.47fF
C55563 VDD AND2X1_LOC_98/Y 0.27fF
C56160 AND2X1_LOC_98/Y OR2X1_LOC_248/Y 0.04fF
C57407 AND2X1_LOC_98/Y VSS 0.32fF
C13360 OR2X1_LOC_779/Y OR2X1_LOC_779/a_36_216# 0.01fF
C4157 OR2X1_LOC_168/a_8_216# OR2X1_LOC_840/A 0.33fF
C18596 OR2X1_LOC_840/A AND2X1_LOC_167/a_8_24# 0.12fF
C30495 OR2X1_LOC_840/A AND2X1_LOC_601/a_8_24# 0.13fF
C43240 OR2X1_LOC_405/A OR2X1_LOC_840/A 0.27fF
C5895 OR2X1_LOC_101/a_8_216# OR2X1_LOC_520/Y 0.02fF
C16638 OR2X1_LOC_520/Y AND2X1_LOC_518/a_8_24# 0.10fF
C22235 OR2X1_LOC_520/Y OR2X1_LOC_520/B 1.08fF
C30125 OR2X1_LOC_520/Y AND2X1_LOC_517/a_8_24# 0.02fF
C1868 OR2X1_LOC_196/Y AND2X1_LOC_754/a_8_24# 0.24fF
C8160 OR2X1_LOC_680/A AND2X1_LOC_631/Y 0.03fF
C45834 VDD AND2X1_LOC_637/Y 0.01fF
C50755 AND2X1_LOC_637/Y AND2X1_LOC_638/a_8_24# 0.13fF
C56638 AND2X1_LOC_637/Y VSS 0.08fF
C477 AND2X1_LOC_831/a_8_24# OR2X1_LOC_416/Y 0.01fF
C3492 OR2X1_LOC_316/Y OR2X1_LOC_416/Y 2.98fF
C4211 AND2X1_LOC_301/a_8_24# OR2X1_LOC_416/Y 0.01fF
C5513 OR2X1_LOC_290/Y OR2X1_LOC_416/Y 0.01fF
C10792 OR2X1_LOC_416/Y AND2X1_LOC_462/a_8_24# 0.01fF
C11186 AND2X1_LOC_334/a_8_24# OR2X1_LOC_416/Y 0.01fF
C12947 OR2X1_LOC_416/Y OR2X1_LOC_75/a_8_216# 0.01fF
C29389 OR2X1_LOC_416/Y AND2X1_LOC_634/a_8_24# 0.01fF
C31117 OR2X1_LOC_462/a_8_216# OR2X1_LOC_416/Y 0.05fF
C33209 OR2X1_LOC_416/Y OR2X1_LOC_27/a_8_216# 0.01fF
C50736 OR2X1_LOC_290/a_8_216# OR2X1_LOC_416/Y 0.01fF
C21039 OR2X1_LOC_318/A OR2X1_LOC_776/Y 0.06fF
C31973 OR2X1_LOC_318/a_8_216# OR2X1_LOC_776/Y 0.02fF
C31582 AND2X1_LOC_437/a_8_24# OR2X1_LOC_168/Y 0.07fF
C49255 AND2X1_LOC_176/a_8_24# OR2X1_LOC_168/Y 0.03fF
C30862 OR2X1_LOC_149/B AND2X1_LOC_525/a_8_24# 0.29fF
C3164 AND2X1_LOC_313/a_36_24# OR2X1_LOC_308/Y 0.01fF
C5660 AND2X1_LOC_423/a_8_24# OR2X1_LOC_308/Y 0.03fF
C6615 AND2X1_LOC_698/a_8_24# OR2X1_LOC_308/Y 0.04fF
C30747 OR2X1_LOC_447/A OR2X1_LOC_308/Y 0.05fF
C39890 OR2X1_LOC_317/B OR2X1_LOC_308/Y 0.06fF
C41785 OR2X1_LOC_447/a_8_216# OR2X1_LOC_308/Y 0.03fF
C43884 OR2X1_LOC_709/B OR2X1_LOC_308/Y 0.04fF
C45518 OR2X1_LOC_704/a_8_216# OR2X1_LOC_308/Y 0.03fF
C48325 AND2X1_LOC_313/a_8_24# OR2X1_LOC_308/Y 0.03fF
C49561 OR2X1_LOC_709/a_8_216# OR2X1_LOC_308/Y 0.04fF
C13854 OR2X1_LOC_708/Y OR2X1_LOC_708/a_8_216# -0.00fF
C13261 OR2X1_LOC_156/Y OR2X1_LOC_160/a_8_216# 0.38fF
C19318 OR2X1_LOC_156/Y VDD 0.06fF
C58028 OR2X1_LOC_156/Y VSS 0.21fF
C22202 OR2X1_LOC_828/Y OR2X1_LOC_198/A 0.17fF
C27775 VDD OR2X1_LOC_828/Y 0.09fF
C36642 OR2X1_LOC_828/a_8_216# OR2X1_LOC_828/Y 0.05fF
C56699 OR2X1_LOC_828/Y VSS 0.13fF
C375 VDD OR2X1_LOC_435/Y 0.12fF
C48081 AND2X1_LOC_594/a_8_24# OR2X1_LOC_435/Y 0.24fF
C53567 OR2X1_LOC_653/B OR2X1_LOC_435/Y 0.16fF
C57156 OR2X1_LOC_435/Y VSS 0.14fF
C18888 OR2X1_LOC_368/a_8_216# AND2X1_LOC_543/Y 0.01fF
C20576 AND2X1_LOC_543/Y AND2X1_LOC_457/a_8_24# 0.01fF
C32407 AND2X1_LOC_543/Y AND2X1_LOC_543/a_8_24# 0.01fF
C2821 AND2X1_LOC_787/A AND2X1_LOC_168/a_8_24# 0.01fF
C4637 AND2X1_LOC_787/A OR2X1_LOC_437/a_8_216# 0.10fF
C8708 AND2X1_LOC_787/A AND2X1_LOC_457/a_8_24# 0.11fF
C15692 AND2X1_LOC_787/A OR2X1_LOC_437/a_36_216# 0.01fF
C40960 AND2X1_LOC_787/A OR2X1_LOC_91/a_8_216# 0.01fF
C50080 OR2X1_LOC_165/a_8_216# AND2X1_LOC_787/A 0.01fF
C1805 AND2X1_LOC_831/Y AND2X1_LOC_138/a_8_24# 0.01fF
C16507 AND2X1_LOC_520/a_8_24# AND2X1_LOC_831/Y 0.02fF
C17957 AND2X1_LOC_831/Y AND2X1_LOC_831/a_36_24# 0.01fF
C18403 AND2X1_LOC_831/Y AND2X1_LOC_138/a_36_24# 0.02fF
C29329 OR2X1_LOC_329/B AND2X1_LOC_831/Y 0.07fF
C39355 OR2X1_LOC_518/a_8_216# AND2X1_LOC_831/Y 0.03fF
C39466 AND2X1_LOC_112/a_8_24# AND2X1_LOC_831/Y 0.01fF
C47710 AND2X1_LOC_332/a_8_24# AND2X1_LOC_831/Y 0.04fF
C52789 AND2X1_LOC_303/A OR2X1_LOC_316/Y -0.00fF
C53897 OR2X1_LOC_464/a_8_216# OR2X1_LOC_471/B -0.00fF
C226 OR2X1_LOC_329/B AND2X1_LOC_112/a_8_24# 0.05fF
C1138 OR2X1_LOC_329/B OR2X1_LOC_674/a_8_216# 0.18fF
C6260 AND2X1_LOC_784/A OR2X1_LOC_329/B 0.07fF
C7178 OR2X1_LOC_329/B OR2X1_LOC_280/Y 0.09fF
C10965 OR2X1_LOC_329/B OR2X1_LOC_237/Y 0.05fF
C11303 OR2X1_LOC_329/B AND2X1_LOC_112/a_36_24# 0.01fF
C11964 OR2X1_LOC_329/B AND2X1_LOC_116/a_8_24# 0.01fF
C14245 OR2X1_LOC_106/Y OR2X1_LOC_329/B 0.17fF
C16492 OR2X1_LOC_329/B OR2X1_LOC_495/a_8_216# 0.02fF
C16606 OR2X1_LOC_329/B OR2X1_LOC_238/a_8_216# 0.02fF
C20496 OR2X1_LOC_329/B AND2X1_LOC_798/A 0.03fF
C23831 OR2X1_LOC_329/B AND2X1_LOC_116/Y 0.01fF
C24897 OR2X1_LOC_329/B OR2X1_LOC_482/Y 0.06fF
C26678 OR2X1_LOC_329/B OR2X1_LOC_316/Y 0.03fF
C27886 OR2X1_LOC_179/a_8_216# OR2X1_LOC_329/B 0.03fF
C28873 OR2X1_LOC_329/B OR2X1_LOC_311/Y 0.03fF
C30377 OR2X1_LOC_329/B OR2X1_LOC_108/a_8_216# 0.03fF
C34755 OR2X1_LOC_329/B AND2X1_LOC_473/a_8_24# 0.01fF
C38886 OR2X1_LOC_179/Y OR2X1_LOC_329/B 0.01fF
C41376 OR2X1_LOC_329/B OR2X1_LOC_108/Y 0.21fF
C44915 OR2X1_LOC_329/B OR2X1_LOC_495/Y 0.03fF
C45306 AND2X1_LOC_776/a_8_24# OR2X1_LOC_329/B 0.13fF
C46794 OR2X1_LOC_329/B OR2X1_LOC_280/a_8_216# 0.03fF
C50063 OR2X1_LOC_329/B AND2X1_LOC_802/Y 0.03fF
C51726 OR2X1_LOC_329/B OR2X1_LOC_312/a_8_216# 0.01fF
C51867 OR2X1_LOC_329/B AND2X1_LOC_114/a_8_24# 0.04fF
C55526 OR2X1_LOC_329/B AND2X1_LOC_809/a_8_24# 0.03fF
C55955 AND2X1_LOC_539/Y OR2X1_LOC_329/B 0.03fF
C56092 OR2X1_LOC_329/B OR2X1_LOC_237/a_8_216# 0.03fF
C17436 OR2X1_LOC_262/Y AND2X1_LOC_266/Y 0.06fF
C43739 OR2X1_LOC_262/Y AND2X1_LOC_266/a_8_24# 0.03fF
C54157 OR2X1_LOC_262/Y OR2X1_LOC_72/a_8_216# 0.09fF
C42025 OR2X1_LOC_117/Y OR2X1_LOC_67/A 0.01fF
C53231 OR2X1_LOC_117/Y OR2X1_LOC_67/a_8_216# 0.01fF
C55176 OR2X1_LOC_117/a_8_216# OR2X1_LOC_117/Y 0.04fF
C1659 OR2X1_LOC_778/Y OR2X1_LOC_778/a_8_216# 0.01fF
C17788 OR2X1_LOC_317/a_8_216# OR2X1_LOC_778/Y 0.33fF
C20639 OR2X1_LOC_778/Y OR2X1_LOC_704/a_8_216# 0.30fF
C41134 OR2X1_LOC_317/A OR2X1_LOC_778/Y 0.08fF
C47734 OR2X1_LOC_405/A OR2X1_LOC_778/Y 0.14fF
C9610 OR2X1_LOC_335/Y AND2X1_LOC_438/a_8_24# 0.03fF
C45563 OR2X1_LOC_335/Y AND2X1_LOC_438/a_36_24# 0.01fF
C14991 OR2X1_LOC_494/a_8_216# AND2X1_LOC_721/A 0.01fF
C33000 AND2X1_LOC_721/A AND2X1_LOC_247/a_8_24# 0.01fF
C43449 AND2X1_LOC_342/a_8_24# AND2X1_LOC_721/A 0.01fF
C51196 AND2X1_LOC_344/a_8_24# AND2X1_LOC_721/A 0.01fF
C52499 AND2X1_LOC_721/A OR2X1_LOC_248/a_8_216# 0.01fF
C320 AND2X1_LOC_83/a_8_24# OR2X1_LOC_624/B 0.02fF
C5094 OR2X1_LOC_624/B AND2X1_LOC_617/a_8_24# 0.01fF
C9883 AND2X1_LOC_393/a_8_24# OR2X1_LOC_624/B 0.02fF
C25441 OR2X1_LOC_621/a_8_216# OR2X1_LOC_624/B 0.01fF
C25884 OR2X1_LOC_624/B AND2X1_LOC_103/a_8_24# 0.02fF
C29249 OR2X1_LOC_624/B AND2X1_LOC_616/a_8_24# 0.01fF
C33856 OR2X1_LOC_673/B OR2X1_LOC_624/B 0.02fF
C42115 OR2X1_LOC_624/B AND2X1_LOC_670/a_8_24# -0.00fF
C52917 OR2X1_LOC_624/B AND2X1_LOC_79/a_8_24# 0.01fF
C377 AND2X1_LOC_266/a_8_24# AND2X1_LOC_266/Y 0.03fF
C16992 AND2X1_LOC_266/a_36_24# AND2X1_LOC_266/Y 0.02fF
C41026 VDD AND2X1_LOC_266/Y 0.04fF
C41155 AND2X1_LOC_266/Y AND2X1_LOC_267/a_8_24# 0.02fF
C51384 AND2X1_LOC_266/Y AND2X1_LOC_249/a_8_24# 0.01fF
C56508 AND2X1_LOC_266/Y VSS 0.22fF
C23621 AND2X1_LOC_101/a_8_24# OR2X1_LOC_813/Y 0.01fF
C24698 OR2X1_LOC_821/a_8_216# OR2X1_LOC_813/Y 0.01fF
C32295 AND2X1_LOC_99/a_8_24# OR2X1_LOC_813/Y 0.01fF
C41666 OR2X1_LOC_316/Y AND2X1_LOC_634/Y 0.03fF
C43804 OR2X1_LOC_290/Y AND2X1_LOC_634/Y 0.15fF
C49583 AND2X1_LOC_334/a_8_24# AND2X1_LOC_634/Y 0.19fF
C33693 OR2X1_LOC_134/a_8_216# AND2X1_LOC_541/Y 0.01fF
C40874 AND2X1_LOC_541/Y AND2X1_LOC_361/a_8_24# 0.04fF
C34421 AND2X1_LOC_633/Y AND2X1_LOC_633/a_36_24# 0.01fF
C36109 OR2X1_LOC_316/Y AND2X1_LOC_633/Y 0.02fF
C4096 OR2X1_LOC_176/a_8_216# AND2X1_LOC_784/A 0.03fF
C14506 AND2X1_LOC_784/A OR2X1_LOC_91/a_8_216# 0.03fF
C20036 AND2X1_LOC_784/A OR2X1_LOC_91/a_36_216# 0.01fF
C37977 AND2X1_LOC_370/a_8_24# AND2X1_LOC_784/A 0.04fF
C45869 AND2X1_LOC_784/A AND2X1_LOC_335/a_8_24# 0.03fF
C52818 OR2X1_LOC_235/a_8_216# OR2X1_LOC_235/Y -0.00fF
C31138 OR2X1_LOC_173/Y OR2X1_LOC_173/a_8_216# -0.00fF
C5680 AND2X1_LOC_383/a_8_24# OR2X1_LOC_292/Y 0.23fF
C3735 OR2X1_LOC_108/Y OR2X1_LOC_680/A 0.05fF
C4453 AND2X1_LOC_778/a_36_24# OR2X1_LOC_680/A 0.01fF
C6265 OR2X1_LOC_187/a_8_216# OR2X1_LOC_680/A 0.01fF
C6445 OR2X1_LOC_680/A OR2X1_LOC_615/Y 0.03fF
C8772 OR2X1_LOC_680/A OR2X1_LOC_525/a_8_216# 0.03fF
C12650 OR2X1_LOC_680/A AND2X1_LOC_778/Y 0.46fF
C16136 OR2X1_LOC_516/a_8_216# OR2X1_LOC_680/A 0.02fF
C16900 AND2X1_LOC_758/a_8_24# OR2X1_LOC_680/A 0.02fF
C19163 OR2X1_LOC_496/Y OR2X1_LOC_680/A 0.12fF
C21288 AND2X1_LOC_186/a_8_24# OR2X1_LOC_680/A 0.02fF
C24700 AND2X1_LOC_778/a_8_24# OR2X1_LOC_680/A 0.03fF
C27232 OR2X1_LOC_680/A OR2X1_LOC_626/a_8_216# 0.03fF
C28193 OR2X1_LOC_680/A OR2X1_LOC_331/a_8_216# 0.09fF
C32123 OR2X1_LOC_680/A AND2X1_LOC_188/a_8_24# 0.07fF
C32552 OR2X1_LOC_680/A OR2X1_LOC_505/Y 0.03fF
C33416 AND2X1_LOC_758/a_36_24# OR2X1_LOC_680/A 0.01fF
C36356 OR2X1_LOC_680/A OR2X1_LOC_627/Y 0.03fF
C39336 VDD OR2X1_LOC_680/A 0.31fF
C39391 OR2X1_LOC_680/A OR2X1_LOC_677/Y 0.01fF
C39442 OR2X1_LOC_680/A OR2X1_LOC_616/Y 0.03fF
C39872 OR2X1_LOC_680/A AND2X1_LOC_834/a_8_24# 0.11fF
C43187 OR2X1_LOC_482/Y OR2X1_LOC_680/A 1.53fF
C47645 AND2X1_LOC_330/a_8_24# OR2X1_LOC_680/A 0.02fF
C55617 OR2X1_LOC_528/Y OR2X1_LOC_680/A 0.25fF
C57575 OR2X1_LOC_680/A VSS -4.91fF
C29397 VDD OR2X1_LOC_152/A 0.21fF
C56288 OR2X1_LOC_152/A VSS -0.04fF
C321 OR2X1_LOC_405/A OR2X1_LOC_317/a_8_216# 0.01fF
C7620 OR2X1_LOC_405/A OR2X1_LOC_539/Y 0.03fF
C8514 OR2X1_LOC_405/A OR2X1_LOC_493/A 0.08fF
C9123 OR2X1_LOC_405/A AND2X1_LOC_406/a_8_24# 0.26fF
C14392 OR2X1_LOC_405/A OR2X1_LOC_174/A 0.13fF
C16239 OR2X1_LOC_405/A AND2X1_LOC_109/a_8_24# 0.01fF
C18241 OR2X1_LOC_405/A AND2X1_LOC_314/a_8_24# 0.02fF
C20179 OR2X1_LOC_405/A AND2X1_LOC_406/a_36_24# 0.06fF
C23813 OR2X1_LOC_405/A OR2X1_LOC_317/A 0.01fF
C24185 OR2X1_LOC_405/A OR2X1_LOC_538/A 0.03fF
C24265 OR2X1_LOC_405/A OR2X1_LOC_802/A 0.02fF
C25015 OR2X1_LOC_405/A OR2X1_LOC_623/B 0.03fF
C26348 OR2X1_LOC_405/A OR2X1_LOC_592/A 0.09fF
C33891 OR2X1_LOC_405/A OR2X1_LOC_475/B 0.09fF
C37967 OR2X1_LOC_653/B OR2X1_LOC_405/A 0.03fF
C39717 OR2X1_LOC_405/A OR2X1_LOC_729/a_8_216# 0.01fF
C40140 OR2X1_LOC_405/A OR2X1_LOC_778/a_8_216# 0.03fF
C40415 OR2X1_LOC_405/A AND2X1_LOC_432/a_8_24# 0.01fF
C40625 OR2X1_LOC_405/A OR2X1_LOC_798/Y 0.03fF
C43692 OR2X1_LOC_405/A OR2X1_LOC_216/A 0.02fF
C44571 OR2X1_LOC_405/A OR2X1_LOC_447/A 0.01fF
C45111 OR2X1_LOC_405/A AND2X1_LOC_491/a_8_24# 0.01fF
C46304 OR2X1_LOC_405/A OR2X1_LOC_802/a_8_216# 0.06fF
C52855 OR2X1_LOC_405/A AND2X1_LOC_680/a_8_24# 0.02fF
C53595 OR2X1_LOC_405/A AND2X1_LOC_492/a_8_24# 0.01fF
C53820 OR2X1_LOC_405/A OR2X1_LOC_317/B 0.03fF
C54813 OR2X1_LOC_405/A OR2X1_LOC_473/a_8_216# 0.01fF
C56207 OR2X1_LOC_405/A OR2X1_LOC_449/B 0.07fF
C8248 OR2X1_LOC_497/a_8_216# OR2X1_LOC_184/Y 0.16fF
C11223 OR2X1_LOC_262/a_8_216# OR2X1_LOC_72/Y 0.01fF
C16739 OR2X1_LOC_262/a_36_216# OR2X1_LOC_72/Y 0.01fF
C10557 AND2X1_LOC_778/a_8_24# AND2X1_LOC_778/Y 0.08fF
C1083 OR2X1_LOC_678/a_8_216# OR2X1_LOC_713/A 0.01fF
C3202 OR2X1_LOC_307/A OR2X1_LOC_713/A 0.03fF
C10373 OR2X1_LOC_308/A OR2X1_LOC_713/A 0.01fF
C36261 OR2X1_LOC_834/a_8_216# OR2X1_LOC_713/A 0.01fF
C36365 AND2X1_LOC_697/a_8_24# OR2X1_LOC_713/A 0.02fF
C46154 OR2X1_LOC_834/A OR2X1_LOC_713/A 0.01fF
C52166 OR2X1_LOC_308/a_8_216# OR2X1_LOC_713/A 0.02fF
C8527 OR2X1_LOC_711/B AND2X1_LOC_698/a_8_24# 0.01fF
C45670 OR2X1_LOC_709/B OR2X1_LOC_711/B 0.83fF
C10394 AND2X1_LOC_832/a_8_24# OR2X1_LOC_589/Y 0.24fF
C15687 OR2X1_LOC_424/Y OR2X1_LOC_589/Y 0.07fF
C48689 VDD OR2X1_LOC_589/Y 0.26fF
C50690 OR2X1_LOC_589/Y AND2X1_LOC_592/a_8_24# -0.01fF
C56248 OR2X1_LOC_589/Y VSS 0.16fF
C13987 OR2X1_LOC_58/Y OR2X1_LOC_32/a_8_216# 0.01fF
C14854 OR2X1_LOC_58/Y OR2X1_LOC_60/a_8_216# 0.01fF
C26080 OR2X1_LOC_316/a_8_216# OR2X1_LOC_58/Y 0.01fF
C52670 OR2X1_LOC_58/Y OR2X1_LOC_316/Y 0.01fF
C3995 OR2X1_LOC_615/Y OR2X1_LOC_754/a_8_216# 0.41fF
C7044 OR2X1_LOC_615/Y AND2X1_LOC_790/a_8_24# 0.03fF
C7767 OR2X1_LOC_252/Y OR2X1_LOC_615/Y 0.02fF
C12445 AND2X1_LOC_631/a_8_24# OR2X1_LOC_615/Y 0.02fF
C23706 OR2X1_LOC_615/Y AND2X1_LOC_790/a_36_24# 0.01fF
C35325 AND2X1_LOC_483/a_8_24# OR2X1_LOC_615/Y -0.00fF
C52179 OR2X1_LOC_615/Y OR2X1_LOC_754/Y 0.02fF
C8399 OR2X1_LOC_497/Y OR2X1_LOC_184/a_8_216# 0.04fF
C10262 OR2X1_LOC_497/a_36_216# OR2X1_LOC_497/Y 0.01fF
C11309 OR2X1_LOC_497/Y AND2X1_LOC_227/a_8_24# 0.01fF
C13903 OR2X1_LOC_497/Y OR2X1_LOC_184/a_36_216# 0.01fF
C45185 OR2X1_LOC_497/Y OR2X1_LOC_224/Y 0.05fF
C55354 OR2X1_LOC_497/a_8_216# OR2X1_LOC_497/Y -0.02fF
C46237 OR2X1_LOC_320/Y OR2X1_LOC_321/a_8_216# 0.46fF
C8367 OR2X1_LOC_396/a_8_216# OR2X1_LOC_396/Y -0.00fF
C50420 OR2X1_LOC_39/Y OR2X1_LOC_39/a_8_216# 0.01fF
C7630 OR2X1_LOC_69/Y OR2X1_LOC_393/a_8_216# 0.04fF
C28884 OR2X1_LOC_69/a_8_216# OR2X1_LOC_69/Y 0.02fF
C16907 OR2X1_LOC_754/Y AND2X1_LOC_790/a_8_24# 0.23fF
C28959 VDD OR2X1_LOC_754/Y 0.16fF
C56494 OR2X1_LOC_754/Y VSS 0.07fF
C9173 OR2X1_LOC_528/Y OR2X1_LOC_627/Y 0.03fF
C19970 OR2X1_LOC_617/a_8_216# OR2X1_LOC_627/Y 0.01fF
C26645 OR2X1_LOC_252/a_8_216# OR2X1_LOC_627/Y 0.01fF
C36781 OR2X1_LOC_626/a_8_216# OR2X1_LOC_627/Y 0.01fF
C37596 OR2X1_LOC_252/Y OR2X1_LOC_627/Y 0.71fF
C49211 VDD OR2X1_LOC_627/Y 0.10fF
C56526 OR2X1_LOC_627/Y VSS 0.08fF
C56060 OR2X1_LOC_674/a_8_216# OR2X1_LOC_495/Y 0.01fF
C45181 OR2X1_LOC_145/a_8_216# OR2X1_LOC_146/Y 0.40fF
C3915 OR2X1_LOC_311/Y OR2X1_LOC_829/a_8_216# 0.01fF
C17152 OR2X1_LOC_311/Y AND2X1_LOC_539/a_8_24# 0.01fF
C22757 OR2X1_LOC_311/Y AND2X1_LOC_538/a_8_24# 0.01fF
C32604 OR2X1_LOC_311/Y AND2X1_LOC_802/Y 0.02fF
C36160 OR2X1_LOC_311/Y AND2X1_LOC_855/a_8_24# 0.01fF
C38062 OR2X1_LOC_311/Y AND2X1_LOC_809/a_8_24# 0.01fF
C45865 OR2X1_LOC_311/Y OR2X1_LOC_13/a_8_216# 0.01fF
C22527 OR2X1_LOC_536/Y OR2X1_LOC_385/Y 0.10fF
C27965 AND2X1_LOC_537/a_8_24# OR2X1_LOC_385/Y 0.05fF
C28460 OR2X1_LOC_385/Y OR2X1_LOC_586/a_8_216# 0.03fF
C33947 OR2X1_LOC_385/Y OR2X1_LOC_586/a_36_216# 0.01fF
C35557 VDD OR2X1_LOC_385/Y 0.17fF
C35695 OR2X1_LOC_385/Y AND2X1_LOC_389/a_8_24# 0.01fF
C57600 OR2X1_LOC_385/Y VSS 0.12fF
C48227 OR2X1_LOC_316/Y OR2X1_LOC_27/Y 0.07fF
C55444 AND2X1_LOC_462/a_8_24# OR2X1_LOC_27/Y 0.01fF
C37443 OR2X1_LOC_316/Y OR2X1_LOC_595/Y 0.02fF
C27614 OR2X1_LOC_669/A AND2X1_LOC_668/a_8_24# 0.11fF
C39057 OR2X1_LOC_669/A OR2X1_LOC_669/a_8_216# 0.47fF
C57335 OR2X1_LOC_669/A VSS 0.26fF
C11522 OR2X1_LOC_280/a_8_216# OR2X1_LOC_237/Y 0.01fF
C20852 OR2X1_LOC_237/a_8_216# OR2X1_LOC_237/Y 0.01fF
C37301 OR2X1_LOC_495/a_8_216# OR2X1_LOC_237/Y 0.01fF
C37407 OR2X1_LOC_237/Y OR2X1_LOC_238/a_8_216# 0.39fF
C52411 OR2X1_LOC_83/Y OR2X1_LOC_81/a_8_216# 0.04fF
C30802 OR2X1_LOC_106/Y OR2X1_LOC_67/A 0.01fF
C33424 OR2X1_LOC_122/a_8_216# OR2X1_LOC_67/A 0.01fF
C35477 OR2X1_LOC_106/a_8_216# OR2X1_LOC_67/A 0.01fF
C55665 OR2X1_LOC_122/Y OR2X1_LOC_67/A 0.01fF
C30759 OR2X1_LOC_680/a_8_216# OR2X1_LOC_677/Y 0.01fF
C31440 OR2X1_LOC_677/Y AND2X1_LOC_678/a_8_24# 0.11fF
C40999 OR2X1_LOC_677/a_8_216# OR2X1_LOC_677/Y 0.01fF
C49694 OR2X1_LOC_526/Y OR2X1_LOC_677/Y 0.44fF
C52183 VDD OR2X1_LOC_677/Y 0.28fF
C52744 OR2X1_LOC_677/Y AND2X1_LOC_834/a_8_24# 0.04fF
C57527 OR2X1_LOC_677/Y VSS 0.20fF
C3704 VDD OR2X1_LOC_290/Y 0.15fF
C9347 OR2X1_LOC_290/Y OR2X1_LOC_316/Y 0.02fF
C17033 OR2X1_LOC_290/Y AND2X1_LOC_334/a_8_24# -0.00fF
C35169 OR2X1_LOC_290/Y AND2X1_LOC_634/a_8_24# 0.24fF
C57694 OR2X1_LOC_290/Y VSS 0.19fF
C19721 OR2X1_LOC_176/Y AND2X1_LOC_799/a_8_24# 0.11fF
C25230 OR2X1_LOC_176/Y AND2X1_LOC_802/B 0.01fF
C9244 AND2X1_LOC_533/a_36_24# OR2X1_LOC_356/A 0.06fF
C54300 AND2X1_LOC_533/a_8_24# OR2X1_LOC_356/A 0.24fF
C3853 OR2X1_LOC_448/Y OR2X1_LOC_779/a_8_216# 0.43fF
C12932 OR2X1_LOC_475/B AND2X1_LOC_406/a_8_24# 0.01fF
C22021 OR2X1_LOC_833/B OR2X1_LOC_629/B 0.07fF
C56691 OR2X1_LOC_629/B VSS 0.19fF
C36794 OR2X1_LOC_489/B OR2X1_LOC_489/a_8_216# 0.05fF
C56792 OR2X1_LOC_489/B VSS 0.22fF
C32619 AND2X1_LOC_314/a_8_24# OR2X1_LOC_447/A 0.20fF
C55607 VDD OR2X1_LOC_447/A 0.21fF
C57164 OR2X1_LOC_447/A VSS 0.15fF
C12278 OR2X1_LOC_837/A OR2X1_LOC_837/a_8_216# 0.02fF
C26605 VDD OR2X1_LOC_837/A 0.21fF
C57484 OR2X1_LOC_837/A VSS 0.14fF
C48751 OR2X1_LOC_128/B OR2X1_LOC_342/a_8_216# 0.47fF
C34926 AND2X1_LOC_178/a_8_24# OR2X1_LOC_192/B 0.21fF
C35265 OR2X1_LOC_98/A OR2X1_LOC_98/a_8_216# 0.47fF
C52176 VDD OR2X1_LOC_98/A -0.00fF
C57592 OR2X1_LOC_98/A VSS 0.15fF
C9149 AND2X1_LOC_183/a_36_24# OR2X1_LOC_190/A 0.01fF
C14377 OR2X1_LOC_190/A OR2X1_LOC_254/B 0.09fF
C37670 AND2X1_LOC_183/a_8_24# OR2X1_LOC_190/A 0.04fF
C42438 OR2X1_LOC_190/A OR2X1_LOC_254/a_8_216# 0.03fF
C48147 OR2X1_LOC_190/A OR2X1_LOC_254/a_36_216# 0.02fF
C10796 AND2X1_LOC_437/a_8_24# OR2X1_LOC_788/B 0.02fF
C13411 AND2X1_LOC_166/a_8_24# OR2X1_LOC_788/B 0.02fF
C26345 OR2X1_LOC_788/B OR2X1_LOC_535/a_8_216# 0.01fF
C19503 OR2X1_LOC_653/B OR2X1_LOC_436/a_8_216# 0.47fF
C14783 OR2X1_LOC_605/B AND2X1_LOC_604/a_8_24# 0.02fF
C28372 OR2X1_LOC_605/B AND2X1_LOC_603/a_8_24# 0.01fF
C29857 OR2X1_LOC_391/A OR2X1_LOC_558/A 0.03fF
C52616 AND2X1_LOC_494/a_8_24# OR2X1_LOC_558/A 0.01fF
C17444 OR2X1_LOC_193/A AND2X1_LOC_16/a_8_24# 0.37fF
C25508 OR2X1_LOC_538/a_8_216# OR2X1_LOC_193/A 0.01fF
C44394 OR2X1_LOC_193/A OR2X1_LOC_789/A 0.02fF
C48288 AND2X1_LOC_135/a_8_24# OR2X1_LOC_193/A 0.14fF
C57909 OR2X1_LOC_318/A VSS 0.21fF
C30848 OR2X1_LOC_678/a_8_216# OR2X1_LOC_678/Y 0.01fF
C9271 VDD OR2X1_LOC_260/Y 0.06fF
C20406 OR2X1_LOC_791/B OR2X1_LOC_260/Y 0.24fF
C54080 OR2X1_LOC_260/Y AND2X1_LOC_261/a_8_24# 0.01fF
C57499 OR2X1_LOC_260/Y VSS 0.10fF
C22667 OR2X1_LOC_140/A OR2X1_LOC_66/Y 0.01fF
C25774 OR2X1_LOC_115/a_8_216# OR2X1_LOC_140/A 0.47fF
C33538 AND2X1_LOC_385/a_8_24# OR2X1_LOC_537/A 0.02fF
C39038 OR2X1_LOC_389/B OR2X1_LOC_537/A 0.16fF
C57680 OR2X1_LOC_537/A VSS -0.01fF
C12494 AND2X1_LOC_229/a_8_24# OR2X1_LOC_231/B 0.01fF
C55548 OR2X1_LOC_440/B AND2X1_LOC_437/a_8_24# 0.01fF
C3801 OR2X1_LOC_254/B OR2X1_LOC_254/A 0.09fF
C19105 OR2X1_LOC_254/B OR2X1_LOC_147/B 0.03fF
C37294 OR2X1_LOC_254/B OR2X1_LOC_483/a_8_216# 0.01fF
C49045 OR2X1_LOC_254/B OR2X1_LOC_254/a_8_216# 0.01fF
C54406 OR2X1_LOC_254/B AND2X1_LOC_253/a_8_24# 0.01fF
C57634 OR2X1_LOC_254/B VSS 0.28fF
C16114 AND2X1_LOC_108/a_8_24# OR2X1_LOC_346/A 0.08fF
C1938 OR2X1_LOC_114/B AND2X1_LOC_184/a_8_24# 0.01fF
C9886 OR2X1_LOC_114/B AND2X1_LOC_497/a_8_24# 0.01fF
C20197 OR2X1_LOC_114/B AND2X1_LOC_248/a_8_24# 0.01fF
C33773 OR2X1_LOC_114/a_8_216# OR2X1_LOC_114/B 0.05fF
C46135 OR2X1_LOC_114/B AND2X1_LOC_295/a_8_24# 0.01fF
C49776 OR2X1_LOC_114/B AND2X1_LOC_292/a_8_24# 0.05fF
C52218 OR2X1_LOC_114/B AND2X1_LOC_297/a_8_24# 0.01fF
C16396 OR2X1_LOC_833/B AND2X1_LOC_626/a_8_24# 0.02fF
C27464 OR2X1_LOC_833/B AND2X1_LOC_626/a_36_24# 0.01fF
C33015 OR2X1_LOC_473/a_8_216# OR2X1_LOC_493/A 0.02fF
C11062 OR2X1_LOC_702/A AND2X1_LOC_173/a_8_24# 0.02fF
C24474 OR2X1_LOC_702/A OR2X1_LOC_332/a_8_216# 0.07fF
C35919 OR2X1_LOC_702/A OR2X1_LOC_138/a_8_216# 0.09fF
C41449 OR2X1_LOC_702/A OR2X1_LOC_138/a_36_216# 0.03fF
C51929 OR2X1_LOC_538/a_8_216# OR2X1_LOC_702/A 0.01fF
C11085 AND2X1_LOC_89/a_8_24# OR2X1_LOC_97/B 0.02fF
C22196 OR2X1_LOC_97/B AND2X1_LOC_89/a_36_24# 0.01fF
C34250 VDD OR2X1_LOC_97/B 0.21fF
C57344 OR2X1_LOC_97/B VSS 0.20fF
C10160 OR2X1_LOC_76/A AND2X1_LOC_604/a_36_24# 0.01fF
C46054 AND2X1_LOC_75/a_8_24# OR2X1_LOC_76/A 0.10fF
C55248 OR2X1_LOC_76/A AND2X1_LOC_604/a_8_24# 0.02fF
C55591 OR2X1_LOC_76/A OR2X1_LOC_301/a_8_216# 0.03fF
C27675 AND2X1_LOC_395/a_8_24# OR2X1_LOC_401/B 0.01fF
C45378 AND2X1_LOC_766/a_8_24# OR2X1_LOC_401/B 0.20fF
C4724 OR2X1_LOC_791/B OR2X1_LOC_287/a_8_216# 0.48fF
C9375 OR2X1_LOC_791/B OR2X1_LOC_260/a_8_216# 0.01fF
C26367 OR2X1_LOC_791/B AND2X1_LOC_281/a_8_24# 0.01fF
C37348 OR2X1_LOC_791/B OR2X1_LOC_285/B 0.01fF
C56201 OR2X1_LOC_791/B AND2X1_LOC_282/a_8_24# 0.01fF
C34953 AND2X1_LOC_744/a_8_24# OR2X1_LOC_712/B 0.01fF
C39966 OR2X1_LOC_450/A OR2X1_LOC_712/B 0.03fF
C46105 AND2X1_LOC_424/a_8_24# OR2X1_LOC_712/B 0.01fF
C17524 OR2X1_LOC_698/a_8_216# AND2X1_LOC_793/B 0.02fF
C23127 OR2X1_LOC_698/a_36_216# AND2X1_LOC_793/B 0.02fF
C50575 AND2X1_LOC_846/a_8_24# AND2X1_LOC_793/B 0.04fF
C31213 OR2X1_LOC_536/Y AND2X1_LOC_537/a_8_24# 0.23fF
C38817 VDD OR2X1_LOC_536/Y 0.16fF
C57619 OR2X1_LOC_536/Y VSS 0.07fF
C21785 OR2X1_LOC_13/Y OR2X1_LOC_311/a_8_216# 0.01fF
C34985 OR2X1_LOC_13/a_8_216# OR2X1_LOC_13/Y 0.01fF
C53383 AND2X1_LOC_195/a_8_24# OR2X1_LOC_13/Y 0.01fF
C54492 OR2X1_LOC_41/a_8_216# OR2X1_LOC_13/Y 0.01fF
C29790 OR2X1_LOC_679/A AND2X1_LOC_147/a_8_24# 0.21fF
C56887 OR2X1_LOC_261/A VSS 0.02fF
C35053 OR2X1_LOC_603/a_8_216# OR2X1_LOC_603/Y -0.00fF
C25398 VDD OR2X1_LOC_380/A 0.03fF
C35531 OR2X1_LOC_380/A OR2X1_LOC_380/a_8_216# 0.08fF
C57536 OR2X1_LOC_380/A VSS 0.16fF
C11833 OR2X1_LOC_494/Y OR2X1_LOC_667/a_8_216# 0.01fF
C1606 VDD OR2X1_LOC_316/Y 0.62fF
C1696 OR2X1_LOC_315/Y OR2X1_LOC_316/Y 0.05fF
C4227 OR2X1_LOC_316/Y AND2X1_LOC_831/a_8_24# 0.01fF
C7995 AND2X1_LOC_301/a_8_24# OR2X1_LOC_316/Y 0.01fF
C12759 OR2X1_LOC_316/Y AND2X1_LOC_318/a_8_24# 0.11fF
C14965 AND2X1_LOC_334/a_8_24# OR2X1_LOC_316/Y 0.01fF
C16662 OR2X1_LOC_316/Y OR2X1_LOC_75/a_8_216# 0.01fF
C33096 OR2X1_LOC_316/Y AND2X1_LOC_634/a_8_24# 0.01fF
C33199 OR2X1_LOC_316/Y OR2X1_LOC_75/Y 0.03fF
C36896 OR2X1_LOC_316/Y OR2X1_LOC_27/a_8_216# 0.01fF
C54396 OR2X1_LOC_290/a_8_216# OR2X1_LOC_316/Y 0.01fF
C57252 OR2X1_LOC_316/Y VSS 0.10fF
C19082 OR2X1_LOC_395/Y OR2X1_LOC_396/a_8_216# 0.40fF
C10505 OR2X1_LOC_755/a_8_216# OR2X1_LOC_755/Y -0.00fF
C1299 OR2X1_LOC_700/Y OR2X1_LOC_701/a_8_216# 0.02fF
C23702 OR2X1_LOC_89/a_8_216# OR2X1_LOC_89/Y 0.01fF
C56754 OR2X1_LOC_89/Y VSS 0.11fF
C42665 OR2X1_LOC_75/a_8_216# OR2X1_LOC_75/Y 0.12fF
C11728 OR2X1_LOC_437/a_8_216# OR2X1_LOC_437/Y 0.05fF
C35647 OR2X1_LOC_81/Y OR2X1_LOC_81/a_8_216# 0.01fF
C698 OR2X1_LOC_528/Y OR2X1_LOC_252/Y 0.12fF
C895 OR2X1_LOC_252/Y AND2X1_LOC_483/a_8_24# 0.09fF
C32079 OR2X1_LOC_252/Y AND2X1_LOC_254/a_8_24# 0.10fF
C34342 OR2X1_LOC_252/Y OR2X1_LOC_627/a_8_216# 0.01fF
C40582 VDD OR2X1_LOC_252/Y -0.00fF
C44467 OR2X1_LOC_482/Y OR2X1_LOC_252/Y 0.01fF
C57309 OR2X1_LOC_252/Y VSS -0.09fF
C4437 OR2X1_LOC_178/a_8_216# OR2X1_LOC_108/Y -0.01fF
C14674 OR2X1_LOC_492/a_8_216# OR2X1_LOC_108/Y 0.06fF
C23273 OR2X1_LOC_179/a_8_216# OR2X1_LOC_108/Y 0.02fF
C25707 OR2X1_LOC_108/a_8_216# OR2X1_LOC_108/Y 0.05fF
C31203 OR2X1_LOC_108/a_36_216# OR2X1_LOC_108/Y 0.01fF
C33734 OR2X1_LOC_491/a_8_216# OR2X1_LOC_108/Y 0.07fF
C39053 OR2X1_LOC_108/Y OR2X1_LOC_224/a_8_216# 0.02fF
C50841 OR2X1_LOC_108/Y OR2X1_LOC_183/a_8_216# 0.03fF
C55804 OR2X1_LOC_108/Y OR2X1_LOC_224/Y 0.01fF
C20648 OR2X1_LOC_482/Y OR2X1_LOC_666/a_8_216# 0.01fF
C35858 OR2X1_LOC_674/a_8_216# OR2X1_LOC_482/Y 0.03fF
C48758 OR2X1_LOC_482/a_8_216# OR2X1_LOC_482/Y 0.01fF
C3622 OR2X1_LOC_492/a_8_216# OR2X1_LOC_492/Y 0.01fF
C31265 OR2X1_LOC_135/Y AND2X1_LOC_138/a_8_24# 0.01fF
C42634 OR2X1_LOC_135/a_8_216# OR2X1_LOC_135/Y -0.01fF
C48344 OR2X1_LOC_135/a_36_216# OR2X1_LOC_135/Y 0.01fF
C48921 OR2X1_LOC_135/Y AND2X1_LOC_307/a_8_24# 0.01fF
C18443 OR2X1_LOC_521/Y OR2X1_LOC_521/a_8_216# -0.00fF
C13735 OR2X1_LOC_315/Y OR2X1_LOC_368/A 0.10fF
C14456 OR2X1_LOC_368/A AND2X1_LOC_457/a_8_24# 0.17fF
C34904 OR2X1_LOC_109/Y OR2X1_LOC_368/A 0.01fF
C47302 OR2X1_LOC_315/a_8_216# OR2X1_LOC_368/A 0.01fF
C13399 OR2X1_LOC_607/a_8_216# OR2X1_LOC_607/Y -0.00fF
C12207 OR2X1_LOC_528/Y OR2X1_LOC_616/Y 0.97fF
C20077 OR2X1_LOC_616/Y AND2X1_LOC_664/a_8_24# 0.03fF
C25577 OR2X1_LOC_616/Y AND2X1_LOC_621/a_8_24# 0.10fF
C29598 AND2X1_LOC_758/a_8_24# OR2X1_LOC_616/Y 0.01fF
C34248 AND2X1_LOC_756/a_8_24# OR2X1_LOC_616/Y 0.01fF
C41105 OR2X1_LOC_616/a_8_216# OR2X1_LOC_616/Y 0.02fF
C57233 OR2X1_LOC_616/Y VSS -0.21fF
C44060 VDD OR2X1_LOC_432/Y 0.16fF
C56625 OR2X1_LOC_432/Y VSS 0.35fF
C17052 OR2X1_LOC_496/Y AND2X1_LOC_778/a_8_24# 0.11fF
C30075 OR2X1_LOC_496/Y OR2X1_LOC_496/a_8_216# 0.01fF
C45384 OR2X1_LOC_482/a_8_216# OR2X1_LOC_666/Y 0.40fF
C26864 OR2X1_LOC_526/Y OR2X1_LOC_526/a_8_216# 0.01fF
C52196 OR2X1_LOC_526/Y OR2X1_LOC_485/a_8_216# 0.01fF
C11705 OR2X1_LOC_583/a_8_216# OR2X1_LOC_583/Y -0.00fF
C46357 OR2X1_LOC_32/Y OR2X1_LOC_58/a_36_216# 0.02fF
C41767 OR2X1_LOC_428/a_8_216# OR2X1_LOC_428/Y 0.01fF
C57012 OR2X1_LOC_428/Y VSS 0.01fF
C35219 VDD OR2X1_LOC_224/Y 0.18fF
C57052 OR2X1_LOC_224/Y VSS 0.08fF
C41058 OR2X1_LOC_298/Y OR2X1_LOC_298/a_8_216# 0.02fF
C57545 OR2X1_LOC_298/Y VSS 0.12fF
C42712 OR2X1_LOC_600/a_8_216# OR2X1_LOC_600/Y -0.00fF
C16409 OR2X1_LOC_368/a_8_216# OR2X1_LOC_109/Y 0.03fF
C18103 OR2X1_LOC_109/Y AND2X1_LOC_457/a_8_24# 0.02fF
C22029 OR2X1_LOC_368/a_36_216# OR2X1_LOC_109/Y 0.01fF
C27549 OR2X1_LOC_109/a_8_216# OR2X1_LOC_109/Y 0.01fF
C30066 AND2X1_LOC_543/a_8_24# OR2X1_LOC_109/Y 0.02fF
C46693 OR2X1_LOC_109/Y AND2X1_LOC_325/a_8_24# 0.01fF
C8890 AND2X1_LOC_543/a_8_24# OR2X1_LOC_315/Y 0.08fF
C29569 OR2X1_LOC_315/a_8_216# OR2X1_LOC_315/Y 0.03fF
C35055 OR2X1_LOC_315/a_36_216# OR2X1_LOC_315/Y 0.03fF
C44601 OR2X1_LOC_399/a_8_216# OR2X1_LOC_399/Y -0.00fF
C33499 OR2X1_LOC_755/a_8_216# OR2X1_LOC_757/Y 0.40fF
C6769 OR2X1_LOC_701/Y OR2X1_LOC_701/a_8_216# 0.05fF
C38782 VDD OR2X1_LOC_744/Y 0.06fF
C46959 OR2X1_LOC_744/Y AND2X1_LOC_780/a_8_24# 0.01fF
C56620 OR2X1_LOC_744/Y VSS 0.10fF
C8139 OR2X1_LOC_45/Y OR2X1_LOC_431/a_8_216# 0.03fF
C16094 OR2X1_LOC_45/Y OR2X1_LOC_45/a_8_216# 0.03fF
C43196 OR2X1_LOC_45/Y AND2X1_LOC_434/a_8_24# 0.11fF
C43908 OR2X1_LOC_45/Y OR2X1_LOC_172/a_8_216# -0.03fF
C54348 OR2X1_LOC_45/Y AND2X1_LOC_434/a_36_24# 0.01fF
C9493 OR2X1_LOC_280/Y OR2X1_LOC_279/Y 0.08fF
C23401 VDD OR2X1_LOC_279/Y 0.18fF
C35078 OR2X1_LOC_279/Y AND2X1_LOC_284/a_8_24# 0.04fF
C39542 OR2X1_LOC_279/a_8_216# OR2X1_LOC_279/Y 0.01fF
C57042 OR2X1_LOC_279/Y VSS 0.27fF
C21297 OR2X1_LOC_424/Y AND2X1_LOC_592/a_8_24# 0.10fF
C15792 OR2X1_LOC_485/Y OR2X1_LOC_526/a_8_216# 0.39fF
C40952 OR2X1_LOC_485/Y OR2X1_LOC_485/a_8_216# 0.01fF
C47544 OR2X1_LOC_485/Y OR2X1_LOC_484/a_8_216# 0.10fF
C23832 VDD OR2X1_LOC_825/Y -0.00fF
C23957 OR2X1_LOC_825/Y OR2X1_LOC_826/a_8_216# 0.41fF
C57551 OR2X1_LOC_825/Y VSS 0.21fF
C11731 OR2X1_LOC_122/Y OR2X1_LOC_106/a_8_216# 0.40fF
C4931 OR2X1_LOC_528/Y AND2X1_LOC_186/a_36_24# 0.01fF
C11692 OR2X1_LOC_528/a_8_216# OR2X1_LOC_528/Y 0.15fF
C24156 OR2X1_LOC_528/Y OR2X1_LOC_406/a_8_216# 0.01fF
C26106 OR2X1_LOC_505/a_8_216# OR2X1_LOC_528/Y 0.14fF
C35081 OR2X1_LOC_528/Y OR2X1_LOC_406/a_36_216# 0.01fF
C41565 OR2X1_LOC_528/Y AND2X1_LOC_621/a_8_24# 0.01fF
C46171 OR2X1_LOC_528/Y AND2X1_LOC_549/a_8_24# 0.04fF
C46183 OR2X1_LOC_528/Y AND2X1_LOC_506/a_8_24# 0.26fF
C50145 OR2X1_LOC_528/Y AND2X1_LOC_186/a_8_24# 0.16fF
C3677 OR2X1_LOC_524/Y OR2X1_LOC_745/a_8_216# 0.09fF
C14605 OR2X1_LOC_524/Y OR2X1_LOC_152/a_8_216# 0.15fF
C14727 OR2X1_LOC_524/Y OR2X1_LOC_745/a_36_216# 0.16fF
C20133 OR2X1_LOC_524/Y OR2X1_LOC_152/a_36_216# 0.17fF
C23718 OR2X1_LOC_524/Y OR2X1_LOC_441/a_8_216# 0.18fF
C29162 OR2X1_LOC_524/Y OR2X1_LOC_441/a_36_216# 0.14fF
C31379 OR2X1_LOC_524/Y OR2X1_LOC_438/a_8_216# 0.12fF
C35953 OR2X1_LOC_524/Y AND2X1_LOC_676/a_8_24# 0.29fF
C47209 OR2X1_LOC_524/Y AND2X1_LOC_676/a_36_24# 0.08fF
C14925 OR2X1_LOC_83/a_8_216# OR2X1_LOC_394/Y 0.01fF
C20328 OR2X1_LOC_394/Y OR2X1_LOC_394/a_8_216# 0.01fF
C33106 AND2X1_LOC_342/a_8_24# OR2X1_LOC_248/Y 0.10fF
C52710 VDD OR2X1_LOC_248/Y 0.23fF
C56954 OR2X1_LOC_248/Y VSS 0.38fF
C39780 OR2X1_LOC_612/a_8_216# OR2X1_LOC_612/B 0.05fF
C52849 AND2X1_LOC_610/a_8_24# OR2X1_LOC_612/B 0.01fF
C56974 OR2X1_LOC_612/B VSS 0.18fF
C4789 OR2X1_LOC_280/Y OR2X1_LOC_224/a_8_216# 0.03fF
C6705 OR2X1_LOC_280/Y AND2X1_LOC_489/a_8_24# 0.17fF
C7723 OR2X1_LOC_280/a_8_216# OR2X1_LOC_280/Y 0.01fF
C15840 OR2X1_LOC_280/Y OR2X1_LOC_224/a_36_216# 0.02fF
C17037 OR2X1_LOC_280/Y OR2X1_LOC_237/a_8_216# 0.01fF
C33677 OR2X1_LOC_280/Y OR2X1_LOC_238/a_8_216# 0.04fF
C50140 OR2X1_LOC_280/Y AND2X1_LOC_284/a_8_24# 0.11fF
C7893 VDD OR2X1_LOC_695/Y 0.16fF
C25322 OR2X1_LOC_695/Y AND2X1_LOC_707/a_8_24# 0.23fF
C57629 OR2X1_LOC_695/Y VSS 0.07fF
C12244 OR2X1_LOC_106/Y AND2X1_LOC_115/a_8_24# 0.09fF
C28601 AND2X1_LOC_361/a_8_24# OR2X1_LOC_106/Y 0.04fF
C36015 OR2X1_LOC_106/Y AND2X1_LOC_116/a_8_24# 0.07fF
C45213 AND2X1_LOC_361/a_36_24# OR2X1_LOC_106/Y 0.01fF
C4917 OR2X1_LOC_107/a_8_216# OR2X1_LOC_103/Y 0.01fF
C13963 OR2X1_LOC_103/Y AND2X1_LOC_113/a_8_24# 0.01fF
C38836 AND2X1_LOC_361/a_8_24# OR2X1_LOC_103/Y 0.01fF
C17274 VDD OR2X1_LOC_330/Y 0.16fF
C44088 OR2X1_LOC_330/Y AND2X1_LOC_331/a_8_24# 0.23fF
C57789 OR2X1_LOC_330/Y VSS 0.07fF
C2825 OR2X1_LOC_450/A OR2X1_LOC_450/a_8_216# 0.01fF
C2913 OR2X1_LOC_450/A AND2X1_LOC_695/a_8_24# 0.24fF
C8883 OR2X1_LOC_450/A OR2X1_LOC_449/B 0.46fF
C17968 OR2X1_LOC_450/A OR2X1_LOC_707/a_8_216# 0.03fF
C19465 OR2X1_LOC_450/A AND2X1_LOC_695/a_36_24# 0.01fF
C50078 VDD OR2X1_LOC_450/A 0.21fF
C57636 OR2X1_LOC_450/A VSS 0.10fF
C14861 OR2X1_LOC_544/A AND2X1_LOC_438/a_8_24# 0.09fF
C9287 OR2X1_LOC_605/A AND2X1_LOC_604/a_8_24# 0.10fF
C20317 OR2X1_LOC_605/A AND2X1_LOC_604/a_36_24# 0.01fF
C34633 OR2X1_LOC_335/a_8_216# OR2X1_LOC_605/A 0.47fF
C44503 OR2X1_LOC_501/B OR2X1_LOC_630/a_8_216# 0.05fF
C5935 VDD OR2X1_LOC_434/A -0.00fF
C35225 OR2X1_LOC_174/A OR2X1_LOC_434/A 0.28fF
C55897 OR2X1_LOC_333/B OR2X1_LOC_434/A 0.01fF
C56849 OR2X1_LOC_434/A VSS 0.31fF
C20334 OR2X1_LOC_633/B AND2X1_LOC_262/a_8_24# 0.01fF
C23490 AND2X1_LOC_118/a_8_24# OR2X1_LOC_633/B 0.01fF
C35157 OR2X1_LOC_633/a_8_216# OR2X1_LOC_633/B 0.02fF
C36531 AND2X1_LOC_117/a_8_24# OR2X1_LOC_633/B 0.01fF
C40668 OR2X1_LOC_633/a_36_216# OR2X1_LOC_633/B 0.02fF
C51570 AND2X1_LOC_81/a_8_24# OR2X1_LOC_633/B 0.01fF
C10699 OR2X1_LOC_835/B AND2X1_LOC_822/a_8_24# 0.04fF
C28143 OR2X1_LOC_835/B AND2X1_LOC_821/a_8_24# 0.01fF
C8681 VDD OR2X1_LOC_317/B 0.03fF
C23991 OR2X1_LOC_317/a_8_216# OR2X1_LOC_317/B 0.07fF
C26743 OR2X1_LOC_317/B OR2X1_LOC_704/a_8_216# 0.10fF
C47468 OR2X1_LOC_317/A OR2X1_LOC_317/B 0.04fF
C56423 OR2X1_LOC_317/B VSS 0.02fF
C1091 OR2X1_LOC_855/a_8_216# OR2X1_LOC_637/A 0.47fF
C8029 OR2X1_LOC_379/Y OR2X1_LOC_637/A 0.01fF
C39655 OR2X1_LOC_637/A AND2X1_LOC_829/a_8_24# 0.05fF
C45272 OR2X1_LOC_637/A OR2X1_LOC_855/A 0.19fF
C57290 OR2X1_LOC_637/A VSS -0.06fF
C7012 VDD OR2X1_LOC_758/Y 0.15fF
C23666 OR2X1_LOC_758/Y AND2X1_LOC_759/a_8_24# 0.23fF
C57827 OR2X1_LOC_758/Y VSS -0.01fF
C3414 OR2X1_LOC_227/a_36_216# OR2X1_LOC_641/A 0.02fF
C36240 AND2X1_LOC_505/a_8_24# OR2X1_LOC_641/A 0.02fF
C52252 OR2X1_LOC_267/a_8_216# OR2X1_LOC_641/A 0.08fF
C54016 OR2X1_LOC_227/a_8_216# OR2X1_LOC_641/A 0.03fF
C20336 AND2X1_LOC_118/a_8_24# OR2X1_LOC_786/A 0.08fF
C40125 OR2X1_LOC_266/a_8_216# OR2X1_LOC_786/A 0.05fF
C48512 AND2X1_LOC_81/a_8_24# OR2X1_LOC_786/A 0.01fF
C1423 OR2X1_LOC_444/B AND2X1_LOC_442/a_8_24# 0.01fF
C39975 OR2X1_LOC_545/B AND2X1_LOC_442/a_8_24# 0.20fF
C52767 AND2X1_LOC_524/a_8_24# OR2X1_LOC_545/B 0.01fF
C19700 AND2X1_LOC_108/a_8_24# OR2X1_LOC_346/B 0.01fF
C27085 OR2X1_LOC_346/B AND2X1_LOC_295/a_8_24# 0.20fF
C17749 OR2X1_LOC_673/B AND2X1_LOC_670/a_8_24# 0.04fF
C26099 OR2X1_LOC_673/B OR2X1_LOC_673/a_8_216# 0.05fF
C57773 OR2X1_LOC_673/B VSS -0.11fF
C22585 AND2X1_LOC_166/a_8_24# OR2X1_LOC_169/B 0.01fF
C8619 OR2X1_LOC_610/Y AND2X1_LOC_612/a_8_24# 0.23fF
C50189 VDD OR2X1_LOC_610/Y 0.12fF
C56870 OR2X1_LOC_610/Y VSS 0.06fF
C20893 AND2X1_LOC_41/Y OR2X1_LOC_195/a_8_216# 0.07fF
C37991 AND2X1_LOC_7/Y AND2X1_LOC_41/Y 0.02fF
C56333 AND2X1_LOC_41/Y VSS 0.36fF
C9663 OR2X1_LOC_333/B OR2X1_LOC_333/a_8_216# 0.03fF
C20705 OR2X1_LOC_333/B OR2X1_LOC_333/a_36_216# 0.02fF
C28527 AND2X1_LOC_171/a_8_24# OR2X1_LOC_333/B 0.01fF
C50416 OR2X1_LOC_333/B AND2X1_LOC_431/a_8_24# 0.01fF
C7150 OR2X1_LOC_848/a_8_216# OR2X1_LOC_391/A 0.03fF
C15322 AND2X1_LOC_494/a_8_24# OR2X1_LOC_391/A 0.23fF
C26358 AND2X1_LOC_494/a_36_24# OR2X1_LOC_391/A -0.01fF
C50524 VDD OR2X1_LOC_391/A 0.21fF
C56705 OR2X1_LOC_391/A VSS -0.56fF
C20117 OR2X1_LOC_549/B OR2X1_LOC_549/a_8_216# 0.07fF
C58130 OR2X1_LOC_549/B VSS 0.27fF
C18485 AND2X1_LOC_745/a_8_24# OR2X1_LOC_781/B 0.01fF
C23054 AND2X1_LOC_393/a_8_24# OR2X1_LOC_400/B 0.01fF
C25335 OR2X1_LOC_769/A VDD 0.21fF
C58083 OR2X1_LOC_769/A VSS 0.20fF
C18202 AND2X1_LOC_751/a_8_24# OR2X1_LOC_789/A 0.01fF
C56267 OR2X1_LOC_789/A VSS 0.14fF
C22656 OR2X1_LOC_846/a_8_216# OR2X1_LOC_846/B 0.02fF
C31915 OR2X1_LOC_846/B AND2X1_LOC_816/a_8_24# 0.21fF
C33590 OR2X1_LOC_846/a_36_216# OR2X1_LOC_846/B 0.01fF
C51732 OR2X1_LOC_846/B OR2X1_LOC_557/a_8_216# 0.12fF
C54832 VDD OR2X1_LOC_846/B 0.27fF
C56879 OR2X1_LOC_846/B VSS 0.36fF
C4662 OR2X1_LOC_285/a_8_216# OR2X1_LOC_285/B 0.03fF
C19204 OR2X1_LOC_285/B AND2X1_LOC_282/a_8_24# 0.20fF
C26295 VDD OR2X1_LOC_285/B 0.21fF
C56941 OR2X1_LOC_285/B VSS 0.21fF
C42999 AND2X1_LOC_7/a_8_24# AND2X1_LOC_7/Y 0.01fF
C1297 AND2X1_LOC_665/a_8_24# OR2X1_LOC_719/B 0.01fF
C28379 AND2X1_LOC_72/a_8_24# OR2X1_LOC_719/B 0.04fF
C44961 AND2X1_LOC_72/a_36_24# OR2X1_LOC_719/B 0.01fF
C53831 OR2X1_LOC_555/A AND2X1_LOC_257/a_8_24# 0.21fF
C6281 AND2X1_LOC_677/a_8_24# OR2X1_LOC_307/A 0.10fF
C10014 VDD OR2X1_LOC_307/A 0.21fF
C10866 OR2X1_LOC_834/A OR2X1_LOC_307/A 0.03fF
C24986 OR2X1_LOC_449/B OR2X1_LOC_307/A 0.03fF
C56615 OR2X1_LOC_307/A VSS 0.39fF
C6591 AND2X1_LOC_397/a_8_24# OR2X1_LOC_402/B 0.01fF
C2094 OR2X1_LOC_590/a_8_216# OR2X1_LOC_593/B 0.02fF
C9450 AND2X1_LOC_591/a_8_24# OR2X1_LOC_593/B 0.01fF
C19719 OR2X1_LOC_832/a_8_216# OR2X1_LOC_593/B 0.14fF
C25294 OR2X1_LOC_831/a_8_216# OR2X1_LOC_593/B 0.01fF
C26971 OR2X1_LOC_593/a_8_216# OR2X1_LOC_593/B 0.06fF
C2054 OR2X1_LOC_147/B OR2X1_LOC_254/A 0.10fF
C31818 OR2X1_LOC_254/a_8_216# OR2X1_LOC_254/A 0.47fF
C56664 OR2X1_LOC_254/A VSS 0.15fF
C2102 OR2X1_LOC_834/a_8_216# OR2X1_LOC_449/B 0.05fF
C11856 OR2X1_LOC_834/A OR2X1_LOC_449/B 0.03fF
C17009 OR2X1_LOC_168/a_8_216# OR2X1_LOC_449/B 0.01fF
C19947 OR2X1_LOC_450/a_8_216# OR2X1_LOC_449/B 0.01fF
C20026 AND2X1_LOC_695/a_8_24# OR2X1_LOC_449/B 0.04fF
C22511 OR2X1_LOC_832/a_8_216# OR2X1_LOC_449/B 0.07fF
C22701 AND2X1_LOC_680/a_8_24# OR2X1_LOC_449/B 0.03fF
C29746 OR2X1_LOC_449/B OR2X1_LOC_593/a_8_216# 0.06fF
C31111 OR2X1_LOC_780/a_8_216# OR2X1_LOC_449/B 0.01fF
C31443 OR2X1_LOC_449/B OR2X1_LOC_592/a_8_216# 0.03fF
C36480 AND2X1_LOC_695/a_36_24# OR2X1_LOC_449/B 0.01fF
C38247 AND2X1_LOC_165/a_8_24# OR2X1_LOC_449/B 0.01fF
C45462 OR2X1_LOC_449/B AND2X1_LOC_423/a_8_24# 0.07fF
C52434 OR2X1_LOC_592/A OR2X1_LOC_449/B 0.05fF
C2832 AND2X1_LOC_586/a_8_24# OR2X1_LOC_855/A 0.05fF
C38766 VDD OR2X1_LOC_855/A 0.21fF
C56697 OR2X1_LOC_855/A VSS 0.01fF
C42688 AND2X1_LOC_250/a_8_24# OR2X1_LOC_343/B 0.01fF
C11642 AND2X1_LOC_134/a_8_24# OR2X1_LOC_720/B 0.01fF
C34515 OR2X1_LOC_709/B OR2X1_LOC_709/a_8_216# 0.06fF
C48125 OR2X1_LOC_709/B AND2X1_LOC_698/a_8_24# 0.01fF
C58093 OR2X1_LOC_709/B VSS 0.10fF
C50564 OR2X1_LOC_113/A OR2X1_LOC_844/B 0.15fF
C57078 OR2X1_LOC_113/A VSS 0.21fF
C8330 OR2X1_LOC_703/B OR2X1_LOC_535/a_8_216# 0.19fF
C51500 OR2X1_LOC_703/B AND2X1_LOC_166/a_8_24# 0.02fF
C26744 VDD OR2X1_LOC_520/B -0.00fF
C51517 OR2X1_LOC_520/B OR2X1_LOC_520/a_8_216# 0.07fF
C52055 AND2X1_LOC_518/a_8_24# OR2X1_LOC_520/B 0.01fF
C57430 OR2X1_LOC_520/B VSS 0.24fF
C50182 OR2X1_LOC_317/a_8_216# OR2X1_LOC_317/A 0.47fF
C57476 OR2X1_LOC_317/A VSS 0.15fF
C5919 OR2X1_LOC_147/a_8_216# OR2X1_LOC_147/B 0.10fF
C19485 AND2X1_LOC_321/a_8_24# OR2X1_LOC_147/B 0.22fF
C23131 OR2X1_LOC_147/B OR2X1_LOC_543/a_8_216# 0.06fF
C25850 OR2X1_LOC_147/B AND2X1_LOC_315/a_8_24# 0.03fF
C27100 OR2X1_LOC_325/a_8_216# OR2X1_LOC_703/A 0.01fF
C11481 AND2X1_LOC_516/a_8_24# OR2X1_LOC_623/B 0.03fF
C36724 OR2X1_LOC_834/A OR2X1_LOC_623/B 0.03fF
C18683 AND2X1_LOC_497/a_8_24# OR2X1_LOC_844/B 0.01fF
C42637 OR2X1_LOC_114/a_8_216# OR2X1_LOC_844/B 0.01fF
C9617 AND2X1_LOC_60/a_8_24# OR2X1_LOC_61/B 0.01fF
C31325 AND2X1_LOC_58/a_8_24# OR2X1_LOC_61/B 0.01fF
C1786 OR2X1_LOC_592/A OR2X1_LOC_592/a_8_216# 0.47fF
C37245 VDD OR2X1_LOC_592/A -0.00fF
C57809 OR2X1_LOC_592/A VSS 0.15fF
C21491 AND2X1_LOC_666/a_8_24# OR2X1_LOC_241/B 0.03fF
C47435 OR2X1_LOC_541/a_8_216# OR2X1_LOC_241/B 0.02fF
C52551 AND2X1_LOC_75/a_8_24# OR2X1_LOC_241/B 0.04fF
C53468 AND2X1_LOC_237/a_8_24# OR2X1_LOC_241/B 0.01fF
C53653 OR2X1_LOC_188/a_8_216# OR2X1_LOC_241/B -0.03fF
C11153 AND2X1_LOC_67/a_8_24# OR2X1_LOC_66/Y 0.11fF
C17060 AND2X1_LOC_131/a_8_24# OR2X1_LOC_66/Y 0.01fF
C27728 OR2X1_LOC_115/a_8_216# OR2X1_LOC_66/Y 0.01fF
C40783 OR2X1_LOC_216/A OR2X1_LOC_66/Y 0.75fF
C49591 OR2X1_LOC_116/a_8_216# OR2X1_LOC_66/Y 0.01fF
C16443 OR2X1_LOC_834/A AND2X1_LOC_305/a_8_24# 0.08fF
C18026 OR2X1_LOC_308/A OR2X1_LOC_834/A 0.04fF
C53048 VDD OR2X1_LOC_834/A 0.21fF
C57461 OR2X1_LOC_834/A VSS 0.40fF
C2473 OR2X1_LOC_334/B OR2X1_LOC_634/a_8_216# 0.08fF
C27376 OR2X1_LOC_334/B OR2X1_LOC_334/a_8_216# 0.07fF
C57454 OR2X1_LOC_334/B VSS -0.03fF
C37438 AND2X1_LOC_27/a_8_24# OR2X1_LOC_34/B 0.01fF
C11911 OR2X1_LOC_668/Y AND2X1_LOC_669/a_8_24# 0.23fF
C29185 VDD OR2X1_LOC_668/Y 0.16fF
C56748 OR2X1_LOC_668/Y VSS 0.07fF
C10390 AND2X1_LOC_437/a_8_24# OR2X1_LOC_180/B 0.01fF
C27860 AND2X1_LOC_176/a_8_24# OR2X1_LOC_180/B 0.09fF
C53381 AND2X1_LOC_177/a_8_24# OR2X1_LOC_180/B 0.01fF
C22058 OR2X1_LOC_319/a_8_216# OR2X1_LOC_538/A 0.01fF
C43946 OR2X1_LOC_538/A OR2X1_LOC_186/a_8_216# 0.01fF
C45367 AND2X1_LOC_173/a_8_24# OR2X1_LOC_538/A 0.01fF
C55214 OR2X1_LOC_325/a_8_216# OR2X1_LOC_538/A 0.01fF
C55596 OR2X1_LOC_538/A AND2X1_LOC_167/a_8_24# 0.01fF
C4342 AND2X1_LOC_394/a_36_24# OR2X1_LOC_84/A 0.01fF
C40396 AND2X1_LOC_393/a_8_24# OR2X1_LOC_84/A 0.20fF
C43875 AND2X1_LOC_394/a_8_24# OR2X1_LOC_84/A 0.03fF
C51644 AND2X1_LOC_393/a_36_24# OR2X1_LOC_84/A 0.01fF
C6823 AND2X1_LOC_385/a_8_24# OR2X1_LOC_389/B 0.02fF
C20291 OR2X1_LOC_389/B OR2X1_LOC_389/a_8_216# 0.01fF
C25302 OR2X1_LOC_389/B OR2X1_LOC_537/a_8_216# 0.47fF
C57847 OR2X1_LOC_389/B VSS 0.23fF
C6173 OR2X1_LOC_113/a_8_216# OR2X1_LOC_643/A 0.01fF
C22673 OR2X1_LOC_643/A AND2X1_LOC_122/a_8_24# 0.05fF
C27725 OR2X1_LOC_643/A AND2X1_LOC_106/a_8_24# 0.01fF
C230 OR2X1_LOC_379/Y OR2X1_LOC_855/a_8_216# 0.01fF
C1588 OR2X1_LOC_379/Y VDD 0.14fF
C21684 OR2X1_LOC_379/Y AND2X1_LOC_586/a_8_24# 0.01fF
C47485 OR2X1_LOC_379/Y OR2X1_LOC_769/a_8_216# 0.01fF
C52076 OR2X1_LOC_379/Y OR2X1_LOC_198/A 0.02fF
C58057 OR2X1_LOC_379/Y VSS 0.08fF
C57921 OR2X1_LOC_308/A VSS 0.18fF
C14097 OR2X1_LOC_198/a_8_216# OR2X1_LOC_198/A 0.13fF
C45117 OR2X1_LOC_855/a_8_216# OR2X1_LOC_198/A 0.14fF
C46069 AND2X1_LOC_52/a_8_24# OR2X1_LOC_198/A 0.23fF
C46497 VDD OR2X1_LOC_198/A 0.48fF
C55451 OR2X1_LOC_828/a_8_216# OR2X1_LOC_198/A 0.12fF
C56244 OR2X1_LOC_198/A VSS 0.46fF
C11633 AND2X1_LOC_635/a_8_24# AND2X1_LOC_639/A 0.05fF
C26546 OR2X1_LOC_451/a_8_216# OR2X1_LOC_452/A -0.00fF
C27522 VDD OR2X1_LOC_593/A -0.00fF
C34350 OR2X1_LOC_799/A OR2X1_LOC_593/A 0.11fF
C46425 OR2X1_LOC_593/A OR2X1_LOC_593/a_8_216# 0.39fF
C48230 OR2X1_LOC_592/a_8_216# OR2X1_LOC_593/A -0.00fF
C56829 OR2X1_LOC_593/A VSS 0.18fF
C2900 VDD OR2X1_LOC_799/A 0.15fF
C21721 OR2X1_LOC_799/A OR2X1_LOC_593/a_8_216# 0.01fF
C23450 OR2X1_LOC_799/A OR2X1_LOC_592/a_8_216# 0.01fF
C29234 OR2X1_LOC_318/Y OR2X1_LOC_799/A 0.03fF
C30206 OR2X1_LOC_799/A AND2X1_LOC_165/a_8_24# 0.23fF
C30640 OR2X1_LOC_799/A OR2X1_LOC_436/Y 0.03fF
C30975 OR2X1_LOC_799/A OR2X1_LOC_799/a_8_216# 0.07fF
C38607 AND2X1_LOC_589/a_8_24# OR2X1_LOC_799/A 0.09fF
C57708 OR2X1_LOC_799/A VSS 0.22fF
C9325 OR2X1_LOC_319/B OR2X1_LOC_319/a_8_216# 0.02fF
C20348 OR2X1_LOC_319/B OR2X1_LOC_319/a_36_216# 0.02fF
C22429 OR2X1_LOC_319/B VDD 0.82fF
C42767 OR2X1_LOC_319/B AND2X1_LOC_167/a_8_24# 0.06fF
C57952 OR2X1_LOC_319/B VSS 0.08fF
C28889 OR2X1_LOC_436/B OR2X1_LOC_436/a_8_216# 0.02fF
C30211 OR2X1_LOC_436/B OR2X1_LOC_436/Y 0.76fF
C42783 OR2X1_LOC_434/a_8_216# OR2X1_LOC_436/B -0.00fF
C57265 OR2X1_LOC_436/B VSS 0.08fF
C13403 VDD AND2X1_LOC_287/B 0.29fF
C43167 OR2X1_LOC_669/a_8_216# AND2X1_LOC_287/B 0.04fF
C56771 AND2X1_LOC_287/B VSS 0.19fF
C17226 AND2X1_LOC_114/Y AND2X1_LOC_116/a_8_24# 0.19fF
C26362 VDD AND2X1_LOC_114/Y 0.21fF
C57170 AND2X1_LOC_114/Y VSS 0.06fF
C20188 AND2X1_LOC_483/Y AND2X1_LOC_483/a_8_24# 0.02fF
C22287 AND2X1_LOC_483/Y AND2X1_LOC_621/Y 0.05fF
C31500 AND2X1_LOC_456/B AND2X1_LOC_483/Y 0.14fF
C28640 AND2X1_LOC_318/Y AND2X1_LOC_319/a_8_24# 0.06fF
C34833 VDD AND2X1_LOC_318/Y 0.51fF
C43384 AND2X1_LOC_335/a_8_24# AND2X1_LOC_318/Y 0.17fF
C57192 AND2X1_LOC_318/Y VSS 0.35fF
C1625 OR2X1_LOC_114/Y VDD 0.12fF
C8955 OR2X1_LOC_114/Y OR2X1_LOC_631/a_8_216# 0.13fF
C12812 OR2X1_LOC_114/Y OR2X1_LOC_116/a_8_216# 0.07fF
C13229 OR2X1_LOC_116/A OR2X1_LOC_114/Y 0.06fF
C19171 OR2X1_LOC_114/Y OR2X1_LOC_631/B 0.10fF
C52668 OR2X1_LOC_114/Y OR2X1_LOC_361/a_8_216# 0.01fF
C53065 OR2X1_LOC_114/Y OR2X1_LOC_267/Y 0.02fF
C57851 OR2X1_LOC_114/Y VSS 0.09fF
C19546 VDD OR2X1_LOC_456/A -0.00fF
C53005 OR2X1_LOC_456/A OR2X1_LOC_344/a_8_216# 0.46fF
C57207 OR2X1_LOC_456/A VSS 0.34fF
C269 OR2X1_LOC_631/B AND2X1_LOC_627/a_8_24# 0.03fF
C1362 OR2X1_LOC_631/B OR2X1_LOC_629/a_8_216# 0.01fF
C4798 OR2X1_LOC_631/B OR2X1_LOC_247/a_8_216# 0.06fF
C6745 OR2X1_LOC_629/Y OR2X1_LOC_631/B 0.01fF
C6847 OR2X1_LOC_631/B OR2X1_LOC_629/a_36_216# 0.01fF
C11609 OR2X1_LOC_631/B AND2X1_LOC_665/a_8_24# 0.04fF
C14498 OR2X1_LOC_483/a_8_216# OR2X1_LOC_631/B 0.03fF
C15846 OR2X1_LOC_631/B OR2X1_LOC_247/a_36_216# 0.01fF
C20855 OR2X1_LOC_631/a_8_216# OR2X1_LOC_631/B 0.02fF
C23430 OR2X1_LOC_630/a_8_216# OR2X1_LOC_631/B 0.01fF
C23442 OR2X1_LOC_664/a_8_216# OR2X1_LOC_631/B 0.03fF
C25533 OR2X1_LOC_483/a_36_216# OR2X1_LOC_631/B 0.01fF
C26319 OR2X1_LOC_631/a_36_216# OR2X1_LOC_631/B 0.01fF
C34339 OR2X1_LOC_664/a_36_216# OR2X1_LOC_631/B 0.01fF
C38634 AND2X1_LOC_72/a_8_24# OR2X1_LOC_631/B 0.04fF
C5624 AND2X1_LOC_172/a_8_24# OR2X1_LOC_539/B 0.17fF
C7860 OR2X1_LOC_539/a_8_216# OR2X1_LOC_539/B 0.40fF
C39170 VDD OR2X1_LOC_539/B 0.31fF
C43639 AND2X1_LOC_431/a_8_24# OR2X1_LOC_539/B 0.18fF
C50876 OR2X1_LOC_539/A OR2X1_LOC_539/B 0.12fF
C56259 OR2X1_LOC_539/B VSS 0.66fF
C58128 OR2X1_LOC_539/A VSS 0.18fF
C549 AND2X1_LOC_537/Y AND2X1_LOC_538/Y 0.11fF
C6046 AND2X1_LOC_537/Y AND2X1_LOC_539/a_8_24# 0.09fF
C7781 AND2X1_LOC_537/Y AND2X1_LOC_307/a_8_24# 0.06fF
C18866 AND2X1_LOC_537/Y AND2X1_LOC_307/a_36_24# 0.01fF
C48979 VDD AND2X1_LOC_537/Y 0.63fF
C57489 AND2X1_LOC_537/Y VSS -0.35fF
C3848 VDD AND2X1_LOC_538/Y 0.23fF
C17157 AND2X1_LOC_538/Y AND2X1_LOC_539/a_8_24# 0.19fF
C22767 AND2X1_LOC_538/a_8_24# AND2X1_LOC_538/Y 0.01fF
C39461 AND2X1_LOC_538/Y AND2X1_LOC_434/Y -0.01fF
C57488 AND2X1_LOC_538/Y VSS 0.07fF
C28937 OR2X1_LOC_802/a_8_216# OR2X1_LOC_436/Y 0.01fF
C37704 OR2X1_LOC_112/a_8_216# OR2X1_LOC_436/Y 0.01fF
C43013 OR2X1_LOC_436/Y OR2X1_LOC_809/a_8_216# 0.01fF
C46044 OR2X1_LOC_436/Y OR2X1_LOC_798/a_8_216# 0.16fF
C50372 OR2X1_LOC_318/Y OR2X1_LOC_436/Y 0.03fF
C52037 OR2X1_LOC_436/Y OR2X1_LOC_799/a_8_216# 0.01fF
C15213 AND2X1_LOC_99/A AND2X1_LOC_99/Y 0.37fF
C27240 AND2X1_LOC_99/Y AND2X1_LOC_101/a_8_24# 0.07fF
C35939 AND2X1_LOC_99/a_8_24# AND2X1_LOC_99/Y 0.02fF
C57406 AND2X1_LOC_99/Y VSS 0.15fF
C57715 OR2X1_LOC_629/Y VSS 0.09fF
C50842 AND2X1_LOC_838/B AND2X1_LOC_838/a_8_24# 0.19fF
C55381 VDD AND2X1_LOC_838/B 0.23fF
C56882 AND2X1_LOC_838/B VSS -0.15fF
C4152 AND2X1_LOC_99/A AND2X1_LOC_99/a_8_24# 0.05fF
C20785 AND2X1_LOC_99/A AND2X1_LOC_99/a_36_24# 0.01fF
C41465 OR2X1_LOC_122/a_8_216# AND2X1_LOC_99/A 0.01fF
C42445 AND2X1_LOC_99/A OR2X1_LOC_67/a_8_216# 0.01fF
C43606 OR2X1_LOC_106/a_8_216# AND2X1_LOC_99/A 0.01fF
C44421 OR2X1_LOC_117/a_8_216# AND2X1_LOC_99/A 0.03fF
C45788 VDD AND2X1_LOC_99/A 0.35fF
C50091 OR2X1_LOC_117/a_36_216# AND2X1_LOC_99/A 0.01fF
C57525 AND2X1_LOC_99/A VSS 0.24fF
C11949 OR2X1_LOC_837/Y AND2X1_LOC_826/a_8_24# 0.01fF
C32922 VDD OR2X1_LOC_837/Y 0.22fF
C35617 OR2X1_LOC_837/Y OR2X1_LOC_20/a_8_216# 0.01fF
C41130 OR2X1_LOC_837/Y OR2X1_LOC_20/a_36_216# 0.02fF
C57417 OR2X1_LOC_837/Y VSS -0.22fF
C50897 VDD OR2X1_LOC_162/Y 0.16fF
C55051 OR2X1_LOC_162/Y AND2X1_LOC_163/a_8_24# 0.23fF
C57638 OR2X1_LOC_162/Y VSS 0.07fF
C2594 OR2X1_LOC_145/a_8_216# AND2X1_LOC_621/Y 0.14fF
C7604 AND2X1_LOC_631/a_8_24# AND2X1_LOC_621/Y 0.02fF
C8105 OR2X1_LOC_627/a_8_216# AND2X1_LOC_621/Y 0.06fF
C12656 OR2X1_LOC_496/a_8_216# AND2X1_LOC_621/Y 0.04fF
C14367 VDD AND2X1_LOC_621/Y 0.98fF
C15244 AND2X1_LOC_621/Y OR2X1_LOC_531/a_8_216# 0.04fF
C30126 AND2X1_LOC_154/a_8_24# AND2X1_LOC_621/Y 0.26fF
C38094 AND2X1_LOC_621/Y AND2X1_LOC_622/a_8_24# 0.03fF
C49406 AND2X1_LOC_621/Y AND2X1_LOC_622/a_36_24# 0.01fF
C49929 AND2X1_LOC_621/Y AND2X1_LOC_678/a_8_24# 0.10fF
C51535 AND2X1_LOC_621/Y OR2X1_LOC_239/a_8_216# 0.04fF
C56914 AND2X1_LOC_621/Y VSS -1.20fF
C3661 VDD AND2X1_LOC_285/Y 0.19fF
C16812 AND2X1_LOC_285/Y AND2X1_LOC_286/a_8_24# 0.11fF
C31261 AND2X1_LOC_456/B AND2X1_LOC_285/Y 0.35fF
C44559 OR2X1_LOC_754/a_8_216# AND2X1_LOC_285/Y 0.14fF
C56665 AND2X1_LOC_285/Y VSS -0.83fF
C4311 AND2X1_LOC_434/Y OR2X1_LOC_311/a_8_216# 0.03fF
C8086 AND2X1_LOC_855/a_8_24# AND2X1_LOC_434/Y 0.02fF
C10008 AND2X1_LOC_809/a_8_24# AND2X1_LOC_434/Y 0.01fF
C12301 AND2X1_LOC_355/a_8_24# AND2X1_LOC_434/Y 0.01fF
C17611 OR2X1_LOC_13/a_8_216# AND2X1_LOC_434/Y 0.03fF
C31725 OR2X1_LOC_829/a_8_216# AND2X1_LOC_434/Y 0.01fF
C35860 AND2X1_LOC_539/a_36_24# AND2X1_LOC_434/Y 0.01fF
C36927 OR2X1_LOC_41/a_8_216# AND2X1_LOC_434/Y 0.04fF
C41364 AND2X1_LOC_538/a_36_24# AND2X1_LOC_434/Y 0.01fF
C42577 AND2X1_LOC_434/Y OR2X1_LOC_331/Y 0.28fF
C45069 AND2X1_LOC_539/a_8_24# AND2X1_LOC_434/Y 0.02fF
C50722 AND2X1_LOC_538/a_8_24# AND2X1_LOC_434/Y 0.03fF
C56573 AND2X1_LOC_434/Y VSS -1.84fF
C15624 AND2X1_LOC_456/B AND2X1_LOC_287/a_8_24# 0.01fF
C16349 OR2X1_LOC_482/a_8_216# AND2X1_LOC_456/B 0.02fF
C23689 VDD AND2X1_LOC_456/B 0.58fF
C36695 AND2X1_LOC_456/B AND2X1_LOC_286/a_8_24# 0.18fF
C41049 AND2X1_LOC_456/B AND2X1_LOC_843/a_8_24# 0.01fF
C41947 AND2X1_LOC_456/B AND2X1_LOC_668/a_8_24# 0.01fF
C44435 AND2X1_LOC_456/B OR2X1_LOC_666/a_8_216# 0.01fF
C53607 AND2X1_LOC_456/B OR2X1_LOC_669/a_8_216# 0.01fF
C57667 AND2X1_LOC_456/B VSS 0.45fF
C20767 VDD OR2X1_LOC_464/B -0.00fF
C28890 OR2X1_LOC_457/a_8_216# OR2X1_LOC_464/B -0.00fF
C44117 OR2X1_LOC_464/a_8_216# OR2X1_LOC_464/B 0.39fF
C57212 OR2X1_LOC_464/B VSS 0.17fF
C9340 OR2X1_LOC_318/Y OR2X1_LOC_319/a_8_216# 0.02fF
C22450 OR2X1_LOC_318/Y VDD 0.15fF
C42873 OR2X1_LOC_318/Y OR2X1_LOC_592/a_8_216# 0.03fF
C48577 OR2X1_LOC_318/Y OR2X1_LOC_592/a_36_216# 0.02fF
C50657 OR2X1_LOC_318/Y OR2X1_LOC_799/a_8_216# 0.04fF
C57864 OR2X1_LOC_318/Y VSS 0.39fF
C23045 OR2X1_LOC_287/A OR2X1_LOC_287/a_8_216# 0.01fF
C25334 VDD OR2X1_LOC_287/A 0.17fF
C57371 OR2X1_LOC_287/A VSS 0.02fF
C3706 AND2X1_LOC_464/a_8_24# AND2X1_LOC_464/A -0.00fF
C56630 AND2X1_LOC_464/A VSS 0.28fF
C12111 AND2X1_LOC_592/Y VDD 0.08fF
C33730 AND2X1_LOC_592/Y AND2X1_LOC_593/a_8_24# 0.01fF
C34632 AND2X1_LOC_592/Y OR2X1_LOC_424/a_8_216# 0.01fF
C55175 AND2X1_LOC_592/Y AND2X1_LOC_593/Y 0.01fF
C58114 AND2X1_LOC_592/Y VSS 0.14fF
C19431 OR2X1_LOC_163/A OR2X1_LOC_163/a_8_216# 0.47fF
C56290 OR2X1_LOC_163/A VSS 0.15fF
C46994 OR2X1_LOC_285/Y OR2X1_LOC_286/a_8_216# 0.39fF
C57258 OR2X1_LOC_285/Y VSS 0.18fF
C527 AND2X1_LOC_319/A AND2X1_LOC_319/a_8_24# 0.03fF
C6667 VDD AND2X1_LOC_319/A 0.29fF
C37124 AND2X1_LOC_319/A OR2X1_LOC_312/a_8_216# 0.18fF
C37339 AND2X1_LOC_319/A OR2X1_LOC_418/a_8_216# 0.47fF
C40969 AND2X1_LOC_319/A AND2X1_LOC_809/a_8_24# 0.13fF
C57298 AND2X1_LOC_319/A VSS 0.54fF
C21185 VDD AND2X1_LOC_113/Y 0.33fF
C51925 AND2X1_LOC_113/Y AND2X1_LOC_114/a_8_24# 0.11fF
C57282 AND2X1_LOC_113/Y VSS 0.15fF
C27089 AND2X1_LOC_593/Y AND2X1_LOC_436/Y 0.02fF
C28746 OR2X1_LOC_600/a_8_216# AND2X1_LOC_593/Y 0.06fF
C38898 VDD AND2X1_LOC_593/Y 0.08fF
C57066 AND2X1_LOC_593/Y VSS 0.32fF
C11055 VDD AND2X1_LOC_629/Y 0.01fF
C31559 AND2X1_LOC_629/Y AND2X1_LOC_630/a_8_24# 0.03fF
C42625 AND2X1_LOC_629/Y AND2X1_LOC_630/a_36_24# 0.01fF
C57070 AND2X1_LOC_629/Y VSS 0.23fF
C3132 AND2X1_LOC_436/a_8_24# OR2X1_LOC_331/Y 0.01fF
C6882 VDD OR2X1_LOC_331/Y 0.12fF
C15001 AND2X1_LOC_330/a_8_24# OR2X1_LOC_331/Y 0.23fF
C19685 OR2X1_LOC_166/a_8_216# OR2X1_LOC_331/Y 0.01fF
C22523 OR2X1_LOC_533/a_8_216# OR2X1_LOC_331/Y 0.05fF
C29390 AND2X1_LOC_535/a_8_24# OR2X1_LOC_331/Y 0.04fF
C43497 AND2X1_LOC_355/a_8_24# OR2X1_LOC_331/Y 0.05fF
C51833 OR2X1_LOC_331/a_8_216# OR2X1_LOC_331/Y 0.03fF
C56387 OR2X1_LOC_331/Y VSS 0.34fF
C9011 OR2X1_LOC_113/Y AND2X1_LOC_106/a_8_24# 0.23fF
C39694 OR2X1_LOC_113/Y VDD 0.12fF
C57937 OR2X1_LOC_113/Y VSS 0.19fF
C7543 OR2X1_LOC_116/A VDD -0.00fF
C18744 OR2X1_LOC_116/A OR2X1_LOC_116/a_8_216# 0.39fF
C53179 OR2X1_LOC_115/a_8_216# OR2X1_LOC_116/A -0.00fF
C57902 OR2X1_LOC_116/A VSS 0.18fF
C45889 VDD OR2X1_LOC_99/B 0.18fF
C56912 OR2X1_LOC_99/B VSS 0.19fF
C36353 VDD OR2X1_LOC_848/B 0.05fF
C45852 OR2X1_LOC_848/B OR2X1_LOC_391/a_8_216# 0.04fF
C57618 OR2X1_LOC_848/B VSS 0.05fF
C25440 OR2X1_LOC_622/A OR2X1_LOC_622/a_8_216# 0.02fF
C57585 OR2X1_LOC_622/A VSS 0.10fF
C7111 AND2X1_LOC_361/a_36_24# AND2X1_LOC_361/A 0.02fF
C7242 AND2X1_LOC_267/a_8_24# AND2X1_LOC_361/A -0.03fF
C11409 OR2X1_LOC_132/a_8_216# AND2X1_LOC_361/A 0.01fF
C32778 OR2X1_LOC_72/a_8_216# AND2X1_LOC_361/A 0.47fF
C33350 AND2X1_LOC_541/a_8_24# AND2X1_LOC_361/A -0.03fF
C36348 AND2X1_LOC_130/a_8_24# AND2X1_LOC_361/A 0.02fF
C39266 OR2X1_LOC_134/a_8_216# AND2X1_LOC_361/A 0.04fF
C46707 AND2X1_LOC_361/a_8_24# AND2X1_LOC_361/A 0.07fF
C53183 OR2X1_LOC_265/a_8_216# AND2X1_LOC_361/A 0.04fF
C5184 AND2X1_LOC_848/A AND2X1_LOC_848/a_8_24# 0.02fF
C23179 OR2X1_LOC_258/a_8_216# AND2X1_LOC_848/A 0.03fF
C30212 AND2X1_LOC_709/a_8_24# AND2X1_LOC_848/A -0.01fF
C31970 OR2X1_LOC_295/a_8_216# AND2X1_LOC_848/A 0.03fF
C41212 AND2X1_LOC_709/a_36_24# AND2X1_LOC_848/A -0.02fF
C56981 AND2X1_LOC_848/A VSS -0.77fF
C11208 OR2X1_LOC_355/A OR2X1_LOC_355/a_8_216# 0.47fF
C56292 OR2X1_LOC_355/A VSS 0.13fF
C8849 OR2X1_LOC_99/Y AND2X1_LOC_607/a_8_24# 0.01fF
C20002 OR2X1_LOC_101/a_8_216# OR2X1_LOC_99/Y 0.03fF
C56816 OR2X1_LOC_99/Y VSS 0.22fF
C11454 OR2X1_LOC_687/Y AND2X1_LOC_615/a_8_24# 0.06fF
C31696 OR2X1_LOC_687/Y OR2X1_LOC_729/a_8_216# 0.05fF
C44975 OR2X1_LOC_687/Y OR2X1_LOC_678/a_8_216# 0.03fF
C50625 OR2X1_LOC_687/Y OR2X1_LOC_678/a_36_216# 0.02fF
C21576 OR2X1_LOC_594/a_8_216# AND2X1_LOC_436/Y -0.00fF
C29897 AND2X1_LOC_799/a_8_24# AND2X1_LOC_436/Y 0.01fF
C38750 AND2X1_LOC_798/a_8_24# AND2X1_LOC_436/Y 0.03fF
C50019 AND2X1_LOC_798/a_36_24# AND2X1_LOC_436/Y 0.01fF
C53050 OR2X1_LOC_166/a_8_216# AND2X1_LOC_436/Y 0.47fF
C8174 OR2X1_LOC_432/a_8_216# AND2X1_LOC_687/Y 0.18fF
C29254 AND2X1_LOC_729/a_8_24# AND2X1_LOC_687/Y 0.09fF
C15462 AND2X1_LOC_116/B AND2X1_LOC_116/a_8_24# 0.01fF
C24662 VDD AND2X1_LOC_116/B 0.04fF
C57224 AND2X1_LOC_116/B VSS -0.15fF
C16404 AND2X1_LOC_798/a_8_24# AND2X1_LOC_798/Y 0.01fF
C56978 AND2X1_LOC_798/Y VSS 0.11fF
C58005 AND2X1_LOC_802/B VSS 0.20fF
C57617 OR2X1_LOC_798/Y VSS 0.28fF
C7108 AND2X1_LOC_539/Y AND2X1_LOC_855/a_8_24# 0.01fF
C11328 AND2X1_LOC_539/Y AND2X1_LOC_355/a_8_24# 0.18fF
C20569 AND2X1_LOC_539/Y AND2X1_LOC_799/a_8_24# 0.01fF
C30712 AND2X1_LOC_539/Y VDD 0.22fF
C58006 AND2X1_LOC_539/Y VSS -0.29fF
C18605 VDD OR2X1_LOC_539/Y 0.27fF
C23804 OR2X1_LOC_802/a_8_216# OR2X1_LOC_539/Y 0.05fF
C32503 OR2X1_LOC_112/a_8_216# OR2X1_LOC_539/Y 0.03fF
C40690 OR2X1_LOC_798/a_8_216# OR2X1_LOC_539/Y 0.01fF
C42196 OR2X1_LOC_539/Y OR2X1_LOC_332/a_8_216# 0.01fF
C12242 OR2X1_LOC_216/A OR2X1_LOC_473/a_8_216# 0.04fF
C47478 OR2X1_LOC_216/A AND2X1_LOC_239/a_8_24# 0.03fF
C54720 VDD OR2X1_LOC_216/A 0.19fF
C45269 AND2X1_LOC_319/a_8_24# AND2X1_LOC_798/A 0.02fF
C51559 VDD AND2X1_LOC_798/A 0.21fF
C54823 VDD AND2X1_LOC_116/Y 0.21fF
C56961 AND2X1_LOC_116/Y VSS 0.25fF
C56336 OR2X1_LOC_319/Y VSS 0.28fF
C56609 OR2X1_LOC_802/A VSS 0.18fF
C14233 AND2X1_LOC_802/Y AND2X1_LOC_809/a_36_24# 0.01fF
C24859 VDD AND2X1_LOC_802/Y 0.01fF
C56585 AND2X1_LOC_802/Y VSS 0.24fF

.ends

* wrdata outputs.out V("OR2X1_LOC_452/A") V("AND2X1_LOC_639/A") V("OR2X1_LOC_460/Y") V("OR2X1_LOC_198/A") V("OR2X1_LOC_308/A") V("OR2X1_LOC_379/Y") V("OR2X1_LOC_643/A") V("OR2X1_LOC_84/A") V("OR2X1_LOC_538/A") V("OR2X1_LOC_180/B") V("OR2X1_LOC_668/Y") V("OR2X1_LOC_34/B") V("OR2X1_LOC_334/B") V("OR2X1_LOC_834/A") V("OR2X1_LOC_241/B") V("OR2X1_LOC_523/A") V("OR2X1_LOC_33/A") V("OR2X1_LOC_61/B") V("OR2X1_LOC_844/B") V("OR2X1_LOC_623/B") V("OR2X1_LOC_770/A") V("OR2X1_LOC_324/A") V("OR2X1_LOC_509/A") V("OR2X1_LOC_703/A") V("OR2X1_LOC_147/B") V("OR2X1_LOC_201/A") V("OR2X1_LOC_520/B") V("OR2X1_LOC_703/B") V("OR2X1_LOC_835/A") V("OR2X1_LOC_709/B") V("OR2X1_LOC_720/B") V("OR2X1_LOC_343/B") V("OR2X1_LOC_855/A") V("OR2X1_LOC_449/B") V("OR2X1_LOC_593/B") V("OR2X1_LOC_773/B") V("OR2X1_LOC_402/B") V("OR2X1_LOC_307/A") V("OR2X1_LOC_128/A") V("OR2X1_LOC_194/B") V("OR2X1_LOC_555/A") V("OR2X1_LOC_719/B") V("AND2X1_LOC_7/Y") V("OR2X1_LOC_789/A") V("OR2X1_LOC_769/A") V("OR2X1_LOC_400/B") V("OR2X1_LOC_781/B") V("OR2X1_LOC_549/B") V("OR2X1_LOC_391/A") V("OR2X1_LOC_333/B") V("OR2X1_LOC_190/B") V("AND2X1_LOC_41/Y") V("OR2X1_LOC_610/Y") V("OR2X1_LOC_191/B") V("OR2X1_LOC_169/B") V("OR2X1_LOC_673/B") V("OR2X1_LOC_346/B") V("OR2X1_LOC_545/B") V("OR2X1_LOC_444/B") V("OR2X1_LOC_620/A") V("OR2X1_LOC_786/A") V("OR2X1_LOC_641/A") V("OR2X1_LOC_758/Y") V("OR2X1_LOC_637/A") V("OR2X1_LOC_174/A") V("AND2X1_LOC_72/Y") V("OR2X1_LOC_175/B") V("OR2X1_LOC_439/B") V("OR2X1_LOC_835/B") V("OR2X1_LOC_123/B") V("OR2X1_LOC_633/B") V("OR2X1_LOC_675/A") V("OR2X1_LOC_501/B") V("OR2X1_LOC_605/A") V("OR2X1_LOC_544/A") V("OR2X1_LOC_450/A") V("OR2X1_LOC_103/Y") V("OR2X1_LOC_106/Y") V("OR2X1_LOC_695/Y") V("OR2X1_LOC_280/Y") V("OR2X1_LOC_601/Y") V("OR2X1_LOC_612/B") V("OR2X1_LOC_248/Y") V("OR2X1_LOC_394/Y") V("OR2X1_LOC_747/Y") V("OR2X1_LOC_524/Y") V("OR2X1_LOC_152/Y") V("OR2X1_LOC_528/Y") V("OR2X1_LOC_122/Y") V("OR2X1_LOC_485/Y") V("OR2X1_LOC_297/Y") V("OR2X1_LOC_424/Y") V("OR2X1_LOC_45/Y") V("OR2X1_LOC_744/Y") V("OR2X1_LOC_701/Y") V("OR2X1_LOC_757/Y") V("OR2X1_LOC_399/Y") V("OR2X1_LOC_517/Y") V("OR2X1_LOC_315/Y") V("OR2X1_LOC_491/Y") V("OR2X1_LOC_109/Y") V("OR2X1_LOC_600/Y") V("OR2X1_LOC_230/Y") V("OR2X1_LOC_298/Y") V("OR2X1_LOC_224/Y") V("OR2X1_LOC_428/Y") V("OR2X1_LOC_74/Y") V("OR2X1_LOC_32/Y") V("OR2X1_LOC_583/Y") V("OR2X1_LOC_526/Y") V("OR2X1_LOC_505/Y") V("OR2X1_LOC_666/Y") V("OR2X1_LOC_496/Y") V("OR2X1_LOC_432/Y") V("OR2X1_LOC_607/Y") V("OR2X1_LOC_257/Y") V("OR2X1_LOC_20/Y") V("OR2X1_LOC_79/Y") V("OR2X1_LOC_521/Y") V("OR2X1_LOC_135/Y") V("OR2X1_LOC_492/Y") V("OR2X1_LOC_482/Y") V("OR2X1_LOC_108/Y") V("OR2X1_LOC_295/Y") V("OR2X1_LOC_81/Y") V("OR2X1_LOC_60/Y") V("OR2X1_LOC_437/Y") V("OR2X1_LOC_609/Y") V("OR2X1_LOC_75/Y") V("OR2X1_LOC_700/Y") V("OR2X1_LOC_755/Y") V("OR2X1_LOC_395/Y") V("OR2X1_LOC_494/Y") V("OR2X1_LOC_380/A") V("OR2X1_LOC_603/Y") V("OR2X1_LOC_261/A") V("OR2X1_LOC_679/A") V("OR2X1_LOC_229/Y") V("OR2X1_LOC_13/Y") V("OR2X1_LOC_765/Y") V("OR2X1_LOC_131/Y") V("AND2X1_LOC_793/B") V("OR2X1_LOC_712/B") V("OR2X1_LOC_791/B") V("OR2X1_LOC_710/B") V("OR2X1_LOC_401/B") V("OR2X1_LOC_84/B") V("OR2X1_LOC_61/A") V("OR2X1_LOC_76/A") V("OR2X1_LOC_702/A") V("OR2X1_LOC_493/A") V("OR2X1_LOC_833/B") V("OR2X1_LOC_114/B") V("OR2X1_LOC_346/A") V("OR2X1_LOC_440/B") V("OR2X1_LOC_646/A") V("OR2X1_LOC_231/B") V("OR2X1_LOC_770/B") V("OR2X1_LOC_140/A") V("OR2X1_LOC_260/Y") V("OR2X1_LOC_678/Y") V("OR2X1_LOC_193/A") V("OR2X1_LOC_558/A") V("OR2X1_LOC_605/B") V("OR2X1_LOC_653/B") V("OR2X1_LOC_788/B") V("OR2X1_LOC_190/A") V("OR2X1_LOC_98/A") V("OR2X1_LOC_137/B") V("OR2X1_LOC_192/B") V("OR2X1_LOC_768/A") V("OR2X1_LOC_128/B") V("OR2X1_LOC_447/A") V("OR2X1_LOC_489/B") V("OR2X1_LOC_475/B") V("OR2X1_LOC_644/B") V("OR2X1_LOC_448/Y") V("OR2X1_LOC_356/A") V("OR2X1_LOC_176/Y") V("OR2X1_LOC_290/Y") V("OR2X1_LOC_677/Y") V("OR2X1_LOC_83/Y") V("OR2X1_LOC_237/Y") V("OR2X1_LOC_669/A") V("OR2X1_LOC_595/Y") V("OR2X1_LOC_27/Y") V("OR2X1_LOC_311/Y") V("OR2X1_LOC_146/Y") V("OR2X1_LOC_179/Y") V("OR2X1_LOC_484/Y") V("OR2X1_LOC_495/Y") V("OR2X1_LOC_754/Y") V("OR2X1_LOC_69/Y") V("OR2X1_LOC_39/Y") V("OR2X1_LOC_396/Y") V("OR2X1_LOC_320/Y") V("OR2X1_LOC_497/Y") V("OR2X1_LOC_615/Y") V("OR2X1_LOC_24/Y") V("OR2X1_LOC_58/Y") V("OR2X1_LOC_522/Y") V("AND2X1_LOC_549/Y") V("OR2X1_LOC_711/B") V("OR2X1_LOC_713/A") V("AND2X1_LOC_335/Y") V("AND2X1_LOC_778/Y") V("AND2X1_LOC_208/B") V("OR2X1_LOC_72/Y") V("OR2X1_LOC_184/Y") V("OR2X1_LOC_152/A") V("OR2X1_LOC_292/Y") V("OR2X1_LOC_173/Y") V("OR2X1_LOC_235/Y") V("AND2X1_LOC_784/A") V("AND2X1_LOC_633/Y") V("AND2X1_LOC_541/Y") V("AND2X1_LOC_634/Y") V("OR2X1_LOC_813/Y") V("OR2X1_LOC_624/B") V("AND2X1_LOC_721/A") V("AND2X1_LOC_69/Y") V("OR2X1_LOC_208/A") V("OR2X1_LOC_335/Y") V("OR2X1_LOC_778/Y") V("OR2X1_LOC_117/Y") V("OR2X1_LOC_262/Y") V("OR2X1_LOC_65/Y") V("OR2X1_LOC_471/B") V("AND2X1_LOC_303/A") V("AND2X1_LOC_831/Y") V("AND2X1_LOC_303/B") V("AND2X1_LOC_787/A") V("AND2X1_LOC_543/Y") V("OR2X1_LOC_841/A") V("OR2X1_LOC_841/B") V("OR2X1_LOC_828/Y") V("OR2X1_LOC_783/A") V("OR2X1_LOC_156/Y") V("OR2X1_LOC_708/Y") V("OR2X1_LOC_308/Y") V("OR2X1_LOC_149/B") V("OR2X1_LOC_168/Y") V("OR2X1_LOC_776/Y") V("OR2X1_LOC_325/Y") V("OR2X1_LOC_463/B") V("OR2X1_LOC_651/B") V("OR2X1_LOC_416/Y") V("AND2X1_LOC_637/Y") V("OR2X1_LOC_481/Y") V("AND2X1_LOC_631/Y") V("OR2X1_LOC_196/Y") V("OR2X1_LOC_520/Y") V("OR2X1_LOC_840/A") V("OR2X1_LOC_779/Y") V("AND2X1_LOC_632/A") V("AND2X1_LOC_448/Y") V("OR2X1_LOC_156/B") V("OR2X1_LOC_636/A") V("OR2X1_LOC_620/B") V("OR2X1_LOC_247/Y") V("OR2X1_LOC_231/A") V("OR2X1_LOC_130/Y") V("AND2X1_LOC_348/A") V("OR2X1_LOC_105/Y") V("OR2X1_LOC_181/A") V("OR2X1_LOC_602/B") V("OR2X1_LOC_345/A") V("OR2X1_LOC_756/Y") V("OR2X1_LOC_401/A") V("OR2X1_LOC_507/A") V("OR2X1_LOC_196/B") V("OR2X1_LOC_707/A") V("OR2X1_LOC_249/Y") V("OR2X1_LOC_776/A") V("OR2X1_LOC_793/B") V("AND2X1_LOC_557/Y") V("AND2X1_LOC_535/Y") V("AND2X1_LOC_199/A") V("AND2X1_LOC_508/A") V("AND2X1_LOC_447/Y") V("AND2X1_LOC_838/Y") V("AND2X1_LOC_139/B") V("OR2X1_LOC_178/Y") V("OR2X1_LOC_613/Y") V("OR2X1_LOC_67/Y") V("OR2X1_LOC_312/Y") V("OR2X1_LOC_647/B") V("OR2X1_LOC_132/Y") V("OR2X1_LOC_305/Y") V("OR2X1_LOC_494/A") V("OR2X1_LOC_91/Y") V("OR2X1_LOC_766/Y") V("OR2X1_LOC_670/Y") V("OR2X1_LOC_533/A") V("OR2X1_LOC_822/Y") V("OR2X1_LOC_420/Y") V("OR2X1_LOC_239/Y") V("OR2X1_LOC_172/Y") V("OR2X1_LOC_591/A") V("OR2X1_LOC_349/B") V("AND2X1_LOC_843/Y") V("AND2X1_LOC_287/Y") V("OR2X1_LOC_608/Y") V("OR2X1_LOC_602/A") V("OR2X1_LOC_78/Y") V("OR2X1_LOC_240/B") V("OR2X1_LOC_446/A") V("OR2X1_LOC_546/A") V("OR2X1_LOC_720/A") V("OR2X1_LOC_546/B") V("OR2X1_LOC_507/B") V("OR2X1_LOC_486/B") V("OR2X1_LOC_859/B") V("AND2X1_LOC_154/Y") V("OR2X1_LOC_189/A") V("OR2X1_LOC_393/Y") V("OR2X1_LOC_595/A") V("AND2X1_LOC_391/Y") V("OR2X1_LOC_823/Y") V("OR2X1_LOC_697/Y") V("OR2X1_LOC_759/Y") V("OR2X1_LOC_34/A") V("OR2X1_LOC_134/Y") V("OR2X1_LOC_427/Y") V("OR2X1_LOC_679/B") V("OR2X1_LOC_754/A") V("OR2X1_LOC_227/Y") V("OR2X1_LOC_446/Y") V("OR2X1_LOC_714/A") V("OR2X1_LOC_338/B") V("OR2X1_LOC_772/B") V("OR2X1_LOC_286/Y") V("OR2X1_LOC_787/B") V("OR2X1_LOC_516/Y") V("OR2X1_LOC_715/B") V("OR2X1_LOC_339/A") V("OR2X1_LOC_550/A") V("OR2X1_LOC_856/A") V("OR2X1_LOC_730/A") V("AND2X1_LOC_462/Y") V("AND2X1_LOC_240/Y") V("AND2X1_LOC_839/B") V("AND2X1_LOC_334/Y") V("OR2X1_LOC_710/A") V("OR2X1_LOC_792/B") V("OR2X1_LOC_836/B") V("OR2X1_LOC_779/A") V("OR2X1_LOC_542/B") V("OR2X1_LOC_383/Y") V("OR2X1_LOC_451/B") V("OR2X1_LOC_636/B") V("OR2X1_LOC_523/B") V("OR2X1_LOC_782/B") V("AND2X1_LOC_52/Y") V("OR2X1_LOC_545/A") V("OR2X1_LOC_676/Y") V("OR2X1_LOC_318/B") V("OR2X1_LOC_614/Y") V("OR2X1_LOC_259/B") V("OR2X1_LOC_131/A") V("OR2X1_LOC_586/Y") V("AND2X1_LOC_789/Y") V("OR2X1_LOC_348/B") V("OR2X1_LOC_423/Y") V("OR2X1_LOC_7/Y") V("OR2X1_LOC_584/Y") V("OR2X1_LOC_248/A") V("OR2X1_LOC_183/Y") V("OR2X1_LOC_33/B") V("OR2X1_LOC_561/B") V("OR2X1_LOC_127/Y") V("OR2X1_LOC_698/Y") V("OR2X1_LOC_764/Y") V("OR2X1_LOC_380/Y") V("OR2X1_LOC_757/A") V("OR2X1_LOC_125/Y") V("OR2X1_LOC_442/Y") V("OR2X1_LOC_261/Y") V("OR2X1_LOC_106/A") V("AND2X1_LOC_216/A") V("OR2X1_LOC_473/Y") V("OR2X1_LOC_362/A") V("OR2X1_LOC_574/A") V("OR2X1_LOC_810/A") V("AND2X1_LOC_79/Y") V("OR2X1_LOC_719/A") V("OR2X1_LOC_778/A") V("OR2X1_LOC_435/B") V("OR2X1_LOC_646/B") V("OR2X1_LOC_790/A") V("OR2X1_LOC_324/B") V("OR2X1_LOC_148/A") V("AND2X1_LOC_39/Y") V("OR2X1_LOC_499/B") V("OR2X1_LOC_781/A") V("OR2X1_LOC_181/B") V("OR2X1_LOC_210/B") V("OR2X1_LOC_462/B") V("OR2X1_LOC_259/A") V("OR2X1_LOC_518/Y") V("OR2X1_LOC_167/Y") V("OR2X1_LOC_667/Y") V("OR2X1_LOC_250/Y") V("OR2X1_LOC_829/Y") V("OR2X1_LOC_591/Y") V("OR2X1_LOC_321/Y") V("OR2X1_LOC_503/Y") V("OR2X1_LOC_142/Y") V("OR2X1_LOC_189/Y") V("OR2X1_LOC_759/A") V("OR2X1_LOC_487/Y") V("OR2X1_LOC_406/Y") V("OR2X1_LOC_96/Y") V("OR2X1_LOC_594/Y") V("OR2X1_LOC_533/Y") V("OR2X1_LOC_165/Y") V("OR2X1_LOC_145/Y") V("OR2X1_LOC_680/Y") V("OR2X1_LOC_251/Y") V("OR2X1_LOC_418/Y") V("OR2X1_LOC_52/Y") V("OR2X1_LOC_238/Y") V("OR2X1_LOC_525/Y") V("OR2X1_LOC_163/Y") V("AND2X1_LOC_451/Y") V("AND2X1_LOC_463/B") V("OR2X1_LOC_771/B") V("OR2X1_LOC_639/B") V("OR2X1_LOC_793/A") V("OR2X1_LOC_400/A") V("OR2X1_LOC_209/A") V("OR2X1_LOC_113/B") V("OR2X1_LOC_115/B") V("OR2X1_LOC_342/A") V("OR2X1_LOC_780/A") V("OR2X1_LOC_791/A") V("OR2X1_LOC_403/B") V("OR2X1_LOC_124/B") V("OR2X1_LOC_705/B") V("OR2X1_LOC_347/B") V("OR2X1_LOC_449/A") V("OR2X1_LOC_76/B") V("OR2X1_LOC_559/B") V("OR2X1_LOC_493/B") V("OR2X1_LOC_112/B") V("OR2X1_LOC_302/B") V("OR2X1_LOC_227/B") V("OR2X1_LOC_97/A") V("OR2X1_LOC_467/B") V("OR2X1_LOC_168/A") V("OR2X1_LOC_148/B") V("OR2X1_LOC_728/A") V("OR2X1_LOC_843/B") V("OR2X1_LOC_506/B") V("AND2X1_LOC_450/Y") V("AND2X1_LOC_707/Y") V("OR2X1_LOC_187/Y") V("OR2X1_LOC_166/Y") V("OR2X1_LOC_441/Y") V("OR2X1_LOC_265/Y") V("OR2X1_LOC_41/Y") V("OR2X1_LOC_745/Y") V("OR2X1_LOC_531/Y") V("OR2X1_LOC_384/Y") V("OR2X1_LOC_171/Y") V("OR2X1_LOC_665/Y") V("OR2X1_LOC_751/Y") V("OR2X1_LOC_767/Y") V("OR2X1_LOC_16/Y") V("OR2X1_LOC_397/Y") V("OR2X1_LOC_177/Y") V("OR2X1_LOC_821/Y") V("OR2X1_LOC_118/Y") V("OR2X1_LOC_674/Y") V("OR2X1_LOC_498/Y") V("OR2X1_LOC_604/Y") V("OR2X1_LOC_438/Y") V("OR2X1_LOC_158/Y") V("OR2X1_LOC_232/Y") V("OR2X1_LOC_258/Y") V("OR2X1_LOC_746/Y") V("OR2X1_LOC_504/Y") V("AND2X1_LOC_197/Y") V("AND2X1_LOC_307/Y") V("AND2X1_LOC_356/B") V("OR2X1_LOC_597/Y") V("AND2X1_LOC_390/B") V("OR2X1_LOC_392/A") V("OR2X1_LOC_549/Y") V("OR2X1_LOC_784/B") V("OR2X1_LOC_633/Y") V("OR2X1_LOC_553/A") V("OR2X1_LOC_640/A") V("OR2X1_LOC_845/A") V("OR2X1_LOC_188/Y") V("OR2X1_LOC_590/Y") V("OR2X1_LOC_460/B") V("OR2X1_LOC_532/Y") V("OR2X1_LOC_243/B") V("OR2X1_LOC_664/Y") V("OR2X1_LOC_151/Y") V("AND2X1_LOC_624/A") V("OR2X1_LOC_79/A") V("OR2X1_LOC_755/A") V("AND2X1_LOC_711/A") V("AND2X1_LOC_706/Y") V("OR2X1_LOC_673/Y") V("AND2X1_LOC_776/Y") V("AND2X1_LOC_168/Y") V("AND2X1_LOC_326/B") V("AND2X1_LOC_459/Y") V("AND2X1_LOC_638/Y") V("AND2X1_LOC_712/B") V("AND2X1_LOC_727/A") V("AND2X1_LOC_147/Y") V("OR2X1_LOC_630/Y") V("OR2X1_LOC_390/A") V("OR2X1_LOC_506/Y") V("OR2X1_LOC_447/Y") V("OR2X1_LOC_852/B") V("OR2X1_LOC_139/A") V("OR2X1_LOC_199/B") V("OR2X1_LOC_854/A") V("AND2X1_LOC_67/Y") V("OR2X1_LOC_612/Y") V("AND2X1_LOC_848/Y") V("OR2X1_LOC_450/Y") V("OR2X1_LOC_303/A") V("OR2X1_LOC_552/A") V("OR2X1_LOC_303/B") V("AND2X1_LOC_227/Y") V("AND2X1_LOC_714/B") V("AND2X1_LOC_454/A") V("AND2X1_LOC_338/A") V("AND2X1_LOC_489/Y") V("AND2X1_LOC_286/Y") V("OR2X1_LOC_632/A") V("OR2X1_LOC_637/Y") V("OR2X1_LOC_850/A") V("OR2X1_LOC_288/A") V("OR2X1_LOC_609/A") V("AND2X1_LOC_342/Y") V("OR2X1_LOC_669/Y") V("AND2X1_LOC_779/Y") V("AND2X1_LOC_840/B") V("AND2X1_LOC_196/Y") V("AND2X1_LOC_769/Y") V("OR2X1_LOC_829/A") V("AND2X1_LOC_520/Y") V("AND2X1_LOC_464/Y") V("AND2X1_LOC_783/B") V("AND2X1_LOC_841/B") V("OR2X1_LOC_158/B") V("AND2X1_LOC_339/B") V("AND2X1_LOC_715/A") V("AND2X1_LOC_547/Y") V("AND2X1_LOC_729/Y") V("AND2X1_LOC_856/B") V("OR2X1_LOC_656/B") V("AND2X1_LOC_362/B") V("AND2X1_LOC_473/Y") V("AND2X1_LOC_810/B") V("OR2X1_LOC_472/B") V("OR2X1_LOC_243/A") V("OR2X1_LOC_836/Y") V("OR2X1_LOC_338/A") V("AND2X1_LOC_687/Y") V("OR2X1_LOC_687/Y") V("AND2X1_LOC_456/B") V("OR2X1_LOC_456/A") V("AND2X1_LOC_99/A") V("OR2X1_LOC_802/A") V("OR2X1_LOC_798/Y") V("OR2X1_LOC_99/B") V("AND2X1_LOC_798/Y") V("AND2X1_LOC_802/B") V("OR2X1_LOC_113/Y") V("OR2X1_LOC_539/Y") V("OR2X1_LOC_319/Y") V("AND2X1_LOC_113/Y") V("AND2X1_LOC_798/A") V("AND2X1_LOC_539/Y") V("OR2X1_LOC_593/A") V("OR2X1_LOC_539/B") V("OR2X1_LOC_436/B") V("AND2X1_LOC_434/Y") V("AND2X1_LOC_537/Y") V("AND2X1_LOC_592/Y") V("AND2X1_LOC_593/Y") V("OR2X1_LOC_799/A") V("OR2X1_LOC_216/A") V("OR2X1_LOC_88/Y") V("AND2X1_LOC_374/Y") V("OR2X1_LOC_599/Y") V("OR2X1_LOC_373/Y") V("OR2X1_LOC_644/A") V("AND2X1_LOC_116/Y") V("AND2X1_LOC_88/Y") V("OR2X1_LOC_374/Y") V("OR2X1_LOC_254/B") V("OR2X1_LOC_252/Y") V("OR2X1_LOC_544/B") V("AND2X1_LOC_361/A") V("AND2X1_LOC_483/Y") V("AND2X1_LOC_436/Y") V("OR2X1_LOC_631/B") V("OR2X1_LOC_436/Y") V("OR2X1_LOC_267/Y") 

* SUBCKT HEAD: NAME;  INPUTS; POWER; OUTPUTS
.subckt AES_SBOX_2
+ OR2X1_LOC_452/A AND2X1_LOC_639/A OR2X1_LOC_460/Y OR2X1_LOC_198/A OR2X1_LOC_308/A OR2X1_LOC_379/Y OR2X1_LOC_643/A OR2X1_LOC_84/A OR2X1_LOC_538/A OR2X1_LOC_180/B OR2X1_LOC_668/Y OR2X1_LOC_34/B OR2X1_LOC_334/B OR2X1_LOC_834/A OR2X1_LOC_241/B OR2X1_LOC_523/A OR2X1_LOC_33/A OR2X1_LOC_61/B OR2X1_LOC_844/B OR2X1_LOC_623/B OR2X1_LOC_770/A OR2X1_LOC_324/A OR2X1_LOC_509/A OR2X1_LOC_703/A OR2X1_LOC_147/B OR2X1_LOC_201/A OR2X1_LOC_520/B OR2X1_LOC_703/B OR2X1_LOC_835/A OR2X1_LOC_709/B OR2X1_LOC_720/B OR2X1_LOC_343/B OR2X1_LOC_855/A OR2X1_LOC_449/B OR2X1_LOC_593/B OR2X1_LOC_773/B OR2X1_LOC_402/B OR2X1_LOC_307/A OR2X1_LOC_128/A OR2X1_LOC_194/B OR2X1_LOC_555/A OR2X1_LOC_719/B AND2X1_LOC_7/Y OR2X1_LOC_789/A OR2X1_LOC_769/A OR2X1_LOC_400/B OR2X1_LOC_781/B OR2X1_LOC_549/B OR2X1_LOC_391/A OR2X1_LOC_333/B OR2X1_LOC_190/B 
+ AND2X1_LOC_41/Y OR2X1_LOC_610/Y OR2X1_LOC_191/B OR2X1_LOC_169/B OR2X1_LOC_673/B OR2X1_LOC_346/B OR2X1_LOC_545/B OR2X1_LOC_444/B OR2X1_LOC_620/A OR2X1_LOC_786/A OR2X1_LOC_641/A OR2X1_LOC_758/Y OR2X1_LOC_637/A OR2X1_LOC_174/A AND2X1_LOC_72/Y OR2X1_LOC_175/B OR2X1_LOC_439/B OR2X1_LOC_835/B OR2X1_LOC_123/B OR2X1_LOC_633/B OR2X1_LOC_675/A OR2X1_LOC_501/B OR2X1_LOC_605/A OR2X1_LOC_544/A OR2X1_LOC_450/A OR2X1_LOC_103/Y OR2X1_LOC_106/Y OR2X1_LOC_695/Y OR2X1_LOC_280/Y OR2X1_LOC_601/Y OR2X1_LOC_612/B OR2X1_LOC_248/Y OR2X1_LOC_394/Y OR2X1_LOC_747/Y OR2X1_LOC_524/Y OR2X1_LOC_152/Y OR2X1_LOC_528/Y OR2X1_LOC_122/Y OR2X1_LOC_485/Y OR2X1_LOC_297/Y OR2X1_LOC_424/Y OR2X1_LOC_45/Y OR2X1_LOC_744/Y OR2X1_LOC_701/Y OR2X1_LOC_757/Y OR2X1_LOC_399/Y OR2X1_LOC_517/Y OR2X1_LOC_315/Y OR2X1_LOC_491/Y OR2X1_LOC_109/Y OR2X1_LOC_600/Y 
+ OR2X1_LOC_230/Y OR2X1_LOC_298/Y OR2X1_LOC_224/Y OR2X1_LOC_428/Y OR2X1_LOC_74/Y OR2X1_LOC_32/Y OR2X1_LOC_583/Y OR2X1_LOC_526/Y OR2X1_LOC_505/Y OR2X1_LOC_666/Y OR2X1_LOC_496/Y OR2X1_LOC_432/Y OR2X1_LOC_607/Y OR2X1_LOC_257/Y OR2X1_LOC_20/Y OR2X1_LOC_79/Y OR2X1_LOC_521/Y OR2X1_LOC_135/Y OR2X1_LOC_492/Y OR2X1_LOC_482/Y OR2X1_LOC_108/Y OR2X1_LOC_295/Y OR2X1_LOC_81/Y OR2X1_LOC_60/Y OR2X1_LOC_437/Y OR2X1_LOC_609/Y OR2X1_LOC_75/Y OR2X1_LOC_700/Y OR2X1_LOC_755/Y OR2X1_LOC_395/Y OR2X1_LOC_494/Y OR2X1_LOC_380/A OR2X1_LOC_603/Y OR2X1_LOC_261/A OR2X1_LOC_679/A OR2X1_LOC_229/Y OR2X1_LOC_13/Y OR2X1_LOC_765/Y OR2X1_LOC_131/Y AND2X1_LOC_793/B OR2X1_LOC_712/B OR2X1_LOC_791/B OR2X1_LOC_710/B OR2X1_LOC_401/B OR2X1_LOC_84/B OR2X1_LOC_61/A OR2X1_LOC_76/A OR2X1_LOC_702/A OR2X1_LOC_493/A OR2X1_LOC_833/B OR2X1_LOC_114/B 
+ OR2X1_LOC_346/A OR2X1_LOC_440/B OR2X1_LOC_646/A OR2X1_LOC_231/B OR2X1_LOC_770/B OR2X1_LOC_140/A OR2X1_LOC_260/Y OR2X1_LOC_678/Y OR2X1_LOC_193/A OR2X1_LOC_558/A OR2X1_LOC_605/B OR2X1_LOC_653/B OR2X1_LOC_788/B OR2X1_LOC_190/A OR2X1_LOC_98/A OR2X1_LOC_137/B OR2X1_LOC_192/B OR2X1_LOC_768/A OR2X1_LOC_128/B OR2X1_LOC_447/A OR2X1_LOC_489/B OR2X1_LOC_475/B OR2X1_LOC_644/B OR2X1_LOC_448/Y OR2X1_LOC_356/A OR2X1_LOC_176/Y OR2X1_LOC_290/Y OR2X1_LOC_677/Y OR2X1_LOC_83/Y OR2X1_LOC_237/Y OR2X1_LOC_669/A OR2X1_LOC_595/Y OR2X1_LOC_27/Y OR2X1_LOC_311/Y OR2X1_LOC_146/Y OR2X1_LOC_179/Y OR2X1_LOC_484/Y OR2X1_LOC_495/Y OR2X1_LOC_754/Y OR2X1_LOC_69/Y OR2X1_LOC_39/Y OR2X1_LOC_396/Y OR2X1_LOC_320/Y OR2X1_LOC_497/Y OR2X1_LOC_615/Y OR2X1_LOC_24/Y OR2X1_LOC_58/Y OR2X1_LOC_522/Y AND2X1_LOC_549/Y OR2X1_LOC_711/B OR2X1_LOC_713/A 
+ AND2X1_LOC_335/Y AND2X1_LOC_778/Y AND2X1_LOC_208/B OR2X1_LOC_72/Y OR2X1_LOC_184/Y OR2X1_LOC_152/A OR2X1_LOC_292/Y OR2X1_LOC_173/Y OR2X1_LOC_235/Y AND2X1_LOC_784/A AND2X1_LOC_633/Y AND2X1_LOC_541/Y AND2X1_LOC_634/Y OR2X1_LOC_813/Y OR2X1_LOC_624/B AND2X1_LOC_721/A AND2X1_LOC_69/Y OR2X1_LOC_208/A OR2X1_LOC_335/Y OR2X1_LOC_778/Y OR2X1_LOC_117/Y OR2X1_LOC_262/Y OR2X1_LOC_65/Y OR2X1_LOC_471/B AND2X1_LOC_303/A AND2X1_LOC_831/Y AND2X1_LOC_303/B AND2X1_LOC_787/A AND2X1_LOC_543/Y OR2X1_LOC_841/A OR2X1_LOC_841/B OR2X1_LOC_828/Y OR2X1_LOC_783/A OR2X1_LOC_156/Y OR2X1_LOC_708/Y OR2X1_LOC_308/Y OR2X1_LOC_149/B OR2X1_LOC_168/Y OR2X1_LOC_776/Y OR2X1_LOC_325/Y OR2X1_LOC_463/B OR2X1_LOC_651/B OR2X1_LOC_416/Y AND2X1_LOC_637/Y OR2X1_LOC_481/Y AND2X1_LOC_631/Y OR2X1_LOC_196/Y OR2X1_LOC_520/Y OR2X1_LOC_840/A OR2X1_LOC_779/Y AND2X1_LOC_632/A 
+ AND2X1_LOC_448/Y OR2X1_LOC_156/B OR2X1_LOC_636/A OR2X1_LOC_620/B OR2X1_LOC_247/Y OR2X1_LOC_231/A OR2X1_LOC_130/Y AND2X1_LOC_348/A OR2X1_LOC_105/Y OR2X1_LOC_181/A OR2X1_LOC_602/B OR2X1_LOC_345/A OR2X1_LOC_756/Y OR2X1_LOC_401/A OR2X1_LOC_507/A OR2X1_LOC_196/B OR2X1_LOC_707/A OR2X1_LOC_249/Y OR2X1_LOC_776/A OR2X1_LOC_793/B AND2X1_LOC_557/Y AND2X1_LOC_535/Y AND2X1_LOC_199/A AND2X1_LOC_508/A AND2X1_LOC_447/Y AND2X1_LOC_838/Y AND2X1_LOC_139/B OR2X1_LOC_178/Y OR2X1_LOC_613/Y OR2X1_LOC_67/Y OR2X1_LOC_312/Y OR2X1_LOC_647/B OR2X1_LOC_132/Y OR2X1_LOC_305/Y OR2X1_LOC_494/A OR2X1_LOC_91/Y OR2X1_LOC_766/Y OR2X1_LOC_670/Y OR2X1_LOC_533/A OR2X1_LOC_822/Y OR2X1_LOC_420/Y OR2X1_LOC_239/Y OR2X1_LOC_172/Y OR2X1_LOC_591/A OR2X1_LOC_349/B AND2X1_LOC_843/Y AND2X1_LOC_287/Y OR2X1_LOC_608/Y OR2X1_LOC_602/A OR2X1_LOC_78/Y OR2X1_LOC_240/B 
+ OR2X1_LOC_446/A OR2X1_LOC_546/A OR2X1_LOC_720/A OR2X1_LOC_546/B OR2X1_LOC_507/B OR2X1_LOC_486/B OR2X1_LOC_859/B AND2X1_LOC_154/Y OR2X1_LOC_189/A OR2X1_LOC_393/Y OR2X1_LOC_595/A AND2X1_LOC_391/Y OR2X1_LOC_823/Y OR2X1_LOC_697/Y OR2X1_LOC_759/Y OR2X1_LOC_34/A OR2X1_LOC_134/Y OR2X1_LOC_427/Y OR2X1_LOC_679/B OR2X1_LOC_754/A OR2X1_LOC_227/Y OR2X1_LOC_446/Y OR2X1_LOC_714/A OR2X1_LOC_338/B OR2X1_LOC_772/B OR2X1_LOC_286/Y OR2X1_LOC_787/B OR2X1_LOC_516/Y OR2X1_LOC_715/B OR2X1_LOC_339/A OR2X1_LOC_550/A OR2X1_LOC_856/A OR2X1_LOC_730/A AND2X1_LOC_462/Y AND2X1_LOC_240/Y AND2X1_LOC_839/B AND2X1_LOC_334/Y OR2X1_LOC_710/A OR2X1_LOC_792/B OR2X1_LOC_836/B OR2X1_LOC_779/A OR2X1_LOC_542/B OR2X1_LOC_383/Y OR2X1_LOC_451/B OR2X1_LOC_636/B OR2X1_LOC_523/B OR2X1_LOC_782/B AND2X1_LOC_52/Y OR2X1_LOC_545/A OR2X1_LOC_676/Y OR2X1_LOC_318/B 
+ OR2X1_LOC_614/Y OR2X1_LOC_259/B OR2X1_LOC_131/A OR2X1_LOC_586/Y AND2X1_LOC_789/Y OR2X1_LOC_348/B OR2X1_LOC_423/Y OR2X1_LOC_7/Y OR2X1_LOC_584/Y OR2X1_LOC_248/A OR2X1_LOC_183/Y OR2X1_LOC_33/B OR2X1_LOC_561/B OR2X1_LOC_127/Y OR2X1_LOC_698/Y OR2X1_LOC_764/Y OR2X1_LOC_380/Y OR2X1_LOC_757/A OR2X1_LOC_125/Y OR2X1_LOC_442/Y OR2X1_LOC_261/Y OR2X1_LOC_106/A AND2X1_LOC_216/A OR2X1_LOC_473/Y OR2X1_LOC_362/A OR2X1_LOC_574/A OR2X1_LOC_810/A AND2X1_LOC_79/Y OR2X1_LOC_719/A OR2X1_LOC_778/A OR2X1_LOC_435/B OR2X1_LOC_646/B OR2X1_LOC_790/A OR2X1_LOC_324/B OR2X1_LOC_148/A AND2X1_LOC_39/Y OR2X1_LOC_499/B OR2X1_LOC_781/A OR2X1_LOC_181/B OR2X1_LOC_210/B OR2X1_LOC_462/B OR2X1_LOC_259/A OR2X1_LOC_518/Y OR2X1_LOC_167/Y OR2X1_LOC_667/Y OR2X1_LOC_250/Y OR2X1_LOC_829/Y OR2X1_LOC_591/Y OR2X1_LOC_321/Y OR2X1_LOC_503/Y OR2X1_LOC_142/Y 
+ OR2X1_LOC_189/Y OR2X1_LOC_759/A OR2X1_LOC_487/Y OR2X1_LOC_406/Y OR2X1_LOC_96/Y OR2X1_LOC_594/Y OR2X1_LOC_533/Y OR2X1_LOC_165/Y OR2X1_LOC_145/Y OR2X1_LOC_680/Y OR2X1_LOC_251/Y OR2X1_LOC_418/Y OR2X1_LOC_52/Y OR2X1_LOC_238/Y OR2X1_LOC_525/Y OR2X1_LOC_163/Y AND2X1_LOC_451/Y AND2X1_LOC_463/B OR2X1_LOC_771/B OR2X1_LOC_639/B OR2X1_LOC_793/A OR2X1_LOC_400/A OR2X1_LOC_209/A OR2X1_LOC_113/B OR2X1_LOC_115/B OR2X1_LOC_342/A OR2X1_LOC_780/A OR2X1_LOC_791/A OR2X1_LOC_403/B OR2X1_LOC_124/B OR2X1_LOC_705/B OR2X1_LOC_347/B OR2X1_LOC_449/A OR2X1_LOC_76/B OR2X1_LOC_559/B OR2X1_LOC_493/B OR2X1_LOC_112/B OR2X1_LOC_302/B OR2X1_LOC_227/B OR2X1_LOC_97/A OR2X1_LOC_467/B OR2X1_LOC_168/A OR2X1_LOC_148/B OR2X1_LOC_728/A OR2X1_LOC_843/B OR2X1_LOC_506/B AND2X1_LOC_450/Y AND2X1_LOC_707/Y OR2X1_LOC_187/Y OR2X1_LOC_166/Y OR2X1_LOC_441/Y 
+ OR2X1_LOC_265/Y OR2X1_LOC_41/Y OR2X1_LOC_745/Y OR2X1_LOC_531/Y OR2X1_LOC_384/Y OR2X1_LOC_171/Y OR2X1_LOC_665/Y OR2X1_LOC_751/Y OR2X1_LOC_767/Y OR2X1_LOC_16/Y OR2X1_LOC_397/Y OR2X1_LOC_177/Y OR2X1_LOC_821/Y OR2X1_LOC_118/Y OR2X1_LOC_674/Y OR2X1_LOC_498/Y OR2X1_LOC_604/Y OR2X1_LOC_438/Y OR2X1_LOC_158/Y OR2X1_LOC_232/Y OR2X1_LOC_258/Y OR2X1_LOC_746/Y OR2X1_LOC_504/Y AND2X1_LOC_197/Y AND2X1_LOC_307/Y AND2X1_LOC_356/B OR2X1_LOC_597/Y AND2X1_LOC_390/B OR2X1_LOC_392/A OR2X1_LOC_549/Y OR2X1_LOC_784/B OR2X1_LOC_633/Y OR2X1_LOC_553/A OR2X1_LOC_640/A OR2X1_LOC_845/A OR2X1_LOC_188/Y OR2X1_LOC_590/Y OR2X1_LOC_460/B OR2X1_LOC_532/Y OR2X1_LOC_243/B OR2X1_LOC_664/Y OR2X1_LOC_151/Y AND2X1_LOC_624/A OR2X1_LOC_79/A OR2X1_LOC_755/A AND2X1_LOC_711/A AND2X1_LOC_706/Y OR2X1_LOC_673/Y AND2X1_LOC_776/Y AND2X1_LOC_168/Y AND2X1_LOC_326/B 
+ AND2X1_LOC_459/Y AND2X1_LOC_638/Y AND2X1_LOC_712/B AND2X1_LOC_727/A AND2X1_LOC_147/Y OR2X1_LOC_630/Y OR2X1_LOC_390/A OR2X1_LOC_506/Y OR2X1_LOC_447/Y OR2X1_LOC_852/B OR2X1_LOC_139/A OR2X1_LOC_199/B OR2X1_LOC_854/A AND2X1_LOC_67/Y OR2X1_LOC_612/Y AND2X1_LOC_848/Y OR2X1_LOC_450/Y OR2X1_LOC_303/A OR2X1_LOC_552/A OR2X1_LOC_303/B AND2X1_LOC_227/Y AND2X1_LOC_714/B AND2X1_LOC_454/A AND2X1_LOC_338/A AND2X1_LOC_489/Y AND2X1_LOC_286/Y OR2X1_LOC_632/A OR2X1_LOC_637/Y OR2X1_LOC_850/A OR2X1_LOC_288/A OR2X1_LOC_609/A AND2X1_LOC_342/Y OR2X1_LOC_669/Y AND2X1_LOC_779/Y AND2X1_LOC_840/B AND2X1_LOC_196/Y AND2X1_LOC_769/Y OR2X1_LOC_829/A AND2X1_LOC_520/Y AND2X1_LOC_464/Y AND2X1_LOC_783/B AND2X1_LOC_841/B OR2X1_LOC_158/B AND2X1_LOC_339/B AND2X1_LOC_715/A AND2X1_LOC_547/Y AND2X1_LOC_729/Y AND2X1_LOC_856/B OR2X1_LOC_656/B AND2X1_LOC_362/B AND2X1_LOC_473/Y 
+ AND2X1_LOC_810/B OR2X1_LOC_472/B OR2X1_LOC_243/A OR2X1_LOC_836/Y OR2X1_LOC_338/A AND2X1_LOC_687/Y OR2X1_LOC_687/Y AND2X1_LOC_456/B OR2X1_LOC_456/A AND2X1_LOC_99/A OR2X1_LOC_802/A OR2X1_LOC_798/Y OR2X1_LOC_99/B AND2X1_LOC_798/Y AND2X1_LOC_802/B OR2X1_LOC_113/Y OR2X1_LOC_539/Y OR2X1_LOC_319/Y AND2X1_LOC_113/Y AND2X1_LOC_798/A AND2X1_LOC_539/Y OR2X1_LOC_593/A OR2X1_LOC_539/B OR2X1_LOC_436/B AND2X1_LOC_434/Y AND2X1_LOC_537/Y AND2X1_LOC_592/Y AND2X1_LOC_593/Y OR2X1_LOC_799/A OR2X1_LOC_216/A OR2X1_LOC_88/Y AND2X1_LOC_374/Y OR2X1_LOC_599/Y OR2X1_LOC_373/Y OR2X1_LOC_644/A AND2X1_LOC_116/Y AND2X1_LOC_88/Y OR2X1_LOC_374/Y OR2X1_LOC_254/B OR2X1_LOC_252/Y OR2X1_LOC_544/B AND2X1_LOC_361/A AND2X1_LOC_483/Y AND2X1_LOC_436/Y OR2X1_LOC_631/B OR2X1_LOC_436/Y OR2X1_LOC_267/Y 
+ VSS VDD 
+ OR2X1_LOC_351/B OR2X1_LOC_852/A OR2X1_LOC_244/A OR2X1_LOC_476/B AND2X1_LOC_810/Y AND2X1_LOC_476/Y AND2X1_LOC_366/A OR2X1_LOC_656/Y OR2X1_LOC_216/Y AND2X1_LOC_863/A AND2X1_LOC_739/B AND2X1_LOC_565/B AND2X1_LOC_715/Y AND2X1_LOC_339/Y AND2X1_LOC_851/B AND2X1_LOC_796/A AND2X1_LOC_471/Y AND2X1_LOC_560/B AND2X1_LOC_642/Y AND2X1_LOC_207/A AND2X1_LOC_851/A AND2X1_LOC_720/Y AND2X1_LOC_359/B OR2X1_LOC_362/B OR2X1_LOC_858/B OR2X1_LOC_632/Y AND2X1_LOC_806/A AND2X1_LOC_772/Y AND2X1_LOC_338/Y AND2X1_LOC_454/Y AND2X1_LOC_724/A AND2X1_LOC_340/Y OR2X1_LOC_566/A OR2X1_LOC_723/B OR2X1_LOC_564/A OR2X1_LOC_467/A AND2X1_LOC_859/Y AND2X1_LOC_647/Y OR2X1_LOC_206/A OR2X1_LOC_856/B OR2X1_LOC_568/A OR2X1_LOC_207/B OR2X1_LOC_141/B OR2X1_LOC_857/B OR2X1_LOC_466/A OR2X1_LOC_392/B AND2X1_LOC_797/A AND2X1_LOC_357/B AND2X1_LOC_727/Y AND2X1_LOC_712/Y AND2X1_LOC_654/B 
+ AND2X1_LOC_472/B AND2X1_LOC_717/Y AND2X1_LOC_170/Y AND2X1_LOC_785/Y OR2X1_LOC_721/Y AND2X1_LOC_713/Y AND2X1_LOC_711/Y AND2X1_LOC_658/A OR2X1_LOC_640/Y OR2X1_LOC_563/B OR2X1_LOC_784/Y OR2X1_LOC_569/A OR2X1_LOC_474/B AND2X1_LOC_392/A AND2X1_LOC_644/Y AND2X1_LOC_365/A AND2X1_LOC_508/B AND2X1_LOC_781/Y AND2X1_LOC_259/Y AND2X1_LOC_213/B AND2X1_LOC_544/Y AND2X1_LOC_675/A AND2X1_LOC_605/Y AND2X1_LOC_501/Y AND2X1_LOC_675/Y AND2X1_LOC_123/Y AND2X1_LOC_839/A AND2X1_LOC_182/A AND2X1_LOC_194/Y AND2X1_LOC_719/Y AND2X1_LOC_175/B AND2X1_LOC_641/Y AND2X1_LOC_551/B AND2X1_LOC_443/Y AND2X1_LOC_170/B AND2X1_LOC_191/Y AND2X1_LOC_452/Y OR2X1_LOC_244/B OR2X1_LOC_349/A OR2X1_LOC_730/B OR2X1_LOC_148/Y OR2X1_LOC_470/A OR2X1_LOC_213/A OR2X1_LOC_443/Y OR2X1_LOC_785/B OR2X1_LOC_493/Y OR2X1_LOC_560/A OR2X1_LOC_453/A OR2X1_LOC_347/Y OR2X1_LOC_486/Y OR2X1_LOC_705/Y 
+ OR2X1_LOC_124/Y OR2X1_LOC_792/A OR2X1_LOC_563/A OR2X1_LOC_772/A OR2X1_LOC_213/B OR2X1_LOC_731/B OR2X1_LOC_403/A OR2X1_LOC_805/A OR2X1_LOC_651/A AND2X1_LOC_470/B AND2X1_LOC_550/A AND2X1_LOC_242/B AND2X1_LOC_228/Y AND2X1_LOC_349/B AND2X1_LOC_728/Y AND2X1_LOC_148/Y AND2X1_LOC_794/B AND2X1_LOC_661/A AND2X1_LOC_734/Y AND2X1_LOC_475/Y AND2X1_LOC_192/Y AND2X1_LOC_842/B AND2X1_LOC_326/A AND2X1_LOC_722/A AND2X1_LOC_703/Y AND2X1_LOC_388/Y OR2X1_LOC_555/B OR2X1_LOC_649/B OR2X1_LOC_553/B OR2X1_LOC_181/Y OR2X1_LOC_781/Y OR2X1_LOC_833/Y OR2X1_LOC_500/A OR2X1_LOC_194/Y OR2X1_LOC_326/B OR2X1_LOC_648/B OR2X1_LOC_647/A OR2X1_LOC_719/Y OR2X1_LOC_204/Y OR2X1_LOC_812/B OR2X1_LOC_575/A OR2X1_LOC_366/B OR2X1_LOC_476/Y AND2X1_LOC_656/Y AND2X1_LOC_216/Y AND2X1_LOC_345/Y AND2X1_LOC_727/B AND2X1_LOC_554/B OR2X1_LOC_561/Y AND2X1_LOC_553/A AND2X1_LOC_191/B 
+ AND2X1_LOC_639/B AND2X1_LOC_193/Y AND2X1_LOC_449/Y OR2X1_LOC_348/Y AND2X1_LOC_793/Y OR2X1_LOC_728/B OR2X1_LOC_551/A OR2X1_LOC_228/Y OR2X1_LOC_797/A OR2X1_LOC_523/Y OR2X1_LOC_639/A OR2X1_LOC_552/B OR2X1_LOC_792/Y OR2X1_LOC_711/A AND2X1_LOC_852/B AND2X1_LOC_243/Y AND2X1_LOC_476/A OR2X1_LOC_739/A OR2X1_LOC_863/B OR2X1_LOC_565/A OR2X1_LOC_339/Y OR2X1_LOC_724/A AND2X1_LOC_574/Y OR2X1_LOC_787/Y OR2X1_LOC_772/Y OR2X1_LOC_714/Y OR2X1_LOC_340/Y OR2X1_LOC_679/Y AND2X1_LOC_772/B AND2X1_LOC_139/A AND2X1_LOC_792/Y AND2X1_LOC_474/A AND2X1_LOC_403/B OR2X1_LOC_862/A OR2X1_LOC_508/A OR2X1_LOC_550/B OR2X1_LOC_720/Y OR2X1_LOC_602/Y AND2X1_LOC_850/Y OR2X1_LOC_359/A AND2X1_LOC_244/A AND2X1_LOC_771/B AND2X1_LOC_785/A OR2X1_LOC_647/Y AND2X1_LOC_552/A AND2X1_LOC_337/B AND2X1_LOC_202/Y AND2X1_LOC_620/Y AND2X1_LOC_181/Y AND2X1_LOC_141/A AND2X1_LOC_852/Y 
+ AND2X1_LOC_568/B AND2X1_LOC_856/A AND2X1_LOC_571/B OR2X1_LOC_241/Y OR2X1_LOC_715/A OR2X1_LOC_401/Y OR2X1_LOC_345/Y AND2X1_LOC_348/Y OR2X1_LOC_641/B OR2X1_LOC_620/Y AND2X1_LOC_453/Y AND2X1_LOC_658/B OR2X1_LOC_796/B OR2X1_LOC_851/B AND2X1_LOC_555/Y OR2X1_LOC_654/A OR2X1_LOC_472/A OR2X1_LOC_723/A OR2X1_LOC_795/B OR2X1_LOC_170/Y OR2X1_LOC_797/B OR2X1_LOC_357/A OR2X1_LOC_731/A OR2X1_LOC_725/B OR2X1_LOC_851/A AND2X1_LOC_564/B AND2X1_LOC_794/A AND2X1_LOC_566/B AND2X1_LOC_716/Y OR2X1_LOC_471/Y AND2X1_LOC_201/Y AND2X1_LOC_786/Y OR2X1_LOC_352/A OR2X1_LOC_214/A AND2X1_LOC_721/Y OR2X1_LOC_624/Y AND2X1_LOC_640/Y AND2X1_LOC_563/A AND2X1_LOC_784/Y AND2X1_LOC_211/B AND2X1_LOC_347/B AND2X1_LOC_850/A AND2X1_LOC_203/Y AND2X1_LOC_208/Y AND2X1_LOC_352/B OR2X1_LOC_725/A OR2X1_LOC_726/A AND2X1_LOC_565/Y AND2X1_LOC_523/Y AND2X1_LOC_61/Y AND2X1_LOC_624/B 
+ AND2X1_LOC_500/Y AND2X1_LOC_401/Y AND2X1_LOC_840/A AND2X1_LOC_500/B AND2X1_LOC_486/Y AND2X1_LOC_649/B AND2X1_LOC_84/Y OR2X1_LOC_365/B OR2X1_LOC_453/Y OR2X1_LOC_475/Y OR2X1_LOC_737/A OR2X1_LOC_140/B OR2X1_LOC_137/Y OR2X1_LOC_739/B OR2X1_LOC_850/B OR2X1_LOC_190/Y OR2X1_LOC_794/A OR2X1_LOC_653/Y OR2X1_LOC_605/Y OR2X1_LOC_561/A OR2X1_LOC_193/Y OR2X1_LOC_140/Y OR2X1_LOC_770/Y OR2X1_LOC_468/A OR2X1_LOC_347/A OR2X1_LOC_842/A OR2X1_LOC_61/Y OR2X1_LOC_84/Y AND2X1_LOC_141/B AND2X1_LOC_231/Y AND2X1_LOC_561/B AND2X1_LOC_792/B AND2X1_LOC_710/Y AND2X1_LOC_647/B AND2X1_LOC_468/B AND2X1_LOC_717/B AND2X1_LOC_702/Y AND2X1_LOC_204/Y AND2X1_LOC_705/Y AND2X1_LOC_645/A AND2X1_LOC_347/Y AND2X1_LOC_572/A AND2X1_LOC_209/Y AND2X1_LOC_726/Y AND2X1_LOC_797/B AND2X1_LOC_554/Y OR2X1_LOC_440/A OR2X1_LOC_551/B OR2X1_LOC_735/B OR2X1_LOC_675/Y OR2X1_LOC_124/A 
+ OR2X1_LOC_835/Y OR2X1_LOC_182/B OR2X1_LOC_175/Y OR2X1_LOC_203/Y OR2X1_LOC_174/Y OR2X1_LOC_641/Y OR2X1_LOC_786/Y OR2X1_LOC_469/B OR2X1_LOC_170/A OR2X1_LOC_192/A OR2X1_LOC_562/B OR2X1_LOC_722/B OR2X1_LOC_703/Y OR2X1_LOC_390/B OR2X1_LOC_201/Y OR2X1_LOC_337/A OR2X1_LOC_624/A OR2X1_LOC_501/A OR2X1_LOC_643/Y AND2X1_LOC_651/B OR2X1_LOC_802/A OR2X1_LOC_798/Y AND2X1_LOC_798/Y AND2X1_LOC_802/B OR2X1_LOC_539/Y AND2X1_LOC_539/Y AND2X1_LOC_810/A OR2X1_LOC_774/Y OR2X1_LOC_510/Y AND2X1_LOC_574/A OR2X1_LOC_35/Y AND2X1_LOC_35/Y AND2X1_LOC_465/A AND2X1_LOC_573/A OR2X1_LOC_465/B OR2X1_LOC_404/Y OR2X1_LOC_799/A AND2X1_LOC_361/A AND2X1_LOC_483/Y AND2X1_LOC_436/Y OR2X1_LOC_631/B OR2X1_LOC_436/Y OR2X1_LOC_319/Y AND2X1_LOC_593/Y OR2X1_LOC_267/Y AND2X1_LOC_798/A 

* NETLIST 
XOR2X1_LOC_338 OR2X1_LOC_338/a_8_216# OR2X1_LOC_338/a_36_216# OR2X1_LOC_351/B VSS VDD OR2X1_LOC_338/A OR2X1_LOC_338/B OR2X1_LOC

XOR2X1_LOC_839 OR2X1_LOC_839/a_8_216# OR2X1_LOC_839/a_36_216# OR2X1_LOC_852/A VSS VDD OR2X1_LOC_836/Y OR2X1_LOC_835/Y OR2X1_LOC

XOR2X1_LOC_243 OR2X1_LOC_243/a_8_216# OR2X1_LOC_243/a_36_216# OR2X1_LOC_244/A VSS VDD OR2X1_LOC_243/A OR2X1_LOC_243/B OR2X1_LOC

XOR2X1_LOC_472 OR2X1_LOC_472/a_8_216# OR2X1_LOC_472/a_36_216# OR2X1_LOC_476/B VSS VDD OR2X1_LOC_472/A OR2X1_LOC_472/B OR2X1_LOC

XAND2X1_LOC_810 AND2X1_LOC_810/a_36_24# AND2X1_LOC_810/Y AND2X1_LOC_810/a_8_24# VSS VDD AND2X1_LOC_810/A AND2X1_LOC_810/B AND2X1_LOC

XAND2X1_LOC_476 AND2X1_LOC_476/a_36_24# AND2X1_LOC_476/Y AND2X1_LOC_476/a_8_24# VSS VDD AND2X1_LOC_476/A AND2X1_LOC_473/Y AND2X1_LOC

XAND2X1_LOC_362 AND2X1_LOC_362/a_36_24# AND2X1_LOC_366/A AND2X1_LOC_362/a_8_24# VSS VDD AND2X1_LOC_806/A AND2X1_LOC_362/B AND2X1_LOC

XOR2X1_LOC_656 OR2X1_LOC_656/a_8_216# OR2X1_LOC_656/a_36_216# OR2X1_LOC_656/Y VSS VDD OR2X1_LOC_647/Y OR2X1_LOC_656/B OR2X1_LOC

XOR2X1_LOC_216 OR2X1_LOC_216/a_8_216# OR2X1_LOC_216/a_36_216# OR2X1_LOC_216/Y VSS VDD OR2X1_LOC_216/A OR2X1_LOC_656/B OR2X1_LOC

XAND2X1_LOC_856 AND2X1_LOC_856/a_36_24# AND2X1_LOC_863/A AND2X1_LOC_856/a_8_24# VSS VDD AND2X1_LOC_856/A AND2X1_LOC_856/B AND2X1_LOC

XAND2X1_LOC_730 AND2X1_LOC_730/a_36_24# AND2X1_LOC_739/B AND2X1_LOC_730/a_8_24# VSS VDD AND2X1_LOC_728/Y AND2X1_LOC_729/Y AND2X1_LOC

XAND2X1_LOC_550 AND2X1_LOC_550/a_36_24# AND2X1_LOC_565/B AND2X1_LOC_550/a_8_24# VSS VDD AND2X1_LOC_550/A AND2X1_LOC_547/Y AND2X1_LOC

XAND2X1_LOC_715 AND2X1_LOC_715/a_36_24# AND2X1_LOC_715/Y AND2X1_LOC_715/a_8_24# VSS VDD AND2X1_LOC_715/A AND2X1_LOC_702/Y AND2X1_LOC

XAND2X1_LOC_339 AND2X1_LOC_339/a_36_24# AND2X1_LOC_339/Y AND2X1_LOC_339/a_8_24# VSS VDD AND2X1_LOC_61/Y AND2X1_LOC_339/B AND2X1_LOC

XAND2X1_LOC_841 AND2X1_LOC_841/a_36_24# AND2X1_LOC_851/B AND2X1_LOC_841/a_8_24# VSS VDD AND2X1_LOC_831/Y AND2X1_LOC_841/B AND2X1_LOC

XAND2X1_LOC_783 AND2X1_LOC_783/a_36_24# AND2X1_LOC_796/A AND2X1_LOC_783/a_8_24# VSS VDD AND2X1_LOC_779/Y AND2X1_LOC_783/B AND2X1_LOC

XAND2X1_LOC_471 AND2X1_LOC_471/a_36_24# AND2X1_LOC_471/Y AND2X1_LOC_471/a_8_24# VSS VDD AND2X1_LOC_464/Y AND2X1_LOC_465/Y AND2X1_LOC

XAND2X1_LOC_559 AND2X1_LOC_559/a_36_24# AND2X1_LOC_560/B AND2X1_LOC_559/a_8_24# VSS VDD OR2X1_LOC_517/Y AND2X1_LOC_520/Y AND2X1_LOC

XAND2X1_LOC_642 AND2X1_LOC_642/a_36_24# AND2X1_LOC_642/Y AND2X1_LOC_642/a_8_24# VSS VDD OR2X1_LOC_416/Y AND2X1_LOC_520/Y AND2X1_LOC

XAND2X1_LOC_771 AND2X1_LOC_771/a_36_24# AND2X1_LOC_774/A AND2X1_LOC_771/a_8_24# VSS VDD AND2X1_LOC_769/Y AND2X1_LOC_771/B AND2X1_LOC

XAND2X1_LOC_199 AND2X1_LOC_199/a_36_24# AND2X1_LOC_207/A AND2X1_LOC_199/a_8_24# VSS VDD AND2X1_LOC_199/A AND2X1_LOC_196/Y AND2X1_LOC

XAND2X1_LOC_840 AND2X1_LOC_840/a_36_24# AND2X1_LOC_851/A AND2X1_LOC_840/a_8_24# VSS VDD AND2X1_LOC_840/A AND2X1_LOC_840/B AND2X1_LOC

XAND2X1_LOC_720 AND2X1_LOC_720/a_36_24# AND2X1_LOC_720/Y AND2X1_LOC_720/a_8_24# VSS VDD OR2X1_LOC_667/Y OR2X1_LOC_669/Y AND2X1_LOC

XAND2X1_LOC_349 AND2X1_LOC_349/a_36_24# AND2X1_LOC_359/B AND2X1_LOC_349/a_8_24# VSS VDD AND2X1_LOC_342/Y AND2X1_LOC_349/B AND2X1_LOC

XOR2X1_LOC_288 OR2X1_LOC_288/a_8_216# OR2X1_LOC_288/a_36_216# OR2X1_LOC_362/B VSS VDD OR2X1_LOC_288/A OR2X1_LOC_286/Y OR2X1_LOC

XOR2X1_LOC_850 OR2X1_LOC_850/a_8_216# OR2X1_LOC_850/a_36_216# OR2X1_LOC_858/B VSS VDD OR2X1_LOC_850/A OR2X1_LOC_850/B OR2X1_LOC

XOR2X1_LOC_632 OR2X1_LOC_632/a_8_216# OR2X1_LOC_632/a_36_216# OR2X1_LOC_632/Y VSS VDD OR2X1_LOC_632/A OR2X1_LOC_630/Y OR2X1_LOC

XAND2X1_LOC_288 AND2X1_LOC_288/a_36_24# AND2X1_LOC_806/A AND2X1_LOC_288/a_8_24# VSS VDD AND2X1_LOC_286/Y AND2X1_LOC_287/Y AND2X1_LOC

XAND2X1_LOC_772 AND2X1_LOC_772/a_36_24# AND2X1_LOC_772/Y AND2X1_LOC_772/a_8_24# VSS VDD AND2X1_LOC_489/Y AND2X1_LOC_772/B AND2X1_LOC

XAND2X1_LOC_338 AND2X1_LOC_338/a_36_24# AND2X1_LOC_338/Y AND2X1_LOC_338/a_8_24# VSS VDD AND2X1_LOC_338/A AND2X1_LOC_334/Y AND2X1_LOC

XAND2X1_LOC_454 AND2X1_LOC_454/a_36_24# AND2X1_LOC_454/Y AND2X1_LOC_454/a_8_24# VSS VDD AND2X1_LOC_454/A AND2X1_LOC_447/Y AND2X1_LOC

XAND2X1_LOC_714 AND2X1_LOC_714/a_36_24# AND2X1_LOC_724/A AND2X1_LOC_714/a_8_24# VSS VDD AND2X1_LOC_703/Y AND2X1_LOC_714/B AND2X1_LOC

XAND2X1_LOC_340 AND2X1_LOC_340/a_36_24# AND2X1_LOC_340/Y AND2X1_LOC_340/a_8_24# VSS VDD OR2X1_LOC_88/Y AND2X1_LOC_227/Y AND2X1_LOC

XAND2X1_LOC_509 AND2X1_LOC_509/a_36_24# AND2X1_LOC_509/Y AND2X1_LOC_509/a_8_24# VSS VDD AND2X1_LOC_227/Y OR2X1_LOC_503/Y AND2X1_LOC

XOR2X1_LOC_303 OR2X1_LOC_303/a_8_216# OR2X1_LOC_303/a_36_216# OR2X1_LOC_566/A VSS VDD OR2X1_LOC_303/A OR2X1_LOC_303/B OR2X1_LOC

XOR2X1_LOC_716 OR2X1_LOC_716/a_8_216# OR2X1_LOC_716/a_36_216# OR2X1_LOC_723/B VSS VDD OR2X1_LOC_303/B OR2X1_LOC_228/Y OR2X1_LOC

XOR2X1_LOC_552 OR2X1_LOC_552/a_8_216# OR2X1_LOC_552/a_36_216# OR2X1_LOC_564/A VSS VDD OR2X1_LOC_552/A OR2X1_LOC_552/B OR2X1_LOC

XOR2X1_LOC_452 OR2X1_LOC_452/a_8_216# OR2X1_LOC_452/a_36_216# OR2X1_LOC_467/A VSS VDD OR2X1_LOC_452/A OR2X1_LOC_450/Y OR2X1_LOC

XAND2X1_LOC_859 AND2X1_LOC_859/a_36_24# AND2X1_LOC_859/Y AND2X1_LOC_859/a_8_24# VSS VDD AND2X1_LOC_848/Y AND2X1_LOC_859/B AND2X1_LOC

XAND2X1_LOC_647 AND2X1_LOC_647/a_36_24# AND2X1_LOC_647/Y AND2X1_LOC_647/a_8_24# VSS VDD OR2X1_LOC_612/Y AND2X1_LOC_647/B AND2X1_LOC

XOR2X1_LOC_202 OR2X1_LOC_202/a_8_216# OR2X1_LOC_202/a_36_216# OR2X1_LOC_206/A VSS VDD AND2X1_LOC_69/Y AND2X1_LOC_67/Y OR2X1_LOC

XOR2X1_LOC_854 OR2X1_LOC_854/a_8_216# OR2X1_LOC_854/a_36_216# OR2X1_LOC_856/B VSS VDD OR2X1_LOC_854/A OR2X1_LOC_354/A OR2X1_LOC

XOR2X1_LOC_567 OR2X1_LOC_567/a_8_216# OR2X1_LOC_567/a_36_216# OR2X1_LOC_568/A VSS VDD OR2X1_LOC_539/Y OR2X1_LOC_854/A OR2X1_LOC

XOR2X1_LOC_199 OR2X1_LOC_199/a_8_216# OR2X1_LOC_199/a_36_216# OR2X1_LOC_207/B VSS VDD OR2X1_LOC_196/Y OR2X1_LOC_199/B OR2X1_LOC

XOR2X1_LOC_139 OR2X1_LOC_139/a_8_216# OR2X1_LOC_139/a_36_216# OR2X1_LOC_141/B VSS VDD OR2X1_LOC_139/A OR2X1_LOC_137/Y OR2X1_LOC

XOR2X1_LOC_852 OR2X1_LOC_852/a_8_216# OR2X1_LOC_852/a_36_216# OR2X1_LOC_857/B VSS VDD OR2X1_LOC_852/A OR2X1_LOC_852/B OR2X1_LOC

XOR2X1_LOC_454 OR2X1_LOC_454/a_8_216# OR2X1_LOC_454/a_36_216# OR2X1_LOC_466/A VSS VDD OR2X1_LOC_447/Y OR2X1_LOC_446/Y OR2X1_LOC

XOR2X1_LOC_508 OR2X1_LOC_508/a_8_216# OR2X1_LOC_508/a_36_216# OR2X1_LOC_508/Y VSS VDD OR2X1_LOC_508/A OR2X1_LOC_506/Y OR2X1_LOC

XOR2X1_LOC_390 OR2X1_LOC_390/a_8_216# OR2X1_LOC_390/a_36_216# OR2X1_LOC_392/B VSS VDD OR2X1_LOC_390/A OR2X1_LOC_390/B OR2X1_LOC

XAND2X1_LOC_149 AND2X1_LOC_149/a_36_24# AND2X1_LOC_797/A AND2X1_LOC_149/a_8_24# VSS VDD AND2X1_LOC_147/Y AND2X1_LOC_148/Y AND2X1_LOC

XAND2X1_LOC_353 AND2X1_LOC_353/a_36_24# AND2X1_LOC_357/B AND2X1_LOC_353/a_8_24# VSS VDD AND2X1_LOC_566/B AND2X1_LOC_727/A AND2X1_LOC

XAND2X1_LOC_727 AND2X1_LOC_727/a_36_24# AND2X1_LOC_727/Y AND2X1_LOC_727/a_8_24# VSS VDD AND2X1_LOC_727/A AND2X1_LOC_727/B AND2X1_LOC

XAND2X1_LOC_712 AND2X1_LOC_712/a_36_24# AND2X1_LOC_712/Y AND2X1_LOC_712/a_8_24# VSS VDD AND2X1_LOC_707/Y AND2X1_LOC_712/B AND2X1_LOC

XAND2X1_LOC_651 AND2X1_LOC_651/a_36_24# AND2X1_LOC_654/B AND2X1_LOC_651/a_8_24# VSS VDD AND2X1_LOC_638/Y AND2X1_LOC_651/B AND2X1_LOC

XAND2X1_LOC_463 AND2X1_LOC_463/a_36_24# AND2X1_LOC_472/B AND2X1_LOC_463/a_8_24# VSS VDD AND2X1_LOC_459/Y AND2X1_LOC_463/B AND2X1_LOC

XAND2X1_LOC_326 AND2X1_LOC_326/a_36_24# AND2X1_LOC_354/B AND2X1_LOC_326/a_8_24# VSS VDD AND2X1_LOC_326/A AND2X1_LOC_326/B AND2X1_LOC

XAND2X1_LOC_717 AND2X1_LOC_717/a_36_24# AND2X1_LOC_717/Y AND2X1_LOC_717/a_8_24# VSS VDD AND2X1_LOC_374/Y AND2X1_LOC_717/B AND2X1_LOC

XAND2X1_LOC_170 AND2X1_LOC_170/a_36_24# AND2X1_LOC_170/Y AND2X1_LOC_170/a_8_24# VSS VDD AND2X1_LOC_168/Y AND2X1_LOC_170/B AND2X1_LOC

XAND2X1_LOC_785 AND2X1_LOC_785/a_36_24# AND2X1_LOC_785/Y AND2X1_LOC_785/a_8_24# VSS VDD AND2X1_LOC_785/A AND2X1_LOC_776/Y AND2X1_LOC

XOR2X1_LOC_845 OR2X1_LOC_845/a_8_216# OR2X1_LOC_845/a_36_216# OR2X1_LOC_849/A VSS VDD OR2X1_LOC_845/A OR2X1_LOC_673/Y OR2X1_LOC

XOR2X1_LOC_721 OR2X1_LOC_721/a_8_216# OR2X1_LOC_721/a_36_216# OR2X1_LOC_721/Y VSS VDD OR2X1_LOC_720/Y OR2X1_LOC_673/Y OR2X1_LOC

XAND2X1_LOC_713 AND2X1_LOC_713/a_36_24# AND2X1_LOC_713/Y AND2X1_LOC_713/a_8_24# VSS VDD AND2X1_LOC_705/Y AND2X1_LOC_706/Y AND2X1_LOC

XAND2X1_LOC_711 AND2X1_LOC_711/a_36_24# AND2X1_LOC_711/Y AND2X1_LOC_711/a_8_24# VSS VDD AND2X1_LOC_711/A AND2X1_LOC_710/Y AND2X1_LOC

XAND2X1_LOC_624 AND2X1_LOC_624/a_36_24# AND2X1_LOC_658/A AND2X1_LOC_624/a_8_24# VSS VDD AND2X1_LOC_624/A AND2X1_LOC_624/B AND2X1_LOC

XOR2X1_LOC_640 OR2X1_LOC_640/a_8_216# OR2X1_LOC_640/a_36_216# OR2X1_LOC_640/Y VSS VDD OR2X1_LOC_640/A OR2X1_LOC_633/Y OR2X1_LOC

XOR2X1_LOC_553 OR2X1_LOC_553/a_8_216# OR2X1_LOC_553/a_36_216# OR2X1_LOC_563/B VSS VDD OR2X1_LOC_553/A OR2X1_LOC_553/B OR2X1_LOC

XOR2X1_LOC_784 OR2X1_LOC_784/a_8_216# OR2X1_LOC_784/a_36_216# OR2X1_LOC_784/Y VSS VDD OR2X1_LOC_778/Y OR2X1_LOC_784/B OR2X1_LOC

XOR2X1_LOC_565 OR2X1_LOC_565/a_8_216# OR2X1_LOC_565/a_36_216# OR2X1_LOC_569/A VSS VDD OR2X1_LOC_565/A OR2X1_LOC_549/Y OR2X1_LOC

XOR2X1_LOC_392 OR2X1_LOC_392/a_8_216# OR2X1_LOC_392/a_36_216# OR2X1_LOC_474/B VSS VDD OR2X1_LOC_392/A OR2X1_LOC_392/B OR2X1_LOC

XAND2X1_LOC_390 AND2X1_LOC_390/a_36_24# AND2X1_LOC_392/A AND2X1_LOC_390/a_8_24# VSS VDD AND2X1_LOC_388/Y AND2X1_LOC_390/B AND2X1_LOC

XAND2X1_LOC_644 AND2X1_LOC_644/a_36_24# AND2X1_LOC_644/Y AND2X1_LOC_644/a_8_24# VSS VDD OR2X1_LOC_597/Y OR2X1_LOC_599/Y AND2X1_LOC

XAND2X1_LOC_356 AND2X1_LOC_356/a_36_24# AND2X1_LOC_365/A AND2X1_LOC_356/a_8_24# VSS VDD AND2X1_LOC_354/Y AND2X1_LOC_356/B AND2X1_LOC

XAND2X1_LOC_507 AND2X1_LOC_507/a_36_24# AND2X1_LOC_508/B AND2X1_LOC_507/a_8_24# VSS VDD OR2X1_LOC_504/Y OR2X1_LOC_505/Y AND2X1_LOC

XAND2X1_LOC_781 AND2X1_LOC_781/a_36_24# AND2X1_LOC_781/Y AND2X1_LOC_781/a_8_24# VSS VDD OR2X1_LOC_745/Y OR2X1_LOC_746/Y AND2X1_LOC

XAND2X1_LOC_259 AND2X1_LOC_259/a_36_24# AND2X1_LOC_259/Y AND2X1_LOC_259/a_8_24# VSS VDD OR2X1_LOC_257/Y OR2X1_LOC_258/Y AND2X1_LOC

XAND2X1_LOC_210 AND2X1_LOC_210/a_36_24# AND2X1_LOC_213/B AND2X1_LOC_210/a_8_24# VSS VDD OR2X1_LOC_158/Y OR2X1_LOC_163/Y AND2X1_LOC

XAND2X1_LOC_544 AND2X1_LOC_544/a_36_24# AND2X1_LOC_544/Y AND2X1_LOC_544/a_8_24# VSS VDD OR2X1_LOC_373/Y OR2X1_LOC_438/Y AND2X1_LOC

XAND2X1_LOC_439 AND2X1_LOC_439/a_36_24# AND2X1_LOC_675/A AND2X1_LOC_439/a_8_24# VSS VDD OR2X1_LOC_177/Y OR2X1_LOC_438/Y AND2X1_LOC

XAND2X1_LOC_605 AND2X1_LOC_605/a_36_24# AND2X1_LOC_605/Y AND2X1_LOC_605/a_8_24# VSS VDD OR2X1_LOC_603/Y OR2X1_LOC_604/Y AND2X1_LOC

XAND2X1_LOC_501 AND2X1_LOC_501/a_36_24# AND2X1_LOC_501/Y AND2X1_LOC_501/a_8_24# VSS VDD OR2X1_LOC_498/Y AND2X1_LOC_500/Y AND2X1_LOC

XAND2X1_LOC_675 AND2X1_LOC_675/a_36_24# AND2X1_LOC_675/Y AND2X1_LOC_675/a_8_24# VSS VDD AND2X1_LOC_675/A OR2X1_LOC_674/Y AND2X1_LOC

XAND2X1_LOC_123 AND2X1_LOC_123/a_36_24# AND2X1_LOC_123/Y AND2X1_LOC_123/a_8_24# VSS VDD OR2X1_LOC_117/Y OR2X1_LOC_118/Y AND2X1_LOC

XAND2X1_LOC_835 AND2X1_LOC_835/a_36_24# AND2X1_LOC_839/A AND2X1_LOC_835/a_8_24# VSS VDD OR2X1_LOC_821/Y OR2X1_LOC_822/Y AND2X1_LOC

XAND2X1_LOC_180 AND2X1_LOC_180/a_36_24# AND2X1_LOC_182/A AND2X1_LOC_180/a_8_24# VSS VDD OR2X1_LOC_176/Y OR2X1_LOC_177/Y AND2X1_LOC

XAND2X1_LOC_402 AND2X1_LOC_402/a_36_24# AND2X1_LOC_404/A AND2X1_LOC_402/a_8_24# VSS VDD OR2X1_LOC_397/Y AND2X1_LOC_401/Y AND2X1_LOC

XAND2X1_LOC_194 AND2X1_LOC_194/a_36_24# AND2X1_LOC_194/Y AND2X1_LOC_194/a_8_24# VSS VDD OR2X1_LOC_16/Y OR2X1_LOC_39/Y AND2X1_LOC

XAND2X1_LOC_773 AND2X1_LOC_773/a_36_24# AND2X1_LOC_773/Y AND2X1_LOC_773/a_8_24# VSS VDD OR2X1_LOC_767/Y AND2X1_LOC_772/Y AND2X1_LOC

XAND2X1_LOC_719 AND2X1_LOC_719/a_36_24# AND2X1_LOC_719/Y AND2X1_LOC_719/a_8_24# VSS VDD OR2X1_LOC_665/Y OR2X1_LOC_666/Y AND2X1_LOC

XAND2X1_LOC_174 AND2X1_LOC_174/a_36_24# AND2X1_LOC_175/B AND2X1_LOC_174/a_8_24# VSS VDD OR2X1_LOC_171/Y OR2X1_LOC_172/Y AND2X1_LOC

XAND2X1_LOC_641 AND2X1_LOC_641/a_36_24# AND2X1_LOC_641/Y AND2X1_LOC_641/a_8_24# VSS VDD AND2X1_LOC_231/Y OR2X1_LOC_265/Y AND2X1_LOC

XAND2X1_LOC_545 AND2X1_LOC_545/a_36_24# AND2X1_LOC_551/B AND2X1_LOC_545/a_8_24# VSS VDD OR2X1_LOC_441/Y OR2X1_LOC_524/Y AND2X1_LOC

XAND2X1_LOC_443 AND2X1_LOC_443/a_36_24# AND2X1_LOC_443/Y AND2X1_LOC_443/a_8_24# VSS VDD OR2X1_LOC_91/Y OR2X1_LOC_441/Y AND2X1_LOC

XAND2X1_LOC_169 AND2X1_LOC_169/a_36_24# AND2X1_LOC_170/B AND2X1_LOC_169/a_8_24# VSS VDD OR2X1_LOC_166/Y OR2X1_LOC_167/Y AND2X1_LOC

XAND2X1_LOC_191 AND2X1_LOC_191/a_36_24# AND2X1_LOC_191/Y AND2X1_LOC_191/a_8_24# VSS VDD OR2X1_LOC_187/Y AND2X1_LOC_191/B AND2X1_LOC

XAND2X1_LOC_452 AND2X1_LOC_452/a_36_24# AND2X1_LOC_452/Y AND2X1_LOC_452/a_8_24# VSS VDD AND2X1_LOC_450/Y AND2X1_LOC_451/Y AND2X1_LOC

XOR2X1_LOC_242 OR2X1_LOC_242/a_8_216# OR2X1_LOC_242/a_36_216# OR2X1_LOC_244/B VSS VDD OR2X1_LOC_241/Y OR2X1_LOC_506/B OR2X1_LOC

XOR2X1_LOC_343 OR2X1_LOC_343/a_8_216# OR2X1_LOC_343/a_36_216# OR2X1_LOC_349/A VSS VDD OR2X1_LOC_843/B OR2X1_LOC_343/B OR2X1_LOC

XOR2X1_LOC_728 OR2X1_LOC_728/a_8_216# OR2X1_LOC_728/a_36_216# OR2X1_LOC_730/B VSS VDD OR2X1_LOC_728/A OR2X1_LOC_728/B OR2X1_LOC

XOR2X1_LOC_148 OR2X1_LOC_148/a_8_216# OR2X1_LOC_148/a_36_216# OR2X1_LOC_148/Y VSS VDD OR2X1_LOC_148/A OR2X1_LOC_148/B OR2X1_LOC

XOR2X1_LOC_467 OR2X1_LOC_467/a_8_216# OR2X1_LOC_467/a_36_216# OR2X1_LOC_470/A VSS VDD OR2X1_LOC_467/A OR2X1_LOC_467/B OR2X1_LOC

XOR2X1_LOC_210 OR2X1_LOC_210/a_8_216# OR2X1_LOC_210/a_36_216# OR2X1_LOC_213/A VSS VDD OR2X1_LOC_467/B OR2X1_LOC_210/B OR2X1_LOC

XOR2X1_LOC_443 OR2X1_LOC_443/a_8_216# OR2X1_LOC_443/a_36_216# OR2X1_LOC_443/Y VSS VDD OR2X1_LOC_545/B OR2X1_LOC_97/A OR2X1_LOC

XOR2X1_LOC_775 OR2X1_LOC_775/a_8_216# OR2X1_LOC_775/a_36_216# OR2X1_LOC_785/B VSS VDD OR2X1_LOC_112/B OR2X1_LOC_97/A OR2X1_LOC

XOR2X1_LOC_493 OR2X1_LOC_493/a_8_216# OR2X1_LOC_493/a_36_216# OR2X1_LOC_493/Y VSS VDD OR2X1_LOC_493/A OR2X1_LOC_493/B OR2X1_LOC

XOR2X1_LOC_559 OR2X1_LOC_559/a_8_216# OR2X1_LOC_559/a_36_216# OR2X1_LOC_560/A VSS VDD OR2X1_LOC_520/Y OR2X1_LOC_559/B OR2X1_LOC

XOR2X1_LOC_76 OR2X1_LOC_76/a_8_216# OR2X1_LOC_76/a_36_216# OR2X1_LOC_76/Y VSS VDD OR2X1_LOC_76/A OR2X1_LOC_76/B OR2X1_LOC

XOR2X1_LOC_449 OR2X1_LOC_449/a_8_216# OR2X1_LOC_449/a_36_216# OR2X1_LOC_453/A VSS VDD OR2X1_LOC_449/A OR2X1_LOC_449/B OR2X1_LOC

XOR2X1_LOC_347 OR2X1_LOC_347/a_8_216# OR2X1_LOC_347/a_36_216# OR2X1_LOC_347/Y VSS VDD OR2X1_LOC_347/A OR2X1_LOC_347/B OR2X1_LOC

XOR2X1_LOC_486 OR2X1_LOC_486/a_8_216# OR2X1_LOC_486/a_36_216# OR2X1_LOC_486/Y VSS VDD OR2X1_LOC_705/B OR2X1_LOC_486/B OR2X1_LOC

XOR2X1_LOC_705 OR2X1_LOC_705/a_8_216# OR2X1_LOC_705/a_36_216# OR2X1_LOC_705/Y VSS VDD OR2X1_LOC_546/A OR2X1_LOC_705/B OR2X1_LOC

XOR2X1_LOC_124 OR2X1_LOC_124/a_8_216# OR2X1_LOC_124/a_36_216# OR2X1_LOC_124/Y VSS VDD OR2X1_LOC_124/A OR2X1_LOC_124/B OR2X1_LOC

XOR2X1_LOC_403 OR2X1_LOC_403/a_8_216# OR2X1_LOC_403/a_36_216# OR2X1_LOC_404/A VSS VDD OR2X1_LOC_403/A OR2X1_LOC_403/B OR2X1_LOC

XOR2X1_LOC_791 OR2X1_LOC_791/a_8_216# OR2X1_LOC_791/a_36_216# OR2X1_LOC_792/A VSS VDD OR2X1_LOC_791/A OR2X1_LOC_791/B OR2X1_LOC

XOR2X1_LOC_554 OR2X1_LOC_554/a_8_216# OR2X1_LOC_554/a_36_216# OR2X1_LOC_563/A VSS VDD OR2X1_LOC_140/B OR2X1_LOC_115/B OR2X1_LOC

XOR2X1_LOC_768 OR2X1_LOC_768/a_8_216# OR2X1_LOC_768/a_36_216# OR2X1_LOC_772/A VSS VDD OR2X1_LOC_768/A OR2X1_LOC_113/B OR2X1_LOC

XOR2X1_LOC_209 OR2X1_LOC_209/a_8_216# OR2X1_LOC_209/a_36_216# OR2X1_LOC_213/B VSS VDD OR2X1_LOC_209/A OR2X1_LOC_797/B OR2X1_LOC

XOR2X1_LOC_726 OR2X1_LOC_726/a_8_216# OR2X1_LOC_726/a_36_216# OR2X1_LOC_731/B VSS VDD OR2X1_LOC_726/A OR2X1_LOC_209/A OR2X1_LOC

XOR2X1_LOC_400 OR2X1_LOC_400/a_8_216# OR2X1_LOC_400/a_36_216# OR2X1_LOC_403/A VSS VDD OR2X1_LOC_400/A OR2X1_LOC_400/B OR2X1_LOC

XOR2X1_LOC_793 OR2X1_LOC_793/a_8_216# OR2X1_LOC_793/a_36_216# OR2X1_LOC_805/A VSS VDD OR2X1_LOC_793/A OR2X1_LOC_793/B OR2X1_LOC

XOR2X1_LOC_639 OR2X1_LOC_639/a_8_216# OR2X1_LOC_639/a_36_216# OR2X1_LOC_651/A VSS VDD OR2X1_LOC_639/A OR2X1_LOC_639/B OR2X1_LOC

XOR2X1_LOC_771 OR2X1_LOC_771/a_8_216# OR2X1_LOC_771/a_36_216# OR2X1_LOC_774/B VSS VDD OR2X1_LOC_770/Y OR2X1_LOC_771/B OR2X1_LOC

XAND2X1_LOC_467 AND2X1_LOC_467/a_36_24# AND2X1_LOC_470/B AND2X1_LOC_467/a_8_24# VSS VDD OR2X1_LOC_163/Y AND2X1_LOC_452/Y AND2X1_LOC

XAND2X1_LOC_546 AND2X1_LOC_546/a_36_24# AND2X1_LOC_550/A AND2X1_LOC_546/a_8_24# VSS VDD OR2X1_LOC_525/Y OR2X1_LOC_526/Y AND2X1_LOC

XAND2X1_LOC_241 AND2X1_LOC_241/a_36_24# AND2X1_LOC_242/B AND2X1_LOC_241/a_8_24# VSS VDD OR2X1_LOC_237/Y OR2X1_LOC_238/Y AND2X1_LOC

XAND2X1_LOC_228 AND2X1_LOC_228/a_36_24# AND2X1_LOC_228/Y AND2X1_LOC_228/a_8_24# VSS VDD OR2X1_LOC_7/Y OR2X1_LOC_52/Y AND2X1_LOC

XAND2X1_LOC_343 AND2X1_LOC_343/a_36_24# AND2X1_LOC_349/B AND2X1_LOC_343/a_8_24# VSS VDD OR2X1_LOC_250/Y OR2X1_LOC_251/Y AND2X1_LOC

XAND2X1_LOC_728 AND2X1_LOC_728/a_36_24# AND2X1_LOC_728/Y AND2X1_LOC_728/a_8_24# VSS VDD OR2X1_LOC_679/Y OR2X1_LOC_680/Y AND2X1_LOC

XAND2X1_LOC_148 AND2X1_LOC_148/a_36_24# AND2X1_LOC_148/Y AND2X1_LOC_148/a_8_24# VSS VDD OR2X1_LOC_145/Y OR2X1_LOC_146/Y AND2X1_LOC

XAND2X1_LOC_788 AND2X1_LOC_788/a_36_24# AND2X1_LOC_794/B AND2X1_LOC_788/a_8_24# VSS VDD OR2X1_LOC_533/Y AND2X1_LOC_645/A AND2X1_LOC

XAND2X1_LOC_653 AND2X1_LOC_653/a_36_24# AND2X1_LOC_661/A AND2X1_LOC_653/a_8_24# VSS VDD OR2X1_LOC_594/Y AND2X1_LOC_653/B AND2X1_LOC

XAND2X1_LOC_734 AND2X1_LOC_734/a_36_24# AND2X1_LOC_734/Y AND2X1_LOC_734/a_8_24# VSS VDD OR2X1_LOC_406/Y AND2X1_LOC_721/Y AND2X1_LOC

XAND2X1_LOC_475 AND2X1_LOC_475/a_36_24# AND2X1_LOC_475/Y AND2X1_LOC_475/a_8_24# VSS VDD OR2X1_LOC_406/Y AND2X1_LOC_474/Y AND2X1_LOC

XAND2X1_LOC_192 AND2X1_LOC_192/a_36_24# AND2X1_LOC_192/Y AND2X1_LOC_192/a_8_24# VSS VDD OR2X1_LOC_189/Y AND2X1_LOC_191/Y AND2X1_LOC

XAND2X1_LOC_830 AND2X1_LOC_830/a_36_24# AND2X1_LOC_842/B AND2X1_LOC_830/a_8_24# VSS VDD OR2X1_LOC_108/Y OR2X1_LOC_142/Y AND2X1_LOC

XAND2X1_LOC_324 AND2X1_LOC_324/a_36_24# AND2X1_LOC_326/A AND2X1_LOC_324/a_8_24# VSS VDD OR2X1_LOC_320/Y OR2X1_LOC_321/Y AND2X1_LOC

XAND2X1_LOC_718 AND2X1_LOC_718/a_36_24# AND2X1_LOC_722/A AND2X1_LOC_718/a_8_24# VSS VDD OR2X1_LOC_591/Y AND2X1_LOC_605/Y AND2X1_LOC

XAND2X1_LOC_703 AND2X1_LOC_703/a_36_24# AND2X1_LOC_703/Y AND2X1_LOC_703/a_8_24# VSS VDD OR2X1_LOC_167/Y OR2X1_LOC_312/Y AND2X1_LOC

XAND2X1_LOC_388 AND2X1_LOC_388/a_36_24# AND2X1_LOC_388/Y AND2X1_LOC_388/a_8_24# VSS VDD OR2X1_LOC_167/Y OR2X1_LOC_176/Y AND2X1_LOC

XOR2X1_LOC_259 OR2X1_LOC_259/a_8_216# OR2X1_LOC_259/a_36_216# OR2X1_LOC_555/B VSS VDD OR2X1_LOC_259/A OR2X1_LOC_259/B OR2X1_LOC

XOR2X1_LOC_642 OR2X1_LOC_642/a_8_216# OR2X1_LOC_642/a_36_216# OR2X1_LOC_649/B VSS VDD OR2X1_LOC_520/Y OR2X1_LOC_462/B OR2X1_LOC

XOR2X1_LOC_540 OR2X1_LOC_540/a_8_216# OR2X1_LOC_540/a_36_216# OR2X1_LOC_553/B VSS VDD OR2X1_LOC_190/B OR2X1_LOC_181/B OR2X1_LOC

XOR2X1_LOC_181 OR2X1_LOC_181/a_8_216# OR2X1_LOC_181/a_36_216# OR2X1_LOC_181/Y VSS VDD OR2X1_LOC_181/A OR2X1_LOC_181/B OR2X1_LOC

XOR2X1_LOC_781 OR2X1_LOC_781/a_8_216# OR2X1_LOC_781/a_36_216# OR2X1_LOC_781/Y VSS VDD OR2X1_LOC_781/A OR2X1_LOC_781/B OR2X1_LOC

XOR2X1_LOC_833 OR2X1_LOC_833/a_8_216# OR2X1_LOC_833/a_36_216# OR2X1_LOC_833/Y VSS VDD OR2X1_LOC_499/B OR2X1_LOC_833/B OR2X1_LOC

XOR2X1_LOC_499 OR2X1_LOC_499/a_8_216# OR2X1_LOC_499/a_36_216# OR2X1_LOC_500/A VSS VDD OR2X1_LOC_778/A OR2X1_LOC_499/B OR2X1_LOC

XOR2X1_LOC_194 OR2X1_LOC_194/a_8_216# OR2X1_LOC_194/a_36_216# OR2X1_LOC_194/Y VSS VDD AND2X1_LOC_39/Y OR2X1_LOC_194/B OR2X1_LOC

XOR2X1_LOC_324 OR2X1_LOC_324/a_8_216# OR2X1_LOC_324/a_36_216# OR2X1_LOC_326/B VSS VDD OR2X1_LOC_324/A OR2X1_LOC_324/B OR2X1_LOC

XOR2X1_LOC_644 OR2X1_LOC_644/a_8_216# OR2X1_LOC_644/a_36_216# OR2X1_LOC_648/B VSS VDD OR2X1_LOC_644/A OR2X1_LOC_644/B OR2X1_LOC

XOR2X1_LOC_646 OR2X1_LOC_646/a_8_216# OR2X1_LOC_646/a_36_216# OR2X1_LOC_647/A VSS VDD OR2X1_LOC_646/A OR2X1_LOC_646/B OR2X1_LOC

XOR2X1_LOC_719 OR2X1_LOC_719/a_8_216# OR2X1_LOC_719/a_36_216# OR2X1_LOC_719/Y VSS VDD OR2X1_LOC_719/A OR2X1_LOC_719/B OR2X1_LOC

XOR2X1_LOC_204 OR2X1_LOC_204/a_8_216# OR2X1_LOC_204/a_36_216# OR2X1_LOC_204/Y VSS VDD OR2X1_LOC_84/Y AND2X1_LOC_79/Y OR2X1_LOC

XOR2X1_LOC_810 OR2X1_LOC_810/a_8_216# OR2X1_LOC_810/a_36_216# OR2X1_LOC_812/B VSS VDD OR2X1_LOC_810/A OR2X1_LOC_774/Y OR2X1_LOC

XOR2X1_LOC_574 OR2X1_LOC_574/a_8_216# OR2X1_LOC_574/a_36_216# OR2X1_LOC_575/A VSS VDD OR2X1_LOC_574/A OR2X1_LOC_510/Y OR2X1_LOC

XOR2X1_LOC_362 OR2X1_LOC_362/a_8_216# OR2X1_LOC_362/a_36_216# OR2X1_LOC_366/B VSS VDD OR2X1_LOC_362/A OR2X1_LOC_362/B OR2X1_LOC

XOR2X1_LOC_476 OR2X1_LOC_476/a_8_216# OR2X1_LOC_476/a_36_216# OR2X1_LOC_476/Y VSS VDD OR2X1_LOC_473/Y OR2X1_LOC_476/B OR2X1_LOC

XAND2X1_LOC_656 AND2X1_LOC_656/a_36_24# AND2X1_LOC_656/Y AND2X1_LOC_656/a_8_24# VSS VDD AND2X1_LOC_216/A AND2X1_LOC_647/Y AND2X1_LOC

XAND2X1_LOC_216 AND2X1_LOC_216/a_36_24# AND2X1_LOC_216/Y AND2X1_LOC_216/a_8_24# VSS VDD AND2X1_LOC_216/A AND2X1_LOC_116/Y AND2X1_LOC

XAND2X1_LOC_345 AND2X1_LOC_345/a_36_24# AND2X1_LOC_345/Y AND2X1_LOC_345/a_8_24# VSS VDD AND2X1_LOC_259/Y OR2X1_LOC_261/Y AND2X1_LOC

XAND2X1_LOC_444 AND2X1_LOC_444/a_36_24# AND2X1_LOC_727/B AND2X1_LOC_444/a_8_24# VSS VDD OR2X1_LOC_442/Y AND2X1_LOC_443/Y AND2X1_LOC

XAND2X1_LOC_128 AND2X1_LOC_128/a_36_24# AND2X1_LOC_554/B AND2X1_LOC_128/a_8_24# VSS VDD OR2X1_LOC_125/Y OR2X1_LOC_127/Y AND2X1_LOC

XOR2X1_LOC_561 OR2X1_LOC_561/a_8_216# OR2X1_LOC_561/a_36_216# OR2X1_LOC_561/Y VSS VDD OR2X1_LOC_561/A OR2X1_LOC_561/B OR2X1_LOC

XOR2X1_LOC_33 OR2X1_LOC_33/a_8_216# OR2X1_LOC_33/a_36_216# OR2X1_LOC_35/B VSS VDD OR2X1_LOC_33/A OR2X1_LOC_33/B OR2X1_LOC

XAND2X1_LOC_540 AND2X1_LOC_540/a_36_24# AND2X1_LOC_553/A AND2X1_LOC_540/a_8_24# VSS VDD OR2X1_LOC_178/Y OR2X1_LOC_183/Y AND2X1_LOC

XAND2X1_LOC_190 AND2X1_LOC_190/a_36_24# AND2X1_LOC_191/B AND2X1_LOC_190/a_8_24# VSS VDD OR2X1_LOC_183/Y OR2X1_LOC_184/Y AND2X1_LOC

XAND2X1_LOC_636 AND2X1_LOC_636/a_36_24# AND2X1_LOC_639/B AND2X1_LOC_636/a_8_24# VSS VDD OR2X1_LOC_583/Y OR2X1_LOC_584/Y AND2X1_LOC

XAND2X1_LOC_193 AND2X1_LOC_193/a_36_24# AND2X1_LOC_193/Y AND2X1_LOC_193/a_8_24# VSS VDD OR2X1_LOC_7/Y OR2X1_LOC_13/Y AND2X1_LOC

XAND2X1_LOC_449 AND2X1_LOC_449/a_36_24# AND2X1_LOC_449/Y AND2X1_LOC_449/a_8_24# VSS VDD OR2X1_LOC_423/Y OR2X1_LOC_424/Y AND2X1_LOC

XOR2X1_LOC_348 OR2X1_LOC_348/a_8_216# OR2X1_LOC_348/a_36_216# OR2X1_LOC_348/Y VSS VDD OR2X1_LOC_345/Y OR2X1_LOC_348/B OR2X1_LOC

XAND2X1_LOC_793 AND2X1_LOC_793/a_36_24# AND2X1_LOC_793/Y AND2X1_LOC_793/a_8_24# VSS VDD AND2X1_LOC_789/Y AND2X1_LOC_793/B AND2X1_LOC

XOR2X1_LOC_445 OR2X1_LOC_445/a_8_216# OR2X1_LOC_445/a_36_216# OR2X1_LOC_455/A VSS VDD OR2X1_LOC_318/B OR2X1_LOC_241/B OR2X1_LOC

XAND2X1_LOC_679 AND2X1_LOC_679/a_36_24# OR2X1_LOC_728/B AND2X1_LOC_679/a_8_24# VSS VDD OR2X1_LOC_676/Y OR2X1_LOC_678/Y AND2X1_LOC

XOR2X1_LOC_545 OR2X1_LOC_545/a_8_216# OR2X1_LOC_545/a_36_216# OR2X1_LOC_551/A VSS VDD OR2X1_LOC_545/A OR2X1_LOC_545/B OR2X1_LOC

XOR2X1_LOC_228 OR2X1_LOC_228/a_8_216# OR2X1_LOC_228/a_36_216# OR2X1_LOC_228/Y VSS VDD AND2X1_LOC_52/Y AND2X1_LOC_7/Y OR2X1_LOC

XOR2X1_LOC_782 OR2X1_LOC_782/a_8_216# OR2X1_LOC_782/a_36_216# OR2X1_LOC_797/A VSS VDD OR2X1_LOC_781/Y OR2X1_LOC_782/B OR2X1_LOC

XOR2X1_LOC_523 OR2X1_LOC_523/a_8_216# OR2X1_LOC_523/a_36_216# OR2X1_LOC_523/Y VSS VDD OR2X1_LOC_523/A OR2X1_LOC_523/B OR2X1_LOC

XOR2X1_LOC_636 OR2X1_LOC_636/a_8_216# OR2X1_LOC_636/a_36_216# OR2X1_LOC_639/A VSS VDD OR2X1_LOC_636/A OR2X1_LOC_636/B OR2X1_LOC

XOR2X1_LOC_542 OR2X1_LOC_542/a_8_216# OR2X1_LOC_542/a_36_216# OR2X1_LOC_552/B VSS VDD OR2X1_LOC_703/A OR2X1_LOC_542/B OR2X1_LOC

XOR2X1_LOC_792 OR2X1_LOC_792/a_8_216# OR2X1_LOC_792/a_36_216# OR2X1_LOC_792/Y VSS VDD OR2X1_LOC_792/A OR2X1_LOC_792/B OR2X1_LOC

XOR2X1_LOC_710 OR2X1_LOC_710/a_8_216# OR2X1_LOC_710/a_36_216# OR2X1_LOC_711/A VSS VDD OR2X1_LOC_710/A OR2X1_LOC_710/B OR2X1_LOC

XAND2X1_LOC_839 AND2X1_LOC_839/a_36_24# AND2X1_LOC_852/B AND2X1_LOC_839/a_8_24# VSS VDD AND2X1_LOC_839/A AND2X1_LOC_839/B AND2X1_LOC

XAND2X1_LOC_243 AND2X1_LOC_243/a_36_24# AND2X1_LOC_243/Y AND2X1_LOC_243/a_8_24# VSS VDD OR2X1_LOC_235/Y AND2X1_LOC_240/Y AND2X1_LOC

XAND2X1_LOC_472 AND2X1_LOC_472/a_36_24# AND2X1_LOC_476/A AND2X1_LOC_472/a_8_24# VSS VDD AND2X1_LOC_462/Y AND2X1_LOC_472/B AND2X1_LOC

XOR2X1_LOC_730 OR2X1_LOC_730/a_8_216# OR2X1_LOC_730/a_36_216# OR2X1_LOC_739/A VSS VDD OR2X1_LOC_730/A OR2X1_LOC_730/B OR2X1_LOC

XOR2X1_LOC_856 OR2X1_LOC_856/a_8_216# OR2X1_LOC_856/a_36_216# OR2X1_LOC_863/B VSS VDD OR2X1_LOC_856/A OR2X1_LOC_856/B OR2X1_LOC

XOR2X1_LOC_550 OR2X1_LOC_550/a_8_216# OR2X1_LOC_550/a_36_216# OR2X1_LOC_565/A VSS VDD OR2X1_LOC_550/A OR2X1_LOC_550/B OR2X1_LOC

XOR2X1_LOC_339 OR2X1_LOC_339/a_8_216# OR2X1_LOC_339/a_36_216# OR2X1_LOC_339/Y VSS VDD OR2X1_LOC_339/A OR2X1_LOC_61/Y OR2X1_LOC

XOR2X1_LOC_715 OR2X1_LOC_715/a_8_216# OR2X1_LOC_715/a_36_216# OR2X1_LOC_724/A VSS VDD OR2X1_LOC_715/A OR2X1_LOC_715/B OR2X1_LOC

XAND2X1_LOC_574 AND2X1_LOC_574/a_36_24# AND2X1_LOC_574/Y AND2X1_LOC_574/a_8_24# VSS VDD AND2X1_LOC_574/A OR2X1_LOC_516/Y AND2X1_LOC

XOR2X1_LOC_787 OR2X1_LOC_787/a_8_216# OR2X1_LOC_787/a_36_216# OR2X1_LOC_787/Y VSS VDD OR2X1_LOC_486/Y OR2X1_LOC_787/B OR2X1_LOC

XOR2X1_LOC_772 OR2X1_LOC_772/a_8_216# OR2X1_LOC_772/a_36_216# OR2X1_LOC_772/Y VSS VDD OR2X1_LOC_772/A OR2X1_LOC_772/B OR2X1_LOC

XOR2X1_LOC_714 OR2X1_LOC_714/a_8_216# OR2X1_LOC_714/a_36_216# OR2X1_LOC_714/Y VSS VDD OR2X1_LOC_714/A OR2X1_LOC_703/Y OR2X1_LOC

XOR2X1_LOC_509 OR2X1_LOC_509/a_8_216# OR2X1_LOC_509/a_36_216# OR2X1_LOC_510/A VSS VDD OR2X1_LOC_509/A OR2X1_LOC_227/Y OR2X1_LOC

XOR2X1_LOC_340 OR2X1_LOC_340/a_8_216# OR2X1_LOC_340/a_36_216# OR2X1_LOC_340/Y VSS VDD OR2X1_LOC_227/Y AND2X1_LOC_88/Y OR2X1_LOC

XOR2X1_LOC_679 OR2X1_LOC_679/a_8_216# OR2X1_LOC_679/a_36_216# OR2X1_LOC_679/Y VSS VDD OR2X1_LOC_679/A OR2X1_LOC_679/B OR2X1_LOC

XAND2X1_LOC_768 AND2X1_LOC_768/a_36_24# AND2X1_LOC_772/B AND2X1_LOC_768/a_8_24# VSS VDD OR2X1_LOC_103/Y OR2X1_LOC_134/Y AND2X1_LOC

XAND2X1_LOC_137 AND2X1_LOC_137/a_36_24# AND2X1_LOC_139/A AND2X1_LOC_137/a_8_24# VSS VDD OR2X1_LOC_132/Y OR2X1_LOC_134/Y AND2X1_LOC

XOR2X1_LOC_34 OR2X1_LOC_34/a_8_216# OR2X1_LOC_34/a_36_216# OR2X1_LOC_35/A VSS VDD OR2X1_LOC_34/A OR2X1_LOC_34/B OR2X1_LOC

XAND2X1_LOC_792 AND2X1_LOC_792/a_36_24# AND2X1_LOC_792/Y AND2X1_LOC_792/a_8_24# VSS VDD OR2X1_LOC_759/Y AND2X1_LOC_792/B AND2X1_LOC

XAND2X1_LOC_392 AND2X1_LOC_392/a_36_24# AND2X1_LOC_474/A AND2X1_LOC_392/a_8_24# VSS VDD AND2X1_LOC_392/A AND2X1_LOC_391/Y AND2X1_LOC

XAND2X1_LOC_400 AND2X1_LOC_400/a_36_24# AND2X1_LOC_403/B AND2X1_LOC_400/a_8_24# VSS VDD OR2X1_LOC_393/Y OR2X1_LOC_394/Y AND2X1_LOC

XOR2X1_LOC_859 OR2X1_LOC_859/a_8_216# OR2X1_LOC_859/a_36_216# OR2X1_LOC_862/A VSS VDD OR2X1_LOC_859/A OR2X1_LOC_859/B OR2X1_LOC

XOR2X1_LOC_507 OR2X1_LOC_507/a_8_216# OR2X1_LOC_507/a_36_216# OR2X1_LOC_508/A VSS VDD OR2X1_LOC_507/A OR2X1_LOC_507/B OR2X1_LOC

XOR2X1_LOC_546 OR2X1_LOC_546/a_8_216# OR2X1_LOC_546/a_36_216# OR2X1_LOC_550/B VSS VDD OR2X1_LOC_546/A OR2X1_LOC_546/B OR2X1_LOC

XOR2X1_LOC_720 OR2X1_LOC_720/a_8_216# OR2X1_LOC_720/a_36_216# OR2X1_LOC_720/Y VSS VDD OR2X1_LOC_720/A OR2X1_LOC_720/B OR2X1_LOC

XOR2X1_LOC_602 OR2X1_LOC_602/a_8_216# OR2X1_LOC_602/a_36_216# OR2X1_LOC_602/Y VSS VDD OR2X1_LOC_602/A OR2X1_LOC_602/B OR2X1_LOC

XAND2X1_LOC_850 AND2X1_LOC_850/a_36_24# AND2X1_LOC_850/Y AND2X1_LOC_850/a_8_24# VSS VDD AND2X1_LOC_850/A AND2X1_LOC_843/Y AND2X1_LOC

XOR2X1_LOC_349 OR2X1_LOC_349/a_8_216# OR2X1_LOC_349/a_36_216# OR2X1_LOC_359/A VSS VDD OR2X1_LOC_349/A OR2X1_LOC_349/B OR2X1_LOC

XAND2X1_LOC_242 AND2X1_LOC_242/a_36_24# AND2X1_LOC_244/A AND2X1_LOC_242/a_8_24# VSS VDD OR2X1_LOC_239/Y AND2X1_LOC_242/B AND2X1_LOC

XAND2X1_LOC_770 AND2X1_LOC_770/a_36_24# AND2X1_LOC_771/B AND2X1_LOC_770/a_8_24# VSS VDD OR2X1_LOC_765/Y OR2X1_LOC_766/Y AND2X1_LOC

XAND2X1_LOC_775 AND2X1_LOC_775/a_36_24# AND2X1_LOC_785/A AND2X1_LOC_775/a_8_24# VSS VDD OR2X1_LOC_91/Y OR2X1_LOC_109/Y AND2X1_LOC

XOR2X1_LOC_647 OR2X1_LOC_647/a_8_216# OR2X1_LOC_647/a_36_216# OR2X1_LOC_647/Y VSS VDD OR2X1_LOC_647/A OR2X1_LOC_647/B OR2X1_LOC

XAND2X1_LOC_542 AND2X1_LOC_542/a_36_24# AND2X1_LOC_552/A AND2X1_LOC_542/a_8_24# VSS VDD OR2X1_LOC_280/Y OR2X1_LOC_312/Y AND2X1_LOC

XAND2X1_LOC_336 AND2X1_LOC_336/a_36_24# AND2X1_LOC_337/B AND2X1_LOC_336/a_8_24# VSS VDD OR2X1_LOC_311/Y OR2X1_LOC_312/Y AND2X1_LOC

XAND2X1_LOC_202 AND2X1_LOC_202/a_36_24# AND2X1_LOC_202/Y AND2X1_LOC_202/a_8_24# VSS VDD OR2X1_LOC_67/Y OR2X1_LOC_69/Y AND2X1_LOC

XAND2X1_LOC_620 AND2X1_LOC_620/a_36_24# AND2X1_LOC_620/Y AND2X1_LOC_620/a_8_24# VSS VDD OR2X1_LOC_528/Y OR2X1_LOC_613/Y AND2X1_LOC

XAND2X1_LOC_181 AND2X1_LOC_181/a_36_24# AND2X1_LOC_181/Y AND2X1_LOC_181/a_8_24# VSS VDD OR2X1_LOC_178/Y OR2X1_LOC_179/Y AND2X1_LOC

XAND2X1_LOC_139 AND2X1_LOC_139/a_36_24# AND2X1_LOC_141/A AND2X1_LOC_139/a_8_24# VSS VDD AND2X1_LOC_139/A AND2X1_LOC_139/B AND2X1_LOC

XAND2X1_LOC_852 AND2X1_LOC_852/a_36_24# AND2X1_LOC_852/Y AND2X1_LOC_852/a_8_24# VSS VDD AND2X1_LOC_838/Y AND2X1_LOC_852/B AND2X1_LOC

XAND2X1_LOC_508 AND2X1_LOC_508/a_36_24# AND2X1_LOC_510/A AND2X1_LOC_508/a_8_24# VSS VDD AND2X1_LOC_508/A AND2X1_LOC_508/B AND2X1_LOC

XAND2X1_LOC_567 AND2X1_LOC_567/a_36_24# AND2X1_LOC_568/B AND2X1_LOC_567/a_8_24# VSS VDD AND2X1_LOC_535/Y AND2X1_LOC_539/Y AND2X1_LOC

XAND2X1_LOC_854 AND2X1_LOC_854/a_36_24# AND2X1_LOC_856/A AND2X1_LOC_854/a_8_24# VSS VDD AND2X1_LOC_354/B AND2X1_LOC_535/Y AND2X1_LOC

XAND2X1_LOC_561 AND2X1_LOC_561/a_36_24# AND2X1_LOC_571/B AND2X1_LOC_561/a_8_24# VSS VDD AND2X1_LOC_557/Y AND2X1_LOC_561/B AND2X1_LOC

XOR2X1_LOC_241 OR2X1_LOC_241/a_8_216# OR2X1_LOC_241/a_36_216# OR2X1_LOC_241/Y VSS VDD OR2X1_LOC_776/A OR2X1_LOC_241/B OR2X1_LOC

XOR2X1_LOC_702 OR2X1_LOC_702/a_8_216# OR2X1_LOC_702/a_36_216# OR2X1_LOC_715/A VSS VDD OR2X1_LOC_702/A OR2X1_LOC_196/B OR2X1_LOC

XOR2X1_LOC_401 OR2X1_LOC_401/a_8_216# OR2X1_LOC_401/a_36_216# OR2X1_LOC_401/Y VSS VDD OR2X1_LOC_401/A OR2X1_LOC_401/B OR2X1_LOC

XOR2X1_LOC_345 OR2X1_LOC_345/a_8_216# OR2X1_LOC_345/a_36_216# OR2X1_LOC_345/Y VSS VDD OR2X1_LOC_345/A OR2X1_LOC_555/B OR2X1_LOC

XAND2X1_LOC_348 AND2X1_LOC_348/a_36_24# AND2X1_LOC_348/Y AND2X1_LOC_348/a_8_24# VSS VDD AND2X1_LOC_348/A AND2X1_LOC_345/Y AND2X1_LOC

XOR2X1_LOC_231 OR2X1_LOC_231/a_8_216# OR2X1_LOC_231/a_36_216# OR2X1_LOC_641/B VSS VDD OR2X1_LOC_231/A OR2X1_LOC_231/B OR2X1_LOC

XOR2X1_LOC_620 OR2X1_LOC_620/a_8_216# OR2X1_LOC_620/a_36_216# OR2X1_LOC_620/Y VSS VDD OR2X1_LOC_620/A OR2X1_LOC_620/B OR2X1_LOC

XAND2X1_LOC_453 AND2X1_LOC_453/a_36_24# AND2X1_LOC_453/Y AND2X1_LOC_453/a_8_24# VSS VDD AND2X1_LOC_448/Y AND2X1_LOC_449/Y AND2X1_LOC

XAND2X1_LOC_632 AND2X1_LOC_632/a_36_24# AND2X1_LOC_658/B AND2X1_LOC_632/a_8_24# VSS VDD AND2X1_LOC_632/A AND2X1_LOC_631/Y AND2X1_LOC

XOR2X1_LOC_783 OR2X1_LOC_783/a_8_216# OR2X1_LOC_783/a_36_216# OR2X1_LOC_796/B VSS VDD OR2X1_LOC_783/A OR2X1_LOC_779/Y OR2X1_LOC

XOR2X1_LOC_840 OR2X1_LOC_840/a_8_216# OR2X1_LOC_840/a_36_216# OR2X1_LOC_851/B VSS VDD OR2X1_LOC_840/A OR2X1_LOC_833/Y OR2X1_LOC

XAND2X1_LOC_555 AND2X1_LOC_555/a_36_24# AND2X1_LOC_555/Y AND2X1_LOC_555/a_8_24# VSS VDD AND2X1_LOC_259/Y OR2X1_LOC_481/Y AND2X1_LOC

XOR2X1_LOC_651 OR2X1_LOC_651/a_8_216# OR2X1_LOC_651/a_36_216# OR2X1_LOC_654/A VSS VDD OR2X1_LOC_651/A OR2X1_LOC_651/B OR2X1_LOC

XOR2X1_LOC_463 OR2X1_LOC_463/a_8_216# OR2X1_LOC_463/a_36_216# OR2X1_LOC_472/A VSS VDD OR2X1_LOC_460/Y OR2X1_LOC_463/B OR2X1_LOC

XOR2X1_LOC_717 OR2X1_LOC_717/a_8_216# OR2X1_LOC_717/a_36_216# OR2X1_LOC_723/A VSS VDD OR2X1_LOC_493/Y OR2X1_LOC_374/Y OR2X1_LOC

XOR2X1_LOC_326 OR2X1_LOC_326/a_8_216# OR2X1_LOC_326/a_36_216# OR2X1_LOC_354/A VSS VDD OR2X1_LOC_325/Y OR2X1_LOC_326/B OR2X1_LOC

XOR2X1_LOC_785 OR2X1_LOC_785/a_8_216# OR2X1_LOC_785/a_36_216# OR2X1_LOC_795/B VSS VDD OR2X1_LOC_776/Y OR2X1_LOC_785/B OR2X1_LOC

XOR2X1_LOC_170 OR2X1_LOC_170/a_8_216# OR2X1_LOC_170/a_36_216# OR2X1_LOC_170/Y VSS VDD OR2X1_LOC_170/A OR2X1_LOC_168/Y OR2X1_LOC

XOR2X1_LOC_149 OR2X1_LOC_149/a_8_216# OR2X1_LOC_149/a_36_216# OR2X1_LOC_797/B VSS VDD OR2X1_LOC_148/Y OR2X1_LOC_149/B OR2X1_LOC

XOR2X1_LOC_353 OR2X1_LOC_353/a_8_216# OR2X1_LOC_353/a_36_216# OR2X1_LOC_357/A VSS VDD OR2X1_LOC_308/Y OR2X1_LOC_566/A OR2X1_LOC

XOR2X1_LOC_727 OR2X1_LOC_727/a_8_216# OR2X1_LOC_727/a_36_216# OR2X1_LOC_731/A VSS VDD OR2X1_LOC_469/B OR2X1_LOC_308/Y OR2X1_LOC

XOR2X1_LOC_712 OR2X1_LOC_712/a_8_216# OR2X1_LOC_712/a_36_216# OR2X1_LOC_725/B VSS VDD OR2X1_LOC_708/Y OR2X1_LOC_712/B OR2X1_LOC

XOR2X1_LOC_841 OR2X1_LOC_841/a_8_216# OR2X1_LOC_841/a_36_216# OR2X1_LOC_851/A VSS VDD OR2X1_LOC_841/A OR2X1_LOC_841/B OR2X1_LOC

XAND2X1_LOC_552 AND2X1_LOC_552/a_36_24# AND2X1_LOC_564/B AND2X1_LOC_552/a_8_24# VSS VDD AND2X1_LOC_552/A AND2X1_LOC_543/Y AND2X1_LOC

XAND2X1_LOC_787 AND2X1_LOC_787/a_36_24# AND2X1_LOC_794/A AND2X1_LOC_787/a_8_24# VSS VDD AND2X1_LOC_787/A AND2X1_LOC_486/Y AND2X1_LOC

XAND2X1_LOC_303 AND2X1_LOC_303/a_36_24# AND2X1_LOC_566/B AND2X1_LOC_303/a_8_24# VSS VDD AND2X1_LOC_303/A AND2X1_LOC_303/B AND2X1_LOC

XAND2X1_LOC_716 AND2X1_LOC_716/a_36_24# AND2X1_LOC_716/Y AND2X1_LOC_716/a_8_24# VSS VDD AND2X1_LOC_228/Y AND2X1_LOC_303/A AND2X1_LOC

XOR2X1_LOC_471 OR2X1_LOC_471/a_8_216# OR2X1_LOC_471/a_36_216# OR2X1_LOC_471/Y VSS VDD OR2X1_LOC_465/Y OR2X1_LOC_471/B OR2X1_LOC

XAND2X1_LOC_201 AND2X1_LOC_201/a_36_24# AND2X1_LOC_201/Y AND2X1_LOC_201/a_8_24# VSS VDD AND2X1_LOC_61/Y OR2X1_LOC_65/Y AND2X1_LOC

XAND2X1_LOC_786 AND2X1_LOC_786/a_36_24# AND2X1_LOC_786/Y AND2X1_LOC_786/a_8_24# VSS VDD AND2X1_LOC_84/Y OR2X1_LOC_262/Y AND2X1_LOC

XOR2X1_LOC_337 OR2X1_LOC_337/a_8_216# OR2X1_LOC_337/a_36_216# OR2X1_LOC_352/A VSS VDD OR2X1_LOC_337/A OR2X1_LOC_335/Y OR2X1_LOC

XOR2X1_LOC_208 OR2X1_LOC_208/a_8_216# OR2X1_LOC_208/a_36_216# OR2X1_LOC_214/A VSS VDD OR2X1_LOC_208/A OR2X1_LOC_35/Y OR2X1_LOC

XAND2X1_LOC_721 AND2X1_LOC_721/a_36_24# AND2X1_LOC_721/Y AND2X1_LOC_721/a_8_24# VSS VDD AND2X1_LOC_721/A AND2X1_LOC_720/Y AND2X1_LOC

XAND2X1_LOC_845 AND2X1_LOC_845/a_36_24# AND2X1_LOC_845/Y AND2X1_LOC_845/a_8_24# VSS VDD AND2X1_LOC_721/A OR2X1_LOC_813/Y AND2X1_LOC

XOR2X1_LOC_624 OR2X1_LOC_624/a_8_216# OR2X1_LOC_624/a_36_216# OR2X1_LOC_624/Y VSS VDD OR2X1_LOC_624/A OR2X1_LOC_624/B OR2X1_LOC

XAND2X1_LOC_640 AND2X1_LOC_640/a_36_24# AND2X1_LOC_640/Y AND2X1_LOC_640/a_8_24# VSS VDD AND2X1_LOC_633/Y AND2X1_LOC_634/Y AND2X1_LOC

XAND2X1_LOC_553 AND2X1_LOC_553/a_36_24# AND2X1_LOC_563/A AND2X1_LOC_553/a_8_24# VSS VDD AND2X1_LOC_553/A AND2X1_LOC_541/Y AND2X1_LOC

XAND2X1_LOC_784 AND2X1_LOC_784/a_36_24# AND2X1_LOC_784/Y AND2X1_LOC_784/a_8_24# VSS VDD AND2X1_LOC_784/A AND2X1_LOC_778/Y AND2X1_LOC

XAND2X1_LOC_175 AND2X1_LOC_175/a_36_24# AND2X1_LOC_211/B AND2X1_LOC_175/a_8_24# VSS VDD OR2X1_LOC_173/Y AND2X1_LOC_175/B AND2X1_LOC

XAND2X1_LOC_346 AND2X1_LOC_346/a_36_24# AND2X1_LOC_347/B AND2X1_LOC_346/a_8_24# VSS VDD OR2X1_LOC_292/Y OR2X1_LOC_295/Y AND2X1_LOC

XAND2X1_LOC_842 AND2X1_LOC_842/a_36_24# AND2X1_LOC_850/A AND2X1_LOC_842/a_8_24# VSS VDD OR2X1_LOC_184/Y AND2X1_LOC_842/B AND2X1_LOC

XAND2X1_LOC_456 AND2X1_LOC_456/a_36_24# AND2X1_LOC_456/Y AND2X1_LOC_456/a_8_24# VSS VDD OR2X1_LOC_184/Y AND2X1_LOC_456/B AND2X1_LOC

XAND2X1_LOC_203 AND2X1_LOC_203/a_36_24# AND2X1_LOC_203/Y AND2X1_LOC_203/a_8_24# VSS VDD OR2X1_LOC_72/Y AND2X1_LOC_76/Y AND2X1_LOC

XAND2X1_LOC_208 AND2X1_LOC_208/a_36_24# AND2X1_LOC_208/Y AND2X1_LOC_208/a_8_24# VSS VDD AND2X1_LOC_35/Y AND2X1_LOC_208/B AND2X1_LOC

XAND2X1_LOC_337 AND2X1_LOC_337/a_36_24# AND2X1_LOC_352/B AND2X1_LOC_337/a_8_24# VSS VDD AND2X1_LOC_335/Y AND2X1_LOC_337/B AND2X1_LOC

XOR2X1_LOC_713 OR2X1_LOC_713/a_8_216# OR2X1_LOC_713/a_36_216# OR2X1_LOC_725/A VSS VDD OR2X1_LOC_713/A OR2X1_LOC_705/Y OR2X1_LOC

XOR2X1_LOC_711 OR2X1_LOC_711/a_8_216# OR2X1_LOC_711/a_36_216# OR2X1_LOC_726/A VSS VDD OR2X1_LOC_711/A OR2X1_LOC_711/B OR2X1_LOC

XAND2X1_LOC_565 AND2X1_LOC_565/a_36_24# AND2X1_LOC_565/Y AND2X1_LOC_565/a_8_24# VSS VDD AND2X1_LOC_549/Y AND2X1_LOC_565/B AND2X1_LOC

XAND2X1_LOC_523 AND2X1_LOC_523/a_36_24# AND2X1_LOC_523/Y AND2X1_LOC_523/a_8_24# VSS VDD OR2X1_LOC_521/Y OR2X1_LOC_522/Y AND2X1_LOC

XAND2X1_LOC_61 AND2X1_LOC_61/a_36_24# AND2X1_LOC_61/Y AND2X1_LOC_61/a_8_24# VSS VDD OR2X1_LOC_58/Y OR2X1_LOC_60/Y AND2X1_LOC

XAND2X1_LOC_33 AND2X1_LOC_33/a_36_24# AND2X1_LOC_33/Y AND2X1_LOC_33/a_8_24# VSS VDD OR2X1_LOC_20/Y OR2X1_LOC_24/Y AND2X1_LOC

XAND2X1_LOC_623 AND2X1_LOC_623/a_36_24# AND2X1_LOC_624/B AND2X1_LOC_623/a_8_24# VSS VDD OR2X1_LOC_615/Y AND2X1_LOC_620/Y AND2X1_LOC

XAND2X1_LOC_500 AND2X1_LOC_500/a_36_24# AND2X1_LOC_500/Y AND2X1_LOC_500/a_8_24# VSS VDD OR2X1_LOC_497/Y AND2X1_LOC_500/B AND2X1_LOC

XAND2X1_LOC_844 AND2X1_LOC_844/a_36_24# AND2X1_LOC_849/A AND2X1_LOC_844/a_8_24# VSS VDD OR2X1_LOC_497/Y AND2X1_LOC_523/Y AND2X1_LOC

XAND2X1_LOC_401 AND2X1_LOC_401/a_36_24# AND2X1_LOC_401/Y AND2X1_LOC_401/a_8_24# VSS VDD OR2X1_LOC_395/Y OR2X1_LOC_396/Y AND2X1_LOC

XAND2X1_LOC_833 AND2X1_LOC_833/a_36_24# AND2X1_LOC_840/A AND2X1_LOC_833/a_8_24# VSS VDD OR2X1_LOC_482/Y OR2X1_LOC_495/Y AND2X1_LOC

XAND2X1_LOC_499 AND2X1_LOC_499/a_36_24# AND2X1_LOC_500/B AND2X1_LOC_499/a_8_24# VSS VDD OR2X1_LOC_495/Y OR2X1_LOC_496/Y AND2X1_LOC

XAND2X1_LOC_486 AND2X1_LOC_486/a_36_24# AND2X1_LOC_486/Y AND2X1_LOC_486/a_8_24# VSS VDD OR2X1_LOC_484/Y OR2X1_LOC_485/Y AND2X1_LOC

XAND2X1_LOC_34 AND2X1_LOC_34/a_36_24# AND2X1_LOC_34/Y AND2X1_LOC_34/a_8_24# VSS VDD OR2X1_LOC_27/Y OR2X1_LOC_32/Y AND2X1_LOC

XAND2X1_LOC_643 AND2X1_LOC_643/a_36_24# AND2X1_LOC_649/B AND2X1_LOC_643/a_8_24# VSS VDD AND2X1_LOC_537/Y OR2X1_LOC_595/Y AND2X1_LOC

XAND2X1_LOC_445 AND2X1_LOC_445/a_36_24# AND2X1_LOC_455/B AND2X1_LOC_445/a_8_24# VSS VDD OR2X1_LOC_237/Y OR2X1_LOC_315/Y AND2X1_LOC

XAND2X1_LOC_84 AND2X1_LOC_84/a_36_24# AND2X1_LOC_84/Y AND2X1_LOC_84/a_8_24# VSS VDD OR2X1_LOC_81/Y OR2X1_LOC_83/Y AND2X1_LOC

XOR2X1_LOC_356 OR2X1_LOC_356/a_8_216# OR2X1_LOC_356/a_36_216# OR2X1_LOC_365/B VSS VDD OR2X1_LOC_356/A OR2X1_LOC_356/B OR2X1_LOC

XOR2X1_LOC_453 OR2X1_LOC_453/a_8_216# OR2X1_LOC_453/a_36_216# OR2X1_LOC_453/Y VSS VDD OR2X1_LOC_453/A OR2X1_LOC_448/Y OR2X1_LOC

XOR2X1_LOC_475 OR2X1_LOC_475/a_8_216# OR2X1_LOC_475/a_36_216# OR2X1_LOC_475/Y VSS VDD OR2X1_LOC_474/Y OR2X1_LOC_475/B OR2X1_LOC

XOR2X1_LOC_734 OR2X1_LOC_734/a_8_216# OR2X1_LOC_734/a_36_216# OR2X1_LOC_737/A VSS VDD OR2X1_LOC_721/Y OR2X1_LOC_475/B OR2X1_LOC

XOR2X1_LOC_128 OR2X1_LOC_128/a_8_216# OR2X1_LOC_128/a_36_216# OR2X1_LOC_140/B VSS VDD OR2X1_LOC_128/A OR2X1_LOC_128/B OR2X1_LOC

XOR2X1_LOC_137 OR2X1_LOC_137/a_8_216# OR2X1_LOC_137/a_36_216# OR2X1_LOC_137/Y VSS VDD OR2X1_LOC_768/A OR2X1_LOC_137/B OR2X1_LOC

XOR2X1_LOC_192 OR2X1_LOC_192/a_8_216# OR2X1_LOC_192/a_36_216# OR2X1_LOC_739/B VSS VDD OR2X1_LOC_192/A OR2X1_LOC_192/B OR2X1_LOC

XOR2X1_LOC_842 OR2X1_LOC_842/a_8_216# OR2X1_LOC_842/a_36_216# OR2X1_LOC_850/B VSS VDD OR2X1_LOC_842/A OR2X1_LOC_190/A OR2X1_LOC

XOR2X1_LOC_456 OR2X1_LOC_456/a_8_216# OR2X1_LOC_456/a_36_216# OR2X1_LOC_456/Y VSS VDD OR2X1_LOC_456/A OR2X1_LOC_190/A OR2X1_LOC

XOR2X1_LOC_190 OR2X1_LOC_190/a_8_216# OR2X1_LOC_190/a_36_216# OR2X1_LOC_190/Y VSS VDD OR2X1_LOC_190/A OR2X1_LOC_190/B OR2X1_LOC

XOR2X1_LOC_788 OR2X1_LOC_788/a_8_216# OR2X1_LOC_788/a_36_216# OR2X1_LOC_794/A VSS VDD OR2X1_LOC_602/Y OR2X1_LOC_788/B OR2X1_LOC

XOR2X1_LOC_653 OR2X1_LOC_653/a_8_216# OR2X1_LOC_653/a_36_216# OR2X1_LOC_653/Y VSS VDD OR2X1_LOC_653/A OR2X1_LOC_653/B OR2X1_LOC

XOR2X1_LOC_605 OR2X1_LOC_605/a_8_216# OR2X1_LOC_605/a_36_216# OR2X1_LOC_605/Y VSS VDD OR2X1_LOC_605/A OR2X1_LOC_605/B OR2X1_LOC

XOR2X1_LOC_558 OR2X1_LOC_558/a_8_216# OR2X1_LOC_558/a_36_216# OR2X1_LOC_561/A VSS VDD OR2X1_LOC_558/A OR2X1_LOC_493/Y OR2X1_LOC

XOR2X1_LOC_193 OR2X1_LOC_193/a_8_216# OR2X1_LOC_193/a_36_216# OR2X1_LOC_193/Y VSS VDD OR2X1_LOC_193/A AND2X1_LOC_7/Y OR2X1_LOC

XOR2X1_LOC_140 OR2X1_LOC_140/a_8_216# OR2X1_LOC_140/a_36_216# OR2X1_LOC_140/Y VSS VDD OR2X1_LOC_140/A OR2X1_LOC_140/B OR2X1_LOC

XOR2X1_LOC_770 OR2X1_LOC_770/a_8_216# OR2X1_LOC_770/a_36_216# OR2X1_LOC_770/Y VSS VDD OR2X1_LOC_770/A OR2X1_LOC_770/B OR2X1_LOC

XOR2X1_LOC_440 OR2X1_LOC_440/a_8_216# OR2X1_LOC_440/a_36_216# OR2X1_LOC_468/A VSS VDD OR2X1_LOC_440/A OR2X1_LOC_440/B OR2X1_LOC

XOR2X1_LOC_346 OR2X1_LOC_346/a_8_216# OR2X1_LOC_346/a_36_216# OR2X1_LOC_347/A VSS VDD OR2X1_LOC_346/A OR2X1_LOC_346/B OR2X1_LOC

XOR2X1_LOC_830 OR2X1_LOC_830/a_8_216# OR2X1_LOC_830/a_36_216# OR2X1_LOC_842/A VSS VDD OR2X1_LOC_147/B OR2X1_LOC_114/B OR2X1_LOC

XOR2X1_LOC_61 OR2X1_LOC_61/a_8_216# OR2X1_LOC_61/a_36_216# OR2X1_LOC_61/Y VSS VDD OR2X1_LOC_61/A OR2X1_LOC_61/B OR2X1_LOC

XOR2X1_LOC_84 OR2X1_LOC_84/a_8_216# OR2X1_LOC_84/a_36_216# OR2X1_LOC_84/Y VSS VDD OR2X1_LOC_84/A OR2X1_LOC_84/B OR2X1_LOC

XAND2X1_LOC_140 AND2X1_LOC_140/a_36_24# AND2X1_LOC_141/B AND2X1_LOC_140/a_8_24# VSS VDD AND2X1_LOC_554/B OR2X1_LOC_131/Y AND2X1_LOC

XAND2X1_LOC_231 AND2X1_LOC_231/a_36_24# AND2X1_LOC_231/Y AND2X1_LOC_231/a_8_24# VSS VDD OR2X1_LOC_229/Y OR2X1_LOC_230/Y AND2X1_LOC

XAND2X1_LOC_558 AND2X1_LOC_558/a_36_24# AND2X1_LOC_561/B AND2X1_LOC_558/a_8_24# VSS VDD AND2X1_LOC_717/B OR2X1_LOC_494/Y AND2X1_LOC

XAND2X1_LOC_791 AND2X1_LOC_791/a_36_24# AND2X1_LOC_792/B AND2X1_LOC_791/a_8_24# VSS VDD OR2X1_LOC_755/Y OR2X1_LOC_757/Y AND2X1_LOC

XAND2X1_LOC_710 AND2X1_LOC_710/a_36_24# AND2X1_LOC_710/Y AND2X1_LOC_710/a_8_24# VSS VDD OR2X1_LOC_700/Y OR2X1_LOC_701/Y AND2X1_LOC

XAND2X1_LOC_76 AND2X1_LOC_76/a_36_24# AND2X1_LOC_76/Y AND2X1_LOC_76/a_8_24# VSS VDD OR2X1_LOC_74/Y OR2X1_LOC_75/Y AND2X1_LOC

XAND2X1_LOC_646 AND2X1_LOC_646/a_36_24# AND2X1_LOC_647/B AND2X1_LOC_646/a_8_24# VSS VDD OR2X1_LOC_607/Y OR2X1_LOC_609/Y AND2X1_LOC

XAND2X1_LOC_440 AND2X1_LOC_440/a_36_24# AND2X1_LOC_468/B AND2X1_LOC_440/a_8_24# VSS VDD OR2X1_LOC_437/Y AND2X1_LOC_675/A AND2X1_LOC

XAND2X1_LOC_493 AND2X1_LOC_493/a_36_24# AND2X1_LOC_717/B AND2X1_LOC_493/a_8_24# VSS VDD OR2X1_LOC_491/Y OR2X1_LOC_492/Y AND2X1_LOC

XAND2X1_LOC_702 AND2X1_LOC_702/a_36_24# AND2X1_LOC_702/Y AND2X1_LOC_702/a_8_24# VSS VDD OR2X1_LOC_45/Y OR2X1_LOC_135/Y AND2X1_LOC

XAND2X1_LOC_204 AND2X1_LOC_204/a_36_24# AND2X1_LOC_204/Y AND2X1_LOC_204/a_8_24# VSS VDD OR2X1_LOC_79/Y AND2X1_LOC_84/Y AND2X1_LOC

XAND2X1_LOC_705 AND2X1_LOC_705/a_36_24# AND2X1_LOC_705/Y AND2X1_LOC_705/a_8_24# VSS VDD OR2X1_LOC_485/Y OR2X1_LOC_526/Y AND2X1_LOC

XAND2X1_LOC_602 AND2X1_LOC_602/a_36_24# AND2X1_LOC_645/A AND2X1_LOC_602/a_8_24# VSS VDD OR2X1_LOC_600/Y OR2X1_LOC_601/Y AND2X1_LOC

XAND2X1_LOC_403 AND2X1_LOC_403/a_36_24# AND2X1_LOC_404/B AND2X1_LOC_403/a_8_24# VSS VDD OR2X1_LOC_399/Y AND2X1_LOC_403/B AND2X1_LOC

XAND2X1_LOC_347 AND2X1_LOC_347/a_36_24# AND2X1_LOC_347/Y AND2X1_LOC_347/a_8_24# VSS VDD OR2X1_LOC_297/Y AND2X1_LOC_347/B AND2X1_LOC

XAND2X1_LOC_124 AND2X1_LOC_124/a_36_24# AND2X1_LOC_572/A AND2X1_LOC_124/a_8_24# VSS VDD OR2X1_LOC_122/Y AND2X1_LOC_123/Y AND2X1_LOC

XAND2X1_LOC_209 AND2X1_LOC_209/a_36_24# AND2X1_LOC_209/Y AND2X1_LOC_209/a_8_24# VSS VDD AND2X1_LOC_797/A OR2X1_LOC_152/Y AND2X1_LOC

XAND2X1_LOC_726 AND2X1_LOC_726/a_36_24# AND2X1_LOC_726/Y AND2X1_LOC_726/a_8_24# VSS VDD OR2X1_LOC_152/Y AND2X1_LOC_711/Y AND2X1_LOC

XAND2X1_LOC_782 AND2X1_LOC_782/a_36_24# AND2X1_LOC_797/B AND2X1_LOC_782/a_8_24# VSS VDD OR2X1_LOC_747/Y AND2X1_LOC_781/Y AND2X1_LOC

XAND2X1_LOC_554 AND2X1_LOC_554/a_36_24# AND2X1_LOC_554/Y AND2X1_LOC_554/a_8_24# VSS VDD OR2X1_LOC_106/Y AND2X1_LOC_554/B AND2X1_LOC

XOR2X1_LOC_439 OR2X1_LOC_439/a_8_216# OR2X1_LOC_439/a_36_216# OR2X1_LOC_440/A VSS VDD OR2X1_LOC_544/A OR2X1_LOC_439/B OR2X1_LOC

XOR2X1_LOC_544 OR2X1_LOC_544/a_8_216# OR2X1_LOC_544/a_36_216# OR2X1_LOC_551/B VSS VDD OR2X1_LOC_544/A OR2X1_LOC_544/B OR2X1_LOC

XOR2X1_LOC_501 OR2X1_LOC_501/a_8_216# OR2X1_LOC_501/a_36_216# OR2X1_LOC_735/B VSS VDD OR2X1_LOC_501/A OR2X1_LOC_501/B OR2X1_LOC

XOR2X1_LOC_675 OR2X1_LOC_675/a_8_216# OR2X1_LOC_675/a_36_216# OR2X1_LOC_675/Y VSS VDD OR2X1_LOC_675/A OR2X1_LOC_440/A OR2X1_LOC

XOR2X1_LOC_123 OR2X1_LOC_123/a_8_216# OR2X1_LOC_123/a_36_216# OR2X1_LOC_124/A VSS VDD OR2X1_LOC_633/B OR2X1_LOC_123/B OR2X1_LOC

XOR2X1_LOC_835 OR2X1_LOC_835/a_8_216# OR2X1_LOC_835/a_36_216# OR2X1_LOC_835/Y VSS VDD OR2X1_LOC_835/A OR2X1_LOC_835/B OR2X1_LOC

XOR2X1_LOC_180 OR2X1_LOC_180/a_8_216# OR2X1_LOC_180/a_36_216# OR2X1_LOC_182/B VSS VDD OR2X1_LOC_439/B OR2X1_LOC_180/B OR2X1_LOC

XOR2X1_LOC_175 OR2X1_LOC_175/a_8_216# OR2X1_LOC_175/a_36_216# OR2X1_LOC_175/Y VSS VDD OR2X1_LOC_174/Y OR2X1_LOC_175/B OR2X1_LOC

XOR2X1_LOC_203 OR2X1_LOC_203/a_8_216# OR2X1_LOC_203/a_36_216# OR2X1_LOC_203/Y VSS VDD OR2X1_LOC_76/Y AND2X1_LOC_72/Y OR2X1_LOC

XOR2X1_LOC_174 OR2X1_LOC_174/a_8_216# OR2X1_LOC_174/a_36_216# OR2X1_LOC_174/Y VSS VDD OR2X1_LOC_174/A OR2X1_LOC_333/B OR2X1_LOC

XOR2X1_LOC_641 OR2X1_LOC_641/a_8_216# OR2X1_LOC_641/a_36_216# OR2X1_LOC_641/Y VSS VDD OR2X1_LOC_641/A OR2X1_LOC_641/B OR2X1_LOC

XOR2X1_LOC_786 OR2X1_LOC_786/a_8_216# OR2X1_LOC_786/a_36_216# OR2X1_LOC_786/Y VSS VDD OR2X1_LOC_786/A OR2X1_LOC_84/Y OR2X1_LOC

XOR2X1_LOC_444 OR2X1_LOC_444/a_8_216# OR2X1_LOC_444/a_36_216# OR2X1_LOC_469/B VSS VDD OR2X1_LOC_443/Y OR2X1_LOC_444/B OR2X1_LOC

XOR2X1_LOC_169 OR2X1_LOC_169/a_8_216# OR2X1_LOC_169/a_36_216# OR2X1_LOC_170/A VSS VDD OR2X1_LOC_703/B OR2X1_LOC_169/B OR2X1_LOC

XOR2X1_LOC_191 OR2X1_LOC_191/a_8_216# OR2X1_LOC_191/a_36_216# OR2X1_LOC_192/A VSS VDD OR2X1_LOC_190/Y OR2X1_LOC_191/B OR2X1_LOC

XOR2X1_LOC_555 OR2X1_LOC_555/a_8_216# OR2X1_LOC_555/a_36_216# OR2X1_LOC_562/B VSS VDD OR2X1_LOC_555/A OR2X1_LOC_555/B OR2X1_LOC

XOR2X1_LOC_402 OR2X1_LOC_402/a_8_216# OR2X1_LOC_402/a_36_216# OR2X1_LOC_402/Y VSS VDD OR2X1_LOC_401/Y OR2X1_LOC_402/B OR2X1_LOC

XOR2X1_LOC_773 OR2X1_LOC_773/a_8_216# OR2X1_LOC_773/a_36_216# OR2X1_LOC_773/Y VSS VDD OR2X1_LOC_772/Y OR2X1_LOC_773/B OR2X1_LOC

XOR2X1_LOC_718 OR2X1_LOC_718/a_8_216# OR2X1_LOC_718/a_36_216# OR2X1_LOC_722/B VSS VDD OR2X1_LOC_605/Y OR2X1_LOC_593/B OR2X1_LOC

XOR2X1_LOC_703 OR2X1_LOC_703/a_8_216# OR2X1_LOC_703/a_36_216# OR2X1_LOC_703/Y VSS VDD OR2X1_LOC_703/A OR2X1_LOC_703/B OR2X1_LOC

XOR2X1_LOC_388 OR2X1_LOC_388/a_8_216# OR2X1_LOC_388/a_36_216# OR2X1_LOC_390/B VSS VDD OR2X1_LOC_180/B OR2X1_LOC_703/B OR2X1_LOC

XOR2X1_LOC_201 OR2X1_LOC_201/a_8_216# OR2X1_LOC_201/a_36_216# OR2X1_LOC_201/Y VSS VDD OR2X1_LOC_201/A OR2X1_LOC_61/Y OR2X1_LOC

XOR2X1_LOC_336 OR2X1_LOC_336/a_8_216# OR2X1_LOC_336/a_36_216# OR2X1_LOC_337/A VSS VDD OR2X1_LOC_703/A OR2X1_LOC_538/A OR2X1_LOC

XOR2X1_LOC_623 OR2X1_LOC_623/a_8_216# OR2X1_LOC_623/a_36_216# OR2X1_LOC_624/A VSS VDD OR2X1_LOC_620/Y OR2X1_LOC_623/B OR2X1_LOC

XOR2X1_LOC_844 OR2X1_LOC_844/a_8_216# OR2X1_LOC_844/a_36_216# OR2X1_LOC_844/Y VSS VDD OR2X1_LOC_523/Y OR2X1_LOC_844/B OR2X1_LOC

XOR2X1_LOC_500 OR2X1_LOC_500/a_8_216# OR2X1_LOC_500/a_36_216# OR2X1_LOC_501/A VSS VDD OR2X1_LOC_500/A OR2X1_LOC_844/B OR2X1_LOC

XOR2X1_LOC_643 OR2X1_LOC_643/a_8_216# OR2X1_LOC_643/a_36_216# OR2X1_LOC_643/Y VSS VDD OR2X1_LOC_643/A OR2X1_LOC_539/B OR2X1_LOC

XAND2X1_LOC_639 AND2X1_LOC_639/a_36_24# AND2X1_LOC_651/B AND2X1_LOC_639/a_8_24# VSS VDD AND2X1_LOC_639/A AND2X1_LOC_639/B AND2X1_LOC

XAND2X1_LOC_774 AND2X1_LOC_774/a_36_24# AND2X1_LOC_810/A AND2X1_LOC_774/a_8_24# VSS VDD AND2X1_LOC_774/A AND2X1_LOC_773/Y AND2X1_LOC

XAND2X1_LOC_465 AND2X1_LOC_465/a_36_24# AND2X1_LOC_465/Y AND2X1_LOC_465/a_8_24# VSS VDD AND2X1_LOC_465/A AND2X1_LOC_456/Y AND2X1_LOC

XAND2X1_LOC_849 AND2X1_LOC_849/a_36_24# AND2X1_LOC_859/B AND2X1_LOC_849/a_8_24# VSS VDD AND2X1_LOC_849/A AND2X1_LOC_845/Y AND2X1_LOC

XAND2X1_LOC_354 AND2X1_LOC_354/a_36_24# AND2X1_LOC_354/Y AND2X1_LOC_354/a_8_24# VSS VDD AND2X1_LOC_798/A AND2X1_LOC_354/B AND2X1_LOC

XAND2X1_LOC_652 AND2X1_LOC_652/a_36_24# AND2X1_LOC_653/B AND2X1_LOC_652/a_8_24# VSS VDD AND2X1_LOC_468/B AND2X1_LOC_593/Y AND2X1_LOC

XAND2X1_LOC_474 AND2X1_LOC_474/a_36_24# AND2X1_LOC_474/Y AND2X1_LOC_474/a_8_24# VSS VDD AND2X1_LOC_474/A AND2X1_LOC_573/A AND2X1_LOC

XOR2X1_LOC_774 OR2X1_LOC_774/a_8_216# OR2X1_LOC_774/a_36_216# OR2X1_LOC_774/Y VSS VDD OR2X1_LOC_773/Y OR2X1_LOC_774/B OR2X1_LOC

XOR2X1_LOC_510 OR2X1_LOC_510/a_8_216# OR2X1_LOC_510/a_36_216# OR2X1_LOC_510/Y VSS VDD OR2X1_LOC_510/A OR2X1_LOC_508/Y OR2X1_LOC

XAND2X1_LOC_510 AND2X1_LOC_510/a_36_24# AND2X1_LOC_574/A AND2X1_LOC_510/a_8_24# VSS VDD AND2X1_LOC_510/A AND2X1_LOC_509/Y AND2X1_LOC

XOR2X1_LOC_849 OR2X1_LOC_849/a_8_216# OR2X1_LOC_849/a_36_216# OR2X1_LOC_859/A VSS VDD OR2X1_LOC_849/A OR2X1_LOC_844/Y OR2X1_LOC

XOR2X1_LOC_465 OR2X1_LOC_465/a_8_216# OR2X1_LOC_465/a_36_216# OR2X1_LOC_465/Y VSS VDD OR2X1_LOC_456/Y OR2X1_LOC_465/B OR2X1_LOC

XOR2X1_LOC_35 OR2X1_LOC_35/a_8_216# OR2X1_LOC_35/a_36_216# OR2X1_LOC_35/Y VSS VDD OR2X1_LOC_35/A OR2X1_LOC_35/B OR2X1_LOC

XAND2X1_LOC_35 AND2X1_LOC_35/a_36_24# AND2X1_LOC_35/Y AND2X1_LOC_35/a_8_24# VSS VDD AND2X1_LOC_33/Y AND2X1_LOC_34/Y AND2X1_LOC

XOR2X1_LOC_354 OR2X1_LOC_354/a_8_216# OR2X1_LOC_354/a_36_216# OR2X1_LOC_356/B VSS VDD OR2X1_LOC_354/A OR2X1_LOC_319/Y OR2X1_LOC

XOR2X1_LOC_474 OR2X1_LOC_474/a_8_216# OR2X1_LOC_474/a_36_216# OR2X1_LOC_474/Y VSS VDD OR2X1_LOC_404/Y OR2X1_LOC_474/B OR2X1_LOC

XOR2X1_LOC_652 OR2X1_LOC_652/a_8_216# OR2X1_LOC_652/a_36_216# OR2X1_LOC_653/A VSS VDD OR2X1_LOC_799/A OR2X1_LOC_468/A OR2X1_LOC

XAND2X1_LOC_455 AND2X1_LOC_455/a_36_24# AND2X1_LOC_465/A AND2X1_LOC_455/a_8_24# VSS VDD AND2X1_LOC_76/Y AND2X1_LOC_455/B AND2X1_LOC

XAND2X1_LOC_404 AND2X1_LOC_404/a_36_24# AND2X1_LOC_573/A AND2X1_LOC_404/a_8_24# VSS VDD AND2X1_LOC_404/A AND2X1_LOC_404/B AND2X1_LOC

XOR2X1_LOC_455 OR2X1_LOC_455/a_8_216# OR2X1_LOC_455/a_36_216# OR2X1_LOC_465/B VSS VDD OR2X1_LOC_455/A OR2X1_LOC_76/Y OR2X1_LOC

XOR2X1_LOC_404 OR2X1_LOC_404/a_8_216# OR2X1_LOC_404/a_36_216# OR2X1_LOC_404/Y VSS VDD OR2X1_LOC_404/A OR2X1_LOC_402/Y OR2X1_LOC

C4377 OR2X1_LOC_338/a_8_216# OR2X1_LOC_338/A 0.06fF
C7371 OR2X1_LOC_34/a_8_216# OR2X1_LOC_338/A 0.01fF
C18412 OR2X1_LOC_338/B OR2X1_LOC_338/A 0.06fF
C18441 OR2X1_LOC_35/A OR2X1_LOC_338/A 0.02fF
C23184 OR2X1_LOC_35/a_8_216# OR2X1_LOC_338/A 0.01fF
C24532 OR2X1_LOC_33/A OR2X1_LOC_338/A 0.01fF
C33419 OR2X1_LOC_34/B OR2X1_LOC_338/A 0.03fF
C35482 OR2X1_LOC_33/B OR2X1_LOC_338/A 0.16fF
C37571 OR2X1_LOC_654/A OR2X1_LOC_338/A 0.07fF
C37880 VDD OR2X1_LOC_338/A 0.12fF
C39626 OR2X1_LOC_35/Y OR2X1_LOC_338/A 0.01fF
C40993 OR2X1_LOC_33/a_8_216# OR2X1_LOC_338/A 0.01fF
C46968 OR2X1_LOC_34/A OR2X1_LOC_338/A 0.01fF
C49936 OR2X1_LOC_771/B OR2X1_LOC_338/A 0.07fF
C52233 OR2X1_LOC_35/B OR2X1_LOC_338/A 0.03fF
C56255 OR2X1_LOC_338/A VSS -0.39fF
C12768 VDD OR2X1_LOC_836/Y -0.00fF
C40423 OR2X1_LOC_836/Y OR2X1_LOC_835/Y 0.14fF
C51677 OR2X1_LOC_836/Y OR2X1_LOC_839/a_8_216# 0.39fF
C57359 OR2X1_LOC_836/Y VSS 0.18fF
C1383 OR2X1_LOC_243/A OR2X1_LOC_244/A 0.01fF
C29178 VDD OR2X1_LOC_243/A 0.12fF
C40769 OR2X1_LOC_243/A OR2X1_LOC_243/B 0.16fF
C57369 OR2X1_LOC_243/A VSS 0.18fF
C103 OR2X1_LOC_476/B OR2X1_LOC_472/B 0.01fF
C1810 OR2X1_LOC_472/B OR2X1_LOC_472/A 0.43fF
C2259 OR2X1_LOC_472/B AND2X1_LOC_34/a_8_24# 0.23fF
C34053 OR2X1_LOC_472/a_8_216# OR2X1_LOC_472/B 0.01fF
C41709 OR2X1_LOC_472/B OR2X1_LOC_27/Y 0.08fF
C51501 VDD OR2X1_LOC_472/B 0.12fF
C52444 OR2X1_LOC_462/B OR2X1_LOC_472/B 0.02fF
C53335 OR2X1_LOC_472/B OR2X1_LOC_416/Y 0.01fF
C57568 OR2X1_LOC_472/B VSS -0.09fF
C3267 AND2X1_LOC_841/B AND2X1_LOC_810/B 0.07fF
C3705 AND2X1_LOC_365/A AND2X1_LOC_810/B 0.07fF
C4406 AND2X1_LOC_388/Y AND2X1_LOC_810/B 0.01fF
C10838 AND2X1_LOC_567/a_8_24# AND2X1_LOC_810/B 0.03fF
C11380 AND2X1_LOC_337/B AND2X1_LOC_810/B 0.03fF
C11773 AND2X1_LOC_388/a_8_24# AND2X1_LOC_810/B 0.02fF
C13791 OR2X1_LOC_176/Y AND2X1_LOC_810/B 0.01fF
C14623 AND2X1_LOC_539/Y AND2X1_LOC_810/B 0.26fF
C16323 AND2X1_LOC_568/B AND2X1_LOC_810/B 0.03fF
C19865 AND2X1_LOC_354/a_8_24# AND2X1_LOC_810/B 0.02fF
C27354 AND2X1_LOC_810/A AND2X1_LOC_810/B 0.16fF
C30121 OR2X1_LOC_167/Y AND2X1_LOC_810/B 0.03fF
C30861 AND2X1_LOC_354/a_36_24# AND2X1_LOC_810/B 0.01fF
C31553 AND2X1_LOC_715/Y AND2X1_LOC_810/B 0.39fF
C32042 AND2X1_LOC_354/Y AND2X1_LOC_810/B 0.15fF
C33383 AND2X1_LOC_661/A AND2X1_LOC_810/B 0.04fF
C35190 AND2X1_LOC_798/A AND2X1_LOC_810/B 0.13fF
C35821 VDD AND2X1_LOC_810/B 0.21fF
C41435 AND2X1_LOC_354/B AND2X1_LOC_810/B 0.01fF
C43704 OR2X1_LOC_311/Y AND2X1_LOC_810/B 0.01fF
C46814 AND2X1_LOC_170/B AND2X1_LOC_810/B 0.07fF
C48833 AND2X1_LOC_356/a_8_24# AND2X1_LOC_810/B 0.20fF
C50995 OR2X1_LOC_312/Y AND2X1_LOC_810/B 0.07fF
C55957 AND2X1_LOC_535/Y AND2X1_LOC_810/B 0.19fF
C56584 AND2X1_LOC_810/B VSS 0.12fF
C13402 VDD AND2X1_LOC_473/Y 0.21fF
C16009 AND2X1_LOC_116/Y AND2X1_LOC_473/Y 0.09fF
C36174 AND2X1_LOC_473/Y AND2X1_LOC_476/a_8_24# 0.11fF
C38990 AND2X1_LOC_476/A AND2X1_LOC_473/Y 0.01fF
C43458 AND2X1_LOC_473/Y AND2X1_LOC_786/Y 0.04fF
C54208 AND2X1_LOC_715/A AND2X1_LOC_473/Y 0.03fF
C55099 AND2X1_LOC_76/Y AND2X1_LOC_473/Y 0.03fF
C56790 AND2X1_LOC_473/Y VSS -0.60fF
C8369 OR2X1_LOC_122/Y AND2X1_LOC_362/B 0.01fF
C12346 AND2X1_LOC_362/B AND2X1_LOC_227/Y 0.01fF
C16442 AND2X1_LOC_362/B AND2X1_LOC_560/B 0.01fF
C18922 AND2X1_LOC_362/B OR2X1_LOC_494/Y 0.07fF
C26960 AND2X1_LOC_362/B AND2X1_LOC_243/Y 0.37fF
C31393 AND2X1_LOC_362/B AND2X1_LOC_845/Y 0.09fF
C32143 AND2X1_LOC_362/B AND2X1_LOC_489/Y 0.03fF
C32507 AND2X1_LOC_554/Y AND2X1_LOC_362/B 0.07fF
C33313 AND2X1_LOC_362/B AND2X1_LOC_474/A 0.03fF
C36713 AND2X1_LOC_362/B AND2X1_LOC_573/A 0.07fF
C37097 AND2X1_LOC_362/B AND2X1_LOC_362/a_8_24# -0.01fF
C42708 AND2X1_LOC_362/B AND2X1_LOC_366/A 0.01fF
C46601 AND2X1_LOC_362/B VDD 0.25fF
C50095 AND2X1_LOC_362/B OR2X1_LOC_103/Y 0.01fF
C52121 AND2X1_LOC_541/Y AND2X1_LOC_362/B 0.03fF
C54328 OR2X1_LOC_91/Y AND2X1_LOC_362/B 0.04fF
C54775 AND2X1_LOC_362/B AND2X1_LOC_806/A 0.04fF
C57944 AND2X1_LOC_362/B VSS 0.28fF
C2995 OR2X1_LOC_656/B OR2X1_LOC_805/A 0.01fF
C7269 OR2X1_LOC_656/B OR2X1_LOC_656/a_8_216# 0.02fF
C10365 OR2X1_LOC_656/B OR2X1_LOC_559/a_8_216# 0.03fF
C24294 OR2X1_LOC_656/B OR2X1_LOC_216/a_8_216# 0.04fF
C26289 OR2X1_LOC_656/B OR2X1_LOC_559/B 0.05fF
C28023 OR2X1_LOC_656/B OR2X1_LOC_520/Y 0.56fF
C28389 OR2X1_LOC_656/B OR2X1_LOC_656/Y 0.40fF
C32531 OR2X1_LOC_656/B VDD 0.09fF
C35122 OR2X1_LOC_656/B OR2X1_LOC_216/A 0.03fF
C37987 OR2X1_LOC_656/B OR2X1_LOC_641/A 0.07fF
C39024 OR2X1_LOC_656/B OR2X1_LOC_643/A 0.07fF
C41683 OR2X1_LOC_656/B OR2X1_LOC_227/Y 0.01fF
C47269 OR2X1_LOC_656/B OR2X1_LOC_340/Y 0.02fF
C47408 OR2X1_LOC_656/B AND2X1_LOC_88/Y 0.81fF
C48958 OR2X1_LOC_656/B OR2X1_LOC_624/A 0.38fF
C49845 OR2X1_LOC_656/B OR2X1_LOC_216/Y 0.10fF
C52904 OR2X1_LOC_656/B OR2X1_LOC_340/a_8_216# 0.02fF
C58025 OR2X1_LOC_656/B VSS 0.53fF
C4765 AND2X1_LOC_856/B AND2X1_LOC_856/a_8_24# 0.01fF
C12664 AND2X1_LOC_539/Y AND2X1_LOC_856/B 0.01fF
C15821 AND2X1_LOC_856/B AND2X1_LOC_863/A 0.05fF
C22808 AND2X1_LOC_856/B OR2X1_LOC_599/Y 0.12fF
C33930 VDD AND2X1_LOC_856/B 0.01fF
C39562 AND2X1_LOC_390/B AND2X1_LOC_856/B 0.03fF
C41718 OR2X1_LOC_311/Y AND2X1_LOC_856/B 0.01fF
C57085 AND2X1_LOC_856/B VSS 0.19fF
C3 AND2X1_LOC_729/Y AND2X1_LOC_191/Y 0.03fF
C299 AND2X1_LOC_729/Y AND2X1_LOC_658/B 0.03fF
C2491 AND2X1_LOC_729/Y AND2X1_LOC_447/Y 0.01fF
C2906 AND2X1_LOC_729/Y AND2X1_LOC_209/a_8_24# 0.01fF
C3108 AND2X1_LOC_729/Y OR2X1_LOC_679/A 0.01fF
C3380 AND2X1_LOC_729/Y AND2X1_LOC_722/A 0.07fF
C4602 AND2X1_LOC_729/Y AND2X1_LOC_841/B 0.07fF
C5514 AND2X1_LOC_729/Y AND2X1_LOC_147/Y 0.01fF
C7474 AND2X1_LOC_729/Y AND2X1_LOC_544/Y 0.03fF
C10639 AND2X1_LOC_729/Y AND2X1_LOC_624/A 0.03fF
C11402 AND2X1_LOC_729/Y OR2X1_LOC_524/Y 0.03fF
C13241 AND2X1_LOC_729/Y OR2X1_LOC_601/Y 0.13fF
C13427 AND2X1_LOC_729/Y OR2X1_LOC_142/Y 0.02fF
C16998 AND2X1_LOC_728/Y AND2X1_LOC_729/Y 0.42fF
C18689 AND2X1_LOC_729/Y AND2X1_LOC_703/a_8_24# 0.03fF
C21295 AND2X1_LOC_729/Y AND2X1_LOC_192/Y 0.03fF
C23735 AND2X1_LOC_729/Y OR2X1_LOC_485/Y 0.39fF
C24290 AND2X1_LOC_729/Y AND2X1_LOC_602/a_8_24# 0.02fF
C26598 AND2X1_LOC_729/Y AND2X1_LOC_705/Y 0.01fF
C30446 AND2X1_LOC_729/Y OR2X1_LOC_679/a_8_216# 0.01fF
C30457 AND2X1_LOC_729/Y AND2X1_LOC_658/A 0.03fF
C31437 AND2X1_LOC_729/Y OR2X1_LOC_680/Y 0.02fF
C31493 AND2X1_LOC_729/Y OR2X1_LOC_167/Y 0.05fF
C32900 AND2X1_LOC_729/Y AND2X1_LOC_715/Y 0.83fF
C34092 AND2X1_LOC_729/Y AND2X1_LOC_796/A 0.03fF
C34655 AND2X1_LOC_729/Y OR2X1_LOC_526/Y 0.03fF
C35208 AND2X1_LOC_729/Y AND2X1_LOC_645/A 0.01fF
C35439 AND2X1_LOC_729/Y AND2X1_LOC_703/Y 0.01fF
C35934 AND2X1_LOC_729/Y OR2X1_LOC_679/a_36_216# 0.01fF
C36657 AND2X1_LOC_729/Y AND2X1_LOC_209/Y 0.01fF
C36890 AND2X1_LOC_729/Y AND2X1_LOC_728/a_8_24# 0.01fF
C37180 AND2X1_LOC_729/Y VDD 0.91fF
C38027 AND2X1_LOC_729/Y OR2X1_LOC_600/Y 0.05fF
C40134 AND2X1_LOC_729/Y AND2X1_LOC_705/a_8_24# 0.01fF
C41469 AND2X1_LOC_729/Y OR2X1_LOC_679/Y 0.01fF
C45083 AND2X1_LOC_729/Y OR2X1_LOC_189/Y 0.03fF
C45093 AND2X1_LOC_729/Y OR2X1_LOC_152/Y 0.32fF
C45849 AND2X1_LOC_729/Y OR2X1_LOC_441/Y 0.03fF
C52191 AND2X1_LOC_729/Y AND2X1_LOC_724/A 0.01fF
C52395 AND2X1_LOC_729/Y OR2X1_LOC_312/Y 0.10fF
C52769 AND2X1_LOC_729/Y OR2X1_LOC_679/B 0.01fF
C58132 AND2X1_LOC_729/Y VSS 0.11fF
C7526 AND2X1_LOC_547/Y AND2X1_LOC_550/A 0.14fF
C11299 AND2X1_LOC_547/Y OR2X1_LOC_524/Y 0.06fF
C21489 AND2X1_LOC_547/Y AND2X1_LOC_564/B 0.02fF
C26125 AND2X1_LOC_547/Y AND2X1_LOC_475/Y 0.23fF
C27825 AND2X1_LOC_547/Y AND2X1_LOC_550/a_8_24# 0.03fF
C31616 AND2X1_LOC_547/Y AND2X1_LOC_476/Y 0.02fF
C33302 AND2X1_LOC_547/Y AND2X1_LOC_565/B 0.15fF
C37089 AND2X1_LOC_547/Y VDD 0.01fF
C38819 AND2X1_LOC_547/Y AND2X1_LOC_550/a_36_24# 0.01fF
C43246 AND2X1_LOC_547/Y AND2X1_LOC_475/a_8_24# 0.01fF
C44972 AND2X1_LOC_547/Y OR2X1_LOC_189/Y 0.03fF
C56119 AND2X1_LOC_547/Y AND2X1_LOC_191/Y 0.03fF
C56138 AND2X1_LOC_547/Y AND2X1_LOC_711/Y 0.09fF
C58074 AND2X1_LOC_547/Y VSS 0.04fF
C6349 AND2X1_LOC_715/A AND2X1_LOC_476/A 0.02fF
C9178 AND2X1_LOC_357/B AND2X1_LOC_715/A 0.10fF
C10092 OR2X1_LOC_521/Y AND2X1_LOC_715/A 0.01fF
C10836 AND2X1_LOC_715/A AND2X1_LOC_786/Y 0.02fF
C15516 AND2X1_LOC_326/B AND2X1_LOC_715/A 0.02fF
C22075 AND2X1_LOC_784/A AND2X1_LOC_715/A 0.02fF
C22461 AND2X1_LOC_76/Y AND2X1_LOC_715/A 0.45fF
C23378 AND2X1_LOC_211/B AND2X1_LOC_715/A 0.12fF
C28234 AND2X1_LOC_810/A AND2X1_LOC_715/A 0.03fF
C32883 AND2X1_LOC_392/A AND2X1_LOC_715/A 0.03fF
C36084 AND2X1_LOC_715/A AND2X1_LOC_798/A 0.20fF
C36655 VDD AND2X1_LOC_715/A 0.22fF
C42366 AND2X1_LOC_715/A AND2X1_LOC_354/B 0.06fF
C48773 AND2X1_LOC_566/B AND2X1_LOC_715/A 0.03fF
C51802 AND2X1_LOC_716/Y AND2X1_LOC_715/A 0.07fF
C54450 AND2X1_LOC_715/A AND2X1_LOC_727/A 0.03fF
C57392 AND2X1_LOC_715/A VSS 0.55fF
C182 AND2X1_LOC_339/B AND2X1_LOC_61/Y 0.23fF
C1035 AND2X1_LOC_339/Y AND2X1_LOC_339/B 0.21fF
C4134 AND2X1_LOC_339/B AND2X1_LOC_339/a_36_24# 0.01fF
C10061 AND2X1_LOC_339/B AND2X1_LOC_649/B 0.01fF
C14474 AND2X1_LOC_339/B AND2X1_LOC_476/A 0.14fF
C20426 AND2X1_LOC_339/B OR2X1_LOC_75/Y 0.01fF
C22898 AND2X1_LOC_339/B OR2X1_LOC_265/Y 0.03fF
C25252 AND2X1_LOC_773/Y AND2X1_LOC_339/B 0.03fF
C26515 OR2X1_LOC_135/Y AND2X1_LOC_339/B 0.03fF
C28613 AND2X1_LOC_340/Y AND2X1_LOC_339/B 1.74fF
C30187 AND2X1_LOC_339/B AND2X1_LOC_643/a_8_24# 0.01fF
C39726 AND2X1_LOC_303/A AND2X1_LOC_339/B 0.03fF
C44814 VDD AND2X1_LOC_339/B 0.39fF
C49318 AND2X1_LOC_339/B AND2X1_LOC_339/a_8_24# 0.04fF
C53198 AND2X1_LOC_339/B AND2X1_LOC_831/Y 0.01fF
C53509 AND2X1_LOC_339/B AND2X1_LOC_139/B 0.01fF
C57725 AND2X1_LOC_339/B VSS 0.23fF
C766 AND2X1_LOC_703/a_8_24# AND2X1_LOC_841/B 0.06fF
C4633 AND2X1_LOC_784/A AND2X1_LOC_841/B 0.07fF
C5476 AND2X1_LOC_356/B AND2X1_LOC_841/B 0.11fF
C5927 AND2X1_LOC_211/B AND2X1_LOC_841/B 0.07fF
C10393 AND2X1_LOC_841/B OR2X1_LOC_423/Y 0.15fF
C10886 AND2X1_LOC_810/A AND2X1_LOC_841/B 0.03fF
C13906 AND2X1_LOC_841/B AND2X1_LOC_476/Y 0.04fF
C14304 AND2X1_LOC_706/Y AND2X1_LOC_841/B 0.02fF
C15112 AND2X1_LOC_715/Y AND2X1_LOC_841/B 0.07fF
C15573 AND2X1_LOC_392/A AND2X1_LOC_841/B 0.07fF
C17000 AND2X1_LOC_841/B AND2X1_LOC_661/A 0.03fF
C17265 AND2X1_LOC_714/B AND2X1_LOC_841/B 0.07fF
C17639 AND2X1_LOC_703/Y AND2X1_LOC_841/B 0.15fF
C19438 VDD AND2X1_LOC_841/B 0.51fF
C25107 AND2X1_LOC_390/B AND2X1_LOC_841/B 0.07fF
C27685 AND2X1_LOC_831/Y AND2X1_LOC_841/B 0.01fF
C28689 AND2X1_LOC_714/a_8_24# AND2X1_LOC_841/B 0.20fF
C30217 AND2X1_LOC_170/B AND2X1_LOC_841/B 0.01fF
C31262 AND2X1_LOC_566/B AND2X1_LOC_841/B 0.03fF
C34257 AND2X1_LOC_716/Y AND2X1_LOC_841/B 0.07fF
C34331 OR2X1_LOC_312/Y AND2X1_LOC_841/B 0.03fF
C36899 AND2X1_LOC_727/A AND2X1_LOC_841/B 0.03fF
C39299 AND2X1_LOC_535/Y AND2X1_LOC_841/B 0.07fF
C39698 AND2X1_LOC_714/a_36_24# AND2X1_LOC_841/B 0.01fF
C40643 OR2X1_LOC_109/Y AND2X1_LOC_841/B 0.02fF
C49941 AND2X1_LOC_841/a_8_24# AND2X1_LOC_841/B 0.09fF
C50554 AND2X1_LOC_567/a_8_24# AND2X1_LOC_841/B 0.02fF
C54245 AND2X1_LOC_539/Y AND2X1_LOC_841/B 0.08fF
C54321 AND2X1_LOC_326/B AND2X1_LOC_841/B 0.23fF
C55408 AND2X1_LOC_851/B AND2X1_LOC_841/B 0.01fF
C56045 AND2X1_LOC_568/B AND2X1_LOC_841/B 0.22fF
C57133 AND2X1_LOC_841/B VSS -0.56fF
C9561 VDD AND2X1_LOC_783/B 0.06fF
C15832 AND2X1_LOC_213/B AND2X1_LOC_783/B 0.10fF
C40268 AND2X1_LOC_783/B AND2X1_LOC_779/Y 0.33fF
C56441 AND2X1_LOC_783/B VSS 0.05fF
C8030 AND2X1_LOC_464/Y AND2X1_LOC_786/Y 0.02fF
C18189 AND2X1_LOC_564/B AND2X1_LOC_464/Y 0.01fF
C33937 VDD AND2X1_LOC_464/Y 0.21fF
C37620 AND2X1_LOC_721/Y AND2X1_LOC_464/Y 0.01fF
C37844 AND2X1_LOC_464/Y AND2X1_LOC_471/a_8_24# 0.18fF
C57048 AND2X1_LOC_464/Y VSS -0.13fF
C3522 AND2X1_LOC_520/Y AND2X1_LOC_476/A 0.04fF
C7916 AND2X1_LOC_520/Y AND2X1_LOC_786/Y 0.05fF
C19515 AND2X1_LOC_76/Y AND2X1_LOC_520/Y 0.02fF
C21235 AND2X1_LOC_520/Y AND2X1_LOC_642/a_8_24# 0.01fF
C33818 VDD AND2X1_LOC_520/Y 0.18fF
C34700 AND2X1_LOC_520/Y AND2X1_LOC_642/Y 0.01fF
C35674 AND2X1_LOC_520/Y OR2X1_LOC_416/Y 0.04fF
C54447 AND2X1_LOC_559/a_8_24# AND2X1_LOC_520/Y 0.11fF
C57007 AND2X1_LOC_520/Y VSS 0.22fF
C9145 VDD AND2X1_LOC_769/Y 0.25fF
C33246 AND2X1_LOC_769/Y AND2X1_LOC_771/a_8_24# 0.19fF
C43933 AND2X1_LOC_771/B AND2X1_LOC_769/Y 0.09fF
C56356 AND2X1_LOC_769/Y VSS 0.10fF
C132 AND2X1_LOC_196/Y AND2X1_LOC_199/a_8_24# 0.03fF
C23444 VDD AND2X1_LOC_196/Y 0.01fF
C27609 AND2X1_LOC_196/Y AND2X1_LOC_199/a_36_24# 0.01fF
C38531 AND2X1_LOC_199/A AND2X1_LOC_196/Y 0.28fF
C57445 AND2X1_LOC_196/Y VSS 0.20fF
C2016 AND2X1_LOC_794/B AND2X1_LOC_840/B 0.10fF
C2052 VDD AND2X1_LOC_840/B 1.59fF
C2568 AND2X1_LOC_486/Y AND2X1_LOC_840/B 0.07fF
C5740 AND2X1_LOC_721/Y AND2X1_LOC_840/B 0.03fF
C5794 OR2X1_LOC_482/Y AND2X1_LOC_840/B 0.02fF
C9825 OR2X1_LOC_91/Y AND2X1_LOC_840/B 0.10fF
C11895 OR2X1_LOC_525/Y AND2X1_LOC_840/B 0.84fF
C14178 AND2X1_LOC_840/B AND2X1_LOC_675/A 0.10fF
C19667 AND2X1_LOC_727/A AND2X1_LOC_840/B 0.05fF
C20998 OR2X1_LOC_437/Y AND2X1_LOC_840/B 0.44fF
C22899 AND2X1_LOC_840/B OR2X1_LOC_373/Y 0.10fF
C23424 OR2X1_LOC_109/Y AND2X1_LOC_840/B 0.05fF
C24657 AND2X1_LOC_794/A AND2X1_LOC_840/B 0.36fF
C25881 OR2X1_LOC_495/Y AND2X1_LOC_840/B 0.19fF
C31384 AND2X1_LOC_833/a_8_24# AND2X1_LOC_840/B 0.01fF
C32068 AND2X1_LOC_840/B AND2X1_LOC_786/Y 0.10fF
C35484 OR2X1_LOC_177/Y AND2X1_LOC_840/B 0.05fF
C36830 AND2X1_LOC_840/A AND2X1_LOC_840/B 0.49fF
C39257 AND2X1_LOC_776/Y AND2X1_LOC_840/B 0.10fF
C42274 AND2X1_LOC_564/B AND2X1_LOC_840/B 0.10fF
C43343 AND2X1_LOC_784/A AND2X1_LOC_840/B 0.10fF
C47699 AND2X1_LOC_840/a_8_24# AND2X1_LOC_840/B 0.05fF
C52671 AND2X1_LOC_840/B AND2X1_LOC_476/Y 0.10fF
C55885 AND2X1_LOC_810/Y AND2X1_LOC_840/B 0.10fF
C57021 AND2X1_LOC_840/B VSS 0.34fF
C18190 AND2X1_LOC_779/Y AND2X1_LOC_783/a_8_24# 0.19fF
C26849 VDD AND2X1_LOC_779/Y 0.25fF
C56310 AND2X1_LOC_779/Y VSS 0.10fF
C5924 AND2X1_LOC_720/a_8_24# OR2X1_LOC_669/Y 0.06fF
C14818 OR2X1_LOC_494/Y OR2X1_LOC_669/Y 0.07fF
C24291 OR2X1_LOC_669/Y AND2X1_LOC_848/Y 0.32fF
C35211 OR2X1_LOC_669/Y AND2X1_LOC_859/a_8_24# 0.23fF
C38519 AND2X1_LOC_366/A OR2X1_LOC_669/Y 0.19fF
C42383 VDD OR2X1_LOC_669/Y 0.12fF
C42514 OR2X1_LOC_251/Y OR2X1_LOC_669/Y 0.01fF
C45901 AND2X1_LOC_720/Y OR2X1_LOC_669/Y 0.03fF
C46223 AND2X1_LOC_721/Y OR2X1_LOC_669/Y 0.01fF
C51099 OR2X1_LOC_667/Y OR2X1_LOC_669/Y 0.04fF
C51498 AND2X1_LOC_721/a_8_24# OR2X1_LOC_669/Y 0.01fF
C53352 OR2X1_LOC_669/Y AND2X1_LOC_721/A 0.06fF
C57334 OR2X1_LOC_669/Y VSS 0.28fF
C2511 AND2X1_LOC_391/Y AND2X1_LOC_342/Y 0.12fF
C6357 AND2X1_LOC_554/B AND2X1_LOC_342/Y 0.02fF
C11080 AND2X1_LOC_342/Y AND2X1_LOC_349/a_36_24# 0.01fF
C12237 VDD AND2X1_LOC_342/Y 0.02fF
C23138 AND2X1_LOC_342/Y AND2X1_LOC_721/A 0.01fF
C45063 AND2X1_LOC_342/Y AND2X1_LOC_349/a_8_24# 0.07fF
C57356 AND2X1_LOC_342/Y VSS -0.23fF
C7293 OR2X1_LOC_792/Y OR2X1_LOC_288/A 0.01fF
C13721 OR2X1_LOC_288/A OR2X1_LOC_286/Y 0.12fF
C15710 VDD OR2X1_LOC_288/A 0.12fF
C26850 OR2X1_LOC_791/B OR2X1_LOC_288/A 0.01fF
C57197 OR2X1_LOC_288/A VSS -0.17fF
C1230 OR2X1_LOC_850/A OR2X1_LOC_362/A 0.02fF
C10576 OR2X1_LOC_850/A OR2X1_LOC_349/A 0.28fF
C27589 OR2X1_LOC_850/a_8_216# OR2X1_LOC_850/A 0.02fF
C36038 OR2X1_LOC_850/B OR2X1_LOC_850/A 0.18fF
C38553 OR2X1_LOC_858/B OR2X1_LOC_850/A 0.03fF
C57801 OR2X1_LOC_850/A VSS 0.16fF
C860 OR2X1_LOC_632/A OR2X1_LOC_574/A 0.04fF
C10859 OR2X1_LOC_632/A OR2X1_LOC_140/B 0.01fF
C14360 VDD OR2X1_LOC_632/A -0.00fF
C16342 OR2X1_LOC_632/A OR2X1_LOC_115/B 0.01fF
C34242 OR2X1_LOC_632/A OR2X1_LOC_630/Y 0.06fF
C37654 OR2X1_LOC_632/A OR2X1_LOC_575/A 0.01fF
C39764 OR2X1_LOC_632/A OR2X1_LOC_632/a_8_216# 0.39fF
C57655 OR2X1_LOC_632/A VSS 0.18fF
C1331 AND2X1_LOC_286/Y AND2X1_LOC_288/a_36_24# 0.01fF
C26646 AND2X1_LOC_719/Y AND2X1_LOC_286/Y 0.04fF
C29726 AND2X1_LOC_286/Y AND2X1_LOC_287/Y 1.01fF
C37313 AND2X1_LOC_859/Y AND2X1_LOC_286/Y 0.02fF
C38172 OR2X1_LOC_251/Y AND2X1_LOC_286/Y 0.01fF
C40717 AND2X1_LOC_286/Y AND2X1_LOC_288/a_8_24# 0.03fF
C45465 AND2X1_LOC_850/Y AND2X1_LOC_286/Y 0.08fF
C56554 AND2X1_LOC_286/Y VSS 0.10fF
C6355 AND2X1_LOC_489/Y AND2X1_LOC_572/A 0.37fF
C6505 AND2X1_LOC_489/Y AND2X1_LOC_772/a_8_24# 0.03fF
C9005 AND2X1_LOC_557/Y AND2X1_LOC_489/Y 0.01fF
C9341 AND2X1_LOC_563/A AND2X1_LOC_489/Y 0.02fF
C9479 AND2X1_LOC_489/Y AND2X1_LOC_717/B 0.09fF
C21241 AND2X1_LOC_489/Y AND2X1_LOC_558/a_8_24# 0.22fF
C23878 AND2X1_LOC_554/Y AND2X1_LOC_489/Y 0.14fF
C23923 AND2X1_LOC_489/Y OR2X1_LOC_280/Y 0.14fF
C26715 AND2X1_LOC_489/Y AND2X1_LOC_561/B 0.65fF
C28066 AND2X1_LOC_489/Y AND2X1_LOC_573/A 0.02fF
C30826 AND2X1_LOC_561/a_8_24# AND2X1_LOC_489/Y 0.02fF
C30851 OR2X1_LOC_106/Y AND2X1_LOC_489/Y 0.21fF
C31883 AND2X1_LOC_489/Y AND2X1_LOC_554/B 0.01fF
C36293 AND2X1_LOC_571/B AND2X1_LOC_489/Y 0.01fF
C37653 VDD AND2X1_LOC_489/Y 0.21fF
C45530 OR2X1_LOC_91/Y AND2X1_LOC_489/Y 0.03fF
C47603 AND2X1_LOC_554/a_8_24# AND2X1_LOC_489/Y 0.01fF
C53996 AND2X1_LOC_772/B AND2X1_LOC_489/Y 0.18fF
C57754 AND2X1_LOC_489/Y VSS 0.28fF
C7439 AND2X1_LOC_338/A AND2X1_LOC_338/a_8_24# 0.01fF
C31188 VDD AND2X1_LOC_338/A -0.00fF
C37864 AND2X1_LOC_338/Y AND2X1_LOC_338/A 0.92fF
C39167 AND2X1_LOC_338/A OR2X1_LOC_171/Y 0.28fF
C52571 AND2X1_LOC_338/A AND2X1_LOC_334/Y 0.06fF
C57663 AND2X1_LOC_338/A VSS 0.10fF
C174 AND2X1_LOC_454/A OR2X1_LOC_423/Y 0.01fF
C20397 AND2X1_LOC_605/Y AND2X1_LOC_454/A 0.02fF
C32426 AND2X1_LOC_454/A OR2X1_LOC_424/Y -0.00fF
C32517 AND2X1_LOC_707/Y AND2X1_LOC_454/A 0.20fF
C35971 AND2X1_LOC_454/a_8_24# AND2X1_LOC_454/A 0.03fF
C36061 AND2X1_LOC_449/Y AND2X1_LOC_454/A 0.09fF
C37305 AND2X1_LOC_452/Y AND2X1_LOC_454/A 0.01fF
C43540 AND2X1_LOC_454/A AND2X1_LOC_449/a_8_24# 0.02fF
C56621 AND2X1_LOC_454/A VSS 0.26fF
C17165 AND2X1_LOC_707/Y AND2X1_LOC_714/B 0.07fF
C22013 AND2X1_LOC_714/B AND2X1_LOC_452/Y 0.01fF
C40777 AND2X1_LOC_714/B OR2X1_LOC_423/Y 0.01fF
C44792 AND2X1_LOC_706/Y AND2X1_LOC_714/B 0.19fF
C48347 AND2X1_LOC_703/Y AND2X1_LOC_714/B 0.01fF
C50061 VDD AND2X1_LOC_714/B 0.35fF
C57819 AND2X1_LOC_714/B VSS 0.22fF
C1692 AND2X1_LOC_340/Y AND2X1_LOC_227/Y 0.10fF
C3266 AND2X1_LOC_227/Y OR2X1_LOC_88/Y 0.24fF
C3660 AND2X1_LOC_227/Y AND2X1_LOC_216/A 0.02fF
C3984 OR2X1_LOC_280/Y AND2X1_LOC_227/Y 0.03fF
C6316 AND2X1_LOC_719/Y AND2X1_LOC_227/Y 0.03fF
C7294 AND2X1_LOC_553/A AND2X1_LOC_227/Y 0.55fF
C8211 AND2X1_LOC_227/Y AND2X1_LOC_573/A 0.01fF
C9091 AND2X1_LOC_456/Y AND2X1_LOC_227/Y 0.02fF
C9420 AND2X1_LOC_340/a_8_24# AND2X1_LOC_227/Y 0.03fF
C10381 AND2X1_LOC_227/Y AND2X1_LOC_842/B 0.29fF
C10593 OR2X1_LOC_134/Y AND2X1_LOC_227/Y 0.02fF
C10989 OR2X1_LOC_106/Y AND2X1_LOC_227/Y 0.03fF
C11121 AND2X1_LOC_227/Y AND2X1_LOC_139/a_8_24# 0.01fF
C14100 AND2X1_LOC_392/A AND2X1_LOC_227/Y 0.03fF
C14669 AND2X1_LOC_227/Y AND2X1_LOC_137/a_8_24# 0.01fF
C16621 AND2X1_LOC_227/Y AND2X1_LOC_842/a_8_24# 0.09fF
C16631 AND2X1_LOC_227/Y AND2X1_LOC_141/A 0.01fF
C17855 VDD AND2X1_LOC_227/Y 0.44fF
C18375 AND2X1_LOC_486/Y AND2X1_LOC_227/Y 0.03fF
C20209 AND2X1_LOC_227/Y AND2X1_LOC_139/A 0.01fF
C20451 AND2X1_LOC_340/a_36_24# AND2X1_LOC_227/Y 0.02fF
C21384 OR2X1_LOC_103/Y AND2X1_LOC_227/Y 0.02fF
C21685 AND2X1_LOC_721/Y AND2X1_LOC_227/Y 0.02fF
C22311 AND2X1_LOC_227/Y AND2X1_LOC_523/Y 0.26fF
C22645 AND2X1_LOC_191/B AND2X1_LOC_227/Y 0.12fF
C23053 AND2X1_LOC_768/a_8_24# AND2X1_LOC_227/Y 0.01fF
C23445 AND2X1_LOC_541/Y AND2X1_LOC_227/Y 0.52fF
C25127 AND2X1_LOC_227/Y AND2X1_LOC_509/a_8_24# 0.10fF
C25616 OR2X1_LOC_91/Y AND2X1_LOC_227/Y 0.03fF
C26433 AND2X1_LOC_227/Y AND2X1_LOC_139/B 0.06fF
C27718 OR2X1_LOC_497/Y AND2X1_LOC_227/Y 0.11fF
C27755 AND2X1_LOC_227/Y AND2X1_LOC_844/a_8_24# 0.01fF
C33975 AND2X1_LOC_772/B AND2X1_LOC_227/Y 0.01fF
C34343 AND2X1_LOC_553/a_8_24# AND2X1_LOC_227/Y 0.01fF
C36636 AND2X1_LOC_227/Y OR2X1_LOC_184/Y 0.98fF
C38622 OR2X1_LOC_132/Y AND2X1_LOC_227/Y 0.02fF
C38744 AND2X1_LOC_227/Y AND2X1_LOC_849/A 0.01fF
C41081 AND2X1_LOC_227/Y AND2X1_LOC_242/B 0.19fF
C43877 AND2X1_LOC_560/B AND2X1_LOC_227/Y 0.12fF
C45508 AND2X1_LOC_563/A AND2X1_LOC_227/Y 0.01fF
C45623 AND2X1_LOC_227/Y AND2X1_LOC_717/B 0.03fF
C48752 AND2X1_LOC_227/Y AND2X1_LOC_656/Y 0.03fF
C48932 AND2X1_LOC_227/Y AND2X1_LOC_772/Y 0.03fF
C50414 OR2X1_LOC_262/Y AND2X1_LOC_227/Y 1.73fF
C50890 AND2X1_LOC_227/Y OR2X1_LOC_503/Y 0.10fF
C52039 AND2X1_LOC_227/Y OR2X1_LOC_265/Y 0.17fF
C57303 AND2X1_LOC_227/Y VSS 0.22fF
C743 OR2X1_LOC_303/B OR2X1_LOC_374/Y 0.57fF
C3142 VDD OR2X1_LOC_303/B 0.08fF
C9254 OR2X1_LOC_440/A OR2X1_LOC_303/B 0.03fF
C9595 OR2X1_LOC_778/Y OR2X1_LOC_303/B 0.05fF
C12372 OR2X1_LOC_303/B OR2X1_LOC_180/B 0.03fF
C14212 OR2X1_LOC_703/A OR2X1_LOC_303/B 0.01fF
C14556 OR2X1_LOC_336/a_8_216# OR2X1_LOC_303/B 0.01fF
C15305 OR2X1_LOC_303/B OR2X1_LOC_593/B 0.03fF
C15344 OR2X1_LOC_303/a_8_216# OR2X1_LOC_303/B 0.01fF
C17746 OR2X1_LOC_303/B OR2X1_LOC_365/B 0.02fF
C20227 OR2X1_LOC_787/Y OR2X1_LOC_303/B 0.08fF
C20546 OR2X1_LOC_439/B OR2X1_LOC_303/B 0.13fF
C25588 OR2X1_LOC_337/A OR2X1_LOC_303/B 0.01fF
C26384 OR2X1_LOC_566/A OR2X1_LOC_303/B 0.77fF
C30805 OR2X1_LOC_76/A OR2X1_LOC_303/B 0.28fF
C33457 OR2X1_LOC_170/Y OR2X1_LOC_303/B 0.20fF
C40901 OR2X1_LOC_605/A OR2X1_LOC_303/B 0.18fF
C41932 OR2X1_LOC_318/B OR2X1_LOC_303/B 0.15fF
C43055 OR2X1_LOC_794/A OR2X1_LOC_303/B 0.03fF
C52026 OR2X1_LOC_97/A OR2X1_LOC_303/B 0.18fF
C54078 OR2X1_LOC_303/B OR2X1_LOC_605/Y 0.81fF
C56369 OR2X1_LOC_303/B VSS 0.28fF
C2690 OR2X1_LOC_542/B OR2X1_LOC_552/A 0.12fF
C3111 OR2X1_LOC_787/B OR2X1_LOC_552/A 0.72fF
C11662 OR2X1_LOC_552/a_8_216# OR2X1_LOC_552/A 0.04fF
C20952 OR2X1_LOC_542/a_8_216# OR2X1_LOC_552/A 0.01fF
C31884 OR2X1_LOC_552/B OR2X1_LOC_552/A 0.15fF
C34060 OR2X1_LOC_147/B OR2X1_LOC_552/A 0.03fF
C51595 VDD OR2X1_LOC_552/A 0.07fF
C56484 OR2X1_LOC_552/A VSS 0.15fF
C13959 OR2X1_LOC_303/A OR2X1_LOC_326/B 0.17fF
C16408 OR2X1_LOC_303/A OR2X1_LOC_703/A 0.03fF
C28628 OR2X1_LOC_303/A OR2X1_LOC_566/A 0.06fF
C36598 OR2X1_LOC_303/A OR2X1_LOC_308/Y 0.20fF
C55632 OR2X1_LOC_303/A OR2X1_LOC_620/Y 0.01fF
C58107 OR2X1_LOC_303/A VSS 0.22fF
C197 VDD OR2X1_LOC_450/Y -0.00fF
C15198 OR2X1_LOC_450/Y OR2X1_LOC_449/B 0.27fF
C15495 OR2X1_LOC_450/Y OR2X1_LOC_452/a_8_216# 0.01fF
C21061 OR2X1_LOC_452/A OR2X1_LOC_450/Y 0.06fF
C37527 OR2X1_LOC_450/Y OR2X1_LOC_467/A 0.73fF
C57505 OR2X1_LOC_450/Y VSS 0.08fF
C10106 AND2X1_LOC_347/B AND2X1_LOC_848/Y 0.04fF
C12701 AND2X1_LOC_711/a_36_24# AND2X1_LOC_848/Y 0.01fF
C16608 OR2X1_LOC_258/Y AND2X1_LOC_848/Y 0.03fF
C18227 AND2X1_LOC_347/Y AND2X1_LOC_848/Y 0.80fF
C21090 AND2X1_LOC_555/Y AND2X1_LOC_848/Y 0.03fF
C26759 AND2X1_LOC_848/Y AND2X1_LOC_859/a_8_24# 0.10fF
C29815 AND2X1_LOC_848/Y AND2X1_LOC_849/a_8_24# 0.01fF
C30072 AND2X1_LOC_366/A AND2X1_LOC_848/Y 0.03fF
C31075 OR2X1_LOC_295/Y AND2X1_LOC_848/Y 0.03fF
C33844 VDD AND2X1_LOC_848/Y 0.15fF
C33964 OR2X1_LOC_251/Y AND2X1_LOC_848/Y 0.03fF
C37547 AND2X1_LOC_721/Y AND2X1_LOC_848/Y 0.03fF
C41032 AND2X1_LOC_710/Y AND2X1_LOC_848/Y 0.10fF
C43094 AND2X1_LOC_848/Y AND2X1_LOC_789/Y 0.08fF
C46744 AND2X1_LOC_711/a_8_24# AND2X1_LOC_848/Y 0.04fF
C52843 AND2X1_LOC_711/Y AND2X1_LOC_848/Y 0.18fF
C55185 AND2X1_LOC_346/a_8_24# AND2X1_LOC_848/Y 0.04fF
C56877 AND2X1_LOC_848/Y VSS 0.16fF
C26200 OR2X1_LOC_612/Y AND2X1_LOC_647/a_8_24# 0.23fF
C30816 VDD OR2X1_LOC_612/Y 0.12fF
C42414 AND2X1_LOC_852/Y OR2X1_LOC_612/Y 0.10fF
C56750 OR2X1_LOC_612/Y VSS -0.10fF
C5161 AND2X1_LOC_67/Y OR2X1_LOC_202/a_36_216# 0.03fF
C6727 OR2X1_LOC_493/B AND2X1_LOC_67/Y 0.16fF
C12319 OR2X1_LOC_493/a_8_216# AND2X1_LOC_67/Y 0.15fF
C12514 AND2X1_LOC_67/Y OR2X1_LOC_493/Y 0.10fF
C20391 VDD AND2X1_LOC_67/Y 0.27fF
C22771 OR2X1_LOC_241/Y AND2X1_LOC_67/Y 0.12fF
C29739 AND2X1_LOC_67/Y OR2X1_LOC_737/A 0.02fF
C43795 OR2X1_LOC_493/A AND2X1_LOC_67/Y 0.18fF
C46880 AND2X1_LOC_67/Y OR2X1_LOC_805/A 0.03fF
C50398 AND2X1_LOC_67/Y OR2X1_LOC_202/a_8_216# 0.02fF
C57055 AND2X1_LOC_67/Y VSS 0.33fF
C1446 OR2X1_LOC_539/Y OR2X1_LOC_854/A 0.20fF
C1710 OR2X1_LOC_854/A OR2X1_LOC_319/Y 0.33fF
C17955 OR2X1_LOC_538/A OR2X1_LOC_854/A 0.02fF
C22738 OR2X1_LOC_354/A OR2X1_LOC_854/A 0.29fF
C23326 OR2X1_LOC_854/A OR2X1_LOC_567/a_8_216# 0.06fF
C26487 OR2X1_LOC_703/B OR2X1_LOC_854/A 0.01fF
C28070 OR2X1_LOC_175/Y OR2X1_LOC_854/A 0.06fF
C29001 OR2X1_LOC_620/Y OR2X1_LOC_854/A 0.02fF
C34246 OR2X1_LOC_854/A OR2X1_LOC_568/A 0.99fF
C36982 OR2X1_LOC_840/A OR2X1_LOC_854/A 0.05fF
C50020 OR2X1_LOC_449/B OR2X1_LOC_854/A 0.03fF
C56397 OR2X1_LOC_854/A VSS 0.38fF
C2705 OR2X1_LOC_207/B OR2X1_LOC_199/B 0.72fF
C47835 OR2X1_LOC_199/a_8_216# OR2X1_LOC_199/B 0.01fF
C56332 OR2X1_LOC_199/B VSS 0.10fF
C1520 OR2X1_LOC_139/A OR2X1_LOC_856/B 0.07fF
C1537 OR2X1_LOC_139/A OR2X1_LOC_793/a_8_216# 0.40fF
C1944 OR2X1_LOC_139/A OR2X1_LOC_175/B 0.27fF
C2413 OR2X1_LOC_139/A OR2X1_LOC_624/A 0.17fF
C3648 OR2X1_LOC_508/A OR2X1_LOC_139/A 0.10fF
C8766 OR2X1_LOC_139/A OR2X1_LOC_475/a_8_216# 0.25fF
C8793 OR2X1_LOC_139/A OR2X1_LOC_539/Y 0.03fF
C10028 OR2X1_LOC_139/A OR2X1_LOC_61/Y 0.07fF
C11339 OR2X1_LOC_139/A OR2X1_LOC_137/Y 0.07fF
C12585 OR2X1_LOC_139/A OR2X1_LOC_805/A 0.10fF
C13681 OR2X1_LOC_139/A OR2X1_LOC_228/Y 0.07fF
C14430 OR2X1_LOC_139/A OR2X1_LOC_244/A 0.02fF
C16871 OR2X1_LOC_139/A OR2X1_LOC_139/a_8_216# 0.08fF
C18820 OR2X1_LOC_139/A OR2X1_LOC_140/Y 0.01fF
C18886 OR2X1_LOC_139/A OR2X1_LOC_390/A 0.06fF
C19692 OR2X1_LOC_139/A OR2X1_LOC_508/Y 0.36fF
C20321 OR2X1_LOC_139/A OR2X1_LOC_473/Y 0.05fF
C21982 OR2X1_LOC_139/A OR2X1_LOC_510/Y 0.11fF
C22886 OR2X1_LOC_139/A OR2X1_LOC_793/A 0.08fF
C23418 OR2X1_LOC_139/A OR2X1_LOC_786/Y 0.23fF
C23694 OR2X1_LOC_139/A OR2X1_LOC_204/Y 0.07fF
C25290 OR2X1_LOC_139/A OR2X1_LOC_538/A 0.03fF
C26559 OR2X1_LOC_139/A OR2X1_LOC_653/Y 0.39fF
C27893 OR2X1_LOC_139/A OR2X1_LOC_141/B 0.01fF
C28999 OR2X1_LOC_139/A OR2X1_LOC_390/a_8_216# 0.05fF
C29140 OR2X1_LOC_139/A OR2X1_LOC_203/Y 0.10fF
C34943 OR2X1_LOC_97/A OR2X1_LOC_139/A 0.03fF
C35015 OR2X1_LOC_139/A OR2X1_LOC_475/B 5.07fF
C35302 OR2X1_LOC_175/Y OR2X1_LOC_139/A 0.12fF
C35356 OR2X1_LOC_124/A OR2X1_LOC_139/A 0.03fF
C36495 OR2X1_LOC_139/A OR2X1_LOC_560/A 0.05fF
C36762 OR2X1_LOC_139/A OR2X1_LOC_476/a_8_216# 0.06fF
C40773 OR2X1_LOC_139/A OR2X1_LOC_174/Y 0.03fF
C42187 OR2X1_LOC_139/A VDD 0.86fF
C44833 OR2X1_LOC_139/A OR2X1_LOC_216/A 0.52fF
C47163 OR2X1_LOC_702/A OR2X1_LOC_139/A 0.02fF
C47207 OR2X1_LOC_139/A OR2X1_LOC_476/B 0.03fF
C47903 OR2X1_LOC_139/A OR2X1_LOC_641/A 0.02fF
C48837 OR2X1_LOC_139/A OR2X1_LOC_643/A 0.07fF
C48841 OR2X1_LOC_139/A OR2X1_LOC_124/Y 0.02fF
C52128 OR2X1_LOC_139/A OR2X1_LOC_244/B 0.01fF
C53854 OR2X1_LOC_139/A OR2X1_LOC_474/Y 0.24fF
C55268 OR2X1_LOC_139/A OR2X1_LOC_720/B 0.60fF
C55732 OR2X1_LOC_139/A OR2X1_LOC_506/B 0.03fF
C57849 OR2X1_LOC_139/A VSS -3.02fF
C5456 OR2X1_LOC_472/A OR2X1_LOC_852/B 0.05fF
C13871 OR2X1_LOC_852/a_8_216# OR2X1_LOC_852/B 0.39fF
C54519 OR2X1_LOC_852/B OR2X1_LOC_852/A 0.12fF
C55162 VDD OR2X1_LOC_852/B -0.00fF
C57416 OR2X1_LOC_852/B VSS 0.17fF
C1493 OR2X1_LOC_447/Y OR2X1_LOC_779/Y 0.10fF
C2462 OR2X1_LOC_447/Y OR2X1_LOC_712/B 0.03fF
C5438 OR2X1_LOC_447/Y OR2X1_LOC_713/A 0.65fF
C6978 OR2X1_LOC_447/Y OR2X1_LOC_783/a_8_216# 0.02fF
C10721 OR2X1_LOC_447/Y OR2X1_LOC_714/Y 0.04fF
C11193 OR2X1_LOC_447/Y OR2X1_LOC_705/Y 0.09fF
C12354 VDD OR2X1_LOC_447/Y 0.08fF
C12540 OR2X1_LOC_447/Y OR2X1_LOC_783/a_36_216# 0.02fF
C16700 OR2X1_LOC_447/Y OR2X1_LOC_713/a_8_216# 0.03fF
C17954 OR2X1_LOC_447/Y OR2X1_LOC_449/A 0.07fF
C18844 OR2X1_LOC_447/Y OR2X1_LOC_778/Y 0.03fF
C20746 OR2X1_LOC_447/Y OR2X1_LOC_714/a_8_216# 0.01fF
C31879 OR2X1_LOC_447/Y OR2X1_LOC_784/Y 0.07fF
C39614 OR2X1_LOC_447/Y OR2X1_LOC_446/Y 1.48fF
C41419 OR2X1_LOC_447/Y OR2X1_LOC_714/A 0.01fF
C42258 OR2X1_LOC_447/Y OR2X1_LOC_724/A 0.24fF
C43499 OR2X1_LOC_447/Y OR2X1_LOC_783/A 0.15fF
C43651 OR2X1_LOC_447/Y OR2X1_LOC_308/Y 0.02fF
C45224 OR2X1_LOC_447/Y OR2X1_LOC_454/a_8_216# 0.02fF
C52752 OR2X1_LOC_447/Y OR2X1_LOC_713/a_36_216# 0.02fF
C53750 OR2X1_LOC_448/Y OR2X1_LOC_447/Y 0.46fF
C57384 OR2X1_LOC_447/Y VSS 0.48fF
C3247 OR2X1_LOC_506/Y OR2X1_LOC_721/Y 0.06fF
C9166 OR2X1_LOC_506/Y OR2X1_LOC_242/a_8_216# 0.41fF
C13780 OR2X1_LOC_506/Y OR2X1_LOC_392/B 0.09fF
C18271 OR2X1_LOC_506/Y OR2X1_LOC_241/Y 0.10fF
C25713 OR2X1_LOC_506/Y OR2X1_LOC_244/B 0.10fF
C29282 OR2X1_LOC_506/Y OR2X1_LOC_506/B 0.26fF
C33315 OR2X1_LOC_508/A OR2X1_LOC_506/Y 0.08fF
C52107 OR2X1_LOC_715/B OR2X1_LOC_506/Y 0.10fF
C58017 OR2X1_LOC_506/Y VSS 0.25fF
C1940 OR2X1_LOC_174/A OR2X1_LOC_390/A 0.03fF
C7335 OR2X1_LOC_339/A OR2X1_LOC_390/A 0.07fF
C13050 OR2X1_LOC_653/Y OR2X1_LOC_390/A 0.01fF
C20163 OR2X1_LOC_174/a_8_216# OR2X1_LOC_390/A 0.03fF
C20581 OR2X1_LOC_390/B OR2X1_LOC_390/A 0.23fF
C21883 OR2X1_LOC_175/Y OR2X1_LOC_390/A 0.01fF
C22502 OR2X1_LOC_333/B OR2X1_LOC_390/A 0.09fF
C25653 OR2X1_LOC_174/a_36_216# OR2X1_LOC_390/A 0.01fF
C28637 VDD OR2X1_LOC_390/A 0.21fF
C44876 OR2X1_LOC_624/A OR2X1_LOC_390/A 0.03fF
C55168 OR2X1_LOC_805/A OR2X1_LOC_390/A 0.03fF
C56246 OR2X1_LOC_390/A VSS -0.53fF
C2554 OR2X1_LOC_630/Y OR2X1_LOC_574/A 0.02fF
C8199 OR2X1_LOC_630/Y OR2X1_LOC_493/Y 0.10fF
C10217 OR2X1_LOC_630/Y OR2X1_LOC_778/A 0.01fF
C12516 OR2X1_LOC_630/Y OR2X1_LOC_140/B 0.07fF
C15947 VDD OR2X1_LOC_630/Y 0.37fF
C18023 OR2X1_LOC_630/Y OR2X1_LOC_115/B 0.12fF
C18627 OR2X1_LOC_630/Y OR2X1_LOC_499/a_8_216# 0.01fF
C29044 OR2X1_LOC_630/Y OR2X1_LOC_554/a_8_216# 0.02fF
C29633 OR2X1_LOC_630/Y OR2X1_LOC_500/A 0.92fF
C39316 OR2X1_LOC_630/Y OR2X1_LOC_575/A 0.01fF
C41407 OR2X1_LOC_630/Y OR2X1_LOC_632/a_8_216# 0.04fF
C45677 OR2X1_LOC_630/Y OR2X1_LOC_563/A 0.02fF
C46209 OR2X1_LOC_630/Y OR2X1_LOC_632/Y 0.03fF
C57584 OR2X1_LOC_630/Y VSS 0.22fF
C10745 AND2X1_LOC_147/Y AND2X1_LOC_149/a_8_24# 0.09fF
C14548 OR2X1_LOC_680/Y AND2X1_LOC_147/Y 0.01fF
C35643 AND2X1_LOC_147/Y OR2X1_LOC_679/B 0.34fF
C39393 AND2X1_LOC_658/B AND2X1_LOC_147/Y 0.03fF
C42137 OR2X1_LOC_679/A AND2X1_LOC_147/Y 0.37fF
C46667 AND2X1_LOC_544/Y AND2X1_LOC_147/Y 0.03fF
C49889 AND2X1_LOC_147/Y AND2X1_LOC_624/A 0.15fF
C50677 OR2X1_LOC_524/Y AND2X1_LOC_147/Y 0.03fF
C55851 AND2X1_LOC_147/Y AND2X1_LOC_148/Y 0.01fF
C56237 AND2X1_LOC_728/Y AND2X1_LOC_147/Y 0.83fF
C57168 AND2X1_LOC_147/Y VSS -0.18fF
C350 AND2X1_LOC_727/A AND2X1_LOC_727/B 0.33fF
C4987 AND2X1_LOC_810/A AND2X1_LOC_727/A 3.08fF
C5565 AND2X1_LOC_727/A AND2X1_LOC_653/a_8_24# 0.01fF
C5982 AND2X1_LOC_727/A AND2X1_LOC_652/a_8_24# 0.01fF
C7418 AND2X1_LOC_727/A AND2X1_LOC_810/a_8_24# 0.01fF
C9801 AND2X1_LOC_392/A AND2X1_LOC_727/A 0.03fF
C9875 AND2X1_LOC_354/Y AND2X1_LOC_727/A 0.01fF
C11148 AND2X1_LOC_727/A AND2X1_LOC_661/A 0.03fF
C11215 AND2X1_LOC_727/A AND2X1_LOC_810/Y 0.01fF
C11564 AND2X1_LOC_727/A AND2X1_LOC_653/B 0.01fF
C12969 AND2X1_LOC_727/A AND2X1_LOC_798/A 0.01fF
C13591 AND2X1_LOC_794/B AND2X1_LOC_727/A 0.03fF
C13624 VDD AND2X1_LOC_727/A 0.60fF
C14117 AND2X1_LOC_486/Y AND2X1_LOC_727/A 0.03fF
C17049 AND2X1_LOC_727/A OR2X1_LOC_594/Y 0.01fF
C19229 AND2X1_LOC_727/A AND2X1_LOC_354/B 0.04fF
C21929 AND2X1_LOC_727/A AND2X1_LOC_486/a_8_24# 0.01fF
C24417 AND2X1_LOC_170/B AND2X1_LOC_727/A 0.03fF
C27694 AND2X1_LOC_702/Y AND2X1_LOC_727/A 0.37fF
C28565 OR2X1_LOC_312/Y AND2X1_LOC_727/A 0.03fF
C31763 AND2X1_LOC_727/a_8_24# AND2X1_LOC_727/A -0.00fF
C33181 AND2X1_LOC_715/a_8_24# AND2X1_LOC_727/A 0.01fF
C33506 AND2X1_LOC_535/Y AND2X1_LOC_727/A 0.01fF
C33544 OR2X1_LOC_484/Y AND2X1_LOC_727/A 0.01fF
C35645 AND2X1_LOC_722/A AND2X1_LOC_727/A 0.03fF
C35715 AND2X1_LOC_727/A AND2X1_LOC_854/a_8_24# 0.01fF
C36417 AND2X1_LOC_353/a_8_24# AND2X1_LOC_727/A 0.11fF
C37363 AND2X1_LOC_365/A AND2X1_LOC_727/A 0.03fF
C38087 AND2X1_LOC_388/Y AND2X1_LOC_727/A 0.01fF
C40403 AND2X1_LOC_727/A AND2X1_LOC_856/a_8_24# 0.01fF
C41227 AND2X1_LOC_727/A AND2X1_LOC_856/A 0.01fF
C44603 AND2X1_LOC_567/a_8_24# AND2X1_LOC_727/A 0.01fF
C45169 AND2X1_LOC_337/B AND2X1_LOC_727/A 0.02fF
C45565 AND2X1_LOC_388/a_8_24# AND2X1_LOC_727/A 0.01fF
C45763 AND2X1_LOC_727/A OR2X1_LOC_142/Y 0.07fF
C47660 OR2X1_LOC_176/Y AND2X1_LOC_727/A 0.02fF
C48509 AND2X1_LOC_539/Y AND2X1_LOC_727/A 0.01fF
C49395 AND2X1_LOC_784/Y AND2X1_LOC_727/A 0.02fF
C50258 AND2X1_LOC_568/B AND2X1_LOC_727/A 0.03fF
C51153 AND2X1_LOC_727/A AND2X1_LOC_468/B 0.04fF
C51651 AND2X1_LOC_727/A AND2X1_LOC_863/A 0.17fF
C53735 AND2X1_LOC_354/a_8_24# AND2X1_LOC_727/A 0.01fF
C57193 AND2X1_LOC_727/A VSS -0.65fF
C9787 AND2X1_LOC_712/Y AND2X1_LOC_712/B 0.06fF
C12326 VDD AND2X1_LOC_712/B 0.05fF
C20830 AND2X1_LOC_713/Y AND2X1_LOC_712/B 0.01fF
C33608 AND2X1_LOC_712/B AND2X1_LOC_448/Y 0.41fF
C46759 AND2X1_LOC_712/a_8_24# AND2X1_LOC_712/B 0.09fF
C57561 AND2X1_LOC_712/B VSS 0.19fF
C2144 AND2X1_LOC_638/Y AND2X1_LOC_651/B 0.01fF
C3282 VDD AND2X1_LOC_638/Y -0.00fF
C21630 AND2X1_LOC_638/Y AND2X1_LOC_651/a_8_24# 0.10fF
C57111 AND2X1_LOC_638/Y VSS -0.03fF
C20443 AND2X1_LOC_459/Y AND2X1_LOC_463/a_8_24# 0.09fF
C56905 AND2X1_LOC_459/Y VSS 0.16fF
C5086 AND2X1_LOC_326/B AND2X1_LOC_841/a_8_24# 0.01fF
C10697 AND2X1_LOC_326/B AND2X1_LOC_851/B 0.83fF
C16065 AND2X1_LOC_784/A AND2X1_LOC_326/B 0.05fF
C17353 AND2X1_LOC_211/B AND2X1_LOC_326/B 0.07fF
C25297 AND2X1_LOC_326/B AND2X1_LOC_476/Y 0.02fF
C26980 AND2X1_LOC_392/A AND2X1_LOC_326/B 0.03fF
C30541 AND2X1_LOC_326/B AND2X1_LOC_326/a_8_24# 0.11fF
C30793 VDD AND2X1_LOC_326/B 0.21fF
C36367 AND2X1_LOC_326/B AND2X1_LOC_354/B 0.01fF
C52231 OR2X1_LOC_109/Y AND2X1_LOC_326/B 0.01fF
C57477 AND2X1_LOC_326/B VSS 0.16fF
C3025 OR2X1_LOC_109/Y AND2X1_LOC_374/Y 0.02fF
C5297 AND2X1_LOC_543/Y AND2X1_LOC_374/Y 0.02fF
C9455 AND2X1_LOC_717/B AND2X1_LOC_374/Y 0.13fF
C11787 AND2X1_LOC_374/Y AND2X1_LOC_786/Y 0.02fF
C15179 OR2X1_LOC_177/Y AND2X1_LOC_374/Y 0.01fF
C21994 AND2X1_LOC_564/B AND2X1_LOC_374/Y 1.23fF
C23911 OR2X1_LOC_280/Y AND2X1_LOC_374/Y 0.01fF
C32105 AND2X1_LOC_476/Y AND2X1_LOC_374/Y 0.05fF
C33526 AND2X1_LOC_717/a_8_24# AND2X1_LOC_374/Y 0.10fF
C37625 VDD AND2X1_LOC_374/Y 0.06fF
C41416 AND2X1_LOC_721/Y AND2X1_LOC_374/Y 0.01fF
C52848 OR2X1_LOC_312/Y AND2X1_LOC_374/Y 0.01fF
C56575 AND2X1_LOC_374/Y VSS 0.26fF
C1706 AND2X1_LOC_784/A AND2X1_LOC_168/Y 0.05fF
C24259 OR2X1_LOC_91/Y AND2X1_LOC_168/Y 0.04fF
C28275 AND2X1_LOC_787/A AND2X1_LOC_168/Y 0.01fF
C31342 AND2X1_LOC_716/Y AND2X1_LOC_168/Y 0.51fF
C50496 OR2X1_LOC_176/Y AND2X1_LOC_168/Y 0.09fF
C53091 AND2X1_LOC_168/Y AND2X1_LOC_568/B 0.02fF
C53604 AND2X1_LOC_168/Y AND2X1_LOC_170/a_8_24# 0.09fF
C57886 AND2X1_LOC_168/Y VSS -0.26fF
C7356 AND2X1_LOC_776/Y AND2X1_LOC_786/Y 0.02fF
C9664 AND2X1_LOC_776/Y OR2X1_LOC_238/Y 0.02fF
C17525 AND2X1_LOC_776/Y AND2X1_LOC_564/B 0.18fF
C20121 AND2X1_LOC_776/Y AND2X1_LOC_785/a_8_24# 0.03fF
C26423 AND2X1_LOC_776/Y AND2X1_LOC_785/A 0.02fF
C31900 OR2X1_LOC_516/Y AND2X1_LOC_776/Y 0.12fF
C33258 AND2X1_LOC_776/Y VDD 0.11fF
C33738 AND2X1_LOC_776/Y AND2X1_LOC_486/Y 0.72fF
C36983 AND2X1_LOC_776/Y AND2X1_LOC_721/Y 0.01fF
C58125 AND2X1_LOC_776/Y VSS -0.35fF
C7144 OR2X1_LOC_768/A OR2X1_LOC_673/Y 0.01fF
C10672 OR2X1_LOC_400/A OR2X1_LOC_673/Y 0.01fF
C15281 OR2X1_LOC_673/Y OR2X1_LOC_137/B 0.03fF
C19266 OR2X1_LOC_673/Y OR2X1_LOC_84/A 0.01fF
C23797 OR2X1_LOC_137/a_8_216# OR2X1_LOC_673/Y 0.01fF
C24738 OR2X1_LOC_673/Y AND2X1_LOC_79/Y 0.07fF
C28826 OR2X1_LOC_673/Y OR2X1_LOC_721/Y 0.01fF
C31258 OR2X1_LOC_673/Y OR2X1_LOC_720/Y 0.06fF
C36481 OR2X1_LOC_673/Y OR2X1_LOC_845/a_8_216# 0.01fF
C41486 VDD OR2X1_LOC_673/Y 0.12fF
C41716 OR2X1_LOC_673/Y OR2X1_LOC_845/A 0.04fF
C47769 OR2X1_LOC_673/Y OR2X1_LOC_849/A 0.01fF
C48018 OR2X1_LOC_673/Y OR2X1_LOC_721/a_8_216# 0.01fF
C53424 OR2X1_LOC_673/Y OR2X1_LOC_771/B 0.07fF
C57673 OR2X1_LOC_673/Y VSS 0.37fF
C139 AND2X1_LOC_706/Y AND2X1_LOC_714/a_8_24# 0.02fF
C1943 AND2X1_LOC_706/Y AND2X1_LOC_605/Y 0.23fF
C5648 AND2X1_LOC_706/Y AND2X1_LOC_724/A 0.02fF
C12101 AND2X1_LOC_706/Y AND2X1_LOC_447/Y 0.02fF
C14167 AND2X1_LOC_706/Y OR2X1_LOC_424/Y 0.01fF
C37799 AND2X1_LOC_706/Y OR2X1_LOC_423/Y 0.03fF
C44933 AND2X1_LOC_706/Y AND2X1_LOC_645/A 0.03fF
C45217 AND2X1_LOC_706/Y AND2X1_LOC_703/Y 0.01fF
C47042 AND2X1_LOC_706/Y VDD 0.57fF
C47484 AND2X1_LOC_706/Y AND2X1_LOC_713/a_8_24# 0.01fF
C55515 AND2X1_LOC_706/Y AND2X1_LOC_713/Y 0.02fF
C57923 AND2X1_LOC_706/Y VSS 0.20fF
C6997 AND2X1_LOC_347/B AND2X1_LOC_711/A 0.05fF
C11209 AND2X1_LOC_711/A AND2X1_LOC_792/a_8_24# 0.05fF
C13587 AND2X1_LOC_711/A OR2X1_LOC_258/Y 0.01fF
C39973 AND2X1_LOC_711/A AND2X1_LOC_789/Y 0.02fF
C50855 AND2X1_LOC_711/A OR2X1_LOC_759/Y 0.24fF
C57494 AND2X1_LOC_711/A VSS 0.29fF
C4683 AND2X1_LOC_148/Y AND2X1_LOC_624/A 0.11fF
C6562 AND2X1_LOC_727/Y AND2X1_LOC_624/A 0.03fF
C8895 AND2X1_LOC_508/A AND2X1_LOC_624/A 0.07fF
C9073 AND2X1_LOC_624/A AND2X1_LOC_620/Y 0.23fF
C9634 AND2X1_LOC_564/B AND2X1_LOC_624/A 0.07fF
C12178 AND2X1_LOC_624/A AND2X1_LOC_727/B 0.03fF
C13937 AND2X1_LOC_719/Y AND2X1_LOC_624/A 0.03fF
C15673 AND2X1_LOC_624/A AND2X1_LOC_573/A 0.03fF
C17438 AND2X1_LOC_624/A OR2X1_LOC_239/Y 0.03fF
C18611 AND2X1_LOC_658/A AND2X1_LOC_624/A 0.10fF
C19623 OR2X1_LOC_680/Y AND2X1_LOC_624/A 0.03fF
C19878 AND2X1_LOC_624/A AND2X1_LOC_476/Y 0.07fF
C20454 OR2X1_LOC_665/Y AND2X1_LOC_624/A 6.13fF
C20455 AND2X1_LOC_624/A AND2X1_LOC_474/Y 0.03fF
C22473 AND2X1_LOC_549/Y AND2X1_LOC_624/A 0.11fF
C22489 AND2X1_LOC_500/Y AND2X1_LOC_624/A 0.12fF
C23673 OR2X1_LOC_406/Y AND2X1_LOC_624/A 0.03fF
C24065 OR2X1_LOC_516/Y AND2X1_LOC_624/A 0.07fF
C24685 AND2X1_LOC_859/Y AND2X1_LOC_624/A 0.07fF
C25386 VDD AND2X1_LOC_624/A 0.39fF
C25548 AND2X1_LOC_624/A AND2X1_LOC_624/a_8_24# 0.10fF
C25637 AND2X1_LOC_624/A AND2X1_LOC_624/B 0.45fF
C25931 OR2X1_LOC_666/Y AND2X1_LOC_624/A 0.03fF
C29116 AND2X1_LOC_721/Y AND2X1_LOC_624/A 0.03fF
C29158 OR2X1_LOC_482/Y AND2X1_LOC_624/A 0.15fF
C29606 AND2X1_LOC_508/B AND2X1_LOC_624/A 0.07fF
C29620 AND2X1_LOC_508/a_8_24# AND2X1_LOC_624/A 0.02fF
C31669 AND2X1_LOC_624/A AND2X1_LOC_213/B 0.03fF
C32631 AND2X1_LOC_850/Y AND2X1_LOC_624/A 0.42fF
C33543 AND2X1_LOC_624/A AND2X1_LOC_806/A 0.03fF
C33893 OR2X1_LOC_441/Y AND2X1_LOC_624/A 17.05fF
C35097 AND2X1_LOC_510/A AND2X1_LOC_624/A 0.03fF
C35550 AND2X1_LOC_734/Y AND2X1_LOC_624/A 0.03fF
C41441 OR2X1_LOC_528/Y AND2X1_LOC_624/A 4.47fF
C42596 AND2X1_LOC_624/A AND2X1_LOC_792/Y 0.07fF
C43703 OR2X1_LOC_438/Y AND2X1_LOC_624/A 0.03fF
C44278 OR2X1_LOC_504/Y AND2X1_LOC_624/A 0.13fF
C44496 AND2X1_LOC_658/B AND2X1_LOC_624/A 26.34fF
C47394 OR2X1_LOC_679/A AND2X1_LOC_624/A 0.03fF
C48687 AND2X1_LOC_624/A OR2X1_LOC_615/Y 0.03fF
C49778 AND2X1_LOC_509/Y AND2X1_LOC_624/A 0.03fF
C51764 AND2X1_LOC_544/Y AND2X1_LOC_624/A 0.03fF
C51909 AND2X1_LOC_550/A AND2X1_LOC_624/A 0.03fF
C52708 AND2X1_LOC_675/Y AND2X1_LOC_624/A 0.18fF
C53786 AND2X1_LOC_624/A AND2X1_LOC_793/Y 0.07fF
C55918 AND2X1_LOC_624/A OR2X1_LOC_746/Y 0.14fF
C56913 AND2X1_LOC_624/A VSS 0.48fF
C7650 VDD OR2X1_LOC_243/B 0.02fF
C24834 OR2X1_LOC_243/B OR2X1_LOC_243/a_8_216# 0.05fF
C35772 OR2X1_LOC_243/B OR2X1_LOC_244/A 0.07fF
C57206 OR2X1_LOC_243/B VSS 0.10fF
C52414 VDD OR2X1_LOC_845/A 0.08fF
C56983 OR2X1_LOC_845/A VSS 0.26fF
C5691 OR2X1_LOC_97/A OR2X1_LOC_640/A 0.09fF
C13068 VDD OR2X1_LOC_640/A 0.06fF
C14024 OR2X1_LOC_462/B OR2X1_LOC_640/A 0.02fF
C17864 OR2X1_LOC_476/B OR2X1_LOC_640/A 0.01fF
C19556 OR2X1_LOC_472/A OR2X1_LOC_640/A 0.11fF
C22526 OR2X1_LOC_633/Y OR2X1_LOC_640/A 0.15fF
C33458 OR2X1_LOC_640/a_8_216# OR2X1_LOC_640/A 0.18fF
C51953 OR2X1_LOC_472/a_8_216# OR2X1_LOC_640/A 0.40fF
C57453 OR2X1_LOC_640/A VSS 0.27fF
C1315 OR2X1_LOC_719/Y OR2X1_LOC_553/A 0.01fF
C2040 OR2X1_LOC_190/A OR2X1_LOC_553/A 0.07fF
C2295 OR2X1_LOC_553/A OR2X1_LOC_241/B 0.15fF
C3851 OR2X1_LOC_456/Y OR2X1_LOC_553/A 0.04fF
C6724 OR2X1_LOC_147/B OR2X1_LOC_553/A 0.07fF
C6928 OR2X1_LOC_553/A OR2X1_LOC_318/B 0.02fF
C8993 OR2X1_LOC_445/a_8_216# OR2X1_LOC_553/A 0.04fF
C10624 OR2X1_LOC_553/B OR2X1_LOC_553/A 0.10fF
C14902 OR2X1_LOC_465/a_8_216# OR2X1_LOC_553/A 0.04fF
C20445 OR2X1_LOC_76/Y OR2X1_LOC_553/A 0.06fF
C20900 OR2X1_LOC_553/A OR2X1_LOC_553/a_8_216# 0.04fF
C20933 OR2X1_LOC_719/A OR2X1_LOC_553/A 0.21fF
C21005 OR2X1_LOC_553/A OR2X1_LOC_675/Y 0.01fF
C23408 OR2X1_LOC_76/B OR2X1_LOC_553/A 0.01fF
C23988 OR2X1_LOC_76/a_8_216# OR2X1_LOC_553/A 0.05fF
C24177 VDD OR2X1_LOC_553/A 0.77fF
C25925 OR2X1_LOC_455/a_8_216# OR2X1_LOC_553/A -0.03fF
C26808 OR2X1_LOC_675/a_8_216# OR2X1_LOC_553/A 0.04fF
C27985 OR2X1_LOC_190/B OR2X1_LOC_553/A 0.17fF
C30246 OR2X1_LOC_440/A OR2X1_LOC_553/A 0.01fF
C31052 OR2X1_LOC_455/A OR2X1_LOC_553/A 0.03fF
C31287 OR2X1_LOC_553/A OR2X1_LOC_719/B 0.02fF
C31315 OR2X1_LOC_542/B OR2X1_LOC_553/A 0.07fF
C31423 OR2X1_LOC_455/a_36_216# OR2X1_LOC_553/A 0.01fF
C36727 OR2X1_LOC_553/A OR2X1_LOC_719/a_8_216# 0.03fF
C36883 OR2X1_LOC_465/B OR2X1_LOC_553/A 0.02fF
C42443 OR2X1_LOC_465/Y OR2X1_LOC_553/A 0.03fF
C45553 OR2X1_LOC_675/A OR2X1_LOC_553/A 0.01fF
C50705 OR2X1_LOC_805/A OR2X1_LOC_553/A 0.94fF
C52010 OR2X1_LOC_76/A OR2X1_LOC_553/A 0.05fF
C55178 OR2X1_LOC_486/Y OR2X1_LOC_553/A 0.07fF
C56591 OR2X1_LOC_553/A VSS -1.03fF
C5338 VDD OR2X1_LOC_633/Y 0.25fF
C24696 OR2X1_LOC_633/Y OR2X1_LOC_633/B 0.16fF
C25886 OR2X1_LOC_633/Y OR2X1_LOC_640/a_8_216# 0.04fF
C31025 OR2X1_LOC_633/Y OR2X1_LOC_647/B 0.07fF
C54271 OR2X1_LOC_97/A OR2X1_LOC_633/Y 0.91fF
C57770 OR2X1_LOC_633/Y VSS 0.02fF
C32008 VDD OR2X1_LOC_784/B -0.00fF
C38488 OR2X1_LOC_778/Y OR2X1_LOC_784/B 0.12fF
C55258 OR2X1_LOC_784/a_8_216# OR2X1_LOC_784/B 0.39fF
C56614 OR2X1_LOC_784/B VSS 0.17fF
C24899 OR2X1_LOC_549/Y OR2X1_LOC_565/a_8_216# 0.07fF
C35668 VDD OR2X1_LOC_549/Y 0.23fF
C43459 OR2X1_LOC_563/B OR2X1_LOC_549/Y 0.17fF
C52404 OR2X1_LOC_565/A OR2X1_LOC_549/Y 0.04fF
C56487 OR2X1_LOC_549/Y VSS 0.35fF
C14263 OR2X1_LOC_392/B OR2X1_LOC_392/A 0.05fF
C24387 OR2X1_LOC_392/A OR2X1_LOC_561/B 0.02fF
C35600 OR2X1_LOC_774/Y OR2X1_LOC_392/A 0.01fF
C56704 OR2X1_LOC_392/A VSS 0.19fF
C1662 VDD AND2X1_LOC_390/B 1.08fF
C6917 AND2X1_LOC_390/B AND2X1_LOC_169/a_8_24# 0.02fF
C9520 AND2X1_LOC_390/B OR2X1_LOC_311/Y 0.06fF
C14508 AND2X1_LOC_356/a_8_24# AND2X1_LOC_390/B 0.01fF
C16637 AND2X1_LOC_390/B OR2X1_LOC_312/Y 0.02fF
C21668 AND2X1_LOC_535/Y AND2X1_LOC_390/B 0.02fF
C22232 AND2X1_LOC_390/B AND2X1_LOC_336/a_8_24# 0.02fF
C25472 OR2X1_LOC_166/Y AND2X1_LOC_390/B 0.02fF
C25538 AND2X1_LOC_365/A AND2X1_LOC_390/B 0.02fF
C26258 AND2X1_LOC_388/Y AND2X1_LOC_390/B 0.07fF
C31318 AND2X1_LOC_390/B AND2X1_LOC_774/A 0.10fF
C33167 AND2X1_LOC_390/B AND2X1_LOC_337/B 0.02fF
C35515 OR2X1_LOC_533/Y AND2X1_LOC_390/B 0.01fF
C36333 AND2X1_LOC_539/Y AND2X1_LOC_390/B 0.02fF
C42837 AND2X1_LOC_390/a_8_24# AND2X1_LOC_390/B 0.05fF
C43841 AND2X1_LOC_356/B AND2X1_LOC_390/B 0.01fF
C46561 AND2X1_LOC_390/B OR2X1_LOC_599/Y 0.08fF
C52050 AND2X1_LOC_390/B OR2X1_LOC_167/Y 0.02fF
C53526 AND2X1_LOC_715/Y AND2X1_LOC_390/B 0.10fF
C53989 AND2X1_LOC_392/A AND2X1_LOC_390/B 0.02fF
C54053 AND2X1_LOC_354/Y AND2X1_LOC_390/B 0.01fF
C54802 AND2X1_LOC_390/B OR2X1_LOC_13/Y 0.16fF
C55849 AND2X1_LOC_390/B AND2X1_LOC_645/A 0.53fF
C57598 AND2X1_LOC_390/B VSS 0.02fF
C24097 OR2X1_LOC_597/Y OR2X1_LOC_599/Y 0.04fF
C35039 OR2X1_LOC_597/Y AND2X1_LOC_644/a_8_24# 0.23fF
C35238 VDD OR2X1_LOC_597/Y 0.12fF
C56917 OR2X1_LOC_597/Y VSS -0.14fF
C2070 AND2X1_LOC_535/Y AND2X1_LOC_356/B 0.01fF
C2673 AND2X1_LOC_356/B AND2X1_LOC_336/a_8_24# 0.01fF
C5949 AND2X1_LOC_356/B AND2X1_LOC_365/A 0.01fF
C13713 AND2X1_LOC_356/B AND2X1_LOC_337/B 0.01fF
C16858 AND2X1_LOC_539/Y AND2X1_LOC_356/B 0.55fF
C38061 VDD AND2X1_LOC_356/B 0.07fF
C46039 AND2X1_LOC_356/B OR2X1_LOC_311/Y 0.01fF
C49106 AND2X1_LOC_356/B AND2X1_LOC_170/B 0.82fF
C51121 AND2X1_LOC_356/B AND2X1_LOC_356/a_8_24# 0.09fF
C53268 AND2X1_LOC_356/B OR2X1_LOC_312/Y 0.03fF
C57660 AND2X1_LOC_356/B VSS 0.16fF
C8103 OR2X1_LOC_504/Y OR2X1_LOC_505/Y 0.01fF
C8113 OR2X1_LOC_504/Y AND2X1_LOC_658/A 0.03fF
C13642 OR2X1_LOC_504/Y AND2X1_LOC_507/a_8_24# 0.01fF
C14907 VDD OR2X1_LOC_504/Y 0.12fF
C19157 OR2X1_LOC_504/Y AND2X1_LOC_508/B 0.01fF
C22237 OR2X1_LOC_504/Y AND2X1_LOC_850/Y 0.18fF
C23120 OR2X1_LOC_504/Y AND2X1_LOC_806/A 0.03fF
C30993 OR2X1_LOC_528/Y OR2X1_LOC_504/Y 0.04fF
C33674 AND2X1_LOC_711/Y OR2X1_LOC_504/Y 0.03fF
C33954 AND2X1_LOC_658/B OR2X1_LOC_504/Y 0.15fF
C57429 OR2X1_LOC_504/Y VSS 0.06fF
C520 OR2X1_LOC_524/Y OR2X1_LOC_746/Y 0.03fF
C26420 VDD OR2X1_LOC_746/Y 0.08fF
C40132 OR2X1_LOC_745/Y OR2X1_LOC_746/Y 0.09fF
C45589 AND2X1_LOC_658/B OR2X1_LOC_746/Y 0.03fF
C52823 AND2X1_LOC_544/Y OR2X1_LOC_746/Y 0.03fF
C56390 OR2X1_LOC_746/Y VSS 0.18fF
C10983 AND2X1_LOC_347/B OR2X1_LOC_258/Y 0.01fF
C31923 OR2X1_LOC_295/Y OR2X1_LOC_258/Y 0.21fF
C32279 AND2X1_LOC_259/Y OR2X1_LOC_258/Y 0.01fF
C34730 VDD OR2X1_LOC_258/Y 0.12fF
C39415 AND2X1_LOC_191/B OR2X1_LOC_258/Y 0.03fF
C40854 OR2X1_LOC_258/Y OR2X1_LOC_257/Y 0.04fF
C48985 OR2X1_LOC_292/Y OR2X1_LOC_258/Y 0.03fF
C52099 OR2X1_LOC_258/Y AND2X1_LOC_259/a_8_24# 0.05fF
C56109 AND2X1_LOC_346/a_8_24# OR2X1_LOC_258/Y 0.01fF
C56997 OR2X1_LOC_258/Y VSS -0.08fF
C41762 VDD OR2X1_LOC_158/Y 0.12fF
C42049 OR2X1_LOC_158/Y OR2X1_LOC_163/Y 0.09fF
C42620 OR2X1_LOC_158/Y AND2X1_LOC_210/a_8_24# 0.23fF
C56606 OR2X1_LOC_158/Y VSS -0.07fF
C7514 OR2X1_LOC_438/Y AND2X1_LOC_658/A 0.11fF
C8785 OR2X1_LOC_438/Y AND2X1_LOC_476/Y 0.02fF
C14322 OR2X1_LOC_438/Y VDD 0.10fF
C24550 OR2X1_LOC_438/Y AND2X1_LOC_734/Y 0.03fF
C25681 OR2X1_LOC_438/Y AND2X1_LOC_439/a_8_24# 0.01fF
C26389 OR2X1_LOC_438/Y AND2X1_LOC_675/A 0.01fF
C33356 AND2X1_LOC_658/B OR2X1_LOC_438/Y 0.14fF
C35021 OR2X1_LOC_438/Y OR2X1_LOC_373/Y 0.33fF
C38024 OR2X1_LOC_438/Y AND2X1_LOC_544/a_8_24# 0.01fF
C40482 AND2X1_LOC_544/Y OR2X1_LOC_438/Y 0.01fF
C40628 OR2X1_LOC_438/Y AND2X1_LOC_550/A 0.04fF
C44480 OR2X1_LOC_438/Y OR2X1_LOC_524/Y 0.08fF
C47973 OR2X1_LOC_177/Y OR2X1_LOC_438/Y 0.41fF
C57867 OR2X1_LOC_438/Y VSS 0.29fF
C1914 VDD OR2X1_LOC_604/Y 0.06fF
C13022 AND2X1_LOC_605/Y OR2X1_LOC_604/Y 0.80fF
C18900 OR2X1_LOC_604/Y AND2X1_LOC_605/a_8_24# 0.01fF
C29993 AND2X1_LOC_452/Y OR2X1_LOC_604/Y 0.05fF
C56636 OR2X1_LOC_604/Y VSS 0.02fF
C330 VDD OR2X1_LOC_498/Y 0.18fF
C18551 AND2X1_LOC_574/Y OR2X1_LOC_498/Y 0.06fF
C51564 OR2X1_LOC_498/Y AND2X1_LOC_474/Y 0.12fF
C53577 AND2X1_LOC_500/Y OR2X1_LOC_498/Y 0.14fF
C57375 OR2X1_LOC_498/Y VSS 0.16fF
C7448 OR2X1_LOC_674/Y AND2X1_LOC_675/a_8_24# 0.01fF
C15309 OR2X1_LOC_674/Y AND2X1_LOC_499/a_8_24# 0.24fF
C20095 OR2X1_LOC_495/Y OR2X1_LOC_674/Y 0.24fF
C20897 OR2X1_LOC_674/Y AND2X1_LOC_500/B 0.01fF
C23489 AND2X1_LOC_675/Y OR2X1_LOC_674/Y 0.15fF
C28374 OR2X1_LOC_674/Y OR2X1_LOC_142/Y 0.03fF
C31929 OR2X1_LOC_496/Y OR2X1_LOC_674/Y 0.02fF
C51029 OR2X1_LOC_516/Y OR2X1_LOC_674/Y 0.12fF
C52410 VDD OR2X1_LOC_674/Y 0.19fF
C56222 OR2X1_LOC_482/Y OR2X1_LOC_674/Y 0.01fF
C57009 OR2X1_LOC_674/Y VSS 0.12fF
C3109 AND2X1_LOC_656/Y OR2X1_LOC_118/Y 0.01fF
C3243 OR2X1_LOC_118/Y AND2X1_LOC_772/Y 0.01fF
C8832 OR2X1_LOC_118/Y AND2X1_LOC_243/Y 0.04fF
C12172 AND2X1_LOC_340/Y OR2X1_LOC_118/Y 0.01fF
C13314 OR2X1_LOC_118/Y AND2X1_LOC_845/Y 0.01fF
C13781 OR2X1_LOC_118/Y OR2X1_LOC_88/Y 1.25fF
C14203 OR2X1_LOC_118/Y AND2X1_LOC_216/A 0.02fF
C18699 OR2X1_LOC_118/Y AND2X1_LOC_573/A 0.04fF
C19718 OR2X1_LOC_118/Y AND2X1_LOC_647/Y 0.02fF
C19886 AND2X1_LOC_340/a_8_24# OR2X1_LOC_118/Y 0.01fF
C22629 AND2X1_LOC_554/B OR2X1_LOC_118/Y 0.61fF
C24539 AND2X1_LOC_392/A OR2X1_LOC_118/Y 0.10fF
C28072 OR2X1_LOC_131/Y OR2X1_LOC_118/Y 0.01fF
C28353 VDD OR2X1_LOC_118/Y 0.38fF
C32668 OR2X1_LOC_117/Y OR2X1_LOC_118/Y 0.03fF
C36178 OR2X1_LOC_118/Y AND2X1_LOC_656/a_8_24# 0.01fF
C39065 AND2X1_LOC_140/a_8_24# OR2X1_LOC_118/Y 0.01fF
C44660 AND2X1_LOC_141/B OR2X1_LOC_118/Y 0.01fF
C49437 AND2X1_LOC_123/a_8_24# OR2X1_LOC_118/Y 0.11fF
C56924 OR2X1_LOC_118/Y VSS 0.23fF
C13837 VDD OR2X1_LOC_821/Y 0.12fF
C35649 OR2X1_LOC_821/Y OR2X1_LOC_813/Y 0.74fF
C53413 OR2X1_LOC_821/Y OR2X1_LOC_822/Y 0.21fF
C57800 OR2X1_LOC_821/Y VSS -0.22fF
C2787 OR2X1_LOC_177/Y AND2X1_LOC_778/Y 0.12fF
C5598 OR2X1_LOC_177/Y OR2X1_LOC_142/Y 0.03fF
C8277 OR2X1_LOC_177/Y AND2X1_LOC_552/a_8_24# 0.01fF
C8351 OR2X1_LOC_177/Y AND2X1_LOC_471/Y 0.03fF
C13787 OR2X1_LOC_177/Y AND2X1_LOC_564/B 0.01fF
C14764 OR2X1_LOC_177/Y AND2X1_LOC_784/A 0.02fF
C18030 OR2X1_LOC_177/Y AND2X1_LOC_719/Y 0.03fF
C22747 AND2X1_LOC_785/A OR2X1_LOC_177/Y 0.01fF
C22831 OR2X1_LOC_177/Y AND2X1_LOC_658/A 0.03fF
C24039 OR2X1_LOC_177/Y AND2X1_LOC_476/Y 0.04fF
C28173 OR2X1_LOC_516/Y OR2X1_LOC_177/Y 0.03fF
C29499 OR2X1_LOC_177/Y VDD 0.41fF
C29960 OR2X1_LOC_177/Y AND2X1_LOC_486/Y 0.03fF
C37146 OR2X1_LOC_91/Y OR2X1_LOC_177/Y 0.04fF
C39674 OR2X1_LOC_177/Y AND2X1_LOC_734/Y 0.03fF
C40812 OR2X1_LOC_177/Y AND2X1_LOC_439/a_8_24# 0.01fF
C41293 OR2X1_LOC_177/Y AND2X1_LOC_787/A 0.63fF
C41570 OR2X1_LOC_177/Y AND2X1_LOC_675/A -0.00fF
C44423 OR2X1_LOC_177/Y AND2X1_LOC_716/Y 0.02fF
C44498 OR2X1_LOC_177/Y OR2X1_LOC_312/Y 0.92fF
C46572 OR2X1_LOC_177/Y AND2X1_LOC_552/A 0.01fF
C48473 AND2X1_LOC_775/a_8_24# OR2X1_LOC_177/Y 0.01fF
C50452 OR2X1_LOC_177/Y OR2X1_LOC_373/Y 0.17fF
C50956 OR2X1_LOC_177/Y OR2X1_LOC_109/Y 0.60fF
C53462 OR2X1_LOC_177/Y AND2X1_LOC_544/a_8_24# 0.01fF
C55057 OR2X1_LOC_177/Y AND2X1_LOC_180/a_8_24# 0.11fF
C55558 OR2X1_LOC_177/Y AND2X1_LOC_717/Y 0.03fF
C55914 OR2X1_LOC_177/Y AND2X1_LOC_544/Y 0.80fF
C56023 OR2X1_LOC_177/Y AND2X1_LOC_550/A 0.04fF
C58053 OR2X1_LOC_177/Y VSS 0.16fF
C2362 AND2X1_LOC_401/Y OR2X1_LOC_397/Y 0.01fF
C7862 AND2X1_LOC_402/a_8_24# OR2X1_LOC_397/Y 0.03fF
C37476 VDD OR2X1_LOC_397/Y 0.12fF
C56385 OR2X1_LOC_397/Y VSS 0.07fF
C4936 OR2X1_LOC_39/Y OR2X1_LOC_16/Y 0.05fF
C39297 VDD OR2X1_LOC_16/Y 0.06fF
C56533 OR2X1_LOC_16/Y VSS 0.22fF
C15866 VDD OR2X1_LOC_767/Y 0.12fF
C46938 OR2X1_LOC_767/Y AND2X1_LOC_772/Y 0.01fF
C52477 OR2X1_LOC_767/Y AND2X1_LOC_773/a_8_24# 0.23fF
C56273 OR2X1_LOC_767/Y VSS 0.06fF
C13805 OR2X1_LOC_262/Y OR2X1_LOC_88/Y 0.01fF
C17930 OR2X1_LOC_88/Y AND2X1_LOC_243/Y 0.01fF
C21373 AND2X1_LOC_340/Y OR2X1_LOC_88/Y 0.84fF
C27754 AND2X1_LOC_573/A OR2X1_LOC_88/Y 0.02fF
C28747 AND2X1_LOC_647/Y OR2X1_LOC_88/Y 0.35fF
C28961 AND2X1_LOC_340/a_8_24# OR2X1_LOC_88/Y 0.01fF
C37399 VDD OR2X1_LOC_88/Y 0.46fF
C37576 OR2X1_LOC_88/Y OR2X1_LOC_67/Y 0.03fF
C56817 OR2X1_LOC_88/Y VSS 0.31fF
C8282 OR2X1_LOC_665/Y AND2X1_LOC_792/Y 0.02fF
C14208 OR2X1_LOC_665/Y OR2X1_LOC_615/Y 0.03fF
C19302 OR2X1_LOC_665/Y AND2X1_LOC_793/Y 0.01fF
C30685 OR2X1_LOC_665/Y AND2X1_LOC_620/Y 3.56fF
C40178 OR2X1_LOC_665/Y AND2X1_LOC_658/A 0.03fF
C46433 OR2X1_LOC_665/Y AND2X1_LOC_859/Y 0.04fF
C47220 VDD OR2X1_LOC_665/Y 0.32fF
C47453 OR2X1_LOC_665/Y AND2X1_LOC_624/B 0.07fF
C47800 OR2X1_LOC_665/Y OR2X1_LOC_666/Y 0.06fF
C51015 OR2X1_LOC_482/Y OR2X1_LOC_665/Y 0.62fF
C57564 OR2X1_LOC_665/Y VSS 0.01fF
C4018 VDD OR2X1_LOC_171/Y 0.27fF
C5751 AND2X1_LOC_640/Y OR2X1_LOC_171/Y 0.02fF
C10781 AND2X1_LOC_338/Y OR2X1_LOC_171/Y 0.16fF
C11337 AND2X1_LOC_641/Y OR2X1_LOC_171/Y 0.13fF
C15543 AND2X1_LOC_852/Y OR2X1_LOC_171/Y 0.02fF
C25255 AND2X1_LOC_334/Y OR2X1_LOC_171/Y 0.02fF
C27738 AND2X1_LOC_231/Y OR2X1_LOC_171/Y 0.10fF
C36207 AND2X1_LOC_338/a_8_24# OR2X1_LOC_171/Y 0.01fF
C36254 AND2X1_LOC_174/a_8_24# OR2X1_LOC_171/Y 0.09fF
C37941 OR2X1_LOC_265/Y OR2X1_LOC_171/Y 0.07fF
C43992 AND2X1_LOC_228/Y OR2X1_LOC_171/Y 0.28fF
C45514 OR2X1_LOC_171/Y OR2X1_LOC_172/Y 0.01fF
C46650 AND2X1_LOC_211/B OR2X1_LOC_171/Y 0.74fF
C56429 OR2X1_LOC_171/Y VSS 0.11fF
C9908 VDD OR2X1_LOC_745/Y 0.12fF
C45806 OR2X1_LOC_745/Y AND2X1_LOC_781/a_8_24# 0.23fF
C56391 OR2X1_LOC_745/Y VSS -0.14fF
C5290 AND2X1_LOC_786/a_8_24# OR2X1_LOC_265/Y 0.03fF
C5591 OR2X1_LOC_75/Y OR2X1_LOC_265/Y 0.15fF
C6338 OR2X1_LOC_262/Y OR2X1_LOC_265/Y 0.02fF
C10203 AND2X1_LOC_76/a_8_24# OR2X1_LOC_265/Y 0.02fF
C11088 AND2X1_LOC_175/a_8_24# OR2X1_LOC_265/Y 0.01fF
C11899 AND2X1_LOC_175/B OR2X1_LOC_265/Y 0.01fF
C13917 AND2X1_LOC_340/Y OR2X1_LOC_265/Y 0.07fF
C14074 AND2X1_LOC_228/Y OR2X1_LOC_265/Y 0.01fF
C15667 AND2X1_LOC_76/Y OR2X1_LOC_265/Y 0.03fF
C16592 AND2X1_LOC_211/B OR2X1_LOC_265/Y 0.19fF
C24012 OR2X1_LOC_265/Y OR2X1_LOC_72/Y 0.52fF
C30041 VDD OR2X1_LOC_265/Y 0.67fF
C31878 OR2X1_LOC_416/Y OR2X1_LOC_265/Y 0.03fF
C37341 AND2X1_LOC_641/Y OR2X1_LOC_265/Y 0.02fF
C44856 AND2X1_LOC_84/Y OR2X1_LOC_265/Y 0.05fF
C47577 OR2X1_LOC_79/Y OR2X1_LOC_265/Y 0.03fF
C49113 AND2X1_LOC_641/a_8_24# OR2X1_LOC_265/Y 0.07fF
C53889 AND2X1_LOC_231/Y OR2X1_LOC_265/Y 0.08fF
C55286 OR2X1_LOC_74/Y OR2X1_LOC_265/Y 0.02fF
C55877 AND2X1_LOC_476/A OR2X1_LOC_265/Y 0.07fF
C56230 OR2X1_LOC_173/Y OR2X1_LOC_265/Y 0.05fF
C56509 OR2X1_LOC_265/Y VSS 0.13fF
C4481 VDD OR2X1_LOC_441/Y 0.48fF
C10863 OR2X1_LOC_441/Y AND2X1_LOC_213/B 0.03fF
C14770 AND2X1_LOC_734/Y OR2X1_LOC_441/Y 0.17fF
C23700 AND2X1_LOC_658/B OR2X1_LOC_441/Y 0.23fF
C26370 OR2X1_LOC_441/Y OR2X1_LOC_679/A 0.03fF
C30752 AND2X1_LOC_544/Y OR2X1_LOC_441/Y 0.03fF
C30921 AND2X1_LOC_550/A OR2X1_LOC_441/Y 0.03fF
C32026 OR2X1_LOC_441/Y AND2X1_LOC_443/a_8_24# 0.01fF
C34640 OR2X1_LOC_524/Y OR2X1_LOC_441/Y 0.09fF
C39732 OR2X1_LOC_441/Y AND2X1_LOC_148/a_8_24# 0.07fF
C41777 AND2X1_LOC_727/Y OR2X1_LOC_441/Y 0.03fF
C47532 OR2X1_LOC_441/Y AND2X1_LOC_727/B 0.03fF
C53904 OR2X1_LOC_441/Y AND2X1_LOC_658/A 0.03fF
C54857 OR2X1_LOC_680/Y OR2X1_LOC_441/Y 0.03fF
C57500 OR2X1_LOC_441/Y VSS 0.33fF
C14108 OR2X1_LOC_166/Y OR2X1_LOC_167/Y 0.20fF
C34726 OR2X1_LOC_166/Y OR2X1_LOC_312/Y 0.09fF
C39678 OR2X1_LOC_166/Y AND2X1_LOC_535/Y 0.80fF
C44404 AND2X1_LOC_388/Y OR2X1_LOC_166/Y 0.29fF
C58059 OR2X1_LOC_166/Y VSS 0.12fF
C5655 OR2X1_LOC_187/Y VDD 0.12fF
C10427 AND2X1_LOC_191/B OR2X1_LOC_187/Y 0.01fF
C24542 OR2X1_LOC_187/Y AND2X1_LOC_711/Y 0.01fF
C26464 OR2X1_LOC_187/Y AND2X1_LOC_191/a_8_24# 0.23fF
C35432 OR2X1_LOC_187/Y OR2X1_LOC_613/Y 0.02fF
C57933 OR2X1_LOC_187/Y VSS -0.14fF
C1057 AND2X1_LOC_707/Y AND2X1_LOC_454/a_36_24# 0.01fF
C10300 AND2X1_LOC_707/Y OR2X1_LOC_423/Y 0.03fF
C19327 AND2X1_LOC_707/Y VDD 0.74fF
C30350 AND2X1_LOC_707/Y AND2X1_LOC_605/Y 0.08fF
C40460 AND2X1_LOC_707/Y AND2X1_LOC_447/Y 0.04fF
C41388 AND2X1_LOC_707/Y AND2X1_LOC_454/Y 0.10fF
C42553 AND2X1_LOC_707/Y OR2X1_LOC_424/Y 0.02fF
C46120 AND2X1_LOC_707/Y AND2X1_LOC_454/a_8_24# 0.07fF
C46192 AND2X1_LOC_707/Y AND2X1_LOC_449/Y 0.01fF
C53752 AND2X1_LOC_707/Y AND2X1_LOC_449/a_8_24# 0.04fF
C53798 AND2X1_LOC_707/Y AND2X1_LOC_712/a_8_24# -0.00fF
C57970 AND2X1_LOC_707/Y VSS 0.06fF
C20214 AND2X1_LOC_450/Y AND2X1_LOC_451/Y 0.10fF
C25698 AND2X1_LOC_450/Y AND2X1_LOC_452/a_8_24# 0.19fF
C30578 VDD AND2X1_LOC_450/Y 0.25fF
C56902 AND2X1_LOC_450/Y VSS 0.05fF
C2658 OR2X1_LOC_506/B OR2X1_LOC_242/a_8_216# 0.06fF
C7179 OR2X1_LOC_506/B OR2X1_LOC_392/B 0.03fF
C11690 OR2X1_LOC_241/Y OR2X1_LOC_506/B 0.09fF
C11972 OR2X1_LOC_216/A OR2X1_LOC_506/B 0.02fF
C19205 OR2X1_LOC_506/B OR2X1_LOC_244/B 0.01fF
C20956 OR2X1_LOC_474/Y OR2X1_LOC_506/B 0.03fF
C25606 OR2X1_LOC_624/A OR2X1_LOC_506/B 0.05fF
C26836 OR2X1_LOC_508/A OR2X1_LOC_506/B 1.00fF
C40252 OR2X1_LOC_508/a_8_216# OR2X1_LOC_506/B 0.01fF
C42820 OR2X1_LOC_506/B OR2X1_LOC_508/Y 0.02fF
C45500 OR2X1_LOC_715/B OR2X1_LOC_506/B 0.01fF
C52876 OR2X1_LOC_506/B OR2X1_LOC_721/Y 0.03fF
C57262 OR2X1_LOC_506/B VSS 0.28fF
C4404 OR2X1_LOC_843/B OR2X1_LOC_349/A 0.03fF
C31835 OR2X1_LOC_843/B OR2X1_LOC_493/Y 0.18fF
C37715 OR2X1_LOC_343/B OR2X1_LOC_843/B 0.30fF
C39634 VDD OR2X1_LOC_843/B 0.28fF
C43539 OR2X1_LOC_561/Y OR2X1_LOC_843/B 0.01fF
C43938 OR2X1_LOC_843/B OR2X1_LOC_343/a_8_216# 0.05fF
C51269 OR2X1_LOC_362/A OR2X1_LOC_843/B 0.01fF
C56344 OR2X1_LOC_843/B VSS 0.24fF
C1495 OR2X1_LOC_449/B OR2X1_LOC_728/A 0.04fF
C8725 OR2X1_LOC_739/A OR2X1_LOC_728/A 0.01fF
C44766 OR2X1_LOC_840/A OR2X1_LOC_728/A 0.40fF
C49851 OR2X1_LOC_728/A OR2X1_LOC_728/a_8_216# 0.47fF
C56324 OR2X1_LOC_728/A VSS 0.13fF
C9292 VDD OR2X1_LOC_148/B -0.00fF
C36944 OR2X1_LOC_148/B OR2X1_LOC_148/A 0.16fF
C52193 OR2X1_LOC_148/a_8_216# OR2X1_LOC_148/B 0.47fF
C57388 OR2X1_LOC_148/B VSS 0.16fF
C5683 VDD OR2X1_LOC_467/B 0.04fF
C8543 OR2X1_LOC_467/B OR2X1_LOC_471/Y 0.09fF
C16036 OR2X1_LOC_467/B OR2X1_LOC_210/B 0.16fF
C43106 OR2X1_LOC_467/B OR2X1_LOC_467/A 0.14fF
C44895 OR2X1_LOC_467/B OR2X1_LOC_467/a_8_216# 0.01fF
C56048 OR2X1_LOC_467/B OR2X1_LOC_470/A 0.01fF
C57637 OR2X1_LOC_467/B VSS -0.48fF
C494 OR2X1_LOC_97/A OR2X1_LOC_771/B 0.05fF
C961 OR2X1_LOC_97/A OR2X1_LOC_593/B 0.02fF
C1516 OR2X1_LOC_97/A OR2X1_LOC_61/a_8_216# 0.01fF
C3449 OR2X1_LOC_97/A OR2X1_LOC_365/B 0.02fF
C4879 OR2X1_LOC_97/A OR2X1_LOC_624/A 0.03fF
C5495 OR2X1_LOC_97/A OR2X1_LOC_551/B 0.08fF
C6064 OR2X1_LOC_97/A OR2X1_LOC_439/B 0.02fF
C9217 OR2X1_LOC_97/A OR2X1_LOC_640/a_8_216# 0.04fF
C12565 OR2X1_LOC_97/A OR2X1_LOC_61/Y 0.04fF
C14700 OR2X1_LOC_97/A OR2X1_LOC_775/a_8_216# 0.03fF
C15139 OR2X1_LOC_97/A OR2X1_LOC_805/A 0.03fF
C16183 OR2X1_LOC_97/A OR2X1_LOC_228/Y 0.02fF
C17628 OR2X1_LOC_97/A OR2X1_LOC_788/a_8_216# 0.01fF
C18057 OR2X1_LOC_97/A OR2X1_LOC_174/A 0.01fF
C19733 OR2X1_LOC_97/A OR2X1_LOC_486/Y 0.03fF
C20237 OR2X1_LOC_97/A OR2X1_LOC_775/a_36_216# 0.03fF
C21008 OR2X1_LOC_97/A OR2X1_LOC_61/A 0.01fF
C22353 OR2X1_LOC_97/A OR2X1_LOC_841/A 0.03fF
C23636 OR2X1_LOC_335/Y OR2X1_LOC_97/A 0.02fF
C24533 OR2X1_LOC_97/A OR2X1_LOC_810/A 0.03fF
C24842 OR2X1_LOC_715/B OR2X1_LOC_97/A 0.05fF
C25725 OR2X1_LOC_97/A OR2X1_LOC_785/B 0.03fF
C26001 OR2X1_LOC_97/A OR2X1_LOC_181/Y 0.06fF
C26580 OR2X1_LOC_97/A OR2X1_LOC_602/A 0.01fF
C27407 OR2X1_LOC_97/A OR2X1_LOC_147/B 0.03fF
C27537 OR2X1_LOC_97/A OR2X1_LOC_545/B 0.17fF
C28673 OR2X1_LOC_97/A OR2X1_LOC_794/A 0.03fF
C28817 OR2X1_LOC_97/A OR2X1_LOC_544/A 0.32fF
C29093 OR2X1_LOC_97/A OR2X1_LOC_653/Y 0.01fF
C30984 OR2X1_LOC_97/A OR2X1_LOC_112/B 0.01fF
C31288 OR2X1_LOC_97/A OR2X1_LOC_574/A 0.03fF
C31543 OR2X1_LOC_97/A OR2X1_LOC_390/a_8_216# 0.01fF
C36570 OR2X1_LOC_97/A OR2X1_LOC_390/B 0.01fF
C36996 OR2X1_LOC_97/A OR2X1_LOC_390/a_36_216# -0.00fF
C37094 OR2X1_LOC_97/A OR2X1_LOC_61/B -0.00fF
C38514 OR2X1_LOC_97/A OR2X1_LOC_443/a_8_216# 0.01fF
C39575 OR2X1_LOC_97/A OR2X1_LOC_605/Y 0.21fF
C39757 OR2X1_LOC_97/A OR2X1_LOC_602/a_8_216# 0.01fF
C39826 OR2X1_LOC_97/A OR2X1_LOC_439/a_8_216# 0.01fF
C42334 OR2X1_LOC_97/A OR2X1_LOC_33/B 0.01fF
C42487 OR2X1_LOC_97/A OR2X1_LOC_374/Y 0.93fF
C42610 OR2X1_LOC_97/A OR2X1_LOC_392/B 0.01fF
C44799 OR2X1_LOC_97/A VDD 0.51fF
C45756 OR2X1_LOC_97/A OR2X1_LOC_462/B 0.03fF
C46119 OR2X1_LOC_97/A OR2X1_LOC_602/Y 0.01fF
C46319 OR2X1_LOC_97/A OR2X1_LOC_602/B 0.01fF
C47073 OR2X1_LOC_97/A OR2X1_LOC_840/A 0.03fF
C48668 OR2X1_LOC_97/A OR2X1_LOC_544/B 0.29fF
C49786 OR2X1_LOC_97/A OR2X1_LOC_476/B 0.02fF
C50723 OR2X1_LOC_97/A OR2X1_LOC_544/a_8_216# 0.02fF
C51075 OR2X1_LOC_97/A OR2X1_LOC_440/A 0.04fF
C51385 OR2X1_LOC_97/A OR2X1_LOC_778/Y 0.05fF
C53796 OR2X1_LOC_97/A OR2X1_LOC_34/A -0.00fF
C55970 OR2X1_LOC_97/A OR2X1_LOC_703/A 0.03fF
C56058 OR2X1_LOC_97/A OR2X1_LOC_653/a_8_216# 0.01fF
C57891 OR2X1_LOC_97/A VSS 0.37fF
C4756 OR2X1_LOC_112/B OR2X1_LOC_539/Y 0.02fF
C8201 OR2X1_LOC_112/B OR2X1_LOC_775/a_8_216# 0.47fF
C18321 OR2X1_LOC_715/B OR2X1_LOC_112/B 0.14fF
C27731 OR2X1_LOC_653/A OR2X1_LOC_112/B 0.26fF
C30098 OR2X1_LOC_112/B OR2X1_LOC_390/B 0.02fF
C38188 VDD OR2X1_LOC_112/B 0.17fF
C54566 OR2X1_LOC_624/A OR2X1_LOC_112/B 0.01fF
C56977 OR2X1_LOC_112/B VSS -0.80fF
C5777 OR2X1_LOC_493/B OR2X1_LOC_493/A 0.02fF
C8851 OR2X1_LOC_493/B OR2X1_LOC_805/A 0.05fF
C30376 OR2X1_LOC_493/B OR2X1_LOC_493/a_8_216# 0.01fF
C30621 OR2X1_LOC_493/B OR2X1_LOC_493/Y 0.79fF
C48035 OR2X1_LOC_493/B OR2X1_LOC_737/A 0.11fF
C57695 OR2X1_LOC_493/B VSS 0.10fF
C4332 OR2X1_LOC_559/B AND2X1_LOC_88/Y 0.03fF
C23563 OR2X1_LOC_559/B OR2X1_LOC_559/a_8_216# 0.50fF
C34474 OR2X1_LOC_559/B OR2X1_LOC_559/a_36_216# 0.02fF
C41114 OR2X1_LOC_520/Y OR2X1_LOC_559/B 0.46fF
C45792 VDD OR2X1_LOC_559/B 0.02fF
C57491 OR2X1_LOC_559/B VSS 0.19fF
C23063 OR2X1_LOC_76/B OR2X1_LOC_76/A 0.04fF
C29409 OR2X1_LOC_76/B OR2X1_LOC_241/B 0.06fF
C34056 OR2X1_LOC_76/B OR2X1_LOC_318/B 0.10fF
C47721 OR2X1_LOC_76/B OR2X1_LOC_76/Y 0.06fF
C51223 OR2X1_LOC_76/B OR2X1_LOC_76/a_8_216# 0.05fF
C57590 OR2X1_LOC_76/B VSS 0.24fF
C334 OR2X1_LOC_466/A OR2X1_LOC_449/A 0.14fF
C7376 OR2X1_LOC_449/A OR2X1_LOC_796/B 0.02fF
C28986 OR2X1_LOC_446/Y OR2X1_LOC_449/A 0.47fF
C32784 OR2X1_LOC_449/A OR2X1_LOC_783/A 0.26fF
C46972 OR2X1_LOC_449/A OR2X1_LOC_779/Y 0.01fF
C47943 OR2X1_LOC_449/A OR2X1_LOC_712/B -0.00fF
C52500 OR2X1_LOC_449/A OR2X1_LOC_783/a_8_216# 0.49fF
C57074 OR2X1_LOC_449/A VSS 0.46fF
C1589 OR2X1_LOC_114/B OR2X1_LOC_347/B 0.03fF
C7609 OR2X1_LOC_347/a_8_216# OR2X1_LOC_347/B 0.01fF
C15422 OR2X1_LOC_347/B OR2X1_LOC_675/Y 0.09fF
C31200 OR2X1_LOC_347/A OR2X1_LOC_347/B 0.06fF
C51842 OR2X1_LOC_347/B OR2X1_LOC_347/Y 0.05fF
C56663 OR2X1_LOC_347/B VSS 0.10fF
C3556 OR2X1_LOC_147/B OR2X1_LOC_705/B 0.02fF
C6835 OR2X1_LOC_705/B OR2X1_LOC_726/A 0.02fF
C7184 OR2X1_LOC_705/B OR2X1_LOC_727/a_8_216# 0.14fF
C9144 OR2X1_LOC_486/B OR2X1_LOC_705/B 0.14fF
C20957 VDD OR2X1_LOC_705/B 0.27fF
C23639 OR2X1_LOC_471/Y OR2X1_LOC_705/B 0.14fF
C29272 OR2X1_LOC_705/B OR2X1_LOC_731/A 0.14fF
C39033 OR2X1_LOC_149/B OR2X1_LOC_705/B 0.01fF
C43027 OR2X1_LOC_705/B OR2X1_LOC_739/A 0.01fF
C43070 OR2X1_LOC_546/B OR2X1_LOC_705/B 0.05fF
C51983 OR2X1_LOC_705/B OR2X1_LOC_486/Y 0.01fF
C52108 OR2X1_LOC_486/a_8_216# OR2X1_LOC_705/B 0.48fF
C52328 OR2X1_LOC_705/B OR2X1_LOC_308/Y 0.14fF
C53144 OR2X1_LOC_705/B OR2X1_LOC_550/B 0.05fF
C56906 OR2X1_LOC_705/B VSS -0.86fF
C29767 OR2X1_LOC_124/B OR2X1_LOC_786/Y -0.00fF
C30053 OR2X1_LOC_124/B OR2X1_LOC_204/Y 0.08fF
C35521 OR2X1_LOC_124/B OR2X1_LOC_203/Y 0.18fF
C41830 OR2X1_LOC_124/A OR2X1_LOC_124/B 0.05fF
C50920 OR2X1_LOC_124/B OR2X1_LOC_124/a_8_216# 0.03fF
C54242 OR2X1_LOC_124/B OR2X1_LOC_641/A 0.07fF
C55250 OR2X1_LOC_124/B OR2X1_LOC_124/Y 0.16fF
C57982 OR2X1_LOC_124/B VSS -0.01fF
C2583 OR2X1_LOC_403/B OR2X1_LOC_403/A 0.07fF
C5575 OR2X1_LOC_403/B OR2X1_LOC_403/a_8_216# 0.05fF
C13252 OR2X1_LOC_400/A OR2X1_LOC_403/B 1.20fF
C27263 OR2X1_LOC_403/B AND2X1_LOC_79/Y 0.04fF
C47372 OR2X1_LOC_403/B OR2X1_LOC_624/B 0.03fF
C47704 OR2X1_LOC_403/B OR2X1_LOC_400/a_8_216# 0.01fF
C55978 OR2X1_LOC_403/B OR2X1_LOC_771/B 0.14fF
C57664 OR2X1_LOC_403/B VSS 0.26fF
C2724 OR2X1_LOC_791/A OR2X1_LOC_345/a_8_216# 0.18fF
C5146 OR2X1_LOC_791/A OR2X1_LOC_792/A 0.95fF
C25109 OR2X1_LOC_791/A OR2X1_LOC_345/A 0.08fF
C26692 OR2X1_LOC_791/A OR2X1_LOC_555/B 0.80fF
C30837 OR2X1_LOC_791/A VDD 0.04fF
C41942 OR2X1_LOC_791/B OR2X1_LOC_791/A 0.03fF
C57928 OR2X1_LOC_791/A VSS 0.18fF
C4471 OR2X1_LOC_643/A OR2X1_LOC_115/B 0.83fF
C9269 OR2X1_LOC_404/Y OR2X1_LOC_115/B 0.02fF
C11167 OR2X1_LOC_115/B OR2X1_LOC_554/a_8_216# 0.18fF
C21528 OR2X1_LOC_575/A OR2X1_LOC_115/B 0.03fF
C23616 OR2X1_LOC_632/a_8_216# OR2X1_LOC_115/B 0.01fF
C28227 OR2X1_LOC_632/Y OR2X1_LOC_115/B 0.68fF
C33757 OR2X1_LOC_510/Y OR2X1_LOC_115/B 0.42fF
C33790 OR2X1_LOC_810/A OR2X1_LOC_115/B 0.01fF
C34086 OR2X1_LOC_715/B OR2X1_LOC_115/B 0.13fF
C37024 OR2X1_LOC_114/B OR2X1_LOC_115/B 0.02fF
C38299 OR2X1_LOC_140/A OR2X1_LOC_115/B 0.03fF
C40548 OR2X1_LOC_574/A OR2X1_LOC_115/B 0.07fF
C40933 OR2X1_LOC_203/Y OR2X1_LOC_115/B 0.07fF
C46026 OR2X1_LOC_115/B OR2X1_LOC_844/B 0.17fF
C48597 OR2X1_LOC_115/B OR2X1_LOC_560/A 0.02fF
C50815 OR2X1_LOC_140/B OR2X1_LOC_115/B 0.59fF
C54196 VDD OR2X1_LOC_115/B 0.07fF
C56489 OR2X1_LOC_115/B VSS -0.21fF
C292 OR2X1_LOC_643/A OR2X1_LOC_113/B 1.62fF
C2428 OR2X1_LOC_523/Y OR2X1_LOC_113/B 0.01fF
C4562 OR2X1_LOC_844/a_8_216# OR2X1_LOC_113/B 0.01fF
C5279 OR2X1_LOC_474/Y OR2X1_LOC_113/B 0.26fF
C10610 OR2X1_LOC_849/a_8_216# OR2X1_LOC_113/B 0.01fF
C14282 OR2X1_LOC_624/a_8_216# OR2X1_LOC_113/B 0.01fF
C15499 OR2X1_LOC_768/A OR2X1_LOC_113/B 0.16fF
C19341 OR2X1_LOC_113/B OR2X1_LOC_772/A 0.01fF
C21693 OR2X1_LOC_849/a_36_216# OR2X1_LOC_113/B -0.00fF
C27168 OR2X1_LOC_474/a_8_216# OR2X1_LOC_113/B 0.01fF
C27183 OR2X1_LOC_859/A OR2X1_LOC_113/B 0.01fF
C29613 OR2X1_LOC_810/A OR2X1_LOC_113/B 0.05fF
C47888 OR2X1_LOC_392/B OR2X1_LOC_113/B 0.05fF
C48395 OR2X1_LOC_624/Y OR2X1_LOC_113/B 0.03fF
C50060 VDD OR2X1_LOC_113/B 0.15fF
C53137 OR2X1_LOC_624/B OR2X1_LOC_113/B 0.89fF
C53392 OR2X1_LOC_113/B OR2X1_LOC_768/a_8_216# 0.49fF
C53811 OR2X1_LOC_474/B OR2X1_LOC_113/B 0.02fF
C55698 OR2X1_LOC_844/Y OR2X1_LOC_113/B 0.03fF
C56065 OR2X1_LOC_849/A OR2X1_LOC_113/B 0.01fF
C56513 OR2X1_LOC_113/B VSS 0.30fF
C7803 VDD OR2X1_LOC_209/A 0.04fF
C10518 OR2X1_LOC_471/Y OR2X1_LOC_209/A 0.09fF
C16214 OR2X1_LOC_209/A OR2X1_LOC_731/A 0.07fF
C22289 OR2X1_LOC_797/B OR2X1_LOC_209/A 0.14fF
C25138 OR2X1_LOC_209/A OR2X1_LOC_726/a_8_216# 0.24fF
C25992 OR2X1_LOC_149/B OR2X1_LOC_209/A 0.03fF
C29912 OR2X1_LOC_739/A OR2X1_LOC_209/A 0.01fF
C32869 OR2X1_LOC_213/A OR2X1_LOC_209/A 0.03fF
C38333 OR2X1_LOC_209/a_8_216# OR2X1_LOC_209/A 0.18fF
C39893 OR2X1_LOC_209/A OR2X1_LOC_550/B 0.88fF
C49986 OR2X1_LOC_726/A OR2X1_LOC_209/A 0.12fF
C52178 OR2X1_LOC_486/B OR2X1_LOC_209/A 0.04fF
C56421 OR2X1_LOC_209/A VSS 0.17fF
C24316 OR2X1_LOC_400/A OR2X1_LOC_624/B 0.01fF
C32860 OR2X1_LOC_400/A OR2X1_LOC_771/B 0.02fF
C37307 OR2X1_LOC_400/B OR2X1_LOC_400/A 0.28fF
C57940 OR2X1_LOC_400/A VSS 0.14fF
C1998 OR2X1_LOC_207/B OR2X1_LOC_793/A 0.02fF
C32578 VDD OR2X1_LOC_793/A 0.08fF
C33423 OR2X1_LOC_676/Y OR2X1_LOC_793/A 0.02fF
C47444 OR2X1_LOC_793/A AND2X1_LOC_39/Y 0.16fF
C48178 OR2X1_LOC_793/A OR2X1_LOC_793/a_8_216# 0.01fF
C57096 OR2X1_LOC_793/A VSS 0.11fF
C4690 OR2X1_LOC_639/B OR2X1_LOC_636/A 0.08fF
C10280 OR2X1_LOC_639/B OR2X1_LOC_636/B 0.06fF
C20542 OR2X1_LOC_639/B OR2X1_LOC_639/a_8_216# 0.07fF
C21365 OR2X1_LOC_639/B OR2X1_LOC_636/a_8_216# 0.06fF
C37772 OR2X1_LOC_639/B OR2X1_LOC_639/A 0.09fF
C45803 VDD OR2X1_LOC_639/B 0.12fF
C57408 OR2X1_LOC_639/B VSS 0.27fF
C943 OR2X1_LOC_175/Y OR2X1_LOC_771/B 0.12fF
C3216 OR2X1_LOC_520/Y OR2X1_LOC_771/B 0.01fF
C4791 OR2X1_LOC_641/Y OR2X1_LOC_771/B 0.10fF
C7468 OR2X1_LOC_654/A OR2X1_LOC_771/B 0.02fF
C7794 VDD OR2X1_LOC_771/B 1.94fF
C8754 OR2X1_LOC_462/B OR2X1_LOC_771/B 0.05fF
C9549 OR2X1_LOC_35/Y OR2X1_LOC_771/B 0.03fF
C10881 OR2X1_LOC_624/B OR2X1_LOC_771/B 0.07fF
C10882 OR2X1_LOC_33/a_8_216# OR2X1_LOC_771/B 0.05fF
C11224 OR2X1_LOC_400/a_8_216# OR2X1_LOC_771/B 0.06fF
C12602 OR2X1_LOC_476/B OR2X1_LOC_771/B 0.10fF
C19772 OR2X1_LOC_402/Y OR2X1_LOC_771/B 0.07fF
C21981 OR2X1_LOC_647/Y OR2X1_LOC_771/B 0.08fF
C23975 OR2X1_LOC_786/A OR2X1_LOC_771/B 0.06fF
C24066 OR2X1_LOC_400/B OR2X1_LOC_771/B 0.01fF
C24207 OR2X1_LOC_84/Y OR2X1_LOC_771/B 0.03fF
C26984 OR2X1_LOC_633/B OR2X1_LOC_771/B 0.05fF
C29842 OR2X1_LOC_786/a_8_216# OR2X1_LOC_771/B 0.26fF
C31081 OR2X1_LOC_770/A OR2X1_LOC_771/B 0.30fF
C33780 OR2X1_LOC_401/A OR2X1_LOC_771/B 0.03fF
C35914 OR2X1_LOC_244/A OR2X1_LOC_771/B 0.07fF
C38395 OR2X1_LOC_656/a_8_216# OR2X1_LOC_771/B 0.35fF
C38495 OR2X1_LOC_770/Y OR2X1_LOC_771/B 0.06fF
C44719 OR2X1_LOC_857/B OR2X1_LOC_771/B 0.03fF
C44871 OR2X1_LOC_401/B OR2X1_LOC_771/B 0.03fF
C45260 OR2X1_LOC_835/B OR2X1_LOC_771/B 0.07fF
C48394 OR2X1_LOC_646/A OR2X1_LOC_771/B 0.43fF
C49651 OR2X1_LOC_84/B OR2X1_LOC_771/B 0.07fF
C49800 OR2X1_LOC_771/a_8_216# OR2X1_LOC_771/B 0.08fF
C56461 OR2X1_LOC_771/B VSS 0.59fF
C18871 AND2X1_LOC_463/B AND2X1_LOC_463/a_8_24# 0.11fF
C54514 VDD AND2X1_LOC_463/B 0.09fF
C57044 AND2X1_LOC_463/B VSS 0.17fF
C41621 VDD AND2X1_LOC_451/Y 0.08fF
C56901 AND2X1_LOC_451/Y VSS 0.02fF
C24402 AND2X1_LOC_452/Y OR2X1_LOC_163/Y 0.08fF
C52447 VDD OR2X1_LOC_163/Y 0.13fF
C56289 OR2X1_LOC_163/Y VSS 0.35fF
C2734 OR2X1_LOC_525/Y AND2X1_LOC_796/A 0.10fF
C3308 OR2X1_LOC_526/Y OR2X1_LOC_525/Y 0.07fF
C5763 VDD OR2X1_LOC_525/Y 0.05fF
C56221 OR2X1_LOC_525/Y OR2X1_LOC_680/Y 0.15fF
C57748 OR2X1_LOC_525/Y VSS 0.19fF
C39 AND2X1_LOC_717/B OR2X1_LOC_238/Y 0.03fF
C1725 AND2X1_LOC_833/a_8_24# OR2X1_LOC_238/Y 0.01fF
C2482 OR2X1_LOC_238/Y AND2X1_LOC_786/Y 0.01fF
C7219 AND2X1_LOC_840/A OR2X1_LOC_238/Y 0.28fF
C8260 AND2X1_LOC_851/B OR2X1_LOC_238/Y 0.04fF
C12619 AND2X1_LOC_564/B OR2X1_LOC_238/Y 0.01fF
C16925 AND2X1_LOC_719/Y OR2X1_LOC_238/Y 0.20fF
C17813 AND2X1_LOC_840/a_8_24# OR2X1_LOC_238/Y 0.01fF
C18326 OR2X1_LOC_237/Y OR2X1_LOC_238/Y 0.06fF
C23436 AND2X1_LOC_851/A OR2X1_LOC_238/Y 0.01fF
C26866 AND2X1_LOC_465/Y OR2X1_LOC_238/Y 0.02fF
C28397 VDD OR2X1_LOC_238/Y 0.27fF
C28855 AND2X1_LOC_486/Y OR2X1_LOC_238/Y 0.10fF
C32077 AND2X1_LOC_721/Y OR2X1_LOC_238/Y 0.06fF
C40551 OR2X1_LOC_238/Y AND2X1_LOC_241/a_8_24# 0.05fF
C51807 OR2X1_LOC_238/Y AND2X1_LOC_242/B 0.01fF
C52360 OR2X1_LOC_495/Y OR2X1_LOC_238/Y 0.85fF
C56713 OR2X1_LOC_238/Y VSS 0.09fF
C5372 OR2X1_LOC_52/Y AND2X1_LOC_208/Y 0.11fF
C28835 VDD OR2X1_LOC_52/Y 0.23fF
C55906 OR2X1_LOC_52/Y OR2X1_LOC_7/Y 0.36fF
C56969 OR2X1_LOC_52/Y VSS 0.19fF
C772 AND2X1_LOC_191/B OR2X1_LOC_251/Y 0.03fF
C4644 OR2X1_LOC_667/Y OR2X1_LOC_251/Y 0.01fF
C5033 AND2X1_LOC_721/a_8_24# OR2X1_LOC_251/Y 0.01fF
C6929 OR2X1_LOC_251/Y AND2X1_LOC_721/A 0.02fF
C15698 AND2X1_LOC_720/a_8_24# OR2X1_LOC_251/Y 0.01fF
C24598 OR2X1_LOC_251/Y OR2X1_LOC_494/Y 0.03fF
C29296 OR2X1_LOC_251/Y OR2X1_LOC_250/Y 1.40fF
C40602 AND2X1_LOC_719/Y OR2X1_LOC_251/Y 0.01fF
C43794 OR2X1_LOC_251/Y AND2X1_LOC_287/Y 0.01fF
C45085 OR2X1_LOC_251/Y AND2X1_LOC_859/a_8_24# -0.00fF
C48552 AND2X1_LOC_366/A OR2X1_LOC_251/Y 0.03fF
C51555 OR2X1_LOC_251/Y AND2X1_LOC_859/Y 0.23fF
C52289 VDD OR2X1_LOC_251/Y 0.42fF
C55740 AND2X1_LOC_720/Y OR2X1_LOC_251/Y 0.01fF
C56038 AND2X1_LOC_721/Y OR2X1_LOC_251/Y 0.01fF
C57729 OR2X1_LOC_251/Y VSS 0.24fF
C9356 AND2X1_LOC_658/B OR2X1_LOC_680/Y 0.03fF
C11083 AND2X1_LOC_546/a_8_24# OR2X1_LOC_680/Y 0.23fF
C12031 OR2X1_LOC_680/Y OR2X1_LOC_679/A 0.01fF
C16407 AND2X1_LOC_544/Y OR2X1_LOC_680/Y 0.09fF
C20409 OR2X1_LOC_524/Y OR2X1_LOC_680/Y 0.03fF
C22391 OR2X1_LOC_680/Y OR2X1_LOC_142/Y 0.02fF
C25943 AND2X1_LOC_728/Y OR2X1_LOC_680/Y 0.01fF
C39408 OR2X1_LOC_680/Y AND2X1_LOC_658/A 0.03fF
C43708 OR2X1_LOC_526/Y OR2X1_LOC_680/Y 0.38fF
C46023 OR2X1_LOC_680/Y AND2X1_LOC_728/a_8_24# 0.11fF
C46320 VDD OR2X1_LOC_680/Y 0.30fF
C57691 OR2X1_LOC_680/Y VSS -0.07fF
C19643 OR2X1_LOC_145/Y AND2X1_LOC_148/a_8_24# 0.23fF
C40284 VDD OR2X1_LOC_145/Y 0.12fF
C45261 OR2X1_LOC_145/Y OR2X1_LOC_146/Y 0.09fF
C46817 OR2X1_LOC_145/Y AND2X1_LOC_213/B 0.01fF
C57223 OR2X1_LOC_145/Y VSS 0.06fF
C15076 AND2X1_LOC_390/a_8_24# OR2X1_LOC_533/Y 0.01fF
C24429 OR2X1_LOC_533/Y AND2X1_LOC_788/a_8_24# 0.01fF
C26113 AND2X1_LOC_392/A OR2X1_LOC_533/Y 0.15fF
C27909 OR2X1_LOC_533/Y AND2X1_LOC_645/A 0.11fF
C29893 OR2X1_LOC_533/Y AND2X1_LOC_794/B 0.79fF
C54647 AND2X1_LOC_388/Y OR2X1_LOC_533/Y 0.28fF
C58004 OR2X1_LOC_533/Y VSS 0.19fF
C36789 AND2X1_LOC_468/B OR2X1_LOC_594/Y 0.23fF
C48119 AND2X1_LOC_652/a_8_24# OR2X1_LOC_594/Y 0.01fF
C53279 AND2X1_LOC_810/Y OR2X1_LOC_594/Y 0.25fF
C53599 AND2X1_LOC_653/B OR2X1_LOC_594/Y 0.10fF
C55557 AND2X1_LOC_794/B OR2X1_LOC_594/Y 0.50fF
C55589 VDD OR2X1_LOC_594/Y 0.12fF
C56710 OR2X1_LOC_594/Y VSS -0.32fF
C278 OR2X1_LOC_406/Y AND2X1_LOC_475/a_8_24# -0.00fF
C2005 OR2X1_LOC_406/Y OR2X1_LOC_189/Y 0.03fF
C3575 OR2X1_LOC_406/Y AND2X1_LOC_734/a_8_24# 0.01fF
C4429 OR2X1_LOC_406/Y AND2X1_LOC_734/Y 0.01fF
C10407 OR2X1_LOC_528/Y OR2X1_LOC_406/Y 0.01fF
C13111 OR2X1_LOC_406/Y AND2X1_LOC_711/Y 0.04fF
C13406 OR2X1_LOC_406/Y AND2X1_LOC_658/B 0.03fF
C29994 OR2X1_LOC_496/Y OR2X1_LOC_406/Y 0.71fF
C34467 AND2X1_LOC_564/B OR2X1_LOC_406/Y 0.02fF
C46569 AND2X1_LOC_565/B OR2X1_LOC_406/Y 0.02fF
C50459 OR2X1_LOC_406/Y VDD -0.00fF
C54173 OR2X1_LOC_406/Y AND2X1_LOC_721/Y 0.01fF
C57963 OR2X1_LOC_406/Y VSS 0.16fF
C3784 OR2X1_LOC_189/Y VDD 0.35fF
C8038 OR2X1_LOC_189/Y OR2X1_LOC_679/Y 0.14fF
C10114 OR2X1_LOC_189/Y AND2X1_LOC_213/B 0.05fF
C11565 OR2X1_LOC_189/Y OR2X1_LOC_152/Y 0.03fF
C19934 OR2X1_LOC_528/Y OR2X1_LOC_189/Y 0.03fF
C22690 OR2X1_LOC_189/Y AND2X1_LOC_711/Y 2.18fF
C33920 OR2X1_LOC_189/Y OR2X1_LOC_524/Y 0.07fF
C35222 OR2X1_LOC_189/Y AND2X1_LOC_565/Y 0.01fF
C35451 AND2X1_LOC_726/Y OR2X1_LOC_189/Y 0.10fF
C38874 OR2X1_LOC_189/Y AND2X1_LOC_192/a_8_24# 0.09fF
C39473 AND2X1_LOC_728/Y OR2X1_LOC_189/Y 0.03fF
C40956 AND2X1_LOC_727/Y OR2X1_LOC_189/Y 0.03fF
C46544 OR2X1_LOC_189/Y AND2X1_LOC_781/Y 0.15fF
C54372 OR2X1_LOC_189/Y AND2X1_LOC_476/Y 1.49fF
C54943 OR2X1_LOC_189/Y AND2X1_LOC_474/Y 1.42fF
C55855 OR2X1_LOC_189/Y AND2X1_LOC_797/A 0.14fF
C56120 AND2X1_LOC_565/B OR2X1_LOC_189/Y 0.26fF
C57885 OR2X1_LOC_189/Y VSS 0.12fF
C1419 AND2X1_LOC_778/Y OR2X1_LOC_142/Y 0.07fF
C2257 AND2X1_LOC_786/Y OR2X1_LOC_142/Y 0.07fF
C2292 AND2X1_LOC_499/a_36_24# OR2X1_LOC_142/Y 0.01fF
C7780 AND2X1_LOC_784/Y OR2X1_LOC_142/Y 0.03fF
C7880 OR2X1_LOC_496/Y OR2X1_LOC_142/Y 0.03fF
C9485 AND2X1_LOC_727/Y OR2X1_LOC_142/Y 0.06fF
C9650 AND2X1_LOC_830/a_8_24# OR2X1_LOC_142/Y 0.03fF
C12440 AND2X1_LOC_564/B OR2X1_LOC_142/Y 0.07fF
C21453 AND2X1_LOC_658/A OR2X1_LOC_142/Y 0.03fF
C22737 AND2X1_LOC_476/Y OR2X1_LOC_142/Y 0.07fF
C25072 AND2X1_LOC_796/A OR2X1_LOC_142/Y 0.55fF
C25794 AND2X1_LOC_810/Y OR2X1_LOC_142/Y 0.37fF
C26184 AND2X1_LOC_830/a_36_24# OR2X1_LOC_142/Y 0.01fF
C26817 OR2X1_LOC_516/Y OR2X1_LOC_142/Y 9.94fF
C28183 VDD OR2X1_LOC_142/Y 0.53fF
C31901 AND2X1_LOC_721/Y OR2X1_LOC_142/Y 0.03fF
C35831 OR2X1_LOC_91/Y OR2X1_LOC_142/Y 0.03fF
C40129 AND2X1_LOC_675/A OR2X1_LOC_142/Y 0.07fF
C46504 AND2X1_LOC_727/a_8_24# OR2X1_LOC_142/Y 0.01fF
C47430 AND2X1_LOC_499/a_8_24# OR2X1_LOC_142/Y 0.03fF
C48710 OR2X1_LOC_108/Y OR2X1_LOC_142/Y 0.14fF
C49090 OR2X1_LOC_373/Y OR2X1_LOC_142/Y 0.07fF
C50142 OR2X1_LOC_679/A OR2X1_LOC_142/Y 0.15fF
C52103 OR2X1_LOC_495/Y OR2X1_LOC_142/Y 0.06fF
C52901 AND2X1_LOC_785/Y OR2X1_LOC_142/Y 0.03fF
C54656 AND2X1_LOC_550/A OR2X1_LOC_142/Y 1.04fF
C56243 OR2X1_LOC_142/Y VSS 0.19fF
C19242 OR2X1_LOC_503/Y AND2X1_LOC_573/A 0.01fF
C28899 VDD OR2X1_LOC_503/Y 0.16fF
C29371 AND2X1_LOC_486/Y OR2X1_LOC_503/Y 0.19fF
C36081 OR2X1_LOC_503/Y AND2X1_LOC_509/a_8_24# 0.23fF
C57302 OR2X1_LOC_503/Y VSS -0.00fF
C7326 OR2X1_LOC_321/Y AND2X1_LOC_324/a_8_24# 0.23fF
C24236 VDD OR2X1_LOC_321/Y 0.16fF
C38206 AND2X1_LOC_702/Y OR2X1_LOC_321/Y 0.01fF
C46924 OR2X1_LOC_320/Y OR2X1_LOC_321/Y 0.19fF
C57541 OR2X1_LOC_321/Y VSS 0.07fF
C1071 OR2X1_LOC_591/Y VDD 0.04fF
C12142 OR2X1_LOC_591/Y AND2X1_LOC_605/Y 0.17fF
C23260 OR2X1_LOC_591/Y AND2X1_LOC_722/A 0.79fF
C58115 OR2X1_LOC_591/Y VSS 0.15fF
C29169 VDD OR2X1_LOC_250/Y 0.03fF
C57434 OR2X1_LOC_250/Y VSS 0.30fF
C4499 OR2X1_LOC_667/Y VDD 0.12fF
C24218 OR2X1_LOC_667/Y AND2X1_LOC_720/a_8_24# 0.23fF
C32957 OR2X1_LOC_667/Y OR2X1_LOC_494/Y 0.01fF
C58090 OR2X1_LOC_667/Y VSS 0.06fF
C5017 AND2X1_LOC_724/A OR2X1_LOC_167/Y 0.05fF
C5167 OR2X1_LOC_312/Y OR2X1_LOC_167/Y 0.09fF
C10238 AND2X1_LOC_535/Y OR2X1_LOC_167/Y 0.02fF
C14886 AND2X1_LOC_388/Y OR2X1_LOC_167/Y 0.07fF
C22250 AND2X1_LOC_388/a_8_24# OR2X1_LOC_167/Y 0.03fF
C24232 OR2X1_LOC_176/Y OR2X1_LOC_167/Y 0.03fF
C25011 AND2X1_LOC_539/Y OR2X1_LOC_167/Y 0.04fF
C27678 AND2X1_LOC_703/a_8_24# OR2X1_LOC_167/Y 0.23fF
C37679 AND2X1_LOC_810/A OR2X1_LOC_167/Y 0.16fF
C38687 AND2X1_LOC_388/a_36_24# OR2X1_LOC_167/Y 0.01fF
C41944 AND2X1_LOC_715/Y OR2X1_LOC_167/Y 0.05fF
C43869 OR2X1_LOC_167/Y AND2X1_LOC_661/A 0.02fF
C46396 VDD OR2X1_LOC_167/Y 0.37fF
C57280 OR2X1_LOC_167/Y VSS 0.27fF
C5270 OR2X1_LOC_259/a_8_216# OR2X1_LOC_259/A 0.47fF
C9001 OR2X1_LOC_259/A OR2X1_LOC_348/B 0.11fF
C56412 OR2X1_LOC_259/A VSS 0.04fF
C8978 OR2X1_LOC_462/B OR2X1_LOC_642/a_8_216# 0.03fF
C14491 OR2X1_LOC_462/B OR2X1_LOC_642/a_36_216# 0.03fF
C17407 OR2X1_LOC_640/a_8_216# OR2X1_LOC_462/B 0.01fF
C48581 OR2X1_LOC_520/Y OR2X1_LOC_462/B 0.01fF
C50173 OR2X1_LOC_641/Y OR2X1_LOC_462/B 0.01fF
C53125 VDD OR2X1_LOC_462/B 0.45fF
C54956 OR2X1_LOC_462/B OR2X1_LOC_416/Y 0.39fF
C55652 OR2X1_LOC_640/Y OR2X1_LOC_462/B 0.01fF
C57653 OR2X1_LOC_462/B VSS 0.36fF
C20449 OR2X1_LOC_210/B OR2X1_LOC_210/a_8_216# 0.47fF
C57277 OR2X1_LOC_210/B VSS 0.16fF
C1139 OR2X1_LOC_181/B OR2X1_LOC_565/A 0.13fF
C1162 OR2X1_LOC_181/B OR2X1_LOC_190/Y 0.06fF
C4978 OR2X1_LOC_181/B OR2X1_LOC_540/a_8_216# 0.02fF
C11923 OR2X1_LOC_181/B OR2X1_LOC_564/A 0.12fF
C16083 OR2X1_LOC_181/B OR2X1_LOC_540/a_36_216# 0.03fF
C16725 OR2X1_LOC_181/B OR2X1_LOC_181/A 0.09fF
C33262 OR2X1_LOC_181/B OR2X1_LOC_181/a_8_216# 0.01fF
C40395 OR2X1_LOC_181/B OR2X1_LOC_192/B 0.11fF
C40568 VDD OR2X1_LOC_181/B 0.10fF
C43385 OR2X1_LOC_181/B OR2X1_LOC_471/Y 0.03fF
C44533 OR2X1_LOC_181/B OR2X1_LOC_190/B 0.05fF
C57391 OR2X1_LOC_181/B VSS 0.14fF
C56987 OR2X1_LOC_781/A VSS 0.13fF
C13844 OR2X1_LOC_499/B OR2X1_LOC_563/A 0.12fF
C22903 OR2X1_LOC_501/B OR2X1_LOC_499/B 0.11fF
C24581 OR2X1_LOC_499/B OR2X1_LOC_833/B 0.05fF
C27166 OR2X1_LOC_499/B OR2X1_LOC_203/Y 0.15fF
C32300 OR2X1_LOC_499/B OR2X1_LOC_493/Y 0.01fF
C34328 OR2X1_LOC_499/B OR2X1_LOC_778/A 1.33fF
C42824 OR2X1_LOC_499/B OR2X1_LOC_499/a_8_216# 0.07fF
C57735 OR2X1_LOC_499/B VSS 0.40fF
C11550 OR2X1_LOC_676/Y AND2X1_LOC_39/Y 0.01fF
C36281 AND2X1_LOC_39/Y OR2X1_LOC_194/a_8_216# 0.47fF
C56382 AND2X1_LOC_39/Y VSS 0.15fF
C23858 VDD OR2X1_LOC_148/A 0.21fF
C57327 OR2X1_LOC_148/A VSS 0.12fF
C4387 OR2X1_LOC_324/B OR2X1_LOC_308/Y 0.14fF
C26642 OR2X1_LOC_324/a_8_216# OR2X1_LOC_324/B 0.01fF
C37593 OR2X1_LOC_326/B OR2X1_LOC_324/B 0.79fF
C51420 OR2X1_LOC_324/B OR2X1_LOC_739/A 0.01fF
C57790 OR2X1_LOC_324/B VSS 0.10fF
C1848 OR2X1_LOC_644/B OR2X1_LOC_644/A 0.04fF
C33152 VDD OR2X1_LOC_644/A 0.05fF
C37907 OR2X1_LOC_644/a_8_216# OR2X1_LOC_644/A 0.47fF
C56312 OR2X1_LOC_644/A VSS 0.29fF
C319 OR2X1_LOC_646/a_8_216# OR2X1_LOC_646/B 0.02fF
C4853 VDD OR2X1_LOC_646/B 0.02fF
C11401 OR2X1_LOC_647/A OR2X1_LOC_646/B 0.67fF
C30468 OR2X1_LOC_647/B OR2X1_LOC_646/B 0.02fF
C45388 OR2X1_LOC_646/A OR2X1_LOC_646/B 0.02fF
C56528 OR2X1_LOC_646/B VSS 0.32fF
C16613 OR2X1_LOC_805/A OR2X1_LOC_778/A 0.01fF
C19907 OR2X1_LOC_778/A OR2X1_LOC_563/A 0.14fF
C33154 OR2X1_LOC_778/A OR2X1_LOC_203/Y 0.01fF
C38312 OR2X1_LOC_778/A OR2X1_LOC_493/Y 0.69fF
C46330 VDD OR2X1_LOC_778/A 0.18fF
C48721 OR2X1_LOC_241/Y OR2X1_LOC_778/A 0.04fF
C52873 OR2X1_LOC_778/A OR2X1_LOC_778/Y 0.11fF
C55790 OR2X1_LOC_778/A OR2X1_LOC_737/A 0.02fF
C56908 OR2X1_LOC_778/A VSS 0.58fF
C19200 OR2X1_LOC_805/A OR2X1_LOC_719/A 0.03fF
C26938 OR2X1_LOC_719/A OR2X1_LOC_241/B 0.41fF
C48965 VDD OR2X1_LOC_719/A 0.21fF
C56921 OR2X1_LOC_719/A VSS 0.12fF
C7346 OR2X1_LOC_244/A AND2X1_LOC_79/Y 0.08fF
C7773 OR2X1_LOC_404/A AND2X1_LOC_79/Y 0.80fF
C23926 AND2X1_LOC_79/Y OR2X1_LOC_204/a_8_216# 0.01fF
C29376 AND2X1_LOC_79/Y OR2X1_LOC_204/a_36_216# 0.02fF
C35131 VDD AND2X1_LOC_79/Y 0.03fF
C38228 OR2X1_LOC_624/B AND2X1_LOC_79/Y 0.01fF
C52914 OR2X1_LOC_403/a_8_216# AND2X1_LOC_79/Y 0.01fF
C56953 AND2X1_LOC_79/Y VSS -0.80fF
C1266 OR2X1_LOC_859/a_8_216# OR2X1_LOC_810/A 0.09fF
C1694 OR2X1_LOC_810/A OR2X1_LOC_775/a_8_216# 0.05fF
C2173 OR2X1_LOC_810/A OR2X1_LOC_805/A 0.15fF
C3187 OR2X1_LOC_810/A OR2X1_LOC_228/Y 0.07fF
C5876 OR2X1_LOC_810/A OR2X1_LOC_632/Y 0.10fF
C9909 OR2X1_LOC_473/Y OR2X1_LOC_810/A 0.01fF
C10257 OR2X1_LOC_652/a_36_216# OR2X1_LOC_810/A 0.02fF
C10657 OR2X1_LOC_810/a_8_216# OR2X1_LOC_810/A 0.06fF
C10700 OR2X1_LOC_859/B OR2X1_LOC_810/A 0.03fF
C11514 OR2X1_LOC_510/Y OR2X1_LOC_810/A 0.03fF
C11826 OR2X1_LOC_715/B OR2X1_LOC_810/A 0.01fF
C12758 OR2X1_LOC_810/A OR2X1_LOC_785/B 0.07fF
C12925 OR2X1_LOC_810/A OR2X1_LOC_786/Y 0.12fF
C17798 OR2X1_LOC_862/A OR2X1_LOC_810/A 0.77fF
C18358 OR2X1_LOC_574/A OR2X1_LOC_810/A 0.19fF
C18781 OR2X1_LOC_810/A OR2X1_LOC_203/Y 0.10fF
C23659 OR2X1_LOC_810/A OR2X1_LOC_844/B 0.38fF
C23685 OR2X1_LOC_810/A OR2X1_LOC_390/B 0.07fF
C27698 OR2X1_LOC_810/A OR2X1_LOC_206/A 0.03fF
C27952 OR2X1_LOC_810/A OR2X1_LOC_776/Y 0.07fF
C28305 OR2X1_LOC_810/A OR2X1_LOC_140/B 0.05fF
C31754 VDD OR2X1_LOC_810/A 2.30fF
C34058 OR2X1_LOC_241/Y OR2X1_LOC_810/A 0.10fF
C34301 OR2X1_LOC_216/A OR2X1_LOC_810/A 0.16fF
C35583 OR2X1_LOC_810/A OR2X1_LOC_561/Y 0.05fF
C38185 OR2X1_LOC_643/A OR2X1_LOC_810/A 0.05fF
C39625 OR2X1_LOC_810/A OR2X1_LOC_561/B 0.20fF
C40254 OR2X1_LOC_810/A OR2X1_LOC_523/Y 0.05fF
C41126 OR2X1_LOC_810/A OR2X1_LOC_737/A 0.10fF
C42538 OR2X1_LOC_844/a_8_216# OR2X1_LOC_810/A 0.13fF
C42975 OR2X1_LOC_404/Y OR2X1_LOC_810/A 0.10fF
C43220 OR2X1_LOC_810/A OR2X1_LOC_362/A 0.05fF
C44168 OR2X1_LOC_810/A OR2X1_LOC_574/a_8_216# 0.20fF
C46769 OR2X1_LOC_468/A OR2X1_LOC_810/A 0.04fF
C48195 OR2X1_LOC_624/A OR2X1_LOC_810/A 0.01fF
C51144 OR2X1_LOC_774/Y OR2X1_LOC_810/A 0.08fF
C53732 OR2X1_LOC_844/a_36_216# OR2X1_LOC_810/A 0.15fF
C55320 OR2X1_LOC_810/A OR2X1_LOC_575/A 0.06fF
C55336 OR2X1_LOC_810/A OR2X1_LOC_493/A 0.18fF
C55350 OR2X1_LOC_652/a_8_216# OR2X1_LOC_810/A 0.03fF
C57195 OR2X1_LOC_810/A VSS -4.69fF
C3363 OR2X1_LOC_574/A OR2X1_LOC_730/A 0.15fF
C5079 OR2X1_LOC_574/A OR2X1_LOC_539/Y 0.15fF
C5287 OR2X1_LOC_574/A OR2X1_LOC_319/Y 0.15fF
C5922 OR2X1_LOC_574/A OR2X1_LOC_575/A 0.01fF
C8061 OR2X1_LOC_632/a_8_216# OR2X1_LOC_574/A 0.02fF
C8986 OR2X1_LOC_574/A OR2X1_LOC_805/A 0.10fF
C9989 OR2X1_LOC_574/A OR2X1_LOC_228/Y 0.10fF
C13392 OR2X1_LOC_574/A AND2X1_LOC_679/a_8_24# 0.20fF
C18328 OR2X1_LOC_574/A OR2X1_LOC_510/Y 0.34fF
C18636 OR2X1_LOC_715/B OR2X1_LOC_574/A 0.01fF
C21248 OR2X1_LOC_574/A OR2X1_LOC_715/A 0.01fF
C21485 OR2X1_LOC_574/A OR2X1_LOC_318/B 0.03fF
C21697 OR2X1_LOC_538/A OR2X1_LOC_574/A 0.03fF
C25545 OR2X1_LOC_574/A OR2X1_LOC_203/Y 0.36fF
C30407 OR2X1_LOC_574/A OR2X1_LOC_390/B 0.10fF
C30695 OR2X1_LOC_574/A OR2X1_LOC_493/Y 0.05fF
C31686 OR2X1_LOC_175/Y OR2X1_LOC_574/A 0.15fF
C32669 OR2X1_LOC_574/A OR2X1_LOC_620/Y 0.07fF
C38503 VDD OR2X1_LOC_574/A 1.98fF
C39380 OR2X1_LOC_676/Y OR2X1_LOC_574/A 0.18fF
C40819 OR2X1_LOC_574/A OR2X1_LOC_241/Y 0.10fF
C48185 OR2X1_LOC_574/A OR2X1_LOC_737/A 0.10fF
C50186 OR2X1_LOC_574/A OR2X1_LOC_362/A 0.08fF
C51095 OR2X1_LOC_574/A OR2X1_LOC_574/a_8_216# 0.02fF
C53588 OR2X1_LOC_468/A OR2X1_LOC_574/A 0.03fF
C53717 OR2X1_LOC_574/A OR2X1_LOC_449/B 0.05fF
C54037 OR2X1_LOC_856/B OR2X1_LOC_574/A 0.07fF
C57556 OR2X1_LOC_574/A VSS 0.95fF
C92 OR2X1_LOC_362/A OR2X1_LOC_349/B 0.02fF
C224 OR2X1_LOC_858/B OR2X1_LOC_362/A 0.02fF
C4004 OR2X1_LOC_362/A OR2X1_LOC_140/B 0.01fF
C5508 OR2X1_LOC_343/B OR2X1_LOC_362/A 0.01fF
C7449 VDD OR2X1_LOC_362/A 0.39fF
C9189 OR2X1_LOC_359/A OR2X1_LOC_362/A 0.02fF
C10087 OR2X1_LOC_362/B OR2X1_LOC_362/A 0.04fF
C11685 OR2X1_LOC_362/A OR2X1_LOC_343/a_8_216# 0.01fF
C13961 OR2X1_LOC_643/A OR2X1_LOC_362/A 0.03fF
C18674 OR2X1_LOC_404/Y OR2X1_LOC_362/A 0.07fF
C19839 OR2X1_LOC_574/a_8_216# OR2X1_LOC_362/A 0.40fF
C28237 OR2X1_LOC_362/A OR2X1_LOC_349/A 0.02fF
C43105 OR2X1_LOC_348/Y OR2X1_LOC_362/A 0.09fF
C43114 OR2X1_LOC_349/a_8_216# OR2X1_LOC_362/A 0.01fF
C45298 OR2X1_LOC_850/a_8_216# OR2X1_LOC_362/A 0.01fF
C46602 OR2X1_LOC_114/B OR2X1_LOC_362/A 0.03fF
C53884 OR2X1_LOC_850/B OR2X1_LOC_362/A 0.01fF
C55455 OR2X1_LOC_362/A OR2X1_LOC_844/B 0.03fF
C55823 OR2X1_LOC_362/A OR2X1_LOC_493/Y 0.03fF
C56542 OR2X1_LOC_362/A VSS 0.45fF
C1497 OR2X1_LOC_473/Y OR2X1_LOC_228/Y 0.01fF
C9062 OR2X1_LOC_473/Y OR2X1_LOC_475/Y 0.02fF
C10188 OR2X1_LOC_715/B OR2X1_LOC_473/Y 0.03fF
C11217 OR2X1_LOC_473/Y OR2X1_LOC_786/Y 0.41fF
C24797 OR2X1_LOC_473/Y OR2X1_LOC_476/a_8_216# 0.04fF
C27926 OR2X1_LOC_473/Y OR2X1_LOC_392/B 0.38fF
C30116 VDD OR2X1_LOC_473/Y 0.22fF
C32682 OR2X1_LOC_216/A OR2X1_LOC_473/Y 0.01fF
C35724 OR2X1_LOC_473/Y OR2X1_LOC_201/Y 0.01fF
C35760 OR2X1_LOC_473/Y OR2X1_LOC_201/a_8_216# 0.01fF
C53698 OR2X1_LOC_473/Y OR2X1_LOC_493/A 0.80fF
C55778 OR2X1_LOC_201/A OR2X1_LOC_473/Y 0.05fF
C57379 OR2X1_LOC_473/Y VSS -0.24fF
C3698 OR2X1_LOC_813/Y AND2X1_LOC_216/A 0.01fF
C12776 AND2X1_LOC_216/A AND2X1_LOC_772/Y 0.01fF
C28180 AND2X1_LOC_573/A AND2X1_LOC_216/A 0.01fF
C29151 AND2X1_LOC_216/A AND2X1_LOC_647/Y 0.71fF
C31102 AND2X1_LOC_139/a_8_24# AND2X1_LOC_216/A 0.17fF
C36555 AND2X1_LOC_141/A AND2X1_LOC_216/A 0.23fF
C37480 OR2X1_LOC_131/Y AND2X1_LOC_216/A 0.10fF
C37787 VDD AND2X1_LOC_216/A 0.54fF
C37968 AND2X1_LOC_216/A OR2X1_LOC_67/Y 0.02fF
C40056 AND2X1_LOC_139/A AND2X1_LOC_216/A 0.02fF
C40447 AND2X1_LOC_116/Y AND2X1_LOC_216/A 0.24fF
C45782 AND2X1_LOC_216/A AND2X1_LOC_656/a_8_24# 0.22fF
C46531 AND2X1_LOC_139/B AND2X1_LOC_216/A 0.14fF
C56872 AND2X1_LOC_216/A VSS -0.28fF
C8371 OR2X1_LOC_261/Y AND2X1_LOC_789/Y 0.02fF
C19060 AND2X1_LOC_555/a_8_24# OR2X1_LOC_261/Y 0.01fF
C40350 OR2X1_LOC_481/Y OR2X1_LOC_261/Y 0.22fF
C42295 AND2X1_LOC_555/Y OR2X1_LOC_261/Y 0.80fF
C52866 AND2X1_LOC_259/Y OR2X1_LOC_261/Y 0.02fF
C55264 VDD OR2X1_LOC_261/Y 0.10fF
C57608 OR2X1_LOC_261/Y VSS 0.14fF
C15557 OR2X1_LOC_442/Y AND2X1_LOC_444/a_8_24# 0.23fF
C28281 VDD OR2X1_LOC_442/Y 0.12fF
C56737 OR2X1_LOC_442/Y VSS 0.06fF
C5457 VDD OR2X1_LOC_125/Y 0.12fF
C26053 OR2X1_LOC_125/Y AND2X1_LOC_128/a_8_24# 0.23fF
C28523 OR2X1_LOC_127/Y OR2X1_LOC_125/Y 0.04fF
C57125 OR2X1_LOC_125/Y VSS 0.06fF
C9305 AND2X1_LOC_391/Y OR2X1_LOC_127/Y 0.06fF
C13265 OR2X1_LOC_127/Y AND2X1_LOC_554/B 0.79fF
C39523 OR2X1_LOC_127/Y AND2X1_LOC_128/a_8_24# 0.05fF
C57852 OR2X1_LOC_127/Y VSS 0.11fF
C3952 VDD OR2X1_LOC_561/B 0.03fF
C5427 OR2X1_LOC_561/B OR2X1_LOC_561/A 0.06fF
C23195 OR2X1_LOC_774/Y OR2X1_LOC_561/B 0.50fF
C29414 OR2X1_LOC_859/a_8_216# OR2X1_LOC_561/B 0.01fF
C34101 OR2X1_LOC_561/a_8_216# OR2X1_LOC_561/B 0.04fF
C37099 OR2X1_LOC_859/A OR2X1_LOC_561/B 0.08fF
C38733 OR2X1_LOC_810/a_8_216# OR2X1_LOC_561/B 0.02fF
C38761 OR2X1_LOC_859/B OR2X1_LOC_561/B 0.04fF
C46070 OR2X1_LOC_862/A OR2X1_LOC_561/B 0.67fF
C50011 OR2X1_LOC_812/B OR2X1_LOC_561/B 0.18fF
C56351 OR2X1_LOC_561/B VSS -0.63fF
C33957 OR2X1_LOC_653/Y OR2X1_LOC_33/B 0.01fF
C36111 OR2X1_LOC_33/A OR2X1_LOC_33/B 0.07fF
C52885 OR2X1_LOC_33/B OR2X1_LOC_33/a_8_216# 0.05fF
C54567 OR2X1_LOC_476/B OR2X1_LOC_33/B 0.02fF
C56814 OR2X1_LOC_33/B VSS -0.20fF
C4169 OR2X1_LOC_184/Y OR2X1_LOC_183/Y 0.14fF
C5623 OR2X1_LOC_108/Y OR2X1_LOC_183/Y 0.01fF
C13038 AND2X1_LOC_717/B OR2X1_LOC_183/Y 0.07fF
C19757 AND2X1_LOC_540/a_8_24# OR2X1_LOC_183/Y 0.04fF
C24010 OR2X1_LOC_178/Y OR2X1_LOC_183/Y 0.18fF
C27425 OR2X1_LOC_280/Y OR2X1_LOC_183/Y 0.03fF
C31087 AND2X1_LOC_465/A OR2X1_LOC_183/Y 0.08fF
C41276 VDD OR2X1_LOC_183/Y 0.14fF
C45162 AND2X1_LOC_721/Y OR2X1_LOC_183/Y 0.02fF
C56378 OR2X1_LOC_183/Y VSS 0.16fF
C37912 VDD OR2X1_LOC_584/Y 0.08fF
C54233 OR2X1_LOC_583/Y OR2X1_LOC_584/Y 0.09fF
C56655 OR2X1_LOC_584/Y VSS 0.12fF
C23033 VDD OR2X1_LOC_7/Y 0.10fF
C48667 AND2X1_LOC_193/a_8_24# OR2X1_LOC_7/Y 0.09fF
C56884 OR2X1_LOC_7/Y VSS 0.33fF
C1796 AND2X1_LOC_724/A OR2X1_LOC_423/Y 0.09fF
C10227 OR2X1_LOC_424/Y OR2X1_LOC_423/Y 0.61fF
C21296 AND2X1_LOC_449/a_8_24# OR2X1_LOC_423/Y 0.23fF
C41205 AND2X1_LOC_703/Y OR2X1_LOC_423/Y 0.02fF
C43009 VDD OR2X1_LOC_423/Y 0.44fF
C52443 AND2X1_LOC_714/a_8_24# OR2X1_LOC_423/Y 0.01fF
C54174 AND2X1_LOC_605/Y OR2X1_LOC_423/Y 0.13fF
C56249 OR2X1_LOC_423/Y VSS 0.39fF
C596 OR2X1_LOC_555/A OR2X1_LOC_348/B 0.28fF
C14122 OR2X1_LOC_563/A OR2X1_LOC_348/B 0.03fF
C20960 OR2X1_LOC_348/a_8_216# OR2X1_LOC_348/B 0.06fF
C40369 VDD OR2X1_LOC_348/B 0.23fF
C51683 OR2X1_LOC_791/B OR2X1_LOC_348/B 0.03fF
C56304 OR2X1_LOC_348/B VSS -0.27fF
C2351 OR2X1_LOC_700/Y AND2X1_LOC_789/Y 0.02fF
C2826 AND2X1_LOC_259/Y AND2X1_LOC_789/Y 0.02fF
C5712 AND2X1_LOC_347/a_8_24# AND2X1_LOC_789/Y 0.02fF
C7736 AND2X1_LOC_792/a_36_24# AND2X1_LOC_789/Y 0.01fF
C7849 OR2X1_LOC_701/Y AND2X1_LOC_789/Y -0.02fF
C9959 AND2X1_LOC_191/B AND2X1_LOC_789/Y 0.07fF
C12486 AND2X1_LOC_710/Y AND2X1_LOC_789/Y 0.01fF
C13031 OR2X1_LOC_757/Y AND2X1_LOC_789/Y 0.02fF
C14124 AND2X1_LOC_791/a_8_24# AND2X1_LOC_789/Y 0.04fF
C16822 AND2X1_LOC_347/a_36_24# AND2X1_LOC_789/Y 0.01fF
C17994 AND2X1_LOC_711/a_8_24# AND2X1_LOC_789/Y 0.01fF
C19395 AND2X1_LOC_345/a_8_24# AND2X1_LOC_789/Y 0.01fF
C19639 AND2X1_LOC_792/B AND2X1_LOC_789/Y 0.03fF
C22531 AND2X1_LOC_792/Y AND2X1_LOC_789/Y 0.07fF
C22827 AND2X1_LOC_710/a_8_24# AND2X1_LOC_789/Y 0.02fF
C24095 AND2X1_LOC_711/Y AND2X1_LOC_789/Y 0.01fF
C25141 AND2X1_LOC_791/a_36_24# AND2X1_LOC_789/Y 0.01fF
C25153 OR2X1_LOC_759/Y AND2X1_LOC_789/Y 0.02fF
C25215 AND2X1_LOC_555/a_8_24# AND2X1_LOC_789/Y 0.01fF
C25550 AND2X1_LOC_789/Y AND2X1_LOC_793/a_8_24# 0.05fF
C26393 AND2X1_LOC_710/a_36_24# AND2X1_LOC_789/Y 0.01fF
C30388 AND2X1_LOC_345/a_36_24# AND2X1_LOC_789/Y 0.01fF
C36168 AND2X1_LOC_555/a_36_24# AND2X1_LOC_789/Y 0.01fF
C37436 AND2X1_LOC_347/B AND2X1_LOC_789/Y 0.02fF
C41656 AND2X1_LOC_792/a_8_24# AND2X1_LOC_789/Y -0.02fF
C45657 AND2X1_LOC_347/Y AND2X1_LOC_789/Y 0.22fF
C46100 OR2X1_LOC_755/Y AND2X1_LOC_789/Y 0.04fF
C46636 OR2X1_LOC_481/Y AND2X1_LOC_789/Y 0.02fF
C48655 AND2X1_LOC_555/Y AND2X1_LOC_789/Y 0.08fF
C50929 OR2X1_LOC_297/Y AND2X1_LOC_789/Y 0.01fF
C50938 AND2X1_LOC_345/Y AND2X1_LOC_789/Y 0.40fF
C56358 AND2X1_LOC_789/Y VSS -2.29fF
C3201 OR2X1_LOC_555/A OR2X1_LOC_259/B 0.09fF
C27746 OR2X1_LOC_259/a_8_216# OR2X1_LOC_259/B 0.06fF
C38734 OR2X1_LOC_555/B OR2X1_LOC_259/B 0.17fF
C55818 OR2X1_LOC_259/B OR2X1_LOC_555/a_8_216# 0.47fF
C56453 OR2X1_LOC_259/B VSS 0.31fF
C6209 OR2X1_LOC_318/B OR2X1_LOC_228/Y 0.01fF
C6513 OR2X1_LOC_76/A OR2X1_LOC_318/B 0.03fF
C8041 OR2X1_LOC_318/B OR2X1_LOC_716/a_8_216# 0.01fF
C9871 OR2X1_LOC_486/Y OR2X1_LOC_318/B 0.12fF
C13069 OR2X1_LOC_318/B OR2X1_LOC_241/B 0.18fF
C16270 OR2X1_LOC_851/A OR2X1_LOC_318/B 0.12fF
C16748 OR2X1_LOC_605/A OR2X1_LOC_318/B 0.21fF
C17997 OR2X1_LOC_841/B OR2X1_LOC_318/B 0.01fF
C22344 OR2X1_LOC_605/B OR2X1_LOC_318/B 0.29fF
C24621 OR2X1_LOC_318/B OR2X1_LOC_723/B 0.02fF
C27785 OR2X1_LOC_605/a_8_216# OR2X1_LOC_318/B 0.01fF
C29701 OR2X1_LOC_318/B OR2X1_LOC_605/Y 0.02fF
C31076 OR2X1_LOC_776/Y OR2X1_LOC_318/B 0.05fF
C31149 OR2X1_LOC_76/Y OR2X1_LOC_318/B 0.11fF
C31864 OR2X1_LOC_787/a_8_216# OR2X1_LOC_318/B 0.48fF
C32499 OR2X1_LOC_318/B OR2X1_LOC_374/Y 0.03fF
C34878 VDD OR2X1_LOC_318/B 0.05fF
C36972 OR2X1_LOC_840/A OR2X1_LOC_318/B 0.03fF
C40917 OR2X1_LOC_440/A OR2X1_LOC_318/B 0.03fF
C41292 OR2X1_LOC_778/Y OR2X1_LOC_318/B 0.05fF
C42552 OR2X1_LOC_787/B OR2X1_LOC_318/B 0.16fF
C46810 OR2X1_LOC_318/B OR2X1_LOC_776/A 0.02fF
C47259 OR2X1_LOC_318/B OR2X1_LOC_593/B 0.03fF
C52096 OR2X1_LOC_787/Y OR2X1_LOC_318/B 0.01fF
C56485 OR2X1_LOC_318/B VSS 0.56fF
C1656 OR2X1_LOC_702/A OR2X1_LOC_676/Y 0.01fF
C2500 OR2X1_LOC_676/Y OR2X1_LOC_194/Y 0.19fF
C18943 OR2X1_LOC_676/Y OR2X1_LOC_702/a_8_216# 0.01fF
C19836 OR2X1_LOC_676/Y OR2X1_LOC_678/Y 0.14fF
C21646 OR2X1_LOC_644/B OR2X1_LOC_676/Y 0.76fF
C22670 OR2X1_LOC_676/Y OR2X1_LOC_194/a_8_216# 0.02fF
C24351 OR2X1_LOC_676/Y OR2X1_LOC_228/Y 0.43fF
C24479 OR2X1_LOC_676/Y OR2X1_LOC_702/a_36_216# 0.01fF
C28111 OR2X1_LOC_676/Y OR2X1_LOC_194/a_36_216# 0.01fF
C31369 OR2X1_LOC_676/Y OR2X1_LOC_193/A 0.03fF
C35418 OR2X1_LOC_676/Y OR2X1_LOC_715/A 0.03fF
C36701 OR2X1_LOC_676/Y OR2X1_LOC_623/B 0.07fF
C39012 OR2X1_LOC_676/Y OR2X1_LOC_196/B 0.08fF
C45350 OR2X1_LOC_676/Y OR2X1_LOC_194/B 0.01fF
C53019 VDD OR2X1_LOC_676/Y 0.67fF
C57594 OR2X1_LOC_676/Y VSS 0.43fF
C2120 OR2X1_LOC_545/A OR2X1_LOC_545/B 0.16fF
C8608 OR2X1_LOC_545/A OR2X1_LOC_545/a_8_216# 0.47fF
C22143 OR2X1_LOC_545/A OR2X1_LOC_471/Y 0.02fF
C36088 OR2X1_LOC_545/A OR2X1_LOC_551/B 0.05fF
C57752 OR2X1_LOC_545/A VSS 0.04fF
C45710 AND2X1_LOC_7/Y AND2X1_LOC_52/Y 0.04fF
C51327 OR2X1_LOC_228/a_8_216# AND2X1_LOC_52/Y 0.47fF
C55116 OR2X1_LOC_651/A AND2X1_LOC_52/Y 0.09fF
C56245 AND2X1_LOC_52/Y VSS 0.26fF
C14560 OR2X1_LOC_782/B OR2X1_LOC_781/Y 0.45fF
C25592 OR2X1_LOC_782/B OR2X1_LOC_782/a_8_216# 0.47fF
C57879 OR2X1_LOC_782/B VSS 0.16fF
C8287 OR2X1_LOC_523/B OR2X1_LOC_392/B 0.04fF
C10450 OR2X1_LOC_523/B VDD -0.00fF
C11168 OR2X1_LOC_523/B OR2X1_LOC_523/A 0.16fF
C21664 OR2X1_LOC_523/B OR2X1_LOC_404/Y 0.01fF
C27730 OR2X1_LOC_523/B OR2X1_LOC_523/a_8_216# 0.47fF
C57914 OR2X1_LOC_523/B VSS 0.16fF
C31494 OR2X1_LOC_636/A OR2X1_LOC_636/B 1.24fF
C48277 OR2X1_LOC_636/B OR2X1_LOC_636/a_8_216# 0.01fF
C57348 OR2X1_LOC_636/B VSS -0.47fF
C3245 VDD OR2X1_LOC_542/B 0.07fF
C16074 OR2X1_LOC_542/B OR2X1_LOC_465/B 0.03fF
C28652 OR2X1_LOC_542/B OR2X1_LOC_542/a_8_216# 0.06fF
C32841 OR2X1_LOC_542/B OR2X1_LOC_563/A 0.07fF
C37101 OR2X1_LOC_190/A OR2X1_LOC_542/B 3.53fF
C41873 OR2X1_LOC_147/B OR2X1_LOC_542/B 13.10fF
C57372 OR2X1_LOC_542/B VSS 0.42fF
C9686 OR2X1_LOC_792/B OR2X1_LOC_792/Y 0.89fF
C25887 OR2X1_LOC_792/B OR2X1_LOC_792/a_8_216# 0.01fF
C29191 OR2X1_LOC_791/B OR2X1_LOC_792/B 0.06fF
C57826 OR2X1_LOC_792/B VSS 0.10fF
C30012 OR2X1_LOC_710/A OR2X1_LOC_705/Y 0.03fF
C30309 OR2X1_LOC_710/B OR2X1_LOC_710/A 0.16fF
C57971 OR2X1_LOC_710/A VSS 0.18fF
C10049 AND2X1_LOC_334/Y AND2X1_LOC_338/a_36_24# 0.01fF
C17238 VDD AND2X1_LOC_334/Y 0.01fF
C19099 AND2X1_LOC_334/Y AND2X1_LOC_640/Y 1.13fF
C19132 AND2X1_LOC_334/Y OR2X1_LOC_416/Y 0.01fF
C42920 AND2X1_LOC_334/Y AND2X1_LOC_476/A 0.04fF
C49674 AND2X1_LOC_334/Y AND2X1_LOC_338/a_8_24# 0.03fF
C57354 AND2X1_LOC_334/Y VSS 0.11fF
C24589 VDD AND2X1_LOC_839/B 0.24fF
C25622 AND2X1_LOC_839/A AND2X1_LOC_839/B 0.10fF
C53190 AND2X1_LOC_839/B AND2X1_LOC_839/a_8_24# 0.19fF
C56932 AND2X1_LOC_839/B VSS 0.07fF
C754 AND2X1_LOC_240/Y AND2X1_LOC_243/Y 0.01fF
C5134 AND2X1_LOC_240/Y AND2X1_LOC_243/a_8_24# 0.11fF
C15815 AND2X1_LOC_835/a_8_24# AND2X1_LOC_240/Y 0.06fF
C20363 VDD AND2X1_LOC_240/Y 0.07fF
C21430 AND2X1_LOC_839/A AND2X1_LOC_240/Y 0.83fF
C56601 AND2X1_LOC_240/Y VSS 0.15fF
C6937 AND2X1_LOC_462/Y OR2X1_LOC_416/Y 0.01fF
C12036 AND2X1_LOC_34/a_8_24# AND2X1_LOC_462/Y 0.11fF
C25279 AND2X1_LOC_462/Y AND2X1_LOC_472/a_8_24# 0.09fF
C30740 AND2X1_LOC_462/Y AND2X1_LOC_476/A 0.04fF
C35718 AND2X1_LOC_34/Y AND2X1_LOC_462/Y 0.89fF
C51670 AND2X1_LOC_462/Y OR2X1_LOC_27/Y 0.30fF
C56991 AND2X1_LOC_462/Y VSS 0.22fF
C22445 OR2X1_LOC_730/a_8_216# OR2X1_LOC_730/A 0.39fF
C34924 OR2X1_LOC_730/B OR2X1_LOC_730/A 0.04fF
C56279 OR2X1_LOC_730/A VSS 0.18fF
C10955 OR2X1_LOC_856/A OR2X1_LOC_856/a_8_216# 0.18fF
C16770 VDD OR2X1_LOC_856/A 0.06fF
C32040 OR2X1_LOC_856/B OR2X1_LOC_856/A 0.14fF
C57731 OR2X1_LOC_856/A VSS 0.17fF
C6078 OR2X1_LOC_550/a_8_216# OR2X1_LOC_550/A 0.39fF
C32761 OR2X1_LOC_550/B OR2X1_LOC_550/A 0.05fF
C56305 OR2X1_LOC_550/A VSS 0.18fF
C4006 OR2X1_LOC_174/A OR2X1_LOC_339/A 0.11fF
C22241 OR2X1_LOC_339/A OR2X1_LOC_174/a_8_216# 0.01fF
C23934 OR2X1_LOC_175/Y OR2X1_LOC_339/A 0.01fF
C24476 OR2X1_LOC_333/B OR2X1_LOC_339/A 0.02fF
C29323 OR2X1_LOC_339/A OR2X1_LOC_174/Y 0.07fF
C30676 VDD OR2X1_LOC_339/A 0.08fF
C53409 OR2X1_LOC_539/Y OR2X1_LOC_339/A 0.73fF
C54645 OR2X1_LOC_61/Y OR2X1_LOC_339/A 0.18fF
C56337 OR2X1_LOC_339/A VSS 0.07fF
C1534 OR2X1_LOC_715/B OR2X1_LOC_201/A 0.08fF
C2468 OR2X1_LOC_715/B OR2X1_LOC_805/A 0.07fF
C3503 OR2X1_LOC_715/B OR2X1_LOC_228/Y 0.10fF
C6838 OR2X1_LOC_715/B AND2X1_LOC_679/a_8_24# 0.02fF
C13259 OR2X1_LOC_715/B OR2X1_LOC_786/Y 0.03fF
C14707 OR2X1_LOC_715/B OR2X1_LOC_715/A 0.21fF
C15121 OR2X1_LOC_715/B OR2X1_LOC_538/A 0.01fF
C15961 OR2X1_LOC_715/B OR2X1_LOC_623/B 0.07fF
C16330 OR2X1_LOC_715/B OR2X1_LOC_140/A 0.17fF
C21620 OR2X1_LOC_715/B OR2X1_LOC_653/A 0.03fF
C23999 OR2X1_LOC_715/B OR2X1_LOC_390/B 0.10fF
C25247 OR2X1_LOC_715/B OR2X1_LOC_175/Y 0.18fF
C26188 OR2X1_LOC_715/B OR2X1_LOC_620/Y 0.33fF
C26411 OR2X1_LOC_715/B OR2X1_LOC_560/A 0.03fF
C27999 OR2X1_LOC_715/B OR2X1_LOC_206/A 0.05fF
C28248 OR2X1_LOC_715/B OR2X1_LOC_776/Y 0.38fF
C28938 OR2X1_LOC_715/B AND2X1_LOC_679/a_36_24# 0.01fF
C31995 OR2X1_LOC_715/B VDD 1.93fF
C34340 OR2X1_LOC_715/B OR2X1_LOC_241/Y 0.98fF
C34587 OR2X1_LOC_715/B OR2X1_LOC_216/A 0.07fF
C36778 OR2X1_LOC_715/B OR2X1_LOC_702/A 0.12fF
C37138 OR2X1_LOC_715/B OR2X1_LOC_623/a_8_216# 0.28fF
C37648 OR2X1_LOC_715/B OR2X1_LOC_201/Y 0.07fF
C37729 OR2X1_LOC_715/B OR2X1_LOC_201/a_8_216# 0.24fF
C41408 OR2X1_LOC_715/B OR2X1_LOC_737/A 0.07fF
C44836 OR2X1_LOC_715/B OR2X1_LOC_785/a_8_216# 0.30fF
C47580 OR2X1_LOC_715/B OR2X1_LOC_856/B 0.10fF
C48460 OR2X1_LOC_715/B OR2X1_LOC_624/A 0.11fF
C51175 OR2X1_LOC_715/B OR2X1_LOC_715/a_8_216# 0.02fF
C54247 OR2X1_LOC_715/B OR2X1_LOC_702/a_8_216# 0.03fF
C54744 OR2X1_LOC_715/B OR2X1_LOC_539/Y 0.41fF
C55112 OR2X1_LOC_715/B OR2X1_LOC_678/Y 0.01fF
C56020 OR2X1_LOC_715/B OR2X1_LOC_61/Y 0.23fF
C58023 OR2X1_LOC_715/B VSS 0.83fF
C2376 OR2X1_LOC_516/Y OR2X1_LOC_91/Y 0.42fF
C2474 OR2X1_LOC_516/Y AND2X1_LOC_574/A 0.01fF
C4449 OR2X1_LOC_516/Y OR2X1_LOC_497/Y 0.02fF
C6673 OR2X1_LOC_516/Y AND2X1_LOC_675/A 0.07fF
C9518 OR2X1_LOC_516/Y AND2X1_LOC_242/a_8_24# 0.02fF
C10797 OR2X1_LOC_516/Y OR2X1_LOC_528/Y 0.03fF
C13774 OR2X1_LOC_516/Y AND2X1_LOC_499/a_8_24# 0.02fF
C13786 OR2X1_LOC_516/Y AND2X1_LOC_658/B 0.05fF
C15023 OR2X1_LOC_516/Y AND2X1_LOC_244/A 0.04fF
C15041 OR2X1_LOC_516/Y OR2X1_LOC_108/Y 0.17fF
C15397 OR2X1_LOC_516/Y OR2X1_LOC_373/Y 0.07fF
C17948 OR2X1_LOC_516/Y AND2X1_LOC_242/B 0.09fF
C18482 OR2X1_LOC_516/Y OR2X1_LOC_495/Y 0.03fF
C19258 OR2X1_LOC_516/Y AND2X1_LOC_785/Y 0.11fF
C19286 OR2X1_LOC_516/Y AND2X1_LOC_500/B 0.04fF
C23986 OR2X1_LOC_516/Y AND2X1_LOC_778/Y 3.05fF
C24798 OR2X1_LOC_516/Y AND2X1_LOC_786/Y 0.07fF
C30282 OR2X1_LOC_516/Y AND2X1_LOC_784/Y 0.37fF
C32061 OR2X1_LOC_516/Y AND2X1_LOC_830/a_8_24# 0.02fF
C34111 OR2X1_LOC_516/Y AND2X1_LOC_508/A 0.05fF
C34911 OR2X1_LOC_516/Y AND2X1_LOC_564/B 0.07fF
C39238 OR2X1_LOC_516/Y AND2X1_LOC_500/a_8_24# 0.04fF
C42722 OR2X1_LOC_516/Y OR2X1_LOC_239/Y 0.04fF
C43177 OR2X1_LOC_516/Y AND2X1_LOC_842/B 0.03fF
C43838 OR2X1_LOC_516/Y AND2X1_LOC_785/A 0.15fF
C43923 OR2X1_LOC_516/Y AND2X1_LOC_658/A 0.07fF
C45193 OR2X1_LOC_516/Y AND2X1_LOC_476/Y 0.07fF
C47882 OR2X1_LOC_516/Y AND2X1_LOC_500/Y 0.24fF
C50854 OR2X1_LOC_516/Y VDD 0.40fF
C54568 OR2X1_LOC_516/Y AND2X1_LOC_721/Y 0.03fF
C54599 OR2X1_LOC_516/Y OR2X1_LOC_482/Y 0.15fF
C58126 OR2X1_LOC_516/Y VSS 0.18fF
C624 OR2X1_LOC_787/a_8_216# OR2X1_LOC_787/B 0.05fF
C3664 VDD OR2X1_LOC_787/B 0.16fF
C34538 OR2X1_LOC_486/Y OR2X1_LOC_787/B 0.22fF
C56650 OR2X1_LOC_787/B VSS -0.15fF
C41510 OR2X1_LOC_792/Y OR2X1_LOC_286/Y 0.04fF
C53606 OR2X1_LOC_286/Y OR2X1_LOC_288/a_8_216# 0.39fF
C57146 OR2X1_LOC_286/Y VSS 0.17fF
C10271 OR2X1_LOC_772/B OR2X1_LOC_772/Y 0.73fF
C22012 VDD OR2X1_LOC_772/B -0.00fF
C41121 OR2X1_LOC_774/Y OR2X1_LOC_772/B 0.04fF
C45456 OR2X1_LOC_772/B OR2X1_LOC_772/a_8_216# 0.01fF
C57268 OR2X1_LOC_772/B VSS 0.15fF
C15440 OR2X1_LOC_351/B OR2X1_LOC_338/B 0.74fF
C55021 OR2X1_LOC_338/a_8_216# OR2X1_LOC_338/B 0.06fF
C56301 OR2X1_LOC_338/B VSS 0.11fF
C442 OR2X1_LOC_714/A OR2X1_LOC_308/Y 0.03fF
C22640 OR2X1_LOC_703/Y OR2X1_LOC_714/A 0.06fF
C25212 VDD OR2X1_LOC_714/A -0.00fF
C33576 OR2X1_LOC_714/a_8_216# OR2X1_LOC_714/A 0.39fF
C55295 OR2X1_LOC_724/A OR2X1_LOC_714/A 0.01fF
C56422 OR2X1_LOC_714/A VSS 0.18fF
C13505 OR2X1_LOC_446/Y OR2X1_LOC_712/B 0.01fF
C23453 VDD OR2X1_LOC_446/Y 0.23fF
C38259 OR2X1_LOC_446/Y OR2X1_LOC_449/B 0.12fF
C54650 OR2X1_LOC_446/Y OR2X1_LOC_783/A 0.03fF
C57383 OR2X1_LOC_446/Y VSS 0.37fF
C5095 VDD OR2X1_LOC_227/Y 0.19fF
C15372 OR2X1_LOC_509/A OR2X1_LOC_227/Y 0.11fF
C19805 OR2X1_LOC_227/Y AND2X1_LOC_88/Y 0.06fF
C25307 OR2X1_LOC_227/Y OR2X1_LOC_340/a_8_216# 0.18fF
C27030 OR2X1_LOC_227/Y OR2X1_LOC_641/B 0.01fF
C38599 OR2X1_LOC_509/a_8_216# OR2X1_LOC_227/Y 0.05fF
C55578 OR2X1_LOC_227/Y OR2X1_LOC_560/A 0.34fF
C56481 OR2X1_LOC_227/Y VSS 0.37fF
C1756 AND2X1_LOC_149/a_8_24# OR2X1_LOC_679/B 0.20fF
C4514 OR2X1_LOC_679/a_8_216# OR2X1_LOC_679/B 0.01fF
C11095 AND2X1_LOC_728/a_8_24# OR2X1_LOC_679/B 0.09fF
C11361 VDD OR2X1_LOC_679/B 0.21fF
C15597 OR2X1_LOC_679/Y OR2X1_LOC_679/B 0.20fF
C17661 OR2X1_LOC_679/B AND2X1_LOC_213/B 0.01fF
C33171 OR2X1_LOC_679/A OR2X1_LOC_679/B 0.33fF
C46869 AND2X1_LOC_148/Y OR2X1_LOC_679/B 0.05fF
C56962 OR2X1_LOC_679/B VSS -0.08fF
C4824 OR2X1_LOC_134/Y AND2X1_LOC_772/B 0.01fF
C9577 OR2X1_LOC_132/Y OR2X1_LOC_134/Y 0.11fF
C14732 OR2X1_LOC_134/Y AND2X1_LOC_560/B 0.15fF
C19500 OR2X1_LOC_134/Y AND2X1_LOC_656/Y 0.03fF
C40853 AND2X1_LOC_392/A OR2X1_LOC_134/Y 0.03fF
C44781 OR2X1_LOC_134/Y VDD 0.11fF
C48377 OR2X1_LOC_134/Y OR2X1_LOC_103/Y 0.10fF
C50022 OR2X1_LOC_134/Y AND2X1_LOC_768/a_8_24# 0.01fF
C50446 OR2X1_LOC_134/Y AND2X1_LOC_541/Y 1.17fF
C58024 OR2X1_LOC_134/Y VSS 0.19fF
C329 OR2X1_LOC_34/B OR2X1_LOC_34/A 0.16fF
C9741 OR2X1_LOC_476/B OR2X1_LOC_34/A -0.00fF
C56753 OR2X1_LOC_34/A VSS -0.08fF
C15849 VDD OR2X1_LOC_759/Y 0.12fF
C28606 AND2X1_LOC_711/a_8_24# OR2X1_LOC_759/Y 0.23fF
C30204 AND2X1_LOC_792/B OR2X1_LOC_759/Y 0.10fF
C34600 AND2X1_LOC_711/Y OR2X1_LOC_759/Y 0.01fF
C56395 OR2X1_LOC_759/Y VSS 0.10fF
C6782 AND2X1_LOC_391/Y AND2X1_LOC_128/a_8_24# 0.01fF
C17852 AND2X1_LOC_391/Y AND2X1_LOC_128/a_36_24# 0.05fF
C29477 AND2X1_LOC_555/Y AND2X1_LOC_391/Y 0.01fF
C36415 AND2X1_LOC_391/Y AND2X1_LOC_554/B 0.29fF
C38369 AND2X1_LOC_392/A AND2X1_LOC_391/Y 0.02fF
C42259 AND2X1_LOC_391/Y VDD 0.08fF
C43601 AND2X1_LOC_391/Y AND2X1_LOC_392/a_8_24# 0.01fF
C53283 AND2X1_LOC_391/Y AND2X1_LOC_721/A 0.03fF
C58022 AND2X1_LOC_391/Y VSS 0.44fF
C19101 OR2X1_LOC_394/Y OR2X1_LOC_393/Y 0.10fF
C32964 VDD OR2X1_LOC_393/Y 0.07fF
C56586 OR2X1_LOC_393/Y VSS 0.22fF
C8213 OR2X1_LOC_859/B OR2X1_LOC_859/A 0.35fF
C30904 VDD OR2X1_LOC_859/B 0.06fF
C50331 OR2X1_LOC_774/Y OR2X1_LOC_859/B 0.04fF
C57486 OR2X1_LOC_859/B VSS 0.18fF
C1550 OR2X1_LOC_486/B OR2X1_LOC_726/a_8_216# 0.47fF
C15390 OR2X1_LOC_486/a_8_216# OR2X1_LOC_486/B 0.05fF
C16355 OR2X1_LOC_486/B OR2X1_LOC_550/B 0.34fF
C26277 OR2X1_LOC_486/B OR2X1_LOC_726/A 0.08fF
C48853 OR2X1_LOC_486/B OR2X1_LOC_731/A 0.01fF
C56949 OR2X1_LOC_486/B VSS -0.05fF
C183 OR2X1_LOC_507/B OR2X1_LOC_508/Y 0.01fF
C2575 OR2X1_LOC_507/B OR2X1_LOC_510/Y 0.01fF
C7090 OR2X1_LOC_507/B OR2X1_LOC_507/A 0.18fF
C11265 OR2X1_LOC_507/B OR2X1_LOC_510/a_8_216# 0.49fF
C11346 OR2X1_LOC_510/A OR2X1_LOC_507/B 0.36fF
C29211 OR2X1_LOC_507/a_8_216# OR2X1_LOC_507/B 0.01fF
C29291 OR2X1_LOC_507/B OR2X1_LOC_643/A 0.03fF
C57626 OR2X1_LOC_507/B VSS 0.20fF
C11702 OR2X1_LOC_546/B OR2X1_LOC_546/A 0.16fF
C36330 OR2X1_LOC_149/B OR2X1_LOC_546/B 0.10fF
C39232 OR2X1_LOC_546/B OR2X1_LOC_546/a_8_216# 0.47fF
C57679 OR2X1_LOC_546/B VSS 0.16fF
C927 OR2X1_LOC_404/Y OR2X1_LOC_720/A 0.01fF
C33045 OR2X1_LOC_720/A OR2X1_LOC_721/Y 0.01fF
C45817 VDD OR2X1_LOC_720/A -0.00fF
C47764 OR2X1_LOC_720/A OR2X1_LOC_720/a_8_216# 0.47fF
C56747 OR2X1_LOC_720/A VSS 0.15fF
C7700 OR2X1_LOC_149/B OR2X1_LOC_546/A 0.13fF
C45603 VDD OR2X1_LOC_546/A 0.21fF
C56374 OR2X1_LOC_546/A VSS 0.02fF
C25732 OR2X1_LOC_602/A OR2X1_LOC_390/B 0.14fF
C28916 OR2X1_LOC_602/a_8_216# OR2X1_LOC_602/A 0.47fF
C56863 OR2X1_LOC_602/A VSS 0.15fF
C32098 AND2X1_LOC_719/Y AND2X1_LOC_287/Y 0.02fF
C43673 VDD AND2X1_LOC_287/Y 0.02fF
C46412 AND2X1_LOC_287/Y AND2X1_LOC_288/a_8_24# 0.01fF
C51964 AND2X1_LOC_287/Y AND2X1_LOC_806/A 0.16fF
C56553 AND2X1_LOC_287/Y VSS 0.13fF
C7049 AND2X1_LOC_719/Y AND2X1_LOC_843/Y -0.05fF
C18575 VDD AND2X1_LOC_843/Y 0.01fF
C19072 AND2X1_LOC_486/Y AND2X1_LOC_843/Y 0.39fF
C22939 AND2X1_LOC_843/Y AND2X1_LOC_850/A 0.31fF
C25856 AND2X1_LOC_843/Y AND2X1_LOC_850/Y 0.01fF
C52310 AND2X1_LOC_843/Y AND2X1_LOC_850/a_8_24# 0.09fF
C57346 AND2X1_LOC_843/Y VSS 0.02fF
C9522 OR2X1_LOC_349/B OR2X1_LOC_349/A 0.10fF
C24381 OR2X1_LOC_348/Y OR2X1_LOC_349/B 0.08fF
C24384 OR2X1_LOC_349/a_8_216# OR2X1_LOC_349/B 0.01fF
C44741 VDD OR2X1_LOC_349/B 0.06fF
C46530 OR2X1_LOC_359/A OR2X1_LOC_349/B 0.04fF
C56386 OR2X1_LOC_349/B VSS 0.08fF
C5183 AND2X1_LOC_654/B OR2X1_LOC_172/Y 0.74fF
C37403 VDD OR2X1_LOC_172/Y 0.35fF
C55019 OR2X1_LOC_45/Y OR2X1_LOC_172/Y 0.20fF
C56381 OR2X1_LOC_172/Y VSS -0.20fF
C27587 AND2X1_LOC_508/A OR2X1_LOC_239/Y 0.01fF
C32726 AND2X1_LOC_500/a_8_24# OR2X1_LOC_239/Y 0.01fF
C37246 AND2X1_LOC_658/A OR2X1_LOC_239/Y 0.03fF
C41078 AND2X1_LOC_500/Y OR2X1_LOC_239/Y 0.01fF
C44122 VDD OR2X1_LOC_239/Y 0.12fF
C54086 OR2X1_LOC_497/Y OR2X1_LOC_239/Y 0.16fF
C56846 OR2X1_LOC_239/Y VSS 0.16fF
C31012 OR2X1_LOC_822/Y AND2X1_LOC_835/a_8_24# 0.23fF
C35395 VDD OR2X1_LOC_822/Y 0.14fF
C57736 OR2X1_LOC_822/Y VSS 0.07fF
C574 OR2X1_LOC_766/Y AND2X1_LOC_770/a_8_24# 0.01fF
C11670 OR2X1_LOC_766/Y AND2X1_LOC_771/B 0.78fF
C32854 VDD OR2X1_LOC_766/Y 0.04fF
C56616 OR2X1_LOC_766/Y VSS 0.08fF
C3744 OR2X1_LOC_91/Y VDD 0.50fF
C3842 OR2X1_LOC_91/Y OR2X1_LOC_315/Y 0.27fF
C4191 OR2X1_LOC_91/Y AND2X1_LOC_486/Y 0.07fF
C7164 OR2X1_LOC_91/Y OR2X1_LOC_103/Y 0.03fF
C8176 OR2X1_LOC_91/Y AND2X1_LOC_523/Y 5.61fF
C15554 OR2X1_LOC_91/Y AND2X1_LOC_787/A 0.85fF
C15799 OR2X1_LOC_91/Y AND2X1_LOC_675/A 0.32fF
C18679 OR2X1_LOC_91/Y AND2X1_LOC_716/Y 0.01fF
C18771 OR2X1_LOC_91/Y OR2X1_LOC_312/Y 0.03fF
C21418 OR2X1_LOC_91/Y AND2X1_LOC_440/a_8_24# 0.03fF
C22749 OR2X1_LOC_91/Y OR2X1_LOC_437/Y 0.40fF
C24167 OR2X1_LOC_91/Y OR2X1_LOC_108/Y 0.07fF
C24515 OR2X1_LOC_91/Y OR2X1_LOC_373/Y 0.14fF
C25070 OR2X1_LOC_91/Y OR2X1_LOC_109/Y 0.18fF
C25854 OR2X1_LOC_91/Y AND2X1_LOC_722/A 0.01fF
C27419 OR2X1_LOC_91/Y AND2X1_LOC_543/Y 0.03fF
C29163 OR2X1_LOC_91/Y AND2X1_LOC_180/a_8_24# 0.02fF
C29561 OR2X1_LOC_91/Y AND2X1_LOC_445/a_8_24# 0.02fF
C29677 OR2X1_LOC_91/Y AND2X1_LOC_717/Y 0.01fF
C29730 OR2X1_LOC_91/Y AND2X1_LOC_560/B 0.07fF
C31285 OR2X1_LOC_91/Y AND2X1_LOC_443/a_8_24# -0.00fF
C32972 OR2X1_LOC_91/Y AND2X1_LOC_778/Y 0.02fF
C33800 OR2X1_LOC_91/Y AND2X1_LOC_786/Y 0.07fF
C34641 OR2X1_LOC_91/Y AND2X1_LOC_182/A 0.02fF
C37553 OR2X1_LOC_176/Y OR2X1_LOC_91/Y 0.01fF
C38459 OR2X1_LOC_91/Y AND2X1_LOC_784/a_8_24# 0.02fF
C38497 OR2X1_LOC_91/Y AND2X1_LOC_471/Y 0.02fF
C39317 AND2X1_LOC_784/Y OR2X1_LOC_91/Y 0.01fF
C39570 OR2X1_LOC_91/Y AND2X1_LOC_851/B 0.07fF
C40123 OR2X1_LOC_91/Y AND2X1_LOC_243/Y 0.02fF
C41113 OR2X1_LOC_91/Y AND2X1_LOC_468/B 0.01fF
C42367 OR2X1_LOC_91/Y OR2X1_LOC_178/Y 0.03fF
C44701 OR2X1_LOC_91/Y AND2X1_LOC_845/Y 0.05fF
C45072 OR2X1_LOC_91/Y AND2X1_LOC_784/A 0.84fF
C46422 OR2X1_LOC_91/Y AND2X1_LOC_211/B 0.58fF
C46767 OR2X1_LOC_91/Y AND2X1_LOC_474/A 0.02fF
C48482 OR2X1_LOC_91/Y AND2X1_LOC_719/Y 0.06fF
C48904 OR2X1_LOC_91/Y AND2X1_LOC_561/B 0.03fF
C49382 OR2X1_LOC_91/Y AND2X1_LOC_553/A 0.03fF
C49679 OR2X1_LOC_91/Y AND2X1_LOC_465/A 0.07fF
C49855 OR2X1_LOC_91/Y OR2X1_LOC_237/Y 0.06fF
C50259 OR2X1_LOC_91/Y AND2X1_LOC_573/A 0.07fF
C54327 OR2X1_LOC_91/Y AND2X1_LOC_476/Y 0.09fF
C58089 OR2X1_LOC_91/Y VSS 0.34fF
C16816 OR2X1_LOC_132/Y VDD 0.17fF
C47772 OR2X1_LOC_132/Y AND2X1_LOC_656/Y 0.01fF
C58098 OR2X1_LOC_132/Y VSS 0.14fF
C5983 OR2X1_LOC_646/A OR2X1_LOC_647/B 0.01fF
C17071 OR2X1_LOC_646/a_8_216# OR2X1_LOC_647/B 0.01fF
C21671 VDD OR2X1_LOC_647/B 0.23fF
C28123 OR2X1_LOC_647/A OR2X1_LOC_647/B 0.25fF
C38689 OR2X1_LOC_647/a_8_216# OR2X1_LOC_647/B 0.04fF
C56869 OR2X1_LOC_647/B VSS 0.30fF
C2480 AND2X1_LOC_810/A OR2X1_LOC_312/Y 0.03fF
C5368 OR2X1_LOC_312/Y AND2X1_LOC_476/Y 0.01fF
C6610 AND2X1_LOC_715/Y OR2X1_LOC_312/Y 0.06fF
C7137 AND2X1_LOC_392/A OR2X1_LOC_312/Y 0.07fF
C8611 OR2X1_LOC_312/Y AND2X1_LOC_661/A 0.03fF
C10978 VDD OR2X1_LOC_312/Y 0.48fF
C16271 OR2X1_LOC_312/Y AND2X1_LOC_169/a_8_24# 0.14fF
C18835 OR2X1_LOC_311/Y OR2X1_LOC_312/Y 0.11fF
C21856 OR2X1_LOC_312/Y AND2X1_LOC_170/B 0.04fF
C22491 AND2X1_LOC_542/a_8_24# OR2X1_LOC_312/Y 0.01fF
C22910 AND2X1_LOC_787/A OR2X1_LOC_312/Y 0.02fF
C22937 AND2X1_LOC_566/B OR2X1_LOC_312/Y 0.03fF
C25897 AND2X1_LOC_716/Y OR2X1_LOC_312/Y 0.07fF
C27932 AND2X1_LOC_552/A OR2X1_LOC_312/Y 0.01fF
C30910 AND2X1_LOC_535/Y OR2X1_LOC_312/Y 0.03fF
C31454 OR2X1_LOC_312/Y AND2X1_LOC_336/a_8_24# 0.01fF
C31708 OR2X1_LOC_312/Y OR2X1_LOC_373/Y 0.56fF
C32218 OR2X1_LOC_109/Y OR2X1_LOC_312/Y 0.41fF
C34611 AND2X1_LOC_543/Y OR2X1_LOC_312/Y 0.63fF
C34810 AND2X1_LOC_365/A OR2X1_LOC_312/Y 0.04fF
C36843 AND2X1_LOC_717/Y OR2X1_LOC_312/Y 0.03fF
C41916 AND2X1_LOC_182/A OR2X1_LOC_312/Y 0.07fF
C42533 OR2X1_LOC_312/Y AND2X1_LOC_337/B 0.01fF
C45759 AND2X1_LOC_539/Y OR2X1_LOC_312/Y 0.07fF
C45766 AND2X1_LOC_552/a_8_24# OR2X1_LOC_312/Y 0.01fF
C47662 AND2X1_LOC_568/B OR2X1_LOC_312/Y 0.07fF
C48579 AND2X1_LOC_703/a_8_24# OR2X1_LOC_312/Y 0.11fF
C51381 AND2X1_LOC_564/B OR2X1_LOC_312/Y 0.01fF
C52415 AND2X1_LOC_784/A OR2X1_LOC_312/Y 0.07fF
C53272 OR2X1_LOC_280/Y OR2X1_LOC_312/Y 0.04fF
C53725 AND2X1_LOC_211/B OR2X1_LOC_312/Y 0.07fF
C55648 AND2X1_LOC_719/Y OR2X1_LOC_312/Y 0.01fF
C57475 OR2X1_LOC_312/Y VSS 0.25fF
C552 OR2X1_LOC_117/Y OR2X1_LOC_67/Y 0.80fF
C7918 AND2X1_LOC_647/B OR2X1_LOC_67/Y 0.06fF
C13061 OR2X1_LOC_67/Y AND2X1_LOC_202/a_8_24# 0.09fF
C30743 AND2X1_LOC_633/Y OR2X1_LOC_67/Y 0.20fF
C32723 AND2X1_LOC_243/Y OR2X1_LOC_67/Y 0.67fF
C42593 AND2X1_LOC_573/A OR2X1_LOC_67/Y 0.07fF
C43593 AND2X1_LOC_647/Y OR2X1_LOC_67/Y 0.80fF
C43976 OR2X1_LOC_607/Y OR2X1_LOC_67/Y 0.03fF
C47551 OR2X1_LOC_609/Y OR2X1_LOC_67/Y 0.12fF
C49119 OR2X1_LOC_69/Y OR2X1_LOC_67/Y 0.01fF
C52430 VDD OR2X1_LOC_67/Y 0.66fF
C53046 AND2X1_LOC_646/a_8_24# OR2X1_LOC_67/Y 0.01fF
C56459 OR2X1_LOC_67/Y VSS 0.31fF
C6347 OR2X1_LOC_613/Y AND2X1_LOC_620/a_8_24# 0.05fF
C9536 OR2X1_LOC_613/Y AND2X1_LOC_620/Y 0.01fF
C19058 OR2X1_LOC_613/Y AND2X1_LOC_658/A 0.01fF
C25812 VDD OR2X1_LOC_613/Y 0.31fF
C25966 OR2X1_LOC_613/Y AND2X1_LOC_624/a_8_24# 0.01fF
C26052 OR2X1_LOC_613/Y AND2X1_LOC_624/B 0.02fF
C30473 AND2X1_LOC_191/B OR2X1_LOC_613/Y 1.38fF
C41900 OR2X1_LOC_528/Y OR2X1_LOC_613/Y 0.87fF
C44670 AND2X1_LOC_191/Y OR2X1_LOC_613/Y 0.01fF
C44679 AND2X1_LOC_711/Y OR2X1_LOC_613/Y 0.03fF
C46649 AND2X1_LOC_191/a_8_24# OR2X1_LOC_613/Y 0.01fF
C52034 OR2X1_LOC_613/Y AND2X1_LOC_632/A 0.04fF
C57402 OR2X1_LOC_613/Y VSS 0.32fF
C13087 AND2X1_LOC_540/a_8_24# OR2X1_LOC_178/Y 0.24fF
C24138 AND2X1_LOC_553/A OR2X1_LOC_178/Y 0.01fF
C24435 OR2X1_LOC_178/Y AND2X1_LOC_465/A 0.02fF
C34571 OR2X1_LOC_178/Y VDD 0.21fF
C39011 OR2X1_LOC_178/Y AND2X1_LOC_523/Y 0.03fF
C52645 OR2X1_LOC_179/Y OR2X1_LOC_178/Y 0.21fF
C55106 OR2X1_LOC_178/Y OR2X1_LOC_108/Y 0.08fF
C57887 OR2X1_LOC_178/Y VSS 0.19fF
C4533 VDD AND2X1_LOC_139/B 0.30fF
C6392 AND2X1_LOC_139/B OR2X1_LOC_416/Y 0.03fF
C6901 AND2X1_LOC_139/A AND2X1_LOC_139/B 0.03fF
C12880 AND2X1_LOC_831/Y AND2X1_LOC_139/B 0.08fF
C25874 AND2X1_LOC_139/B AND2X1_LOC_649/B 0.46fF
C30249 AND2X1_LOC_139/B AND2X1_LOC_476/A 0.07fF
C34609 AND2X1_LOC_139/B AND2X1_LOC_786/Y 0.07fF
C40945 AND2X1_LOC_773/Y AND2X1_LOC_139/B 0.41fF
C42303 OR2X1_LOC_135/Y AND2X1_LOC_139/B 0.01fF
C46344 AND2X1_LOC_76/Y AND2X1_LOC_139/B 0.03fF
C53985 AND2X1_LOC_139/B AND2X1_LOC_139/a_8_24# 0.03fF
C57169 AND2X1_LOC_139/B VSS -0.31fF
C18688 AND2X1_LOC_838/Y AND2X1_LOC_852/B 0.26fF
C34797 AND2X1_LOC_838/Y AND2X1_LOC_852/a_8_24# 0.11fF
C35088 VDD AND2X1_LOC_838/Y 0.20fF
C57241 AND2X1_LOC_838/Y VSS -0.06fF
C4161 AND2X1_LOC_602/a_8_24# AND2X1_LOC_447/Y 0.04fF
C6523 AND2X1_LOC_705/Y AND2X1_LOC_447/Y 0.18fF
C12972 AND2X1_LOC_715/Y AND2X1_LOC_447/Y 0.02fF
C15222 AND2X1_LOC_645/A AND2X1_LOC_447/Y 0.07fF
C17235 VDD AND2X1_LOC_447/Y 0.19fF
C18090 OR2X1_LOC_600/Y AND2X1_LOC_447/Y 0.05fF
C20792 AND2X1_LOC_602/a_36_24# AND2X1_LOC_447/Y 0.01fF
C28309 AND2X1_LOC_605/Y AND2X1_LOC_447/Y 0.02fF
C31978 AND2X1_LOC_724/A AND2X1_LOC_447/Y 0.13fF
C40402 AND2X1_LOC_447/Y OR2X1_LOC_424/Y 0.04fF
C43993 AND2X1_LOC_447/Y AND2X1_LOC_454/a_8_24# 0.11fF
C49350 OR2X1_LOC_601/Y AND2X1_LOC_447/Y 0.05fF
C56788 AND2X1_LOC_447/Y VSS 0.44fF
C28714 AND2X1_LOC_508/A AND2X1_LOC_658/A 0.03fF
C30518 AND2X1_LOC_508/A AND2X1_LOC_474/Y 0.02fF
C32483 AND2X1_LOC_500/Y AND2X1_LOC_508/A 0.05fF
C35436 VDD AND2X1_LOC_508/A 0.21fF
C39709 AND2X1_LOC_508/A AND2X1_LOC_508/B 0.01fF
C39716 AND2X1_LOC_508/A AND2X1_LOC_508/a_8_24# 0.10fF
C43349 AND2X1_LOC_508/A AND2X1_LOC_574/A 0.12fF
C45335 AND2X1_LOC_508/A AND2X1_LOC_510/A 0.27fF
C45347 AND2X1_LOC_574/a_8_24# AND2X1_LOC_508/A 0.20fF
C51774 OR2X1_LOC_528/Y AND2X1_LOC_508/A 0.06fF
C57493 AND2X1_LOC_508/A VSS -0.18fF
C8317 AND2X1_LOC_199/A OR2X1_LOC_13/Y 0.01fF
C11256 VDD AND2X1_LOC_199/A 0.25fF
C44157 AND2X1_LOC_199/A AND2X1_LOC_199/a_8_24# 0.19fF
C57700 AND2X1_LOC_199/A VSS -0.11fF
C7423 AND2X1_LOC_810/A AND2X1_LOC_535/Y 0.01fF
C11659 AND2X1_LOC_715/Y AND2X1_LOC_535/Y 0.13fF
C12195 AND2X1_LOC_535/Y AND2X1_LOC_354/Y 0.03fF
C13536 AND2X1_LOC_535/Y AND2X1_LOC_661/A 0.02fF
C15920 VDD AND2X1_LOC_535/Y 0.01fF
C21313 AND2X1_LOC_535/Y AND2X1_LOC_169/a_8_24# 0.01fF
C21633 AND2X1_LOC_535/Y AND2X1_LOC_354/B 0.27fF
C26773 AND2X1_LOC_535/Y AND2X1_LOC_170/B 0.35fF
C36373 AND2X1_LOC_535/Y AND2X1_LOC_336/a_8_24# 0.01fF
C38037 AND2X1_LOC_535/Y AND2X1_LOC_854/a_8_24# 0.03fF
C39736 AND2X1_LOC_535/Y AND2X1_LOC_365/A 0.02fF
C40478 AND2X1_LOC_388/Y AND2X1_LOC_535/Y 0.03fF
C47069 AND2X1_LOC_535/Y AND2X1_LOC_567/a_8_24# 0.10fF
C47663 AND2X1_LOC_535/Y AND2X1_LOC_337/B 0.02fF
C49341 AND2X1_LOC_535/Y AND2X1_LOC_854/a_36_24# 0.01fF
C50867 AND2X1_LOC_539/Y AND2X1_LOC_535/Y 0.47fF
C53145 AND2X1_LOC_535/Y AND2X1_LOC_336/a_36_24# -0.00fF
C57807 AND2X1_LOC_535/Y VSS 0.34fF
C9397 AND2X1_LOC_557/Y AND2X1_LOC_554/Y 0.20fF
C12259 AND2X1_LOC_557/Y AND2X1_LOC_561/B 0.15fF
C13629 AND2X1_LOC_557/Y AND2X1_LOC_573/A 0.03fF
C16344 AND2X1_LOC_557/Y AND2X1_LOC_561/a_8_24# -0.00fF
C23334 AND2X1_LOC_557/Y VDD 0.21fF
C51008 AND2X1_LOC_557/Y AND2X1_LOC_563/A 0.09fF
C58078 AND2X1_LOC_557/Y VSS 0.11fF
C9344 VDD OR2X1_LOC_793/B -0.00fF
C24702 OR2X1_LOC_793/a_8_216# OR2X1_LOC_793/B 0.01fF
C35650 OR2X1_LOC_805/A OR2X1_LOC_793/B 0.74fF
C56564 OR2X1_LOC_793/B VSS 0.08fF
C7812 VDD OR2X1_LOC_776/A 0.16fF
C10141 OR2X1_LOC_241/Y OR2X1_LOC_776/A 0.01fF
C17197 OR2X1_LOC_737/A OR2X1_LOC_776/A 0.07fF
C23191 OR2X1_LOC_841/a_8_216# OR2X1_LOC_776/A 0.06fF
C34142 OR2X1_LOC_805/A OR2X1_LOC_776/A 0.07fF
C35182 OR2X1_LOC_228/Y OR2X1_LOC_776/A 0.01fF
C41284 OR2X1_LOC_841/A OR2X1_LOC_776/A 0.16fF
C41962 OR2X1_LOC_241/B OR2X1_LOC_776/A 0.09fF
C47085 OR2X1_LOC_841/B OR2X1_LOC_776/A 0.05fF
C55087 OR2X1_LOC_241/a_8_216# OR2X1_LOC_776/A 0.01fF
C56164 OR2X1_LOC_493/Y OR2X1_LOC_776/A 0.15fF
C56322 OR2X1_LOC_776/A VSS 0.23fF
C4222 OR2X1_LOC_196/B OR2X1_LOC_702/a_8_216# 0.02fF
C9817 OR2X1_LOC_196/B OR2X1_LOC_702/a_36_216# 0.02fF
C38111 VDD OR2X1_LOC_196/B 0.26fF
C43007 OR2X1_LOC_702/A OR2X1_LOC_196/B 0.01fF
C57341 OR2X1_LOC_196/B VSS 0.48fF
C13779 OR2X1_LOC_507/A OR2X1_LOC_508/Y 0.02fF
C16026 OR2X1_LOC_507/A OR2X1_LOC_510/Y 0.09fF
C24829 OR2X1_LOC_507/A OR2X1_LOC_510/a_8_216# 0.01fF
C24888 OR2X1_LOC_510/A OR2X1_LOC_507/A 0.30fF
C30639 OR2X1_LOC_507/A OR2X1_LOC_560/A 0.04fF
C36255 VDD OR2X1_LOC_507/A 0.25fF
C42731 OR2X1_LOC_507/a_8_216# OR2X1_LOC_507/A 0.04fF
C42804 OR2X1_LOC_643/A OR2X1_LOC_507/A 0.03fF
C57560 OR2X1_LOC_507/A VSS 0.13fF
C3143 OR2X1_LOC_401/A OR2X1_LOC_401/B 0.08fF
C22139 VDD OR2X1_LOC_401/A 0.21fF
C33991 OR2X1_LOC_401/A OR2X1_LOC_402/Y 0.03fF
C45379 OR2X1_LOC_770/A OR2X1_LOC_401/A 0.16fF
C57276 OR2X1_LOC_401/A VSS 0.18fF
C18064 OR2X1_LOC_345/A OR2X1_LOC_345/a_8_216# 0.47fF
C46348 VDD OR2X1_LOC_345/A -0.00fF
C56835 OR2X1_LOC_345/A VSS 0.15fF
C48706 OR2X1_LOC_602/a_8_216# OR2X1_LOC_602/B 0.05fF
C54875 OR2X1_LOC_602/Y OR2X1_LOC_602/B 0.81fF
C56920 OR2X1_LOC_602/B VSS -0.16fF
C20842 OR2X1_LOC_181/A OR2X1_LOC_181/a_8_216# 0.47fF
C56473 OR2X1_LOC_181/A VSS 0.15fF
C23708 OR2X1_LOC_494/Y AND2X1_LOC_348/A 0.81fF
C36011 AND2X1_LOC_348/A AND2X1_LOC_348/Y 0.04fF
C38994 AND2X1_LOC_348/A AND2X1_LOC_359/B 0.01fF
C40705 AND2X1_LOC_348/A AND2X1_LOC_345/Y 0.01fF
C46398 AND2X1_LOC_348/A AND2X1_LOC_348/a_8_24# 0.10fF
C57665 AND2X1_LOC_348/A VSS 0.24fF
C3365 OR2X1_LOC_231/A OR2X1_LOC_475/B 0.13fF
C10514 VDD OR2X1_LOC_231/A 0.21fF
C17001 OR2X1_LOC_643/A OR2X1_LOC_231/A 0.03fF
C26712 OR2X1_LOC_624/A OR2X1_LOC_231/A 0.06fF
C32333 OR2X1_LOC_231/A OR2X1_LOC_641/B 0.26fF
C34266 OR2X1_LOC_231/A OR2X1_LOC_61/Y 0.03fF
C36815 OR2X1_LOC_231/A OR2X1_LOC_805/A 0.03fF
C41526 OR2X1_LOC_231/A OR2X1_LOC_231/a_8_216# 0.01fF
C49676 OR2X1_LOC_231/B OR2X1_LOC_231/A 0.16fF
C57260 OR2X1_LOC_231/A VSS 0.13fF
C9182 OR2X1_LOC_620/B OR2X1_LOC_550/B 0.04fF
C12241 OR2X1_LOC_620/a_8_216# OR2X1_LOC_620/B 0.05fF
C35735 OR2X1_LOC_620/B OR2X1_LOC_471/Y 0.02fF
C36997 OR2X1_LOC_620/B OR2X1_LOC_620/A 0.11fF
C57490 OR2X1_LOC_620/B VSS -0.01fF
C57349 OR2X1_LOC_636/A VSS -0.13fF
C14756 AND2X1_LOC_712/Y AND2X1_LOC_448/Y 0.01fF
C25782 AND2X1_LOC_713/Y AND2X1_LOC_448/Y 0.01fF
C33933 AND2X1_LOC_448/Y AND2X1_LOC_453/Y 0.18fF
C39434 AND2X1_LOC_448/Y AND2X1_LOC_454/Y 0.37fF
C44167 AND2X1_LOC_448/Y AND2X1_LOC_449/Y 0.13fF
C45459 AND2X1_LOC_448/Y AND2X1_LOC_452/Y 0.02fF
C49841 AND2X1_LOC_448/Y AND2X1_LOC_453/a_8_24# 0.03fF
C56848 AND2X1_LOC_448/Y VSS 0.31fF
C5673 AND2X1_LOC_632/A AND2X1_LOC_620/Y 0.01fF
C11250 AND2X1_LOC_632/A AND2X1_LOC_623/a_8_24# 0.01fF
C22172 VDD AND2X1_LOC_632/A 0.06fF
C22365 AND2X1_LOC_632/A AND2X1_LOC_624/B 0.01fF
C40800 AND2X1_LOC_191/Y AND2X1_LOC_632/A 0.03fF
C40807 AND2X1_LOC_711/Y AND2X1_LOC_632/A 0.03fF
C45237 AND2X1_LOC_632/A OR2X1_LOC_615/Y 0.16fF
C46964 AND2X1_LOC_632/A AND2X1_LOC_631/Y 0.19fF
C57069 AND2X1_LOC_632/A VSS 0.05fF
C4747 OR2X1_LOC_779/Y OR2X1_LOC_784/Y 0.11fF
C22715 OR2X1_LOC_779/Y OR2X1_LOC_725/B 0.72fF
C31328 OR2X1_LOC_779/Y OR2X1_LOC_712/B 0.05fF
C35855 OR2X1_LOC_779/Y OR2X1_LOC_783/a_8_216# 0.02fF
C41184 VDD OR2X1_LOC_779/Y 0.07fF
C41370 OR2X1_LOC_779/Y OR2X1_LOC_783/a_36_216# 0.03fF
C56897 OR2X1_LOC_779/Y VSS 0.18fF
C1109 OR2X1_LOC_851/B OR2X1_LOC_840/A 0.25fF
C10410 OR2X1_LOC_840/A OR2X1_LOC_593/B 0.01fF
C13074 OR2X1_LOC_840/A OR2X1_LOC_468/A 0.03fF
C13203 OR2X1_LOC_840/A OR2X1_LOC_449/B 0.79fF
C20355 OR2X1_LOC_840/A OR2X1_LOC_739/A 0.05fF
C20794 OR2X1_LOC_840/A OR2X1_LOC_539/Y 0.16fF
C25633 OR2X1_LOC_840/A OR2X1_LOC_228/Y 0.10fF
C28181 OR2X1_LOC_840/A OR2X1_LOC_724/A 0.10fF
C29472 OR2X1_LOC_840/A OR2X1_LOC_308/Y 1.77fF
C35524 OR2X1_LOC_851/A OR2X1_LOC_840/A 0.17fF
C37163 OR2X1_LOC_840/A OR2X1_LOC_538/A 0.03fF
C37493 OR2X1_LOC_840/A OR2X1_LOC_356/B 0.10fF
C40518 OR2X1_LOC_833/Y OR2X1_LOC_840/A 0.04fF
C41906 OR2X1_LOC_354/A OR2X1_LOC_840/A 0.05fF
C42594 OR2X1_LOC_840/A OR2X1_LOC_567/a_8_216# 0.31fF
C43935 OR2X1_LOC_840/A OR2X1_LOC_723/B 1.25fF
C46132 OR2X1_LOC_840/A OR2X1_LOC_390/B 0.10fF
C46179 OR2X1_LOC_840/a_8_216# OR2X1_LOC_840/A 0.05fF
C47520 OR2X1_LOC_175/Y OR2X1_LOC_840/A 0.10fF
C47546 OR2X1_LOC_840/A OR2X1_LOC_713/A 0.02fF
C48520 OR2X1_LOC_840/A OR2X1_LOC_620/Y 0.10fF
C54294 VDD OR2X1_LOC_840/A 2.44fF
C57675 OR2X1_LOC_840/A VSS -4.67fF
C3443 OR2X1_LOC_520/Y OR2X1_LOC_642/a_8_216# 0.01fF
C6031 OR2X1_LOC_520/Y AND2X1_LOC_88/Y 0.14fF
C14492 OR2X1_LOC_520/Y OR2X1_LOC_649/B 0.01fF
C25240 OR2X1_LOC_520/Y OR2X1_LOC_559/a_8_216# 0.10fF
C43269 OR2X1_LOC_656/Y OR2X1_LOC_520/Y 0.10fF
C44510 OR2X1_LOC_641/Y OR2X1_LOC_520/Y 0.13fF
C47634 VDD OR2X1_LOC_520/Y 0.03fF
C57654 OR2X1_LOC_520/Y VSS 0.53fF
C55504 OR2X1_LOC_196/Y VDD 0.12fF
C58062 OR2X1_LOC_196/Y VSS 0.14fF
C4385 AND2X1_LOC_631/Y AND2X1_LOC_620/Y 0.01fF
C20813 VDD AND2X1_LOC_631/Y 0.04fF
C36799 OR2X1_LOC_528/Y AND2X1_LOC_631/Y 0.16fF
C39828 AND2X1_LOC_658/B AND2X1_LOC_631/Y 0.01fF
C43922 AND2X1_LOC_631/Y OR2X1_LOC_615/Y 0.01fF
C51204 AND2X1_LOC_631/Y AND2X1_LOC_632/a_8_24# 0.01fF
C56973 AND2X1_LOC_631/Y VSS 0.12fF
C1236 AND2X1_LOC_555/a_8_24# OR2X1_LOC_481/Y 0.04fF
C26856 OR2X1_LOC_481/Y AND2X1_LOC_345/Y 0.82fF
C34887 OR2X1_LOC_481/Y AND2X1_LOC_259/Y 0.03fF
C37251 VDD OR2X1_LOC_481/Y 0.05fF
C51602 OR2X1_LOC_481/Y AND2X1_LOC_345/a_8_24# 0.01fF
C57764 OR2X1_LOC_481/Y VSS 0.14fF
C2251 AND2X1_LOC_339/a_8_24# OR2X1_LOC_416/Y 0.01fF
C4741 AND2X1_LOC_34/a_8_24# OR2X1_LOC_416/Y 0.01fF
C6056 AND2X1_LOC_831/Y OR2X1_LOC_416/Y 0.01fF
C9390 AND2X1_LOC_61/Y OR2X1_LOC_416/Y 0.03fF
C9496 AND2X1_LOC_852/Y OR2X1_LOC_416/Y 0.03fF
C10158 AND2X1_LOC_339/Y OR2X1_LOC_416/Y 0.01fF
C19192 AND2X1_LOC_649/B OR2X1_LOC_416/Y 0.04fF
C23591 AND2X1_LOC_476/A OR2X1_LOC_416/Y 0.03fF
C27961 OR2X1_LOC_416/Y AND2X1_LOC_786/Y 0.15fF
C28521 AND2X1_LOC_34/Y OR2X1_LOC_416/Y 0.01fF
C29454 OR2X1_LOC_416/Y OR2X1_LOC_75/Y 0.23fF
C32335 AND2X1_LOC_633/Y OR2X1_LOC_416/Y 0.02fF
C33725 OR2X1_LOC_595/Y OR2X1_LOC_416/Y 0.02fF
C34263 AND2X1_LOC_773/Y OR2X1_LOC_416/Y 0.03fF
C37642 AND2X1_LOC_340/Y OR2X1_LOC_416/Y 0.03fF
C37846 AND2X1_LOC_634/Y OR2X1_LOC_416/Y 0.58fF
C43454 AND2X1_LOC_640/a_8_24# OR2X1_LOC_416/Y 0.01fF
C44303 OR2X1_LOC_416/Y OR2X1_LOC_27/Y 0.02fF
C49952 OR2X1_LOC_32/Y OR2X1_LOC_416/Y 0.02fF
C54022 VDD OR2X1_LOC_416/Y 0.64fF
C54914 OR2X1_LOC_416/Y AND2X1_LOC_642/Y 0.16fF
C55876 AND2X1_LOC_640/Y OR2X1_LOC_416/Y 0.01fF
C56959 OR2X1_LOC_416/Y VSS -0.01fF
C2579 OR2X1_LOC_651/a_8_216# OR2X1_LOC_651/B 0.06fF
C24671 OR2X1_LOC_654/A OR2X1_LOC_651/B 0.76fF
C24942 VDD OR2X1_LOC_651/B -0.00fF
C57242 OR2X1_LOC_651/B VSS 0.11fF
C17414 OR2X1_LOC_460/Y OR2X1_LOC_463/B 0.07fF
C33956 OR2X1_LOC_463/a_8_216# OR2X1_LOC_463/B 0.03fF
C49754 VDD OR2X1_LOC_463/B 0.12fF
C57118 OR2X1_LOC_463/B VSS -0.00fF
C127 OR2X1_LOC_778/Y OR2X1_LOC_374/Y 0.02fF
C3141 OR2X1_LOC_737/A OR2X1_LOC_374/Y 0.10fF
C5873 OR2X1_LOC_374/Y OR2X1_LOC_593/B 0.03fF
C7969 OR2X1_LOC_374/Y OR2X1_LOC_723/A 0.02fF
C10812 OR2X1_LOC_787/Y OR2X1_LOC_374/Y 0.68fF
C15074 OR2X1_LOC_675/A OR2X1_LOC_374/Y 0.26fF
C20147 OR2X1_LOC_805/A OR2X1_LOC_374/Y 0.10fF
C33666 OR2X1_LOC_794/A OR2X1_LOC_374/Y 0.10fF
C36078 OR2X1_LOC_833/Y OR2X1_LOC_374/Y 0.16fF
C39392 OR2X1_LOC_723/B OR2X1_LOC_374/Y 0.32fF
C41860 OR2X1_LOC_493/Y OR2X1_LOC_374/Y 0.08fF
C44594 OR2X1_LOC_374/Y OR2X1_LOC_605/Y 0.04fF
C49922 VDD OR2X1_LOC_374/Y 0.10fF
C53077 OR2X1_LOC_374/Y OR2X1_LOC_717/a_8_216# 0.02fF
C56326 OR2X1_LOC_374/Y VSS 0.20fF
C22879 OR2X1_LOC_325/Y OR2X1_LOC_538/A 0.01fF
C33822 OR2X1_LOC_325/Y OR2X1_LOC_620/Y 0.02fF
C39679 OR2X1_LOC_325/Y VDD -0.00fF
C48472 OR2X1_LOC_326/B OR2X1_LOC_325/Y 0.06fF
C49686 OR2X1_LOC_325/Y OR2X1_LOC_326/a_8_216# 0.39fF
C50957 OR2X1_LOC_325/Y OR2X1_LOC_703/A 0.03fF
C58038 OR2X1_LOC_325/Y VSS 0.18fF
C4872 OR2X1_LOC_776/Y OR2X1_LOC_785/a_8_216# 0.02fF
C19676 OR2X1_LOC_776/Y OR2X1_LOC_228/Y 0.01fF
C27003 OR2X1_LOC_776/Y OR2X1_LOC_795/B 0.02fF
C29150 OR2X1_LOC_776/Y OR2X1_LOC_785/B 0.16fF
C29339 OR2X1_LOC_786/Y OR2X1_LOC_776/Y 0.03fF
C56781 OR2X1_LOC_776/Y VSS 0.20fF
C12004 OR2X1_LOC_168/Y OR2X1_LOC_170/a_8_216# 0.02fF
C18074 OR2X1_LOC_703/B OR2X1_LOC_168/Y 0.04fF
C18397 OR2X1_LOC_168/Y OR2X1_LOC_390/B 0.71fF
C19693 OR2X1_LOC_175/Y OR2X1_LOC_168/Y 0.01fF
C23113 OR2X1_LOC_168/Y OR2X1_LOC_170/a_36_216# 0.03fF
C24831 OR2X1_LOC_440/B OR2X1_LOC_168/Y 0.01fF
C25916 OR2X1_LOC_168/Y OR2X1_LOC_568/A 0.06fF
C26494 VDD OR2X1_LOC_168/Y 0.24fF
C30298 OR2X1_LOC_440/a_8_216# OR2X1_LOC_168/Y 0.01fF
C32902 OR2X1_LOC_778/Y OR2X1_LOC_168/Y 0.19fF
C35699 OR2X1_LOC_168/Y OR2X1_LOC_180/B 0.03fF
C36093 OR2X1_LOC_168/Y OR2X1_LOC_788/B 0.03fF
C40059 OR2X1_LOC_170/A OR2X1_LOC_168/Y 0.06fF
C41290 OR2X1_LOC_468/A OR2X1_LOC_168/Y 0.03fF
C41383 OR2X1_LOC_449/B OR2X1_LOC_168/Y 0.12fF
C52450 OR2X1_LOC_168/Y OR2X1_LOC_388/a_8_216# 0.02fF
C56472 OR2X1_LOC_168/Y VSS 0.24fF
C6466 OR2X1_LOC_149/B OR2X1_LOC_148/Y 0.14fF
C14238 OR2X1_LOC_149/B VDD 0.12fF
C16934 OR2X1_LOC_149/B OR2X1_LOC_471/Y 0.12fF
C35248 OR2X1_LOC_149/B OR2X1_LOC_546/a_8_216# 0.03fF
C39258 OR2X1_LOC_149/B OR2X1_LOC_213/A 1.83fF
C46473 OR2X1_LOC_149/B OR2X1_LOC_550/B 0.03fF
C57945 OR2X1_LOC_149/B VSS -0.05fF
C1301 OR2X1_LOC_724/A OR2X1_LOC_308/Y 0.21fF
C2289 OR2X1_LOC_711/a_8_216# OR2X1_LOC_308/Y 0.04fF
C4356 OR2X1_LOC_711/B OR2X1_LOC_308/Y 0.04fF
C9994 OR2X1_LOC_147/B OR2X1_LOC_308/Y 0.10fF
C13362 OR2X1_LOC_726/A OR2X1_LOC_308/Y 0.01fF
C13709 OR2X1_LOC_308/Y OR2X1_LOC_727/a_8_216# 0.05fF
C15123 OR2X1_LOC_711/A OR2X1_LOC_308/Y 0.02fF
C20566 OR2X1_LOC_308/Y OR2X1_LOC_713/A 0.02fF
C21506 OR2X1_LOC_620/Y OR2X1_LOC_308/Y 0.03fF
C24747 OR2X1_LOC_703/Y OR2X1_LOC_308/Y 0.03fF
C27344 VDD OR2X1_LOC_308/Y 0.12fF
C33756 OR2X1_LOC_778/Y OR2X1_LOC_308/Y 0.10fF
C35687 OR2X1_LOC_714/a_8_216# OR2X1_LOC_308/Y 0.03fF
C35809 OR2X1_LOC_326/B OR2X1_LOC_308/Y 0.03fF
C38307 OR2X1_LOC_703/A OR2X1_LOC_308/Y 0.12fF
C42236 OR2X1_LOC_449/B OR2X1_LOC_308/Y 2.67fF
C47789 OR2X1_LOC_469/B OR2X1_LOC_308/Y 0.20fF
C49641 OR2X1_LOC_739/A OR2X1_LOC_308/Y 0.03fF
C50796 OR2X1_LOC_566/A OR2X1_LOC_308/Y 0.07fF
C56372 OR2X1_LOC_308/Y VSS 1.05fF
C247 VDD OR2X1_LOC_708/Y -0.00fF
C21192 OR2X1_LOC_708/Y OR2X1_LOC_712/a_8_216# 0.39fF
C41508 OR2X1_LOC_448/Y OR2X1_LOC_708/Y 0.03fF
C46555 OR2X1_LOC_708/Y OR2X1_LOC_712/B 0.06fF
C56572 OR2X1_LOC_708/Y VSS 0.18fF
C4032 OR2X1_LOC_454/a_8_216# OR2X1_LOC_783/A 0.39fF
C8606 OR2X1_LOC_467/A OR2X1_LOC_783/A 0.01fF
C57039 OR2X1_LOC_783/A VSS 0.30fF
C6486 OR2X1_LOC_841/B OR2X1_LOC_228/Y 0.02fF
C12692 OR2X1_LOC_841/B OR2X1_LOC_841/A 0.20fF
C16540 OR2X1_LOC_851/A OR2X1_LOC_841/B 0.86fF
C47527 OR2X1_LOC_841/B OR2X1_LOC_593/B 0.01fF
C50670 OR2X1_LOC_841/a_8_216# OR2X1_LOC_841/B 0.06fF
C57860 OR2X1_LOC_841/B VSS 0.08fF
C953 OR2X1_LOC_841/A OR2X1_LOC_228/Y 0.01fF
C10922 OR2X1_LOC_851/A OR2X1_LOC_841/A 0.01fF
C21479 OR2X1_LOC_841/A OR2X1_LOC_390/B 0.03fF
C29531 VDD OR2X1_LOC_841/A 0.23fF
C41735 OR2X1_LOC_841/A OR2X1_LOC_593/B 0.49fF
C44889 OR2X1_LOC_841/a_8_216# OR2X1_LOC_841/A 0.02fF
C56037 OR2X1_LOC_841/a_36_216# OR2X1_LOC_841/A 0.03fF
C57799 OR2X1_LOC_841/A VSS 0.06fF
C3973 AND2X1_LOC_543/Y AND2X1_LOC_564/B 0.02fF
C5754 AND2X1_LOC_543/Y OR2X1_LOC_280/Y 0.01fF
C14220 AND2X1_LOC_543/Y AND2X1_LOC_476/Y 0.04fF
C19745 AND2X1_LOC_543/Y VDD 0.10fF
C31538 AND2X1_LOC_787/A AND2X1_LOC_543/Y 0.03fF
C36587 AND2X1_LOC_543/Y AND2X1_LOC_552/A 0.09fF
C40411 AND2X1_LOC_543/Y OR2X1_LOC_373/Y 0.14fF
C40907 AND2X1_LOC_543/Y OR2X1_LOC_109/Y 0.04fF
C45700 AND2X1_LOC_543/Y AND2X1_LOC_717/Y 0.01fF
C54583 AND2X1_LOC_543/Y AND2X1_LOC_552/a_8_24# 0.02fF
C57993 AND2X1_LOC_543/Y VSS 0.14fF
C2319 AND2X1_LOC_787/A AND2X1_LOC_476/Y 0.02fF
C7825 AND2X1_LOC_787/A AND2X1_LOC_794/B 0.01fF
C7841 AND2X1_LOC_787/A VDD 0.28fF
C8359 AND2X1_LOC_486/Y AND2X1_LOC_787/A 0.05fF
C19384 AND2X1_LOC_787/a_8_24# AND2X1_LOC_787/A 0.03fF
C19979 AND2X1_LOC_787/A AND2X1_LOC_675/A 0.08fF
C22847 AND2X1_LOC_787/A AND2X1_LOC_716/Y 0.01fF
C25466 AND2X1_LOC_787/A AND2X1_LOC_440/a_8_24# 0.01fF
C26765 AND2X1_LOC_787/A OR2X1_LOC_437/Y 0.06fF
C29109 AND2X1_LOC_787/A OR2X1_LOC_109/Y 0.02fF
C33257 AND2X1_LOC_787/A AND2X1_LOC_180/a_8_24# 0.04fF
C33752 AND2X1_LOC_787/A AND2X1_LOC_717/Y 0.12fF
C35864 AND2X1_LOC_787/a_36_24# AND2X1_LOC_787/A 0.01fF
C38755 AND2X1_LOC_787/A AND2X1_LOC_182/A 0.01fF
C42679 AND2X1_LOC_787/A AND2X1_LOC_471/Y 0.02fF
C45299 AND2X1_LOC_787/A AND2X1_LOC_468/B 0.01fF
C49260 AND2X1_LOC_787/A AND2X1_LOC_784/A 0.19fF
C50561 AND2X1_LOC_787/A AND2X1_LOC_211/B 0.03fF
C52537 AND2X1_LOC_787/A AND2X1_LOC_719/Y 0.10fF
C58018 AND2X1_LOC_787/A VSS 0.08fF
C2934 VDD AND2X1_LOC_303/B 0.02fF
C14765 AND2X1_LOC_566/B AND2X1_LOC_303/B 0.14fF
C17778 AND2X1_LOC_716/Y AND2X1_LOC_303/B 0.52fF
C31352 AND2X1_LOC_303/B AND2X1_LOC_303/a_8_24# 0.01fF
C45528 AND2X1_LOC_211/B AND2X1_LOC_303/B 0.21fF
C54041 AND2X1_LOC_303/A AND2X1_LOC_303/B 0.03fF
C57543 AND2X1_LOC_303/B VSS 0.08fF
C421 AND2X1_LOC_392/A AND2X1_LOC_831/Y 0.07fF
C25587 OR2X1_LOC_109/Y AND2X1_LOC_831/Y 0.02fF
C29906 AND2X1_LOC_831/Y AND2X1_LOC_476/A 0.08fF
C34296 AND2X1_LOC_831/Y AND2X1_LOC_786/Y 0.01fF
C34519 AND2X1_LOC_831/Y AND2X1_LOC_841/a_8_24# 0.03fF
C40660 AND2X1_LOC_773/Y AND2X1_LOC_831/Y 0.21fF
C41983 OR2X1_LOC_135/Y AND2X1_LOC_831/Y 0.10fF
C54861 AND2X1_LOC_831/Y AND2X1_LOC_476/Y 0.09fF
C57238 AND2X1_LOC_831/Y VSS -2.49fF
C2896 AND2X1_LOC_566/B AND2X1_LOC_303/A 0.01fF
C5884 AND2X1_LOC_716/Y AND2X1_LOC_303/A 0.01fF
C16676 AND2X1_LOC_303/A AND2X1_LOC_476/A 0.03fF
C19502 AND2X1_LOC_303/A AND2X1_LOC_303/a_8_24# 0.01fF
C21137 AND2X1_LOC_303/A AND2X1_LOC_786/Y -0.03fF
C28724 AND2X1_LOC_303/A OR2X1_LOC_135/Y 0.09fF
C33572 AND2X1_LOC_303/A AND2X1_LOC_211/B 0.14fF
C47188 VDD AND2X1_LOC_303/A 0.06fF
C47741 AND2X1_LOC_303/A AND2X1_LOC_716/a_8_24# 0.05fF
C57758 AND2X1_LOC_303/A VSS 0.29fF
C9302 OR2X1_LOC_471/a_8_216# OR2X1_LOC_471/B 0.39fF
C30390 VDD OR2X1_LOC_471/B -0.00fF
C48887 OR2X1_LOC_465/Y OR2X1_LOC_471/B 0.12fF
C57439 OR2X1_LOC_471/B VSS 0.17fF
C2713 OR2X1_LOC_65/Y AND2X1_LOC_201/a_8_24# 0.01fF
C4544 AND2X1_LOC_84/Y OR2X1_LOC_65/Y 0.01fF
C14789 OR2X1_LOC_65/Y AND2X1_LOC_201/Y 0.80fF
C24393 AND2X1_LOC_633/Y OR2X1_LOC_65/Y 0.16fF
C39657 OR2X1_LOC_65/Y OR2X1_LOC_72/Y 0.07fF
C45904 VDD OR2X1_LOC_65/Y 0.06fF
C56875 OR2X1_LOC_65/Y VSS 0.10fF
C3710 AND2X1_LOC_786/a_8_24# OR2X1_LOC_262/Y 0.11fF
C12209 AND2X1_LOC_340/Y OR2X1_LOC_262/Y 0.46fF
C18746 OR2X1_LOC_262/Y AND2X1_LOC_573/A 0.02fF
C19927 AND2X1_LOC_340/a_8_24# OR2X1_LOC_262/Y 0.02fF
C22335 OR2X1_LOC_262/Y OR2X1_LOC_72/Y 0.78fF
C28388 VDD OR2X1_LOC_262/Y 0.19fF
C45781 OR2X1_LOC_262/Y OR2X1_LOC_79/Y 0.03fF
C57368 OR2X1_LOC_262/Y VSS 0.22fF
C326 VDD OR2X1_LOC_117/Y 0.04fF
C36751 OR2X1_LOC_117/Y AND2X1_LOC_243/Y 0.02fF
C41237 OR2X1_LOC_117/Y AND2X1_LOC_845/Y 0.08fF
C50763 AND2X1_LOC_554/B OR2X1_LOC_117/Y 0.04fF
C52702 AND2X1_LOC_392/A OR2X1_LOC_117/Y 0.43fF
C57390 OR2X1_LOC_117/Y VSS 0.17fF
C1880 OR2X1_LOC_778/Y OR2X1_LOC_568/A 0.10fF
C2517 VDD OR2X1_LOC_778/Y 2.81fF
C3776 OR2X1_LOC_602/Y OR2X1_LOC_778/Y 0.23fF
C5081 OR2X1_LOC_169/a_8_216# OR2X1_LOC_778/Y 0.35fF
C5354 OR2X1_LOC_851/B OR2X1_LOC_778/Y 0.19fF
C5634 OR2X1_LOC_778/Y OR2X1_LOC_717/a_8_216# 0.01fF
C11727 OR2X1_LOC_778/Y OR2X1_LOC_180/B 0.05fF
C11904 OR2X1_LOC_778/Y OR2X1_LOC_737/A 0.54fF
C12112 OR2X1_LOC_778/Y OR2X1_LOC_788/B 0.03fF
C13595 OR2X1_LOC_703/A OR2X1_LOC_778/Y 0.14fF
C14703 OR2X1_LOC_778/Y OR2X1_LOC_593/B 0.03fF
C16728 OR2X1_LOC_778/Y OR2X1_LOC_723/A 0.03fF
C17161 OR2X1_LOC_778/Y OR2X1_LOC_365/B 0.05fF
C17343 OR2X1_LOC_468/A OR2X1_LOC_778/Y 0.47fF
C21330 OR2X1_LOC_169/B OR2X1_LOC_778/Y 0.05fF
C24120 OR2X1_LOC_778/Y OR2X1_LOC_703/a_8_216# 0.33fF
C24688 OR2X1_LOC_778/Y OR2X1_LOC_739/A 0.05fF
C25554 OR2X1_LOC_778/Y OR2X1_LOC_784/a_8_216# 0.01fF
C28883 OR2X1_LOC_805/A OR2X1_LOC_778/Y 0.11fF
C32387 OR2X1_LOC_778/Y OR2X1_LOC_724/A 0.10fF
C37599 OR2X1_LOC_778/Y OR2X1_LOC_356/A 0.10fF
C41533 OR2X1_LOC_538/A OR2X1_LOC_778/Y 0.03fF
C46351 OR2X1_LOC_354/A OR2X1_LOC_778/Y 0.10fF
C48386 OR2X1_LOC_778/Y OR2X1_LOC_723/B 0.16fF
C50305 OR2X1_LOC_703/B OR2X1_LOC_778/Y 0.22fF
C50858 OR2X1_LOC_778/Y OR2X1_LOC_493/Y 0.45fF
C51799 OR2X1_LOC_175/Y OR2X1_LOC_778/Y 0.10fF
C51835 OR2X1_LOC_778/Y OR2X1_LOC_713/A 0.10fF
C52785 OR2X1_LOC_620/Y OR2X1_LOC_778/Y 0.10fF
C56842 OR2X1_LOC_778/Y VSS 1.13fF
C14941 OR2X1_LOC_335/Y OR2X1_LOC_544/A 0.02fF
C15163 OR2X1_LOC_335/Y OR2X1_LOC_337/a_8_216# 0.07fF
C30823 OR2X1_LOC_335/Y VDD 0.31fF
C45594 OR2X1_LOC_335/Y OR2X1_LOC_365/B 0.03fF
C53436 OR2X1_LOC_337/A OR2X1_LOC_335/Y 0.14fF
C58030 OR2X1_LOC_335/Y VSS 0.05fF
C1450 OR2X1_LOC_208/A OR2X1_LOC_648/B 0.04fF
C23965 OR2X1_LOC_208/A OR2X1_LOC_175/Y 0.04fF
C46144 OR2X1_LOC_208/A OR2X1_LOC_856/B 0.05fF
C58096 OR2X1_LOC_208/A VSS 0.14fF
C39123 AND2X1_LOC_69/Y OR2X1_LOC_202/a_8_216# 0.47fF
C57056 AND2X1_LOC_69/Y VSS 0.13fF
C1024 AND2X1_LOC_554/B AND2X1_LOC_721/A 0.02fF
C3070 AND2X1_LOC_392/A AND2X1_LOC_721/A 0.15fF
C3099 AND2X1_LOC_366/A AND2X1_LOC_721/A 0.08fF
C6833 VDD AND2X1_LOC_721/A 0.60fF
C10322 AND2X1_LOC_720/Y AND2X1_LOC_721/A 0.11fF
C15794 AND2X1_LOC_721/a_8_24# AND2X1_LOC_721/A -0.00fF
C23577 AND2X1_LOC_349/B AND2X1_LOC_721/A 0.10fF
C28692 AND2X1_LOC_721/A OR2X1_LOC_813/Y 0.04fF
C35240 OR2X1_LOC_494/Y AND2X1_LOC_721/A 0.57fF
C39588 AND2X1_LOC_349/a_8_24# AND2X1_LOC_721/A 0.01fF
C50844 AND2X1_LOC_359/B AND2X1_LOC_721/A 0.20fF
C57033 AND2X1_LOC_721/A VSS -2.03fF
C2521 OR2X1_LOC_624/B OR2X1_LOC_768/a_8_216# 0.01fF
C2609 OR2X1_LOC_624/B OR2X1_LOC_400/a_8_216# 0.01fF
C5544 OR2X1_LOC_643/A OR2X1_LOC_624/B 0.03fF
C10328 OR2X1_LOC_624/B OR2X1_LOC_404/Y 0.03fF
C11096 OR2X1_LOC_624/B OR2X1_LOC_402/Y 0.07fF
C13644 OR2X1_LOC_624/B OR2X1_LOC_403/A 0.02fF
C15350 OR2X1_LOC_400/B OR2X1_LOC_624/B 0.05fF
C16681 OR2X1_LOC_624/B OR2X1_LOC_403/a_8_216# 0.01fF
C19565 OR2X1_LOC_624/B OR2X1_LOC_624/a_8_216# 0.01fF
C22206 OR2X1_LOC_624/B OR2X1_LOC_404/a_8_216# 0.05fF
C24609 OR2X1_LOC_624/B OR2X1_LOC_772/A 0.01fF
C27729 OR2X1_LOC_624/B OR2X1_LOC_404/A 0.07fF
C32807 OR2X1_LOC_624/B OR2X1_LOC_84/A 0.01fF
C53639 OR2X1_LOC_624/B OR2X1_LOC_624/Y 0.02fF
C57523 OR2X1_LOC_624/B VSS 0.26fF
C2804 OR2X1_LOC_813/Y AND2X1_LOC_845/Y 0.01fF
C45313 OR2X1_LOC_813/Y AND2X1_LOC_845/a_8_24# 0.05fF
C57032 OR2X1_LOC_813/Y VSS 0.15fF
C5653 AND2X1_LOC_634/Y AND2X1_LOC_476/A 0.03fF
C14628 AND2X1_LOC_633/Y AND2X1_LOC_634/Y 0.19fF
C36037 VDD AND2X1_LOC_634/Y 0.45fF
C37826 AND2X1_LOC_640/Y AND2X1_LOC_634/Y 0.03fF
C47733 AND2X1_LOC_61/Y AND2X1_LOC_634/Y 0.04fF
C47829 AND2X1_LOC_634/Y AND2X1_LOC_852/Y 0.03fF
C57112 AND2X1_LOC_634/Y VSS -0.16fF
C1507 AND2X1_LOC_541/Y VDD 0.19fF
C4884 AND2X1_LOC_541/Y OR2X1_LOC_103/Y 0.19fF
C6545 AND2X1_LOC_541/Y AND2X1_LOC_768/a_8_24# 0.02fF
C17617 AND2X1_LOC_541/Y AND2X1_LOC_772/B 0.01fF
C18050 AND2X1_LOC_541/Y AND2X1_LOC_553/a_8_24# 0.05fF
C27491 AND2X1_LOC_541/Y AND2X1_LOC_560/B 0.24fF
C29069 AND2X1_LOC_541/Y AND2X1_LOC_563/A 0.02fF
C47115 AND2X1_LOC_553/A AND2X1_LOC_541/Y 0.04fF
C50861 AND2X1_LOC_541/Y OR2X1_LOC_106/Y 0.07fF
C53849 AND2X1_LOC_392/A AND2X1_LOC_541/Y 0.03fF
C57957 AND2X1_LOC_541/Y VSS 0.14fF
C143 AND2X1_LOC_633/Y AND2X1_LOC_476/A 0.01fF
C4970 AND2X1_LOC_633/Y AND2X1_LOC_202/Y 0.16fF
C16198 AND2X1_LOC_76/Y AND2X1_LOC_633/Y 0.06fF
C20165 AND2X1_LOC_633/Y AND2X1_LOC_640/a_8_24# 0.11fF
C24465 AND2X1_LOC_633/Y OR2X1_LOC_72/Y 0.02fF
C30539 VDD AND2X1_LOC_633/Y 0.41fF
C35393 AND2X1_LOC_633/Y AND2X1_LOC_203/a_8_24# 0.17fF
C42005 AND2X1_LOC_61/Y AND2X1_LOC_633/Y 0.07fF
C43434 AND2X1_LOC_633/Y AND2X1_LOC_201/a_8_24# 0.17fF
C45396 AND2X1_LOC_84/Y AND2X1_LOC_633/Y 0.02fF
C47510 AND2X1_LOC_633/Y AND2X1_LOC_202/a_8_24# 0.17fF
C55660 AND2X1_LOC_633/Y AND2X1_LOC_201/Y 0.06fF
C57113 AND2X1_LOC_633/Y VSS -0.10fF
C108 AND2X1_LOC_784/A OR2X1_LOC_437/Y 0.31fF
C1454 AND2X1_LOC_784/A AND2X1_LOC_784/a_36_24# 0.01fF
C3406 AND2X1_LOC_784/A AND2X1_LOC_722/A 0.07fF
C3844 AND2X1_LOC_794/A AND2X1_LOC_784/A -0.01fF
C6640 AND2X1_LOC_784/A AND2X1_LOC_180/a_8_24# 0.01fF
C9726 AND2X1_LOC_784/A AND2X1_LOC_357/B 0.02fF
C10549 AND2X1_LOC_784/A AND2X1_LOC_778/Y 0.02fF
C12232 AND2X1_LOC_784/A AND2X1_LOC_182/A 0.04fF
C15155 OR2X1_LOC_176/Y AND2X1_LOC_784/A 0.06fF
C16047 AND2X1_LOC_784/A AND2X1_LOC_784/a_8_24# 0.01fF
C16086 AND2X1_LOC_784/A AND2X1_LOC_471/Y 0.03fF
C17683 AND2X1_LOC_773/Y AND2X1_LOC_784/A 0.10fF
C17741 AND2X1_LOC_784/A AND2X1_LOC_568/B 0.02fF
C18288 AND2X1_LOC_784/A AND2X1_LOC_170/a_8_24# 0.03fF
C18733 AND2X1_LOC_784/A AND2X1_LOC_468/B 0.12fF
C21183 AND2X1_LOC_784/A AND2X1_LOC_181/Y 0.05fF
C23902 AND2X1_LOC_784/A AND2X1_LOC_211/B 1.36fF
C31473 AND2X1_LOC_784/A AND2X1_LOC_326/A 0.02fF
C33427 AND2X1_LOC_392/A AND2X1_LOC_784/A 0.17fF
C36946 AND2X1_LOC_784/A AND2X1_LOC_326/a_8_24# 0.03fF
C37170 AND2X1_LOC_784/A AND2X1_LOC_794/B 0.01fF
C37207 AND2X1_LOC_784/A VDD 0.88fF
C37685 AND2X1_LOC_486/Y AND2X1_LOC_784/A 0.08fF
C40269 AND2X1_LOC_784/A AND2X1_LOC_170/a_36_24# 0.01fF
C42911 AND2X1_LOC_784/A AND2X1_LOC_354/B 0.03fF
C48305 AND2X1_LOC_784/A AND2X1_LOC_170/B 0.02fF
C48604 AND2X1_LOC_784/A AND2X1_LOC_170/Y 0.02fF
C48977 AND2X1_LOC_787/a_8_24# AND2X1_LOC_784/A 0.02fF
C49313 AND2X1_LOC_784/A AND2X1_LOC_566/B 0.03fF
C49550 AND2X1_LOC_784/A AND2X1_LOC_675/A 0.02fF
C50184 AND2X1_LOC_784/A AND2X1_LOC_335/Y 0.02fF
C51544 AND2X1_LOC_784/A AND2X1_LOC_702/Y 0.01fF
C52340 AND2X1_LOC_784/A AND2X1_LOC_716/Y 0.18fF
C58007 AND2X1_LOC_784/A VSS 0.56fF
C4556 VDD OR2X1_LOC_235/Y 0.12fF
C45554 OR2X1_LOC_235/Y AND2X1_LOC_243/a_8_24# 0.23fF
C57057 OR2X1_LOC_235/Y VSS -0.14fF
C3068 OR2X1_LOC_173/Y AND2X1_LOC_175/a_8_24# 0.23fF
C8617 OR2X1_LOC_173/Y AND2X1_LOC_211/B 0.01fF
C22080 VDD OR2X1_LOC_173/Y 0.12fF
C57574 OR2X1_LOC_173/Y VSS 0.06fF
C7240 OR2X1_LOC_292/Y OR2X1_LOC_295/Y 0.04fF
C7625 AND2X1_LOC_259/Y OR2X1_LOC_292/Y 0.14fF
C10068 VDD OR2X1_LOC_292/Y 0.31fF
C53399 AND2X1_LOC_555/Y OR2X1_LOC_292/Y 0.01fF
C57565 OR2X1_LOC_292/Y VSS 0.15fF
C1704 OR2X1_LOC_184/Y AND2X1_LOC_456/a_8_24# 0.10fF
C3455 AND2X1_LOC_719/Y OR2X1_LOC_184/Y 0.31fF
C4615 OR2X1_LOC_184/Y AND2X1_LOC_465/A 0.06fF
C5163 OR2X1_LOC_184/Y AND2X1_LOC_573/A 0.02fF
C6049 AND2X1_LOC_456/Y OR2X1_LOC_184/Y 0.60fF
C8618 AND2X1_LOC_190/a_8_24# OR2X1_LOC_184/Y 0.11fF
C14945 VDD OR2X1_LOC_184/Y 0.36fF
C15376 AND2X1_LOC_486/Y OR2X1_LOC_184/Y 0.25fF
C19645 AND2X1_LOC_191/B OR2X1_LOC_184/Y 0.11fF
C24814 OR2X1_LOC_497/Y OR2X1_LOC_184/Y 0.03fF
C38102 OR2X1_LOC_184/Y AND2X1_LOC_242/B 0.06fF
C57181 OR2X1_LOC_184/Y VSS 0.32fF
C1391 AND2X1_LOC_61/Y OR2X1_LOC_72/Y 0.01fF
C2799 AND2X1_LOC_201/a_8_24# OR2X1_LOC_72/Y 0.06fF
C4673 AND2X1_LOC_84/Y OR2X1_LOC_72/Y 0.03fF
C6624 AND2X1_LOC_202/a_8_24# OR2X1_LOC_72/Y 0.05fF
C14929 OR2X1_LOC_72/Y AND2X1_LOC_201/Y 0.12fF
C20463 OR2X1_LOC_72/Y AND2X1_LOC_202/Y 0.04fF
C42640 OR2X1_LOC_69/Y OR2X1_LOC_72/Y 0.02fF
C46029 VDD OR2X1_LOC_72/Y 0.22fF
C51019 OR2X1_LOC_72/Y AND2X1_LOC_203/a_8_24# 0.09fF
C55144 AND2X1_LOC_201/a_36_24# OR2X1_LOC_72/Y 0.01fF
C56415 OR2X1_LOC_72/Y VSS 0.31fF
C26697 AND2X1_LOC_208/B AND2X1_LOC_34/Y 0.03fF
C28449 AND2X1_LOC_208/B OR2X1_LOC_24/Y 0.05fF
C43266 AND2X1_LOC_208/B AND2X1_LOC_35/Y 0.41fF
C52187 VDD AND2X1_LOC_208/B 0.04fF
C57508 AND2X1_LOC_208/B VSS 0.20fF
C4052 AND2X1_LOC_778/Y AND2X1_LOC_784/a_8_24# 0.11fF
C4948 OR2X1_LOC_496/Y AND2X1_LOC_778/Y 0.01fF
C9562 AND2X1_LOC_564/B AND2X1_LOC_778/Y 0.02fF
C12058 AND2X1_LOC_785/a_8_24# AND2X1_LOC_778/Y 0.01fF
C19787 AND2X1_LOC_476/Y AND2X1_LOC_778/Y 0.07fF
C25306 VDD AND2X1_LOC_778/Y 0.30fF
C29028 AND2X1_LOC_721/Y AND2X1_LOC_778/Y 0.01fF
C37298 AND2X1_LOC_675/A AND2X1_LOC_778/Y 0.07fF
C44076 AND2X1_LOC_775/a_8_24# AND2X1_LOC_778/Y 0.12fF
C46114 OR2X1_LOC_373/Y AND2X1_LOC_778/Y 0.07fF
C50031 AND2X1_LOC_785/Y AND2X1_LOC_778/Y 0.41fF
C55503 AND2X1_LOC_786/Y AND2X1_LOC_778/Y 0.02fF
C56269 AND2X1_LOC_778/Y VSS 0.21fF
C4867 AND2X1_LOC_392/A AND2X1_LOC_335/Y 0.01fF
C20649 AND2X1_LOC_566/B AND2X1_LOC_335/Y 0.02fF
C23704 AND2X1_LOC_716/Y AND2X1_LOC_335/Y 0.04fF
C32445 AND2X1_LOC_335/Y AND2X1_LOC_337/a_8_24# 0.09fF
C57411 AND2X1_LOC_335/Y VSS 0.08fF
C4119 OR2X1_LOC_449/B OR2X1_LOC_713/A 0.07fF
C12131 OR2X1_LOC_678/Y OR2X1_LOC_713/A 0.73fF
C29104 OR2X1_LOC_623/B OR2X1_LOC_713/A 0.15fF
C44103 OR2X1_LOC_705/Y OR2X1_LOC_713/A 0.10fF
C56328 OR2X1_LOC_713/A VSS -0.72fF
C4039 OR2X1_LOC_711/B OR2X1_LOC_711/a_8_216# 0.04fF
C16919 OR2X1_LOC_711/B OR2X1_LOC_711/A 0.48fF
C29066 OR2X1_LOC_711/B VDD 0.06fF
C49562 OR2X1_LOC_711/B OR2X1_LOC_469/B 0.01fF
C58092 OR2X1_LOC_711/B VSS 0.17fF
C1087 AND2X1_LOC_549/Y AND2X1_LOC_565/a_8_24# 0.19fF
C12136 AND2X1_LOC_658/B AND2X1_LOC_549/Y 0.03fF
C45279 AND2X1_LOC_565/B AND2X1_LOC_549/Y 0.09fF
C49202 AND2X1_LOC_549/Y VDD 0.25fF
C57913 AND2X1_LOC_549/Y VSS 0.10fF
C2795 VDD OR2X1_LOC_522/Y 0.04fF
C7143 AND2X1_LOC_523/Y OR2X1_LOC_522/Y 0.79fF
C38564 AND2X1_LOC_851/B OR2X1_LOC_522/Y 0.01fF
C44429 AND2X1_LOC_76/Y OR2X1_LOC_522/Y 0.21fF
C48827 AND2X1_LOC_523/a_8_24# OR2X1_LOC_522/Y 0.01fF
C56445 OR2X1_LOC_522/Y VSS 0.08fF
C42818 OR2X1_LOC_58/Y OR2X1_LOC_32/Y 0.80fF
C47080 VDD OR2X1_LOC_58/Y 0.11fF
C47530 OR2X1_LOC_58/Y OR2X1_LOC_60/Y 0.21fF
C57718 OR2X1_LOC_58/Y VSS 0.13fF
C3052 AND2X1_LOC_34/Y OR2X1_LOC_24/Y 0.04fF
C4923 OR2X1_LOC_24/Y AND2X1_LOC_208/Y 0.80fF
C8603 AND2X1_LOC_35/a_8_24# OR2X1_LOC_24/Y 0.01fF
C24223 AND2X1_LOC_33/a_8_24# OR2X1_LOC_24/Y -0.01fF
C28399 VDD OR2X1_LOC_24/Y 0.07fF
C48973 AND2X1_LOC_208/a_8_24# OR2X1_LOC_24/Y 0.01fF
C53690 AND2X1_LOC_33/Y OR2X1_LOC_24/Y 0.01fF
C56693 OR2X1_LOC_24/Y VSS 0.06fF
C2822 OR2X1_LOC_615/Y AND2X1_LOC_620/Y 1.01fF
C8357 OR2X1_LOC_615/Y AND2X1_LOC_623/a_8_24# 0.03fF
C12393 AND2X1_LOC_658/A OR2X1_LOC_615/Y 0.19fF
C19678 AND2X1_LOC_486/Y OR2X1_LOC_615/Y 0.01fF
C35210 OR2X1_LOC_528/Y OR2X1_LOC_615/Y 0.03fF
C49598 AND2X1_LOC_632/a_8_24# OR2X1_LOC_615/Y 0.02fF
C56866 OR2X1_LOC_615/Y VSS 0.41fF
C4596 OR2X1_LOC_497/Y AND2X1_LOC_842/a_8_24# 0.02fF
C5829 VDD OR2X1_LOC_497/Y 0.39fF
C6284 AND2X1_LOC_486/Y OR2X1_LOC_497/Y 0.10fF
C9669 AND2X1_LOC_721/Y OR2X1_LOC_497/Y 0.04fF
C9712 OR2X1_LOC_482/Y OR2X1_LOC_497/Y 0.01fF
C10192 OR2X1_LOC_497/Y AND2X1_LOC_850/A 0.01fF
C10304 OR2X1_LOC_497/Y AND2X1_LOC_523/Y 0.19fF
C10580 AND2X1_LOC_191/B OR2X1_LOC_497/Y 0.07fF
C15775 OR2X1_LOC_497/Y AND2X1_LOC_844/a_8_24# 0.04fF
C20707 OR2X1_LOC_497/Y AND2X1_LOC_242/a_8_24# 0.05fF
C26195 OR2X1_LOC_497/Y AND2X1_LOC_244/A 0.01fF
C26844 OR2X1_LOC_497/Y AND2X1_LOC_849/A 0.01fF
C29135 OR2X1_LOC_497/Y AND2X1_LOC_242/B 0.51fF
C30460 OR2X1_LOC_497/Y AND2X1_LOC_500/B 0.01fF
C33591 OR2X1_LOC_497/Y AND2X1_LOC_717/B 0.07fF
C48228 OR2X1_LOC_280/Y OR2X1_LOC_497/Y 0.15fF
C50584 AND2X1_LOC_719/Y OR2X1_LOC_497/Y 0.10fF
C53255 AND2X1_LOC_456/Y OR2X1_LOC_497/Y 0.03fF
C54535 OR2X1_LOC_497/Y AND2X1_LOC_842/B 0.03fF
C57437 OR2X1_LOC_497/Y VSS 0.26fF
C519 OR2X1_LOC_320/Y AND2X1_LOC_863/A 0.10fF
C18673 VDD OR2X1_LOC_320/Y 0.04fF
C32731 AND2X1_LOC_702/Y OR2X1_LOC_320/Y 0.01fF
C55223 AND2X1_LOC_773/Y OR2X1_LOC_320/Y 0.56fF
C57542 OR2X1_LOC_320/Y VSS 0.24fF
C30652 AND2X1_LOC_401/a_8_24# OR2X1_LOC_396/Y 0.05fF
C41082 OR2X1_LOC_395/Y OR2X1_LOC_396/Y 0.11fF
C56436 OR2X1_LOC_396/Y VSS 0.24fF
C7341 OR2X1_LOC_599/Y AND2X1_LOC_644/Y 0.79fF
C19568 AND2X1_LOC_539/Y OR2X1_LOC_599/Y 0.03fF
C40531 OR2X1_LOC_599/Y AND2X1_LOC_644/a_8_24# 0.05fF
C40756 VDD OR2X1_LOC_599/Y 0.04fF
C48756 OR2X1_LOC_311/Y OR2X1_LOC_599/Y 0.03fF
C56916 OR2X1_LOC_599/Y VSS -0.03fF
C17665 VDD OR2X1_LOC_39/Y 0.07fF
C34579 OR2X1_LOC_39/Y AND2X1_LOC_194/Y 0.01fF
C44913 OR2X1_LOC_39/Y AND2X1_LOC_194/a_8_24# 0.01fF
C57767 OR2X1_LOC_39/Y VSS -0.02fF
C4266 AND2X1_LOC_852/Y OR2X1_LOC_69/Y 0.03fF
C7493 AND2X1_LOC_84/Y OR2X1_LOC_69/Y 0.80fF
C48907 VDD OR2X1_LOC_69/Y 0.26fF
C56644 OR2X1_LOC_69/Y VSS 0.07fF
C8398 AND2X1_LOC_719/Y OR2X1_LOC_495/Y 0.01fF
C9319 AND2X1_LOC_840/a_8_24# OR2X1_LOC_495/Y 0.01fF
C9782 OR2X1_LOC_495/Y OR2X1_LOC_237/Y 0.24fF
C14806 AND2X1_LOC_851/A OR2X1_LOC_495/Y 0.01fF
C18346 OR2X1_LOC_495/Y AND2X1_LOC_465/Y 0.02fF
C19867 VDD OR2X1_LOC_495/Y 0.26fF
C20338 AND2X1_LOC_486/Y OR2X1_LOC_495/Y 0.03fF
C23687 OR2X1_LOC_482/Y OR2X1_LOC_495/Y 0.04fF
C31997 OR2X1_LOC_495/Y AND2X1_LOC_241/a_8_24# 0.23fF
C43118 OR2X1_LOC_495/Y AND2X1_LOC_242/B 0.01fF
C49352 OR2X1_LOC_495/Y AND2X1_LOC_833/a_8_24# 0.01fF
C54805 OR2X1_LOC_495/Y AND2X1_LOC_840/A 0.03fF
C55747 OR2X1_LOC_496/Y OR2X1_LOC_495/Y 0.05fF
C55858 AND2X1_LOC_851/B OR2X1_LOC_495/Y 0.35fF
C57091 OR2X1_LOC_495/Y VSS 0.13fF
C2406 OR2X1_LOC_485/Y OR2X1_LOC_484/Y 0.29fF
C13690 OR2X1_LOC_484/Y AND2X1_LOC_810/Y 0.26fF
C16425 AND2X1_LOC_486/Y OR2X1_LOC_484/Y 0.78fF
C24352 OR2X1_LOC_484/Y AND2X1_LOC_486/a_8_24# 0.02fF
C57571 OR2X1_LOC_484/Y VSS 0.24fF
C3639 OR2X1_LOC_179/Y AND2X1_LOC_465/A 0.06fF
C13102 OR2X1_LOC_179/Y AND2X1_LOC_181/a_8_24# 0.23fF
C13907 OR2X1_LOC_179/Y VDD 0.16fF
C34183 OR2X1_LOC_179/Y OR2X1_LOC_108/Y 0.01fF
C57981 OR2X1_LOC_179/Y VSS -0.09fF
C892 VDD OR2X1_LOC_146/Y 0.08fF
C7210 OR2X1_LOC_146/Y AND2X1_LOC_213/B 0.31fF
C50336 AND2X1_LOC_658/A OR2X1_LOC_146/Y 0.03fF
C57222 OR2X1_LOC_146/Y VSS 0.22fF
C797 OR2X1_LOC_311/Y OR2X1_LOC_13/Y 1.09fF
C3837 VDD OR2X1_LOC_311/Y 0.11fF
C16628 AND2X1_LOC_356/a_8_24# OR2X1_LOC_311/Y 0.01fF
C27674 AND2X1_LOC_365/A OR2X1_LOC_311/Y 0.15fF
C33456 OR2X1_LOC_311/Y AND2X1_LOC_774/A 0.03fF
C38478 AND2X1_LOC_539/Y OR2X1_LOC_311/Y 0.01fF
C55651 AND2X1_LOC_715/Y OR2X1_LOC_311/Y 0.01fF
C57555 OR2X1_LOC_311/Y VSS 0.32fF
C5215 AND2X1_LOC_719/Y OR2X1_LOC_373/Y 0.03fF
C9941 AND2X1_LOC_785/A OR2X1_LOC_373/Y 0.01fF
C11235 AND2X1_LOC_476/Y OR2X1_LOC_373/Y 0.05fF
C16765 VDD OR2X1_LOC_373/Y 0.39fF
C17245 AND2X1_LOC_486/Y OR2X1_LOC_373/Y 0.19fF
C28164 OR2X1_LOC_373/Y AND2X1_LOC_439/a_8_24# 0.24fF
C28214 AND2X1_LOC_542/a_8_24# OR2X1_LOC_373/Y 0.01fF
C28839 AND2X1_LOC_675/A OR2X1_LOC_373/Y 0.11fF
C33707 AND2X1_LOC_552/A OR2X1_LOC_373/Y 0.03fF
C35462 AND2X1_LOC_775/a_8_24# OR2X1_LOC_373/Y 0.03fF
C37958 OR2X1_LOC_109/Y OR2X1_LOC_373/Y 0.45fF
C51752 AND2X1_LOC_471/Y OR2X1_LOC_373/Y 0.03fF
C56475 OR2X1_LOC_373/Y VSS 0.19fF
C12054 AND2X1_LOC_476/A OR2X1_LOC_27/Y 0.04fF
C17056 AND2X1_LOC_34/Y OR2X1_LOC_27/Y 0.01fF
C42433 VDD OR2X1_LOC_27/Y 0.12fF
C49523 AND2X1_LOC_34/a_8_24# OR2X1_LOC_27/Y 0.01fF
C56530 OR2X1_LOC_27/Y VSS 0.16fF
C5950 OR2X1_LOC_595/Y AND2X1_LOC_786/Y 0.02fF
C8247 OR2X1_LOC_595/Y AND2X1_LOC_643/a_36_24# 0.01fF
C13675 OR2X1_LOC_135/Y OR2X1_LOC_595/Y 0.02fF
C17279 OR2X1_LOC_595/Y AND2X1_LOC_643/a_8_24# 0.07fF
C17529 AND2X1_LOC_76/Y OR2X1_LOC_595/Y 0.01fF
C31877 VDD OR2X1_LOC_595/Y 0.06fF
C56967 OR2X1_LOC_595/Y VSS 0.06fF
C13667 AND2X1_LOC_717/B OR2X1_LOC_237/Y 0.03fF
C21840 AND2X1_LOC_851/B OR2X1_LOC_237/Y 0.06fF
C28081 OR2X1_LOC_280/Y OR2X1_LOC_237/Y 0.72fF
C41904 VDD OR2X1_LOC_237/Y 0.11fF
C41993 OR2X1_LOC_315/Y OR2X1_LOC_237/Y 0.05fF
C45744 AND2X1_LOC_721/Y OR2X1_LOC_237/Y 0.02fF
C46460 AND2X1_LOC_523/Y OR2X1_LOC_237/Y 0.03fF
C56950 OR2X1_LOC_237/Y VSS 0.34fF
C2652 OR2X1_LOC_81/Y OR2X1_LOC_83/Y 0.01fF
C7585 VDD OR2X1_LOC_83/Y 0.24fF
C10250 OR2X1_LOC_83/Y AND2X1_LOC_403/B 0.81fF
C49865 OR2X1_LOC_83/Y OR2X1_LOC_394/Y 0.01fF
C55342 OR2X1_LOC_83/Y AND2X1_LOC_400/a_8_24# 0.01fF
C57657 OR2X1_LOC_83/Y VSS -0.10fF
C10425 OR2X1_LOC_176/Y AND2X1_LOC_568/B 0.03fF
C10888 OR2X1_LOC_176/Y AND2X1_LOC_170/a_8_24# 0.29fF
C21467 AND2X1_LOC_810/A OR2X1_LOC_176/Y 0.17fF
C23849 OR2X1_LOC_176/Y AND2X1_LOC_810/a_8_24# 0.01fF
C26108 AND2X1_LOC_392/A OR2X1_LOC_176/Y 0.03fF
C27570 OR2X1_LOC_176/Y AND2X1_LOC_810/Y 0.01fF
C29901 OR2X1_LOC_176/Y VDD 0.32fF
C40657 OR2X1_LOC_176/Y AND2X1_LOC_170/B 0.02fF
C40961 OR2X1_LOC_176/Y AND2X1_LOC_170/Y 0.25fF
C41754 OR2X1_LOC_176/Y AND2X1_LOC_566/B 0.51fF
C44844 OR2X1_LOC_176/Y AND2X1_LOC_716/Y 0.05fF
C55483 OR2X1_LOC_176/Y AND2X1_LOC_180/a_8_24# 0.09fF
C58095 OR2X1_LOC_176/Y VSS -0.33fF
C9997 OR2X1_LOC_356/A OR2X1_LOC_356/a_8_216# 0.17fF
C14621 OR2X1_LOC_356/B OR2X1_LOC_356/A 0.78fF
C18945 OR2X1_LOC_354/A OR2X1_LOC_356/A 0.37fF
C22905 OR2X1_LOC_703/B OR2X1_LOC_356/A 0.01fF
C25346 OR2X1_LOC_620/Y OR2X1_LOC_356/A 0.27fF
C28577 OR2X1_LOC_703/Y OR2X1_LOC_356/A 0.15fF
C31194 VDD OR2X1_LOC_356/A 0.48fF
C40788 OR2X1_LOC_788/B OR2X1_LOC_356/A 0.04fF
C42241 OR2X1_LOC_703/A OR2X1_LOC_356/A 0.11fF
C45978 OR2X1_LOC_356/A OR2X1_LOC_365/B 0.05fF
C52950 OR2X1_LOC_703/a_8_216# OR2X1_LOC_356/A 0.02fF
C53498 OR2X1_LOC_739/A OR2X1_LOC_356/A 0.03fF
C56291 OR2X1_LOC_356/A VSS 0.20fF
C806 OR2X1_LOC_448/Y OR2X1_LOC_784/Y 0.18fF
C2082 OR2X1_LOC_448/Y OR2X1_LOC_712/a_8_216# 0.03fF
C8985 OR2X1_LOC_448/Y OR2X1_LOC_453/A 0.06fF
C18680 OR2X1_LOC_448/Y OR2X1_LOC_725/B 0.01fF
C27375 OR2X1_LOC_448/Y OR2X1_LOC_712/B 0.02fF
C33521 OR2X1_LOC_448/Y OR2X1_LOC_453/a_8_216# 0.07fF
C35937 OR2X1_LOC_448/Y OR2X1_LOC_466/A 0.03fF
C37177 VDD OR2X1_LOC_448/Y 0.24fF
C57442 OR2X1_LOC_448/Y VSS 0.53fF
C25602 OR2X1_LOC_644/B OR2X1_LOC_644/a_8_216# 0.07fF
C48345 OR2X1_LOC_644/B OR2X1_LOC_228/Y 0.10fF
C57950 OR2X1_LOC_644/B VSS 0.20fF
C4985 OR2X1_LOC_624/A OR2X1_LOC_475/B 0.03fF
C11385 OR2X1_LOC_475/a_8_216# OR2X1_LOC_475/B 0.03fF
C12688 OR2X1_LOC_61/Y OR2X1_LOC_475/B 0.10fF
C15236 OR2X1_LOC_805/A OR2X1_LOC_475/B 5.79fF
C16280 OR2X1_LOC_475/B OR2X1_LOC_228/Y 0.08fF
C16924 OR2X1_LOC_475/a_36_216# OR2X1_LOC_475/B 0.01fF
C17401 OR2X1_LOC_643/a_8_216# OR2X1_LOC_475/B 0.47fF
C23872 OR2X1_LOC_475/Y OR2X1_LOC_475/B 0.01fF
C36456 OR2X1_LOC_216/a_8_216# OR2X1_LOC_475/B 0.05fF
C42692 OR2X1_LOC_392/B OR2X1_LOC_475/B 0.05fF
C44888 VDD OR2X1_LOC_475/B 0.09fF
C47639 OR2X1_LOC_216/A OR2X1_LOC_475/B 0.01fF
C51484 OR2X1_LOC_643/A OR2X1_LOC_475/B 0.08fF
C56566 OR2X1_LOC_475/B VSS 0.46fF
C31381 OR2X1_LOC_128/A OR2X1_LOC_128/B 0.05fF
C42454 OR2X1_LOC_128/B OR2X1_LOC_128/a_8_216# 0.08fF
C55613 OR2X1_LOC_114/B OR2X1_LOC_128/B 0.39fF
C57787 OR2X1_LOC_128/B VSS 0.11fF
C17644 OR2X1_LOC_768/A VDD -0.00fF
C23798 OR2X1_LOC_768/A OR2X1_LOC_849/A 0.02fF
C28850 OR2X1_LOC_768/A OR2X1_LOC_404/Y 0.03fF
C30574 OR2X1_LOC_768/A OR2X1_LOC_720/B 0.01fF
C56028 OR2X1_LOC_768/A OR2X1_LOC_137/a_8_216# 0.47fF
C57894 OR2X1_LOC_768/A VSS 0.26fF
C6612 OR2X1_LOC_192/B OR2X1_LOC_192/a_8_216# 0.07fF
C12399 OR2X1_LOC_565/A OR2X1_LOC_192/B 0.03fF
C12423 OR2X1_LOC_190/Y OR2X1_LOC_192/B 0.35fF
C23168 OR2X1_LOC_564/A OR2X1_LOC_192/B 0.13fF
C34424 OR2X1_LOC_192/A OR2X1_LOC_192/B 0.06fF
C52020 VDD OR2X1_LOC_192/B 0.21fF
C56474 OR2X1_LOC_192/B VSS 0.22fF
C8022 OR2X1_LOC_137/a_8_216# OR2X1_LOC_137/B 0.02fF
C19074 OR2X1_LOC_137/a_36_216# OR2X1_LOC_137/B 0.02fF
C25791 VDD OR2X1_LOC_137/B 0.03fF
C36903 OR2X1_LOC_137/B OR2X1_LOC_404/Y 0.01fF
C38667 OR2X1_LOC_137/B OR2X1_LOC_720/B 0.09fF
C51116 OR2X1_LOC_137/Y OR2X1_LOC_137/B 0.80fF
C57515 OR2X1_LOC_137/B VSS 0.14fF
C3623 OR2X1_LOC_190/A OR2X1_LOC_563/A 0.07fF
C3693 OR2X1_LOC_842/a_8_216# OR2X1_LOC_190/A 0.05fF
C9721 OR2X1_LOC_190/A OR2X1_LOC_456/Y 0.03fF
C12620 OR2X1_LOC_190/A OR2X1_LOC_147/B 0.03fF
C13018 OR2X1_LOC_190/A OR2X1_LOC_190/a_8_216# 0.03fF
C13019 OR2X1_LOC_114/B OR2X1_LOC_190/A 0.03fF
C18523 OR2X1_LOC_830/a_8_216# OR2X1_LOC_190/A 0.01fF
C29532 OR2X1_LOC_842/A OR2X1_LOC_190/A 1.19fF
C29942 VDD OR2X1_LOC_190/A 0.10fF
C32665 OR2X1_LOC_190/A OR2X1_LOC_471/Y 0.08fF
C33799 OR2X1_LOC_190/A OR2X1_LOC_190/B 0.03fF
C44073 OR2X1_LOC_190/A OR2X1_LOC_456/a_8_216# 0.03fF
C49742 OR2X1_LOC_190/A OR2X1_LOC_456/a_36_216# 0.01fF
C57703 OR2X1_LOC_190/A VSS -0.35fF
C458 OR2X1_LOC_788/B OR2X1_LOC_605/Y 0.02fF
C3058 OR2X1_LOC_703/Y OR2X1_LOC_788/B 0.81fF
C3975 OR2X1_LOC_440/B OR2X1_LOC_788/B 0.10fF
C5016 OR2X1_LOC_568/A OR2X1_LOC_788/B 0.13fF
C5612 VDD OR2X1_LOC_788/B 0.02fF
C6915 OR2X1_LOC_602/Y OR2X1_LOC_788/B 0.06fF
C8331 OR2X1_LOC_169/a_8_216# OR2X1_LOC_788/B 0.02fF
C11805 OR2X1_LOC_440/A OR2X1_LOC_788/B 0.11fF
C14938 OR2X1_LOC_788/B OR2X1_LOC_180/B 0.03fF
C16717 OR2X1_LOC_703/A OR2X1_LOC_788/B 0.03fF
C19352 OR2X1_LOC_170/A OR2X1_LOC_788/B 0.03fF
C20360 OR2X1_LOC_788/B OR2X1_LOC_365/B 0.16fF
C24443 OR2X1_LOC_169/B OR2X1_LOC_788/B 0.01fF
C34501 OR2X1_LOC_788/a_8_216# OR2X1_LOC_788/B 0.07fF
C44764 OR2X1_LOC_538/A OR2X1_LOC_788/B 0.02fF
C47365 OR2X1_LOC_170/a_8_216# OR2X1_LOC_788/B 0.06fF
C49600 OR2X1_LOC_354/A OR2X1_LOC_788/B 0.01fF
C53407 OR2X1_LOC_703/B OR2X1_LOC_788/B 0.85fF
C54959 OR2X1_LOC_175/Y OR2X1_LOC_788/B 0.14fF
C55939 OR2X1_LOC_620/Y OR2X1_LOC_788/B 0.03fF
C56346 OR2X1_LOC_788/B VSS 0.40fF
C4140 OR2X1_LOC_653/B OR2X1_LOC_653/a_8_216# 0.05fF
C33335 OR2X1_LOC_653/B OR2X1_LOC_653/Y 0.03fF
C38433 OR2X1_LOC_653/B OR2X1_LOC_653/A 0.11fF
C40827 OR2X1_LOC_653/B OR2X1_LOC_390/B 0.05fF
C58075 OR2X1_LOC_653/B VSS 0.29fF
C480 OR2X1_LOC_605/B OR2X1_LOC_787/Y 0.01fF
C11159 OR2X1_LOC_76/A OR2X1_LOC_605/B 1.93fF
C21404 OR2X1_LOC_605/A OR2X1_LOC_605/B 0.61fF
C32293 OR2X1_LOC_605/B OR2X1_LOC_605/a_8_216# 0.05fF
C45636 OR2X1_LOC_605/B OR2X1_LOC_440/A 0.03fF
C57230 OR2X1_LOC_605/B VSS -0.17fF
C21475 OR2X1_LOC_812/B OR2X1_LOC_558/A 0.03fF
C23758 OR2X1_LOC_493/Y OR2X1_LOC_558/A 0.08fF
C56308 OR2X1_LOC_558/A VSS 0.12fF
C6919 OR2X1_LOC_193/A AND2X1_LOC_7/Y 0.14fF
C23059 OR2X1_LOC_193/A OR2X1_LOC_194/B 0.13fF
C23649 OR2X1_LOC_193/A OR2X1_LOC_193/a_8_216# 0.18fF
C30511 VDD OR2X1_LOC_193/A 0.71fF
C35266 OR2X1_LOC_702/A OR2X1_LOC_193/A 0.15fF
C36096 OR2X1_LOC_193/A OR2X1_LOC_194/Y 0.37fF
C41654 OR2X1_LOC_193/A OR2X1_LOC_193/Y 0.06fF
C45952 OR2X1_LOC_856/B OR2X1_LOC_193/A 0.02fF
C56094 OR2X1_LOC_207/B OR2X1_LOC_193/A 0.02fF
C57291 OR2X1_LOC_193/A VSS 0.51fF
C2910 OR2X1_LOC_678/Y OR2X1_LOC_623/B 0.03fF
C18960 VDD OR2X1_LOC_678/Y 0.14fF
C49957 OR2X1_LOC_678/Y AND2X1_LOC_679/a_8_24# 0.10fF
C57460 OR2X1_LOC_678/Y VSS -0.13fF
C16023 OR2X1_LOC_140/A OR2X1_LOC_510/Y 0.03fF
C17448 OR2X1_LOC_140/A OR2X1_LOC_786/Y 0.01fF
C23332 OR2X1_LOC_140/A OR2X1_LOC_203/Y 0.02fF
C30637 OR2X1_LOC_140/A OR2X1_LOC_560/A 0.14fF
C57578 OR2X1_LOC_140/A VSS 0.29fF
C5295 OR2X1_LOC_770/B OR2X1_LOC_402/Y 0.03fF
C16710 OR2X1_LOC_770/B OR2X1_LOC_770/A 0.22fF
C37175 OR2X1_LOC_770/B OR2X1_LOC_401/Y 0.86fF
C58048 OR2X1_LOC_770/B VSS 0.18fF
C907 OR2X1_LOC_231/B OR2X1_LOC_641/B 0.01fF
C10057 OR2X1_LOC_231/B OR2X1_LOC_231/a_8_216# 0.47fF
C41433 OR2X1_LOC_231/B OR2X1_LOC_643/A 0.05fF
C58139 OR2X1_LOC_231/B VSS 0.10fF
C42956 OR2X1_LOC_646/A OR2X1_LOC_647/A 0.01fF
C50792 OR2X1_LOC_647/Y OR2X1_LOC_646/A 0.95fF
C53756 OR2X1_LOC_646/A OR2X1_LOC_647/a_8_216# 0.01fF
C57395 OR2X1_LOC_646/A VSS 0.08fF
C429 OR2X1_LOC_440/B OR2X1_LOC_440/A 0.16fF
C3577 OR2X1_LOC_440/B OR2X1_LOC_180/B 0.01fF
C54246 OR2X1_LOC_440/B OR2X1_LOC_440/a_8_216# 0.47fF
C57567 OR2X1_LOC_440/B VSS 0.16fF
C3309 OR2X1_LOC_346/a_8_216# OR2X1_LOC_346/A 0.05fF
C25219 OR2X1_LOC_347/A OR2X1_LOC_346/A 0.01fF
C32551 OR2X1_LOC_346/B OR2X1_LOC_346/A 0.05fF
C51731 OR2X1_LOC_114/B OR2X1_LOC_346/A 0.03fF
C56769 OR2X1_LOC_346/A VSS 0.20fF
C2449 OR2X1_LOC_114/B OR2X1_LOC_575/A 0.02fF
C2711 OR2X1_LOC_114/B OR2X1_LOC_735/B 0.03fF
C4929 OR2X1_LOC_114/B OR2X1_LOC_128/a_8_216# 0.01fF
C5340 OR2X1_LOC_114/B OR2X1_LOC_805/A 0.03fF
C9203 OR2X1_LOC_114/B OR2X1_LOC_632/Y 0.01fF
C17676 OR2X1_LOC_114/B OR2X1_LOC_147/B 0.14fF
C23644 OR2X1_LOC_114/B OR2X1_LOC_830/a_8_216# 0.05fF
C25349 OR2X1_LOC_114/B OR2X1_LOC_850/B 0.81fF
C26901 OR2X1_LOC_114/B OR2X1_LOC_844/B 0.92fF
C27264 OR2X1_LOC_114/B OR2X1_LOC_493/Y 0.03fF
C31568 OR2X1_LOC_114/B OR2X1_LOC_140/B 0.01fF
C31881 OR2X1_LOC_114/B OR2X1_LOC_675/Y 0.02fF
C32343 OR2X1_LOC_114/B OR2X1_LOC_500/a_8_216# 0.01fF
C34559 OR2X1_LOC_114/B OR2X1_LOC_842/A 0.02fF
C47847 OR2X1_LOC_114/B OR2X1_LOC_501/a_8_216# 0.01fF
C50144 OR2X1_LOC_114/B OR2X1_LOC_128/A 0.03fF
C54616 OR2X1_LOC_114/B OR2X1_LOC_501/A 0.01fF
C55244 OR2X1_LOC_114/B OR2X1_LOC_346/B 0.03fF
C57908 OR2X1_LOC_114/B VSS 0.53fF
C6733 OR2X1_LOC_833/B OR2X1_LOC_805/A 0.03fF
C10039 OR2X1_LOC_833/B OR2X1_LOC_563/A 0.01fF
C22877 OR2X1_LOC_833/Y OR2X1_LOC_833/B 0.02fF
C23421 OR2X1_LOC_833/B OR2X1_LOC_203/Y 0.45fF
C33229 OR2X1_LOC_833/B OR2X1_LOC_675/Y 0.02fF
C41052 OR2X1_LOC_833/a_8_216# OR2X1_LOC_833/B 0.08fF
C43276 OR2X1_LOC_833/B AND2X1_LOC_72/Y 0.03fF
C43598 OR2X1_LOC_833/B OR2X1_LOC_719/B 0.02fF
C54436 OR2X1_LOC_833/B OR2X1_LOC_203/a_8_216# 0.01fF
C57051 OR2X1_LOC_833/B VSS 0.07fF
C507 OR2X1_LOC_493/A OR2X1_LOC_786/Y 0.01fF
C11356 OR2X1_LOC_493/a_8_216# OR2X1_LOC_493/A 0.01fF
C19440 VDD OR2X1_LOC_493/A 0.02fF
C22079 OR2X1_LOC_216/A OR2X1_LOC_493/A 0.13fF
C28806 OR2X1_LOC_493/A OR2X1_LOC_737/A 0.23fF
C45881 OR2X1_LOC_493/A OR2X1_LOC_805/A 0.15fF
C57104 OR2X1_LOC_493/A VSS 0.22fF
C779 OR2X1_LOC_702/A VDD 0.23fF
C16156 OR2X1_LOC_702/A OR2X1_LOC_856/B 0.03fF
C17032 OR2X1_LOC_702/A OR2X1_LOC_624/A 0.05fF
C27246 OR2X1_LOC_702/A OR2X1_LOC_805/A 0.08fF
C39841 OR2X1_LOC_702/A OR2X1_LOC_538/A 0.02fF
C50143 OR2X1_LOC_175/Y OR2X1_LOC_702/A 0.10fF
C57850 OR2X1_LOC_702/A VSS 0.56fF
C1887 OR2X1_LOC_76/A OR2X1_LOC_241/B 0.23fF
C5584 OR2X1_LOC_76/A OR2X1_LOC_605/A 0.19fF
C16671 OR2X1_LOC_76/A OR2X1_LOC_605/a_8_216# 0.01fF
C18583 OR2X1_LOC_76/A OR2X1_LOC_605/Y 0.01fF
C20088 OR2X1_LOC_76/A OR2X1_LOC_76/Y 0.01fF
C20635 OR2X1_LOC_76/A OR2X1_LOC_675/Y 0.81fF
C23834 VDD OR2X1_LOC_76/A 0.02fF
C26435 OR2X1_LOC_675/a_8_216# OR2X1_LOC_76/A 0.03fF
C29876 OR2X1_LOC_76/A OR2X1_LOC_440/A 4.41fF
C33121 OR2X1_LOC_76/A OR2X1_LOC_737/A 0.07fF
C40780 OR2X1_LOC_76/A OR2X1_LOC_787/Y 0.01fF
C57533 OR2X1_LOC_76/A VSS -0.02fF
C12572 OR2X1_LOC_653/Y OR2X1_LOC_61/A 0.02fF
C20669 OR2X1_LOC_61/A OR2X1_LOC_61/B 0.07fF
C33013 OR2X1_LOC_61/A OR2X1_LOC_476/B 0.04fF
C40913 OR2X1_LOC_61/A OR2X1_LOC_61/a_8_216# 0.47fF
C57775 OR2X1_LOC_61/A VSS 0.15fF
C9936 OR2X1_LOC_84/B OR2X1_LOC_244/A 0.01fF
C15419 OR2X1_LOC_84/B OR2X1_LOC_84/A 0.04fF
C19176 OR2X1_LOC_84/B OR2X1_LOC_204/Y 0.01fF
C26396 OR2X1_LOC_84/B OR2X1_LOC_204/a_8_216# 0.03fF
C31938 OR2X1_LOC_84/B OR2X1_LOC_84/a_8_216# 0.05fF
C53957 OR2X1_LOC_84/B OR2X1_LOC_786/A 1.10fF
C54186 OR2X1_LOC_84/B OR2X1_LOC_84/Y 0.03fF
C57841 OR2X1_LOC_84/B VSS 0.03fF
C307 OR2X1_LOC_770/A OR2X1_LOC_401/B 0.05fF
C33059 VDD OR2X1_LOC_401/B 0.21fF
C45114 OR2X1_LOC_401/B OR2X1_LOC_402/Y 0.03fF
C57275 OR2X1_LOC_401/B VSS 0.14fF
C27959 OR2X1_LOC_710/B OR2X1_LOC_710/a_8_216# 0.05fF
C50237 OR2X1_LOC_710/B OR2X1_LOC_705/Y 0.39fF
C51329 OR2X1_LOC_710/B VDD 0.21fF
C58002 OR2X1_LOC_710/B VSS 0.14fF
C2997 OR2X1_LOC_791/B OR2X1_LOC_555/B 0.06fF
C7106 OR2X1_LOC_791/B VDD 0.09fF
C14947 OR2X1_LOC_791/B OR2X1_LOC_792/a_8_216# 0.03fF
C32478 OR2X1_LOC_345/Y OR2X1_LOC_791/B 0.01fF
C34958 OR2X1_LOC_791/B OR2X1_LOC_345/a_8_216# 0.03fF
C37434 OR2X1_LOC_791/B OR2X1_LOC_792/A 0.44fF
C40431 OR2X1_LOC_791/B OR2X1_LOC_345/a_36_216# 0.01fF
C42771 OR2X1_LOC_348/Y OR2X1_LOC_791/B 0.01fF
C43602 OR2X1_LOC_348/a_8_216# OR2X1_LOC_791/B 0.01fF
C53585 OR2X1_LOC_791/B OR2X1_LOC_850/B 0.16fF
C58015 OR2X1_LOC_791/B VSS 0.32fF
C5656 OR2X1_LOC_784/Y OR2X1_LOC_712/B 0.05fF
C6955 OR2X1_LOC_712/a_8_216# OR2X1_LOC_712/B 0.02fF
C18011 OR2X1_LOC_712/a_36_216# OR2X1_LOC_712/B 0.03fF
C36769 OR2X1_LOC_783/a_8_216# OR2X1_LOC_712/B 0.01fF
C42150 VDD OR2X1_LOC_712/B 0.33fF
C56282 OR2X1_LOC_712/B VSS 0.28fF
C12203 AND2X1_LOC_792/Y AND2X1_LOC_793/B 0.02fF
C15273 AND2X1_LOC_793/B AND2X1_LOC_793/a_8_24# 0.01fF
C23304 AND2X1_LOC_793/Y AND2X1_LOC_793/B 0.01fF
C51198 VDD AND2X1_LOC_793/B 0.06fF
C51656 AND2X1_LOC_486/Y AND2X1_LOC_793/B 0.17fF
C56493 AND2X1_LOC_793/B VSS 0.22fF
C3624 OR2X1_LOC_131/Y AND2X1_LOC_656/a_8_24# 0.24fF
C11997 OR2X1_LOC_131/Y AND2X1_LOC_141/B 0.28fF
C20468 OR2X1_LOC_131/Y AND2X1_LOC_572/A 0.13fF
C26463 OR2X1_LOC_131/Y AND2X1_LOC_656/Y 0.16fF
C26607 OR2X1_LOC_131/Y AND2X1_LOC_772/Y 0.07fF
C42048 OR2X1_LOC_131/Y AND2X1_LOC_573/A 0.11fF
C43074 OR2X1_LOC_131/Y AND2X1_LOC_647/Y 0.02fF
C46017 AND2X1_LOC_554/B OR2X1_LOC_131/Y 0.17fF
C51896 VDD OR2X1_LOC_131/Y 0.25fF
C57705 OR2X1_LOC_131/Y VSS -0.31fF
C12553 VDD OR2X1_LOC_765/Y -0.00fF
C36219 OR2X1_LOC_765/Y AND2X1_LOC_770/a_8_24# 0.10fF
C40558 AND2X1_LOC_452/Y OR2X1_LOC_765/Y 0.78fF
C56670 OR2X1_LOC_765/Y VSS 0.15fF
C4418 OR2X1_LOC_13/Y AND2X1_LOC_193/Y 0.01fF
C9999 OR2X1_LOC_13/Y AND2X1_LOC_194/Y 0.01fF
C16824 AND2X1_LOC_654/B OR2X1_LOC_13/Y 0.02fF
C18590 AND2X1_LOC_193/a_8_24# OR2X1_LOC_13/Y 0.01fF
C25894 AND2X1_LOC_199/a_8_24# OR2X1_LOC_13/Y 0.01fF
C42213 AND2X1_LOC_207/A OR2X1_LOC_13/Y 0.01fF
C49192 VDD OR2X1_LOC_13/Y 0.20fF
C56696 OR2X1_LOC_13/Y VSS -0.27fF
C5866 VDD OR2X1_LOC_229/Y 0.12fF
C45968 AND2X1_LOC_228/Y OR2X1_LOC_229/Y 0.01fF
C51827 OR2X1_LOC_229/Y AND2X1_LOC_231/a_8_24# 0.23fF
C56661 OR2X1_LOC_229/Y VSS -0.13fF
C17533 AND2X1_LOC_728/a_8_24# OR2X1_LOC_679/A 0.09fF
C17836 VDD OR2X1_LOC_679/A 0.21fF
C22178 OR2X1_LOC_679/A OR2X1_LOC_679/Y 0.07fF
C36864 AND2X1_LOC_658/B OR2X1_LOC_679/A 0.03fF
C44107 AND2X1_LOC_544/Y OR2X1_LOC_679/A 0.03fF
C48215 OR2X1_LOC_524/Y OR2X1_LOC_679/A 0.03fF
C53749 AND2X1_LOC_728/Y OR2X1_LOC_679/A 0.01fF
C7830 OR2X1_LOC_603/Y AND2X1_LOC_605/a_8_24# 0.23fF
C18973 AND2X1_LOC_452/Y OR2X1_LOC_603/Y 0.02fF
C47039 VDD OR2X1_LOC_603/Y 0.12fF
C56637 OR2X1_LOC_603/Y VSS 0.06fF
C4862 OR2X1_LOC_494/Y AND2X1_LOC_243/Y 0.07fF
C7901 OR2X1_LOC_494/Y AND2X1_LOC_558/a_8_24# 0.09fF
C9310 OR2X1_LOC_494/Y AND2X1_LOC_348/Y 0.01fF
C9416 OR2X1_LOC_494/Y AND2X1_LOC_845/Y 0.12fF
C11306 OR2X1_LOC_494/Y AND2X1_LOC_474/A 0.05fF
C12258 OR2X1_LOC_494/Y AND2X1_LOC_359/B 0.01fF
C14773 OR2X1_LOC_494/Y AND2X1_LOC_573/A 0.02fF
C15133 AND2X1_LOC_362/a_8_24# OR2X1_LOC_494/Y 0.11fF
C20685 AND2X1_LOC_366/A OR2X1_LOC_494/Y 0.03fF
C24471 VDD OR2X1_LOC_494/Y 0.25fF
C26171 AND2X1_LOC_362/a_36_24# OR2X1_LOC_494/Y 0.01fF
C27877 AND2X1_LOC_720/Y OR2X1_LOC_494/Y 0.01fF
C32588 OR2X1_LOC_494/Y AND2X1_LOC_806/A 0.10fF
C33361 AND2X1_LOC_721/a_8_24# OR2X1_LOC_494/Y 0.04fF
C44055 AND2X1_LOC_720/a_8_24# OR2X1_LOC_494/Y 0.01fF
C57687 OR2X1_LOC_494/Y VSS 0.02fF
C24000 VDD OR2X1_LOC_395/Y 0.08fF
C56476 OR2X1_LOC_395/Y VSS 0.24fF
C36680 VDD OR2X1_LOC_755/Y 0.12fF
C41410 AND2X1_LOC_191/B OR2X1_LOC_755/Y 0.01fF
C44593 OR2X1_LOC_755/Y OR2X1_LOC_757/Y 0.05fF
C45655 OR2X1_LOC_755/Y AND2X1_LOC_791/a_8_24# 0.23fF
C55752 AND2X1_LOC_711/Y OR2X1_LOC_755/Y 0.01fF
C56612 OR2X1_LOC_755/Y VSS 0.06fF
C49294 OR2X1_LOC_700/Y VDD 0.04fF
C51907 OR2X1_LOC_700/Y OR2X1_LOC_701/Y 0.94fF
C58051 OR2X1_LOC_700/Y VSS 0.26fF
C1700 OR2X1_LOC_75/Y AND2X1_LOC_786/Y 0.01fF
C11483 AND2X1_LOC_340/Y OR2X1_LOC_75/Y 0.01fF
C13318 AND2X1_LOC_76/Y OR2X1_LOC_75/Y 0.04fF
C27637 VDD OR2X1_LOC_75/Y 0.21fF
C39840 AND2X1_LOC_339/Y OR2X1_LOC_75/Y 0.81fF
C52882 OR2X1_LOC_74/Y OR2X1_LOC_75/Y 0.08fF
C53412 AND2X1_LOC_476/A OR2X1_LOC_75/Y 0.03fF
C56911 OR2X1_LOC_75/Y VSS 0.19fF
C2831 OR2X1_LOC_609/Y AND2X1_LOC_647/B 0.78fF
C38385 AND2X1_LOC_647/Y OR2X1_LOC_609/Y 0.03fF
C47352 VDD OR2X1_LOC_609/Y 0.04fF
C47963 OR2X1_LOC_609/Y AND2X1_LOC_646/a_8_24# 0.01fF
C56811 OR2X1_LOC_609/Y VSS 0.08fF
C14956 VDD OR2X1_LOC_437/Y 0.12fF
C15386 AND2X1_LOC_486/Y OR2X1_LOC_437/Y 0.23fF
C26969 OR2X1_LOC_437/Y AND2X1_LOC_675/A 0.19fF
C49905 OR2X1_LOC_437/Y AND2X1_LOC_784/a_8_24# 0.23fF
C57106 OR2X1_LOC_437/Y VSS 0.26fF
C2385 OR2X1_LOC_60/Y AND2X1_LOC_61/a_8_24# 0.23fF
C52595 VDD OR2X1_LOC_60/Y 0.16fF
C57717 OR2X1_LOC_60/Y VSS 0.07fF
C47206 VDD OR2X1_LOC_81/Y 0.12fF
C57658 OR2X1_LOC_81/Y VSS 0.08fF
C14450 AND2X1_LOC_346/a_8_24# OR2X1_LOC_295/Y 0.01fF
C25475 AND2X1_LOC_347/B OR2X1_LOC_295/Y 0.79fF
C49409 VDD OR2X1_LOC_295/Y 0.04fF
C57373 OR2X1_LOC_295/Y VSS 0.08fF
C176 AND2X1_LOC_181/Y OR2X1_LOC_108/Y 0.81fF
C2530 OR2X1_LOC_108/Y OR2X1_LOC_280/Y 0.07fF
C4852 AND2X1_LOC_719/Y OR2X1_LOC_108/Y 0.10fF
C6066 OR2X1_LOC_108/Y AND2X1_LOC_465/A 0.15fF
C10027 AND2X1_LOC_190/a_8_24# OR2X1_LOC_108/Y 0.01fF
C15531 AND2X1_LOC_181/a_8_24# OR2X1_LOC_108/Y 0.01fF
C16339 VDD OR2X1_LOC_108/Y 0.06fF
C16466 OR2X1_LOC_108/Y OR2X1_LOC_491/Y 0.02fF
C16847 AND2X1_LOC_486/Y OR2X1_LOC_108/Y 0.07fF
C18658 AND2X1_LOC_465/a_8_24# OR2X1_LOC_108/Y 0.04fF
C20191 AND2X1_LOC_721/Y OR2X1_LOC_108/Y 0.02fF
C20221 OR2X1_LOC_482/Y OR2X1_LOC_108/Y 0.11fF
C20822 OR2X1_LOC_108/Y AND2X1_LOC_523/Y 0.07fF
C25701 OR2X1_LOC_492/Y OR2X1_LOC_108/Y 0.13fF
C33009 OR2X1_LOC_108/Y AND2X1_LOC_493/a_8_24# 0.05fF
C44109 OR2X1_LOC_108/Y AND2X1_LOC_717/B 0.07fF
C50949 AND2X1_LOC_540/a_8_24# OR2X1_LOC_108/Y 0.01fF
C54005 OR2X1_LOC_108/Y AND2X1_LOC_830/a_8_24# 0.03fF
C57659 OR2X1_LOC_108/Y VSS 0.43fF
C235 AND2X1_LOC_486/Y OR2X1_LOC_482/Y 0.07fF
C317 OR2X1_LOC_482/Y OR2X1_LOC_666/Y 0.02fF
C5830 OR2X1_LOC_482/Y AND2X1_LOC_719/a_8_24# 0.23fF
C7056 OR2X1_LOC_482/Y AND2X1_LOC_850/Y 0.07fF
C7999 OR2X1_LOC_482/Y AND2X1_LOC_806/A 0.03fF
C9152 OR2X1_LOC_492/Y OR2X1_LOC_482/Y 0.19fF
C14652 OR2X1_LOC_482/Y AND2X1_LOC_242/a_8_24# 0.04fF
C16460 OR2X1_LOC_482/Y AND2X1_LOC_493/a_8_24# 0.12fF
C18914 OR2X1_LOC_482/Y AND2X1_LOC_499/a_8_24# 0.04fF
C23166 OR2X1_LOC_482/Y AND2X1_LOC_242/B 0.07fF
C24083 AND2X1_LOC_509/Y OR2X1_LOC_482/Y 0.03fF
C25673 OR2X1_LOC_482/Y AND2X1_LOC_242/a_36_24# 0.01fF
C27505 OR2X1_LOC_482/Y AND2X1_LOC_717/B 0.05fF
C29130 OR2X1_LOC_482/Y AND2X1_LOC_833/a_8_24# 0.10fF
C33003 OR2X1_LOC_482/Y AND2X1_LOC_493/a_36_24# 0.06fF
C34604 OR2X1_LOC_482/Y AND2X1_LOC_840/A 0.17fF
C37235 OR2X1_LOC_482/Y AND2X1_LOC_830/a_8_24# 0.06fF
C40090 OR2X1_LOC_482/Y AND2X1_LOC_833/a_36_24# 0.07fF
C44383 AND2X1_LOC_719/Y OR2X1_LOC_482/Y 0.03fF
C46220 OR2X1_LOC_482/Y AND2X1_LOC_573/A 0.03fF
C48548 OR2X1_LOC_482/Y AND2X1_LOC_842/B 0.03fF
C49199 OR2X1_LOC_482/Y AND2X1_LOC_658/A 0.33fF
C51812 OR2X1_LOC_482/Y AND2X1_LOC_474/a_8_24# 0.06fF
C55216 OR2X1_LOC_482/Y AND2X1_LOC_859/Y 0.01fF
C55968 VDD OR2X1_LOC_482/Y 0.60fF
C56074 OR2X1_LOC_482/Y OR2X1_LOC_491/Y 0.15fF
C57696 OR2X1_LOC_482/Y VSS 0.60fF
C5241 VDD OR2X1_LOC_492/Y 0.17fF
C5720 AND2X1_LOC_486/Y OR2X1_LOC_492/Y 0.03fF
C22056 OR2X1_LOC_492/Y AND2X1_LOC_493/a_8_24# 0.01fF
C32993 OR2X1_LOC_492/Y AND2X1_LOC_717/B 0.01fF
C42836 OR2X1_LOC_492/Y AND2X1_LOC_830/a_8_24# 0.23fF
C57763 OR2X1_LOC_492/Y VSS 0.10fF
C6133 OR2X1_LOC_135/Y AND2X1_LOC_303/a_8_24# 0.15fF
C6163 AND2X1_LOC_702/a_8_24# OR2X1_LOC_135/Y 0.01fF
C14228 AND2X1_LOC_773/Y OR2X1_LOC_135/Y 0.03fF
C19180 OR2X1_LOC_135/Y AND2X1_LOC_643/a_8_24# 0.03fF
C20307 OR2X1_LOC_135/Y AND2X1_LOC_211/B 0.10fF
C33727 VDD OR2X1_LOC_135/Y 1.34fF
C45666 AND2X1_LOC_566/B OR2X1_LOC_135/Y 0.01fF
C48039 AND2X1_LOC_702/Y OR2X1_LOC_135/Y 0.79fF
C48804 AND2X1_LOC_716/Y OR2X1_LOC_135/Y 0.10fF
C51354 OR2X1_LOC_45/Y OR2X1_LOC_135/Y 0.10fF
C55127 OR2X1_LOC_135/Y AND2X1_LOC_649/B 0.19fF
C57726 OR2X1_LOC_135/Y VSS 0.34fF
C5139 OR2X1_LOC_521/Y AND2X1_LOC_851/B 0.01fF
C10981 OR2X1_LOC_521/Y AND2X1_LOC_76/Y 0.01fF
C18506 OR2X1_LOC_106/Y OR2X1_LOC_521/Y 0.18fF
C57817 OR2X1_LOC_521/Y VSS 0.09fF
C13415 VDD OR2X1_LOC_79/Y 0.06fF
C28187 AND2X1_LOC_84/Y OR2X1_LOC_79/Y 0.42fF
C43468 OR2X1_LOC_79/Y AND2X1_LOC_786/Y 0.79fF
C44761 AND2X1_LOC_786/a_8_24# OR2X1_LOC_79/Y 0.01fF
C53368 AND2X1_LOC_340/Y OR2X1_LOC_79/Y 0.14fF
C56684 OR2X1_LOC_79/Y VSS 0.11fF
C26987 OR2X1_LOC_20/Y AND2X1_LOC_33/a_8_24# 0.23fF
C31215 VDD OR2X1_LOC_20/Y 0.12fF
C57404 OR2X1_LOC_20/Y VSS 0.06fF
C2220 VDD OR2X1_LOC_257/Y 0.12fF
C19411 OR2X1_LOC_257/Y AND2X1_LOC_259/a_8_24# 0.23fF
C55925 AND2X1_LOC_259/Y OR2X1_LOC_257/Y 0.01fF
C56363 OR2X1_LOC_257/Y VSS 0.06fF
C35024 OR2X1_LOC_607/Y AND2X1_LOC_647/Y 0.02fF
C43781 VDD OR2X1_LOC_607/Y 0.12fF
C44396 OR2X1_LOC_607/Y AND2X1_LOC_646/a_8_24# 0.23fF
C57131 OR2X1_LOC_607/Y VSS 0.06fF
C273 OR2X1_LOC_496/Y AND2X1_LOC_785/Y 0.27fF
C5771 OR2X1_LOC_496/Y AND2X1_LOC_786/Y 0.04fF
C15972 AND2X1_LOC_564/B OR2X1_LOC_496/Y 0.02fF
C25007 OR2X1_LOC_496/Y AND2X1_LOC_658/A 0.03fF
C31746 OR2X1_LOC_496/Y VDD 0.14fF
C35457 OR2X1_LOC_496/Y AND2X1_LOC_721/Y 0.03fF
C41970 OR2X1_LOC_496/Y AND2X1_LOC_734/Y 0.01fF
C43881 OR2X1_LOC_496/Y AND2X1_LOC_675/A 0.02fF
C51011 OR2X1_LOC_496/Y AND2X1_LOC_499/a_8_24# 0.11fF
C57964 OR2X1_LOC_496/Y VSS 0.19fF
C45854 OR2X1_LOC_666/Y AND2X1_LOC_658/A 0.40fF
C51989 OR2X1_LOC_666/Y AND2X1_LOC_859/Y 0.02fF
C52727 VDD OR2X1_LOC_666/Y 0.05fF
C57563 OR2X1_LOC_666/Y VSS 0.18fF
C5248 OR2X1_LOC_528/Y OR2X1_LOC_505/Y 0.04fF
C8047 AND2X1_LOC_711/Y OR2X1_LOC_505/Y 0.08fF
C8358 AND2X1_LOC_658/B OR2X1_LOC_505/Y 0.13fF
C16356 AND2X1_LOC_675/Y OR2X1_LOC_505/Y 0.02fF
C43980 OR2X1_LOC_505/Y AND2X1_LOC_507/a_8_24# 0.01fF
C45280 VDD OR2X1_LOC_505/Y 0.19fF
C49654 OR2X1_LOC_505/Y AND2X1_LOC_508/B 0.01fF
C53562 OR2X1_LOC_505/Y AND2X1_LOC_806/A 0.25fF
C57428 OR2X1_LOC_505/Y VSS 0.12fF
C35847 OR2X1_LOC_485/Y OR2X1_LOC_526/Y 0.42fF
C42709 OR2X1_LOC_526/Y AND2X1_LOC_658/A 0.03fF
C46499 OR2X1_LOC_526/Y AND2X1_LOC_796/A 0.28fF
C49658 VDD OR2X1_LOC_526/Y 0.31fF
C52596 OR2X1_LOC_526/Y AND2X1_LOC_705/a_8_24# 0.08fF
C57761 OR2X1_LOC_526/Y VSS -0.09fF
C6966 AND2X1_LOC_636/a_8_24# OR2X1_LOC_583/Y 0.23fF
C12127 VDD OR2X1_LOC_583/Y 0.12fF
C56711 OR2X1_LOC_583/Y VSS 0.06fF
C48094 VDD OR2X1_LOC_32/Y 0.11fF
C54941 OR2X1_LOC_32/Y AND2X1_LOC_34/a_8_24# 0.11fF
C57351 OR2X1_LOC_32/Y VSS 0.12fF
C1223 OR2X1_LOC_74/Y AND2X1_LOC_76/a_8_24# 0.23fF
C6695 OR2X1_LOC_74/Y AND2X1_LOC_76/Y 0.01fF
C21145 VDD OR2X1_LOC_74/Y 0.12fF
C57467 OR2X1_LOC_74/Y VSS 0.06fF
C3991 AND2X1_LOC_231/Y OR2X1_LOC_230/Y 0.79fF
C20255 AND2X1_LOC_228/Y OR2X1_LOC_230/Y 0.01fF
C26045 OR2X1_LOC_230/Y AND2X1_LOC_231/a_8_24# 0.01fF
C36212 VDD OR2X1_LOC_230/Y 0.04fF
C56660 OR2X1_LOC_230/Y VSS 0.08fF
C39804 OR2X1_LOC_600/Y AND2X1_LOC_602/a_8_24# 0.23fF
C42215 AND2X1_LOC_705/Y OR2X1_LOC_600/Y 0.03fF
C53032 VDD OR2X1_LOC_600/Y 0.12fF
C57528 OR2X1_LOC_600/Y VSS -0.33fF
C1136 AND2X1_LOC_181/Y OR2X1_LOC_109/Y 0.04fF
C3448 OR2X1_LOC_280/Y OR2X1_LOC_109/Y 0.02fF
C5753 AND2X1_LOC_719/Y OR2X1_LOC_109/Y 0.10fF
C11777 OR2X1_LOC_109/Y AND2X1_LOC_476/Y 0.19fF
C17300 VDD OR2X1_LOC_109/Y 0.62fF
C17388 OR2X1_LOC_109/Y OR2X1_LOC_315/Y 0.01fF
C17761 AND2X1_LOC_486/Y OR2X1_LOC_109/Y 0.03fF
C28715 AND2X1_LOC_542/a_8_24# OR2X1_LOC_109/Y 0.01fF
C34196 AND2X1_LOC_552/A OR2X1_LOC_109/Y 0.01fF
C43256 AND2X1_LOC_717/Y OR2X1_LOC_109/Y 0.07fF
C47823 OR2X1_LOC_109/Y AND2X1_LOC_841/a_8_24# 0.01fF
C52158 AND2X1_LOC_552/a_8_24# OR2X1_LOC_109/Y 0.02fF
C52265 OR2X1_LOC_109/Y AND2X1_LOC_471/Y 0.03fF
C53301 OR2X1_LOC_109/Y AND2X1_LOC_851/B 0.01fF
C57611 OR2X1_LOC_109/Y VSS 0.27fF
C12829 OR2X1_LOC_491/Y AND2X1_LOC_493/a_8_24# 0.23fF
C23910 OR2X1_LOC_491/Y AND2X1_LOC_717/B 0.01fF
C52277 VDD OR2X1_LOC_491/Y 0.12fF
C57050 OR2X1_LOC_491/Y VSS 0.06fF
C457 OR2X1_LOC_315/Y AND2X1_LOC_523/Y 0.02fF
C21979 OR2X1_LOC_315/Y AND2X1_LOC_445/a_8_24# 0.11fF
C26176 OR2X1_LOC_315/Y AND2X1_LOC_786/Y 0.07fF
C31909 OR2X1_LOC_315/Y AND2X1_LOC_851/B 0.04fF
C35900 AND2X1_LOC_181/Y OR2X1_LOC_315/Y 1.82fF
C46674 OR2X1_LOC_315/Y AND2X1_LOC_476/Y 0.09fF
C52237 VDD OR2X1_LOC_315/Y 0.20fF
C57253 OR2X1_LOC_315/Y VSS 0.38fF
C5363 VDD OR2X1_LOC_517/Y 0.12fF
C25922 OR2X1_LOC_517/Y AND2X1_LOC_559/a_8_24# 0.23fF
C47278 OR2X1_LOC_517/Y AND2X1_LOC_76/Y 0.01fF
C57625 OR2X1_LOC_517/Y VSS 0.06fF
C530 VDD OR2X1_LOC_399/Y 0.12fF
C3189 AND2X1_LOC_403/B OR2X1_LOC_399/Y 0.13fF
C22739 AND2X1_LOC_403/a_8_24# OR2X1_LOC_399/Y 0.23fF
C47014 AND2X1_LOC_573/A OR2X1_LOC_399/Y 0.01fF
C56295 OR2X1_LOC_399/Y VSS -0.33fF
C8524 AND2X1_LOC_191/B OR2X1_LOC_757/Y 0.38fF
C12574 OR2X1_LOC_757/Y AND2X1_LOC_791/a_8_24# 0.04fF
C22696 AND2X1_LOC_711/Y OR2X1_LOC_757/Y 0.01fF
C56514 OR2X1_LOC_757/Y VSS 0.22fF
C54763 OR2X1_LOC_701/Y VDD 0.08fF
C58050 OR2X1_LOC_701/Y VSS 0.12fF
C13503 OR2X1_LOC_45/Y VDD 0.26fF
C37218 OR2X1_LOC_45/Y AND2X1_LOC_654/B 0.14fF
C57927 OR2X1_LOC_45/Y VSS 0.39fF
C19268 VDD OR2X1_LOC_424/Y 0.09fF
C30295 AND2X1_LOC_605/Y OR2X1_LOC_424/Y 0.07fF
C53685 OR2X1_LOC_424/Y AND2X1_LOC_449/a_8_24# 0.09fF
C56465 OR2X1_LOC_424/Y VSS -0.02fF
C25895 AND2X1_LOC_347/Y OR2X1_LOC_297/Y 0.06fF
C41513 VDD OR2X1_LOC_297/Y 0.12fF
C42094 OR2X1_LOC_297/Y AND2X1_LOC_347/a_8_24# 0.23fF
C48954 AND2X1_LOC_710/Y OR2X1_LOC_297/Y 0.01fF
C57482 OR2X1_LOC_297/Y VSS 0.06fF
C36057 OR2X1_LOC_485/Y AND2X1_LOC_810/Y 0.02fF
C38350 VDD OR2X1_LOC_485/Y 0.31fF
C41357 OR2X1_LOC_485/Y AND2X1_LOC_705/a_8_24# 0.07fF
C46894 OR2X1_LOC_485/Y AND2X1_LOC_486/a_8_24# 0.05fF
C57762 OR2X1_LOC_485/Y VSS 0.47fF
C690 OR2X1_LOC_122/Y AND2X1_LOC_474/A 0.01fF
C6974 OR2X1_LOC_122/Y OR2X1_LOC_106/Y 0.15fF
C50502 OR2X1_LOC_122/Y AND2X1_LOC_243/Y 0.03fF
C54919 OR2X1_LOC_122/Y AND2X1_LOC_845/Y 0.03fF
C58064 OR2X1_LOC_122/Y VSS 0.20fF
C1062 OR2X1_LOC_528/Y AND2X1_LOC_475/Y 0.05fF
C2461 OR2X1_LOC_528/Y AND2X1_LOC_573/A 0.03fF
C5265 OR2X1_LOC_528/Y AND2X1_LOC_658/A 0.03fF
C7126 OR2X1_LOC_528/Y AND2X1_LOC_474/Y 0.14fF
C8345 OR2X1_LOC_528/Y AND2X1_LOC_565/B 0.02fF
C9180 OR2X1_LOC_528/Y AND2X1_LOC_500/Y 0.03fF
C11379 OR2X1_LOC_528/Y AND2X1_LOC_859/Y 0.14fF
C12116 OR2X1_LOC_528/Y VDD 0.90fF
C12294 OR2X1_LOC_528/Y AND2X1_LOC_624/a_8_24# 0.01fF
C12391 OR2X1_LOC_528/Y AND2X1_LOC_624/B 0.05fF
C15875 OR2X1_LOC_528/Y AND2X1_LOC_721/Y 0.06fF
C16334 OR2X1_LOC_528/Y AND2X1_LOC_508/B 0.02fF
C18207 OR2X1_LOC_528/Y AND2X1_LOC_475/a_8_24# 0.01fF
C19995 OR2X1_LOC_528/Y AND2X1_LOC_574/A 0.09fF
C20320 OR2X1_LOC_528/Y AND2X1_LOC_806/A 0.02fF
C21490 OR2X1_LOC_528/Y AND2X1_LOC_734/a_8_24# 0.01fF
C22404 OR2X1_LOC_528/Y AND2X1_LOC_734/Y 0.01fF
C29344 OR2X1_LOC_528/Y AND2X1_LOC_792/Y 0.07fF
C30925 OR2X1_LOC_528/Y AND2X1_LOC_191/Y 0.03fF
C30937 OR2X1_LOC_528/Y AND2X1_LOC_711/Y 0.03fF
C31209 OR2X1_LOC_528/Y AND2X1_LOC_658/B 0.57fF
C39243 OR2X1_LOC_528/Y AND2X1_LOC_675/Y 0.06fF
C40305 OR2X1_LOC_528/Y AND2X1_LOC_793/Y 0.19fF
C48896 OR2X1_LOC_528/Y AND2X1_LOC_620/a_8_24# 0.01fF
C51975 OR2X1_LOC_528/Y AND2X1_LOC_620/Y 0.04fF
C52531 OR2X1_LOC_528/Y AND2X1_LOC_564/B 0.19fF
C58081 OR2X1_LOC_528/Y VSS -0.77fF
C3300 OR2X1_LOC_152/Y AND2X1_LOC_209/Y 0.01fF
C3798 VDD OR2X1_LOC_152/Y 0.39fF
C8051 OR2X1_LOC_152/Y OR2X1_LOC_679/Y 0.01fF
C22689 AND2X1_LOC_191/Y OR2X1_LOC_152/Y 0.03fF
C25434 AND2X1_LOC_209/a_8_24# OR2X1_LOC_152/Y 0.01fF
C40973 AND2X1_LOC_727/Y OR2X1_LOC_152/Y 0.01fF
C53100 OR2X1_LOC_152/Y AND2X1_LOC_726/a_8_24# 0.25fF
C53156 OR2X1_LOC_152/Y OR2X1_LOC_679/a_8_216# 0.03fF
C57821 OR2X1_LOC_152/Y VSS -0.33fF
C5447 OR2X1_LOC_524/Y AND2X1_LOC_148/Y 0.03fF
C5757 OR2X1_LOC_524/Y AND2X1_LOC_545/a_8_24# 0.07fF
C5835 AND2X1_LOC_728/Y OR2X1_LOC_524/Y 0.06fF
C7426 AND2X1_LOC_727/Y OR2X1_LOC_524/Y 0.03fF
C15116 OR2X1_LOC_524/Y AND2X1_LOC_475/Y 0.01fF
C16823 AND2X1_LOC_550/a_8_24# OR2X1_LOC_524/Y 0.03fF
C16876 OR2X1_LOC_524/Y AND2X1_LOC_545/a_36_24# 0.01fF
C20671 OR2X1_LOC_524/Y AND2X1_LOC_476/Y 0.15fF
C22411 AND2X1_LOC_565/B OR2X1_LOC_524/Y 0.01fF
C25890 OR2X1_LOC_524/Y AND2X1_LOC_728/a_8_24# 0.13fF
C26168 VDD OR2X1_LOC_524/Y 2.11fF
C32425 OR2X1_LOC_524/Y AND2X1_LOC_213/B 0.03fF
C45032 AND2X1_LOC_191/Y OR2X1_LOC_524/Y 0.07fF
C45042 AND2X1_LOC_711/Y OR2X1_LOC_524/Y 0.07fF
C45315 AND2X1_LOC_658/B OR2X1_LOC_524/Y 0.39fF
C52562 AND2X1_LOC_544/Y OR2X1_LOC_524/Y 0.43fF
C52696 OR2X1_LOC_524/Y AND2X1_LOC_550/A 0.02fF
C57805 OR2X1_LOC_524/Y VSS 0.66fF
C17141 AND2X1_LOC_192/Y OR2X1_LOC_747/Y 0.02fF
C19831 OR2X1_LOC_747/Y AND2X1_LOC_781/Y 0.09fF
C25341 OR2X1_LOC_747/Y AND2X1_LOC_782/a_8_24# 0.23fF
C33147 VDD OR2X1_LOC_747/Y 0.12fF
C56354 OR2X1_LOC_747/Y VSS 0.06fF
C29669 OR2X1_LOC_394/Y AND2X1_LOC_400/a_8_24# 0.01fF
C37997 VDD OR2X1_LOC_394/Y 0.05fF
C40655 OR2X1_LOC_394/Y AND2X1_LOC_403/B 0.01fF
C56745 OR2X1_LOC_394/Y VSS 0.22fF
C14942 OR2X1_LOC_601/Y AND2X1_LOC_602/a_8_24# -0.00fF
C23699 AND2X1_LOC_715/Y OR2X1_LOC_601/Y 0.14fF
C25953 OR2X1_LOC_601/Y AND2X1_LOC_645/A 0.01fF
C27947 VDD OR2X1_LOC_601/Y 0.18fF
C42763 AND2X1_LOC_724/A OR2X1_LOC_601/Y 0.12fF
C56807 OR2X1_LOC_601/Y VSS 0.11fF
C7990 OR2X1_LOC_280/Y AND2X1_LOC_445/a_8_24# 0.23fF
C9898 OR2X1_LOC_280/Y AND2X1_LOC_717/B 0.10fF
C10153 AND2X1_LOC_542/a_36_24# OR2X1_LOC_280/Y 0.02fF
C12228 OR2X1_LOC_280/Y AND2X1_LOC_786/Y 0.07fF
C14175 OR2X1_LOC_280/Y AND2X1_LOC_844/a_36_24# 0.01fF
C16869 AND2X1_LOC_552/a_8_24# OR2X1_LOC_280/Y 0.03fF
C17979 OR2X1_LOC_280/Y AND2X1_LOC_851/B 0.16fF
C18649 OR2X1_LOC_280/Y AND2X1_LOC_243/Y 0.02fF
C22459 AND2X1_LOC_564/B OR2X1_LOC_280/Y 1.43fF
C23132 OR2X1_LOC_280/Y AND2X1_LOC_845/Y 0.02fF
C25058 OR2X1_LOC_280/Y AND2X1_LOC_474/A 0.02fF
C26684 AND2X1_LOC_719/Y OR2X1_LOC_280/Y 0.10fF
C27888 OR2X1_LOC_280/Y AND2X1_LOC_465/A 0.07fF
C27892 AND2X1_LOC_552/a_36_24# OR2X1_LOC_280/Y 0.01fF
C28486 OR2X1_LOC_280/Y AND2X1_LOC_573/A 0.02fF
C32585 OR2X1_LOC_280/Y AND2X1_LOC_476/Y 0.21fF
C33961 AND2X1_LOC_717/a_8_24# OR2X1_LOC_280/Y 0.04fF
C38065 VDD OR2X1_LOC_280/Y 0.39fF
C41890 AND2X1_LOC_721/Y OR2X1_LOC_280/Y 1.54fF
C42566 OR2X1_LOC_280/Y AND2X1_LOC_523/Y 0.92fF
C45079 AND2X1_LOC_717/a_36_24# OR2X1_LOC_280/Y 0.01fF
C46456 OR2X1_LOC_280/Y AND2X1_LOC_806/A 0.02fF
C48278 OR2X1_LOC_280/Y AND2X1_LOC_844/a_8_24# 0.03fF
C49771 AND2X1_LOC_542/a_8_24# OR2X1_LOC_280/Y 0.03fF
C55237 AND2X1_LOC_552/A OR2X1_LOC_280/Y 0.02fF
C57631 OR2X1_LOC_280/Y VSS 0.33fF
C8378 OR2X1_LOC_106/Y AND2X1_LOC_124/a_8_24# 0.23fF
C13883 OR2X1_LOC_106/Y AND2X1_LOC_572/A 0.27fF
C15141 OR2X1_LOC_106/Y AND2X1_LOC_560/B 0.07fF
C25663 OR2X1_LOC_106/Y AND2X1_LOC_243/Y 0.05fF
C30078 OR2X1_LOC_106/Y AND2X1_LOC_845/Y -0.01fF
C31225 AND2X1_LOC_554/Y OR2X1_LOC_106/Y 0.02fF
C31967 OR2X1_LOC_106/Y AND2X1_LOC_474/A 0.03fF
C35398 OR2X1_LOC_106/Y AND2X1_LOC_573/A 0.04fF
C39303 OR2X1_LOC_106/Y AND2X1_LOC_554/B 0.14fF
C45222 OR2X1_LOC_106/Y VDD 0.51fF
C48765 OR2X1_LOC_106/Y OR2X1_LOC_103/Y 0.03fF
C55000 OR2X1_LOC_106/Y AND2X1_LOC_554/a_8_24# 0.03fF
C57916 OR2X1_LOC_106/Y VSS 0.20fF
C3870 OR2X1_LOC_103/Y AND2X1_LOC_523/Y 0.16fF
C15963 AND2X1_LOC_553/a_8_24# OR2X1_LOC_103/Y 0.01fF
C25467 AND2X1_LOC_560/B OR2X1_LOC_103/Y 0.23fF
C27039 AND2X1_LOC_563/A OR2X1_LOC_103/Y 0.01fF
C44938 AND2X1_LOC_553/A OR2X1_LOC_103/Y 0.02fF
C55582 VDD OR2X1_LOC_103/Y 0.24fF
C57331 OR2X1_LOC_103/Y VSS 0.26fF
C31170 OR2X1_LOC_544/A OR2X1_LOC_439/a_8_216# 0.47fF
C39729 OR2X1_LOC_544/A OR2X1_LOC_544/B 0.07fF
C53643 OR2X1_LOC_544/A OR2X1_LOC_439/B 0.04fF
C57002 OR2X1_LOC_544/A VSS 0.21fF
C26855 OR2X1_LOC_605/A OR2X1_LOC_605/a_8_216# 0.03fF
C28716 OR2X1_LOC_605/A OR2X1_LOC_605/Y 0.16fF
C39974 OR2X1_LOC_605/A OR2X1_LOC_440/A 0.07fF
C51172 OR2X1_LOC_605/A OR2X1_LOC_787/Y 0.02fF
C57231 OR2X1_LOC_605/A VSS 0.30fF
C2026 OR2X1_LOC_501/B OR2X1_LOC_575/A 0.07fF
C8328 OR2X1_LOC_501/B OR2X1_LOC_563/A 0.46fF
C8811 OR2X1_LOC_501/B OR2X1_LOC_632/Y 0.08fF
C21666 OR2X1_LOC_501/B OR2X1_LOC_203/Y 0.01fF
C31174 OR2X1_LOC_501/B OR2X1_LOC_140/B 0.03fF
C34584 VDD OR2X1_LOC_501/B 0.03fF
C54201 OR2X1_LOC_501/B OR2X1_LOC_501/A 0.11fF
C56795 OR2X1_LOC_501/B VSS -0.22fF
C23571 OR2X1_LOC_675/A OR2X1_LOC_440/A 0.42fF
C26793 OR2X1_LOC_675/A OR2X1_LOC_737/A 0.01fF
C43819 OR2X1_LOC_675/A OR2X1_LOC_805/A 0.03fF
C50777 OR2X1_LOC_675/A OR2X1_LOC_719/Y 0.43fF
C51701 OR2X1_LOC_675/A OR2X1_LOC_241/B 0.03fF
C57072 OR2X1_LOC_675/A VSS 0.32fF
C8515 OR2X1_LOC_124/A OR2X1_LOC_633/B 0.26fF
C15224 VDD OR2X1_LOC_633/B 0.16fF
C28155 OR2X1_LOC_633/B OR2X1_LOC_720/B 0.08fF
C31331 OR2X1_LOC_633/B OR2X1_LOC_786/A 0.01fF
C37205 OR2X1_LOC_633/B OR2X1_LOC_786/a_8_216# 0.01fF
C42099 OR2X1_LOC_123/B OR2X1_LOC_633/B 0.05fF
C48116 OR2X1_LOC_123/a_8_216# OR2X1_LOC_633/B 0.14fF
C52506 OR2X1_LOC_633/B OR2X1_LOC_786/Y 0.93fF
C57079 OR2X1_LOC_633/B VSS -0.12fF
C4011 OR2X1_LOC_123/B OR2X1_LOC_786/Y 0.01fF
C16106 OR2X1_LOC_124/A OR2X1_LOC_123/B 0.81fF
C22992 VDD OR2X1_LOC_123/B -0.00fF
C55719 OR2X1_LOC_123/a_8_216# OR2X1_LOC_123/B 0.06fF
C57126 OR2X1_LOC_123/B VSS 0.12fF
C9415 OR2X1_LOC_835/A OR2X1_LOC_835/B 0.14fF
C33129 OR2X1_LOC_654/A OR2X1_LOC_835/B 0.07fF
C33417 VDD OR2X1_LOC_835/B 0.02fF
C57615 OR2X1_LOC_835/B VSS 0.24fF
C8556 OR2X1_LOC_439/a_8_216# OR2X1_LOC_439/B 0.08fF
C13434 VDD OR2X1_LOC_439/B 0.23fF
C17114 OR2X1_LOC_439/B OR2X1_LOC_544/B 0.49fF
C19580 OR2X1_LOC_440/A OR2X1_LOC_439/B 0.50fF
C22746 OR2X1_LOC_439/B OR2X1_LOC_180/B 0.76fF
C41766 OR2X1_LOC_439/B OR2X1_LOC_180/a_8_216# 0.16fF
C56537 OR2X1_LOC_439/B VSS 0.02fF
C4866 OR2X1_LOC_175/Y OR2X1_LOC_175/B 0.09fF
C10414 OR2X1_LOC_175/B OR2X1_LOC_174/Y 0.04fF
C21495 OR2X1_LOC_175/B OR2X1_LOC_175/a_8_216# 0.06fF
C27136 OR2X1_LOC_856/B OR2X1_LOC_175/B 0.02fF
C27981 OR2X1_LOC_175/B OR2X1_LOC_624/A 0.01fF
C50997 OR2X1_LOC_175/B OR2X1_LOC_538/A 0.03fF
C57702 OR2X1_LOC_175/B VSS 0.23fF
C10080 AND2X1_LOC_72/Y OR2X1_LOC_719/B 1.05fF
C20831 AND2X1_LOC_72/Y OR2X1_LOC_203/a_8_216# 0.05fF
C32449 AND2X1_LOC_72/Y OR2X1_LOC_563/A 0.01fF
C55330 OR2X1_LOC_76/Y AND2X1_LOC_72/Y 0.17fF
C56994 AND2X1_LOC_72/Y VSS 0.14fF
C16768 OR2X1_LOC_174/A OR2X1_LOC_174/a_8_216# 0.01fF
C19125 OR2X1_LOC_333/B OR2X1_LOC_174/A 0.08fF
C24013 OR2X1_LOC_174/A OR2X1_LOC_174/Y 0.20fF
C41491 OR2X1_LOC_624/A OR2X1_LOC_174/A 0.03fF
C49316 OR2X1_LOC_174/A OR2X1_LOC_61/Y 0.01fF
C57266 OR2X1_LOC_174/A VSS 0.38fF
C1510 VDD OR2X1_LOC_641/A 0.14fF
C3646 OR2X1_LOC_124/a_8_216# OR2X1_LOC_641/A 0.06fF
C9181 OR2X1_LOC_124/a_36_216# OR2X1_LOC_641/A 0.01fF
C16005 OR2X1_LOC_641/A OR2X1_LOC_340/Y 1.22fF
C23517 OR2X1_LOC_641/A OR2X1_LOC_641/B 0.25fF
C29708 OR2X1_LOC_244/A OR2X1_LOC_641/A 0.01fF
C38529 OR2X1_LOC_643/Y OR2X1_LOC_641/A 0.03fF
C38611 OR2X1_LOC_786/Y OR2X1_LOC_641/A 0.03fF
C38908 OR2X1_LOC_204/Y OR2X1_LOC_641/A 0.39fF
C46143 OR2X1_LOC_510/A OR2X1_LOC_641/A 0.03fF
C52030 OR2X1_LOC_641/A OR2X1_LOC_560/A 0.03fF
C56603 OR2X1_LOC_641/A VSS 0.28fF
C28503 OR2X1_LOC_84/Y OR2X1_LOC_786/A 0.16fF
C34129 OR2X1_LOC_786/A OR2X1_LOC_786/a_8_216# 0.01fF
C40248 OR2X1_LOC_244/A OR2X1_LOC_786/A 0.02fF
C49460 OR2X1_LOC_786/Y OR2X1_LOC_786/A 0.02fF
C56774 OR2X1_LOC_786/A VSS 0.34fF
C0 VDD OR2X1_LOC_620/A -0.00fF
C2774 OR2X1_LOC_471/Y OR2X1_LOC_620/A 0.12fF
C32089 OR2X1_LOC_620/A OR2X1_LOC_550/B 0.02fF
C35185 OR2X1_LOC_620/a_8_216# OR2X1_LOC_620/A 0.47fF
C56809 OR2X1_LOC_620/A VSS -0.01fF
C1847 OR2X1_LOC_444/B OR2X1_LOC_444/a_8_216# 0.47fF
C46974 OR2X1_LOC_443/Y OR2X1_LOC_444/B 0.16fF
C57311 OR2X1_LOC_444/B VSS 0.16fF
C15991 OR2X1_LOC_545/B OR2X1_LOC_181/Y 0.17fF
C24059 OR2X1_LOC_545/B OR2X1_LOC_545/a_8_216# 0.05fF
C28609 OR2X1_LOC_545/B OR2X1_LOC_443/a_8_216# 0.01fF
C29436 OR2X1_LOC_545/B OR2X1_LOC_443/Y 0.03fF
C34799 VDD OR2X1_LOC_545/B 0.21fF
C37464 OR2X1_LOC_545/B OR2X1_LOC_471/Y 0.16fF
C45971 OR2X1_LOC_703/A OR2X1_LOC_545/B 0.05fF
C51751 OR2X1_LOC_545/B OR2X1_LOC_551/B 0.07fF
C57378 OR2X1_LOC_545/B VSS 0.04fF
C16069 VDD OR2X1_LOC_346/B 0.21fF
C56942 OR2X1_LOC_346/B VSS 0.20fF
C6302 OR2X1_LOC_703/B OR2X1_LOC_169/B 0.24fF
C7917 OR2X1_LOC_175/Y OR2X1_LOC_169/B 0.01fF
C14226 OR2X1_LOC_169/B OR2X1_LOC_568/A 0.06fF
C17411 OR2X1_LOC_169/a_8_216# OR2X1_LOC_169/B 0.47fF
C29421 OR2X1_LOC_169/B OR2X1_LOC_365/B 0.01fF
C57446 OR2X1_LOC_169/B VSS 0.15fF
C25003 VDD OR2X1_LOC_191/B 0.30fF
C41478 OR2X1_LOC_191/B OR2X1_LOC_565/A 0.34fF
C41745 OR2X1_LOC_191/B OR2X1_LOC_551/B 0.04fF
C52731 OR2X1_LOC_191/B OR2X1_LOC_191/a_8_216# 0.10fF
C57514 OR2X1_LOC_191/B VSS 0.25fF
C16387 OR2X1_LOC_190/B OR2X1_LOC_190/Y 0.10fF
C38857 OR2X1_LOC_190/B OR2X1_LOC_190/a_8_216# 0.01fF
C52771 OR2X1_LOC_190/B OR2X1_LOC_553/a_8_216# 0.47fF
C56658 OR2X1_LOC_190/B VSS 0.35fF
C5869 OR2X1_LOC_339/a_8_216# OR2X1_LOC_333/B 0.01fF
C16482 OR2X1_LOC_333/B OR2X1_LOC_648/B 0.03fF
C17187 OR2X1_LOC_333/B OR2X1_LOC_228/Y 0.16fF
C28784 OR2X1_LOC_351/B OR2X1_LOC_333/B 0.03fF
C37149 OR2X1_LOC_333/B OR2X1_LOC_174/a_8_216# 0.03fF
C42759 OR2X1_LOC_333/B OR2X1_LOC_174/a_36_216# 0.03fF
C45851 OR2X1_LOC_333/B VDD 0.11fF
C54195 OR2X1_LOC_333/B OR2X1_LOC_339/Y 0.11fF
C57834 OR2X1_LOC_333/B VSS 0.39fF
C2035 OR2X1_LOC_781/B OR2X1_LOC_781/a_8_216# 0.01fF
C10009 OR2X1_LOC_781/B VDD -0.00fF
C36817 OR2X1_LOC_781/B OR2X1_LOC_781/Y 0.80fF
C57961 OR2X1_LOC_781/B VSS 0.10fF
C15668 OR2X1_LOC_400/B OR2X1_LOC_400/a_8_216# 0.47fF
C57979 OR2X1_LOC_400/B VSS 0.16fF
C10406 AND2X1_LOC_7/Y OR2X1_LOC_228/a_8_216# 0.07fF
C14243 OR2X1_LOC_651/A AND2X1_LOC_7/Y 0.12fF
C21565 AND2X1_LOC_7/Y OR2X1_LOC_193/a_8_216# 0.07fF
C28467 VDD AND2X1_LOC_7/Y 0.21fF
C34037 OR2X1_LOC_194/Y AND2X1_LOC_7/Y 0.03fF
C39555 OR2X1_LOC_193/Y AND2X1_LOC_7/Y 0.03fF
C56854 AND2X1_LOC_7/Y VSS -0.03fF
C3227 VDD OR2X1_LOC_719/B 0.17fF
C15903 OR2X1_LOC_719/B OR2X1_LOC_719/a_8_216# 0.02fF
C21152 OR2X1_LOC_203/a_8_216# OR2X1_LOC_719/B 0.14fF
C21515 OR2X1_LOC_719/B OR2X1_LOC_719/a_36_216# 0.03fF
C32821 OR2X1_LOC_563/A OR2X1_LOC_719/B 0.02fF
C37338 OR2X1_LOC_241/B OR2X1_LOC_719/B 0.03fF
C46247 OR2X1_LOC_203/Y OR2X1_LOC_719/B 0.17fF
C56239 OR2X1_LOC_719/B VSS 0.17fF
C8117 OR2X1_LOC_555/A OR2X1_LOC_555/B 0.04fF
C12287 VDD OR2X1_LOC_555/A 0.21fF
C57103 OR2X1_LOC_555/A VSS 0.12fF
C14189 OR2X1_LOC_194/B OR2X1_LOC_194/a_8_216# 0.06fF
C44475 VDD OR2X1_LOC_194/B -0.00fF
C50252 OR2X1_LOC_194/Y OR2X1_LOC_194/B 0.86fF
C57136 OR2X1_LOC_194/B VSS 0.12fF
C36827 OR2X1_LOC_128/A OR2X1_LOC_128/a_8_216# 0.47fF
C57788 OR2X1_LOC_128/A VSS 0.15fF
C4901 AND2X1_LOC_88/Y OR2X1_LOC_560/A 0.01fF
C6410 OR2X1_LOC_656/Y AND2X1_LOC_88/Y 0.01fF
C44446 AND2X1_LOC_88/Y OR2X1_LOC_559/a_8_216# 0.01fF
C56480 AND2X1_LOC_88/Y VSS 0.32fF
C4081 VDD OR2X1_LOC_402/B 0.04fF
C8539 OR2X1_LOC_402/B OR2X1_LOC_402/a_8_216# 0.02fF
C16043 OR2X1_LOC_402/B OR2X1_LOC_402/Y 0.17fF
C19548 OR2X1_LOC_402/B OR2X1_LOC_402/a_36_216# 0.01fF
C57783 OR2X1_LOC_402/B VSS -0.16fF
C1319 OR2X1_LOC_773/B OR2X1_LOC_774/Y 0.09fF
C24907 OR2X1_LOC_773/B OR2X1_LOC_773/Y 0.16fF
C26394 OR2X1_LOC_773/B OR2X1_LOC_772/Y 0.06fF
C38011 OR2X1_LOC_773/B VDD 0.21fF
C48652 OR2X1_LOC_773/B OR2X1_LOC_773/a_8_216# 0.06fF
C57965 OR2X1_LOC_773/B VSS 0.19fF
C49 OR2X1_LOC_593/B OR2X1_LOC_390/B 0.02fF
C3090 OR2X1_LOC_593/B OR2X1_LOC_605/Y 0.08fF
C8262 VDD OR2X1_LOC_593/B 0.38fF
C19659 OR2X1_LOC_593/B OR2X1_LOC_718/a_8_216# 0.01fF
C23237 OR2X1_LOC_449/B OR2X1_LOC_593/B 0.66fF
C23604 OR2X1_LOC_841/a_8_216# OR2X1_LOC_593/B 0.03fF
C25329 OR2X1_LOC_787/Y OR2X1_LOC_593/B 0.05fF
C37326 OR2X1_LOC_716/a_8_216# OR2X1_LOC_593/B 0.01fF
C45665 OR2X1_LOC_851/A OR2X1_LOC_593/B 0.01fF
C54074 OR2X1_LOC_723/B OR2X1_LOC_593/B 0.01fF
C56297 OR2X1_LOC_593/B VSS 0.42fF
C2630 OR2X1_LOC_703/B OR2X1_LOC_449/B 0.15fF
C2846 OR2X1_LOC_449/B OR2X1_LOC_390/B 0.05fF
C4095 OR2X1_LOC_175/Y OR2X1_LOC_449/B 0.07fF
C5044 OR2X1_LOC_620/Y OR2X1_LOC_449/B 0.07fF
C9750 OR2X1_LOC_466/A OR2X1_LOC_449/B 0.21fF
C10415 OR2X1_LOC_449/B OR2X1_LOC_568/A 0.55fF
C10969 VDD OR2X1_LOC_449/B 0.27fF
C25829 OR2X1_LOC_468/A OR2X1_LOC_449/B 0.03fF
C26251 OR2X1_LOC_452/a_8_216# OR2X1_LOC_449/B 0.04fF
C33081 OR2X1_LOC_449/B OR2X1_LOC_739/A 0.03fF
C40866 OR2X1_LOC_449/B OR2X1_LOC_724/A 0.87fF
C43879 OR2X1_LOC_454/a_8_216# OR2X1_LOC_449/B 0.01fF
C48533 OR2X1_LOC_467/A OR2X1_LOC_449/B 1.26fF
C50229 OR2X1_LOC_538/A OR2X1_LOC_449/B 0.03fF
C50504 OR2X1_LOC_449/B OR2X1_LOC_356/B 0.07fF
C54839 OR2X1_LOC_354/A OR2X1_LOC_449/B 0.46fF
C56830 OR2X1_LOC_449/B VSS 0.54fF
C42251 OR2X1_LOC_343/B OR2X1_LOC_493/Y 0.01fF
C50329 VDD OR2X1_LOC_343/B -0.00fF
C54465 OR2X1_LOC_343/B OR2X1_LOC_343/a_8_216# 0.47fF
C56832 OR2X1_LOC_343/B VSS 0.15fF
C2169 OR2X1_LOC_124/A OR2X1_LOC_720/B 0.09fF
C8969 VDD OR2X1_LOC_720/B 0.09fF
C10767 OR2X1_LOC_720/B OR2X1_LOC_720/a_8_216# 0.02fF
C15229 OR2X1_LOC_720/B OR2X1_LOC_721/a_8_216# 0.01fF
C15382 OR2X1_LOC_643/A OR2X1_LOC_720/B 0.03fF
C16251 OR2X1_LOC_720/B OR2X1_LOC_720/a_36_216# 0.03fF
C34045 OR2X1_LOC_137/Y OR2X1_LOC_720/B 0.05fF
C37025 OR2X1_LOC_244/A OR2X1_LOC_720/B 0.07fF
C39567 OR2X1_LOC_139/a_8_216# OR2X1_LOC_720/B 0.02fF
C41590 OR2X1_LOC_123/a_8_216# OR2X1_LOC_720/B 0.47fF
C45176 OR2X1_LOC_139/a_36_216# OR2X1_LOC_720/B 0.02fF
C46491 OR2X1_LOC_204/Y OR2X1_LOC_720/B 0.03fF
C47337 OR2X1_LOC_137/a_8_216# OR2X1_LOC_720/B 0.02fF
C52422 OR2X1_LOC_720/B OR2X1_LOC_721/Y 0.39fF
C56867 OR2X1_LOC_720/B VSS 0.45fF
C20444 OR2X1_LOC_835/A OR2X1_LOC_835/a_8_216# 0.47fF
C57616 OR2X1_LOC_835/A VSS 0.15fF
C2302 OR2X1_LOC_703/B OR2X1_LOC_365/B 0.17fF
C2496 OR2X1_LOC_703/B OR2X1_LOC_468/A 0.02fF
C9205 OR2X1_LOC_703/B OR2X1_LOC_703/a_8_216# 0.07fF
C13444 OR2X1_LOC_703/B OR2X1_LOC_388/a_8_216# 0.18fF
C26689 OR2X1_LOC_703/B OR2X1_LOC_538/A 0.04fF
C31359 OR2X1_LOC_703/B OR2X1_LOC_354/A 0.01fF
C36677 OR2X1_LOC_703/B OR2X1_LOC_175/Y 0.03fF
C37681 OR2X1_LOC_703/B OR2X1_LOC_620/Y 0.01fF
C43052 OR2X1_LOC_703/B OR2X1_LOC_568/A 0.16fF
C43660 OR2X1_LOC_703/B VDD 0.24fF
C46385 OR2X1_LOC_703/B OR2X1_LOC_169/a_8_216# 0.05fF
C53007 OR2X1_LOC_703/B OR2X1_LOC_180/B 0.07fF
C54818 OR2X1_LOC_703/B OR2X1_LOC_703/A 0.16fF
C57936 OR2X1_LOC_703/B VSS 0.59fF
C413 OR2X1_LOC_201/A OR2X1_LOC_475/Y 0.02fF
C17424 OR2X1_LOC_201/A OR2X1_LOC_206/A 0.34fF
C19357 OR2X1_LOC_201/A OR2X1_LOC_392/B 0.03fF
C27203 OR2X1_LOC_201/A OR2X1_LOC_201/Y 0.07fF
C45381 OR2X1_LOC_201/A OR2X1_LOC_61/Y 0.22fF
C57473 OR2X1_LOC_201/A VSS 0.15fF
C777 OR2X1_LOC_147/B OR2X1_LOC_739/A 0.10fF
C8349 OR2X1_LOC_147/B OR2X1_LOC_563/A 0.07fF
C9642 OR2X1_LOC_147/B OR2X1_LOC_486/Y 0.08fF
C9651 OR2X1_LOC_147/B OR2X1_LOC_711/a_8_216# 0.14fF
C15876 OR2X1_LOC_147/B OR2X1_LOC_181/Y 0.05fF
C20695 OR2X1_LOC_147/B OR2X1_LOC_726/A 0.05fF
C23288 OR2X1_LOC_830/a_8_216# OR2X1_LOC_147/B 0.09fF
C28793 OR2X1_LOC_147/B OR2X1_LOC_620/Y 0.03fF
C34625 VDD OR2X1_LOC_147/B 0.80fF
C45808 OR2X1_LOC_703/A OR2X1_LOC_147/B 10.54fF
C47722 OR2X1_LOC_147/B OR2X1_LOC_465/B 0.14fF
C51635 OR2X1_LOC_147/B OR2X1_LOC_551/B 0.07fF
C55055 OR2X1_LOC_147/B OR2X1_LOC_469/B 6.63fF
C57576 OR2X1_LOC_147/B VSS -0.99fF
C901 OR2X1_LOC_703/A OR2X1_LOC_443/a_8_216# 0.04fF
C1196 OR2X1_LOC_703/A OR2X1_LOC_620/Y 0.07fF
C4399 OR2X1_LOC_703/A OR2X1_LOC_703/Y 0.01fF
C7038 VDD OR2X1_LOC_703/A 0.06fF
C16864 OR2X1_LOC_326/a_8_216# OR2X1_LOC_703/A 0.01fF
C18510 OR2X1_LOC_336/a_8_216# OR2X1_LOC_703/A 0.01fF
C19334 OR2X1_LOC_303/a_8_216# OR2X1_LOC_703/A 0.01fF
C20567 OR2X1_LOC_703/A OR2X1_LOC_353/a_8_216# 0.01fF
C21831 OR2X1_LOC_703/A OR2X1_LOC_365/B 0.35fF
C23950 OR2X1_LOC_703/A OR2X1_LOC_551/B 0.07fF
C27355 OR2X1_LOC_703/A OR2X1_LOC_469/B 0.67fF
C28635 OR2X1_LOC_703/A OR2X1_LOC_703/a_8_216# 0.01fF
C29519 OR2X1_LOC_337/A OR2X1_LOC_703/A 0.01fF
C30342 OR2X1_LOC_566/A OR2X1_LOC_703/A 0.01fF
C37937 OR2X1_LOC_703/A OR2X1_LOC_486/Y 0.03fF
C42601 OR2X1_LOC_703/A OR2X1_LOC_357/A 0.01fF
C44345 OR2X1_LOC_703/A OR2X1_LOC_181/Y 0.15fF
C46224 OR2X1_LOC_538/A OR2X1_LOC_703/A 1.36fF
C50991 OR2X1_LOC_354/A OR2X1_LOC_703/A 0.28fF
C57612 OR2X1_LOC_703/A VSS -0.23fF
C546 OR2X1_LOC_509/A OR2X1_LOC_560/A 0.04fF
C39710 OR2X1_LOC_509/a_8_216# OR2X1_LOC_509/A 0.47fF
C57684 OR2X1_LOC_509/A VSS -0.07fF
C8520 OR2X1_LOC_324/A OR2X1_LOC_739/A 0.01fF
C39789 OR2X1_LOC_324/a_8_216# OR2X1_LOC_324/A 0.47fF
C57721 OR2X1_LOC_324/A VSS 0.05fF
C5815 OR2X1_LOC_770/A OR2X1_LOC_401/a_8_216# 0.47fF
C8915 OR2X1_LOC_770/A OR2X1_LOC_770/a_8_216# 0.01fF
C31233 OR2X1_LOC_770/A OR2X1_LOC_402/Y 0.01fF
C50268 OR2X1_LOC_770/A OR2X1_LOC_770/Y 0.01fF
C58012 OR2X1_LOC_770/A VSS 0.33fF
C18589 OR2X1_LOC_623/B OR2X1_LOC_715/A 0.04fF
C35893 VDD OR2X1_LOC_623/B 0.64fF
C41060 OR2X1_LOC_623/a_8_216# OR2X1_LOC_623/B 0.08fF
C51436 OR2X1_LOC_856/B OR2X1_LOC_623/B 0.01fF
C52303 OR2X1_LOC_624/A OR2X1_LOC_623/B 0.08fF
C56688 OR2X1_LOC_623/B VSS 0.22fF
C1504 OR2X1_LOC_500/A OR2X1_LOC_844/B 0.14fF
C18004 OR2X1_LOC_632/Y OR2X1_LOC_844/B 0.02fF
C35990 OR2X1_LOC_844/B OR2X1_LOC_493/Y 0.01fF
C41191 OR2X1_LOC_844/B OR2X1_LOC_500/a_8_216# 0.08fF
C52560 OR2X1_LOC_523/Y OR2X1_LOC_844/B 0.16fF
C54709 OR2X1_LOC_844/a_8_216# OR2X1_LOC_844/B 0.07fF
C55152 OR2X1_LOC_404/Y OR2X1_LOC_844/B 0.19fF
C56447 OR2X1_LOC_844/B VSS 0.43fF
C1209 OR2X1_LOC_61/B OR2X1_LOC_61/a_8_216# 0.05fF
C15823 OR2X1_LOC_61/B OR2X1_LOC_228/Y 0.06fF
C28790 OR2X1_LOC_653/Y OR2X1_LOC_61/B -0.01fF
C49466 OR2X1_LOC_476/B OR2X1_LOC_61/B 0.01fF
C57245 OR2X1_LOC_61/B VSS 0.24fF
C41673 OR2X1_LOC_33/A OR2X1_LOC_33/a_8_216# 0.47fF
C56815 OR2X1_LOC_33/A VSS 0.15fF
C5216 OR2X1_LOC_523/Y OR2X1_LOC_523/A 0.95fF
C7933 OR2X1_LOC_404/Y OR2X1_LOC_523/A 0.16fF
C14123 OR2X1_LOC_523/A OR2X1_LOC_523/a_8_216# 0.01fF
C26917 OR2X1_LOC_632/Y OR2X1_LOC_523/A 0.05fF
C47283 OR2X1_LOC_523/A OR2X1_LOC_560/A 0.10fF
C56402 OR2X1_LOC_523/A VSS 0.13fF
C537 OR2X1_LOC_805/A OR2X1_LOC_241/B 0.07fF
C7373 OR2X1_LOC_719/Y OR2X1_LOC_241/B 0.02fF
C16589 OR2X1_LOC_833/Y OR2X1_LOC_241/B 0.01fF
C21448 OR2X1_LOC_241/a_8_216# OR2X1_LOC_241/B 0.05fF
C22416 OR2X1_LOC_241/B OR2X1_LOC_493/Y 0.10fF
C26479 OR2X1_LOC_76/Y OR2X1_LOC_241/B 0.03fF
C27041 OR2X1_LOC_675/Y OR2X1_LOC_241/B 0.01fF
C29984 OR2X1_LOC_76/a_8_216# OR2X1_LOC_241/B 0.03fF
C32435 OR2X1_LOC_241/Y OR2X1_LOC_241/B 0.23fF
C32822 OR2X1_LOC_675/a_8_216# OR2X1_LOC_241/B 0.01fF
C36249 OR2X1_LOC_440/A OR2X1_LOC_241/B 0.03fF
C42926 OR2X1_LOC_241/B OR2X1_LOC_719/a_8_216# 0.51fF
C56366 OR2X1_LOC_241/B VSS 0.46fF
C16953 OR2X1_LOC_34/B OR2X1_LOC_34/a_8_216# 0.47fF
C47716 VDD OR2X1_LOC_34/B -0.00fF
C57134 OR2X1_LOC_34/B VSS 0.16fF
C5192 VDD OR2X1_LOC_180/B 0.09fF
C8999 OR2X1_LOC_544/B OR2X1_LOC_180/B 0.01fF
C9109 OR2X1_LOC_440/a_8_216# OR2X1_LOC_180/B 0.01fF
C20160 OR2X1_LOC_468/A OR2X1_LOC_180/B 0.83fF
C33675 OR2X1_LOC_180/a_8_216# OR2X1_LOC_180/B 0.02fF
C39158 OR2X1_LOC_180/a_36_216# OR2X1_LOC_180/B 0.02fF
C56294 OR2X1_LOC_180/B VSS 0.36fF
C1873 OR2X1_LOC_538/A OR2X1_LOC_319/Y 0.22fF
C2350 OR2X1_LOC_566/A OR2X1_LOC_538/A 0.03fF
C5387 OR2X1_LOC_538/A OR2X1_LOC_805/A 0.03fF
C7407 OR2X1_LOC_538/A OR2X1_LOC_354/a_8_216# 0.01fF
C13886 OR2X1_LOC_538/A OR2X1_LOC_356/a_8_216# 0.01fF
C18468 OR2X1_LOC_538/A OR2X1_LOC_356/B 0.09fF
C22914 OR2X1_LOC_354/A OR2X1_LOC_538/A 0.37fF
C29188 OR2X1_LOC_538/A OR2X1_LOC_620/Y 0.27fF
C33835 OR2X1_LOC_854/a_8_216# OR2X1_LOC_538/A -0.00fF
C35038 VDD OR2X1_LOC_538/A 0.21fF
C40143 OR2X1_LOC_538/A OR2X1_LOC_623/a_8_216# 0.01fF
C44884 OR2X1_LOC_326/a_8_216# OR2X1_LOC_538/A 0.01fF
C46605 OR2X1_LOC_336/a_8_216# OR2X1_LOC_538/A 0.07fF
C49953 OR2X1_LOC_538/A OR2X1_LOC_365/B 1.62fF
C50582 OR2X1_LOC_856/B OR2X1_LOC_538/A 0.16fF
C51426 OR2X1_LOC_538/A OR2X1_LOC_624/A 0.18fF
C57661 OR2X1_LOC_538/A VSS 0.52fF
C1896 OR2X1_LOC_244/A OR2X1_LOC_84/A 0.04fF
C24068 OR2X1_LOC_84/A OR2X1_LOC_84/a_8_216# 0.18fF
C29761 VDD OR2X1_LOC_84/A 0.36fF
C57014 OR2X1_LOC_84/A VSS -0.02fF
C5392 OR2X1_LOC_544/a_8_216# OR2X1_LOC_544/B 0.03fF
C5787 OR2X1_LOC_440/A OR2X1_LOC_544/B 0.88fF
C28154 OR2X1_LOC_180/a_8_216# OR2X1_LOC_544/B 0.47fF
C50979 OR2X1_LOC_439/a_8_216# OR2X1_LOC_544/B 0.04fF
C56433 OR2X1_LOC_544/B VSS 0.51fF
C254 OR2X1_LOC_643/A OR2X1_LOC_392/B 0.05fF
C778 OR2X1_LOC_643/A OR2X1_LOC_624/Y 0.03fF
C1962 OR2X1_LOC_643/A OR2X1_LOC_510/a_36_216# 0.01fF
C2508 VDD OR2X1_LOC_643/A 0.29fF
C4268 OR2X1_LOC_643/A OR2X1_LOC_720/a_8_216# 0.02fF
C6176 OR2X1_LOC_643/A OR2X1_LOC_474/B 0.02fF
C8198 OR2X1_LOC_643/A OR2X1_LOC_844/Y 0.67fF
C8607 OR2X1_LOC_849/A OR2X1_LOC_643/A 0.03fF
C8997 OR2X1_LOC_643/A OR2X1_LOC_124/Y 0.03fF
C11039 OR2X1_LOC_643/A OR2X1_LOC_523/Y 0.01fF
C13297 OR2X1_LOC_844/a_8_216# OR2X1_LOC_643/A 0.01fF
C13718 OR2X1_LOC_643/A OR2X1_LOC_404/Y 0.03fF
C14044 OR2X1_LOC_643/A OR2X1_LOC_474/Y 0.01fF
C19231 OR2X1_LOC_643/A OR2X1_LOC_849/a_8_216# 0.01fF
C19612 OR2X1_LOC_216/Y OR2X1_LOC_643/A 0.48fF
C22981 OR2X1_LOC_643/A OR2X1_LOC_624/a_8_216# 0.01fF
C24425 OR2X1_LOC_643/A OR2X1_LOC_641/B 0.03fF
C29888 OR2X1_LOC_643/A OR2X1_LOC_228/Y 0.01fF
C30233 OR2X1_LOC_643/A OR2X1_LOC_849/a_36_216# -0.00fF
C30654 OR2X1_LOC_643/A OR2X1_LOC_244/A 0.07fF
C31050 OR2X1_LOC_643/A OR2X1_LOC_643/a_8_216# 0.02fF
C33530 OR2X1_LOC_643/A OR2X1_LOC_231/a_8_216# 0.03fF
C35711 OR2X1_LOC_643/A OR2X1_LOC_474/a_8_216# 0.01fF
C35717 OR2X1_LOC_643/A OR2X1_LOC_859/A 0.01fF
C35859 OR2X1_LOC_643/A OR2X1_LOC_508/Y 0.09fF
C39587 OR2X1_LOC_643/A OR2X1_LOC_786/Y 0.07fF
C44245 OR2X1_LOC_141/B OR2X1_LOC_643/A 0.03fF
C44625 OR2X1_LOC_643/A OR2X1_LOC_231/a_36_216# 0.02fF
C45520 OR2X1_LOC_643/A OR2X1_LOC_203/Y 0.07fF
C45884 OR2X1_LOC_643/A OR2X1_LOC_721/Y 0.03fF
C47094 OR2X1_LOC_643/A OR2X1_LOC_510/a_8_216# 0.02fF
C47193 OR2X1_LOC_510/A OR2X1_LOC_643/A 0.23fF
C52971 OR2X1_LOC_643/A OR2X1_LOC_560/A 0.03fF
C57583 OR2X1_LOC_643/A VSS 0.16fF
C4249 OR2X1_LOC_460/Y OR2X1_LOC_463/a_8_216# 0.39fF
C57503 OR2X1_LOC_460/Y VSS 0.18fF
C25201 AND2X1_LOC_639/A AND2X1_LOC_639/a_8_24# 0.03fF
C36154 AND2X1_LOC_639/A AND2X1_LOC_651/B 0.03fF
C41710 AND2X1_LOC_639/A AND2X1_LOC_639/a_36_24# 0.01fF
C43258 AND2X1_LOC_639/A AND2X1_LOC_639/B 0.24fF
C56803 AND2X1_LOC_639/A VSS 0.27fF
C16786 VDD OR2X1_LOC_452/A -0.00fF
C31999 OR2X1_LOC_452/A OR2X1_LOC_452/a_8_216# 0.39fF
C57572 OR2X1_LOC_452/A VSS 0.18fF
C1575 AND2X1_LOC_810/A AND2X1_LOC_702/Y 0.02fF
C15176 AND2X1_LOC_810/A AND2X1_LOC_856/A 0.01fF
C24045 AND2X1_LOC_810/A AND2X1_LOC_568/B 0.03fF
C19031 AND2X1_LOC_810/A AND2X1_LOC_337/B 0.02fF
C12077 AND2X1_LOC_810/A AND2X1_LOC_388/Y 0.01fF
C40981 AND2X1_LOC_810/A AND2X1_LOC_661/A 0.02fF
C54443 AND2X1_LOC_810/A AND2X1_LOC_170/B 0.05fF
C24014 AND2X1_LOC_773/Y AND2X1_LOC_810/A 0.30fF
C11318 AND2X1_LOC_810/A AND2X1_LOC_365/A 0.03fF
C39632 AND2X1_LOC_810/A AND2X1_LOC_392/A 0.02fF
C49270 AND2X1_LOC_810/A AND2X1_LOC_354/B 0.04fF
C39179 AND2X1_LOC_810/A AND2X1_LOC_715/Y -0.00fF
C25433 AND2X1_LOC_810/A AND2X1_LOC_863/A 0.01fF
C39696 AND2X1_LOC_810/A AND2X1_LOC_354/Y 0.01fF
C7081 AND2X1_LOC_810/A AND2X1_LOC_715/a_8_24# 0.01fF
C18484 AND2X1_LOC_810/A AND2X1_LOC_567/a_8_24# 0.01fF
C22269 AND2X1_LOC_717/B AND2X1_LOC_465/Y 0.03fF
C54386 AND2X1_LOC_721/Y AND2X1_LOC_465/Y 0.02fF
C24612 AND2X1_LOC_465/Y AND2X1_LOC_786/Y 0.01fF
C34682 AND2X1_LOC_564/B AND2X1_LOC_465/Y 0.01fF
C45538 AND2X1_LOC_851/A AND2X1_LOC_465/Y 0.04fF
C30315 AND2X1_LOC_851/B AND2X1_LOC_465/Y 0.09fF
C40149 AND2X1_LOC_465/Y AND2X1_LOC_465/A 0.16fF
C50702 VDD AND2X1_LOC_465/Y 0.16fF
C57047 AND2X1_LOC_465/Y VSS 0.28fF
C45981 AND2X1_LOC_474/A AND2X1_LOC_859/B 0.01fF
C7684 AND2X1_LOC_191/B AND2X1_LOC_859/B 0.02fF
C47735 AND2X1_LOC_719/Y AND2X1_LOC_859/B 0.05fF
C2273 AND2X1_LOC_859/Y AND2X1_LOC_859/B 0.01fF
C11169 AND2X1_LOC_859/B AND2X1_LOC_806/A 0.01fF
C3048 VDD AND2X1_LOC_859/B 0.01fF
C56827 AND2X1_LOC_859/B VSS 0.26fF
C43987 AND2X1_LOC_715/Y AND2X1_LOC_354/Y 0.01fF
C5007 AND2X1_LOC_354/Y AND2X1_LOC_356/a_8_24# 0.10fF
C48478 VDD AND2X1_LOC_354/Y 0.21fF
C36826 AND2X1_LOC_593/Y AND2X1_LOC_653/B 0.01fF
C47830 AND2X1_LOC_653/B AND2X1_LOC_810/Y 0.05fF
C42013 AND2X1_LOC_653/B AND2X1_LOC_653/a_8_24# 0.19fF
C57065 AND2X1_LOC_653/B VSS 0.07fF
C22651 AND2X1_LOC_565/Y AND2X1_LOC_474/Y 0.03fF
C10174 AND2X1_LOC_658/B AND2X1_LOC_474/Y 0.03fF
C780 AND2X1_LOC_510/A AND2X1_LOC_474/Y 0.89fF
C9238 AND2X1_LOC_574/Y AND2X1_LOC_474/Y 0.05fF
C9895 AND2X1_LOC_191/Y AND2X1_LOC_474/Y 9.02fF
C18254 AND2X1_LOC_675/Y AND2X1_LOC_474/Y 0.02fF
C4578 AND2X1_LOC_501/Y AND2X1_LOC_474/Y 0.02fF
C40179 AND2X1_LOC_658/A AND2X1_LOC_474/Y 0.03fF
C9901 AND2X1_LOC_711/Y AND2X1_LOC_474/Y 0.03fF
C15246 AND2X1_LOC_509/Y AND2X1_LOC_474/Y 0.01fF
C26294 AND2X1_LOC_510/a_8_24# AND2X1_LOC_474/Y 0.01fF
C37309 AND2X1_LOC_573/A AND2X1_LOC_474/Y 0.01fF
C47221 VDD AND2X1_LOC_474/Y 0.18fF
C51456 AND2X1_LOC_508/a_8_24# AND2X1_LOC_474/Y -0.00fF
C54982 AND2X1_LOC_474/Y AND2X1_LOC_574/A 0.39fF
C1987 OR2X1_LOC_774/Y OR2X1_LOC_773/Y 0.74fF
C1278 OR2X1_LOC_774/Y OR2X1_LOC_862/A 0.14fF
C3531 OR2X1_LOC_774/Y OR2X1_LOC_772/Y 0.17fF
C25619 OR2X1_LOC_774/Y OR2X1_LOC_773/a_8_216# 0.01fF
C38616 OR2X1_LOC_774/Y OR2X1_LOC_772/a_8_216# 0.01fF
C40663 OR2X1_LOC_774/Y OR2X1_LOC_859/a_8_216# 0.01fF
C57863 OR2X1_LOC_774/Y VSS 0.24fF
C48157 OR2X1_LOC_624/A OR2X1_LOC_510/Y 0.03fF
C12903 OR2X1_LOC_510/Y OR2X1_LOC_786/Y 0.03fF
C18742 OR2X1_LOC_510/Y OR2X1_LOC_203/Y 0.18fF
C38151 OR2X1_LOC_510/Y OR2X1_LOC_124/Y 0.18fF
C26082 OR2X1_LOC_510/Y OR2X1_LOC_560/A 0.04fF
C41501 OR2X1_LOC_510/Y OR2X1_LOC_244/B 0.05fF
C19094 OR2X1_LOC_510/Y OR2X1_LOC_721/Y 0.03fF
C29542 OR2X1_LOC_510/Y OR2X1_LOC_392/B 0.01fF
C9172 OR2X1_LOC_510/Y OR2X1_LOC_508/Y 0.01fF
C3944 OR2X1_LOC_510/Y OR2X1_LOC_244/A 0.01fF
C43259 OR2X1_LOC_474/Y OR2X1_LOC_510/Y 0.03fF
C31721 VDD OR2X1_LOC_510/Y 0.18fF
C23030 AND2X1_LOC_658/B AND2X1_LOC_574/A 0.20fF
C31014 AND2X1_LOC_675/Y AND2X1_LOC_574/A 0.43fF
C3845 VDD AND2X1_LOC_574/A 0.01fF
C13649 AND2X1_LOC_574/a_8_24# AND2X1_LOC_574/A 0.09fF
C50365 AND2X1_LOC_573/A AND2X1_LOC_574/A 0.01fF
C34937 OR2X1_LOC_844/Y OR2X1_LOC_859/A 0.01fF
C27629 OR2X1_LOC_859/A OR2X1_LOC_624/Y 0.03fF
C33097 OR2X1_LOC_859/A OR2X1_LOC_561/Y 0.10fF
C27135 OR2X1_LOC_859/A OR2X1_LOC_392/B 0.06fF
C48683 OR2X1_LOC_774/Y OR2X1_LOC_859/A 0.05fF
C29287 VDD OR2X1_LOC_859/A 0.08fF
C54907 OR2X1_LOC_859/a_8_216# OR2X1_LOC_859/A 0.05fF
C57420 OR2X1_LOC_859/A VSS -1.35fF
C27206 OR2X1_LOC_465/Y OR2X1_LOC_465/B 0.01fF
C14346 VDD OR2X1_LOC_465/Y 0.12fF
C57697 OR2X1_LOC_465/Y VSS 0.19fF
C47024 OR2X1_LOC_175/Y OR2X1_LOC_35/Y 0.02fF
C11886 OR2X1_LOC_35/B OR2X1_LOC_35/Y 0.73fF
C24469 OR2X1_LOC_648/B OR2X1_LOC_35/Y 0.03fF
C34545 OR2X1_LOC_857/B OR2X1_LOC_35/Y 0.30fF
C44127 OR2X1_LOC_208/a_8_216# OR2X1_LOC_35/Y 0.03fF
C53870 VDD OR2X1_LOC_35/Y 0.13fF
C19840 AND2X1_LOC_35/Y AND2X1_LOC_208/Y 0.01fF
C29748 AND2X1_LOC_211/B AND2X1_LOC_35/Y 0.01fF
C7598 AND2X1_LOC_208/a_8_24# AND2X1_LOC_35/Y 0.26fF
C43206 VDD AND2X1_LOC_35/Y 0.21fF
C57293 AND2X1_LOC_35/Y VSS 0.43fF
C23208 OR2X1_LOC_354/A OR2X1_LOC_356/B 0.08fF
C29505 OR2X1_LOC_620/Y OR2X1_LOC_356/B 0.02fF
C7749 OR2X1_LOC_354/a_8_216# OR2X1_LOC_356/B 0.03fF
C14219 OR2X1_LOC_356/B OR2X1_LOC_356/a_8_216# 0.08fF
C23782 OR2X1_LOC_624/A OR2X1_LOC_474/Y 0.15fF
C44695 OR2X1_LOC_474/Y OR2X1_LOC_786/Y 0.42fF
C50656 OR2X1_LOC_474/Y OR2X1_LOC_203/Y 0.07fF
C39990 OR2X1_LOC_474/Y OR2X1_LOC_140/Y 0.11fF
C5778 OR2X1_LOC_474/Y OR2X1_LOC_624/Y 0.01fF
C24979 OR2X1_LOC_508/A OR2X1_LOC_474/Y 0.07fF
C33896 OR2X1_LOC_474/Y OR2X1_LOC_805/A 0.01fF
C1829 OR2X1_LOC_474/Y OR2X1_LOC_560/A 0.03fF
C17299 OR2X1_LOC_474/Y OR2X1_LOC_244/B 0.05fF
C11268 OR2X1_LOC_474/Y OR2X1_LOC_474/B 0.03fF
C51007 OR2X1_LOC_474/Y OR2X1_LOC_721/Y 0.10fF
C13611 OR2X1_LOC_849/A OR2X1_LOC_474/Y 0.17fF
C7504 VDD OR2X1_LOC_474/Y 1.02fF
C30047 OR2X1_LOC_474/Y OR2X1_LOC_475/a_8_216# 0.01fF
C38361 OR2X1_LOC_508/a_8_216# OR2X1_LOC_474/Y 0.05fF
C51972 OR2X1_LOC_474/a_36_216# OR2X1_LOC_474/Y 0.01fF
C33318 OR2X1_LOC_653/A OR2X1_LOC_390/B 0.16fF
C25885 OR2X1_LOC_653/Y OR2X1_LOC_653/A 0.01fF
C39272 OR2X1_LOC_653/A OR2X1_LOC_392/B 0.12fF
C57707 OR2X1_LOC_653/A VSS 0.13fF
C13489 AND2X1_LOC_717/B AND2X1_LOC_465/A 0.21fF
C17146 AND2X1_LOC_465/A AND2X1_LOC_455/B 0.83fF
C46253 AND2X1_LOC_523/Y AND2X1_LOC_465/A 0.08fF
C32940 AND2X1_LOC_456/Y AND2X1_LOC_465/A 0.09fF
C45626 AND2X1_LOC_721/Y AND2X1_LOC_465/A 0.02fF
C46570 AND2X1_LOC_191/B AND2X1_LOC_465/A 0.09fF
C9083 AND2X1_LOC_465/A AND2X1_LOC_242/B 0.06fF
C30299 AND2X1_LOC_719/Y AND2X1_LOC_465/A 0.10fF
C21682 AND2X1_LOC_851/B AND2X1_LOC_465/A 0.03fF
C4506 AND2X1_LOC_465/a_36_24# AND2X1_LOC_465/A 0.01fF
C41757 VDD AND2X1_LOC_465/A 0.34fF
C28436 AND2X1_LOC_554/Y AND2X1_LOC_573/A 0.01fF
C11035 AND2X1_LOC_572/A AND2X1_LOC_573/A 0.06fF
C19458 AND2X1_LOC_573/A AND2X1_LOC_404/B 0.91fF
C14103 AND2X1_LOC_717/B AND2X1_LOC_573/A 0.01fF
C31312 AND2X1_LOC_561/B AND2X1_LOC_573/A 0.03fF
C2649 AND2X1_LOC_141/B AND2X1_LOC_573/A 0.03fF
C42842 AND2X1_LOC_486/Y AND2X1_LOC_573/A 0.03fF
C7278 AND2X1_LOC_849/A AND2X1_LOC_573/A 0.02fF
C33558 AND2X1_LOC_456/Y AND2X1_LOC_573/A 0.03fF
C46761 AND2X1_LOC_850/A AND2X1_LOC_573/A 0.03fF
C13949 AND2X1_LOC_563/A AND2X1_LOC_573/A 0.01fF
C46184 AND2X1_LOC_721/Y AND2X1_LOC_573/A 0.02fF
C5343 AND2X1_LOC_658/B AND2X1_LOC_573/A 0.36fF
C40894 AND2X1_LOC_571/B AND2X1_LOC_573/A 0.03fF
C52255 AND2X1_LOC_510/A AND2X1_LOC_573/A 0.01fF
C54040 AND2X1_LOC_852/Y AND2X1_LOC_573/A 0.07fF
C41062 AND2X1_LOC_141/A AND2X1_LOC_573/A 0.01fF
C6584 AND2X1_LOC_573/A AND2X1_LOC_244/A 0.03fF
C45031 AND2X1_LOC_573/A AND2X1_LOC_403/B 0.09fF
C29202 AND2X1_LOC_474/A AND2X1_LOC_573/A 0.16fF
C2493 AND2X1_LOC_772/B AND2X1_LOC_573/A 0.01fF
C13988 AND2X1_LOC_456/B AND2X1_LOC_573/A 0.04fF
C47181 AND2X1_LOC_191/B AND2X1_LOC_573/A 0.07fF
C36484 AND2X1_LOC_554/B AND2X1_LOC_573/A 0.15fF
C17095 AND2X1_LOC_656/Y AND2X1_LOC_573/A 0.03fF
C30857 AND2X1_LOC_719/Y AND2X1_LOC_573/A 0.10fF
C13543 AND2X1_LOC_675/Y AND2X1_LOC_573/A 0.02fF
C56056 AND2X1_LOC_501/Y AND2X1_LOC_573/A 0.27fF
C46704 AND2X1_LOC_508/B AND2X1_LOC_573/A 0.02fF
C38445 AND2X1_LOC_392/A AND2X1_LOC_573/A 0.07fF
C35500 AND2X1_LOC_658/A AND2X1_LOC_573/A 0.03fF
C33681 AND2X1_LOC_573/A AND2X1_LOC_647/Y 0.02fF
C10559 AND2X1_LOC_509/Y AND2X1_LOC_573/A 0.57fF
C26174 AND2X1_LOC_340/Y AND2X1_LOC_573/A 0.02fF
C17231 AND2X1_LOC_573/A AND2X1_LOC_772/Y 0.02fF
C8447 AND2X1_LOC_573/A AND2X1_LOC_403/a_8_24# 0.01fF
C11203 AND2X1_LOC_573/A AND2X1_LOC_772/a_8_24# 0.01fF
C25796 AND2X1_LOC_558/a_8_24# AND2X1_LOC_573/A 0.01fF
C29111 AND2X1_LOC_573/A AND2X1_LOC_456/a_8_24# 0.04fF
C33820 AND2X1_LOC_340/a_8_24# AND2X1_LOC_573/A 0.01fF
C46719 AND2X1_LOC_508/a_8_24# AND2X1_LOC_573/A 0.01fF
C50433 AND2X1_LOC_573/A AND2X1_LOC_656/a_8_24# 0.01fF
C44647 OR2X1_LOC_456/Y OR2X1_LOC_465/B 0.04fF
C8892 VDD OR2X1_LOC_465/B -0.00fF
C57314 OR2X1_LOC_465/B VSS 0.10fF
C26609 OR2X1_LOC_404/Y OR2X1_LOC_501/A 0.03fF
C23483 OR2X1_LOC_404/Y OR2X1_LOC_624/A 0.03fF
C30806 OR2X1_LOC_404/Y OR2X1_LOC_735/B 0.14fF
C32285 OR2X1_LOC_137/Y OR2X1_LOC_404/Y -0.00fF
C53120 OR2X1_LOC_404/Y OR2X1_LOC_720/Y 0.01fF
C15727 OR2X1_LOC_404/Y OR2X1_LOC_523/Y 0.14fF
C30580 OR2X1_LOC_404/Y OR2X1_LOC_575/A 0.03fF
C1503 OR2X1_LOC_404/Y OR2X1_LOC_560/A 0.03fF
C55506 OR2X1_LOC_404/Y OR2X1_LOC_493/Y 0.10fF
C10947 OR2X1_LOC_404/Y OR2X1_LOC_474/B 0.07fF
C13312 OR2X1_LOC_849/A OR2X1_LOC_404/Y 2.15fF
C4939 OR2X1_LOC_404/Y OR2X1_LOC_392/B 0.05fF
C37283 OR2X1_LOC_404/Y OR2X1_LOC_632/Y 0.19fF
C18754 OR2X1_LOC_404/Y OR2X1_LOC_474/Y 0.05fF
C9036 OR2X1_LOC_404/Y OR2X1_LOC_720/a_8_216# 0.01fF
C13541 OR2X1_LOC_404/Y OR2X1_LOC_721/a_8_216# 0.01fF
C19821 OR2X1_LOC_404/Y OR2X1_LOC_501/a_8_216# 0.02fF
C671 VDD OR2X1_LOC_833/a_8_216# 0.21fF
C1783 VDD OR2X1_LOC_544/a_8_216# 0.21fF
C5218 AND2X1_LOC_734/a_8_24# VDD -0.00fF
C8009 VDD OR2X1_LOC_642/a_8_216# 0.21fF
C8450 AND2X1_LOC_730/a_8_24# AND2X1_LOC_209/a_8_24# 0.23fF
C10241 OR2X1_LOC_475/a_8_216# OR2X1_LOC_216/a_8_216# 0.47fF
C10834 OR2X1_LOC_852/a_8_216# VDD -0.00fF
C12140 OR2X1_LOC_339/a_8_216# VDD 0.21fF
C13228 VDD OR2X1_LOC_243/a_8_216# 0.21fF
C13468 OR2X1_LOC_349/a_8_216# OR2X1_LOC_850/a_8_216# 0.47fF
C13527 AND2X1_LOC_710/a_8_24# VDD -0.00fF
C14805 AND2X1_LOC_840/a_8_24# AND2X1_LOC_833/a_8_24# 0.23fF
C15451 AND2X1_LOC_632/a_8_24# AND2X1_LOC_623/a_8_24# 0.23fF
C16439 VDD OR2X1_LOC_640/a_8_216# 0.21fF
C18061 VDD OR2X1_LOC_786/a_8_216# 0.21fF
C18501 OR2X1_LOC_338/a_8_216# VDD 0.21fF
C19021 VDD OR2X1_LOC_404/a_8_216# 0.21fF
C19456 VDD OR2X1_LOC_652/a_8_216# 0.21fF
C21527 AND2X1_LOC_180/a_8_24# VDD -0.00fF
C21759 OR2X1_LOC_303/a_8_216# OR2X1_LOC_353/a_8_216# 0.47fF
C21850 AND2X1_LOC_388/a_8_24# AND2X1_LOC_810/a_8_24# 0.23fF
C21880 VDD OR2X1_LOC_388/a_8_216# 0.21fF
C23172 OR2X1_LOC_791/a_8_216# OR2X1_LOC_792/a_8_216# 0.47fF
C23207 OR2X1_LOC_854/a_8_216# OR2X1_LOC_354/a_8_216# 0.47fF
C23280 VDD AND2X1_LOC_194/a_8_24# -0.00fF
C24517 VDD AND2X1_LOC_839/a_8_24# -0.00fF
C24768 AND2X1_LOC_392/a_8_24# AND2X1_LOC_845/a_8_24# 0.23fF
C25188 AND2X1_LOC_786/a_8_24# AND2X1_LOC_204/a_8_24# 0.23fF
C26737 VDD OR2X1_LOC_656/a_8_216# 0.21fF
C27556 VDD OR2X1_LOC_636/a_8_216# 0.21fF
C29643 VDD OR2X1_LOC_651/a_8_216# 0.21fF
C30076 AND2X1_LOC_555/a_8_24# AND2X1_LOC_345/a_8_24# 0.23fF
C30414 AND2X1_LOC_540/a_8_24# VDD -0.00fF
C35443 AND2X1_LOC_510/a_8_24# AND2X1_LOC_508/a_8_24# 0.23fF
C39819 VDD AND2X1_LOC_639/a_8_24# -0.00fF
C42388 VDD OR2X1_LOC_208/a_8_216# 0.21fF
C42588 VDD OR2X1_LOC_558/a_8_216# 0.21fF
C42794 OR2X1_LOC_346/a_8_216# VDD 0.21fF
C42796 VDD OR2X1_LOC_465/a_8_216# 0.21fF
C45008 VDD OR2X1_LOC_605/a_8_216# 0.21fF
C45283 VDD OR2X1_LOC_679/a_8_216# 0.21fF
C46072 OR2X1_LOC_474/a_8_216# OR2X1_LOC_849/a_8_216# 0.47fF
C47021 VDD AND2X1_LOC_636/a_8_24# -0.00fF
C47202 VDD OR2X1_LOC_845/a_8_216# 0.21fF
C47672 VDD OR2X1_LOC_646/a_8_216# 0.21fF
C50007 VDD AND2X1_LOC_204/a_8_24# -0.00fF
C52021 VDD OR2X1_LOC_76/a_8_216# 0.21fF
C54252 OR2X1_LOC_124/a_8_216# VDD 0.21fF
C55590 AND2X1_LOC_500/a_8_24# AND2X1_LOC_242/a_8_24# 0.23fF
C55782 AND2X1_LOC_715/a_8_24# AND2X1_LOC_354/a_8_24# 0.23fF
C56275 AND2X1_LOC_228/a_8_24# VSS 0.10fF
C56357 AND2X1_LOC_793/a_8_24# VSS 0.10fF
C56393 AND2X1_LOC_770/a_8_24# VSS 0.10fF
C56394 AND2X1_LOC_792/a_8_24# VSS 0.10fF
C56458 AND2X1_LOC_202/a_8_24# VSS 0.10fF
C56743 AND2X1_LOC_455/a_8_24# VSS 0.10fF
C56789 AND2X1_LOC_476/a_8_24# VSS 0.10fF
C56957 AND2X1_LOC_440/a_8_24# VSS 0.10fF
C57008 AND2X1_LOC_675/a_8_24# VSS 0.10fF
C57010 AND2X1_LOC_620/a_8_24# VSS 0.10fF
C57094 AND2X1_LOC_844/a_8_24# VSS 0.10fF
C57180 AND2X1_LOC_842/a_8_24# VSS 0.10fF
C57227 AND2X1_LOC_137/a_8_24# VSS 0.10fF
C57237 AND2X1_LOC_841/a_8_24# VSS 0.10fF
C57240 AND2X1_LOC_852/a_8_24# VSS 0.10fF
C57353 AND2X1_LOC_338/a_8_24# VSS 0.10fF
C57389 AND2X1_LOC_123/a_8_24# VSS 0.10fF
C57412 AND2X1_LOC_326/a_8_24# VSS 0.10fF
C57427 AND2X1_LOC_507/a_8_24# VSS 0.10fF
C57643 AND2X1_LOC_174/a_8_24# VSS 0.10fF
C57656 AND2X1_LOC_84/a_8_24# VSS 0.10fF
C57690 AND2X1_LOC_728/a_8_24# VSS 0.10fF
C57728 AND2X1_LOC_343/a_8_24# VSS 0.10fF
C57757 AND2X1_LOC_716/a_8_24# VSS 0.10fF
C57760 AND2X1_LOC_705/a_8_24# VSS 0.10fF
C57926 AND2X1_LOC_702/a_8_24# VSS 0.10fF
C57954 AND2X1_LOC_542/a_8_24# VSS 0.10fF
C57976 AND2X1_LOC_190/a_8_24# VSS 0.10fF
C58049 AND2X1_LOC_710/a_8_24# VSS 0.10fF
C58073 AND2X1_LOC_550/a_8_24# VSS 0.10fF
C58102 AND2X1_LOC_390/a_8_24# VSS 0.10fF
C58123 AND2X1_LOC_774/a_8_24# VSS 0.10fF
C14820 OR2X1_LOC_216/A OR2X1_LOC_624/A 0.33fF
C35706 OR2X1_LOC_216/A OR2X1_LOC_786/Y 0.14fF
C41534 OR2X1_LOC_216/A OR2X1_LOC_203/Y 0.01fF
C8014 OR2X1_LOC_216/A OR2X1_LOC_737/A 0.01fF
C16041 OR2X1_LOC_508/A OR2X1_LOC_216/A 0.03fF
C25027 OR2X1_LOC_216/A OR2X1_LOC_805/A 0.03fF
C49110 OR2X1_LOC_216/A OR2X1_LOC_560/A 0.02fF
C41911 OR2X1_LOC_216/A OR2X1_LOC_721/Y 0.03fF
C52581 OR2X1_LOC_216/A OR2X1_LOC_392/B 0.10fF
C31963 OR2X1_LOC_216/A OR2X1_LOC_508/Y 0.06fF
C10123 OR2X1_LOC_216/A OR2X1_LOC_474/Y 0.21fF
C46379 OR2X1_LOC_216/A OR2X1_LOC_216/a_8_216# 0.08fF
C53126 OR2X1_LOC_216/A OR2X1_LOC_734/a_8_216# 0.03fF
C36784 AND2X1_LOC_216/Y AND2X1_LOC_116/Y 0.02fF
C51039 AND2X1_LOC_392/A AND2X1_LOC_116/Y 0.03fF
C24743 AND2X1_LOC_560/B AND2X1_LOC_116/Y 0.03fF
C34754 OR2X1_LOC_624/A OR2X1_LOC_539/Y 0.03fF
C17204 OR2X1_LOC_539/Y OR2X1_LOC_174/Y 0.02fF
C11741 OR2X1_LOC_175/Y OR2X1_LOC_539/Y 0.10fF
C33409 OR2X1_LOC_468/A OR2X1_LOC_539/Y 0.27fF
C45046 OR2X1_LOC_805/A OR2X1_LOC_539/Y 0.03fF
C28240 OR2X1_LOC_539/Y OR2X1_LOC_175/a_8_216# 0.01fF
C12016 OR2X1_LOC_175/Y OR2X1_LOC_319/Y 0.03fF
C6498 OR2X1_LOC_354/A OR2X1_LOC_319/Y 0.13fF
C12991 OR2X1_LOC_620/Y OR2X1_LOC_319/Y 0.01fF
C34123 OR2X1_LOC_856/B OR2X1_LOC_319/Y 0.83fF
C19251 AND2X1_LOC_365/A AND2X1_LOC_798/A 0.26fF
C47833 AND2X1_LOC_354/Y AND2X1_LOC_798/A 0.01fF
C42878 AND2X1_LOC_810/A AND2X1_LOC_798/A 0.01fF
C35288 AND2X1_LOC_354/a_8_24# AND2X1_LOC_798/A 0.01fF
C6184 AND2X1_LOC_539/Y AND2X1_LOC_337/B 0.01fF
C55476 AND2X1_LOC_388/Y AND2X1_LOC_539/Y 0.01fF
C28306 AND2X1_LOC_539/Y AND2X1_LOC_661/A 0.53fF
C41515 AND2X1_LOC_539/Y AND2X1_LOC_170/B 0.12fF
C54694 AND2X1_LOC_539/Y AND2X1_LOC_365/A 0.01fF
C26457 AND2X1_LOC_539/Y AND2X1_LOC_715/Y 0.03fF
C28408 AND2X1_LOC_539/Y AND2X1_LOC_810/Y 0.20fF
C22302 AND2X1_LOC_810/A AND2X1_LOC_539/Y 0.03fF
C6570 AND2X1_LOC_539/Y AND2X1_LOC_388/a_8_24# 0.01fF
C22337 AND2X1_LOC_539/Y AND2X1_LOC_567/a_36_24# 0.01fF
C43558 AND2X1_LOC_539/Y AND2X1_LOC_356/a_8_24# 0.01fF
C51380 AND2X1_LOC_539/Y AND2X1_LOC_336/a_8_24# 0.01fF
C51057 VDD AND2X1_LOC_651/B 0.17fF
C56578 AND2X1_LOC_651/B VSS 0.21fF
C14060 OR2X1_LOC_641/a_8_216# OR2X1_LOC_643/Y 0.01fF
C12853 OR2X1_LOC_500/a_8_216# OR2X1_LOC_501/A -0.00fF
C15443 VDD OR2X1_LOC_501/A -0.00fF
C28086 OR2X1_LOC_501/A OR2X1_LOC_501/a_8_216# 0.39fF
C38794 OR2X1_LOC_575/A OR2X1_LOC_501/A 0.19fF
C45663 OR2X1_LOC_632/Y OR2X1_LOC_501/A 0.03fF
C56446 OR2X1_LOC_501/A VSS 0.18fF
C1693 VDD OR2X1_LOC_844/Y 0.05fF
C10279 OR2X1_LOC_844/Y OR2X1_LOC_523/Y 0.01fF
C18423 OR2X1_LOC_844/Y OR2X1_LOC_849/a_8_216# 0.02fF
C29420 OR2X1_LOC_844/Y OR2X1_LOC_849/a_36_216# 0.02fF
C52141 OR2X1_LOC_844/Y OR2X1_LOC_560/A 0.09fF
C55646 OR2X1_LOC_844/Y OR2X1_LOC_392/B 0.07fF
C56214 OR2X1_LOC_844/Y OR2X1_LOC_624/Y 0.33fF
C57421 OR2X1_LOC_844/Y VSS 0.03fF
C3878 OR2X1_LOC_624/A OR2X1_LOC_216/a_8_216# 0.14fF
C5275 OR2X1_LOC_175/Y OR2X1_LOC_624/A 0.29fF
C6271 OR2X1_LOC_620/Y OR2X1_LOC_624/A 0.52fF
C6470 OR2X1_LOC_624/A OR2X1_LOC_560/A 0.05fF
C9443 OR2X1_LOC_624/A OR2X1_LOC_216/a_36_216# 0.15fF
C10830 OR2X1_LOC_624/A OR2X1_LOC_174/Y 0.04fF
C12216 VDD OR2X1_LOC_624/A 2.15fF
C15944 OR2X1_LOC_624/A OR2X1_LOC_474/B 0.02fF
C17061 OR2X1_LOC_476/B OR2X1_LOC_624/A 0.01fF
C17373 OR2X1_LOC_623/a_8_216# OR2X1_LOC_624/A 0.02fF
C18296 OR2X1_LOC_849/A OR2X1_LOC_624/A 0.01fF
C21921 OR2X1_LOC_624/A OR2X1_LOC_175/a_8_216# 0.03fF
C22071 OR2X1_LOC_624/A OR2X1_LOC_244/B 0.07fF
C27539 OR2X1_LOC_856/B OR2X1_LOC_624/A 0.13fF
C29653 OR2X1_LOC_508/A OR2X1_LOC_624/A 0.10fF
C35982 OR2X1_LOC_624/A OR2X1_LOC_61/Y 0.10fF
C38541 OR2X1_LOC_624/A OR2X1_LOC_805/A 3.90fF
C39601 OR2X1_LOC_624/A OR2X1_LOC_228/Y 0.10fF
C44785 OR2X1_LOC_624/A OR2X1_LOC_140/Y 0.05fF
C45555 OR2X1_LOC_474/a_8_216# OR2X1_LOC_624/A 0.13fF
C45692 OR2X1_LOC_624/A OR2X1_LOC_508/Y 0.05fF
C49545 OR2X1_LOC_624/A OR2X1_LOC_786/Y 0.10fF
C52743 OR2X1_LOC_653/Y OR2X1_LOC_624/A 0.10fF
C55326 OR2X1_LOC_624/A OR2X1_LOC_203/Y 0.10fF
C55678 OR2X1_LOC_624/A OR2X1_LOC_721/Y 0.10fF
C57451 OR2X1_LOC_624/A VSS 1.10fF
C1889 OR2X1_LOC_337/A OR2X1_LOC_182/B 0.02fF
C2818 OR2X1_LOC_337/A OR2X1_LOC_337/a_8_216# 0.18fF
C13862 OR2X1_LOC_337/A OR2X1_LOC_352/A 0.37fF
C18488 OR2X1_LOC_337/A VDD 0.06fF
C33115 OR2X1_LOC_337/A OR2X1_LOC_365/B 0.44fF
C41733 OR2X1_LOC_566/A OR2X1_LOC_337/A 0.74fF
C58068 OR2X1_LOC_337/A VSS 0.17fF
C7378 OR2X1_LOC_201/a_8_216# OR2X1_LOC_201/Y 0.02fF
C25521 OR2X1_LOC_61/Y OR2X1_LOC_201/Y 0.13fF
C13829 OR2X1_LOC_775/a_8_216# OR2X1_LOC_390/B -0.02fF
C28244 OR2X1_LOC_653/Y OR2X1_LOC_390/B 0.04fF
C30660 OR2X1_LOC_390/a_8_216# OR2X1_LOC_390/B 0.13fF
C48870 OR2X1_LOC_476/B OR2X1_LOC_390/B 0.05fF
C55159 OR2X1_LOC_653/a_8_216# OR2X1_LOC_390/B 0.05fF
C56293 OR2X1_LOC_390/B VSS 0.43fF
C1785 OR2X1_LOC_703/Y OR2X1_LOC_714/a_8_216# 0.06fF
C15480 OR2X1_LOC_739/A OR2X1_LOC_703/Y 0.02fF
C23440 OR2X1_LOC_703/Y OR2X1_LOC_724/A 0.01fF
C37044 OR2X1_LOC_354/A OR2X1_LOC_703/Y 0.02fF
C43511 OR2X1_LOC_620/Y OR2X1_LOC_703/Y 0.01fF
C49587 VDD OR2X1_LOC_703/Y 0.16fF
C56463 OR2X1_LOC_703/Y VSS 0.44fF
C17703 OR2X1_LOC_799/A OR2X1_LOC_468/A 0.11fF
C52162 OR2X1_LOC_175/Y OR2X1_LOC_799/A 0.14fF
C35622 OR2X1_LOC_774/B OR2X1_LOC_773/Y 0.08fF
C42142 OR2X1_LOC_773/Y OR2X1_LOC_774/a_8_216# 0.08fF
C56783 OR2X1_LOC_773/Y VSS 0.11fF
C5546 OR2X1_LOC_401/a_36_216# OR2X1_LOC_402/Y 0.01fF
C7984 VDD OR2X1_LOC_402/Y 0.62fF
C12373 OR2X1_LOC_402/a_8_216# OR2X1_LOC_402/Y 0.01fF
C23468 OR2X1_LOC_402/a_36_216# OR2X1_LOC_402/Y -0.00fF
C30972 OR2X1_LOC_402/Y OR2X1_LOC_404/a_8_216# 0.03fF
C36521 OR2X1_LOC_404/A OR2X1_LOC_402/Y 0.18fF
C50761 OR2X1_LOC_401/a_8_216# OR2X1_LOC_402/Y 0.05fF
C51960 OR2X1_LOC_401/Y OR2X1_LOC_402/Y 0.03fF
C57109 OR2X1_LOC_402/Y VSS 0.24fF
C32365 OR2X1_LOC_555/a_8_216# OR2X1_LOC_562/B -0.00fF
C6161 OR2X1_LOC_191/a_8_216# OR2X1_LOC_192/A -0.00fF
C34574 VDD OR2X1_LOC_192/A -0.00fF
C45586 OR2X1_LOC_192/A OR2X1_LOC_192/a_8_216# 0.39fF
C51323 OR2X1_LOC_565/A OR2X1_LOC_192/A 0.05fF
C56534 OR2X1_LOC_192/A VSS 0.18fF
C2858 OR2X1_LOC_170/A OR2X1_LOC_175/Y 0.07fF
C9128 OR2X1_LOC_170/A OR2X1_LOC_568/A 0.05fF
C9730 OR2X1_LOC_170/A VDD -0.00fF
C24415 OR2X1_LOC_170/A OR2X1_LOC_365/B 0.01fF
C51344 OR2X1_LOC_170/A OR2X1_LOC_170/a_8_216# 0.39fF
C57935 OR2X1_LOC_170/A VSS 0.18fF
C2290 OR2X1_LOC_726/A OR2X1_LOC_469/B 0.09fF
C4071 OR2X1_LOC_711/A OR2X1_LOC_469/B 0.04fF
C10429 OR2X1_LOC_620/Y OR2X1_LOC_469/B 0.03fF
C47425 OR2X1_LOC_711/a_8_216# OR2X1_LOC_469/B 0.02fF
C9872 OR2X1_LOC_123/a_8_216# OR2X1_LOC_786/Y 0.01fF
C14161 OR2X1_LOC_786/Y OR2X1_LOC_785/B 0.03fF
C20526 OR2X1_LOC_786/Y OR2X1_LOC_721/Y 0.03fF
C26382 OR2X1_LOC_124/A OR2X1_LOC_786/Y 0.01fF
C30978 OR2X1_LOC_786/Y OR2X1_LOC_392/B 0.01fF
C35228 OR2X1_LOC_124/a_8_216# OR2X1_LOC_786/Y 0.01fF
C35369 OR2X1_LOC_241/Y OR2X1_LOC_786/Y 0.10fF
C4959 OR2X1_LOC_641/Y OR2X1_LOC_642/a_8_216# 0.03fF
C4269 OR2X1_LOC_174/Y OR2X1_LOC_175/a_8_216# 0.18fF
C21046 OR2X1_LOC_805/A OR2X1_LOC_174/Y 0.03fF
C50839 VDD OR2X1_LOC_174/Y 0.04fF
C56241 OR2X1_LOC_174/Y VSS 0.10fF
C25373 OR2X1_LOC_833/Y OR2X1_LOC_203/Y 0.01fF
C26290 OR2X1_LOC_203/Y OR2X1_LOC_721/Y 0.10fF
C31136 OR2X1_LOC_203/Y OR2X1_LOC_493/Y 0.10fF
C36690 OR2X1_LOC_203/Y OR2X1_LOC_392/B 0.10fF
C43727 OR2X1_LOC_833/a_8_216# OR2X1_LOC_203/Y 0.04fF
C30664 OR2X1_LOC_175/Y OR2X1_LOC_170/a_8_216# 0.05fF
C32292 OR2X1_LOC_175/Y OR2X1_LOC_539/B 0.01fF
C33570 OR2X1_LOC_175/Y OR2X1_LOC_567/a_8_216# 0.05fF
C35461 OR2X1_LOC_175/Y OR2X1_LOC_208/a_8_216# 0.01fF
C47993 OR2X1_LOC_169/a_8_216# OR2X1_LOC_175/Y 0.04fF
C54971 OR2X1_LOC_175/Y OR2X1_LOC_175/a_8_216# 0.01fF
C19829 OR2X1_LOC_337/a_8_216# OR2X1_LOC_182/B 0.01fF
C23852 VDD OR2X1_LOC_835/Y 0.04fF
C57358 OR2X1_LOC_835/Y VSS 0.14fF
C21963 OR2X1_LOC_123/a_8_216# OR2X1_LOC_124/A 0.01fF
C45297 OR2X1_LOC_124/A VDD 0.05fF
C58027 OR2X1_LOC_124/A VSS 0.22fF
C37839 OR2X1_LOC_347/a_8_216# OR2X1_LOC_675/Y 0.04fF
C39143 OR2X1_LOC_850/B OR2X1_LOC_675/Y 0.03fF
C43436 OR2X1_LOC_347/a_36_216# OR2X1_LOC_675/Y 0.02fF
C45216 OR2X1_LOC_76/Y OR2X1_LOC_675/Y 0.01fF
C1981 OR2X1_LOC_551/B OR2X1_LOC_545/a_8_216# 0.01fF
C6546 OR2X1_LOC_443/a_8_216# OR2X1_LOC_551/B 0.05fF
C7437 OR2X1_LOC_443/Y OR2X1_LOC_551/B 0.01fF
C2183 VDD OR2X1_LOC_440/A 0.10fF
C4795 OR2X1_LOC_675/a_8_216# OR2X1_LOC_440/A 0.07fF
C11573 OR2X1_LOC_440/A OR2X1_LOC_737/A 0.02fF
C19274 OR2X1_LOC_440/A OR2X1_LOC_787/Y 0.07fF
C30553 OR2X1_LOC_440/A OR2X1_LOC_180/a_8_216# 0.02fF
C53391 OR2X1_LOC_439/a_8_216# OR2X1_LOC_440/A 0.01fF
C57001 OR2X1_LOC_440/A VSS 0.57fF
C6935 AND2X1_LOC_554/Y AND2X1_LOC_772/a_8_24# 0.20fF
C32233 AND2X1_LOC_554/Y AND2X1_LOC_554/B 0.02fF
C47976 AND2X1_LOC_554/Y AND2X1_LOC_554/a_8_24# 0.03fF
C54347 AND2X1_LOC_554/Y AND2X1_LOC_772/B 0.39fF
C31221 AND2X1_LOC_728/Y AND2X1_LOC_209/Y 0.01fF
C55934 OR2X1_LOC_679/Y AND2X1_LOC_209/Y 0.80fF
C5571 AND2X1_LOC_572/A AND2X1_LOC_845/Y 0.01fF
C14939 AND2X1_LOC_554/B AND2X1_LOC_572/A 0.34fF
C16901 AND2X1_LOC_392/A AND2X1_LOC_572/A 0.03fF
C30391 AND2X1_LOC_554/a_8_24# AND2X1_LOC_572/A 0.15fF
C31448 AND2X1_LOC_140/a_8_24# AND2X1_LOC_572/A 0.01fF
C34318 AND2X1_LOC_123/Y AND2X1_LOC_572/A 0.81fF
C36756 AND2X1_LOC_772/B AND2X1_LOC_572/A 0.28fF
C45654 AND2X1_LOC_572/A AND2X1_LOC_772/a_8_24# 0.01fF
C51767 AND2X1_LOC_572/A AND2X1_LOC_772/Y 0.01fF
C12580 AND2X1_LOC_347/Y AND2X1_LOC_347/B 0.11fF
C33935 AND2X1_LOC_347/Y AND2X1_LOC_259/Y 0.03fF
C36838 AND2X1_LOC_347/Y AND2X1_LOC_347/a_8_24# 0.06fF
C43612 AND2X1_LOC_710/Y AND2X1_LOC_347/Y 0.17fF
C29094 VDD AND2X1_LOC_404/B 0.02fF
C34690 AND2X1_LOC_404/B AND2X1_LOC_404/a_8_24# 0.01fF
C51333 AND2X1_LOC_403/a_8_24# AND2X1_LOC_404/B 0.01fF
C56577 AND2X1_LOC_404/B VSS 0.08fF
C18630 AND2X1_LOC_388/Y AND2X1_LOC_645/A 0.09fF
C35116 AND2X1_LOC_390/a_8_24# AND2X1_LOC_645/A 0.03fF
C36868 AND2X1_LOC_593/Y AND2X1_LOC_645/A 0.12fF
C44500 AND2X1_LOC_788/a_8_24# AND2X1_LOC_645/A 0.03fF
C7465 AND2X1_LOC_705/Y AND2X1_LOC_722/A 0.15fF
C28313 AND2X1_LOC_705/Y AND2X1_LOC_593/Y 0.07fF
C28356 AND2X1_LOC_705/Y AND2X1_LOC_602/a_8_24# 0.10fF
C41326 AND2X1_LOC_705/Y VDD 0.21fF
C41759 AND2X1_LOC_705/Y AND2X1_LOC_713/a_8_24# 0.09fF
C57924 AND2X1_LOC_705/Y VSS -0.59fF
C10340 AND2X1_LOC_76/Y AND2X1_LOC_204/Y 0.03fF
C39446 AND2X1_LOC_84/Y AND2X1_LOC_204/Y 0.01fF
C4306 AND2X1_LOC_702/Y AND2X1_LOC_326/A 0.01fF
C6880 AND2X1_LOC_702/Y AND2X1_LOC_537/Y 0.03fF
C10140 VDD AND2X1_LOC_702/Y 0.28fF
C15719 AND2X1_LOC_702/Y AND2X1_LOC_354/B 0.06fF
C29745 AND2X1_LOC_702/Y AND2X1_LOC_715/a_8_24# 0.11fF
C32984 AND2X1_LOC_702/Y AND2X1_LOC_353/a_8_24# 0.01fF
C46666 AND2X1_LOC_773/Y AND2X1_LOC_702/Y 0.03fF
C48259 AND2X1_LOC_702/Y AND2X1_LOC_863/A 0.02fF
C49508 AND2X1_LOC_702/Y AND2X1_LOC_324/a_8_24# 0.01fF
C57822 AND2X1_LOC_702/Y VSS 0.05fF
C3573 AND2X1_LOC_851/B AND2X1_LOC_717/B 0.07fF
C7972 AND2X1_LOC_564/B AND2X1_LOC_717/B 0.10fF
C12257 AND2X1_LOC_719/Y AND2X1_LOC_717/B 0.03fF
C17360 AND2X1_LOC_190/a_8_24# AND2X1_LOC_717/B 0.03fF
C23796 VDD AND2X1_LOC_717/B 0.19fF
C24272 AND2X1_LOC_486/Y AND2X1_LOC_717/B 0.18fF
C25982 AND2X1_LOC_465/a_8_24# AND2X1_LOC_717/B 0.01fF
C27471 AND2X1_LOC_721/Y AND2X1_LOC_717/B 0.06fF
C44707 AND2X1_LOC_849/A AND2X1_LOC_717/B 0.03fF
C47145 AND2X1_LOC_717/B AND2X1_LOC_242/B 0.02fF
C53930 AND2X1_LOC_717/B AND2X1_LOC_786/Y 0.09fF
C57049 AND2X1_LOC_717/B VSS -0.59fF
C20396 AND2X1_LOC_468/B AND2X1_LOC_593/Y 0.04fF
C3107 AND2X1_LOC_647/B AND2X1_LOC_647/a_8_24# 0.01fF
C7711 VDD AND2X1_LOC_647/B 0.03fF
C8377 AND2X1_LOC_646/a_8_24# AND2X1_LOC_647/B 0.01fF
C55147 AND2X1_LOC_647/Y AND2X1_LOC_647/B 1.20fF
C56810 AND2X1_LOC_647/B VSS 0.17fF
C2129 AND2X1_LOC_559/a_8_24# AND2X1_LOC_76/Y 0.01fF
C4758 AND2X1_LOC_76/Y AND2X1_LOC_203/Y 0.03fF
C7638 AND2X1_LOC_560/B AND2X1_LOC_76/Y 0.01fF
C11740 AND2X1_LOC_76/Y AND2X1_LOC_786/Y 0.34fF
C13036 AND2X1_LOC_76/Y AND2X1_LOC_455/B 0.04fF
C17509 AND2X1_LOC_76/Y AND2X1_LOC_851/B 0.14fF
C17758 AND2X1_LOC_76/a_8_24# AND2X1_LOC_76/Y 0.02fF
C18094 AND2X1_LOC_773/Y AND2X1_LOC_76/Y 0.03fF
C21556 AND2X1_LOC_340/Y AND2X1_LOC_76/Y 0.03fF
C21566 AND2X1_LOC_181/Y AND2X1_LOC_76/Y 0.03fF
C27534 AND2X1_LOC_523/a_8_24# AND2X1_LOC_76/Y 0.01fF
C33808 AND2X1_LOC_392/A AND2X1_LOC_76/Y 0.03fF
C37577 VDD AND2X1_LOC_76/Y 0.26fF
C42055 AND2X1_LOC_76/Y AND2X1_LOC_523/Y 0.32fF
C42615 AND2X1_LOC_76/Y AND2X1_LOC_203/a_8_24# 0.01fF
C57466 AND2X1_LOC_76/Y VSS 0.25fF
C3259 AND2X1_LOC_710/Y VDD 0.11fF
C3821 AND2X1_LOC_710/Y AND2X1_LOC_347/a_8_24# 0.05fF
C15960 AND2X1_LOC_710/Y AND2X1_LOC_711/a_8_24# 0.01fF
C20762 AND2X1_LOC_710/a_8_24# AND2X1_LOC_710/Y 0.01fF
C22137 AND2X1_LOC_710/Y AND2X1_LOC_711/Y 0.01fF
C35390 AND2X1_LOC_710/Y AND2X1_LOC_347/B 0.03fF
C58016 AND2X1_LOC_710/Y VSS 0.11fF
C10372 VDD AND2X1_LOC_792/B 0.01fF
C15050 AND2X1_LOC_191/B AND2X1_LOC_792/B 0.18fF
C19197 AND2X1_LOC_791/a_8_24# AND2X1_LOC_792/B 0.01fF
C27531 AND2X1_LOC_792/Y AND2X1_LOC_792/B 0.83fF
C29120 AND2X1_LOC_711/Y AND2X1_LOC_792/B 0.01fF
C46901 AND2X1_LOC_792/B AND2X1_LOC_792/a_8_24# 0.01fF
C56443 AND2X1_LOC_792/B VSS 0.10fF
C24485 AND2X1_LOC_558/a_8_24# AND2X1_LOC_561/B 0.01fF
C39610 AND2X1_LOC_571/B AND2X1_LOC_561/B 0.01fF
C40921 VDD AND2X1_LOC_561/B 0.02fF
C57686 AND2X1_LOC_561/B VSS 0.08fF
C38582 AND2X1_LOC_231/Y AND2X1_LOC_641/a_8_24# 0.11fF
C6412 AND2X1_LOC_554/B AND2X1_LOC_141/B 0.02fF
C23110 AND2X1_LOC_140/a_8_24# AND2X1_LOC_141/B -0.06fF
C43186 AND2X1_LOC_141/B AND2X1_LOC_772/Y 1.03fF
C12404 VDD OR2X1_LOC_84/Y 0.12fF
C34377 OR2X1_LOC_84/Y OR2X1_LOC_786/a_8_216# 0.07fF
C40487 OR2X1_LOC_244/A OR2X1_LOC_84/Y 0.05fF
C57013 OR2X1_LOC_84/Y VSS 0.20fF
C4162 OR2X1_LOC_653/Y OR2X1_LOC_61/Y 0.01fF
C6964 OR2X1_LOC_61/Y OR2X1_LOC_539/B 0.02fF
C15731 OR2X1_LOC_61/Y OR2X1_LOC_206/A 0.11fF
C17619 OR2X1_LOC_61/Y OR2X1_LOC_392/B 0.10fF
C19871 VDD OR2X1_LOC_61/Y 0.23fF
C24726 OR2X1_LOC_476/B OR2X1_LOC_61/Y 0.10fF
C25582 OR2X1_LOC_201/a_8_216# OR2X1_LOC_61/Y 0.05fF
C35908 OR2X1_LOC_339/a_8_216# OR2X1_LOC_61/Y 0.05fF
C46328 OR2X1_LOC_61/Y OR2X1_LOC_805/A 0.07fF
C47442 OR2X1_LOC_61/Y OR2X1_LOC_228/Y 0.07fF
C54886 OR2X1_LOC_475/Y OR2X1_LOC_61/Y 0.02fF
C57075 OR2X1_LOC_61/Y VSS 0.30fF
C57907 OR2X1_LOC_842/A VSS 0.11fF
C53840 OR2X1_LOC_347/A OR2X1_LOC_347/a_8_216# 0.39fF
C58111 OR2X1_LOC_347/A VSS 0.02fF
C49321 OR2X1_LOC_456/A OR2X1_LOC_563/A 0.04fF
C34235 OR2X1_LOC_652/a_8_216# OR2X1_LOC_468/A 0.18fF
C47889 OR2X1_LOC_468/A OR2X1_LOC_388/a_36_216# -0.00fF
C12584 OR2X1_LOC_770/Y OR2X1_LOC_771/a_8_216# 0.39fF
C26819 VDD OR2X1_LOC_770/Y -0.00fF
C56945 OR2X1_LOC_770/Y VSS 0.18fF
C10630 OR2X1_LOC_228/Y OR2X1_LOC_539/B 0.02fF
C11726 OR2X1_LOC_643/a_8_216# OR2X1_LOC_539/B 0.02fF
C17240 OR2X1_LOC_643/a_36_216# OR2X1_LOC_539/B 0.03fF
C23618 OR2X1_LOC_653/Y OR2X1_LOC_539/B 0.02fF
C44023 OR2X1_LOC_476/B OR2X1_LOC_539/B 0.02fF
C15856 OR2X1_LOC_721/Y OR2X1_LOC_140/Y 0.34fF
C26400 OR2X1_LOC_392/B OR2X1_LOC_140/Y 0.03fF
C150 OR2X1_LOC_193/Y OR2X1_LOC_193/a_8_216# 0.01fF
C27798 OR2X1_LOC_561/a_8_216# OR2X1_LOC_561/A 0.39fF
C43490 OR2X1_LOC_812/B OR2X1_LOC_561/A 0.01fF
C45833 OR2X1_LOC_493/Y OR2X1_LOC_561/A 0.10fF
C56307 OR2X1_LOC_561/A VSS 0.18fF
C19786 OR2X1_LOC_788/a_8_216# OR2X1_LOC_605/Y 0.01fF
C23235 OR2X1_LOC_653/Y OR2X1_LOC_390/a_8_216# 0.02fF
C34152 OR2X1_LOC_653/Y OR2X1_LOC_392/B 0.02fF
C41178 OR2X1_LOC_653/Y OR2X1_LOC_476/B 0.04fF
C47746 OR2X1_LOC_653/Y OR2X1_LOC_653/a_8_216# 0.02fF
C49351 OR2X1_LOC_653/Y OR2X1_LOC_61/a_8_216# 0.03fF
C12566 VDD OR2X1_LOC_190/Y 0.07fF
C32949 OR2X1_LOC_540/a_8_216# OR2X1_LOC_190/Y 0.40fF
C39808 OR2X1_LOC_564/A OR2X1_LOC_190/Y 0.02fF
C56535 OR2X1_LOC_190/Y VSS 0.43fF
C22608 OR2X1_LOC_456/Y OR2X1_LOC_465/a_8_216# 0.18fF
C31726 VDD OR2X1_LOC_456/Y 0.10fF
C45910 OR2X1_LOC_456/Y OR2X1_LOC_456/a_8_216# 0.01fF
C57381 OR2X1_LOC_456/Y VSS 0.09fF
C7024 OR2X1_LOC_850/B OR2X1_LOC_349/A 0.03fF
C12716 OR2X1_LOC_850/B OR2X1_LOC_805/A 0.23fF
C21996 OR2X1_LOC_348/Y OR2X1_LOC_850/B 0.02fF
C22005 OR2X1_LOC_349/a_8_216# OR2X1_LOC_850/B 0.01fF
C24154 OR2X1_LOC_850/a_8_216# OR2X1_LOC_850/B 0.05fF
C38343 OR2X1_LOC_850/B OR2X1_LOC_362/a_8_216# 0.01fF
C42294 OR2X1_LOC_850/B VDD 0.06fF
C44039 OR2X1_LOC_359/A OR2X1_LOC_850/B 0.03fF
C44974 OR2X1_LOC_850/B OR2X1_LOC_362/B 0.02fF
C49650 OR2X1_LOC_850/B OR2X1_LOC_366/B 0.01fF
C57861 OR2X1_LOC_850/B VSS 0.18fF
C2641 OR2X1_LOC_137/Y OR2X1_LOC_204/Y 0.02fF
C21217 VDD OR2X1_LOC_137/Y 0.06fF
C51992 OR2X1_LOC_137/Y OR2X1_LOC_139/a_8_216# 0.18fF
C57786 OR2X1_LOC_137/Y VSS 0.18fF
C4847 OR2X1_LOC_574/a_8_216# OR2X1_LOC_140/B 0.01fF
C5601 OR2X1_LOC_140/B OR2X1_LOC_554/a_8_216# 0.03fF
C6140 OR2X1_LOC_500/A OR2X1_LOC_140/B 0.01fF
C15912 OR2X1_LOC_575/A OR2X1_LOC_140/B 0.03fF
C16682 OR2X1_LOC_140/B OR2X1_LOC_554/a_36_216# 0.02fF
C18024 OR2X1_LOC_632/a_8_216# OR2X1_LOC_140/B 0.01fF
C22284 OR2X1_LOC_140/B OR2X1_LOC_563/A 0.01fF
C22807 OR2X1_LOC_632/Y OR2X1_LOC_140/B 0.09fF
C40682 OR2X1_LOC_140/B OR2X1_LOC_493/Y 0.03fF
C42901 OR2X1_LOC_140/B OR2X1_LOC_560/A 0.02fF
C48740 VDD OR2X1_LOC_140/B 0.19fF
C48991 OR2X1_LOC_140/B OR2X1_LOC_140/a_8_216# 0.03fF
C51326 OR2X1_LOC_499/a_8_216# OR2X1_LOC_140/B 0.01fF
C54463 OR2X1_LOC_140/B OR2X1_LOC_140/a_36_216# 0.02fF
C56490 OR2X1_LOC_140/B VSS -0.01fF
C3774 OR2X1_LOC_734/a_8_216# OR2X1_LOC_737/A 0.03fF
C8685 OR2X1_LOC_737/A OR2X1_LOC_717/a_8_216# 0.03fF
C47985 OR2X1_LOC_833/Y OR2X1_LOC_737/A 0.02fF
C53521 OR2X1_LOC_493/a_8_216# OR2X1_LOC_737/A 0.01fF
C53773 OR2X1_LOC_737/A OR2X1_LOC_493/Y 0.04fF
C18305 OR2X1_LOC_475/Y OR2X1_LOC_721/Y 0.09fF
C28749 OR2X1_LOC_475/Y OR2X1_LOC_392/B 0.08fF
C29310 OR2X1_LOC_475/Y OR2X1_LOC_734/a_8_216# 0.41fF
C3812 OR2X1_LOC_467/A OR2X1_LOC_453/Y 0.01fF
C18785 OR2X1_LOC_453/a_8_216# OR2X1_LOC_453/Y 0.01fF
C505 OR2X1_LOC_337/a_36_216# OR2X1_LOC_365/B 0.02fF
C22195 OR2X1_LOC_336/a_8_216# OR2X1_LOC_365/B 0.14fF
C32208 OR2X1_LOC_703/a_8_216# OR2X1_LOC_365/B 0.39fF
C52354 OR2X1_LOC_170/a_8_216# OR2X1_LOC_365/B 0.01fF
C8656 AND2X1_LOC_84/Y AND2X1_LOC_204/a_8_24# 0.01fF
C10815 AND2X1_LOC_84/Y VDD 0.01fF
C22338 AND2X1_LOC_84/Y AND2X1_LOC_61/Y 0.09fF
C22424 AND2X1_LOC_84/Y AND2X1_LOC_852/Y 0.03fF
C23737 AND2X1_LOC_84/Y AND2X1_LOC_201/a_8_24# 0.01fF
C27876 AND2X1_LOC_84/Y AND2X1_LOC_84/a_8_24# 0.01fF
C35740 AND2X1_LOC_84/Y AND2X1_LOC_201/Y 0.01fF
C58080 AND2X1_LOC_84/Y VSS 0.07fF
C7199 AND2X1_LOC_851/B AND2X1_LOC_455/B 0.05fF
C11624 AND2X1_LOC_455/a_8_24# AND2X1_LOC_455/B -0.01fF
C27371 VDD AND2X1_LOC_455/B 0.03fF
C31743 AND2X1_LOC_523/Y AND2X1_LOC_455/B 0.01fF
C53357 AND2X1_LOC_445/a_8_24# AND2X1_LOC_455/B 0.01fF
C56679 AND2X1_LOC_455/B VSS 0.08fF
C42981 AND2X1_LOC_476/A AND2X1_LOC_649/B 0.02fF
C53874 AND2X1_LOC_773/Y AND2X1_LOC_649/B 0.10fF
C2165 AND2X1_LOC_34/Y AND2X1_LOC_472/B 0.14fF
C6749 AND2X1_LOC_34/Y AND2X1_LOC_35/a_8_24# 0.06fF
C26650 VDD AND2X1_LOC_34/Y 0.24fF
C46935 AND2X1_LOC_34/Y AND2X1_LOC_472/a_8_24# 0.17fF
C52469 AND2X1_LOC_34/Y AND2X1_LOC_476/A 0.19fF
C57294 AND2X1_LOC_34/Y VSS 0.27fF
C4604 AND2X1_LOC_566/B AND2X1_LOC_537/Y 0.16fF
C21334 AND2X1_LOC_537/Y AND2X1_LOC_303/a_8_24# 0.17fF
C22540 AND2X1_LOC_537/Y AND2X1_LOC_774/A 0.17fF
C35271 AND2X1_LOC_211/B AND2X1_LOC_537/Y 0.02fF
C201 AND2X1_LOC_486/Y AND2X1_LOC_721/Y 0.03fF
C723 AND2X1_LOC_486/Y AND2X1_LOC_850/A 0.23fF
C8026 AND2X1_LOC_486/Y AND2X1_LOC_787/a_8_24# 0.05fF
C8631 AND2X1_LOC_486/Y AND2X1_LOC_675/A 0.07fF
C13217 AND2X1_LOC_486/Y AND2X1_LOC_493/a_8_24# 0.08fF
C19810 AND2X1_LOC_486/Y AND2X1_LOC_242/B 0.03fF
C24172 AND2X1_LOC_486/Y AND2X1_LOC_456/B 0.03fF
C25825 AND2X1_LOC_486/Y AND2X1_LOC_833/a_8_24# 0.06fF
C30088 AND2X1_LOC_486/Y AND2X1_LOC_850/a_8_24# 0.13fF
C31338 AND2X1_LOC_486/Y AND2X1_LOC_840/A 0.03fF
C13194 AND2X1_LOC_842/B AND2X1_LOC_500/B 0.53fF
C20658 VDD AND2X1_LOC_500/B 0.17fF
C47974 AND2X1_LOC_675/Y AND2X1_LOC_500/B 0.82fF
C56731 AND2X1_LOC_500/B VSS 0.19fF
C4164 AND2X1_LOC_833/a_8_24# AND2X1_LOC_840/A 0.01fF
C30864 VDD AND2X1_LOC_840/A 0.11fF
C57090 AND2X1_LOC_840/A VSS 0.21fF
C16838 VDD AND2X1_LOC_401/Y 0.38fF
C56635 AND2X1_LOC_401/Y VSS 0.15fF
C1849 AND2X1_LOC_849/A AND2X1_LOC_845/Y 0.02fF
C3864 AND2X1_LOC_474/A AND2X1_LOC_849/A 0.02fF
C16997 VDD AND2X1_LOC_849/A 0.38fF
C20764 AND2X1_LOC_721/Y AND2X1_LOC_849/A 1.01fF
C25172 AND2X1_LOC_849/A AND2X1_LOC_806/A 0.02fF
C37212 AND2X1_LOC_849/A AND2X1_LOC_244/A 0.28fF
C53621 AND2X1_LOC_849/A AND2X1_LOC_243/Y 0.09fF
C57093 AND2X1_LOC_849/A VSS 0.19fF
C2852 AND2X1_LOC_574/a_8_24# AND2X1_LOC_500/Y 0.01fF
C6560 AND2X1_LOC_501/Y AND2X1_LOC_500/Y 0.01fF
C11228 AND2X1_LOC_574/Y AND2X1_LOC_500/Y 0.24fF
C11875 AND2X1_LOC_711/Y AND2X1_LOC_500/Y 0.08fF
C12145 AND2X1_LOC_658/B AND2X1_LOC_500/Y 0.03fF
C20264 AND2X1_LOC_675/Y AND2X1_LOC_500/Y 0.02fF
C42253 AND2X1_LOC_500/Y AND2X1_LOC_658/A 0.03fF
C49214 VDD AND2X1_LOC_500/Y 0.07fF
C51772 AND2X1_LOC_500/Y AND2X1_LOC_501/a_8_24# 0.01fF
C57818 AND2X1_LOC_500/Y VSS 0.09fF
C929 AND2X1_LOC_191/B AND2X1_LOC_624/B 0.03fF
C13457 AND2X1_LOC_624/B AND2X1_LOC_792/Y 0.02fF
C15061 AND2X1_LOC_711/Y AND2X1_LOC_624/B 0.03fF
C18471 AND2X1_LOC_624/B AND2X1_LOC_624/a_36_24# 0.01fF
C23940 AND2X1_LOC_456/B AND2X1_LOC_624/B 0.01fF
C24490 AND2X1_LOC_624/B AND2X1_LOC_793/Y 0.02fF
C35863 AND2X1_LOC_620/Y AND2X1_LOC_624/B 0.05fF
C52429 VDD AND2X1_LOC_624/B 0.46fF
C52541 AND2X1_LOC_624/B AND2X1_LOC_624/a_8_24# 0.03fF
C56864 AND2X1_LOC_624/B VSS 0.24fF
C1279 AND2X1_LOC_33/Y AND2X1_LOC_35/a_8_24# 0.18fF
C21182 VDD AND2X1_LOC_33/Y 0.21fF
C57295 AND2X1_LOC_33/Y VSS 0.06fF
C7471 VDD AND2X1_LOC_61/Y 0.15fF
C11855 AND2X1_LOC_61/Y AND2X1_LOC_339/a_8_24# -0.00fF
C12452 AND2X1_LOC_61/Y AND2X1_LOC_203/a_8_24# 0.01fF
C19070 AND2X1_LOC_61/Y AND2X1_LOC_852/Y 0.06fF
C32384 AND2X1_LOC_61/Y AND2X1_LOC_201/Y 0.22fF
C33116 AND2X1_LOC_61/Y AND2X1_LOC_476/A 0.02fF
C53219 AND2X1_LOC_61/Y AND2X1_LOC_640/a_8_24# 0.02fF
C57716 AND2X1_LOC_61/Y VSS -0.47fF
C4131 AND2X1_LOC_721/Y AND2X1_LOC_523/Y 0.37fF
C10341 AND2X1_LOC_523/Y AND2X1_LOC_844/a_8_24# 0.09fF
C26249 AND2X1_LOC_523/Y AND2X1_LOC_445/a_8_24# 0.01fF
C40581 AND2X1_LOC_523/Y AND2X1_LOC_455/a_8_24# -0.00fF
C45947 AND2X1_LOC_553/A AND2X1_LOC_523/Y 0.14fF
C23759 AND2X1_LOC_565/B AND2X1_LOC_565/Y 0.21fF
C35519 AND2X1_LOC_565/a_8_24# AND2X1_LOC_565/Y 0.01fF
C46436 AND2X1_LOC_191/Y AND2X1_LOC_565/Y 0.07fF
C46454 AND2X1_LOC_711/Y AND2X1_LOC_565/Y 0.03fF
C14182 OR2X1_LOC_726/A OR2X1_LOC_550/B 0.11fF
C24394 OR2X1_LOC_726/A OR2X1_LOC_727/a_8_216# 0.39fF
C37918 VDD OR2X1_LOC_726/A 0.06fF
C40673 OR2X1_LOC_471/Y OR2X1_LOC_726/A 0.99fF
C46537 OR2X1_LOC_726/A OR2X1_LOC_731/A 0.09fF
C55448 OR2X1_LOC_726/A OR2X1_LOC_726/a_8_216# 0.02fF
C56619 OR2X1_LOC_726/A VSS 0.26fF
C46297 OR2X1_LOC_705/Y OR2X1_LOC_725/A 0.02fF
C788 AND2X1_LOC_337/B AND2X1_LOC_352/B 0.15fF
C21538 AND2X1_LOC_392/A AND2X1_LOC_352/B 0.05fF
C49221 AND2X1_LOC_337/a_8_24# AND2X1_LOC_352/B 0.01fF
C10513 AND2X1_LOC_456/Y AND2X1_LOC_242/B 0.02fF
C30014 AND2X1_LOC_456/Y AND2X1_LOC_456/a_8_24# 0.01fF
C43252 VDD AND2X1_LOC_456/Y 0.27fF
C45564 AND2X1_LOC_456/Y AND2X1_LOC_465/a_8_24# 0.06fF
C56791 AND2X1_LOC_456/Y VSS 0.37fF
C241 VDD AND2X1_LOC_850/A 0.17fF
C7511 AND2X1_LOC_509/a_8_24# AND2X1_LOC_850/A 0.03fF
C8529 AND2X1_LOC_850/A AND2X1_LOC_806/A 0.03fF
C20654 AND2X1_LOC_850/A AND2X1_LOC_244/A 1.35fF
C23633 AND2X1_LOC_850/A AND2X1_LOC_242/B 0.01fF
C24530 AND2X1_LOC_509/Y AND2X1_LOC_850/A 0.08fF
C43184 AND2X1_LOC_474/A AND2X1_LOC_850/A 0.03fF
C49004 AND2X1_LOC_842/B AND2X1_LOC_850/A 0.01fF
C57179 AND2X1_LOC_850/A VSS -0.13fF
C28253 VDD AND2X1_LOC_347/B 0.01fF
C28795 AND2X1_LOC_347/B AND2X1_LOC_347/a_8_24# 0.04fF
C39807 AND2X1_LOC_347/B AND2X1_LOC_347/a_36_24# 0.01fF
C40912 AND2X1_LOC_711/a_8_24# AND2X1_LOC_347/B 0.05fF
C47224 AND2X1_LOC_711/Y AND2X1_LOC_347/B 0.01fF
C57547 AND2X1_LOC_347/B VSS 0.24fF
C1457 AND2X1_LOC_211/B AND2X1_LOC_641/a_8_24# 0.01fF
C11017 AND2X1_LOC_211/B AND2X1_LOC_303/a_8_24# 0.01fF
C19012 AND2X1_LOC_773/Y AND2X1_LOC_211/B 0.10fF
C19646 AND2X1_LOC_175/a_8_24# AND2X1_LOC_211/B 0.01fF
C20447 AND2X1_LOC_175/B AND2X1_LOC_211/B 0.36fF
C32753 AND2X1_LOC_211/B AND2X1_LOC_326/A 0.02fF
C34698 AND2X1_LOC_392/A AND2X1_LOC_211/B 0.10fF
C38255 AND2X1_LOC_211/B AND2X1_LOC_326/a_8_24# 0.03fF
C39067 AND2X1_LOC_716/a_8_24# AND2X1_LOC_211/B 0.01fF
C44233 AND2X1_LOC_211/B AND2X1_LOC_354/B 0.03fF
C43761 AND2X1_LOC_784/Y AND2X1_LOC_675/A 0.01fF
C3978 AND2X1_LOC_640/Y AND2X1_LOC_640/a_36_24# 0.01fF
C23561 AND2X1_LOC_640/Y AND2X1_LOC_476/A 0.21fF
C43422 AND2X1_LOC_640/Y AND2X1_LOC_640/a_8_24# 0.01fF
C367 OR2X1_LOC_849/A OR2X1_LOC_624/Y 0.01fF
C11069 OR2X1_LOC_849/a_8_216# OR2X1_LOC_624/Y 0.01fF
C14752 OR2X1_LOC_624/a_8_216# OR2X1_LOC_624/Y 0.01fF
C25773 OR2X1_LOC_624/a_36_216# OR2X1_LOC_624/Y 0.01fF
C27615 OR2X1_LOC_474/a_8_216# OR2X1_LOC_624/Y 0.01fF
C48370 OR2X1_LOC_624/Y OR2X1_LOC_392/B 0.05fF
C65 AND2X1_LOC_124/a_8_24# AND2X1_LOC_845/Y 0.03fF
C1252 AND2X1_LOC_845/Y AND2X1_LOC_244/A 0.03fF
C1820 AND2X1_LOC_123/a_8_24# AND2X1_LOC_845/Y 0.02fF
C17408 AND2X1_LOC_845/Y AND2X1_LOC_243/Y 1.38fF
C23889 AND2X1_LOC_474/A AND2X1_LOC_845/Y 0.07fF
C25490 AND2X1_LOC_719/Y AND2X1_LOC_845/Y 0.50fF
C27639 AND2X1_LOC_362/a_8_24# AND2X1_LOC_845/Y -0.00fF
C31115 AND2X1_LOC_554/B AND2X1_LOC_845/Y 0.02fF
C32831 AND2X1_LOC_845/Y AND2X1_LOC_849/a_8_24# 0.07fF
C33075 AND2X1_LOC_392/A AND2X1_LOC_845/Y 0.07fF
C33117 AND2X1_LOC_366/A AND2X1_LOC_845/Y 0.03fF
C36860 VDD AND2X1_LOC_845/Y 0.68fF
C40639 AND2X1_LOC_721/Y AND2X1_LOC_845/Y 0.02fF
C41608 AND2X1_LOC_191/B AND2X1_LOC_845/Y 0.65fF
C45171 AND2X1_LOC_845/Y AND2X1_LOC_806/A 0.15fF
C50789 AND2X1_LOC_123/Y AND2X1_LOC_845/Y 0.01fF
C56828 AND2X1_LOC_845/Y VSS -4.38fF
C3777 AND2X1_LOC_721/Y AND2X1_LOC_471/a_8_24# 0.01fF
C7956 AND2X1_LOC_721/Y AND2X1_LOC_806/A 0.02fF
C9105 AND2X1_LOC_721/Y AND2X1_LOC_734/a_8_24# 0.09fF
C9728 AND2X1_LOC_721/Y AND2X1_LOC_844/a_8_24# 0.17fF
C10010 AND2X1_LOC_721/Y AND2X1_LOC_734/Y 0.01fF
C11873 AND2X1_LOC_721/Y AND2X1_LOC_675/A 0.02fF
C18902 AND2X1_LOC_721/Y AND2X1_LOC_658/B 0.03fF
C24410 AND2X1_LOC_721/Y AND2X1_LOC_785/Y 0.01fF
C27392 AND2X1_LOC_721/Y AND2X1_LOC_456/B 0.01fF
C29868 AND2X1_LOC_721/Y AND2X1_LOC_786/Y 0.19fF
C34530 AND2X1_LOC_721/Y AND2X1_LOC_471/Y 0.01fF
C35590 AND2X1_LOC_721/Y AND2X1_LOC_851/B 0.02fF
C36205 AND2X1_LOC_721/Y AND2X1_LOC_243/Y 0.02fF
C39968 AND2X1_LOC_564/B AND2X1_LOC_721/Y 0.05fF
C42598 AND2X1_LOC_785/a_8_24# AND2X1_LOC_721/Y 0.01fF
C42676 AND2X1_LOC_721/Y AND2X1_LOC_474/A 0.02fF
C44357 AND2X1_LOC_719/Y AND2X1_LOC_721/Y 0.01fF
C46589 AND2X1_LOC_721/Y AND2X1_LOC_362/a_8_24# 0.05fF
C49167 AND2X1_LOC_721/Y AND2X1_LOC_658/A 0.03fF
C51765 AND2X1_LOC_721/Y AND2X1_LOC_717/a_8_24# 0.05fF
C55943 AND2X1_LOC_721/Y VDD 1.02fF
C57962 AND2X1_LOC_721/Y VSS -2.77fF
C31694 OR2X1_LOC_337/a_8_216# OR2X1_LOC_352/A 0.01fF
C6475 AND2X1_LOC_773/Y AND2X1_LOC_786/Y 0.21fF
C12922 AND2X1_LOC_785/a_8_24# AND2X1_LOC_786/Y 0.02fF
C13458 AND2X1_LOC_642/a_8_24# AND2X1_LOC_786/Y 0.06fF
C19260 AND2X1_LOC_785/A AND2X1_LOC_786/Y 0.01fF
C21974 AND2X1_LOC_717/a_8_24# AND2X1_LOC_786/Y 0.04fF
C22352 AND2X1_LOC_392/A AND2X1_LOC_786/Y 0.07fF
C30092 AND2X1_LOC_471/a_8_24# AND2X1_LOC_786/Y 0.02fF
C49125 AND2X1_LOC_476/a_8_24# AND2X1_LOC_786/Y 0.05fF
C51924 AND2X1_LOC_476/A AND2X1_LOC_786/Y 0.02fF
C33843 AND2X1_LOC_201/a_8_24# AND2X1_LOC_201/Y 0.01fF
C12860 OR2X1_LOC_471/Y OR2X1_LOC_210/a_8_216# 0.14fF
C16004 OR2X1_LOC_471/Y OR2X1_LOC_726/a_8_216# 0.04fF
C19843 OR2X1_LOC_471/Y OR2X1_LOC_546/a_8_216# 0.10fF
C29373 OR2X1_LOC_471/Y OR2X1_LOC_209/a_8_216# 0.04fF
C30839 OR2X1_LOC_471/Y OR2X1_LOC_550/B 6.13fF
C37705 OR2X1_LOC_471/Y OR2X1_LOC_190/a_8_216# 0.40fF
C41529 OR2X1_LOC_148/a_8_216# OR2X1_LOC_471/Y 0.14fF
C43961 OR2X1_LOC_471/Y OR2X1_LOC_545/a_8_216# 0.06fF
C47264 OR2X1_LOC_148/Y OR2X1_LOC_471/Y 0.13fF
C7051 AND2X1_LOC_392/A AND2X1_LOC_716/Y 0.07fF
C10703 AND2X1_LOC_716/Y AND2X1_LOC_326/a_8_24# 0.01fF
C16524 AND2X1_LOC_716/Y AND2X1_LOC_354/B 0.08fF
C21792 AND2X1_LOC_716/Y AND2X1_LOC_326/a_36_24# 0.01fF
C36283 AND2X1_LOC_716/Y AND2X1_LOC_180/a_8_24# 0.03fF
C39325 AND2X1_LOC_716/Y AND2X1_LOC_303/a_8_24# 0.01fF
C47537 AND2X1_LOC_773/Y AND2X1_LOC_716/Y 0.10fF
C47567 AND2X1_LOC_716/Y AND2X1_LOC_180/a_36_24# 0.01fF
C50581 AND2X1_LOC_716/Y AND2X1_LOC_303/a_36_24# 0.01fF
C2083 AND2X1_LOC_566/B AND2X1_LOC_326/A 0.02fF
C4051 AND2X1_LOC_392/A AND2X1_LOC_566/B 0.07fF
C13520 AND2X1_LOC_566/B AND2X1_LOC_354/B 0.04fF
C30750 AND2X1_LOC_566/B AND2X1_LOC_353/a_8_24# 0.10fF
C36263 AND2X1_LOC_566/B AND2X1_LOC_303/a_8_24# 0.01fF
C44364 AND2X1_LOC_773/Y AND2X1_LOC_566/B 0.03fF
C23130 AND2X1_LOC_785/a_8_24# AND2X1_LOC_564/B 0.02fF
C29403 AND2X1_LOC_785/A AND2X1_LOC_564/B 0.01fF
C32015 AND2X1_LOC_564/B AND2X1_LOC_717/a_8_24# 0.02fF
C32380 AND2X1_LOC_565/B AND2X1_LOC_564/B 0.14fF
C40160 AND2X1_LOC_564/B AND2X1_LOC_471/a_8_24# 0.02fF
C45631 AND2X1_LOC_564/B AND2X1_LOC_734/a_8_24# 0.01fF
C55198 AND2X1_LOC_564/B AND2X1_LOC_711/Y 0.13fF
C32231 OR2X1_LOC_725/B OR2X1_LOC_705/Y 0.02fF
C21809 OR2X1_LOC_726/a_8_216# OR2X1_LOC_731/A 0.03fF
C36508 OR2X1_LOC_731/A OR2X1_LOC_550/B 0.03fF
C40983 OR2X1_LOC_797/B OR2X1_LOC_209/a_8_216# 0.08fF
C11802 OR2X1_LOC_795/B OR2X1_LOC_785/B 0.01fF
C43579 OR2X1_LOC_785/a_8_216# OR2X1_LOC_795/B -0.00fF
C5240 OR2X1_LOC_354/A OR2X1_LOC_703/a_8_216# 0.04fF
C12082 OR2X1_LOC_354/A OR2X1_LOC_354/a_8_216# 0.01fF
C18550 OR2X1_LOC_354/A OR2X1_LOC_356/a_8_216# 0.03fF
C33864 OR2X1_LOC_354/A OR2X1_LOC_620/Y 0.01fF
C39715 VDD OR2X1_LOC_354/A 0.12fF
C57798 OR2X1_LOC_354/A VSS 0.19fF
C13497 OR2X1_LOC_717/a_8_216# OR2X1_LOC_723/A -0.00fF
C1825 OR2X1_LOC_472/A OR2X1_LOC_852/A 0.01fF
C2524 VDD OR2X1_LOC_472/A 0.34fF
C7319 OR2X1_LOC_476/B OR2X1_LOC_472/A 0.01fF
C17303 OR2X1_LOC_852/a_8_216# OR2X1_LOC_472/A 0.03fF
C28358 OR2X1_LOC_852/a_36_216# OR2X1_LOC_472/A 0.02fF
C41216 OR2X1_LOC_472/a_8_216# OR2X1_LOC_472/A 0.02fF
C41244 OR2X1_LOC_472/A OR2X1_LOC_839/a_8_216# 0.06fF
C57502 OR2X1_LOC_472/A VSS -1.25fF
C501 OR2X1_LOC_654/A OR2X1_LOC_476/B 0.01fF
C9914 OR2X1_LOC_654/A OR2X1_LOC_35/B 0.03fF
C36797 OR2X1_LOC_654/A OR2X1_LOC_35/a_8_216# 0.02fF
C3169 AND2X1_LOC_555/Y AND2X1_LOC_555/a_8_24# 0.02fF
C28726 AND2X1_LOC_555/Y AND2X1_LOC_345/Y 0.68fF
C34204 AND2X1_LOC_555/Y AND2X1_LOC_348/a_8_24# 0.01fF
C36696 AND2X1_LOC_555/Y AND2X1_LOC_259/Y 0.05fF
C43940 AND2X1_LOC_555/Y AND2X1_LOC_191/B 0.03fF
C53506 AND2X1_LOC_555/Y AND2X1_LOC_345/a_8_24# 0.03fF
C41306 OR2X1_LOC_833/Y OR2X1_LOC_851/B 0.02fF
C47019 OR2X1_LOC_840/a_8_216# OR2X1_LOC_851/B 0.03fF
C19382 AND2X1_LOC_658/B AND2X1_LOC_508/B 0.03fF
C23245 AND2X1_LOC_658/B AND2X1_LOC_565/a_8_24# 0.03fF
C24926 AND2X1_LOC_574/a_8_24# AND2X1_LOC_658/B 0.02fF
C33901 AND2X1_LOC_658/B AND2X1_LOC_191/Y 0.03fF
C33909 AND2X1_LOC_658/B AND2X1_LOC_711/Y 0.03fF
C41454 AND2X1_LOC_658/B AND2X1_LOC_550/A 0.03fF
C50652 AND2X1_LOC_658/B AND2X1_LOC_148/Y 0.05fF
C50947 AND2X1_LOC_658/B AND2X1_LOC_545/a_8_24# 0.03fF
C50999 AND2X1_LOC_728/Y AND2X1_LOC_658/B 0.14fF
C54932 AND2X1_LOC_658/B AND2X1_LOC_620/Y 0.01fF
C39435 AND2X1_LOC_449/Y AND2X1_LOC_453/Y 0.03fF
C40670 AND2X1_LOC_453/Y AND2X1_LOC_452/Y 0.03fF
C45043 AND2X1_LOC_453/a_8_24# AND2X1_LOC_453/Y 0.02fF
C5396 OR2X1_LOC_856/B OR2X1_LOC_620/Y 0.41fF
C11714 OR2X1_LOC_620/Y OR2X1_LOC_703/a_8_216# 0.01fF
C18497 OR2X1_LOC_620/Y OR2X1_LOC_354/a_8_216# 0.01fF
C21111 OR2X1_LOC_620/Y OR2X1_LOC_486/Y 0.03fF
C24948 OR2X1_LOC_620/Y OR2X1_LOC_356/a_8_216# 0.01fF
C44962 OR2X1_LOC_854/a_8_216# OR2X1_LOC_620/Y -0.03fF
C51458 OR2X1_LOC_620/Y OR2X1_LOC_623/a_8_216# 0.01fF
C56063 OR2X1_LOC_326/a_8_216# OR2X1_LOC_620/Y 0.02fF
C57452 OR2X1_LOC_620/Y VSS 0.52fF
C49117 OR2X1_LOC_231/a_8_216# OR2X1_LOC_641/B 0.01fF
C8516 AND2X1_LOC_456/B AND2X1_LOC_348/Y 0.37fF
C58033 OR2X1_LOC_345/Y VSS 0.14fF
C57221 OR2X1_LOC_401/Y VSS 0.19fF
C9498 AND2X1_LOC_679/a_8_24# OR2X1_LOC_715/A 0.02fF
C20537 OR2X1_LOC_728/B OR2X1_LOC_715/A 0.14fF
C34576 VDD OR2X1_LOC_715/A 0.12fF
C56517 OR2X1_LOC_715/A VSS 0.15fF
C45602 OR2X1_LOC_241/a_8_216# OR2X1_LOC_241/Y 0.02fF
C46616 OR2X1_LOC_241/Y OR2X1_LOC_493/Y 0.03fF
C57263 OR2X1_LOC_241/Y VSS 0.15fF
C23775 VDD AND2X1_LOC_856/A 0.21fF
C50788 AND2X1_LOC_856/A AND2X1_LOC_856/a_8_24# 0.19fF
C57127 AND2X1_LOC_856/A VSS 0.06fF
C13510 AND2X1_LOC_170/a_8_24# AND2X1_LOC_568/B 0.02fF
C28656 AND2X1_LOC_392/A AND2X1_LOC_568/B 0.07fF
C43337 AND2X1_LOC_568/B AND2X1_LOC_170/B 0.20fF
C29980 AND2X1_LOC_509/Y AND2X1_LOC_510/A 0.02fF
C40949 AND2X1_LOC_510/a_8_24# AND2X1_LOC_510/A 0.03fF
C57363 AND2X1_LOC_510/A VSS 0.04fF
C7241 AND2X1_LOC_852/a_8_24# AND2X1_LOC_852/Y 0.03fF
C23890 AND2X1_LOC_852/a_36_24# AND2X1_LOC_852/Y 0.01fF
C33217 AND2X1_LOC_476/A AND2X1_LOC_852/Y 0.07fF
C47290 AND2X1_LOC_852/Y AND2X1_LOC_852/B 0.05fF
C25699 AND2X1_LOC_141/A AND2X1_LOC_772/Y 0.01fF
C53274 AND2X1_LOC_139/A AND2X1_LOC_141/A 0.83fF
C7306 AND2X1_LOC_456/B AND2X1_LOC_620/Y 0.39fF
C7915 AND2X1_LOC_620/Y AND2X1_LOC_793/Y 0.07fF
C9974 AND2X1_LOC_632/a_8_24# AND2X1_LOC_620/Y 0.01fF
C24902 AND2X1_LOC_620/Y AND2X1_LOC_623/a_8_24# 0.04fF
C28924 AND2X1_LOC_658/A AND2X1_LOC_620/Y 1.09fF
C35675 VDD AND2X1_LOC_620/Y 0.10fF
C40323 AND2X1_LOC_191/B AND2X1_LOC_620/Y 0.01fF
C47102 AND2X1_LOC_620/Y AND2X1_LOC_623/a_36_24# 0.01fF
C53039 AND2X1_LOC_620/Y AND2X1_LOC_792/Y 0.07fF
C54626 AND2X1_LOC_711/Y AND2X1_LOC_620/Y 0.01fF
C56865 AND2X1_LOC_620/Y VSS -0.16fF
C43324 AND2X1_LOC_202/a_8_24# AND2X1_LOC_202/Y 0.01fF
C23794 AND2X1_LOC_392/A AND2X1_LOC_337/B 0.01fF
C25142 AND2X1_LOC_337/B AND2X1_LOC_661/A 0.14fF
C27529 VDD AND2X1_LOC_337/B 0.39fF
C51461 AND2X1_LOC_337/B AND2X1_LOC_337/a_8_24# 0.01fF
C51548 AND2X1_LOC_365/A AND2X1_LOC_337/B 0.03fF
C57474 AND2X1_LOC_337/B VSS 0.27fF
C1490 AND2X1_LOC_719/Y AND2X1_LOC_552/A 0.03fF
C7428 AND2X1_LOC_552/A AND2X1_LOC_476/Y 0.04fF
C12999 AND2X1_LOC_552/A VDD 0.25fF
C47880 AND2X1_LOC_552/a_8_24# AND2X1_LOC_552/A 0.19fF
C57953 AND2X1_LOC_552/A VSS 0.10fF
C57458 OR2X1_LOC_647/Y VSS 0.16fF
C13748 AND2X1_LOC_785/A AND2X1_LOC_785/Y 0.51fF
C31903 AND2X1_LOC_785/a_8_24# AND2X1_LOC_785/A 0.01fF
C39591 AND2X1_LOC_785/A AND2X1_LOC_476/Y 0.04fF
C58088 AND2X1_LOC_785/A VSS 0.04fF
C4401 AND2X1_LOC_771/B AND2X1_LOC_774/A -0.00fF
C30756 VDD AND2X1_LOC_771/B 0.14fF
C55045 AND2X1_LOC_771/B AND2X1_LOC_771/a_8_24# 0.11fF
C56392 AND2X1_LOC_771/B VSS 0.19fF
C8876 AND2X1_LOC_842/B AND2X1_LOC_244/A 0.01fF
C12166 AND2X1_LOC_474/a_8_24# AND2X1_LOC_244/A 0.10fF
C12310 AND2X1_LOC_849/a_8_24# AND2X1_LOC_244/A 0.01fF
C18994 AND2X1_LOC_244/A AND2X1_LOC_288/a_8_24# 0.01fF
C21045 AND2X1_LOC_191/B AND2X1_LOC_244/A 0.03fF
C39592 AND2X1_LOC_242/B AND2X1_LOC_244/A 0.01fF
C40486 AND2X1_LOC_509/Y AND2X1_LOC_244/A 0.03fF
C43973 AND2X1_LOC_456/B AND2X1_LOC_244/A 0.02fF
C50087 AND2X1_LOC_850/a_8_24# AND2X1_LOC_244/A 0.01fF
C5921 AND2X1_LOC_850/Y AND2X1_LOC_288/a_8_24# 0.20fF
C36808 AND2X1_LOC_850/a_8_24# AND2X1_LOC_850/Y -0.05fF
C48132 AND2X1_LOC_850/a_36_24# AND2X1_LOC_850/Y 0.01fF
C48553 OR2X1_LOC_602/Y OR2X1_LOC_602/a_8_216# 0.01fF
C29074 OR2X1_LOC_720/Y OR2X1_LOC_721/Y -0.01fF
C43610 OR2X1_LOC_720/a_8_216# OR2X1_LOC_720/Y -0.00fF
C48324 OR2X1_LOC_720/Y OR2X1_LOC_721/a_8_216# 0.39fF
C56671 OR2X1_LOC_720/Y VSS 0.10fF
C2783 OR2X1_LOC_209/a_8_216# OR2X1_LOC_550/B 0.40fF
C3257 OR2X1_LOC_486/a_8_216# OR2X1_LOC_550/B 0.06fF
C7323 OR2X1_LOC_620/a_8_216# OR2X1_LOC_550/B 0.06fF
C28169 VDD OR2X1_LOC_550/B 0.09fF
C33649 OR2X1_LOC_550/a_8_216# OR2X1_LOC_550/B 0.08fF
C50460 OR2X1_LOC_739/A OR2X1_LOC_550/B 0.03fF
C53402 OR2X1_LOC_213/A OR2X1_LOC_550/B 0.04fF
C56359 OR2X1_LOC_550/B VSS 0.40fF
C729 OR2X1_LOC_508/A OR2X1_LOC_721/Y 0.45fF
C11269 OR2X1_LOC_508/A OR2X1_LOC_392/B 0.10fF
C23307 OR2X1_LOC_508/A OR2X1_LOC_244/B 0.13fF
C44415 OR2X1_LOC_508/A OR2X1_LOC_508/a_8_216# -0.04fF
C47025 OR2X1_LOC_508/A OR2X1_LOC_508/Y 0.01fF
C58041 OR2X1_LOC_508/A VSS 0.01fF
C7541 OR2X1_LOC_859/a_8_216# OR2X1_LOC_862/A 0.04fF
C16930 OR2X1_LOC_810/a_8_216# OR2X1_LOC_862/A 0.41fF
C20737 AND2X1_LOC_403/B AND2X1_LOC_403/a_8_24# 0.04fF
C54762 VDD AND2X1_LOC_403/B 0.04fF
C56744 AND2X1_LOC_403/B VSS 0.02fF
C2069 AND2X1_LOC_474/A AND2X1_LOC_124/a_8_24# 0.01fF
C7060 AND2X1_LOC_509/Y AND2X1_LOC_474/A 0.15fF
C10515 AND2X1_LOC_456/B AND2X1_LOC_474/A 0.02fF
C16457 AND2X1_LOC_474/A AND2X1_LOC_850/a_8_24# 0.01fF
C29571 AND2X1_LOC_362/a_8_24# AND2X1_LOC_474/A 0.01fF
C33056 AND2X1_LOC_554/B AND2X1_LOC_474/A 0.23fF
C34685 AND2X1_LOC_474/A AND2X1_LOC_474/a_8_24# -0.00fF
C34841 AND2X1_LOC_474/A AND2X1_LOC_849/a_8_24# 0.01fF
C41521 AND2X1_LOC_474/A AND2X1_LOC_288/a_8_24# 0.01fF
C43591 AND2X1_LOC_191/B AND2X1_LOC_474/A 0.03fF
C52711 AND2X1_LOC_474/A AND2X1_LOC_123/Y 0.14fF
C17913 AND2X1_LOC_191/B AND2X1_LOC_792/Y 0.01fF
C31952 AND2X1_LOC_711/Y AND2X1_LOC_792/Y 0.01fF
C33468 AND2X1_LOC_792/Y AND2X1_LOC_793/a_8_24# 0.04fF
C17595 OR2X1_LOC_35/A OR2X1_LOC_35/a_8_216# 0.39fF
C46749 OR2X1_LOC_35/B OR2X1_LOC_35/A 0.06fF
C56752 OR2X1_LOC_35/A VSS 0.18fF
C47805 AND2X1_LOC_139/A AND2X1_LOC_139/a_8_24# 0.01fF
C51284 AND2X1_LOC_137/a_8_24# AND2X1_LOC_139/A 0.01fF
C54486 VDD AND2X1_LOC_139/A -0.00fF
C57226 AND2X1_LOC_139/A VSS -0.23fF
C12143 AND2X1_LOC_772/B VDD 0.04fF
C21911 AND2X1_LOC_772/B AND2X1_LOC_554/a_8_24# 0.03fF
C38052 AND2X1_LOC_772/B AND2X1_LOC_560/B 0.01fF
C57922 AND2X1_LOC_772/B VSS 0.35fF
C10456 AND2X1_LOC_456/B AND2X1_LOC_456/a_8_24# 0.11fF
C11450 AND2X1_LOC_456/B AND2X1_LOC_359/B 0.02fF
C16493 AND2X1_LOC_456/B AND2X1_LOC_859/a_8_24# 0.01fF
C16842 AND2X1_LOC_456/B AND2X1_LOC_658/A 0.03fF
C19879 AND2X1_LOC_366/A AND2X1_LOC_456/B 0.03fF
C22987 AND2X1_LOC_456/B AND2X1_LOC_859/Y 0.10fF
C26287 AND2X1_LOC_456/B AND2X1_LOC_288/a_8_24# 0.17fF
C27087 AND2X1_LOC_720/Y AND2X1_LOC_456/B 0.01fF
C28325 AND2X1_LOC_191/B AND2X1_LOC_456/B 0.03fF
C31777 AND2X1_LOC_456/B AND2X1_LOC_806/A 0.06fF
C32553 AND2X1_LOC_721/a_8_24# AND2X1_LOC_456/B 0.01fF
C43223 AND2X1_LOC_720/a_8_24# AND2X1_LOC_456/B 0.01fF
C208 VDD OR2X1_LOC_679/Y -0.00fF
C35935 AND2X1_LOC_728/Y OR2X1_LOC_679/Y 0.21fF
C49664 OR2X1_LOC_679/a_8_216# OR2X1_LOC_679/Y 0.01fF
C57400 OR2X1_LOC_679/Y VSS 0.07fF
C17981 OR2X1_LOC_510/A OR2X1_LOC_508/Y 0.01fF
C29010 OR2X1_LOC_510/A OR2X1_LOC_510/a_8_216# 0.06fF
C34892 OR2X1_LOC_510/A OR2X1_LOC_560/A 0.04fF
C40496 OR2X1_LOC_510/A VDD 0.19fF
C57969 OR2X1_LOC_510/A VSS -0.62fF
C40230 VDD OR2X1_LOC_772/Y 0.10fF
C56841 OR2X1_LOC_772/Y VSS 0.16fF
C6000 OR2X1_LOC_605/a_8_216# OR2X1_LOC_787/Y 0.01fF
C11580 OR2X1_LOC_605/a_36_216# OR2X1_LOC_787/Y 0.01fF
C16746 AND2X1_LOC_574/Y AND2X1_LOC_501/a_8_24# 0.01fF
C24042 AND2X1_LOC_574/a_8_24# AND2X1_LOC_574/Y 0.01fF
C32945 AND2X1_LOC_574/Y AND2X1_LOC_191/Y 0.04fF
C32958 AND2X1_LOC_574/Y AND2X1_LOC_711/Y 0.03fF
C34336 OR2X1_LOC_714/a_8_216# OR2X1_LOC_724/A 0.01fF
C44965 OR2X1_LOC_715/a_8_216# OR2X1_LOC_724/A 0.03fF
C12550 VDD OR2X1_LOC_565/A 0.16fF
C39771 OR2X1_LOC_565/A OR2X1_LOC_564/A 0.68fF
C55157 OR2X1_LOC_565/A OR2X1_LOC_553/B 0.18fF
C56707 OR2X1_LOC_565/A VSS 0.45fF
C3990 OR2X1_LOC_728/B OR2X1_LOC_739/A 0.12fF
C15643 OR2X1_LOC_324/a_8_216# OR2X1_LOC_739/A 0.01fF
C25267 OR2X1_LOC_739/A OR2X1_LOC_728/a_8_216# 0.01fF
C26705 OR2X1_LOC_326/B OR2X1_LOC_739/A 0.03fF
C36215 OR2X1_LOC_739/A OR2X1_LOC_730/B 0.78fF
C49478 OR2X1_LOC_486/a_8_216# OR2X1_LOC_739/A 0.01fF
C2124 AND2X1_LOC_773/Y AND2X1_LOC_476/A 0.10fF
C5458 AND2X1_LOC_340/Y AND2X1_LOC_476/A 0.07fF
C9050 AND2X1_LOC_642/a_8_24# AND2X1_LOC_476/A 0.01fF
C11233 AND2X1_LOC_640/a_8_24# AND2X1_LOC_476/A 0.03fF
C16149 AND2X1_LOC_476/A AND2X1_LOC_476/Y 0.19fF
C17862 AND2X1_LOC_392/A AND2X1_LOC_476/A 0.07fF
C21769 VDD AND2X1_LOC_476/A -0.00fF
C22693 AND2X1_LOC_476/A AND2X1_LOC_642/Y 0.04fF
C25609 AND2X1_LOC_642/a_36_24# AND2X1_LOC_476/A 0.01fF
C26046 AND2X1_LOC_339/a_8_24# AND2X1_LOC_476/A 0.03fF
C27786 AND2X1_LOC_640/a_36_24# AND2X1_LOC_476/A 0.01fF
C33934 AND2X1_LOC_339/Y AND2X1_LOC_476/A 0.04fF
C44584 AND2X1_LOC_476/A AND2X1_LOC_476/a_8_24# 0.11fF
C56990 AND2X1_LOC_476/A VSS 0.79fF
C2769 AND2X1_LOC_243/a_36_24# AND2X1_LOC_243/Y 0.01fF
C23257 AND2X1_LOC_362/a_8_24# AND2X1_LOC_243/Y 0.01fF
C26693 AND2X1_LOC_554/B AND2X1_LOC_243/Y 0.03fF
C28649 AND2X1_LOC_392/A AND2X1_LOC_243/Y 0.07fF
C46234 AND2X1_LOC_123/Y AND2X1_LOC_243/Y 0.04fF
C51829 AND2X1_LOC_124/a_8_24# AND2X1_LOC_243/Y 0.04fF
C53565 AND2X1_LOC_123/a_8_24# AND2X1_LOC_243/Y 0.03fF
C35161 AND2X1_LOC_852/a_8_24# AND2X1_LOC_852/B 0.04fF
C35463 VDD AND2X1_LOC_852/B 0.01fF
C51919 AND2X1_LOC_852/a_36_24# AND2X1_LOC_852/B 0.01fF
C56762 AND2X1_LOC_852/B VSS -0.41fF
C38663 OR2X1_LOC_711/A OR2X1_LOC_705/Y 0.74fF
C39796 VDD OR2X1_LOC_711/A 0.18fF
C56672 OR2X1_LOC_711/A VSS -0.13fF
C47239 OR2X1_LOC_792/Y OR2X1_LOC_288/a_8_216# 0.01fF
C32433 VDD OR2X1_LOC_552/B -0.00fF
C48908 OR2X1_LOC_552/a_8_216# OR2X1_LOC_552/B 0.39fF
C56544 OR2X1_LOC_552/B VSS 0.17fF
C18878 OR2X1_LOC_639/A OR2X1_LOC_639/a_8_216# 0.39fF
C57347 OR2X1_LOC_639/A VSS 0.18fF
C15302 OR2X1_LOC_844/a_8_216# OR2X1_LOC_523/Y 0.01fF
C9214 OR2X1_LOC_651/A OR2X1_LOC_228/Y 0.03fF
C18060 OR2X1_LOC_476/a_8_216# OR2X1_LOC_228/Y 0.01fF
C21344 OR2X1_LOC_392/B OR2X1_LOC_228/Y 0.07fF
C28250 OR2X1_LOC_476/B OR2X1_LOC_228/Y 0.04fF
C28259 OR2X1_LOC_644/a_8_216# OR2X1_LOC_228/Y 0.02fF
C36129 OR2X1_LOC_785/a_8_216# OR2X1_LOC_228/Y 0.01fF
C38711 OR2X1_LOC_841/a_8_216# OR2X1_LOC_228/Y 0.02fF
C38728 OR2X1_LOC_856/B OR2X1_LOC_228/Y 0.07fF
C44690 OR2X1_LOC_644/a_36_216# OR2X1_LOC_228/Y 0.02fF
C52104 OR2X1_LOC_643/a_8_216# OR2X1_LOC_228/Y 0.02fF
C52754 OR2X1_LOC_228/Y OR2X1_LOC_716/a_8_216# 0.05fF
C720 OR2X1_LOC_728/B OR2X1_LOC_715/a_8_216# 0.47fF
C44990 OR2X1_LOC_728/B OR2X1_LOC_728/a_8_216# 0.01fF
C56144 OR2X1_LOC_728/B OR2X1_LOC_730/B 0.01fF
C56808 OR2X1_LOC_728/B VSS 0.26fF
C4710 OR2X1_LOC_455/a_8_216# OR2X1_LOC_455/A 0.39fF
C33866 OR2X1_LOC_455/A OR2X1_LOC_486/Y 0.11fF
C55389 OR2X1_LOC_76/Y OR2X1_LOC_455/A 0.12fF
C57267 OR2X1_LOC_455/A VSS -0.05fF
C44566 AND2X1_LOC_793/Y AND2X1_LOC_793/a_8_24# 0.01fF
C12098 OR2X1_LOC_348/a_8_216# OR2X1_LOC_348/Y -0.00fF
C27777 OR2X1_LOC_348/Y OR2X1_LOC_362/a_8_216# 0.01fF
C15697 AND2X1_LOC_449/Y AND2X1_LOC_453/a_36_24# 0.01fF
C22928 VDD AND2X1_LOC_449/Y 0.21fF
C33883 AND2X1_LOC_605/Y AND2X1_LOC_449/Y 0.01fF
C39724 AND2X1_LOC_449/Y AND2X1_LOC_605/a_8_24# 0.01fF
C45045 AND2X1_LOC_449/Y AND2X1_LOC_454/Y 0.20fF
C49755 AND2X1_LOC_449/Y AND2X1_LOC_454/a_8_24# 0.20fF
C51081 AND2X1_LOC_449/Y AND2X1_LOC_452/Y 0.03fF
C55318 AND2X1_LOC_449/Y AND2X1_LOC_453/a_8_24# 0.03fF
C56847 AND2X1_LOC_449/Y VSS 0.12fF
C1898 VDD AND2X1_LOC_639/B 0.06fF
C45804 AND2X1_LOC_639/B AND2X1_LOC_639/a_8_24# 0.03fF
C56746 AND2X1_LOC_639/B VSS 0.31fF
C641 AND2X1_LOC_191/B VDD 0.58fF
C812 AND2X1_LOC_191/B AND2X1_LOC_624/a_8_24# 0.01fF
C2980 AND2X1_LOC_191/B AND2X1_LOC_465/a_8_24# 0.19fF
C8899 AND2X1_LOC_191/B AND2X1_LOC_806/A 0.03fF
C9554 AND2X1_LOC_191/B AND2X1_LOC_791/a_8_24# 0.01fF
C24040 AND2X1_LOC_191/B AND2X1_LOC_242/B 0.29fF
C37027 AND2X1_LOC_191/B AND2X1_LOC_792/a_8_24# 0.05fF
C37224 AND2X1_LOC_191/B AND2X1_LOC_620/a_8_24# 0.01fF
C45278 AND2X1_LOC_719/Y AND2X1_LOC_191/B 0.07fF
C49774 AND2X1_LOC_191/B AND2X1_LOC_859/a_8_24# 0.03fF
C50092 AND2X1_LOC_191/B AND2X1_LOC_658/A 0.01fF
C52827 AND2X1_LOC_191/B AND2X1_LOC_849/a_8_24# 0.04fF
C56110 AND2X1_LOC_191/B AND2X1_LOC_859/Y 0.39fF
C57975 AND2X1_LOC_191/B VSS -0.86fF
C11466 AND2X1_LOC_553/A AND2X1_LOC_560/B 0.02fF
C41418 AND2X1_LOC_553/A VDD 0.17fF
C58036 AND2X1_LOC_553/A VSS 0.28fF
C51476 OR2X1_LOC_35/B OR2X1_LOC_35/a_8_216# 0.05fF
C56813 OR2X1_LOC_35/B VSS 0.11fF
C942 AND2X1_LOC_554/B AND2X1_LOC_140/a_8_24# 0.01fF
C3883 AND2X1_LOC_554/B AND2X1_LOC_123/Y 0.04fF
C11125 AND2X1_LOC_554/B AND2X1_LOC_123/a_8_24# 0.17fF
C15081 AND2X1_LOC_554/B AND2X1_LOC_772/a_8_24# 0.11fF
C21146 AND2X1_LOC_554/B AND2X1_LOC_772/Y 0.01fF
C42404 AND2X1_LOC_392/A AND2X1_LOC_554/B 0.03fF
C46316 VDD AND2X1_LOC_554/B 0.50fF
C47702 AND2X1_LOC_392/a_8_24# AND2X1_LOC_554/B 0.17fF
C56051 AND2X1_LOC_554/a_8_24# AND2X1_LOC_554/B 0.01fF
C57706 AND2X1_LOC_554/B VSS -0.06fF
C1031 AND2X1_LOC_727/a_8_24# AND2X1_LOC_727/B 0.11fF
C9221 AND2X1_LOC_550/A AND2X1_LOC_727/B 0.03fF
C26136 AND2X1_LOC_444/a_8_24# AND2X1_LOC_727/B 0.01fF
C36533 AND2X1_LOC_345/Y AND2X1_LOC_348/a_8_24# 0.03fF
C39090 AND2X1_LOC_259/Y AND2X1_LOC_345/Y 0.13fF
C41527 VDD AND2X1_LOC_345/Y 0.05fF
C57413 AND2X1_LOC_345/Y VSS -0.32fF
C1644 AND2X1_LOC_656/Y AND2X1_LOC_772/Y 0.09fF
C20118 OR2X1_LOC_476/a_8_216# OR2X1_LOC_476/Y -0.00fF
C23310 OR2X1_LOC_476/Y OR2X1_LOC_392/B 0.01fF
C11604 OR2X1_LOC_575/A OR2X1_LOC_493/Y 0.01fF
C16756 OR2X1_LOC_575/A OR2X1_LOC_500/a_8_216# 0.01fF
C32427 OR2X1_LOC_575/A OR2X1_LOC_554/a_8_216# 0.03fF
C33040 OR2X1_LOC_500/A OR2X1_LOC_575/A 0.02fF
C43541 OR2X1_LOC_575/A OR2X1_LOC_554/a_36_216# 0.01fF
C50577 OR2X1_LOC_632/a_36_216# OR2X1_LOC_575/A 0.01fF
C16115 OR2X1_LOC_812/B OR2X1_LOC_561/a_8_216# 0.02fF
C32374 OR2X1_LOC_812/B OR2X1_LOC_558/a_8_216# 0.02fF
C34051 OR2X1_LOC_812/B OR2X1_LOC_493/Y 0.09fF
C31865 OR2X1_LOC_675/a_8_216# OR2X1_LOC_719/Y 0.39fF
C2544 VDD OR2X1_LOC_647/A 0.06fF
C19690 OR2X1_LOC_647/A OR2X1_LOC_647/a_8_216# 0.08fF
C54104 OR2X1_LOC_646/a_8_216# OR2X1_LOC_647/A 0.01fF
C57394 OR2X1_LOC_647/A VSS 0.23fF
C13148 OR2X1_LOC_648/B OR2X1_LOC_208/a_8_216# 0.33fF
C27564 OR2X1_LOC_476/B OR2X1_LOC_648/B 0.02fF
C37976 OR2X1_LOC_856/B OR2X1_LOC_648/B 0.10fF
C4498 OR2X1_LOC_326/B VDD 0.08fF
C58106 OR2X1_LOC_326/B VSS 0.08fF
C6993 OR2X1_LOC_500/A OR2X1_LOC_500/a_8_216# 0.18fF
C9710 VDD OR2X1_LOC_500/A 0.07fF
C39263 OR2X1_LOC_500/A OR2X1_LOC_563/A 0.01fF
C39781 OR2X1_LOC_500/A OR2X1_LOC_632/Y 0.01fF
C57316 OR2X1_LOC_500/A VSS 0.18fF
C8815 OR2X1_LOC_833/Y OR2X1_LOC_805/A 0.02fF
C28151 OR2X1_LOC_833/Y OR2X1_LOC_723/B 0.07fF
C30319 OR2X1_LOC_833/Y OR2X1_LOC_840/a_8_216# 0.10fF
C38330 OR2X1_LOC_833/Y VDD 0.48fF
C41632 OR2X1_LOC_833/Y OR2X1_LOC_717/a_8_216# 0.14fF
C57948 OR2X1_LOC_833/Y VSS 0.15fF
C4801 OR2X1_LOC_781/Y OR2X1_LOC_782/a_8_216# 0.02fF
C23023 VDD OR2X1_LOC_781/Y 0.08fF
C56948 OR2X1_LOC_781/Y VSS 0.12fF
C27063 OR2X1_LOC_443/a_8_216# OR2X1_LOC_181/Y 0.18fF
C27713 OR2X1_LOC_553/B OR2X1_LOC_565/a_8_216# 0.39fF
C35188 OR2X1_LOC_553/B OR2X1_LOC_553/a_8_216# 0.03fF
C46394 OR2X1_LOC_553/B OR2X1_LOC_563/B 0.09fF
C56657 OR2X1_LOC_553/B VSS 0.28fF
C4469 OR2X1_LOC_555/B OR2X1_LOC_555/a_8_216# 0.07fF
C19731 OR2X1_LOC_555/B OR2X1_LOC_345/a_8_216# 0.02fF
C25238 OR2X1_LOC_555/B OR2X1_LOC_345/a_36_216# 0.03fF
C48052 VDD OR2X1_LOC_555/B 0.26fF
C56955 OR2X1_LOC_555/B VSS 0.46fF
C5681 AND2X1_LOC_388/Y AND2X1_LOC_390/a_8_24# 0.01fF
C16777 AND2X1_LOC_388/Y AND2X1_LOC_392/A 0.01fF
C18175 AND2X1_LOC_388/Y AND2X1_LOC_661/A 0.03fF
C20651 AND2X1_LOC_388/Y VDD 0.06fF
C58103 AND2X1_LOC_388/Y VSS -0.09fF
C3595 AND2X1_LOC_703/Y AND2X1_LOC_714/a_8_24# 0.09fF
C46078 AND2X1_LOC_715/Y AND2X1_LOC_703/Y 0.02fF
C50465 AND2X1_LOC_703/Y VDD 0.21fF
C57876 AND2X1_LOC_703/Y VSS 0.08fF
C30998 AND2X1_LOC_593/Y AND2X1_LOC_653/a_8_24# 0.01fF
C31380 AND2X1_LOC_593/Y AND2X1_LOC_652/a_8_24# 0.04fF
C35069 AND2X1_LOC_392/A AND2X1_LOC_593/Y 0.03fF
C36452 AND2X1_LOC_593/Y AND2X1_LOC_661/A 0.01fF
C36539 AND2X1_LOC_593/Y AND2X1_LOC_810/Y 0.08fF
C42453 AND2X1_LOC_593/Y AND2X1_LOC_652/a_36_24# 0.01fF
C50187 AND2X1_LOC_605/Y AND2X1_LOC_593/Y 0.01fF
C28167 AND2X1_LOC_326/A AND2X1_LOC_863/A 0.09fF
C46066 AND2X1_LOC_326/A AND2X1_LOC_326/a_8_24# 0.10fF
C46346 VDD AND2X1_LOC_326/A 0.21fF
C52019 AND2X1_LOC_326/A AND2X1_LOC_354/B 0.06fF
C57540 AND2X1_LOC_326/A VSS 0.15fF
C3349 AND2X1_LOC_842/B AND2X1_LOC_242/a_8_24# 0.01fF
C11820 AND2X1_LOC_842/B AND2X1_LOC_242/B 0.33fF
C43325 AND2X1_LOC_842/B AND2X1_LOC_842/a_8_24# 0.05fF
C44589 VDD AND2X1_LOC_842/B 0.18fF
C57239 AND2X1_LOC_842/B VSS 0.24fF
C15689 AND2X1_LOC_728/Y AND2X1_LOC_192/Y 0.06fF
C22753 AND2X1_LOC_192/Y AND2X1_LOC_781/Y 0.05fF
C26762 AND2X1_LOC_730/a_8_24# AND2X1_LOC_192/Y 0.03fF
C28188 AND2X1_LOC_192/Y AND2X1_LOC_782/a_8_24# 0.10fF
C3760 AND2X1_LOC_191/Y AND2X1_LOC_475/Y 0.03fF
C37070 AND2X1_LOC_565/B AND2X1_LOC_475/Y 0.31fF
C47199 AND2X1_LOC_475/a_8_24# AND2X1_LOC_475/Y 0.02fF
C32589 AND2X1_LOC_734/Y AND2X1_LOC_550/A 3.04fF
C4335 AND2X1_LOC_170/B AND2X1_LOC_661/A 0.11fF
C24579 AND2X1_LOC_567/a_8_24# AND2X1_LOC_661/A 0.17fF
C25514 AND2X1_LOC_388/a_8_24# AND2X1_LOC_661/A 0.01fF
C43446 AND2X1_LOC_810/a_8_24# AND2X1_LOC_661/A 0.01fF
C45824 AND2X1_LOC_392/A AND2X1_LOC_661/A 0.16fF
C7491 AND2X1_LOC_787/a_8_24# AND2X1_LOC_794/B 0.02fF
C1576 AND2X1_LOC_544/Y AND2X1_LOC_148/Y 0.03fF
C31360 VDD AND2X1_LOC_148/Y 0.29fF
C37606 AND2X1_LOC_148/Y AND2X1_LOC_213/B 0.26fF
C57167 AND2X1_LOC_148/Y VSS 0.14fF
C1954 AND2X1_LOC_728/Y AND2X1_LOC_544/Y 0.03fF
C24972 AND2X1_LOC_728/Y OR2X1_LOC_679/a_8_216# 0.01fF
C27654 AND2X1_LOC_728/Y AND2X1_LOC_797/A 0.18fF
C31436 AND2X1_LOC_728/Y AND2X1_LOC_728/a_8_24# 0.02fF
C50740 AND2X1_LOC_728/Y AND2X1_LOC_191/Y 0.03fF
C53529 AND2X1_LOC_728/Y AND2X1_LOC_209/a_8_24# 0.01fF
C58133 AND2X1_LOC_728/Y VSS 0.08fF
C453 AND2X1_LOC_349/B AND2X1_LOC_359/B 0.31fF
C12710 VDD AND2X1_LOC_349/B 0.08fF
C45536 AND2X1_LOC_349/B AND2X1_LOC_349/a_8_24# 0.01fF
C57727 AND2X1_LOC_349/B VSS 0.15fF
C17801 AND2X1_LOC_228/Y AND2X1_LOC_175/B 0.02fF
C25744 AND2X1_LOC_228/Y AND2X1_LOC_231/a_8_24# 0.01fF
C36453 AND2X1_LOC_228/Y AND2X1_LOC_716/a_8_24# 0.10fF
C18047 AND2X1_LOC_842/a_8_24# AND2X1_LOC_242/B 0.01fF
C19319 VDD AND2X1_LOC_242/B 0.23fF
C34068 AND2X1_LOC_242/B AND2X1_LOC_242/a_8_24# 0.01fF
C55289 AND2X1_LOC_851/B AND2X1_LOC_242/B 0.01fF
C56712 AND2X1_LOC_242/B VSS -0.51fF
C3655 AND2X1_LOC_727/Y AND2X1_LOC_550/A 0.01fF
C9725 AND2X1_LOC_550/A AND2X1_LOC_444/a_8_24# 0.07fF
C13106 AND2X1_LOC_550/a_8_24# AND2X1_LOC_550/A 0.03fF
C15596 AND2X1_LOC_550/A AND2X1_LOC_658/A 9.73fF
C16856 AND2X1_LOC_550/A AND2X1_LOC_476/Y 0.02fF
C20104 AND2X1_LOC_550/A AND2X1_LOC_810/Y 0.03fF
C22468 VDD AND2X1_LOC_550/A 0.16fF
C40527 AND2X1_LOC_727/a_8_24# AND2X1_LOC_550/A 0.07fF
C46306 AND2X1_LOC_544/a_8_24# AND2X1_LOC_550/A 0.02fF
C48795 AND2X1_LOC_544/Y AND2X1_LOC_550/A 0.01fF
C57747 AND2X1_LOC_550/A VSS 0.35fF
C7194 AND2X1_LOC_452/Y AND2X1_LOC_470/B 0.23fF
C12755 AND2X1_LOC_467/a_8_24# AND2X1_LOC_470/B 0.01fF
C49051 VDD OR2X1_LOC_774/B 0.30fF
C52381 OR2X1_LOC_774/B OR2X1_LOC_774/a_8_216# 0.06fF
C56944 OR2X1_LOC_774/B VSS 0.27fF
C19761 OR2X1_LOC_651/A OR2X1_LOC_228/a_8_216# 0.03fF
C37744 VDD OR2X1_LOC_651/A 0.14fF
C57182 OR2X1_LOC_651/A VSS -1.01fF
C9772 OR2X1_LOC_805/A OR2X1_LOC_721/Y 0.02fF
C14116 OR2X1_LOC_805/A OR2X1_LOC_216/a_8_216# 0.01fF
C14375 OR2X1_LOC_493/a_8_216# OR2X1_LOC_805/A 0.04fF
C14618 OR2X1_LOC_805/A OR2X1_LOC_493/Y 0.05fF
C18540 OR2X1_LOC_805/A OR2X1_LOC_362/a_8_216# 0.02fF
C19632 OR2X1_LOC_805/A OR2X1_LOC_216/a_36_216# 0.02fF
C19918 OR2X1_LOC_493/a_36_216# OR2X1_LOC_805/A 0.01fF
C20254 OR2X1_LOC_805/A OR2X1_LOC_392/B 0.10fF
C20808 OR2X1_LOC_805/A OR2X1_LOC_734/a_8_216# 0.06fF
C24103 OR2X1_LOC_805/A OR2X1_LOC_362/a_36_216# 0.02fF
C25647 OR2X1_LOC_805/A OR2X1_LOC_717/a_8_216# 0.06fF
C26288 OR2X1_LOC_805/A OR2X1_LOC_734/a_36_216# 0.01fF
C27269 OR2X1_LOC_476/B OR2X1_LOC_805/A 0.03fF
C31131 OR2X1_LOC_805/A OR2X1_LOC_717/a_36_216# 0.01fF
C37673 OR2X1_LOC_856/B OR2X1_LOC_805/A 0.07fF
C45000 OR2X1_LOC_475/a_8_216# OR2X1_LOC_805/A 0.03fF
C50650 OR2X1_LOC_475/a_36_216# OR2X1_LOC_805/A -0.01fF
C10503 VDD OR2X1_LOC_403/A -0.00fF
C28094 OR2X1_LOC_403/A OR2X1_LOC_403/a_8_216# 0.39fF
C57317 OR2X1_LOC_403/A VSS 0.18fF
C41650 OR2X1_LOC_726/a_8_216# OR2X1_LOC_731/B -0.00fF
C21533 VDD OR2X1_LOC_772/A 0.08fF
C56512 OR2X1_LOC_772/A VSS 0.24fF
C17834 OR2X1_LOC_563/A OR2X1_LOC_493/Y 0.03fF
C28285 OR2X1_LOC_499/a_8_216# OR2X1_LOC_563/A 0.40fF
C45730 OR2X1_LOC_791/a_8_216# OR2X1_LOC_792/A 0.05fF
C57038 OR2X1_LOC_792/A VSS 0.38fF
C24677 VDD OR2X1_LOC_404/A 0.04fF
C57159 OR2X1_LOC_404/A VSS 0.14fF
C27684 OR2X1_LOC_710/a_8_216# OR2X1_LOC_705/Y 0.01fF
C55422 OR2X1_LOC_705/Y OR2X1_LOC_713/a_8_216# 0.03fF
C56519 OR2X1_LOC_705/Y VSS 0.12fF
C23308 OR2X1_LOC_76/Y OR2X1_LOC_486/Y 0.03fF
C4992 OR2X1_LOC_467/A OR2X1_LOC_453/A 0.01fF
C20035 OR2X1_LOC_453/a_8_216# OR2X1_LOC_453/A 0.39fF
C22538 OR2X1_LOC_466/A OR2X1_LOC_453/A 0.01fF
C23792 VDD OR2X1_LOC_453/A -0.00fF
C40316 OR2X1_LOC_449/a_8_216# OR2X1_LOC_453/A -0.00fF
C57073 OR2X1_LOC_453/A VSS 0.18fF
C33144 OR2X1_LOC_76/Y OR2X1_LOC_445/a_8_216# 0.40fF
C48333 OR2X1_LOC_76/Y OR2X1_LOC_76/a_8_216# 0.01fF
C48522 VDD OR2X1_LOC_76/Y 0.13fF
C50328 OR2X1_LOC_76/Y OR2X1_LOC_455/a_8_216# 0.08fF
C51155 OR2X1_LOC_675/a_8_216# OR2X1_LOC_76/Y 0.13fF
C57315 OR2X1_LOC_76/Y VSS 0.37fF
C10499 OR2X1_LOC_340/a_8_216# OR2X1_LOC_560/A 0.39fF
C23928 OR2X1_LOC_509/a_8_216# OR2X1_LOC_560/A 0.01fF
C33676 OR2X1_LOC_721/Y OR2X1_LOC_560/A 0.05fF
C44229 OR2X1_LOC_392/B OR2X1_LOC_560/A 0.03fF
C18387 OR2X1_LOC_632/Y OR2X1_LOC_493/Y 0.10fF
C34681 OR2X1_LOC_493/Y OR2X1_LOC_558/a_8_216# 0.05fF
C44259 VDD OR2X1_LOC_493/Y 1.69fF
C46962 OR2X1_LOC_499/a_8_216# OR2X1_LOC_493/Y 0.28fF
C48611 OR2X1_LOC_343/a_8_216# OR2X1_LOC_493/Y 0.29fF
C56327 OR2X1_LOC_493/Y VSS 0.73fF
C32939 VDD OR2X1_LOC_785/B 0.33fF
C45775 OR2X1_LOC_785/a_8_216# OR2X1_LOC_785/B 0.03fF
C56721 OR2X1_LOC_785/B VSS 0.08fF
C46823 VDD OR2X1_LOC_443/Y 0.12fF
C57312 OR2X1_LOC_443/Y VSS 0.19fF
C13499 OR2X1_LOC_148/Y OR2X1_LOC_213/A 0.28fF
C51934 OR2X1_LOC_213/A OR2X1_LOC_209/a_8_216# 0.01fF
C29284 OR2X1_LOC_467/a_8_216# OR2X1_LOC_470/A -0.00fF
C47912 OR2X1_LOC_148/Y OR2X1_LOC_149/a_8_216# 0.39fF
C57857 OR2X1_LOC_148/Y VSS 0.18fF
C14200 VDD OR2X1_LOC_730/B 0.05fF
C19755 OR2X1_LOC_730/a_8_216# OR2X1_LOC_730/B 0.01fF
C56323 OR2X1_LOC_730/B VSS 0.11fF
C9631 OR2X1_LOC_858/B OR2X1_LOC_349/A 0.02fF
C54690 OR2X1_LOC_850/a_8_216# OR2X1_LOC_349/A 0.01fF
C56343 OR2X1_LOC_349/A VSS 0.26fF
C3635 OR2X1_LOC_244/B OR2X1_LOC_392/B 0.03fF
C36651 OR2X1_LOC_508/a_8_216# OR2X1_LOC_244/B 0.40fF
C49295 OR2X1_LOC_244/B OR2X1_LOC_721/Y 1.26fF
C395 AND2X1_LOC_453/a_8_24# AND2X1_LOC_452/Y 0.02fF
C1689 AND2X1_LOC_452/Y AND2X1_LOC_467/a_8_24# 0.05fF
C24159 VDD AND2X1_LOC_452/Y 0.89fF
C35117 AND2X1_LOC_605/Y AND2X1_LOC_452/Y 0.01fF
C40967 AND2X1_LOC_452/Y AND2X1_LOC_605/a_8_24# 0.02fF
C46359 AND2X1_LOC_454/Y AND2X1_LOC_452/Y 0.07fF
C56674 AND2X1_LOC_452/Y VSS 0.14fF
C1460 AND2X1_LOC_191/Y AND2X1_LOC_781/Y 0.03fF
C4919 AND2X1_LOC_191/Y AND2X1_LOC_192/a_36_24# 0.01fF
C9321 AND2X1_LOC_191/Y AND2X1_LOC_476/Y 1.50fF
C10749 AND2X1_LOC_191/Y AND2X1_LOC_797/A 0.03fF
C14829 AND2X1_LOC_191/Y VDD 0.69fF
C20959 AND2X1_LOC_191/Y AND2X1_LOC_475/a_8_24# 0.05fF
C21187 AND2X1_LOC_191/Y AND2X1_LOC_213/B 0.04fF
C28404 AND2X1_LOC_501/Y AND2X1_LOC_191/Y 0.03fF
C31888 AND2X1_LOC_191/Y AND2X1_LOC_475/a_36_24# 0.01fF
C36389 AND2X1_LOC_209/a_8_24# AND2X1_LOC_191/Y 0.06fF
C50135 AND2X1_LOC_191/Y AND2X1_LOC_192/a_8_24# 0.01fF
C52200 AND2X1_LOC_727/Y AND2X1_LOC_191/Y 0.04fF
C57884 AND2X1_LOC_191/Y VSS -1.39fF
C3040 AND2X1_LOC_392/A AND2X1_LOC_170/B 0.03fF
C6794 VDD AND2X1_LOC_170/B 0.12fF
C17959 AND2X1_LOC_170/Y AND2X1_LOC_170/B 0.01fF
C43855 AND2X1_LOC_170/a_8_24# AND2X1_LOC_170/B -0.00fF
C57279 AND2X1_LOC_170/B VSS 0.19fF
C21126 AND2X1_LOC_443/Y AND2X1_LOC_444/a_8_24# 0.03fF
C27022 AND2X1_LOC_658/A AND2X1_LOC_443/Y 0.09fF
C32059 AND2X1_LOC_443/Y AND2X1_LOC_444/a_36_24# 0.01fF
C33767 VDD AND2X1_LOC_443/Y 0.21fF
C56736 AND2X1_LOC_443/Y VSS -0.09fF
C22329 AND2X1_LOC_641/Y AND2X1_LOC_641/a_8_24# 0.01fF
C1651 AND2X1_LOC_175/B AND2X1_LOC_654/B 0.01fF
C14912 AND2X1_LOC_175/B AND2X1_LOC_175/a_8_24# 0.01fF
C33834 VDD AND2X1_LOC_175/B 0.23fF
C13387 AND2X1_LOC_719/Y AND2X1_LOC_241/a_36_24# 0.06fF
C34145 AND2X1_LOC_719/Y AND2X1_LOC_190/a_8_24# 0.29fF
C36443 AND2X1_LOC_719/Y AND2X1_LOC_849/a_8_24# 0.23fF
C44490 AND2X1_LOC_719/Y AND2X1_LOC_859/a_36_24# 0.06fF
C46751 AND2X1_LOC_719/Y AND2X1_LOC_719/a_8_24# 0.01fF
C50917 AND2X1_LOC_719/Y AND2X1_LOC_190/a_36_24# 0.06fF
C52111 AND2X1_LOC_719/Y AND2X1_LOC_542/a_8_24# 0.11fF
C52959 AND2X1_LOC_719/Y AND2X1_LOC_241/a_8_24# 0.25fF
C53220 AND2X1_LOC_719/Y AND2X1_LOC_849/a_36_24# 0.08fF
C6058 AND2X1_LOC_773/Y AND2X1_LOC_774/A 0.01fF
C7357 AND2X1_LOC_773/Y AND2X1_LOC_772/Y 0.17fF
C18451 AND2X1_LOC_773/Y AND2X1_LOC_774/a_8_24# 0.11fF
C32402 AND2X1_LOC_773/Y VDD 1.46fF
C58124 AND2X1_LOC_773/Y VSS 0.35fF
C38452 AND2X1_LOC_193/a_8_24# AND2X1_LOC_194/Y 0.01fF
C40075 AND2X1_LOC_194/a_8_24# AND2X1_LOC_194/Y 0.02fF
C33359 VDD AND2X1_LOC_404/A 0.21fF
C38993 AND2X1_LOC_404/A AND2X1_LOC_404/a_8_24# 0.18fF
C56634 AND2X1_LOC_404/A VSS 0.06fF
C25563 AND2X1_LOC_839/A AND2X1_LOC_839/a_8_24# 0.10fF
C56984 AND2X1_LOC_839/A VSS 0.16fF
C9708 VDD AND2X1_LOC_123/Y 0.02fF
C28847 AND2X1_LOC_123/Y AND2X1_LOC_124/a_8_24# 0.01fF
C30573 AND2X1_LOC_123/a_8_24# AND2X1_LOC_123/Y 0.01fF
C57330 AND2X1_LOC_123/Y VSS 0.08fF
C27429 AND2X1_LOC_675/Y AND2X1_LOC_508/B 0.02fF
C32938 AND2X1_LOC_574/a_8_24# AND2X1_LOC_675/Y 0.18fF
C34400 AND2X1_LOC_675/Y AND2X1_LOC_675/a_8_24# 0.01fF
C35226 AND2X1_LOC_675/Y AND2X1_LOC_675/A 0.02fF
C28412 AND2X1_LOC_501/Y AND2X1_LOC_711/Y 0.03fF
C33792 AND2X1_LOC_605/Y AND2X1_LOC_454/a_8_24# 0.01fF
C41287 AND2X1_LOC_605/Y AND2X1_LOC_449/a_8_24# 0.11fF
C41346 AND2X1_LOC_712/a_8_24# AND2X1_LOC_605/Y 0.01fF
C2601 AND2X1_LOC_675/A AND2X1_LOC_476/Y 0.05fF
C8120 VDD AND2X1_LOC_675/A 0.82fF
C19473 AND2X1_LOC_675/A AND2X1_LOC_439/a_8_24# 0.01fF
C31871 AND2X1_LOC_544/a_8_24# AND2X1_LOC_675/A 0.20fF
C42887 AND2X1_LOC_675/A AND2X1_LOC_784/a_8_24# 0.04fF
C42929 AND2X1_LOC_675/A AND2X1_LOC_471/Y 0.04fF
C56958 AND2X1_LOC_675/A VSS 0.07fF
C1903 AND2X1_LOC_544/Y AND2X1_LOC_545/a_8_24# 0.04fF
C22028 AND2X1_LOC_544/Y AND2X1_LOC_728/a_8_24# 0.03fF
C32963 AND2X1_LOC_544/Y AND2X1_LOC_728/a_36_24# 0.01fF
C37514 AND2X1_LOC_148/a_8_24# AND2X1_LOC_213/B 0.01fF
C48895 AND2X1_LOC_149/a_8_24# AND2X1_LOC_213/B 0.01fF
C49913 AND2X1_LOC_213/B AND2X1_LOC_783/a_8_24# 0.01fF
C7732 AND2X1_LOC_259/Y AND2X1_LOC_345/a_8_24# 0.10fF
C10809 AND2X1_LOC_259/Y AND2X1_LOC_259/a_8_24# 0.01fF
C14791 AND2X1_LOC_259/Y AND2X1_LOC_346/a_8_24# 0.20fF
C49802 VDD AND2X1_LOC_259/Y 0.21fF
C57609 AND2X1_LOC_259/Y VSS 0.49fF
C18577 AND2X1_LOC_781/a_8_24# AND2X1_LOC_781/Y 0.01fF
C38642 VDD AND2X1_LOC_781/Y 0.06fF
C56353 AND2X1_LOC_781/Y VSS 0.18fF
C206 VDD AND2X1_LOC_508/B 0.27fF
C24487 AND2X1_LOC_509/Y AND2X1_LOC_508/B 0.12fF
C49668 AND2X1_LOC_508/B AND2X1_LOC_658/A 0.03fF
C57426 AND2X1_LOC_508/B VSS 0.16fF
C16019 AND2X1_LOC_392/A AND2X1_LOC_365/A 0.02fF
C40282 AND2X1_LOC_365/A AND2X1_LOC_336/a_8_24# 0.20fF
C3346 AND2X1_LOC_392/A AND2X1_LOC_170/Y 0.17fF
C13160 AND2X1_LOC_392/A AND2X1_LOC_123/a_8_24# 0.03fF
C15550 AND2X1_LOC_392/A AND2X1_LOC_392/a_36_24# 0.01fF
C15933 AND2X1_LOC_392/A AND2X1_LOC_337/a_8_24# 0.02fF
C17097 AND2X1_LOC_392/A AND2X1_LOC_772/a_8_24# 0.06fF
C18192 AND2X1_LOC_392/A AND2X1_LOC_560/B 0.07fF
C29655 AND2X1_LOC_392/A AND2X1_LOC_123/a_36_24# 0.01fF
C45946 AND2X1_LOC_392/A AND2X1_LOC_810/Y 0.07fF
C48389 AND2X1_LOC_392/A VDD 0.49fF
C49681 AND2X1_LOC_392/A AND2X1_LOC_392/a_8_24# 0.05fF
C58101 AND2X1_LOC_392/A VSS 0.61fF
C33002 OR2X1_LOC_474/a_8_216# OR2X1_LOC_474/B 0.18fF
C53789 OR2X1_LOC_392/B OR2X1_LOC_474/B 0.16fF
C19035 OR2X1_LOC_640/Y OR2X1_LOC_640/a_8_216# -0.00fF
C6275 AND2X1_LOC_719/a_36_24# AND2X1_LOC_658/A 0.01fF
C7436 AND2X1_LOC_727/a_8_24# AND2X1_LOC_658/A 0.03fF
C8064 AND2X1_LOC_711/Y AND2X1_LOC_658/A 0.01fF
C10112 AND2X1_LOC_546/a_8_24# AND2X1_LOC_658/A 0.04fF
C13085 AND2X1_LOC_544/a_8_24# AND2X1_LOC_658/A 0.04fF
C13471 AND2X1_LOC_509/Y AND2X1_LOC_658/A 0.03fF
C24058 AND2X1_LOC_727/a_36_24# AND2X1_LOC_658/A 0.01fF
C24137 AND2X1_LOC_544/a_36_24# AND2X1_LOC_658/A 0.01fF
C24499 AND2X1_LOC_510/a_8_24# AND2X1_LOC_658/A 0.05fF
C26657 AND2X1_LOC_546/a_36_24# AND2X1_LOC_658/A 0.01fF
C32469 AND2X1_LOC_658/A AND2X1_LOC_444/a_8_24# 0.04fF
C40955 AND2X1_LOC_510/a_36_24# AND2X1_LOC_658/A 0.01fF
C43590 AND2X1_LOC_658/A AND2X1_LOC_444/a_36_24# 0.01fF
C51462 AND2X1_LOC_719/a_8_24# AND2X1_LOC_658/A 0.02fF
C4012 AND2X1_LOC_711/Y AND2X1_LOC_623/a_8_24# 0.07fF
C5416 AND2X1_LOC_550/a_8_24# AND2X1_LOC_711/Y 0.04fF
C7988 AND2X1_LOC_711/Y AND2X1_LOC_726/a_8_24# 0.04fF
C9336 AND2X1_LOC_711/Y AND2X1_LOC_476/Y 0.07fF
C10999 AND2X1_LOC_565/B AND2X1_LOC_711/Y 0.08fF
C13584 AND2X1_LOC_711/Y AND2X1_LOC_507/a_8_24# 0.05fF
C14839 VDD AND2X1_LOC_711/Y 0.92fF
C15005 AND2X1_LOC_711/Y AND2X1_LOC_624/a_8_24# 0.01fF
C16509 AND2X1_LOC_550/a_36_24# AND2X1_LOC_711/Y 0.01fF
C17381 AND2X1_LOC_711/Y AND2X1_LOC_501/a_8_24# 0.05fF
C23678 AND2X1_LOC_711/Y AND2X1_LOC_791/a_8_24# 0.01fF
C24629 AND2X1_LOC_711/Y AND2X1_LOC_507/a_36_24# 0.01fF
C27578 AND2X1_LOC_711/a_8_24# AND2X1_LOC_711/Y 0.01fF
C35495 AND2X1_LOC_191/a_8_24# AND2X1_LOC_711/Y 0.08fF
C39427 AND2X1_LOC_711/Y AND2X1_LOC_501/a_36_24# 0.01fF
C51377 AND2X1_LOC_711/Y AND2X1_LOC_792/a_8_24# 0.01fF
C51581 AND2X1_LOC_711/Y AND2X1_LOC_620/a_8_24# 0.01fF
C52214 AND2X1_LOC_727/Y AND2X1_LOC_711/Y 0.03fF
C57820 AND2X1_LOC_711/Y VSS 0.27fF
C578 OR2X1_LOC_721/Y OR2X1_LOC_523/a_8_216# 0.29fF
C37079 OR2X1_LOC_392/B OR2X1_LOC_721/Y 0.10fF
C37614 OR2X1_LOC_721/Y OR2X1_LOC_734/a_8_216# 0.02fF
C39291 VDD OR2X1_LOC_721/Y 1.36fF
C41106 OR2X1_LOC_720/a_8_216# OR2X1_LOC_721/Y 0.01fF
C45708 OR2X1_LOC_721/a_8_216# OR2X1_LOC_721/Y 0.01fF
C56567 OR2X1_LOC_721/Y VSS 0.66fF
C2065 VDD OR2X1_LOC_849/A 0.12fF
C5353 OR2X1_LOC_849/A OR2X1_LOC_768/a_8_216# 0.01fF
C22561 OR2X1_LOC_849/A OR2X1_LOC_624/a_8_216# 0.01fF
C57672 OR2X1_LOC_849/A VSS -0.41fF
C7355 AND2X1_LOC_785/a_8_24# AND2X1_LOC_785/Y 0.11fF
C44181 AND2X1_LOC_170/a_8_24# AND2X1_LOC_170/Y 0.01fF
C1387 AND2X1_LOC_326/a_8_24# AND2X1_LOC_354/B 0.04fF
C1624 VDD AND2X1_LOC_354/B 0.10fF
C21338 AND2X1_LOC_715/a_8_24# AND2X1_LOC_354/B 0.01fF
C23884 AND2X1_LOC_354/B AND2X1_LOC_854/a_8_24# 0.04fF
C53482 AND2X1_LOC_715/Y AND2X1_LOC_354/B 0.09fF
C57128 AND2X1_LOC_354/B VSS 0.16fF
C27511 VDD AND2X1_LOC_472/B 0.21fF
C56904 AND2X1_LOC_472/B VSS 0.30fF
C52302 AND2X1_LOC_174/a_8_24# AND2X1_LOC_654/B 0.01fF
C26458 AND2X1_LOC_727/Y AND2X1_LOC_726/a_8_24# 0.01fF
C51658 AND2X1_LOC_727/Y AND2X1_LOC_727/a_8_24# 0.01fF
C13585 AND2X1_LOC_209/a_8_24# AND2X1_LOC_797/A 0.03fF
C38243 AND2X1_LOC_149/a_8_24# AND2X1_LOC_797/A 0.01fF
C38636 AND2X1_LOC_730/a_8_24# AND2X1_LOC_797/A 0.09fF
C4924 OR2X1_LOC_653/a_8_216# OR2X1_LOC_392/B 0.40fF
C10566 OR2X1_LOC_849/a_8_216# OR2X1_LOC_392/B 0.10fF
C16335 OR2X1_LOC_475/a_8_216# OR2X1_LOC_392/B 0.12fF
C24830 OR2X1_LOC_508/a_8_216# OR2X1_LOC_392/B 0.13fF
C31699 OR2X1_LOC_392/B OR2X1_LOC_392/a_8_216# 0.08fF
C35767 OR2X1_LOC_508/a_36_216# OR2X1_LOC_392/B 0.13fF
C44516 OR2X1_LOC_476/a_8_216# OR2X1_LOC_392/B 0.04fF
C50030 VDD OR2X1_LOC_392/B 2.02fF
C56764 OR2X1_LOC_392/B VSS 0.65fF
C17928 OR2X1_LOC_508/Y OR2X1_LOC_510/a_8_216# 0.02fF
C28962 OR2X1_LOC_508/Y OR2X1_LOC_510/a_36_216# 0.02fF
C29439 VDD OR2X1_LOC_508/Y 0.19fF
C35798 OR2X1_LOC_507/a_8_216# OR2X1_LOC_508/Y 0.01fF
C56498 OR2X1_LOC_508/Y VSS -0.12fF
C11417 OR2X1_LOC_466/A OR2X1_LOC_449/a_8_216# 0.40fF
C27626 OR2X1_LOC_454/a_8_216# OR2X1_LOC_466/A -0.00fF
C32022 OR2X1_LOC_467/A OR2X1_LOC_466/A 0.01fF
C47189 OR2X1_LOC_453/a_8_216# OR2X1_LOC_466/A 0.01fF
C14547 OR2X1_LOC_207/B OR2X1_LOC_193/a_8_216# 0.05fF
C36869 OR2X1_LOC_170/a_8_216# OR2X1_LOC_568/A 0.03fF
C39769 OR2X1_LOC_567/a_8_216# OR2X1_LOC_568/A 0.13fF
C54193 OR2X1_LOC_169/a_8_216# OR2X1_LOC_568/A 0.03fF
C5490 OR2X1_LOC_856/B OR2X1_LOC_856/a_8_216# 0.05fF
C10151 OR2X1_LOC_854/a_8_216# OR2X1_LOC_856/B 0.01fF
C11342 VDD OR2X1_LOC_856/B 0.27fF
C16494 OR2X1_LOC_856/B OR2X1_LOC_623/a_8_216# 0.02fF
C57797 OR2X1_LOC_856/B VSS 0.30fF
C53807 OR2X1_LOC_201/a_8_216# OR2X1_LOC_206/A 0.01fF
C18290 AND2X1_LOC_647/Y AND2X1_LOC_772/Y 0.01fF
C43396 VDD AND2X1_LOC_647/Y 0.41fF
C44008 AND2X1_LOC_647/Y AND2X1_LOC_646/a_8_24# 0.04fF
C51393 AND2X1_LOC_647/Y AND2X1_LOC_656/a_8_24# 0.11fF
C56871 AND2X1_LOC_647/Y VSS -0.25fF
C1347 AND2X1_LOC_719/a_8_24# AND2X1_LOC_859/Y 0.03fF
C10256 OR2X1_LOC_467/A OR2X1_LOC_454/a_8_216# 0.01fF
C16453 OR2X1_LOC_467/A OR2X1_LOC_467/a_8_216# 0.04fF
C29625 OR2X1_LOC_467/A OR2X1_LOC_453/a_8_216# 0.01fF
C33316 VDD OR2X1_LOC_467/A 0.20fF
C50209 OR2X1_LOC_467/A OR2X1_LOC_449/a_8_216# 0.01fF
C57504 OR2X1_LOC_467/A VSS -0.19fF
C33656 OR2X1_LOC_840/a_8_216# OR2X1_LOC_723/B 0.03fF
C39144 OR2X1_LOC_840/a_36_216# OR2X1_LOC_723/B 0.02fF
C44999 OR2X1_LOC_723/B OR2X1_LOC_717/a_8_216# 0.01fF
C50648 OR2X1_LOC_723/B OR2X1_LOC_717/a_36_216# 0.02fF
C30678 OR2X1_LOC_566/A OR2X1_LOC_336/a_8_216# 0.01fF
C31527 OR2X1_LOC_303/a_8_216# OR2X1_LOC_566/A 0.01fF
C16059 AND2X1_LOC_509/Y AND2X1_LOC_474/a_8_24# 0.20fF
C20256 AND2X1_LOC_509/Y VDD 0.27fF
C24494 AND2X1_LOC_509/Y AND2X1_LOC_508/a_8_24# 0.01fF
C27440 AND2X1_LOC_509/Y AND2X1_LOC_509/a_8_24# 0.01fF
C57919 AND2X1_LOC_509/Y VSS 0.03fF
C48426 AND2X1_LOC_703/a_8_24# AND2X1_LOC_724/A 0.01fF
C52622 AND2X1_LOC_712/a_8_24# AND2X1_LOC_454/Y 0.21fF
C7339 AND2X1_LOC_772/Y AND2X1_LOC_773/a_8_24# 0.07fF
C20241 AND2X1_LOC_656/a_36_24# AND2X1_LOC_772/Y 0.01fF
C26928 VDD AND2X1_LOC_772/Y 0.75fF
C34804 AND2X1_LOC_656/a_8_24# AND2X1_LOC_772/Y 0.02fF
C37578 AND2X1_LOC_140/a_8_24# AND2X1_LOC_772/Y -0.00fF
C56272 AND2X1_LOC_772/Y VSS 0.29fF
C83 AND2X1_LOC_849/a_8_24# AND2X1_LOC_806/A 0.01fF
C6814 AND2X1_LOC_288/a_8_24# AND2X1_LOC_806/A 0.01fF
C37709 AND2X1_LOC_850/a_8_24# AND2X1_LOC_806/A 0.01fF
C23593 OR2X1_LOC_632/Y OR2X1_LOC_500/a_8_216# 0.02fF
C34502 OR2X1_LOC_632/Y OR2X1_LOC_500/a_36_216# 0.01fF
C38730 OR2X1_LOC_632/Y OR2X1_LOC_501/a_8_216# 0.02fF
C39209 OR2X1_LOC_632/Y OR2X1_LOC_554/a_8_216# 0.40fF
C44335 OR2X1_LOC_632/Y OR2X1_LOC_501/a_36_216# 0.01fF
C26616 OR2X1_LOC_850/a_8_216# OR2X1_LOC_858/B -0.00fF
C50927 OR2X1_LOC_362/B OR2X1_LOC_362/a_8_216# 0.07fF
C8464 AND2X1_LOC_720/Y AND2X1_LOC_721/a_8_24# 0.19fF
C55583 AND2X1_LOC_720/Y VDD 0.24fF
C58052 AND2X1_LOC_720/Y VSS 0.07fF
C11652 AND2X1_LOC_774/a_8_24# AND2X1_LOC_774/A 0.04fF
C22786 AND2X1_LOC_774/a_36_24# AND2X1_LOC_774/A 0.01fF
C25695 VDD AND2X1_LOC_774/A 0.75fF
C56355 AND2X1_LOC_774/A VSS -1.63fF
C40170 AND2X1_LOC_642/a_8_24# AND2X1_LOC_642/Y 0.02fF
C27127 AND2X1_LOC_768/a_8_24# AND2X1_LOC_560/B 0.02fF
C38475 AND2X1_LOC_553/a_8_24# AND2X1_LOC_560/B 0.02fF
C34812 AND2X1_LOC_471/a_8_24# AND2X1_LOC_471/Y 0.04fF
C48630 AND2X1_LOC_440/a_8_24# AND2X1_LOC_471/Y 0.20fF
C1695 AND2X1_LOC_851/B AND2X1_LOC_445/a_8_24# 0.04fF
C16092 AND2X1_LOC_851/B AND2X1_LOC_455/a_8_24# 0.03fF
C21829 AND2X1_LOC_523/a_8_24# AND2X1_LOC_851/B 0.01fF
C44135 AND2X1_LOC_851/B AND2X1_LOC_241/a_8_24# 0.02fF
C13914 AND2X1_LOC_715/Y AND2X1_LOC_854/a_8_24# 0.20fF
C29083 AND2X1_LOC_715/Y AND2X1_LOC_703/a_8_24# 0.03fF
C205 AND2X1_LOC_565/B AND2X1_LOC_565/a_8_24# 0.01fF
C42685 AND2X1_LOC_565/B AND2X1_LOC_476/Y 0.04fF
C48396 AND2X1_LOC_565/B VDD 0.48fF
C58072 AND2X1_LOC_565/B VSS 0.28fF
C4773 AND2X1_LOC_856/a_8_24# AND2X1_LOC_863/A 0.02fF
C17131 AND2X1_LOC_324/a_8_24# AND2X1_LOC_863/A 0.11fF
C4699 OR2X1_LOC_216/Y OR2X1_LOC_216/a_8_216# 0.02fF
C1168 AND2X1_LOC_721/a_8_24# AND2X1_LOC_366/A 0.04fF
C1834 AND2X1_LOC_476/Y AND2X1_LOC_439/a_8_24# 0.04fF
C1895 AND2X1_LOC_542/a_8_24# AND2X1_LOC_476/Y 0.01fF
C9274 AND2X1_LOC_775/a_8_24# AND2X1_LOC_476/Y 0.03fF
C14300 AND2X1_LOC_544/a_8_24# AND2X1_LOC_476/Y 0.02fF
C18489 AND2X1_LOC_542/a_36_24# AND2X1_LOC_476/Y -0.02fF
C25244 AND2X1_LOC_552/a_8_24# AND2X1_LOC_476/Y 0.03fF
C36192 AND2X1_LOC_552/a_36_24# AND2X1_LOC_476/Y 0.01fF
C37069 AND2X1_LOC_550/a_8_24# AND2X1_LOC_476/Y 0.03fF
C1949 AND2X1_LOC_810/Y AND2X1_LOC_486/a_8_24# 0.03fF
C11892 AND2X1_LOC_727/a_8_24# AND2X1_LOC_810/Y 0.02fF
C41705 AND2X1_LOC_810/Y AND2X1_LOC_653/a_8_24# 0.09fF
C42111 AND2X1_LOC_652/a_8_24# AND2X1_LOC_810/Y 0.07fF
C43529 AND2X1_LOC_810/a_8_24# AND2X1_LOC_810/Y 0.01fF
C52926 AND2X1_LOC_810/Y AND2X1_LOC_653/a_36_24# 0.01fF
C819 VDD OR2X1_LOC_476/B 1.07fF
C1002 OR2X1_LOC_476/B OR2X1_LOC_476/a_36_216# 0.03fF
C13671 OR2X1_LOC_476/B OR2X1_LOC_61/a_8_216# 0.04fF
C19179 OR2X1_LOC_476/B OR2X1_LOC_61/a_36_216# 0.01fF
C39576 OR2X1_LOC_472/a_8_216# OR2X1_LOC_476/B 0.01fF
C43666 OR2X1_LOC_476/B OR2X1_LOC_390/a_8_216# 0.01fF
C49325 OR2X1_LOC_476/B OR2X1_LOC_390/a_36_216# 0.03fF
C50824 OR2X1_LOC_472/a_36_216# OR2X1_LOC_476/B -0.01fF
C51640 OR2X1_LOC_476/B OR2X1_LOC_476/a_8_216# 0.02fF
C57632 OR2X1_LOC_476/B VSS -1.86fF
C12914 OR2X1_LOC_244/A OR2X1_LOC_204/a_8_216# 0.04fF
C18493 OR2X1_LOC_244/A OR2X1_LOC_84/a_8_216# 0.04fF
C41294 OR2X1_LOC_243/a_8_216# OR2X1_LOC_244/A 0.05fF
C47002 OR2X1_LOC_243/a_36_216# OR2X1_LOC_244/A 0.01fF
C54991 OR2X1_LOC_139/a_8_216# OR2X1_LOC_244/A -0.05fF
C51534 VDD OR2X1_LOC_852/A 0.12fF
C57357 OR2X1_LOC_852/A VSS 0.18fF
C57602 AND2X1_LOC_354/Y VSS 0.08fF
C24296 OR2X1_LOC_474/Y OR2X1_LOC_849/a_8_216# 0.06fF
C27900 OR2X1_LOC_474/Y OR2X1_LOC_624/a_8_216# 0.39fF
C40721 OR2X1_LOC_474/a_8_216# OR2X1_LOC_474/Y 0.02fF
C57438 OR2X1_LOC_474/Y VSS -1.48fF
C9684 AND2X1_LOC_810/A AND2X1_LOC_854/a_8_24# 0.01fF
C14410 AND2X1_LOC_810/A AND2X1_LOC_856/a_8_24# 0.01fF
C19419 AND2X1_LOC_810/A AND2X1_LOC_388/a_8_24# 0.01fF
C27454 AND2X1_LOC_810/A AND2X1_LOC_354/a_8_24# 0.01fF
C55806 OR2X1_LOC_465/a_8_216# OR2X1_LOC_465/B 0.01fF
C38066 OR2X1_LOC_507/a_8_216# OR2X1_LOC_510/Y 0.40fF
C44132 OR2X1_LOC_510/Y OR2X1_LOC_574/a_8_216# 0.07fF
C49813 OR2X1_LOC_208/a_36_216# OR2X1_LOC_35/Y 0.03fF
C56851 AND2X1_LOC_474/Y VSS -0.28fF
C35330 VDD OR2X1_LOC_356/B 0.27fF
C56335 OR2X1_LOC_356/B VSS 0.36fF
C54608 AND2X1_LOC_465/Y AND2X1_LOC_471/a_8_24# 0.11fF
C52040 AND2X1_LOC_859/a_8_24# AND2X1_LOC_859/B 0.12fF
C5644 AND2X1_LOC_539/Y AND2X1_LOC_567/a_8_24# 0.04fF
C24646 AND2X1_LOC_539/Y AND2X1_LOC_810/a_8_24# 0.01fF
C21200 OR2X1_LOC_216/A OR2X1_LOC_475/a_8_216# 0.03fF
C20220 AND2X1_LOC_540/a_8_24# AND2X1_LOC_465/A 0.01fF
C40869 AND2X1_LOC_181/a_8_24# AND2X1_LOC_465/A 0.01fF
C44038 AND2X1_LOC_465/a_8_24# AND2X1_LOC_465/A 0.08fF
C56742 AND2X1_LOC_465/A VSS 0.28fF
C50156 VDD AND2X1_LOC_653/B 0.22fF
C37494 AND2X1_LOC_116/Y AND2X1_LOC_216/a_8_24# 0.02fF
C21648 AND2X1_LOC_510/a_8_24# AND2X1_LOC_573/A 0.01fF
C35373 AND2X1_LOC_561/a_8_24# AND2X1_LOC_573/A 0.01fF
C38096 AND2X1_LOC_573/A AND2X1_LOC_474/a_8_24# 0.01fF
C49750 AND2X1_LOC_509/a_8_24# AND2X1_LOC_573/A 0.01fF
C52165 AND2X1_LOC_554/a_8_24# AND2X1_LOC_573/A 0.01fF
C53244 AND2X1_LOC_140/a_8_24# AND2X1_LOC_573/A 0.01fF
C17588 OR2X1_LOC_854/a_8_216# OR2X1_LOC_319/Y 0.06fF
C4491 OR2X1_LOC_404/Y OR2X1_LOC_500/a_8_216# 0.02fF
C24508 OR2X1_LOC_404/Y OR2X1_LOC_523/a_8_216# 0.02fF
C52853 OR2X1_LOC_653/A OR2X1_LOC_653/a_8_216# 0.01fF

.ends

* wrdata outputs.out V("OR2X1_LOC_351/B") V("OR2X1_LOC_852/A") V("OR2X1_LOC_244/A") V("OR2X1_LOC_476/B") V("AND2X1_LOC_810/Y") V("AND2X1_LOC_476/Y") V("AND2X1_LOC_366/A") V("OR2X1_LOC_656/Y") V("OR2X1_LOC_216/Y") V("AND2X1_LOC_863/A") V("AND2X1_LOC_739/B") V("AND2X1_LOC_565/B") V("AND2X1_LOC_715/Y") V("AND2X1_LOC_339/Y") V("AND2X1_LOC_851/B") V("AND2X1_LOC_796/A") V("AND2X1_LOC_471/Y") V("AND2X1_LOC_560/B") V("AND2X1_LOC_642/Y") V("AND2X1_LOC_207/A") V("AND2X1_LOC_851/A") V("AND2X1_LOC_720/Y") V("AND2X1_LOC_359/B") V("OR2X1_LOC_362/B") V("OR2X1_LOC_858/B") V("OR2X1_LOC_632/Y") V("AND2X1_LOC_806/A") V("AND2X1_LOC_772/Y") V("AND2X1_LOC_338/Y") V("AND2X1_LOC_454/Y") V("AND2X1_LOC_724/A") V("AND2X1_LOC_340/Y") V("OR2X1_LOC_566/A") V("OR2X1_LOC_723/B") V("OR2X1_LOC_564/A") V("OR2X1_LOC_467/A") V("AND2X1_LOC_859/Y") V("AND2X1_LOC_647/Y") V("OR2X1_LOC_206/A") V("OR2X1_LOC_856/B") V("OR2X1_LOC_568/A") V("OR2X1_LOC_207/B") V("OR2X1_LOC_141/B") V("OR2X1_LOC_857/B") V("OR2X1_LOC_466/A") V("OR2X1_LOC_392/B") V("AND2X1_LOC_797/A") V("AND2X1_LOC_357/B") V("AND2X1_LOC_727/Y") V("AND2X1_LOC_712/Y") V("AND2X1_LOC_654/B") V("AND2X1_LOC_472/B") V("AND2X1_LOC_717/Y") V("AND2X1_LOC_170/Y") V("AND2X1_LOC_785/Y") V("OR2X1_LOC_721/Y") V("AND2X1_LOC_713/Y") V("AND2X1_LOC_711/Y") V("AND2X1_LOC_658/A") V("OR2X1_LOC_640/Y") V("OR2X1_LOC_563/B") V("OR2X1_LOC_784/Y") V("OR2X1_LOC_569/A") V("OR2X1_LOC_474/B") V("AND2X1_LOC_392/A") V("AND2X1_LOC_644/Y") V("AND2X1_LOC_365/A") V("AND2X1_LOC_508/B") V("AND2X1_LOC_781/Y") V("AND2X1_LOC_259/Y") V("AND2X1_LOC_213/B") V("AND2X1_LOC_544/Y") V("AND2X1_LOC_675/A") V("AND2X1_LOC_605/Y") V("AND2X1_LOC_501/Y") V("AND2X1_LOC_675/Y") V("AND2X1_LOC_123/Y") V("AND2X1_LOC_839/A") V("AND2X1_LOC_182/A") V("AND2X1_LOC_194/Y") V("AND2X1_LOC_719/Y") V("AND2X1_LOC_175/B") V("AND2X1_LOC_641/Y") V("AND2X1_LOC_551/B") V("AND2X1_LOC_443/Y") V("AND2X1_LOC_170/B") V("AND2X1_LOC_191/Y") V("AND2X1_LOC_452/Y") V("OR2X1_LOC_244/B") V("OR2X1_LOC_349/A") V("OR2X1_LOC_730/B") V("OR2X1_LOC_148/Y") V("OR2X1_LOC_470/A") V("OR2X1_LOC_213/A") V("OR2X1_LOC_443/Y") V("OR2X1_LOC_785/B") V("OR2X1_LOC_493/Y") V("OR2X1_LOC_560/A") V("OR2X1_LOC_453/A") V("OR2X1_LOC_347/Y") V("OR2X1_LOC_486/Y") V("OR2X1_LOC_705/Y") V("OR2X1_LOC_124/Y") V("OR2X1_LOC_792/A") V("OR2X1_LOC_563/A") V("OR2X1_LOC_772/A") V("OR2X1_LOC_213/B") V("OR2X1_LOC_731/B") V("OR2X1_LOC_403/A") V("OR2X1_LOC_805/A") V("OR2X1_LOC_651/A") V("AND2X1_LOC_470/B") V("AND2X1_LOC_550/A") V("AND2X1_LOC_242/B") V("AND2X1_LOC_228/Y") V("AND2X1_LOC_349/B") V("AND2X1_LOC_728/Y") V("AND2X1_LOC_148/Y") V("AND2X1_LOC_794/B") V("AND2X1_LOC_661/A") V("AND2X1_LOC_734/Y") V("AND2X1_LOC_475/Y") V("AND2X1_LOC_192/Y") V("AND2X1_LOC_842/B") V("AND2X1_LOC_326/A") V("AND2X1_LOC_722/A") V("AND2X1_LOC_703/Y") V("AND2X1_LOC_388/Y") V("OR2X1_LOC_555/B") V("OR2X1_LOC_649/B") V("OR2X1_LOC_553/B") V("OR2X1_LOC_181/Y") V("OR2X1_LOC_781/Y") V("OR2X1_LOC_833/Y") V("OR2X1_LOC_500/A") V("OR2X1_LOC_194/Y") V("OR2X1_LOC_326/B") V("OR2X1_LOC_648/B") V("OR2X1_LOC_647/A") V("OR2X1_LOC_719/Y") V("OR2X1_LOC_204/Y") V("OR2X1_LOC_812/B") V("OR2X1_LOC_575/A") V("OR2X1_LOC_366/B") V("OR2X1_LOC_476/Y") V("AND2X1_LOC_656/Y") V("AND2X1_LOC_216/Y") V("AND2X1_LOC_345/Y") V("AND2X1_LOC_727/B") V("AND2X1_LOC_554/B") V("OR2X1_LOC_561/Y") V("AND2X1_LOC_553/A") V("AND2X1_LOC_191/B") V("AND2X1_LOC_639/B") V("AND2X1_LOC_193/Y") V("AND2X1_LOC_449/Y") V("OR2X1_LOC_348/Y") V("AND2X1_LOC_793/Y") V("OR2X1_LOC_728/B") V("OR2X1_LOC_551/A") V("OR2X1_LOC_228/Y") V("OR2X1_LOC_797/A") V("OR2X1_LOC_523/Y") V("OR2X1_LOC_639/A") V("OR2X1_LOC_552/B") V("OR2X1_LOC_792/Y") V("OR2X1_LOC_711/A") V("AND2X1_LOC_852/B") V("AND2X1_LOC_243/Y") V("AND2X1_LOC_476/A") V("OR2X1_LOC_739/A") V("OR2X1_LOC_863/B") V("OR2X1_LOC_565/A") V("OR2X1_LOC_339/Y") V("OR2X1_LOC_724/A") V("AND2X1_LOC_574/Y") V("OR2X1_LOC_787/Y") V("OR2X1_LOC_772/Y") V("OR2X1_LOC_714/Y") V("OR2X1_LOC_340/Y") V("OR2X1_LOC_679/Y") V("AND2X1_LOC_772/B") V("AND2X1_LOC_139/A") V("AND2X1_LOC_792/Y") V("AND2X1_LOC_474/A") V("AND2X1_LOC_403/B") V("OR2X1_LOC_862/A") V("OR2X1_LOC_508/A") V("OR2X1_LOC_550/B") V("OR2X1_LOC_720/Y") V("OR2X1_LOC_602/Y") V("AND2X1_LOC_850/Y") V("OR2X1_LOC_359/A") V("AND2X1_LOC_244/A") V("AND2X1_LOC_771/B") V("AND2X1_LOC_785/A") V("OR2X1_LOC_647/Y") V("AND2X1_LOC_552/A") V("AND2X1_LOC_337/B") V("AND2X1_LOC_202/Y") V("AND2X1_LOC_620/Y") V("AND2X1_LOC_181/Y") V("AND2X1_LOC_141/A") V("AND2X1_LOC_852/Y") V("AND2X1_LOC_568/B") V("AND2X1_LOC_856/A") V("AND2X1_LOC_571/B") V("OR2X1_LOC_241/Y") V("OR2X1_LOC_715/A") V("OR2X1_LOC_401/Y") V("OR2X1_LOC_345/Y") V("AND2X1_LOC_348/Y") V("OR2X1_LOC_641/B") V("OR2X1_LOC_620/Y") V("AND2X1_LOC_453/Y") V("AND2X1_LOC_658/B") V("OR2X1_LOC_796/B") V("OR2X1_LOC_851/B") V("AND2X1_LOC_555/Y") V("OR2X1_LOC_654/A") V("OR2X1_LOC_472/A") V("OR2X1_LOC_723/A") V("OR2X1_LOC_795/B") V("OR2X1_LOC_170/Y") V("OR2X1_LOC_797/B") V("OR2X1_LOC_357/A") V("OR2X1_LOC_731/A") V("OR2X1_LOC_725/B") V("OR2X1_LOC_851/A") V("AND2X1_LOC_564/B") V("AND2X1_LOC_794/A") V("AND2X1_LOC_566/B") V("AND2X1_LOC_716/Y") V("OR2X1_LOC_471/Y") V("AND2X1_LOC_201/Y") V("AND2X1_LOC_786/Y") V("OR2X1_LOC_352/A") V("OR2X1_LOC_214/A") V("AND2X1_LOC_721/Y") V("OR2X1_LOC_624/Y") V("AND2X1_LOC_640/Y") V("AND2X1_LOC_563/A") V("AND2X1_LOC_784/Y") V("AND2X1_LOC_211/B") V("AND2X1_LOC_347/B") V("AND2X1_LOC_850/A") V("AND2X1_LOC_203/Y") V("AND2X1_LOC_208/Y") V("AND2X1_LOC_352/B") V("OR2X1_LOC_725/A") V("OR2X1_LOC_726/A") V("AND2X1_LOC_565/Y") V("AND2X1_LOC_523/Y") V("AND2X1_LOC_61/Y") V("AND2X1_LOC_624/B") V("AND2X1_LOC_500/Y") V("AND2X1_LOC_401/Y") V("AND2X1_LOC_840/A") V("AND2X1_LOC_500/B") V("AND2X1_LOC_486/Y") V("AND2X1_LOC_649/B") V("AND2X1_LOC_84/Y") V("OR2X1_LOC_365/B") V("OR2X1_LOC_453/Y") V("OR2X1_LOC_475/Y") V("OR2X1_LOC_737/A") V("OR2X1_LOC_140/B") V("OR2X1_LOC_137/Y") V("OR2X1_LOC_739/B") V("OR2X1_LOC_850/B") V("OR2X1_LOC_190/Y") V("OR2X1_LOC_794/A") V("OR2X1_LOC_653/Y") V("OR2X1_LOC_605/Y") V("OR2X1_LOC_561/A") V("OR2X1_LOC_193/Y") V("OR2X1_LOC_140/Y") V("OR2X1_LOC_770/Y") V("OR2X1_LOC_468/A") V("OR2X1_LOC_347/A") V("OR2X1_LOC_842/A") V("OR2X1_LOC_61/Y") V("OR2X1_LOC_84/Y") V("AND2X1_LOC_141/B") V("AND2X1_LOC_231/Y") V("AND2X1_LOC_561/B") V("AND2X1_LOC_792/B") V("AND2X1_LOC_710/Y") V("AND2X1_LOC_647/B") V("AND2X1_LOC_468/B") V("AND2X1_LOC_717/B") V("AND2X1_LOC_702/Y") V("AND2X1_LOC_204/Y") V("AND2X1_LOC_705/Y") V("AND2X1_LOC_645/A") V("AND2X1_LOC_347/Y") V("AND2X1_LOC_572/A") V("AND2X1_LOC_209/Y") V("AND2X1_LOC_726/Y") V("AND2X1_LOC_797/B") V("AND2X1_LOC_554/Y") V("OR2X1_LOC_440/A") V("OR2X1_LOC_551/B") V("OR2X1_LOC_735/B") V("OR2X1_LOC_675/Y") V("OR2X1_LOC_124/A") V("OR2X1_LOC_835/Y") V("OR2X1_LOC_182/B") V("OR2X1_LOC_175/Y") V("OR2X1_LOC_203/Y") V("OR2X1_LOC_174/Y") V("OR2X1_LOC_641/Y") V("OR2X1_LOC_786/Y") V("OR2X1_LOC_469/B") V("OR2X1_LOC_170/A") V("OR2X1_LOC_192/A") V("OR2X1_LOC_562/B") V("OR2X1_LOC_722/B") V("OR2X1_LOC_703/Y") V("OR2X1_LOC_390/B") V("OR2X1_LOC_201/Y") V("OR2X1_LOC_337/A") V("OR2X1_LOC_624/A") V("OR2X1_LOC_501/A") V("OR2X1_LOC_643/Y") V("AND2X1_LOC_651/B") V("OR2X1_LOC_802/A") V("OR2X1_LOC_798/Y") V("AND2X1_LOC_798/Y") V("AND2X1_LOC_802/B") V("OR2X1_LOC_539/Y") V("AND2X1_LOC_539/Y") V("AND2X1_LOC_810/A") V("OR2X1_LOC_774/Y") V("OR2X1_LOC_510/Y") V("AND2X1_LOC_574/A") V("OR2X1_LOC_35/Y") V("AND2X1_LOC_35/Y") V("AND2X1_LOC_465/A") V("AND2X1_LOC_573/A") V("OR2X1_LOC_465/B") V("OR2X1_LOC_404/Y") V("OR2X1_LOC_799/A") V("AND2X1_LOC_361/A") V("AND2X1_LOC_483/Y") V("AND2X1_LOC_436/Y") V("OR2X1_LOC_631/B") V("OR2X1_LOC_436/Y") V("OR2X1_LOC_319/Y") V("AND2X1_LOC_593/Y") V("OR2X1_LOC_267/Y") V("AND2X1_LOC_798/A") 

* SUBCKT HEAD: NAME;  INPUTS; POWER; OUTPUTS
.subckt AES_SBOX_3
+ OR2X1_LOC_351/B OR2X1_LOC_852/A OR2X1_LOC_244/A OR2X1_LOC_476/B AND2X1_LOC_810/Y AND2X1_LOC_476/Y AND2X1_LOC_366/A OR2X1_LOC_656/Y OR2X1_LOC_216/Y AND2X1_LOC_863/A AND2X1_LOC_739/B AND2X1_LOC_565/B AND2X1_LOC_715/Y AND2X1_LOC_339/Y AND2X1_LOC_851/B AND2X1_LOC_796/A AND2X1_LOC_471/Y AND2X1_LOC_560/B AND2X1_LOC_642/Y AND2X1_LOC_207/A AND2X1_LOC_851/A AND2X1_LOC_720/Y AND2X1_LOC_359/B OR2X1_LOC_362/B OR2X1_LOC_858/B OR2X1_LOC_632/Y AND2X1_LOC_806/A AND2X1_LOC_772/Y AND2X1_LOC_338/Y AND2X1_LOC_454/Y AND2X1_LOC_724/A AND2X1_LOC_340/Y OR2X1_LOC_566/A OR2X1_LOC_723/B OR2X1_LOC_564/A OR2X1_LOC_467/A AND2X1_LOC_859/Y AND2X1_LOC_647/Y OR2X1_LOC_206/A OR2X1_LOC_856/B OR2X1_LOC_568/A OR2X1_LOC_207/B OR2X1_LOC_141/B OR2X1_LOC_857/B OR2X1_LOC_466/A OR2X1_LOC_392/B AND2X1_LOC_797/A AND2X1_LOC_357/B AND2X1_LOC_727/Y AND2X1_LOC_712/Y AND2X1_LOC_654/B 
+ AND2X1_LOC_472/B AND2X1_LOC_717/Y AND2X1_LOC_170/Y AND2X1_LOC_785/Y OR2X1_LOC_721/Y AND2X1_LOC_713/Y AND2X1_LOC_711/Y AND2X1_LOC_658/A OR2X1_LOC_640/Y OR2X1_LOC_563/B OR2X1_LOC_784/Y OR2X1_LOC_569/A OR2X1_LOC_474/B AND2X1_LOC_392/A AND2X1_LOC_644/Y AND2X1_LOC_365/A AND2X1_LOC_508/B AND2X1_LOC_781/Y AND2X1_LOC_259/Y AND2X1_LOC_213/B AND2X1_LOC_544/Y AND2X1_LOC_675/A AND2X1_LOC_605/Y AND2X1_LOC_501/Y AND2X1_LOC_675/Y AND2X1_LOC_123/Y AND2X1_LOC_839/A AND2X1_LOC_182/A AND2X1_LOC_194/Y AND2X1_LOC_719/Y AND2X1_LOC_175/B AND2X1_LOC_641/Y AND2X1_LOC_551/B AND2X1_LOC_443/Y AND2X1_LOC_170/B AND2X1_LOC_191/Y AND2X1_LOC_452/Y OR2X1_LOC_244/B OR2X1_LOC_349/A OR2X1_LOC_730/B OR2X1_LOC_148/Y OR2X1_LOC_470/A OR2X1_LOC_213/A OR2X1_LOC_443/Y OR2X1_LOC_785/B OR2X1_LOC_493/Y OR2X1_LOC_560/A OR2X1_LOC_453/A OR2X1_LOC_347/Y OR2X1_LOC_486/Y OR2X1_LOC_705/Y 
+ OR2X1_LOC_124/Y OR2X1_LOC_792/A OR2X1_LOC_563/A OR2X1_LOC_772/A OR2X1_LOC_213/B OR2X1_LOC_731/B OR2X1_LOC_403/A OR2X1_LOC_805/A OR2X1_LOC_651/A AND2X1_LOC_470/B AND2X1_LOC_550/A AND2X1_LOC_242/B AND2X1_LOC_228/Y AND2X1_LOC_349/B AND2X1_LOC_728/Y AND2X1_LOC_148/Y AND2X1_LOC_794/B AND2X1_LOC_661/A AND2X1_LOC_734/Y AND2X1_LOC_475/Y AND2X1_LOC_192/Y AND2X1_LOC_842/B AND2X1_LOC_326/A AND2X1_LOC_722/A AND2X1_LOC_703/Y AND2X1_LOC_388/Y OR2X1_LOC_555/B OR2X1_LOC_649/B OR2X1_LOC_553/B OR2X1_LOC_181/Y OR2X1_LOC_781/Y OR2X1_LOC_833/Y OR2X1_LOC_500/A OR2X1_LOC_194/Y OR2X1_LOC_326/B OR2X1_LOC_648/B OR2X1_LOC_647/A OR2X1_LOC_719/Y OR2X1_LOC_204/Y OR2X1_LOC_812/B OR2X1_LOC_575/A OR2X1_LOC_366/B OR2X1_LOC_476/Y AND2X1_LOC_656/Y AND2X1_LOC_216/Y AND2X1_LOC_345/Y AND2X1_LOC_727/B AND2X1_LOC_554/B OR2X1_LOC_561/Y AND2X1_LOC_553/A AND2X1_LOC_191/B 
+ AND2X1_LOC_639/B AND2X1_LOC_193/Y AND2X1_LOC_449/Y OR2X1_LOC_348/Y AND2X1_LOC_793/Y OR2X1_LOC_728/B OR2X1_LOC_551/A OR2X1_LOC_228/Y OR2X1_LOC_797/A OR2X1_LOC_523/Y OR2X1_LOC_639/A OR2X1_LOC_552/B OR2X1_LOC_792/Y OR2X1_LOC_711/A AND2X1_LOC_852/B AND2X1_LOC_243/Y AND2X1_LOC_476/A OR2X1_LOC_739/A OR2X1_LOC_863/B OR2X1_LOC_565/A OR2X1_LOC_339/Y OR2X1_LOC_724/A AND2X1_LOC_574/Y OR2X1_LOC_787/Y OR2X1_LOC_772/Y OR2X1_LOC_714/Y OR2X1_LOC_340/Y OR2X1_LOC_679/Y AND2X1_LOC_772/B AND2X1_LOC_139/A AND2X1_LOC_792/Y AND2X1_LOC_474/A AND2X1_LOC_403/B OR2X1_LOC_862/A OR2X1_LOC_508/A OR2X1_LOC_550/B OR2X1_LOC_720/Y OR2X1_LOC_602/Y AND2X1_LOC_850/Y OR2X1_LOC_359/A AND2X1_LOC_244/A AND2X1_LOC_771/B AND2X1_LOC_785/A OR2X1_LOC_647/Y AND2X1_LOC_552/A AND2X1_LOC_337/B AND2X1_LOC_202/Y AND2X1_LOC_620/Y AND2X1_LOC_181/Y AND2X1_LOC_141/A AND2X1_LOC_852/Y 
+ AND2X1_LOC_568/B AND2X1_LOC_856/A AND2X1_LOC_571/B OR2X1_LOC_241/Y OR2X1_LOC_715/A OR2X1_LOC_401/Y OR2X1_LOC_345/Y AND2X1_LOC_348/Y OR2X1_LOC_641/B OR2X1_LOC_620/Y AND2X1_LOC_453/Y AND2X1_LOC_658/B OR2X1_LOC_796/B OR2X1_LOC_851/B AND2X1_LOC_555/Y OR2X1_LOC_654/A OR2X1_LOC_472/A OR2X1_LOC_723/A OR2X1_LOC_795/B OR2X1_LOC_170/Y OR2X1_LOC_797/B OR2X1_LOC_357/A OR2X1_LOC_731/A OR2X1_LOC_725/B OR2X1_LOC_851/A AND2X1_LOC_564/B AND2X1_LOC_794/A AND2X1_LOC_566/B AND2X1_LOC_716/Y OR2X1_LOC_471/Y AND2X1_LOC_201/Y AND2X1_LOC_786/Y OR2X1_LOC_352/A OR2X1_LOC_214/A AND2X1_LOC_721/Y OR2X1_LOC_624/Y AND2X1_LOC_640/Y AND2X1_LOC_563/A AND2X1_LOC_784/Y AND2X1_LOC_211/B AND2X1_LOC_347/B AND2X1_LOC_850/A AND2X1_LOC_203/Y AND2X1_LOC_208/Y AND2X1_LOC_352/B OR2X1_LOC_725/A OR2X1_LOC_726/A AND2X1_LOC_565/Y AND2X1_LOC_523/Y AND2X1_LOC_61/Y AND2X1_LOC_624/B 
+ AND2X1_LOC_500/Y AND2X1_LOC_401/Y AND2X1_LOC_840/A AND2X1_LOC_500/B AND2X1_LOC_486/Y AND2X1_LOC_649/B AND2X1_LOC_84/Y OR2X1_LOC_365/B OR2X1_LOC_453/Y OR2X1_LOC_475/Y OR2X1_LOC_737/A OR2X1_LOC_140/B OR2X1_LOC_137/Y OR2X1_LOC_739/B OR2X1_LOC_850/B OR2X1_LOC_190/Y OR2X1_LOC_794/A OR2X1_LOC_653/Y OR2X1_LOC_605/Y OR2X1_LOC_561/A OR2X1_LOC_193/Y OR2X1_LOC_140/Y OR2X1_LOC_770/Y OR2X1_LOC_468/A OR2X1_LOC_347/A OR2X1_LOC_842/A OR2X1_LOC_61/Y OR2X1_LOC_84/Y AND2X1_LOC_141/B AND2X1_LOC_231/Y AND2X1_LOC_561/B AND2X1_LOC_792/B AND2X1_LOC_710/Y AND2X1_LOC_647/B AND2X1_LOC_468/B AND2X1_LOC_717/B AND2X1_LOC_702/Y AND2X1_LOC_204/Y AND2X1_LOC_705/Y AND2X1_LOC_645/A AND2X1_LOC_347/Y AND2X1_LOC_572/A AND2X1_LOC_209/Y AND2X1_LOC_726/Y AND2X1_LOC_797/B AND2X1_LOC_554/Y OR2X1_LOC_440/A OR2X1_LOC_551/B OR2X1_LOC_735/B OR2X1_LOC_675/Y OR2X1_LOC_124/A 
+ OR2X1_LOC_835/Y OR2X1_LOC_182/B OR2X1_LOC_175/Y OR2X1_LOC_203/Y OR2X1_LOC_174/Y OR2X1_LOC_641/Y OR2X1_LOC_786/Y OR2X1_LOC_469/B OR2X1_LOC_170/A OR2X1_LOC_192/A OR2X1_LOC_562/B OR2X1_LOC_722/B OR2X1_LOC_703/Y OR2X1_LOC_390/B OR2X1_LOC_201/Y OR2X1_LOC_337/A OR2X1_LOC_624/A OR2X1_LOC_501/A OR2X1_LOC_643/Y AND2X1_LOC_651/B OR2X1_LOC_802/A OR2X1_LOC_798/Y AND2X1_LOC_798/Y AND2X1_LOC_802/B OR2X1_LOC_539/Y AND2X1_LOC_539/Y AND2X1_LOC_810/A OR2X1_LOC_774/Y OR2X1_LOC_510/Y AND2X1_LOC_574/A OR2X1_LOC_35/Y AND2X1_LOC_35/Y AND2X1_LOC_465/A AND2X1_LOC_573/A OR2X1_LOC_465/B OR2X1_LOC_404/Y OR2X1_LOC_799/A AND2X1_LOC_361/A AND2X1_LOC_483/Y AND2X1_LOC_436/Y OR2X1_LOC_631/B OR2X1_LOC_436/Y OR2X1_LOC_319/Y AND2X1_LOC_593/Y OR2X1_LOC_267/Y AND2X1_LOC_798/A 
+ VSS VDD 
+ GATE_222 GATE_366 GATE_479 GATE_579 GATE_662 GATE_741 GATE_811 GATE_865 D_GATE_222 D_GATE_366 D_GATE_479 D_GATE_579 D_GATE_662 D_GATE_741 D_GATE_811 D_GATE_865 

* NETLIST 
XOR2X1_LOC_649 OR2X1_LOC_649/a_8_216# OR2X1_LOC_649/a_36_216# OR2X1_LOC_655/A VSS VDD OR2X1_LOC_643/Y OR2X1_LOC_649/B OR2X1_LOC

XOR2X1_LOC_206 OR2X1_LOC_206/a_8_216# OR2X1_LOC_206/a_36_216# OR2X1_LOC_215/A VSS VDD OR2X1_LOC_206/A OR2X1_LOC_201/Y OR2X1_LOC

XOR2X1_LOC_722 OR2X1_LOC_722/a_8_216# OR2X1_LOC_722/a_36_216# OR2X1_LOC_733/B VSS VDD OR2X1_LOC_719/Y OR2X1_LOC_722/B OR2X1_LOC

XOR2X1_LOC_562 OR2X1_LOC_562/a_8_216# OR2X1_LOC_562/a_36_216# OR2X1_LOC_562/Y VSS VDD OR2X1_LOC_562/A OR2X1_LOC_562/B OR2X1_LOC

XOR2X1_LOC_469 OR2X1_LOC_469/a_8_216# OR2X1_LOC_469/a_36_216# OR2X1_LOC_469/Y VSS VDD OR2X1_LOC_468/Y OR2X1_LOC_469/B OR2X1_LOC

XOR2X1_LOC_795 OR2X1_LOC_795/a_8_216# OR2X1_LOC_795/a_36_216# OR2X1_LOC_804/A VSS VDD OR2X1_LOC_786/Y OR2X1_LOC_795/B OR2X1_LOC

XOR2X1_LOC_650 OR2X1_LOC_650/a_8_216# OR2X1_LOC_650/a_36_216# OR2X1_LOC_650/Y VSS VDD OR2X1_LOC_641/Y OR2X1_LOC_640/Y OR2X1_LOC

XOR2X1_LOC_205 OR2X1_LOC_205/a_8_216# OR2X1_LOC_205/a_36_216# OR2X1_LOC_205/Y VSS VDD OR2X1_LOC_204/Y OR2X1_LOC_203/Y OR2X1_LOC

XOR2X1_LOC_853 OR2X1_LOC_853/a_8_216# OR2X1_LOC_853/a_36_216# OR2X1_LOC_857/A VSS VDD OR2X1_LOC_175/Y OR2X1_LOC_35/Y OR2X1_LOC

XOR2X1_LOC_211 OR2X1_LOC_211/a_8_216# OR2X1_LOC_211/a_36_216# OR2X1_LOC_212/A VSS VDD OR2X1_LOC_175/Y OR2X1_LOC_170/Y OR2X1_LOC

XOR2X1_LOC_182 OR2X1_LOC_182/a_8_216# OR2X1_LOC_182/a_36_216# OR2X1_LOC_212/B VSS VDD OR2X1_LOC_181/Y OR2X1_LOC_182/B OR2X1_LOC

XOR2X1_LOC_806 OR2X1_LOC_806/a_8_216# OR2X1_LOC_806/a_36_216# OR2X1_LOC_807/A VSS VDD OR2X1_LOC_675/Y OR2X1_LOC_362/B OR2X1_LOC

XOR2X1_LOC_736 OR2X1_LOC_736/a_8_216# OR2X1_LOC_736/a_36_216# OR2X1_LOC_736/Y VSS VDD OR2X1_LOC_736/A OR2X1_LOC_675/Y OR2X1_LOC

XOR2X1_LOC_573 OR2X1_LOC_573/a_8_216# OR2X1_LOC_573/a_36_216# OR2X1_LOC_573/Y VSS VDD OR2X1_LOC_735/B OR2X1_LOC_404/Y OR2X1_LOC

XOR2X1_LOC_735 OR2X1_LOC_735/a_8_216# OR2X1_LOC_735/a_36_216# OR2X1_LOC_736/A VSS VDD OR2X1_LOC_632/Y OR2X1_LOC_735/B OR2X1_LOC

XOR2X1_LOC_551 OR2X1_LOC_551/a_8_216# OR2X1_LOC_551/a_36_216# OR2X1_LOC_564/B VSS VDD OR2X1_LOC_551/A OR2X1_LOC_551/B OR2X1_LOC

XAND2X1_LOC_563 AND2X1_LOC_563/a_36_24# AND2X1_LOC_563/Y AND2X1_LOC_563/a_8_24# VSS VDD AND2X1_LOC_563/A AND2X1_LOC_554/Y AND2X1_LOC

XAND2X1_LOC_797 AND2X1_LOC_797/a_36_24# AND2X1_LOC_803/B AND2X1_LOC_797/a_8_24# VSS VDD AND2X1_LOC_797/A AND2X1_LOC_797/B AND2X1_LOC

XAND2X1_LOC_731 AND2X1_LOC_731/a_36_24# AND2X1_LOC_731/Y AND2X1_LOC_731/a_8_24# VSS VDD AND2X1_LOC_726/Y AND2X1_LOC_727/Y AND2X1_LOC

XAND2X1_LOC_213 AND2X1_LOC_213/a_36_24# AND2X1_LOC_220/B AND2X1_LOC_213/a_8_24# VSS VDD AND2X1_LOC_209/Y AND2X1_LOC_213/B AND2X1_LOC

XAND2X1_LOC_572 AND2X1_LOC_572/a_36_24# AND2X1_LOC_572/Y AND2X1_LOC_572/a_8_24# VSS VDD AND2X1_LOC_572/A AND2X1_LOC_361/A AND2X1_LOC

XAND2X1_LOC_217 AND2X1_LOC_217/a_36_24# AND2X1_LOC_217/Y AND2X1_LOC_217/a_8_24# VSS VDD AND2X1_LOC_572/A AND2X1_LOC_657/A AND2X1_LOC

XAND2X1_LOC_360 AND2X1_LOC_360/a_36_24# AND2X1_LOC_363/B AND2X1_LOC_360/a_8_24# VSS VDD AND2X1_LOC_860/A AND2X1_LOC_347/Y AND2X1_LOC

XAND2X1_LOC_645 AND2X1_LOC_645/a_36_24# AND2X1_LOC_648/B AND2X1_LOC_645/a_8_24# VSS VDD AND2X1_LOC_645/A AND2X1_LOC_605/Y AND2X1_LOC

XAND2X1_LOC_205 AND2X1_LOC_205/a_36_24# AND2X1_LOC_215/A AND2X1_LOC_205/a_8_24# VSS VDD AND2X1_LOC_203/Y AND2X1_LOC_204/Y AND2X1_LOC

XAND2X1_LOC_556 AND2X1_LOC_556/a_36_24# AND2X1_LOC_562/B AND2X1_LOC_556/a_8_24# VSS VDD AND2X1_LOC_483/Y AND2X1_LOC_486/Y AND2X1_LOC

XAND2X1_LOC_468 AND2X1_LOC_468/a_36_24# AND2X1_LOC_469/B AND2X1_LOC_468/a_8_24# VSS VDD AND2X1_LOC_436/Y AND2X1_LOC_468/B AND2X1_LOC

XAND2X1_LOC_341 AND2X1_LOC_341/a_36_24# AND2X1_LOC_350/B AND2X1_LOC_341/a_8_24# VSS VDD AND2X1_LOC_228/Y AND2X1_LOC_231/Y AND2X1_LOC

XAND2X1_LOC_141 AND2X1_LOC_141/a_36_24# AND2X1_LOC_657/A AND2X1_LOC_141/a_8_24# VSS VDD AND2X1_LOC_141/A AND2X1_LOC_141/B AND2X1_LOC

XOR2X1_LOC_556 OR2X1_LOC_556/a_8_216# OR2X1_LOC_556/a_36_216# OR2X1_LOC_562/A VSS VDD OR2X1_LOC_486/Y OR2X1_LOC_631/B OR2X1_LOC

XOR2X1_LOC_468 OR2X1_LOC_468/a_8_216# OR2X1_LOC_468/a_36_216# OR2X1_LOC_468/Y VSS VDD OR2X1_LOC_468/A OR2X1_LOC_436/Y OR2X1_LOC

XOR2X1_LOC_141 OR2X1_LOC_141/a_8_216# OR2X1_LOC_141/a_36_216# OR2X1_LOC_217/A VSS VDD OR2X1_LOC_140/Y OR2X1_LOC_141/B OR2X1_LOC

XOR2X1_LOC_200 OR2X1_LOC_200/a_8_216# OR2X1_LOC_200/a_36_216# OR2X1_LOC_200/Y VSS VDD OR2X1_LOC_194/Y OR2X1_LOC_193/Y OR2X1_LOC

XOR2X1_LOC_645 OR2X1_LOC_645/a_8_216# OR2X1_LOC_645/a_36_216# OR2X1_LOC_648/A VSS VDD OR2X1_LOC_605/Y OR2X1_LOC_602/Y OR2X1_LOC

XOR2X1_LOC_661 OR2X1_LOC_661/a_8_216# OR2X1_LOC_661/a_36_216# OR2X1_LOC_662/A VSS VDD OR2X1_LOC_661/A OR2X1_LOC_653/Y OR2X1_LOC

XOR2X1_LOC_794 OR2X1_LOC_794/a_8_216# OR2X1_LOC_794/a_36_216# OR2X1_LOC_804/B VSS VDD OR2X1_LOC_794/A OR2X1_LOC_787/Y OR2X1_LOC

XOR2X1_LOC_221 OR2X1_LOC_221/a_8_216# OR2X1_LOC_221/a_36_216# OR2X1_LOC_223/B VSS VDD OR2X1_LOC_221/A OR2X1_LOC_739/B OR2X1_LOC

XOR2X1_LOC_739 OR2X1_LOC_739/a_8_216# OR2X1_LOC_739/a_36_216# OR2X1_LOC_739/Y VSS VDD OR2X1_LOC_739/A OR2X1_LOC_739/B OR2X1_LOC

XOR2X1_LOC_737 OR2X1_LOC_737/a_8_216# OR2X1_LOC_737/a_36_216# OR2X1_LOC_741/A VSS VDD OR2X1_LOC_737/A OR2X1_LOC_733/Y OR2X1_LOC

XOR2X1_LOC_479 OR2X1_LOC_479/a_8_216# OR2X1_LOC_479/a_36_216# OR2X1_LOC_479/Y VSS VDD OR2X1_LOC_476/Y OR2X1_LOC_475/Y OR2X1_LOC

XOR2X1_LOC_466 OR2X1_LOC_466/a_8_216# OR2X1_LOC_466/a_36_216# OR2X1_LOC_470/B VSS VDD OR2X1_LOC_466/A OR2X1_LOC_453/Y OR2X1_LOC

XOR2X1_LOC_365 OR2X1_LOC_365/a_8_216# OR2X1_LOC_365/a_36_216# OR2X1_LOC_367/B VSS VDD OR2X1_LOC_364/Y OR2X1_LOC_365/B OR2X1_LOC

XAND2X1_LOC_649 AND2X1_LOC_649/a_36_24# AND2X1_LOC_649/Y AND2X1_LOC_649/a_8_24# VSS VDD AND2X1_LOC_642/Y AND2X1_LOC_649/B AND2X1_LOC

XAND2X1_LOC_560 AND2X1_LOC_560/a_36_24# AND2X1_LOC_571/A AND2X1_LOC_560/a_8_24# VSS VDD AND2X1_LOC_523/Y AND2X1_LOC_560/B AND2X1_LOC

XAND2X1_LOC_569 AND2X1_LOC_569/a_36_24# AND2X1_LOC_577/A AND2X1_LOC_569/a_8_24# VSS VDD AND2X1_LOC_569/A AND2X1_LOC_565/Y AND2X1_LOC

XOR2X1_LOC_725 OR2X1_LOC_725/a_8_216# OR2X1_LOC_725/a_36_216# OR2X1_LOC_732/A VSS VDD OR2X1_LOC_725/A OR2X1_LOC_725/B OR2X1_LOC

XAND2X1_LOC_352 AND2X1_LOC_352/a_36_24# AND2X1_LOC_357/A AND2X1_LOC_352/a_8_24# VSS VDD AND2X1_LOC_212/A AND2X1_LOC_352/B AND2X1_LOC

XAND2X1_LOC_214 AND2X1_LOC_214/a_36_24# AND2X1_LOC_219/A AND2X1_LOC_214/a_8_24# VSS VDD AND2X1_LOC_214/A AND2X1_LOC_208/Y AND2X1_LOC

XAND2X1_LOC_853 AND2X1_LOC_853/a_36_24# AND2X1_LOC_853/Y AND2X1_LOC_853/a_8_24# VSS VDD AND2X1_LOC_35/Y AND2X1_LOC_211/B AND2X1_LOC

XAND2X1_LOC_211 AND2X1_LOC_211/a_36_24# AND2X1_LOC_212/B AND2X1_LOC_211/a_8_24# VSS VDD AND2X1_LOC_170/Y AND2X1_LOC_211/B AND2X1_LOC

XAND2X1_LOC_796 AND2X1_LOC_796/a_36_24# AND2X1_LOC_796/Y AND2X1_LOC_796/a_8_24# VSS VDD AND2X1_LOC_796/A AND2X1_LOC_784/Y AND2X1_LOC

XAND2X1_LOC_650 AND2X1_LOC_650/a_36_24# AND2X1_LOC_650/Y AND2X1_LOC_650/a_8_24# VSS VDD AND2X1_LOC_640/Y AND2X1_LOC_641/Y AND2X1_LOC

XOR2X1_LOC_861 OR2X1_LOC_861/a_8_216# OR2X1_LOC_861/a_36_216# OR2X1_LOC_865/B VSS VDD OR2X1_LOC_860/Y OR2X1_LOC_624/Y OR2X1_LOC

XOR2X1_LOC_658 OR2X1_LOC_658/a_8_216# OR2X1_LOC_658/a_36_216# OR2X1_LOC_659/A VSS VDD OR2X1_LOC_632/Y OR2X1_LOC_624/Y OR2X1_LOC

XOR2X1_LOC_214 OR2X1_LOC_214/a_8_216# OR2X1_LOC_214/a_36_216# OR2X1_LOC_219/B VSS VDD OR2X1_LOC_214/A OR2X1_LOC_214/B OR2X1_LOC

XOR2X1_LOC_352 OR2X1_LOC_352/a_8_216# OR2X1_LOC_352/a_36_216# OR2X1_LOC_357/B VSS VDD OR2X1_LOC_352/A OR2X1_LOC_212/B OR2X1_LOC

XAND2X1_LOC_795 AND2X1_LOC_795/a_36_24# AND2X1_LOC_795/Y AND2X1_LOC_795/a_8_24# VSS VDD AND2X1_LOC_785/Y AND2X1_LOC_786/Y AND2X1_LOC

XAND2X1_LOC_206 AND2X1_LOC_206/a_36_24# AND2X1_LOC_206/Y AND2X1_LOC_206/a_8_24# VSS VDD AND2X1_LOC_201/Y AND2X1_LOC_202/Y AND2X1_LOC

XOR2X1_LOC_477 OR2X1_LOC_477/a_8_216# OR2X1_LOC_477/a_36_216# OR2X1_LOC_477/Y VSS VDD OR2X1_LOC_471/Y OR2X1_LOC_477/B OR2X1_LOC

XAND2X1_LOC_723 AND2X1_LOC_723/a_36_24# AND2X1_LOC_723/Y AND2X1_LOC_723/a_8_24# VSS VDD AND2X1_LOC_716/Y AND2X1_LOC_717/Y AND2X1_LOC

XAND2X1_LOC_566 AND2X1_LOC_566/a_36_24# AND2X1_LOC_566/Y AND2X1_LOC_566/a_8_24# VSS VDD AND2X1_LOC_170/Y AND2X1_LOC_566/B AND2X1_LOC

XAND2X1_LOC_794 AND2X1_LOC_794/a_36_24# AND2X1_LOC_804/A AND2X1_LOC_794/a_8_24# VSS VDD AND2X1_LOC_794/A AND2X1_LOC_794/B AND2X1_LOC

XAND2X1_LOC_564 AND2X1_LOC_564/a_36_24# AND2X1_LOC_569/A AND2X1_LOC_564/a_8_24# VSS VDD AND2X1_LOC_564/A AND2X1_LOC_564/B AND2X1_LOC

XOR2X1_LOC_851 OR2X1_LOC_851/a_8_216# OR2X1_LOC_851/a_36_216# OR2X1_LOC_858/A VSS VDD OR2X1_LOC_851/A OR2X1_LOC_851/B OR2X1_LOC

XOR2X1_LOC_731 OR2X1_LOC_731/a_8_216# OR2X1_LOC_731/a_36_216# OR2X1_LOC_738/B VSS VDD OR2X1_LOC_731/A OR2X1_LOC_731/B OR2X1_LOC

XOR2X1_LOC_357 OR2X1_LOC_357/a_8_216# OR2X1_LOC_357/a_36_216# OR2X1_LOC_364/B VSS VDD OR2X1_LOC_357/A OR2X1_LOC_357/B OR2X1_LOC

XOR2X1_LOC_797 OR2X1_LOC_797/a_8_216# OR2X1_LOC_797/a_36_216# OR2X1_LOC_803/A VSS VDD OR2X1_LOC_797/A OR2X1_LOC_797/B OR2X1_LOC

XOR2X1_LOC_566 OR2X1_LOC_566/a_8_216# OR2X1_LOC_566/a_36_216# OR2X1_LOC_566/Y VSS VDD OR2X1_LOC_566/A OR2X1_LOC_170/Y OR2X1_LOC

XOR2X1_LOC_723 OR2X1_LOC_723/a_8_216# OR2X1_LOC_723/a_36_216# OR2X1_LOC_733/A VSS VDD OR2X1_LOC_723/A OR2X1_LOC_723/B OR2X1_LOC

XOR2X1_LOC_654 OR2X1_LOC_654/a_8_216# OR2X1_LOC_654/a_36_216# OR2X1_LOC_661/A VSS VDD OR2X1_LOC_654/A OR2X1_LOC_650/Y OR2X1_LOC

XAND2X1_LOC_562 AND2X1_LOC_562/a_36_24# AND2X1_LOC_562/Y AND2X1_LOC_562/a_8_24# VSS VDD AND2X1_LOC_555/Y AND2X1_LOC_562/B AND2X1_LOC

XOR2X1_LOC_796 OR2X1_LOC_796/a_8_216# OR2X1_LOC_796/a_36_216# OR2X1_LOC_803/B VSS VDD OR2X1_LOC_784/Y OR2X1_LOC_796/B OR2X1_LOC

XAND2X1_LOC_735 AND2X1_LOC_735/a_36_24# AND2X1_LOC_735/Y AND2X1_LOC_735/a_8_24# VSS VDD AND2X1_LOC_501/Y AND2X1_LOC_658/B AND2X1_LOC

XAND2X1_LOC_658 AND2X1_LOC_658/a_36_24# AND2X1_LOC_658/Y AND2X1_LOC_658/a_8_24# VSS VDD AND2X1_LOC_658/A AND2X1_LOC_658/B AND2X1_LOC

XAND2X1_LOC_466 AND2X1_LOC_466/a_36_24# AND2X1_LOC_470/A AND2X1_LOC_466/a_8_24# VSS VDD AND2X1_LOC_453/Y AND2X1_LOC_454/Y AND2X1_LOC

XOR2X1_LOC_341 OR2X1_LOC_341/a_8_216# OR2X1_LOC_341/a_36_216# OR2X1_LOC_341/Y VSS VDD OR2X1_LOC_641/B OR2X1_LOC_228/Y OR2X1_LOC

XAND2X1_LOC_359 AND2X1_LOC_359/a_36_24# AND2X1_LOC_363/A AND2X1_LOC_359/a_8_24# VSS VDD AND2X1_LOC_348/Y AND2X1_LOC_359/B AND2X1_LOC

XAND2X1_LOC_571 AND2X1_LOC_571/a_36_24# AND2X1_LOC_571/Y AND2X1_LOC_571/a_8_24# VSS VDD AND2X1_LOC_571/A AND2X1_LOC_571/B AND2X1_LOC

XAND2X1_LOC_568 AND2X1_LOC_568/a_36_24# AND2X1_LOC_578/A AND2X1_LOC_568/a_8_24# VSS VDD AND2X1_LOC_566/Y AND2X1_LOC_568/B AND2X1_LOC

XAND2X1_LOC_857 AND2X1_LOC_857/a_36_24# AND2X1_LOC_857/Y AND2X1_LOC_857/a_8_24# VSS VDD AND2X1_LOC_852/Y AND2X1_LOC_853/Y AND2X1_LOC

XAND2X1_LOC_182 AND2X1_LOC_182/a_36_24# AND2X1_LOC_212/A AND2X1_LOC_182/a_8_24# VSS VDD AND2X1_LOC_182/A AND2X1_LOC_181/Y AND2X1_LOC

XAND2X1_LOC_244 AND2X1_LOC_244/a_36_24# AND2X1_LOC_860/A AND2X1_LOC_244/a_8_24# VSS VDD AND2X1_LOC_244/A AND2X1_LOC_243/Y AND2X1_LOC

XOR2X1_LOC_359 OR2X1_LOC_359/a_8_216# OR2X1_LOC_359/a_36_216# OR2X1_LOC_363/B VSS VDD OR2X1_LOC_359/A OR2X1_LOC_348/Y OR2X1_LOC

XAND2X1_LOC_858 AND2X1_LOC_858/a_36_24# AND2X1_LOC_862/A AND2X1_LOC_858/a_8_24# VSS VDD AND2X1_LOC_850/Y AND2X1_LOC_858/B AND2X1_LOC

XOR2X1_LOC_862 OR2X1_LOC_862/a_8_216# OR2X1_LOC_862/a_36_216# OR2X1_LOC_865/A VSS VDD OR2X1_LOC_862/A OR2X1_LOC_862/B OR2X1_LOC

XAND2X1_LOC_860 AND2X1_LOC_860/a_36_24# AND2X1_LOC_861/B AND2X1_LOC_860/a_8_24# VSS VDD AND2X1_LOC_860/A AND2X1_LOC_474/A AND2X1_LOC

XAND2X1_LOC_805 AND2X1_LOC_805/a_36_24# AND2X1_LOC_805/Y AND2X1_LOC_805/a_8_24# VSS VDD AND2X1_LOC_792/Y AND2X1_LOC_793/Y AND2X1_LOC

XOR2X1_LOC_350 OR2X1_LOC_350/a_8_216# OR2X1_LOC_350/a_36_216# OR2X1_LOC_358/B VSS VDD OR2X1_LOC_341/Y OR2X1_LOC_340/Y OR2X1_LOC

XOR2X1_LOC_724 OR2X1_LOC_724/a_8_216# OR2X1_LOC_724/a_36_216# OR2X1_LOC_732/B VSS VDD OR2X1_LOC_724/A OR2X1_LOC_714/Y OR2X1_LOC

XAND2X1_LOC_575 AND2X1_LOC_575/a_36_24# AND2X1_LOC_575/Y AND2X1_LOC_575/a_8_24# VSS VDD AND2X1_LOC_573/Y AND2X1_LOC_574/Y AND2X1_LOC

XOR2X1_LOC_351 OR2X1_LOC_351/a_8_216# OR2X1_LOC_351/a_36_216# OR2X1_LOC_358/A VSS VDD OR2X1_LOC_339/Y OR2X1_LOC_351/B OR2X1_LOC

XOR2X1_LOC_863 OR2X1_LOC_863/a_8_216# OR2X1_LOC_863/a_36_216# OR2X1_LOC_864/A VSS VDD OR2X1_LOC_863/A OR2X1_LOC_863/B OR2X1_LOC

XOR2X1_LOC_805 OR2X1_LOC_805/a_8_216# OR2X1_LOC_805/a_36_216# OR2X1_LOC_807/B VSS VDD OR2X1_LOC_805/A OR2X1_LOC_792/Y OR2X1_LOC

XOR2X1_LOC_560 OR2X1_LOC_560/a_8_216# OR2X1_LOC_560/a_36_216# OR2X1_LOC_571/B VSS VDD OR2X1_LOC_560/A OR2X1_LOC_523/Y OR2X1_LOC

XAND2X1_LOC_200 AND2X1_LOC_200/a_36_24# AND2X1_LOC_207/B AND2X1_LOC_200/a_8_24# VSS VDD AND2X1_LOC_193/Y AND2X1_LOC_194/Y AND2X1_LOC

XOR2X1_LOC_571 OR2X1_LOC_571/a_8_216# OR2X1_LOC_571/a_36_216# OR2X1_LOC_571/Y VSS VDD OR2X1_LOC_561/Y OR2X1_LOC_571/B OR2X1_LOC

XAND2X1_LOC_469 AND2X1_LOC_469/a_36_24# AND2X1_LOC_469/Y AND2X1_LOC_469/a_8_24# VSS VDD AND2X1_LOC_727/B AND2X1_LOC_469/B AND2X1_LOC

XAND2X1_LOC_218 AND2X1_LOC_218/a_36_24# AND2X1_LOC_218/Y AND2X1_LOC_218/a_8_24# VSS VDD AND2X1_LOC_216/Y AND2X1_LOC_217/Y AND2X1_LOC

XAND2X1_LOC_660 AND2X1_LOC_660/a_36_24# AND2X1_LOC_660/Y AND2X1_LOC_660/a_8_24# VSS VDD AND2X1_LOC_660/A AND2X1_LOC_656/Y AND2X1_LOC

XOR2X1_LOC_366 OR2X1_LOC_366/a_8_216# OR2X1_LOC_366/a_36_216# OR2X1_LOC_366/Y VSS VDD OR2X1_LOC_366/A OR2X1_LOC_366/B OR2X1_LOC

XOR2X1_LOC_575 OR2X1_LOC_575/a_8_216# OR2X1_LOC_575/a_36_216# OR2X1_LOC_579/B VSS VDD OR2X1_LOC_575/A OR2X1_LOC_573/Y OR2X1_LOC

XOR2X1_LOC_812 OR2X1_LOC_812/a_8_216# OR2X1_LOC_812/a_36_216# D_GATE_811 VSS VDD OR2X1_LOC_812/A OR2X1_LOC_812/B OR2X1_LOC

XOR2X1_LOC_648 OR2X1_LOC_648/a_8_216# OR2X1_LOC_648/a_36_216# OR2X1_LOC_655/B VSS VDD OR2X1_LOC_648/A OR2X1_LOC_648/B OR2X1_LOC

XAND2X1_LOC_722 AND2X1_LOC_722/a_36_24# AND2X1_LOC_722/Y AND2X1_LOC_722/a_8_24# VSS VDD AND2X1_LOC_722/A AND2X1_LOC_719/Y AND2X1_LOC

XAND2X1_LOC_739 AND2X1_LOC_739/a_36_24# AND2X1_LOC_740/B AND2X1_LOC_739/a_8_24# VSS VDD AND2X1_LOC_192/Y AND2X1_LOC_739/B AND2X1_LOC

XAND2X1_LOC_221 AND2X1_LOC_221/a_36_24# AND2X1_LOC_223/A AND2X1_LOC_221/a_8_24# VSS VDD AND2X1_LOC_192/Y AND2X1_LOC_220/Y AND2X1_LOC

XAND2X1_LOC_479 AND2X1_LOC_479/a_36_24# AND2X1_LOC_479/Y AND2X1_LOC_479/a_8_24# VSS VDD AND2X1_LOC_475/Y AND2X1_LOC_476/Y AND2X1_LOC

XAND2X1_LOC_737 AND2X1_LOC_737/a_36_24# AND2X1_LOC_737/Y AND2X1_LOC_737/a_8_24# VSS VDD AND2X1_LOC_733/Y AND2X1_LOC_734/Y AND2X1_LOC

XAND2X1_LOC_661 AND2X1_LOC_661/a_36_24# AND2X1_LOC_662/B AND2X1_LOC_661/a_8_24# VSS VDD AND2X1_LOC_661/A AND2X1_LOC_654/Y AND2X1_LOC

XAND2X1_LOC_470 AND2X1_LOC_470/a_36_24# AND2X1_LOC_477/A AND2X1_LOC_470/a_8_24# VSS VDD AND2X1_LOC_470/A AND2X1_LOC_470/B AND2X1_LOC

XOR2X1_LOC_213 OR2X1_LOC_213/a_8_216# OR2X1_LOC_213/a_36_216# OR2X1_LOC_220/A VSS VDD OR2X1_LOC_213/A OR2X1_LOC_213/B OR2X1_LOC

XOR2X1_LOC_563 OR2X1_LOC_563/a_8_216# OR2X1_LOC_563/a_36_216# OR2X1_LOC_570/A VSS VDD OR2X1_LOC_563/A OR2X1_LOC_563/B OR2X1_LOC

XOR2X1_LOC_217 OR2X1_LOC_217/a_8_216# OR2X1_LOC_217/a_36_216# OR2X1_LOC_217/Y VSS VDD OR2X1_LOC_217/A OR2X1_LOC_124/Y OR2X1_LOC

XOR2X1_LOC_572 OR2X1_LOC_572/a_8_216# OR2X1_LOC_572/a_36_216# OR2X1_LOC_576/A VSS VDD OR2X1_LOC_267/Y OR2X1_LOC_124/Y OR2X1_LOC

XOR2X1_LOC_360 OR2X1_LOC_360/a_8_216# OR2X1_LOC_360/a_36_216# OR2X1_LOC_363/A VSS VDD OR2X1_LOC_347/Y OR2X1_LOC_244/Y OR2X1_LOC

XOR2X1_LOC_470 OR2X1_LOC_470/a_8_216# OR2X1_LOC_470/a_36_216# OR2X1_LOC_477/B VSS VDD OR2X1_LOC_470/A OR2X1_LOC_470/B OR2X1_LOC

XOR2X1_LOC_244 OR2X1_LOC_244/a_8_216# OR2X1_LOC_244/a_36_216# OR2X1_LOC_244/Y VSS VDD OR2X1_LOC_244/A OR2X1_LOC_244/B OR2X1_LOC

XAND2X1_LOC_551 AND2X1_LOC_551/a_36_24# AND2X1_LOC_564/A AND2X1_LOC_551/a_8_24# VSS VDD AND2X1_LOC_544/Y AND2X1_LOC_551/B AND2X1_LOC

XAND2X1_LOC_736 AND2X1_LOC_736/a_36_24# AND2X1_LOC_736/Y AND2X1_LOC_736/a_8_24# VSS VDD AND2X1_LOC_675/Y AND2X1_LOC_735/Y AND2X1_LOC

XAND2X1_LOC_806 AND2X1_LOC_806/a_36_24# AND2X1_LOC_807/B AND2X1_LOC_806/a_8_24# VSS VDD AND2X1_LOC_806/A AND2X1_LOC_675/Y AND2X1_LOC

XAND2X1_LOC_573 AND2X1_LOC_573/a_36_24# AND2X1_LOC_573/Y AND2X1_LOC_573/a_8_24# VSS VDD AND2X1_LOC_573/A AND2X1_LOC_501/Y AND2X1_LOC

XAND2X1_LOC_365 AND2X1_LOC_365/a_36_24# AND2X1_LOC_367/A AND2X1_LOC_365/a_8_24# VSS VDD AND2X1_LOC_365/A AND2X1_LOC_364/Y AND2X1_LOC

XAND2X1_LOC_648 AND2X1_LOC_648/a_36_24# AND2X1_LOC_655/A AND2X1_LOC_648/a_8_24# VSS VDD AND2X1_LOC_644/Y AND2X1_LOC_648/B AND2X1_LOC

XOR2X1_LOC_860 OR2X1_LOC_860/a_8_216# OR2X1_LOC_860/a_36_216# OR2X1_LOC_860/Y VSS VDD OR2X1_LOC_474/B OR2X1_LOC_244/Y OR2X1_LOC

XOR2X1_LOC_569 OR2X1_LOC_569/a_8_216# OR2X1_LOC_569/a_36_216# OR2X1_LOC_577/B VSS VDD OR2X1_LOC_569/A OR2X1_LOC_569/B OR2X1_LOC

XAND2X1_LOC_861 AND2X1_LOC_861/a_36_24# AND2X1_LOC_865/A AND2X1_LOC_861/a_8_24# VSS VDD AND2X1_LOC_658/A AND2X1_LOC_861/B AND2X1_LOC

XAND2X1_LOC_725 AND2X1_LOC_725/a_36_24# AND2X1_LOC_732/B AND2X1_LOC_725/a_8_24# VSS VDD AND2X1_LOC_712/Y AND2X1_LOC_713/Y AND2X1_LOC

XAND2X1_LOC_654 AND2X1_LOC_654/a_36_24# AND2X1_LOC_654/Y AND2X1_LOC_654/a_8_24# VSS VDD AND2X1_LOC_650/Y AND2X1_LOC_654/B AND2X1_LOC

XAND2X1_LOC_357 AND2X1_LOC_357/a_36_24# AND2X1_LOC_364/A AND2X1_LOC_357/a_8_24# VSS VDD AND2X1_LOC_357/A AND2X1_LOC_357/B AND2X1_LOC

XOR2X1_LOC_857 OR2X1_LOC_857/a_8_216# OR2X1_LOC_857/a_36_216# OR2X1_LOC_863/A VSS VDD OR2X1_LOC_857/A OR2X1_LOC_857/B OR2X1_LOC

XOR2X1_LOC_207 OR2X1_LOC_207/a_8_216# OR2X1_LOC_207/a_36_216# OR2X1_LOC_214/B VSS VDD OR2X1_LOC_200/Y OR2X1_LOC_207/B OR2X1_LOC

XOR2X1_LOC_568 OR2X1_LOC_568/a_8_216# OR2X1_LOC_568/a_36_216# OR2X1_LOC_578/B VSS VDD OR2X1_LOC_568/A OR2X1_LOC_566/Y OR2X1_LOC

XAND2X1_LOC_862 AND2X1_LOC_862/a_36_24# AND2X1_LOC_862/Y AND2X1_LOC_862/a_8_24# VSS VDD AND2X1_LOC_862/A AND2X1_LOC_859/Y AND2X1_LOC

XOR2X1_LOC_564 OR2X1_LOC_564/a_8_216# OR2X1_LOC_564/a_36_216# OR2X1_LOC_569/B VSS VDD OR2X1_LOC_564/A OR2X1_LOC_564/B OR2X1_LOC

XAND2X1_LOC_350 AND2X1_LOC_350/a_36_24# AND2X1_LOC_350/Y AND2X1_LOC_350/a_8_24# VSS VDD AND2X1_LOC_340/Y AND2X1_LOC_350/B AND2X1_LOC

XAND2X1_LOC_724 AND2X1_LOC_724/a_36_24# AND2X1_LOC_724/Y AND2X1_LOC_724/a_8_24# VSS VDD AND2X1_LOC_724/A AND2X1_LOC_715/Y AND2X1_LOC

XAND2X1_LOC_351 AND2X1_LOC_351/a_36_24# AND2X1_LOC_351/Y AND2X1_LOC_351/a_8_24# VSS VDD AND2X1_LOC_338/Y AND2X1_LOC_339/Y AND2X1_LOC

XOR2X1_LOC_858 OR2X1_LOC_858/a_8_216# OR2X1_LOC_858/a_36_216# OR2X1_LOC_862/B VSS VDD OR2X1_LOC_858/A OR2X1_LOC_858/B OR2X1_LOC

XAND2X1_LOC_851 AND2X1_LOC_851/a_36_24# AND2X1_LOC_858/B AND2X1_LOC_851/a_8_24# VSS VDD AND2X1_LOC_851/A AND2X1_LOC_851/B AND2X1_LOC

XAND2X1_LOC_207 AND2X1_LOC_207/a_36_24# AND2X1_LOC_214/A AND2X1_LOC_207/a_8_24# VSS VDD AND2X1_LOC_207/A AND2X1_LOC_207/B AND2X1_LOC

XAND2X1_LOC_477 AND2X1_LOC_477/a_36_24# AND2X1_LOC_477/Y AND2X1_LOC_477/a_8_24# VSS VDD AND2X1_LOC_477/A AND2X1_LOC_471/Y AND2X1_LOC

XAND2X1_LOC_863 AND2X1_LOC_863/a_36_24# AND2X1_LOC_863/Y AND2X1_LOC_863/a_8_24# VSS VDD AND2X1_LOC_863/A AND2X1_LOC_857/Y AND2X1_LOC

XOR2X1_LOC_218 OR2X1_LOC_218/a_8_216# OR2X1_LOC_218/a_36_216# OR2X1_LOC_218/Y VSS VDD OR2X1_LOC_217/Y OR2X1_LOC_216/Y OR2X1_LOC

XOR2X1_LOC_660 OR2X1_LOC_660/a_8_216# OR2X1_LOC_660/a_36_216# OR2X1_LOC_660/Y VSS VDD OR2X1_LOC_656/Y OR2X1_LOC_660/B OR2X1_LOC

XAND2X1_LOC_366 AND2X1_LOC_366/a_36_24# AND2X1_LOC_367/B AND2X1_LOC_366/a_8_24# VSS VDD AND2X1_LOC_366/A AND2X1_LOC_363/Y AND2X1_LOC

XAND2X1_LOC_812 AND2X1_LOC_812/a_36_24# GATE_811 AND2X1_LOC_812/a_8_24# VSS VDD AND2X1_LOC_810/Y AND2X1_LOC_811/Y AND2X1_LOC

XAND2X1_LOC_367 AND2X1_LOC_367/a_36_24# GATE_366 AND2X1_LOC_367/a_8_24# VSS VDD AND2X1_LOC_367/A AND2X1_LOC_367/B AND2X1_LOC

XOR2X1_LOC_662 OR2X1_LOC_662/a_8_216# OR2X1_LOC_662/a_36_216# OR2X1_LOC_663/A VSS VDD OR2X1_LOC_662/A OR2X1_LOC_660/Y OR2X1_LOC

XOR2X1_LOC_222 OR2X1_LOC_222/a_8_216# OR2X1_LOC_222/a_36_216# OR2X1_LOC_223/A VSS VDD OR2X1_LOC_222/A OR2X1_LOC_218/Y OR2X1_LOC

XAND2X1_LOC_864 AND2X1_LOC_864/a_36_24# AND2X1_LOC_866/A AND2X1_LOC_864/a_8_24# VSS VDD AND2X1_LOC_810/A AND2X1_LOC_863/Y AND2X1_LOC

XAND2X1_LOC_478 AND2X1_LOC_478/a_36_24# AND2X1_LOC_480/A AND2X1_LOC_478/a_8_24# VSS VDD AND2X1_LOC_469/Y AND2X1_LOC_477/Y AND2X1_LOC

XAND2X1_LOC_358 AND2X1_LOC_358/a_36_24# AND2X1_LOC_358/Y AND2X1_LOC_358/a_8_24# VSS VDD AND2X1_LOC_350/Y AND2X1_LOC_351/Y AND2X1_LOC

XAND2X1_LOC_732 AND2X1_LOC_732/a_36_24# AND2X1_LOC_738/B AND2X1_LOC_732/a_8_24# VSS VDD AND2X1_LOC_724/Y AND2X1_LOC_732/B AND2X1_LOC

XAND2X1_LOC_865 AND2X1_LOC_865/a_36_24# AND2X1_LOC_866/B AND2X1_LOC_865/a_8_24# VSS VDD AND2X1_LOC_865/A AND2X1_LOC_862/Y AND2X1_LOC

XOR2X1_LOC_578 OR2X1_LOC_578/a_8_216# OR2X1_LOC_578/a_36_216# OR2X1_LOC_580/B VSS VDD OR2X1_LOC_577/Y OR2X1_LOC_578/B OR2X1_LOC

XAND2X1_LOC_364 AND2X1_LOC_364/a_36_24# AND2X1_LOC_364/Y AND2X1_LOC_364/a_8_24# VSS VDD AND2X1_LOC_364/A AND2X1_LOC_358/Y AND2X1_LOC

XOR2X1_LOC_577 OR2X1_LOC_577/a_8_216# OR2X1_LOC_577/a_36_216# OR2X1_LOC_577/Y VSS VDD OR2X1_LOC_570/Y OR2X1_LOC_577/B OR2X1_LOC

XAND2X1_LOC_655 AND2X1_LOC_655/a_36_24# AND2X1_LOC_660/A AND2X1_LOC_655/a_8_24# VSS VDD AND2X1_LOC_655/A AND2X1_LOC_649/Y AND2X1_LOC

XAND2X1_LOC_807 AND2X1_LOC_807/a_36_24# AND2X1_LOC_807/Y AND2X1_LOC_807/a_8_24# VSS VDD AND2X1_LOC_805/Y AND2X1_LOC_807/B AND2X1_LOC

XAND2X1_LOC_741 AND2X1_LOC_741/a_36_24# AND2X1_LOC_741/Y AND2X1_LOC_741/a_8_24# VSS VDD AND2X1_LOC_736/Y AND2X1_LOC_737/Y AND2X1_LOC

XOR2X1_LOC_363 OR2X1_LOC_363/a_8_216# OR2X1_LOC_363/a_36_216# OR2X1_LOC_366/A VSS VDD OR2X1_LOC_363/A OR2X1_LOC_363/B OR2X1_LOC

XOR2X1_LOC_576 OR2X1_LOC_576/a_8_216# OR2X1_LOC_576/a_36_216# OR2X1_LOC_579/A VSS VDD OR2X1_LOC_576/A OR2X1_LOC_571/Y OR2X1_LOC

XOR2X1_LOC_570 OR2X1_LOC_570/a_8_216# OR2X1_LOC_570/a_36_216# OR2X1_LOC_570/Y VSS VDD OR2X1_LOC_570/A OR2X1_LOC_562/Y OR2X1_LOC

XOR2X1_LOC_220 OR2X1_LOC_220/a_8_216# OR2X1_LOC_220/a_36_216# OR2X1_LOC_221/A VSS VDD OR2X1_LOC_220/A OR2X1_LOC_220/B OR2X1_LOC

XAND2X1_LOC_662 AND2X1_LOC_662/a_36_24# AND2X1_LOC_663/B AND2X1_LOC_662/a_8_24# VSS VDD AND2X1_LOC_660/Y AND2X1_LOC_662/B AND2X1_LOC

XAND2X1_LOC_480 AND2X1_LOC_480/a_36_24# GATE_479 AND2X1_LOC_480/a_8_24# VSS VDD AND2X1_LOC_480/A AND2X1_LOC_479/Y AND2X1_LOC

XAND2X1_LOC_223 AND2X1_LOC_223/a_36_24# GATE_222 AND2X1_LOC_223/a_8_24# VSS VDD AND2X1_LOC_223/A AND2X1_LOC_222/Y AND2X1_LOC

XAND2X1_LOC_740 AND2X1_LOC_740/a_36_24# AND2X1_LOC_742/A AND2X1_LOC_740/a_8_24# VSS VDD AND2X1_LOC_738/Y AND2X1_LOC_740/B AND2X1_LOC

XAND2X1_LOC_733 AND2X1_LOC_733/a_36_24# AND2X1_LOC_733/Y AND2X1_LOC_733/a_8_24# VSS VDD AND2X1_LOC_722/Y AND2X1_LOC_723/Y AND2X1_LOC

XOR2X1_LOC_655 OR2X1_LOC_655/a_8_216# OR2X1_LOC_655/a_36_216# OR2X1_LOC_660/B VSS VDD OR2X1_LOC_655/A OR2X1_LOC_655/B OR2X1_LOC

XOR2X1_LOC_579 OR2X1_LOC_579/a_8_216# OR2X1_LOC_579/a_36_216# OR2X1_LOC_580/A VSS VDD OR2X1_LOC_579/A OR2X1_LOC_579/B OR2X1_LOC

XOR2X1_LOC_367 OR2X1_LOC_367/a_8_216# OR2X1_LOC_367/a_36_216# D_GATE_366 VSS VDD OR2X1_LOC_366/Y OR2X1_LOC_367/B OR2X1_LOC

XAND2X1_LOC_222 AND2X1_LOC_222/a_36_24# AND2X1_LOC_222/Y AND2X1_LOC_222/a_8_24# VSS VDD AND2X1_LOC_218/Y AND2X1_LOC_219/Y AND2X1_LOC

XOR2X1_LOC_807 OR2X1_LOC_807/a_8_216# OR2X1_LOC_807/a_36_216# OR2X1_LOC_807/Y VSS VDD OR2X1_LOC_807/A OR2X1_LOC_807/B OR2X1_LOC

XOR2X1_LOC_864 OR2X1_LOC_864/a_8_216# OR2X1_LOC_864/a_36_216# OR2X1_LOC_866/B VSS VDD OR2X1_LOC_864/A OR2X1_LOC_774/Y OR2X1_LOC

XOR2X1_LOC_358 OR2X1_LOC_358/a_8_216# OR2X1_LOC_358/a_36_216# OR2X1_LOC_364/A VSS VDD OR2X1_LOC_358/A OR2X1_LOC_358/B OR2X1_LOC

XAND2X1_LOC_579 AND2X1_LOC_579/a_36_24# AND2X1_LOC_580/B AND2X1_LOC_579/a_8_24# VSS VDD AND2X1_LOC_575/Y AND2X1_LOC_576/Y AND2X1_LOC

XOR2X1_LOC_732 OR2X1_LOC_732/a_8_216# OR2X1_LOC_732/a_36_216# OR2X1_LOC_738/A VSS VDD OR2X1_LOC_732/A OR2X1_LOC_732/B OR2X1_LOC

XOR2X1_LOC_657 OR2X1_LOC_657/a_8_216# OR2X1_LOC_657/a_36_216# OR2X1_LOC_659/B VSS VDD OR2X1_LOC_510/Y OR2X1_LOC_217/A OR2X1_LOC

XOR2X1_LOC_865 OR2X1_LOC_865/a_8_216# OR2X1_LOC_865/a_36_216# OR2X1_LOC_865/Y VSS VDD OR2X1_LOC_865/A OR2X1_LOC_865/B OR2X1_LOC

XAND2X1_LOC_212 AND2X1_LOC_212/a_36_24# AND2X1_LOC_212/Y AND2X1_LOC_212/a_8_24# VSS VDD AND2X1_LOC_212/A AND2X1_LOC_212/B AND2X1_LOC

XAND2X1_LOC_657 AND2X1_LOC_657/a_36_24# AND2X1_LOC_657/Y AND2X1_LOC_657/a_8_24# VSS VDD AND2X1_LOC_657/A AND2X1_LOC_574/A AND2X1_LOC

XAND2X1_LOC_578 AND2X1_LOC_578/a_36_24# AND2X1_LOC_580/A AND2X1_LOC_578/a_8_24# VSS VDD AND2X1_LOC_578/A AND2X1_LOC_577/Y AND2X1_LOC

XAND2X1_LOC_576 AND2X1_LOC_576/a_36_24# AND2X1_LOC_576/Y AND2X1_LOC_576/a_8_24# VSS VDD AND2X1_LOC_571/Y AND2X1_LOC_572/Y AND2X1_LOC

XAND2X1_LOC_363 AND2X1_LOC_363/a_36_24# AND2X1_LOC_363/Y AND2X1_LOC_363/a_8_24# VSS VDD AND2X1_LOC_363/A AND2X1_LOC_363/B AND2X1_LOC

XAND2X1_LOC_659 AND2X1_LOC_659/a_36_24# AND2X1_LOC_663/A AND2X1_LOC_659/a_8_24# VSS VDD AND2X1_LOC_657/Y AND2X1_LOC_658/Y AND2X1_LOC

XOR2X1_LOC_803 OR2X1_LOC_803/a_8_216# OR2X1_LOC_803/a_36_216# OR2X1_LOC_808/B VSS VDD OR2X1_LOC_803/A OR2X1_LOC_803/B OR2X1_LOC

XAND2X1_LOC_570 AND2X1_LOC_570/a_36_24# AND2X1_LOC_570/Y AND2X1_LOC_570/a_8_24# VSS VDD AND2X1_LOC_562/Y AND2X1_LOC_563/Y AND2X1_LOC

XOR2X1_LOC_733 OR2X1_LOC_733/a_8_216# OR2X1_LOC_733/a_36_216# OR2X1_LOC_733/Y VSS VDD OR2X1_LOC_733/A OR2X1_LOC_733/B OR2X1_LOC

XOR2X1_LOC_364 OR2X1_LOC_364/a_8_216# OR2X1_LOC_364/a_36_216# OR2X1_LOC_364/Y VSS VDD OR2X1_LOC_364/A OR2X1_LOC_364/B OR2X1_LOC

XOR2X1_LOC_738 OR2X1_LOC_738/a_8_216# OR2X1_LOC_738/a_36_216# OR2X1_LOC_740/B VSS VDD OR2X1_LOC_738/A OR2X1_LOC_738/B OR2X1_LOC

XAND2X1_LOC_804 AND2X1_LOC_804/a_36_24# AND2X1_LOC_804/Y AND2X1_LOC_804/a_8_24# VSS VDD AND2X1_LOC_804/A AND2X1_LOC_795/Y AND2X1_LOC

XOR2X1_LOC_478 OR2X1_LOC_478/a_8_216# OR2X1_LOC_478/a_36_216# OR2X1_LOC_478/Y VSS VDD OR2X1_LOC_477/Y OR2X1_LOC_469/Y OR2X1_LOC

XAND2X1_LOC_215 AND2X1_LOC_215/a_36_24# AND2X1_LOC_215/Y AND2X1_LOC_215/a_8_24# VSS VDD AND2X1_LOC_215/A AND2X1_LOC_206/Y AND2X1_LOC

XOR2X1_LOC_219 OR2X1_LOC_219/a_8_216# OR2X1_LOC_219/a_36_216# OR2X1_LOC_222/A VSS VDD OR2X1_LOC_215/Y OR2X1_LOC_219/B OR2X1_LOC

XOR2X1_LOC_659 OR2X1_LOC_659/a_8_216# OR2X1_LOC_659/a_36_216# OR2X1_LOC_659/Y VSS VDD OR2X1_LOC_659/A OR2X1_LOC_659/B OR2X1_LOC

XAND2X1_LOC_803 AND2X1_LOC_803/a_36_24# AND2X1_LOC_808/A AND2X1_LOC_803/a_8_24# VSS VDD AND2X1_LOC_796/Y AND2X1_LOC_803/B AND2X1_LOC

XAND2X1_LOC_219 AND2X1_LOC_219/a_36_24# AND2X1_LOC_219/Y AND2X1_LOC_219/a_8_24# VSS VDD AND2X1_LOC_219/A AND2X1_LOC_215/Y AND2X1_LOC

XAND2X1_LOC_577 AND2X1_LOC_577/a_36_24# AND2X1_LOC_577/Y AND2X1_LOC_577/a_8_24# VSS VDD AND2X1_LOC_577/A AND2X1_LOC_570/Y AND2X1_LOC

XOR2X1_LOC_480 OR2X1_LOC_480/a_8_216# OR2X1_LOC_480/a_36_216# D_GATE_479 VSS VDD OR2X1_LOC_479/Y OR2X1_LOC_478/Y OR2X1_LOC

XOR2X1_LOC_741 OR2X1_LOC_741/a_8_216# OR2X1_LOC_741/a_36_216# OR2X1_LOC_741/Y VSS VDD OR2X1_LOC_741/A OR2X1_LOC_736/Y OR2X1_LOC

XOR2X1_LOC_740 OR2X1_LOC_740/a_8_216# OR2X1_LOC_740/a_36_216# OR2X1_LOC_742/B VSS VDD OR2X1_LOC_739/Y OR2X1_LOC_740/B OR2X1_LOC

XOR2X1_LOC_223 OR2X1_LOC_223/a_8_216# OR2X1_LOC_223/a_36_216# D_GATE_222 VSS VDD OR2X1_LOC_223/A OR2X1_LOC_223/B OR2X1_LOC

XOR2X1_LOC_804 OR2X1_LOC_804/a_8_216# OR2X1_LOC_804/a_36_216# OR2X1_LOC_808/A VSS VDD OR2X1_LOC_804/A OR2X1_LOC_804/B OR2X1_LOC

XAND2X1_LOC_220 AND2X1_LOC_220/a_36_24# AND2X1_LOC_220/Y AND2X1_LOC_220/a_8_24# VSS VDD AND2X1_LOC_212/Y AND2X1_LOC_220/B AND2X1_LOC

XAND2X1_LOC_738 AND2X1_LOC_738/a_36_24# AND2X1_LOC_738/Y AND2X1_LOC_738/a_8_24# VSS VDD AND2X1_LOC_731/Y AND2X1_LOC_738/B AND2X1_LOC

XOR2X1_LOC_212 OR2X1_LOC_212/a_8_216# OR2X1_LOC_212/a_36_216# OR2X1_LOC_220/B VSS VDD OR2X1_LOC_212/A OR2X1_LOC_212/B OR2X1_LOC

XOR2X1_LOC_215 OR2X1_LOC_215/a_8_216# OR2X1_LOC_215/a_36_216# OR2X1_LOC_215/Y VSS VDD OR2X1_LOC_215/A OR2X1_LOC_205/Y OR2X1_LOC

XOR2X1_LOC_808 OR2X1_LOC_808/a_8_216# OR2X1_LOC_808/a_36_216# OR2X1_LOC_811/A VSS VDD OR2X1_LOC_808/A OR2X1_LOC_808/B OR2X1_LOC

XOR2X1_LOC_742 OR2X1_LOC_742/a_8_216# OR2X1_LOC_742/a_36_216# D_GATE_741 VSS VDD OR2X1_LOC_741/Y OR2X1_LOC_742/B OR2X1_LOC

XAND2X1_LOC_808 AND2X1_LOC_808/a_36_24# AND2X1_LOC_811/B AND2X1_LOC_808/a_8_24# VSS VDD AND2X1_LOC_808/A AND2X1_LOC_804/Y AND2X1_LOC

XOR2X1_LOC_663 OR2X1_LOC_663/a_8_216# OR2X1_LOC_663/a_36_216# D_GATE_662 VSS VDD OR2X1_LOC_663/A OR2X1_LOC_659/Y OR2X1_LOC

XAND2X1_LOC_663 AND2X1_LOC_663/a_36_24# GATE_662 AND2X1_LOC_663/a_8_24# VSS VDD AND2X1_LOC_663/A AND2X1_LOC_663/B AND2X1_LOC

XAND2X1_LOC_580 AND2X1_LOC_580/a_36_24# GATE_579 AND2X1_LOC_580/a_8_24# VSS VDD AND2X1_LOC_580/A AND2X1_LOC_580/B AND2X1_LOC

XOR2X1_LOC_866 OR2X1_LOC_866/a_8_216# OR2X1_LOC_866/a_36_216# D_GATE_865 VSS VDD OR2X1_LOC_865/Y OR2X1_LOC_866/B OR2X1_LOC

XOR2X1_LOC_811 OR2X1_LOC_811/a_8_216# OR2X1_LOC_811/a_36_216# OR2X1_LOC_812/A VSS VDD OR2X1_LOC_811/A OR2X1_LOC_807/Y OR2X1_LOC

XOR2X1_LOC_580 OR2X1_LOC_580/a_8_216# OR2X1_LOC_580/a_36_216# D_GATE_579 VSS VDD OR2X1_LOC_580/A OR2X1_LOC_580/B OR2X1_LOC

XAND2X1_LOC_742 AND2X1_LOC_742/a_36_24# GATE_741 AND2X1_LOC_742/a_8_24# VSS VDD AND2X1_LOC_742/A AND2X1_LOC_741/Y AND2X1_LOC

XAND2X1_LOC_811 AND2X1_LOC_811/a_36_24# AND2X1_LOC_811/Y AND2X1_LOC_811/a_8_24# VSS VDD AND2X1_LOC_807/Y AND2X1_LOC_811/B AND2X1_LOC

XAND2X1_LOC_866 AND2X1_LOC_866/a_36_24# GATE_865 AND2X1_LOC_866/a_8_24# VSS VDD AND2X1_LOC_866/A AND2X1_LOC_866/B AND2X1_LOC

C4433 OR2X1_LOC_643/Y OR2X1_LOC_228/Y 0.02fF
C13305 OR2X1_LOC_643/Y OR2X1_LOC_215/Y 0.09fF
C15500 OR2X1_LOC_643/Y OR2X1_LOC_341/a_8_216# 0.01fF
C24337 OR2X1_LOC_643/Y OR2X1_LOC_219/a_8_216# 0.39fF
C30136 OR2X1_LOC_641/Y OR2X1_LOC_643/Y 0.26fF
C35255 OR2X1_LOC_643/Y OR2X1_LOC_222/A 0.01fF
C42082 OR2X1_LOC_643/Y OR2X1_LOC_341/Y 0.01fF
C47804 OR2X1_LOC_643/Y OR2X1_LOC_340/Y 0.02fF
C50768 OR2X1_LOC_662/A OR2X1_LOC_643/Y 0.06fF
C52458 OR2X1_LOC_864/A OR2X1_LOC_643/Y 0.03fF
C55083 OR2X1_LOC_643/Y OR2X1_LOC_641/B 0.72fF
C57229 OR2X1_LOC_643/Y VSS 0.19fF
C1668 VDD OR2X1_LOC_201/Y 0.12fF
C53769 OR2X1_LOC_206/A OR2X1_LOC_201/Y 0.04fF
C56856 OR2X1_LOC_201/Y VSS 0.15fF
C1119 OR2X1_LOC_719/Y OR2X1_LOC_722/B 0.07fF
C17673 OR2X1_LOC_722/a_8_216# OR2X1_LOC_722/B 0.18fF
C21056 OR2X1_LOC_808/B OR2X1_LOC_722/B 0.02fF
C21518 OR2X1_LOC_808/A OR2X1_LOC_722/B 0.10fF
C24030 VDD OR2X1_LOC_722/B 0.06fF
C33297 OR2X1_LOC_737/A OR2X1_LOC_722/B 0.02fF
C35840 OR2X1_LOC_808/a_8_216# OR2X1_LOC_722/B 0.40fF
C39722 OR2X1_LOC_733/B OR2X1_LOC_722/B 0.21fF
C56280 OR2X1_LOC_722/B VSS 0.28fF
C13428 OR2X1_LOC_562/a_8_216# OR2X1_LOC_562/B 0.39fF
C19781 VDD OR2X1_LOC_562/B -0.00fF
C47448 OR2X1_LOC_562/B OR2X1_LOC_562/A 0.14fF
C56440 OR2X1_LOC_562/B VSS 0.17fF
C7022 OR2X1_LOC_479/Y OR2X1_LOC_469/B 0.09fF
C8609 OR2X1_LOC_182/a_8_216# OR2X1_LOC_469/B 0.40fF
C16290 VDD OR2X1_LOC_469/B 0.14fF
C18928 OR2X1_LOC_468/Y OR2X1_LOC_469/B 0.05fF
C29937 OR2X1_LOC_469/a_8_216# OR2X1_LOC_469/B 0.03fF
C35830 OR2X1_LOC_738/A OR2X1_LOC_469/B 0.01fF
C38329 OR2X1_LOC_739/A OR2X1_LOC_469/B 0.03fF
C42660 OR2X1_LOC_212/a_8_216# OR2X1_LOC_469/B 0.02fF
C47422 OR2X1_LOC_486/Y OR2X1_LOC_469/B 4.61fF
C53697 OR2X1_LOC_181/Y OR2X1_LOC_469/B 0.08fF
C53836 OR2X1_LOC_220/B OR2X1_LOC_469/B 0.07fF
C56373 OR2X1_LOC_469/B VSS 0.18fF
C3553 OR2X1_LOC_805/A OR2X1_LOC_786/Y 0.10fF
C4485 OR2X1_LOC_786/Y OR2X1_LOC_228/Y 0.01fF
C11957 OR2X1_LOC_786/Y OR2X1_LOC_795/B 0.12fF
C25641 OR2X1_LOC_205/a_8_216# OR2X1_LOC_786/Y 0.01fF
C27453 OR2X1_LOC_786/Y OR2X1_LOC_560/A 0.16fF
C29030 OR2X1_LOC_206/A OR2X1_LOC_786/Y 0.13fF
C30794 OR2X1_LOC_786/Y OR2X1_LOC_795/a_8_216# 0.02fF
C32282 OR2X1_LOC_663/A OR2X1_LOC_786/Y 0.03fF
C33130 VDD OR2X1_LOC_786/Y 1.70fF
C35856 OR2X1_LOC_205/Y OR2X1_LOC_786/Y 0.14fF
C37194 OR2X1_LOC_786/Y OR2X1_LOC_217/A 0.02fF
C39589 OR2X1_LOC_124/Y OR2X1_LOC_786/Y 0.03fF
C42571 OR2X1_LOC_786/Y OR2X1_LOC_737/A 0.10fF
C42955 OR2X1_LOC_244/B OR2X1_LOC_786/Y 0.02fF
C44733 OR2X1_LOC_217/Y OR2X1_LOC_786/Y 0.23fF
C45196 OR2X1_LOC_217/a_8_216# OR2X1_LOC_786/Y 0.04fF
C50846 OR2X1_LOC_217/a_36_216# OR2X1_LOC_786/Y 0.01fF
C52496 OR2X1_LOC_864/A OR2X1_LOC_786/Y 0.03fF
C56840 OR2X1_LOC_786/Y VSS -2.78fF
C1105 OR2X1_LOC_641/Y OR2X1_LOC_650/a_8_216# 0.03fF
C10541 OR2X1_LOC_641/Y OR2X1_LOC_662/A 0.30fF
C16068 OR2X1_LOC_641/Y OR2X1_LOC_649/B 0.01fF
C28742 OR2X1_LOC_641/Y OR2X1_LOC_655/a_8_216# 0.02fF
C41133 OR2X1_LOC_641/Y OR2X1_LOC_649/a_8_216# 0.40fF
C45371 OR2X1_LOC_641/Y OR2X1_LOC_660/B 0.01fF
C51766 OR2X1_LOC_641/Y OR2X1_LOC_640/Y 0.12fF
C51950 OR2X1_LOC_641/Y OR2X1_LOC_655/B 0.12fF
C52373 OR2X1_LOC_641/Y OR2X1_LOC_655/A 0.03fF
C54031 OR2X1_LOC_641/Y OR2X1_LOC_650/Y 0.02fF
C57838 OR2X1_LOC_641/Y VSS 0.49fF
C9409 OR2X1_LOC_805/A OR2X1_LOC_203/Y 0.07fF
C20448 OR2X1_LOC_204/Y OR2X1_LOC_203/Y 0.29fF
C31427 OR2X1_LOC_203/Y OR2X1_LOC_205/a_8_216# 0.10fF
C41727 OR2X1_LOC_205/Y OR2X1_LOC_203/Y 0.02fF
C45523 OR2X1_LOC_203/Y OR2X1_LOC_124/Y 0.30fF
C48939 OR2X1_LOC_244/B OR2X1_LOC_203/Y 0.02fF
C50730 OR2X1_LOC_217/Y OR2X1_LOC_203/Y 0.01fF
C51132 OR2X1_LOC_203/Y OR2X1_LOC_217/a_8_216# 0.02fF
C56898 OR2X1_LOC_203/Y VSS 0.70fF
C4026 OR2X1_LOC_175/Y OR2X1_LOC_468/A 0.07fF
C4365 OR2X1_LOC_175/Y OR2X1_LOC_857/A 0.18fF
C6175 OR2X1_LOC_175/Y OR2X1_LOC_214/a_8_216# 0.01fF
C8409 OR2X1_LOC_864/A OR2X1_LOC_175/Y 0.03fF
C12466 OR2X1_LOC_566/A OR2X1_LOC_175/Y 0.27fF
C15400 OR2X1_LOC_175/Y OR2X1_LOC_214/A 0.01fF
C15536 OR2X1_LOC_175/Y OR2X1_LOC_805/A 0.03fF
C15872 OR2X1_LOC_175/Y OR2X1_LOC_648/B 0.10fF
C16595 OR2X1_LOC_175/Y OR2X1_LOC_228/Y 0.22fF
C16973 OR2X1_LOC_175/Y OR2X1_LOC_436/Y 0.13fF
C17036 OR2X1_LOC_175/Y OR2X1_LOC_566/Y 0.09fF
C17280 OR2X1_LOC_175/Y OR2X1_LOC_219/B 0.01fF
C19613 OR2X1_LOC_175/Y OR2X1_LOC_170/Y 0.09fF
C22564 OR2X1_LOC_175/Y OR2X1_LOC_468/a_8_216# 0.05fF
C22639 OR2X1_LOC_175/Y OR2X1_LOC_568/a_8_216# 0.03fF
C23425 OR2X1_LOC_175/Y OR2X1_LOC_214/B 0.02fF
C24988 OR2X1_LOC_175/Y OR2X1_LOC_857/a_8_216# 0.04fF
C26075 OR2X1_LOC_857/B OR2X1_LOC_175/Y 0.08fF
C30582 OR2X1_LOC_175/Y OR2X1_LOC_566/a_8_216# 0.08fF
C42218 OR2X1_LOC_175/Y OR2X1_LOC_808/B 0.09fF
C44658 OR2X1_LOC_175/Y OR2X1_LOC_568/A 0.80fF
C44665 OR2X1_LOC_175/Y OR2X1_LOC_578/B 0.01fF
C48000 OR2X1_LOC_863/a_8_216# OR2X1_LOC_175/Y 0.04fF
C48001 OR2X1_LOC_175/Y OR2X1_LOC_468/Y 0.03fF
C49576 OR2X1_LOC_175/Y OR2X1_LOC_853/a_8_216# 0.01fF
C50573 OR2X1_LOC_175/Y OR2X1_LOC_863/B 0.06fF
C52523 OR2X1_LOC_175/Y OR2X1_LOC_863/A 0.04fF
C57859 OR2X1_LOC_175/Y VSS -1.06fF
C9137 OR2X1_LOC_182/B OR2X1_LOC_357/B 0.01fF
C10434 OR2X1_LOC_486/Y OR2X1_LOC_182/B 0.03fF
C15003 OR2X1_LOC_182/B OR2X1_LOC_357/A 0.02fF
C26266 OR2X1_LOC_479/Y OR2X1_LOC_182/B 0.03fF
C27734 OR2X1_LOC_182/B OR2X1_LOC_182/a_8_216# 0.02fF
C30815 OR2X1_LOC_352/A OR2X1_LOC_182/B 0.96fF
C34897 OR2X1_LOC_182/B OR2X1_LOC_578/B 0.04fF
C35346 OR2X1_LOC_357/a_8_216# OR2X1_LOC_182/B 0.01fF
C35376 VDD OR2X1_LOC_182/B 0.10fF
C38721 OR2X1_LOC_182/B OR2X1_LOC_212/B 0.44fF
C46576 OR2X1_LOC_364/B OR2X1_LOC_182/B 0.01fF
C48743 OR2X1_LOC_182/B OR2X1_LOC_352/a_8_216# 0.01fF
C50353 OR2X1_LOC_182/B OR2X1_LOC_365/B 0.25fF
C56536 OR2X1_LOC_182/B VSS 0.18fF
C84 OR2X1_LOC_736/A OR2X1_LOC_675/Y 0.04fF
C706 OR2X1_LOC_675/Y OR2X1_LOC_736/a_8_216# 0.14fF
C5400 OR2X1_LOC_675/Y OR2X1_LOC_580/A 0.07fF
C10396 OR2X1_LOC_631/B OR2X1_LOC_675/Y 0.02fF
C15822 OR2X1_LOC_811/A OR2X1_LOC_675/Y 2.04fF
C17550 OR2X1_LOC_807/A OR2X1_LOC_675/Y 0.16fF
C28532 OR2X1_LOC_348/Y OR2X1_LOC_675/Y 0.07fF
C30716 OR2X1_LOC_807/a_8_216# OR2X1_LOC_675/Y 0.02fF
C40394 OR2X1_LOC_792/Y OR2X1_LOC_675/Y 0.01fF
C44027 OR2X1_LOC_675/Y OR2X1_LOC_366/a_8_216# 0.05fF
C45982 OR2X1_LOC_736/Y OR2X1_LOC_675/Y 0.04fF
C49062 VDD OR2X1_LOC_675/Y 0.46fF
C51653 OR2X1_LOC_362/B OR2X1_LOC_675/Y 0.32fF
C56462 OR2X1_LOC_675/Y VSS -1.69fF
C2291 OR2X1_LOC_244/Y OR2X1_LOC_735/B 0.02fF
C10374 OR2X1_LOC_735/a_8_216# OR2X1_LOC_735/B 0.39fF
C38275 OR2X1_LOC_858/A OR2X1_LOC_735/B 0.02fF
C50005 OR2X1_LOC_632/Y OR2X1_LOC_735/B 0.23fF
C56403 OR2X1_LOC_735/B VSS -0.05fF
C3614 OR2X1_LOC_479/Y OR2X1_LOC_551/B 0.03fF
C12047 OR2X1_LOC_364/A OR2X1_LOC_551/B 0.10fF
C12230 OR2X1_LOC_551/B OR2X1_LOC_578/B 0.68fF
C12844 VDD OR2X1_LOC_551/B 0.05fF
C13073 OR2X1_LOC_551/B OR2X1_LOC_551/A 0.08fF
C15486 OR2X1_LOC_471/Y OR2X1_LOC_551/B 0.19fF
C19635 OR2X1_LOC_551/B OR2X1_LOC_364/a_8_216# 0.40fF
C26230 OR2X1_LOC_551/B OR2X1_LOC_364/Y 0.07fF
C27455 OR2X1_LOC_551/B OR2X1_LOC_365/B 0.06fF
C37188 OR2X1_LOC_551/B OR2X1_LOC_365/a_8_216# 0.03fF
C43803 OR2X1_LOC_486/Y OR2X1_LOC_551/B 0.07fF
C45794 OR2X1_LOC_742/B OR2X1_LOC_551/B 0.09fF
C48510 OR2X1_LOC_551/B OR2X1_LOC_367/B 0.20fF
C50214 OR2X1_LOC_551/B OR2X1_LOC_181/Y 0.02fF
C56444 OR2X1_LOC_551/B VSS 0.37fF
C6747 AND2X1_LOC_554/Y AND2X1_LOC_572/A 0.17fF
C9688 AND2X1_LOC_554/Y AND2X1_LOC_563/A 0.01fF
C29206 AND2X1_LOC_554/Y AND2X1_LOC_367/A 0.10fF
C30380 AND2X1_LOC_572/a_8_24# AND2X1_LOC_554/Y 0.03fF
C37857 AND2X1_LOC_554/Y AND2X1_LOC_657/A 0.47fF
C38004 AND2X1_LOC_554/Y VDD 0.23fF
C49429 AND2X1_LOC_554/Y AND2X1_LOC_361/A 0.05fF
C49832 AND2X1_LOC_554/Y AND2X1_LOC_572/Y 0.17fF
C57994 AND2X1_LOC_554/Y VSS -0.32fF
C12405 AND2X1_LOC_797/a_8_24# AND2X1_LOC_797/B 0.01fF
C23498 AND2X1_LOC_803/B AND2X1_LOC_797/B 0.01fF
C49919 VDD AND2X1_LOC_797/B 0.13fF
C56352 AND2X1_LOC_797/B VSS 0.19fF
C9071 AND2X1_LOC_726/Y AND2X1_LOC_727/Y 0.11fF
C11220 AND2X1_LOC_726/Y AND2X1_LOC_731/Y 0.02fF
C14599 AND2X1_LOC_726/Y AND2X1_LOC_731/a_8_24# 0.18fF
C27769 AND2X1_LOC_726/Y VDD 0.21fF
C58087 AND2X1_LOC_726/Y VSS 0.06fF
C1832 AND2X1_LOC_213/B AND2X1_LOC_209/Y 0.01fF
C11608 AND2X1_LOC_209/Y AND2X1_LOC_213/a_8_24# 0.09fF
C25249 AND2X1_LOC_803/B AND2X1_LOC_209/Y 0.01fF
C47602 AND2X1_LOC_797/A AND2X1_LOC_209/Y 0.09fF
C56450 AND2X1_LOC_209/Y VSS 0.08fF
C1169 AND2X1_LOC_572/A AND2X1_LOC_243/Y 0.02fF
C7589 AND2X1_LOC_474/A AND2X1_LOC_572/A 0.03fF
C16626 AND2X1_LOC_572/A AND2X1_LOC_663/B 0.06fF
C20596 AND2X1_LOC_572/A AND2X1_LOC_657/A 0.14fF
C20749 VDD AND2X1_LOC_572/A 0.15fF
C31821 AND2X1_LOC_572/A AND2X1_LOC_361/A 0.14fF
C36900 AND2X1_LOC_141/B AND2X1_LOC_572/A 0.11fF
C57329 AND2X1_LOC_572/A VSS 0.23fF
C2672 AND2X1_LOC_347/Y AND2X1_LOC_866/A 0.07fF
C23629 AND2X1_LOC_555/Y AND2X1_LOC_347/Y 0.02fF
C31716 AND2X1_LOC_347/Y AND2X1_LOC_360/a_8_24# 0.11fF
C32220 AND2X1_LOC_347/Y AND2X1_LOC_663/B 0.04fF
C36300 AND2X1_LOC_347/Y VDD 0.12fF
C57985 AND2X1_LOC_347/Y VSS 0.20fF
C1245 AND2X1_LOC_738/B AND2X1_LOC_645/A 0.01fF
C2514 AND2X1_LOC_713/Y AND2X1_LOC_645/A 0.09fF
C34067 AND2X1_LOC_645/a_8_24# AND2X1_LOC_645/A 0.10fF
C40633 AND2X1_LOC_724/Y AND2X1_LOC_645/A 1.03fF
C48293 AND2X1_LOC_477/A AND2X1_LOC_645/A 0.07fF
C50200 VDD AND2X1_LOC_645/A 0.24fF
C56806 AND2X1_LOC_645/A VSS 0.22fF
C2860 AND2X1_LOC_204/Y AND2X1_LOC_205/a_8_24# 0.03fF
C13911 AND2X1_LOC_204/Y AND2X1_LOC_205/a_36_24# 0.01fF
C24748 VDD AND2X1_LOC_204/Y 0.01fF
C47991 AND2X1_LOC_203/Y AND2X1_LOC_204/Y 0.28fF
C56319 AND2X1_LOC_204/Y VSS 0.32fF
C3924 VDD AND2X1_LOC_483/Y -0.00fF
C53273 AND2X1_LOC_658/A AND2X1_LOC_483/Y 0.03fF
C57011 AND2X1_LOC_483/Y VSS 0.15fF
C2457 AND2X1_LOC_468/B AND2X1_LOC_477/Y 0.01fF
C11313 AND2X1_LOC_468/B AND2X1_LOC_212/Y 0.07fF
C12248 AND2X1_LOC_468/B AND2X1_LOC_471/Y 0.23fF
C21622 AND2X1_LOC_468/B AND2X1_LOC_436/Y 0.01fF
C24399 AND2X1_LOC_468/B AND2X1_LOC_222/Y 0.01fF
C31086 AND2X1_LOC_468/B AND2X1_LOC_810/Y 0.02fF
C31464 AND2X1_LOC_477/A AND2X1_LOC_468/B 0.03fF
C32555 AND2X1_LOC_468/B AND2X1_LOC_468/a_8_24# 0.01fF
C33353 AND2X1_LOC_794/B AND2X1_LOC_468/B 0.10fF
C33391 VDD AND2X1_LOC_468/B 0.10fF
C38020 AND2X1_LOC_468/B AND2X1_LOC_469/B 0.04fF
C38041 AND2X1_LOC_733/Y AND2X1_LOC_468/B 0.91fF
C55668 AND2X1_LOC_722/A AND2X1_LOC_468/B 0.94fF
C57067 AND2X1_LOC_468/B VSS 0.29fF
C681 AND2X1_LOC_231/Y AND2X1_LOC_650/Y 0.26fF
C3690 AND2X1_LOC_231/Y AND2X1_LOC_228/Y 0.07fF
C4062 AND2X1_LOC_231/Y AND2X1_LOC_857/Y 0.01fF
C6201 AND2X1_LOC_231/Y AND2X1_LOC_211/B 0.26fF
C19765 AND2X1_LOC_231/Y VDD 0.06fF
C27090 AND2X1_LOC_231/Y AND2X1_LOC_641/Y 0.07fF
C57846 AND2X1_LOC_231/Y VSS 0.18fF
C8223 AND2X1_LOC_141/B AND2X1_LOC_663/B 0.10fF
C11061 AND2X1_LOC_141/B AND2X1_LOC_141/A 0.14fF
C12100 AND2X1_LOC_141/B AND2X1_LOC_657/A 0.18fF
C12308 VDD AND2X1_LOC_141/B 0.01fF
C23223 AND2X1_LOC_141/B AND2X1_LOC_217/a_8_24# 0.07fF
C39658 AND2X1_LOC_141/B AND2X1_LOC_217/a_36_24# 0.01fF
C43035 AND2X1_LOC_141/B AND2X1_LOC_656/Y 0.15fF
C46349 AND2X1_LOC_141/B AND2X1_LOC_141/a_8_24# 0.06fF
C56146 AND2X1_LOC_217/Y AND2X1_LOC_141/B 0.01fF
C57704 AND2X1_LOC_141/B VSS 0.36fF
C10526 OR2X1_LOC_631/B OR2X1_LOC_736/Y 0.19fF
C13553 VDD OR2X1_LOC_631/B 0.63fF
C29966 OR2X1_LOC_631/B OR2X1_LOC_556/a_8_216# 0.41fF
C32156 OR2X1_LOC_858/A OR2X1_LOC_631/B 0.03fF
C35429 OR2X1_LOC_631/B OR2X1_LOC_556/a_36_216# 0.01fF
C36436 OR2X1_LOC_631/B OR2X1_LOC_811/A 0.07fF
C39874 OR2X1_LOC_631/B OR2X1_LOC_805/A 0.07fF
C43166 OR2X1_LOC_631/B OR2X1_LOC_563/A 0.03fF
C43705 OR2X1_LOC_631/B OR2X1_LOC_632/Y 0.01fF
C44485 OR2X1_LOC_631/B OR2X1_LOC_486/Y 0.09fF
C57633 OR2X1_LOC_631/B VSS 0.42fF
C10868 VDD OR2X1_LOC_468/A 0.26fF
C13550 OR2X1_LOC_468/A OR2X1_LOC_468/Y 0.02fF
C38609 OR2X1_LOC_468/A OR2X1_LOC_436/Y 0.52fF
C44219 OR2X1_LOC_468/A OR2X1_LOC_468/a_8_216# 0.18fF
C57566 OR2X1_LOC_468/A VSS -0.01fF
C679 OR2X1_LOC_244/A OR2X1_LOC_140/Y 0.20fF
C11183 OR2X1_LOC_244/Y OR2X1_LOC_140/Y 0.01fF
C18879 OR2X1_LOC_244/a_8_216# OR2X1_LOC_140/Y 0.01fF
C23920 OR2X1_LOC_267/Y OR2X1_LOC_140/Y 0.01fF
C38283 OR2X1_LOC_244/B OR2X1_LOC_140/Y 0.11fF
C56287 OR2X1_LOC_140/Y VSS 0.10fF
C7119 VDD OR2X1_LOC_193/Y 0.12fF
C12801 OR2X1_LOC_194/Y OR2X1_LOC_193/Y 0.12fF
C32506 OR2X1_LOC_207/B OR2X1_LOC_193/Y 0.21fF
C57149 OR2X1_LOC_193/Y VSS 0.07fF
C7936 OR2X1_LOC_787/Y OR2X1_LOC_605/Y 0.01fF
C15644 OR2X1_LOC_223/A OR2X1_LOC_605/Y 0.15fF
C30757 OR2X1_LOC_794/A OR2X1_LOC_605/Y -0.00fF
C37560 OR2X1_LOC_479/Y OR2X1_LOC_605/Y 0.12fF
C44372 OR2X1_LOC_808/A OR2X1_LOC_605/Y 0.01fF
C46170 OR2X1_LOC_364/A OR2X1_LOC_605/Y 0.01fF
C46998 VDD OR2X1_LOC_605/Y 0.23fF
C48336 OR2X1_LOC_602/Y OR2X1_LOC_605/Y 0.15fF
C56281 OR2X1_LOC_605/Y VSS 0.27fF
C6725 OR2X1_LOC_653/Y OR2X1_LOC_805/A 0.46fF
C7052 OR2X1_LOC_653/Y OR2X1_LOC_648/B 0.18fF
C7800 OR2X1_LOC_653/Y OR2X1_LOC_228/Y 0.02fF
C8560 OR2X1_LOC_653/Y OR2X1_LOC_219/B 0.07fF
C10782 OR2X1_LOC_653/Y OR2X1_LOC_358/A 0.01fF
C24641 OR2X1_LOC_358/a_8_216# OR2X1_LOC_653/Y 0.03fF
C28104 OR2X1_LOC_653/Y OR2X1_LOC_648/a_8_216# 0.03fF
C35597 OR2X1_LOC_364/A OR2X1_LOC_653/Y 0.23fF
C36326 OR2X1_LOC_653/Y VDD 0.12fF
C37240 OR2X1_LOC_653/Y OR2X1_LOC_661/a_8_216# 0.03fF
C37559 OR2X1_LOC_653/Y OR2X1_LOC_661/A 0.04fF
C39087 OR2X1_LOC_653/Y OR2X1_LOC_655/B 0.01fF
C53998 OR2X1_LOC_653/Y OR2X1_LOC_662/A 0.01fF
C54332 OR2X1_LOC_653/Y OR2X1_LOC_648/A 0.75fF
C55756 OR2X1_LOC_864/A OR2X1_LOC_653/Y 0.07fF
C57836 OR2X1_LOC_653/Y VSS 0.17fF
C4737 OR2X1_LOC_223/A OR2X1_LOC_794/A 0.02fF
C8110 OR2X1_LOC_794/a_8_216# OR2X1_LOC_794/A 0.18fF
C26784 OR2X1_LOC_479/Y OR2X1_LOC_794/A 0.01fF
C33422 OR2X1_LOC_808/A OR2X1_LOC_794/A 0.01fF
C35166 OR2X1_LOC_364/A OR2X1_LOC_794/A 0.03fF
C35906 VDD OR2X1_LOC_794/A 0.18fF
C53222 OR2X1_LOC_787/Y OR2X1_LOC_794/A 0.44fF
C56611 OR2X1_LOC_794/A VSS 0.07fF
C1684 OR2X1_LOC_739/B OR2X1_LOC_739/A 0.14fF
C14510 OR2X1_LOC_221/A OR2X1_LOC_739/B 0.90fF
C16982 OR2X1_LOC_739/B OR2X1_LOC_220/B 0.14fF
C17327 OR2X1_LOC_739/B D_GATE_741 0.01fF
C24649 OR2X1_LOC_739/B OR2X1_LOC_221/a_8_216# 0.09fF
C25757 OR2X1_LOC_739/B OR2X1_LOC_740/B 0.07fF
C30127 OR2X1_LOC_739/B OR2X1_LOC_221/a_36_216# 0.03fF
C33180 OR2X1_LOC_739/B OR2X1_LOC_223/a_8_216# 0.14fF
C35493 VDD OR2X1_LOC_739/B 0.37fF
C35601 OR2X1_LOC_739/B OR2X1_LOC_223/B 0.23fF
C37862 OR2X1_LOC_739/B OR2X1_LOC_739/a_8_216# 0.07fF
C44284 OR2X1_LOC_739/B D_GATE_222 0.05fF
C54057 OR2X1_LOC_220/a_8_216# OR2X1_LOC_739/B 0.14fF
C57200 OR2X1_LOC_739/B VSS 0.17fF
C5318 VDD OR2X1_LOC_737/A 0.12fF
C10915 OR2X1_LOC_733/A OR2X1_LOC_737/A 0.04fF
C17349 OR2X1_LOC_733/a_8_216# OR2X1_LOC_737/A 0.01fF
C19711 OR2X1_LOC_737/A OR2X1_LOC_723/A 0.04fF
C21312 OR2X1_LOC_733/B OR2X1_LOC_737/A 0.12fF
C24158 OR2X1_LOC_858/A OR2X1_LOC_737/A 0.03fF
C28396 OR2X1_LOC_811/A OR2X1_LOC_737/A 0.14fF
C31778 OR2X1_LOC_805/A OR2X1_LOC_737/A 0.08fF
C38551 OR2X1_LOC_719/Y OR2X1_LOC_737/A 0.01fF
C45172 OR2X1_LOC_737/A OR2X1_LOC_733/Y 0.16fF
C51265 OR2X1_LOC_737/A OR2X1_LOC_723/B 0.09fF
C55323 OR2X1_LOC_722/a_8_216# OR2X1_LOC_737/A 0.02fF
C56033 OR2X1_LOC_723/a_8_216# OR2X1_LOC_737/A 0.03fF
C56565 OR2X1_LOC_737/A VSS -1.19fF
C1344 OR2X1_LOC_475/Y OR2X1_LOC_805/A 0.01fF
C2358 OR2X1_LOC_475/Y OR2X1_LOC_228/Y 0.01fF
C4328 OR2X1_LOC_476/Y OR2X1_LOC_475/Y 0.06fF
C26440 OR2X1_LOC_475/Y OR2X1_LOC_479/a_8_216# 0.07fF
C26872 OR2X1_LOC_475/Y OR2X1_LOC_206/A 0.23fF
C30960 VDD OR2X1_LOC_475/Y 0.22fF
C42119 OR2X1_LOC_475/Y OR2X1_LOC_206/a_8_216# 0.14fF
C53311 OR2X1_LOC_475/Y OR2X1_LOC_215/A 0.14fF
C57210 OR2X1_LOC_475/Y VSS 0.45fF
C3936 OR2X1_LOC_453/Y OR2X1_LOC_466/a_8_216# 0.39fF
C21237 OR2X1_LOC_466/A OR2X1_LOC_453/Y 0.15fF
C46249 D_GATE_479 OR2X1_LOC_453/Y 0.01fF
C57323 OR2X1_LOC_453/Y VSS 0.17fF
C1472 OR2X1_LOC_479/Y OR2X1_LOC_365/B 0.03fF
C2968 OR2X1_LOC_182/a_8_216# OR2X1_LOC_365/B 0.12fF
C7766 OR2X1_LOC_808/B OR2X1_LOC_365/B 0.03fF
C10126 OR2X1_LOC_578/B OR2X1_LOC_365/B 0.06fF
C10691 OR2X1_LOC_357/a_8_216# OR2X1_LOC_365/B 0.01fF
C10730 VDD OR2X1_LOC_365/B 0.30fF
C13378 OR2X1_LOC_468/Y OR2X1_LOC_365/B 0.02fF
C14030 OR2X1_LOC_212/B OR2X1_LOC_365/B 0.36fF
C21779 OR2X1_LOC_364/B OR2X1_LOC_365/B 0.01fF
C23869 OR2X1_LOC_352/a_8_216# OR2X1_LOC_365/B 0.01fF
C24175 OR2X1_LOC_364/Y OR2X1_LOC_365/B 0.06fF
C31120 OR2X1_LOC_211/a_8_216# OR2X1_LOC_365/B 0.01fF
C33951 OR2X1_LOC_566/A OR2X1_LOC_365/B 0.02fF
C35096 OR2X1_LOC_365/a_8_216# OR2X1_LOC_365/B 0.07fF
C38442 OR2X1_LOC_566/Y OR2X1_LOC_365/B 0.01fF
C40276 OR2X1_LOC_357/B OR2X1_LOC_365/B 0.02fF
C41638 OR2X1_LOC_486/Y OR2X1_LOC_365/B 0.13fF
C44063 OR2X1_LOC_568/a_8_216# OR2X1_LOC_365/B 0.01fF
C46269 OR2X1_LOC_357/A OR2X1_LOC_365/B 0.02fF
C46282 OR2X1_LOC_367/B OR2X1_LOC_365/B 0.05fF
C47861 OR2X1_LOC_212/A OR2X1_LOC_365/B 0.02fF
C52228 OR2X1_LOC_566/a_8_216# OR2X1_LOC_365/B 0.01fF
C56253 OR2X1_LOC_365/B VSS 0.59fF
C17291 VDD AND2X1_LOC_649/B 0.23fF
C18213 AND2X1_LOC_649/B AND2X1_LOC_642/Y 0.01fF
C34713 AND2X1_LOC_649/B AND2X1_LOC_649/a_8_24# 0.01fF
C35412 AND2X1_LOC_358/Y AND2X1_LOC_649/B 0.01fF
C47555 AND2X1_LOC_649/B AND2X1_LOC_786/Y 0.01fF
C53115 AND2X1_LOC_649/B AND2X1_LOC_219/Y 0.01fF
C56966 AND2X1_LOC_649/B VSS 0.18fF
C1153 AND2X1_LOC_486/Y AND2X1_LOC_469/B 0.22fF
C1185 AND2X1_LOC_486/Y AND2X1_LOC_733/Y 0.42fF
C3783 AND2X1_LOC_486/Y AND2X1_LOC_850/Y 0.10fF
C4620 AND2X1_LOC_486/Y AND2X1_LOC_806/A 0.01fF
C10097 AND2X1_LOC_486/Y AND2X1_LOC_570/Y 0.03fF
C16529 AND2X1_LOC_486/Y AND2X1_LOC_576/Y 0.10fF
C16802 AND2X1_LOC_486/Y AND2X1_LOC_244/A 0.03fF
C21563 AND2X1_LOC_486/Y AND2X1_LOC_477/Y 0.13fF
C23747 AND2X1_LOC_486/Y AND2X1_LOC_556/a_8_24# 0.06fF
C26561 AND2X1_LOC_486/Y AND2X1_LOC_786/Y 0.07fF
C26776 AND2X1_LOC_486/Y AND2X1_LOC_578/A 0.07fF
C30381 AND2X1_LOC_486/Y AND2X1_LOC_212/Y 0.07fF
C31298 AND2X1_LOC_486/Y AND2X1_LOC_471/Y 0.09fF
C34665 AND2X1_LOC_486/Y AND2X1_LOC_562/B 0.03fF
C36647 AND2X1_LOC_486/Y AND2X1_LOC_564/B 0.07fF
C39324 AND2X1_LOC_486/Y AND2X1_LOC_474/A 0.03fF
C40941 AND2X1_LOC_486/Y AND2X1_LOC_719/Y 0.10fF
C42766 AND2X1_LOC_486/Y AND2X1_LOC_858/B 0.10fF
C43432 AND2X1_LOC_486/Y AND2X1_LOC_222/Y 0.03fF
C44025 AND2X1_LOC_486/Y AND2X1_LOC_860/A 0.10fF
C47114 AND2X1_LOC_486/Y AND2X1_LOC_476/Y 0.07fF
C50758 AND2X1_LOC_486/Y AND2X1_LOC_477/A 0.06fF
C51916 AND2X1_LOC_486/Y AND2X1_LOC_859/Y 0.10fF
C52497 AND2X1_LOC_486/Y AND2X1_LOC_657/A 0.10fF
C52615 AND2X1_LOC_486/Y AND2X1_LOC_794/B 0.01fF
C52643 AND2X1_LOC_486/Y VDD 1.60fF
C58047 AND2X1_LOC_486/Y VSS 0.35fF
C387 VDD AND2X1_LOC_523/Y 0.37fF
C7085 AND2X1_LOC_560/a_8_24# AND2X1_LOC_523/Y 0.01fF
C12634 AND2X1_LOC_571/A AND2X1_LOC_523/Y 0.03fF
C20505 AND2X1_LOC_576/Y AND2X1_LOC_523/Y 0.01fF
C22776 AND2X1_LOC_866/A AND2X1_LOC_523/Y 0.03fF
C26407 AND2X1_LOC_560/B AND2X1_LOC_523/Y 1.20fF
C36190 AND2X1_LOC_851/B AND2X1_LOC_523/Y 0.09fF
C40177 AND2X1_LOC_181/Y AND2X1_LOC_523/Y 0.03fF
C47738 AND2X1_LOC_367/A AND2X1_LOC_523/Y 0.46fF
C57095 AND2X1_LOC_523/Y VSS -0.64fF
C1770 AND2X1_LOC_578/A AND2X1_LOC_565/Y 0.01fF
C8065 AND2X1_LOC_736/Y AND2X1_LOC_565/Y 0.14fF
C27502 VDD AND2X1_LOC_565/Y 0.04fF
C29740 AND2X1_LOC_569/A AND2X1_LOC_565/Y 0.06fF
C53226 AND2X1_LOC_580/A AND2X1_LOC_565/Y 0.01fF
C57683 AND2X1_LOC_565/Y VSS 0.12fF
C12428 OR2X1_LOC_725/A OR2X1_LOC_725/a_8_216# 0.39fF
C28694 OR2X1_LOC_725/B OR2X1_LOC_725/A 0.07fF
C47501 VDD OR2X1_LOC_725/A -0.00fF
C56518 OR2X1_LOC_725/A VSS 0.18fF
C713 AND2X1_LOC_352/B AND2X1_LOC_662/B 0.82fF
C5299 AND2X1_LOC_364/Y AND2X1_LOC_352/B 0.04fF
C25324 VDD AND2X1_LOC_352/B 0.11fF
C31030 AND2X1_LOC_352/B AND2X1_LOC_863/Y 0.02fF
C37085 AND2X1_LOC_566/B AND2X1_LOC_352/B 0.01fF
C40116 AND2X1_LOC_352/B AND2X1_LOC_654/Y 0.09fF
C42691 AND2X1_LOC_212/A AND2X1_LOC_352/B 0.05fF
C49317 AND2X1_LOC_365/A AND2X1_LOC_352/B 0.11fF
C57410 AND2X1_LOC_352/B VSS 0.14fF
C10801 AND2X1_LOC_208/Y AND2X1_LOC_214/a_8_24# 0.02fF
C21879 AND2X1_LOC_208/Y AND2X1_LOC_219/A 0.16fF
C26545 AND2X1_LOC_214/A AND2X1_LOC_208/Y 0.04fF
C28622 VDD AND2X1_LOC_208/Y 0.02fF
C32812 AND2X1_LOC_208/Y AND2X1_LOC_214/a_36_24# 0.01fF
C56406 AND2X1_LOC_208/Y VSS 0.10fF
C2859 AND2X1_LOC_203/Y AND2X1_LOC_215/A 0.01fF
C19206 VDD AND2X1_LOC_203/Y 0.25fF
C53480 AND2X1_LOC_203/Y AND2X1_LOC_205/a_8_24# 0.19fF
C56320 AND2X1_LOC_203/Y VSS 0.10fF
C704 AND2X1_LOC_358/Y AND2X1_LOC_211/B 0.04fF
C936 AND2X1_LOC_211/B AND2X1_LOC_650/a_8_24# 0.01fF
C1720 AND2X1_LOC_211/B AND2X1_LOC_357/a_8_24# 0.04fF
C4779 AND2X1_LOC_211/B AND2X1_LOC_866/A 0.07fF
C5112 AND2X1_LOC_211/B AND2X1_LOC_857/a_8_24# 0.01fF
C6205 AND2X1_LOC_364/a_8_24# AND2X1_LOC_211/B 0.01fF
C7215 AND2X1_LOC_211/B AND2X1_LOC_364/A 0.31fF
C10968 AND2X1_LOC_357/B AND2X1_LOC_211/B 0.07fF
C11985 AND2X1_LOC_211/B AND2X1_LOC_853/a_8_24# 0.01fF
C13539 AND2X1_LOC_182/A AND2X1_LOC_211/B 0.11fF
C14094 AND2X1_LOC_211/B AND2X1_LOC_662/B 0.07fF
C14982 AND2X1_LOC_211/B AND2X1_LOC_211/a_36_24# 0.01fF
C17302 AND2X1_LOC_350/B AND2X1_LOC_211/B 0.89fF
C19079 AND2X1_LOC_568/B AND2X1_LOC_211/B 0.01fF
C19633 AND2X1_LOC_211/B AND2X1_LOC_650/Y 0.01fF
C22076 AND2X1_LOC_357/A AND2X1_LOC_211/B 0.02fF
C22498 AND2X1_LOC_181/Y AND2X1_LOC_211/B 0.03fF
C22633 AND2X1_LOC_228/Y AND2X1_LOC_211/B 0.01fF
C23013 AND2X1_LOC_211/B AND2X1_LOC_857/Y 0.04fF
C27234 AND2X1_LOC_211/B AND2X1_LOC_655/A 0.10fF
C29684 AND2X1_LOC_367/A AND2X1_LOC_211/B 0.07fF
C33425 AND2X1_LOC_182/a_8_24# AND2X1_LOC_211/B 0.02fF
C38501 VDD AND2X1_LOC_211/B 0.94fF
C40338 AND2X1_LOC_211/B AND2X1_LOC_640/Y 0.11fF
C46010 AND2X1_LOC_211/B AND2X1_LOC_641/Y 0.01fF
C50338 AND2X1_LOC_211/B AND2X1_LOC_852/Y 0.02fF
C50598 AND2X1_LOC_566/B AND2X1_LOC_211/B 0.03fF
C54529 AND2X1_LOC_211/B AND2X1_LOC_211/a_8_24# 0.03fF
C55826 AND2X1_LOC_211/B AND2X1_LOC_853/Y 0.44fF
C57573 AND2X1_LOC_211/B VSS 0.20fF
C16773 AND2X1_LOC_784/Y AND2X1_LOC_796/a_8_24# 0.11fF
C22679 AND2X1_LOC_784/Y AND2X1_LOC_222/Y 0.01fF
C28543 AND2X1_LOC_784/Y AND2X1_LOC_796/A 0.02fF
C29298 AND2X1_LOC_784/Y AND2X1_LOC_810/Y 0.01fF
C31623 AND2X1_LOC_784/Y VDD 0.40fF
C36259 AND2X1_LOC_784/Y AND2X1_LOC_469/B 0.02fF
C36602 AND2X1_LOC_784/Y AND2X1_LOC_804/A 0.26fF
C48629 AND2X1_LOC_784/Y AND2X1_LOC_804/a_8_24# 0.20fF
C58121 AND2X1_LOC_784/Y VSS -0.03fF
C20736 AND2X1_LOC_563/a_8_24# AND2X1_LOC_563/A 0.10fF
C23530 AND2X1_LOC_563/A AND2X1_LOC_657/A 0.07fF
C49772 AND2X1_LOC_563/A AND2X1_LOC_560/B 0.01fF
C57956 AND2X1_LOC_563/A VSS 0.15fF
C5136 AND2X1_LOC_640/Y AND2X1_LOC_641/Y 0.23fF
C9467 AND2X1_LOC_640/Y AND2X1_LOC_852/Y 2.74fF
C13579 AND2X1_LOC_215/Y AND2X1_LOC_640/Y 0.01fF
C16231 AND2X1_LOC_640/Y AND2X1_LOC_650/a_8_24# 0.04fF
C47179 AND2X1_LOC_640/Y AND2X1_LOC_219/A 0.17fF
C53990 VDD AND2X1_LOC_640/Y 0.13fF
C57161 AND2X1_LOC_640/Y VSS 0.37fF
C3716 OR2X1_LOC_624/Y OR2X1_LOC_658/a_36_216# 0.03fF
C9251 OR2X1_LOC_624/Y OR2X1_LOC_659/A 0.14fF
C11703 OR2X1_LOC_624/Y OR2X1_LOC_576/A 0.03fF
C31309 OR2X1_LOC_861/a_8_216# OR2X1_LOC_624/Y 0.02fF
C32920 OR2X1_LOC_624/Y OR2X1_LOC_244/Y 0.02fF
C36744 OR2X1_LOC_861/a_36_216# OR2X1_LOC_624/Y 0.03fF
C38940 OR2X1_LOC_624/Y OR2X1_LOC_659/a_8_216# 0.40fF
C42346 OR2X1_LOC_865/B OR2X1_LOC_624/Y 0.02fF
C50507 VDD OR2X1_LOC_624/Y 0.14fF
C54227 OR2X1_LOC_624/Y OR2X1_LOC_474/B 0.02fF
C54303 OR2X1_LOC_624/Y OR2X1_LOC_658/a_8_216# 0.02fF
C57338 OR2X1_LOC_624/Y VSS 0.34fF
C392 OR2X1_LOC_214/B OR2X1_LOC_214/A 0.06fF
C39279 OR2X1_LOC_214/a_8_216# OR2X1_LOC_214/A 0.39fF
C49885 OR2X1_LOC_214/A OR2X1_LOC_228/Y 0.10fF
C56733 OR2X1_LOC_214/A VSS 0.02fF
C46960 OR2X1_LOC_352/A OR2X1_LOC_578/B 0.01fF
C47571 OR2X1_LOC_352/A VDD -0.00fF
C50872 OR2X1_LOC_352/A OR2X1_LOC_212/B 0.19fF
C58029 OR2X1_LOC_352/A VSS 0.11fF
C181 AND2X1_LOC_218/Y AND2X1_LOC_786/Y 0.04fF
C302 AND2X1_LOC_578/A AND2X1_LOC_786/Y 0.07fF
C1543 AND2X1_LOC_662/B AND2X1_LOC_786/Y 0.07fF
C4858 AND2X1_LOC_471/Y AND2X1_LOC_786/Y 0.01fF
C5636 AND2X1_LOC_786/Y AND2X1_LOC_795/a_8_24# 0.08fF
C5685 AND2X1_LOC_219/Y AND2X1_LOC_786/Y 0.02fF
C5918 AND2X1_LOC_851/B AND2X1_LOC_786/Y 0.07fF
C9971 AND2X1_LOC_340/Y AND2X1_LOC_786/Y 2.01fF
C9981 AND2X1_LOC_181/Y AND2X1_LOC_786/Y 0.07fF
C10370 AND2X1_LOC_564/B AND2X1_LOC_786/Y 0.02fF
C11264 AND2X1_LOC_222/a_8_24# AND2X1_LOC_786/Y 0.05fF
C14659 AND2X1_LOC_719/Y AND2X1_LOC_786/Y 0.10fF
C15678 AND2X1_LOC_649/Y AND2X1_LOC_786/Y 0.01fF
C17055 AND2X1_LOC_222/Y AND2X1_LOC_786/Y 0.04fF
C17219 AND2X1_LOC_367/A AND2X1_LOC_786/Y 0.10fF
C20607 AND2X1_LOC_476/Y AND2X1_LOC_786/Y 0.04fF
C26111 VDD AND2X1_LOC_786/Y 1.35fF
C26750 AND2X1_LOC_660/A AND2X1_LOC_786/Y 0.07fF
C26993 AND2X1_LOC_642/Y AND2X1_LOC_786/Y 0.04fF
C37310 AND2X1_LOC_795/Y AND2X1_LOC_786/Y 0.01fF
C43566 AND2X1_LOC_649/a_8_24# AND2X1_LOC_786/Y 0.03fF
C48566 AND2X1_LOC_866/A AND2X1_LOC_786/Y 0.07fF
C50860 AND2X1_LOC_785/Y AND2X1_LOC_786/Y 0.02fF
C52163 AND2X1_LOC_717/Y AND2X1_LOC_786/Y 0.02fF
C56270 AND2X1_LOC_786/Y VSS -3.08fF
C6459 AND2X1_LOC_201/Y AND2X1_LOC_206/a_8_24# 0.07fF
C56277 AND2X1_LOC_201/Y VSS 0.13fF
C7115 OR2X1_LOC_471/Y OR2X1_LOC_731/A 0.07fF
C8975 OR2X1_LOC_471/Y OR2X1_LOC_741/Y 0.02fF
C18383 OR2X1_LOC_471/Y OR2X1_LOC_738/A 0.07fF
C20961 OR2X1_LOC_471/Y OR2X1_LOC_739/A 0.03fF
C23589 OR2X1_LOC_471/Y OR2X1_LOC_477/a_8_216# 0.07fF
C23614 OR2X1_LOC_471/Y OR2X1_LOC_223/A 0.03fF
C23936 OR2X1_LOC_471/Y OR2X1_LOC_213/A 0.80fF
C25518 OR2X1_LOC_471/Y OR2X1_LOC_742/a_8_216# 0.06fF
C26026 OR2X1_LOC_471/Y OR2X1_LOC_564/A 0.04fF
C36103 OR2X1_LOC_471/Y OR2X1_LOC_220/B 0.03fF
C40785 OR2X1_LOC_477/B OR2X1_LOC_471/Y 0.03fF
C48197 OR2X1_LOC_471/Y OR2X1_LOC_803/A 0.02fF
C54867 VDD OR2X1_LOC_471/Y 0.50fF
C57321 OR2X1_LOC_471/Y VSS -0.77fF
C2029 AND2X1_LOC_716/Y AND2X1_LOC_367/A 0.03fF
C5726 AND2X1_LOC_716/Y AND2X1_LOC_182/a_8_24# 0.02fF
C8496 AND2X1_LOC_716/Y AND2X1_LOC_723/a_36_24# 0.01fF
C10912 AND2X1_LOC_716/Y VDD -0.00fF
C22421 AND2X1_LOC_716/Y AND2X1_LOC_182/a_36_24# 0.01fF
C22870 AND2X1_LOC_716/Y AND2X1_LOC_566/B 1.18fF
C28290 AND2X1_LOC_716/Y AND2X1_LOC_212/A 0.04fF
C30065 AND2X1_LOC_716/Y AND2X1_LOC_357/a_8_24# 0.02fF
C33164 AND2X1_LOC_716/Y AND2X1_LOC_866/A 0.02fF
C34562 AND2X1_LOC_716/Y AND2X1_LOC_364/a_8_24# 0.01fF
C35537 AND2X1_LOC_716/Y AND2X1_LOC_364/A -0.03fF
C36763 AND2X1_LOC_716/Y AND2X1_LOC_717/Y 0.02fF
C39281 AND2X1_LOC_716/Y AND2X1_LOC_357/B 0.03fF
C41844 AND2X1_LOC_716/Y AND2X1_LOC_182/A 0.14fF
C42371 AND2X1_LOC_716/Y AND2X1_LOC_723/a_8_24# 0.11fF
C42390 AND2X1_LOC_716/Y AND2X1_LOC_662/B 0.02fF
C42782 AND2X1_LOC_723/Y AND2X1_LOC_716/Y 0.03fF
C47160 AND2X1_LOC_716/Y AND2X1_LOC_364/Y 0.03fF
C50528 AND2X1_LOC_716/Y AND2X1_LOC_357/A 0.02fF
C50940 AND2X1_LOC_716/Y AND2X1_LOC_181/Y 0.02fF
C55701 AND2X1_LOC_716/Y AND2X1_LOC_655/A 0.10fF
C57974 AND2X1_LOC_716/Y VSS -5.02fF
C7868 VDD AND2X1_LOC_566/B 0.01fF
C13633 AND2X1_LOC_566/B AND2X1_LOC_863/Y 0.09fF
C19023 AND2X1_LOC_170/Y AND2X1_LOC_566/B 0.17fF
C22884 AND2X1_LOC_566/B AND2X1_LOC_654/Y 0.02fF
C23779 AND2X1_LOC_566/B AND2X1_LOC_211/a_8_24# 0.01fF
C24679 AND2X1_LOC_566/B AND2X1_LOC_864/a_8_24# 0.01fF
C25281 AND2X1_LOC_212/A AND2X1_LOC_566/B 0.02fF
C28317 AND2X1_LOC_566/B AND2X1_LOC_661/a_8_24# 0.01fF
C30152 AND2X1_LOC_566/B AND2X1_LOC_866/A 0.02fF
C31588 AND2X1_LOC_364/a_8_24# AND2X1_LOC_566/B 0.01fF
C32477 AND2X1_LOC_566/B AND2X1_LOC_364/A 0.01fF
C34707 AND2X1_LOC_566/B AND2X1_LOC_212/B 0.01fF
C35509 AND2X1_LOC_566/a_8_24# AND2X1_LOC_566/B 0.04fF
C36234 AND2X1_LOC_566/B AND2X1_LOC_357/B 0.02fF
C38788 AND2X1_LOC_182/A AND2X1_LOC_566/B 0.53fF
C39296 AND2X1_LOC_566/B AND2X1_LOC_662/B 0.02fF
C41761 AND2X1_LOC_566/B AND2X1_LOC_212/Y 0.02fF
C41775 AND2X1_LOC_352/a_8_24# AND2X1_LOC_566/B 0.01fF
C43990 AND2X1_LOC_566/B AND2X1_LOC_364/Y 0.12fF
C44397 AND2X1_LOC_568/B AND2X1_LOC_566/B 0.01fF
C46735 AND2X1_LOC_566/a_36_24# AND2X1_LOC_566/B 0.01fF
C47507 AND2X1_LOC_357/A AND2X1_LOC_566/B 0.02fF
C49666 AND2X1_LOC_566/B AND2X1_LOC_365/a_8_24# 0.01fF
C52653 AND2X1_LOC_566/B AND2X1_LOC_655/A 0.03fF
C55109 AND2X1_LOC_566/B AND2X1_LOC_367/A 0.02fF
C57793 AND2X1_LOC_566/B VSS -1.48fF
C18079 AND2X1_LOC_794/A AND2X1_LOC_794/a_8_24# 0.19fF
C18552 AND2X1_LOC_794/A AND2X1_LOC_794/B 0.11fF
C18582 AND2X1_LOC_794/A VDD 0.25fF
C23314 AND2X1_LOC_794/A AND2X1_LOC_469/B 0.01fF
C43599 AND2X1_LOC_794/A AND2X1_LOC_477/Y 0.02fF
C52619 AND2X1_LOC_794/A AND2X1_LOC_212/Y 0.03fF
C58046 AND2X1_LOC_794/A VSS -0.02fF
C4797 AND2X1_LOC_564/B AND2X1_LOC_785/Y 0.01fF
C6971 AND2X1_LOC_564/B AND2X1_LOC_663/A 0.10fF
C10524 AND2X1_LOC_564/B AND2X1_LOC_578/A 0.07fF
C15843 AND2X1_LOC_564/B AND2X1_LOC_795/a_8_24# 0.02fF
C16783 AND2X1_LOC_736/Y AND2X1_LOC_564/B 0.19fF
C23142 AND2X1_LOC_564/A AND2X1_LOC_564/B 0.02fF
C24837 AND2X1_LOC_719/Y AND2X1_LOC_564/B 0.10fF
C29479 AND2X1_LOC_564/B AND2X1_LOC_658/A 0.07fF
C30692 AND2X1_LOC_564/B AND2X1_LOC_476/Y 0.04fF
C36209 AND2X1_LOC_564/B VDD 0.70fF
C40865 AND2X1_LOC_564/B AND2X1_LOC_657/Y 0.10fF
C47728 AND2X1_LOC_564/B AND2X1_LOC_795/Y -0.00fF
C55494 AND2X1_LOC_564/B AND2X1_LOC_658/B 0.07fF
C57992 AND2X1_LOC_564/B VSS 0.19fF
C1055 OR2X1_LOC_436/Y OR2X1_LOC_468/a_8_216# 0.02fF
C12092 OR2X1_LOC_436/Y OR2X1_LOC_468/a_36_216# 0.03fF
C23877 VDD OR2X1_LOC_436/Y 0.19fF
C26446 OR2X1_LOC_436/Y OR2X1_LOC_468/Y 0.15fF
C57209 OR2X1_LOC_436/Y VSS 0.37fF
C2246 OR2X1_LOC_851/A OR2X1_LOC_223/A 0.01fF
C4783 OR2X1_LOC_851/A OR2X1_LOC_228/Y 0.02fF
C24283 OR2X1_LOC_851/A OR2X1_LOC_479/Y 0.03fF
C36288 OR2X1_LOC_851/B OR2X1_LOC_851/A 0.19fF
C47840 OR2X1_LOC_851/A OR2X1_LOC_804/A 0.01fF
C57906 OR2X1_LOC_851/A VSS 0.20fF
C54617 OR2X1_LOC_725/B OR2X1_LOC_725/a_8_216# 0.05fF
C56571 OR2X1_LOC_725/B VSS 0.21fF
C4383 VDD OR2X1_LOC_731/A 0.12fF
C24076 OR2X1_LOC_738/A OR2X1_LOC_731/A 0.40fF
C32748 OR2X1_LOC_731/B OR2X1_LOC_731/A 0.16fF
C56371 OR2X1_LOC_731/A VSS 0.36fF
C1852 OR2X1_LOC_212/a_8_216# OR2X1_LOC_357/A 0.40fF
C5119 OR2X1_LOC_357/B OR2X1_LOC_357/A 0.15fF
C12498 OR2X1_LOC_212/A OR2X1_LOC_357/A 0.14fF
C31466 OR2X1_LOC_357/a_8_216# OR2X1_LOC_357/A 0.18fF
C31517 VDD OR2X1_LOC_357/A 0.06fF
C34792 OR2X1_LOC_212/B OR2X1_LOC_357/A 0.85fF
C56384 OR2X1_LOC_357/A VSS 0.01fF
C3422 OR2X1_LOC_797/B OR2X1_LOC_797/A 0.11fF
C7104 OR2X1_LOC_797/B OR2X1_LOC_213/B 0.01fF
C10457 OR2X1_LOC_797/B VDD 0.19fF
C35488 OR2X1_LOC_797/B OR2X1_LOC_213/A 0.02fF
C43104 OR2X1_LOC_797/B OR2X1_LOC_797/a_8_216# 0.18fF
C57856 OR2X1_LOC_797/B VSS 0.38fF
C3739 OR2X1_LOC_170/Y OR2X1_LOC_568/a_8_216# 0.40fF
C11817 OR2X1_LOC_170/Y OR2X1_LOC_566/a_8_216# 0.01fF
C23543 OR2X1_LOC_808/B OR2X1_LOC_170/Y 0.02fF
C25805 OR2X1_LOC_170/Y OR2X1_LOC_568/A 0.22fF
C25814 OR2X1_LOC_170/Y OR2X1_LOC_578/B 0.01fF
C26414 VDD OR2X1_LOC_170/Y -0.00fF
C29022 OR2X1_LOC_468/Y OR2X1_LOC_170/Y 0.01fF
C49880 OR2X1_LOC_566/A OR2X1_LOC_170/Y 0.17fF
C54344 OR2X1_LOC_170/Y OR2X1_LOC_566/Y 0.34fF
C56438 OR2X1_LOC_170/Y VSS 0.30fF
C2261 OR2X1_LOC_795/B OR2X1_LOC_228/Y 0.01fF
C21701 OR2X1_LOC_479/Y OR2X1_LOC_795/B 0.02fF
C28528 OR2X1_LOC_795/a_8_216# OR2X1_LOC_795/B 0.39fF
C30810 VDD OR2X1_LOC_795/B -0.00fF
C55831 OR2X1_LOC_223/A OR2X1_LOC_795/B 0.01fF
C56780 OR2X1_LOC_795/B VSS 0.17fF
C4713 OR2X1_LOC_723/a_8_216# OR2X1_LOC_723/A 0.39fF
C10306 VDD OR2X1_LOC_723/A -0.00fF
C36583 OR2X1_LOC_805/A OR2X1_LOC_723/A 0.03fF
C56152 OR2X1_LOC_723/B OR2X1_LOC_723/A 0.08fF
C56325 OR2X1_LOC_723/A VSS 0.18fF
C32568 OR2X1_LOC_857/B OR2X1_LOC_654/A 0.03fF
C51887 VDD OR2X1_LOC_654/A 0.22fF
C57774 OR2X1_LOC_654/A VSS -0.15fF
C5402 AND2X1_LOC_555/Y AND2X1_LOC_866/A 0.05fF
C11660 AND2X1_LOC_555/Y AND2X1_LOC_363/Y 0.01fF
C21510 AND2X1_LOC_555/Y AND2X1_LOC_562/B 0.07fF
C23156 AND2X1_LOC_555/Y AND2X1_LOC_363/a_8_24# 0.01fF
C24101 AND2X1_LOC_555/Y AND2X1_LOC_348/Y 0.01fF
C31017 AND2X1_LOC_555/Y AND2X1_LOC_562/Y 0.01fF
C34528 AND2X1_LOC_555/Y AND2X1_LOC_360/a_8_24# 0.01fF
C35073 AND2X1_LOC_555/Y AND2X1_LOC_663/B 0.01fF
C39191 AND2X1_LOC_555/Y VDD 0.27fF
C43011 AND2X1_LOC_555/Y AND2X1_LOC_562/a_8_24# 0.01fF
C45690 AND2X1_LOC_555/Y AND2X1_LOC_363/B 0.01fF
C54275 AND2X1_LOC_555/Y GATE_366 0.03fF
C58037 AND2X1_LOC_555/Y VSS -0.36fF
C17613 OR2X1_LOC_851/B OR2X1_LOC_858/A 0.03fF
C44723 OR2X1_LOC_851/B OR2X1_LOC_723/B 0.17fF
C51747 OR2X1_LOC_851/B OR2X1_LOC_851/a_8_216# 0.05fF
C55080 OR2X1_LOC_851/B VDD 0.12fF
C57947 OR2X1_LOC_851/B VSS 0.16fF
C1773 VDD OR2X1_LOC_796/B -0.00fF
C21425 OR2X1_LOC_796/B OR2X1_LOC_784/Y 0.21fF
C32318 OR2X1_LOC_796/B OR2X1_LOC_796/a_8_216# 0.39fF
C56896 OR2X1_LOC_796/B VSS 0.17fF
C1144 AND2X1_LOC_737/Y AND2X1_LOC_658/B 0.03fF
C1348 AND2X1_LOC_658/B AND2X1_LOC_808/A 0.03fF
C1907 AND2X1_LOC_658/B AND2X1_LOC_727/B 0.06fF
C6004 AND2X1_LOC_658/B AND2X1_LOC_222/Y 0.03fF
C6635 AND2X1_LOC_573/a_8_24# AND2X1_LOC_658/B 0.01fF
C8375 AND2X1_LOC_658/B AND2X1_LOC_658/A 0.28fF
C9606 AND2X1_LOC_658/B AND2X1_LOC_476/Y 0.07fF
C15008 AND2X1_LOC_658/B AND2X1_LOC_657/A 0.37fF
C15115 AND2X1_LOC_658/B VDD 0.87fF
C18500 AND2X1_LOC_658/B AND2X1_LOC_469/a_8_24# 0.03fF
C19826 AND2X1_LOC_658/B AND2X1_LOC_657/Y 0.44fF
C19830 AND2X1_LOC_658/B AND2X1_LOC_469/B 0.03fF
C21512 AND2X1_LOC_658/B AND2X1_LOC_213/B 0.03fF
C22330 AND2X1_LOC_573/Y AND2X1_LOC_658/B 0.01fF
C22393 AND2X1_LOC_738/B AND2X1_LOC_658/B 0.07fF
C23363 AND2X1_LOC_658/B AND2X1_LOC_806/A 0.03fF
C24916 AND2X1_LOC_658/B AND2X1_LOC_865/A 0.23fF
C25331 AND2X1_LOC_658/B AND2X1_LOC_658/Y 0.37fF
C25352 AND2X1_LOC_658/B AND2X1_LOC_734/Y 0.14fF
C27871 AND2X1_LOC_658/B AND2X1_LOC_862/Y 0.06fF
C28670 AND2X1_LOC_501/Y AND2X1_LOC_658/B 0.03fF
C28676 AND2X1_LOC_658/B AND2X1_LOC_570/Y 0.03fF
C29757 AND2X1_LOC_658/B AND2X1_LOC_796/Y 0.07fF
C32554 AND2X1_LOC_658/B AND2X1_LOC_807/Y 0.02fF
C33358 AND2X1_LOC_658/B AND2X1_LOC_865/a_8_24# 0.18fF
C33949 AND2X1_LOC_658/B AND2X1_LOC_657/a_8_24# 0.04fF
C35107 AND2X1_LOC_658/B AND2X1_LOC_576/Y 0.07fF
C36279 AND2X1_LOC_658/B AND2X1_LOC_659/a_8_24# 0.01fF
C38873 AND2X1_LOC_658/B AND2X1_LOC_866/B 0.45fF
C39682 AND2X1_LOC_658/B AND2X1_LOC_735/a_8_24# 0.01fF
C40041 AND2X1_LOC_658/B AND2X1_LOC_477/Y 0.07fF
C40297 AND2X1_LOC_658/B GATE_811 0.03fF
C40604 AND2X1_LOC_658/B AND2X1_LOC_580/A 0.03fF
C41302 AND2X1_LOC_544/Y AND2X1_LOC_658/B 0.03fF
C41839 AND2X1_LOC_658/B AND2X1_LOC_663/A 0.01fF
C42269 AND2X1_LOC_658/B AND2X1_LOC_675/Y 0.09fF
C45442 AND2X1_LOC_658/B AND2X1_LOC_578/A 0.07fF
C46435 AND2X1_LOC_658/B AND2X1_LOC_803/a_8_24# 0.02fF
C47961 AND2X1_LOC_658/B AND2X1_LOC_658/a_8_24# 0.01fF
C47989 AND2X1_LOC_658/B AND2X1_LOC_735/Y 0.01fF
C49183 AND2X1_LOC_658/B AND2X1_LOC_212/Y 0.07fF
C52543 AND2X1_LOC_727/Y AND2X1_LOC_658/B 0.03fF
C57930 AND2X1_LOC_658/B VSS 0.41fF
C12654 VDD AND2X1_LOC_453/Y -0.00fF
C34759 AND2X1_LOC_453/Y AND2X1_LOC_454/Y 0.14fF
C56729 AND2X1_LOC_453/Y VSS 0.16fF
C20711 OR2X1_LOC_205/Y OR2X1_LOC_641/B 0.04fF
C26198 OR2X1_LOC_215/a_8_216# OR2X1_LOC_641/B 0.39fF
C32349 OR2X1_LOC_340/Y OR2X1_LOC_641/B 0.02fF
C37032 OR2X1_LOC_864/A OR2X1_LOC_641/B 0.01fF
C40027 OR2X1_LOC_215/A OR2X1_LOC_641/B 0.08fF
C45380 OR2X1_LOC_641/B OR2X1_LOC_228/Y 0.09fF
C56435 OR2X1_LOC_641/B VSS 0.31fF
C3138 AND2X1_LOC_348/Y AND2X1_LOC_866/A 0.68fF
C9318 AND2X1_LOC_363/Y AND2X1_LOC_348/Y 1.02fF
C20733 AND2X1_LOC_363/a_8_24# AND2X1_LOC_348/Y 0.01fF
C24706 AND2X1_LOC_348/Y AND2X1_LOC_359/B 0.47fF
C27986 AND2X1_LOC_367/A AND2X1_LOC_348/Y 0.08fF
C28373 AND2X1_LOC_348/Y AND2X1_LOC_860/A 0.03fF
C36759 VDD AND2X1_LOC_348/Y 0.04fF
C57415 AND2X1_LOC_348/Y VSS -0.03fF
C524 AND2X1_LOC_571/a_8_24# AND2X1_LOC_571/B 0.19fF
C6126 AND2X1_LOC_571/B AND2X1_LOC_572/Y 0.02fF
C6887 AND2X1_LOC_571/A AND2X1_LOC_571/B 0.10fF
C48187 AND2X1_LOC_571/B AND2X1_LOC_563/Y 0.01fF
C50719 AND2X1_LOC_571/B AND2X1_LOC_657/A 0.02fF
C50859 AND2X1_LOC_571/B VDD 0.24fF
C58077 AND2X1_LOC_571/B VSS 0.07fF
C3400 AND2X1_LOC_568/B AND2X1_LOC_212/B 0.01fF
C4155 AND2X1_LOC_566/a_8_24# AND2X1_LOC_568/B 0.01fF
C10444 AND2X1_LOC_568/B AND2X1_LOC_212/Y 0.01fF
C12583 AND2X1_LOC_568/B AND2X1_LOC_364/Y 0.09fF
C18108 AND2X1_LOC_568/B AND2X1_LOC_365/a_8_24# 0.01fF
C23686 AND2X1_LOC_568/B AND2X1_LOC_367/A 0.03fF
C30064 AND2X1_LOC_568/B AND2X1_LOC_661/A 0.67fF
C30545 AND2X1_LOC_568/B AND2X1_LOC_477/A 0.19fF
C32442 VDD AND2X1_LOC_568/B 0.59fF
C33659 AND2X1_LOC_568/B AND2X1_LOC_212/a_8_24# 0.02fF
C38149 AND2X1_LOC_568/B AND2X1_LOC_863/Y 0.01fF
C43682 AND2X1_LOC_170/Y AND2X1_LOC_568/B 0.02fF
C46313 AND2X1_LOC_568/B AND2X1_LOC_566/Y 0.04fF
C48546 AND2X1_LOC_568/B AND2X1_LOC_211/a_8_24# 0.01fF
C49449 AND2X1_LOC_568/B AND2X1_LOC_864/a_8_24# 0.02fF
C50062 AND2X1_LOC_212/A AND2X1_LOC_568/B 0.02fF
C54891 AND2X1_LOC_568/B AND2X1_LOC_866/A 0.02fF
C695 AND2X1_LOC_852/Y AND2X1_LOC_219/A 0.46fF
C7579 VDD AND2X1_LOC_852/Y 0.61fF
C23361 AND2X1_LOC_215/Y AND2X1_LOC_852/Y 0.13fF
C24731 AND2X1_LOC_852/Y AND2X1_LOC_853/Y 0.23fF
C56980 AND2X1_LOC_852/Y VSS -0.73fF
C5897 AND2X1_LOC_141/A AND2X1_LOC_361/A 0.04fF
C25561 AND2X1_LOC_656/Y AND2X1_LOC_141/A 0.09fF
C28723 AND2X1_LOC_141/a_8_24# AND2X1_LOC_141/A 0.10fF
C57123 AND2X1_LOC_141/A VSS 0.16fF
C15700 AND2X1_LOC_181/Y AND2X1_LOC_851/B 0.07fF
C26823 AND2X1_LOC_181/Y AND2X1_LOC_222/Y 0.02fF
C30336 AND2X1_LOC_181/Y AND2X1_LOC_476/Y 0.51fF
C30738 AND2X1_LOC_181/Y AND2X1_LOC_182/a_8_24# 0.11fF
C35835 AND2X1_LOC_181/Y VDD 0.21fF
C57833 AND2X1_LOC_181/Y VSS 0.25fF
C12044 AND2X1_LOC_202/Y AND2X1_LOC_206/a_8_24# 0.11fF
C26517 VDD AND2X1_LOC_202/Y 0.31fF
C56276 AND2X1_LOC_202/Y VSS 0.15fF
C2335 AND2X1_LOC_244/A AND2X1_LOC_244/a_8_24# 0.10fF
C3224 AND2X1_LOC_474/A AND2X1_LOC_244/A 1.37fF
C4817 AND2X1_LOC_719/Y AND2X1_LOC_244/A 0.05fF
C6529 AND2X1_LOC_858/B AND2X1_LOC_244/A 0.03fF
C7839 AND2X1_LOC_244/A AND2X1_LOC_860/A 0.05fF
C8148 AND2X1_LOC_244/A AND2X1_LOC_562/Y 0.06fF
C16194 AND2X1_LOC_244/A AND2X1_LOC_657/A 0.07fF
C16313 VDD AND2X1_LOC_244/A 0.28fF
C24525 AND2X1_LOC_244/A AND2X1_LOC_806/A 0.03fF
C36309 AND2X1_LOC_576/Y AND2X1_LOC_244/A 0.01fF
C52977 AND2X1_LOC_244/A AND2X1_LOC_243/Y 0.14fF
C56667 AND2X1_LOC_244/A VSS 0.30fF
C10360 OR2X1_LOC_359/A OR2X1_LOC_580/A 0.05fF
C38833 OR2X1_LOC_359/a_8_216# OR2X1_LOC_359/A 0.39fF
C53873 OR2X1_LOC_359/A VDD -0.00fF
C57998 OR2X1_LOC_359/A VSS 0.18fF
C3314 VDD AND2X1_LOC_850/Y 0.21fF
C11494 AND2X1_LOC_850/Y AND2X1_LOC_806/A 0.01fF
C46272 AND2X1_LOC_474/A AND2X1_LOC_850/Y 0.01fF
C49751 AND2X1_LOC_858/B AND2X1_LOC_850/Y 0.02fF
C50972 AND2X1_LOC_850/Y AND2X1_LOC_860/A 0.09fF
C51858 AND2X1_LOC_860/a_8_24# AND2X1_LOC_850/Y 0.02fF
C56935 AND2X1_LOC_850/Y VSS 0.20fF
C4076 OR2X1_LOC_602/Y OR2X1_LOC_645/a_8_216# 0.01fF
C15129 OR2X1_LOC_602/Y OR2X1_LOC_648/A 0.40fF
C52697 OR2X1_LOC_364/A OR2X1_LOC_602/Y 0.35fF
C57457 OR2X1_LOC_602/Y VSS 0.40fF
C16397 OR2X1_LOC_862/B OR2X1_LOC_862/A 0.56fF
C25296 OR2X1_LOC_862/a_8_216# OR2X1_LOC_862/A 0.08fF
C27956 OR2X1_LOC_812/B OR2X1_LOC_862/A 0.14fF
C30767 OR2X1_LOC_862/a_36_216# OR2X1_LOC_862/A 0.01fF
C36245 OR2X1_LOC_865/A OR2X1_LOC_862/A 0.03fF
C37975 VDD OR2X1_LOC_862/A 0.13fF
C41894 OR2X1_LOC_862/A OR2X1_LOC_561/Y 0.19fF
C57487 OR2X1_LOC_862/A VSS 0.08fF
C5107 AND2X1_LOC_474/A AND2X1_LOC_866/A 0.03fF
C19393 AND2X1_LOC_474/A AND2X1_LOC_243/Y 0.07fF
C24914 AND2X1_LOC_474/A AND2X1_LOC_244/a_8_24# 0.01fF
C27412 AND2X1_LOC_719/Y AND2X1_LOC_474/A 0.05fF
C29147 AND2X1_LOC_474/A AND2X1_LOC_858/B 0.05fF
C30003 AND2X1_LOC_367/A AND2X1_LOC_474/A 0.05fF
C30387 AND2X1_LOC_474/A AND2X1_LOC_860/A 0.01fF
C30658 AND2X1_LOC_474/A AND2X1_LOC_562/Y 0.03fF
C31276 AND2X1_LOC_474/A AND2X1_LOC_860/a_8_24# 0.08fF
C35056 AND2X1_LOC_366/A AND2X1_LOC_474/A 0.01fF
C38704 AND2X1_LOC_474/A AND2X1_LOC_657/A 0.01fF
C38841 VDD AND2X1_LOC_474/A 0.48fF
C47247 AND2X1_LOC_474/A AND2X1_LOC_806/A 1.73fF
C57399 AND2X1_LOC_474/A VSS -0.42fF
C6388 AND2X1_LOC_658/A AND2X1_LOC_792/Y 0.07fF
C9138 AND2X1_LOC_663/B AND2X1_LOC_792/Y 0.01fF
C10773 AND2X1_LOC_792/Y AND2X1_LOC_805/Y 0.01fF
C35378 AND2X1_LOC_866/A AND2X1_LOC_792/Y 0.01fF
C36950 AND2X1_LOC_866/B AND2X1_LOC_792/Y 0.06fF
C38726 AND2X1_LOC_580/A AND2X1_LOC_792/Y 0.07fF
C39924 AND2X1_LOC_792/Y AND2X1_LOC_663/A 0.10fF
C41391 AND2X1_LOC_792/Y AND2X1_LOC_793/Y 0.72fF
C44338 AND2X1_LOC_580/B AND2X1_LOC_792/Y 0.04fF
C47110 AND2X1_LOC_792/Y AND2X1_LOC_805/a_8_24# 0.04fF
C56826 AND2X1_LOC_792/Y VSS -2.90fF
C10539 VDD OR2X1_LOC_340/Y 0.20fF
C19555 OR2X1_LOC_341/Y OR2X1_LOC_340/Y 0.06fF
C36032 OR2X1_LOC_340/Y OR2X1_LOC_350/a_8_216# 0.07fF
C37854 OR2X1_LOC_340/Y OR2X1_LOC_228/Y 0.01fF
C38597 OR2X1_LOC_219/B OR2X1_LOC_340/Y 0.03fF
C56540 OR2X1_LOC_340/Y VSS 0.36fF
C24406 OR2X1_LOC_714/Y OR2X1_LOC_724/A 0.14fF
C54398 OR2X1_LOC_714/Y OR2X1_LOC_724/a_8_216# 0.39fF
C56516 OR2X1_LOC_714/Y VSS 0.17fF
C3934 OR2X1_LOC_479/Y OR2X1_LOC_787/Y 0.19fF
C10222 OR2X1_LOC_808/B OR2X1_LOC_787/Y 0.10fF
C13173 VDD OR2X1_LOC_787/Y 0.35fF
C37848 OR2X1_LOC_223/A OR2X1_LOC_787/Y 0.29fF
C41210 OR2X1_LOC_787/Y OR2X1_LOC_794/a_8_216# 0.02fF
C46910 OR2X1_LOC_787/Y OR2X1_LOC_794/a_36_216# 0.02fF
C56895 OR2X1_LOC_787/Y VSS 0.13fF
C14236 AND2X1_LOC_574/Y VDD 0.05fF
C21424 AND2X1_LOC_573/Y AND2X1_LOC_574/Y 0.01fF
C27773 AND2X1_LOC_574/Y AND2X1_LOC_501/Y 0.83fF
C27779 AND2X1_LOC_574/Y AND2X1_LOC_570/Y 0.01fF
C34175 AND2X1_LOC_574/Y AND2X1_LOC_576/Y 0.03fF
C41318 AND2X1_LOC_574/Y AND2X1_LOC_675/Y 0.05fF
C47032 AND2X1_LOC_574/Y AND2X1_LOC_735/Y 0.02fF
C57958 AND2X1_LOC_574/Y VSS 0.06fF
C56425 OR2X1_LOC_724/A VSS 0.40fF
C4300 VDD OR2X1_LOC_339/Y 0.12fF
C32364 OR2X1_LOC_219/B OR2X1_LOC_339/Y 0.03fF
C34626 OR2X1_LOC_339/Y OR2X1_LOC_358/A 0.06fF
C56479 OR2X1_LOC_339/Y VSS 0.14fF
C1256 VDD OR2X1_LOC_863/B 0.12fF
C3922 OR2X1_LOC_863/a_8_216# OR2X1_LOC_863/B 0.05fF
C8481 OR2X1_LOC_863/B OR2X1_LOC_863/A 0.07fF
C57671 OR2X1_LOC_863/B VSS 0.21fF
C8405 OR2X1_LOC_739/A OR2X1_LOC_740/B 0.03fF
C8991 OR2X1_LOC_479/Y OR2X1_LOC_739/A 0.03fF
C15215 OR2X1_LOC_808/B OR2X1_LOC_739/A 0.05fF
C18165 VDD OR2X1_LOC_739/A 0.49fF
C20594 OR2X1_LOC_739/A OR2X1_LOC_739/a_8_216# 0.18fF
C20859 OR2X1_LOC_468/Y OR2X1_LOC_739/A 0.03fF
C39387 OR2X1_LOC_220/A OR2X1_LOC_739/A 0.03fF
C49247 OR2X1_LOC_739/A OR2X1_LOC_486/Y 0.12fF
C56779 OR2X1_LOC_739/A VSS 0.34fF
C23671 AND2X1_LOC_367/A AND2X1_LOC_243/Y 0.10fF
C28420 AND2X1_LOC_663/B AND2X1_LOC_243/Y 0.10fF
C28680 AND2X1_LOC_366/A AND2X1_LOC_243/Y 0.02fF
C32431 VDD AND2X1_LOC_243/Y 1.16fF
C40601 AND2X1_LOC_243/Y AND2X1_LOC_806/A 0.03fF
C54880 AND2X1_LOC_866/A AND2X1_LOC_243/Y 0.07fF
C56563 AND2X1_LOC_243/Y VSS -2.09fF
C136 OR2X1_LOC_792/Y OR2X1_LOC_580/A 0.01fF
C1242 OR2X1_LOC_792/Y OR2X1_LOC_807/B 0.04fF
C10584 OR2X1_LOC_792/Y OR2X1_LOC_811/A 0.02fF
C12307 OR2X1_LOC_792/Y OR2X1_LOC_807/A 0.04fF
C14293 OR2X1_LOC_792/Y OR2X1_LOC_580/B 0.26fF
C15036 OR2X1_LOC_792/Y D_GATE_579 0.01fF
C25502 OR2X1_LOC_792/Y OR2X1_LOC_807/a_8_216# 0.02fF
C39375 OR2X1_LOC_807/Y OR2X1_LOC_792/Y 0.42fF
C46307 OR2X1_LOC_792/Y OR2X1_LOC_805/a_8_216# 0.02fF
C46315 OR2X1_LOC_792/Y OR2X1_LOC_362/B 0.05fF
C51895 OR2X1_LOC_792/Y OR2X1_LOC_806/a_8_216# 0.02fF
C54586 OR2X1_LOC_792/Y OR2X1_LOC_580/a_8_216# 0.02fF
C57425 OR2X1_LOC_792/Y VSS 0.10fF
C18664 OR2X1_LOC_523/Y OR2X1_LOC_560/a_8_216# 0.08fF
C34658 OR2X1_LOC_523/Y OR2X1_LOC_632/Y 0.13fF
C43189 OR2X1_LOC_523/Y OR2X1_LOC_244/Y 0.53fF
C55014 OR2X1_LOC_523/Y OR2X1_LOC_560/A 0.44fF
C56766 OR2X1_LOC_523/Y VSS 0.13fF
C21735 OR2X1_LOC_797/A OR2X1_LOC_797/a_8_216# 0.39fF
C56947 OR2X1_LOC_797/A VSS 0.18fF
C3589 OR2X1_LOC_215/Y OR2X1_LOC_228/Y 0.01fF
C5816 OR2X1_LOC_228/Y OR2X1_LOC_341/a_8_216# 0.03fF
C6402 OR2X1_LOC_351/B OR2X1_LOC_228/Y 0.33fF
C9558 OR2X1_LOC_358/B OR2X1_LOC_228/Y 0.02fF
C11391 OR2X1_LOC_228/Y OR2X1_LOC_341/a_36_216# 0.03fF
C13201 OR2X1_LOC_228/Y OR2X1_LOC_723/B 0.01fF
C14250 OR2X1_LOC_479/Y OR2X1_LOC_228/Y 0.01fF
C14638 OR2X1_LOC_219/a_8_216# OR2X1_LOC_228/Y 0.01fF
C18919 OR2X1_LOC_479/a_8_216# OR2X1_LOC_228/Y 0.01fF
C20679 OR2X1_LOC_218/Y OR2X1_LOC_228/Y 0.01fF
C21144 OR2X1_LOC_795/a_8_216# OR2X1_LOC_228/Y 0.01fF
C23528 VDD OR2X1_LOC_228/Y 0.62fF
C25662 OR2X1_LOC_222/A OR2X1_LOC_228/Y 0.01fF
C26165 OR2X1_LOC_222/a_8_216# OR2X1_LOC_228/Y 0.01fF
C32350 OR2X1_LOC_341/Y OR2X1_LOC_228/Y 0.03fF
C37575 OR2X1_LOC_804/A OR2X1_LOC_228/Y 1.17fF
C41233 OR2X1_LOC_648/A OR2X1_LOC_228/Y 0.02fF
C42768 OR2X1_LOC_351/a_8_216# OR2X1_LOC_228/Y 0.13fF
C48445 OR2X1_LOC_223/A OR2X1_LOC_228/Y 0.01fF
C49140 OR2X1_LOC_350/a_8_216# OR2X1_LOC_228/Y 0.01fF
C50014 OR2X1_LOC_805/A OR2X1_LOC_228/Y 0.07fF
C51700 OR2X1_LOC_219/B OR2X1_LOC_228/Y 0.02fF
C52988 OR2X1_LOC_476/Y OR2X1_LOC_228/Y 0.01fF
C53932 OR2X1_LOC_358/A OR2X1_LOC_228/Y 0.05fF
C56434 OR2X1_LOC_228/Y VSS 0.57fF
C4002 OR2X1_LOC_551/a_8_216# OR2X1_LOC_551/A 0.39fF
C52437 VDD OR2X1_LOC_551/A -0.00fF
C56398 OR2X1_LOC_551/A VSS 0.18fF
C1980 AND2X1_LOC_793/Y AND2X1_LOC_805/a_8_24# 0.05fF
C17483 AND2X1_LOC_658/A AND2X1_LOC_793/Y 0.07fF
C21847 AND2X1_LOC_793/Y AND2X1_LOC_805/Y 0.01fF
C24330 VDD AND2X1_LOC_793/Y 0.24fF
C48284 AND2X1_LOC_866/B AND2X1_LOC_793/Y 0.10fF
C50003 AND2X1_LOC_580/A AND2X1_LOC_793/Y 0.07fF
C51177 AND2X1_LOC_793/Y AND2X1_LOC_663/A 0.10fF
C55470 AND2X1_LOC_580/B AND2X1_LOC_793/Y 0.02fF
C56825 AND2X1_LOC_793/Y VSS 0.16fF
C2033 OR2X1_LOC_348/Y OR2X1_LOC_805/A 0.07fF
C2346 OR2X1_LOC_348/Y OR2X1_LOC_580/B 0.10fF
C14640 OR2X1_LOC_348/Y OR2X1_LOC_363/a_8_216# 0.02fF
C16796 OR2X1_LOC_348/Y OR2X1_LOC_359/a_8_216# 0.05fF
C26824 OR2X1_LOC_348/Y OR2X1_LOC_366/a_8_216# 0.03fF
C27839 OR2X1_LOC_348/Y OR2X1_LOC_363/B 0.12fF
C30808 OR2X1_LOC_348/Y OR2X1_LOC_363/A 0.01fF
C31155 OR2X1_LOC_348/Y OR2X1_LOC_366/A 0.03fF
C34213 OR2X1_LOC_348/Y OR2X1_LOC_362/B 0.01fF
C38767 OR2X1_LOC_348/Y OR2X1_LOC_366/B 0.27fF
C44308 OR2X1_LOC_348/Y OR2X1_LOC_580/A 0.59fF
C54737 OR2X1_LOC_348/Y OR2X1_LOC_811/A 0.10fF
C58032 OR2X1_LOC_348/Y VSS 0.24fF
C7447 VDD AND2X1_LOC_193/Y 0.25fF
C24451 AND2X1_LOC_193/Y AND2X1_LOC_194/Y 0.21fF
C35368 AND2X1_LOC_193/Y AND2X1_LOC_200/a_8_24# 0.19fF
C56557 AND2X1_LOC_193/Y VSS 0.10fF
C12483 OR2X1_LOC_561/Y OR2X1_LOC_580/A 0.35fF
C34185 OR2X1_LOC_862/B OR2X1_LOC_561/Y 0.01fF
C43089 OR2X1_LOC_862/a_8_216# OR2X1_LOC_561/Y 0.39fF
C45818 OR2X1_LOC_812/B OR2X1_LOC_561/Y 0.01fF
C47890 OR2X1_LOC_561/Y OR2X1_LOC_579/A 0.01fF
C52062 OR2X1_LOC_561/Y OR2X1_LOC_579/a_8_216# 0.01fF
C56767 OR2X1_LOC_561/Y VSS 0.28fF
C7832 AND2X1_LOC_477/Y AND2X1_LOC_727/B 0.11fF
C9602 AND2X1_LOC_663/A AND2X1_LOC_727/B 0.73fF
C16736 AND2X1_LOC_212/Y AND2X1_LOC_727/B 0.08fF
C20150 AND2X1_LOC_727/Y AND2X1_LOC_727/B 0.01fF
C25095 AND2X1_LOC_808/A AND2X1_LOC_727/B 0.53fF
C28286 AND2X1_LOC_804/Y AND2X1_LOC_727/B 0.03fF
C31980 AND2X1_LOC_658/A AND2X1_LOC_727/B 0.09fF
C33769 AND2X1_LOC_808/a_8_24# AND2X1_LOC_727/B 0.19fF
C38786 VDD AND2X1_LOC_727/B 0.31fF
C39265 AND2X1_LOC_811/B AND2X1_LOC_727/B 0.09fF
C41991 AND2X1_LOC_811/Y AND2X1_LOC_727/B 0.02fF
C43523 AND2X1_LOC_657/Y AND2X1_LOC_727/B 0.01fF
C43528 AND2X1_LOC_469/B AND2X1_LOC_727/B 0.03fF
C56574 AND2X1_LOC_727/B VSS 0.16fF
C21940 AND2X1_LOC_216/Y AND2X1_LOC_217/Y 0.01fF
C27395 AND2X1_LOC_216/Y AND2X1_LOC_218/a_8_24# 0.18fF
C34146 AND2X1_LOC_216/Y VDD 0.21fF
C34818 AND2X1_LOC_216/Y AND2X1_LOC_660/A 0.01fF
C58138 AND2X1_LOC_216/Y VSS 0.06fF
C880 AND2X1_LOC_656/Y AND2X1_LOC_218/Y 0.01fF
C4678 AND2X1_LOC_141/a_8_24# AND2X1_LOC_656/Y 0.23fF
C6965 AND2X1_LOC_656/Y AND2X1_LOC_660/a_8_24# 0.04fF
C14480 AND2X1_LOC_217/Y AND2X1_LOC_656/Y 3.33fF
C20022 AND2X1_LOC_218/a_8_24# AND2X1_LOC_656/Y 0.01fF
C22769 AND2X1_LOC_656/Y AND2X1_LOC_663/B 0.08fF
C26574 AND2X1_LOC_656/Y AND2X1_LOC_657/A 0.11fF
C26782 VDD AND2X1_LOC_656/Y 0.40fF
C37823 AND2X1_LOC_656/Y AND2X1_LOC_361/A 0.07fF
C52910 AND2X1_LOC_560/B AND2X1_LOC_656/Y 0.03fF
C57216 AND2X1_LOC_656/Y VSS 0.08fF
C20981 OR2X1_LOC_476/Y OR2X1_LOC_479/a_8_216# 0.39fF
C50442 OR2X1_LOC_476/Y OR2X1_LOC_223/A 0.01fF
C57211 OR2X1_LOC_476/Y VSS 0.18fF
C2355 OR2X1_LOC_363/A OR2X1_LOC_366/B 0.27fF
C2719 OR2X1_LOC_366/B OR2X1_LOC_366/A 0.08fF
C3198 VDD OR2X1_LOC_366/B 0.06fF
C15774 OR2X1_LOC_366/B OR2X1_LOC_580/A 0.02fF
C26154 OR2X1_LOC_811/A OR2X1_LOC_366/B 0.03fF
C42131 OR2X1_LOC_366/B OR2X1_LOC_363/a_8_216# 0.40fF
C55511 OR2X1_LOC_363/B OR2X1_LOC_366/B 0.11fF
C56482 OR2X1_LOC_366/B VSS 0.32fF
C2010 OR2X1_LOC_575/A OR2X1_LOC_244/Y 0.02fF
C11445 OR2X1_LOC_575/A OR2X1_LOC_573/Y 0.12fF
C19430 VDD OR2X1_LOC_575/A 0.33fF
C49203 OR2X1_LOC_575/A OR2X1_LOC_563/A 0.02fF
C49736 OR2X1_LOC_575/A OR2X1_LOC_632/Y 0.40fF
C56593 OR2X1_LOC_575/A VSS -0.05fF
C20299 OR2X1_LOC_812/B OR2X1_LOC_862/B 0.12fF
C29089 OR2X1_LOC_862/a_8_216# OR2X1_LOC_812/B 0.01fF
C29137 OR2X1_LOC_812/B OR2X1_LOC_812/a_8_216# 0.04fF
C40055 OR2X1_LOC_865/A OR2X1_LOC_812/B 0.71fF
C40096 OR2X1_LOC_812/B D_GATE_811 0.03fF
C41888 VDD OR2X1_LOC_812/B 0.07fF
C54429 OR2X1_LOC_812/B OR2X1_LOC_812/A 0.06fF
C57803 OR2X1_LOC_812/B VSS -0.51fF
C5577 OR2X1_LOC_244/A OR2X1_LOC_204/Y 0.03fF
C19187 OR2X1_LOC_141/B OR2X1_LOC_204/Y 0.20fF
C28703 OR2X1_LOC_204/Y OR2X1_LOC_267/Y 0.05fF
C32618 OR2X1_LOC_663/A OR2X1_LOC_204/Y 0.03fF
C39894 OR2X1_LOC_204/Y OR2X1_LOC_124/Y 0.24fF
C52829 OR2X1_LOC_864/A OR2X1_LOC_204/Y 0.03fF
C56899 OR2X1_LOC_204/Y VSS 0.44fF
C34670 OR2X1_LOC_719/Y OR2X1_LOC_733/A 0.21fF
C56618 OR2X1_LOC_719/Y VSS 0.29fF
C5678 OR2X1_LOC_351/B OR2X1_LOC_648/B 0.10fF
C14467 OR2X1_LOC_648/B OR2X1_LOC_648/a_8_216# 0.01fF
C22841 VDD OR2X1_LOC_648/B 0.88fF
C25494 OR2X1_LOC_648/B OR2X1_LOC_655/B 0.15fF
C40507 OR2X1_LOC_648/B OR2X1_LOC_648/A 0.19fF
C57520 OR2X1_LOC_648/B VSS 0.62fF
C1617 VDD OR2X1_LOC_194/Y 0.11fF
C23875 OR2X1_LOC_194/Y OR2X1_LOC_200/a_8_216# 0.06fF
C27046 OR2X1_LOC_207/B OR2X1_LOC_194/Y 0.03fF
C57150 OR2X1_LOC_194/Y VSS 0.05fF
C2042 OR2X1_LOC_223/A OR2X1_LOC_181/Y 0.01fF
C12770 OR2X1_LOC_181/Y OR2X1_LOC_367/B 0.80fF
C33228 VDD OR2X1_LOC_181/Y 0.19fF
C56431 OR2X1_LOC_181/Y VSS 0.10fF
C11152 OR2X1_LOC_649/B OR2X1_LOC_649/a_8_216# 0.06fF
C15286 OR2X1_LOC_649/B OR2X1_LOC_660/B 0.72fF
C21835 OR2X1_LOC_649/B OR2X1_LOC_655/B 0.04fF
C22260 OR2X1_LOC_649/B OR2X1_LOC_655/A 0.03fF
C36457 OR2X1_LOC_662/A OR2X1_LOC_649/B 0.16fF
C54862 OR2X1_LOC_649/B OR2X1_LOC_655/a_8_216# 0.02fF
C57652 OR2X1_LOC_649/B VSS 0.14fF
C6174 AND2X1_LOC_722/A AND2X1_LOC_436/Y 0.03fF
C15758 AND2X1_LOC_722/A AND2X1_LOC_810/Y 0.07fF
C16181 AND2X1_LOC_722/A AND2X1_LOC_477/A 0.03fF
C18089 AND2X1_LOC_794/B AND2X1_LOC_722/A 0.07fF
C18119 VDD AND2X1_LOC_722/A 0.10fF
C25359 AND2X1_LOC_738/B AND2X1_LOC_722/A 0.07fF
C38891 AND2X1_LOC_722/Y AND2X1_LOC_722/A 0.04fF
C48578 AND2X1_LOC_578/A AND2X1_LOC_722/A 0.10fF
C50152 AND2X1_LOC_723/Y AND2X1_LOC_722/A 0.01fF
C52156 AND2X1_LOC_722/A AND2X1_LOC_212/Y 0.07fF
C57627 AND2X1_LOC_722/A VSS 0.29fF
C5175 AND2X1_LOC_192/Y GATE_811 0.09fF
C7247 AND2X1_LOC_192/Y AND2X1_LOC_220/Y 0.12fF
C9727 AND2X1_LOC_803/B AND2X1_LOC_192/Y 0.03fF
C16028 AND2X1_LOC_192/Y AND2X1_LOC_480/A 0.08fF
C16395 AND2X1_LOC_741/Y AND2X1_LOC_192/Y 0.14fF
C22018 AND2X1_LOC_742/a_8_24# AND2X1_LOC_192/Y 0.02fF
C31018 AND2X1_LOC_192/Y AND2X1_LOC_739/a_8_24# 0.03fF
C31859 AND2X1_LOC_192/Y AND2X1_LOC_797/A 0.09fF
C35946 VDD AND2X1_LOC_192/Y 0.35fF
C36476 AND2X1_LOC_192/Y AND2X1_LOC_740/B 0.03fF
C49173 AND2X1_LOC_192/Y AND2X1_LOC_742/A 0.13fF
C54777 AND2X1_LOC_797/a_8_24# AND2X1_LOC_192/Y 0.02fF
C57693 AND2X1_LOC_192/Y VSS 0.24fF
C35355 AND2X1_LOC_475/Y AND2X1_LOC_476/Y 0.05fF
C40875 AND2X1_LOC_475/Y AND2X1_LOC_479/a_8_24# 0.09fF
C40884 VDD AND2X1_LOC_475/Y 0.21fF
C56629 AND2X1_LOC_475/Y VSS 0.20fF
C643 AND2X1_LOC_734/Y AND2X1_LOC_476/Y 0.07fF
C6166 VDD AND2X1_LOC_734/Y 0.05fF
C10907 AND2X1_LOC_734/Y AND2X1_LOC_657/Y 0.03fF
C23786 AND2X1_LOC_734/Y AND2X1_LOC_807/Y 0.09fF
C27486 AND2X1_LOC_734/Y AND2X1_LOC_737/a_8_24# 0.01fF
C32411 AND2X1_LOC_544/Y AND2X1_LOC_734/Y 0.14fF
C32946 AND2X1_LOC_734/Y AND2X1_LOC_663/A 1.17fF
C48500 AND2X1_LOC_737/Y AND2X1_LOC_734/Y 0.07fF
C53318 AND2X1_LOC_734/Y AND2X1_LOC_222/Y 0.18fF
C55580 AND2X1_LOC_734/Y AND2X1_LOC_658/A 0.07fF
C57824 AND2X1_LOC_734/Y VSS 0.27fF
C8552 AND2X1_LOC_654/Y AND2X1_LOC_661/A 0.09fF
C10936 AND2X1_LOC_212/A AND2X1_LOC_661/A 0.02fF
C17417 AND2X1_LOC_365/A AND2X1_LOC_661/A 0.18fF
C29663 AND2X1_LOC_364/Y AND2X1_LOC_661/A 0.02fF
C35139 AND2X1_LOC_365/a_8_24# AND2X1_LOC_661/A 0.09fF
C37633 AND2X1_LOC_661/A AND2X1_LOC_436/Y 1.09fF
C47419 AND2X1_LOC_810/Y AND2X1_LOC_661/A 0.02fF
C49779 VDD AND2X1_LOC_661/A 0.42fF
C55426 AND2X1_LOC_863/Y AND2X1_LOC_661/A 0.02fF
C57006 AND2X1_LOC_661/A VSS 0.33fF
C623 AND2X1_LOC_794/B AND2X1_LOC_469/B 0.22fF
C3234 AND2X1_LOC_738/B AND2X1_LOC_794/B 0.03fF
C21038 AND2X1_LOC_794/B AND2X1_LOC_477/Y 0.01fF
C26255 AND2X1_LOC_794/B AND2X1_LOC_578/A 0.05fF
C29895 AND2X1_LOC_794/B AND2X1_LOC_212/Y 0.01fF
C30787 AND2X1_LOC_794/B AND2X1_LOC_471/Y 0.01fF
C40040 AND2X1_LOC_794/B AND2X1_LOC_436/Y 0.05fF
C41822 AND2X1_LOC_794/B AND2X1_LOC_477/a_8_24# 0.01fF
C49854 AND2X1_LOC_794/B AND2X1_LOC_810/Y 0.07fF
C50240 AND2X1_LOC_794/B AND2X1_LOC_477/A 0.01fF
C51681 AND2X1_LOC_794/B AND2X1_LOC_794/a_8_24# 0.02fF
C52129 AND2X1_LOC_794/B VDD 0.38fF
C58003 AND2X1_LOC_794/B VSS 0.19fF
C9232 AND2X1_LOC_341/a_8_24# AND2X1_LOC_228/Y 0.03fF
C17018 AND2X1_LOC_228/Y AND2X1_LOC_650/Y 0.46fF
C20270 AND2X1_LOC_341/a_36_24# AND2X1_LOC_228/Y 0.01fF
C20366 AND2X1_LOC_228/Y AND2X1_LOC_857/Y 0.03fF
C33553 AND2X1_LOC_228/Y AND2X1_LOC_654/a_8_24# 0.01fF
C35936 VDD AND2X1_LOC_228/Y -0.00fF
C43361 AND2X1_LOC_228/Y AND2X1_LOC_641/Y 0.08fF
C57759 AND2X1_LOC_228/Y VSS 0.38fF
C17815 AND2X1_LOC_470/A AND2X1_LOC_470/B 0.09fF
C22234 AND2X1_LOC_470/a_8_24# AND2X1_LOC_470/B 0.01fF
C33168 AND2X1_LOC_477/A AND2X1_LOC_470/B 0.83fF
C35086 VDD AND2X1_LOC_470/B 0.02fF
C56673 AND2X1_LOC_470/B VSS 0.08fF
C4943 OR2X1_LOC_805/A OR2X1_LOC_244/Y 0.03fF
C10651 OR2X1_LOC_358/a_8_216# OR2X1_LOC_805/A 0.05fF
C12096 OR2X1_LOC_805/A OR2X1_LOC_723/B 0.09fF
C16883 OR2X1_LOC_805/A OR2X1_LOC_723/a_8_216# 0.04fF
C18256 OR2X1_LOC_807/Y OR2X1_LOC_805/A 0.02fF
C18616 OR2X1_LOC_363/B OR2X1_LOC_805/A 0.03fF
C19686 OR2X1_LOC_218/Y OR2X1_LOC_805/A 0.09fF
C22474 OR2X1_LOC_805/A OR2X1_LOC_723/a_36_216# 0.01fF
C22482 VDD OR2X1_LOC_805/A 1.20fF
C25061 OR2X1_LOC_362/B OR2X1_LOC_805/A 0.30fF
C25191 OR2X1_LOC_222/a_8_216# OR2X1_LOC_805/A 0.04fF
C27907 OR2X1_LOC_805/A OR2X1_LOC_733/A 0.03fF
C29659 OR2X1_LOC_805/A OR2X1_LOC_736/A 0.03fF
C34983 OR2X1_LOC_805/A OR2X1_LOC_580/A 0.07fF
C39451 OR2X1_LOC_216/Y OR2X1_LOC_805/A 0.12fF
C40144 OR2X1_LOC_648/A OR2X1_LOC_805/A 0.07fF
C41031 OR2X1_LOC_858/A OR2X1_LOC_805/A 0.03fF
C44676 OR2X1_LOC_805/A OR2X1_LOC_215/A 0.03fF
C45450 OR2X1_LOC_811/A OR2X1_LOC_805/A 0.30fF
C52170 OR2X1_LOC_805/A OR2X1_LOC_563/A 0.07fF
C56943 OR2X1_LOC_805/A VSS -2.11fF
C24409 VDD OR2X1_LOC_731/B -0.00fF
C38778 OR2X1_LOC_731/a_8_216# OR2X1_LOC_731/B 0.39fF
C43966 OR2X1_LOC_738/A OR2X1_LOC_731/B 0.04fF
C56420 OR2X1_LOC_731/B VSS 0.17fF
C17844 OR2X1_LOC_213/A OR2X1_LOC_213/B 0.13fF
C23144 OR2X1_LOC_213/a_8_216# OR2X1_LOC_213/B 0.39fF
C48898 VDD OR2X1_LOC_213/B -0.00fF
C56680 OR2X1_LOC_213/B VSS 0.17fF
C560 OR2X1_LOC_486/Y OR2X1_LOC_563/A 0.01fF
C22778 OR2X1_LOC_736/Y OR2X1_LOC_563/A 0.07fF
C41655 OR2X1_LOC_563/A OR2X1_LOC_366/Y 0.07fF
C42136 OR2X1_LOC_563/A OR2X1_LOC_556/a_8_216# 0.01fF
C44377 OR2X1_LOC_858/A OR2X1_LOC_563/A 0.07fF
C48793 OR2X1_LOC_811/A OR2X1_LOC_563/A 0.07fF
C52510 OR2X1_LOC_563/A OR2X1_LOC_580/B 0.07fF
C53327 OR2X1_LOC_563/A OR2X1_LOC_562/A 0.02fF
C56488 OR2X1_LOC_563/A VSS -1.40fF
C5189 OR2X1_LOC_205/Y OR2X1_LOC_124/Y 0.01fF
C6543 OR2X1_LOC_124/Y OR2X1_LOC_217/A 0.16fF
C8818 OR2X1_LOC_124/Y OR2X1_LOC_572/a_8_216# 0.07fF
C14516 OR2X1_LOC_124/Y OR2X1_LOC_217/a_8_216# 0.05fF
C30656 OR2X1_LOC_244/A OR2X1_LOC_124/Y 0.01fF
C51131 OR2X1_LOC_205/a_8_216# OR2X1_LOC_124/Y 0.39fF
C53902 OR2X1_LOC_124/Y OR2X1_LOC_267/Y 0.14fF
C56857 OR2X1_LOC_124/Y VSS 0.44fF
C939 OR2X1_LOC_486/Y OR2X1_LOC_365/a_36_216# 0.02fF
C2854 OR2X1_LOC_212/a_36_216# OR2X1_LOC_486/Y 0.02fF
C6411 OR2X1_LOC_486/Y OR2X1_LOC_367/B 0.39fF
C19254 OR2X1_LOC_486/Y OR2X1_LOC_182/a_8_216# 0.03fF
C26403 OR2X1_LOC_486/Y OR2X1_LOC_578/B 9.76fF
C26962 VDD OR2X1_LOC_486/Y 0.56fF
C30257 OR2X1_LOC_486/Y OR2X1_LOC_212/B 0.05fF
C37071 OR2X1_LOC_741/Y OR2X1_LOC_486/Y 0.03fF
C43456 OR2X1_LOC_486/Y OR2X1_LOC_556/a_8_216# 0.01fF
C51593 OR2X1_LOC_486/Y OR2X1_LOC_365/a_8_216# 0.02fF
C51946 OR2X1_LOC_223/A OR2X1_LOC_486/Y 0.03fF
C53479 OR2X1_LOC_212/a_8_216# OR2X1_LOC_486/Y 0.03fF
C53824 OR2X1_LOC_486/Y OR2X1_LOC_580/B 0.18fF
C54612 OR2X1_LOC_486/Y OR2X1_LOC_562/A 0.01fF
C56668 OR2X1_LOC_486/Y VSS 0.17fF
C11735 OR2X1_LOC_347/Y OR2X1_LOC_244/Y 0.06fF
C17252 OR2X1_LOC_347/Y OR2X1_LOC_360/a_8_216# 0.39fF
C56589 OR2X1_LOC_347/Y VSS 0.18fF
C89 OR2X1_LOC_244/B OR2X1_LOC_560/A 0.02fF
C1869 OR2X1_LOC_217/Y OR2X1_LOC_560/A 0.46fF
C2334 OR2X1_LOC_217/a_8_216# OR2X1_LOC_560/A 0.01fF
C9571 OR2X1_LOC_864/A OR2X1_LOC_560/A 0.14fF
C28979 OR2X1_LOC_244/Y OR2X1_LOC_560/A 0.02fF
C41629 OR2X1_LOC_267/Y OR2X1_LOC_560/A 0.09fF
C45616 OR2X1_LOC_663/A OR2X1_LOC_560/A 0.03fF
C46494 VDD OR2X1_LOC_560/A 0.41fF
C49273 OR2X1_LOC_205/Y OR2X1_LOC_560/A 0.04fF
C56260 OR2X1_LOC_560/A VSS -0.12fF
C14396 OR2X1_LOC_213/A OR2X1_LOC_803/A 0.73fF
C21198 VDD OR2X1_LOC_213/A 0.08fF
C57208 OR2X1_LOC_213/A VSS 0.04fF
C19096 OR2X1_LOC_477/Y OR2X1_LOC_470/A 0.01fF
C21326 OR2X1_LOC_470/a_8_216# OR2X1_LOC_470/A 0.39fF
C44252 OR2X1_LOC_470/B OR2X1_LOC_470/A 0.08fF
C46262 VDD OR2X1_LOC_470/A -0.00fF
C57271 OR2X1_LOC_470/A VSS 0.18fF
C1066 OR2X1_LOC_244/B OR2X1_LOC_267/Y 0.47fF
C5723 VDD OR2X1_LOC_244/B 0.12fF
C33981 OR2X1_LOC_244/B OR2X1_LOC_244/A 0.29fF
C44443 OR2X1_LOC_244/B OR2X1_LOC_244/Y 0.01fF
C52221 OR2X1_LOC_244/B OR2X1_LOC_244/a_8_216# 0.02fF
C57261 OR2X1_LOC_244/B VSS 0.22fF
C7435 AND2X1_LOC_544/Y AND2X1_LOC_551/B 0.10fF
C18498 AND2X1_LOC_551/a_8_24# AND2X1_LOC_551/B 0.19fF
C37123 VDD AND2X1_LOC_551/B 0.23fF
C57804 AND2X1_LOC_551/B VSS 0.07fF
C3096 AND2X1_LOC_663/B AND2X1_LOC_361/A 0.10fF
C6959 AND2X1_LOC_361/A AND2X1_LOC_657/A 0.02fF
C7128 VDD AND2X1_LOC_361/A 0.01fF
C10497 AND2X1_LOC_572/a_36_24# AND2X1_LOC_361/A 0.01fF
C33110 AND2X1_LOC_560/B AND2X1_LOC_361/A 0.01fF
C47148 AND2X1_LOC_340/Y AND2X1_LOC_361/A 0.25fF
C51014 AND2X1_LOC_217/Y AND2X1_LOC_361/A 0.02fF
C55575 AND2X1_LOC_572/a_8_24# AND2X1_LOC_361/A 0.03fF
C56507 AND2X1_LOC_361/A VSS 0.68fF
C3391 VDD AND2X1_LOC_641/Y 0.21fF
C21827 AND2X1_LOC_641/Y AND2X1_LOC_650/a_8_24# 0.04fF
C32557 AND2X1_LOC_341/a_8_24# AND2X1_LOC_641/Y 0.20fF
C32763 AND2X1_LOC_641/Y AND2X1_LOC_650/a_36_24# 0.01fF
C40317 AND2X1_LOC_641/Y AND2X1_LOC_650/Y 0.04fF
C57160 AND2X1_LOC_641/Y VSS 0.18fF
C4527 AND2X1_LOC_719/Y AND2X1_LOC_576/Y 0.10fF
C10110 AND2X1_LOC_719/Y AND2X1_LOC_580/A 0.03fF
C11282 AND2X1_LOC_719/Y AND2X1_LOC_663/A 0.52fF
C13932 AND2X1_LOC_719/Y AND2X1_LOC_862/A 0.25fF
C14821 AND2X1_LOC_719/Y AND2X1_LOC_578/A 0.10fF
C16358 AND2X1_LOC_719/Y AND2X1_LOC_723/Y 0.15fF
C20441 AND2X1_LOC_719/Y AND2X1_LOC_851/B 0.10fF
C31462 AND2X1_LOC_719/Y AND2X1_LOC_222/Y 0.03fF
C31988 AND2X1_LOC_719/Y AND2X1_LOC_860/A 0.10fF
C32278 AND2X1_LOC_719/Y AND2X1_LOC_562/Y 0.10fF
C33747 AND2X1_LOC_719/Y AND2X1_LOC_658/A 0.04fF
C34992 AND2X1_LOC_719/Y AND2X1_LOC_476/Y 0.10fF
C37789 AND2X1_LOC_719/Y AND2X1_LOC_563/Y 0.03fF
C38367 AND2X1_LOC_719/Y AND2X1_LOC_861/B 0.03fF
C39754 AND2X1_LOC_719/Y AND2X1_LOC_859/Y 0.06fF
C40030 AND2X1_LOC_719/Y AND2X1_LOC_722/a_8_24# 0.25fF
C40345 AND2X1_LOC_719/Y AND2X1_LOC_657/A 0.10fF
C40493 AND2X1_LOC_719/Y VDD 1.87fF
C45375 AND2X1_LOC_719/Y AND2X1_LOC_862/a_8_24# 0.20fF
C48886 AND2X1_LOC_719/Y AND2X1_LOC_806/A 0.01fF
C58011 AND2X1_LOC_719/Y VSS 1.03fF
C13006 VDD AND2X1_LOC_194/Y 0.01fF
C56556 AND2X1_LOC_194/Y VSS -0.02fF
C17908 AND2X1_LOC_182/A AND2X1_LOC_222/Y 0.01fF
C21920 AND2X1_LOC_182/A AND2X1_LOC_182/a_8_24# 0.10fF
C49424 AND2X1_LOC_182/A AND2X1_LOC_866/A 0.25fF
C57932 AND2X1_LOC_182/A VSS 0.30fF
C13888 AND2X1_LOC_675/Y AND2X1_LOC_806/a_8_24# 0.11fF
C16371 AND2X1_LOC_675/Y AND2X1_LOC_658/A 0.03fF
C23270 AND2X1_LOC_675/Y VDD 0.73fF
C27859 AND2X1_LOC_675/Y AND2X1_LOC_657/Y 0.18fF
C31357 AND2X1_LOC_675/Y AND2X1_LOC_806/A 0.23fF
C36675 AND2X1_LOC_501/Y AND2X1_LOC_675/Y 0.05fF
C36682 AND2X1_LOC_675/Y AND2X1_LOC_570/Y 0.16fF
C40616 AND2X1_LOC_675/Y AND2X1_LOC_807/Y 0.22fF
C42035 AND2X1_LOC_675/Y AND2X1_LOC_657/a_8_24# 0.18fF
C43253 AND2X1_LOC_675/Y AND2X1_LOC_576/Y 0.03fF
C48923 AND2X1_LOC_675/Y AND2X1_LOC_580/A 0.03fF
C50111 AND2X1_LOC_675/Y AND2X1_LOC_663/A 0.19fF
C53636 AND2X1_LOC_675/Y AND2X1_LOC_578/A 0.12fF
C56036 AND2X1_LOC_675/Y AND2X1_LOC_735/Y 0.61fF
C57881 AND2X1_LOC_675/Y VSS -1.14fF
C1165 AND2X1_LOC_573/a_8_24# AND2X1_LOC_501/Y 0.15fF
C9618 AND2X1_LOC_501/Y VDD 0.01fF
C14287 AND2X1_LOC_501/Y AND2X1_LOC_657/Y 0.04fF
C16733 AND2X1_LOC_573/Y AND2X1_LOC_501/Y 0.01fF
C29629 AND2X1_LOC_501/Y AND2X1_LOC_576/Y 0.03fF
C34161 AND2X1_LOC_501/Y AND2X1_LOC_735/a_8_24# 0.01fF
C42268 AND2X1_LOC_501/Y AND2X1_LOC_735/Y 0.38fF
C57931 AND2X1_LOC_501/Y VSS -0.05fF
C5085 AND2X1_LOC_605/Y AND2X1_LOC_477/A 0.03fF
C7036 VDD AND2X1_LOC_605/Y 0.29fF
C8802 AND2X1_LOC_732/a_8_24# AND2X1_LOC_605/Y 0.01fF
C14321 AND2X1_LOC_738/B AND2X1_LOC_605/Y 0.01fF
C26578 AND2X1_LOC_732/B AND2X1_LOC_605/Y 0.04fF
C29210 AND2X1_LOC_605/Y AND2X1_LOC_454/Y 0.01fF
C47373 AND2X1_LOC_605/Y AND2X1_LOC_645/a_8_24# 0.11fF
C57628 AND2X1_LOC_605/Y VSS 0.19fF
C111 AND2X1_LOC_544/Y AND2X1_LOC_212/Y 0.19fF
C2805 AND2X1_LOC_736/Y AND2X1_LOC_544/Y 1.68fF
C3555 AND2X1_LOC_727/Y AND2X1_LOC_544/Y 0.03fF
C8343 AND2X1_LOC_737/Y AND2X1_LOC_544/Y 0.05fF
C8545 AND2X1_LOC_544/Y AND2X1_LOC_808/A 3.01fF
C13247 AND2X1_LOC_544/Y AND2X1_LOC_222/Y 0.03fF
C16718 AND2X1_LOC_544/Y AND2X1_LOC_476/Y 0.02fF
C22332 AND2X1_LOC_544/Y VDD 0.38fF
C25651 AND2X1_LOC_544/Y AND2X1_LOC_469/a_8_24# 0.03fF
C26937 AND2X1_LOC_544/Y AND2X1_LOC_657/Y 0.03fF
C28593 AND2X1_LOC_544/Y AND2X1_LOC_213/B 0.03fF
C29473 AND2X1_LOC_738/B AND2X1_LOC_544/Y 0.07fF
C39683 AND2X1_LOC_544/Y AND2X1_LOC_807/Y 0.20fF
C47460 AND2X1_LOC_544/Y AND2X1_LOC_477/Y 0.07fF
C47695 AND2X1_LOC_544/Y GATE_811 0.05fF
C49166 AND2X1_LOC_544/Y AND2X1_LOC_663/A 0.41fF
C52100 AND2X1_LOC_803/B AND2X1_LOC_544/Y 0.03fF
C53620 AND2X1_LOC_544/Y AND2X1_LOC_803/a_8_24# 0.07fF
C58035 AND2X1_LOC_544/Y VSS 0.17fF
C2348 VDD AND2X1_LOC_213/B 0.19fF
C6980 AND2X1_LOC_657/Y AND2X1_LOC_213/B 0.03fF
C29062 AND2X1_LOC_663/A AND2X1_LOC_213/B 0.05fF
C45204 AND2X1_LOC_564/A AND2X1_LOC_213/B 0.03fF
C51727 AND2X1_LOC_658/A AND2X1_LOC_213/B 0.03fF
C54367 AND2X1_LOC_797/A AND2X1_LOC_213/B 0.12fF
C55387 AND2X1_LOC_213/B AND2X1_LOC_796/A 0.01fF
C56605 AND2X1_LOC_213/B VSS 0.21fF
C5383 AND2X1_LOC_365/a_8_24# AND2X1_LOC_365/A 0.03fF
C19909 VDD AND2X1_LOC_365/A 0.24fF
C25597 AND2X1_LOC_365/A AND2X1_LOC_863/Y 0.25fF
C34736 AND2X1_LOC_365/A AND2X1_LOC_654/Y 0.08fF
C37144 AND2X1_LOC_212/A AND2X1_LOC_365/A 0.12fF
C40208 AND2X1_LOC_365/A AND2X1_LOC_661/a_8_24# -0.01fF
C56103 AND2X1_LOC_364/Y AND2X1_LOC_365/A 0.04fF
C57601 AND2X1_LOC_365/A VSS 0.20fF
C1685 AND2X1_LOC_644/Y AND2X1_LOC_648/a_8_24# 0.09fF
C56687 AND2X1_LOC_644/Y VSS 0.08fF
C17154 OR2X1_LOC_576/A OR2X1_LOC_474/B 0.15fF
C25721 OR2X1_LOC_860/Y OR2X1_LOC_474/B 0.89fF
C47970 OR2X1_LOC_865/B OR2X1_LOC_474/B 0.04fF
C55948 VDD OR2X1_LOC_474/B 0.06fF
C56654 OR2X1_LOC_474/B VSS 0.29fF
C33549 OR2X1_LOC_569/B OR2X1_LOC_569/A 0.43fF
C56486 OR2X1_LOC_569/A VSS 0.18fF
C15582 VDD OR2X1_LOC_784/Y 0.08fF
C56786 OR2X1_LOC_784/Y VSS -0.05fF
C3786 VDD OR2X1_LOC_563/B 0.21fF
C4465 OR2X1_LOC_563/B OR2X1_LOC_577/B 0.88fF
C8439 OR2X1_LOC_563/B OR2X1_LOC_577/Y 0.02fF
C16975 OR2X1_LOC_563/a_8_216# OR2X1_LOC_563/B 0.06fF
C41803 OR2X1_LOC_563/B D_GATE_366 0.02fF
C56546 OR2X1_LOC_563/B VSS 0.21fF
C6575 OR2X1_LOC_640/Y OR2X1_LOC_650/a_8_216# 0.39fF
C57837 OR2X1_LOC_640/Y VSS 0.17fF
C8704 OR2X1_LOC_267/Y OR2X1_LOC_576/A 0.74fF
C19511 OR2X1_LOC_244/A OR2X1_LOC_267/Y 0.13fF
C29900 OR2X1_LOC_267/Y OR2X1_LOC_244/Y 0.01fF
C32952 OR2X1_LOC_141/B OR2X1_LOC_267/Y 0.67fF
C37511 OR2X1_LOC_244/a_8_216# OR2X1_LOC_267/Y 0.01fF
C40344 OR2X1_LOC_267/Y OR2X1_LOC_141/a_8_216# 0.01fF
C43587 OR2X1_LOC_657/a_8_216# OR2X1_LOC_267/Y 0.01fF
C47487 VDD OR2X1_LOC_267/Y -0.00fF
C51596 OR2X1_LOC_267/Y OR2X1_LOC_217/A 0.01fF
C53791 OR2X1_LOC_267/Y OR2X1_LOC_572/a_8_216# 0.01fF
C54717 OR2X1_LOC_659/B OR2X1_LOC_267/Y 0.09fF
C56709 OR2X1_LOC_267/Y VSS 0.32fF
C1993 AND2X1_LOC_658/A AND2X1_LOC_862/Y 0.21fF
C2840 AND2X1_LOC_570/Y AND2X1_LOC_658/A 0.03fF
C3894 AND2X1_LOC_658/A AND2X1_LOC_796/Y 0.03fF
C7515 AND2X1_LOC_658/A AND2X1_LOC_865/a_8_24# 0.01fF
C9322 AND2X1_LOC_576/Y AND2X1_LOC_658/A 0.07fF
C10501 AND2X1_LOC_737/a_8_24# AND2X1_LOC_658/A 0.04fF
C11532 AND2X1_LOC_658/A AND2X1_LOC_866/A 0.01fF
C13088 AND2X1_LOC_658/A AND2X1_LOC_866/B 0.01fF
C13122 AND2X1_LOC_658/A AND2X1_LOC_858/a_8_24# 0.04fF
C14272 AND2X1_LOC_658/A AND2X1_LOC_477/Y 0.07fF
C14795 AND2X1_LOC_580/A AND2X1_LOC_658/A 11.83fF
C15952 AND2X1_LOC_658/A AND2X1_LOC_663/A 0.03fF
C19526 AND2X1_LOC_578/A AND2X1_LOC_658/A 0.07fF
C21591 AND2X1_LOC_737/a_36_24# AND2X1_LOC_658/A 0.01fF
C21956 AND2X1_LOC_658/A AND2X1_LOC_658/a_8_24# 0.01fF
C23219 AND2X1_LOC_658/A AND2X1_LOC_212/Y 0.07fF
C24181 AND2X1_LOC_658/A AND2X1_LOC_858/a_36_24# 0.01fF
C34639 AND2X1_LOC_658/A AND2X1_LOC_804/Y 0.03fF
C35428 AND2X1_LOC_658/A AND2X1_LOC_858/B 0.08fF
C36125 AND2X1_LOC_658/A AND2X1_LOC_222/Y 0.03fF
C39659 AND2X1_LOC_658/A AND2X1_LOC_476/Y 0.07fF
C41110 AND2X1_LOC_658/A AND2X1_LOC_663/B 0.01fF
C41372 AND2X1_LOC_658/A AND2X1_LOC_807/B 0.10fF
C42916 AND2X1_LOC_658/A AND2X1_LOC_810/Y 0.03fF
C43163 AND2X1_LOC_861/B AND2X1_LOC_658/A 0.31fF
C44535 AND2X1_LOC_658/A AND2X1_LOC_859/Y 0.07fF
C45161 AND2X1_LOC_658/A AND2X1_LOC_657/A 0.07fF
C45291 VDD AND2X1_LOC_658/A 0.32fF
C50093 AND2X1_LOC_658/A AND2X1_LOC_469/B 0.03fF
C50195 AND2X1_LOC_658/A AND2X1_LOC_862/a_8_24# 0.01fF
C52607 AND2X1_LOC_738/B AND2X1_LOC_658/A 0.07fF
C53572 AND2X1_LOC_658/A AND2X1_LOC_806/A 0.03fF
C55128 AND2X1_LOC_658/A AND2X1_LOC_865/A 0.16fF
C57333 AND2X1_LOC_658/A VSS -1.46fF
C1917 AND2X1_LOC_712/Y AND2X1_LOC_713/Y 0.08fF
C4436 AND2X1_LOC_713/Y VDD 0.38fF
C44646 AND2X1_LOC_713/Y AND2X1_LOC_645/a_8_24# 0.19fF
C57873 AND2X1_LOC_713/Y VSS 0.15fF
C130 AND2X1_LOC_785/Y AND2X1_LOC_795/a_8_24# -0.00fF
C20621 VDD AND2X1_LOC_785/Y 0.21fF
C56271 AND2X1_LOC_785/Y VSS 0.16fF
C20925 AND2X1_LOC_170/Y AND2X1_LOC_566/Y 0.83fF
C34837 AND2X1_LOC_170/Y AND2X1_LOC_566/a_8_24# 0.01fF
C40985 AND2X1_LOC_170/Y AND2X1_LOC_212/Y 0.06fF
C57866 AND2X1_LOC_170/Y VSS 0.12fF
C12915 AND2X1_LOC_717/Y AND2X1_LOC_222/Y 0.03fF
C16377 AND2X1_LOC_717/Y AND2X1_LOC_476/Y 0.07fF
C22019 AND2X1_LOC_717/Y VDD 0.09fF
C53571 AND2X1_LOC_717/Y AND2X1_LOC_723/a_8_24# -0.01fF
C53944 AND2X1_LOC_723/Y AND2X1_LOC_717/Y 0.13fF
C57973 AND2X1_LOC_717/Y VSS -0.04fF
C4128 AND2X1_LOC_857/Y AND2X1_LOC_654/B 0.34fF
C19860 VDD AND2X1_LOC_654/B 0.24fF
C57110 AND2X1_LOC_654/B VSS 0.30fF
C7440 AND2X1_LOC_712/Y AND2X1_LOC_725/a_8_24# 0.18fF
C15583 AND2X1_LOC_712/Y AND2X1_LOC_454/Y 0.01fF
C49648 AND2X1_LOC_712/Y VDD 0.21fF
C57874 AND2X1_LOC_712/Y VSS 0.06fF
C2565 AND2X1_LOC_727/Y GATE_811 0.01fF
C4028 AND2X1_LOC_727/Y AND2X1_LOC_663/A 0.45fF
C16737 AND2X1_LOC_727/Y AND2X1_LOC_731/Y 0.26fF
C19544 AND2X1_LOC_727/Y AND2X1_LOC_808/A 0.03fF
C20132 AND2X1_LOC_727/Y AND2X1_LOC_564/A 0.03fF
C30946 AND2X1_LOC_727/Y AND2X1_LOC_810/Y 0.09fF
C33263 AND2X1_LOC_727/Y VDD 0.24fF
C37882 AND2X1_LOC_727/Y AND2X1_LOC_657/Y 0.03fF
C47687 AND2X1_LOC_727/Y AND2X1_LOC_812/a_8_24# 0.20fF
C58086 AND2X1_LOC_727/Y VSS 0.10fF
C4459 AND2X1_LOC_357/B AND2X1_LOC_364/Y 0.01fF
C7865 AND2X1_LOC_357/A AND2X1_LOC_357/B 1.32fF
C24459 VDD AND2X1_LOC_357/B 0.01fF
C30153 AND2X1_LOC_357/B AND2X1_LOC_863/Y 0.01fF
C39295 AND2X1_LOC_357/B AND2X1_LOC_654/Y 0.02fF
C43597 AND2X1_LOC_357/B AND2X1_LOC_357/a_8_24# 0.04fF
C54731 AND2X1_LOC_357/B AND2X1_LOC_357/a_36_24# 0.01fF
C57792 AND2X1_LOC_357/B VSS 0.19fF
C7980 AND2X1_LOC_797/A AND2X1_LOC_213/a_8_24# 0.20fF
C10607 AND2X1_LOC_797/a_8_24# AND2X1_LOC_797/A 0.09fF
C13511 AND2X1_LOC_797/A AND2X1_LOC_220/B 0.45fF
C48134 VDD AND2X1_LOC_797/A 0.21fF
C57166 AND2X1_LOC_797/A VSS 0.26fF
C57382 OR2X1_LOC_466/A VSS 0.21fF
C32859 OR2X1_LOC_857/B VDD 0.05fF
C37019 OR2X1_LOC_857/B OR2X1_LOC_853/a_8_216# 0.04fF
C48341 OR2X1_LOC_857/B OR2X1_LOC_857/A 0.14fF
C57904 OR2X1_LOC_857/B VSS 0.26fF
C9939 OR2X1_LOC_141/B OR2X1_LOC_244/A 0.18fF
C30780 OR2X1_LOC_141/B OR2X1_LOC_141/a_8_216# 0.02fF
C33982 OR2X1_LOC_141/B OR2X1_LOC_657/a_8_216# 0.01fF
C37646 VDD OR2X1_LOC_141/B 0.10fF
C41817 OR2X1_LOC_141/B OR2X1_LOC_217/A 0.01fF
C44049 OR2X1_LOC_141/B OR2X1_LOC_572/a_8_216# 0.01fF
C45099 OR2X1_LOC_141/B OR2X1_LOC_659/B 0.01fF
C55200 OR2X1_LOC_141/B OR2X1_LOC_576/A 0.01fF
C57785 OR2X1_LOC_141/B VSS 0.29fF
C22597 OR2X1_LOC_207/B OR2X1_LOC_200/Y 0.07fF
C43622 OR2X1_LOC_207/B OR2X1_LOC_200/a_8_216# 0.01fF
C58061 OR2X1_LOC_207/B VSS -0.44fF
C23337 OR2X1_LOC_568/A OR2X1_LOC_566/Y 0.10fF
C54198 OR2X1_LOC_468/Y OR2X1_LOC_568/A 0.01fF
C56396 OR2X1_LOC_568/A VSS -0.26fF
C3136 OR2X1_LOC_206/A OR2X1_LOC_206/a_8_216# 0.08fF
C57054 OR2X1_LOC_206/A VSS 0.12fF
C12790 AND2X1_LOC_859/Y AND2X1_LOC_807/Y 0.02fF
C20886 AND2X1_LOC_580/A AND2X1_LOC_859/Y 0.07fF
C22098 AND2X1_LOC_859/Y AND2X1_LOC_663/A 0.10fF
C43062 AND2X1_LOC_859/Y AND2X1_LOC_562/Y 0.10fF
C49380 AND2X1_LOC_861/B AND2X1_LOC_859/Y 0.01fF
C51429 VDD AND2X1_LOC_859/Y 0.71fF
C57288 AND2X1_LOC_859/Y VSS -1.05fF
C23377 VDD OR2X1_LOC_564/A 0.12fF
C33463 OR2X1_LOC_741/Y OR2X1_LOC_564/A 0.02fF
C47792 OR2X1_LOC_564/B OR2X1_LOC_564/A 0.13fF
C49729 OR2X1_LOC_564/A OR2X1_LOC_564/a_8_216# 0.01fF
C56590 OR2X1_LOC_564/A VSS -0.01fF
C10554 OR2X1_LOC_223/A OR2X1_LOC_723/B 0.01fF
C32452 OR2X1_LOC_479/Y OR2X1_LOC_723/B 0.03fF
C41725 VDD OR2X1_LOC_723/B 0.02fF
C56121 OR2X1_LOC_804/A OR2X1_LOC_723/B 0.07fF
C56368 OR2X1_LOC_723/B VSS 0.35fF
C209 OR2X1_LOC_566/A OR2X1_LOC_212/A 0.02fF
C10103 OR2X1_LOC_566/A OR2X1_LOC_479/Y 0.05fF
C16326 OR2X1_LOC_566/A OR2X1_LOC_808/B 0.05fF
C21978 OR2X1_LOC_566/A OR2X1_LOC_468/Y 0.02fF
C39664 OR2X1_LOC_566/A OR2X1_LOC_211/a_8_216# 0.01fF
C58069 OR2X1_LOC_566/A VSS 0.22fF
C15487 AND2X1_LOC_340/Y AND2X1_LOC_219/Y 0.07fF
C24599 AND2X1_LOC_340/Y AND2X1_LOC_350/Y 0.03fF
C30085 AND2X1_LOC_340/Y AND2X1_LOC_351/Y 0.20fF
C35815 AND2X1_LOC_340/Y VDD 0.09fF
C57938 AND2X1_LOC_340/Y VSS -0.29fF
C6465 AND2X1_LOC_715/Y AND2X1_LOC_724/A 0.01fF
C10840 AND2X1_LOC_724/A VDD 0.21fF
C12052 AND2X1_LOC_724/a_8_24# AND2X1_LOC_724/A 0.03fF
C57875 AND2X1_LOC_724/A VSS 0.21fF
C11916 AND2X1_LOC_454/Y AND2X1_LOC_466/a_36_24# 0.01fF
C18172 VDD AND2X1_LOC_454/Y 0.21fF
C51507 AND2X1_LOC_454/Y AND2X1_LOC_466/a_8_24# 0.03fF
C56728 AND2X1_LOC_454/Y VSS 0.11fF
C15043 AND2X1_LOC_338/Y AND2X1_LOC_339/Y 0.14fF
C26073 AND2X1_LOC_338/Y AND2X1_LOC_351/a_8_24# 0.03fF
C57898 AND2X1_LOC_338/Y VSS 0.14fF
C2093 AND2X1_LOC_861/B AND2X1_LOC_806/A 0.01fF
C4150 VDD AND2X1_LOC_806/A 0.31fF
C21740 AND2X1_LOC_807/Y AND2X1_LOC_806/A 0.03fF
C28047 AND2X1_LOC_858/a_8_24# AND2X1_LOC_806/A 0.01fF
C29736 AND2X1_LOC_580/A AND2X1_LOC_806/A 0.03fF
C30944 AND2X1_LOC_663/A AND2X1_LOC_806/A 0.05fF
C33541 AND2X1_LOC_862/A AND2X1_LOC_806/A 0.01fF
C46279 AND2X1_LOC_244/a_8_24# AND2X1_LOC_806/A 0.01fF
C50637 AND2X1_LOC_858/B AND2X1_LOC_806/A 0.38fF
C51863 AND2X1_LOC_860/A AND2X1_LOC_806/A 0.02fF
C52091 AND2X1_LOC_806/A AND2X1_LOC_562/Y 0.01fF
C52745 AND2X1_LOC_860/a_8_24# AND2X1_LOC_806/A 0.01fF
C56552 AND2X1_LOC_806/A VSS -0.43fF
C8794 OR2X1_LOC_244/Y OR2X1_LOC_632/Y 0.06fF
C26164 VDD OR2X1_LOC_632/Y 0.47fF
C44874 OR2X1_LOC_858/A OR2X1_LOC_632/Y 0.23fF
C51417 OR2X1_LOC_571/B OR2X1_LOC_632/Y 0.08fF
C56511 OR2X1_LOC_632/Y VSS 0.48fF
C1444 OR2X1_LOC_858/B OR2X1_LOC_580/A 0.02fF
C6597 OR2X1_LOC_858/B OR2X1_LOC_858/a_8_216# 0.39fF
C7512 OR2X1_LOC_858/B OR2X1_LOC_858/A 0.46fF
C57988 OR2X1_LOC_858/B VSS 0.09fF
C1250 OR2X1_LOC_805/a_8_216# OR2X1_LOC_362/B 0.01fF
C6729 OR2X1_LOC_362/B OR2X1_LOC_806/a_8_216# 0.09fF
C9537 OR2X1_LOC_362/B OR2X1_LOC_580/a_8_216# 0.01fF
C11231 OR2X1_LOC_362/B OR2X1_LOC_580/A 0.01fF
C12306 OR2X1_LOC_807/B OR2X1_LOC_362/B 0.01fF
C21678 OR2X1_LOC_362/B OR2X1_LOC_811/A 0.12fF
C23411 OR2X1_LOC_362/B OR2X1_LOC_807/A 0.25fF
C25344 OR2X1_LOC_362/B OR2X1_LOC_580/B 0.12fF
C26054 OR2X1_LOC_362/B D_GATE_579 0.73fF
C36472 OR2X1_LOC_362/B OR2X1_LOC_807/a_8_216# 0.01fF
C50647 OR2X1_LOC_807/Y OR2X1_LOC_362/B 0.01fF
C50993 OR2X1_LOC_363/B OR2X1_LOC_362/B 0.12fF
C57362 OR2X1_LOC_362/B VSS 0.42fF
C6029 AND2X1_LOC_359/B AND2X1_LOC_866/A 0.08fF
C12264 AND2X1_LOC_363/Y AND2X1_LOC_359/B 0.02fF
C30950 AND2X1_LOC_367/A AND2X1_LOC_359/B 0.19fF
C31321 AND2X1_LOC_359/B AND2X1_LOC_860/A 0.03fF
C39776 VDD AND2X1_LOC_359/B 0.02fF
C57355 AND2X1_LOC_359/B VSS 0.19fF
C21327 AND2X1_LOC_578/A AND2X1_LOC_851/A 0.06fF
C26843 AND2X1_LOC_851/A AND2X1_LOC_851/B 0.09fF
C31704 AND2X1_LOC_851/a_8_24# AND2X1_LOC_851/A 0.19fF
C47139 VDD AND2X1_LOC_851/A 0.25fF
C57285 AND2X1_LOC_851/A VSS 0.10fF
C22843 AND2X1_LOC_207/A AND2X1_LOC_207/B 0.19fF
C37543 AND2X1_LOC_207/a_8_24# AND2X1_LOC_207/A 0.19fF
C45277 VDD AND2X1_LOC_207/A 0.25fF
C57444 AND2X1_LOC_207/A VSS 0.10fF
C14406 AND2X1_LOC_642/Y AND2X1_LOC_649/a_8_24# 0.03fF
C32535 AND2X1_LOC_642/Y AND2X1_LOC_219/Y 0.03fF
C43886 AND2X1_LOC_642/Y AND2X1_LOC_222/Y 0.88fF
C53748 AND2X1_LOC_660/A AND2X1_LOC_642/Y 0.15fF
C56640 AND2X1_LOC_642/Y VSS 0.13fF
C2272 AND2X1_LOC_560/B AND2X1_LOC_660/a_8_24# 0.02fF
C13178 AND2X1_LOC_367/A AND2X1_LOC_560/B 0.10fF
C17917 AND2X1_LOC_560/B AND2X1_LOC_663/B 4.54fF
C22074 VDD AND2X1_LOC_560/B 0.55fF
C22744 AND2X1_LOC_560/B AND2X1_LOC_660/A 0.06fF
C28685 AND2X1_LOC_560/a_8_24# AND2X1_LOC_560/B 0.11fF
C34167 AND2X1_LOC_571/A AND2X1_LOC_560/B 0.01fF
C44302 AND2X1_LOC_560/B AND2X1_LOC_866/A 0.07fF
C52301 AND2X1_LOC_560/B AND2X1_LOC_218/Y 0.18fF
C57624 AND2X1_LOC_560/B VSS 0.18fF
C8765 AND2X1_LOC_471/Y AND2X1_LOC_212/Y 0.01fF
C20721 AND2X1_LOC_471/Y AND2X1_LOC_477/a_8_24# 0.06fF
C21838 AND2X1_LOC_471/Y AND2X1_LOC_222/Y 0.11fF
C25319 AND2X1_LOC_471/Y AND2X1_LOC_476/Y 0.21fF
C28894 AND2X1_LOC_477/A AND2X1_LOC_471/Y 0.16fF
C30819 VDD AND2X1_LOC_471/Y 0.10fF
C35472 AND2X1_LOC_733/Y AND2X1_LOC_471/Y 0.02fF
C55990 AND2X1_LOC_471/Y AND2X1_LOC_477/Y 0.04fF
C56730 AND2X1_LOC_471/Y VSS 0.34fF
C78 AND2X1_LOC_738/B AND2X1_LOC_796/A 0.10fF
C7501 AND2X1_LOC_796/Y AND2X1_LOC_796/A 0.23fF
C34023 AND2X1_LOC_796/a_8_24# AND2X1_LOC_796/A 0.03fF
C46641 AND2X1_LOC_810/Y AND2X1_LOC_796/A 0.11fF
C49078 VDD AND2X1_LOC_796/A 0.75fF
C56309 AND2X1_LOC_796/A VSS 0.65fF
C6048 AND2X1_LOC_578/A AND2X1_LOC_851/B 0.08fF
C16615 AND2X1_LOC_851/a_8_24# AND2X1_LOC_851/B 0.01fF
C22217 AND2X1_LOC_858/B AND2X1_LOC_851/B 0.24fF
C23083 AND2X1_LOC_367/A AND2X1_LOC_851/B 0.10fF
C26336 AND2X1_LOC_851/B AND2X1_LOC_476/Y 0.02fF
C31838 VDD AND2X1_LOC_851/B 0.58fF
C54218 AND2X1_LOC_851/B AND2X1_LOC_866/A 0.07fF
C57236 AND2X1_LOC_851/B VSS 0.21fF
C37749 AND2X1_LOC_810/Y AND2X1_LOC_436/Y 0.02fF
C38135 AND2X1_LOC_477/A AND2X1_LOC_436/Y 0.03fF
C39254 AND2X1_LOC_436/Y AND2X1_LOC_468/a_8_24# 0.10fF
C40053 VDD AND2X1_LOC_436/Y 0.01fF
C56627 AND2X1_LOC_436/Y VSS -0.28fF
C8319 AND2X1_LOC_339/Y VDD 0.01fF
C31561 AND2X1_LOC_339/Y AND2X1_LOC_351/a_8_24# 0.03fF
C42623 AND2X1_LOC_339/Y AND2X1_LOC_351/a_36_24# 0.01fF
C43963 AND2X1_LOC_339/Y AND2X1_LOC_219/Y 0.03fF
C57897 AND2X1_LOC_339/Y VSS 0.23fF
C47905 AND2X1_LOC_715/Y VDD 1.06fF
C57925 AND2X1_LOC_715/Y VSS -5.71fF
C12135 AND2X1_LOC_739/B AND2X1_LOC_739/a_8_24# 0.01fF
C17156 AND2X1_LOC_739/B VDD 0.13fF
C17625 AND2X1_LOC_739/B AND2X1_LOC_740/B 0.05fF
C46982 AND2X1_LOC_739/B AND2X1_LOC_803/B 0.35fF
C58131 AND2X1_LOC_739/B VSS 0.19fF
C14090 AND2X1_LOC_364/Y AND2X1_LOC_863/A 0.16fF
C18322 AND2X1_LOC_857/Y AND2X1_LOC_863/A 0.06fF
C33939 VDD AND2X1_LOC_863/A 0.38fF
C49035 AND2X1_LOC_654/Y AND2X1_LOC_863/A 0.02fF
C57029 AND2X1_LOC_863/A VSS 0.05fF
C10337 OR2X1_LOC_216/Y OR2X1_LOC_218/Y 0.03fF
C13141 VDD OR2X1_LOC_216/Y 0.34fF
C15833 OR2X1_LOC_216/Y OR2X1_LOC_205/Y 0.07fF
C46865 OR2X1_LOC_216/Y OR2X1_LOC_218/a_8_216# 0.05fF
C56798 OR2X1_LOC_216/Y VSS -0.13fF
C4132 OR2X1_LOC_656/Y OR2X1_LOC_660/a_8_216# 0.18fF
C44113 OR2X1_LOC_656/Y OR2X1_LOC_660/B 0.17fF
C48009 OR2X1_LOC_656/Y VDD 0.27fF
C57889 OR2X1_LOC_656/Y VSS -0.61fF
C1647 AND2X1_LOC_366/A AND2X1_LOC_367/a_8_24# 0.01fF
C7154 AND2X1_LOC_366/A GATE_366 0.01fF
C20689 AND2X1_LOC_366/A AND2X1_LOC_363/Y 0.19fF
C26173 AND2X1_LOC_366/A AND2X1_LOC_366/a_8_24# 0.01fF
C31668 AND2X1_LOC_366/A AND2X1_LOC_367/B 0.23fF
C39306 AND2X1_LOC_366/A AND2X1_LOC_367/A 0.49fF
C39692 AND2X1_LOC_366/A AND2X1_LOC_860/A 0.07fF
C48433 AND2X1_LOC_366/A VDD 0.11fF
C57901 AND2X1_LOC_366/A VSS 0.19fF
C1758 AND2X1_LOC_795/Y AND2X1_LOC_476/Y 0.12fF
C7975 AND2X1_LOC_807/Y AND2X1_LOC_476/Y 0.02fF
C12781 AND2X1_LOC_866/A AND2X1_LOC_476/Y 0.07fF
C17228 AND2X1_LOC_663/A AND2X1_LOC_476/Y 0.10fF
C20777 AND2X1_LOC_578/A AND2X1_LOC_476/Y 0.07fF
C22008 AND2X1_LOC_662/B AND2X1_LOC_476/Y 0.08fF
C27023 AND2X1_LOC_736/Y AND2X1_LOC_476/Y 0.07fF
C33255 AND2X1_LOC_564/A AND2X1_LOC_476/Y 0.07fF
C37537 AND2X1_LOC_367/A AND2X1_LOC_476/Y 0.09fF
C46584 AND2X1_LOC_476/Y AND2X1_LOC_479/a_8_24# 0.03fF
C46600 VDD AND2X1_LOC_476/Y 0.47fF
C51311 AND2X1_LOC_657/Y AND2X1_LOC_476/Y 0.10fF
C56628 AND2X1_LOC_476/Y VSS -1.73fF
C7851 AND2X1_LOC_810/Y AND2X1_LOC_812/a_8_24# 0.03fF
C8327 AND2X1_LOC_810/Y AND2X1_LOC_796/Y 0.01fF
C20473 AND2X1_LOC_810/Y AND2X1_LOC_663/A 0.03fF
C34805 AND2X1_LOC_796/a_8_24# AND2X1_LOC_810/Y 0.07fF
C47900 AND2X1_LOC_477/A AND2X1_LOC_810/Y 0.07fF
C49029 AND2X1_LOC_810/Y AND2X1_LOC_468/a_8_24# 0.04fF
C54495 AND2X1_LOC_810/Y AND2X1_LOC_469/B 0.01fF
C57028 AND2X1_LOC_810/Y VSS 0.32fF
C14524 OR2X1_LOC_244/A OR2X1_LOC_244/a_8_216# 0.06fF
C17286 OR2X1_LOC_244/A OR2X1_LOC_141/a_8_216# 0.03fF
C20543 OR2X1_LOC_657/a_8_216# OR2X1_LOC_244/A 0.03fF
C23482 OR2X1_LOC_663/A OR2X1_LOC_244/A 0.07fF
C24281 VDD OR2X1_LOC_244/A 0.99fF
C26015 OR2X1_LOC_657/a_36_216# OR2X1_LOC_244/A 0.01fF
C28345 OR2X1_LOC_244/A OR2X1_LOC_217/A 0.01fF
C30498 OR2X1_LOC_244/A OR2X1_LOC_572/a_8_216# 0.03fF
C31513 OR2X1_LOC_659/B OR2X1_LOC_244/A 0.01fF
C35985 OR2X1_LOC_244/A OR2X1_LOC_572/a_36_216# 0.01fF
C41531 OR2X1_LOC_244/A OR2X1_LOC_576/A 0.02fF
C43416 OR2X1_LOC_864/A OR2X1_LOC_244/A 0.07fF
C57205 OR2X1_LOC_244/A VSS -1.70fF
C3918 OR2X1_LOC_351/B OR2X1_LOC_351/a_36_216# 0.02fF
C7118 OR2X1_LOC_351/B OR2X1_LOC_219/B 0.10fF
C9468 OR2X1_LOC_351/B OR2X1_LOC_358/A 0.08fF
C35008 OR2X1_LOC_351/B VDD 0.18fF
C54351 OR2X1_LOC_351/B OR2X1_LOC_864/A 0.79fF
C54512 OR2X1_LOC_351/B OR2X1_LOC_351/a_8_216# 0.03fF
C57995 OR2X1_LOC_351/B VSS 0.33fF
C4689 AND2X1_LOC_731/Y GATE_811 0.02fF
C7214 AND2X1_LOC_742/a_8_24# GATE_811 0.05fF
C7457 GATE_811 AND2X1_LOC_808/A 0.09fF
C8074 AND2X1_LOC_564/A GATE_811 0.03fF
C12782 GATE_741 GATE_811 0.28fF
C16276 AND2X1_LOC_739/a_8_24# GATE_811 0.01fF
C17694 GATE_811 AND2X1_LOC_738/Y 0.01fF
C25952 GATE_811 AND2X1_LOC_657/Y 0.39fF
C28745 GATE_811 AND2X1_LOC_740/a_8_24# 0.01fF
C34225 GATE_811 AND2X1_LOC_742/A 0.29fF
C35837 GATE_811 AND2X1_LOC_796/Y 0.09fF
C42861 GATE_811 AND2X1_LOC_220/B 0.03fF
C57026 GATE_811 VSS 0.19fF
C7905 AND2X1_LOC_363/Y AND2X1_LOC_367/B 0.21fF
C26589 AND2X1_LOC_367/A AND2X1_LOC_367/B 0.29fF
C35406 VDD AND2X1_LOC_367/B 0.05fF
C44958 AND2X1_LOC_367/B AND2X1_LOC_367/a_8_24# 0.05fF
C50614 AND2X1_LOC_367/B GATE_366 0.83fF
C57668 AND2X1_LOC_367/B VSS 0.02fF
C675 OR2X1_LOC_660/Y OR2X1_LOC_662/a_8_216# 0.01fF
C22902 OR2X1_LOC_660/Y OR2X1_LOC_663/A 0.74fF
C23674 VDD OR2X1_LOC_660/Y -0.00fF
C41035 OR2X1_LOC_662/A OR2X1_LOC_660/Y 0.01fF
C57772 OR2X1_LOC_660/Y VSS 0.10fF
C15433 OR2X1_LOC_218/Y OR2X1_LOC_215/A 0.24fF
C49451 VDD OR2X1_LOC_218/Y 0.20fF
C51625 OR2X1_LOC_218/Y OR2X1_LOC_222/A 0.04fF
C52112 OR2X1_LOC_218/Y OR2X1_LOC_222/a_8_216# 0.06fF
C52139 OR2X1_LOC_218/Y OR2X1_LOC_205/Y 0.03fF
C57141 OR2X1_LOC_218/Y VSS 0.59fF
C1739 VDD AND2X1_LOC_863/Y 0.21fF
C2871 AND2X1_LOC_863/Y AND2X1_LOC_212/a_8_24# 0.04fF
C16643 AND2X1_LOC_863/Y AND2X1_LOC_654/Y 0.04fF
C18473 AND2X1_LOC_863/Y AND2X1_LOC_864/a_8_24# 0.04fF
C19136 AND2X1_LOC_212/A AND2X1_LOC_863/Y 0.13fF
C22239 AND2X1_LOC_863/Y AND2X1_LOC_661/a_8_24# -0.01fF
C24037 AND2X1_LOC_863/Y AND2X1_LOC_866/A 0.03fF
C28589 AND2X1_LOC_863/Y AND2X1_LOC_212/B 0.02fF
C35598 AND2X1_LOC_863/Y AND2X1_LOC_212/Y 0.13fF
C35623 AND2X1_LOC_352/a_8_24# AND2X1_LOC_863/Y 0.02fF
C37757 AND2X1_LOC_364/Y AND2X1_LOC_863/Y 0.38fF
C41140 AND2X1_LOC_357/A AND2X1_LOC_863/Y 0.01fF
C43365 AND2X1_LOC_365/a_8_24# AND2X1_LOC_863/Y 0.01fF
C47797 AND2X1_LOC_863/a_8_24# AND2X1_LOC_863/Y 0.01fF
C49036 AND2X1_LOC_367/A AND2X1_LOC_863/Y 0.01fF
C57175 AND2X1_LOC_863/Y VSS 0.15fF
C7244 AND2X1_LOC_808/A AND2X1_LOC_477/Y 0.01fF
C7824 AND2X1_LOC_564/A AND2X1_LOC_477/Y 0.07fF
C9995 AND2X1_LOC_477/Y AND2X1_LOC_220/a_8_24# 0.01fF
C10489 AND2X1_LOC_477/Y AND2X1_LOC_804/Y 0.01fF
C10879 AND2X1_LOC_477/a_8_24# AND2X1_LOC_477/Y 0.02fF
C15971 AND2X1_LOC_477/Y AND2X1_LOC_808/a_8_24# 0.01fF
C19124 AND2X1_LOC_477/A AND2X1_LOC_477/Y 0.23fF
C20599 AND2X1_LOC_477/Y AND2X1_LOC_794/a_8_24# 0.02fF
C21064 VDD AND2X1_LOC_477/Y 0.03fF
C24442 AND2X1_LOC_477/Y AND2X1_LOC_469/a_8_24# 0.03fF
C25715 AND2X1_LOC_657/Y AND2X1_LOC_477/Y 0.10fF
C25723 AND2X1_LOC_477/Y AND2X1_LOC_469/B 0.17fF
C26089 AND2X1_LOC_477/Y AND2X1_LOC_804/A 0.01fF
C40467 AND2X1_LOC_469/Y AND2X1_LOC_477/Y 0.23fF
C42626 AND2X1_LOC_477/Y AND2X1_LOC_220/B 0.01fF
C47958 AND2X1_LOC_663/A AND2X1_LOC_477/Y 0.10fF
C48511 AND2X1_LOC_477/Y AND2X1_LOC_220/Y 0.21fF
C51733 AND2X1_LOC_477/Y AND2X1_LOC_478/a_8_24# 0.03fF
C55060 AND2X1_LOC_477/Y AND2X1_LOC_212/Y 0.93fF
C56677 AND2X1_LOC_477/Y VSS 0.21fF
C27426 AND2X1_LOC_214/A AND2X1_LOC_207/B 0.83fF
C50097 AND2X1_LOC_214/A VDD 0.19fF
C58136 AND2X1_LOC_214/A VSS -0.31fF
C6256 AND2X1_LOC_576/Y AND2X1_LOC_858/B 0.10fF
C16538 AND2X1_LOC_578/A AND2X1_LOC_858/B 0.08fF
C27036 AND2X1_LOC_851/a_8_24# AND2X1_LOC_858/B 0.01fF
C33760 AND2X1_LOC_858/B AND2X1_LOC_860/A 0.01fF
C34043 AND2X1_LOC_858/B AND2X1_LOC_562/Y 0.10fF
C34622 AND2X1_LOC_860/a_8_24# AND2X1_LOC_858/B 0.02fF
C39563 AND2X1_LOC_858/B AND2X1_LOC_563/Y 0.01fF
C40100 AND2X1_LOC_861/B AND2X1_LOC_858/B 0.01fF
C42128 AND2X1_LOC_858/B AND2X1_LOC_657/A 0.10fF
C42260 VDD AND2X1_LOC_858/B 0.95fF
C57286 AND2X1_LOC_858/B VSS 0.38fF
C57550 OR2X1_LOC_862/B VSS 0.20fF
C13568 AND2X1_LOC_351/a_8_24# AND2X1_LOC_351/Y 0.01fF
C25005 AND2X1_LOC_350/B AND2X1_LOC_351/Y 0.01fF
C34928 AND2X1_LOC_350/Y AND2X1_LOC_351/Y 0.91fF
C46361 VDD AND2X1_LOC_351/Y 0.04fF
C46780 AND2X1_LOC_350/a_8_24# AND2X1_LOC_351/Y 0.01fF
C57480 AND2X1_LOC_351/Y VSS 0.26fF
C6135 AND2X1_LOC_724/Y AND2X1_LOC_732/B 0.01fF
C44410 AND2X1_LOC_724/Y AND2X1_LOC_732/a_8_24# 0.09fF
C58043 AND2X1_LOC_724/Y VSS 0.03fF
C19482 AND2X1_LOC_350/B AND2X1_LOC_350/Y 0.01fF
C41069 AND2X1_LOC_350/a_8_24# AND2X1_LOC_350/Y 0.02fF
C57481 AND2X1_LOC_350/Y VSS 0.12fF
C23123 OR2X1_LOC_569/B OR2X1_LOC_569/a_8_216# 0.07fF
C33280 VDD OR2X1_LOC_569/B 0.20fF
C56545 OR2X1_LOC_569/B VSS 0.16fF
C6631 AND2X1_LOC_861/B AND2X1_LOC_862/Y 0.01fF
C8804 VDD AND2X1_LOC_862/Y 0.02fF
C13601 AND2X1_LOC_862/a_8_24# AND2X1_LOC_862/Y 0.01fF
C18570 AND2X1_LOC_865/A AND2X1_LOC_862/Y 0.02fF
C26269 AND2X1_LOC_862/Y AND2X1_LOC_807/Y 0.02fF
C27095 AND2X1_LOC_862/Y AND2X1_LOC_865/a_8_24# 0.01fF
C32561 AND2X1_LOC_862/Y AND2X1_LOC_866/B 0.86fF
C57130 AND2X1_LOC_862/Y VSS 0.08fF
C926 OR2X1_LOC_357/a_36_216# OR2X1_LOC_578/B 0.02fF
C2233 OR2X1_LOC_364/a_8_216# OR2X1_LOC_578/B 0.05fF
C5585 OR2X1_LOC_741/Y OR2X1_LOC_578/B 0.03fF
C8613 OR2X1_LOC_352/a_8_216# OR2X1_LOC_578/B 0.01fF
C11119 OR2X1_LOC_578/a_8_216# OR2X1_LOC_578/B 0.02fF
C20274 OR2X1_LOC_223/A OR2X1_LOC_578/B 0.03fF
C23352 OR2X1_LOC_566/Y OR2X1_LOC_578/B 0.74fF
C25145 OR2X1_LOC_357/B OR2X1_LOC_578/B 0.09fF
C42212 OR2X1_LOC_479/Y OR2X1_LOC_578/B 5.87fF
C48709 OR2X1_LOC_808/B OR2X1_LOC_578/B 0.05fF
C51577 OR2X1_LOC_357/a_8_216# OR2X1_LOC_578/B 0.03fF
C51618 VDD OR2X1_LOC_578/B 0.39fF
C54202 OR2X1_LOC_468/Y OR2X1_LOC_578/B 0.01fF
C54858 OR2X1_LOC_212/B OR2X1_LOC_578/B 0.03fF
C56347 OR2X1_LOC_578/B VSS 0.39fF
C30194 VDD OR2X1_LOC_214/B 0.15fF
C47450 OR2X1_LOC_214/a_8_216# OR2X1_LOC_214/B 0.06fF
C56801 OR2X1_LOC_214/B VSS 0.22fF
C5779 OR2X1_LOC_863/a_8_216# OR2X1_LOC_863/A 0.39fF
C38967 OR2X1_LOC_857/a_8_216# OR2X1_LOC_863/A 0.01fF
C57614 OR2X1_LOC_863/A VSS 0.18fF
C9369 AND2X1_LOC_364/A AND2X1_LOC_655/A 0.10fF
C20723 VDD AND2X1_LOC_364/A 0.03fF
C38830 AND2X1_LOC_358/Y AND2X1_LOC_364/A 0.02fF
C39794 AND2X1_LOC_357/a_8_24# AND2X1_LOC_364/A 0.01fF
C44417 AND2X1_LOC_364/a_8_24# AND2X1_LOC_364/A 0.04fF
C57537 AND2X1_LOC_364/A VSS 0.32fF
C740 AND2X1_LOC_863/a_8_24# AND2X1_LOC_654/Y 0.04fF
C10921 VDD AND2X1_LOC_654/Y 0.80fF
C28310 AND2X1_LOC_212/A AND2X1_LOC_654/Y 0.02fF
C31349 AND2X1_LOC_654/Y AND2X1_LOC_661/a_8_24# 0.11fF
C42411 AND2X1_LOC_654/Y AND2X1_LOC_662/B 0.02fF
C44880 AND2X1_LOC_352/a_8_24# AND2X1_LOC_654/Y 0.04fF
C47178 AND2X1_LOC_364/Y AND2X1_LOC_654/Y 0.04fF
C50543 AND2X1_LOC_357/A AND2X1_LOC_654/Y 0.03fF
C51427 AND2X1_LOC_857/Y AND2X1_LOC_654/Y 0.18fF
C55716 AND2X1_LOC_654/Y AND2X1_LOC_655/A 0.10fF
C57154 AND2X1_LOC_654/Y VSS -1.24fF
C15504 AND2X1_LOC_732/B VDD 0.41fF
C57872 AND2X1_LOC_732/B VSS -0.02fF
C1959 AND2X1_LOC_865/A AND2X1_LOC_807/B 0.24fF
C3327 AND2X1_LOC_865/A AND2X1_LOC_805/Y 0.08fF
C3709 AND2X1_LOC_861/B AND2X1_LOC_865/A 0.01fF
C10062 AND2X1_LOC_861/a_8_24# AND2X1_LOC_865/A 0.01fF
C23342 AND2X1_LOC_865/A AND2X1_LOC_807/Y 1.19fF
C24141 AND2X1_LOC_865/A AND2X1_LOC_865/a_8_24# 0.04fF
C35065 AND2X1_LOC_865/A AND2X1_LOC_865/a_36_24# 0.01fF
C57332 AND2X1_LOC_865/A VSS -0.05fF
C33482 OR2X1_LOC_577/a_8_216# OR2X1_LOC_577/B 0.05fF
C34839 OR2X1_LOC_577/B D_GATE_366 0.03fF
C52948 VDD OR2X1_LOC_577/B 0.10fF
C56306 OR2X1_LOC_577/B VSS 0.16fF
C13997 OR2X1_LOC_860/Y OR2X1_LOC_865/B 0.14fF
C22016 OR2X1_LOC_860/Y VDD -0.00fF
C57987 OR2X1_LOC_860/Y VSS -0.10fF
C20772 AND2X1_LOC_364/Y AND2X1_LOC_655/A 0.48fF
C25025 AND2X1_LOC_857/Y AND2X1_LOC_655/A 0.05fF
C30245 AND2X1_LOC_649/Y AND2X1_LOC_655/A 0.27fF
C35728 AND2X1_LOC_655/a_8_24# AND2X1_LOC_655/A 0.27fF
C40590 VDD AND2X1_LOC_655/A 1.21fF
C56685 AND2X1_LOC_655/A VSS -3.03fF
C4450 AND2X1_LOC_212/A AND2X1_LOC_367/A 0.42fF
C9461 AND2X1_LOC_367/A AND2X1_LOC_866/A 0.10fF
C15552 AND2X1_LOC_367/A AND2X1_LOC_363/Y 0.11fF
C34047 AND2X1_LOC_367/A AND2X1_LOC_222/Y 0.03fF
C34588 AND2X1_LOC_367/A AND2X1_LOC_860/A 0.07fF
C38981 AND2X1_LOC_367/A AND2X1_LOC_359/a_8_24# 0.01fF
C43016 AND2X1_LOC_367/A AND2X1_LOC_657/A 0.10fF
C43154 VDD AND2X1_LOC_367/A 3.16fF
C44332 AND2X1_LOC_367/A AND2X1_LOC_212/a_8_24# 0.20fF
C44573 AND2X1_LOC_367/A AND2X1_LOC_363/A 0.14fF
C54800 AND2X1_LOC_572/Y AND2X1_LOC_367/A 0.09fF
C57722 AND2X1_LOC_367/A VSS 0.43fF
C23266 AND2X1_LOC_573/Y AND2X1_LOC_576/Y 0.02fF
C35804 AND2X1_LOC_573/Y AND2X1_LOC_735/Y 0.91fF
C57959 AND2X1_LOC_573/Y VSS 0.08fF
C6203 AND2X1_LOC_807/B AND2X1_LOC_807/a_8_24# 0.01fF
C9709 AND2X1_LOC_807/Y AND2X1_LOC_807/B 0.13fF
C10490 AND2X1_LOC_865/a_8_24# AND2X1_LOC_807/B 0.09fF
C45783 AND2X1_LOC_807/B AND2X1_LOC_805/Y 0.03fF
C46198 AND2X1_LOC_861/B AND2X1_LOC_807/B 0.52fF
C48397 VDD AND2X1_LOC_807/B 0.03fF
C52602 AND2X1_LOC_861/a_8_24# AND2X1_LOC_807/B 0.03fF
C56763 AND2X1_LOC_807/B VSS -0.17fF
C2096 AND2X1_LOC_736/Y AND2X1_LOC_580/A 0.29fF
C6776 AND2X1_LOC_736/Y AND2X1_LOC_578/A 0.07fF
C14772 AND2X1_LOC_736/Y AND2X1_LOC_736/a_8_24# 0.01fF
C18634 AND2X1_LOC_736/Y AND2X1_LOC_737/Y 0.05fF
C23550 AND2X1_LOC_736/Y AND2X1_LOC_222/Y 0.03fF
C32494 AND2X1_LOC_736/Y VDD 0.11fF
C58135 AND2X1_LOC_736/Y VSS -0.41fF
C43516 AND2X1_LOC_810/A VDD 0.50fF
C58122 AND2X1_LOC_810/A VSS -0.56fF
C2315 AND2X1_LOC_564/A AND2X1_LOC_469/Y 0.03fF
C4352 AND2X1_LOC_564/A AND2X1_LOC_220/B 0.03fF
C12519 AND2X1_LOC_803/B AND2X1_LOC_564/A 0.03fF
C22339 AND2X1_LOC_564/A AND2X1_LOC_731/Y 0.03fF
C27761 AND2X1_LOC_564/A AND2X1_LOC_220/a_8_24# 0.07fF
C29741 AND2X1_LOC_564/A AND2X1_LOC_222/Y 0.03fF
C29983 AND2X1_LOC_564/A AND2X1_LOC_564/a_8_24# 0.05fF
C30366 AND2X1_LOC_741/a_8_24# AND2X1_LOC_564/A 0.07fF
C38764 AND2X1_LOC_564/A VDD 0.56fF
C38777 AND2X1_LOC_564/A AND2X1_LOC_738/a_8_24# 0.03fF
C46117 AND2X1_LOC_738/B AND2X1_LOC_564/A 0.12fF
C58034 AND2X1_LOC_564/A VSS -0.59fF
C18156 OR2X1_LOC_860/a_8_216# OR2X1_LOC_244/Y 0.02fF
C22864 OR2X1_LOC_244/Y OR2X1_LOC_360/a_8_216# 0.08fF
C23732 OR2X1_LOC_860/a_36_216# OR2X1_LOC_244/Y 0.03fF
C26643 OR2X1_LOC_865/B OR2X1_LOC_244/Y 0.02fF
C26664 OR2X1_LOC_244/Y OR2X1_LOC_573/Y 0.01fF
C32121 OR2X1_LOC_244/Y OR2X1_LOC_575/a_8_216# 0.01fF
C34567 VDD OR2X1_LOC_244/Y 0.38fF
C38394 OR2X1_LOC_658/a_8_216# OR2X1_LOC_244/Y 0.01fF
C41845 OR2X1_LOC_573/a_8_216# OR2X1_LOC_244/Y 0.01fF
C49697 OR2X1_LOC_659/A OR2X1_LOC_244/Y 0.36fF
C52119 OR2X1_LOC_576/A OR2X1_LOC_244/Y 0.05fF
C53473 OR2X1_LOC_858/A OR2X1_LOC_244/Y 0.03fF
C56588 OR2X1_LOC_244/Y VSS 0.47fF
C6906 OR2X1_LOC_477/B OR2X1_LOC_477/a_8_216# 0.02fF
C11023 OR2X1_LOC_477/B OR2X1_LOC_477/Y 0.72fF
C38045 VDD OR2X1_LOC_477/B 0.05fF
C57766 OR2X1_LOC_477/B VSS 0.11fF
C7799 OR2X1_LOC_363/A OR2X1_LOC_580/A 0.04fF
C34108 OR2X1_LOC_363/A OR2X1_LOC_363/a_8_216# 0.19fF
C47563 OR2X1_LOC_363/B OR2X1_LOC_363/A 0.18fF
C51345 VDD OR2X1_LOC_363/A 0.19fF
C56587 OR2X1_LOC_363/A VSS 0.19fF
C3647 OR2X1_LOC_244/a_8_216# OR2X1_LOC_576/A 0.01fF
C5277 OR2X1_LOC_865/B OR2X1_LOC_576/A 0.02fF
C6415 OR2X1_LOC_576/A OR2X1_LOC_141/a_8_216# 0.01fF
C9667 OR2X1_LOC_657/a_8_216# OR2X1_LOC_576/A 0.01fF
C13413 VDD OR2X1_LOC_576/A 0.19fF
C17513 OR2X1_LOC_576/A OR2X1_LOC_217/A 0.01fF
C19725 OR2X1_LOC_572/a_8_216# OR2X1_LOC_576/A 0.01fF
C20708 OR2X1_LOC_659/B OR2X1_LOC_576/A 0.02fF
C28251 OR2X1_LOC_659/A OR2X1_LOC_576/A 0.50fF
C33635 OR2X1_LOC_576/A OR2X1_LOC_571/Y 0.15fF
C39112 OR2X1_LOC_576/A OR2X1_LOC_576/a_8_216# 0.16fF
C53038 OR2X1_LOC_860/a_8_216# OR2X1_LOC_576/A 0.01fF
C56708 OR2X1_LOC_576/A VSS 0.35fF
C7561 VDD OR2X1_LOC_217/Y 0.06fF
C10357 OR2X1_LOC_217/Y OR2X1_LOC_205/Y 0.03fF
C19616 OR2X1_LOC_217/Y OR2X1_LOC_217/a_8_216# 0.01fF
C56799 OR2X1_LOC_217/Y VSS 0.20fF
C11162 OR2X1_LOC_562/Y OR2X1_LOC_570/A 0.06fF
C20258 VDD OR2X1_LOC_570/A -0.00fF
C41492 OR2X1_LOC_570/a_8_216# OR2X1_LOC_570/A 0.39fF
C56594 OR2X1_LOC_570/A VSS 0.18fF
C7479 OR2X1_LOC_220/A OR2X1_LOC_740/B 0.03fF
C11607 OR2X1_LOC_220/A OR2X1_LOC_739/Y 0.02fF
C17276 VDD OR2X1_LOC_220/A 0.26fF
C28163 OR2X1_LOC_220/A OR2X1_LOC_740/a_8_216# 0.06fF
C36804 OR2X1_LOC_220/A OR2X1_LOC_738/A 0.42fF
C53980 OR2X1_LOC_220/A OR2X1_LOC_738/B 0.12fF
C57058 OR2X1_LOC_220/A VSS -0.06fF
C1311 AND2X1_LOC_738/B AND2X1_LOC_477/A 1.00fF
C18856 AND2X1_LOC_568/a_8_24# AND2X1_LOC_477/A 0.01fF
C24379 AND2X1_LOC_578/A AND2X1_LOC_477/A 0.01fF
C28001 AND2X1_LOC_477/A AND2X1_LOC_212/Y 0.01fF
C39896 AND2X1_LOC_477/A AND2X1_LOC_477/a_8_24# 0.01fF
C50275 VDD AND2X1_LOC_477/A 0.14fF
C57102 AND2X1_LOC_477/A VSS 0.23fF
C7562 AND2X1_LOC_364/Y AND2X1_LOC_662/B 0.01fF
C17881 AND2X1_LOC_662/B AND2X1_LOC_662/a_8_24# 0.08fF
C18432 AND2X1_LOC_662/B AND2X1_LOC_222/Y 0.03fF
C27476 VDD AND2X1_LOC_662/B 0.21fF
C44881 AND2X1_LOC_212/A AND2X1_LOC_662/B 0.01fF
C57153 AND2X1_LOC_662/B VSS 0.23fF
C8839 AND2X1_LOC_737/Y AND2X1_LOC_663/A 0.30fF
C10613 AND2X1_LOC_737/Y AND2X1_LOC_811/a_8_24# 0.19fF
C28993 AND2X1_LOC_737/Y AND2X1_LOC_222/Y 0.48fF
C37982 AND2X1_LOC_737/Y VDD 0.34fF
C41213 AND2X1_LOC_737/Y AND2X1_LOC_811/Y 0.01fF
C42752 AND2X1_LOC_737/Y AND2X1_LOC_657/Y 0.03fF
C55704 AND2X1_LOC_737/Y AND2X1_LOC_807/Y 0.33fF
C58134 AND2X1_LOC_737/Y VSS 0.05fF
C23267 AND2X1_LOC_479/Y AND2X1_LOC_222/Y 0.02fF
C29057 AND2X1_LOC_479/Y AND2X1_LOC_480/a_8_24# 0.11fF
C32217 AND2X1_LOC_479/Y AND2X1_LOC_479/a_8_24# 0.02fF
C32234 VDD AND2X1_LOC_479/Y 0.09fF
C57148 AND2X1_LOC_479/Y VSS 0.15fF
C14403 AND2X1_LOC_480/A AND2X1_LOC_223/A 0.10fF
C25266 AND2X1_LOC_223/A AND2X1_LOC_222/Y 0.01fF
C30724 AND2X1_LOC_223/A AND2X1_LOC_223/a_8_24# 0.01fF
C36214 AND2X1_LOC_223/A GATE_222 0.27fF
C36584 GATE_479 AND2X1_LOC_223/A 0.10fF
C56607 AND2X1_LOC_223/A VSS 0.21fF
C4048 AND2X1_LOC_740/B AND2X1_LOC_740/a_8_24# 0.05fF
C9588 AND2X1_LOC_740/B AND2X1_LOC_742/A 0.01fF
C18118 AND2X1_LOC_740/B AND2X1_LOC_220/B 0.03fF
C47762 AND2X1_LOC_739/a_8_24# AND2X1_LOC_740/B 0.01fF
C49174 AND2X1_LOC_740/B AND2X1_LOC_738/Y 0.09fF
C52704 VDD AND2X1_LOC_740/B 0.07fF
C57692 AND2X1_LOC_740/B VSS 0.13fF
C3728 AND2X1_LOC_722/Y AND2X1_LOC_733/a_8_24# 0.18fF
C7768 AND2X1_LOC_722/Y AND2X1_LOC_222/Y 0.01fF
C16357 AND2X1_LOC_722/a_8_24# AND2X1_LOC_722/Y 0.01fF
C16831 AND2X1_LOC_722/Y VDD 0.21fF
C48861 AND2X1_LOC_722/Y AND2X1_LOC_723/Y 0.02fF
C58010 AND2X1_LOC_722/Y VSS -0.13fF
C1862 OR2X1_LOC_655/B OR2X1_LOC_655/A 0.07fF
C16227 OR2X1_LOC_662/A OR2X1_LOC_655/B 0.24fF
C17953 OR2X1_LOC_864/A OR2X1_LOC_655/B 0.02fF
C34412 OR2X1_LOC_655/a_8_216# OR2X1_LOC_655/B 0.08fF
C46993 OR2X1_LOC_655/B OR2X1_LOC_649/a_8_216# 0.04fF
C54873 VDD OR2X1_LOC_655/B 0.26fF
C57283 OR2X1_LOC_655/B VSS 0.11fF
C50477 VDD D_GATE_811 0.06fF
C57678 D_GATE_811 VSS 0.18fF
C585 OR2X1_LOC_579/B OR2X1_LOC_579/a_8_216# 0.04fF
C4543 VDD OR2X1_LOC_579/B 0.06fF
C11682 OR2X1_LOC_579/B OR2X1_LOC_579/a_36_216# 0.02fF
C17195 OR2X1_LOC_579/B OR2X1_LOC_580/A 0.01fF
C56547 OR2X1_LOC_579/B VSS 0.18fF
C12023 VDD OR2X1_LOC_366/Y 0.65fF
C16645 OR2X1_LOC_577/Y OR2X1_LOC_366/Y 0.47fF
C24667 OR2X1_LOC_580/A OR2X1_LOC_366/Y 0.01fF
C34964 OR2X1_LOC_811/A OR2X1_LOC_366/Y 0.08fF
C38669 OR2X1_LOC_580/B OR2X1_LOC_366/Y 0.10fF
C39018 OR2X1_LOC_366/Y OR2X1_LOC_367/a_8_216# 0.01fF
C39510 OR2X1_LOC_562/A OR2X1_LOC_366/Y 0.03fF
C47703 OR2X1_LOC_367/B OR2X1_LOC_366/Y 0.23fF
C56258 OR2X1_LOC_366/Y VSS 0.41fF
C21833 AND2X1_LOC_660/Y AND2X1_LOC_662/a_8_24# 0.09fF
C31367 VDD AND2X1_LOC_660/Y 0.21fF
C57115 AND2X1_LOC_660/Y VSS 0.08fF
C5732 AND2X1_LOC_218/Y AND2X1_LOC_219/Y 0.11fF
C6354 AND2X1_LOC_660/a_8_24# AND2X1_LOC_218/Y 0.20fF
C11317 AND2X1_LOC_218/Y AND2X1_LOC_222/a_8_24# 0.11fF
C22161 AND2X1_LOC_663/B AND2X1_LOC_218/Y 0.23fF
C26159 VDD AND2X1_LOC_218/Y 0.38fF
C26816 AND2X1_LOC_660/A AND2X1_LOC_218/Y 0.09fF
C56561 AND2X1_LOC_218/Y VSS -0.06fF
C1747 AND2X1_LOC_808/A AND2X1_LOC_469/Y 0.02fF
C4412 AND2X1_LOC_469/Y AND2X1_LOC_220/a_8_24# 0.20fF
C15488 VDD AND2X1_LOC_469/Y 0.21fF
C18903 AND2X1_LOC_469/Y AND2X1_LOC_469/a_8_24# 0.01fF
C37017 AND2X1_LOC_469/Y AND2X1_LOC_220/B 0.01fF
C42799 AND2X1_LOC_469/Y AND2X1_LOC_220/Y 0.16fF
C49626 AND2X1_LOC_469/Y AND2X1_LOC_212/Y 0.23fF
C56678 AND2X1_LOC_469/Y VSS 0.11fF
C8131 OR2X1_LOC_571/Y OR2X1_LOC_579/A 0.89fF
C8308 OR2X1_LOC_865/B OR2X1_LOC_571/Y 0.07fF
C16281 VDD OR2X1_LOC_571/Y -0.00fF
C41308 OR2X1_LOC_571/B OR2X1_LOC_571/Y 0.01fF
C42032 OR2X1_LOC_571/Y OR2X1_LOC_576/a_8_216# 0.03fF
C56492 OR2X1_LOC_571/Y VSS 0.11fF
C1509 AND2X1_LOC_200/a_8_24# AND2X1_LOC_207/B 0.01fF
C21967 AND2X1_LOC_207/a_8_24# AND2X1_LOC_207/B 0.01fF
C29521 VDD AND2X1_LOC_207/B 0.01fF
C56555 AND2X1_LOC_207/B VSS 0.10fF
C12985 OR2X1_LOC_571/B OR2X1_LOC_579/A 0.02fF
C13183 OR2X1_LOC_865/B OR2X1_LOC_571/B 0.02fF
C21173 VDD OR2X1_LOC_571/B 0.20fF
C24991 OR2X1_LOC_658/a_8_216# OR2X1_LOC_571/B 0.40fF
C35957 OR2X1_LOC_571/a_8_216# OR2X1_LOC_571/B 0.10fF
C56765 OR2X1_LOC_571/B VSS 0.28fF
C5415 OR2X1_LOC_807/Y OR2X1_LOC_807/B 0.84fF
C9687 VDD OR2X1_LOC_807/B -0.00fF
C32612 OR2X1_LOC_807/B OR2X1_LOC_811/A 0.05fF
C34298 OR2X1_LOC_807/B OR2X1_LOC_807/A 0.19fF
C47748 OR2X1_LOC_807/B OR2X1_LOC_807/a_8_216# 0.01fF
C57424 OR2X1_LOC_807/B VSS -0.02fF
C7321 OR2X1_LOC_864/A OR2X1_LOC_649/a_8_216# 0.01fF
C14447 OR2X1_LOC_864/A OR2X1_LOC_663/A 14.17fF
C15205 OR2X1_LOC_864/A VDD 0.37fF
C18405 OR2X1_LOC_864/A OR2X1_LOC_655/A 0.01fF
C57905 OR2X1_LOC_864/A VSS -0.59fF
C26410 VDD OR2X1_LOC_358/A 0.25fF
C44279 OR2X1_LOC_648/A OR2X1_LOC_358/A 0.01fF
C45777 OR2X1_LOC_351/a_8_216# OR2X1_LOC_358/A 0.01fF
C54637 OR2X1_LOC_219/B OR2X1_LOC_358/A 0.07fF
C56478 OR2X1_LOC_358/A VSS -0.48fF
C10552 VDD AND2X1_LOC_575/Y 0.25fF
C24199 AND2X1_LOC_570/Y AND2X1_LOC_575/Y 0.01fF
C30568 AND2X1_LOC_575/Y AND2X1_LOC_576/Y 0.27fF
C36062 AND2X1_LOC_575/Y AND2X1_LOC_579/a_8_24# 0.19fF
C57746 AND2X1_LOC_575/Y VSS 0.10fF
C9133 OR2X1_LOC_732/B OR2X1_LOC_732/A 0.13fF
C19075 OR2X1_LOC_808/B OR2X1_LOC_732/B 0.10fF
C19525 OR2X1_LOC_732/a_8_216# OR2X1_LOC_732/B 0.04fF
C22040 VDD OR2X1_LOC_732/B 0.04fF
C56515 OR2X1_LOC_732/B VSS 0.14fF
C28045 OR2X1_LOC_510/Y OR2X1_LOC_657/a_8_216# 0.01fF
C34462 OR2X1_LOC_510/Y OR2X1_LOC_205/Y 0.25fF
C57397 OR2X1_LOC_510/Y VSS 0.05fF
C10268 OR2X1_LOC_219/B OR2X1_LOC_358/B 0.01fF
C26333 OR2X1_LOC_358/a_8_216# OR2X1_LOC_358/B 0.02fF
C31812 OR2X1_LOC_358/a_36_216# OR2X1_LOC_358/B 0.03fF
C38036 VDD OR2X1_LOC_358/B 0.15fF
C40267 OR2X1_LOC_222/A OR2X1_LOC_358/B 0.72fF
C56105 OR2X1_LOC_648/A OR2X1_LOC_358/B 0.01fF
C56539 OR2X1_LOC_358/B VSS 0.24fF
C1900 OR2X1_LOC_853/a_8_216# OR2X1_LOC_35/Y 0.03fF
C12986 OR2X1_LOC_857/A OR2X1_LOC_35/Y 0.04fF
C56695 OR2X1_LOC_35/Y VSS 0.24fF
C7613 AND2X1_LOC_805/Y AND2X1_LOC_807/a_8_24# 0.01fF
C11011 AND2X1_LOC_807/Y AND2X1_LOC_805/Y 0.01fF
C17340 AND2X1_LOC_866/B AND2X1_LOC_805/Y 0.02fF
C24664 AND2X1_LOC_580/B AND2X1_LOC_805/Y 0.03fF
C49717 VDD AND2X1_LOC_805/Y 0.36fF
C56703 AND2X1_LOC_805/Y VSS -0.00fF
C12220 AND2X1_LOC_861/B AND2X1_LOC_865/a_8_24# 0.01fF
C19513 AND2X1_LOC_580/A AND2X1_LOC_861/B 0.07fF
C20712 AND2X1_LOC_861/B AND2X1_LOC_663/A 0.10fF
C23365 AND2X1_LOC_861/B AND2X1_LOC_862/A 0.01fF
C50104 VDD AND2X1_LOC_861/B 0.01fF
C54298 AND2X1_LOC_861/B AND2X1_LOC_861/a_8_24# 0.01fF
C54831 AND2X1_LOC_861/B AND2X1_LOC_862/a_8_24# 0.01fF
C57398 AND2X1_LOC_861/B VSS 0.27fF
C6870 OR2X1_LOC_865/A OR2X1_LOC_580/A 0.09fF
C33788 OR2X1_LOC_865/A OR2X1_LOC_865/a_8_216# 0.14fF
C42245 OR2X1_LOC_865/B OR2X1_LOC_865/A 2.15fF
C50461 OR2X1_LOC_865/A VDD 0.07fF
C57949 OR2X1_LOC_865/A VSS 0.15fF
C30157 AND2X1_LOC_862/a_8_24# AND2X1_LOC_862/A 0.10fF
C52267 AND2X1_LOC_862/A AND2X1_LOC_663/A 0.45fF
C56934 AND2X1_LOC_862/A VSS 0.25fF
C4778 OR2X1_LOC_363/B OR2X1_LOC_580/A 0.01fF
C58031 OR2X1_LOC_363/B VSS 0.23fF
C15928 AND2X1_LOC_363/Y AND2X1_LOC_860/A 0.03fF
C35258 AND2X1_LOC_860/A AND2X1_LOC_562/Y 0.10fF
C35869 AND2X1_LOC_860/a_8_24# AND2X1_LOC_860/A 0.08fF
C38860 AND2X1_LOC_360/a_8_24# AND2X1_LOC_860/A 0.06fF
C43547 VDD AND2X1_LOC_860/A 0.58fF
C44956 AND2X1_LOC_363/A AND2X1_LOC_860/A 0.03fF
C56562 AND2X1_LOC_860/A VSS 0.24fF
C4295 AND2X1_LOC_212/A AND2X1_LOC_222/Y 0.01fF
C14576 AND2X1_LOC_212/A AND2X1_LOC_212/a_8_24# 0.09fF
C49660 AND2X1_LOC_212/A AND2X1_LOC_364/Y 0.59fF
C55101 AND2X1_LOC_212/A AND2X1_LOC_365/a_8_24# 0.01fF
C57844 AND2X1_LOC_212/A VSS 0.29fF
C16416 AND2X1_LOC_364/Y AND2X1_LOC_857/Y 0.12fF
C33925 AND2X1_LOC_857/Y AND2X1_LOC_654/a_8_24# 0.01fF
C36303 VDD AND2X1_LOC_857/Y 0.29fF
C53623 AND2X1_LOC_857/Y AND2X1_LOC_853/Y 0.13fF
C57235 AND2X1_LOC_857/Y VSS 0.08fF
C3656 AND2X1_LOC_574/A AND2X1_LOC_657/A 0.16fF
C8565 AND2X1_LOC_574/A AND2X1_LOC_657/Y 0.15fF
C21389 AND2X1_LOC_807/Y AND2X1_LOC_574/A 0.03fF
C23937 AND2X1_LOC_576/Y AND2X1_LOC_574/A 0.02fF
C39184 AND2X1_LOC_574/A AND2X1_LOC_657/a_36_24# 0.01fF
C56812 AND2X1_LOC_574/A VSS 0.17fF
C2139 AND2X1_LOC_723/Y AND2X1_LOC_578/A 0.07fF
C4144 AND2X1_LOC_578/A AND2X1_LOC_212/Y 0.01fF
C11025 AND2X1_LOC_578/A AND2X1_LOC_851/a_8_24# 0.03fF
C12837 AND2X1_LOC_578/A AND2X1_LOC_569/a_8_24# 0.03fF
C17190 AND2X1_LOC_578/A AND2X1_LOC_222/Y 0.03fF
C18364 AND2X1_LOC_578/A AND2X1_LOC_577/A 0.11fF
C26283 VDD AND2X1_LOC_578/A 0.14fF
C28522 AND2X1_LOC_569/A AND2X1_LOC_578/A 0.06fF
C29763 AND2X1_LOC_577/Y AND2X1_LOC_578/A 0.04fF
C30964 AND2X1_LOC_578/A AND2X1_LOC_657/Y 0.10fF
C43800 AND2X1_LOC_578/A AND2X1_LOC_807/Y 0.07fF
C53185 AND2X1_LOC_578/A AND2X1_LOC_663/A 0.10fF
C57741 AND2X1_LOC_578/A VSS 0.26fF
C8071 AND2X1_LOC_571/Y AND2X1_LOC_572/Y 0.12fF
C8764 AND2X1_LOC_571/A AND2X1_LOC_571/Y 0.26fF
C13614 AND2X1_LOC_571/Y AND2X1_LOC_576/a_8_24# 0.18fF
C50010 AND2X1_LOC_571/Y AND2X1_LOC_563/Y 0.01fF
C52514 AND2X1_LOC_571/Y AND2X1_LOC_657/A 0.02fF
C52661 AND2X1_LOC_571/Y VDD 0.25fF
C57918 AND2X1_LOC_571/Y VSS 0.10fF
C3832 AND2X1_LOC_363/B AND2X1_LOC_363/A 0.10fF
C6808 AND2X1_LOC_367/a_8_24# AND2X1_LOC_363/A 0.20fF
C25831 AND2X1_LOC_363/Y AND2X1_LOC_363/A 0.10fF
C37179 AND2X1_LOC_363/a_8_24# AND2X1_LOC_363/A 0.03fF
C48968 AND2X1_LOC_360/a_8_24# AND2X1_LOC_363/A 0.02fF
C49470 AND2X1_LOC_359/a_8_24# AND2X1_LOC_363/A 0.01fF
C53568 VDD AND2X1_LOC_363/A 0.21fF
C57414 AND2X1_LOC_363/A VSS 0.24fF
C30531 OR2X1_LOC_341/Y OR2X1_LOC_350/a_8_216# 0.39fF
C43465 OR2X1_LOC_341/Y OR2X1_LOC_341/a_8_216# -0.00fF
C56541 OR2X1_LOC_341/Y VSS 0.18fF
C21815 AND2X1_LOC_470/a_8_24# AND2X1_LOC_470/A 0.19fF
C34664 VDD AND2X1_LOC_470/A 0.25fF
C56727 AND2X1_LOC_470/A VSS 0.10fF
C6144 VDD AND2X1_LOC_658/Y 0.26fF
C27432 AND2X1_LOC_658/Y AND2X1_LOC_659/a_8_24# 0.01fF
C32912 AND2X1_LOC_658/Y AND2X1_LOC_663/A 0.01fF
C38829 AND2X1_LOC_658/a_8_24# AND2X1_LOC_658/Y 0.01fF
C56682 AND2X1_LOC_658/Y VSS 0.12fF
C10916 AND2X1_LOC_735/Y AND2X1_LOC_736/a_8_24# 0.11fF
C28698 AND2X1_LOC_735/Y VDD 0.16fF
C42276 AND2X1_LOC_735/Y AND2X1_LOC_570/Y 0.02fF
C42378 AND2X1_LOC_573/a_36_24# AND2X1_LOC_735/Y 0.01fF
C48936 AND2X1_LOC_735/Y AND2X1_LOC_576/Y 0.03fF
C57880 AND2X1_LOC_735/Y VSS -0.04fF
C12689 OR2X1_LOC_803/a_8_216# OR2X1_LOC_803/B 0.02fF
C34706 OR2X1_LOC_808/B OR2X1_LOC_803/B 0.73fF
C37590 VDD OR2X1_LOC_803/B 0.05fF
C56785 OR2X1_LOC_803/B VSS -0.02fF
C41027 AND2X1_LOC_562/Y AND2X1_LOC_563/Y 0.16fF
C43679 AND2X1_LOC_657/A AND2X1_LOC_562/Y 0.06fF
C43850 VDD AND2X1_LOC_562/Y 0.72fF
C46733 AND2X1_LOC_562/Y AND2X1_LOC_570/a_8_24# 0.17fF
C47760 AND2X1_LOC_562/a_8_24# AND2X1_LOC_562/Y 0.01fF
C56252 AND2X1_LOC_562/Y VSS 0.70fF
C54304 OR2X1_LOC_661/a_8_216# OR2X1_LOC_661/A 0.39fF
C57581 OR2X1_LOC_661/A VSS 0.18fF
C1514 VDD OR2X1_LOC_733/A 0.12fF
C17350 OR2X1_LOC_733/B OR2X1_LOC_733/A 0.08fF
C51431 OR2X1_LOC_722/a_8_216# OR2X1_LOC_733/A 0.01fF
C56569 OR2X1_LOC_733/A VSS 0.24fF
C1189 OR2X1_LOC_566/Y OR2X1_LOC_568/a_8_216# 0.03fF
C26508 OR2X1_LOC_468/Y OR2X1_LOC_566/Y 0.01fF
C56348 OR2X1_LOC_566/Y VSS 0.11fF
C23714 OR2X1_LOC_469/Y OR2X1_LOC_803/A 0.03fF
C36004 OR2X1_LOC_479/Y OR2X1_LOC_803/A 0.03fF
C45296 VDD OR2X1_LOC_803/A -0.00fF
C6191 OR2X1_LOC_364/B OR2X1_LOC_364/A 0.18fF
C10339 OR2X1_LOC_364/B OR2X1_LOC_212/B 0.01fF
C13808 OR2X1_LOC_364/B OR2X1_LOC_364/a_8_216# 0.05fF
C36595 OR2X1_LOC_364/B OR2X1_LOC_357/B 0.75fF
C53954 OR2X1_LOC_364/B OR2X1_LOC_479/Y 0.06fF
C58109 OR2X1_LOC_364/B VSS 0.21fF
C6153 OR2X1_LOC_738/B OR2X1_LOC_738/a_8_216# 0.39fF
C32525 VDD OR2X1_LOC_738/B -0.00fF
C47225 OR2X1_LOC_731/a_8_216# OR2X1_LOC_738/B -0.00fF
C52329 OR2X1_LOC_738/B OR2X1_LOC_738/A 0.15fF
C56725 OR2X1_LOC_738/B VSS 0.17fF
C5312 OR2X1_LOC_858/A OR2X1_LOC_735/a_8_216# 0.27fF
C14714 OR2X1_LOC_858/A VDD 1.33fF
C27329 OR2X1_LOC_858/A OR2X1_LOC_580/A 0.18fF
C57946 OR2X1_LOC_858/A VSS -1.81fF
C54378 AND2X1_LOC_569/A VDD 0.51fF
C57955 AND2X1_LOC_569/A VSS 0.05fF
C5674 AND2X1_LOC_469/B AND2X1_LOC_804/A 0.01fF
C5686 AND2X1_LOC_733/Y AND2X1_LOC_804/A 0.02fF
C17840 AND2X1_LOC_804/a_8_24# AND2X1_LOC_804/A -0.00fF
C34954 AND2X1_LOC_212/Y AND2X1_LOC_804/A 0.01fF
C56313 AND2X1_LOC_804/A VSS 0.26fF
C34418 AND2X1_LOC_566/Y AND2X1_LOC_568/a_8_24# 0.06fF
C43665 AND2X1_LOC_566/Y AND2X1_LOC_212/Y 0.34fF
C45577 AND2X1_LOC_566/Y AND2X1_LOC_568/a_36_24# 0.01fF
C57743 AND2X1_LOC_566/Y VSS 0.20fF
C3341 AND2X1_LOC_723/Y AND2X1_LOC_723/a_8_24# 0.04fF
C18849 AND2X1_LOC_723/Y AND2X1_LOC_222/Y 0.01fF
C27430 AND2X1_LOC_722/a_8_24# AND2X1_LOC_723/Y -0.00fF
C27866 AND2X1_LOC_723/Y VDD 0.52fF
C58009 AND2X1_LOC_723/Y VSS 0.05fF
C3339 OR2X1_LOC_477/Y OR2X1_LOC_469/Y 0.19fF
C23040 OR2X1_LOC_470/B OR2X1_LOC_477/Y 0.01fF
C56168 OR2X1_LOC_470/a_8_216# OR2X1_LOC_477/Y 0.01fF
C57273 OR2X1_LOC_477/Y VSS 0.11fF
C963 VDD AND2X1_LOC_206/Y 0.01fF
C11428 AND2X1_LOC_206/Y AND2X1_LOC_215/a_8_24# 0.03fF
C33483 AND2X1_LOC_206/Y AND2X1_LOC_215/a_36_24# 0.01fF
C40588 AND2X1_LOC_206/Y AND2X1_LOC_215/A 0.23fF
C56365 AND2X1_LOC_206/Y VSS 0.18fF
C7283 VDD AND2X1_LOC_795/Y 0.06fF
C24112 AND2X1_LOC_795/Y AND2X1_LOC_804/a_8_24# 0.11fF
C42903 AND2X1_LOC_795/Y AND2X1_LOC_795/a_8_24# 0.10fF
C54061 AND2X1_LOC_795/Y AND2X1_LOC_795/a_36_24# 0.01fF
C54306 AND2X1_LOC_795/Y AND2X1_LOC_222/Y 0.02fF
C56878 AND2X1_LOC_795/Y VSS 0.31fF
C16441 OR2X1_LOC_479/Y OR2X1_LOC_357/B 0.03fF
C25657 OR2X1_LOC_357/a_8_216# OR2X1_LOC_357/B 0.03fF
C25682 VDD OR2X1_LOC_357/B -0.00fF
C28978 OR2X1_LOC_357/B OR2X1_LOC_212/B 0.01fF
C56432 OR2X1_LOC_357/B VSS 0.11fF
C4246 OR2X1_LOC_219/B OR2X1_LOC_215/Y 0.05fF
C15312 OR2X1_LOC_219/B OR2X1_LOC_219/a_8_216# 0.02fF
C20902 OR2X1_LOC_219/B OR2X1_LOC_219/a_36_216# 0.01fF
C24204 VDD OR2X1_LOC_219/B 0.13fF
C26349 OR2X1_LOC_219/B OR2X1_LOC_222/A 0.17fF
C41948 OR2X1_LOC_648/A OR2X1_LOC_219/B 0.07fF
C43481 OR2X1_LOC_219/B OR2X1_LOC_351/a_8_216# 0.13fF
C55364 OR2X1_LOC_219/B OR2X1_LOC_350/a_36_216# 0.02fF
C56993 OR2X1_LOC_219/B VSS 0.47fF
C57337 OR2X1_LOC_659/A VSS 0.25fF
C2935 OR2X1_LOC_865/B OR2X1_LOC_571/a_8_216# 0.06fF
C13812 OR2X1_LOC_865/B OR2X1_LOC_576/a_8_216# 0.04fF
C25021 OR2X1_LOC_861/a_8_216# OR2X1_LOC_865/B 0.04fF
C27532 OR2X1_LOC_860/a_8_216# OR2X1_LOC_865/B 0.06fF
C27588 OR2X1_LOC_865/B OR2X1_LOC_865/a_8_216# 0.04fF
C33062 OR2X1_LOC_865/B OR2X1_LOC_865/a_36_216# 0.02fF
C35811 OR2X1_LOC_865/B OR2X1_LOC_579/A 0.16fF
C44051 OR2X1_LOC_865/B VDD 0.01fF
C57986 OR2X1_LOC_865/B VSS 0.36fF
C30586 AND2X1_LOC_650/Y AND2X1_LOC_654/a_8_24# 0.07fF
C32997 VDD AND2X1_LOC_650/Y 0.21fF
C51575 AND2X1_LOC_650/a_8_24# AND2X1_LOC_650/Y 0.01fF
C56965 AND2X1_LOC_650/Y VSS 0.13fF
C10694 VDD AND2X1_LOC_796/Y 0.21fF
C15332 AND2X1_LOC_796/Y AND2X1_LOC_657/Y 0.03fF
C17883 AND2X1_LOC_738/B AND2X1_LOC_796/Y 0.02fF
C37351 AND2X1_LOC_796/Y AND2X1_LOC_663/A 0.03fF
C41795 AND2X1_LOC_796/Y AND2X1_LOC_803/a_8_24# 0.10fF
C56937 AND2X1_LOC_796/Y VSS 0.02fF
C741 AND2X1_LOC_212/Y AND2X1_LOC_212/B 0.02fF
C22988 VDD AND2X1_LOC_212/B 0.26fF
C24070 AND2X1_LOC_212/B AND2X1_LOC_212/a_8_24# 0.05fF
C39594 AND2X1_LOC_864/a_8_24# AND2X1_LOC_212/B 0.20fF
C45199 AND2X1_LOC_866/A AND2X1_LOC_212/B 0.01fF
C56558 AND2X1_LOC_212/B VSS 0.13fF
C13158 VDD AND2X1_LOC_853/Y 0.05fF
C35673 AND2X1_LOC_853/Y AND2X1_LOC_857/a_8_24# 0.05fF
C56979 AND2X1_LOC_853/Y VSS 0.19fF
C10436 AND2X1_LOC_219/a_8_24# AND2X1_LOC_219/A 0.07fF
C45245 VDD AND2X1_LOC_219/A 0.29fF
C56405 AND2X1_LOC_219/A VSS 0.22fF
C15528 AND2X1_LOC_357/A AND2X1_LOC_364/Y 0.01fF
C35380 AND2X1_LOC_357/A VDD -0.00fF
C54721 AND2X1_LOC_357/A AND2X1_LOC_357/a_8_24# 0.07fF
C57843 AND2X1_LOC_357/A VSS 0.22fF
C36185 OR2X1_LOC_808/B OR2X1_LOC_732/A 0.72fF
C36601 OR2X1_LOC_732/a_8_216# OR2X1_LOC_732/A 0.04fF
C39147 VDD OR2X1_LOC_732/A 0.30fF
C56464 OR2X1_LOC_732/A VSS 0.21fF
C2622 AND2X1_LOC_578/a_8_24# AND2X1_LOC_577/A 0.20fF
C12708 AND2X1_LOC_577/a_8_24# AND2X1_LOC_577/A 0.07fF
C13653 AND2X1_LOC_580/A AND2X1_LOC_577/A 0.02fF
C44099 VDD AND2X1_LOC_577/A 0.21fF
C57682 AND2X1_LOC_577/A VSS 0.22fF
C8116 AND2X1_LOC_571/A AND2X1_LOC_657/A 0.03fF
C19813 AND2X1_LOC_571/A AND2X1_LOC_572/Y 0.20fF
C25314 AND2X1_LOC_571/A AND2X1_LOC_576/a_8_24# 0.09fF
C58116 AND2X1_LOC_571/A VSS 0.29fF
C16622 AND2X1_LOC_35/Y AND2X1_LOC_853/a_8_24# 0.06fF
C36631 AND2X1_LOC_649/Y AND2X1_LOC_655/a_8_24# 0.13fF
C41618 VDD AND2X1_LOC_649/Y 0.01fF
C56919 AND2X1_LOC_649/Y VSS -0.17fF
C279 OR2X1_LOC_223/A OR2X1_LOC_367/B 0.03fF
C2582 OR2X1_LOC_367/B OR2X1_LOC_367/a_8_216# 0.33fF
C31522 VDD OR2X1_LOC_367/B 1.52fF
C41706 OR2X1_LOC_741/Y OR2X1_LOC_367/B 0.03fF
C56157 OR2X1_LOC_365/a_8_216# OR2X1_LOC_367/B 0.09fF
C56339 OR2X1_LOC_367/B VSS 0.81fF
C1181 OR2X1_LOC_478/Y OR2X1_LOC_470/B 0.02fF
C6657 OR2X1_LOC_480/a_8_216# OR2X1_LOC_470/B 0.01fF
C17729 D_GATE_479 OR2X1_LOC_470/B 0.75fF
C28476 OR2X1_LOC_470/B OR2X1_LOC_469/Y 0.03fF
C31502 OR2X1_LOC_466/a_8_216# OR2X1_LOC_470/B -0.00fF
C33959 OR2X1_LOC_470/B OR2X1_LOC_478/a_8_216# 0.01fF
C57322 OR2X1_LOC_470/B VSS 0.14fF
C463 OR2X1_LOC_479/Y OR2X1_LOC_469/a_8_216# 0.03fF
C1040 OR2X1_LOC_479/Y OR2X1_LOC_804/A 0.02fF
C5980 OR2X1_LOC_479/Y OR2X1_LOC_469/a_36_216# 0.02fF
C6356 OR2X1_LOC_479/Y OR2X1_LOC_738/A 0.07fF
C11644 OR2X1_LOC_479/Y OR2X1_LOC_223/A 1.05fF
C14984 OR2X1_LOC_479/Y OR2X1_LOC_794/a_8_216# -0.03fF
C21308 OR2X1_LOC_479/Y OR2X1_LOC_469/Y 7.71fF
C23887 OR2X1_LOC_479/Y OR2X1_LOC_212/A 0.03fF
C24017 OR2X1_LOC_479/Y OR2X1_LOC_364/a_36_216# 0.02fF
C25999 OR2X1_LOC_479/Y OR2X1_LOC_804/B 0.17fF
C29271 OR2X1_LOC_479/Y OR2X1_LOC_804/a_8_216# 0.02fF
C34777 OR2X1_LOC_479/Y OR2X1_LOC_804/a_36_216# 0.01fF
C39863 OR2X1_LOC_479/Y OR2X1_LOC_808/B 0.10fF
C40244 OR2X1_LOC_479/Y OR2X1_LOC_808/A 0.12fF
C40433 OR2X1_LOC_479/Y OR2X1_LOC_795/a_8_216# 0.01fF
C42072 OR2X1_LOC_364/A OR2X1_LOC_479/Y 0.39fF
C42793 OR2X1_LOC_357/a_8_216# OR2X1_LOC_479/Y 0.05fF
C42851 OR2X1_LOC_479/Y VDD 1.06fF
C45549 OR2X1_LOC_479/Y OR2X1_LOC_468/Y 5.32fF
C46189 OR2X1_LOC_479/Y OR2X1_LOC_212/B 0.03fF
C49788 OR2X1_LOC_479/Y OR2X1_LOC_364/a_8_216# 0.02fF
C50151 OR2X1_LOC_479/Y OR2X1_LOC_478/Y 0.13fF
C57831 OR2X1_LOC_479/Y VSS 0.60fF
C1788 VDD OR2X1_LOC_741/A -0.00fF
C4270 OR2X1_LOC_741/a_8_216# OR2X1_LOC_741/A 0.39fF
C52630 OR2X1_LOC_737/a_8_216# OR2X1_LOC_741/A -0.00fF
C54918 OR2X1_LOC_736/Y OR2X1_LOC_741/A 0.06fF
C56416 OR2X1_LOC_741/A VSS 0.18fF
C1149 OR2X1_LOC_739/Y OR2X1_LOC_740/a_8_216# 0.39fF
C36493 OR2X1_LOC_739/Y OR2X1_LOC_740/B 0.08fF
C46479 VDD OR2X1_LOC_739/Y -0.00fF
C48881 OR2X1_LOC_739/Y OR2X1_LOC_739/a_8_216# -0.00fF
C56844 OR2X1_LOC_739/Y VSS 0.18fF
C20988 OR2X1_LOC_223/B OR2X1_LOC_223/A 0.17fF
C49955 OR2X1_LOC_223/B OR2X1_LOC_223/a_8_216# 0.05fF
C57199 OR2X1_LOC_223/B VSS 0.21fF
C4001 OR2X1_LOC_223/A OR2X1_LOC_804/B 0.09fF
C7314 OR2X1_LOC_794/a_8_216# OR2X1_LOC_804/B 0.01fF
C21717 OR2X1_LOC_804/a_8_216# OR2X1_LOC_804/B 0.01fF
C32657 OR2X1_LOC_808/A OR2X1_LOC_804/B 0.93fF
C35142 VDD OR2X1_LOC_804/B 0.27fF
C49610 OR2X1_LOC_804/B OR2X1_LOC_804/A 0.07fF
C56894 OR2X1_LOC_804/B VSS -0.01fF
C9794 OR2X1_LOC_662/A OR2X1_LOC_660/B 0.03fF
C12704 OR2X1_LOC_662/A OR2X1_LOC_663/A 0.01fF
C13519 OR2X1_LOC_662/A VDD 0.09fF
C46746 OR2X1_LOC_662/A OR2X1_LOC_662/a_8_216# 0.01fF
C49390 OR2X1_LOC_662/A OR2X1_LOC_655/a_8_216# 0.02fF
C57835 OR2X1_LOC_662/A VSS 0.12fF
C2057 OR2X1_LOC_358/a_8_216# OR2X1_LOC_648/A 0.03fF
C13152 OR2X1_LOC_364/A OR2X1_LOC_648/A 0.02fF
C13876 VDD OR2X1_LOC_648/A 0.12fF
C57456 OR2X1_LOC_648/A VSS 0.33fF
C14691 OR2X1_LOC_200/Y OR2X1_LOC_207/a_8_216# 0.39fF
C56802 OR2X1_LOC_200/Y VSS 0.18fF
C52574 OR2X1_LOC_657/a_8_216# OR2X1_LOC_217/A 0.39fF
C56286 OR2X1_LOC_217/A VSS 0.36fF
C18292 OR2X1_LOC_468/Y OR2X1_LOC_738/A 0.01fF
C19131 OR2X1_LOC_468/Y OR2X1_LOC_211/a_8_216# 0.01fF
C31921 OR2X1_LOC_468/a_8_216# OR2X1_LOC_468/Y 0.01fF
C31951 OR2X1_LOC_468/Y OR2X1_LOC_568/a_8_216# 0.01fF
C35620 OR2X1_LOC_468/Y OR2X1_LOC_212/A 0.57fF
C40001 OR2X1_LOC_468/Y OR2X1_LOC_566/a_8_216# 0.01fF
C51902 OR2X1_LOC_808/B OR2X1_LOC_468/Y 0.05fF
C54787 VDD OR2X1_LOC_468/Y 0.25fF
C57162 OR2X1_LOC_468/Y VSS 0.53fF
C14502 OR2X1_LOC_562/Y OR2X1_LOC_562/A 0.14fF
C17176 OR2X1_LOC_562/a_8_216# OR2X1_LOC_562/A 0.18fF
C23601 VDD OR2X1_LOC_562/A 0.28fF
C36616 OR2X1_LOC_563/a_8_216# OR2X1_LOC_562/A 0.02fF
C44852 OR2X1_LOC_570/a_8_216# OR2X1_LOC_562/A 0.01fF
C50432 OR2X1_LOC_562/A OR2X1_LOC_580/B 0.03fF
C56401 OR2X1_LOC_562/A VSS 0.30fF
C506 AND2X1_LOC_657/Y AND2X1_LOC_657/A 0.01fF
C1762 AND2X1_LOC_571/a_8_24# AND2X1_LOC_657/A 0.01fF
C6690 AND2X1_LOC_657/A AND2X1_LOC_217/a_8_24# 0.02fF
C12950 AND2X1_LOC_576/a_8_24# AND2X1_LOC_657/A 0.02fF
C13380 AND2X1_LOC_807/Y AND2X1_LOC_657/A 0.10fF
C15874 AND2X1_LOC_576/Y AND2X1_LOC_657/A 0.01fF
C18111 AND2X1_LOC_866/A AND2X1_LOC_657/A 0.07fF
C21481 AND2X1_LOC_580/A AND2X1_LOC_657/A 0.07fF
C22733 AND2X1_LOC_663/A AND2X1_LOC_657/A 0.10fF
C39538 AND2X1_LOC_217/Y AND2X1_LOC_657/A 0.83fF
C44224 AND2X1_LOC_572/a_8_24# AND2X1_LOC_657/A 0.01fF
C47939 AND2X1_LOC_663/B AND2X1_LOC_657/A 0.10fF
C49143 AND2X1_LOC_563/a_8_24# AND2X1_LOC_657/A 0.04fF
C49335 AND2X1_LOC_657/A AND2X1_LOC_563/Y 0.02fF
C52032 VDD AND2X1_LOC_657/A 0.05fF
C54795 AND2X1_LOC_657/A AND2X1_LOC_570/a_8_24# 0.01fF
C56278 AND2X1_LOC_657/A VSS 0.26fF
C4003 AND2X1_LOC_341/a_8_24# AND2X1_LOC_350/B 0.04fF
C30739 AND2X1_LOC_350/B VDD 0.19fF
C31158 AND2X1_LOC_350/a_8_24# AND2X1_LOC_350/B 0.01fF
C54188 AND2X1_LOC_351/a_8_24# AND2X1_LOC_350/B 0.01fF
C57845 AND2X1_LOC_350/B VSS -0.25fF
C161 AND2X1_LOC_469/B AND2X1_LOC_794/a_8_24# 0.01fF
C644 VDD AND2X1_LOC_469/B 0.27fF
C1173 AND2X1_LOC_811/B AND2X1_LOC_469/B 0.01fF
C3899 AND2X1_LOC_811/Y AND2X1_LOC_469/B 0.02fF
C5285 AND2X1_LOC_657/Y AND2X1_LOC_469/B 0.03fF
C27441 AND2X1_LOC_663/A AND2X1_LOC_469/B 0.05fF
C34544 AND2X1_LOC_212/Y AND2X1_LOC_469/B 0.01fF
C42947 AND2X1_LOC_808/A AND2X1_LOC_469/B 0.02fF
C46656 AND2X1_LOC_477/a_8_24# AND2X1_LOC_469/B 0.01fF
C51838 AND2X1_LOC_808/a_8_24# AND2X1_LOC_469/B 0.01fF
C56626 AND2X1_LOC_469/B VSS 0.05fF
C34186 VDD AND2X1_LOC_562/B 0.04fF
C57813 AND2X1_LOC_562/B VSS 0.19fF
C13912 AND2X1_LOC_205/a_8_24# AND2X1_LOC_215/A 0.01fF
C35691 VDD AND2X1_LOC_215/A 0.06fF
C56318 AND2X1_LOC_215/A VSS 0.21fF
C24785 AND2X1_LOC_648/B AND2X1_LOC_648/a_8_24# 0.11fF
C41627 VDD AND2X1_LOC_648/B 0.30fF
C56861 AND2X1_LOC_648/B VSS 0.25fF
C3415 AND2X1_LOC_576/a_8_24# AND2X1_LOC_573/A 0.02fF
C5131 AND2X1_LOC_573/A AND2X1_LOC_657/a_8_24# 0.01fF
C8659 AND2X1_LOC_866/A AND2X1_LOC_573/A 0.07fF
C11903 AND2X1_LOC_580/A AND2X1_LOC_573/A 0.03fF
C13138 AND2X1_LOC_573/A AND2X1_LOC_663/A 0.05fF
C34570 AND2X1_LOC_572/a_8_24# AND2X1_LOC_573/A 0.03fF
C39430 AND2X1_LOC_563/a_8_24# AND2X1_LOC_573/A 0.03fF
C42330 VDD AND2X1_LOC_573/A 1.84fF
C45206 AND2X1_LOC_573/A AND2X1_LOC_570/a_8_24# 0.03fF
C47175 AND2X1_LOC_573/A AND2X1_LOC_657/Y 0.09fF
C54017 AND2X1_LOC_572/Y AND2X1_LOC_573/A 0.08fF
C56909 AND2X1_LOC_573/A VSS 0.05fF
C2455 AND2X1_LOC_363/B VDD 0.24fF
C30852 AND2X1_LOC_363/B AND2X1_LOC_363/Y 0.03fF
C42262 AND2X1_LOC_363/B AND2X1_LOC_363/a_8_24# 0.19fF
C57984 AND2X1_LOC_363/B VSS -0.09fF
C32876 AND2X1_LOC_217/Y AND2X1_LOC_218/a_8_24# 0.03fF
C39663 AND2X1_LOC_217/Y VDD 0.05fF
C58137 AND2X1_LOC_217/Y VSS -0.01fF
C4626 AND2X1_LOC_563/a_8_24# AND2X1_LOC_572/Y 0.02fF
C4806 AND2X1_LOC_572/Y AND2X1_LOC_563/Y 0.54fF
C7540 AND2X1_LOC_572/Y VDD 0.33fF
C13460 AND2X1_LOC_571/a_8_24# AND2X1_LOC_572/Y 0.01fF
C29819 AND2X1_LOC_572/Y AND2X1_LOC_866/A 0.03fF
C57917 AND2X1_LOC_572/Y VSS 0.05fF
C1045 AND2X1_LOC_731/Y AND2X1_LOC_220/B 0.03fF
C4346 AND2X1_LOC_731/a_8_24# AND2X1_LOC_220/B 0.07fF
C6471 AND2X1_LOC_220/a_8_24# AND2X1_LOC_220/B 0.01fF
C17573 VDD AND2X1_LOC_220/B 0.40fF
C25159 AND2X1_LOC_220/B AND2X1_LOC_740/a_8_24# 0.07fF
C36204 AND2X1_LOC_797/a_8_24# AND2X1_LOC_220/B 0.20fF
C44887 AND2X1_LOC_220/Y AND2X1_LOC_220/B 0.15fF
C47483 AND2X1_LOC_803/B AND2X1_LOC_220/B 0.03fF
C48339 AND2X1_LOC_478/a_8_24# AND2X1_LOC_220/B 0.02fF
C56449 AND2X1_LOC_220/B VSS -0.20fF
C21509 AND2X1_LOC_742/a_8_24# AND2X1_LOC_731/Y 0.19fF
C21788 AND2X1_LOC_731/Y AND2X1_LOC_808/A 0.32fF
C22331 AND2X1_LOC_731/a_8_24# AND2X1_LOC_731/Y 0.02fF
C35389 VDD AND2X1_LOC_731/Y 0.21fF
C35401 AND2X1_LOC_731/Y AND2X1_LOC_738/a_8_24# 0.09fF
C42711 AND2X1_LOC_738/B AND2X1_LOC_731/Y 0.02fF
C48694 AND2X1_LOC_731/Y AND2X1_LOC_742/A 0.23fF
C57756 AND2X1_LOC_731/Y VSS -0.20fF
C898 AND2X1_LOC_803/B AND2X1_LOC_803/a_8_24# 0.11fF
C25729 AND2X1_LOC_803/B VDD 0.18fF
C32892 AND2X1_LOC_803/B AND2X1_LOC_738/B 0.06fF
C58079 AND2X1_LOC_803/B VSS 0.22fF
C10389 AND2X1_LOC_576/a_8_24# AND2X1_LOC_563/Y 0.01fF
C13389 AND2X1_LOC_576/Y AND2X1_LOC_563/Y 0.01fF
C15539 AND2X1_LOC_866/A AND2X1_LOC_563/Y 0.03fF
C49528 VDD AND2X1_LOC_563/Y 0.38fF
C55372 AND2X1_LOC_571/a_8_24# AND2X1_LOC_563/Y 0.01fF
C56251 AND2X1_LOC_563/Y VSS 0.05fF
C2091 D_GATE_741 OR2X1_LOC_564/B 0.02fF
C17966 OR2X1_LOC_223/a_8_216# OR2X1_LOC_564/B 0.40fF
C20353 VDD OR2X1_LOC_564/B 0.08fF
C45195 OR2X1_LOC_223/A OR2X1_LOC_564/B 0.62fF
C56656 OR2X1_LOC_564/B VSS 0.40fF
C3287 VDD OR2X1_LOC_736/A 0.03fF
C11174 OR2X1_LOC_736/A OR2X1_LOC_736/a_8_216# 0.04fF
C50147 OR2X1_LOC_735/a_8_216# OR2X1_LOC_736/A -0.00fF
C56510 OR2X1_LOC_736/A VSS 0.22fF
C41573 OR2X1_LOC_573/Y OR2X1_LOC_575/a_8_216# 0.39fF
C56548 OR2X1_LOC_573/Y VSS 0.17fF
C49182 VDD OR2X1_LOC_736/Y 0.18fF
C51702 OR2X1_LOC_736/Y OR2X1_LOC_741/a_8_216# 0.03fF
C56782 OR2X1_LOC_736/Y VSS 0.42fF
C20742 VDD OR2X1_LOC_807/A 0.04fF
C28841 OR2X1_LOC_806/a_8_216# OR2X1_LOC_807/A 0.01fF
C31549 OR2X1_LOC_807/A OR2X1_LOC_580/a_8_216# 0.39fF
C33272 OR2X1_LOC_807/A OR2X1_LOC_580/A 0.08fF
C57361 OR2X1_LOC_807/A VSS 0.10fF
C12449 OR2X1_LOC_352/a_8_216# OR2X1_LOC_212/B 0.01fF
C25684 OR2X1_LOC_212/a_8_216# OR2X1_LOC_212/B 0.18fF
C36228 OR2X1_LOC_212/A OR2X1_LOC_212/B 0.07fF
C55423 OR2X1_LOC_357/a_8_216# OR2X1_LOC_212/B 0.41fF
C55464 VDD OR2X1_LOC_212/B 0.08fF
C56430 OR2X1_LOC_212/B VSS 0.36fF
C32971 VDD OR2X1_LOC_212/A 0.08fF
C57139 OR2X1_LOC_212/A VSS -0.28fF
C15430 OR2X1_LOC_853/a_8_216# OR2X1_LOC_857/A 0.01fF
C57858 OR2X1_LOC_857/A VSS 0.09fF
C7019 OR2X1_LOC_205/Y OR2X1_LOC_215/a_8_216# 0.06fF
C10800 OR2X1_LOC_205/Y OR2X1_LOC_217/a_8_216# 0.07fF
C21025 OR2X1_LOC_205/Y OR2X1_LOC_215/A 0.31fF
C54935 VDD OR2X1_LOC_205/Y 0.12fF
C56951 OR2X1_LOC_205/Y VSS 0.30fF
C831 VDD OR2X1_LOC_650/Y 0.39fF
C8966 OR2X1_LOC_650/a_8_216# OR2X1_LOC_650/Y 0.01fF
C35998 OR2X1_LOC_650/Y OR2X1_LOC_654/a_8_216# 0.03fF
C47265 OR2X1_LOC_650/Y OR2X1_LOC_654/a_36_216# 0.02fF
C57582 OR2X1_LOC_650/Y VSS 0.25fF
C10295 VDD OR2X1_LOC_804/A 0.30fF
C35025 OR2X1_LOC_223/A OR2X1_LOC_804/A 0.01fF
C56839 OR2X1_LOC_804/A VSS 0.51fF
C14390 OR2X1_LOC_469/Y OR2X1_LOC_478/a_8_216# 0.06fF
C30420 VDD OR2X1_LOC_469/Y 0.18fF
C50218 OR2X1_LOC_469/Y OR2X1_LOC_738/A 0.01fF
C57272 OR2X1_LOC_469/Y VSS -0.35fF
C8283 OR2X1_LOC_562/Y OR2X1_LOC_570/a_8_216# 0.02fF
C13790 OR2X1_LOC_562/Y OR2X1_LOC_570/a_36_216# 0.03fF
C42986 VDD OR2X1_LOC_562/Y 0.09fF
C56831 OR2X1_LOC_562/Y VSS 0.18fF
C6324 OR2X1_LOC_663/A OR2X1_LOC_404/Y 0.03fF
C14470 OR2X1_LOC_404/Y OR2X1_LOC_573/a_8_216# 0.05fF
C57501 OR2X1_LOC_404/Y VSS -0.73fF
C8000 OR2X1_LOC_774/Y D_GATE_662 0.25fF
C15214 OR2X1_LOC_774/Y VDD 0.11fF
C26805 OR2X1_LOC_774/Y D_GATE_865 0.01fF
C36313 OR2X1_LOC_774/Y OR2X1_LOC_866/B 0.20fF
C54908 OR2X1_LOC_774/Y OR2X1_LOC_865/a_8_216# 0.01fF
C5540 OR2X1_LOC_722/a_8_216# OR2X1_LOC_733/B 0.01fF
C11854 VDD OR2X1_LOC_733/B -0.00fF
C56617 OR2X1_LOC_733/B VSS 0.13fF
C26516 OR2X1_LOC_215/a_8_216# OR2X1_LOC_215/A 0.02fF
C54511 OR2X1_LOC_215/A OR2X1_LOC_215/Y 0.01fF
C56855 OR2X1_LOC_215/A VSS 0.08fF
C34864 OR2X1_LOC_655/a_8_216# OR2X1_LOC_655/A 0.39fF
C47451 OR2X1_LOC_649/a_8_216# OR2X1_LOC_655/A -0.00fF
C55329 VDD OR2X1_LOC_655/A -0.00fF
C57228 OR2X1_LOC_655/A VSS 0.18fF
C32100 VDD OR2X1_LOC_215/Y 0.12fF
C34323 OR2X1_LOC_215/Y OR2X1_LOC_222/A 0.05fF
C56735 OR2X1_LOC_215/Y VSS 0.12fF
C10369 OR2X1_LOC_220/B OR2X1_LOC_742/B 0.03fF
C57097 OR2X1_LOC_220/B VSS 0.18fF
C48688 VDD AND2X1_LOC_738/Y 0.25fF
C56192 AND2X1_LOC_738/Y AND2X1_LOC_740/a_8_24# 0.19fF
C56266 AND2X1_LOC_738/Y VSS 0.10fF
C3353 AND2X1_LOC_480/A AND2X1_LOC_220/Y 0.05fF
C3727 AND2X1_LOC_741/Y AND2X1_LOC_220/Y 0.11fF
C23372 VDD AND2X1_LOC_220/Y 0.29fF
C53955 AND2X1_LOC_478/a_8_24# AND2X1_LOC_220/Y 0.20fF
C56608 AND2X1_LOC_220/Y VSS 0.14fF
C252 OR2X1_LOC_808/A OR2X1_LOC_645/a_8_216# 0.01fF
C18379 OR2X1_LOC_808/A OR2X1_LOC_223/A 0.20fF
C21716 OR2X1_LOC_808/A OR2X1_LOC_794/a_8_216# 0.03fF
C35915 OR2X1_LOC_804/a_8_216# OR2X1_LOC_808/A 0.12fF
C46705 OR2X1_LOC_808/B OR2X1_LOC_808/A 0.05fF
C49692 VDD OR2X1_LOC_808/A 0.27fF
C57485 OR2X1_LOC_808/A VSS -0.64fF
C4669 VDD D_GATE_222 0.04fF
C57099 D_GATE_222 VSS 0.02fF
C10772 OR2X1_LOC_742/B D_GATE_741 0.18fF
C28964 VDD OR2X1_LOC_742/B 0.17fF
C36607 OR2X1_LOC_742/B OR2X1_LOC_551/a_8_216# 0.03fF
C39118 OR2X1_LOC_742/B OR2X1_LOC_741/Y 0.03fF
C47907 OR2X1_LOC_742/B OR2X1_LOC_551/a_36_216# 0.02fF
C53895 OR2X1_LOC_223/A OR2X1_LOC_742/B 0.03fF
C55874 OR2X1_LOC_742/B OR2X1_LOC_742/a_8_216# 0.01fF
C56843 OR2X1_LOC_742/B VSS 0.24fF
C6141 VDD OR2X1_LOC_741/Y 0.06fF
C32904 OR2X1_LOC_741/Y OR2X1_LOC_742/a_8_216# 0.07fF
C56723 OR2X1_LOC_741/Y VSS -0.10fF
C1180 D_GATE_479 OR2X1_LOC_466/a_8_216# 0.01fF
C19767 D_GATE_479 VDD 0.11fF
C57829 D_GATE_479 VSS 0.04fF
C14068 AND2X1_LOC_577/Y AND2X1_LOC_578/a_8_24# 0.03fF
C25083 AND2X1_LOC_577/Y AND2X1_LOC_580/A 0.20fF
C30546 AND2X1_LOC_577/Y AND2X1_LOC_578/a_36_24# 0.01fF
C55626 VDD AND2X1_LOC_577/Y 0.01fF
C57812 AND2X1_LOC_577/Y VSS 0.23fF
C16841 AND2X1_LOC_219/Y AND2X1_LOC_222/a_8_24# 0.01fF
C22716 AND2X1_LOC_219/Y AND2X1_LOC_222/Y 0.02fF
C31653 VDD AND2X1_LOC_219/Y 0.78fF
C32264 AND2X1_LOC_660/A AND2X1_LOC_219/Y 0.07fF
C49307 AND2X1_LOC_649/a_8_24# AND2X1_LOC_219/Y 0.01fF
C56560 AND2X1_LOC_219/Y VSS -1.06fF
C16157 AND2X1_LOC_808/A AND2X1_LOC_212/Y 0.06fF
C27706 AND2X1_LOC_808/A AND2X1_LOC_804/Y 0.24fF
C33196 AND2X1_LOC_808/A AND2X1_LOC_808/a_8_24# 0.01fF
C38196 VDD AND2X1_LOC_808/A 0.36fF
C38203 AND2X1_LOC_738/a_8_24# AND2X1_LOC_808/A 0.20fF
C38692 AND2X1_LOC_808/A AND2X1_LOC_811/B 0.01fF
C41342 AND2X1_LOC_811/Y AND2X1_LOC_808/A 0.05fF
C41598 AND2X1_LOC_808/A AND2X1_LOC_469/a_8_24# 0.01fF
C42936 AND2X1_LOC_808/A AND2X1_LOC_657/Y 0.03fF
C45551 AND2X1_LOC_738/B AND2X1_LOC_808/A 0.03fF
C56936 AND2X1_LOC_808/A VSS 0.29fF
C9980 OR2X1_LOC_659/Y OR2X1_LOC_663/a_8_216# 0.03fF
C21030 OR2X1_LOC_659/Y D_GATE_662 0.74fF
C27405 OR2X1_LOC_663/A OR2X1_LOC_659/Y 0.10fF
C28235 VDD OR2X1_LOC_659/Y -0.00fF
C35478 OR2X1_LOC_659/Y OR2X1_LOC_659/B 0.13fF
C57711 OR2X1_LOC_659/Y VSS -0.00fF
C976 OR2X1_LOC_222/a_8_216# OR2X1_LOC_222/A 0.04fF
C45485 OR2X1_LOC_219/a_8_216# OR2X1_LOC_222/A 0.01fF
C54357 VDD OR2X1_LOC_222/A 0.07fF
C56734 OR2X1_LOC_222/A VSS 0.17fF
C11723 AND2X1_LOC_215/Y VDD 0.19fF
C58091 AND2X1_LOC_215/Y VSS 0.15fF
C3194 OR2X1_LOC_478/Y VDD -0.00fF
C15835 OR2X1_LOC_478/Y OR2X1_LOC_480/a_8_216# 0.39fF
C43122 OR2X1_LOC_478/Y OR2X1_LOC_478/a_8_216# -0.00fF
C57830 OR2X1_LOC_478/Y VSS 0.17fF
C12224 AND2X1_LOC_663/A AND2X1_LOC_804/Y 0.05fF
C19399 AND2X1_LOC_212/Y AND2X1_LOC_804/Y 0.02fF
C32330 AND2X1_LOC_804/Y AND2X1_LOC_222/Y 0.01fF
C36391 AND2X1_LOC_804/Y AND2X1_LOC_808/a_8_24# 0.04fF
C41431 VDD AND2X1_LOC_804/Y 0.21fF
C44696 AND2X1_LOC_811/Y AND2X1_LOC_804/Y 0.59fF
C46270 AND2X1_LOC_733/Y AND2X1_LOC_804/Y 0.01fF
C53161 AND2X1_LOC_804/Y AND2X1_LOC_808/a_36_24# 0.01fF
C56648 AND2X1_LOC_804/Y VSS 0.02fF
C42207 VDD OR2X1_LOC_740/B 0.03fF
C44685 OR2X1_LOC_740/B OR2X1_LOC_739/a_8_216# 0.02fF
C50368 OR2X1_LOC_740/B OR2X1_LOC_739/a_36_216# 0.02fF
C56370 OR2X1_LOC_740/B VSS 0.17fF
C33899 OR2X1_LOC_364/Y OR2X1_LOC_365/a_8_216# 0.39fF
C56340 OR2X1_LOC_364/Y VSS 0.02fF
C2706 OR2X1_LOC_811/A OR2X1_LOC_733/Y 0.17fF
C30392 OR2X1_LOC_733/Y OR2X1_LOC_737/a_8_216# 0.39fF
C47841 OR2X1_LOC_733/a_8_216# OR2X1_LOC_733/Y 0.01fF
C56417 OR2X1_LOC_733/Y VSS 0.17fF
C9625 AND2X1_LOC_570/Y VDD 0.52fF
C14295 AND2X1_LOC_570/Y AND2X1_LOC_657/Y 0.05fF
C27107 AND2X1_LOC_570/Y AND2X1_LOC_807/Y 0.03fF
C34171 AND2X1_LOC_570/Y AND2X1_LOC_577/a_8_24# 0.11fF
C35108 AND2X1_LOC_570/Y AND2X1_LOC_580/A 0.03fF
C35121 AND2X1_LOC_570/Y AND2X1_LOC_579/a_8_24# 0.02fF
C36286 AND2X1_LOC_570/Y AND2X1_LOC_663/A 0.05fF
C38773 AND2X1_LOC_575/a_8_24# AND2X1_LOC_570/Y 0.01fF
C57869 AND2X1_LOC_570/Y VSS -0.24fF
C13556 OR2X1_LOC_808/B OR2X1_LOC_211/a_8_216# 0.35fF
C17923 OR2X1_LOC_808/B OR2X1_LOC_223/A 0.03fF
C46756 OR2X1_LOC_808/B OR2X1_LOC_732/a_8_216# 0.30fF
C48551 OR2X1_LOC_364/A OR2X1_LOC_808/B 0.22fF
C49242 VDD OR2X1_LOC_808/B 2.03fF
C57553 OR2X1_LOC_808/B VSS 0.90fF
C618 AND2X1_LOC_663/A AND2X1_LOC_212/Y 0.10fF
C13738 AND2X1_LOC_663/A AND2X1_LOC_222/Y 0.03fF
C22362 AND2X1_LOC_663/A GATE_579 0.38fF
C22863 VDD AND2X1_LOC_663/A 5.74fF
C29970 AND2X1_LOC_738/B AND2X1_LOC_663/A 0.10fF
C40152 AND2X1_LOC_807/Y AND2X1_LOC_663/A 1.20fF
C42516 AND2X1_LOC_663/a_8_24# AND2X1_LOC_663/A 0.07fF
C42831 AND2X1_LOC_576/Y AND2X1_LOC_663/A 0.10fF
C45101 AND2X1_LOC_866/A AND2X1_LOC_663/A 0.05fF
C48532 AND2X1_LOC_580/A AND2X1_LOC_663/A 0.03fF
C53986 AND2X1_LOC_580/B AND2X1_LOC_663/A 0.03fF
C56681 AND2X1_LOC_663/A VSS 0.56fF
C2405 AND2X1_LOC_363/Y AND2X1_LOC_366/a_8_24# 0.09fF
C8339 AND2X1_LOC_363/a_8_24# AND2X1_LOC_363/Y 0.02fF
C19365 AND2X1_LOC_363/a_36_24# AND2X1_LOC_363/Y 0.02fF
C20344 AND2X1_LOC_363/Y AND2X1_LOC_359/a_8_24# 0.01fF
C24475 VDD AND2X1_LOC_363/Y 0.19fF
C33859 AND2X1_LOC_363/Y AND2X1_LOC_367/a_8_24# 0.01fF
C39356 AND2X1_LOC_363/Y GATE_366 0.01fF
C46867 AND2X1_LOC_363/Y AND2X1_LOC_866/A 0.06fF
C57669 AND2X1_LOC_363/Y VSS -0.22fF
C16051 VDD AND2X1_LOC_576/Y 0.02fF
C20769 AND2X1_LOC_576/Y AND2X1_LOC_657/Y 0.10fF
C33532 AND2X1_LOC_576/Y AND2X1_LOC_807/Y 0.10fF
C41597 AND2X1_LOC_580/A AND2X1_LOC_576/Y 0.07fF
C45321 AND2X1_LOC_575/a_8_24# AND2X1_LOC_576/Y 0.04fF
C57745 AND2X1_LOC_576/Y VSS -1.59fF
C8119 AND2X1_LOC_580/A AND2X1_LOC_569/a_8_24# 0.01fF
C10060 AND2X1_LOC_580/A AND2X1_LOC_580/a_8_24# 0.10fF
C21116 AND2X1_LOC_580/A GATE_579 0.05fF
C21637 VDD AND2X1_LOC_580/A 0.31fF
C26247 AND2X1_LOC_580/A AND2X1_LOC_657/Y 0.03fF
C36043 AND2X1_LOC_578/a_8_24# AND2X1_LOC_580/A 0.01fF
C39027 AND2X1_LOC_580/A AND2X1_LOC_807/Y 1.46fF
C43871 AND2X1_LOC_580/A AND2X1_LOC_866/A 0.03fF
C45473 AND2X1_LOC_580/A AND2X1_LOC_858/a_8_24# 0.04fF
C52819 AND2X1_LOC_580/A AND2X1_LOC_580/B 0.47fF
C57811 AND2X1_LOC_580/A VSS -0.49fF
C636 VDD AND2X1_LOC_657/Y 3.89fF
C1163 AND2X1_LOC_657/Y AND2X1_LOC_811/B 0.42fF
C3884 AND2X1_LOC_811/Y AND2X1_LOC_657/Y 0.34fF
C7912 AND2X1_LOC_738/B AND2X1_LOC_657/Y 0.10fF
C19591 AND2X1_LOC_657/a_8_24# AND2X1_LOC_657/Y 0.01fF
C21972 AND2X1_LOC_657/Y AND2X1_LOC_659/a_8_24# 0.29fF
C34534 AND2X1_LOC_657/Y AND2X1_LOC_212/Y 0.10fF
C47819 AND2X1_LOC_657/Y AND2X1_LOC_222/Y 0.03fF
C48490 AND2X1_LOC_573/a_8_24# AND2X1_LOC_657/Y 0.20fF
C56683 AND2X1_LOC_657/Y VSS 0.91fF
C1599 AND2X1_LOC_566/a_8_24# AND2X1_LOC_212/Y 0.01fF
C19815 AND2X1_LOC_477/a_8_24# AND2X1_LOC_212/Y 0.01fF
C24924 AND2X1_LOC_212/Y AND2X1_LOC_808/a_8_24# 0.03fF
C29447 AND2X1_LOC_212/Y AND2X1_LOC_794/a_8_24# 0.02fF
C30400 AND2X1_LOC_212/Y AND2X1_LOC_811/B 0.01fF
C31080 AND2X1_LOC_212/Y AND2X1_LOC_212/a_8_24# 0.01fF
C33068 AND2X1_LOC_811/Y AND2X1_LOC_212/Y 0.02fF
C33268 AND2X1_LOC_212/Y AND2X1_LOC_469/a_8_24# 0.03fF
C45822 AND2X1_LOC_212/Y AND2X1_LOC_211/a_8_24# 0.03fF
C46818 AND2X1_LOC_864/a_8_24# AND2X1_LOC_212/Y 0.01fF
C52351 AND2X1_LOC_866/A AND2X1_LOC_212/Y 0.83fF
C54784 AND2X1_LOC_568/a_8_24# AND2X1_LOC_212/Y 0.02fF
C56659 AND2X1_LOC_212/Y VSS 0.16fF
C6588 OR2X1_LOC_866/B OR2X1_LOC_865/Y 0.06fF
C42021 OR2X1_LOC_865/Y OR2X1_LOC_866/a_8_216# 0.39fF
C57738 OR2X1_LOC_865/Y VSS 0.18fF
C3350 VDD OR2X1_LOC_659/B 0.18fF
C9666 OR2X1_LOC_659/B OR2X1_LOC_572/a_8_216# 0.40fF
C48191 OR2X1_LOC_659/B OR2X1_LOC_659/a_8_216# 0.06fF
C57396 OR2X1_LOC_659/B VSS 0.47fF
C15599 VDD OR2X1_LOC_738/A 0.05fF
C29297 OR2X1_LOC_469/a_8_216# OR2X1_LOC_738/A 0.02fF
C30097 OR2X1_LOC_731/a_8_216# OR2X1_LOC_738/A 0.03fF
C56669 OR2X1_LOC_738/A VSS 0.57fF
C4805 AND2X1_LOC_580/B AND2X1_LOC_805/a_8_24# 0.01fF
C15561 AND2X1_LOC_580/B AND2X1_LOC_580/a_8_24# 0.03fF
C27124 VDD AND2X1_LOC_580/B 0.61fF
C32064 AND2X1_LOC_580/B AND2X1_LOC_580/a_36_24# 0.01fF
C49556 AND2X1_LOC_580/B AND2X1_LOC_866/A 0.02fF
C51078 AND2X1_LOC_580/B AND2X1_LOC_866/B 0.02fF
C57744 AND2X1_LOC_580/B VSS 0.36fF
C2058 OR2X1_LOC_364/A OR2X1_LOC_645/a_8_216# 0.01fF
C58070 OR2X1_LOC_364/A VSS -1.40fF
C9968 OR2X1_LOC_866/B D_GATE_662 0.14fF
C17177 OR2X1_LOC_866/B VDD 0.08fF
C17664 OR2X1_LOC_866/B OR2X1_LOC_866/a_8_216# 0.06fF
C28711 OR2X1_LOC_866/B D_GATE_865 0.02fF
C57862 OR2X1_LOC_866/B VSS 0.38fF
C14825 OR2X1_LOC_807/Y OR2X1_LOC_811/A 0.04fF
C48036 VDD OR2X1_LOC_807/Y 0.05fF
C50634 OR2X1_LOC_807/Y OR2X1_LOC_805/a_8_216# 0.05fF
C57740 OR2X1_LOC_807/Y VSS 0.27fF
C3718 AND2X1_LOC_804/a_8_24# AND2X1_LOC_222/Y 0.01fF
C4371 AND2X1_LOC_807/Y AND2X1_LOC_222/Y 0.16fF
C6038 AND2X1_LOC_357/a_8_24# AND2X1_LOC_222/Y 0.01fF
C8242 AND2X1_LOC_737/a_8_24# AND2X1_LOC_222/Y 0.01fF
C9204 AND2X1_LOC_866/A AND2X1_LOC_222/Y 0.03fF
C15437 AND2X1_LOC_811/a_8_24# AND2X1_LOC_222/Y 0.01fF
C18424 AND2X1_LOC_723/a_8_24# AND2X1_LOC_222/Y 0.01fF
C23481 AND2X1_LOC_741/Y AND2X1_LOC_222/Y 0.01fF
C29840 AND2X1_LOC_733/a_8_24# AND2X1_LOC_222/Y 0.01fF
C34463 AND2X1_LOC_741/a_8_24# AND2X1_LOC_222/Y 0.01fF
C37782 AND2X1_LOC_182/a_8_24# AND2X1_LOC_222/Y 0.01fF
C39329 AND2X1_LOC_222/Y AND2X1_LOC_223/a_8_24# 0.04fF
C39702 AND2X1_LOC_480/a_8_24# AND2X1_LOC_222/Y 0.01fF
C42544 AND2X1_LOC_722/a_8_24# AND2X1_LOC_222/Y 0.01fF
C42977 VDD AND2X1_LOC_222/Y 0.57fF
C45323 GATE_479 AND2X1_LOC_222/Y 0.01fF
C46188 AND2X1_LOC_811/Y AND2X1_LOC_222/Y 0.01fF
C47845 AND2X1_LOC_733/Y AND2X1_LOC_222/Y 0.01fF
C56500 AND2X1_LOC_222/Y VSS -0.64fF
C14800 OR2X1_LOC_577/a_8_216# D_GATE_366 0.01fF
C34059 VDD D_GATE_366 0.10fF
C38671 OR2X1_LOC_577/Y D_GATE_366 0.02fF
C56257 D_GATE_366 VSS 0.02fF
C3767 OR2X1_LOC_580/A OR2X1_LOC_366/a_8_216# 0.03fF
C8169 OR2X1_LOC_366/A OR2X1_LOC_580/A 0.04fF
C8690 VDD OR2X1_LOC_580/A 0.12fF
C26456 OR2X1_LOC_858/a_8_216# OR2X1_LOC_580/A 0.03fF
C31578 OR2X1_LOC_811/A OR2X1_LOC_580/A 0.10fF
C47784 OR2X1_LOC_363/a_8_216# OR2X1_LOC_580/A 0.04fF
C49984 OR2X1_LOC_359/a_8_216# OR2X1_LOC_580/A 0.04fF
C56350 OR2X1_LOC_580/A VSS -0.80fF
C4590 OR2X1_LOC_660/a_8_216# OR2X1_LOC_660/B 0.05fF
C57522 OR2X1_LOC_660/B VSS 0.21fF
C17512 AND2X1_LOC_733/Y AND2X1_LOC_804/a_8_24# 0.03fF
C22044 AND2X1_LOC_733/Y AND2X1_LOC_737/a_8_24# -0.00fF
C57825 AND2X1_LOC_733/Y VSS -0.27fF
C4047 AND2X1_LOC_739/a_8_24# AND2X1_LOC_742/A 0.20fF
C9078 VDD AND2X1_LOC_742/A 0.21fF
C51190 AND2X1_LOC_742/a_8_24# AND2X1_LOC_742/A 0.03fF
C56265 AND2X1_LOC_742/A VSS 0.16fF
C248 GATE_479 GATE_222 0.03fF
C56499 GATE_222 VSS 0.04fF
C34362 GATE_479 AND2X1_LOC_480/A 0.24fF
C34790 AND2X1_LOC_741/Y GATE_479 0.15fF
C50950 GATE_479 AND2X1_LOC_223/a_8_24# 0.20fF
C51308 AND2X1_LOC_480/a_8_24# GATE_479 0.01fF
C54496 VDD GATE_479 0.22fF
C57147 GATE_479 VSS 0.03fF
C2812 AND2X1_LOC_663/B AND2X1_LOC_217/a_8_24# 0.13fF
C6858 GATE_366 AND2X1_LOC_663/B 0.03fF
C14216 AND2X1_LOC_866/A AND2X1_LOC_663/B 0.02fF
C28196 AND2X1_LOC_660/a_8_24# AND2X1_LOC_663/B 0.08fF
C36352 AND2X1_LOC_663/B AND2X1_LOC_580/a_8_24# 0.01fF
C39182 AND2X1_LOC_660/a_36_24# AND2X1_LOC_663/B 0.01fF
C47641 AND2X1_LOC_663/B GATE_579 0.01fF
C48142 VDD AND2X1_LOC_663/B 1.66fF
C48736 AND2X1_LOC_663/B AND2X1_LOC_660/A 0.07fF
C57114 AND2X1_LOC_663/B VSS -3.54fF
C20042 OR2X1_LOC_221/A OR2X1_LOC_221/a_8_216# 0.18fF
C30955 VDD OR2X1_LOC_221/A 0.06fF
C57259 OR2X1_LOC_221/A VSS 0.16fF
C56439 OR2X1_LOC_570/Y VSS 0.19fF
C2759 OR2X1_LOC_571/a_8_216# OR2X1_LOC_579/A 0.03fF
C8301 OR2X1_LOC_571/a_36_216# OR2X1_LOC_579/A 0.01fF
C13673 OR2X1_LOC_576/a_8_216# OR2X1_LOC_579/A 0.01fF
C43905 VDD OR2X1_LOC_579/A 0.18fF
C56491 OR2X1_LOC_579/A VSS 0.36fF
C34438 OR2X1_LOC_363/a_8_216# OR2X1_LOC_366/A -0.00fF
C46822 OR2X1_LOC_366/A OR2X1_LOC_366/a_8_216# 0.39fF
C51692 VDD OR2X1_LOC_366/A -0.00fF
C56437 OR2X1_LOC_366/A VSS 0.18fF
C9277 AND2X1_LOC_741/Y AND2X1_LOC_221/a_8_24# 0.14fF
C12521 AND2X1_LOC_741/Y AND2X1_LOC_480/A 0.10fF
C18455 AND2X1_LOC_741/Y AND2X1_LOC_742/a_8_24# 0.11fF
C20309 AND2X1_LOC_741/Y AND2X1_LOC_221/a_36_24# 0.01fF
C29286 AND2X1_LOC_741/Y AND2X1_LOC_480/a_8_24# 0.21fF
C32405 AND2X1_LOC_741/Y VDD 0.29fF
C58085 AND2X1_LOC_741/Y VSS -0.08fF
C13524 VDD AND2X1_LOC_807/Y 1.36fF
C14040 AND2X1_LOC_807/Y AND2X1_LOC_811/B 0.04fF
C16667 AND2X1_LOC_807/Y AND2X1_LOC_811/Y 0.03fF
C17730 AND2X1_LOC_861/a_8_24# AND2X1_LOC_807/Y 0.04fF
C31768 AND2X1_LOC_865/a_8_24# AND2X1_LOC_807/Y 0.02fF
C37241 AND2X1_LOC_866/B AND2X1_LOC_807/Y 0.03fF
C41998 AND2X1_LOC_807/Y AND2X1_LOC_811/a_8_24# 0.05fF
C45951 AND2X1_LOC_862/a_36_24# AND2X1_LOC_807/Y 0.05fF
C57089 AND2X1_LOC_807/Y VSS 0.60fF
C14160 AND2X1_LOC_660/A AND2X1_LOC_649/a_8_24# 0.05fF
C32850 AND2X1_LOC_660/a_8_24# AND2X1_LOC_660/A 0.02fF
C45954 AND2X1_LOC_218/a_8_24# AND2X1_LOC_660/A 0.02fF
C52837 VDD AND2X1_LOC_660/A 0.26fF
C56918 AND2X1_LOC_660/A VSS 0.23fF
C27690 OR2X1_LOC_577/Y OR2X1_LOC_367/a_8_216# 0.01fF
C56400 OR2X1_LOC_577/Y VSS 0.25fF
C10041 AND2X1_LOC_352/a_8_24# AND2X1_LOC_364/Y 0.01fF
C22035 AND2X1_LOC_364/Y AND2X1_LOC_863/a_8_24# 0.01fF
C32037 VDD AND2X1_LOC_364/Y 0.29fF
C57723 AND2X1_LOC_364/Y VSS -0.85fF
C22818 VDD OR2X1_LOC_580/B 0.70fF
C33575 OR2X1_LOC_580/a_8_216# OR2X1_LOC_580/B 0.06fF
C50333 D_GATE_579 OR2X1_LOC_580/B 0.02fF
C56399 OR2X1_LOC_580/B VSS -2.43fF
C19369 AND2X1_LOC_866/B GATE_579 0.03fF
C19857 VDD AND2X1_LOC_866/B 0.39fF
C42088 AND2X1_LOC_866/A AND2X1_LOC_866/B 0.07fF
C45140 AND2X1_LOC_866/B GATE_662 0.03fF
C57129 AND2X1_LOC_866/B VSS 0.11fF
C3251 AND2X1_LOC_738/B VDD 1.29fF
C34389 AND2X1_LOC_738/B AND2X1_LOC_803/a_8_24# 0.03fF
C58042 AND2X1_LOC_738/B VSS 0.54fF
C14247 VDD AND2X1_LOC_358/Y 0.46fF
C57795 AND2X1_LOC_358/Y VSS 0.15fF
C8879 AND2X1_LOC_480/A AND2X1_LOC_221/a_8_24# 0.20fF
C28893 AND2X1_LOC_480/a_8_24# AND2X1_LOC_480/A 0.01fF
C32000 VDD AND2X1_LOC_480/A 0.21fF
C56676 AND2X1_LOC_480/A VSS 0.19fF
C2141 AND2X1_LOC_363/a_8_24# AND2X1_LOC_866/A 0.17fF
C6722 AND2X1_LOC_866/A AND2X1_LOC_580/a_8_24# 0.02fF
C17785 AND2X1_LOC_866/A GATE_579 0.01fF
C18320 VDD AND2X1_LOC_866/A 0.62fF
C21049 AND2X1_LOC_866/A AND2X1_LOC_866/a_8_24# -0.00fF
C33210 GATE_366 AND2X1_LOC_866/A 0.07fF
C37902 AND2X1_LOC_866/A AND2X1_LOC_663/a_8_24# 0.04fF
C43522 AND2X1_LOC_866/A GATE_662 0.03fF
C57174 AND2X1_LOC_866/A VSS 0.30fF
C2670 OR2X1_LOC_223/A D_GATE_741 0.01fF
C7292 OR2X1_LOC_804/a_8_216# OR2X1_LOC_223/A 0.01fF
C16303 OR2X1_LOC_479/a_8_216# OR2X1_LOC_223/A 0.01fF
C18487 OR2X1_LOC_223/A OR2X1_LOC_223/a_8_216# 0.18fF
C18520 OR2X1_LOC_223/A OR2X1_LOC_795/a_8_216# 0.01fF
C20915 VDD OR2X1_LOC_223/A 0.41fF
C47787 OR2X1_LOC_223/A OR2X1_LOC_742/a_8_216# 0.01fF
C57140 OR2X1_LOC_223/A VSS -0.45fF
C28343 OR2X1_LOC_662/a_8_216# OR2X1_LOC_663/A 0.01fF
C51367 VDD OR2X1_LOC_663/A 0.11fF
C57771 OR2X1_LOC_663/A VSS -0.17fF
C10954 VDD GATE_366 0.17fF
C57610 GATE_366 VSS 0.14fF
C57092 GATE_865 VSS 0.02fF
C13430 AND2X1_LOC_811/Y AND2X1_LOC_812/a_8_24# 0.06fF
C27715 AND2X1_LOC_811/a_8_24# AND2X1_LOC_811/Y 0.10fF
C50379 AND2X1_LOC_811/Y AND2X1_LOC_808/a_8_24# 0.25fF
C55361 VDD AND2X1_LOC_811/Y 0.24fF
C55863 AND2X1_LOC_811/Y AND2X1_LOC_811/B 0.29fF
C57027 AND2X1_LOC_811/Y VSS 0.29fF
C58084 GATE_741 VSS 0.12fF
C23522 VDD D_GATE_579 0.06fF
C56886 D_GATE_579 VSS 0.09fF
C51796 OR2X1_LOC_812/A OR2X1_LOC_812/a_8_216# 0.39fF
C57739 OR2X1_LOC_812/A VSS 0.18fF
C7575 VDD D_GATE_865 0.06fF
C57737 D_GATE_865 VSS 0.08fF
C15255 AND2X1_LOC_663/a_8_24# GATE_579 0.20fF
C20839 GATE_662 GATE_579 0.02fF
C29300 AND2X1_LOC_805/a_8_24# GATE_579 0.01fF
C51707 VDD GATE_579 0.21fF
C56296 GATE_579 VSS 0.09fF
C21351 VDD GATE_662 0.07fF
C57068 GATE_662 VSS 0.24fF
C24574 OR2X1_LOC_864/a_8_216# D_GATE_662 0.14fF
C44818 VDD D_GATE_662 0.24fF
C57710 D_GATE_662 VSS 0.21fF
C25055 AND2X1_LOC_811/a_8_24# AND2X1_LOC_811/B 0.04fF
C36026 AND2X1_LOC_811/a_36_24# AND2X1_LOC_811/B 0.01fF
C52654 VDD AND2X1_LOC_811/B 0.21fF
C56014 AND2X1_LOC_811/B AND2X1_LOC_469/a_8_24# 0.20fF
C56647 AND2X1_LOC_811/B VSS 0.23fF
C56722 D_GATE_741 VSS 0.12fF
C845 OR2X1_LOC_807/a_8_216# OR2X1_LOC_811/A 0.14fF
C14184 OR2X1_LOC_811/A OR2X1_LOC_366/a_8_216# 0.11fF
C19002 VDD OR2X1_LOC_811/A 0.64fF
C21667 OR2X1_LOC_805/a_8_216# OR2X1_LOC_811/A 0.06fF
C26886 OR2X1_LOC_811/A OR2X1_LOC_736/a_8_216# 0.02fF
C30935 OR2X1_LOC_811/A OR2X1_LOC_733/a_8_216# 0.04fF
C57254 OR2X1_LOC_811/A VSS -1.96fF
C1713 OR2X1_LOC_733/a_8_216# OR2X1_LOC_722/a_8_216# 0.47fF
C1840 OR2X1_LOC_211/a_8_216# OR2X1_LOC_566/a_8_216# 0.47fF
C2041 AND2X1_LOC_365/a_8_24# AND2X1_LOC_661/a_8_24# 0.23fF
C3265 VDD OR2X1_LOC_573/a_8_216# 0.21fF
C5211 OR2X1_LOC_860/a_8_216# OR2X1_LOC_576/a_8_216# 0.47fF
C8027 VDD OR2X1_LOC_217/a_8_216# 0.21fF
C9736 VDD OR2X1_LOC_469/a_8_216# 0.21fF
C18569 AND2X1_LOC_861/a_8_24# AND2X1_LOC_865/a_8_24# 0.23fF
C22857 VDD OR2X1_LOC_742/a_8_216# 0.21fF
C31196 VDD OR2X1_LOC_654/a_8_216# 0.21fF
C35329 OR2X1_LOC_244/a_8_216# OR2X1_LOC_141/a_8_216# 0.47fF
C35954 OR2X1_LOC_853/a_8_216# OR2X1_LOC_857/a_8_216# 0.47fF
C36925 AND2X1_LOC_650/a_8_24# AND2X1_LOC_857/a_8_24# 0.23fF
C37485 VDD AND2X1_LOC_206/a_8_24# -0.00fF
C38670 OR2X1_LOC_578/a_8_216# OR2X1_LOC_367/a_8_216# 0.47fF
C39519 AND2X1_LOC_566/a_8_24# AND2X1_LOC_211/a_8_24# 0.23fF
C42033 OR2X1_LOC_806/a_8_216# OR2X1_LOC_807/a_8_216# 0.47fF
C49721 VDD OR2X1_LOC_732/a_8_216# 0.21fF
C51340 VDD AND2X1_LOC_468/a_8_24# -0.00fF
C54896 VDD OR2X1_LOC_222/a_8_216# 0.21fF
C55937 AND2X1_LOC_562/a_8_24# VDD -0.00fF
C56135 OR2X1_LOC_811/a_8_216# OR2X1_LOC_805/a_8_216# 0.47fF
C56250 AND2X1_LOC_570/a_8_24# VSS 0.10fF
C56559 AND2X1_LOC_222/a_8_24# VSS 0.10fF
C56686 AND2X1_LOC_648/a_8_24# VSS 0.10fF
C57176 AND2X1_LOC_853/a_8_24# VSS 0.10fF
C57479 AND2X1_LOC_358/a_8_24# VSS 0.10fF
C57538 AND2X1_LOC_357/a_8_24# VSS 0.10fF
C57742 AND2X1_LOC_568/a_8_24# VSS 0.10fF
C57794 AND2X1_LOC_364/a_8_24# VSS 0.10fF
C57814 AND2X1_LOC_556/a_8_24# VSS 0.10fF
C57868 AND2X1_LOC_577/a_8_24# VSS 0.10fF
C57972 AND2X1_LOC_723/a_8_24# VSS 0.10fF
C31608 AND2X1_LOC_810/A AND2X1_LOC_436/Y 0.01fF
C49398 AND2X1_LOC_810/A AND2X1_LOC_863/Y 0.14fF
C32051 AND2X1_LOC_810/A AND2X1_LOC_655/A 0.05fF
C14388 AND2X1_LOC_810/A AND2X1_LOC_212/B 0.15fF
C21484 AND2X1_LOC_810/A AND2X1_LOC_212/Y 0.05fF
C13496 OR2X1_LOC_865/A OR2X1_LOC_774/Y 0.06fF
C7218 OR2X1_LOC_865/B OR2X1_LOC_774/Y 0.06fF
C4676 OR2X1_LOC_774/Y OR2X1_LOC_865/Y 0.01fF
C15728 OR2X1_LOC_774/Y OR2X1_LOC_866/a_8_216# 0.01fF
C51154 OR2X1_LOC_774/Y OR2X1_LOC_864/a_8_216# 0.03fF
C43315 OR2X1_LOC_217/Y OR2X1_LOC_510/Y 0.02fF
C35820 OR2X1_LOC_510/Y OR2X1_LOC_217/A 0.14fF
C43777 OR2X1_LOC_510/Y OR2X1_LOC_217/a_8_216# 0.01fF
C22770 AND2X1_LOC_574/A AND2X1_LOC_657/a_8_24# 0.08fF
C30561 AND2X1_LOC_574/A AND2X1_LOC_663/A 0.50fF
C4857 OR2X1_LOC_863/A OR2X1_LOC_35/Y 0.01fF
C16956 OR2X1_LOC_864/A OR2X1_LOC_35/Y 0.03fF
C332 OR2X1_LOC_863/a_8_216# OR2X1_LOC_35/Y 0.01fF
C7432 OR2X1_LOC_853/a_36_216# OR2X1_LOC_35/Y 0.03fF
C33519 OR2X1_LOC_857/a_8_216# OR2X1_LOC_35/Y 0.01fF
C36305 AND2X1_LOC_35/Y AND2X1_LOC_219/A 0.07fF
C53669 AND2X1_LOC_573/A AND2X1_LOC_361/A 0.02fF
C32577 AND2X1_LOC_858/B AND2X1_LOC_573/A 0.10fF
C33436 AND2X1_LOC_367/A AND2X1_LOC_573/A 0.10fF
C42858 AND2X1_LOC_571/Y AND2X1_LOC_573/A 0.01fF
C34076 AND2X1_LOC_573/A AND2X1_LOC_562/Y 0.01fF
C54678 AND2X1_LOC_571/A AND2X1_LOC_573/A 0.01fF
C42169 AND2X1_LOC_573/A AND2X1_LOC_657/A 0.16fF
C3829 AND2X1_LOC_807/Y AND2X1_LOC_573/A 0.03fF
C6308 AND2X1_LOC_576/Y AND2X1_LOC_573/A 0.02fF
C20313 AND2X1_LOC_141/a_8_24# AND2X1_LOC_573/A 0.03fF
C38198 AND2X1_LOC_663/B AND2X1_LOC_573/A 0.10fF
C39603 AND2X1_LOC_573/A AND2X1_LOC_563/Y 0.19fF
C48424 AND2X1_LOC_571/a_8_24# AND2X1_LOC_573/A 0.01fF
C53369 AND2X1_LOC_573/A AND2X1_LOC_217/a_8_24# 0.01fF
C56069 AND2X1_LOC_570/Y AND2X1_LOC_573/A 0.02fF
C45895 OR2X1_LOC_404/Y OR2X1_LOC_244/Y 0.43fF
C24578 OR2X1_LOC_404/Y OR2X1_LOC_576/A 0.03fF
C26409 OR2X1_LOC_864/A OR2X1_LOC_404/Y 0.03fF
C22175 OR2X1_LOC_404/Y OR2X1_LOC_659/A 0.02fF
C14542 OR2X1_LOC_404/Y OR2X1_LOC_659/B 0.02fF

.ends

* wrdata outputs.out V("GATE_222") V("GATE_366") V("GATE_479") V("GATE_579") V("GATE_662") V("GATE_741") V("GATE_811") V("GATE_865") V("D_GATE_222") V("D_GATE_366") V("D_GATE_479") V("D_GATE_579") V("D_GATE_662") V("D_GATE_741") V("D_GATE_811") V("D_GATE_865") 

