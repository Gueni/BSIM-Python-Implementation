* SPICE3 file created from PAND2X1_NOCTRL_UP.ext - technology: scmos

.subckt PAND2X1 VDD GND B A Y
X0 Y O VDD VDD PMOS_MAGIC ad=1.95p pd=8.8u as=3.47p ps=16.6u w=3.9u l=0.2u
**devattr s=S d=D
X1 O GND GND GND NMOS_MAGIC ad=0.9p pd=4.2u as=2.61p ps=14u w=1.5u l=0.2u
**devattr s=S d=D
X2 Y O GND GND NMOS_MAGIC ad=1.1p pd=5.4u as=0p ps=0u w=2.2u l=0.2u
**devattr s=S d=D
X3 O GND a_48_324# VDD PMOS_MAGIC ad=0.96p pd=4.4u as=1.52p ps=7.8u w=1.6u l=0.2u
**devattr s=S d=D
X4 a_8_28# B a_36_28# GND NMOS_MAGIC ad=0.99p pd=6u as=0.12p ps=1.4u w=0.4u l=0.2u
**devattr s=S d=D
X5 a_8_28# A a_88_28# GND NMOS_MAGIC ad=0p pd=0u as=0.12p ps=1.4u w=0.4u l=0.2u
**devattr s=S d=D
X6 a_88_28# B GND GND NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X7 a_48_324# A VDD VDD PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=1.2u l=0.2u
**devattr s=S d=D
X8 a_36_28# A GND GND NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X9 a_48_324# B VDD VDD PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=1.2u l=0.2u
**devattr s=S d=D
X10 O VDD VDD VDD PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=1.6u l=0.2u
**devattr s=S d=D
X11 O VDD a_8_28# GND NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=1.5u l=0.2u
**devattr s=S d=D
C0 A a_8_28# 0.01fF
C1 O a_48_324# 0.22fF
C2 O a_8_28# 0.15fF
C3 VDD B 0.39fF
C4 VDD A 0.37fF
C5 a_8_28# a_36_28# 0.00fF
C6 B A 0.83fF
C7 VDD Y 0.54fF
C8 a_8_28# a_88_28# 0.00fF
C9 VDD O 0.61fF
C10 B O 0.03fF
C11 VDD a_48_324# 0.40fF
C12 A O 0.07fF
C13 B a_48_324# 0.01fF
C14 A a_48_324# 0.01fF
C15 B a_8_28# 0.01fF
C16 Y O 0.05fF
.ends

