magic
tech scmos
magscale 1 2
timestamp 1612251229
<< metal1 >>
rect 4984 7537 5075 7543
rect 920 7516 924 7524
rect 1597 7517 1683 7523
rect 2045 7517 2060 7523
rect 2509 7517 2524 7523
rect 2788 7517 2796 7523
rect 2940 7523 2948 7524
rect 2940 7517 3027 7523
rect 3924 7516 3932 7524
rect 4285 7517 4300 7523
rect 4356 7517 4371 7523
rect 4748 7517 4835 7523
rect 5069 7517 5075 7537
rect 5860 7537 5891 7543
rect 6332 7537 6355 7543
rect 5885 7523 5891 7537
rect 5885 7517 5955 7523
rect 6349 7523 6355 7537
rect 6349 7517 6408 7523
rect 6612 7517 6627 7523
rect 6804 7517 6852 7523
rect 7005 7517 7052 7523
rect 7076 7517 7091 7523
rect 7453 7517 7468 7523
rect 9197 7517 9244 7523
rect 76 7504 84 7514
rect 316 7484 324 7490
rect 908 7484 916 7490
rect 4604 7484 4612 7490
rect 461 7477 524 7483
rect 685 7477 748 7483
rect 932 7477 980 7483
rect 1368 7477 1459 7483
rect 2068 7477 2131 7483
rect 2292 7477 2360 7483
rect 2532 7477 2579 7483
rect 2740 7477 2803 7483
rect 3389 7477 3452 7483
rect 3613 7477 3708 7483
rect 4524 7477 4588 7483
rect 5437 7477 5523 7483
rect 6412 7483 6420 7490
rect 6388 7477 6420 7483
rect 7548 7483 7556 7490
rect 8204 7484 8212 7490
rect 7540 7477 7556 7483
rect 7901 7477 7987 7483
rect 1844 7457 1907 7463
rect 234 7437 300 7443
rect 3176 7436 3180 7444
rect 3236 7437 3251 7443
rect 3476 7436 3478 7444
rect 4077 7437 4092 7443
rect 5658 7436 5660 7444
rect 6557 7437 6572 7443
rect 6776 7436 6780 7444
rect 7229 7437 7244 7443
rect 7693 7437 7708 7443
rect 8124 7437 8140 7443
rect 8568 7436 8572 7444
rect 9044 7437 9059 7443
rect 9421 7437 9436 7443
rect 9852 7437 9868 7443
rect 676 7377 739 7383
rect 2244 7377 2296 7383
rect 3124 7377 3187 7383
rect 4468 7377 4516 7383
rect 5140 7377 5190 7383
rect 5588 7377 5651 7383
rect 7188 7377 7235 7383
rect 7860 7377 7907 7383
rect 8068 7377 8132 7383
rect 8308 7377 8371 7383
rect 10061 7377 10268 7383
rect 1348 7357 1411 7363
rect 4020 7357 4072 7363
rect 6728 7357 6796 7363
rect 1548 7337 1580 7343
rect 876 7330 884 7336
rect 1548 7330 1556 7337
rect 2020 7337 2083 7343
rect 3981 7337 3996 7343
rect 4964 7337 4979 7343
rect 6324 7337 6356 7343
rect 2748 7330 2756 7336
rect 4444 7330 4452 7336
rect 6348 7330 6356 7337
rect 6797 7343 6803 7356
rect 6797 7337 6819 7343
rect 7468 7330 7476 7336
rect 8044 7330 8052 7336
rect 5117 7317 5164 7323
rect 205 7297 268 7303
rect 2020 7297 2070 7303
rect 2445 7297 2460 7303
rect 2740 7296 2744 7304
rect 4884 7297 4924 7303
rect 5341 7297 5356 7303
rect 5565 7297 5580 7303
rect 5860 7297 5891 7303
rect 7821 7297 7836 7303
rect 8733 7297 8819 7303
rect 9261 7283 9267 7303
rect 9194 7277 9267 7283
rect 2221 7237 2236 7243
rect 2893 7237 2908 7243
rect 3396 7236 3398 7244
rect 5380 7237 5427 7243
rect 6957 7237 6972 7243
rect 7165 7237 7180 7243
rect 8957 7237 8972 7243
rect 9405 7237 9420 7243
rect 7028 7176 7030 7184
rect 221 7117 268 7123
rect 669 7117 684 7123
rect 1140 7117 1203 7123
rect 2013 7117 2035 7123
rect 908 7097 940 7103
rect 429 7077 520 7083
rect 1101 7077 1148 7083
rect 1581 7077 1652 7083
rect 2029 7083 2035 7117
rect 2924 7123 2932 7124
rect 2924 7117 3011 7123
rect 3373 7117 3459 7123
rect 4461 7117 4476 7123
rect 5357 7117 5443 7123
rect 9005 7117 9052 7123
rect 2029 7077 2099 7083
rect 2237 7077 2252 7083
rect 2780 7083 2788 7090
rect 2477 7077 2563 7083
rect 2700 7077 2788 7083
rect 3188 7077 3235 7083
rect 5812 7077 5880 7083
rect 6940 7083 6948 7090
rect 8172 7084 8180 7090
rect 6940 7077 6956 7083
rect 7476 7077 7491 7083
rect 7629 7077 7718 7083
rect 7876 7077 7955 7083
rect 9212 7077 9299 7083
rect 9869 7077 9940 7083
rect 3834 7057 3868 7063
rect 68 7037 83 7043
rect 1352 7036 1356 7044
rect 5594 7036 5596 7044
rect 6268 7037 6284 7043
rect 6728 7037 6780 7043
rect 8317 7037 8332 7043
rect 8552 7036 8556 7044
rect 8781 7037 8796 7043
rect 9684 7037 9731 7043
rect 276 6977 291 6983
rect 2010 6977 2028 6983
rect 2221 6977 2252 6983
rect 2468 6977 2515 6983
rect 3348 6977 3398 6983
rect 4452 6977 4484 6983
rect 6020 6977 6083 6983
rect 6484 6977 6547 6983
rect 7396 6977 7427 6983
rect 9140 6977 9203 6983
rect 10029 6977 10060 6983
rect 676 6957 739 6963
rect 3796 6957 3843 6963
rect 7604 6957 7640 6963
rect 8708 6957 8742 6963
rect 9581 6957 9644 6963
rect 429 6937 518 6943
rect 876 6930 884 6936
rect 1548 6937 1612 6943
rect 972 6930 980 6936
rect 1548 6930 1556 6937
rect 6308 6937 6324 6943
rect 2652 6930 2660 6936
rect 6220 6930 6228 6936
rect 6316 6930 6324 6937
rect 7565 6937 7580 6943
rect 8012 6930 8020 6936
rect 8669 6937 8684 6943
rect 8900 6937 8979 6943
rect 9341 6937 9372 6943
rect 8108 6930 8116 6936
rect 1773 6917 1860 6923
rect 2877 6917 2940 6923
rect 1852 6906 1860 6917
rect 7133 6917 7220 6923
rect 7212 6906 7220 6917
rect 221 6897 268 6903
rect 2664 6897 2684 6903
rect 3549 6897 3635 6903
rect 4861 6897 4876 6903
rect 5325 6897 5411 6903
rect 5629 6883 5635 6903
rect 6740 6897 6772 6903
rect 7364 6897 7404 6903
rect 7789 6897 7876 6903
rect 8252 6897 8323 6903
rect 8252 6896 8260 6897
rect 9814 6897 9891 6903
rect 10068 6897 10099 6903
rect 5562 6877 5635 6883
rect 4708 6837 4723 6843
rect 8472 6836 8476 6844
rect 8516 6837 8531 6843
rect 6316 6777 6364 6783
rect 10045 6777 10060 6783
rect 10084 6777 10115 6783
rect 669 6717 755 6723
rect 1821 6717 1852 6723
rect 4493 6717 4508 6723
rect 4772 6717 4803 6723
rect 6077 6717 6092 6723
rect 6524 6723 6532 6724
rect 6310 6717 6387 6723
rect 6524 6717 6611 6723
rect 7044 6717 7059 6723
rect 9814 6717 9868 6723
rect 1132 6704 1140 6714
rect 316 6683 324 6690
rect 4588 6684 4596 6690
rect 308 6677 324 6683
rect 1368 6677 1459 6683
rect 2084 6677 2131 6683
rect 2269 6677 2284 6683
rect 2964 6677 3027 6683
rect 3162 6677 3251 6683
rect 3389 6677 3452 6683
rect 3820 6677 3907 6683
rect 4733 6677 4808 6683
rect 5860 6677 5928 6683
rect 6340 6677 6387 6683
rect 6836 6677 6851 6683
rect 7924 6677 7939 6683
rect 8100 6677 8132 6683
rect 8292 6677 8355 6683
rect 9162 6677 9196 6683
rect 9900 6683 9908 6690
rect 9844 6677 9908 6683
rect 7645 6657 7676 6663
rect 461 6637 476 6643
rect 908 6637 924 6643
rect 1652 6637 1670 6643
rect 2058 6636 2060 6644
rect 3613 6637 3628 6643
rect 4068 6637 4136 6643
rect 5405 6637 5420 6643
rect 5444 6637 5491 6643
rect 6760 6636 6764 6644
rect 6989 6637 7020 6643
rect 7197 6637 7212 6643
rect 7434 6636 7436 6644
rect 8076 6637 8092 6643
rect 8717 6637 8732 6643
rect 9396 6637 9432 6643
rect 10045 6637 10060 6643
rect 676 6577 739 6583
rect 1124 6577 1171 6583
rect 1994 6577 2060 6583
rect 2900 6577 2963 6583
rect 6712 6577 6748 6583
rect 7188 6577 7235 6583
rect 7844 6577 7891 6583
rect 8068 6577 8116 6583
rect 8932 6577 8995 6583
rect 452 6557 504 6563
rect 5124 6557 5174 6563
rect 6948 6557 6998 6563
rect 68 6537 83 6543
rect 413 6537 428 6543
rect 1533 6537 1548 6543
rect 2052 6537 2083 6543
rect 5085 6537 5100 6543
rect 5773 6537 5788 6543
rect 6276 6537 6340 6543
rect 876 6530 884 6536
rect 6332 6530 6340 6537
rect 6909 6537 6924 6543
rect 8276 6537 8344 6543
rect 8488 6537 8563 6543
rect 8740 6537 8772 6543
rect 9204 6537 9219 6543
rect 3101 6497 3116 6503
rect 3325 6497 3411 6503
rect 3757 6497 3772 6503
rect 4861 6497 4892 6503
rect 5549 6497 5564 6503
rect 6084 6497 6099 6503
rect 7149 6497 7164 6503
rect 7821 6497 7868 6503
rect 8029 6497 8044 6503
rect 6013 6477 6092 6483
rect 9213 6483 9219 6503
rect 9581 6497 9612 6503
rect 10052 6497 10115 6503
rect 9156 6477 9219 6483
rect 2221 6437 2236 6443
rect 8701 6437 8732 6443
rect 9357 6437 9388 6443
rect 9428 6436 9432 6444
rect 9146 6376 9148 6384
rect 4500 6337 4548 6343
rect 5165 6337 5212 6343
rect 7418 6337 7491 6343
rect 1604 6317 1651 6323
rect 1789 6317 1875 6323
rect 2712 6317 2764 6323
rect 2948 6317 3011 6323
rect 4269 6317 4316 6323
rect 4477 6317 4492 6323
rect 4980 6317 5012 6323
rect 7181 6317 7267 6323
rect 7485 6317 7491 6337
rect 7837 6317 7852 6323
rect 8045 6317 8060 6323
rect 8324 6317 8339 6323
rect 8925 6317 8940 6323
rect 10012 6317 10060 6323
rect 892 6283 900 6290
rect 892 6277 980 6283
rect 1133 6283 1139 6314
rect 2700 6284 2708 6290
rect 6364 6284 6372 6290
rect 1133 6277 1203 6283
rect 3160 6277 3251 6283
rect 4964 6277 5027 6283
rect 6772 6277 6819 6283
rect 6957 6277 7020 6283
rect 9172 6277 9219 6283
rect 9604 6277 9651 6283
rect 9997 6277 10012 6283
rect 2052 6257 2099 6263
rect 5188 6257 5238 6263
rect 6744 6257 6780 6263
rect 234 6236 236 6244
rect 260 6237 307 6243
rect 724 6237 755 6243
rect 2516 6237 2563 6243
rect 3620 6237 3683 6243
rect 3844 6237 3907 6243
rect 4740 6237 4787 6243
rect 6509 6237 6524 6243
rect 7652 6237 7688 6243
rect 7892 6237 7907 6243
rect 8084 6237 8116 6243
rect 8724 6237 8774 6243
rect 9581 6237 9596 6243
rect 9828 6237 9860 6243
rect 10084 6237 10099 6243
rect 244 6177 307 6183
rect 1332 6177 1395 6183
rect 1556 6177 1622 6183
rect 2004 6177 2067 6183
rect 2668 6177 2684 6183
rect 3588 6177 3635 6183
rect 4476 6177 4524 6183
rect 5149 6177 5212 6183
rect 6712 6177 6748 6183
rect 7412 6177 7443 6183
rect 9172 6177 9203 6183
rect 10052 6177 10099 6183
rect 3124 6157 3187 6163
rect 5828 6157 5864 6163
rect 6036 6157 6099 6163
rect 445 6137 492 6143
rect 1533 6137 1596 6143
rect 2500 6137 2531 6143
rect 3325 6137 3388 6143
rect 4324 6137 4339 6143
rect 4996 6137 5011 6143
rect 5580 6137 5596 6143
rect 6236 6130 6244 6136
rect 6932 6137 7014 6143
rect 7386 6137 7420 6143
rect 7581 6137 7628 6143
rect 9788 6137 9836 6143
rect 6332 6130 6340 6136
rect 8108 6130 8116 6136
rect 9788 6130 9796 6137
rect 9844 6137 9852 6143
rect 9884 6130 9892 6136
rect 221 6097 252 6103
rect 2900 6097 2963 6103
rect 4237 6097 4300 6103
rect 4333 6083 4339 6103
rect 4548 6097 4563 6103
rect 9565 6097 9580 6103
rect 9800 6096 9804 6104
rect 4260 6077 4339 6083
rect 9146 6077 9180 6083
rect 7805 6037 7820 6043
rect 7860 6037 7875 6043
rect 8340 5977 8387 5983
rect 685 5917 700 5923
rect 1357 5917 1372 5923
rect 2045 5917 2060 5923
rect 2996 5917 3011 5923
rect 6781 5917 6796 5923
rect 7028 5917 7075 5923
rect 7660 5923 7668 5924
rect 7660 5917 7731 5923
rect 8086 5917 8163 5923
rect 8973 5917 8988 5923
rect 9428 5917 9475 5923
rect 9830 5917 9907 5923
rect 4476 5884 4484 5890
rect 468 5877 536 5883
rect 1124 5877 1219 5883
rect 1581 5877 1628 5883
rect 2068 5877 2131 5883
rect 2269 5877 2284 5883
rect 4500 5877 4564 5883
rect 4717 5883 4723 5914
rect 7292 5903 7300 5914
rect 7213 5897 7300 5903
rect 8749 5897 8796 5903
rect 6316 5884 6324 5890
rect 4717 5877 4803 5883
rect 4938 5877 5043 5883
rect 6852 5877 6867 5883
rect 7450 5877 7523 5883
rect 7869 5877 7955 5883
rect 9028 5877 9059 5883
rect 9194 5877 9244 5883
rect 9613 5877 9676 5883
rect 1396 5857 1443 5863
rect 1604 5857 1670 5863
rect 6340 5857 6404 5863
rect 2340 5837 2360 5843
rect 3444 5836 3446 5844
rect 3652 5837 3667 5843
rect 4292 5837 4339 5843
rect 5869 5837 5884 5843
rect 5940 5836 5944 5844
rect 6164 5837 6179 5843
rect 6580 5837 6643 5843
rect 7005 5837 7020 5843
rect 8356 5837 8387 5843
rect 8788 5837 8822 5843
rect 9405 5837 9420 5843
rect 637 5777 684 5783
rect 1336 5777 1404 5783
rect 2253 5777 2268 5783
rect 2724 5777 2772 5783
rect 3160 5777 3180 5783
rect 4029 5777 4044 5783
rect 5373 5777 5388 5783
rect 5610 5777 5660 5783
rect 6744 5777 6812 5783
rect 7181 5777 7196 5783
rect 7418 5776 7420 5784
rect 7645 5777 7692 5783
rect 8301 5777 8316 5783
rect 9162 5776 9164 5784
rect 9188 5777 9235 5783
rect 2700 5757 2748 5763
rect 1085 5737 1100 5743
rect 1565 5737 1628 5743
rect 2026 5737 2115 5743
rect 2477 5737 2563 5743
rect 5133 5737 5180 5743
rect 7028 5737 7044 5743
rect 7869 5737 7916 5743
rect 3372 5730 3380 5736
rect 708 5717 724 5723
rect 716 5706 724 5717
rect 3188 5717 3235 5723
rect 1124 5697 1187 5703
rect 2925 5697 2940 5703
rect 3386 5696 3388 5704
rect 3805 5697 3884 5703
rect 4260 5697 4340 5703
rect 5172 5697 5235 5703
rect 5396 5697 5459 5703
rect 5837 5697 5900 5703
rect 6116 5697 6132 5703
rect 7012 5697 7043 5703
rect 8077 5697 8092 5703
rect 8148 5697 8163 5703
rect 8717 5683 8723 5703
rect 8788 5697 8803 5703
rect 9892 5697 9907 5703
rect 8717 5677 8780 5683
rect 9613 5677 9692 5683
rect 5373 5637 5404 5643
rect 6744 5636 6748 5644
rect 8941 5637 8956 5643
rect 4340 5577 4355 5583
rect 8317 5577 8332 5583
rect 6532 5537 6595 5543
rect 1357 5517 1372 5523
rect 2509 5517 2524 5523
rect 2744 5516 2748 5524
rect 5428 5517 5491 5523
rect 6285 5517 6300 5523
rect 6733 5517 6748 5523
rect 7028 5517 7043 5523
rect 8356 5517 8387 5523
rect 9181 5517 9196 5523
rect 1844 5497 1907 5503
rect 3188 5497 3251 5503
rect 908 5484 916 5490
rect 468 5477 536 5483
rect 1156 5477 1219 5483
rect 1380 5477 1443 5483
rect 1581 5477 1596 5483
rect 1805 5477 1836 5483
rect 2084 5477 2147 5483
rect 2732 5483 2740 5490
rect 2532 5477 2595 5483
rect 2732 5477 2748 5483
rect 2756 5477 2804 5483
rect 2941 5477 2956 5483
rect 3388 5483 3396 5490
rect 3388 5477 3404 5483
rect 4492 5483 4500 5490
rect 4588 5484 4596 5490
rect 8172 5484 8180 5490
rect 4492 5477 4508 5483
rect 5642 5477 5708 5483
rect 6340 5477 6371 5483
rect 6756 5477 6819 5483
rect 6957 5477 7020 5483
rect 9180 5477 9267 5483
rect 9624 5477 9699 5483
rect 9860 5477 9908 5483
rect 7645 5457 7692 5463
rect 8772 5457 8822 5463
rect 68 5437 83 5443
rect 708 5437 771 5443
rect 1133 5437 1148 5443
rect 2285 5437 2300 5443
rect 2356 5436 2360 5444
rect 4733 5437 4748 5443
rect 4968 5436 4972 5444
rect 6132 5437 6147 5443
rect 6509 5437 6524 5443
rect 7181 5437 7196 5443
rect 8564 5437 8595 5443
rect 9476 5436 9480 5444
rect 1620 5377 1670 5383
rect 2068 5377 2131 5383
rect 2532 5377 2595 5383
rect 3012 5377 3059 5383
rect 3908 5377 3971 5383
rect 5508 5377 5571 5383
rect 6884 5377 6931 5383
rect 7309 5377 7372 5383
rect 8468 5377 8531 5383
rect 8948 5376 8950 5384
rect 10012 5377 10060 5383
rect 532 5356 536 5364
rect 1844 5357 1907 5363
rect 3444 5357 3510 5363
rect 4372 5357 4435 5363
rect 4589 5357 4660 5363
rect 316 5330 324 5336
rect 908 5330 916 5336
rect 2732 5330 2740 5336
rect 4589 5343 4595 5357
rect 7332 5357 7395 5363
rect 4572 5337 4595 5343
rect 2828 5330 2836 5336
rect 4572 5330 4580 5337
rect 4868 5337 4883 5343
rect 6380 5330 6388 5336
rect 8740 5337 8755 5343
rect 10036 5337 10100 5343
rect 6476 5330 6484 5336
rect 7628 5330 7636 5336
rect 10092 5330 10100 5337
rect 1148 5306 1156 5316
rect 221 5297 284 5303
rect 685 5297 772 5303
rect 1821 5297 1852 5303
rect 2045 5297 2060 5303
rect 2356 5297 2371 5303
rect 3661 5297 3747 5303
rect 3885 5297 3948 5303
rect 4349 5297 4412 5303
rect 7156 5297 7171 5303
rect 7772 5297 7859 5303
rect 7772 5296 7780 5297
rect 7997 5277 8044 5283
rect 3268 5237 3283 5243
rect 5732 5237 5779 5243
rect 6856 5237 6908 5243
rect 4093 5177 4124 5183
rect 7661 5177 7708 5183
rect 68 5117 83 5123
rect 1346 5117 1428 5123
rect 1652 5117 1667 5123
rect 2029 5117 2044 5123
rect 3165 5117 3212 5123
rect 3700 5117 3715 5123
rect 3940 5116 3942 5124
rect 4973 5117 4988 5123
rect 5284 5117 5299 5123
rect 5645 5117 5660 5123
rect 4396 5104 4404 5114
rect 892 5084 900 5090
rect 260 5077 307 5083
rect 1380 5077 1443 5083
rect 2716 5083 2724 5090
rect 2516 5077 2579 5083
rect 2716 5077 2796 5083
rect 2964 5077 3027 5083
rect 4580 5077 4612 5083
rect 4749 5077 4764 5083
rect 4970 5077 5059 5083
rect 5869 5077 5884 5083
rect 5908 5077 5958 5083
rect 6792 5077 6844 5083
rect 7508 5077 7523 5083
rect 9852 5077 9884 5083
rect 3405 5057 3452 5063
rect 234 5036 236 5044
rect 692 5037 755 5043
rect 1117 5037 1132 5043
rect 1805 5037 1820 5043
rect 2269 5037 2284 5043
rect 2324 5037 2344 5043
rect 3476 5036 3478 5044
rect 6093 5037 6108 5043
rect 7076 5036 7078 5044
rect 8333 5037 8348 5043
rect 8596 5037 8611 5043
rect 9194 5036 9196 5044
rect 20 4977 83 4983
rect 260 4977 307 4983
rect 1805 4977 1836 4983
rect 2042 4976 2044 4984
rect 3405 4977 3420 4983
rect 3629 4977 3644 4983
rect 4772 4977 4819 4983
rect 4996 4977 5043 4983
rect 6493 4977 6540 4983
rect 7620 4977 7640 4983
rect 8456 4976 8460 4984
rect 8484 4977 8531 4983
rect 461 4957 536 4963
rect 2269 4957 2344 4963
rect 461 4943 467 4957
rect 445 4937 467 4943
rect 2269 4943 2275 4957
rect 3652 4957 3715 4963
rect 2253 4937 2275 4943
rect 5389 4937 5452 4943
rect 9114 4937 9164 4943
rect 9533 4937 9580 4943
rect 9965 4937 10040 4943
rect 908 4930 916 4936
rect 4604 4930 4612 4936
rect 6348 4930 6356 4936
rect 2732 4917 2764 4923
rect 6925 4917 6972 4923
rect 7868 4906 7876 4916
rect 221 4897 252 4903
rect 460 4897 508 4903
rect 685 4897 772 4903
rect 920 4897 940 4903
rect 2268 4897 2316 4903
rect 2493 4897 2508 4903
rect 2532 4897 2579 4903
rect 3853 4897 3868 4903
rect 4509 4897 4524 4903
rect 5405 4897 5475 4903
rect 5613 4897 5628 4903
rect 6045 4897 6116 4903
rect 7172 4897 7219 4903
rect 8893 4897 8963 4903
rect 9750 4897 9827 4903
rect 6268 4877 6332 4883
rect 6516 4877 6563 4883
rect 1412 4857 1427 4863
rect 4301 4857 4348 4863
rect 7370 4836 7372 4844
rect 9325 4837 9340 4843
rect 3236 4777 3251 4783
rect 5853 4777 5916 4783
rect 8324 4777 8355 4783
rect 7821 4737 7836 4743
rect 532 4716 542 4724
rect 1357 4717 1372 4723
rect 2052 4717 2102 4723
rect 2788 4717 2796 4723
rect 3165 4717 3196 4723
rect 3402 4716 3404 4724
rect 6285 4717 6300 4723
rect 6980 4717 7027 4723
rect 8029 4717 8044 4723
rect 9830 4717 9907 4723
rect 10100 4717 10115 4723
rect 908 4684 916 4690
rect 2700 4684 2708 4690
rect 708 4677 771 4683
rect 2100 4677 2115 4683
rect 2724 4677 2803 4683
rect 3388 4683 3396 4690
rect 3388 4677 3462 4683
rect 4045 4677 4136 4683
rect 4308 4677 4355 4683
rect 4964 4677 5027 4683
rect 5165 4677 5180 4683
rect 6077 4677 6124 4683
rect 6308 4677 6356 4683
rect 6493 4677 6508 4683
rect 6941 4677 6972 4683
rect 8029 4677 8116 4683
rect 9220 4677 9235 4683
rect 9396 4677 9448 4683
rect 10045 4677 10120 4683
rect 1604 4657 1654 4663
rect 2964 4657 3027 4663
rect 234 4636 236 4644
rect 292 4637 307 4643
rect 932 4637 996 4643
rect 2276 4637 2328 4643
rect 2532 4637 2563 4643
rect 2941 4637 2956 4643
rect 3892 4637 3907 4643
rect 4740 4637 4803 4643
rect 5405 4637 5468 4643
rect 5642 4636 5644 4644
rect 6744 4636 6748 4644
rect 7844 4637 7891 4643
rect 8292 4637 8355 4643
rect 8948 4637 9011 4643
rect 9373 4637 9388 4643
rect 20 4577 83 4583
rect 1412 4577 1459 4583
rect 2058 4577 2092 4583
rect 2116 4577 2131 4583
rect 2308 4577 2360 4583
rect 3204 4577 3251 4583
rect 3476 4576 3478 4584
rect 4308 4577 4371 4583
rect 6324 4577 6356 4583
rect 7012 4577 7030 4583
rect 8292 4577 8339 4583
rect 8701 4577 8732 4583
rect 461 4557 524 4563
rect 8269 4557 8316 4563
rect 8724 4557 8758 4563
rect 9588 4557 9651 4563
rect 4061 4537 4076 4543
rect 4717 4537 4732 4543
rect 4968 4537 5043 4543
rect 7172 4537 7212 4543
rect 7460 4537 7475 4543
rect 8916 4537 8995 4543
rect 9412 4536 9416 4544
rect 9860 4537 9892 4543
rect 316 4530 324 4536
rect 908 4530 916 4536
rect 1596 4530 1604 4536
rect 3388 4530 3396 4536
rect 4508 4530 4516 4536
rect 8124 4530 8132 4536
rect 9788 4530 9796 4536
rect 9884 4530 9892 4537
rect 1148 4517 1180 4523
rect 1148 4506 1156 4517
rect 3628 4517 3676 4523
rect 3628 4506 3636 4517
rect 6300 4517 6332 4523
rect 7402 4517 7436 4523
rect 8044 4517 8067 4523
rect 221 4497 252 4503
rect 484 4497 547 4503
rect 920 4497 1002 4503
rect 2509 4497 2524 4503
rect 2717 4497 2764 4503
rect 4520 4496 4524 4504
rect 4756 4497 4819 4503
rect 7612 4497 7683 4503
rect 7612 4496 7620 4497
rect 8061 4503 8067 4517
rect 8061 4497 8120 4503
rect 9796 4497 9852 4503
rect 10237 4497 10252 4503
rect 756 4457 771 4463
rect 3012 4457 3027 4463
rect 6061 4457 6140 4463
rect 3668 4437 3715 4443
rect 5460 4437 5475 4443
rect 6744 4436 6748 4444
rect 7821 4437 7836 4443
rect 10084 4437 10099 4443
rect 1149 4377 1164 4383
rect 1652 4376 1654 4384
rect 3188 4377 3235 4383
rect 8765 4377 8812 4383
rect 8557 4337 8620 4343
rect 460 4317 492 4323
rect 2029 4317 2044 4323
rect 3597 4317 3612 4323
rect 4877 4317 4924 4323
rect 7901 4317 7916 4323
rect 9405 4317 9420 4323
rect 9908 4317 9923 4323
rect 908 4284 916 4290
rect 445 4277 460 4283
rect 1004 4284 1012 4290
rect 2700 4284 2708 4290
rect 1354 4277 1443 4283
rect 1812 4277 1891 4283
rect 2796 4283 2804 4290
rect 2724 4277 2804 4283
rect 3373 4277 3446 4283
rect 4013 4277 4060 4283
rect 5530 4277 5603 4283
rect 5764 4277 5800 4283
rect 7037 4277 7052 4283
rect 9428 4277 9475 4283
rect 2941 4257 3004 4263
rect 4692 4257 4739 4263
rect 6196 4257 6244 4263
rect 20 4237 83 4243
rect 244 4237 307 4243
rect 1204 4237 1219 4243
rect 2084 4237 2115 4243
rect 2964 4237 3027 4243
rect 3428 4237 3446 4243
rect 4460 4237 4476 4243
rect 4932 4237 4947 4243
rect 5741 4237 5756 4243
rect 6468 4237 6483 4243
rect 6676 4237 6691 4243
rect 6900 4236 6902 4244
rect 7748 4237 7763 4243
rect 8986 4236 8988 4244
rect 932 4177 980 4183
rect 1620 4177 1670 4183
rect 2500 4177 2563 4183
rect 2724 4177 2788 4183
rect 2964 4177 3027 4183
rect 3236 4177 3251 4183
rect 3428 4177 3478 4183
rect 3652 4177 3699 4183
rect 4301 4177 4316 4183
rect 5885 4177 5932 4183
rect 6776 4176 6780 4184
rect 8116 4177 8148 4183
rect 8532 4177 8595 4183
rect 8820 4176 8822 4184
rect 9194 4177 9212 4183
rect 9852 4177 9884 4183
rect 10061 4177 10268 4183
rect 908 4157 940 4163
rect 1844 4157 1891 4163
rect 4772 4157 4835 4163
rect 5268 4156 5270 4164
rect 8324 4157 8371 4163
rect 1396 4137 1443 4143
rect 1581 4137 1596 4143
rect 2237 4137 2328 4143
rect 3388 4137 3404 4143
rect 316 4130 324 4136
rect 2700 4130 2708 4136
rect 3388 4130 3396 4137
rect 4061 4137 4124 4143
rect 4372 4137 4387 4143
rect 4524 4137 4540 4143
rect 4524 4130 4532 4137
rect 4733 4137 4748 4143
rect 6557 4137 6632 4143
rect 8076 4137 8124 4143
rect 9700 4137 9715 4143
rect 8732 4130 8740 4136
rect 9276 4130 9284 4136
rect 3668 4117 3699 4123
rect 3860 4117 3923 4123
rect 7629 4117 7676 4123
rect 8300 4117 8348 4123
rect 1820 4106 1828 4116
rect 8300 4106 8308 4117
rect 9421 4117 9468 4123
rect 221 4097 236 4103
rect 1362 4097 1420 4103
rect 2029 4097 2076 4103
rect 2941 4097 2956 4103
rect 4148 4097 4163 4103
rect 5645 4097 5660 4103
rect 6989 4097 7059 4103
rect 6109 4057 6188 4063
rect 5492 4037 5507 4043
rect 3460 3976 3462 3984
rect 6541 3977 6588 3983
rect 6996 3977 7030 3983
rect 221 3917 236 3923
rect 904 3916 908 3924
rect 2685 3917 2732 3923
rect 3149 3917 3196 3923
rect 3837 3917 3852 3923
rect 4301 3917 4332 3923
rect 5268 3917 5283 3923
rect 8100 3917 8115 3923
rect 8461 3917 8476 3923
rect 9117 3917 9132 3923
rect 9860 3917 9875 3923
rect 3612 3904 3620 3914
rect 1565 3897 1612 3903
rect 429 3877 520 3883
rect 892 3883 900 3890
rect 3372 3884 3380 3890
rect 892 3877 964 3883
rect 1101 3877 1116 3883
rect 1336 3877 1427 3883
rect 2237 3877 2328 3883
rect 2964 3877 3011 3883
rect 5421 3877 5484 3883
rect 6332 3877 6403 3883
rect 8484 3877 8547 3883
rect 8877 3877 8979 3883
rect 2724 3857 2772 3863
rect 5658 3857 5708 3863
rect 740 3837 755 3843
rect 1636 3836 1638 3844
rect 2532 3837 2547 3843
rect 3652 3837 3699 3843
rect 4749 3837 4764 3843
rect 4984 3836 4988 3844
rect 5213 3837 5260 3843
rect 6596 3837 6611 3843
rect 7821 3837 7836 3843
rect 8253 3837 8300 3843
rect 8685 3837 8700 3843
rect 8740 3836 8742 3844
rect 9804 3837 9820 3843
rect 10232 3836 10236 3844
rect 20 3777 83 3783
rect 260 3777 307 3783
rect 708 3777 771 3783
rect 932 3777 980 3783
rect 1156 3777 1219 3783
rect 2052 3777 2115 3783
rect 2756 3777 2804 3783
rect 3428 3777 3494 3783
rect 4148 3776 4152 3784
rect 4564 3777 4596 3783
rect 4804 3777 4835 3783
rect 5284 3776 5286 3784
rect 7012 3777 7046 3783
rect 7220 3777 7267 3783
rect 7684 3777 7720 3783
rect 7924 3777 7939 3783
rect 8317 3777 8364 3783
rect 8749 3777 8764 3783
rect 8996 3777 9043 3783
rect 9836 3777 9852 3783
rect 10045 3777 10076 3783
rect 10100 3777 10115 3783
rect 1844 3757 1891 3763
rect 2276 3757 2344 3763
rect 2980 3757 3043 3763
rect 7645 3757 7692 3763
rect 9405 3757 9452 3763
rect 468 3737 536 3743
rect 908 3737 940 3743
rect 908 3730 916 3737
rect 1117 3737 1132 3743
rect 1581 3737 1628 3743
rect 3716 3737 3731 3743
rect 6332 3737 6403 3743
rect 7476 3737 7507 3743
rect 8077 3737 8108 3743
rect 6972 3730 6980 3736
rect 8172 3730 8180 3736
rect 6541 3717 6588 3723
rect 8973 3717 9020 3723
rect 221 3697 236 3703
rect 685 3697 700 3703
rect 1357 3697 1443 3703
rect 1821 3697 1852 3703
rect 2493 3697 2540 3703
rect 2726 3697 2780 3703
rect 3181 3697 3228 3703
rect 3645 3697 3692 3703
rect 4973 3697 4988 3703
rect 5885 3697 5955 3703
rect 7869 3697 7884 3703
rect 8077 3697 8140 3703
rect 3188 3677 3267 3683
rect 6093 3677 6172 3683
rect 8605 3683 8611 3703
rect 9613 3697 9684 3703
rect 9860 3697 9907 3703
rect 10253 3697 10268 3703
rect 8536 3677 8611 3683
rect 5674 3657 5756 3663
rect 5012 3637 5059 3643
rect 6760 3636 6764 3644
rect 68 3577 83 3583
rect 4996 3577 5011 3583
rect 6948 3557 6998 3563
rect 1204 3517 1219 3523
rect 2941 3517 2956 3523
rect 3165 3517 3180 3523
rect 3821 3517 3836 3523
rect 4516 3517 4568 3523
rect 5396 3517 5459 3523
rect 6340 3517 6355 3523
rect 7149 3517 7164 3523
rect 8054 3517 8124 3523
rect 8788 3517 8803 3523
rect 1132 3504 1140 3514
rect 1668 3496 1670 3504
rect 1820 3503 1828 3514
rect 1820 3497 1843 3503
rect 6493 3497 6540 3503
rect 244 3477 307 3483
rect 892 3483 900 3490
rect 664 3477 755 3483
rect 892 3477 956 3483
rect 1444 3477 1459 3483
rect 1837 3483 1843 3497
rect 2700 3484 2708 3490
rect 4476 3484 4484 3490
rect 1837 3477 1891 3483
rect 2276 3477 2328 3483
rect 2724 3477 2788 3483
rect 3844 3477 3891 3483
rect 4572 3484 4580 3490
rect 5148 3484 5156 3490
rect 6284 3477 6355 3483
rect 6712 3477 6787 3483
rect 8116 3477 8124 3483
rect 9836 3477 9900 3483
rect 1597 3457 1644 3463
rect 3620 3457 3683 3463
rect 2052 3437 2115 3443
rect 4324 3437 4339 3443
rect 5220 3436 5222 3444
rect 5610 3436 5612 3444
rect 6045 3437 6060 3443
rect 7386 3436 7388 3444
rect 8941 3437 8988 3443
rect 9162 3436 9164 3444
rect 9373 3437 9388 3443
rect 9597 3437 9612 3443
rect 68 3377 83 3383
rect 1149 3377 1180 3383
rect 1444 3377 1459 3383
rect 3652 3377 3715 3383
rect 4340 3377 4371 3383
rect 5658 3377 5692 3383
rect 6093 3377 6108 3383
rect 6340 3377 6388 3383
rect 7005 3377 7068 3383
rect 8108 3377 8124 3383
rect 8333 3377 8348 3383
rect 8989 3377 9036 3383
rect 2509 3357 2556 3363
rect 2980 3357 3043 3363
rect 3204 3357 3267 3363
rect 3421 3357 3478 3363
rect 445 3337 508 3343
rect 908 3337 940 3343
rect 908 3330 916 3337
rect 2058 3337 2124 3343
rect 2717 3337 2796 3343
rect 3421 3343 3427 3357
rect 4756 3357 4819 3363
rect 9652 3357 9699 3363
rect 3405 3337 3427 3343
rect 4061 3337 4076 3343
rect 4717 3337 4732 3343
rect 6116 3337 6140 3343
rect 6852 3337 6867 3343
rect 7450 3337 7484 3343
rect 7645 3337 7708 3343
rect 9252 3337 9283 3343
rect 9421 3337 9494 3343
rect 1004 3330 1012 3336
rect 1596 3330 1604 3336
rect 2140 3330 2148 3336
rect 2812 3330 2820 3336
rect 4508 3330 4516 3336
rect 8188 3330 8196 3336
rect 685 3297 772 3303
rect 1378 3297 1436 3303
rect 2132 3296 2134 3304
rect 2717 3297 2732 3303
rect 3181 3297 3228 3303
rect 3853 3297 3923 3303
rect 4100 3297 4147 3303
rect 4520 3296 4524 3304
rect 4957 3297 5043 3303
rect 5220 3297 5283 3303
rect 7076 3297 7091 3303
rect 7716 3297 7731 3303
rect 7229 3277 7308 3283
rect 8637 3283 8643 3303
rect 8781 3297 8851 3303
rect 9277 3283 9283 3303
rect 9908 3297 9923 3303
rect 8568 3277 8643 3283
rect 9210 3277 9283 3283
rect 5421 3237 5436 3243
rect 5869 3237 5884 3243
rect 708 3177 739 3183
rect 8580 3176 8582 3184
rect 8996 3137 9027 3143
rect 205 3117 284 3123
rect 1330 3117 1372 3123
rect 1620 3117 1635 3123
rect 2429 3117 2476 3123
rect 2500 3117 2515 3123
rect 3164 3123 3172 3124
rect 3156 3117 3172 3123
rect 5917 3117 5988 3123
rect 6164 3117 6211 3123
rect 7450 3117 7523 3123
rect 7869 3117 7884 3123
rect 8733 3117 8803 3123
rect 9021 3117 9027 3137
rect 9165 3117 9212 3123
rect 9389 3117 9452 3123
rect 10045 3117 10060 3123
rect 429 3077 492 3083
rect 876 3083 884 3090
rect 876 3077 948 3083
rect 1533 3077 1548 3083
rect 1773 3077 1852 3083
rect 3308 3083 3316 3090
rect 3308 3077 3324 3083
rect 3348 3077 3398 3083
rect 3981 3077 4056 3083
rect 7869 3077 7916 3083
rect 8116 3077 8163 3083
rect 8717 3077 8732 3083
rect 9628 3077 9699 3083
rect 653 3057 716 3063
rect 2010 3057 2044 3063
rect 4660 3057 4707 3063
rect 5709 3037 5724 3043
rect 6568 3036 6572 3044
rect 6797 3037 6812 3043
rect 7028 3037 7091 3043
rect 7716 3037 7731 3043
rect 8954 3036 8956 3044
rect 1332 2977 1395 2983
rect 1556 2977 1622 2983
rect 1796 2977 1859 2983
rect 2724 2977 2756 2983
rect 2932 2977 2995 2983
rect 3172 2977 3219 2983
rect 3380 2977 3446 2983
rect 4492 2977 4524 2983
rect 4756 2977 4787 2983
rect 7354 2977 7404 2983
rect 8701 2977 8716 2983
rect 8740 2977 8774 2983
rect 8996 2977 9011 2983
rect 4052 2957 4104 2963
rect 5828 2957 5880 2963
rect 948 2937 964 2943
rect 956 2930 964 2937
rect 1533 2937 1548 2943
rect 3357 2937 3420 2943
rect 4013 2937 4028 2943
rect 5156 2937 5222 2943
rect 5789 2937 5804 2943
rect 6260 2937 6340 2943
rect 2684 2930 2692 2936
rect 6332 2930 6340 2937
rect 8012 2930 8020 2936
rect 9916 2930 9924 2936
rect 876 2917 899 2923
rect 76 2906 84 2916
rect 893 2903 899 2917
rect 3596 2917 3667 2923
rect 6696 2917 6748 2923
rect 3596 2904 3604 2917
rect 9668 2917 9684 2923
rect 9676 2904 9684 2917
rect 893 2897 952 2903
rect 1546 2897 1596 2903
rect 1773 2897 1836 2903
rect 2696 2896 2700 2904
rect 3133 2897 3196 2903
rect 4548 2897 4563 2903
rect 5373 2897 5443 2903
rect 6029 2897 6060 2903
rect 6980 2897 6995 2903
rect 7580 2897 7596 2903
rect 8084 2897 8099 2903
rect 8925 2897 8940 2903
rect 9597 2897 9612 2903
rect 234 2837 268 2843
rect 6477 2837 6492 2843
rect 6756 2837 6771 2843
rect 7133 2837 7164 2843
rect 9444 2836 9448 2844
rect 1821 2777 1836 2783
rect 1860 2777 1891 2783
rect 6413 2777 6444 2783
rect 7069 2777 7100 2783
rect 9869 2777 9916 2783
rect 221 2717 236 2723
rect 685 2717 700 2723
rect 1149 2717 1180 2723
rect 1668 2717 1683 2723
rect 3133 2717 3148 2723
rect 3357 2717 3404 2723
rect 3805 2717 3836 2723
rect 5757 2717 5827 2723
rect 6900 2717 6931 2723
rect 9421 2717 9436 2723
rect 9668 2717 9720 2723
rect 6036 2697 6051 2703
rect 9644 2697 9692 2703
rect 244 2677 307 2683
rect 468 2677 536 2683
rect 908 2683 916 2690
rect 708 2677 771 2683
rect 908 2677 996 2683
rect 1428 2677 1459 2683
rect 2700 2683 2708 2690
rect 6188 2684 6196 2690
rect 9724 2684 9732 2690
rect 2700 2677 2748 2683
rect 6660 2677 6723 2683
rect 7290 2677 7363 2683
rect 7709 2677 7795 2683
rect 8628 2676 8630 2684
rect 9220 2677 9272 2683
rect 1597 2657 1660 2663
rect 2500 2657 2563 2663
rect 68 2637 83 2643
rect 2084 2637 2115 2643
rect 2756 2637 2772 2643
rect 3428 2636 3430 2644
rect 3652 2637 3667 2643
rect 4460 2637 4476 2643
rect 4516 2637 4532 2643
rect 5117 2637 5148 2643
rect 5965 2637 5980 2643
rect 6484 2637 6499 2643
rect 6861 2637 6876 2643
rect 9002 2636 9004 2644
rect 234 2576 236 2584
rect 260 2577 307 2583
rect 685 2577 700 2583
rect 924 2577 940 2583
rect 1581 2577 1596 2583
rect 3204 2577 3251 2583
rect 3444 2577 3478 2583
rect 3668 2577 3715 2583
rect 3876 2577 3939 2583
rect 5453 2577 5484 2583
rect 7012 2577 7046 2583
rect 7668 2577 7720 2583
rect 8116 2577 8148 2583
rect 8733 2577 8764 2583
rect 4100 2557 4168 2563
rect 7220 2557 7283 2563
rect 7892 2557 7939 2563
rect 1428 2537 1443 2543
rect 1828 2537 1891 2543
rect 2500 2537 2563 2543
rect 2700 2537 2764 2543
rect 2700 2530 2708 2537
rect 4388 2537 4403 2543
rect 4540 2537 4556 2543
rect 2796 2530 2804 2536
rect 4540 2530 4548 2537
rect 6348 2537 6419 2543
rect 7181 2537 7196 2543
rect 9012 2537 9027 2543
rect 9892 2537 9940 2543
rect 5756 2530 5764 2536
rect 9932 2530 9940 2537
rect 5674 2517 5699 2523
rect 68 2497 83 2503
rect 500 2497 547 2503
rect 708 2497 771 2503
rect 2029 2497 2044 2503
rect 2477 2497 2540 2503
rect 2712 2497 2748 2503
rect 3853 2497 3884 2503
rect 4092 2497 4108 2503
rect 4781 2497 4851 2503
rect 5309 2484 5315 2503
rect 5693 2503 5699 2517
rect 5693 2497 5750 2503
rect 6404 2497 6419 2503
rect 6765 2497 6780 2503
rect 7869 2497 7884 2503
rect 8788 2497 8803 2503
rect 9876 2497 9928 2503
rect 5229 2477 5308 2483
rect 516 2376 520 2384
rect 7274 2376 7276 2384
rect 4173 2337 4236 2343
rect 7916 2337 7980 2343
rect 444 2317 492 2323
rect 1562 2317 1596 2323
rect 1997 2317 2012 2323
rect 3085 2317 3100 2323
rect 4845 2317 4860 2323
rect 5300 2317 5347 2323
rect 5524 2317 5574 2323
rect 7485 2317 7555 2323
rect 7972 2317 7987 2323
rect 204 2277 291 2283
rect 429 2277 492 2283
rect 692 2277 739 2283
rect 1117 2283 1123 2314
rect 1548 2284 1556 2290
rect 4396 2284 4404 2290
rect 1117 2277 1187 2283
rect 2861 2277 2876 2283
rect 3724 2277 3788 2283
rect 4492 2283 4500 2290
rect 4420 2277 4500 2283
rect 4868 2277 4931 2283
rect 5498 2277 5587 2283
rect 6252 2283 6260 2290
rect 6244 2277 6260 2283
rect 6397 2277 6472 2283
rect 6845 2277 6892 2283
rect 8404 2277 8419 2283
rect 8788 2277 8851 2283
rect 8986 2276 8988 2284
rect 8557 2257 8604 2263
rect 1396 2237 1411 2243
rect 4196 2237 4259 2243
rect 5933 2237 5948 2243
rect 6616 2236 6620 2244
rect 7053 2237 7068 2243
rect 7693 2237 7708 2243
rect 8180 2237 8195 2243
rect 9405 2237 9420 2243
rect 9460 2237 9475 2243
rect 10056 2236 10060 2244
rect 234 2176 236 2184
rect 724 2177 739 2183
rect 1812 2177 1875 2183
rect 2500 2177 2547 2183
rect 3428 2177 3462 2183
rect 3636 2177 3699 2183
rect 4084 2177 4136 2183
rect 4980 2177 5027 2183
rect 6957 2177 6972 2183
rect 7629 2177 7660 2183
rect 7837 2177 7852 2183
rect 8269 2177 8300 2183
rect 1565 2157 1638 2163
rect 2701 2157 2772 2163
rect 5181 2157 5254 2163
rect 6300 2157 6364 2163
rect 877 2137 956 2143
rect 1565 2143 1571 2157
rect 1548 2137 1571 2143
rect 316 2130 324 2136
rect 972 2130 980 2136
rect 1548 2130 1556 2137
rect 2237 2137 2312 2143
rect 2701 2143 2707 2157
rect 2684 2137 2707 2143
rect 2684 2130 2692 2137
rect 3160 2137 3251 2143
rect 4308 2137 4355 2143
rect 5181 2143 5187 2157
rect 5165 2137 5187 2143
rect 6077 2137 6163 2143
rect 6744 2137 6819 2143
rect 8996 2137 9011 2143
rect 6380 2130 6388 2136
rect 68 2117 84 2123
rect 76 2106 84 2117
rect 1788 2117 1836 2123
rect 1788 2106 1796 2117
rect 308 2096 310 2104
rect 877 2097 892 2103
rect 964 2096 968 2104
rect 2013 2097 2044 2103
rect 2052 2097 2060 2103
rect 2252 2097 2284 2103
rect 2461 2097 2476 2103
rect 3613 2097 3628 2103
rect 3837 2097 3852 2103
rect 4285 2097 4300 2103
rect 4716 2097 4803 2103
rect 5405 2097 5420 2103
rect 5629 2097 5644 2103
rect 5892 2097 5939 2103
rect 8772 2097 8787 2103
rect 9188 2097 9238 2103
rect 9388 2097 9459 2103
rect 9388 2096 9396 2097
rect 9597 2097 9668 2103
rect 9814 2097 9891 2103
rect 10028 2097 10099 2103
rect 1117 2077 1164 2083
rect 1396 2037 1411 2043
rect 5853 1977 5884 1983
rect 6941 1977 6956 1983
rect 7386 1976 7388 1984
rect 8269 1977 8284 1983
rect 6061 1937 6108 1943
rect 6964 1937 7020 1943
rect 7188 1937 7244 1943
rect 7412 1937 7459 1943
rect 1325 1917 1340 1923
rect 1396 1917 1412 1923
rect 2696 1916 2700 1924
rect 3613 1917 3628 1923
rect 3837 1917 3852 1923
rect 4756 1917 4803 1923
rect 5188 1917 5228 1923
rect 5236 1917 5251 1923
rect 5389 1917 5475 1923
rect 6269 1917 6284 1923
rect 6980 1917 7027 1923
rect 7188 1917 7235 1923
rect 7453 1917 7459 1937
rect 8996 1917 9011 1923
rect 9597 1917 9628 1923
rect 10028 1917 10099 1923
rect 956 1884 964 1890
rect 2684 1884 2692 1890
rect 204 1877 291 1883
rect 1796 1877 1868 1883
rect 2237 1877 2268 1883
rect 2276 1877 2326 1883
rect 2780 1883 2788 1890
rect 3372 1884 3380 1890
rect 5708 1884 5716 1890
rect 2724 1877 2788 1883
rect 3860 1877 3923 1883
rect 4061 1877 4076 1883
rect 6292 1877 6356 1883
rect 6509 1883 6515 1914
rect 8124 1884 8132 1890
rect 6509 1877 6579 1883
rect 7165 1877 7251 1883
rect 8580 1877 8595 1883
rect 9389 1877 9420 1883
rect 9668 1877 9683 1883
rect 9820 1877 9891 1883
rect 1101 1857 1164 1863
rect 1565 1857 1612 1863
rect 2484 1857 2547 1863
rect 2925 1857 2972 1863
rect 3160 1857 3180 1863
rect 1588 1837 1638 1843
rect 3444 1837 3462 1843
rect 3684 1837 3699 1843
rect 4308 1837 4355 1843
rect 4532 1837 4580 1843
rect 5626 1836 5628 1844
rect 6084 1837 6131 1843
rect 6941 1837 6956 1843
rect 8504 1837 8540 1843
rect 8733 1837 8748 1843
rect 8941 1837 8956 1843
rect 9444 1836 9448 1844
rect 10248 1836 10252 1844
rect 260 1777 307 1783
rect 1581 1777 1628 1783
rect 1652 1776 1654 1784
rect 3176 1777 3212 1783
rect 3613 1777 3628 1783
rect 3834 1776 3836 1784
rect 4045 1777 4076 1783
rect 4100 1777 4120 1783
rect 4936 1777 4956 1783
rect 6292 1777 6324 1783
rect 6925 1777 6972 1783
rect 7149 1777 7180 1783
rect 7597 1777 7644 1783
rect 8285 1777 8316 1783
rect 3220 1757 3235 1763
rect 892 1737 980 1743
rect 972 1730 980 1737
rect 2052 1737 2115 1743
rect 2276 1737 2344 1743
rect 3373 1737 3404 1743
rect 4996 1737 5011 1743
rect 6268 1737 6284 1743
rect 8520 1737 8595 1743
rect 8733 1737 8804 1743
rect 9162 1737 9235 1743
rect 9620 1737 9667 1743
rect 10013 1737 10088 1743
rect 2796 1730 2804 1736
rect 5148 1730 5156 1736
rect 8140 1730 8148 1736
rect 7844 1717 7908 1723
rect 76 1706 84 1716
rect 7900 1706 7908 1717
rect 932 1697 968 1703
rect 1412 1697 1428 1703
rect 1805 1697 1868 1703
rect 2493 1697 2564 1703
rect 4269 1697 4340 1703
rect 4548 1697 4563 1703
rect 5162 1696 5164 1704
rect 5188 1697 5251 1703
rect 5389 1697 5459 1703
rect 5677 1683 5683 1703
rect 6029 1697 6115 1703
rect 6476 1697 6492 1703
rect 6996 1697 7011 1703
rect 7357 1697 7372 1703
rect 8308 1697 8371 1703
rect 8756 1697 8803 1703
rect 8964 1697 9011 1703
rect 9372 1697 9443 1703
rect 9581 1697 9652 1703
rect 9372 1696 9380 1697
rect 5610 1677 5683 1683
rect 892 1657 940 1663
rect 6452 1657 6563 1663
rect 4717 1577 4764 1583
rect 5149 1577 5180 1583
rect 6029 1577 6044 1583
rect 6500 1577 6563 1583
rect 1404 1523 1412 1524
rect 1341 1517 1412 1523
rect 1844 1517 1859 1523
rect 2925 1517 2940 1523
rect 3613 1517 3660 1523
rect 3837 1517 3868 1523
rect 4084 1517 4147 1523
rect 5581 1517 5596 1523
rect 6964 1517 7011 1523
rect 7612 1523 7620 1524
rect 7612 1517 7683 1523
rect 8029 1517 8044 1523
rect 9828 1517 9843 1523
rect 8972 1504 8980 1514
rect 892 1497 924 1503
rect 972 1484 980 1490
rect 1156 1477 1203 1483
rect 1549 1477 1612 1483
rect 1773 1477 1852 1483
rect 2092 1483 2100 1490
rect 2010 1477 2100 1483
rect 2237 1477 2300 1483
rect 2461 1477 2540 1483
rect 2932 1477 3011 1483
rect 3372 1483 3380 1490
rect 7468 1484 7476 1490
rect 3172 1477 3235 1483
rect 3372 1477 3436 1483
rect 3460 1476 3462 1484
rect 5364 1477 5443 1483
rect 5604 1477 5651 1483
rect 6237 1477 6324 1483
rect 8260 1477 8323 1483
rect 8516 1477 8547 1483
rect 8877 1477 8940 1483
rect 9549 1477 9596 1483
rect 9780 1477 9843 1483
rect 9981 1477 10056 1483
rect 7821 1457 7868 1463
rect 9572 1457 9619 1463
rect 68 1437 83 1443
rect 2010 1437 2044 1443
rect 2724 1437 2772 1443
rect 3636 1437 3699 1443
rect 4308 1437 4355 1443
rect 7149 1437 7164 1443
rect 7386 1437 7404 1443
rect 7876 1437 7891 1443
rect 8685 1437 8700 1443
rect 8740 1436 8742 1444
rect 9130 1436 9132 1444
rect 1380 1377 1427 1383
rect 1805 1377 1836 1383
rect 3357 1377 3388 1383
rect 4324 1377 4339 1383
rect 5357 1377 5372 1383
rect 5594 1377 5644 1383
rect 6493 1377 6508 1383
rect 6712 1376 6716 1384
rect 7386 1376 7388 1384
rect 7821 1377 7852 1383
rect 8504 1376 8508 1384
rect 8532 1377 8563 1383
rect 9162 1376 9164 1384
rect 9860 1377 9892 1383
rect 3812 1357 3875 1363
rect 932 1337 980 1343
rect 972 1330 980 1337
rect 1565 1337 1580 1343
rect 3204 1337 3219 1343
rect 4013 1337 4060 1343
rect 4906 1337 5011 1343
rect 6100 1337 6131 1343
rect 7188 1337 7251 1343
rect 8060 1337 8131 1343
rect 8941 1337 9027 1343
rect 9389 1337 9462 1343
rect 9836 1337 9868 1343
rect 6348 1330 6356 1336
rect 444 1297 531 1303
rect 444 1296 452 1297
rect 2052 1297 2108 1303
rect 2461 1297 2476 1303
rect 3156 1297 3204 1303
rect 3789 1297 3804 1303
rect 4028 1297 4044 1303
rect 4253 1297 4284 1303
rect 4477 1297 4524 1303
rect 4909 1297 4924 1303
rect 6045 1297 6116 1303
rect 6548 1297 6563 1303
rect 7012 1297 7027 1303
rect 7165 1297 7235 1303
rect 7668 1297 7683 1303
rect 8701 1283 8707 1303
rect 8788 1297 8803 1303
rect 9412 1297 9459 1303
rect 8701 1277 8796 1283
rect 234 1236 236 1244
rect 1352 1236 1356 1244
rect 1844 1237 1891 1243
rect 4068 1237 4104 1243
rect 5149 1177 5164 1183
rect 6525 1177 6556 1183
rect 5172 1157 5222 1163
rect 669 1117 684 1123
rect 916 1117 940 1123
rect 948 1117 963 1123
rect 1124 1117 1187 1123
rect 1364 1117 1412 1123
rect 1789 1117 1836 1123
rect 2461 1117 2476 1123
rect 3101 1117 3164 1123
rect 4300 1123 4308 1124
rect 4244 1117 4308 1123
rect 4532 1117 4547 1123
rect 5917 1117 5923 1136
rect 7044 1117 7059 1123
rect 7405 1117 7452 1123
rect 8045 1117 8060 1123
rect 9165 1117 9180 1123
rect 9388 1123 9396 1124
rect 9388 1117 9459 1123
rect 892 1097 940 1103
rect 1101 1097 1164 1103
rect 1336 1097 1388 1103
rect 244 1077 307 1083
rect 445 1077 460 1083
rect 1364 1077 1427 1083
rect 1828 1077 1875 1083
rect 2484 1077 2531 1083
rect 2877 1077 2892 1083
rect 3325 1077 3340 1083
rect 4445 1077 4460 1083
rect 5610 1077 5699 1083
rect 5837 1077 5900 1083
rect 6084 1077 6140 1083
rect 6380 1083 6388 1090
rect 9820 1084 9828 1090
rect 6324 1077 6388 1083
rect 7404 1077 7491 1083
rect 8045 1077 8116 1083
rect 8253 1077 8284 1083
rect 8724 1077 8790 1083
rect 9916 1084 9924 1090
rect 3549 1057 3580 1063
rect 7197 1057 7244 1063
rect 7860 1057 7907 1063
rect 1636 1036 1638 1044
rect 2260 1037 2312 1043
rect 2932 1037 2963 1043
rect 3124 1037 3187 1043
rect 6760 1036 6764 1044
rect 7220 1037 7267 1043
rect 7629 1037 7644 1043
rect 8516 1037 8563 1043
rect 8964 1037 9027 1043
rect 9668 1037 9683 1043
rect 468 977 520 983
rect 692 977 755 983
rect 932 977 980 983
rect 2010 977 2060 983
rect 2260 977 2312 983
rect 3325 977 3340 983
rect 3780 977 3827 983
rect 4052 976 4056 984
rect 5588 977 5651 983
rect 6477 977 6524 983
rect 6712 977 6748 983
rect 8044 977 8060 983
rect 8084 977 8100 983
rect 8724 977 8774 983
rect 9389 977 9404 983
rect 9428 977 9448 983
rect 6029 957 6092 963
rect 9620 957 9683 963
rect 2221 937 2284 943
rect 3965 937 4056 943
rect 4429 937 4460 943
rect 6268 937 6339 943
rect 6932 937 6998 943
rect 8237 937 8328 943
rect 9172 937 9251 943
rect 892 930 900 936
rect 9820 930 9828 936
rect 1852 906 1860 916
rect 221 897 291 903
rect 669 897 684 903
rect 2461 897 2476 903
rect 2948 897 2963 903
rect 3757 897 3772 903
rect 4877 897 4892 903
rect 5188 897 5203 903
rect 5565 897 5580 903
rect 5588 897 5596 903
rect 6548 897 6563 903
rect 7597 897 7683 903
rect 7821 897 7892 903
rect 8308 897 8323 903
rect 9597 897 9660 903
rect 9876 897 9907 903
rect 68 837 83 843
rect 7386 836 7388 844
rect 8701 837 8716 843
rect 234 776 236 784
rect 669 777 684 783
rect 1604 776 1606 784
rect 2484 777 2499 783
rect 4724 777 4739 783
rect 5876 776 5880 784
rect 6268 777 6284 783
rect 68 717 83 723
rect 484 717 531 723
rect 1325 717 1340 723
rect 2413 717 2476 723
rect 2877 717 2892 723
rect 3741 717 3756 723
rect 4189 717 4204 723
rect 4877 717 4940 723
rect 5140 717 5203 723
rect 5565 717 5580 723
rect 5588 717 5654 723
rect 6029 717 6044 723
rect 6052 717 6115 723
rect 4436 697 4476 703
rect 8988 703 8996 714
rect 8932 697 8996 703
rect 2636 684 2644 690
rect 8028 684 8036 690
rect 9884 684 9892 690
rect 877 677 963 683
rect 1348 677 1395 683
rect 2884 677 2947 683
rect 4874 677 4963 683
rect 5636 677 5667 683
rect 6772 677 6803 683
rect 7828 677 7891 683
rect 8052 677 8115 683
rect 8893 677 8956 683
rect 9364 677 9416 683
rect 276 637 291 643
rect 724 637 739 643
rect 1172 637 1187 643
rect 2189 637 2204 643
rect 6292 637 6340 643
rect 6941 637 6956 643
rect 7165 637 7180 643
rect 7396 637 7443 643
rect 8500 637 8547 643
rect 8708 637 8758 643
rect 9146 636 9148 644
rect 9804 637 9820 643
rect 10248 637 10268 643
rect 445 577 476 583
rect 516 576 520 584
rect 1364 577 1427 583
rect 1588 577 1654 583
rect 2068 577 2099 583
rect 3828 577 3875 583
rect 4724 577 4787 583
rect 4948 577 5011 583
rect 6077 577 6092 583
rect 6760 577 6796 583
rect 8100 577 8148 583
rect 8324 577 8371 583
rect 9162 576 9164 584
rect 9188 577 9219 583
rect 9860 577 9876 583
rect 10248 576 10252 584
rect 692 557 739 563
rect 1140 557 1203 563
rect 5389 557 5452 563
rect 9396 557 9432 563
rect 3188 537 3203 543
rect 3341 537 3356 543
rect 3428 536 3430 544
rect 4276 537 4323 543
rect 4461 537 4540 543
rect 5149 537 5180 543
rect 5684 537 5716 543
rect 5708 530 5716 537
rect 9357 537 9372 543
rect 6396 530 6404 536
rect 6972 530 6980 536
rect 9804 530 9812 536
rect 7236 517 7284 523
rect 3580 506 3588 516
rect 7276 506 7284 517
rect 8300 506 8308 516
rect 221 497 268 503
rect 669 497 716 503
rect 877 497 892 503
rect 1117 497 1132 503
rect 1341 497 1372 503
rect 2252 497 2300 503
rect 2484 497 2547 503
rect 3117 497 3132 503
rect 3604 497 3651 503
rect 4028 497 4092 503
rect 4109 483 4115 503
rect 4548 497 4563 503
rect 4925 497 4940 503
rect 5188 497 5244 503
rect 5876 497 5939 503
rect 6310 497 6392 503
rect 6540 497 6611 503
rect 7501 483 7507 503
rect 7668 497 7715 503
rect 7853 497 7924 503
rect 8509 497 8579 503
rect 8788 497 8803 503
rect 8964 497 9011 503
rect 9581 497 9668 503
rect 4052 477 4115 483
rect 7434 477 7507 483
rect 8076 477 8124 483
rect 5546 376 5548 384
rect 5773 377 5788 383
rect 6220 337 6284 343
rect 205 317 220 323
rect 1530 316 1532 324
rect 2429 317 2444 323
rect 3741 317 3772 323
rect 4388 317 4396 323
rect 4850 317 4932 323
rect 5085 317 5171 323
rect 6244 317 6291 323
rect 8468 317 8484 323
rect 10173 317 10268 323
rect 1756 304 1764 314
rect 860 283 868 290
rect 860 277 892 283
rect 1516 283 1524 290
rect 2652 284 2660 290
rect 1516 277 1532 283
rect 2189 277 2280 283
rect 3124 277 3171 283
rect 3540 277 3603 283
rect 3740 277 3820 283
rect 4168 277 4243 283
rect 4420 277 4468 283
rect 5309 277 5388 283
rect 5628 283 5636 290
rect 7948 284 7956 290
rect 9740 284 9748 290
rect 5546 277 5636 283
rect 6676 277 6707 283
rect 7076 277 7155 283
rect 7524 277 7576 283
rect 8408 277 8499 283
rect 9082 277 9155 283
rect 9293 277 9308 283
rect 9965 277 10012 283
rect 708 237 723 243
rect 1364 237 1379 243
rect 1556 237 1606 243
rect 1978 236 1980 244
rect 2452 237 2515 243
rect 3380 236 3382 244
rect 5997 237 6028 243
rect 6429 237 6444 243
rect 6916 236 6918 244
rect 7748 237 7811 243
rect 8660 237 8710 243
rect 9364 236 9368 244
rect 9540 237 9603 243
rect 685 177 748 183
rect 1204 177 1235 183
rect 1613 177 1628 183
rect 1860 177 1923 183
rect 2301 177 2348 183
rect 4317 177 4364 183
rect 4556 177 4620 183
rect 5016 177 5036 183
rect 5706 177 5772 183
rect 7268 177 7299 183
rect 8301 177 8348 183
rect 8733 177 8780 183
rect 9389 177 9436 183
rect 1636 157 1686 163
rect 2548 157 2595 163
rect 3444 157 3478 163
rect 4781 157 4844 163
rect 6589 157 6636 163
rect 308 137 324 143
rect 316 130 324 137
rect 908 137 924 143
rect 908 130 916 137
rect 1460 137 1475 143
rect 2980 137 3059 143
rect 3405 137 3420 143
rect 3613 137 3692 143
rect 3876 137 3939 143
rect 4077 137 4092 143
rect 6157 137 6243 143
rect 7005 137 7052 143
rect 7213 137 7228 143
rect 7661 137 7692 143
rect 8077 137 8108 143
rect 8132 137 8163 143
rect 8356 137 8371 143
rect 9204 137 9251 143
rect 1004 130 1012 136
rect 4636 130 4644 136
rect 5788 130 5796 136
rect 68 117 84 123
rect 76 106 84 117
rect 1836 117 1900 123
rect 1836 106 1844 117
rect 7684 117 7720 123
rect 8956 117 8972 123
rect 8956 106 8964 117
rect 228 97 310 103
rect 460 97 547 103
rect 920 97 940 103
rect 460 96 468 97
rect 996 96 1000 104
rect 1148 97 1212 103
rect 1148 96 1156 97
rect 1373 97 1388 103
rect 2061 97 2076 103
rect 2525 97 2572 103
rect 3197 97 3219 103
rect 3213 83 3219 97
rect 4612 97 4632 103
rect 5245 97 5331 103
rect 6374 97 6451 103
rect 6797 97 6844 103
rect 7016 97 7084 103
rect 7229 97 7244 103
rect 7437 97 7516 103
rect 7869 97 7940 103
rect 8148 97 8163 103
rect 8509 97 8524 103
rect 8756 97 8812 103
rect 3213 77 3267 83
rect 5933 77 6012 83
<< m2contact >>
rect 1820 7576 1828 7584
rect 6092 7556 6100 7564
rect 316 7516 324 7524
rect 554 7516 562 7524
rect 924 7516 932 7524
rect 1116 7516 1124 7524
rect 1212 7516 1220 7524
rect 1452 7516 1460 7524
rect 2060 7516 2068 7524
rect 2284 7516 2292 7524
rect 2524 7516 2532 7524
rect 2716 7516 2724 7524
rect 2780 7516 2788 7524
rect 2796 7516 2804 7524
rect 3388 7516 3396 7524
rect 3612 7516 3620 7524
rect 3708 7516 3716 7524
rect 3916 7516 3924 7524
rect 3932 7516 3940 7524
rect 4300 7516 4308 7524
rect 4348 7516 4356 7524
rect 4604 7516 4612 7524
rect 5708 7536 5716 7544
rect 5852 7536 5860 7544
rect 5292 7516 5300 7524
rect 5500 7516 5508 7524
rect 5852 7516 5860 7524
rect 6188 7516 6196 7524
rect 6604 7516 6612 7524
rect 6796 7516 6804 7524
rect 7052 7516 7060 7524
rect 7068 7516 7076 7524
rect 7468 7516 7476 7524
rect 7548 7516 7556 7524
rect 7756 7516 7764 7524
rect 7980 7516 7988 7524
rect 8204 7516 8212 7524
rect 8412 7516 8420 7524
rect 8620 7516 8628 7524
rect 8764 7516 8772 7524
rect 8844 7516 8852 7524
rect 9244 7516 9252 7524
rect 9276 7516 9284 7524
rect 9484 7516 9492 7524
rect 9708 7516 9716 7524
rect 9916 7516 9924 7524
rect 76 7496 84 7504
rect 92 7476 100 7484
rect 316 7476 324 7484
rect 524 7476 532 7484
rect 556 7476 564 7484
rect 748 7476 756 7484
rect 908 7476 916 7484
rect 924 7476 932 7484
rect 1116 7476 1124 7484
rect 1228 7476 1236 7484
rect 1692 7476 1700 7484
rect 2028 7476 2036 7484
rect 2060 7476 2068 7484
rect 2268 7476 2276 7484
rect 2284 7476 2292 7484
rect 2492 7476 2500 7484
rect 2524 7476 2532 7484
rect 2716 7476 2724 7484
rect 2732 7476 2740 7484
rect 3036 7476 3044 7484
rect 3452 7476 3460 7484
rect 3708 7476 3716 7484
rect 3724 7476 3732 7484
rect 3740 7476 3748 7484
rect 3948 7476 3956 7484
rect 4140 7476 4148 7484
rect 4268 7476 4276 7484
rect 4380 7476 4388 7484
rect 4588 7476 4596 7484
rect 4604 7476 4612 7484
rect 4844 7476 4852 7484
rect 5084 7476 5092 7484
rect 5308 7476 5316 7484
rect 5852 7476 5860 7484
rect 5964 7476 5972 7484
rect 6188 7476 6196 7484
rect 6380 7476 6388 7484
rect 6652 7476 6660 7484
rect 6860 7476 6868 7484
rect 7100 7476 7108 7484
rect 7436 7476 7444 7484
rect 7532 7476 7540 7484
rect 7788 7476 7796 7484
rect 8204 7476 8212 7484
rect 8444 7476 8452 7484
rect 8748 7476 8756 7484
rect 8860 7476 8868 7484
rect 9180 7476 9188 7484
rect 9292 7476 9300 7484
rect 9500 7476 9508 7484
rect 9708 7476 9716 7484
rect 9932 7476 9940 7484
rect 1836 7456 1844 7464
rect 3854 7456 3862 7464
rect 300 7436 308 7444
rect 764 7436 772 7444
rect 3180 7436 3188 7444
rect 3228 7436 3236 7444
rect 3468 7436 3476 7444
rect 4092 7436 4100 7444
rect 5212 7436 5220 7444
rect 5660 7436 5668 7444
rect 6572 7436 6580 7444
rect 6780 7436 6788 7444
rect 7244 7436 7252 7444
rect 7308 7436 7316 7444
rect 7708 7436 7716 7444
rect 8140 7436 8148 7444
rect 8348 7436 8356 7444
rect 8572 7436 8580 7444
rect 8988 7436 8996 7444
rect 9036 7436 9044 7444
rect 9436 7436 9444 7444
rect 9628 7436 9636 7444
rect 9868 7436 9876 7444
rect 10060 7436 10068 7444
rect 60 7376 68 7384
rect 284 7376 292 7384
rect 508 7376 516 7384
rect 668 7376 676 7384
rect 940 7376 948 7384
rect 2236 7376 2244 7384
rect 2508 7376 2516 7384
rect 2956 7376 2964 7384
rect 3116 7376 3124 7384
rect 4300 7376 4308 7384
rect 4460 7376 4468 7384
rect 5132 7376 5140 7384
rect 5580 7376 5588 7384
rect 6028 7376 6036 7384
rect 6492 7376 6500 7384
rect 7180 7376 7188 7384
rect 7852 7376 7860 7384
rect 8060 7376 8068 7384
rect 8300 7376 8308 7384
rect 8732 7376 8740 7384
rect 10268 7376 10276 7384
rect 1340 7356 1348 7364
rect 1772 7356 1780 7364
rect 3836 7356 3844 7364
rect 4012 7356 4020 7364
rect 4732 7356 4740 7364
rect 6796 7356 6804 7364
rect 188 7336 196 7344
rect 428 7336 436 7344
rect 636 7336 644 7344
rect 876 7336 884 7344
rect 1084 7336 1092 7344
rect 1308 7336 1316 7344
rect 1580 7336 1588 7344
rect 1644 7336 1652 7344
rect 1868 7336 1876 7344
rect 2012 7336 2020 7344
rect 2428 7336 2436 7344
rect 2636 7336 2644 7344
rect 2748 7336 2756 7344
rect 3084 7336 3092 7344
rect 3324 7336 3332 7344
rect 3516 7336 3524 7344
rect 3644 7336 3652 7344
rect 3996 7336 4004 7344
rect 4204 7336 4212 7344
rect 4444 7336 4452 7344
rect 4652 7336 4660 7344
rect 4844 7336 4852 7344
rect 4956 7336 4964 7344
rect 5324 7336 5332 7344
rect 5548 7336 5556 7344
rect 5788 7336 5796 7344
rect 5900 7336 5908 7344
rect 6124 7336 6132 7344
rect 6316 7336 6324 7344
rect 6588 7336 6596 7344
rect 7036 7336 7044 7344
rect 7356 7336 7364 7344
rect 7468 7336 7476 7344
rect 7788 7336 7796 7344
rect 8044 7336 8052 7344
rect 8268 7336 8276 7344
rect 8492 7336 8500 7344
rect 8604 7336 8612 7344
rect 8828 7336 8836 7344
rect 9052 7336 9060 7344
rect 9260 7336 9268 7344
rect 9580 7336 9588 7344
rect 9708 7336 9716 7344
rect 9916 7336 9924 7344
rect 5164 7316 5172 7324
rect 268 7296 276 7304
rect 428 7296 436 7304
rect 652 7296 660 7304
rect 876 7296 884 7304
rect 1084 7296 1092 7304
rect 1324 7296 1332 7304
rect 1548 7296 1556 7304
rect 1628 7296 1636 7304
rect 1852 7296 1860 7304
rect 2012 7296 2020 7304
rect 2460 7296 2468 7304
rect 2652 7296 2660 7304
rect 2732 7296 2740 7304
rect 3100 7296 3108 7304
rect 3324 7296 3332 7304
rect 3532 7296 3540 7304
rect 3628 7296 3636 7304
rect 3980 7296 3988 7304
rect 4204 7296 4212 7304
rect 4444 7296 4452 7304
rect 4652 7296 4660 7304
rect 4876 7296 4884 7304
rect 4924 7296 4932 7304
rect 4972 7296 4980 7304
rect 5356 7296 5364 7304
rect 5580 7296 5588 7304
rect 5788 7296 5796 7304
rect 5852 7296 5860 7304
rect 6124 7296 6132 7304
rect 6348 7296 6356 7304
rect 6572 7296 6580 7304
rect 6812 7296 6820 7304
rect 7020 7296 7028 7304
rect 7372 7296 7380 7304
rect 7468 7296 7476 7304
rect 7836 7296 7844 7304
rect 8044 7296 8052 7304
rect 8268 7296 8276 7304
rect 8494 7296 8502 7304
rect 8588 7296 8596 7304
rect 9036 7296 9044 7304
rect 1982 7276 1990 7284
rect 9612 7296 9620 7304
rect 9692 7296 9700 7304
rect 9916 7296 9924 7304
rect 1180 7236 1188 7244
rect 2236 7236 2244 7244
rect 2908 7236 2916 7244
rect 3388 7236 3396 7244
rect 3774 7236 3782 7244
rect 5372 7236 5380 7244
rect 6268 7236 6276 7244
rect 6972 7236 6980 7244
rect 7180 7236 7188 7244
rect 7612 7236 7620 7244
rect 7676 7236 7684 7244
rect 8972 7236 8980 7244
rect 9420 7236 9428 7244
rect 9468 7236 9476 7244
rect 9852 7236 9860 7244
rect 7020 7176 7028 7184
rect 8092 7176 8100 7184
rect 268 7116 276 7124
rect 428 7116 436 7124
rect 684 7116 692 7124
rect 764 7116 772 7124
rect 1100 7116 1108 7124
rect 1132 7116 1140 7124
rect 1420 7116 1428 7124
rect 1644 7116 1652 7124
rect 940 7096 948 7104
rect 204 7076 212 7084
rect 652 7076 660 7084
rect 764 7076 772 7084
rect 1148 7076 1156 7084
rect 1212 7076 1220 7084
rect 1436 7076 1444 7084
rect 1996 7076 2004 7084
rect 2236 7116 2244 7124
rect 2332 7116 2340 7124
rect 2556 7116 2564 7124
rect 2780 7116 2788 7124
rect 3228 7116 3236 7124
rect 3692 7116 3700 7124
rect 4028 7116 4036 7124
rect 4252 7116 4260 7124
rect 4476 7116 4484 7124
rect 4540 7116 4548 7124
rect 4892 7116 4900 7124
rect 4988 7116 4996 7124
rect 5212 7116 5220 7124
rect 5788 7116 5796 7124
rect 6012 7116 6020 7124
rect 6124 7116 6132 7124
rect 6476 7116 6484 7124
rect 6572 7116 6580 7124
rect 6940 7116 6948 7124
rect 7164 7116 7172 7124
rect 7388 7116 7396 7124
rect 7484 7116 7492 7124
rect 7708 7116 7716 7124
rect 7948 7116 7956 7124
rect 8172 7116 8180 7124
rect 8396 7116 8404 7124
rect 8636 7116 8644 7124
rect 8860 7116 8868 7124
rect 9052 7116 9060 7124
rect 9212 7116 9220 7124
rect 9436 7116 9444 7124
rect 9644 7116 9652 7124
rect 9868 7116 9876 7124
rect 10076 7116 10084 7124
rect 6332 7096 6340 7104
rect 2252 7076 2260 7084
rect 2348 7076 2356 7084
rect 3020 7076 3028 7084
rect 3180 7076 3188 7084
rect 3468 7076 3476 7084
rect 3692 7076 3700 7084
rect 4012 7076 4020 7084
rect 4236 7076 4244 7084
rect 4316 7076 4324 7084
rect 4460 7076 4468 7084
rect 4540 7076 4548 7084
rect 4876 7076 4884 7084
rect 4988 7076 4996 7084
rect 5132 7076 5140 7084
rect 5228 7076 5236 7084
rect 5452 7076 5460 7084
rect 5788 7076 5796 7084
rect 5804 7076 5812 7084
rect 6012 7076 6020 7084
rect 6124 7076 6132 7084
rect 6460 7076 6468 7084
rect 6588 7076 6596 7084
rect 6956 7076 6964 7084
rect 7164 7076 7172 7084
rect 7244 7076 7252 7084
rect 7388 7076 7396 7084
rect 7468 7076 7476 7084
rect 7868 7076 7876 7084
rect 7964 7076 7972 7084
rect 8172 7076 8180 7084
rect 8412 7076 8420 7084
rect 8636 7076 8644 7084
rect 8876 7076 8884 7084
rect 9436 7076 9444 7084
rect 9628 7076 9636 7084
rect 10060 7076 10068 7084
rect 3868 7056 3876 7064
rect 4108 7056 4116 7064
rect 60 7036 68 7044
rect 284 7036 292 7044
rect 956 7036 964 7044
rect 1356 7036 1364 7044
rect 1788 7036 1796 7044
rect 1868 7036 1876 7044
rect 3148 7036 3156 7044
rect 3596 7036 3604 7044
rect 3884 7036 3892 7044
rect 4684 7036 4692 7044
rect 4748 7036 4756 7044
rect 5596 7036 5604 7044
rect 5644 7036 5652 7044
rect 6284 7036 6292 7044
rect 6780 7036 6788 7044
rect 6796 7036 6804 7044
rect 7852 7036 7860 7044
rect 8332 7036 8340 7044
rect 8556 7036 8564 7044
rect 8796 7036 8804 7044
rect 9068 7036 9076 7044
rect 9516 7036 9524 7044
rect 9676 7036 9684 7044
rect 268 6976 276 6984
rect 652 6976 660 6984
rect 1116 6976 1124 6984
rect 1404 6976 1412 6984
rect 2028 6976 2036 6984
rect 2252 6976 2260 6984
rect 2284 6976 2292 6984
rect 2460 6976 2468 6984
rect 3100 6976 3108 6984
rect 3164 6976 3172 6984
rect 3340 6976 3348 6984
rect 4444 6976 4452 6984
rect 6012 6976 6020 6984
rect 6460 6976 6468 6984
rect 6476 6976 6484 6984
rect 6924 6976 6932 6984
rect 7388 6976 7396 6984
rect 9132 6976 9140 6984
rect 10060 6976 10068 6984
rect 10236 6976 10244 6984
rect 668 6956 676 6964
rect 3788 6956 3796 6964
rect 4204 6956 4212 6964
rect 7596 6956 7604 6964
rect 8700 6956 8708 6964
rect 9644 6956 9652 6964
rect 204 6936 212 6944
rect 540 6936 548 6944
rect 876 6936 884 6944
rect 972 6936 980 6944
rect 1196 6936 1204 6944
rect 1324 6936 1332 6944
rect 1612 6936 1620 6944
rect 1644 6936 1652 6944
rect 1868 6936 1876 6944
rect 2092 6936 2100 6944
rect 2412 6936 2420 6944
rect 2652 6936 2660 6944
rect 2748 6936 2756 6944
rect 2972 6936 2980 6944
rect 3308 6936 3316 6944
rect 3532 6936 3540 6944
rect 3756 6936 3764 6944
rect 3980 6936 3988 6944
rect 4092 6936 4100 6944
rect 4412 6936 4420 6944
rect 4604 6936 4612 6944
rect 4828 6936 4836 6944
rect 5068 6936 5076 6944
rect 5196 6936 5204 6944
rect 5420 6936 5428 6944
rect 5644 6936 5652 6944
rect 5980 6936 5988 6944
rect 6220 6936 6228 6944
rect 6300 6936 6308 6944
rect 6668 6936 6676 6944
rect 6780 6936 6788 6944
rect 7004 6936 7012 6944
rect 7228 6936 7236 6944
rect 7580 6936 7588 6944
rect 7772 6936 7780 6944
rect 8012 6936 8020 6944
rect 8108 6936 8116 6944
rect 8332 6936 8340 6944
rect 8684 6936 8692 6944
rect 8860 6936 8868 6944
rect 8892 6936 8900 6944
rect 9100 6936 9108 6944
rect 9372 6936 9380 6944
rect 9452 6936 9460 6944
rect 9676 6936 9684 6944
rect 9884 6936 9892 6944
rect 10108 6936 10116 6944
rect 2940 6916 2948 6924
rect 268 6896 276 6904
rect 428 6896 436 6904
rect 508 6896 516 6904
rect 876 6896 884 6904
rect 972 6896 980 6904
rect 1180 6896 1188 6904
rect 1548 6896 1556 6904
rect 1628 6896 1636 6904
rect 2076 6896 2084 6904
rect 2428 6896 2436 6904
rect 2684 6896 2692 6904
rect 2732 6896 2740 6904
rect 2956 6896 2964 6904
rect 3308 6896 3316 6904
rect 3772 6896 3780 6904
rect 3980 6896 3988 6904
rect 4074 6896 4082 6904
rect 4412 6896 4420 6904
rect 4620 6896 4628 6904
rect 4876 6896 4884 6904
rect 5084 6896 5092 6904
rect 5180 6896 5188 6904
rect 5996 6896 6004 6904
rect 6220 6896 6228 6904
rect 6316 6896 6324 6904
rect 6684 6896 6692 6904
rect 6732 6896 6740 6904
rect 6988 6896 6996 6904
rect 7404 6896 7412 6904
rect 7564 6896 7572 6904
rect 8012 6896 8020 6904
rect 8108 6896 8116 6904
rect 8668 6896 8676 6904
rect 8892 6896 8900 6904
rect 9116 6896 9124 6904
rect 9340 6896 9348 6904
rect 9436 6896 9444 6904
rect 9660 6896 9668 6904
rect 10060 6896 10068 6904
rect 76 6836 84 6844
rect 1324 6836 1332 6844
rect 3164 6836 3172 6844
rect 4204 6836 4212 6844
rect 4268 6836 4276 6844
rect 4700 6836 4708 6844
rect 4940 6836 4948 6844
rect 5772 6836 5780 6844
rect 5852 6836 5860 6844
rect 8476 6836 8484 6844
rect 8508 6836 8516 6844
rect 972 6776 980 6784
rect 2572 6776 2580 6784
rect 6364 6776 6372 6784
rect 10060 6776 10068 6784
rect 10076 6776 10084 6784
rect 76 6716 84 6724
rect 316 6716 324 6724
rect 524 6716 532 6724
rect 1212 6716 1220 6724
rect 1436 6716 1444 6724
rect 1852 6716 1860 6724
rect 1900 6716 1908 6724
rect 2268 6716 2276 6724
rect 2364 6716 2372 6724
rect 2716 6716 2724 6724
rect 2940 6716 2948 6724
rect 3164 6716 3172 6724
rect 3244 6716 3252 6724
rect 3468 6716 3476 6724
rect 3820 6716 3828 6724
rect 4044 6716 4052 6724
rect 4268 6716 4276 6724
rect 4508 6716 4516 6724
rect 4588 6716 4596 6724
rect 4764 6716 4772 6724
rect 5036 6716 5044 6724
rect 5260 6716 5268 6724
rect 5628 6716 5636 6724
rect 5836 6716 5844 6724
rect 6092 6716 6100 6724
rect 6172 6716 6180 6724
rect 6844 6716 6852 6724
rect 7036 6716 7044 6724
rect 7292 6716 7300 6724
rect 7500 6716 7508 6724
rect 7708 6716 7716 6724
rect 7932 6716 7940 6724
rect 8284 6716 8292 6724
rect 8492 6716 8500 6724
rect 8572 6716 8580 6724
rect 8924 6716 8932 6724
rect 9004 6716 9012 6724
rect 9356 6716 9364 6724
rect 9564 6716 9572 6724
rect 9660 6716 9668 6724
rect 9868 6716 9876 6724
rect 9900 6716 9908 6724
rect 10252 6716 10260 6724
rect 1132 6696 1140 6704
rect 92 6676 100 6684
rect 300 6676 308 6684
rect 556 6676 564 6684
rect 764 6676 772 6684
rect 1116 6676 1124 6684
rect 1244 6676 1252 6684
rect 1804 6676 1812 6684
rect 1932 6676 1940 6684
rect 2076 6676 2084 6684
rect 2284 6676 2292 6684
rect 2380 6676 2388 6684
rect 2700 6676 2708 6684
rect 2940 6676 2948 6684
rect 2956 6676 2964 6684
rect 3132 6676 3140 6684
rect 3452 6676 3460 6684
rect 3484 6676 3492 6684
rect 4044 6676 4052 6684
rect 4268 6676 4276 6684
rect 4492 6676 4500 6684
rect 4588 6676 4596 6684
rect 5036 6676 5044 6684
rect 5276 6676 5284 6684
rect 5612 6676 5620 6684
rect 5820 6676 5828 6684
rect 5852 6676 5860 6684
rect 6060 6676 6068 6684
rect 6172 6676 6180 6684
rect 6332 6676 6340 6684
rect 6620 6676 6628 6684
rect 6828 6676 6836 6684
rect 7068 6676 7076 6684
rect 7292 6676 7300 6684
rect 7516 6676 7524 6684
rect 7724 6676 7732 6684
rect 7916 6676 7924 6684
rect 8092 6676 8100 6684
rect 8268 6676 8276 6684
rect 8284 6676 8292 6684
rect 8460 6676 8468 6684
rect 8572 6676 8580 6684
rect 8908 6676 8916 6684
rect 9020 6676 9028 6684
rect 9196 6676 9204 6684
rect 9340 6676 9348 6684
rect 9564 6676 9572 6684
rect 9676 6676 9684 6684
rect 9836 6676 9844 6684
rect 10236 6676 10244 6684
rect 7676 6656 7684 6664
rect 222 6636 230 6644
rect 476 6636 484 6644
rect 924 6636 932 6644
rect 1596 6636 1604 6644
rect 1644 6636 1652 6644
rect 2060 6636 2068 6644
rect 2508 6636 2516 6644
rect 2796 6636 2804 6644
rect 3628 6636 3636 6644
rect 3676 6636 3684 6644
rect 4060 6636 4068 6644
rect 4348 6636 4356 6644
rect 4940 6636 4948 6644
rect 5180 6636 5188 6644
rect 5420 6636 5428 6644
rect 5436 6636 5444 6644
rect 5692 6636 5700 6644
rect 6764 6636 6772 6644
rect 7020 6636 7028 6644
rect 7212 6636 7220 6644
rect 7436 6636 7444 6644
rect 7852 6636 7860 6644
rect 8092 6636 8100 6644
rect 8732 6636 8740 6644
rect 8778 6636 8786 6644
rect 9212 6636 9220 6644
rect 9388 6636 9396 6644
rect 10060 6636 10068 6644
rect 268 6576 276 6584
rect 668 6576 676 6584
rect 1100 6576 1108 6584
rect 1116 6576 1124 6584
rect 1388 6576 1396 6584
rect 1756 6576 1764 6584
rect 2060 6576 2068 6584
rect 2284 6576 2292 6584
rect 2492 6576 2500 6584
rect 2716 6576 2724 6584
rect 2892 6576 2900 6584
rect 3612 6576 3620 6584
rect 3820 6576 3828 6584
rect 4044 6576 4052 6584
rect 4252 6576 4260 6584
rect 5404 6576 5412 6584
rect 5628 6576 5636 6584
rect 6476 6576 6484 6584
rect 6748 6576 6756 6584
rect 7180 6576 7188 6584
rect 7676 6576 7684 6584
rect 7836 6576 7844 6584
rect 8060 6576 8068 6584
rect 8908 6576 8916 6584
rect 8924 6576 8932 6584
rect 9804 6576 9812 6584
rect 10252 6576 10260 6584
rect 206 6556 214 6564
rect 444 6556 452 6564
rect 4716 6556 4724 6564
rect 5116 6556 5124 6564
rect 6940 6556 6948 6564
rect 60 6536 68 6544
rect 428 6536 436 6544
rect 636 6536 644 6544
rect 876 6536 884 6544
rect 972 6536 980 6544
rect 1292 6536 1300 6544
rect 1516 6536 1524 6544
rect 1548 6536 1556 6544
rect 1628 6536 1636 6544
rect 1852 6536 1860 6544
rect 2044 6536 2052 6544
rect 2396 6536 2404 6544
rect 2620 6536 2628 6544
rect 2844 6536 2852 6544
rect 3084 6536 3092 6544
rect 3180 6536 3188 6544
rect 3420 6536 3428 6544
rect 3740 6536 3748 6544
rect 3964 6536 3972 6544
rect 4172 6536 4180 6544
rect 4380 6536 4388 6544
rect 4508 6536 4516 6544
rect 4828 6536 4836 6544
rect 5100 6536 5108 6544
rect 5292 6536 5300 6544
rect 5532 6536 5540 6544
rect 5788 6536 5796 6544
rect 5884 6536 5892 6544
rect 6108 6536 6116 6544
rect 6268 6536 6276 6544
rect 6572 6536 6580 6544
rect 6924 6536 6932 6544
rect 7132 6536 7140 6544
rect 7356 6536 7364 6544
rect 7596 6536 7604 6544
rect 7788 6536 7796 6544
rect 8028 6536 8036 6544
rect 8252 6536 8260 6544
rect 8268 6536 8276 6544
rect 8732 6536 8740 6544
rect 9116 6536 9124 6544
rect 9196 6536 9204 6544
rect 9564 6536 9572 6544
rect 9676 6536 9684 6544
rect 10012 6536 10020 6544
rect 10124 6536 10132 6544
rect 76 6496 84 6504
rect 412 6496 420 6504
rect 636 6496 644 6504
rect 876 6496 884 6504
rect 956 6496 964 6504
rect 1308 6496 1316 6504
rect 1532 6496 1540 6504
rect 1612 6496 1620 6504
rect 1852 6496 1860 6504
rect 2076 6496 2084 6504
rect 2428 6496 2436 6504
rect 2636 6496 2644 6504
rect 2860 6496 2868 6504
rect 3116 6496 3124 6504
rect 3180 6496 3188 6504
rect 3772 6496 3780 6504
rect 3964 6496 3972 6504
rect 4172 6496 4180 6504
rect 4396 6496 4404 6504
rect 4492 6496 4500 6504
rect 4892 6496 4900 6504
rect 5084 6496 5092 6504
rect 5324 6496 5332 6504
rect 5564 6496 5572 6504
rect 5772 6496 5780 6504
rect 5868 6496 5876 6504
rect 6076 6496 6084 6504
rect 6332 6496 6340 6504
rect 6572 6496 6580 6504
rect 6908 6496 6916 6504
rect 7164 6496 7172 6504
rect 7372 6496 7380 6504
rect 7596 6496 7604 6504
rect 7868 6496 7876 6504
rect 8044 6496 8052 6504
rect 8252 6496 8260 6504
rect 8348 6496 8356 6504
rect 8556 6496 8564 6504
rect 8764 6496 8772 6504
rect 9132 6496 9140 6504
rect 6092 6476 6100 6484
rect 9148 6476 9156 6484
rect 9612 6496 9620 6504
rect 9644 6496 9652 6504
rect 10012 6496 10020 6504
rect 10044 6496 10052 6504
rect 2236 6436 2244 6444
rect 3548 6436 3556 6444
rect 4636 6436 4644 6444
rect 4940 6436 4948 6444
rect 6012 6436 6020 6444
rect 6252 6436 6260 6444
rect 6764 6436 6772 6444
rect 7452 6436 7460 6444
rect 8732 6436 8740 6444
rect 9388 6436 9396 6444
rect 9420 6436 9428 6444
rect 9868 6436 9876 6444
rect 6284 6376 6292 6384
rect 9148 6376 9156 6384
rect 9644 6376 9652 6384
rect 4492 6336 4500 6344
rect 5212 6336 5220 6344
rect 92 6316 100 6324
rect 460 6316 468 6324
rect 668 6316 676 6324
rect 892 6316 900 6324
rect 1340 6316 1348 6324
rect 1420 6316 1428 6324
rect 1596 6316 1604 6324
rect 2252 6316 2260 6324
rect 2476 6316 2484 6324
rect 2764 6316 2772 6324
rect 2780 6316 2788 6324
rect 2940 6316 2948 6324
rect 3244 6316 3252 6324
rect 3596 6316 3604 6324
rect 3820 6316 3828 6324
rect 4044 6316 4052 6324
rect 4316 6316 4324 6324
rect 4492 6316 4500 6324
rect 4684 6316 4692 6324
rect 4910 6316 4918 6324
rect 4972 6316 4980 6324
rect 5372 6316 5380 6324
rect 5452 6316 5460 6324
rect 5820 6316 5828 6324
rect 5900 6316 5908 6324
rect 6124 6316 6132 6324
rect 6364 6316 6372 6324
rect 6588 6316 6596 6324
rect 6812 6316 6820 6324
rect 7036 6316 7044 6324
rect 7852 6316 7860 6324
rect 8060 6316 8068 6324
rect 8252 6316 8260 6324
rect 8316 6316 8324 6324
rect 8476 6316 8484 6324
rect 8556 6316 8564 6324
rect 8908 6316 8916 6324
rect 8940 6316 8948 6324
rect 8988 6316 8996 6324
rect 9356 6316 9364 6324
rect 9436 6316 9444 6324
rect 9788 6316 9796 6324
rect 10060 6316 10068 6324
rect 10222 6316 10230 6324
rect 92 6276 100 6284
rect 444 6276 452 6284
rect 652 6276 660 6284
rect 1116 6276 1124 6284
rect 1324 6276 1332 6284
rect 1436 6276 1444 6284
rect 1660 6276 1668 6284
rect 1884 6276 1892 6284
rect 2236 6276 2244 6284
rect 2460 6276 2468 6284
rect 2700 6276 2708 6284
rect 2796 6276 2804 6284
rect 2924 6276 2932 6284
rect 3020 6276 3028 6284
rect 3564 6276 3572 6284
rect 3804 6276 3812 6284
rect 4044 6276 4052 6284
rect 4236 6276 4244 6284
rect 4476 6276 4484 6284
rect 4684 6276 4692 6284
rect 4908 6276 4916 6284
rect 4956 6276 4964 6284
rect 5372 6276 5380 6284
rect 5484 6276 5492 6284
rect 5804 6276 5812 6284
rect 5916 6276 5924 6284
rect 6140 6276 6148 6284
rect 6364 6276 6372 6284
rect 6604 6276 6612 6284
rect 6764 6276 6772 6284
rect 7020 6276 7028 6284
rect 7052 6276 7060 6284
rect 7276 6276 7284 6284
rect 7500 6276 7508 6284
rect 7804 6276 7812 6284
rect 8028 6276 8036 6284
rect 8252 6276 8260 6284
rect 8444 6276 8452 6284
rect 8572 6276 8580 6284
rect 8908 6276 8916 6284
rect 9020 6276 9028 6284
rect 9164 6276 9172 6284
rect 9356 6276 9364 6284
rect 9468 6276 9476 6284
rect 9596 6276 9604 6284
rect 9788 6276 9796 6284
rect 10012 6276 10020 6284
rect 10220 6276 10228 6284
rect 524 6256 532 6264
rect 2044 6256 2052 6264
rect 3450 6256 3458 6264
rect 5180 6256 5188 6264
rect 6780 6256 6788 6264
rect 236 6236 244 6244
rect 252 6236 260 6244
rect 716 6236 724 6244
rect 1564 6236 1572 6244
rect 2014 6236 2022 6244
rect 2332 6236 2340 6244
rect 2508 6236 2516 6244
rect 3388 6236 3396 6244
rect 3612 6236 3620 6244
rect 3836 6236 3844 6244
rect 4124 6236 4132 6244
rect 4332 6236 4340 6244
rect 4732 6236 4740 6244
rect 5598 6236 5606 6244
rect 5676 6236 5684 6244
rect 6044 6236 6052 6244
rect 6524 6236 6532 6244
rect 7180 6236 7188 6244
rect 7628 6236 7636 6244
rect 7644 6236 7652 6244
rect 7884 6236 7892 6244
rect 8076 6236 8084 6244
rect 8700 6236 8708 6244
rect 8716 6236 8724 6244
rect 9596 6236 9604 6244
rect 9820 6236 9828 6244
rect 10076 6236 10084 6244
rect 76 6176 84 6184
rect 236 6176 244 6184
rect 940 6176 948 6184
rect 1164 6176 1172 6184
rect 1324 6176 1332 6184
rect 1548 6176 1556 6184
rect 1836 6176 1844 6184
rect 1996 6176 2004 6184
rect 2444 6176 2452 6184
rect 2684 6176 2692 6184
rect 2716 6176 2724 6184
rect 3418 6176 3426 6184
rect 3580 6176 3588 6184
rect 4524 6176 4532 6184
rect 4700 6176 4708 6184
rect 4908 6176 4916 6184
rect 5212 6176 5220 6184
rect 5372 6176 5380 6184
rect 5804 6176 5812 6184
rect 6748 6176 6756 6184
rect 7404 6176 7412 6184
rect 8252 6176 8260 6184
rect 8460 6176 8468 6184
rect 8684 6176 8692 6184
rect 8762 6176 8770 6184
rect 9164 6176 9172 6184
rect 9644 6176 9652 6184
rect 10028 6176 10036 6184
rect 10044 6176 10052 6184
rect 3116 6156 3124 6164
rect 5820 6156 5828 6164
rect 6028 6156 6036 6164
rect 204 6136 212 6144
rect 492 6136 500 6144
rect 652 6136 660 6144
rect 876 6136 884 6144
rect 1084 6136 1092 6144
rect 1292 6136 1300 6144
rect 1596 6136 1604 6144
rect 1756 6136 1764 6144
rect 1964 6136 1972 6144
rect 2204 6136 2212 6144
rect 2316 6136 2324 6144
rect 2492 6136 2500 6144
rect 2844 6136 2852 6144
rect 3084 6136 3092 6144
rect 3388 6136 3396 6144
rect 3548 6136 3556 6144
rect 3756 6136 3764 6144
rect 3852 6136 3860 6144
rect 3996 6136 4004 6144
rect 4220 6136 4228 6144
rect 4316 6136 4324 6144
rect 4572 6136 4580 6144
rect 4780 6136 4788 6144
rect 4988 6136 4996 6144
rect 5244 6136 5252 6144
rect 5436 6136 5444 6144
rect 5596 6136 5604 6144
rect 5660 6136 5668 6144
rect 5996 6136 6004 6144
rect 6236 6136 6244 6144
rect 6332 6136 6340 6144
rect 6572 6136 6580 6144
rect 6924 6136 6932 6144
rect 7148 6136 7156 6144
rect 7244 6136 7252 6144
rect 7420 6136 7428 6144
rect 7628 6136 7636 6144
rect 7676 6136 7684 6144
rect 8012 6136 8020 6144
rect 8108 6136 8116 6144
rect 8332 6136 8340 6144
rect 8556 6136 8564 6144
rect 8892 6136 8900 6144
rect 9004 6136 9012 6144
rect 9340 6136 9348 6144
rect 9532 6136 9540 6144
rect 9836 6136 9844 6144
rect 9852 6136 9860 6144
rect 9884 6136 9892 6144
rect 10204 6136 10212 6144
rect 252 6096 260 6104
rect 460 6096 468 6104
rect 652 6096 660 6104
rect 876 6096 884 6104
rect 1084 6096 1092 6104
rect 1308 6096 1316 6104
rect 1532 6096 1540 6104
rect 1772 6096 1780 6104
rect 1980 6096 1988 6104
rect 2204 6096 2212 6104
rect 2300 6096 2308 6104
rect 2524 6096 2532 6104
rect 2860 6096 2868 6104
rect 2892 6096 2900 6104
rect 3100 6096 3108 6104
rect 3324 6096 3332 6104
rect 3564 6096 3572 6104
rect 3772 6096 3780 6104
rect 4012 6096 4020 6104
rect 4300 6096 4308 6104
rect 524 6076 532 6084
rect 4252 6076 4260 6084
rect 4540 6096 4548 6104
rect 4764 6096 4772 6104
rect 5004 6096 5012 6104
rect 5228 6096 5236 6104
rect 5580 6096 5588 6104
rect 5660 6096 5668 6104
rect 6012 6096 6020 6104
rect 6236 6096 6244 6104
rect 6332 6096 6340 6104
rect 6556 6096 6564 6104
rect 6924 6096 6932 6104
rect 7148 6096 7156 6104
rect 7228 6096 7236 6104
rect 7580 6096 7588 6104
rect 7674 6096 7682 6104
rect 8012 6096 8020 6104
rect 8108 6096 8116 6104
rect 8332 6096 8340 6104
rect 8540 6096 8548 6104
rect 8892 6096 8900 6104
rect 9004 6096 9012 6104
rect 9340 6096 9348 6104
rect 9580 6096 9588 6104
rect 9804 6096 9812 6104
rect 9884 6096 9892 6104
rect 10222 6096 10230 6104
rect 9180 6076 9188 6084
rect 6780 6056 6788 6064
rect 732 6036 740 6044
rect 4092 6036 4100 6044
rect 6476 6036 6484 6044
rect 7820 6036 7828 6044
rect 7852 6036 7860 6044
rect 9420 6036 9428 6044
rect 5258 5976 5266 5984
rect 5630 5976 5638 5984
rect 8332 5976 8340 5984
rect 220 5916 228 5924
rect 460 5916 468 5924
rect 700 5916 708 5924
rect 764 5916 772 5924
rect 1116 5916 1124 5924
rect 1372 5916 1380 5924
rect 1580 5916 1588 5924
rect 1804 5916 1812 5924
rect 2060 5916 2068 5924
rect 2268 5916 2276 5924
rect 2508 5916 2516 5924
rect 2716 5916 2724 5924
rect 2924 5916 2932 5924
rect 2988 5916 2996 5924
rect 3356 5916 3364 5924
rect 3596 5916 3604 5924
rect 3804 5916 3812 5924
rect 4044 5916 4052 5924
rect 4252 5916 4260 5924
rect 4476 5916 4484 5924
rect 4940 5916 4948 5924
rect 5036 5916 5044 5924
rect 5404 5916 5412 5924
rect 5500 5916 5508 5924
rect 5724 5916 5732 5924
rect 6076 5916 6084 5924
rect 6316 5916 6324 5924
rect 6556 5916 6564 5924
rect 6796 5916 6804 5924
rect 6860 5916 6868 5924
rect 7020 5916 7028 5924
rect 7516 5916 7524 5924
rect 7948 5916 7956 5924
rect 8524 5916 8532 5924
rect 8604 5916 8612 5924
rect 8988 5916 8996 5924
rect 9036 5916 9044 5924
rect 9260 5916 9268 5924
rect 9420 5916 9428 5924
rect 9692 5916 9700 5924
rect 204 5876 212 5884
rect 444 5876 452 5884
rect 460 5876 468 5884
rect 668 5876 676 5884
rect 780 5876 788 5884
rect 1116 5876 1124 5884
rect 1340 5876 1348 5884
rect 1628 5876 1636 5884
rect 1804 5876 1812 5884
rect 2028 5876 2036 5884
rect 2060 5876 2068 5884
rect 2284 5876 2292 5884
rect 2492 5876 2500 5884
rect 2700 5876 2708 5884
rect 2908 5876 2916 5884
rect 3020 5876 3028 5884
rect 3356 5876 3364 5884
rect 3580 5876 3588 5884
rect 3788 5876 3796 5884
rect 4028 5876 4036 5884
rect 4236 5876 4244 5884
rect 4476 5876 4484 5884
rect 4492 5876 4500 5884
rect 4700 5876 4708 5884
rect 8796 5896 8804 5904
rect 4908 5876 4916 5884
rect 5372 5876 5380 5884
rect 5500 5876 5508 5884
rect 5724 5876 5732 5884
rect 6076 5876 6084 5884
rect 6316 5876 6324 5884
rect 6540 5876 6548 5884
rect 6764 5876 6772 5884
rect 6844 5876 6852 5884
rect 7084 5876 7092 5884
rect 7308 5876 7316 5884
rect 7740 5876 7748 5884
rect 8156 5876 8164 5884
rect 8508 5876 8516 5884
rect 8604 5876 8612 5884
rect 8956 5876 8964 5884
rect 9020 5876 9028 5884
rect 9244 5876 9252 5884
rect 9260 5876 9268 5884
rect 9484 5876 9492 5884
rect 9676 5876 9684 5884
rect 9692 5876 9700 5884
rect 9900 5876 9908 5884
rect 1388 5856 1396 5864
rect 1596 5856 1604 5864
rect 6332 5856 6340 5864
rect 76 5836 84 5844
rect 300 5836 308 5844
rect 924 5836 932 5844
rect 972 5836 980 5844
rect 1900 5836 1908 5844
rect 2332 5836 2340 5844
rect 2572 5836 2580 5844
rect 2780 5836 2788 5844
rect 3148 5836 3156 5844
rect 3212 5836 3220 5844
rect 3436 5836 3444 5844
rect 3644 5836 3652 5844
rect 3884 5836 3892 5844
rect 4108 5836 4116 5844
rect 4284 5836 4292 5844
rect 5180 5836 5188 5844
rect 5884 5836 5892 5844
rect 5932 5836 5940 5844
rect 6156 5836 6164 5844
rect 6572 5836 6580 5844
rect 7020 5836 7028 5844
rect 8300 5836 8308 5844
rect 8348 5836 8356 5844
rect 8780 5836 8788 5844
rect 9420 5836 9428 5844
rect 10044 5836 10052 5844
rect 684 5776 692 5784
rect 876 5776 884 5784
rect 1404 5776 1412 5784
rect 2268 5776 2276 5784
rect 2716 5776 2724 5784
rect 3180 5776 3188 5784
rect 3450 5776 3458 5784
rect 3660 5776 3668 5784
rect 4044 5776 4052 5784
rect 4492 5776 4500 5784
rect 4716 5776 4724 5784
rect 4924 5776 4932 5784
rect 4988 5776 4996 5784
rect 5388 5776 5396 5784
rect 5660 5776 5668 5784
rect 6812 5776 6820 5784
rect 6972 5776 6980 5784
rect 7196 5776 7204 5784
rect 7420 5776 7428 5784
rect 7692 5776 7700 5784
rect 7932 5776 7940 5784
rect 8316 5776 8324 5784
rect 8364 5776 8372 5784
rect 8572 5776 8580 5784
rect 9164 5776 9172 5784
rect 9180 5776 9188 5784
rect 9836 5776 9844 5784
rect 10044 5776 10052 5784
rect 2748 5756 2756 5764
rect 188 5736 196 5744
rect 412 5736 420 5744
rect 508 5736 516 5744
rect 732 5736 740 5744
rect 1068 5736 1076 5744
rect 1100 5736 1108 5744
rect 1196 5736 1204 5744
rect 1420 5736 1428 5744
rect 1628 5736 1636 5744
rect 1660 5736 1668 5744
rect 1884 5736 1892 5744
rect 2348 5736 2356 5744
rect 2908 5736 2916 5744
rect 3020 5736 3028 5744
rect 3372 5736 3380 5744
rect 3580 5736 3588 5744
rect 3788 5736 3796 5744
rect 3900 5736 3908 5744
rect 4108 5736 4116 5744
rect 4220 5736 4228 5744
rect 4364 5736 4372 5744
rect 4572 5736 4580 5744
rect 4796 5736 4804 5744
rect 5180 5736 5188 5744
rect 5244 5736 5252 5744
rect 5468 5736 5476 5744
rect 5692 5736 5700 5744
rect 5932 5736 5940 5744
rect 6156 5736 6164 5744
rect 6492 5736 6500 5744
rect 6604 5736 6612 5744
rect 6828 5736 6836 5744
rect 7020 5736 7028 5744
rect 7276 5736 7284 5744
rect 7500 5736 7508 5744
rect 7740 5736 7748 5744
rect 7916 5736 7924 5744
rect 8060 5736 8068 5744
rect 8156 5736 8164 5744
rect 8492 5736 8500 5744
rect 8700 5736 8708 5744
rect 8812 5736 8820 5744
rect 9036 5736 9044 5744
rect 9372 5736 9380 5744
rect 9484 5736 9492 5744
rect 9708 5736 9716 5744
rect 9900 5736 9908 5744
rect 700 5716 708 5724
rect 3180 5716 3188 5724
rect 204 5696 212 5704
rect 412 5696 420 5704
rect 492 5696 500 5704
rect 1084 5696 1092 5704
rect 1116 5696 1124 5704
rect 1420 5696 1428 5704
rect 1644 5696 1652 5704
rect 1884 5696 1892 5704
rect 2108 5696 2116 5704
rect 2332 5696 2340 5704
rect 2556 5696 2564 5704
rect 2940 5696 2948 5704
rect 3004 5696 3012 5704
rect 3388 5696 3396 5704
rect 3596 5696 3604 5704
rect 3884 5696 3892 5704
rect 4252 5696 4260 5704
rect 4348 5696 4356 5704
rect 4572 5696 4580 5704
rect 4780 5696 4788 5704
rect 5132 5696 5140 5704
rect 5164 5696 5172 5704
rect 5388 5696 5396 5704
rect 5692 5696 5700 5704
rect 5900 5696 5908 5704
rect 5916 5696 5924 5704
rect 6108 5696 6116 5704
rect 6492 5696 6500 5704
rect 6588 5696 6596 5704
rect 6828 5696 6836 5704
rect 7004 5696 7012 5704
rect 7276 5696 7284 5704
rect 7500 5696 7508 5704
rect 7724 5696 7732 5704
rect 8092 5696 8100 5704
rect 8140 5696 8148 5704
rect 8508 5696 8516 5704
rect 8780 5696 8788 5704
rect 9004 5696 9012 5704
rect 9372 5696 9380 5704
rect 9468 5696 9476 5704
rect 9692 5696 9700 5704
rect 9884 5696 9892 5704
rect 8780 5676 8788 5684
rect 9692 5676 9700 5684
rect 940 5656 948 5664
rect 60 5636 68 5644
rect 268 5636 276 5644
rect 1788 5636 1796 5644
rect 2700 5636 2708 5644
rect 3228 5636 3236 5644
rect 4924 5636 4932 5644
rect 5404 5636 5412 5644
rect 6060 5636 6068 5644
rect 6284 5636 6292 5644
rect 6348 5636 6356 5644
rect 6748 5636 6756 5644
rect 8956 5636 8964 5644
rect 4332 5576 4340 5584
rect 8332 5576 8340 5584
rect 9036 5576 9044 5584
rect 1674 5556 1682 5564
rect 8092 5556 8100 5564
rect 6524 5536 6532 5544
rect 220 5516 228 5524
rect 460 5516 468 5524
rect 684 5516 692 5524
rect 908 5516 916 5524
rect 988 5516 996 5524
rect 1372 5516 1380 5524
rect 1580 5516 1588 5524
rect 1804 5516 1812 5524
rect 2044 5516 2052 5524
rect 2140 5516 2148 5524
rect 2524 5516 2532 5524
rect 2748 5516 2756 5524
rect 2940 5516 2948 5524
rect 3164 5516 3172 5524
rect 3388 5516 3396 5524
rect 3468 5516 3476 5524
rect 3820 5516 3828 5524
rect 3916 5516 3924 5524
rect 4268 5516 4276 5524
rect 4492 5516 4500 5524
rect 4588 5516 4596 5524
rect 4812 5516 4820 5524
rect 5180 5516 5188 5524
rect 5404 5516 5412 5524
rect 5420 5516 5428 5524
rect 5724 5516 5732 5524
rect 6076 5516 6084 5524
rect 6300 5516 6308 5524
rect 6364 5516 6372 5524
rect 6748 5516 6756 5524
rect 6812 5516 6820 5524
rect 7020 5516 7028 5524
rect 7404 5516 7412 5524
rect 7500 5516 7508 5524
rect 7708 5516 7716 5524
rect 7932 5516 7940 5524
rect 8172 5516 8180 5524
rect 8348 5516 8356 5524
rect 8732 5516 8740 5524
rect 8956 5516 8964 5524
rect 9196 5516 9204 5524
rect 9404 5516 9412 5524
rect 9420 5516 9428 5524
rect 9628 5516 9636 5524
rect 9836 5516 9844 5524
rect 10060 5516 10068 5524
rect 1836 5496 1844 5504
rect 3180 5496 3188 5504
rect 204 5476 212 5484
rect 444 5476 452 5484
rect 460 5476 468 5484
rect 668 5476 676 5484
rect 908 5476 916 5484
rect 1004 5476 1012 5484
rect 1148 5476 1156 5484
rect 1340 5476 1348 5484
rect 1372 5476 1380 5484
rect 1596 5476 1604 5484
rect 1836 5476 1844 5484
rect 2028 5476 2036 5484
rect 2076 5476 2084 5484
rect 2492 5476 2500 5484
rect 2524 5476 2532 5484
rect 2748 5476 2756 5484
rect 2956 5476 2964 5484
rect 3148 5476 3156 5484
rect 3404 5476 3412 5484
rect 3484 5476 3492 5484
rect 3804 5476 3812 5484
rect 3916 5476 3924 5484
rect 4252 5476 4260 5484
rect 4508 5476 4516 5484
rect 4588 5476 4596 5484
rect 4828 5476 4836 5484
rect 5180 5476 5188 5484
rect 5388 5476 5396 5484
rect 5500 5476 5508 5484
rect 5708 5476 5716 5484
rect 5724 5476 5732 5484
rect 6060 5476 6068 5484
rect 6284 5476 6292 5484
rect 6332 5476 6340 5484
rect 6716 5476 6724 5484
rect 6748 5476 6756 5484
rect 7020 5476 7028 5484
rect 7052 5476 7060 5484
rect 7388 5476 7396 5484
rect 7500 5476 7508 5484
rect 7724 5476 7732 5484
rect 7948 5476 7956 5484
rect 8172 5476 8180 5484
rect 8412 5476 8420 5484
rect 8716 5476 8724 5484
rect 8956 5476 8964 5484
rect 9404 5476 9412 5484
rect 9820 5476 9828 5484
rect 9852 5476 9860 5484
rect 10028 5476 10036 5484
rect 5258 5456 5266 5464
rect 7692 5456 7700 5464
rect 8764 5456 8772 5464
rect 60 5436 68 5444
rect 300 5436 308 5444
rect 700 5436 708 5444
rect 1148 5436 1156 5444
rect 2300 5436 2308 5444
rect 2348 5436 2356 5444
rect 3020 5436 3028 5444
rect 3612 5436 3620 5444
rect 3676 5436 3684 5444
rect 4060 5436 4068 5444
rect 4124 5436 4132 5444
rect 4748 5436 4756 5444
rect 4972 5436 4980 5444
rect 5036 5436 5044 5444
rect 5868 5436 5876 5444
rect 5932 5436 5940 5444
rect 6124 5436 6132 5444
rect 6524 5436 6532 5444
rect 7196 5436 7204 5444
rect 7260 5436 7268 5444
rect 7852 5436 7860 5444
rect 8524 5436 8532 5444
rect 8556 5436 8564 5444
rect 9036 5436 9044 5444
rect 9468 5436 9476 5444
rect 988 5376 996 5384
rect 1612 5376 1620 5384
rect 2060 5376 2068 5384
rect 2508 5376 2516 5384
rect 2524 5376 2532 5384
rect 3004 5376 3012 5384
rect 3900 5376 3908 5384
rect 5100 5376 5108 5384
rect 5500 5376 5508 5384
rect 6236 5376 6244 5384
rect 6620 5376 6628 5384
rect 6844 5376 6852 5384
rect 6876 5376 6884 5384
rect 7372 5376 7380 5384
rect 8060 5376 8068 5384
rect 8460 5376 8468 5384
rect 8892 5376 8900 5384
rect 8940 5376 8948 5384
rect 9326 5376 9334 5384
rect 10060 5376 10068 5384
rect 524 5356 532 5364
rect 1836 5356 1844 5364
rect 3436 5356 3444 5364
rect 4364 5356 4372 5364
rect 204 5336 212 5344
rect 316 5336 324 5344
rect 668 5336 676 5344
rect 908 5336 916 5344
rect 1132 5336 1140 5344
rect 1356 5336 1364 5344
rect 1436 5336 1444 5344
rect 1580 5336 1588 5344
rect 1804 5336 1812 5344
rect 2028 5336 2036 5344
rect 2268 5336 2276 5344
rect 2380 5336 2388 5344
rect 2732 5336 2740 5344
rect 2828 5336 2836 5344
rect 2972 5336 2980 5344
rect 3180 5336 3188 5344
rect 3420 5336 3428 5344
rect 3644 5336 3652 5344
rect 3868 5336 3876 5344
rect 4108 5336 4116 5344
rect 4220 5336 4228 5344
rect 6012 5356 6020 5364
rect 7324 5356 7332 5364
rect 8284 5356 8292 5364
rect 9644 5356 9652 5364
rect 10236 5356 10244 5364
rect 4796 5336 4804 5344
rect 4860 5336 4868 5344
rect 4988 5336 4996 5344
rect 5228 5336 5236 5344
rect 5356 5336 5364 5344
rect 5692 5336 5700 5344
rect 5900 5336 5908 5344
rect 6124 5336 6132 5344
rect 6380 5336 6388 5344
rect 6476 5336 6484 5344
rect 6716 5336 6724 5344
rect 7068 5336 7076 5344
rect 7180 5336 7188 5344
rect 7516 5336 7524 5344
rect 7628 5336 7636 5344
rect 7868 5336 7876 5344
rect 8188 5336 8196 5344
rect 8428 5336 8436 5344
rect 8652 5336 8660 5344
rect 8732 5336 8740 5344
rect 9068 5336 9076 5344
rect 9196 5336 9204 5344
rect 9548 5336 9556 5344
rect 9772 5336 9780 5344
rect 9868 5336 9876 5344
rect 10028 5336 10036 5344
rect 1148 5316 1156 5324
rect 284 5296 292 5304
rect 316 5296 324 5304
rect 908 5296 916 5304
rect 1372 5296 1380 5304
rect 1580 5296 1588 5304
rect 1852 5296 1860 5304
rect 2060 5296 2068 5304
rect 2268 5296 2276 5304
rect 2348 5296 2356 5304
rect 2732 5296 2740 5304
rect 2828 5296 2836 5304
rect 3196 5296 3204 5304
rect 3420 5296 3428 5304
rect 3948 5296 3956 5304
rect 4108 5296 4116 5304
rect 4204 5296 4212 5304
rect 4412 5296 4420 5304
rect 4572 5296 4580 5304
rect 4796 5296 4804 5304
rect 5020 5296 5028 5304
rect 5244 5296 5252 5304
rect 5340 5296 5348 5304
rect 5484 5296 5492 5304
rect 5708 5296 5716 5304
rect 5916 5296 5924 5304
rect 6140 5296 6148 5304
rect 6380 5296 6388 5304
rect 6476 5296 6484 5304
rect 6700 5296 6708 5304
rect 7068 5296 7076 5304
rect 7148 5296 7156 5304
rect 7532 5296 7540 5304
rect 7628 5296 7636 5304
rect 8204 5296 8212 5304
rect 8428 5296 8436 5304
rect 8654 5296 8662 5304
rect 8748 5296 8756 5304
rect 9084 5296 9092 5304
rect 9180 5296 9188 5304
rect 9548 5296 9556 5304
rect 9772 5296 9780 5304
rect 9868 5296 9876 5304
rect 10092 5296 10100 5304
rect 8044 5276 8052 5284
rect 76 5236 84 5244
rect 460 5236 468 5244
rect 1228 5236 1236 5244
rect 3260 5236 3268 5244
rect 5724 5236 5732 5244
rect 6908 5236 6916 5244
rect 7308 5236 7316 5244
rect 7772 5236 7780 5244
rect 8524 5236 8532 5244
rect 9404 5236 9412 5244
rect 1580 5176 1588 5184
rect 4124 5176 4132 5184
rect 6332 5176 6340 5184
rect 7708 5176 7716 5184
rect 60 5116 68 5124
rect 444 5116 452 5124
rect 668 5116 676 5124
rect 892 5116 900 5124
rect 972 5116 980 5124
rect 1212 5116 1220 5124
rect 1644 5116 1652 5124
rect 2044 5116 2052 5124
rect 2124 5116 2132 5124
rect 2476 5116 2484 5124
rect 2716 5116 2724 5124
rect 2940 5116 2948 5124
rect 3212 5116 3220 5124
rect 3244 5116 3252 5124
rect 3612 5116 3620 5124
rect 3692 5116 3700 5124
rect 3932 5116 3940 5124
rect 4300 5116 4308 5124
rect 4748 5116 4756 5124
rect 4988 5116 4996 5124
rect 5196 5116 5204 5124
rect 5276 5116 5284 5124
rect 5660 5116 5668 5124
rect 5868 5116 5876 5124
rect 5948 5116 5956 5124
rect 6188 5116 6196 5124
rect 6556 5116 6564 5124
rect 6652 5116 6660 5124
rect 7004 5116 7012 5124
rect 7212 5116 7220 5124
rect 7436 5116 7444 5124
rect 7516 5116 7524 5124
rect 7868 5116 7876 5124
rect 7964 5116 7972 5124
rect 8188 5116 8196 5124
rect 8540 5116 8548 5124
rect 8748 5116 8756 5124
rect 8828 5116 8836 5124
rect 9036 5116 9044 5124
rect 9388 5116 9396 5124
rect 9468 5116 9476 5124
rect 9692 5116 9700 5124
rect 10044 5116 10052 5124
rect 1884 5096 1892 5104
rect 4396 5096 4404 5104
rect 5500 5096 5508 5104
rect 92 5076 100 5084
rect 252 5076 260 5084
rect 444 5076 452 5084
rect 652 5076 660 5084
rect 892 5076 900 5084
rect 988 5076 996 5084
rect 1212 5076 1220 5084
rect 1372 5076 1380 5084
rect 1676 5076 1684 5084
rect 2012 5076 2020 5084
rect 2124 5076 2132 5084
rect 2476 5076 2484 5084
rect 2508 5076 2516 5084
rect 2796 5076 2804 5084
rect 2940 5076 2948 5084
rect 2956 5076 2964 5084
rect 3148 5076 3156 5084
rect 3260 5076 3268 5084
rect 3612 5076 3620 5084
rect 3724 5076 3732 5084
rect 3948 5076 3956 5084
rect 4172 5076 4180 5084
rect 4300 5076 4308 5084
rect 4412 5076 4420 5084
rect 4572 5076 4580 5084
rect 4764 5076 4772 5084
rect 5196 5076 5204 5084
rect 5308 5076 5316 5084
rect 5628 5076 5636 5084
rect 5884 5076 5892 5084
rect 5900 5076 5908 5084
rect 6188 5076 6196 5084
rect 6540 5076 6548 5084
rect 6652 5076 6660 5084
rect 6844 5076 6852 5084
rect 7004 5076 7012 5084
rect 7212 5076 7220 5084
rect 7404 5076 7412 5084
rect 7500 5076 7508 5084
rect 7868 5076 7876 5084
rect 7980 5076 7988 5084
rect 8204 5076 8212 5084
rect 8524 5076 8532 5084
rect 8748 5076 8756 5084
rect 8844 5076 8852 5084
rect 9052 5076 9060 5084
rect 9388 5076 9396 5084
rect 9500 5076 9508 5084
rect 9612 5076 9620 5084
rect 9708 5076 9716 5084
rect 9884 5076 9892 5084
rect 10028 5076 10036 5084
rect 524 5056 532 5064
rect 3452 5056 3460 5064
rect 8972 5056 8980 5064
rect 236 5036 244 5044
rect 684 5036 692 5044
rect 1132 5036 1140 5044
rect 1820 5036 1828 5044
rect 2284 5036 2292 5044
rect 2316 5036 2324 5044
rect 3468 5036 3476 5044
rect 3854 5036 3862 5044
rect 4092 5036 4100 5044
rect 4556 5036 4564 5044
rect 4828 5036 4836 5044
rect 5436 5036 5444 5044
rect 5724 5036 5732 5044
rect 6108 5036 6116 5044
rect 6396 5036 6404 5044
rect 6860 5036 6868 5044
rect 7068 5036 7076 5044
rect 7292 5036 7300 5044
rect 7740 5036 7748 5044
rect 8124 5036 8132 5044
rect 8348 5036 8356 5044
rect 8396 5036 8404 5044
rect 8588 5036 8596 5044
rect 9196 5036 9204 5044
rect 9244 5036 9252 5044
rect 9900 5036 9908 5044
rect 12 4976 20 4984
rect 252 4976 260 4984
rect 972 4976 980 4984
rect 1340 4976 1348 4984
rect 1836 4976 1844 4984
rect 2044 4976 2052 4984
rect 2940 4976 2948 4984
rect 3164 4976 3172 4984
rect 3420 4976 3428 4984
rect 3644 4976 3652 4984
rect 3932 4976 3940 4984
rect 4364 4976 4372 4984
rect 4748 4976 4756 4984
rect 4764 4976 4772 4984
rect 4988 4976 4996 4984
rect 5836 4976 5844 4984
rect 6540 4976 6548 4984
rect 7132 4976 7140 4984
rect 7358 4976 7366 4984
rect 7612 4976 7620 4984
rect 8460 4976 8468 4984
rect 8476 4976 8484 4984
rect 10172 4976 10180 4984
rect 204 4936 212 4944
rect 668 4936 676 4944
rect 908 4936 916 4944
rect 1116 4936 1124 4944
rect 1228 4936 1236 4944
rect 1564 4936 1572 4944
rect 1676 4936 1684 4944
rect 1900 4936 1908 4944
rect 3644 4956 3652 4964
rect 8076 4956 8084 4964
rect 2476 4936 2484 4944
rect 2588 4936 2596 4944
rect 2796 4936 2804 4944
rect 3036 4936 3044 4944
rect 3260 4936 3268 4944
rect 3500 4936 3508 4944
rect 3836 4936 3844 4944
rect 4076 4936 4084 4944
rect 4172 4936 4180 4944
rect 4492 4936 4500 4944
rect 4604 4936 4612 4944
rect 4940 4936 4948 4944
rect 5180 4936 5188 4944
rect 5452 4936 5460 4944
rect 5596 4936 5604 4944
rect 5692 4936 5700 4944
rect 5916 4936 5924 4944
rect 6140 4936 6148 4944
rect 6348 4936 6356 4944
rect 6684 4936 6692 4944
rect 6796 4936 6804 4944
rect 7004 4936 7012 4944
rect 7228 4936 7236 4944
rect 7436 4936 7444 4944
rect 7772 4936 7780 4944
rect 7884 4936 7892 4944
rect 8204 4936 8212 4944
rect 8316 4936 8324 4944
rect 8668 4936 8676 4944
rect 8764 4936 8772 4944
rect 8972 4936 8980 4944
rect 9164 4936 9172 4944
rect 9196 4936 9204 4944
rect 9404 4936 9412 4944
rect 9580 4936 9588 4944
rect 9612 4936 9620 4944
rect 9820 4936 9828 4944
rect 2764 4916 2772 4924
rect 6972 4916 6980 4924
rect 7868 4916 7876 4924
rect 252 4896 260 4904
rect 508 4896 516 4904
rect 940 4896 948 4904
rect 1116 4896 1124 4904
rect 1196 4896 1204 4904
rect 1564 4896 1572 4904
rect 1660 4896 1668 4904
rect 1900 4896 1908 4904
rect 2316 4896 2324 4904
rect 2508 4896 2516 4904
rect 2524 4896 2532 4904
rect 2796 4896 2804 4904
rect 3020 4896 3028 4904
rect 3260 4896 3268 4904
rect 3484 4896 3492 4904
rect 3868 4896 3876 4904
rect 4076 4896 4084 4904
rect 4156 4896 4164 4904
rect 4524 4896 4532 4904
rect 4604 4896 4612 4904
rect 4956 4896 4964 4904
rect 5180 4896 5188 4904
rect 5628 4896 5636 4904
rect 5692 4896 5700 4904
rect 5900 4896 5908 4904
rect 6348 4896 6356 4904
rect 6700 4896 6708 4904
rect 6780 4896 6788 4904
rect 6988 4896 6996 4904
rect 7164 4896 7172 4904
rect 7436 4896 7444 4904
rect 7772 4896 7780 4904
rect 8220 4896 8228 4904
rect 8300 4896 8308 4904
rect 8668 4896 8676 4904
rect 8748 4896 8756 4904
rect 9180 4896 9188 4904
rect 9388 4896 9396 4904
rect 9612 4896 9620 4904
rect 10028 4896 10036 4904
rect 6332 4876 6340 4884
rect 6508 4876 6516 4884
rect 7580 4876 7588 4884
rect 1404 4856 1412 4864
rect 4348 4856 4356 4864
rect 2108 4836 2116 4844
rect 5258 4836 5266 4844
rect 7372 4836 7380 4844
rect 8028 4836 8036 4844
rect 9340 4836 9348 4844
rect 3228 4776 3236 4784
rect 4140 4776 4148 4784
rect 5916 4776 5924 4784
rect 6140 4776 6148 4784
rect 8316 4776 8324 4784
rect 2014 4736 2022 4744
rect 7836 4736 7844 4744
rect 76 4716 84 4724
rect 444 4716 452 4724
rect 524 4716 532 4724
rect 684 4716 692 4724
rect 908 4716 916 4724
rect 1148 4716 1156 4724
rect 1212 4716 1220 4724
rect 1372 4716 1380 4724
rect 1564 4716 1572 4724
rect 1788 4716 1796 4724
rect 1884 4716 1892 4724
rect 2044 4716 2052 4724
rect 2476 4716 2484 4724
rect 2700 4716 2708 4724
rect 2780 4716 2788 4724
rect 2796 4716 2804 4724
rect 3196 4716 3204 4724
rect 3404 4716 3412 4724
rect 3596 4716 3604 4724
rect 3820 4716 3828 4724
rect 4060 4716 4068 4724
rect 4284 4716 4292 4724
rect 4492 4716 4500 4724
rect 4572 4716 4580 4724
rect 4940 4716 4948 4724
rect 5164 4716 5172 4724
rect 5260 4716 5268 4724
rect 5484 4716 5492 4724
rect 5708 4716 5716 4724
rect 5932 4716 5940 4724
rect 5946 4716 5954 4724
rect 6300 4716 6308 4724
rect 6492 4716 6500 4724
rect 6588 4716 6596 4724
rect 6940 4716 6948 4724
rect 6972 4716 6980 4724
rect 7260 4716 7268 4724
rect 7596 4716 7604 4724
rect 7676 4716 7684 4724
rect 8044 4716 8052 4724
rect 8252 4716 8260 4724
rect 8492 4716 8500 4724
rect 8572 4716 8580 4724
rect 8780 4716 8788 4724
rect 9148 4716 9156 4724
rect 9228 4716 9236 4724
rect 9580 4716 9588 4724
rect 9692 4716 9700 4724
rect 10092 4716 10100 4724
rect 92 4676 100 4684
rect 444 4676 452 4684
rect 668 4676 676 4684
rect 700 4676 708 4684
rect 908 4676 916 4684
rect 1132 4676 1140 4684
rect 1340 4676 1348 4684
rect 1548 4676 1556 4684
rect 1788 4676 1796 4684
rect 1900 4676 1908 4684
rect 2092 4676 2100 4684
rect 2460 4676 2468 4684
rect 2700 4676 2708 4684
rect 2716 4676 2724 4684
rect 2812 4676 2820 4684
rect 3148 4676 3156 4684
rect 3580 4676 3588 4684
rect 3804 4676 3812 4684
rect 4268 4676 4276 4684
rect 4300 4676 4308 4684
rect 4476 4676 4484 4684
rect 4588 4676 4596 4684
rect 4924 4676 4932 4684
rect 4956 4676 4964 4684
rect 5180 4676 5188 4684
rect 5276 4676 5284 4684
rect 5500 4676 5508 4684
rect 5724 4676 5732 4684
rect 5948 4676 5956 4684
rect 6124 4676 6132 4684
rect 6284 4676 6292 4684
rect 6300 4676 6308 4684
rect 6508 4676 6516 4684
rect 6604 4676 6612 4684
rect 6972 4676 6980 4684
rect 7036 4676 7044 4684
rect 7260 4676 7268 4684
rect 7580 4676 7588 4684
rect 7692 4676 7700 4684
rect 8252 4676 8260 4684
rect 8476 4676 8484 4684
rect 8588 4676 8596 4684
rect 8796 4676 8804 4684
rect 9132 4676 9140 4684
rect 9212 4676 9220 4684
rect 9388 4676 9396 4684
rect 9580 4676 9588 4684
rect 9692 4676 9700 4684
rect 9916 4676 9924 4684
rect 1596 4656 1604 4664
rect 2956 4656 2964 4664
rect 236 4636 244 4644
rect 284 4636 292 4644
rect 924 4636 932 4644
rect 1420 4636 1428 4644
rect 2252 4636 2260 4644
rect 2268 4636 2276 4644
rect 2524 4636 2532 4644
rect 2956 4636 2964 4644
rect 3676 4636 3684 4644
rect 3884 4636 3892 4644
rect 4716 4636 4724 4644
rect 4732 4636 4740 4644
rect 5468 4636 5476 4644
rect 5644 4636 5652 4644
rect 6748 4636 6756 4644
rect 6796 4636 6804 4644
rect 7164 4636 7172 4644
rect 7390 4636 7398 4644
rect 7452 4636 7460 4644
rect 7836 4636 7844 4644
rect 8284 4636 8292 4644
rect 8716 4636 8724 4644
rect 8924 4636 8932 4644
rect 8940 4636 8948 4644
rect 9388 4636 9396 4644
rect 10252 4636 10260 4644
rect 12 4576 20 4584
rect 684 4576 692 4584
rect 1372 4576 1380 4584
rect 1404 4576 1412 4584
rect 1836 4576 1844 4584
rect 2092 4576 2100 4584
rect 2108 4576 2116 4584
rect 2300 4576 2308 4584
rect 3196 4576 3204 4584
rect 3468 4576 3476 4584
rect 3916 4576 3924 4584
rect 4140 4576 4148 4584
rect 4300 4576 4308 4584
rect 4572 4576 4580 4584
rect 5180 4576 5188 4584
rect 5242 4576 5250 4584
rect 5692 4576 5700 4584
rect 6316 4576 6324 4584
rect 6972 4576 6980 4584
rect 7004 4576 7012 4584
rect 8284 4576 8292 4584
rect 8732 4576 8740 4584
rect 10028 4576 10036 4584
rect 524 4556 532 4564
rect 2572 4556 2580 4564
rect 2940 4556 2948 4564
rect 8316 4556 8324 4564
rect 8716 4556 8724 4564
rect 9580 4556 9588 4564
rect 204 4536 212 4544
rect 316 4536 324 4544
rect 556 4536 564 4544
rect 908 4536 916 4544
rect 988 4536 996 4544
rect 1132 4536 1140 4544
rect 1244 4536 1252 4544
rect 1596 4536 1604 4544
rect 1708 4536 1716 4544
rect 1932 4536 1940 4544
rect 2268 4536 2276 4544
rect 2492 4536 2500 4544
rect 2716 4536 2724 4544
rect 2812 4536 2820 4544
rect 3148 4536 3156 4544
rect 3388 4536 3396 4544
rect 3612 4536 3620 4544
rect 3836 4536 3844 4544
rect 4076 4536 4084 4544
rect 4268 4536 4276 4544
rect 4508 4536 4516 4544
rect 4732 4536 4740 4544
rect 4828 4536 4836 4544
rect 5356 4536 5364 4544
rect 5596 4536 5604 4544
rect 5836 4536 5844 4544
rect 5948 4536 5956 4544
rect 6156 4536 6164 4544
rect 6476 4536 6484 4544
rect 6604 4536 6612 4544
rect 6828 4536 6836 4544
rect 7164 4536 7172 4544
rect 7212 4536 7220 4544
rect 7276 4536 7284 4544
rect 7452 4536 7460 4544
rect 7708 4536 7716 4544
rect 7900 4536 7908 4544
rect 8124 4536 8132 4544
rect 8444 4536 8452 4544
rect 8572 4536 8580 4544
rect 8892 4536 8900 4544
rect 8908 4536 8916 4544
rect 9116 4536 9124 4544
rect 9228 4536 9236 4544
rect 9404 4536 9412 4544
rect 9548 4536 9556 4544
rect 9788 4536 9796 4544
rect 9852 4536 9860 4544
rect 10204 4536 10212 4544
rect 1180 4516 1188 4524
rect 3676 4516 3684 4524
rect 6332 4516 6340 4524
rect 7436 4516 7444 4524
rect 252 4496 260 4504
rect 316 4496 324 4504
rect 476 4496 484 4504
rect 1244 4496 1252 4504
rect 1596 4496 1604 4504
rect 1692 4496 1700 4504
rect 1900 4496 1908 4504
rect 2284 4496 2292 4504
rect 2524 4496 2532 4504
rect 2764 4496 2772 4504
rect 2796 4496 2804 4504
rect 3164 4496 3172 4504
rect 3388 4496 3396 4504
rect 3852 4496 3860 4504
rect 4060 4496 4068 4504
rect 4268 4496 4276 4504
rect 4524 4496 4532 4504
rect 4716 4496 4724 4504
rect 4748 4496 4756 4504
rect 5036 4496 5044 4504
rect 5372 4496 5380 4504
rect 5612 4496 5620 4504
rect 5836 4496 5844 4504
rect 5916 4496 5924 4504
rect 6140 4496 6148 4504
rect 6492 4496 6500 4504
rect 6588 4496 6596 4504
rect 6828 4496 6836 4504
rect 7164 4496 7172 4504
rect 7260 4496 7268 4504
rect 7468 4496 7476 4504
rect 7900 4496 7908 4504
rect 8476 4496 8484 4504
rect 8556 4496 8564 4504
rect 8908 4496 8916 4504
rect 9132 4496 9140 4504
rect 9212 4496 9220 4504
rect 9548 4496 9556 4504
rect 9788 4496 9796 4504
rect 9852 4496 9860 4504
rect 9884 4496 9892 4504
rect 10252 4496 10260 4504
rect 748 4456 756 4464
rect 3004 4456 3012 4464
rect 6140 4456 6148 4464
rect 1452 4436 1460 4444
rect 3660 4436 3668 4444
rect 5452 4436 5460 4444
rect 6748 4436 6756 4444
rect 7836 4436 7844 4444
rect 9356 4436 9364 4444
rect 10076 4436 10084 4444
rect 684 4376 692 4384
rect 1164 4376 1172 4384
rect 1644 4376 1652 4384
rect 3180 4376 3188 4384
rect 8812 4376 8820 4384
rect 8620 4336 8628 4344
rect 220 4316 228 4324
rect 492 4316 500 4324
rect 554 4316 562 4324
rect 908 4316 916 4324
rect 1004 4316 1012 4324
rect 1356 4316 1364 4324
rect 1436 4316 1444 4324
rect 1804 4316 1812 4324
rect 2044 4316 2052 4324
rect 2252 4316 2260 4324
rect 2332 4316 2340 4324
rect 2700 4316 2708 4324
rect 2796 4316 2804 4324
rect 3164 4316 3172 4324
rect 3372 4316 3380 4324
rect 3612 4316 3620 4324
rect 3804 4316 3812 4324
rect 4012 4316 4020 4324
rect 4236 4316 4244 4324
rect 4316 4316 4324 4324
rect 4524 4316 4532 4324
rect 4924 4316 4932 4324
rect 5084 4316 5092 4324
rect 5308 4316 5316 4324
rect 5388 4316 5396 4324
rect 5596 4316 5604 4324
rect 5932 4316 5940 4324
rect 6156 4316 6164 4324
rect 6380 4316 6388 4324
rect 6620 4316 6628 4324
rect 6828 4316 6836 4324
rect 7036 4316 7044 4324
rect 7260 4316 7268 4324
rect 7468 4316 7476 4324
rect 7548 4316 7556 4324
rect 7916 4316 7924 4324
rect 8108 4316 8116 4324
rect 8188 4316 8196 4324
rect 8412 4316 8420 4324
rect 8620 4316 8628 4324
rect 8828 4316 8836 4324
rect 9180 4316 9188 4324
rect 9420 4316 9428 4324
rect 9612 4316 9620 4324
rect 9852 4316 9860 4324
rect 9900 4316 9908 4324
rect 2556 4296 2564 4304
rect 7324 4296 7332 4304
rect 204 4276 212 4284
rect 460 4276 468 4284
rect 556 4276 564 4284
rect 908 4276 916 4284
rect 1004 4276 1012 4284
rect 1452 4276 1460 4284
rect 1788 4276 1796 4284
rect 1804 4276 1812 4284
rect 2012 4276 2020 4284
rect 2252 4276 2260 4284
rect 2348 4276 2356 4284
rect 2476 4276 2484 4284
rect 2700 4276 2708 4284
rect 2716 4276 2724 4284
rect 3148 4276 3156 4284
rect 3580 4276 3588 4284
rect 3788 4276 3796 4284
rect 3996 4276 4004 4284
rect 4060 4276 4068 4284
rect 4220 4276 4228 4284
rect 4316 4276 4324 4284
rect 4540 4276 4548 4284
rect 4860 4276 4868 4284
rect 5068 4276 5076 4284
rect 5276 4276 5284 4284
rect 5388 4276 5396 4284
rect 5756 4276 5764 4284
rect 5916 4276 5924 4284
rect 6156 4276 6164 4284
rect 6380 4276 6388 4284
rect 6604 4276 6612 4284
rect 6812 4276 6820 4284
rect 7052 4276 7060 4284
rect 7244 4276 7252 4284
rect 7468 4276 7476 4284
rect 7564 4276 7572 4284
rect 7692 4276 7700 4284
rect 7884 4276 7892 4284
rect 8092 4276 8100 4284
rect 8220 4276 8228 4284
rect 8428 4276 8436 4284
rect 8636 4276 8644 4284
rect 8844 4276 8852 4284
rect 9164 4276 9172 4284
rect 9372 4276 9380 4284
rect 9420 4276 9428 4284
rect 9612 4276 9620 4284
rect 9836 4276 9844 4284
rect 9932 4276 9940 4284
rect 3004 4256 3012 4264
rect 4684 4256 4692 4264
rect 6188 4256 6196 4264
rect 12 4236 20 4244
rect 236 4236 244 4244
rect 764 4236 772 4244
rect 1196 4236 1204 4244
rect 1580 4236 1588 4244
rect 2076 4236 2084 4244
rect 2956 4236 2964 4244
rect 3420 4236 3428 4244
rect 3660 4236 3668 4244
rect 3868 4236 3876 4244
rect 4092 4236 4100 4244
rect 4476 4236 4484 4244
rect 4668 4236 4676 4244
rect 4924 4236 4932 4244
rect 5162 4236 5170 4244
rect 5756 4236 5764 4244
rect 6012 4236 6020 4244
rect 6460 4236 6468 4244
rect 6668 4236 6676 4244
rect 6892 4236 6900 4244
rect 7116 4236 7124 4244
rect 7740 4236 7748 4244
rect 7964 4236 7972 4244
rect 8332 4236 8340 4244
rect 8988 4236 8996 4244
rect 9036 4236 9044 4244
rect 9260 4236 9268 4244
rect 9692 4236 9700 4244
rect 10060 4236 10068 4244
rect 76 4176 84 4184
rect 460 4176 468 4184
rect 668 4176 676 4184
rect 924 4176 932 4184
rect 1612 4176 1620 4184
rect 2092 4176 2100 4184
rect 2332 4176 2340 4184
rect 2492 4176 2500 4184
rect 2716 4176 2724 4184
rect 2956 4176 2964 4184
rect 3228 4176 3236 4184
rect 3420 4176 3428 4184
rect 3644 4176 3652 4184
rect 4316 4176 4324 4184
rect 5212 4176 5220 4184
rect 5932 4176 5940 4184
rect 6348 4176 6356 4184
rect 6780 4176 6788 4184
rect 7196 4176 7204 4184
rect 7708 4176 7716 4184
rect 8108 4176 8116 4184
rect 8524 4176 8532 4184
rect 8812 4176 8820 4184
rect 9212 4176 9220 4184
rect 9628 4176 9636 4184
rect 9884 4176 9892 4184
rect 10268 4176 10276 4184
rect 940 4156 948 4164
rect 1836 4156 1844 4164
rect 4764 4156 4772 4164
rect 5260 4156 5268 4164
rect 8316 4156 8324 4164
rect 204 4136 212 4144
rect 316 4136 324 4144
rect 540 4136 548 4144
rect 764 4136 772 4144
rect 1116 4136 1124 4144
rect 1228 4136 1236 4144
rect 1388 4136 1396 4144
rect 1596 4136 1604 4144
rect 1804 4136 1812 4144
rect 2012 4136 2020 4144
rect 2460 4136 2468 4144
rect 2700 4136 2708 4144
rect 2924 4136 2932 4144
rect 3132 4136 3140 4144
rect 3404 4136 3412 4144
rect 3612 4136 3620 4144
rect 3820 4136 3828 4144
rect 4124 4136 4132 4144
rect 4172 4136 4180 4144
rect 4364 4136 4372 4144
rect 4540 4136 4548 4144
rect 4748 4136 4756 4144
rect 4956 4136 4964 4144
rect 5068 4136 5076 4144
rect 5388 4136 5396 4144
rect 5628 4136 5636 4144
rect 5740 4136 5748 4144
rect 5980 4136 5988 4144
rect 6204 4136 6212 4144
rect 6428 4136 6436 4144
rect 6860 4136 6868 4144
rect 7068 4136 7076 4144
rect 7388 4136 7396 4144
rect 7484 4136 7492 4144
rect 7836 4136 7844 4144
rect 7948 4136 7956 4144
rect 8124 4136 8132 4144
rect 8284 4136 8292 4144
rect 8492 4136 8500 4144
rect 8732 4136 8740 4144
rect 8956 4136 8964 4144
rect 9068 4136 9076 4144
rect 9276 4136 9284 4144
rect 9500 4136 9508 4144
rect 9692 4136 9700 4144
rect 9916 4136 9924 4144
rect 1820 4116 1828 4124
rect 3660 4116 3668 4124
rect 3852 4116 3860 4124
rect 7676 4116 7684 4124
rect 8348 4116 8356 4124
rect 9468 4116 9476 4124
rect 236 4096 244 4104
rect 316 4096 324 4104
rect 524 4096 532 4104
rect 764 4096 772 4104
rect 1116 4096 1124 4104
rect 1212 4096 1220 4104
rect 1420 4096 1428 4104
rect 1580 4096 1588 4104
rect 2076 4096 2084 4104
rect 2236 4096 2244 4104
rect 2476 4096 2484 4104
rect 2700 4096 2708 4104
rect 2956 4096 2964 4104
rect 3150 4096 3158 4104
rect 3388 4096 3396 4104
rect 3612 4096 3620 4104
rect 3836 4096 3844 4104
rect 4060 4096 4068 4104
rect 4140 4096 4148 4104
rect 4524 4096 4532 4104
rect 4732 4096 4740 4104
rect 4972 4096 4980 4104
rect 5052 4096 5060 4104
rect 5420 4096 5428 4104
rect 5660 4096 5668 4104
rect 5740 4096 5748 4104
rect 5964 4096 5972 4104
rect 6188 4096 6196 4104
rect 6412 4096 6420 4104
rect 6636 4096 6644 4104
rect 6844 4096 6852 4104
rect 7404 4096 7412 4104
rect 7484 4096 7492 4104
rect 7836 4096 7844 4104
rect 7932 4096 7940 4104
rect 8494 4096 8502 4104
rect 8732 4096 8740 4104
rect 8956 4096 8964 4104
rect 9036 4096 9044 4104
rect 9276 4096 9284 4104
rect 9484 4096 9492 4104
rect 9708 4096 9716 4104
rect 9916 4096 9924 4104
rect 4588 4056 4596 4064
rect 6188 4056 6196 4064
rect 5484 4036 5492 4044
rect 7260 4036 7268 4044
rect 76 3976 84 3984
rect 524 3976 532 3984
rect 3452 3976 3460 3984
rect 4076 3976 4084 3984
rect 6588 3976 6596 3984
rect 6972 3976 6980 3984
rect 6988 3976 6996 3984
rect 9580 3976 9588 3984
rect 5724 3936 5732 3944
rect 236 3916 244 3924
rect 428 3916 436 3924
rect 668 3916 676 3924
rect 908 3916 916 3924
rect 1100 3916 1108 3924
rect 1196 3916 1204 3924
rect 1420 3916 1428 3924
rect 1772 3916 1780 3924
rect 1868 3916 1876 3924
rect 2236 3916 2244 3924
rect 2476 3916 2484 3924
rect 2732 3916 2740 3924
rect 2924 3916 2932 3924
rect 3196 3916 3204 3924
rect 3372 3916 3380 3924
rect 3852 3916 3860 3924
rect 3932 3916 3940 3924
rect 4332 3916 4340 3924
rect 4380 3916 4388 3924
rect 4604 3916 4612 3924
rect 4844 3916 4852 3924
rect 5068 3916 5076 3924
rect 5260 3916 5268 3924
rect 5500 3916 5508 3924
rect 5868 3916 5876 3924
rect 6092 3916 6100 3924
rect 6172 3916 6180 3924
rect 6396 3916 6404 3924
rect 6748 3916 6756 3924
rect 6828 3916 6836 3924
rect 7180 3916 7188 3924
rect 7388 3916 7396 3924
rect 7468 3916 7476 3924
rect 7676 3916 7684 3924
rect 7900 3916 7908 3924
rect 8092 3916 8100 3924
rect 8476 3916 8484 3924
rect 8540 3916 8548 3924
rect 8892 3916 8900 3924
rect 9132 3916 9140 3924
rect 9212 3916 9220 3924
rect 9436 3916 9444 3924
rect 9660 3916 9668 3924
rect 9852 3916 9860 3924
rect 10076 3916 10084 3924
rect 1612 3896 1620 3904
rect 3612 3896 3620 3904
rect 204 3876 212 3884
rect 652 3876 660 3884
rect 1116 3876 1124 3884
rect 1212 3876 1220 3884
rect 1772 3876 1780 3884
rect 1884 3876 1892 3884
rect 2460 3876 2468 3884
rect 2668 3876 2676 3884
rect 2908 3876 2916 3884
rect 2956 3876 2964 3884
rect 3132 3876 3140 3884
rect 3372 3876 3380 3884
rect 3596 3876 3604 3884
rect 3820 3876 3828 3884
rect 3948 3876 3956 3884
rect 4284 3876 4292 3884
rect 4396 3876 4404 3884
rect 4620 3876 4628 3884
rect 4844 3876 4852 3884
rect 5068 3876 5076 3884
rect 5292 3876 5300 3884
rect 5484 3876 5492 3884
rect 5516 3876 5524 3884
rect 5868 3876 5876 3884
rect 6060 3876 6068 3884
rect 6188 3876 6196 3884
rect 6412 3876 6420 3884
rect 6732 3876 6740 3884
rect 6828 3876 6836 3884
rect 7164 3876 7172 3884
rect 7372 3876 7380 3884
rect 7468 3876 7476 3884
rect 7484 3876 7492 3884
rect 7612 3876 7620 3884
rect 7692 3876 7700 3884
rect 7916 3876 7924 3884
rect 8124 3876 8132 3884
rect 8444 3876 8452 3884
rect 8476 3876 8484 3884
rect 9100 3876 9108 3884
rect 9212 3876 9220 3884
rect 9452 3876 9460 3884
rect 9660 3876 9668 3884
rect 9884 3876 9892 3884
rect 10092 3876 10100 3884
rect 2716 3856 2724 3864
rect 5708 3856 5716 3864
rect 7244 3856 7252 3864
rect 8044 3856 8052 3864
rect 284 3836 292 3844
rect 732 3836 740 3844
rect 1628 3836 1636 3844
rect 2014 3836 2022 3844
rect 2092 3836 2100 3844
rect 2524 3836 2532 3844
rect 3228 3836 3236 3844
rect 3644 3836 3652 3844
rect 4156 3836 4164 3844
rect 4540 3836 4548 3844
rect 4764 3836 4772 3844
rect 4988 3836 4996 3844
rect 5260 3836 5268 3844
rect 5948 3836 5956 3844
rect 6588 3836 6596 3844
rect 7836 3836 7844 3844
rect 8300 3836 8308 3844
rect 8316 3836 8324 3844
rect 8700 3836 8708 3844
rect 8732 3836 8740 3844
rect 8972 3836 8980 3844
rect 9356 3836 9364 3844
rect 9820 3836 9828 3844
rect 10012 3836 10020 3844
rect 10236 3836 10244 3844
rect 12 3776 20 3784
rect 252 3776 260 3784
rect 700 3776 708 3784
rect 924 3776 932 3784
rect 1148 3776 1156 3784
rect 2044 3776 2052 3784
rect 2748 3776 2756 3784
rect 3260 3776 3268 3784
rect 3420 3776 3428 3784
rect 3854 3776 3862 3784
rect 4140 3776 4148 3784
rect 4364 3776 4372 3784
rect 4556 3776 4564 3784
rect 4796 3776 4804 3784
rect 5276 3776 5284 3784
rect 6828 3776 6836 3784
rect 7004 3776 7012 3784
rect 7212 3776 7220 3784
rect 7676 3776 7684 3784
rect 7916 3776 7924 3784
rect 8364 3776 8372 3784
rect 8764 3776 8772 3784
rect 8988 3776 8996 3784
rect 9852 3776 9860 3784
rect 10076 3776 10084 3784
rect 10092 3776 10100 3784
rect 1674 3756 1682 3764
rect 1836 3756 1844 3764
rect 2268 3756 2276 3764
rect 2972 3756 2980 3764
rect 7692 3756 7700 3764
rect 9452 3756 9460 3764
rect 204 3736 212 3744
rect 444 3736 452 3744
rect 460 3736 468 3744
rect 668 3736 676 3744
rect 940 3736 948 3744
rect 1132 3736 1140 3744
rect 1340 3736 1348 3744
rect 1628 3736 1636 3744
rect 1804 3736 1812 3744
rect 2012 3736 2020 3744
rect 2252 3736 2260 3744
rect 2476 3736 2484 3744
rect 2588 3736 2596 3744
rect 2940 3736 2948 3744
rect 3164 3736 3172 3744
rect 3404 3736 3412 3744
rect 3628 3736 3636 3744
rect 3708 3736 3716 3744
rect 4044 3736 4052 3744
rect 4284 3736 4292 3744
rect 4492 3736 4500 3744
rect 4732 3736 4740 3744
rect 4956 3736 4964 3744
rect 5196 3736 5204 3744
rect 5420 3736 5428 3744
rect 5532 3736 5540 3744
rect 5756 3736 5764 3744
rect 5964 3736 5972 3744
rect 6188 3736 6196 3744
rect 6636 3736 6644 3744
rect 6972 3736 6980 3744
rect 7180 3736 7188 3744
rect 7388 3736 7396 3744
rect 7468 3736 7476 3744
rect 7852 3736 7860 3744
rect 8108 3736 8116 3744
rect 8172 3736 8180 3744
rect 8396 3736 8404 3744
rect 8604 3736 8612 3744
rect 8844 3736 8852 3744
rect 9164 3736 9172 3744
rect 9276 3736 9284 3744
rect 9500 3736 9508 3744
rect 9692 3736 9700 3744
rect 9916 3736 9924 3744
rect 10236 3736 10244 3744
rect 6588 3716 6596 3724
rect 9020 3716 9028 3724
rect 236 3696 244 3704
rect 460 3696 468 3704
rect 700 3696 708 3704
rect 908 3696 916 3704
rect 1116 3696 1124 3704
rect 1580 3696 1588 3704
rect 1852 3696 1860 3704
rect 2028 3696 2036 3704
rect 2252 3696 2260 3704
rect 2540 3696 2548 3704
rect 2588 3696 2596 3704
rect 2780 3696 2788 3704
rect 2940 3696 2948 3704
rect 3228 3696 3236 3704
rect 3404 3696 3412 3704
rect 3692 3696 3700 3704
rect 3724 3696 3732 3704
rect 4060 3696 4068 3704
rect 4300 3696 4308 3704
rect 4508 3696 4516 3704
rect 4748 3696 4756 3704
rect 4988 3696 4996 3704
rect 5196 3696 5204 3704
rect 5420 3696 5428 3704
rect 5532 3696 5540 3704
rect 5740 3696 5748 3704
rect 6172 3696 6180 3704
rect 6396 3696 6404 3704
rect 6604 3696 6612 3704
rect 6972 3696 6980 3704
rect 7196 3696 7204 3704
rect 7404 3696 7412 3704
rect 7500 3696 7508 3704
rect 7884 3696 7892 3704
rect 8140 3696 8148 3704
rect 8172 3696 8180 3704
rect 8380 3696 8388 3704
rect 3180 3676 3188 3684
rect 3916 3676 3924 3684
rect 6172 3676 6180 3684
rect 8828 3696 8836 3704
rect 9180 3696 9188 3704
rect 9260 3696 9268 3704
rect 9468 3696 9476 3704
rect 9852 3696 9860 3704
rect 10268 3696 10276 3704
rect 5756 3656 5764 3664
rect 5004 3636 5012 3644
rect 6764 3636 6772 3644
rect 60 3576 68 3584
rect 2556 3576 2564 3584
rect 3020 3576 3028 3584
rect 4988 3576 4996 3584
rect 8348 3576 8356 3584
rect 6940 3556 6948 3564
rect 4924 3536 4932 3544
rect 220 3516 228 3524
rect 444 3516 452 3524
rect 668 3516 676 3524
rect 892 3516 900 3524
rect 1196 3516 1204 3524
rect 1342 3516 1350 3524
rect 1452 3516 1460 3524
rect 2028 3516 2036 3524
rect 2268 3516 2276 3524
rect 2476 3516 2484 3524
rect 2700 3516 2708 3524
rect 2956 3516 2964 3524
rect 3180 3516 3188 3524
rect 3372 3516 3380 3524
rect 3596 3516 3604 3524
rect 3836 3516 3844 3524
rect 4028 3516 4036 3524
rect 4108 3516 4116 3524
rect 4476 3516 4484 3524
rect 4508 3516 4516 3524
rect 4780 3516 4788 3524
rect 5148 3516 5156 3524
rect 5372 3516 5380 3524
rect 5388 3516 5396 3524
rect 5804 3516 5812 3524
rect 5900 3516 5908 3524
rect 6124 3516 6132 3524
rect 6332 3516 6340 3524
rect 6572 3516 6580 3524
rect 6780 3516 6788 3524
rect 7164 3516 7172 3524
rect 7228 3516 7236 3524
rect 7580 3516 7588 3524
rect 7676 3516 7684 3524
rect 7900 3516 7908 3524
rect 8124 3516 8132 3524
rect 8492 3516 8500 3524
rect 8572 3516 8580 3524
rect 8780 3516 8788 3524
rect 9020 3516 9028 3524
rect 9228 3516 9236 3524
rect 9452 3516 9460 3524
rect 9676 3516 9684 3524
rect 9900 3516 9908 3524
rect 10108 3516 10116 3524
rect 1132 3496 1140 3504
rect 1660 3496 1668 3504
rect 204 3476 212 3484
rect 236 3476 244 3484
rect 444 3476 452 3484
rect 956 3476 964 3484
rect 1116 3476 1124 3484
rect 1340 3476 1348 3484
rect 1436 3476 1444 3484
rect 1804 3476 1812 3484
rect 6540 3496 6548 3504
rect 2012 3476 2020 3484
rect 2252 3476 2260 3484
rect 2268 3476 2276 3484
rect 2444 3476 2452 3484
rect 2700 3476 2708 3484
rect 2716 3476 2724 3484
rect 2924 3476 2932 3484
rect 3148 3476 3156 3484
rect 3372 3476 3380 3484
rect 3580 3476 3588 3484
rect 3804 3476 3812 3484
rect 3836 3476 3844 3484
rect 4012 3476 4020 3484
rect 4124 3476 4132 3484
rect 4476 3476 4484 3484
rect 4572 3476 4580 3484
rect 4796 3476 4804 3484
rect 5148 3476 5156 3484
rect 5340 3476 5348 3484
rect 5468 3476 5476 3484
rect 5804 3476 5812 3484
rect 5916 3476 5924 3484
rect 6140 3476 6148 3484
rect 6572 3476 6580 3484
rect 7132 3476 7140 3484
rect 7244 3476 7252 3484
rect 7564 3476 7572 3484
rect 7692 3476 7700 3484
rect 7916 3476 7924 3484
rect 8108 3476 8116 3484
rect 8124 3476 8132 3484
rect 8476 3476 8484 3484
rect 8572 3476 8580 3484
rect 8812 3476 8820 3484
rect 9020 3476 9028 3484
rect 9244 3476 9252 3484
rect 9468 3476 9476 3484
rect 9692 3476 9700 3484
rect 9900 3476 9908 3484
rect 10124 3476 10132 3484
rect 10252 3476 10260 3484
rect 1644 3456 1652 3464
rect 3612 3456 3620 3464
rect 524 3436 532 3444
rect 972 3436 980 3444
rect 2044 3436 2052 3444
rect 3228 3436 3236 3444
rect 3450 3436 3458 3444
rect 4252 3436 4260 3444
rect 4316 3436 4324 3444
rect 4716 3436 4724 3444
rect 5212 3436 5220 3444
rect 5612 3436 5620 3444
rect 5660 3436 5668 3444
rect 6060 3436 6068 3444
rect 6924 3436 6932 3444
rect 7388 3436 7396 3444
rect 7436 3436 7444 3444
rect 7820 3436 7828 3444
rect 8268 3436 8276 3444
rect 8716 3436 8724 3444
rect 8988 3436 8996 3444
rect 9164 3436 9172 3444
rect 9388 3436 9396 3444
rect 9612 3436 9620 3444
rect 10044 3436 10052 3444
rect 60 3376 68 3384
rect 300 3376 308 3384
rect 540 3376 548 3384
rect 1180 3376 1188 3384
rect 1436 3376 1444 3384
rect 1836 3376 1844 3384
rect 2284 3376 2292 3384
rect 2572 3376 2580 3384
rect 2956 3376 2964 3384
rect 3644 3376 3652 3384
rect 4284 3376 4292 3384
rect 4332 3376 4340 3384
rect 5692 3376 5700 3384
rect 6108 3376 6116 3384
rect 6156 3376 6164 3384
rect 6332 3376 6340 3384
rect 6764 3376 6772 3384
rect 7068 3376 7076 3384
rect 7500 3376 7508 3384
rect 8124 3376 8132 3384
rect 8348 3376 8356 3384
rect 9036 3376 9044 3384
rect 9628 3376 9636 3384
rect 2556 3356 2564 3364
rect 2972 3356 2980 3364
rect 3196 3356 3204 3364
rect 204 3336 212 3344
rect 508 3336 516 3344
rect 668 3336 676 3344
rect 940 3336 948 3344
rect 1004 3336 1012 3344
rect 1244 3336 1252 3344
rect 1596 3336 1604 3344
rect 1708 3336 1716 3344
rect 1932 3336 1940 3344
rect 2124 3336 2132 3344
rect 2140 3336 2148 3344
rect 2380 3336 2388 3344
rect 2796 3336 2804 3344
rect 2812 3336 2820 3344
rect 3164 3336 3172 3344
rect 4748 3356 4756 3364
rect 9644 3356 9652 3364
rect 10060 3356 10068 3364
rect 3596 3336 3604 3344
rect 3836 3336 3844 3344
rect 4076 3336 4084 3344
rect 4156 3336 4164 3344
rect 4508 3336 4516 3344
rect 4732 3336 4740 3344
rect 4940 3336 4948 3344
rect 5180 3336 5188 3344
rect 5292 3336 5300 3344
rect 5516 3336 5524 3344
rect 5740 3336 5748 3344
rect 5964 3336 5972 3344
rect 6108 3336 6116 3344
rect 6140 3336 6148 3344
rect 6284 3336 6292 3344
rect 6524 3336 6532 3344
rect 6636 3336 6644 3344
rect 6844 3336 6852 3344
rect 7100 3336 7108 3344
rect 7324 3336 7332 3344
rect 7484 3336 7492 3344
rect 7708 3336 7716 3344
rect 7740 3336 7748 3344
rect 7964 3336 7972 3344
rect 8188 3336 8196 3344
rect 8428 3336 8436 3344
rect 8652 3336 8660 3344
rect 8860 3336 8868 3344
rect 9068 3336 9076 3344
rect 9244 3336 9252 3344
rect 9836 3336 9844 3344
rect 9916 3336 9924 3344
rect 220 3296 228 3304
rect 444 3296 452 3304
rect 908 3296 916 3304
rect 1004 3296 1012 3304
rect 1244 3296 1252 3304
rect 1436 3296 1444 3304
rect 1596 3296 1604 3304
rect 1692 3296 1700 3304
rect 1916 3296 1924 3304
rect 2124 3296 2132 3304
rect 2378 3296 2386 3304
rect 2732 3296 2740 3304
rect 2812 3296 2820 3304
rect 3228 3296 3236 3304
rect 3404 3296 3412 3304
rect 3612 3296 3620 3304
rect 4060 3296 4068 3304
rect 4092 3296 4100 3304
rect 4524 3296 4532 3304
rect 4716 3296 4724 3304
rect 5180 3296 5188 3304
rect 5212 3296 5220 3304
rect 5500 3296 5508 3304
rect 5724 3296 5732 3304
rect 5948 3296 5956 3304
rect 6300 3296 6308 3304
rect 6540 3296 6548 3304
rect 6620 3296 6628 3304
rect 6860 3296 6868 3304
rect 7068 3296 7076 3304
rect 7308 3296 7316 3304
rect 7644 3296 7652 3304
rect 7708 3296 7716 3304
rect 7948 3296 7956 3304
rect 8188 3296 8196 3304
rect 8428 3296 8436 3304
rect 7308 3276 7316 3284
rect 9052 3296 9060 3304
rect 9484 3296 9492 3304
rect 9836 3296 9844 3304
rect 9900 3296 9908 3304
rect 4572 3236 4580 3244
rect 5436 3236 5444 3244
rect 5884 3236 5892 3244
rect 7868 3236 7876 3244
rect 700 3176 708 3184
rect 3612 3176 3620 3184
rect 3836 3176 3844 3184
rect 8572 3176 8580 3184
rect 9836 3176 9844 3184
rect 2284 3156 2292 3164
rect 5130 3136 5138 3144
rect 5486 3136 5494 3144
rect 8988 3136 8996 3144
rect 284 3116 292 3124
rect 508 3116 516 3124
rect 876 3116 884 3124
rect 1084 3116 1092 3124
rect 1196 3116 1204 3124
rect 1372 3116 1380 3124
rect 1532 3116 1540 3124
rect 1612 3116 1620 3124
rect 1852 3116 1860 3124
rect 2076 3116 2084 3124
rect 2476 3116 2484 3124
rect 2492 3116 2500 3124
rect 2860 3116 2868 3124
rect 3084 3116 3092 3124
rect 3148 3116 3156 3124
rect 3308 3116 3316 3124
rect 3532 3116 3540 3124
rect 3756 3116 3764 3124
rect 3980 3116 3988 3124
rect 4204 3116 4212 3124
rect 4284 3116 4292 3124
rect 4620 3116 4628 3124
rect 4830 3116 4838 3124
rect 5052 3116 5060 3124
rect 5260 3116 5268 3124
rect 5356 3116 5364 3124
rect 5564 3116 5572 3124
rect 5772 3116 5780 3124
rect 6156 3116 6164 3124
rect 6412 3116 6420 3124
rect 6652 3116 6660 3124
rect 6860 3116 6868 3124
rect 7228 3116 7236 3124
rect 7436 3116 7444 3124
rect 7884 3116 7892 3124
rect 8076 3116 8084 3124
rect 8300 3116 8308 3124
rect 8380 3116 8388 3124
rect 8716 3116 8724 3124
rect 9212 3116 9220 3124
rect 9244 3116 9252 3124
rect 9452 3116 9460 3124
rect 9484 3116 9492 3124
rect 9692 3116 9700 3124
rect 10060 3116 10068 3124
rect 188 3076 196 3084
rect 300 3076 308 3084
rect 492 3076 500 3084
rect 524 3076 532 3084
rect 1084 3076 1092 3084
rect 1196 3076 1204 3084
rect 1548 3076 1556 3084
rect 1644 3076 1652 3084
rect 1852 3076 1860 3084
rect 1868 3076 1876 3084
rect 2092 3076 2100 3084
rect 2412 3076 2420 3084
rect 2524 3076 2532 3084
rect 2844 3076 2852 3084
rect 3052 3076 3060 3084
rect 3324 3076 3332 3084
rect 3340 3076 3348 3084
rect 3532 3076 3540 3084
rect 3740 3076 3748 3084
rect 4188 3076 4196 3084
rect 4284 3076 4292 3084
rect 4620 3076 4628 3084
rect 4828 3076 4836 3084
rect 5036 3076 5044 3084
rect 5244 3076 5252 3084
rect 5372 3076 5380 3084
rect 5564 3076 5572 3084
rect 5788 3076 5796 3084
rect 5996 3076 6004 3084
rect 6204 3076 6212 3084
rect 6428 3076 6436 3084
rect 6652 3076 6660 3084
rect 6876 3076 6884 3084
rect 7212 3076 7220 3084
rect 7420 3076 7428 3084
rect 7532 3076 7540 3084
rect 7916 3076 7924 3084
rect 8060 3076 8068 3084
rect 8108 3076 8116 3084
rect 8284 3076 8292 3084
rect 8396 3076 8404 3084
rect 8732 3076 8740 3084
rect 8812 3076 8820 3084
rect 9020 3076 9028 3084
rect 9260 3076 9268 3084
rect 9484 3076 9492 3084
rect 10028 3076 10036 3084
rect 716 3056 724 3064
rect 1388 3056 1396 3064
rect 2044 3056 2052 3064
rect 2668 3056 2676 3064
rect 4652 3056 4660 3064
rect 60 3036 68 3044
rect 940 3036 948 3044
rect 2220 3036 2228 3044
rect 2716 3036 2724 3044
rect 2940 3036 2948 3044
rect 4428 3036 4436 3044
rect 4476 3036 4484 3044
rect 4908 3036 4916 3044
rect 5724 3036 5732 3044
rect 6140 3036 6148 3044
rect 6348 3036 6356 3044
rect 6572 3036 6580 3044
rect 6812 3036 6820 3044
rect 7004 3036 7012 3044
rect 7020 3036 7028 3044
rect 7292 3036 7300 3044
rect 7660 3036 7668 3044
rect 7708 3036 7716 3044
rect 7932 3036 7940 3044
rect 8524 3036 8532 3044
rect 8956 3036 8964 3044
rect 9628 3036 9636 3044
rect 9900 3036 9908 3044
rect 508 2976 516 2984
rect 1164 2976 1172 2984
rect 1324 2976 1332 2984
rect 1548 2976 1556 2984
rect 1788 2976 1796 2984
rect 2236 2976 2244 2984
rect 2460 2976 2468 2984
rect 2540 2976 2548 2984
rect 2716 2976 2724 2984
rect 2924 2976 2932 2984
rect 3164 2976 3172 2984
rect 3372 2976 3380 2984
rect 3868 2976 3876 2984
rect 4524 2976 4532 2984
rect 4700 2976 4708 2984
rect 4748 2976 4756 2984
rect 4988 2976 4996 2984
rect 5644 2976 5652 2984
rect 7404 2976 7412 2984
rect 7420 2976 7428 2984
rect 7788 2976 7796 2984
rect 8236 2976 8244 2984
rect 8460 2976 8468 2984
rect 8716 2976 8724 2984
rect 8732 2976 8740 2984
rect 8988 2976 8996 2984
rect 9228 2976 9236 2984
rect 9836 2976 9844 2984
rect 10060 2976 10068 2984
rect 284 2956 292 2964
rect 4044 2956 4052 2964
rect 5820 2956 5828 2964
rect 92 2936 100 2944
rect 428 2936 436 2944
rect 636 2936 644 2944
rect 732 2936 740 2944
rect 748 2936 756 2944
rect 940 2936 948 2944
rect 1292 2936 1300 2944
rect 1548 2936 1556 2944
rect 1756 2936 1764 2944
rect 1980 2936 1988 2944
rect 2092 2936 2100 2944
rect 2332 2936 2340 2944
rect 2684 2936 2692 2944
rect 2892 2936 2900 2944
rect 3116 2936 3124 2944
rect 3420 2936 3428 2944
rect 3580 2936 3588 2944
rect 3788 2936 3796 2944
rect 4028 2936 4036 2944
rect 4236 2936 4244 2944
rect 4348 2936 4356 2944
rect 4572 2936 4580 2944
rect 4908 2936 4916 2944
rect 5132 2936 5140 2944
rect 5148 2936 5156 2944
rect 5356 2936 5364 2944
rect 5564 2936 5572 2944
rect 5804 2936 5812 2944
rect 6012 2936 6020 2944
rect 6092 2936 6100 2944
rect 6236 2936 6244 2944
rect 6252 2936 6260 2944
rect 6572 2936 6580 2944
rect 6908 2936 6916 2944
rect 7004 2936 7012 2944
rect 7228 2936 7236 2944
rect 7564 2936 7572 2944
rect 7676 2936 7684 2944
rect 8012 2936 8020 2944
rect 8092 2936 8100 2944
rect 8332 2936 8340 2944
rect 8556 2936 8564 2944
rect 8908 2936 8916 2944
rect 9132 2936 9140 2944
rect 9372 2936 9380 2944
rect 9580 2936 9588 2944
rect 9692 2936 9700 2944
rect 9916 2936 9924 2944
rect 76 2916 84 2924
rect 428 2896 436 2904
rect 652 2896 660 2904
rect 732 2896 740 2904
rect 6748 2916 6756 2924
rect 9660 2916 9668 2924
rect 1308 2896 1316 2904
rect 1596 2896 1604 2904
rect 1836 2896 1844 2904
rect 1996 2896 2004 2904
rect 2092 2896 2100 2904
rect 2316 2896 2324 2904
rect 2700 2896 2708 2904
rect 2892 2896 2900 2904
rect 3196 2896 3204 2904
rect 3356 2896 3364 2904
rect 3596 2896 3604 2904
rect 3804 2896 3812 2904
rect 4012 2896 4020 2904
rect 4236 2896 4244 2904
rect 4332 2896 4340 2904
rect 4540 2896 4548 2904
rect 4924 2896 4932 2904
rect 5132 2896 5140 2904
rect 5580 2896 5588 2904
rect 5788 2896 5796 2904
rect 6060 2896 6068 2904
rect 6236 2896 6244 2904
rect 6332 2896 6340 2904
rect 6540 2896 6548 2904
rect 6908 2896 6916 2904
rect 6972 2896 6980 2904
rect 7196 2896 7204 2904
rect 7596 2896 7604 2904
rect 7644 2896 7652 2904
rect 7868 2896 7876 2904
rect 8012 2896 8020 2904
rect 8076 2896 8084 2904
rect 8332 2896 8340 2904
rect 8556 2896 8564 2904
rect 8940 2896 8948 2904
rect 9148 2896 9156 2904
rect 9372 2896 9380 2904
rect 9612 2896 9620 2904
rect 9676 2896 9684 2904
rect 9916 2896 9924 2904
rect 268 2836 276 2844
rect 1100 2836 1108 2844
rect 2236 2836 2244 2844
rect 6492 2836 6500 2844
rect 6748 2836 6756 2844
rect 7164 2836 7172 2844
rect 9436 2836 9444 2844
rect 1836 2776 1844 2784
rect 1852 2776 1860 2784
rect 2332 2776 2340 2784
rect 2988 2776 2996 2784
rect 6444 2776 6452 2784
rect 7100 2776 7108 2784
rect 9916 2776 9924 2784
rect 4092 2756 4100 2764
rect 236 2716 244 2724
rect 460 2716 468 2724
rect 700 2716 708 2724
rect 908 2716 916 2724
rect 1180 2716 1188 2724
rect 1228 2716 1236 2724
rect 1452 2716 1460 2724
rect 1660 2716 1668 2724
rect 2028 2716 2036 2724
rect 2252 2716 2260 2724
rect 2476 2716 2484 2724
rect 2700 2716 2708 2724
rect 2908 2716 2916 2724
rect 3148 2716 3156 2724
rect 3212 2716 3220 2724
rect 3404 2716 3412 2724
rect 3564 2716 3572 2724
rect 3836 2716 3844 2724
rect 4012 2716 4020 2724
rect 4220 2716 4228 2724
rect 4316 2716 4324 2724
rect 4668 2716 4676 2724
rect 4892 2716 4900 2724
rect 4972 2716 4980 2724
rect 5180 2716 5188 2724
rect 5532 2716 5540 2724
rect 5612 2716 5620 2724
rect 6188 2716 6196 2724
rect 6268 2716 6276 2724
rect 6636 2716 6644 2724
rect 6716 2716 6724 2724
rect 6892 2716 6900 2724
rect 7132 2716 7140 2724
rect 7356 2716 7364 2724
rect 7564 2716 7572 2724
rect 7788 2716 7796 2724
rect 8124 2716 8132 2724
rect 8204 2716 8212 2724
rect 8428 2716 8436 2724
rect 8764 2716 8772 2724
rect 8844 2716 8852 2724
rect 9196 2716 9204 2724
rect 9436 2716 9444 2724
rect 9500 2716 9508 2724
rect 9660 2716 9668 2724
rect 9948 2716 9956 2724
rect 10076 2716 10084 2724
rect 6028 2696 6036 2704
rect 9692 2696 9700 2704
rect 204 2676 212 2684
rect 236 2676 244 2684
rect 444 2676 452 2684
rect 460 2676 468 2684
rect 668 2676 676 2684
rect 700 2676 708 2684
rect 1132 2676 1140 2684
rect 1244 2676 1252 2684
rect 1420 2676 1428 2684
rect 1692 2676 1700 2684
rect 2012 2676 2020 2684
rect 2252 2676 2260 2684
rect 2460 2676 2468 2684
rect 2748 2676 2756 2684
rect 2892 2676 2900 2684
rect 3100 2676 3108 2684
rect 3212 2676 3220 2684
rect 3564 2676 3572 2684
rect 3788 2676 3796 2684
rect 3996 2676 4004 2684
rect 4204 2676 4212 2684
rect 4316 2676 4324 2684
rect 4668 2676 4676 2684
rect 4876 2676 4884 2684
rect 4972 2676 4980 2684
rect 5196 2676 5204 2684
rect 5516 2676 5524 2684
rect 5628 2676 5636 2684
rect 5836 2676 5844 2684
rect 6188 2676 6196 2684
rect 6268 2676 6276 2684
rect 6620 2676 6628 2684
rect 6652 2676 6660 2684
rect 6940 2676 6948 2684
rect 7148 2676 7156 2684
rect 7580 2676 7588 2684
rect 8108 2676 8116 2684
rect 8236 2676 8244 2684
rect 8444 2676 8452 2684
rect 8572 2676 8580 2684
rect 8620 2676 8628 2684
rect 8748 2676 8756 2684
rect 8860 2676 8868 2684
rect 9196 2676 9204 2684
rect 9212 2676 9220 2684
rect 9388 2676 9396 2684
rect 9516 2676 9524 2684
rect 9724 2676 9732 2684
rect 9948 2676 9956 2684
rect 1660 2656 1668 2664
rect 2492 2656 2500 2664
rect 3868 2656 3876 2664
rect 60 2636 68 2644
rect 1356 2636 1364 2644
rect 2076 2636 2084 2644
rect 2748 2636 2756 2644
rect 3420 2636 3428 2644
rect 3644 2636 3652 2644
rect 4476 2636 4484 2644
rect 4508 2636 4516 2644
rect 4748 2636 4756 2644
rect 5148 2636 5156 2644
rect 5324 2636 5332 2644
rect 5388 2636 5396 2644
rect 5980 2636 5988 2644
rect 6476 2636 6484 2644
rect 6876 2636 6884 2644
rect 7500 2636 7508 2644
rect 7932 2636 7940 2644
rect 7980 2636 7988 2644
rect 8348 2636 8356 2644
rect 9004 2636 9012 2644
rect 9052 2636 9060 2644
rect 236 2576 244 2584
rect 252 2576 260 2584
rect 700 2576 708 2584
rect 940 2576 948 2584
rect 1132 2576 1140 2584
rect 1340 2576 1348 2584
rect 1596 2576 1604 2584
rect 1658 2576 1666 2584
rect 2092 2576 2100 2584
rect 2940 2576 2948 2584
rect 3196 2576 3204 2584
rect 3436 2576 3444 2584
rect 3660 2576 3668 2584
rect 3868 2576 3876 2584
rect 5484 2576 5492 2584
rect 5900 2576 5908 2584
rect 6556 2576 6564 2584
rect 6620 2576 6628 2584
rect 6828 2576 6836 2584
rect 7004 2576 7012 2584
rect 7500 2576 7508 2584
rect 7660 2576 7668 2584
rect 8108 2576 8116 2584
rect 8764 2576 8772 2584
rect 9150 2576 9158 2584
rect 9388 2576 9396 2584
rect 9852 2576 9860 2584
rect 10076 2576 10084 2584
rect 4092 2556 4100 2564
rect 4620 2556 4628 2564
rect 7212 2556 7220 2564
rect 7884 2556 7892 2564
rect 8508 2556 8516 2564
rect 8940 2556 8948 2564
rect 92 2536 100 2544
rect 444 2536 452 2544
rect 556 2536 564 2544
rect 780 2536 788 2544
rect 1004 2536 1012 2544
rect 1228 2536 1236 2544
rect 1420 2536 1428 2544
rect 1788 2536 1796 2544
rect 1820 2536 1828 2544
rect 2012 2536 2020 2544
rect 2220 2536 2228 2544
rect 2348 2536 2356 2544
rect 2492 2536 2500 2544
rect 2764 2536 2772 2544
rect 2796 2536 2804 2544
rect 3036 2536 3044 2544
rect 3372 2536 3380 2544
rect 3612 2536 3620 2544
rect 3836 2536 3844 2544
rect 4076 2536 4084 2544
rect 4300 2536 4308 2544
rect 4380 2536 4388 2544
rect 4556 2536 4564 2544
rect 4764 2536 4772 2544
rect 4972 2536 4980 2544
rect 5084 2536 5092 2544
rect 5324 2536 5332 2544
rect 5548 2536 5556 2544
rect 5756 2536 5764 2544
rect 5980 2536 5988 2544
rect 6204 2536 6212 2544
rect 6748 2536 6756 2544
rect 6956 2536 6964 2544
rect 7196 2536 7204 2544
rect 7404 2536 7412 2544
rect 7644 2536 7652 2544
rect 7852 2536 7860 2544
rect 8076 2536 8084 2544
rect 8284 2536 8292 2544
rect 8396 2536 8404 2544
rect 8588 2536 8596 2544
rect 8812 2536 8820 2544
rect 9004 2536 9012 2544
rect 9244 2536 9252 2544
rect 9596 2536 9604 2544
rect 9708 2536 9716 2544
rect 9884 2536 9892 2544
rect 60 2496 68 2504
rect 444 2496 452 2504
rect 492 2496 500 2504
rect 700 2496 708 2504
rect 988 2496 996 2504
rect 1212 2496 1220 2504
rect 1436 2496 1444 2504
rect 1804 2496 1812 2504
rect 2044 2496 2052 2504
rect 2236 2496 2244 2504
rect 2332 2496 2340 2504
rect 2540 2496 2548 2504
rect 2748 2496 2756 2504
rect 2796 2496 2804 2504
rect 3020 2496 3028 2504
rect 3388 2496 3396 2504
rect 3628 2496 3636 2504
rect 3884 2496 3892 2504
rect 4108 2496 4116 2504
rect 4316 2496 4324 2504
rect 4540 2496 4548 2504
rect 4974 2496 4982 2504
rect 5084 2496 5092 2504
rect 5532 2496 5540 2504
rect 5964 2496 5972 2504
rect 6188 2496 6196 2504
rect 6396 2496 6404 2504
rect 6780 2496 6788 2504
rect 6972 2496 6980 2504
rect 7180 2496 7188 2504
rect 7420 2496 7428 2504
rect 7644 2496 7652 2504
rect 7884 2496 7892 2504
rect 8076 2496 8084 2504
rect 8284 2496 8292 2504
rect 8380 2496 8388 2504
rect 8588 2496 8596 2504
rect 8780 2496 8788 2504
rect 9020 2496 9028 2504
rect 9244 2496 9252 2504
rect 9596 2496 9604 2504
rect 9692 2496 9700 2504
rect 9868 2496 9876 2504
rect 5308 2476 5316 2484
rect 1132 2436 1140 2444
rect 3164 2436 3172 2444
rect 6108 2436 6116 2444
rect 9468 2436 9476 2444
rect 508 2376 516 2384
rect 2284 2376 2292 2384
rect 7276 2376 7284 2384
rect 8124 2376 8132 2384
rect 8764 2376 8772 2384
rect 4700 2356 4708 2364
rect 4236 2336 4244 2344
rect 5276 2336 5284 2344
rect 7980 2336 7988 2344
rect 204 2316 212 2324
rect 492 2316 500 2324
rect 652 2316 660 2324
rect 876 2316 884 2324
rect 1324 2316 1332 2324
rect 1596 2316 1604 2324
rect 1772 2316 1780 2324
rect 2012 2316 2020 2324
rect 2204 2316 2212 2324
rect 2428 2316 2436 2324
rect 2508 2316 2516 2324
rect 2860 2316 2868 2324
rect 3100 2316 3108 2324
rect 3164 2316 3172 2324
rect 3500 2316 3508 2324
rect 3724 2316 3732 2324
rect 3932 2316 3940 2324
rect 4028 2316 4036 2324
rect 4396 2316 4404 2324
rect 4492 2316 4500 2324
rect 4860 2316 4868 2324
rect 4924 2316 4932 2324
rect 5132 2316 5140 2324
rect 5292 2316 5300 2324
rect 5516 2316 5524 2324
rect 5788 2316 5796 2324
rect 6028 2316 6036 2324
rect 6252 2316 6260 2324
rect 6476 2316 6484 2324
rect 6700 2316 6708 2324
rect 6908 2316 6916 2324
rect 7132 2316 7140 2324
rect 7340 2316 7348 2324
rect 7772 2316 7780 2324
rect 7964 2316 7972 2324
rect 8332 2316 8340 2324
rect 8412 2316 8420 2324
rect 8620 2316 8628 2324
rect 8844 2316 8852 2324
rect 9180 2316 9188 2324
rect 9274 2316 9282 2324
rect 9612 2316 9620 2324
rect 9820 2316 9828 2324
rect 9900 2316 9908 2324
rect 492 2276 500 2284
rect 652 2276 660 2284
rect 684 2276 692 2284
rect 876 2276 884 2284
rect 1100 2276 1108 2284
rect 1308 2276 1316 2284
rect 1548 2276 1556 2284
rect 1756 2276 1764 2284
rect 1980 2276 1988 2284
rect 2188 2276 2196 2284
rect 2412 2276 2420 2284
rect 2524 2276 2532 2284
rect 2876 2276 2884 2284
rect 3068 2276 3076 2284
rect 3180 2276 3188 2284
rect 3484 2276 3492 2284
rect 3788 2276 3796 2284
rect 3932 2276 3940 2284
rect 4044 2276 4052 2284
rect 4396 2276 4404 2284
rect 4412 2276 4420 2284
rect 4812 2276 4820 2284
rect 4860 2276 4868 2284
rect 4940 2276 4948 2284
rect 5148 2276 5156 2284
rect 5356 2276 5364 2284
rect 5804 2276 5812 2284
rect 6028 2276 6036 2284
rect 6236 2276 6244 2284
rect 6700 2276 6708 2284
rect 6892 2276 6900 2284
rect 6924 2276 6932 2284
rect 7132 2276 7140 2284
rect 7356 2276 7364 2284
rect 7564 2276 7572 2284
rect 7788 2276 7796 2284
rect 7996 2276 8004 2284
rect 8316 2276 8324 2284
rect 8396 2276 8404 2284
rect 8636 2276 8644 2284
rect 8780 2276 8788 2284
rect 8988 2276 8996 2284
rect 9164 2276 9172 2284
rect 9276 2276 9284 2284
rect 9596 2276 9604 2284
rect 9820 2276 9828 2284
rect 9916 2276 9924 2284
rect 3308 2256 3316 2264
rect 3370 2256 3378 2264
rect 8604 2256 8612 2264
rect 60 2236 68 2244
rect 956 2236 964 2244
rect 1388 2236 1396 2244
rect 1626 2236 1634 2244
rect 1852 2236 1860 2244
rect 2060 2236 2068 2244
rect 2284 2236 2292 2244
rect 2668 2236 2676 2244
rect 2716 2236 2724 2244
rect 2940 2236 2948 2244
rect 3580 2236 3588 2244
rect 4188 2236 4196 2244
rect 4636 2236 4644 2244
rect 5068 2236 5076 2244
rect 5724 2236 5732 2244
rect 5948 2236 5956 2244
rect 6172 2236 6180 2244
rect 6620 2236 6628 2244
rect 7068 2236 7076 2244
rect 7708 2236 7716 2244
rect 8172 2236 8180 2244
rect 9036 2236 9044 2244
rect 9420 2236 9428 2244
rect 9452 2236 9460 2244
rect 9676 2236 9684 2244
rect 10060 2236 10068 2244
rect 236 2176 244 2184
rect 460 2176 468 2184
rect 716 2176 724 2184
rect 1180 2176 1188 2184
rect 1804 2176 1812 2184
rect 2092 2176 2100 2184
rect 2492 2176 2500 2184
rect 3420 2176 3428 2184
rect 3628 2176 3636 2184
rect 4060 2176 4068 2184
rect 4076 2176 4084 2184
rect 4940 2176 4948 2184
rect 4972 2176 4980 2184
rect 5484 2176 5492 2184
rect 5868 2176 5876 2184
rect 6524 2176 6532 2184
rect 6972 2176 6980 2184
rect 7180 2176 7188 2184
rect 7406 2176 7414 2184
rect 7660 2176 7668 2184
rect 7852 2176 7860 2184
rect 8060 2176 8068 2184
rect 8300 2176 8308 2184
rect 8492 2176 8500 2184
rect 8556 2176 8564 2184
rect 10236 2176 10244 2184
rect 524 2156 532 2164
rect 92 2136 100 2144
rect 316 2136 324 2144
rect 652 2136 660 2144
rect 956 2136 964 2144
rect 972 2136 980 2144
rect 1292 2136 1300 2144
rect 1772 2136 1780 2144
rect 1996 2136 2004 2144
rect 2428 2136 2436 2144
rect 2908 2136 2916 2144
rect 3020 2136 3028 2144
rect 3596 2136 3604 2144
rect 3820 2136 3828 2144
rect 3932 2136 3940 2144
rect 4268 2136 4276 2144
rect 4300 2136 4308 2144
rect 4492 2136 4500 2144
rect 4572 2136 4580 2144
rect 4812 2136 4820 2144
rect 6364 2156 6372 2164
rect 8924 2156 8932 2164
rect 5388 2136 5396 2144
rect 5612 2136 5620 2144
rect 5724 2136 5732 2144
rect 5964 2136 5972 2144
rect 6380 2136 6388 2144
rect 6620 2136 6628 2144
rect 7052 2136 7060 2144
rect 7276 2136 7284 2144
rect 7484 2136 7492 2144
rect 7708 2136 7716 2144
rect 7932 2136 7940 2144
rect 8124 2136 8132 2144
rect 8364 2136 8372 2144
rect 8684 2136 8692 2144
rect 8796 2136 8804 2144
rect 8988 2136 8996 2144
rect 9132 2136 9140 2144
rect 9244 2136 9252 2144
rect 9468 2136 9476 2144
rect 9676 2136 9684 2144
rect 9884 2136 9892 2144
rect 10108 2136 10116 2144
rect 60 2116 68 2124
rect 1836 2116 1844 2124
rect 300 2096 308 2104
rect 668 2096 676 2104
rect 892 2096 900 2104
rect 956 2096 964 2104
rect 1324 2096 1332 2104
rect 1548 2096 1556 2104
rect 2044 2096 2052 2104
rect 2060 2096 2068 2104
rect 2284 2096 2292 2104
rect 2316 2096 2324 2104
rect 2476 2096 2484 2104
rect 2684 2096 2692 2104
rect 2908 2096 2916 2104
rect 3004 2096 3012 2104
rect 3244 2096 3252 2104
rect 3628 2096 3636 2104
rect 3852 2096 3860 2104
rect 3916 2096 3924 2104
rect 4300 2096 4308 2104
rect 4492 2096 4500 2104
rect 4572 2096 4580 2104
rect 5164 2096 5172 2104
rect 5420 2096 5428 2104
rect 5644 2096 5652 2104
rect 5724 2096 5732 2104
rect 5884 2096 5892 2104
rect 6156 2096 6164 2104
rect 6380 2096 6388 2104
rect 6588 2096 6596 2104
rect 6812 2096 6820 2104
rect 7036 2096 7044 2104
rect 7260 2096 7268 2104
rect 7484 2096 7492 2104
rect 7692 2096 7700 2104
rect 7916 2096 7924 2104
rect 8124 2096 8132 2104
rect 8364 2096 8372 2104
rect 8700 2096 8708 2104
rect 8764 2096 8772 2104
rect 9148 2096 9156 2104
rect 9180 2096 9188 2104
rect 9466 2096 9474 2104
rect 1164 2076 1172 2084
rect 1388 2036 1396 2044
rect 3388 2036 3396 2044
rect 508 1976 516 1984
rect 5884 1976 5892 1984
rect 6956 1976 6964 1984
rect 7388 1976 7396 1984
rect 8284 1976 8292 1984
rect 8492 1976 8500 1984
rect 2014 1956 2022 1964
rect 6108 1936 6116 1944
rect 6956 1936 6964 1944
rect 7020 1936 7028 1944
rect 7180 1936 7188 1944
rect 7244 1936 7252 1944
rect 7404 1936 7412 1944
rect 204 1916 212 1924
rect 284 1916 292 1924
rect 652 1916 660 1924
rect 860 1916 868 1924
rect 956 1916 964 1924
rect 1340 1916 1348 1924
rect 1388 1916 1396 1924
rect 1788 1916 1796 1924
rect 1884 1916 1892 1924
rect 2236 1916 2244 1924
rect 2330 1916 2338 1924
rect 2700 1916 2708 1924
rect 2780 1916 2788 1924
rect 3004 1916 3012 1924
rect 3372 1916 3380 1924
rect 3628 1916 3636 1924
rect 3852 1916 3860 1924
rect 4076 1916 4084 1924
rect 4284 1916 4292 1924
rect 4492 1916 4500 1924
rect 4732 1916 4740 1924
rect 4748 1916 4756 1924
rect 5020 1916 5028 1924
rect 5180 1916 5188 1924
rect 5228 1916 5236 1924
rect 5708 1916 5716 1924
rect 5916 1916 5924 1924
rect 6284 1916 6292 1924
rect 6702 1916 6710 1924
rect 6796 1916 6804 1924
rect 6972 1916 6980 1924
rect 7180 1916 7188 1924
rect 7660 1916 7668 1924
rect 7884 1916 7892 1924
rect 8124 1916 8132 1924
rect 8348 1916 8356 1924
rect 8588 1916 8596 1924
rect 8796 1916 8804 1924
rect 8988 1916 8996 1924
rect 9148 1916 9156 1924
rect 9244 1916 9252 1924
rect 9628 1916 9636 1924
rect 9676 1916 9684 1924
rect 9884 1916 9892 1924
rect 300 1876 308 1884
rect 636 1876 644 1884
rect 860 1876 868 1884
rect 956 1876 964 1884
rect 1308 1876 1316 1884
rect 1420 1876 1428 1884
rect 1772 1876 1780 1884
rect 1788 1876 1796 1884
rect 1868 1876 1876 1884
rect 1884 1876 1892 1884
rect 2268 1876 2276 1884
rect 2684 1876 2692 1884
rect 2716 1876 2724 1884
rect 3020 1876 3028 1884
rect 3372 1876 3380 1884
rect 3596 1876 3604 1884
rect 3820 1876 3828 1884
rect 3852 1876 3860 1884
rect 4076 1876 4084 1884
rect 4268 1876 4276 1884
rect 4476 1876 4484 1884
rect 4716 1876 4724 1884
rect 4812 1876 4820 1884
rect 5020 1876 5028 1884
rect 5260 1876 5268 1884
rect 5484 1876 5492 1884
rect 5708 1876 5716 1884
rect 5932 1876 5940 1884
rect 6268 1876 6276 1884
rect 6284 1876 6292 1884
rect 6492 1876 6500 1884
rect 6684 1876 6692 1884
rect 6812 1876 6820 1884
rect 7036 1876 7044 1884
rect 7468 1876 7476 1884
rect 7676 1876 7684 1884
rect 7900 1876 7908 1884
rect 8124 1876 8132 1884
rect 8364 1876 8372 1884
rect 8572 1876 8580 1884
rect 8812 1876 8820 1884
rect 9132 1876 9140 1884
rect 9244 1876 9252 1884
rect 9420 1876 9428 1884
rect 9564 1876 9572 1884
rect 9660 1876 9668 1884
rect 10108 1876 10116 1884
rect 1164 1856 1172 1864
rect 1612 1856 1620 1864
rect 2476 1856 2484 1864
rect 2972 1856 2980 1864
rect 3180 1856 3188 1864
rect 60 1836 68 1844
rect 428 1836 436 1844
rect 716 1836 724 1844
rect 1180 1836 1188 1844
rect 1580 1836 1588 1844
rect 2092 1836 2100 1844
rect 2460 1836 2468 1844
rect 3228 1836 3236 1844
rect 3436 1836 3444 1844
rect 3676 1836 3684 1844
rect 4140 1836 4148 1844
rect 4300 1836 4308 1844
rect 4524 1836 4532 1844
rect 4940 1836 4948 1844
rect 5164 1836 5172 1844
rect 5628 1836 5636 1844
rect 6076 1836 6084 1844
rect 6956 1836 6964 1844
rect 7596 1836 7604 1844
rect 7804 1836 7812 1844
rect 8044 1836 8052 1844
rect 8268 1836 8276 1844
rect 8540 1836 8548 1844
rect 8748 1836 8756 1844
rect 8956 1836 8964 1844
rect 9436 1836 9444 1844
rect 10252 1836 10260 1844
rect 222 1776 230 1784
rect 252 1776 260 1784
rect 1116 1776 1124 1784
rect 1340 1776 1348 1784
rect 1628 1776 1636 1784
rect 1644 1776 1652 1784
rect 1884 1776 1892 1784
rect 2940 1776 2948 1784
rect 3212 1776 3220 1784
rect 3628 1776 3636 1784
rect 3836 1776 3844 1784
rect 4076 1776 4084 1784
rect 4092 1776 4100 1784
rect 4700 1776 4708 1784
rect 4956 1776 4964 1784
rect 5820 1776 5828 1784
rect 6284 1776 6292 1784
rect 6972 1776 6980 1784
rect 7180 1776 7188 1784
rect 7212 1776 7220 1784
rect 7644 1776 7652 1784
rect 7676 1776 7684 1784
rect 8316 1776 8324 1784
rect 8940 1776 8948 1784
rect 9804 1776 9812 1784
rect 10220 1776 10228 1784
rect 3212 1756 3220 1764
rect 92 1736 100 1744
rect 444 1736 452 1744
rect 524 1736 532 1744
rect 652 1736 660 1744
rect 764 1736 772 1744
rect 1212 1736 1220 1744
rect 1436 1736 1444 1744
rect 1788 1736 1796 1744
rect 2012 1736 2020 1744
rect 2044 1736 2052 1744
rect 2252 1736 2260 1744
rect 2268 1736 2276 1744
rect 2476 1736 2484 1744
rect 2700 1736 2708 1744
rect 2796 1736 2804 1744
rect 3036 1736 3044 1744
rect 3404 1736 3412 1744
rect 3484 1736 3492 1744
rect 3692 1736 3700 1744
rect 3900 1736 3908 1744
rect 4252 1736 4260 1744
rect 4460 1736 4468 1744
rect 4556 1736 4564 1744
rect 4796 1736 4804 1744
rect 4988 1736 4996 1744
rect 5148 1736 5156 1744
rect 5260 1736 5268 1744
rect 5484 1736 5492 1744
rect 5676 1736 5684 1744
rect 5900 1736 5908 1744
rect 6124 1736 6132 1744
rect 6284 1736 6292 1744
rect 6444 1736 6452 1744
rect 6684 1736 6692 1744
rect 6780 1736 6788 1744
rect 6796 1736 6804 1744
rect 7020 1736 7028 1744
rect 7340 1736 7348 1744
rect 7452 1736 7460 1744
rect 7804 1736 7812 1744
rect 7916 1736 7924 1744
rect 8140 1736 8148 1744
rect 8380 1736 8388 1744
rect 9020 1736 9028 1744
rect 9452 1736 9460 1744
rect 9612 1736 9620 1744
rect 9868 1736 9876 1744
rect 76 1716 84 1724
rect 7836 1716 7844 1724
rect 444 1696 452 1704
rect 668 1696 676 1704
rect 748 1696 756 1704
rect 924 1696 932 1704
rect 1212 1696 1220 1704
rect 1404 1696 1412 1704
rect 1868 1696 1876 1704
rect 2028 1696 2036 1704
rect 2268 1696 2276 1704
rect 2700 1696 2708 1704
rect 2796 1696 2804 1704
rect 3020 1696 3028 1704
rect 3372 1696 3380 1704
rect 3468 1696 3476 1704
rect 3692 1696 3700 1704
rect 3900 1696 3908 1704
rect 4476 1696 4484 1704
rect 4540 1696 4548 1704
rect 4796 1696 4804 1704
rect 5164 1696 5172 1704
rect 5180 1696 5188 1704
rect 5884 1696 5892 1704
rect 6492 1696 6500 1704
rect 6700 1696 6708 1704
rect 6780 1696 6788 1704
rect 6988 1696 6996 1704
rect 7372 1696 7380 1704
rect 7452 1696 7460 1704
rect 7804 1696 7812 1704
rect 8140 1696 8148 1704
rect 8300 1696 8308 1704
rect 8588 1696 8596 1704
rect 8748 1696 8756 1704
rect 8956 1696 8964 1704
rect 9228 1696 9236 1704
rect 9868 1696 9876 1704
rect 10076 1696 10084 1704
rect 940 1656 948 1664
rect 6444 1656 6452 1664
rect 8060 1636 8068 1644
rect 1116 1576 1124 1584
rect 1404 1576 1412 1584
rect 4764 1576 4772 1584
rect 4924 1576 4932 1584
rect 5180 1576 5188 1584
rect 5210 1576 5218 1584
rect 6044 1576 6052 1584
rect 6492 1576 6500 1584
rect 284 1556 292 1564
rect 220 1516 228 1524
rect 428 1516 436 1524
rect 524 1516 532 1524
rect 748 1516 756 1524
rect 972 1516 980 1524
rect 1548 1516 1556 1524
rect 1628 1516 1636 1524
rect 1836 1516 1844 1524
rect 2092 1516 2100 1524
rect 2330 1516 2338 1524
rect 2540 1516 2548 1524
rect 2940 1516 2948 1524
rect 3148 1516 3156 1524
rect 3372 1516 3380 1524
rect 3660 1516 3668 1524
rect 3868 1516 3876 1524
rect 3916 1516 3924 1524
rect 4076 1516 4084 1524
rect 4492 1516 4500 1524
rect 4572 1516 4580 1524
rect 4780 1516 4788 1524
rect 5004 1516 5012 1524
rect 5356 1516 5364 1524
rect 5596 1516 5604 1524
rect 5788 1516 5796 1524
rect 5884 1516 5892 1524
rect 6236 1516 6244 1524
rect 6476 1516 6484 1524
rect 6700 1516 6708 1524
rect 6780 1516 6788 1524
rect 6956 1516 6964 1524
rect 7244 1516 7252 1524
rect 7468 1516 7476 1524
rect 8044 1516 8052 1524
rect 8252 1516 8260 1524
rect 8460 1516 8468 1524
rect 8540 1516 8548 1524
rect 8892 1516 8900 1524
rect 9324 1516 9332 1524
rect 9404 1516 9412 1524
rect 9756 1516 9764 1524
rect 9820 1516 9828 1524
rect 10060 1516 10068 1524
rect 924 1496 932 1504
rect 8972 1496 8980 1504
rect 9980 1496 9988 1504
rect 204 1476 212 1484
rect 428 1476 436 1484
rect 540 1476 548 1484
rect 764 1476 772 1484
rect 972 1476 980 1484
rect 1148 1476 1156 1484
rect 1324 1476 1332 1484
rect 1612 1476 1620 1484
rect 1644 1476 1652 1484
rect 1852 1476 1860 1484
rect 1868 1476 1876 1484
rect 2300 1476 2308 1484
rect 2332 1476 2340 1484
rect 2540 1476 2548 1484
rect 2556 1476 2564 1484
rect 2908 1476 2916 1484
rect 2924 1476 2932 1484
rect 3132 1476 3140 1484
rect 3164 1476 3172 1484
rect 3436 1476 3444 1484
rect 3452 1476 3460 1484
rect 3596 1476 3604 1484
rect 3820 1476 3828 1484
rect 3932 1476 3940 1484
rect 4156 1476 4164 1484
rect 4476 1476 4484 1484
rect 4588 1476 4596 1484
rect 4812 1476 4820 1484
rect 5020 1476 5028 1484
rect 5340 1476 5348 1484
rect 5356 1476 5364 1484
rect 5564 1476 5572 1484
rect 5596 1476 5604 1484
rect 5788 1476 5796 1484
rect 5900 1476 5908 1484
rect 6460 1476 6468 1484
rect 6684 1476 6692 1484
rect 6796 1476 6804 1484
rect 7020 1476 7028 1484
rect 7244 1476 7252 1484
rect 7468 1476 7476 1484
rect 7692 1476 7700 1484
rect 8012 1476 8020 1484
rect 8236 1476 8244 1484
rect 8252 1476 8260 1484
rect 8444 1476 8452 1484
rect 8508 1476 8516 1484
rect 8940 1476 8948 1484
rect 8988 1476 8996 1484
rect 9308 1476 9316 1484
rect 9420 1476 9428 1484
rect 9596 1476 9604 1484
rect 9740 1476 9748 1484
rect 9772 1476 9780 1484
rect 7868 1456 7876 1464
rect 9564 1456 9572 1464
rect 60 1436 68 1444
rect 668 1436 676 1444
rect 2044 1436 2052 1444
rect 2700 1436 2708 1444
rect 2716 1436 2724 1444
rect 3628 1436 3636 1444
rect 4060 1436 4068 1444
rect 4284 1436 4292 1444
rect 4300 1436 4308 1444
rect 6092 1436 6100 1444
rect 6924 1436 6932 1444
rect 7164 1436 7172 1444
rect 7404 1436 7412 1444
rect 7868 1436 7876 1444
rect 8092 1436 8100 1444
rect 8700 1436 8708 1444
rect 8732 1436 8740 1444
rect 9132 1436 9140 1444
rect 9180 1436 9188 1444
rect 10188 1436 10196 1444
rect 668 1376 676 1384
rect 1116 1376 1124 1384
rect 1372 1376 1380 1384
rect 1836 1376 1844 1384
rect 2252 1376 2260 1384
rect 2316 1376 2324 1384
rect 2700 1376 2708 1384
rect 2908 1376 2916 1384
rect 3388 1376 3396 1384
rect 3418 1376 3426 1384
rect 3644 1376 3652 1384
rect 4316 1376 4324 1384
rect 4540 1376 4548 1384
rect 4764 1376 4772 1384
rect 5148 1376 5156 1384
rect 5372 1376 5380 1384
rect 5644 1376 5652 1384
rect 5660 1376 5668 1384
rect 6508 1376 6516 1384
rect 6716 1376 6724 1384
rect 6940 1376 6948 1384
rect 7388 1376 7396 1384
rect 7852 1376 7860 1384
rect 8508 1376 8516 1384
rect 8524 1376 8532 1384
rect 9164 1376 9172 1384
rect 9596 1376 9604 1384
rect 9852 1376 9860 1384
rect 3804 1356 3812 1364
rect 92 1336 100 1344
rect 316 1336 324 1344
rect 540 1336 548 1344
rect 732 1336 740 1344
rect 876 1336 884 1344
rect 924 1336 932 1344
rect 1212 1336 1220 1344
rect 1580 1336 1588 1344
rect 1676 1336 1684 1344
rect 2012 1336 2020 1344
rect 2108 1336 2116 1344
rect 2444 1336 2452 1344
rect 2556 1336 2564 1344
rect 2780 1336 2788 1344
rect 2988 1336 2996 1344
rect 3196 1336 3204 1344
rect 3532 1336 3540 1344
rect 3772 1336 3780 1344
rect 4060 1336 4068 1344
rect 4236 1336 4244 1344
rect 4460 1336 4468 1344
rect 4668 1336 4676 1344
rect 5020 1336 5028 1344
rect 5228 1336 5236 1344
rect 5452 1336 5460 1344
rect 5804 1336 5812 1344
rect 5916 1336 5924 1344
rect 6092 1336 6100 1344
rect 6348 1336 6356 1344
rect 6572 1336 6580 1344
rect 6796 1336 6804 1344
rect 7036 1336 7044 1344
rect 7180 1336 7188 1344
rect 7596 1336 7604 1344
rect 7692 1336 7700 1344
rect 7916 1336 7924 1344
rect 8364 1336 8372 1344
rect 8684 1336 8692 1344
rect 8812 1336 8820 1344
rect 9244 1336 9252 1344
rect 9692 1336 9700 1344
rect 9868 1336 9876 1344
rect 10012 1336 10020 1344
rect 92 1296 100 1304
rect 300 1296 308 1304
rect 876 1296 884 1304
rect 972 1296 980 1304
rect 1196 1296 1204 1304
rect 1564 1296 1572 1304
rect 1660 1296 1668 1304
rect 2028 1296 2036 1304
rect 2044 1296 2052 1304
rect 2108 1296 2116 1304
rect 2476 1296 2484 1304
rect 2556 1296 2564 1304
rect 2764 1296 2772 1304
rect 2972 1296 2980 1304
rect 3148 1296 3156 1304
rect 3564 1296 3572 1304
rect 3804 1296 3812 1304
rect 4044 1296 4052 1304
rect 4284 1296 4292 1304
rect 4524 1296 4532 1304
rect 4684 1296 4692 1304
rect 4924 1296 4932 1304
rect 5004 1296 5012 1304
rect 5212 1296 5220 1304
rect 5452 1296 5460 1304
rect 5804 1296 5812 1304
rect 5900 1296 5908 1304
rect 6348 1296 6356 1304
rect 6540 1296 6548 1304
rect 6796 1296 6804 1304
rect 7004 1296 7012 1304
rect 7596 1296 7604 1304
rect 7660 1296 7668 1304
rect 7900 1296 7908 1304
rect 8124 1296 8132 1304
rect 8348 1296 8356 1304
rect 3116 1276 3124 1284
rect 8780 1296 8788 1304
rect 9004 1296 9012 1304
rect 9244 1296 9252 1304
rect 9404 1296 9412 1304
rect 9676 1296 9684 1304
rect 10028 1296 10036 1304
rect 8796 1276 8804 1284
rect 6268 1256 6276 1264
rect 236 1236 244 1244
rect 1356 1236 1364 1244
rect 1836 1236 1844 1244
rect 4060 1236 4068 1244
rect 7452 1236 7460 1244
rect 8268 1236 8276 1244
rect 76 1176 84 1184
rect 892 1176 900 1184
rect 3774 1176 3782 1184
rect 3852 1176 3860 1184
rect 4076 1176 4084 1184
rect 4908 1176 4916 1184
rect 5164 1176 5172 1184
rect 6060 1176 6068 1184
rect 6300 1176 6308 1184
rect 6556 1176 6564 1184
rect 6812 1176 6820 1184
rect 10060 1176 10068 1184
rect 5164 1156 5172 1164
rect 1564 1136 1572 1144
rect 5916 1136 5924 1144
rect 220 1116 228 1124
rect 444 1116 452 1124
rect 684 1116 692 1124
rect 748 1116 756 1124
rect 908 1116 916 1124
rect 940 1116 948 1124
rect 1116 1116 1124 1124
rect 1356 1116 1364 1124
rect 1836 1116 1844 1124
rect 2012 1116 2020 1124
rect 2092 1116 2100 1124
rect 2476 1116 2484 1124
rect 2668 1116 2676 1124
rect 2876 1116 2884 1124
rect 3164 1116 3172 1124
rect 3324 1116 3332 1124
rect 3404 1116 3412 1124
rect 3628 1116 3636 1124
rect 4012 1116 4020 1124
rect 4204 1116 4212 1124
rect 4236 1116 4244 1124
rect 4444 1116 4452 1124
rect 4524 1116 4532 1124
rect 4780 1116 4788 1124
rect 5004 1116 5012 1124
rect 5356 1116 5364 1124
rect 5452 1116 5460 1124
rect 5692 1116 5700 1124
rect 6140 1116 6148 1124
rect 6380 1116 6388 1124
rect 6620 1116 6628 1124
rect 6956 1116 6964 1124
rect 7036 1116 7044 1124
rect 7452 1116 7460 1124
rect 7484 1116 7492 1124
rect 7706 1116 7714 1124
rect 8060 1116 8068 1124
rect 8268 1116 8276 1124
rect 8492 1116 8500 1124
rect 8700 1116 8708 1124
rect 8924 1116 8932 1124
rect 9180 1116 9188 1124
rect 9244 1116 9252 1124
rect 9820 1116 9828 1124
rect 9916 1116 9924 1124
rect 940 1096 948 1104
rect 1164 1096 1172 1104
rect 1388 1096 1396 1104
rect 4684 1096 4692 1104
rect 204 1076 212 1084
rect 236 1076 244 1084
rect 460 1076 468 1084
rect 652 1076 660 1084
rect 764 1076 772 1084
rect 956 1076 964 1084
rect 972 1076 980 1084
rect 1196 1076 1204 1084
rect 1356 1076 1364 1084
rect 1772 1076 1780 1084
rect 1820 1076 1828 1084
rect 1996 1076 2004 1084
rect 2108 1076 2116 1084
rect 2444 1076 2452 1084
rect 2476 1076 2484 1084
rect 2668 1076 2676 1084
rect 2892 1076 2900 1084
rect 3084 1076 3092 1084
rect 3340 1076 3348 1084
rect 3420 1076 3428 1084
rect 3644 1076 3652 1084
rect 3996 1076 4004 1084
rect 4188 1076 4196 1084
rect 4428 1076 4436 1084
rect 4460 1076 4468 1084
rect 4556 1076 4564 1084
rect 4796 1076 4804 1084
rect 5020 1076 5028 1084
rect 5356 1076 5364 1084
rect 5468 1076 5476 1084
rect 5900 1076 5908 1084
rect 5932 1076 5940 1084
rect 6076 1076 6084 1084
rect 6140 1076 6148 1084
rect 6156 1076 6164 1084
rect 6316 1076 6324 1084
rect 6620 1076 6628 1084
rect 6956 1076 6964 1084
rect 7068 1076 7076 1084
rect 7388 1076 7396 1084
rect 7708 1076 7716 1084
rect 8236 1076 8244 1084
rect 8284 1076 8292 1084
rect 8476 1076 8484 1084
rect 8700 1076 8708 1084
rect 8716 1076 8724 1084
rect 8924 1076 8932 1084
rect 9148 1076 9156 1084
rect 9260 1076 9268 1084
rect 9468 1076 9476 1084
rect 9820 1076 9828 1084
rect 9916 1076 9924 1084
rect 3580 1056 3588 1064
rect 7244 1056 7252 1064
rect 7852 1056 7860 1064
rect 524 1036 532 1044
rect 1628 1036 1636 1044
rect 2236 1036 2244 1044
rect 2252 1036 2260 1044
rect 2732 1036 2740 1044
rect 2924 1036 2932 1044
rect 3116 1036 3124 1044
rect 5598 1036 5606 1044
rect 6764 1036 6772 1044
rect 7212 1036 7220 1044
rect 7644 1036 7652 1044
rect 7836 1036 7844 1044
rect 8348 1036 8356 1044
rect 8508 1036 8516 1044
rect 8956 1036 8964 1044
rect 9388 1036 9396 1044
rect 9596 1036 9604 1044
rect 9660 1036 9668 1044
rect 460 976 468 984
rect 684 976 692 984
rect 924 976 932 984
rect 1196 976 1204 984
rect 1404 976 1412 984
rect 1772 976 1780 984
rect 2060 976 2068 984
rect 2076 976 2084 984
rect 2252 976 2260 984
rect 3340 976 3348 984
rect 3532 976 3540 984
rect 3612 976 3620 984
rect 3772 976 3780 984
rect 4044 976 4052 984
rect 4284 976 4292 984
rect 4508 976 4516 984
rect 4732 976 4740 984
rect 4956 976 4964 984
rect 5340 976 5348 984
rect 5420 976 5428 984
rect 5580 976 5588 984
rect 6524 976 6532 984
rect 6748 976 6756 984
rect 8060 976 8068 984
rect 8076 976 8084 984
rect 8716 976 8724 984
rect 9004 976 9012 984
rect 9404 976 9412 984
rect 9420 976 9428 984
rect 2524 956 2532 964
rect 6092 956 6100 964
rect 9612 956 9620 964
rect 204 936 212 944
rect 428 936 436 944
rect 652 936 660 944
rect 892 936 900 944
rect 1116 936 1124 944
rect 1324 936 1332 944
rect 1532 936 1540 944
rect 1644 936 1652 944
rect 1868 936 1876 944
rect 2284 936 2292 944
rect 2444 936 2452 944
rect 2652 936 2660 944
rect 2764 936 2772 944
rect 2972 936 2980 944
rect 3196 936 3204 944
rect 3404 936 3412 944
rect 3740 936 3748 944
rect 3948 936 3956 944
rect 4188 936 4196 944
rect 4412 936 4420 944
rect 4460 936 4468 944
rect 4636 936 4644 944
rect 4860 936 4868 944
rect 5100 936 5108 944
rect 5212 936 5220 944
rect 5548 936 5556 944
rect 5788 936 5796 944
rect 5900 936 5908 944
rect 6124 936 6132 944
rect 6572 936 6580 944
rect 6892 936 6900 944
rect 6924 936 6932 944
rect 7132 936 7140 944
rect 7244 936 7252 944
rect 7452 936 7460 944
rect 7692 936 7700 944
rect 7916 936 7924 944
rect 8348 936 8356 944
rect 8556 936 8564 944
rect 8908 936 8916 944
rect 9132 936 9140 944
rect 9164 936 9172 944
rect 9580 936 9588 944
rect 9820 936 9828 944
rect 9900 936 9908 944
rect 1852 916 1860 924
rect 428 896 436 904
rect 684 896 692 904
rect 892 896 900 904
rect 1116 896 1124 904
rect 1340 896 1348 904
rect 1548 896 1556 904
rect 1628 896 1636 904
rect 2236 896 2244 904
rect 2476 896 2484 904
rect 2668 896 2676 904
rect 2748 896 2756 904
rect 2940 896 2948 904
rect 3180 896 3188 904
rect 3388 896 3396 904
rect 3772 896 3780 904
rect 3964 896 3972 904
rect 4188 896 4196 904
rect 4428 896 4436 904
rect 4652 896 4660 904
rect 4892 896 4900 904
rect 5100 896 5108 904
rect 5180 896 5188 904
rect 5580 896 5588 904
rect 5596 896 5604 904
rect 5788 896 5796 904
rect 5884 896 5892 904
rect 6124 896 6132 904
rect 6332 896 6340 904
rect 6540 896 6548 904
rect 6908 896 6916 904
rect 7148 896 7156 904
rect 7244 896 7252 904
rect 7452 896 7460 904
rect 8236 896 8244 904
rect 8300 896 8308 904
rect 8556 896 8564 904
rect 8908 896 8916 904
rect 9148 896 9156 904
rect 9244 896 9252 904
rect 9660 896 9668 904
rect 9820 896 9828 904
rect 9868 896 9876 904
rect 60 836 68 844
rect 2892 836 2900 844
rect 3100 836 3108 844
rect 6764 836 6772 844
rect 7388 836 7396 844
rect 8460 836 8468 844
rect 8716 836 8724 844
rect 10044 836 10052 844
rect 236 776 244 784
rect 684 776 692 784
rect 1596 776 1604 784
rect 2476 776 2484 784
rect 3596 776 3604 784
rect 4044 776 4052 784
rect 4268 776 4276 784
rect 4716 776 4724 784
rect 5340 776 5348 784
rect 5420 776 5428 784
rect 5804 776 5812 784
rect 5868 776 5876 784
rect 6284 776 6292 784
rect 60 716 68 724
rect 428 716 436 724
rect 476 716 484 724
rect 876 716 884 724
rect 956 716 964 724
rect 1340 716 1348 724
rect 1532 716 1540 724
rect 1740 716 1748 724
rect 1964 716 1972 724
rect 2044 716 2052 724
rect 2476 716 2484 724
rect 2636 716 2644 724
rect 2892 716 2900 724
rect 3084 716 3092 724
rect 3164 716 3172 724
rect 3372 716 3380 724
rect 3756 716 3764 724
rect 3820 716 3828 724
rect 4204 716 4212 724
rect 4412 716 4420 724
rect 4636 716 4644 724
rect 4732 716 4740 724
rect 4940 716 4948 724
rect 5100 716 5108 724
rect 5132 716 5140 724
rect 5580 716 5588 724
rect 6044 716 6052 724
rect 6492 716 6500 724
rect 6716 716 6724 724
rect 6796 716 6804 724
rect 7020 716 7028 724
rect 7372 716 7380 724
rect 7580 716 7588 724
rect 7660 716 7668 724
rect 8028 716 8036 724
rect 8108 716 8116 724
rect 8316 716 8324 724
rect 8684 716 8692 724
rect 8892 716 8900 724
rect 9340 716 9348 724
rect 9548 716 9556 724
rect 9644 716 9652 724
rect 9884 716 9892 724
rect 10092 716 10100 724
rect 4428 696 4436 704
rect 4476 696 4484 704
rect 4492 696 4500 704
rect 8924 696 8932 704
rect 92 676 100 684
rect 428 676 436 684
rect 540 676 548 684
rect 972 676 980 684
rect 1100 676 1108 684
rect 1308 676 1316 684
rect 1340 676 1348 684
rect 1532 676 1540 684
rect 1740 676 1748 684
rect 1948 676 1956 684
rect 2044 676 2052 684
rect 2396 676 2404 684
rect 2636 676 2644 684
rect 2860 676 2868 684
rect 2876 676 2884 684
rect 3068 676 3076 684
rect 3180 676 3188 684
rect 3388 676 3396 684
rect 3724 676 3732 684
rect 3820 676 3828 684
rect 4172 676 4180 684
rect 4396 676 4404 684
rect 4636 676 4644 684
rect 4860 676 4868 684
rect 5084 676 5092 684
rect 5212 676 5220 684
rect 5548 676 5556 684
rect 5628 676 5636 684
rect 6012 676 6020 684
rect 6124 676 6132 684
rect 6476 676 6484 684
rect 6700 676 6708 684
rect 6764 676 6772 684
rect 7036 676 7044 684
rect 7356 676 7364 684
rect 7580 676 7588 684
rect 7692 676 7700 684
rect 7820 676 7828 684
rect 8028 676 8036 684
rect 8044 676 8052 684
rect 8332 676 8340 684
rect 8460 676 8468 684
rect 8684 676 8692 684
rect 8956 676 8964 684
rect 9004 676 9012 684
rect 9324 676 9332 684
rect 9356 676 9364 684
rect 9532 676 9540 684
rect 9660 676 9668 684
rect 9884 676 9892 684
rect 10108 676 10116 684
rect 268 636 276 644
rect 716 636 724 644
rect 1164 636 1172 644
rect 1820 636 1828 644
rect 2204 636 2212 644
rect 2268 636 2276 644
rect 2716 636 2724 644
rect 3308 636 3316 644
rect 3516 636 3524 644
rect 3596 636 3604 644
rect 3964 636 3972 644
rect 6284 636 6292 644
rect 6572 636 6580 644
rect 6956 636 6964 644
rect 7180 636 7188 644
rect 7228 636 7236 644
rect 7388 636 7396 644
rect 7804 636 7812 644
rect 8252 636 8260 644
rect 8492 636 8500 644
rect 8700 636 8708 644
rect 9148 636 9156 644
rect 9196 636 9204 644
rect 9820 636 9828 644
rect 10028 636 10036 644
rect 10268 636 10276 644
rect 76 576 84 584
rect 476 576 484 584
rect 508 576 516 584
rect 956 576 964 584
rect 1356 576 1364 584
rect 1580 576 1588 584
rect 2060 576 2068 584
rect 2460 576 2468 584
rect 2700 576 2708 584
rect 2748 576 2756 584
rect 3790 576 3798 584
rect 3820 576 3828 584
rect 4252 576 4260 584
rect 4700 576 4708 584
rect 4716 576 4724 584
rect 4940 576 4948 584
rect 5468 576 5476 584
rect 5852 576 5860 584
rect 6092 576 6100 584
rect 6796 576 6804 584
rect 8092 576 8100 584
rect 8316 576 8324 584
rect 9164 576 9172 584
rect 9180 576 9188 584
rect 9852 576 9860 584
rect 10252 576 10260 584
rect 684 556 692 564
rect 1132 556 1140 564
rect 2014 556 2022 564
rect 2972 556 2980 564
rect 5452 556 5460 564
rect 9388 556 9396 564
rect 204 536 212 544
rect 316 536 324 544
rect 652 536 660 544
rect 860 536 868 544
rect 1100 536 1108 544
rect 1324 536 1332 544
rect 1564 536 1572 544
rect 1788 536 1796 544
rect 1884 536 1892 544
rect 2236 536 2244 544
rect 2332 536 2340 544
rect 2556 536 2564 544
rect 2876 536 2884 544
rect 3100 536 3108 544
rect 3180 536 3188 544
rect 3356 536 3364 544
rect 3420 536 3428 544
rect 3564 536 3572 544
rect 3676 536 3684 544
rect 4012 536 4020 544
rect 4124 536 4132 544
rect 4268 536 4276 544
rect 4444 536 4452 544
rect 4540 536 4548 544
rect 4556 536 4564 544
rect 4908 536 4916 544
rect 5132 536 5140 544
rect 5180 536 5188 544
rect 5260 536 5268 544
rect 5596 536 5604 544
rect 5676 536 5684 544
rect 5948 536 5956 544
rect 6172 536 6180 544
rect 6396 536 6404 544
rect 6620 536 6628 544
rect 6972 536 6980 544
rect 7068 536 7076 544
rect 7292 536 7300 544
rect 7500 536 7508 544
rect 7740 536 7748 544
rect 7932 536 7940 544
rect 8284 536 8292 544
rect 8476 536 8484 544
rect 8716 536 8724 544
rect 8812 536 8820 544
rect 9036 536 9044 544
rect 9372 536 9380 544
rect 9564 536 9572 544
rect 9804 536 9812 544
rect 9996 536 10004 544
rect 10108 536 10116 544
rect 3580 516 3588 524
rect 7228 516 7236 524
rect 8300 516 8308 524
rect 268 496 276 504
rect 300 496 308 504
rect 716 496 724 504
rect 892 496 900 504
rect 1132 496 1140 504
rect 1372 496 1380 504
rect 1564 496 1572 504
rect 1804 496 1812 504
rect 1868 496 1876 504
rect 2300 496 2308 504
rect 2330 496 2338 504
rect 2476 496 2484 504
rect 2892 496 2900 504
rect 3132 496 3140 504
rect 3340 496 3348 504
rect 3596 496 3604 504
rect 4092 496 4100 504
rect 4044 476 4052 484
rect 4460 496 4468 504
rect 4540 496 4548 504
rect 4940 496 4948 504
rect 5148 496 5156 504
rect 5180 496 5188 504
rect 5244 496 5252 504
rect 5612 496 5620 504
rect 5708 496 5716 504
rect 5868 496 5876 504
rect 6156 496 6164 504
rect 6972 496 6980 504
rect 7052 496 7060 504
rect 7660 496 7668 504
rect 8716 496 8724 504
rect 8780 496 8788 504
rect 8956 496 8964 504
rect 9356 496 9364 504
rect 9804 496 9812 504
rect 10028 496 10036 504
rect 10108 496 10116 504
rect 8124 476 8132 484
rect 6828 436 6836 444
rect 7196 436 7204 444
rect 7644 436 7652 444
rect 8940 436 8948 444
rect 4028 376 4036 384
rect 4460 376 4468 384
rect 5548 376 5556 384
rect 5788 376 5796 384
rect 6636 376 6644 384
rect 6284 336 6292 344
rect 220 316 228 324
rect 412 316 420 324
rect 620 316 628 324
rect 860 316 868 324
rect 1068 316 1076 324
rect 1292 316 1300 324
rect 1532 316 1540 324
rect 1836 316 1844 324
rect 2188 316 2196 324
rect 2444 316 2452 324
rect 2652 316 2660 324
rect 2860 316 2868 324
rect 3100 316 3108 324
rect 3308 316 3316 324
rect 3532 316 3540 324
rect 3772 316 3780 324
rect 3820 316 3828 324
rect 4156 316 4164 324
rect 4380 316 4388 324
rect 4396 316 4404 324
rect 4604 316 4612 324
rect 4716 316 4724 324
rect 4940 316 4948 324
rect 5388 316 5396 324
rect 5628 316 5636 324
rect 5852 316 5860 324
rect 6076 316 6084 324
rect 6236 316 6244 324
rect 6492 316 6500 324
rect 6844 316 6852 324
rect 7068 316 7076 324
rect 7292 316 7300 324
rect 7500 316 7508 324
rect 7708 316 7716 324
rect 7948 316 7956 324
rect 8172 316 8180 324
rect 8268 316 8276 324
rect 8460 316 8468 324
rect 8860 316 8868 324
rect 8924 316 8932 324
rect 9148 316 9156 324
rect 9500 316 9508 324
rect 9740 316 9748 324
rect 9820 316 9828 324
rect 10268 316 10276 324
rect 1756 296 1764 304
rect 3964 296 3972 304
rect 188 276 196 284
rect 412 276 420 284
rect 620 276 628 284
rect 892 276 900 284
rect 1068 276 1076 284
rect 1260 276 1268 284
rect 1532 276 1540 284
rect 1740 276 1748 284
rect 1836 276 1844 284
rect 2412 276 2420 284
rect 2652 276 2660 284
rect 2844 276 2852 284
rect 3084 276 3092 284
rect 3116 276 3124 284
rect 3308 276 3316 284
rect 3500 276 3508 284
rect 3532 276 3540 284
rect 3820 276 3828 284
rect 4364 276 4372 284
rect 4412 276 4420 284
rect 4604 276 4612 284
rect 4716 276 4724 284
rect 4940 276 4948 284
rect 5180 276 5188 284
rect 5388 276 5396 284
rect 5404 276 5412 284
rect 5868 276 5876 284
rect 6076 276 6084 284
rect 6284 276 6292 284
rect 6524 276 6532 284
rect 6668 276 6676 284
rect 6828 276 6836 284
rect 7036 276 7044 284
rect 7068 276 7076 284
rect 7276 276 7284 284
rect 7484 276 7492 284
rect 7516 276 7524 284
rect 7708 276 7716 284
rect 7948 276 7956 284
rect 8172 276 8180 284
rect 8268 276 8276 284
rect 8844 276 8852 284
rect 8940 276 8948 284
rect 9308 276 9316 284
rect 9500 276 9508 284
rect 9740 276 9748 284
rect 9820 276 9828 284
rect 9836 276 9844 284
rect 10012 276 10020 284
rect 10140 276 10148 284
rect 2956 256 2964 264
rect 60 236 68 244
rect 268 236 276 244
rect 492 236 500 244
rect 700 236 708 244
rect 924 236 932 244
rect 1148 236 1156 244
rect 1356 236 1364 244
rect 1548 236 1556 244
rect 1980 236 1988 244
rect 2044 236 2052 244
rect 2444 236 2452 244
rect 2716 236 2724 244
rect 3372 236 3380 244
rect 6028 236 6036 244
rect 6444 236 6452 244
rect 6908 236 6916 244
rect 7356 236 7364 244
rect 7740 236 7748 244
rect 8028 236 8036 244
rect 8636 236 8644 244
rect 8652 236 8660 244
rect 9356 236 9364 244
rect 9532 236 9540 244
rect 10028 236 10036 244
rect 748 176 756 184
rect 764 176 772 184
rect 1196 176 1204 184
rect 1628 176 1636 184
rect 1852 176 1860 184
rect 2348 176 2356 184
rect 2380 176 2388 184
rect 3708 176 3716 184
rect 4364 176 4372 184
rect 4620 176 4628 184
rect 5036 176 5044 184
rect 5468 176 5476 184
rect 5772 176 5780 184
rect 6860 176 6868 184
rect 7260 176 7268 184
rect 8348 176 8356 184
rect 8780 176 8788 184
rect 9166 176 9174 184
rect 9436 176 9444 184
rect 9596 176 9604 184
rect 9836 176 9844 184
rect 9884 176 9892 184
rect 1628 156 1636 164
rect 2540 156 2548 164
rect 2812 156 2820 164
rect 3436 156 3444 164
rect 4844 156 4852 164
rect 6636 156 6644 164
rect 92 136 100 144
rect 300 136 308 144
rect 556 136 564 144
rect 924 136 932 144
rect 1004 136 1012 144
rect 1356 136 1364 144
rect 1452 136 1460 144
rect 1820 136 1828 144
rect 2044 136 2052 144
rect 2156 136 2164 144
rect 2508 136 2516 144
rect 2732 136 2740 144
rect 2956 136 2964 144
rect 2972 136 2980 144
rect 3180 136 3188 144
rect 3420 136 3428 144
rect 3692 136 3700 144
rect 3836 136 3844 144
rect 3868 136 3876 144
rect 4092 136 4100 144
rect 4188 136 4196 144
rect 4412 136 4420 144
rect 4636 136 4644 144
rect 4876 136 4884 144
rect 5100 136 5108 144
rect 5340 136 5348 144
rect 5564 136 5572 144
rect 5788 136 5796 144
rect 6028 136 6036 144
rect 6444 136 6452 144
rect 6780 136 6788 144
rect 7052 136 7060 144
rect 7228 136 7236 144
rect 7420 136 7428 144
rect 7532 136 7540 144
rect 7692 136 7700 144
rect 7852 136 7860 144
rect 8108 136 8116 144
rect 8124 136 8132 144
rect 8348 136 8356 144
rect 8492 136 8500 144
rect 8588 136 8596 144
rect 8940 136 8948 144
rect 9036 136 9044 144
rect 9196 136 9204 144
rect 9484 136 9492 144
rect 9692 136 9700 144
rect 10012 136 10020 144
rect 60 116 68 124
rect 1900 116 1908 124
rect 7676 116 7684 124
rect 8972 116 8980 124
rect 940 96 948 104
rect 988 96 996 104
rect 1212 96 1220 104
rect 1388 96 1396 104
rect 1468 96 1476 104
rect 2076 96 2084 104
rect 2156 96 2164 104
rect 2572 96 2580 104
rect 2732 96 2740 104
rect 2972 96 2980 104
rect 3404 96 3412 104
rect 3628 96 3636 104
rect 3852 96 3860 104
rect 4076 96 4084 104
rect 4172 96 4180 104
rect 4396 96 4404 104
rect 4604 96 4612 104
rect 4860 96 4868 104
rect 5100 96 5108 104
rect 5548 96 5556 104
rect 5788 96 5796 104
rect 6026 96 6034 104
rect 6236 96 6244 104
rect 6844 96 6852 104
rect 7244 96 7252 104
rect 7516 96 7524 104
rect 8076 96 8084 104
rect 8140 96 8148 104
rect 8524 96 8532 104
rect 8588 96 8596 104
rect 8748 96 8756 104
rect 9020 96 9028 104
rect 9244 96 9252 104
rect 9466 96 9474 104
rect 9676 96 9684 104
rect 10028 96 10036 104
rect 6012 76 6020 84
rect 6652 36 6660 44
<< metal2 >>
rect 1101 7524 1107 7683
rect 1773 7604 1779 7683
rect 1821 7584 1827 7596
rect 2781 7524 2787 7683
rect 3357 7544 3363 7683
rect 3581 7624 3587 7683
rect 3389 7524 3395 7536
rect 3613 7524 3619 7616
rect 1108 7517 1116 7523
rect 317 7504 323 7516
rect 77 7464 83 7496
rect 925 7484 931 7516
rect 93 7464 99 7476
rect 909 7464 915 7476
rect 1117 7444 1123 7476
rect 1213 7464 1219 7516
rect 2061 7484 2067 7516
rect 2285 7484 2291 7516
rect 2797 7504 2803 7516
rect 1700 7477 1708 7483
rect 2029 7464 2035 7476
rect 285 7384 291 7416
rect 301 7344 307 7436
rect 669 7384 675 7396
rect 765 7344 771 7436
rect 941 7384 947 7416
rect 2525 7383 2531 7436
rect 2717 7404 2723 7476
rect 2733 7444 2739 7476
rect 3037 7464 3043 7476
rect 2516 7377 2531 7383
rect 877 7344 883 7356
rect 1085 7344 1091 7356
rect 2013 7344 2019 7356
rect 2429 7344 2435 7356
rect 644 7337 652 7343
rect 189 7324 195 7336
rect 269 7284 275 7296
rect 429 7264 435 7296
rect 877 7264 883 7296
rect 269 7124 275 7136
rect 765 7124 771 7136
rect 205 7064 211 7076
rect 61 6544 67 7036
rect 285 6963 291 7036
rect 269 6957 291 6963
rect 205 6944 211 6956
rect 269 6904 275 6957
rect 541 6944 547 6956
rect 436 6897 444 6903
rect 509 6884 515 6896
rect 77 6824 83 6836
rect 77 6724 83 6736
rect 317 6724 323 6756
rect 525 6704 531 6716
rect 93 6664 99 6676
rect 221 6636 222 6643
rect 221 6584 227 6636
rect 269 6584 275 6616
rect 301 6564 307 6676
rect 429 6557 444 6563
rect 429 6544 435 6557
rect 413 6484 419 6496
rect 445 6284 451 6296
rect 93 6264 99 6276
rect 461 6264 467 6316
rect 228 6237 236 6243
rect 77 6184 83 6196
rect 237 6184 243 6216
rect 253 6104 259 6236
rect 477 6164 483 6636
rect 669 6584 675 6596
rect 685 6564 691 7116
rect 1085 7104 1091 7296
rect 1309 7284 1315 7336
rect 1581 7284 1587 7336
rect 1629 7284 1635 7296
rect 1101 7124 1107 7136
rect 1133 7103 1139 7116
rect 1124 7097 1139 7103
rect 765 7084 771 7096
rect 1149 7084 1155 7096
rect 1117 6984 1123 7036
rect 884 6937 892 6943
rect 1181 6943 1187 7236
rect 1645 7204 1651 7336
rect 1869 7324 1875 7336
rect 1853 7304 1859 7316
rect 2013 7284 2019 7296
rect 2237 7224 2243 7236
rect 2461 7184 2467 7296
rect 2637 7124 2643 7336
rect 2733 7304 2739 7436
rect 2957 7384 2963 7456
rect 3181 7404 3187 7436
rect 3117 7384 3123 7396
rect 3229 7344 3235 7436
rect 3092 7337 3100 7343
rect 3325 7324 3331 7336
rect 2653 7284 2659 7296
rect 3101 7264 3107 7296
rect 2909 7124 2915 7236
rect 3229 7124 3235 7296
rect 3325 7264 3331 7296
rect 3517 7284 3523 7336
rect 3533 7264 3539 7296
rect 2772 7117 2780 7123
rect 1421 7104 1427 7116
rect 1220 7077 1251 7083
rect 1245 7044 1251 7077
rect 1421 7063 1427 7096
rect 1437 7084 1443 7096
rect 2237 7084 2243 7116
rect 2333 7104 2339 7116
rect 3389 7104 3395 7236
rect 3613 7164 3619 7516
rect 3709 7504 3715 7516
rect 3725 7484 3731 7683
rect 3917 7524 3923 7683
rect 4349 7524 4355 7683
rect 5165 7624 5171 7683
rect 6093 7564 6099 7576
rect 5716 7537 5852 7543
rect 4605 7524 4611 7536
rect 6189 7524 6195 7536
rect 9277 7524 9283 7536
rect 4589 7517 4604 7523
rect 3917 7484 3923 7516
rect 4132 7477 4140 7483
rect 3741 7384 3747 7476
rect 3949 7464 3955 7476
rect 4093 7364 4099 7436
rect 4269 7424 4275 7476
rect 4301 7384 4307 7516
rect 4589 7484 4595 7517
rect 6596 7517 6604 7523
rect 4605 7464 4611 7476
rect 4845 7464 4851 7476
rect 4461 7384 4467 7416
rect 5085 7404 5091 7476
rect 5133 7384 5139 7396
rect 5213 7364 5219 7436
rect 5357 7404 5363 7476
rect 5501 7424 5507 7516
rect 5853 7504 5859 7516
rect 6381 7484 6387 7516
rect 3997 7357 4012 7363
rect 3645 7344 3651 7356
rect 3997 7344 4003 7357
rect 4205 7344 4211 7356
rect 5325 7344 5331 7356
rect 4852 7337 4860 7343
rect 4445 7324 4451 7336
rect 4653 7324 4659 7336
rect 3629 7304 3635 7316
rect 4205 7304 4211 7316
rect 3981 7284 3987 7296
rect 3773 7236 3774 7243
rect 3773 7124 3779 7236
rect 4877 7144 4883 7296
rect 4957 7264 4963 7336
rect 5357 7304 5363 7396
rect 5581 7384 5587 7416
rect 5661 7384 5667 7436
rect 5837 7384 5843 7436
rect 5853 7384 5859 7476
rect 6189 7464 6195 7476
rect 6573 7424 6579 7436
rect 6029 7384 6035 7396
rect 6653 7384 6659 7476
rect 6493 7364 6499 7376
rect 5853 7304 5859 7316
rect 5901 7304 5907 7336
rect 6125 7324 6131 7336
rect 6141 7324 6147 7356
rect 6317 7304 6323 7336
rect 6356 7297 6364 7303
rect 4973 7284 4979 7296
rect 5581 7284 5587 7296
rect 5853 7284 5859 7296
rect 6589 7284 6595 7336
rect 4253 7124 4259 7136
rect 4548 7117 4556 7123
rect 4980 7117 4988 7123
rect 5220 7117 5228 7123
rect 3469 7084 3475 7096
rect 2004 7077 2035 7083
rect 1405 7057 1427 7063
rect 1181 6937 1196 6943
rect 877 6904 883 6916
rect 973 6884 979 6896
rect 1181 6884 1187 6896
rect 973 6784 979 6796
rect 1357 6724 1363 7036
rect 1405 6984 1411 7057
rect 1645 6944 1651 7056
rect 1796 7037 1804 7043
rect 1869 7024 1875 7036
rect 2029 6984 2035 7077
rect 2340 7077 2348 7083
rect 3028 7077 3036 7083
rect 2253 6984 2259 7076
rect 2285 6984 2291 6996
rect 2461 6984 2467 7076
rect 2093 6944 2099 6956
rect 1549 6864 1555 6896
rect 1613 6744 1619 6936
rect 1140 6697 1148 6703
rect 877 6524 883 6536
rect 877 6464 883 6496
rect 925 6324 931 6636
rect 1117 6584 1123 6596
rect 973 6544 979 6556
rect 1293 6484 1299 6536
rect 1309 6524 1315 6676
rect 1437 6624 1443 6716
rect 1389 6584 1395 6616
rect 1309 6504 1315 6516
rect 1325 6284 1331 6556
rect 1549 6544 1555 6636
rect 1517 6524 1523 6536
rect 1117 6264 1123 6276
rect 653 6144 659 6216
rect 221 5864 227 5916
rect 77 5744 83 5836
rect 205 5704 211 5716
rect 61 5544 67 5636
rect 221 5524 227 5536
rect 205 5484 211 5516
rect 61 5124 67 5436
rect 253 5364 259 6096
rect 445 5884 451 5956
rect 461 5884 467 5916
rect 301 5764 307 5836
rect 413 5744 419 5756
rect 413 5684 419 5696
rect 269 5524 275 5636
rect 461 5484 467 5516
rect 205 5344 211 5356
rect 301 5344 307 5436
rect 317 5344 323 5356
rect 301 5323 307 5336
rect 285 5317 307 5323
rect 285 5304 291 5317
rect 333 5303 339 5356
rect 324 5297 339 5303
rect 77 5224 83 5236
rect 461 5224 467 5236
rect 445 5124 451 5136
rect 452 5077 460 5083
rect 93 5064 99 5076
rect 205 4944 211 4956
rect 237 4804 243 5036
rect 77 4724 83 4736
rect 253 4724 259 4896
rect 445 4724 451 4736
rect 237 4564 243 4636
rect 205 4544 211 4556
rect 205 4284 211 4336
rect 221 4284 227 4316
rect 93 4203 99 4276
rect 77 4197 99 4203
rect 77 4184 83 4197
rect 237 4164 243 4236
rect 205 4144 211 4156
rect 237 4064 243 4096
rect 77 3984 83 4016
rect 237 3884 243 3916
rect 212 3877 220 3883
rect 253 3844 259 4496
rect 285 4344 291 4636
rect 477 4504 483 6136
rect 525 6084 531 6096
rect 653 6084 659 6096
rect 669 5884 675 5896
rect 701 5803 707 5916
rect 717 5904 723 6236
rect 877 6144 883 6156
rect 1085 6144 1091 6196
rect 1325 6184 1331 6196
rect 1293 6144 1299 6156
rect 1085 6104 1091 6116
rect 1309 6104 1315 6116
rect 877 6084 883 6096
rect 1309 6084 1315 6096
rect 765 5924 771 5936
rect 781 5884 787 5896
rect 685 5797 707 5803
rect 685 5784 691 5797
rect 877 5784 883 5876
rect 493 5704 499 5716
rect 493 5124 499 5696
rect 509 5264 515 5736
rect 701 5724 707 5776
rect 733 5724 739 5736
rect 925 5624 931 5836
rect 973 5784 979 5836
rect 1101 5744 1107 6076
rect 1117 5924 1123 5936
rect 1373 5924 1379 6516
rect 1533 6504 1539 6516
rect 1421 6324 1427 6336
rect 1533 6324 1539 6496
rect 1597 6324 1603 6636
rect 1613 6504 1619 6736
rect 1629 6724 1635 6896
rect 2077 6884 2083 6896
rect 2413 6864 2419 6936
rect 2733 6924 2739 7056
rect 3101 6984 3107 7076
rect 2733 6904 2739 6916
rect 2749 6904 2755 6936
rect 2973 6924 2979 6936
rect 2948 6917 2956 6923
rect 1853 6724 1859 6756
rect 2685 6744 2691 6896
rect 1901 6724 1907 6736
rect 2269 6704 2275 6716
rect 1933 6684 1939 6696
rect 2365 6684 2371 6716
rect 2381 6684 2387 6736
rect 2717 6724 2723 6736
rect 2749 6704 2755 6896
rect 2957 6884 2963 6896
rect 2941 6724 2947 6756
rect 2948 6677 2956 6683
rect 1652 6637 1660 6643
rect 1757 6584 1763 6636
rect 1933 6584 1939 6676
rect 2045 6637 2060 6643
rect 2045 6544 2051 6637
rect 2285 6584 2291 6676
rect 2701 6664 2707 6676
rect 2404 6537 2412 6543
rect 1629 6504 1635 6536
rect 2429 6504 2435 6656
rect 2493 6584 2499 6616
rect 2509 6564 2515 6636
rect 2717 6584 2723 6596
rect 2797 6544 2803 6636
rect 2845 6544 2851 6556
rect 1437 6264 1443 6276
rect 1613 6244 1619 6496
rect 1629 6324 1635 6496
rect 2637 6464 2643 6496
rect 2861 6484 2867 6496
rect 2237 6424 2243 6436
rect 3117 6364 3123 6496
rect 3149 6404 3155 7036
rect 3181 7023 3187 7076
rect 3693 7064 3699 7076
rect 4013 7064 4019 7076
rect 3165 7017 3187 7023
rect 3165 6984 3171 7017
rect 3341 6984 3347 6996
rect 3309 6884 3315 6896
rect 3533 6864 3539 6936
rect 3165 6844 3171 6856
rect 3165 6823 3171 6836
rect 3165 6817 3187 6823
rect 3181 6544 3187 6817
rect 3245 6724 3251 6736
rect 3597 6724 3603 7036
rect 3885 7024 3891 7036
rect 3757 6904 3763 6936
rect 3789 6904 3795 6956
rect 3981 6944 3987 7036
rect 4029 6904 4035 7116
rect 4477 7084 4483 7116
rect 4541 7084 4547 7096
rect 4100 7057 4108 7063
rect 4237 6944 4243 7076
rect 4317 6944 4323 7076
rect 4461 7064 4467 7076
rect 4413 6944 4419 6976
rect 4100 6937 4227 6943
rect 4077 6904 4083 6916
rect 3773 6864 3779 6896
rect 4221 6884 4227 6937
rect 4196 6837 4204 6843
rect 4045 6724 4051 6736
rect 4237 6724 4243 6936
rect 4269 6824 4275 6836
rect 4269 6724 4275 6756
rect 4413 6744 4419 6896
rect 4461 6823 4467 7056
rect 4541 6944 4547 7076
rect 4557 6964 4563 7116
rect 4989 7084 4995 7096
rect 5236 7077 5244 7083
rect 4605 6944 4611 6956
rect 4621 6904 4627 6916
rect 4461 6817 4483 6823
rect 3245 6544 3251 6716
rect 4061 6684 4067 6696
rect 4477 6684 4483 6817
rect 4685 6724 4691 7036
rect 4989 6944 4995 7076
rect 5373 7064 5379 7236
rect 5796 7117 5811 7123
rect 5805 7084 5811 7117
rect 5197 6924 5203 6936
rect 4877 6884 4883 6896
rect 4701 6824 4707 6836
rect 4941 6824 4947 6836
rect 5037 6724 5043 6756
rect 5085 6724 5091 6896
rect 5597 6824 5603 7036
rect 5645 6944 5651 7036
rect 5789 7004 5795 7076
rect 6125 7064 6131 7076
rect 5901 6944 5907 7036
rect 6013 6984 6019 6996
rect 6269 6924 6275 7236
rect 6573 7124 6579 7136
rect 6285 6944 6291 7036
rect 6461 6984 6467 7076
rect 6477 6984 6483 7116
rect 6589 7084 6595 7096
rect 6781 7064 6787 7436
rect 6797 7364 6803 7516
rect 7037 7344 7043 7436
rect 7069 7404 7075 7516
rect 7101 7464 7107 7476
rect 7245 7384 7251 7436
rect 7309 7363 7315 7436
rect 7469 7424 7475 7516
rect 7549 7504 7555 7516
rect 7533 7384 7539 7476
rect 7309 7357 7363 7363
rect 7357 7344 7363 7357
rect 7709 7344 7715 7436
rect 7789 7384 7795 7476
rect 7981 7404 7987 7516
rect 8205 7504 8211 7516
rect 8413 7504 8419 7516
rect 8452 7477 8460 7483
rect 8740 7477 8748 7483
rect 8205 7464 8211 7476
rect 8765 7444 8771 7516
rect 9485 7504 9491 7516
rect 9709 7504 9715 7516
rect 9917 7504 9923 7516
rect 9940 7477 9948 7483
rect 9293 7464 9299 7476
rect 9501 7464 9507 7476
rect 9709 7464 9715 7476
rect 7821 7397 7859 7403
rect 7821 7384 7827 7397
rect 7853 7384 7859 7397
rect 8141 7384 8147 7436
rect 8301 7384 8307 7396
rect 7780 7337 7788 7343
rect 7469 7324 7475 7336
rect 7837 7304 7843 7376
rect 8349 7364 8355 7436
rect 8045 7344 8051 7356
rect 8269 7344 8275 7356
rect 8493 7324 8499 7336
rect 8573 7324 8579 7436
rect 8733 7384 8739 7396
rect 8589 7304 8595 7316
rect 8052 7297 8060 7303
rect 6957 7064 6963 7076
rect 6797 7024 6803 7036
rect 6925 6984 6931 6996
rect 6781 6944 6787 6956
rect 6212 6897 6220 6903
rect 6301 6864 6307 6936
rect 6957 6904 6963 7056
rect 6317 6884 6323 6896
rect 6685 6884 6691 6896
rect 5773 6764 5779 6836
rect 5853 6743 5859 6836
rect 6365 6784 6371 6856
rect 6733 6744 6739 6896
rect 6973 6744 6979 7236
rect 7021 7184 7027 7296
rect 7373 7264 7379 7296
rect 7469 7284 7475 7296
rect 8269 7264 8275 7296
rect 7181 7224 7187 7236
rect 7389 7124 7395 7136
rect 7613 7124 7619 7236
rect 7165 7084 7171 7096
rect 7389 6984 7395 7076
rect 7469 6964 7475 7076
rect 7677 6964 7683 7236
rect 8173 7124 8179 7156
rect 7949 7104 7955 7116
rect 8397 7104 8403 7116
rect 8173 7084 8179 7096
rect 8413 7084 8419 7156
rect 7869 7064 7875 7076
rect 7581 6957 7596 6963
rect 7469 6944 7475 6956
rect 7581 6944 7587 6957
rect 7236 6937 7244 6943
rect 7005 6924 7011 6936
rect 7773 6904 7779 6936
rect 6989 6884 6995 6896
rect 6989 6844 6995 6876
rect 7853 6803 7859 7036
rect 7965 6964 7971 7076
rect 8333 6944 8339 7036
rect 8557 6984 8563 7036
rect 8589 6944 8595 7296
rect 8605 7104 8611 7336
rect 8829 7264 8835 7336
rect 8637 7124 8643 7136
rect 8973 7124 8979 7236
rect 8989 7124 8995 7436
rect 9037 7424 9043 7436
rect 9261 7344 9267 7376
rect 9053 7324 9059 7336
rect 9421 7224 9427 7236
rect 9437 7224 9443 7436
rect 9581 7344 9587 7356
rect 8868 7117 8876 7123
rect 9437 7104 9443 7116
rect 8637 7084 8643 7096
rect 8884 7077 8892 7083
rect 8685 6957 8700 6963
rect 8685 6944 8691 6957
rect 8797 6944 8803 7036
rect 8861 6924 8867 6936
rect 8893 6904 8899 6936
rect 8669 6864 8675 6896
rect 7853 6797 7875 6803
rect 5853 6737 5875 6743
rect 5261 6724 5267 6736
rect 4756 6717 4764 6723
rect 4052 6677 4060 6683
rect 4484 6677 4492 6683
rect 3629 6584 3635 6636
rect 4349 6624 4355 6636
rect 4045 6584 4051 6596
rect 4253 6584 4259 6596
rect 4509 6544 4515 6716
rect 4589 6704 4595 6716
rect 4589 6664 4595 6676
rect 4829 6544 4835 6556
rect 4180 6537 4195 6543
rect 3181 6504 3187 6516
rect 3549 6324 3555 6436
rect 3236 6317 3244 6323
rect 2237 6284 2243 6296
rect 1661 6264 1667 6276
rect 1885 6264 1891 6276
rect 2013 6236 2014 6243
rect 1549 6184 1555 6196
rect 1997 6184 2003 6216
rect 1748 6137 1756 6143
rect 1773 6104 1779 6136
rect 1117 5784 1123 5876
rect 989 5524 995 5536
rect 916 5517 931 5523
rect 685 5504 691 5516
rect 669 5484 675 5496
rect 925 5484 931 5517
rect 909 5464 915 5476
rect 989 5384 995 5496
rect 1005 5484 1011 5696
rect 1069 5544 1075 5736
rect 1197 5724 1203 5736
rect 1373 5724 1379 5916
rect 1405 5784 1411 6096
rect 1533 6064 1539 6096
rect 1588 5917 1603 5923
rect 1597 5864 1603 5917
rect 1629 5884 1635 6096
rect 1965 6084 1971 6136
rect 2013 6024 2019 6236
rect 2253 6204 2259 6316
rect 2461 6284 2467 6296
rect 2477 6264 2483 6316
rect 2333 6224 2339 6236
rect 2445 6184 2451 6196
rect 2205 6144 2211 6156
rect 2493 6144 2499 6316
rect 2765 6284 2771 6316
rect 2797 6284 2803 6296
rect 2701 6264 2707 6276
rect 2685 6184 2691 6196
rect 2717 6184 2723 6196
rect 1805 5904 1811 5916
rect 2029 5884 2035 5896
rect 2061 5884 2067 5916
rect 1805 5864 1811 5876
rect 1885 5744 1891 5756
rect 1085 5704 1091 5716
rect 1901 5704 1907 5836
rect 1117 5664 1123 5696
rect 1421 5664 1427 5696
rect 1645 5664 1651 5696
rect 1885 5684 1891 5696
rect 1373 5484 1379 5516
rect 1005 5464 1011 5476
rect 1149 5424 1155 5436
rect 669 5324 675 5336
rect 1149 5324 1155 5356
rect 1357 5344 1363 5356
rect 1581 5304 1587 5316
rect 909 5284 915 5296
rect 1229 5244 1235 5276
rect 1229 5224 1235 5236
rect 669 5124 675 5136
rect 893 5124 899 5156
rect 1565 5124 1571 5256
rect 1581 5184 1587 5276
rect 964 5117 972 5123
rect 989 5084 995 5096
rect 1220 5077 1228 5083
rect 893 5064 899 5076
rect 509 4904 515 5036
rect 909 4944 915 4956
rect 1117 4944 1123 4956
rect 669 4904 675 4936
rect 941 4724 947 4896
rect 1133 4884 1139 5036
rect 1341 4984 1347 5076
rect 1517 4964 1523 5036
rect 1517 4944 1523 4956
rect 1565 4944 1571 4956
rect 1197 4904 1203 4916
rect 1373 4724 1379 4936
rect 1597 4924 1603 5476
rect 1789 5424 1795 5636
rect 1805 5524 1811 5676
rect 2029 5484 2035 5496
rect 2077 5484 2083 6096
rect 2205 6084 2211 6096
rect 2205 6064 2211 6076
rect 2317 6064 2323 6136
rect 2493 6084 2499 6136
rect 2861 6104 2867 6236
rect 3101 6157 3116 6163
rect 3101 6143 3107 6157
rect 3389 6144 3395 6236
rect 3565 6144 3571 6276
rect 3581 6184 3587 6536
rect 3965 6524 3971 6536
rect 3773 6324 3779 6496
rect 3965 6464 3971 6496
rect 4189 6344 4195 6537
rect 3821 6324 3827 6336
rect 4045 6324 4051 6336
rect 4317 6324 4323 6336
rect 3092 6137 3107 6143
rect 3549 6104 3555 6136
rect 3316 6097 3324 6103
rect 2509 5924 2515 5936
rect 2269 5904 2275 5916
rect 2509 5904 2515 5916
rect 2285 5864 2291 5876
rect 2493 5864 2499 5876
rect 2525 5864 2531 6096
rect 2724 5917 2732 5923
rect 2701 5884 2707 5896
rect 2909 5884 2915 5956
rect 2925 5924 2931 6056
rect 2285 5844 2291 5856
rect 2333 5824 2339 5836
rect 2269 5784 2275 5796
rect 2349 5744 2355 5756
rect 2525 5744 2531 5856
rect 2116 5697 2124 5703
rect 2340 5697 2348 5703
rect 2493 5484 2499 5496
rect 2525 5484 2531 5516
rect 1613 5384 1619 5396
rect 1805 5344 1811 5356
rect 1853 5304 1859 5376
rect 2029 5344 2035 5356
rect 1645 5124 1651 5296
rect 1677 5064 1683 5076
rect 1821 4964 1827 5036
rect 1837 4984 1843 5116
rect 2045 4984 2051 5116
rect 1901 4944 1907 4956
rect 1677 4924 1683 4936
rect 2061 4924 2067 5296
rect 2013 4736 2014 4743
rect 916 4717 924 4723
rect 685 4663 691 4716
rect 909 4664 915 4676
rect 1149 4664 1155 4716
rect 685 4657 707 4663
rect 685 4584 691 4596
rect 308 4497 316 4503
rect 461 4184 467 4276
rect 429 3904 435 3916
rect 205 3664 211 3736
rect 237 3704 243 3816
rect 253 3784 259 3796
rect 285 3764 291 3836
rect 445 3744 451 3756
rect 461 3704 467 3736
rect 61 3584 67 3656
rect 61 3384 67 3496
rect 221 3464 227 3516
rect 445 3464 451 3476
rect 301 3384 307 3416
rect 205 3324 211 3336
rect 61 2964 67 3036
rect 189 3004 195 3076
rect 93 2944 99 2956
rect 301 2944 307 3076
rect 77 2924 83 2936
rect 237 2684 243 2716
rect 461 2684 467 2716
rect 205 2664 211 2676
rect 61 2504 67 2636
rect 237 2584 243 2656
rect 253 2584 259 2616
rect 205 2324 211 2476
rect 61 2124 67 2236
rect 237 2184 243 2336
rect 461 2184 467 2396
rect 301 2104 307 2156
rect 205 1904 211 1916
rect 61 1764 67 1836
rect 221 1784 227 2016
rect 301 1864 307 1876
rect 429 1824 435 1836
rect 253 1784 259 1816
rect 221 1777 222 1784
rect 93 1744 99 1756
rect 445 1744 451 1756
rect 77 1724 83 1736
rect 445 1664 451 1696
rect 205 1484 211 1556
rect 429 1524 435 1536
rect 429 1464 435 1476
rect 61 1344 67 1436
rect 100 1297 108 1303
rect 77 1184 83 1196
rect 237 1124 243 1236
rect 221 1104 227 1116
rect 461 984 467 1076
rect 477 1004 483 4496
rect 493 4324 499 4456
rect 685 4384 691 4496
rect 669 4184 675 4256
rect 525 4084 531 4096
rect 541 4063 547 4136
rect 525 4057 547 4063
rect 525 3984 531 4057
rect 653 3864 659 3876
rect 669 3864 675 3916
rect 701 3784 707 4657
rect 909 4544 915 4556
rect 1181 4524 1187 4636
rect 1341 4584 1347 4676
rect 1373 4604 1379 4716
rect 1549 4684 1555 4736
rect 1789 4724 1795 4736
rect 1885 4724 1891 4736
rect 2013 4724 2019 4736
rect 1789 4664 1795 4676
rect 1901 4664 1907 4676
rect 1917 4604 1923 4676
rect 1405 4584 1411 4596
rect 1837 4584 1843 4596
rect 1613 4544 1619 4556
rect 1604 4537 1612 4543
rect 1700 4537 1708 4543
rect 1245 4524 1251 4536
rect 2077 4524 2083 5476
rect 2221 5344 2227 5436
rect 2301 5324 2307 5436
rect 2349 5304 2355 5436
rect 2532 5377 2540 5383
rect 2269 5284 2275 5296
rect 2349 5264 2355 5296
rect 2125 5124 2131 5136
rect 2557 5103 2563 5696
rect 2573 5664 2579 5836
rect 2781 5804 2787 5836
rect 2909 5744 2915 5756
rect 2941 5704 2947 5956
rect 2989 5944 2995 6096
rect 3101 6084 3107 6096
rect 3565 6084 3571 6096
rect 3581 6024 3587 6176
rect 3597 6124 3603 6316
rect 4477 6284 4483 6536
rect 3805 6264 3811 6276
rect 4045 6264 4051 6276
rect 4477 6264 4483 6276
rect 3613 5964 3619 6236
rect 3757 6144 3763 6156
rect 2989 5924 2995 5936
rect 3597 5924 3603 5936
rect 2573 5644 2579 5656
rect 2749 5524 2755 5536
rect 2749 5424 2755 5476
rect 2740 5337 2748 5343
rect 2733 5284 2739 5296
rect 2717 5124 2723 5156
rect 2541 5097 2563 5103
rect 2125 5084 2131 5096
rect 2477 5064 2483 5076
rect 2109 4824 2115 4836
rect 2093 4584 2099 4676
rect 2269 4624 2275 4636
rect 2285 4624 2291 5036
rect 2317 4904 2323 5036
rect 2477 4924 2483 4936
rect 2509 4624 2515 4896
rect 2525 4724 2531 4896
rect 2525 4644 2531 4656
rect 2301 4584 2307 4596
rect 2253 4537 2268 4543
rect 1245 4484 1251 4496
rect 1165 4384 1171 4396
rect 909 4324 915 4336
rect 1437 4324 1443 4516
rect 1597 4464 1603 4496
rect 1693 4464 1699 4496
rect 2253 4464 2259 4537
rect 2285 4504 2291 4576
rect 2461 4544 2467 4576
rect 900 4277 908 4283
rect 772 4237 780 4243
rect 925 4184 931 4216
rect 941 4164 947 4316
rect 1437 4304 1443 4316
rect 1453 4284 1459 4436
rect 2045 4324 2051 4436
rect 2461 4324 2467 4476
rect 2260 4317 2268 4323
rect 1805 4284 1811 4316
rect 2260 4277 2268 4283
rect 2333 4277 2348 4283
rect 1197 4164 1203 4236
rect 1581 4224 1587 4236
rect 1821 4224 1827 4276
rect 2013 4264 2019 4276
rect 1613 4184 1619 4196
rect 1229 4144 1235 4156
rect 1597 4144 1603 4176
rect 1805 4144 1811 4156
rect 2020 4137 2028 4143
rect 765 4104 771 4116
rect 2077 4104 2083 4236
rect 2333 4184 2339 4277
rect 2525 4224 2531 4496
rect 2493 4184 2499 4216
rect 2461 4144 2467 4156
rect 1220 4097 1228 4103
rect 2237 4084 2243 4096
rect 2477 4064 2483 4096
rect 2541 4084 2547 5097
rect 2669 4984 2675 5076
rect 2589 4924 2595 4936
rect 2781 4724 2787 5676
rect 2957 5484 2963 5736
rect 2836 5337 2844 5343
rect 2829 5304 2835 5316
rect 2948 5117 2956 5123
rect 2948 5077 2956 5083
rect 2941 4984 2947 4996
rect 2797 4944 2803 4956
rect 2989 4944 2995 5916
rect 3805 5904 3811 5916
rect 3357 5884 3363 5896
rect 3021 5864 3027 5876
rect 3149 5804 3155 5836
rect 3181 5784 3187 5876
rect 3021 5744 3027 5756
rect 3005 5664 3011 5696
rect 3165 5524 3171 5536
rect 3149 5464 3155 5476
rect 3005 5384 3011 5396
rect 3021 5304 3027 5436
rect 3181 5324 3187 5336
rect 3197 5284 3203 5296
rect 3213 5203 3219 5836
rect 3437 5804 3443 5836
rect 3373 5724 3379 5736
rect 3389 5704 3395 5776
rect 3581 5744 3587 5756
rect 3645 5724 3651 5836
rect 3661 5784 3667 5796
rect 3789 5724 3795 5736
rect 3645 5664 3651 5716
rect 3229 5584 3235 5636
rect 3389 5524 3395 5556
rect 3469 5524 3475 5536
rect 3485 5484 3491 5656
rect 3837 5624 3843 6236
rect 4125 6224 4131 6236
rect 3997 6124 4003 6136
rect 4013 6104 4019 6176
rect 4221 6144 4227 6176
rect 4493 6084 4499 6316
rect 4509 6304 4515 6536
rect 4941 6503 4947 6636
rect 5181 6624 5187 6636
rect 5101 6557 5116 6563
rect 5101 6544 5107 6557
rect 5284 6537 5292 6543
rect 5325 6504 5331 6636
rect 5405 6604 5411 6736
rect 5844 6717 5859 6723
rect 5629 6684 5635 6716
rect 5821 6684 5827 6696
rect 5853 6684 5859 6717
rect 5869 6704 5875 6737
rect 6173 6724 6179 6736
rect 7501 6724 7507 6736
rect 7300 6717 7308 6723
rect 6068 6677 6076 6683
rect 5405 6584 5411 6596
rect 5421 6544 5427 6636
rect 5533 6544 5539 6676
rect 5613 6664 5619 6676
rect 5565 6544 5571 6656
rect 5629 6584 5635 6596
rect 5693 6564 5699 6636
rect 5789 6544 5795 6636
rect 5533 6504 5539 6536
rect 5565 6504 5571 6536
rect 4941 6497 4963 6503
rect 4509 6104 4515 6296
rect 4525 6184 4531 6356
rect 4637 6344 4643 6436
rect 4909 6324 4915 6356
rect 4909 6317 4910 6324
rect 4685 6304 4691 6316
rect 4909 6264 4915 6276
rect 4941 6264 4947 6436
rect 4957 6284 4963 6497
rect 5764 6497 5772 6503
rect 5085 6484 5091 6496
rect 5533 6344 5539 6496
rect 4573 6144 4579 6156
rect 4548 6097 4556 6103
rect 4253 5924 4259 6076
rect 4029 5884 4035 5896
rect 3885 5724 3891 5836
rect 4045 5784 4051 5916
rect 4253 5904 4259 5916
rect 4244 5877 4252 5883
rect 4093 5837 4108 5843
rect 3885 5684 3891 5696
rect 3901 5644 3907 5736
rect 4093 5644 4099 5837
rect 4228 5737 4236 5743
rect 3805 5484 3811 5596
rect 3917 5524 3923 5556
rect 3821 5484 3827 5516
rect 3917 5484 3923 5496
rect 4253 5484 4259 5696
rect 4269 5524 4275 6076
rect 4484 5917 4499 5923
rect 4493 5884 4499 5917
rect 4733 5884 4739 6236
rect 4973 6204 4979 6316
rect 4909 6184 4915 6196
rect 4989 6144 4995 6336
rect 5373 6324 5379 6336
rect 5453 6304 5459 6316
rect 5485 6284 5491 6296
rect 5373 6264 5379 6276
rect 5805 6264 5811 6276
rect 5597 6236 5598 6243
rect 5373 6184 5379 6196
rect 5597 6144 5603 6236
rect 5661 6144 5667 6156
rect 4788 6137 4796 6143
rect 5229 6104 5235 6136
rect 4756 6097 4764 6103
rect 5005 6064 5011 6096
rect 5245 6064 5251 6136
rect 5677 6124 5683 6236
rect 5805 6184 5811 6236
rect 5405 6044 5411 6096
rect 5581 6084 5587 6096
rect 5629 6044 5635 6056
rect 5261 5984 5267 5996
rect 5266 5977 5267 5984
rect 5037 5924 5043 5936
rect 5405 5924 5411 6036
rect 5629 5984 5635 6036
rect 5629 5977 5630 5984
rect 4701 5864 4707 5876
rect 4493 5784 4499 5816
rect 4717 5784 4723 5796
rect 4909 5764 4915 5876
rect 4989 5784 4995 5916
rect 5380 5877 5388 5883
rect 5181 5744 5187 5836
rect 5389 5784 5395 5856
rect 4349 5684 4355 5696
rect 4333 5664 4339 5676
rect 4333 5584 4339 5656
rect 4365 5524 4371 5736
rect 4573 5724 4579 5736
rect 5165 5704 5171 5716
rect 4781 5684 4787 5696
rect 4925 5624 4931 5636
rect 4493 5524 4499 5556
rect 4269 5504 4275 5516
rect 4509 5484 4515 5516
rect 4589 5484 4595 5496
rect 4829 5484 4835 5556
rect 5405 5544 5411 5636
rect 5181 5524 5187 5536
rect 5421 5524 5427 5936
rect 5501 5864 5507 5876
rect 5661 5784 5667 6096
rect 5837 6084 5843 6656
rect 6093 6624 6099 6716
rect 6333 6684 6339 6696
rect 6173 6664 6179 6676
rect 6621 6664 6627 6676
rect 6269 6544 6275 6556
rect 5885 6524 5891 6536
rect 5869 6504 5875 6516
rect 6013 6344 6019 6436
rect 5917 6244 5923 6276
rect 6077 6264 6083 6496
rect 6093 6484 6099 6496
rect 6253 6344 6259 6436
rect 6285 6384 6291 6656
rect 6829 6644 6835 6676
rect 6765 6604 6771 6636
rect 6477 6584 6483 6596
rect 6925 6557 6940 6563
rect 6925 6544 6931 6557
rect 7021 6544 7027 6636
rect 7037 6604 7043 6716
rect 7069 6644 7075 6676
rect 7293 6664 7299 6676
rect 7181 6584 7187 6596
rect 6573 6524 6579 6536
rect 6909 6504 6915 6536
rect 7165 6504 7171 6576
rect 7165 6484 7171 6496
rect 6365 6324 6371 6356
rect 6589 6324 6595 6336
rect 6125 6304 6131 6316
rect 6141 6264 6147 6276
rect 6365 6264 6371 6276
rect 5997 6144 6003 6156
rect 6045 5964 6051 6236
rect 6253 6104 6259 6256
rect 6333 6144 6339 6156
rect 6244 6097 6252 6103
rect 5725 5924 5731 5936
rect 5725 5884 5731 5896
rect 6077 5884 6083 5896
rect 6157 5864 6163 6096
rect 6333 6064 6339 6096
rect 6477 5944 6483 6036
rect 6525 6024 6531 6236
rect 6749 6184 6755 6336
rect 6765 6284 6771 6436
rect 6813 6324 6819 6336
rect 7213 6284 7219 6636
rect 7357 6544 7363 6556
rect 7437 6504 7443 6636
rect 7517 6604 7523 6676
rect 7725 6664 7731 6676
rect 7668 6657 7676 6663
rect 7837 6584 7843 6596
rect 7853 6564 7859 6636
rect 7796 6537 7804 6543
rect 7869 6504 7875 6797
rect 7933 6684 7939 6716
rect 8269 6684 8275 6816
rect 8477 6723 8483 6836
rect 8477 6717 8492 6723
rect 8580 6717 8588 6723
rect 8285 6684 8291 6716
rect 8909 6684 8915 6716
rect 7917 6664 7923 6676
rect 8461 6664 8467 6676
rect 8786 6636 8787 6643
rect 8061 6584 8067 6616
rect 8093 6544 8099 6636
rect 8733 6544 8739 6636
rect 8781 6604 8787 6636
rect 8925 6584 8931 6716
rect 8228 6537 8243 6543
rect 7364 6497 7372 6503
rect 7597 6484 7603 6496
rect 7869 6484 7875 6496
rect 7277 6284 7283 6296
rect 7012 6277 7020 6283
rect 7181 6184 7187 6236
rect 6925 6144 6931 6156
rect 7245 6144 7251 6216
rect 7341 6144 7347 6236
rect 7453 6224 7459 6436
rect 7501 6284 7507 6436
rect 8029 6324 8035 6536
rect 8045 6504 8051 6536
rect 8237 6523 8243 6537
rect 8269 6523 8275 6536
rect 8237 6517 8275 6523
rect 8356 6497 8364 6503
rect 8253 6484 8259 6496
rect 8253 6324 8259 6336
rect 7629 6144 7635 6236
rect 6557 6104 6563 6136
rect 6573 6124 6579 6136
rect 7645 6124 7651 6236
rect 7853 6224 7859 6316
rect 8020 6277 8028 6283
rect 8061 6264 8067 6316
rect 8436 6277 8444 6283
rect 7677 6144 7683 6176
rect 7885 6144 7891 6236
rect 8013 6144 8019 6236
rect 8253 6184 8259 6276
rect 8461 6184 8467 6496
rect 8477 6324 8483 6356
rect 8557 6244 8563 6316
rect 8573 6284 8579 6356
rect 8109 6144 8115 6156
rect 8333 6124 8339 6136
rect 7149 6104 7155 6116
rect 7581 6104 7587 6116
rect 7677 6104 7683 6116
rect 8541 6104 8547 6236
rect 8685 6184 8691 6276
rect 7220 6097 7228 6103
rect 7682 6097 7683 6104
rect 6925 6084 6931 6096
rect 8013 6084 8019 6096
rect 8109 6064 8115 6096
rect 6781 6044 6787 6056
rect 6797 5924 6803 6036
rect 7821 5944 7827 6036
rect 7853 5944 7859 6036
rect 8333 5984 8339 6096
rect 7949 5924 7955 5936
rect 6541 5884 6547 5896
rect 6756 5877 6764 5883
rect 5693 5744 5699 5756
rect 5469 5724 5475 5736
rect 5693 5664 5699 5696
rect 5709 5517 5724 5523
rect 5181 5484 5187 5496
rect 5389 5484 5395 5496
rect 5709 5484 5715 5517
rect 3405 5424 3411 5476
rect 3485 5464 3491 5476
rect 3805 5464 3811 5476
rect 4132 5437 4147 5443
rect 3613 5424 3619 5436
rect 4061 5384 4067 5436
rect 3636 5337 3644 5343
rect 3421 5324 3427 5336
rect 3869 5324 3875 5336
rect 3949 5304 3955 5316
rect 3412 5297 3420 5303
rect 3268 5237 3276 5243
rect 3197 5197 3219 5203
rect 3149 5084 3155 5096
rect 3181 4983 3187 5156
rect 3172 4977 3187 4983
rect 2797 4884 2803 4896
rect 3037 4744 3043 4936
rect 3197 4724 3203 5197
rect 3213 5124 3219 5136
rect 2708 4717 2716 4723
rect 2797 4704 2803 4716
rect 2820 4677 2828 4683
rect 2701 4664 2707 4676
rect 2717 4544 2723 4676
rect 3149 4664 3155 4676
rect 2957 4544 2963 4636
rect 3149 4544 3155 4556
rect 2765 4484 2771 4496
rect 2797 4484 2803 4496
rect 3165 4464 3171 4496
rect 3181 4384 3187 4656
rect 3197 4584 3203 4596
rect 2797 4324 2803 4336
rect 2701 4304 2707 4316
rect 3149 4284 3155 4296
rect 2701 4264 2707 4276
rect 3165 4264 3171 4316
rect 2717 4184 2723 4196
rect 2701 4144 2707 4156
rect 3133 4144 3139 4156
rect 3149 4104 3155 4116
rect 3149 4097 3150 4104
rect 2701 4084 2707 4096
rect 1197 3924 1203 3936
rect 1773 3924 1779 3956
rect 2237 3924 2243 3936
rect 2653 3923 2659 4076
rect 2733 3924 2739 3936
rect 2653 3917 2675 3923
rect 733 3744 739 3836
rect 909 3823 915 3916
rect 1421 3904 1427 3916
rect 1869 3904 1875 3916
rect 2461 3884 2467 3896
rect 1773 3864 1779 3876
rect 2477 3864 2483 3916
rect 2669 3884 2675 3917
rect 2916 3917 2924 3923
rect 2957 3884 2963 4096
rect 3197 3924 3203 4376
rect 2013 3836 2014 3843
rect 909 3817 931 3823
rect 925 3784 931 3817
rect 1629 3744 1635 3836
rect 1805 3757 1836 3763
rect 1805 3744 1811 3757
rect 509 3437 524 3443
rect 509 3344 515 3437
rect 541 3384 547 3456
rect 701 3184 707 3696
rect 893 3504 899 3516
rect 941 3464 947 3736
rect 957 3504 963 3696
rect 1117 3684 1123 3696
rect 1133 3664 1139 3736
rect 1853 3704 1859 3776
rect 2013 3764 2019 3836
rect 2093 3824 2099 3836
rect 2045 3784 2051 3796
rect 2477 3724 2483 3736
rect 2029 3704 2035 3716
rect 2253 3664 2259 3696
rect 1117 3484 1123 3556
rect 1341 3524 1347 3536
rect 1341 3517 1342 3524
rect 1197 3504 1203 3516
rect 1133 3464 1139 3496
rect 1341 3484 1347 3496
rect 973 3344 979 3436
rect 1181 3384 1187 3456
rect 1437 3384 1443 3476
rect 1453 3464 1459 3516
rect 1805 3464 1811 3476
rect 1837 3384 1843 3576
rect 2484 3517 2492 3523
rect 2029 3504 2035 3516
rect 2269 3484 2275 3516
rect 2013 3464 2019 3476
rect 2013 3384 2019 3456
rect 1245 3344 1251 3356
rect 1588 3337 1596 3343
rect 909 3304 915 3336
rect 941 3164 947 3336
rect 1709 3324 1715 3336
rect 1933 3324 1939 3336
rect 1005 3304 1011 3316
rect 1245 3264 1251 3296
rect 1597 3284 1603 3296
rect 509 3124 515 3136
rect 877 3124 883 3136
rect 1092 3117 1100 3123
rect 509 3083 515 3116
rect 500 3077 515 3083
rect 525 3064 531 3076
rect 509 2984 515 2996
rect 637 2944 643 2956
rect 941 2944 947 3036
rect 1165 2984 1171 3256
rect 1533 3124 1539 3136
rect 1533 3104 1539 3116
rect 1197 3064 1203 3076
rect 1325 2984 1331 2996
rect 1549 2984 1555 3076
rect 653 2884 659 2896
rect 701 2724 707 2836
rect 669 2664 675 2676
rect 701 2584 707 2596
rect 749 2544 755 2936
rect 1101 2823 1107 2836
rect 1085 2817 1107 2823
rect 909 2684 915 2716
rect 941 2584 947 2756
rect 1085 2724 1091 2817
rect 1181 2724 1187 2796
rect 1293 2764 1299 2936
rect 1309 2904 1315 2916
rect 1549 2864 1555 2936
rect 1597 2904 1603 3196
rect 1613 3004 1619 3116
rect 2093 3084 2099 3476
rect 2269 3404 2275 3436
rect 2285 3384 2291 3476
rect 2125 3344 2131 3376
rect 2141 3344 2147 3356
rect 2381 3344 2387 3356
rect 2125 3304 2131 3336
rect 2386 3296 2387 3303
rect 2381 3284 2387 3296
rect 1860 3077 1868 3083
rect 1645 3064 1651 3076
rect 2093 3064 2099 3076
rect 1789 2984 1795 2996
rect 2237 2984 2243 3276
rect 2525 3224 2531 3836
rect 2541 3704 2547 3796
rect 2669 3744 2675 3876
rect 2909 3864 2915 3876
rect 2957 3864 2963 3876
rect 2749 3784 2755 3816
rect 2957 3757 2972 3763
rect 2957 3743 2963 3757
rect 2948 3737 2963 3743
rect 2589 3724 2595 3736
rect 2557 3584 2563 3596
rect 3021 3584 3027 3876
rect 3133 3864 3139 3876
rect 3172 3737 3180 3743
rect 2708 3517 2723 3523
rect 2717 3484 2723 3517
rect 2692 3477 2700 3483
rect 2573 3384 2579 3416
rect 2957 3384 2963 3516
rect 3156 3477 3164 3483
rect 3181 3424 3187 3516
rect 2733 3304 2739 3376
rect 2781 3323 2787 3356
rect 2797 3344 2803 3356
rect 2813 3323 2819 3336
rect 2781 3317 2819 3323
rect 3165 3304 3171 3336
rect 2813 3284 2819 3296
rect 3213 3284 3219 5116
rect 3245 5084 3251 5116
rect 3261 5064 3267 5076
rect 3421 4984 3427 5196
rect 3565 5123 3571 5176
rect 3565 5117 3612 5123
rect 3604 5077 3612 5083
rect 3469 5024 3475 5036
rect 3645 4984 3651 5196
rect 3693 5124 3699 5236
rect 4125 5184 4131 5196
rect 3933 5124 3939 5156
rect 3725 5064 3731 5076
rect 3853 5036 3854 5043
rect 3853 5024 3859 5036
rect 3261 4944 3267 4956
rect 3261 4904 3267 4916
rect 3485 4904 3491 4956
rect 3501 4864 3507 4936
rect 3837 4864 3843 4936
rect 3869 4904 3875 5016
rect 4077 4944 4083 4956
rect 4141 4884 4147 5437
rect 4221 5344 4227 5356
rect 4253 5344 4259 5476
rect 5709 5464 5715 5476
rect 4749 5344 4755 5436
rect 4973 5343 4979 5436
rect 4973 5337 4988 5343
rect 4205 5304 4211 5336
rect 4797 5324 4803 5336
rect 4861 5324 4867 5336
rect 5012 5297 5020 5303
rect 4797 5284 4803 5296
rect 4301 5084 4307 5096
rect 4397 5084 4403 5096
rect 4413 5064 4419 5076
rect 4365 4984 4371 4996
rect 4164 4897 4172 4903
rect 4493 4864 4499 4936
rect 4525 4904 4531 4956
rect 3229 4784 3235 4856
rect 4141 4784 4147 4836
rect 3597 4724 3603 4736
rect 3405 4684 3411 4716
rect 3597 4704 3603 4716
rect 3581 4664 3587 4676
rect 3469 4584 3475 4636
rect 3613 4524 3619 4536
rect 3677 4524 3683 4636
rect 3805 4564 3811 4676
rect 3837 4524 3843 4536
rect 3869 4524 3875 4636
rect 3613 4324 3619 4336
rect 3581 4264 3587 4276
rect 3229 4184 3235 4236
rect 3405 4144 3411 4256
rect 3421 4184 3427 4196
rect 3645 4184 3651 4516
rect 3860 4497 3868 4503
rect 3661 4364 3667 4436
rect 3885 4384 3891 4636
rect 4061 4584 4067 4716
rect 4285 4663 4291 4716
rect 4477 4664 4483 4676
rect 4285 4657 4307 4663
rect 4301 4624 4307 4657
rect 4269 4544 4275 4576
rect 4013 4324 4019 4336
rect 3805 4304 3811 4316
rect 3789 4244 3795 4276
rect 3661 4224 3667 4236
rect 3821 4144 3827 4316
rect 4061 4284 4067 4496
rect 3997 4264 4003 4276
rect 4077 4264 4083 4536
rect 4269 4504 4275 4516
rect 4525 4504 4531 4876
rect 4557 4744 4563 5036
rect 4749 4984 4755 5116
rect 4765 4984 4771 5076
rect 4829 4984 4835 5036
rect 4989 4984 4995 5116
rect 4605 4944 4611 4956
rect 4948 4937 4956 4943
rect 4605 4884 4611 4896
rect 4573 4743 4579 4856
rect 5037 4744 5043 5436
rect 5101 5384 5107 5396
rect 5229 5324 5235 5336
rect 5245 5284 5251 5296
rect 5197 5124 5203 5136
rect 5277 5124 5283 5456
rect 5501 5384 5507 5396
rect 5357 5344 5363 5376
rect 5581 5344 5587 5436
rect 5837 5344 5843 5476
rect 5869 5343 5875 5436
rect 5885 5384 5891 5836
rect 5933 5824 5939 5836
rect 6157 5744 6163 5836
rect 6493 5744 6499 5756
rect 6493 5724 6499 5736
rect 5917 5704 5923 5716
rect 6061 5544 6067 5636
rect 5869 5337 5900 5343
rect 5693 5264 5699 5336
rect 5197 5064 5203 5076
rect 5181 4904 5187 4916
rect 5266 4836 5267 4843
rect 5261 4824 5267 4836
rect 4573 4737 4595 4743
rect 4237 4324 4243 4496
rect 4237 4304 4243 4316
rect 4541 4284 4547 4716
rect 4589 4684 4595 4737
rect 4941 4724 4947 4736
rect 5261 4724 5267 4736
rect 5165 4664 5171 4716
rect 5277 4684 5283 4696
rect 4701 4637 4716 4643
rect 4573 4584 4579 4616
rect 4317 4244 4323 4276
rect 4701 4244 4707 4637
rect 5181 4584 5187 4676
rect 5245 4584 5251 4596
rect 5250 4577 5251 4584
rect 4829 4544 4835 4556
rect 5348 4537 5356 4543
rect 4733 4523 4739 4536
rect 4733 4517 4755 4523
rect 4749 4504 4755 4517
rect 4717 4324 4723 4496
rect 4925 4324 4931 4336
rect 5309 4324 5315 4496
rect 5373 4484 5379 4496
rect 5389 4324 5395 4356
rect 5437 4324 5443 5036
rect 5453 4944 5459 5116
rect 5629 5084 5635 5156
rect 5725 5124 5731 5236
rect 5933 5164 5939 5436
rect 6077 5404 6083 5516
rect 6285 5484 6291 5636
rect 6125 5364 6131 5436
rect 6301 5384 6307 5516
rect 6333 5464 6339 5476
rect 6349 5424 6355 5636
rect 6365 5524 6371 5536
rect 6525 5343 6531 5436
rect 6573 5384 6579 5836
rect 6861 5824 6867 5916
rect 7021 5904 7027 5916
rect 7085 5864 7091 5876
rect 6973 5784 6979 5816
rect 7021 5744 7027 5836
rect 7517 5824 7523 5916
rect 8157 5884 8163 5896
rect 7421 5784 7427 5816
rect 7693 5784 7699 5856
rect 7741 5824 7747 5876
rect 7933 5784 7939 5816
rect 7188 5777 7196 5783
rect 7741 5744 7747 5756
rect 8148 5737 8156 5743
rect 7021 5704 7027 5736
rect 7277 5724 7283 5736
rect 7492 5697 7500 5703
rect 6589 5684 6595 5696
rect 6749 5524 6755 5636
rect 6813 5524 6819 5536
rect 7005 5484 7011 5696
rect 7725 5664 7731 5696
rect 8093 5684 8099 5696
rect 7021 5524 7027 5536
rect 7405 5524 7411 5556
rect 7501 5524 7507 5536
rect 7709 5524 7715 5556
rect 7933 5504 7939 5516
rect 7053 5484 7059 5496
rect 7725 5484 7731 5496
rect 7949 5484 7955 5496
rect 6740 5477 6748 5483
rect 6621 5404 6627 5476
rect 6717 5464 6723 5476
rect 6621 5384 6627 5396
rect 6845 5384 6851 5476
rect 7197 5424 7203 5436
rect 6717 5344 6723 5356
rect 6493 5337 6531 5343
rect 6477 5324 6483 5336
rect 6141 5304 6147 5316
rect 6381 5304 6387 5316
rect 5949 5124 5955 5216
rect 6285 5124 6291 5276
rect 6493 5263 6499 5337
rect 6717 5324 6723 5336
rect 6701 5304 6707 5316
rect 7149 5304 7155 5376
rect 7325 5364 7331 5476
rect 7389 5464 7395 5476
rect 7853 5424 7859 5436
rect 8141 5404 8147 5696
rect 8301 5524 8307 5836
rect 8333 5584 8339 5956
rect 8701 5924 8707 6236
rect 8733 5924 8739 6436
rect 8941 6324 8947 7076
rect 9069 6984 9075 7036
rect 9469 7024 9475 7236
rect 9629 7124 9635 7436
rect 9693 7264 9699 7296
rect 9629 7064 9635 7076
rect 9133 6984 9139 7016
rect 9453 6944 9459 6956
rect 9517 6944 9523 7036
rect 9645 7004 9651 7116
rect 9853 7104 9859 7236
rect 9869 7144 9875 7436
rect 9917 7324 9923 7336
rect 9924 7297 9932 7303
rect 9684 7037 9692 7043
rect 10061 6984 10067 7076
rect 9885 6944 9891 6956
rect 9373 6904 9379 6936
rect 9117 6884 9123 6896
rect 9341 6884 9347 6896
rect 9437 6884 9443 6896
rect 9661 6884 9667 6896
rect 10061 6784 10067 6896
rect 10077 6784 10083 7116
rect 10237 6984 10243 6996
rect 10109 6924 10115 6936
rect 9565 6724 9571 6736
rect 9005 6704 9011 6716
rect 9901 6704 9907 6716
rect 10244 6677 10259 6683
rect 9021 6664 9027 6676
rect 9188 6537 9196 6543
rect 9133 6504 9139 6516
rect 9149 6384 9155 6476
rect 8989 6324 8995 6376
rect 9149 6344 9155 6376
rect 8909 6304 8915 6316
rect 8909 6264 8915 6276
rect 8765 6184 8771 6236
rect 9165 6184 9171 6216
rect 8770 6177 8771 6184
rect 9213 6144 9219 6636
rect 9565 6624 9571 6676
rect 9677 6664 9683 6676
rect 9805 6584 9811 6616
rect 9565 6544 9571 6556
rect 9677 6524 9683 6536
rect 8996 6137 9004 6143
rect 8893 6124 8899 6136
rect 9341 6084 9347 6096
rect 8989 5924 8995 5996
rect 9389 5984 9395 6436
rect 9421 6364 9427 6436
rect 9437 6324 9443 6436
rect 9645 6384 9651 6496
rect 9789 6324 9795 6356
rect 9533 6144 9539 6156
rect 9037 5924 9043 5936
rect 9261 5924 9267 5976
rect 9421 5924 9427 6036
rect 9581 5924 9587 6096
rect 9597 5924 9603 6236
rect 9789 6224 9795 6276
rect 9821 6264 9827 6456
rect 9645 6184 9651 6196
rect 9837 6144 9843 6556
rect 10013 6524 10019 6536
rect 10013 6484 10019 6496
rect 9869 6364 9875 6436
rect 10061 6324 10067 6636
rect 10253 6584 10259 6677
rect 10125 6544 10131 6556
rect 10221 6284 10227 6296
rect 10013 6184 10019 6276
rect 10077 6244 10083 6276
rect 10029 6184 10035 6196
rect 10077 6144 10083 6236
rect 9805 6064 9811 6096
rect 8509 5864 8515 5876
rect 8349 5524 8355 5836
rect 8365 5784 8371 5796
rect 8493 5744 8499 5796
rect 8573 5784 8579 5916
rect 8605 5864 8611 5876
rect 8493 5544 8499 5736
rect 8509 5684 8515 5696
rect 8701 5564 8707 5736
rect 8781 5704 8787 5836
rect 8813 5744 8819 5776
rect 8781 5684 8787 5696
rect 8957 5624 8963 5636
rect 8733 5524 8739 5536
rect 8957 5504 8963 5516
rect 8605 5477 8716 5483
rect 8173 5464 8179 5476
rect 8413 5424 8419 5476
rect 8605 5464 8611 5477
rect 8061 5384 8067 5396
rect 8461 5384 8467 5396
rect 7181 5344 7187 5356
rect 7517 5344 7523 5356
rect 8420 5337 8428 5343
rect 8525 5343 8531 5436
rect 8557 5344 8563 5436
rect 8893 5384 8899 5396
rect 8941 5384 8947 5396
rect 8733 5344 8739 5356
rect 8509 5337 8531 5343
rect 7629 5324 7635 5336
rect 7869 5324 7875 5336
rect 7069 5264 7075 5296
rect 7149 5284 7155 5296
rect 7629 5284 7635 5296
rect 6493 5257 6531 5263
rect 6333 5184 6339 5256
rect 6525 5224 6531 5257
rect 6557 5124 6563 5136
rect 6909 5124 6915 5236
rect 7213 5124 7219 5176
rect 7309 5124 7315 5236
rect 7709 5184 7715 5216
rect 8189 5184 8195 5336
rect 8205 5284 8211 5296
rect 8429 5264 8435 5296
rect 7869 5124 7875 5136
rect 7965 5124 7971 5156
rect 8196 5117 8204 5123
rect 8509 5123 8515 5337
rect 8749 5304 8755 5376
rect 8989 5344 8995 5916
rect 9261 5884 9267 5896
rect 9005 5664 9011 5696
rect 9021 5404 9027 5876
rect 9165 5784 9171 5856
rect 9037 5584 9043 5736
rect 9373 5724 9379 5736
rect 9421 5624 9427 5836
rect 9581 5804 9587 5876
rect 9693 5864 9699 5876
rect 9716 5737 9724 5743
rect 9853 5724 9859 6136
rect 9885 6124 9891 6136
rect 10221 6096 10222 6103
rect 9869 6064 9875 6096
rect 9885 6084 9891 6096
rect 10045 5824 10051 5836
rect 10045 5784 10051 5796
rect 9901 5724 9907 5736
rect 9885 5704 9891 5716
rect 9460 5697 9468 5703
rect 10221 5684 10227 6096
rect 9837 5524 9843 5536
rect 9037 5344 9043 5436
rect 9197 5424 9203 5516
rect 9396 5477 9404 5483
rect 9325 5384 9331 5396
rect 9325 5377 9326 5384
rect 9197 5344 9203 5356
rect 9421 5344 9427 5516
rect 10029 5484 10035 5496
rect 9469 5364 9475 5436
rect 9821 5384 9827 5476
rect 9645 5364 9651 5376
rect 10045 5364 10051 5396
rect 10061 5384 10067 5516
rect 9869 5344 9875 5356
rect 10029 5344 10035 5356
rect 8525 5204 8531 5236
rect 8541 5124 8547 5256
rect 9069 5204 9075 5336
rect 9085 5304 9091 5336
rect 9549 5324 9555 5336
rect 9181 5284 9187 5296
rect 9773 5284 9779 5296
rect 8509 5117 8531 5123
rect 5661 5004 5667 5116
rect 5869 5104 5875 5116
rect 6653 5104 6659 5116
rect 5853 5063 5859 5096
rect 5885 5084 5891 5096
rect 5901 5063 5907 5076
rect 6541 5064 6547 5076
rect 7005 5064 7011 5076
rect 7213 5064 7219 5076
rect 5853 5057 5907 5063
rect 5597 4944 5603 4976
rect 5597 4904 5603 4936
rect 5629 4904 5635 4976
rect 5725 4964 5731 5036
rect 5837 4984 5843 4996
rect 6109 4964 6115 5036
rect 6397 4984 6403 5036
rect 7069 5024 7075 5036
rect 6541 4984 6547 4996
rect 5693 4944 5699 4956
rect 5693 4884 5699 4896
rect 5917 4784 5923 4936
rect 6141 4784 6147 4936
rect 6685 4924 6691 4936
rect 6781 4904 6787 4976
rect 6797 4944 6803 5016
rect 7133 4984 7139 5036
rect 7293 4944 7299 5036
rect 7357 4984 7363 5056
rect 7357 4977 7358 4984
rect 6509 4884 6515 4896
rect 6989 4884 6995 4896
rect 6509 4844 6515 4876
rect 5492 4717 5500 4723
rect 5693 4717 5708 4723
rect 5613 4464 5619 4496
rect 5453 4364 5459 4436
rect 5645 4344 5651 4636
rect 5693 4584 5699 4717
rect 5933 4684 5939 4716
rect 6301 4684 6307 4716
rect 6509 4684 6515 4736
rect 6589 4724 6595 4736
rect 6948 4717 6956 4723
rect 6973 4684 6979 4716
rect 5956 4677 5964 4683
rect 5725 4664 5731 4676
rect 6285 4624 6291 4676
rect 6317 4584 6323 4616
rect 5949 4544 5955 4556
rect 6157 4544 6163 4556
rect 6157 4524 6163 4536
rect 6477 4524 6483 4536
rect 5917 4504 5923 4516
rect 5837 4464 5843 4496
rect 6141 4484 6147 4496
rect 6493 4484 6499 4496
rect 6749 4484 6755 4636
rect 6749 4343 6755 4436
rect 6797 4364 6803 4636
rect 6973 4584 6979 4676
rect 7005 4584 7011 4936
rect 7405 4884 7411 5076
rect 7501 5044 7507 5076
rect 7517 5004 7523 5116
rect 7981 5084 7987 5096
rect 8525 5084 8531 5117
rect 9037 5104 9043 5116
rect 7869 5064 7875 5076
rect 7437 4924 7443 4936
rect 7444 4897 7452 4903
rect 7261 4724 7267 4736
rect 7373 4724 7379 4836
rect 7597 4724 7603 5036
rect 7613 4984 7619 4996
rect 7741 4944 7747 5036
rect 7885 4944 7891 4956
rect 8125 4944 8131 5036
rect 8205 4984 8211 5076
rect 8749 5064 8755 5076
rect 7780 4937 7788 4943
rect 7869 4924 7875 4936
rect 8221 4904 8227 4976
rect 8349 4964 8355 5036
rect 8397 4944 8403 5036
rect 8429 4944 8435 5056
rect 8461 4984 8467 5056
rect 8589 4964 8595 5036
rect 8765 4944 8771 4976
rect 9037 4944 9043 5096
rect 9053 5084 9059 5156
rect 9405 5123 9411 5236
rect 9693 5124 9699 5136
rect 10045 5124 10051 5356
rect 9396 5117 9411 5123
rect 9476 5117 9484 5123
rect 9149 4984 9155 5076
rect 9501 5064 9507 5076
rect 9197 4944 9203 5036
rect 9245 4964 9251 5036
rect 9901 4944 9907 5036
rect 10173 4984 10179 4996
rect 9572 4937 9580 4943
rect 9604 4937 9612 4943
rect 8301 4904 8307 4916
rect 7652 4897 7772 4903
rect 7844 4737 7852 4743
rect 7037 4684 7043 4696
rect 7693 4684 7699 4696
rect 7389 4636 7390 4643
rect 7165 4544 7171 4636
rect 7389 4604 7395 4636
rect 7277 4544 7283 4596
rect 7453 4544 7459 4636
rect 7581 4604 7587 4676
rect 7709 4544 7715 4636
rect 8029 4544 8035 4836
rect 8317 4784 8323 4936
rect 8564 4717 8572 4723
rect 8045 4604 8051 4716
rect 8477 4684 8483 4716
rect 8493 4704 8499 4716
rect 8253 4664 8259 4676
rect 8589 4664 8595 4676
rect 8573 4564 8579 4596
rect 8717 4584 8723 4636
rect 8733 4584 8739 4756
rect 8749 4644 8755 4896
rect 8781 4724 8787 4876
rect 8973 4784 8979 4936
rect 9181 4904 9187 4916
rect 10020 4897 10028 4903
rect 9613 4884 9619 4896
rect 9149 4724 9155 4736
rect 9341 4724 9347 4836
rect 9581 4724 9587 4736
rect 9693 4724 9699 4756
rect 10093 4724 10099 4736
rect 8797 4684 8803 4696
rect 9229 4684 9235 4716
rect 9693 4704 9699 4716
rect 9684 4677 9692 4683
rect 9213 4664 9219 4676
rect 9917 4664 9923 4676
rect 10253 4644 10259 4676
rect 8445 4544 8451 4556
rect 8573 4544 8579 4556
rect 8893 4544 8899 4636
rect 6829 4524 6835 4536
rect 7156 4497 7164 4503
rect 6829 4464 6835 4496
rect 6749 4337 6803 4343
rect 6157 4324 6163 4336
rect 6621 4324 6627 4336
rect 5092 4317 5100 4323
rect 5604 4317 5612 4323
rect 6797 4323 6803 4337
rect 7037 4324 7043 4356
rect 6797 4317 6828 4323
rect 4861 4284 4867 4296
rect 5069 4284 5075 4296
rect 5170 4236 5171 4243
rect 3604 4097 3612 4103
rect 3389 4064 3395 4096
rect 3453 4044 3459 4096
rect 3453 3984 3459 4036
rect 3373 3924 3379 3936
rect 3229 3704 3235 3836
rect 3261 3784 3267 3876
rect 3645 3824 3651 3836
rect 3661 3744 3667 4116
rect 3837 4084 3843 4096
rect 3821 3884 3827 3896
rect 3853 3784 3859 3916
rect 3869 3904 3875 4236
rect 4061 4104 4067 4136
rect 3949 3784 3955 3876
rect 3853 3777 3854 3784
rect 3709 3744 3715 3756
rect 4045 3744 4051 3756
rect 3412 3737 3420 3743
rect 3405 3704 3411 3716
rect 3693 3684 3699 3696
rect 3725 3624 3731 3696
rect 4029 3524 4035 3696
rect 3597 3504 3603 3516
rect 3805 3484 3811 3516
rect 3837 3484 3843 3516
rect 3581 3464 3587 3476
rect 3620 3457 3628 3463
rect 4013 3444 4019 3476
rect 3458 3436 3459 3443
rect 3453 3404 3459 3436
rect 3405 3264 3411 3296
rect 2493 3124 2499 3156
rect 3085 3124 3091 3136
rect 3453 3124 3459 3396
rect 3597 3344 3603 3436
rect 3837 3344 3843 3356
rect 4077 3344 4083 3696
rect 4093 3484 4099 4236
rect 4317 4184 4323 4236
rect 4477 4144 4483 4236
rect 4541 4144 4547 4236
rect 4669 4144 4675 4236
rect 4749 4157 4764 4163
rect 4749 4144 4755 4157
rect 4109 3524 4115 3736
rect 4125 3584 4131 4136
rect 4173 4064 4179 4136
rect 4525 4104 4531 4116
rect 4333 3924 4339 4056
rect 4381 3924 4387 3936
rect 4605 3904 4611 3916
rect 4621 3884 4627 3896
rect 4141 3784 4147 3836
rect 4157 3764 4163 3836
rect 4365 3784 4371 3796
rect 4285 3744 4291 3756
rect 4493 3724 4499 3736
rect 4509 3504 4515 3516
rect 4541 3504 4547 3836
rect 4557 3784 4563 3856
rect 4765 3764 4771 3836
rect 4733 3744 4739 3756
rect 4749 3684 4755 3696
rect 4125 3464 4131 3476
rect 4244 3437 4252 3443
rect 4285 3384 4291 3436
rect 4077 3324 4083 3336
rect 3613 3284 3619 3296
rect 4061 3284 4067 3296
rect 3613 3184 3619 3256
rect 2477 3104 2483 3116
rect 2861 3104 2867 3116
rect 2413 3084 2419 3096
rect 2461 2984 2467 3016
rect 2093 2944 2099 2956
rect 1757 2924 1763 2936
rect 1229 2724 1235 2736
rect 1140 2677 1148 2683
rect 1357 2644 1363 2656
rect 1133 2584 1139 2596
rect 1005 2544 1011 2556
rect 564 2537 572 2543
rect 493 2344 499 2496
rect 701 2484 707 2496
rect 653 2324 659 2336
rect 877 2304 883 2316
rect 493 2264 499 2276
rect 653 2144 659 2156
rect 669 2104 675 2116
rect 509 1984 515 2016
rect 653 1884 659 1916
rect 637 1864 643 1876
rect 653 1744 659 1756
rect 669 1704 675 1716
rect 532 1517 540 1523
rect 653 1403 659 1476
rect 669 1424 675 1436
rect 653 1397 675 1403
rect 669 1384 675 1397
rect 653 1144 659 1296
rect 653 1084 659 1136
rect 685 1124 691 2256
rect 708 2177 716 2183
rect 893 2104 899 2496
rect 989 2484 995 2496
rect 1005 2324 1011 2536
rect 1101 2264 1107 2276
rect 1133 2264 1139 2436
rect 1309 2284 1315 2336
rect 1309 2264 1315 2276
rect 957 2184 963 2236
rect 957 2144 963 2156
rect 1293 2144 1299 2256
rect 957 2064 963 2096
rect 861 1924 867 1936
rect 957 1924 963 1956
rect 717 1764 723 1836
rect 765 1744 771 1876
rect 861 1864 867 1876
rect 1309 1864 1315 1876
rect 1341 1844 1347 1916
rect 1117 1784 1123 1796
rect 1181 1744 1187 1836
rect 1341 1784 1347 1796
rect 925 1504 931 1696
rect 1213 1684 1219 1696
rect 941 1564 947 1656
rect 1117 1584 1123 1656
rect 973 1524 979 1556
rect 733 1344 739 1356
rect 877 1344 883 1436
rect 925 1344 931 1496
rect 1149 1484 1155 1496
rect 980 1477 988 1483
rect 1117 1384 1123 1416
rect 1357 1403 1363 2616
rect 1421 2584 1427 2676
rect 1597 2584 1603 2876
rect 1837 2784 1843 2876
rect 1997 2864 2003 2896
rect 1853 2784 1859 2796
rect 2029 2724 2035 2916
rect 2317 2904 2323 2916
rect 2333 2864 2339 2936
rect 2237 2824 2243 2836
rect 2253 2724 2259 2756
rect 1661 2704 1667 2716
rect 2253 2684 2259 2696
rect 1693 2664 1699 2676
rect 1661 2584 1667 2616
rect 1666 2577 1667 2584
rect 1421 2544 1427 2576
rect 1796 2537 1804 2543
rect 1828 2537 1836 2543
rect 2020 2537 2028 2543
rect 1812 2497 1820 2503
rect 1597 2324 1603 2336
rect 2013 2324 2019 2396
rect 1773 2304 1779 2316
rect 1757 2284 1763 2296
rect 1981 2284 1987 2316
rect 1389 2164 1395 2236
rect 1645 2164 1651 2256
rect 1805 2184 1811 2196
rect 1773 2144 1779 2156
rect 1837 2124 1843 2236
rect 1549 2084 1555 2096
rect 1389 1924 1395 2036
rect 1796 1917 1804 1923
rect 1757 1897 1795 1903
rect 1421 1864 1427 1876
rect 1757 1864 1763 1897
rect 1789 1884 1795 1897
rect 1773 1864 1779 1876
rect 1629 1784 1635 1816
rect 1645 1784 1651 1796
rect 1437 1744 1443 1756
rect 1789 1724 1795 1736
rect 1821 1724 1827 1856
rect 1405 1584 1411 1696
rect 1629 1524 1635 1596
rect 1613 1484 1619 1496
rect 1357 1397 1379 1403
rect 1373 1384 1379 1397
rect 1213 1344 1219 1356
rect 1581 1344 1587 1396
rect 1677 1344 1683 1356
rect 877 1324 883 1336
rect 1197 1304 1203 1336
rect 893 1184 899 1236
rect 909 1124 915 1136
rect 941 1124 947 1276
rect 973 1264 979 1296
rect 1661 1264 1667 1296
rect 1357 1124 1363 1236
rect 1117 1104 1123 1116
rect 1197 1084 1203 1096
rect 1357 1084 1363 1096
rect 765 1064 771 1076
rect 685 984 691 996
rect 205 944 211 956
rect 653 944 659 956
rect 893 924 899 936
rect 61 724 67 836
rect 237 784 243 796
rect 429 724 435 736
rect 436 677 444 683
rect 93 664 99 676
rect 77 584 83 596
rect 205 544 211 556
rect 269 504 275 636
rect 477 584 483 716
rect 509 584 515 916
rect 909 903 915 1036
rect 900 897 915 903
rect 685 784 691 896
rect 957 744 963 1076
rect 1117 924 1123 936
rect 1341 884 1347 896
rect 884 717 892 723
rect 957 664 963 716
rect 973 684 979 696
rect 1341 684 1347 716
rect 653 544 659 556
rect 317 524 323 536
rect 717 504 723 636
rect 957 584 963 616
rect 861 544 867 556
rect 1101 544 1107 556
rect 1149 543 1155 596
rect 1133 537 1155 543
rect 893 504 899 536
rect 1133 504 1139 537
rect 221 324 227 396
rect 621 324 627 496
rect 1165 484 1171 636
rect 1357 584 1363 596
rect 1325 544 1331 556
rect 1373 504 1379 1176
rect 1565 1144 1571 1156
rect 1821 1084 1827 1716
rect 1853 1624 1859 2236
rect 1997 2104 2003 2136
rect 2045 2104 2051 2496
rect 2077 2404 2083 2636
rect 2093 2584 2099 2656
rect 2093 2504 2099 2576
rect 2228 2537 2236 2543
rect 2244 2497 2259 2503
rect 2205 2324 2211 2336
rect 2180 2277 2188 2283
rect 2093 2184 2099 2276
rect 2253 2124 2259 2497
rect 2285 2384 2291 2856
rect 2324 2777 2332 2783
rect 2317 2764 2323 2776
rect 2477 2724 2483 3096
rect 2845 3084 2851 3096
rect 3309 3084 3315 3116
rect 3748 3077 3756 3083
rect 2717 3044 2723 3076
rect 2717 3003 2723 3036
rect 2701 2997 2723 3003
rect 2541 2984 2547 2996
rect 2701 2904 2707 2997
rect 2925 2984 2931 2996
rect 2941 2824 2947 3036
rect 3165 2984 3171 3016
rect 3117 2944 3123 2956
rect 2701 2724 2707 2756
rect 2477 2704 2483 2716
rect 2893 2684 2899 2816
rect 2916 2717 2924 2723
rect 2749 2664 2755 2676
rect 2893 2664 2899 2676
rect 3101 2664 3107 2676
rect 2356 2537 2364 2543
rect 2749 2504 2755 2636
rect 2941 2584 2947 2656
rect 3133 2624 3139 2656
rect 3149 2604 3155 2716
rect 3181 2603 3187 3036
rect 3325 3024 3331 3076
rect 3373 2984 3379 2996
rect 3789 2944 3795 3256
rect 4205 3124 4211 3136
rect 4301 3123 4307 3496
rect 4573 3484 4579 3556
rect 4781 3524 4787 4236
rect 4925 4144 4931 4236
rect 5165 4184 5171 4236
rect 5213 4184 5219 4276
rect 5277 4264 5283 4276
rect 4948 4137 4956 4143
rect 4973 4104 4979 4116
rect 5053 4104 5059 4156
rect 5309 4144 5315 4316
rect 5917 4264 5923 4276
rect 5389 4124 5395 4136
rect 5629 4124 5635 4136
rect 5661 4104 5667 4236
rect 5757 4224 5763 4236
rect 5933 4184 5939 4316
rect 6381 4284 6387 4296
rect 7053 4284 7059 4456
rect 7213 4324 7219 4536
rect 7901 4524 7907 4536
rect 8125 4524 8131 4536
rect 8477 4504 8483 4516
rect 8909 4504 8915 4536
rect 8541 4497 8556 4503
rect 7469 4484 7475 4496
rect 7837 4364 7843 4436
rect 7901 4364 7907 4496
rect 7460 4317 7468 4323
rect 7325 4304 7331 4316
rect 7549 4304 7555 4316
rect 7469 4284 7475 4296
rect 6605 4264 6611 4276
rect 6349 4184 6355 4196
rect 5748 4137 5756 4143
rect 5965 4104 5971 4156
rect 5981 4144 5987 4156
rect 5741 4084 5747 4096
rect 5965 4084 5971 4096
rect 5485 4004 5491 4036
rect 5069 3924 5075 3936
rect 5069 3884 5075 3896
rect 4836 3877 4844 3883
rect 5261 3863 5267 3916
rect 5293 3884 5299 3996
rect 5501 3864 5507 3916
rect 5517 3884 5523 3936
rect 5869 3924 5875 3936
rect 6093 3924 6099 3936
rect 6061 3864 6067 3876
rect 6157 3864 6163 4176
rect 6205 4144 6211 4156
rect 6461 4144 6467 4236
rect 6669 4224 6675 4236
rect 6413 4104 6419 4136
rect 6429 4064 6435 4136
rect 6589 3984 6595 4196
rect 6781 4184 6787 4256
rect 6813 4244 6819 4276
rect 7117 4164 7123 4236
rect 7197 4184 7203 4196
rect 7069 4144 7075 4156
rect 7245 4144 7251 4276
rect 7565 4224 7571 4276
rect 7389 4144 7395 4156
rect 7485 4144 7491 4156
rect 6637 3944 6643 4096
rect 6173 3924 6179 3936
rect 6388 3917 6396 3923
rect 6733 3884 6739 4096
rect 6861 3984 6867 4136
rect 6973 3984 6979 4056
rect 6749 3924 6755 3976
rect 7261 3924 7267 4036
rect 6829 3904 6835 3916
rect 7165 3884 7171 3896
rect 5261 3857 5283 3863
rect 4957 3744 4963 3756
rect 4989 3724 4995 3836
rect 5277 3784 5283 3857
rect 5197 3744 5203 3756
rect 5421 3744 5427 3756
rect 5949 3743 5955 3836
rect 6413 3784 6419 3876
rect 6589 3764 6595 3836
rect 6637 3744 6643 3856
rect 6829 3784 6835 3796
rect 7012 3777 7020 3783
rect 5949 3737 5964 3743
rect 6180 3737 6188 3743
rect 5197 3704 5203 3716
rect 5421 3704 5427 3716
rect 4989 3584 4995 3696
rect 5533 3684 5539 3696
rect 5757 3664 5763 3736
rect 6973 3724 6979 3736
rect 6173 3704 6179 3716
rect 6989 3703 6995 3776
rect 7101 3744 7107 3836
rect 7181 3784 7187 3916
rect 7373 3884 7379 4096
rect 7405 4064 7411 4096
rect 7485 4084 7491 4096
rect 7469 3924 7475 4076
rect 7389 3904 7395 3916
rect 7485 3884 7491 3916
rect 6980 3697 6995 3703
rect 5757 3644 5763 3656
rect 4797 3484 4803 3496
rect 4468 3477 4476 3483
rect 4573 3464 4579 3476
rect 4317 3344 4323 3436
rect 4333 3384 4339 3396
rect 4621 3344 4627 3436
rect 4733 3357 4748 3363
rect 4733 3344 4739 3357
rect 4941 3344 4947 3356
rect 5005 3304 5011 3636
rect 6397 3564 6403 3696
rect 6605 3684 6611 3696
rect 5149 3524 5155 3536
rect 5373 3524 5379 3536
rect 5805 3524 5811 3536
rect 5901 3524 5907 3536
rect 6125 3524 6131 3536
rect 6573 3524 6579 3556
rect 5332 3477 5340 3483
rect 6132 3477 6140 3483
rect 5149 3464 5155 3476
rect 5469 3464 5475 3476
rect 5917 3464 5923 3476
rect 5181 3324 5187 3336
rect 5213 3304 5219 3436
rect 5613 3384 5619 3436
rect 5725 3384 5731 3396
rect 6061 3384 6067 3436
rect 6100 3377 6108 3383
rect 6164 3377 6172 3383
rect 5501 3304 5507 3356
rect 5517 3344 5523 3356
rect 5725 3304 5731 3376
rect 5741 3344 5747 3376
rect 6285 3344 6291 3396
rect 6333 3384 6339 3516
rect 6765 3424 6771 3636
rect 6781 3504 6787 3516
rect 7165 3504 7171 3516
rect 7124 3477 7132 3483
rect 6765 3384 6771 3396
rect 6637 3344 6643 3356
rect 6845 3344 6851 3436
rect 6925 3344 6931 3436
rect 7069 3384 7075 3456
rect 7181 3384 7187 3736
rect 7197 3704 7203 3816
rect 7469 3744 7475 3756
rect 7229 3464 7235 3516
rect 7325 3344 7331 3436
rect 7389 3344 7395 3436
rect 7405 3384 7411 3696
rect 7437 3344 7443 3436
rect 7501 3384 7507 3476
rect 7565 3464 7571 3476
rect 5972 3337 6108 3343
rect 6148 3337 6204 3343
rect 6532 3337 6540 3343
rect 5188 3297 5196 3303
rect 6292 3297 6300 3303
rect 5501 3284 5507 3296
rect 6621 3264 6627 3296
rect 6845 3264 6851 3336
rect 4573 3144 4579 3236
rect 4621 3124 4627 3176
rect 5437 3164 5443 3236
rect 5476 3137 5486 3143
rect 5357 3124 5363 3136
rect 5773 3124 5779 3176
rect 5885 3144 5891 3236
rect 6157 3124 6163 3156
rect 6413 3124 6419 3156
rect 6653 3124 6659 3136
rect 6861 3124 6867 3136
rect 4292 3117 4307 3123
rect 4829 3116 4830 3123
rect 3981 3064 3987 3116
rect 4829 3104 4835 3116
rect 5053 3104 5059 3116
rect 5565 3104 5571 3116
rect 4285 3084 4291 3096
rect 6429 3084 6435 3096
rect 4196 3077 4204 3083
rect 4628 3077 4636 3083
rect 3869 2984 3875 3056
rect 4477 3024 4483 3036
rect 4525 2984 4531 3016
rect 4029 2957 4044 2963
rect 4029 2944 4035 2957
rect 4237 2944 4243 2956
rect 3421 2924 3427 2936
rect 3357 2864 3363 2896
rect 3581 2864 3587 2936
rect 3789 2924 3795 2936
rect 3597 2904 3603 2916
rect 4541 2904 4547 3036
rect 4573 2944 4579 3076
rect 4701 2984 4707 2996
rect 4749 2984 4755 3076
rect 5037 3064 5043 3076
rect 5245 3064 5251 3076
rect 5373 3064 5379 3076
rect 6205 3064 6211 3076
rect 6877 3064 6883 3076
rect 4916 3037 4924 3043
rect 4909 2944 4915 2956
rect 4573 2924 4579 2936
rect 4324 2897 4332 2903
rect 3597 2764 3603 2796
rect 3837 2724 3843 2756
rect 4013 2744 4019 2896
rect 4541 2884 4547 2896
rect 4317 2724 4323 2776
rect 4669 2724 4675 2756
rect 3220 2717 3228 2723
rect 3412 2717 3564 2723
rect 3181 2597 3203 2603
rect 3197 2584 3203 2597
rect 2765 2544 2771 2556
rect 2804 2537 2812 2543
rect 3021 2504 3027 2556
rect 3373 2544 3379 2716
rect 4221 2704 4227 2716
rect 3565 2664 3571 2676
rect 3645 2644 3651 2696
rect 4308 2677 4316 2683
rect 3789 2664 3795 2676
rect 3421 2564 3427 2636
rect 3437 2584 3443 2596
rect 3613 2544 3619 2556
rect 3645 2544 3651 2636
rect 3661 2584 3667 2596
rect 3869 2584 3875 2616
rect 3837 2544 3843 2556
rect 3373 2524 3379 2536
rect 3885 2504 3891 2636
rect 4301 2544 4307 2556
rect 4084 2537 4092 2543
rect 4109 2504 4115 2536
rect 4317 2504 4323 2556
rect 4477 2544 4483 2636
rect 4493 2584 4499 2696
rect 4877 2684 4883 2756
rect 4973 2744 4979 3036
rect 4989 2984 4995 3036
rect 5645 2984 5651 3056
rect 7069 3044 7075 3296
rect 7213 3084 7219 3096
rect 7277 3084 7283 3316
rect 7309 3304 7315 3336
rect 7661 3323 7667 4276
rect 7709 4184 7715 4316
rect 7885 4304 7891 4356
rect 8477 4344 8483 4496
rect 7885 4284 7891 4296
rect 7917 4264 7923 4316
rect 7741 4224 7747 4236
rect 7837 4144 7843 4156
rect 7949 4144 7955 4256
rect 7965 4144 7971 4236
rect 8109 4184 8115 4316
rect 8413 4304 8419 4316
rect 8429 4284 8435 4336
rect 8541 4324 8547 4497
rect 8333 4204 8339 4236
rect 8285 4157 8316 4163
rect 8285 4144 8291 4157
rect 8493 4144 8499 4196
rect 8525 4184 8531 4196
rect 8605 4184 8611 4496
rect 8813 4384 8819 4496
rect 8813 4184 8819 4356
rect 8829 4324 8835 4336
rect 8925 4324 8931 4636
rect 9229 4544 9235 4556
rect 9213 4504 9219 4536
rect 9133 4484 9139 4496
rect 9181 4324 9187 4436
rect 8845 4284 8851 4296
rect 8957 4144 8963 4156
rect 7837 4124 7843 4136
rect 8733 4124 8739 4136
rect 7933 4104 7939 4116
rect 7837 4084 7843 4096
rect 8733 4084 8739 4096
rect 8989 3964 8995 4236
rect 9133 4184 9139 4276
rect 9165 4264 9171 4276
rect 9149 4184 9155 4256
rect 9213 4184 9219 4336
rect 9357 4324 9363 4436
rect 9389 4304 9395 4636
rect 10029 4584 10035 4596
rect 9549 4544 9555 4556
rect 10205 4544 10211 4636
rect 9780 4537 9788 4543
rect 9853 4504 9859 4536
rect 10253 4504 10259 4636
rect 9549 4364 9555 4496
rect 9885 4464 9891 4496
rect 9613 4324 9619 4336
rect 9853 4324 9859 4336
rect 9421 4284 9427 4316
rect 9828 4277 9836 4283
rect 9037 4124 9043 4156
rect 9037 4104 9043 4116
rect 9069 3964 9075 4136
rect 7901 3924 7907 3936
rect 8541 3924 8547 3936
rect 8893 3924 8899 3956
rect 9133 3924 9139 4096
rect 9261 4064 9267 4236
rect 9613 4203 9619 4276
rect 9901 4243 9907 4316
rect 9933 4284 9939 4296
rect 9885 4237 9907 4243
rect 9613 4197 9635 4203
rect 9629 4184 9635 4197
rect 9501 4144 9507 4176
rect 9693 4144 9699 4236
rect 9885 4184 9891 4237
rect 10061 4204 10067 4236
rect 9908 4137 9916 4143
rect 9277 4124 9283 4136
rect 9476 4117 9484 4123
rect 9485 4104 9491 4116
rect 9709 4104 9715 4116
rect 9917 4084 9923 4096
rect 9581 3984 9587 4076
rect 9437 3924 9443 3936
rect 7677 3864 7683 3916
rect 7693 3884 7699 3896
rect 8093 3884 8099 3916
rect 8477 3884 8483 3916
rect 9101 3884 9107 3896
rect 8452 3877 8460 3883
rect 7828 3837 7836 3843
rect 7917 3784 7923 3876
rect 7860 3737 7868 3743
rect 7885 3684 7891 3696
rect 7677 3524 7683 3556
rect 8109 3484 8115 3736
rect 8125 3663 8131 3876
rect 8317 3784 8323 3836
rect 8477 3824 8483 3876
rect 8365 3784 8371 3816
rect 8173 3744 8179 3756
rect 8605 3744 8611 3756
rect 8701 3744 8707 3836
rect 8733 3804 8739 3836
rect 8765 3784 8771 3876
rect 8141 3684 8147 3696
rect 8125 3657 8147 3663
rect 8125 3524 8131 3616
rect 7693 3464 7699 3476
rect 7821 3384 7827 3436
rect 8125 3384 8131 3476
rect 7709 3344 7715 3376
rect 7661 3317 7683 3323
rect 7645 3284 7651 3296
rect 7437 3063 7443 3116
rect 7677 3084 7683 3317
rect 7709 3304 7715 3336
rect 7741 3244 7747 3336
rect 7965 3324 7971 3336
rect 7949 3284 7955 3296
rect 7524 3077 7532 3083
rect 7421 3057 7443 3063
rect 5565 2944 5571 2956
rect 5725 2944 5731 3036
rect 5805 2957 5820 2963
rect 5805 2944 5811 2957
rect 5149 2903 5155 2936
rect 5140 2897 5155 2903
rect 4973 2724 4979 2736
rect 4893 2704 4899 2716
rect 4973 2684 4979 2696
rect 4596 2677 4668 2683
rect 4557 2544 4563 2636
rect 4749 2624 4755 2636
rect 5133 2564 5139 2836
rect 5165 2704 5171 2936
rect 5357 2924 5363 2936
rect 6061 2904 6067 3036
rect 6141 2984 6147 3036
rect 6573 2964 6579 3036
rect 6253 2944 6259 2956
rect 6813 2944 6819 3036
rect 6925 2903 6931 3036
rect 7005 3004 7011 3036
rect 7021 3024 7027 3036
rect 6973 2904 6979 2976
rect 7229 2944 7235 2996
rect 7293 2984 7299 3036
rect 7005 2924 7011 2936
rect 6916 2897 6931 2903
rect 5181 2724 5187 2736
rect 5197 2664 5203 2676
rect 5613 2664 5619 2716
rect 5380 2637 5388 2643
rect 5149 2604 5155 2636
rect 5485 2584 5491 2656
rect 5789 2624 5795 2896
rect 6061 2884 6067 2896
rect 6445 2784 6451 2896
rect 6493 2724 6499 2836
rect 6637 2724 6643 2736
rect 6717 2724 6723 2776
rect 6749 2724 6755 2836
rect 7101 2784 7107 2896
rect 6621 2684 6627 2696
rect 5837 2664 5843 2676
rect 6269 2664 6275 2676
rect 5901 2584 5907 2596
rect 5981 2564 5987 2636
rect 4765 2544 4771 2556
rect 6205 2544 6211 2556
rect 6477 2544 6483 2636
rect 6557 2584 6563 2656
rect 6653 2584 6659 2676
rect 6941 2664 6947 2676
rect 6829 2584 6835 2596
rect 6756 2537 6764 2543
rect 5085 2524 5091 2536
rect 5757 2524 5763 2536
rect 4541 2504 4547 2516
rect 6189 2504 6195 2516
rect 6397 2504 6403 2536
rect 6781 2504 6787 2576
rect 6877 2544 6883 2636
rect 7133 2604 7139 2716
rect 7149 2684 7155 2796
rect 7165 2704 7171 2836
rect 7357 2724 7363 3056
rect 7421 2984 7427 3057
rect 7565 2944 7571 2956
rect 7597 2904 7603 2996
rect 7661 2764 7667 3036
rect 7677 2964 7683 3076
rect 7709 3024 7715 3036
rect 7789 2984 7795 2996
rect 7869 2984 7875 3236
rect 7885 3124 7891 3236
rect 8084 3117 8092 3123
rect 7917 3064 7923 3076
rect 7693 2943 7699 2956
rect 7684 2937 7699 2943
rect 7997 2937 8012 2943
rect 7876 2897 7884 2903
rect 7997 2884 8003 2937
rect 8013 2904 8019 2916
rect 7565 2724 7571 2756
rect 7789 2724 7795 2736
rect 8061 2724 8067 3076
rect 8093 3064 8099 3116
rect 8141 3004 8147 3657
rect 8381 3584 8387 3696
rect 8573 3524 8579 3576
rect 8781 3524 8787 3876
rect 9133 3844 9139 3916
rect 9213 3864 9219 3876
rect 8973 3804 8979 3836
rect 9357 3764 9363 3836
rect 9277 3744 9283 3756
rect 8829 3704 8835 3716
rect 9181 3704 9187 3716
rect 9261 3704 9267 3716
rect 9469 3704 9475 3716
rect 9021 3524 9027 3556
rect 8493 3504 8499 3516
rect 9229 3504 9235 3516
rect 8269 3384 8275 3436
rect 8349 3384 8355 3476
rect 8477 3464 8483 3476
rect 8573 3464 8579 3476
rect 9021 3464 9027 3476
rect 8429 3344 8435 3356
rect 8429 3304 8435 3316
rect 8381 3124 8387 3296
rect 8589 3223 8595 3436
rect 8717 3344 8723 3436
rect 9037 3384 9043 3496
rect 9245 3484 9251 3496
rect 9069 3344 9075 3436
rect 9165 3344 9171 3436
rect 9389 3344 9395 3436
rect 9613 3344 9619 3436
rect 9629 3384 9635 4016
rect 10077 3964 10083 4436
rect 9652 3897 9667 3903
rect 9661 3884 9667 3897
rect 9693 3744 9699 3756
rect 9821 3744 9827 3836
rect 9853 3784 9859 3916
rect 9885 3884 9891 3956
rect 10013 3744 10019 3836
rect 10077 3784 10083 3916
rect 10093 3784 10099 3796
rect 10237 3744 10243 3836
rect 9853 3704 9859 3716
rect 9677 3524 9683 3536
rect 9901 3524 9907 3536
rect 9917 3484 9923 3736
rect 10100 3517 10108 3523
rect 9837 3344 9843 3356
rect 8653 3324 8659 3336
rect 8653 3304 8659 3316
rect 9901 3304 9907 3476
rect 10045 3344 10051 3436
rect 8573 3217 8595 3223
rect 8573 3184 8579 3217
rect 8989 3144 8995 3156
rect 8285 3084 8291 3116
rect 8301 3004 8307 3116
rect 8237 2984 8243 2996
rect 8461 2984 8467 2996
rect 8077 2904 8083 2976
rect 8093 2924 8099 2936
rect 8333 2924 8339 2936
rect 8125 2684 8131 2716
rect 8205 2704 8211 2716
rect 7197 2557 7212 2563
rect 7197 2544 7203 2557
rect 6957 2524 6963 2536
rect 3636 2497 3644 2503
rect 5972 2497 5980 2503
rect 6964 2497 6972 2503
rect 2413 2264 2419 2276
rect 2285 2104 2291 2236
rect 2477 2104 2483 2316
rect 2493 2184 2499 2496
rect 2852 2317 2860 2323
rect 2509 2304 2515 2316
rect 2877 2284 2883 2496
rect 3389 2484 3395 2496
rect 5533 2484 5539 2496
rect 7405 2484 7411 2536
rect 7421 2504 7427 2556
rect 5309 2464 5315 2476
rect 3101 2324 3107 2436
rect 3165 2343 3171 2436
rect 4692 2357 4700 2363
rect 3149 2337 3171 2343
rect 2941 2244 2947 2276
rect 2669 2224 2675 2236
rect 2061 2084 2067 2096
rect 1885 1924 1891 1936
rect 2237 1924 2243 1956
rect 2477 1944 2483 2096
rect 2685 2064 2691 2096
rect 2333 1924 2339 1936
rect 2338 1917 2339 1924
rect 2269 1884 2275 1916
rect 2685 1903 2691 1956
rect 2701 1924 2707 1936
rect 2685 1897 2707 1903
rect 1876 1877 1884 1883
rect 2685 1864 2691 1876
rect 1885 1784 1891 1796
rect 1869 1704 1875 1736
rect 2093 1724 2099 1836
rect 2461 1824 2467 1836
rect 2701 1803 2707 1897
rect 2717 1884 2723 2236
rect 2909 2144 2915 2156
rect 2941 1884 2947 2236
rect 3021 2144 3027 2156
rect 3149 2143 3155 2337
rect 3725 2324 3731 2356
rect 3933 2324 3939 2336
rect 4029 2324 4035 2336
rect 4397 2324 4403 2336
rect 3172 2317 3180 2323
rect 3492 2317 3500 2323
rect 4477 2317 4492 2323
rect 3149 2137 3171 2143
rect 2685 1797 2707 1803
rect 2477 1744 2483 1756
rect 2269 1704 2275 1736
rect 2029 1684 2035 1696
rect 2685 1683 2691 1797
rect 2941 1784 2947 1816
rect 2701 1744 2707 1756
rect 2797 1744 2803 1756
rect 2797 1704 2803 1716
rect 2685 1677 2707 1683
rect 2093 1524 2099 1536
rect 2333 1524 2339 1536
rect 2541 1524 2547 1536
rect 2338 1517 2339 1524
rect 1837 1384 1843 1516
rect 1860 1477 1868 1483
rect 2548 1477 2556 1483
rect 2701 1483 2707 1677
rect 2941 1524 2947 1696
rect 2685 1477 2707 1483
rect 2020 1337 2028 1343
rect 2045 1323 2051 1436
rect 2253 1384 2259 1416
rect 2685 1383 2691 1477
rect 2916 1477 2924 1483
rect 2701 1404 2707 1436
rect 2685 1377 2700 1383
rect 2916 1377 2924 1383
rect 2109 1344 2115 1356
rect 2445 1344 2451 1356
rect 2989 1344 2995 2096
rect 3005 2084 3011 2096
rect 3165 2084 3171 2137
rect 3181 1904 3187 2276
rect 3485 2264 3491 2276
rect 3572 2237 3580 2243
rect 3245 2084 3251 2096
rect 3389 2024 3395 2036
rect 3021 1864 3027 1876
rect 3037 1744 3043 1756
rect 3021 1664 3027 1696
rect 3149 1464 3155 1516
rect 3197 1344 3203 1876
rect 3213 1784 3219 1936
rect 3373 1924 3379 1956
rect 3373 1864 3379 1876
rect 3229 1724 3235 1836
rect 3405 1764 3411 2236
rect 3421 2184 3427 2236
rect 3629 2184 3635 2276
rect 3933 2264 3939 2276
rect 3597 2144 3603 2156
rect 3828 2137 3836 2143
rect 3629 1944 3635 2096
rect 3853 1964 3859 2096
rect 3405 1744 3411 1756
rect 3380 1697 3388 1703
rect 3373 1484 3379 1516
rect 3437 1484 3443 1836
rect 3629 1784 3635 1916
rect 3821 1884 3827 1956
rect 3853 1884 3859 1916
rect 3485 1724 3491 1736
rect 3476 1697 3484 1703
rect 3661 1524 3667 1776
rect 3677 1664 3683 1836
rect 3837 1784 3843 1796
rect 3693 1724 3699 1736
rect 3693 1684 3699 1696
rect 3869 1524 3875 2216
rect 4077 2184 4083 2276
rect 4397 2263 4403 2276
rect 4397 2257 4419 2263
rect 4413 2244 4419 2257
rect 4189 2224 4195 2236
rect 4061 2144 4067 2176
rect 4477 2144 4483 2317
rect 4861 2284 4867 2316
rect 4925 2304 4931 2316
rect 4941 2284 4947 2296
rect 5149 2284 5155 2356
rect 5517 2324 5523 2336
rect 5357 2284 5363 2296
rect 4573 2144 4579 2156
rect 4308 2137 4316 2143
rect 4493 2104 4499 2116
rect 4077 1924 4083 1956
rect 4285 1924 4291 1936
rect 4077 1784 4083 1876
rect 4269 1824 4275 1876
rect 4301 1844 4307 2096
rect 4493 1924 4499 1936
rect 4509 1884 4515 2096
rect 4301 1764 4307 1836
rect 3901 1744 3907 1756
rect 4253 1744 4259 1756
rect 3901 1704 3907 1716
rect 3933 1484 3939 1536
rect 4077 1524 4083 1536
rect 3389 1384 3395 1456
rect 3469 1404 3475 1436
rect 3421 1384 3427 1396
rect 3426 1377 3427 1384
rect 3533 1344 3539 1476
rect 3597 1464 3603 1476
rect 3629 1424 3635 1436
rect 3645 1384 3651 1476
rect 4301 1444 4307 1476
rect 2029 1317 2051 1323
rect 2029 1304 2035 1317
rect 1837 1184 1843 1236
rect 1837 1124 1843 1156
rect 2013 1104 2019 1116
rect 1764 1077 1772 1083
rect 2004 1077 2012 1083
rect 1629 1024 1635 1036
rect 1773 984 1779 996
rect 1405 924 1411 976
rect 1773 964 1779 976
rect 1837 963 1843 976
rect 1837 957 1859 963
rect 1533 944 1539 956
rect 1645 924 1651 936
rect 1853 924 1859 957
rect 1869 944 1875 956
rect 1629 904 1635 916
rect 1597 784 1603 836
rect 1533 724 1539 736
rect 1741 724 1747 876
rect 2045 724 2051 1296
rect 2093 1124 2099 1336
rect 2445 1324 2451 1336
rect 2477 1304 2483 1336
rect 2557 1324 2563 1336
rect 2564 1297 2572 1303
rect 2973 1284 2979 1296
rect 3117 1284 3123 1296
rect 2669 1124 2675 1156
rect 2877 1124 2883 1136
rect 3165 1124 3171 1156
rect 3325 1124 3331 1156
rect 2093 1104 2099 1116
rect 2477 1084 2483 1116
rect 2669 1084 2675 1096
rect 2893 1084 2899 1096
rect 3085 1084 3091 1096
rect 2109 1064 2115 1076
rect 2077 984 2083 1016
rect 1741 684 1747 696
rect 1949 684 1955 696
rect 2036 677 2044 683
rect 1565 544 1571 556
rect 1565 464 1571 496
rect 1789 484 1795 536
rect 1805 504 1811 516
rect 1821 484 1827 636
rect 420 317 428 323
rect 868 317 876 323
rect 189 284 195 296
rect 893 284 899 456
rect 1069 324 1075 336
rect 1533 324 1539 356
rect 1837 324 1843 516
rect 1869 504 1875 636
rect 2061 584 2067 956
rect 2237 904 2243 1036
rect 2260 977 2268 983
rect 2285 944 2291 956
rect 2477 943 2483 996
rect 2925 984 2931 1036
rect 3117 1004 3123 1036
rect 3341 984 3347 1076
rect 2452 937 2483 943
rect 2477 784 2483 896
rect 2493 763 2499 976
rect 2941 944 2947 976
rect 2973 944 2979 956
rect 3197 944 3203 956
rect 2653 924 2659 936
rect 2765 924 2771 936
rect 2653 883 2659 916
rect 2669 904 2675 916
rect 2749 904 2755 916
rect 2941 904 2947 936
rect 2653 877 2675 883
rect 2477 757 2499 763
rect 2477 724 2483 757
rect 2637 724 2643 736
rect 2669 684 2675 877
rect 2893 844 2899 856
rect 2893 724 2899 836
rect 3085 724 3091 896
rect 3181 884 3187 896
rect 3101 824 3107 836
rect 3373 724 3379 1136
rect 3421 1084 3427 1216
rect 3565 1144 3571 1296
rect 3533 984 3539 996
rect 3389 724 3395 896
rect 3597 784 3603 1376
rect 3773 1324 3779 1336
rect 3805 1304 3811 1356
rect 4061 1344 4067 1436
rect 4237 1344 4243 1356
rect 4285 1304 4291 1436
rect 3773 1184 3779 1196
rect 4045 1184 4051 1296
rect 3773 1177 3774 1184
rect 4013 1124 4019 1156
rect 3629 1064 3635 1116
rect 3997 1064 4003 1076
rect 3613 984 3619 996
rect 3773 984 3779 1016
rect 4045 984 4051 1036
rect 4061 944 4067 1236
rect 4205 1124 4211 1136
rect 4285 984 4291 1136
rect 4301 1124 4307 1436
rect 4317 1384 4323 1856
rect 4477 1684 4483 1696
rect 4493 1524 4499 1856
rect 4477 1464 4483 1476
rect 4445 1124 4451 1156
rect 4461 1084 4467 1336
rect 4429 1044 4435 1076
rect 4509 984 4515 1876
rect 4541 1704 4547 2136
rect 4573 2084 4579 2096
rect 4733 1924 4739 1936
rect 4749 1924 4755 2256
rect 4941 2184 4947 2256
rect 4973 2184 4979 2196
rect 5053 1923 5059 2096
rect 5229 1924 5235 2256
rect 5389 2064 5395 2136
rect 5421 2104 5427 2236
rect 5485 2184 5491 2196
rect 5533 2184 5539 2476
rect 5789 2204 5795 2316
rect 5805 2284 5811 2456
rect 6029 2324 6035 2336
rect 7469 2324 7475 2636
rect 7501 2584 7507 2616
rect 7581 2564 7587 2676
rect 8237 2664 8243 2676
rect 7933 2604 7939 2636
rect 7661 2584 7667 2596
rect 7853 2544 7859 2556
rect 7981 2544 7987 2636
rect 8077 2544 8083 2596
rect 8109 2584 8115 2596
rect 7885 2504 7891 2536
rect 8285 2504 8291 2516
rect 8077 2404 8083 2496
rect 8125 2384 8131 2396
rect 6692 2317 6700 2323
rect 7332 2317 7340 2323
rect 6237 2284 6243 2316
rect 6253 2304 6259 2316
rect 6029 2264 6035 2276
rect 5869 2184 5875 2196
rect 5613 2144 5619 2156
rect 5725 2124 5731 2136
rect 5949 2104 5955 2236
rect 5965 2144 5971 2236
rect 6477 2204 6483 2316
rect 7133 2304 7139 2316
rect 7565 2284 7571 2296
rect 7773 2284 7779 2316
rect 7789 2284 7795 2336
rect 7965 2324 7971 2336
rect 8004 2277 8012 2283
rect 6925 2264 6931 2276
rect 7133 2264 7139 2276
rect 6525 2184 6531 2196
rect 6621 2144 6627 2236
rect 6973 2184 6979 2256
rect 7069 2224 7075 2236
rect 7181 2184 7187 2256
rect 7357 2204 7363 2276
rect 7405 2184 7411 2196
rect 7661 2184 7667 2276
rect 7709 2224 7715 2236
rect 7405 2177 7406 2184
rect 7277 2144 7283 2156
rect 7709 2144 7715 2196
rect 7853 2184 7859 2256
rect 7485 2124 7491 2136
rect 6589 2104 6595 2116
rect 5732 2097 5740 2103
rect 5037 1917 5059 1923
rect 4717 1864 4723 1876
rect 4701 1784 4707 1796
rect 4557 1744 4563 1756
rect 4541 1644 4547 1696
rect 4580 1517 4588 1523
rect 4548 1377 4556 1383
rect 4589 1364 4595 1476
rect 4749 1424 4755 1916
rect 4813 1884 4819 1916
rect 4941 1764 4947 1836
rect 5037 1784 5043 1917
rect 5181 1904 5187 1916
rect 5476 1877 5484 1883
rect 5149 1744 5155 1756
rect 4797 1704 4803 1716
rect 5165 1704 5171 1836
rect 5629 1804 5635 1836
rect 5485 1744 5491 1796
rect 4765 1584 4771 1636
rect 5181 1584 5187 1696
rect 5213 1584 5219 1656
rect 5218 1577 5219 1584
rect 4781 1504 4787 1516
rect 4525 1304 4531 1316
rect 4692 1297 4700 1303
rect 4532 1117 4540 1123
rect 4557 1084 4563 1156
rect 4189 924 4195 936
rect 3085 704 3091 716
rect 2868 677 2876 683
rect 3076 677 3084 683
rect 2397 664 2403 676
rect 2205 624 2211 636
rect 1885 544 1891 556
rect 2237 544 2243 556
rect 1869 484 1875 496
rect 2269 364 2275 636
rect 2461 584 2467 596
rect 2701 584 2707 616
rect 2333 544 2339 556
rect 2557 544 2563 556
rect 2301 504 2307 516
rect 2477 444 2483 496
rect 2189 324 2195 356
rect 2445 324 2451 436
rect 2717 324 2723 636
rect 3309 624 3315 636
rect 2877 544 2883 596
rect 2964 557 2972 563
rect 3101 544 3107 556
rect 3357 544 3363 576
rect 3517 544 3523 636
rect 3565 544 3571 556
rect 3188 537 3196 543
rect 3133 504 3139 536
rect 3341 504 3347 536
rect 3597 504 3603 636
rect 3757 564 3763 716
rect 3677 544 3683 556
rect 3773 544 3779 896
rect 4189 884 4195 896
rect 4029 783 4035 876
rect 4029 777 4044 783
rect 3821 724 3827 736
rect 3821 664 3827 676
rect 3789 584 3795 596
rect 3789 577 3790 584
rect 3965 544 3971 636
rect 4205 544 4211 716
rect 4253 584 4259 836
rect 4269 784 4275 956
rect 4637 944 4643 1036
rect 4413 743 4419 936
rect 4653 904 4659 936
rect 4429 884 4435 896
rect 4397 737 4419 743
rect 4397 684 4403 737
rect 4413 684 4419 716
rect 4429 704 4435 876
rect 4637 724 4643 736
rect 4445 544 4451 556
rect 2893 484 2899 496
rect 1741 284 1747 296
rect 1268 277 1276 283
rect 413 264 419 276
rect 1069 264 1075 276
rect 932 237 947 243
rect 61 124 67 236
rect 493 204 499 236
rect 93 144 99 156
rect 301 144 307 196
rect 701 144 707 236
rect 749 184 755 236
rect 925 144 931 216
rect 941 104 947 237
rect 989 104 995 256
rect 1149 224 1155 236
rect 1197 184 1203 276
rect 1357 224 1363 236
rect 1005 144 1011 156
rect 1357 144 1363 156
rect 1005 124 1011 136
rect 1389 104 1395 156
rect 1453 144 1459 196
rect 1533 144 1539 276
rect 1757 264 1763 296
rect 1837 284 1843 296
rect 2413 284 2419 296
rect 2845 284 2851 336
rect 3101 324 3107 356
rect 3309 324 3315 396
rect 3533 324 3539 356
rect 3773 324 3779 336
rect 3821 324 3827 516
rect 4125 484 4131 536
rect 4477 524 4483 696
rect 4637 604 4643 676
rect 4701 584 4707 796
rect 4717 784 4723 1416
rect 4765 1384 4771 1396
rect 4813 1384 4819 1476
rect 4781 1104 4787 1116
rect 4797 1064 4803 1076
rect 4733 984 4739 996
rect 4861 684 4867 936
rect 4893 904 4899 916
rect 4925 904 4931 1296
rect 4893 704 4899 896
rect 4941 724 4947 1096
rect 4957 984 4963 1516
rect 5005 1504 5011 1516
rect 5021 1364 5027 1476
rect 5149 1384 5155 1416
rect 5005 1124 5011 1296
rect 5021 1164 5027 1336
rect 5165 1184 5171 1536
rect 5357 1484 5363 1516
rect 5341 1464 5347 1476
rect 5373 1384 5379 1696
rect 5213 1284 5219 1296
rect 5005 1104 5011 1116
rect 5021 984 5027 1076
rect 5341 1063 5347 1296
rect 5357 1104 5363 1116
rect 5364 1077 5372 1083
rect 5341 1057 5363 1063
rect 5341 984 5347 1036
rect 5357 1024 5363 1057
rect 5421 984 5427 1716
rect 5597 1484 5603 1516
rect 5645 1384 5651 2096
rect 5885 1984 5891 2096
rect 6381 2084 6387 2096
rect 7261 2084 7267 2096
rect 6957 1984 6963 2016
rect 7389 1984 7395 2096
rect 7485 2084 7491 2096
rect 7693 2084 7699 2096
rect 6804 1937 6956 1943
rect 7028 1937 7180 1943
rect 7252 1937 7404 1943
rect 5716 1917 5724 1923
rect 6788 1917 6796 1923
rect 5933 1884 5939 1896
rect 6285 1884 6291 1916
rect 5789 1744 5795 1856
rect 5821 1784 5827 1816
rect 5901 1744 5907 1756
rect 5677 1664 5683 1736
rect 5789 1464 5795 1476
rect 5661 1384 5667 1416
rect 5821 1344 5827 1476
rect 5812 1337 5820 1343
rect 5453 1284 5459 1296
rect 5805 1264 5811 1296
rect 5677 1123 5683 1156
rect 5677 1117 5692 1123
rect 5581 984 5587 1016
rect 5101 864 5107 896
rect 5181 824 5187 896
rect 5213 884 5219 936
rect 5597 904 5603 1036
rect 5677 964 5683 1117
rect 5789 924 5795 936
rect 5869 924 5875 1736
rect 5885 1684 5891 1696
rect 6045 1584 6051 1856
rect 6269 1823 6275 1876
rect 6269 1817 6291 1823
rect 6285 1784 6291 1817
rect 6237 1524 6243 1656
rect 5885 1504 5891 1516
rect 6301 1464 6307 1876
rect 6685 1864 6691 1876
rect 6685 1744 6691 1756
rect 6781 1744 6787 1896
rect 6813 1884 6819 1896
rect 6685 1724 6691 1736
rect 6493 1584 6499 1696
rect 6484 1517 6492 1523
rect 6061 1344 6067 1456
rect 6093 1344 6099 1436
rect 5901 1264 5907 1296
rect 6061 1184 6067 1336
rect 6301 1184 6307 1456
rect 6509 1384 6515 1636
rect 6701 1524 6707 1536
rect 6797 1524 6803 1736
rect 6788 1517 6796 1523
rect 6797 1484 6803 1496
rect 6685 1464 6691 1476
rect 6717 1384 6723 1456
rect 6925 1444 6931 1536
rect 6957 1524 6963 1836
rect 6973 1784 6979 1916
rect 7037 1864 7043 1876
rect 7181 1784 7187 1916
rect 7469 1884 7475 1976
rect 7661 1924 7667 1956
rect 7677 1884 7683 1896
rect 6989 1704 6995 1776
rect 7341 1744 7347 1876
rect 7021 1724 7027 1736
rect 7373 1704 7379 1876
rect 7245 1524 7251 1536
rect 7597 1524 7603 1836
rect 7805 1824 7811 1836
rect 7645 1784 7651 1796
rect 7844 1717 7852 1723
rect 7805 1704 7811 1716
rect 7869 1703 7875 2156
rect 7933 2144 7939 2216
rect 8061 2184 8067 2236
rect 8173 2224 8179 2236
rect 8301 2184 8307 2276
rect 8349 2223 8355 2636
rect 8381 2504 8387 2836
rect 8525 2744 8531 3036
rect 8541 2904 8547 3136
rect 9053 3124 9059 3296
rect 9837 3184 9843 3296
rect 9204 3117 9212 3123
rect 8717 2984 8723 3116
rect 8813 3044 8819 3076
rect 8557 2924 8563 2936
rect 8941 2904 8947 3036
rect 8941 2884 8947 2896
rect 8429 2704 8435 2716
rect 8621 2684 8627 2856
rect 8957 2724 8963 3036
rect 8989 2984 8995 3116
rect 9245 3104 9251 3116
rect 9485 3104 9491 3116
rect 9252 3077 9260 3083
rect 9021 3044 9027 3076
rect 9485 3064 9491 3076
rect 9629 3004 9635 3036
rect 9133 2944 9139 2956
rect 9373 2944 9379 2956
rect 9581 2944 9587 2996
rect 9373 2904 9379 2916
rect 9613 2904 9619 2976
rect 9661 2924 9667 3096
rect 10036 3077 10044 3083
rect 9901 2944 9907 3036
rect 10061 2984 10067 3116
rect 9917 2924 9923 2936
rect 9677 2884 9683 2896
rect 8845 2684 8851 2716
rect 8445 2564 8451 2676
rect 8589 2544 8595 2556
rect 8413 2284 8419 2316
rect 8397 2264 8403 2276
rect 8333 2217 8355 2223
rect 8285 1984 8291 2096
rect 8333 1984 8339 2217
rect 8493 2184 8499 2276
rect 8589 2164 8595 2496
rect 8749 2444 8755 2676
rect 8765 2584 8771 2676
rect 8861 2644 8867 2676
rect 8765 2384 8771 2516
rect 8781 2504 8787 2576
rect 8957 2484 8963 2636
rect 9005 2544 9011 2636
rect 9053 2544 9059 2636
rect 9149 2584 9155 2596
rect 9149 2577 9150 2584
rect 9037 2503 9043 2516
rect 9028 2497 9043 2503
rect 8621 2324 8627 2336
rect 8781 2284 8787 2436
rect 8957 2324 8963 2476
rect 9181 2324 9187 2876
rect 9437 2724 9443 2836
rect 9204 2717 9219 2723
rect 9213 2684 9219 2717
rect 9197 2644 9203 2676
rect 9213 2664 9219 2676
rect 9389 2584 9395 2676
rect 9437 2664 9443 2716
rect 9517 2704 9523 2796
rect 9661 2724 9667 2736
rect 9517 2684 9523 2696
rect 9245 2524 9251 2536
rect 9597 2524 9603 2536
rect 9229 2503 9235 2516
rect 9229 2497 9244 2503
rect 9597 2484 9603 2496
rect 9277 2324 9283 2336
rect 9469 2324 9475 2436
rect 9282 2317 9283 2324
rect 9165 2284 9171 2316
rect 9181 2304 9187 2316
rect 9268 2277 9276 2283
rect 8637 2184 8643 2276
rect 8676 2137 8684 2143
rect 8365 2124 8371 2136
rect 8701 2104 8707 2156
rect 9037 2144 9043 2236
rect 9133 2144 9139 2156
rect 8765 2104 8771 2136
rect 8493 1984 8499 2016
rect 8125 1884 8131 1896
rect 8365 1884 8371 1956
rect 8797 1944 8803 2136
rect 9421 2124 9427 2236
rect 9453 2164 9459 2236
rect 9469 2144 9475 2156
rect 9181 2104 9187 2116
rect 9156 2097 9164 2103
rect 9474 2096 9475 2103
rect 9469 1984 9475 2096
rect 8589 1924 8595 1936
rect 9149 1924 9155 1936
rect 9245 1924 9251 1956
rect 9629 1924 9635 2576
rect 9885 2544 9891 2916
rect 9908 2897 9916 2903
rect 9917 2784 9923 2796
rect 9949 2684 9955 2696
rect 10125 2684 10131 3476
rect 10077 2584 10083 2596
rect 9869 2484 9875 2496
rect 9821 2304 9827 2316
rect 9677 2144 9683 2236
rect 9885 2164 9891 2536
rect 9901 2324 9907 2336
rect 9917 2244 9923 2276
rect 10061 2144 10067 2236
rect 10237 2184 10243 2196
rect 9885 2124 9891 2136
rect 9661 1884 9667 1896
rect 8573 1864 8579 1876
rect 8269 1744 8275 1836
rect 8317 1784 8323 1836
rect 8381 1744 8387 1756
rect 7917 1724 7923 1736
rect 7853 1697 7875 1703
rect 7460 1517 7468 1523
rect 7469 1484 7475 1496
rect 7693 1484 7699 1496
rect 7021 1464 7027 1476
rect 7245 1464 7251 1476
rect 6925 1384 6931 1436
rect 6941 1384 6947 1396
rect 6349 1324 6355 1336
rect 6573 1324 6579 1336
rect 6797 1324 6803 1336
rect 7005 1304 7011 1376
rect 7165 1343 7171 1436
rect 7380 1377 7388 1383
rect 7165 1337 7180 1343
rect 7037 1324 7043 1336
rect 6349 1284 6355 1296
rect 6541 1284 6547 1296
rect 6797 1284 6803 1296
rect 6557 1184 6563 1276
rect 7405 1264 7411 1436
rect 7853 1384 7859 1697
rect 8148 1697 8156 1703
rect 8301 1684 8307 1696
rect 8061 1644 8067 1656
rect 8061 1623 8067 1636
rect 8045 1617 8067 1623
rect 8045 1524 8051 1617
rect 8461 1524 8467 1536
rect 8541 1524 8547 1836
rect 8749 1764 8755 1836
rect 8813 1824 8819 1876
rect 8941 1784 8947 1816
rect 8957 1763 8963 1836
rect 9133 1824 9139 1876
rect 9437 1764 9443 1836
rect 9677 1824 9683 1916
rect 9805 1784 9811 1816
rect 8941 1757 8963 1763
rect 8589 1704 8595 1736
rect 8749 1664 8755 1696
rect 8237 1484 8243 1496
rect 8253 1484 8259 1516
rect 8893 1504 8899 1516
rect 8941 1484 8947 1757
rect 9021 1744 9027 1756
rect 9869 1744 9875 1936
rect 9885 1904 9891 1916
rect 10100 1877 10108 1883
rect 10269 1823 10275 3696
rect 10253 1817 10275 1823
rect 10221 1784 10227 1796
rect 9444 1737 9452 1743
rect 8957 1704 8963 1736
rect 8973 1484 8979 1496
rect 9412 1477 9420 1483
rect 7869 1384 7875 1436
rect 8013 1384 8019 1476
rect 7597 1304 7603 1316
rect 7661 1304 7667 1376
rect 7693 1324 7699 1336
rect 7917 1324 7923 1336
rect 7597 1284 7603 1296
rect 6813 1184 6819 1196
rect 5924 1137 5955 1143
rect 5949 1124 5955 1137
rect 6381 1124 6387 1136
rect 6621 1124 6627 1136
rect 7453 1124 7459 1236
rect 7485 1124 7491 1136
rect 6148 1117 6156 1123
rect 5917 1063 5923 1116
rect 5933 1084 5939 1116
rect 6957 1104 6963 1116
rect 6317 1084 6323 1096
rect 6148 1077 6156 1083
rect 6077 1063 6083 1076
rect 5917 1057 6083 1063
rect 6525 984 6531 1096
rect 7709 1084 7715 1096
rect 6957 1044 6963 1076
rect 7069 1064 7075 1076
rect 7389 1064 7395 1076
rect 6765 964 6771 1036
rect 6893 944 6899 956
rect 7133 944 7139 956
rect 7453 944 7459 976
rect 5892 937 5900 943
rect 6132 937 6140 943
rect 6564 937 6572 943
rect 5421 784 5427 816
rect 5101 724 5107 736
rect 5581 724 5587 896
rect 5789 884 5795 896
rect 5805 784 5811 796
rect 5869 784 5875 916
rect 6541 904 6547 936
rect 6925 903 6931 936
rect 7453 904 7459 916
rect 6916 897 6931 903
rect 5885 884 5891 896
rect 4717 584 4723 596
rect 4909 544 4915 696
rect 4941 584 4947 716
rect 5085 664 5091 676
rect 5101 664 5107 716
rect 5133 704 5139 716
rect 5549 684 5555 696
rect 6013 684 6019 696
rect 5213 664 5219 676
rect 5469 584 5475 676
rect 5629 664 5635 676
rect 5853 584 5859 616
rect 6045 584 6051 716
rect 6093 664 6099 876
rect 6285 784 6291 896
rect 6125 664 6131 676
rect 6093 584 6099 656
rect 5588 537 5596 543
rect 4045 383 4051 476
rect 4036 377 4051 383
rect 3805 317 3820 323
rect 2861 284 2867 316
rect 3501 284 3507 296
rect 2653 264 2659 276
rect 2957 264 2963 276
rect 3309 244 3315 276
rect 1549 204 1555 236
rect 1629 184 1635 236
rect 1853 184 1859 196
rect 1821 144 1827 156
rect 1981 144 1987 236
rect 2045 144 2051 156
rect 1901 124 1907 136
rect 2077 104 2083 236
rect 2381 184 2387 236
rect 2445 204 2451 236
rect 2509 157 2540 163
rect 2173 103 2179 156
rect 2509 144 2515 157
rect 2573 104 2579 236
rect 2733 144 2739 236
rect 3373 224 3379 236
rect 3805 204 3811 317
rect 3709 184 3715 196
rect 3421 157 3436 163
rect 2957 144 2963 156
rect 3181 144 3187 156
rect 3421 144 3427 157
rect 3837 144 3843 336
rect 4365 284 4371 496
rect 4461 444 4467 496
rect 4381 324 4387 436
rect 4477 423 4483 516
rect 4541 504 4547 536
rect 4557 524 4563 536
rect 4941 504 4947 536
rect 4941 444 4947 496
rect 4461 417 4483 423
rect 4461 384 4467 417
rect 4605 324 4611 436
rect 4717 324 4723 336
rect 4941 324 4947 356
rect 4397 243 4403 316
rect 5133 304 5139 536
rect 5149 504 5155 516
rect 5181 504 5187 536
rect 5245 484 5251 496
rect 5613 464 5619 496
rect 5677 484 5683 536
rect 5949 524 5955 536
rect 6157 504 6163 536
rect 6173 524 6179 536
rect 5709 464 5715 496
rect 5549 384 5555 456
rect 5629 324 5635 356
rect 4605 284 4611 296
rect 4941 284 4947 296
rect 5405 284 5411 296
rect 4381 237 4403 243
rect 4189 144 4195 156
rect 2733 104 2739 116
rect 2973 104 2979 136
rect 2164 97 2179 103
rect 2685 -37 2691 16
rect 2653 -43 2691 -37
rect 3597 -43 3603 96
rect 3837 -37 3843 136
rect 4077 104 4083 136
rect 4093 124 4099 136
rect 4180 97 4188 103
rect 3853 84 3859 96
rect 4077 84 4083 96
rect 4077 24 4083 76
rect 3821 -43 3843 -37
rect 4045 -43 4051 16
rect 4381 -43 4387 237
rect 5037 184 5043 276
rect 5389 263 5395 276
rect 5421 263 5427 276
rect 5389 257 5427 263
rect 5469 184 5475 236
rect 5773 184 5779 436
rect 5789 384 5795 496
rect 5869 484 5875 496
rect 6333 444 6339 896
rect 7245 884 7251 896
rect 6493 724 6499 736
rect 6717 724 6723 756
rect 6701 684 6707 696
rect 6765 684 6771 836
rect 7389 764 7395 836
rect 7021 724 7027 736
rect 7373 724 7379 756
rect 7581 724 7587 776
rect 6397 544 6403 556
rect 6573 544 6579 636
rect 6797 584 6803 716
rect 7037 684 7043 696
rect 7364 677 7372 683
rect 6957 624 6963 636
rect 7181 564 7187 636
rect 6973 524 6979 536
rect 7229 524 7235 636
rect 7389 544 7395 636
rect 7581 604 7587 676
rect 7501 544 7507 556
rect 7284 537 7292 543
rect 7645 503 7651 1036
rect 7837 844 7843 1036
rect 8061 984 8067 1116
rect 8077 984 8083 1016
rect 8093 1004 8099 1436
rect 8445 1404 8451 1476
rect 8509 1384 8515 1476
rect 9309 1464 9315 1476
rect 8525 1384 8531 1396
rect 8365 1344 8371 1356
rect 8365 1324 8371 1336
rect 8125 1264 8131 1296
rect 8349 1284 8355 1296
rect 8685 1264 8691 1336
rect 8269 1244 8275 1256
rect 8237 1084 8243 1156
rect 8269 1124 8275 1236
rect 8701 1144 8707 1436
rect 8493 1124 8499 1136
rect 8708 1117 8723 1123
rect 8717 1084 8723 1117
rect 8468 1077 8476 1083
rect 8285 1044 8291 1076
rect 8701 1063 8707 1076
rect 8701 1057 8723 1063
rect 8301 904 8307 956
rect 8349 944 8355 1036
rect 8717 984 8723 1057
rect 8557 944 8563 956
rect 8468 837 8476 843
rect 7661 724 7667 756
rect 8317 724 8323 836
rect 8717 724 8723 836
rect 8692 717 8700 723
rect 8029 684 8035 696
rect 8045 684 8051 696
rect 8477 683 8483 696
rect 8468 677 8483 683
rect 8333 644 8339 676
rect 8244 637 8252 643
rect 7805 584 7811 636
rect 8317 584 8323 596
rect 7741 544 7747 576
rect 8285 544 8291 556
rect 8468 537 8476 543
rect 8301 524 8307 536
rect 7645 497 7660 503
rect 7053 484 7059 496
rect 6637 384 6643 396
rect 5869 284 5875 336
rect 6237 324 6243 336
rect 6285 324 6291 336
rect 6829 284 6835 436
rect 6845 284 6851 316
rect 6077 244 6083 276
rect 7037 244 7043 276
rect 6029 224 6035 236
rect 4852 157 4867 163
rect 4861 143 4867 157
rect 4861 137 4876 143
rect 4413 124 4419 136
rect 4877 124 4883 136
rect 4605 104 4611 116
rect 4404 97 4412 103
rect 4605 -43 4611 96
rect 4685 -37 4691 16
rect 4669 -43 4691 -37
rect 5069 -37 5075 156
rect 5101 144 5107 156
rect 5341 124 5347 136
rect 5101 104 5107 116
rect 5549 104 5555 156
rect 5789 144 5795 156
rect 6445 144 6451 236
rect 6020 137 6028 143
rect 5565 124 5571 136
rect 6029 104 6035 116
rect 6845 104 6851 216
rect 6861 184 6867 236
rect 6909 224 6915 236
rect 7053 144 7059 376
rect 7197 344 7203 436
rect 7197 324 7203 336
rect 7508 317 7523 323
rect 7485 284 7491 296
rect 7517 284 7523 317
rect 7229 144 7235 176
rect 7245 104 7251 236
rect 7357 144 7363 236
rect 7533 144 7539 436
rect 7709 324 7715 336
rect 7949 324 7955 356
rect 8173 324 8179 336
rect 8269 324 8275 336
rect 7709 284 7715 296
rect 7949 284 7955 296
rect 8260 277 8268 283
rect 7853 144 7859 176
rect 8029 144 8035 236
rect 8109 144 8115 236
rect 8429 144 8435 496
rect 8461 324 8467 496
rect 8493 424 8499 636
rect 8701 324 8707 636
rect 8717 544 8723 576
rect 8717 484 8723 496
rect 8733 384 8739 1436
rect 8781 1304 8787 1436
rect 9133 1344 9139 1436
rect 9165 1384 9171 1416
rect 9597 1384 9603 1396
rect 9613 1384 9619 1736
rect 9869 1544 9875 1696
rect 9741 1484 9747 1536
rect 10061 1524 10067 1776
rect 9773 1484 9779 1496
rect 9821 1464 9827 1516
rect 9853 1384 9859 1456
rect 8820 1337 8828 1343
rect 9236 1337 9244 1343
rect 8797 1284 8803 1296
rect 8925 1124 8931 1136
rect 8925 1064 8931 1076
rect 8909 944 8915 956
rect 8957 684 8963 1036
rect 9005 984 9011 1296
rect 9181 1124 9187 1336
rect 9245 1304 9251 1316
rect 9677 1284 9683 1296
rect 10029 1204 10035 1296
rect 10061 1184 10067 1196
rect 9245 1124 9251 1156
rect 9917 1124 9923 1136
rect 9469 1084 9475 1096
rect 9149 1064 9155 1076
rect 9261 1024 9267 1076
rect 9821 1064 9827 1076
rect 9389 1044 9395 1056
rect 9405 984 9411 1056
rect 9421 984 9427 996
rect 9133 944 9139 956
rect 9149 904 9155 956
rect 9165 924 9171 936
rect 9245 904 9251 956
rect 9581 944 9587 956
rect 9597 924 9603 1036
rect 9661 904 9667 1036
rect 9869 904 9875 916
rect 9901 884 9907 936
rect 9645 724 9651 736
rect 9348 717 9363 723
rect 9325 684 9331 716
rect 9357 684 9363 717
rect 9540 717 9548 723
rect 8781 524 8787 636
rect 8813 544 8819 636
rect 9149 604 9155 636
rect 9037 544 9043 596
rect 9165 584 9171 676
rect 9661 664 9667 676
rect 9197 624 9203 636
rect 9373 557 9388 563
rect 9373 544 9379 557
rect 9565 544 9571 576
rect 9805 544 9811 556
rect 9821 544 9827 636
rect 8781 504 8787 516
rect 9357 504 9363 516
rect 8957 444 8963 496
rect 8941 344 8947 436
rect 8925 324 8931 336
rect 9149 324 9155 336
rect 9501 324 9507 336
rect 9732 317 9740 323
rect 8861 264 8867 316
rect 9821 304 9827 316
rect 9837 284 9843 716
rect 9885 684 9891 696
rect 10029 504 10035 636
rect 10045 324 10051 836
rect 10093 724 10099 736
rect 10109 684 10115 896
rect 10189 724 10195 1436
rect 10253 584 10259 1817
rect 10100 537 10108 543
rect 10109 504 10115 516
rect 10269 324 10275 636
rect 8932 277 8940 283
rect 9821 264 9827 276
rect 8493 144 8499 196
rect 8637 164 8643 236
rect 8749 204 8755 236
rect 8781 184 8787 236
rect 8125 124 8131 136
rect 7517 104 7523 116
rect 8077 104 8083 116
rect 8141 104 8147 136
rect 8525 104 8531 156
rect 8589 124 8595 136
rect 8973 124 8979 236
rect 9357 184 9363 236
rect 9533 224 9539 236
rect 9597 184 9603 196
rect 9837 184 9843 216
rect 9156 177 9166 183
rect 9037 144 9043 156
rect 9021 104 9027 136
rect 9197 104 9203 136
rect 9245 104 9251 176
rect 9485 144 9491 156
rect 9677 104 9683 116
rect 10020 97 10028 103
rect 6237 84 6243 96
rect 5149 -37 5155 16
rect 5069 -43 5107 -37
rect 5133 -43 5155 -37
rect 6653 -37 6659 36
rect 7357 -37 7363 16
rect 6653 -43 6675 -37
rect 7341 -43 7363 -37
<< m3contact >>
rect 1772 7596 1780 7604
rect 1820 7596 1828 7604
rect 3580 7616 3588 7624
rect 3612 7616 3620 7624
rect 3356 7536 3364 7544
rect 3388 7536 3396 7544
rect 556 7516 562 7524
rect 562 7516 564 7524
rect 1100 7516 1108 7524
rect 1452 7516 1460 7524
rect 2524 7516 2532 7524
rect 2716 7516 2724 7524
rect 316 7496 324 7504
rect 316 7476 324 7484
rect 524 7476 532 7484
rect 556 7476 564 7484
rect 748 7476 756 7484
rect 76 7456 84 7464
rect 92 7456 100 7464
rect 908 7456 916 7464
rect 2796 7496 2804 7504
rect 1228 7476 1236 7484
rect 1708 7476 1716 7484
rect 2268 7476 2276 7484
rect 2492 7476 2500 7484
rect 2524 7476 2532 7484
rect 3452 7476 3460 7484
rect 1212 7456 1220 7464
rect 1836 7456 1844 7464
rect 2028 7456 2036 7464
rect 1116 7436 1124 7444
rect 2524 7436 2532 7444
rect 284 7416 292 7424
rect 60 7376 68 7384
rect 668 7396 676 7404
rect 508 7376 516 7384
rect 940 7416 948 7424
rect 2236 7376 2244 7384
rect 2956 7456 2964 7464
rect 3036 7456 3044 7464
rect 2732 7436 2740 7444
rect 2716 7396 2724 7404
rect 876 7356 884 7364
rect 1084 7356 1092 7364
rect 1340 7356 1348 7364
rect 1772 7356 1780 7364
rect 2012 7356 2020 7364
rect 2428 7356 2436 7364
rect 300 7336 308 7344
rect 428 7336 436 7344
rect 652 7336 660 7344
rect 764 7336 772 7344
rect 188 7316 196 7324
rect 652 7296 660 7304
rect 1084 7296 1092 7304
rect 268 7276 276 7284
rect 428 7256 436 7264
rect 876 7256 884 7264
rect 268 7136 276 7144
rect 764 7136 772 7144
rect 428 7116 436 7124
rect 652 7076 660 7084
rect 204 7056 212 7064
rect 268 6976 276 6984
rect 204 6956 212 6964
rect 652 6976 660 6984
rect 540 6956 548 6964
rect 668 6956 676 6964
rect 444 6896 452 6904
rect 508 6876 516 6884
rect 76 6816 84 6824
rect 316 6756 324 6764
rect 76 6736 84 6744
rect 524 6696 532 6704
rect 556 6676 564 6684
rect 92 6656 100 6664
rect 268 6616 276 6624
rect 220 6576 228 6584
rect 204 6556 206 6564
rect 206 6556 212 6564
rect 300 6556 308 6564
rect 76 6496 84 6504
rect 412 6476 420 6484
rect 92 6316 100 6324
rect 444 6296 452 6304
rect 92 6256 100 6264
rect 460 6256 468 6264
rect 220 6236 228 6244
rect 236 6216 244 6224
rect 76 6196 84 6204
rect 204 6136 212 6144
rect 668 6596 676 6604
rect 1324 7296 1332 7304
rect 1548 7296 1556 7304
rect 1308 7276 1316 7284
rect 1580 7276 1588 7284
rect 1628 7276 1636 7284
rect 1100 7136 1108 7144
rect 764 7096 772 7104
rect 940 7096 948 7104
rect 1084 7096 1092 7104
rect 1116 7096 1124 7104
rect 1148 7096 1156 7104
rect 956 7036 964 7044
rect 1116 7036 1124 7044
rect 892 6936 900 6944
rect 972 6936 980 6944
rect 1852 7316 1860 7324
rect 1868 7316 1876 7324
rect 1852 7296 1860 7304
rect 1980 7276 1982 7284
rect 1982 7276 1988 7284
rect 2012 7276 2020 7284
rect 2236 7216 2244 7224
rect 1644 7196 1652 7204
rect 2460 7176 2468 7184
rect 3468 7436 3476 7444
rect 3116 7396 3124 7404
rect 3180 7396 3188 7404
rect 2748 7336 2756 7344
rect 3100 7336 3108 7344
rect 3228 7336 3236 7344
rect 3324 7316 3332 7324
rect 3228 7296 3236 7304
rect 2652 7276 2660 7284
rect 3100 7256 3108 7264
rect 3516 7276 3524 7284
rect 3324 7256 3332 7264
rect 3532 7256 3540 7264
rect 1644 7116 1652 7124
rect 2556 7116 2564 7124
rect 2636 7116 2644 7124
rect 2764 7116 2772 7124
rect 2908 7116 2916 7124
rect 1420 7096 1428 7104
rect 1436 7096 1444 7104
rect 3708 7496 3716 7504
rect 5164 7616 5172 7624
rect 6092 7576 6100 7584
rect 4604 7536 4612 7544
rect 6188 7536 6196 7544
rect 9276 7536 9284 7544
rect 3932 7516 3940 7524
rect 4348 7516 4356 7524
rect 3708 7476 3716 7484
rect 3916 7476 3924 7484
rect 4124 7476 4132 7484
rect 3852 7456 3854 7464
rect 3854 7456 3860 7464
rect 3948 7456 3956 7464
rect 3740 7376 3748 7384
rect 4268 7416 4276 7424
rect 5292 7516 5300 7524
rect 6380 7516 6388 7524
rect 6588 7516 6596 7524
rect 7052 7516 7060 7524
rect 7756 7516 7764 7524
rect 8620 7516 8628 7524
rect 8844 7516 8852 7524
rect 9244 7516 9252 7524
rect 4380 7476 4388 7484
rect 5308 7476 5316 7484
rect 5356 7476 5364 7484
rect 4604 7456 4612 7464
rect 4844 7456 4852 7464
rect 4460 7416 4468 7424
rect 5084 7396 5092 7404
rect 5132 7396 5140 7404
rect 5852 7496 5860 7504
rect 5964 7476 5972 7484
rect 5836 7436 5844 7444
rect 5500 7416 5508 7424
rect 5580 7416 5588 7424
rect 5356 7396 5364 7404
rect 3644 7356 3652 7364
rect 3836 7356 3844 7364
rect 4092 7356 4100 7364
rect 4204 7356 4212 7364
rect 4732 7356 4740 7364
rect 5212 7356 5220 7364
rect 5324 7356 5332 7364
rect 4204 7336 4212 7344
rect 4860 7336 4868 7344
rect 3628 7316 3636 7324
rect 4204 7316 4212 7324
rect 4444 7316 4452 7324
rect 4652 7316 4660 7324
rect 4444 7296 4452 7304
rect 4652 7296 4660 7304
rect 4924 7296 4932 7304
rect 3980 7276 3988 7284
rect 3612 7156 3620 7164
rect 5164 7316 5172 7324
rect 6188 7456 6196 7464
rect 6572 7416 6580 7424
rect 6028 7396 6036 7404
rect 5660 7376 5668 7384
rect 5836 7376 5844 7384
rect 5852 7376 5860 7384
rect 6492 7376 6500 7384
rect 6652 7376 6660 7384
rect 6140 7356 6148 7364
rect 6492 7356 6500 7364
rect 5548 7336 5556 7344
rect 5788 7336 5796 7344
rect 5852 7316 5860 7324
rect 6124 7316 6132 7324
rect 6140 7316 6148 7324
rect 5788 7296 5796 7304
rect 5900 7296 5908 7304
rect 6124 7296 6132 7304
rect 6316 7296 6324 7304
rect 6364 7296 6372 7304
rect 6572 7296 6580 7304
rect 4972 7276 4980 7284
rect 5580 7276 5588 7284
rect 5852 7276 5860 7284
rect 6588 7276 6596 7284
rect 4956 7256 4964 7264
rect 4252 7136 4260 7144
rect 4876 7136 4884 7144
rect 3692 7116 3700 7124
rect 3772 7116 3780 7124
rect 4556 7116 4564 7124
rect 4892 7116 4900 7124
rect 4972 7116 4980 7124
rect 5228 7116 5236 7124
rect 2332 7096 2340 7104
rect 3388 7096 3396 7104
rect 3468 7096 3476 7104
rect 1244 7036 1252 7044
rect 1324 6936 1332 6944
rect 876 6916 884 6924
rect 972 6876 980 6884
rect 1180 6876 1188 6884
rect 1324 6836 1332 6844
rect 972 6796 980 6804
rect 1644 7056 1652 7064
rect 1804 7036 1812 7044
rect 1868 7016 1876 7024
rect 2236 7076 2244 7084
rect 2332 7076 2340 7084
rect 2460 7076 2468 7084
rect 3036 7076 3044 7084
rect 3100 7076 3108 7084
rect 2284 6996 2292 7004
rect 2732 7056 2740 7064
rect 2460 6976 2468 6984
rect 2092 6956 2100 6964
rect 1868 6936 1876 6944
rect 2652 6936 2660 6944
rect 1548 6856 1556 6864
rect 1628 6896 1636 6904
rect 1612 6736 1620 6744
rect 1212 6716 1220 6724
rect 1356 6716 1364 6724
rect 1148 6696 1156 6704
rect 764 6676 772 6684
rect 1116 6676 1124 6684
rect 1244 6676 1252 6684
rect 1308 6676 1316 6684
rect 684 6556 692 6564
rect 636 6536 644 6544
rect 876 6516 884 6524
rect 636 6496 644 6504
rect 876 6456 884 6464
rect 1116 6596 1124 6604
rect 1100 6576 1108 6584
rect 972 6556 980 6564
rect 956 6496 964 6504
rect 1548 6636 1556 6644
rect 1388 6616 1396 6624
rect 1436 6616 1444 6624
rect 1324 6556 1332 6564
rect 1308 6516 1316 6524
rect 1292 6476 1300 6484
rect 668 6316 676 6324
rect 892 6316 900 6324
rect 924 6316 932 6324
rect 1372 6516 1380 6524
rect 1516 6516 1524 6524
rect 1532 6516 1540 6524
rect 1340 6316 1348 6324
rect 652 6276 660 6284
rect 524 6256 532 6264
rect 1116 6256 1124 6264
rect 652 6216 660 6224
rect 476 6156 484 6164
rect 476 6136 484 6144
rect 492 6136 500 6144
rect 460 6096 468 6104
rect 204 5876 212 5884
rect 220 5856 228 5864
rect 76 5736 84 5744
rect 188 5736 196 5744
rect 204 5716 212 5724
rect 60 5536 68 5544
rect 220 5536 228 5544
rect 204 5516 212 5524
rect 444 5956 452 5964
rect 300 5756 308 5764
rect 412 5756 420 5764
rect 412 5676 420 5684
rect 268 5516 276 5524
rect 444 5476 452 5484
rect 204 5356 212 5364
rect 252 5356 260 5364
rect 316 5356 324 5364
rect 332 5356 340 5364
rect 300 5336 308 5344
rect 76 5216 84 5224
rect 460 5216 468 5224
rect 444 5136 452 5144
rect 252 5076 260 5084
rect 460 5076 468 5084
rect 92 5056 100 5064
rect 12 4976 20 4984
rect 204 4956 212 4964
rect 252 4976 260 4984
rect 236 4796 244 4804
rect 76 4736 84 4744
rect 444 4736 452 4744
rect 252 4716 260 4724
rect 92 4676 100 4684
rect 444 4676 452 4684
rect 12 4576 20 4584
rect 204 4556 212 4564
rect 236 4556 244 4564
rect 204 4336 212 4344
rect 92 4276 100 4284
rect 220 4276 228 4284
rect 12 4236 20 4244
rect 204 4156 212 4164
rect 236 4156 244 4164
rect 236 4056 244 4064
rect 76 4016 84 4024
rect 220 3876 228 3884
rect 236 3876 244 3884
rect 316 4536 324 4544
rect 524 6096 532 6104
rect 652 6076 660 6084
rect 668 5896 676 5904
rect 1084 6196 1092 6204
rect 1324 6196 1332 6204
rect 940 6176 948 6184
rect 876 6156 884 6164
rect 1164 6176 1172 6184
rect 1292 6156 1300 6164
rect 1084 6116 1092 6124
rect 1308 6116 1316 6124
rect 876 6076 884 6084
rect 1100 6076 1108 6084
rect 1308 6076 1316 6084
rect 732 6036 740 6044
rect 764 5936 772 5944
rect 716 5896 724 5904
rect 780 5896 788 5904
rect 876 5876 884 5884
rect 700 5776 708 5784
rect 492 5716 500 5724
rect 732 5716 740 5724
rect 972 5776 980 5784
rect 1116 5936 1124 5944
rect 1420 6336 1428 6344
rect 2076 6876 2084 6884
rect 2732 6916 2740 6924
rect 2956 6916 2964 6924
rect 2972 6916 2980 6924
rect 2428 6896 2436 6904
rect 2748 6896 2756 6904
rect 2412 6856 2420 6864
rect 2572 6776 2580 6784
rect 1852 6756 1860 6764
rect 1900 6736 1908 6744
rect 2380 6736 2388 6744
rect 2684 6736 2692 6744
rect 2716 6736 2724 6744
rect 1628 6716 1636 6724
rect 1932 6696 1940 6704
rect 2268 6696 2276 6704
rect 2716 6716 2724 6724
rect 2956 6876 2964 6884
rect 2940 6756 2948 6764
rect 2748 6696 2756 6704
rect 1804 6676 1812 6684
rect 2076 6676 2084 6684
rect 2364 6676 2372 6684
rect 3132 6676 3140 6684
rect 1660 6636 1668 6644
rect 1756 6636 1764 6644
rect 1932 6576 1940 6584
rect 2428 6656 2436 6664
rect 2700 6656 2708 6664
rect 2060 6576 2068 6584
rect 1852 6536 1860 6544
rect 2412 6536 2420 6544
rect 2508 6636 2516 6644
rect 2492 6616 2500 6624
rect 2716 6596 2724 6604
rect 2508 6556 2516 6564
rect 2892 6576 2900 6584
rect 2844 6556 2852 6564
rect 2620 6536 2628 6544
rect 2796 6536 2804 6544
rect 3084 6536 3092 6544
rect 1628 6496 1636 6504
rect 1852 6496 1860 6504
rect 2076 6496 2084 6504
rect 2428 6496 2436 6504
rect 1532 6316 1540 6324
rect 1436 6256 1444 6264
rect 2860 6476 2868 6484
rect 2636 6456 2644 6464
rect 2236 6416 2244 6424
rect 3692 7056 3700 7064
rect 3868 7056 3876 7064
rect 4012 7056 4020 7064
rect 3980 7036 3988 7044
rect 3340 6996 3348 7004
rect 3308 6936 3316 6944
rect 3308 6876 3316 6884
rect 3164 6856 3172 6864
rect 3532 6856 3540 6864
rect 3164 6716 3172 6724
rect 3244 6736 3252 6744
rect 3884 7016 3892 7024
rect 4540 7096 4548 7104
rect 4316 7076 4324 7084
rect 4476 7076 4484 7084
rect 4092 7056 4100 7064
rect 4204 6956 4212 6964
rect 4460 7056 4468 7064
rect 4412 6976 4420 6984
rect 4444 6976 4452 6984
rect 4076 6916 4084 6924
rect 3756 6896 3764 6904
rect 3788 6896 3796 6904
rect 3980 6896 3988 6904
rect 4028 6896 4036 6904
rect 4076 6896 4082 6904
rect 4082 6896 4084 6904
rect 4236 6936 4244 6944
rect 4316 6936 4324 6944
rect 4220 6876 4228 6884
rect 3772 6856 3780 6864
rect 4188 6836 4196 6844
rect 4044 6736 4052 6744
rect 4268 6816 4276 6824
rect 4268 6756 4276 6764
rect 4988 7096 4996 7104
rect 4876 7076 4884 7084
rect 5132 7076 5140 7084
rect 5244 7076 5252 7084
rect 4748 7036 4756 7044
rect 4556 6956 4564 6964
rect 4604 6956 4612 6964
rect 4540 6936 4548 6944
rect 4620 6916 4628 6924
rect 4412 6736 4420 6744
rect 3468 6716 3476 6724
rect 3596 6716 3604 6724
rect 3820 6716 3828 6724
rect 4236 6716 4244 6724
rect 4060 6696 4068 6704
rect 6012 7116 6020 7124
rect 6124 7116 6132 7124
rect 5452 7076 5460 7084
rect 6012 7076 6020 7084
rect 5372 7056 5380 7064
rect 4828 6936 4836 6944
rect 4988 6936 4996 6944
rect 5068 6936 5076 6944
rect 5420 6936 5428 6944
rect 5196 6916 5204 6924
rect 5180 6896 5188 6904
rect 4876 6876 4884 6884
rect 4700 6816 4708 6824
rect 4940 6816 4948 6824
rect 5036 6756 5044 6764
rect 6124 7056 6132 7064
rect 5900 7036 5908 7044
rect 5788 6996 5796 7004
rect 6012 6996 6020 7004
rect 5900 6936 5908 6944
rect 5980 6936 5988 6944
rect 6220 6936 6228 6944
rect 6572 7136 6580 7144
rect 6332 7096 6340 7104
rect 6588 7096 6596 7104
rect 6860 7476 6868 7484
rect 7036 7436 7044 7444
rect 7436 7476 7444 7484
rect 7100 7456 7108 7464
rect 7068 7396 7076 7404
rect 7180 7376 7188 7384
rect 7244 7376 7252 7384
rect 7548 7496 7556 7504
rect 7468 7416 7476 7424
rect 7532 7376 7540 7384
rect 8204 7496 8212 7504
rect 8412 7496 8420 7504
rect 8460 7476 8468 7484
rect 8732 7476 8740 7484
rect 8204 7456 8212 7464
rect 9484 7496 9492 7504
rect 9708 7496 9716 7504
rect 9916 7496 9924 7504
rect 8860 7476 8868 7484
rect 9180 7476 9188 7484
rect 9948 7476 9956 7484
rect 9292 7456 9300 7464
rect 9500 7456 9508 7464
rect 9708 7456 9716 7464
rect 8764 7436 8772 7444
rect 10060 7436 10068 7444
rect 7980 7396 7988 7404
rect 8300 7396 8308 7404
rect 7788 7376 7796 7384
rect 7820 7376 7828 7384
rect 7836 7376 7844 7384
rect 8060 7376 8068 7384
rect 8140 7376 8148 7384
rect 7708 7336 7716 7344
rect 7772 7336 7780 7344
rect 7468 7316 7476 7324
rect 8044 7356 8052 7364
rect 8268 7356 8276 7364
rect 8348 7356 8356 7364
rect 8732 7396 8740 7404
rect 8492 7316 8500 7324
rect 8572 7316 8580 7324
rect 8588 7316 8596 7324
rect 6812 7296 6820 7304
rect 8060 7296 8068 7304
rect 8492 7296 8494 7304
rect 8494 7296 8500 7304
rect 6940 7116 6948 7124
rect 6780 7056 6788 7064
rect 6956 7056 6964 7064
rect 6780 7036 6788 7044
rect 6796 7016 6804 7024
rect 6924 6996 6932 7004
rect 6780 6956 6788 6964
rect 6284 6936 6292 6944
rect 6668 6936 6676 6944
rect 6268 6916 6276 6924
rect 5996 6896 6004 6904
rect 6204 6896 6212 6904
rect 6956 6896 6964 6904
rect 6316 6876 6324 6884
rect 6684 6876 6692 6884
rect 6300 6856 6308 6864
rect 6364 6856 6372 6864
rect 5596 6816 5604 6824
rect 5772 6756 5780 6764
rect 5260 6736 5268 6744
rect 5404 6736 5412 6744
rect 7468 7276 7476 7284
rect 7372 7256 7380 7264
rect 8268 7256 8276 7264
rect 7180 7216 7188 7224
rect 7388 7136 7396 7144
rect 7164 7116 7172 7124
rect 7484 7116 7492 7124
rect 7612 7116 7620 7124
rect 7164 7096 7172 7104
rect 7244 7076 7252 7084
rect 8092 7176 8100 7184
rect 8172 7156 8180 7164
rect 8412 7156 8420 7164
rect 7708 7116 7716 7124
rect 7948 7116 7956 7124
rect 7948 7096 7956 7104
rect 8172 7096 8180 7104
rect 8396 7096 8404 7104
rect 7868 7056 7876 7064
rect 7468 6956 7476 6964
rect 7676 6956 7684 6964
rect 7244 6936 7252 6944
rect 7468 6936 7476 6944
rect 7004 6916 7012 6924
rect 7404 6896 7412 6904
rect 7564 6896 7572 6904
rect 7772 6896 7780 6904
rect 6988 6876 6996 6884
rect 6988 6836 6996 6844
rect 7964 6956 7972 6964
rect 8556 6976 8564 6984
rect 8828 7256 8836 7264
rect 8636 7136 8644 7144
rect 9036 7416 9044 7424
rect 9260 7376 9268 7384
rect 9052 7316 9060 7324
rect 9036 7296 9044 7304
rect 9580 7356 9588 7364
rect 9612 7296 9620 7304
rect 9420 7216 9428 7224
rect 9436 7216 9444 7224
rect 8876 7116 8884 7124
rect 8972 7116 8980 7124
rect 8988 7116 8996 7124
rect 9052 7116 9060 7124
rect 9212 7116 9220 7124
rect 8604 7096 8612 7104
rect 8636 7096 8644 7104
rect 9436 7096 9444 7104
rect 8636 7076 8644 7084
rect 8892 7076 8900 7084
rect 8940 7076 8948 7084
rect 9436 7076 9444 7084
rect 8012 6936 8020 6944
rect 8108 6936 8116 6944
rect 8588 6936 8596 6944
rect 8796 6936 8804 6944
rect 8860 6916 8868 6924
rect 8012 6896 8020 6904
rect 8108 6896 8116 6904
rect 8668 6856 8676 6864
rect 8508 6836 8516 6844
rect 8268 6816 8276 6824
rect 4508 6716 4516 6724
rect 4684 6716 4692 6724
rect 4748 6716 4756 6724
rect 5084 6716 5092 6724
rect 3452 6676 3460 6684
rect 3484 6676 3492 6684
rect 4060 6676 4068 6684
rect 4268 6676 4276 6684
rect 4476 6676 4484 6684
rect 3676 6636 3684 6644
rect 4060 6636 4068 6644
rect 4348 6616 4356 6624
rect 4044 6596 4052 6604
rect 4252 6596 4260 6604
rect 3612 6576 3620 6584
rect 3628 6576 3636 6584
rect 3820 6576 3828 6584
rect 4588 6696 4596 6704
rect 5036 6676 5044 6684
rect 5276 6676 5284 6684
rect 4588 6656 4596 6664
rect 5324 6636 5332 6644
rect 4716 6556 4724 6564
rect 4828 6556 4836 6564
rect 3244 6536 3252 6544
rect 3420 6536 3428 6544
rect 3580 6536 3588 6544
rect 3740 6536 3748 6544
rect 3180 6516 3188 6524
rect 3148 6396 3156 6404
rect 3116 6356 3124 6364
rect 1628 6316 1636 6324
rect 2492 6316 2500 6324
rect 2780 6316 2788 6324
rect 2940 6316 2948 6324
rect 3228 6316 3236 6324
rect 3548 6316 3556 6324
rect 2236 6296 2244 6304
rect 1660 6256 1668 6264
rect 1884 6256 1892 6264
rect 2044 6256 2052 6264
rect 1564 6236 1572 6244
rect 1612 6236 1620 6244
rect 1996 6216 2004 6224
rect 1548 6196 1556 6204
rect 1836 6176 1844 6184
rect 1596 6136 1604 6144
rect 1740 6136 1748 6144
rect 1772 6136 1780 6144
rect 1404 6096 1412 6104
rect 1628 6096 1636 6104
rect 1340 5876 1348 5884
rect 1116 5776 1124 5784
rect 1004 5696 1012 5704
rect 940 5656 948 5664
rect 924 5616 932 5624
rect 988 5536 996 5544
rect 668 5496 676 5504
rect 684 5496 692 5504
rect 988 5496 996 5504
rect 924 5476 932 5484
rect 908 5456 916 5464
rect 700 5436 708 5444
rect 1388 5856 1396 5864
rect 1532 6056 1540 6064
rect 1980 6096 1988 6104
rect 1964 6076 1972 6084
rect 2460 6296 2468 6304
rect 2476 6256 2484 6264
rect 2332 6216 2340 6224
rect 2252 6196 2260 6204
rect 2444 6196 2452 6204
rect 2204 6156 2212 6164
rect 2796 6296 2804 6304
rect 2764 6276 2772 6284
rect 2924 6276 2932 6284
rect 3020 6276 3028 6284
rect 3564 6276 3572 6284
rect 2700 6256 2708 6264
rect 3452 6256 3458 6264
rect 3458 6256 3460 6264
rect 2508 6236 2516 6244
rect 2860 6236 2868 6244
rect 2684 6196 2692 6204
rect 2716 6196 2724 6204
rect 2844 6136 2852 6144
rect 2076 6096 2084 6104
rect 2300 6096 2308 6104
rect 2012 6016 2020 6024
rect 1804 5896 1812 5904
rect 2028 5896 2036 5904
rect 1804 5856 1812 5864
rect 1884 5756 1892 5764
rect 1420 5736 1428 5744
rect 1628 5736 1636 5744
rect 1660 5736 1668 5744
rect 1084 5716 1092 5724
rect 1196 5716 1204 5724
rect 1372 5716 1380 5724
rect 1900 5696 1908 5704
rect 1804 5676 1812 5684
rect 1884 5676 1892 5684
rect 1116 5656 1124 5664
rect 1420 5656 1428 5664
rect 1644 5656 1652 5664
rect 1676 5556 1682 5564
rect 1682 5556 1684 5564
rect 1068 5536 1076 5544
rect 1580 5516 1588 5524
rect 1148 5476 1156 5484
rect 1340 5476 1348 5484
rect 1004 5456 1012 5464
rect 1148 5416 1156 5424
rect 524 5356 532 5364
rect 1148 5356 1156 5364
rect 1356 5356 1364 5364
rect 908 5336 916 5344
rect 1132 5336 1140 5344
rect 1436 5336 1444 5344
rect 1580 5336 1588 5344
rect 668 5316 676 5324
rect 1580 5316 1588 5324
rect 1372 5296 1380 5304
rect 908 5276 916 5284
rect 1228 5276 1236 5284
rect 1580 5276 1588 5284
rect 508 5256 516 5264
rect 1564 5256 1572 5264
rect 1228 5216 1236 5224
rect 892 5156 900 5164
rect 668 5136 676 5144
rect 492 5116 500 5124
rect 956 5116 964 5124
rect 1212 5116 1220 5124
rect 1564 5116 1572 5124
rect 988 5096 996 5104
rect 652 5076 660 5084
rect 1228 5076 1236 5084
rect 1340 5076 1348 5084
rect 1372 5076 1380 5084
rect 524 5056 532 5064
rect 892 5056 900 5064
rect 508 5036 516 5044
rect 684 5036 692 5044
rect 972 4976 980 4984
rect 908 4956 916 4964
rect 1116 4956 1124 4964
rect 668 4896 676 4904
rect 1116 4896 1124 4904
rect 1516 5036 1524 5044
rect 1516 4956 1524 4964
rect 1564 4956 1572 4964
rect 1228 4936 1236 4944
rect 1372 4936 1380 4944
rect 1516 4936 1524 4944
rect 1196 4916 1204 4924
rect 1132 4876 1140 4884
rect 2044 5516 2052 5524
rect 1836 5496 1844 5504
rect 2028 5496 2036 5504
rect 2204 6076 2212 6084
rect 3420 6176 3426 6184
rect 3426 6176 3428 6184
rect 3964 6516 3972 6524
rect 4172 6496 4180 6504
rect 3964 6456 3972 6464
rect 4380 6536 4388 6544
rect 4476 6536 4484 6544
rect 4396 6496 4404 6504
rect 3820 6336 3828 6344
rect 4044 6336 4052 6344
rect 4188 6336 4196 6344
rect 4316 6336 4324 6344
rect 3772 6316 3780 6324
rect 3564 6136 3572 6144
rect 2892 6096 2900 6104
rect 2988 6096 2996 6104
rect 3308 6096 3316 6104
rect 3548 6096 3556 6104
rect 2492 6076 2500 6084
rect 2204 6056 2212 6064
rect 2316 6056 2324 6064
rect 2508 5936 2516 5944
rect 2268 5896 2276 5904
rect 2508 5896 2516 5904
rect 2924 6056 2932 6064
rect 2908 5956 2916 5964
rect 2732 5916 2740 5924
rect 2700 5896 2708 5904
rect 2940 5956 2948 5964
rect 2284 5856 2292 5864
rect 2492 5856 2500 5864
rect 2524 5856 2532 5864
rect 2284 5836 2292 5844
rect 2332 5816 2340 5824
rect 2268 5796 2276 5804
rect 2348 5756 2356 5764
rect 2524 5736 2532 5744
rect 2124 5696 2132 5704
rect 2348 5696 2356 5704
rect 2556 5696 2564 5704
rect 2140 5516 2148 5524
rect 2492 5496 2500 5504
rect 1836 5476 1844 5484
rect 1788 5416 1796 5424
rect 1612 5396 1620 5404
rect 1852 5376 1860 5384
rect 2060 5376 2068 5384
rect 1804 5356 1812 5364
rect 1836 5356 1844 5364
rect 2028 5356 2036 5364
rect 1644 5296 1652 5304
rect 1836 5116 1844 5124
rect 1676 5056 1684 5064
rect 1884 5096 1892 5104
rect 2012 5076 2020 5084
rect 1820 4956 1828 4964
rect 1900 4956 1908 4964
rect 1596 4916 1604 4924
rect 1676 4916 1684 4924
rect 2060 4916 2068 4924
rect 1564 4896 1572 4904
rect 1660 4896 1668 4904
rect 1900 4896 1908 4904
rect 1404 4856 1412 4864
rect 1548 4736 1556 4744
rect 1788 4736 1796 4744
rect 1884 4736 1892 4744
rect 524 4716 532 4724
rect 924 4716 932 4724
rect 940 4716 948 4724
rect 1212 4716 1220 4724
rect 668 4676 676 4684
rect 700 4676 708 4684
rect 1132 4676 1140 4684
rect 684 4596 692 4604
rect 524 4556 532 4564
rect 556 4536 564 4544
rect 300 4496 308 4504
rect 684 4496 692 4504
rect 284 4336 292 4344
rect 316 4136 324 4144
rect 316 4096 324 4104
rect 428 3896 436 3904
rect 252 3836 260 3844
rect 236 3816 244 3824
rect 12 3776 20 3784
rect 252 3796 260 3804
rect 284 3756 292 3764
rect 444 3756 452 3764
rect 60 3656 68 3664
rect 204 3656 212 3664
rect 444 3516 452 3524
rect 60 3496 68 3504
rect 204 3476 212 3484
rect 236 3476 244 3484
rect 220 3456 228 3464
rect 444 3456 452 3464
rect 300 3416 308 3424
rect 204 3316 212 3324
rect 220 3296 228 3304
rect 444 3296 452 3304
rect 284 3116 292 3124
rect 188 2996 196 3004
rect 60 2956 68 2964
rect 92 2956 100 2964
rect 284 2956 292 2964
rect 76 2936 84 2944
rect 300 2936 308 2944
rect 428 2936 436 2944
rect 428 2896 436 2904
rect 268 2836 276 2844
rect 444 2676 452 2684
rect 204 2656 212 2664
rect 236 2656 244 2664
rect 252 2616 260 2624
rect 92 2536 100 2544
rect 444 2536 452 2544
rect 444 2496 452 2504
rect 204 2476 212 2484
rect 460 2396 468 2404
rect 236 2336 244 2344
rect 300 2156 308 2164
rect 92 2136 100 2144
rect 316 2136 324 2144
rect 220 2016 228 2024
rect 204 1896 212 1904
rect 284 1916 292 1924
rect 300 1856 308 1864
rect 252 1816 260 1824
rect 428 1816 436 1824
rect 60 1756 68 1764
rect 92 1756 100 1764
rect 444 1756 452 1764
rect 76 1736 84 1744
rect 444 1656 452 1664
rect 204 1556 212 1564
rect 284 1556 292 1564
rect 428 1536 436 1544
rect 220 1516 228 1524
rect 428 1456 436 1464
rect 60 1336 68 1344
rect 92 1336 100 1344
rect 316 1336 324 1344
rect 108 1296 116 1304
rect 300 1296 308 1304
rect 76 1196 84 1204
rect 236 1116 244 1124
rect 444 1116 452 1124
rect 220 1096 228 1104
rect 204 1076 212 1084
rect 236 1076 244 1084
rect 492 4456 500 4464
rect 556 4316 562 4324
rect 562 4316 564 4324
rect 556 4276 564 4284
rect 668 4256 676 4264
rect 524 4076 532 4084
rect 652 3856 660 3864
rect 668 3856 676 3864
rect 908 4656 916 4664
rect 1148 4656 1156 4664
rect 924 4636 932 4644
rect 1180 4636 1188 4644
rect 908 4556 916 4564
rect 988 4536 996 4544
rect 1132 4536 1140 4544
rect 1564 4716 1572 4724
rect 2012 4716 2020 4724
rect 2044 4716 2052 4724
rect 1916 4676 1924 4684
rect 1596 4656 1604 4664
rect 1788 4656 1796 4664
rect 1900 4656 1908 4664
rect 1420 4636 1428 4644
rect 1372 4596 1380 4604
rect 1404 4596 1412 4604
rect 1836 4596 1844 4604
rect 1916 4596 1924 4604
rect 1340 4576 1348 4584
rect 1372 4576 1380 4584
rect 1612 4556 1620 4564
rect 1612 4536 1620 4544
rect 1692 4536 1700 4544
rect 1932 4536 1940 4544
rect 2220 5436 2228 5444
rect 2220 5336 2228 5344
rect 2268 5336 2276 5344
rect 2300 5316 2308 5324
rect 2508 5376 2516 5384
rect 2540 5376 2548 5384
rect 2380 5336 2388 5344
rect 2268 5276 2276 5284
rect 2348 5256 2356 5264
rect 2124 5136 2132 5144
rect 2476 5116 2484 5124
rect 2124 5096 2132 5104
rect 2780 5796 2788 5804
rect 2716 5776 2724 5784
rect 2748 5756 2756 5764
rect 2908 5756 2916 5764
rect 3100 6076 3108 6084
rect 3564 6076 3572 6084
rect 4492 6496 4500 6504
rect 4492 6336 4500 6344
rect 4236 6276 4244 6284
rect 3804 6256 3812 6264
rect 4044 6256 4052 6264
rect 4476 6256 4484 6264
rect 4332 6236 4340 6244
rect 3596 6116 3604 6124
rect 3580 6016 3588 6024
rect 3756 6156 3764 6164
rect 3772 6096 3780 6104
rect 3612 5956 3620 5964
rect 2988 5936 2996 5944
rect 3596 5936 3604 5944
rect 3356 5916 3364 5924
rect 2956 5736 2964 5744
rect 2780 5676 2788 5684
rect 2572 5656 2580 5664
rect 2572 5636 2580 5644
rect 2700 5636 2708 5644
rect 2748 5536 2756 5544
rect 2748 5416 2756 5424
rect 2748 5336 2756 5344
rect 2732 5276 2740 5284
rect 2716 5156 2724 5164
rect 2508 5076 2516 5084
rect 2476 5056 2484 5064
rect 2108 4816 2116 4824
rect 2252 4636 2260 4644
rect 2476 4916 2484 4924
rect 2476 4716 2484 4724
rect 2460 4676 2468 4684
rect 2524 4716 2532 4724
rect 2524 4656 2532 4664
rect 2268 4616 2276 4624
rect 2284 4616 2292 4624
rect 2508 4616 2516 4624
rect 2300 4596 2308 4604
rect 2108 4576 2116 4584
rect 2284 4576 2292 4584
rect 2460 4576 2468 4584
rect 1244 4516 1252 4524
rect 1436 4516 1444 4524
rect 2076 4516 2084 4524
rect 1244 4476 1252 4484
rect 748 4456 756 4464
rect 1164 4396 1172 4404
rect 908 4336 916 4344
rect 1900 4496 1908 4504
rect 2460 4536 2468 4544
rect 2492 4536 2500 4544
rect 2460 4476 2468 4484
rect 1596 4456 1604 4464
rect 1692 4456 1700 4464
rect 2252 4456 2260 4464
rect 2044 4436 2052 4444
rect 940 4316 948 4324
rect 1004 4316 1012 4324
rect 1356 4316 1364 4324
rect 892 4276 900 4284
rect 780 4236 788 4244
rect 924 4216 932 4224
rect 1436 4296 1444 4304
rect 1644 4376 1652 4384
rect 2268 4316 2276 4324
rect 2332 4316 2340 4324
rect 2460 4316 2468 4324
rect 1004 4276 1012 4284
rect 1788 4276 1796 4284
rect 1820 4276 1828 4284
rect 2268 4276 2276 4284
rect 2012 4256 2020 4264
rect 1580 4216 1588 4224
rect 1820 4216 1828 4224
rect 1612 4196 1620 4204
rect 1596 4176 1604 4184
rect 1196 4156 1204 4164
rect 1228 4156 1236 4164
rect 1804 4156 1812 4164
rect 1836 4156 1844 4164
rect 764 4136 772 4144
rect 1116 4136 1124 4144
rect 1388 4136 1396 4144
rect 2028 4136 2036 4144
rect 764 4116 772 4124
rect 1820 4116 1828 4124
rect 2476 4276 2484 4284
rect 2492 4216 2500 4224
rect 2524 4216 2532 4224
rect 2092 4176 2100 4184
rect 2460 4156 2468 4164
rect 1116 4096 1124 4104
rect 1228 4096 1236 4104
rect 1420 4096 1428 4104
rect 1580 4096 1588 4104
rect 2476 4096 2484 4104
rect 2236 4076 2244 4084
rect 2668 5076 2676 5084
rect 2668 4976 2676 4984
rect 2588 4916 2596 4924
rect 2764 4916 2772 4924
rect 2940 5516 2948 5524
rect 2844 5336 2852 5344
rect 2972 5336 2980 5344
rect 2828 5316 2836 5324
rect 2956 5116 2964 5124
rect 2796 5076 2804 5084
rect 2940 4996 2948 5004
rect 2796 4956 2804 4964
rect 3356 5896 3364 5904
rect 3804 5896 3812 5904
rect 3180 5876 3188 5884
rect 3580 5876 3588 5884
rect 3788 5876 3796 5884
rect 3020 5856 3028 5864
rect 3148 5796 3156 5804
rect 3020 5756 3028 5764
rect 3180 5716 3188 5724
rect 3004 5656 3012 5664
rect 3164 5536 3172 5544
rect 3180 5496 3188 5504
rect 3148 5456 3156 5464
rect 3004 5396 3012 5404
rect 3180 5316 3188 5324
rect 3020 5296 3028 5304
rect 3196 5276 3204 5284
rect 3436 5796 3444 5804
rect 3388 5776 3396 5784
rect 3452 5776 3458 5784
rect 3458 5776 3460 5784
rect 3372 5716 3380 5724
rect 3580 5756 3588 5764
rect 3660 5796 3668 5804
rect 3644 5716 3652 5724
rect 3788 5716 3796 5724
rect 3596 5696 3604 5704
rect 3484 5656 3492 5664
rect 3644 5656 3652 5664
rect 3228 5576 3236 5584
rect 3388 5556 3396 5564
rect 3468 5536 3476 5544
rect 4124 6216 4132 6224
rect 4012 6176 4020 6184
rect 4220 6176 4228 6184
rect 3852 6136 3860 6144
rect 3996 6116 4004 6124
rect 4316 6136 4324 6144
rect 4300 6096 4308 6104
rect 4892 6496 4900 6504
rect 5180 6616 5188 6624
rect 5276 6536 5284 6544
rect 5820 6696 5828 6704
rect 6172 6736 6180 6744
rect 6732 6736 6740 6744
rect 6972 6736 6980 6744
rect 7500 6736 7508 6744
rect 6844 6716 6852 6724
rect 7308 6716 7316 6724
rect 7708 6716 7716 6724
rect 5868 6696 5876 6704
rect 5532 6676 5540 6684
rect 5628 6676 5636 6684
rect 6076 6676 6084 6684
rect 5436 6636 5444 6644
rect 5404 6596 5412 6604
rect 5564 6656 5572 6664
rect 5612 6656 5620 6664
rect 5836 6656 5844 6664
rect 5788 6636 5796 6644
rect 5628 6596 5636 6604
rect 5692 6556 5700 6564
rect 5420 6536 5428 6544
rect 5564 6536 5572 6544
rect 4524 6356 4532 6364
rect 4508 6296 4516 6304
rect 4908 6356 4916 6364
rect 4636 6336 4644 6344
rect 4684 6296 4692 6304
rect 4684 6276 4692 6284
rect 5532 6496 5540 6504
rect 5756 6496 5764 6504
rect 5084 6476 5092 6484
rect 4988 6336 4996 6344
rect 5212 6336 5220 6344
rect 5372 6336 5380 6344
rect 5532 6336 5540 6344
rect 4908 6256 4916 6264
rect 4940 6256 4948 6264
rect 4700 6176 4708 6184
rect 4572 6156 4580 6164
rect 4508 6096 4516 6104
rect 4556 6096 4564 6104
rect 4268 6076 4276 6084
rect 4492 6076 4500 6084
rect 4092 6036 4100 6044
rect 4028 5896 4036 5904
rect 4252 5896 4260 5904
rect 4252 5876 4260 5884
rect 3884 5716 3892 5724
rect 3884 5676 3892 5684
rect 4108 5736 4116 5744
rect 4236 5736 4244 5744
rect 3900 5636 3908 5644
rect 4092 5636 4100 5644
rect 3836 5616 3844 5624
rect 3804 5596 3812 5604
rect 3916 5556 3924 5564
rect 3916 5496 3924 5504
rect 4908 6196 4916 6204
rect 4972 6196 4980 6204
rect 5820 6316 5828 6324
rect 5452 6296 5460 6304
rect 5484 6296 5492 6304
rect 5180 6256 5188 6264
rect 5372 6256 5380 6264
rect 5804 6256 5812 6264
rect 5804 6236 5812 6244
rect 5372 6196 5380 6204
rect 5212 6176 5220 6184
rect 5660 6156 5668 6164
rect 4796 6136 4804 6144
rect 5228 6136 5236 6144
rect 5436 6136 5444 6144
rect 4748 6096 4756 6104
rect 5004 6096 5012 6104
rect 5820 6156 5828 6164
rect 5676 6116 5684 6124
rect 5404 6096 5412 6104
rect 5004 6056 5012 6064
rect 5244 6056 5252 6064
rect 5580 6076 5588 6084
rect 5628 6056 5636 6064
rect 5404 6036 5412 6044
rect 5628 6036 5636 6044
rect 5260 5996 5268 6004
rect 5036 5936 5044 5944
rect 5420 5936 5428 5944
rect 4940 5916 4948 5924
rect 4988 5916 4996 5924
rect 4476 5876 4484 5884
rect 4732 5876 4740 5884
rect 4700 5856 4708 5864
rect 4284 5836 4292 5844
rect 4492 5816 4500 5824
rect 4716 5796 4724 5804
rect 5388 5876 5396 5884
rect 5388 5856 5396 5864
rect 4924 5776 4932 5784
rect 4908 5756 4916 5764
rect 4364 5736 4372 5744
rect 4796 5736 4804 5744
rect 5244 5736 5252 5744
rect 4332 5676 4340 5684
rect 4348 5676 4356 5684
rect 4332 5656 4340 5664
rect 4572 5716 4580 5724
rect 5164 5716 5172 5724
rect 4572 5696 4580 5704
rect 5132 5696 5140 5704
rect 5388 5696 5396 5704
rect 4780 5676 4788 5684
rect 4924 5616 4932 5624
rect 4492 5556 4500 5564
rect 4828 5556 4836 5564
rect 4364 5516 4372 5524
rect 4508 5516 4516 5524
rect 4588 5516 4596 5524
rect 4812 5516 4820 5524
rect 4268 5496 4276 5504
rect 4588 5496 4596 5504
rect 5180 5536 5188 5544
rect 5404 5536 5412 5544
rect 5500 5916 5508 5924
rect 5500 5856 5508 5864
rect 6332 6696 6340 6704
rect 6172 6656 6180 6664
rect 6284 6656 6292 6664
rect 6620 6656 6628 6664
rect 6092 6616 6100 6624
rect 6268 6556 6276 6564
rect 5884 6536 5892 6544
rect 6108 6536 6116 6544
rect 5868 6516 5876 6524
rect 5884 6516 5892 6524
rect 6076 6496 6084 6504
rect 6092 6496 6100 6504
rect 6012 6336 6020 6344
rect 5900 6316 5908 6324
rect 6828 6636 6836 6644
rect 6476 6596 6484 6604
rect 6764 6596 6772 6604
rect 6748 6576 6756 6584
rect 7292 6656 7300 6664
rect 7068 6636 7076 6644
rect 7036 6596 7044 6604
rect 7180 6596 7188 6604
rect 7164 6576 7172 6584
rect 6908 6536 6916 6544
rect 7020 6536 7028 6544
rect 7132 6536 7140 6544
rect 6572 6516 6580 6524
rect 6332 6496 6340 6504
rect 6572 6496 6580 6504
rect 7164 6476 7172 6484
rect 6364 6356 6372 6364
rect 6252 6336 6260 6344
rect 6588 6336 6596 6344
rect 6748 6336 6756 6344
rect 6124 6296 6132 6304
rect 6604 6276 6612 6284
rect 6076 6256 6084 6264
rect 6140 6256 6148 6264
rect 6252 6256 6260 6264
rect 6364 6256 6372 6264
rect 5916 6236 5924 6244
rect 5996 6156 6004 6164
rect 6028 6156 6036 6164
rect 6012 6096 6020 6104
rect 5836 6076 5844 6084
rect 6236 6136 6244 6144
rect 6332 6156 6340 6164
rect 6156 6096 6164 6104
rect 6252 6096 6260 6104
rect 6044 5956 6052 5964
rect 5724 5936 5732 5944
rect 6076 5916 6084 5924
rect 5724 5896 5732 5904
rect 6076 5896 6084 5904
rect 6332 6056 6340 6064
rect 6812 6336 6820 6344
rect 7036 6316 7044 6324
rect 7356 6556 7364 6564
rect 7660 6656 7668 6664
rect 7724 6656 7732 6664
rect 7516 6596 7524 6604
rect 7836 6596 7844 6604
rect 7676 6576 7684 6584
rect 7852 6556 7860 6564
rect 7596 6536 7604 6544
rect 7804 6536 7812 6544
rect 8588 6716 8596 6724
rect 8908 6716 8916 6724
rect 7932 6676 7940 6684
rect 8092 6676 8100 6684
rect 8572 6676 8580 6684
rect 7916 6656 7924 6664
rect 8460 6656 8468 6664
rect 8060 6616 8068 6624
rect 8780 6596 8788 6604
rect 8908 6576 8916 6584
rect 8044 6536 8052 6544
rect 8092 6536 8100 6544
rect 8220 6536 8228 6544
rect 7356 6496 7364 6504
rect 7436 6496 7444 6504
rect 7596 6476 7604 6484
rect 7868 6476 7876 6484
rect 7500 6436 7508 6444
rect 7276 6296 7284 6304
rect 7004 6276 7012 6284
rect 7052 6276 7060 6284
rect 7212 6276 7220 6284
rect 6780 6256 6788 6264
rect 7340 6236 7348 6244
rect 7244 6216 7252 6224
rect 7180 6176 7188 6184
rect 6924 6156 6932 6164
rect 8252 6536 8260 6544
rect 8252 6496 8260 6504
rect 8364 6496 8372 6504
rect 8460 6496 8468 6504
rect 8556 6496 8564 6504
rect 8764 6496 8772 6504
rect 8252 6476 8260 6484
rect 8252 6336 8260 6344
rect 8028 6316 8036 6324
rect 8316 6316 8324 6324
rect 7804 6276 7812 6284
rect 7452 6216 7460 6224
rect 7404 6176 7412 6184
rect 6556 6136 6564 6144
rect 7148 6136 7156 6144
rect 7340 6136 7348 6144
rect 7420 6136 7428 6144
rect 8012 6276 8020 6284
rect 8428 6276 8436 6284
rect 8060 6256 8068 6264
rect 8012 6236 8020 6244
rect 8076 6236 8084 6244
rect 7852 6216 7860 6224
rect 7676 6176 7684 6184
rect 8476 6356 8484 6364
rect 8572 6356 8580 6364
rect 8684 6276 8692 6284
rect 8540 6236 8548 6244
rect 8556 6236 8564 6244
rect 8108 6156 8116 6164
rect 7884 6136 7892 6144
rect 6572 6116 6580 6124
rect 7148 6116 7156 6124
rect 7580 6116 7588 6124
rect 7644 6116 7652 6124
rect 7676 6116 7684 6124
rect 8332 6116 8340 6124
rect 8716 6236 8724 6244
rect 8556 6136 8564 6144
rect 7212 6096 7220 6104
rect 6924 6076 6932 6084
rect 8012 6076 8020 6084
rect 8108 6056 8116 6064
rect 6780 6036 6788 6044
rect 6796 6036 6804 6044
rect 6524 6016 6532 6024
rect 6476 5936 6484 5944
rect 8332 5956 8340 5964
rect 7820 5936 7828 5944
rect 7852 5936 7860 5944
rect 7948 5936 7956 5944
rect 6316 5916 6324 5924
rect 6556 5916 6564 5924
rect 6540 5896 6548 5904
rect 6316 5876 6324 5884
rect 6748 5876 6756 5884
rect 6844 5876 6852 5884
rect 6156 5856 6164 5864
rect 6332 5856 6340 5864
rect 5884 5836 5892 5844
rect 5692 5756 5700 5764
rect 5468 5716 5476 5724
rect 5692 5656 5700 5664
rect 5404 5516 5412 5524
rect 5180 5496 5188 5504
rect 5388 5496 5396 5504
rect 3820 5476 3828 5484
rect 5500 5476 5508 5484
rect 5724 5476 5732 5484
rect 5836 5476 5844 5484
rect 3484 5456 3492 5464
rect 3804 5456 3812 5464
rect 3676 5436 3684 5444
rect 3404 5416 3412 5424
rect 3612 5416 3620 5424
rect 3900 5376 3908 5384
rect 4060 5376 4068 5384
rect 3436 5356 3444 5364
rect 3628 5336 3636 5344
rect 4108 5336 4116 5344
rect 3420 5316 3428 5324
rect 3868 5316 3876 5324
rect 3948 5316 3956 5324
rect 3404 5296 3412 5304
rect 4108 5296 4116 5304
rect 3276 5236 3284 5244
rect 3692 5236 3700 5244
rect 3180 5156 3188 5164
rect 3148 5096 3156 5104
rect 2988 4936 2996 4944
rect 3020 4896 3028 4904
rect 2796 4876 2804 4884
rect 3036 4736 3044 4744
rect 3420 5196 3428 5204
rect 3644 5196 3652 5204
rect 3212 5136 3220 5144
rect 2716 4716 2724 4724
rect 2796 4696 2804 4704
rect 2828 4676 2836 4684
rect 2700 4656 2708 4664
rect 2572 4556 2580 4564
rect 2956 4656 2964 4664
rect 3148 4656 3156 4664
rect 3180 4656 3188 4664
rect 2940 4556 2948 4564
rect 3148 4556 3156 4564
rect 2812 4536 2820 4544
rect 2956 4536 2964 4544
rect 2764 4476 2772 4484
rect 2796 4476 2804 4484
rect 3004 4456 3012 4464
rect 3164 4456 3172 4464
rect 3196 4596 3204 4604
rect 3196 4376 3204 4384
rect 2796 4336 2804 4344
rect 2556 4296 2564 4304
rect 2700 4296 2708 4304
rect 3148 4296 3156 4304
rect 2716 4276 2724 4284
rect 2700 4256 2708 4264
rect 3004 4256 3012 4264
rect 3164 4256 3172 4264
rect 2956 4236 2964 4244
rect 2716 4196 2724 4204
rect 2956 4176 2964 4184
rect 2700 4156 2708 4164
rect 3132 4156 3140 4164
rect 2924 4136 2932 4144
rect 3148 4116 3156 4124
rect 2540 4076 2548 4084
rect 2652 4076 2660 4084
rect 2700 4076 2708 4084
rect 2476 4056 2484 4064
rect 1772 3956 1780 3964
rect 1196 3936 1204 3944
rect 2236 3936 2244 3944
rect 1100 3916 1108 3924
rect 2732 3936 2740 3944
rect 732 3836 740 3844
rect 1420 3896 1428 3904
rect 1612 3896 1620 3904
rect 1868 3896 1876 3904
rect 2460 3896 2468 3904
rect 1116 3876 1124 3884
rect 1212 3876 1220 3884
rect 1884 3876 1892 3884
rect 2908 3916 2916 3924
rect 3020 3876 3028 3884
rect 1772 3856 1780 3864
rect 2476 3856 2484 3864
rect 1148 3776 1156 3784
rect 1852 3776 1860 3784
rect 1676 3756 1682 3764
rect 1682 3756 1684 3764
rect 668 3736 676 3744
rect 732 3736 740 3744
rect 1340 3736 1348 3744
rect 908 3696 916 3704
rect 668 3516 676 3524
rect 540 3456 548 3464
rect 668 3336 676 3344
rect 892 3496 900 3504
rect 956 3696 964 3704
rect 1116 3676 1124 3684
rect 2092 3816 2100 3824
rect 2044 3796 2052 3804
rect 2012 3756 2020 3764
rect 2268 3756 2276 3764
rect 2012 3736 2020 3744
rect 2252 3736 2260 3744
rect 2028 3716 2036 3724
rect 2476 3716 2484 3724
rect 1580 3696 1588 3704
rect 1132 3656 1140 3664
rect 2252 3656 2260 3664
rect 1836 3576 1844 3584
rect 1116 3556 1124 3564
rect 956 3496 964 3504
rect 1340 3536 1348 3544
rect 1196 3496 1204 3504
rect 1340 3496 1348 3504
rect 956 3476 964 3484
rect 940 3456 948 3464
rect 1132 3456 1140 3464
rect 1180 3456 1188 3464
rect 1660 3496 1668 3504
rect 1452 3456 1460 3464
rect 1644 3456 1652 3464
rect 1804 3456 1812 3464
rect 2492 3516 2500 3524
rect 2028 3496 2036 3504
rect 2092 3476 2100 3484
rect 2252 3476 2260 3484
rect 2284 3476 2292 3484
rect 2444 3476 2452 3484
rect 2012 3456 2020 3464
rect 2044 3436 2052 3444
rect 2012 3376 2020 3384
rect 1244 3356 1252 3364
rect 908 3336 916 3344
rect 972 3336 980 3344
rect 1004 3336 1012 3344
rect 1580 3336 1588 3344
rect 1004 3316 1012 3324
rect 1708 3316 1716 3324
rect 1932 3316 1940 3324
rect 1436 3296 1444 3304
rect 1692 3296 1700 3304
rect 1916 3296 1924 3304
rect 1596 3276 1604 3284
rect 1164 3256 1172 3264
rect 1244 3256 1252 3264
rect 940 3156 948 3164
rect 508 3136 516 3144
rect 876 3136 884 3144
rect 1100 3116 1108 3124
rect 1084 3076 1092 3084
rect 524 3056 532 3064
rect 716 3056 724 3064
rect 508 2996 516 3004
rect 636 2956 644 2964
rect 1596 3196 1604 3204
rect 1532 3136 1540 3144
rect 1196 3116 1204 3124
rect 1372 3116 1380 3124
rect 1532 3096 1540 3104
rect 1196 3056 1204 3064
rect 1388 3056 1396 3064
rect 1324 2996 1332 3004
rect 732 2936 740 2944
rect 732 2896 740 2904
rect 652 2876 660 2884
rect 700 2836 708 2844
rect 700 2676 708 2684
rect 668 2656 676 2664
rect 700 2596 708 2604
rect 940 2756 948 2764
rect 908 2676 916 2684
rect 1180 2796 1188 2804
rect 1308 2916 1316 2924
rect 1852 3116 1860 3124
rect 2076 3116 2084 3124
rect 2268 3436 2276 3444
rect 2268 3396 2276 3404
rect 2124 3376 2132 3384
rect 2140 3356 2148 3364
rect 2380 3356 2388 3364
rect 2236 3276 2244 3284
rect 2380 3276 2388 3284
rect 1644 3056 1652 3064
rect 2044 3056 2052 3064
rect 2092 3056 2100 3064
rect 2220 3036 2228 3044
rect 1612 2996 1620 3004
rect 1788 2996 1796 3004
rect 2540 3796 2548 3804
rect 2716 3856 2724 3864
rect 2908 3856 2916 3864
rect 2956 3856 2964 3864
rect 2748 3816 2756 3824
rect 2668 3736 2676 3744
rect 2588 3716 2596 3724
rect 2588 3696 2596 3704
rect 2780 3696 2788 3704
rect 2940 3696 2948 3704
rect 2556 3596 2564 3604
rect 3132 3856 3140 3864
rect 3180 3736 3188 3744
rect 3180 3676 3188 3684
rect 2684 3476 2692 3484
rect 2924 3476 2932 3484
rect 2572 3416 2580 3424
rect 3164 3476 3172 3484
rect 3180 3416 3188 3424
rect 2732 3376 2740 3384
rect 2556 3356 2564 3364
rect 2780 3356 2788 3364
rect 2796 3356 2804 3364
rect 2972 3356 2980 3364
rect 3196 3356 3204 3364
rect 3164 3296 3172 3304
rect 3244 5076 3252 5084
rect 3260 5056 3268 5064
rect 3564 5176 3572 5184
rect 3596 5076 3604 5084
rect 3452 5056 3460 5064
rect 3468 5016 3476 5024
rect 4124 5196 4132 5204
rect 3932 5156 3940 5164
rect 3948 5076 3956 5084
rect 3724 5056 3732 5064
rect 4092 5036 4100 5044
rect 3852 5016 3860 5024
rect 3868 5016 3876 5024
rect 3260 4956 3268 4964
rect 3484 4956 3492 4964
rect 3644 4956 3652 4964
rect 3260 4916 3268 4924
rect 3932 4976 3940 4984
rect 4076 4956 4084 4964
rect 4076 4896 4084 4904
rect 4220 5356 4228 5364
rect 5260 5456 5266 5464
rect 5266 5456 5268 5464
rect 5276 5456 5284 5464
rect 5708 5456 5716 5464
rect 4364 5356 4372 5364
rect 4204 5336 4212 5344
rect 4252 5336 4260 5344
rect 4748 5336 4756 5344
rect 4796 5316 4804 5324
rect 4860 5316 4868 5324
rect 4412 5296 4420 5304
rect 4572 5296 4580 5304
rect 5004 5296 5012 5304
rect 4796 5276 4804 5284
rect 4300 5116 4308 5124
rect 4300 5096 4308 5104
rect 4172 5076 4180 5084
rect 4396 5076 4404 5084
rect 4572 5076 4580 5084
rect 4412 5056 4420 5064
rect 4364 4996 4372 5004
rect 4524 4956 4532 4964
rect 4172 4936 4180 4944
rect 4172 4896 4180 4904
rect 4140 4876 4148 4884
rect 4524 4876 4532 4884
rect 3228 4856 3236 4864
rect 3500 4856 3508 4864
rect 3836 4856 3844 4864
rect 4348 4856 4356 4864
rect 4492 4856 4500 4864
rect 4140 4836 4148 4844
rect 3596 4736 3604 4744
rect 3820 4716 3828 4724
rect 4492 4716 4500 4724
rect 3596 4696 3604 4704
rect 3404 4676 3412 4684
rect 3580 4656 3588 4664
rect 3468 4636 3476 4644
rect 3388 4536 3396 4544
rect 3868 4636 3876 4644
rect 3804 4556 3812 4564
rect 3612 4516 3620 4524
rect 3644 4516 3652 4524
rect 3836 4516 3844 4524
rect 3868 4516 3876 4524
rect 3388 4496 3396 4504
rect 3612 4336 3620 4344
rect 3372 4316 3380 4324
rect 3612 4316 3620 4324
rect 3404 4256 3412 4264
rect 3580 4256 3588 4264
rect 3228 4236 3236 4244
rect 3420 4236 3428 4244
rect 3420 4196 3428 4204
rect 3868 4496 3876 4504
rect 4268 4676 4276 4684
rect 4300 4676 4308 4684
rect 4476 4656 4484 4664
rect 4300 4616 4308 4624
rect 3916 4576 3924 4584
rect 4060 4576 4068 4584
rect 4140 4576 4148 4584
rect 4268 4576 4276 4584
rect 4300 4576 4308 4584
rect 4508 4536 4516 4544
rect 4060 4496 4068 4504
rect 3884 4376 3892 4384
rect 3660 4356 3668 4364
rect 4012 4336 4020 4344
rect 3820 4316 3828 4324
rect 3804 4296 3812 4304
rect 3788 4236 3796 4244
rect 3660 4216 3668 4224
rect 4268 4516 4276 4524
rect 4828 4976 4836 4984
rect 4604 4956 4612 4964
rect 4956 4936 4964 4944
rect 4956 4896 4964 4904
rect 4604 4876 4612 4884
rect 4572 4856 4580 4864
rect 4556 4736 4564 4744
rect 5100 5396 5108 5404
rect 5228 5316 5236 5324
rect 5244 5276 5252 5284
rect 5196 5136 5204 5144
rect 5580 5436 5588 5444
rect 5500 5396 5508 5404
rect 5356 5376 5364 5384
rect 5580 5336 5588 5344
rect 5836 5336 5844 5344
rect 5932 5816 5940 5824
rect 6492 5756 6500 5764
rect 5932 5736 5940 5744
rect 5916 5716 5924 5724
rect 6492 5716 6500 5724
rect 5900 5696 5908 5704
rect 6108 5696 6116 5704
rect 6492 5696 6500 5704
rect 6060 5536 6068 5544
rect 6060 5476 6068 5484
rect 5884 5376 5892 5384
rect 5340 5296 5348 5304
rect 5484 5296 5492 5304
rect 5708 5296 5716 5304
rect 5916 5296 5924 5304
rect 5692 5256 5700 5264
rect 5628 5156 5636 5164
rect 5452 5116 5460 5124
rect 5308 5076 5316 5084
rect 5196 5056 5204 5064
rect 5180 4936 5188 4944
rect 5180 4916 5188 4924
rect 5260 4816 5268 4824
rect 4540 4716 4548 4724
rect 4572 4716 4580 4724
rect 4236 4496 4244 4504
rect 4316 4316 4324 4324
rect 4524 4316 4532 4324
rect 4236 4296 4244 4304
rect 4940 4736 4948 4744
rect 5036 4736 5044 4744
rect 5260 4736 5268 4744
rect 4924 4676 4932 4684
rect 4956 4676 4964 4684
rect 5276 4696 5284 4704
rect 5164 4656 5172 4664
rect 4572 4616 4580 4624
rect 4220 4276 4228 4284
rect 4540 4276 4548 4284
rect 3996 4256 4004 4264
rect 4076 4256 4084 4264
rect 4684 4256 4692 4264
rect 4732 4636 4740 4644
rect 5244 4596 5252 4604
rect 4828 4556 4836 4564
rect 4732 4536 4740 4544
rect 5340 4536 5348 4544
rect 5036 4496 5044 4504
rect 5308 4496 5316 4504
rect 4924 4336 4932 4344
rect 5372 4476 5380 4484
rect 5388 4356 5396 4364
rect 5500 5096 5508 5104
rect 6076 5396 6084 5404
rect 6332 5456 6340 5464
rect 6364 5536 6372 5544
rect 6524 5536 6532 5544
rect 6348 5416 6356 5424
rect 6236 5376 6244 5384
rect 6300 5376 6308 5384
rect 6012 5356 6020 5364
rect 6124 5356 6132 5364
rect 6124 5336 6132 5344
rect 6380 5336 6388 5344
rect 7020 5896 7028 5904
rect 7308 5876 7316 5884
rect 7084 5856 7092 5864
rect 6860 5816 6868 5824
rect 6972 5816 6980 5824
rect 6812 5776 6820 5784
rect 8156 5896 8164 5904
rect 7692 5856 7700 5864
rect 7420 5816 7428 5824
rect 7516 5816 7524 5824
rect 7740 5816 7748 5824
rect 7932 5816 7940 5824
rect 7180 5776 7188 5784
rect 7740 5756 7748 5764
rect 6604 5736 6612 5744
rect 6828 5736 6836 5744
rect 7500 5736 7508 5744
rect 7916 5736 7924 5744
rect 8060 5736 8068 5744
rect 8140 5736 8148 5744
rect 7276 5716 7284 5724
rect 6828 5696 6836 5704
rect 7020 5696 7028 5704
rect 7276 5696 7284 5704
rect 7484 5696 7492 5704
rect 6588 5676 6596 5684
rect 6812 5536 6820 5544
rect 8092 5676 8100 5684
rect 7724 5656 7732 5664
rect 7404 5556 7412 5564
rect 7708 5556 7716 5564
rect 8092 5556 8100 5564
rect 7020 5536 7028 5544
rect 7500 5536 7508 5544
rect 7052 5496 7060 5504
rect 7724 5496 7732 5504
rect 7932 5496 7940 5504
rect 7948 5496 7956 5504
rect 6620 5476 6628 5484
rect 6732 5476 6740 5484
rect 6844 5476 6852 5484
rect 7004 5476 7012 5484
rect 7020 5476 7028 5484
rect 7324 5476 7332 5484
rect 7500 5476 7508 5484
rect 6716 5456 6724 5464
rect 6620 5396 6628 5404
rect 7260 5436 7268 5444
rect 7196 5416 7204 5424
rect 6572 5376 6580 5384
rect 6876 5376 6884 5384
rect 7148 5376 7156 5384
rect 6716 5356 6724 5364
rect 6140 5316 6148 5324
rect 6380 5316 6388 5324
rect 6476 5316 6484 5324
rect 6476 5296 6484 5304
rect 6284 5276 6292 5284
rect 5948 5216 5956 5224
rect 5932 5156 5940 5164
rect 6332 5256 6340 5264
rect 7068 5336 7076 5344
rect 6700 5316 6708 5324
rect 6716 5316 6724 5324
rect 7388 5456 7396 5464
rect 7692 5456 7700 5464
rect 7852 5416 7860 5424
rect 8316 5776 8324 5784
rect 9708 7336 9716 7344
rect 9692 7256 9700 7264
rect 9628 7116 9636 7124
rect 9628 7056 9636 7064
rect 9132 7016 9140 7024
rect 9468 7016 9476 7024
rect 9068 6976 9076 6984
rect 9452 6956 9460 6964
rect 10268 7376 10276 7384
rect 9916 7316 9924 7324
rect 9932 7296 9940 7304
rect 9868 7136 9876 7144
rect 9868 7116 9876 7124
rect 9852 7096 9860 7104
rect 9692 7036 9700 7044
rect 9644 6996 9652 7004
rect 9644 6956 9652 6964
rect 9884 6956 9892 6964
rect 9100 6936 9108 6944
rect 9516 6936 9524 6944
rect 9676 6936 9684 6944
rect 9372 6896 9380 6904
rect 9116 6876 9124 6884
rect 9340 6876 9348 6884
rect 9436 6876 9444 6884
rect 9660 6876 9668 6884
rect 10236 6996 10244 7004
rect 10108 6916 10116 6924
rect 9564 6736 9572 6744
rect 9356 6716 9364 6724
rect 9660 6716 9668 6724
rect 9868 6716 9876 6724
rect 10252 6716 10260 6724
rect 9004 6696 9012 6704
rect 9900 6696 9908 6704
rect 9196 6676 9204 6684
rect 9340 6676 9348 6684
rect 9836 6676 9844 6684
rect 9020 6656 9028 6664
rect 9388 6636 9396 6644
rect 9116 6536 9124 6544
rect 9180 6536 9188 6544
rect 9132 6516 9140 6524
rect 8988 6376 8996 6384
rect 9148 6336 9156 6344
rect 8908 6296 8916 6304
rect 9020 6276 9028 6284
rect 9164 6276 9172 6284
rect 8908 6256 8916 6264
rect 8764 6236 8772 6244
rect 9164 6216 9172 6224
rect 9676 6656 9684 6664
rect 9564 6616 9572 6624
rect 9804 6616 9812 6624
rect 9564 6556 9572 6564
rect 9836 6556 9844 6564
rect 9676 6516 9684 6524
rect 9612 6496 9620 6504
rect 9436 6436 9444 6444
rect 9356 6316 9364 6324
rect 9356 6276 9364 6284
rect 8988 6136 8996 6144
rect 9212 6136 9220 6144
rect 9340 6136 9348 6144
rect 8892 6116 8900 6124
rect 8892 6096 8900 6104
rect 9004 6096 9012 6104
rect 9180 6076 9188 6084
rect 9340 6076 9348 6084
rect 8988 5996 8996 6004
rect 9420 6356 9428 6364
rect 9820 6456 9828 6464
rect 9788 6356 9796 6364
rect 9468 6276 9476 6284
rect 9596 6276 9604 6284
rect 9532 6156 9540 6164
rect 9260 5976 9268 5984
rect 9388 5976 9396 5984
rect 9036 5936 9044 5944
rect 9820 6256 9828 6264
rect 9820 6236 9828 6244
rect 9788 6216 9796 6224
rect 9644 6196 9652 6204
rect 10012 6516 10020 6524
rect 10044 6496 10052 6504
rect 10012 6476 10020 6484
rect 9868 6356 9876 6364
rect 10124 6556 10132 6564
rect 10220 6316 10222 6324
rect 10222 6316 10228 6324
rect 10220 6296 10228 6304
rect 10076 6276 10084 6284
rect 10028 6196 10036 6204
rect 10012 6176 10020 6184
rect 10044 6176 10052 6184
rect 10076 6136 10084 6144
rect 10204 6136 10212 6144
rect 9804 6056 9812 6064
rect 8524 5916 8532 5924
rect 8572 5916 8580 5924
rect 8604 5916 8612 5924
rect 8700 5916 8708 5924
rect 8732 5916 8740 5924
rect 9580 5916 9588 5924
rect 9596 5916 9604 5924
rect 9692 5916 9700 5924
rect 8508 5856 8516 5864
rect 8364 5796 8372 5804
rect 8492 5796 8500 5804
rect 8796 5896 8804 5904
rect 8956 5876 8964 5884
rect 8604 5856 8612 5864
rect 8508 5676 8516 5684
rect 8812 5776 8820 5784
rect 8956 5616 8964 5624
rect 8700 5556 8708 5564
rect 8492 5536 8500 5544
rect 8732 5536 8740 5544
rect 8172 5516 8180 5524
rect 8300 5516 8308 5524
rect 8956 5496 8964 5504
rect 8172 5456 8180 5464
rect 8956 5476 8964 5484
rect 8604 5456 8612 5464
rect 8764 5456 8772 5464
rect 8412 5416 8420 5424
rect 8060 5396 8068 5404
rect 8140 5396 8148 5404
rect 8460 5396 8468 5404
rect 7372 5376 7380 5384
rect 7180 5356 7188 5364
rect 7516 5356 7524 5364
rect 8284 5356 8292 5364
rect 8412 5336 8420 5344
rect 8892 5396 8900 5404
rect 8940 5396 8948 5404
rect 8748 5376 8756 5384
rect 8732 5356 8740 5364
rect 7628 5316 7636 5324
rect 7868 5316 7876 5324
rect 7532 5296 7540 5304
rect 7148 5276 7156 5284
rect 7628 5276 7636 5284
rect 8044 5276 8052 5284
rect 7068 5256 7076 5264
rect 7772 5236 7780 5244
rect 6524 5216 6532 5224
rect 6556 5136 6564 5144
rect 7212 5176 7220 5184
rect 7708 5216 7716 5224
rect 8204 5276 8212 5284
rect 8428 5256 8436 5264
rect 8188 5176 8196 5184
rect 7964 5156 7972 5164
rect 7868 5136 7876 5144
rect 5724 5116 5732 5124
rect 6188 5116 6196 5124
rect 6284 5116 6292 5124
rect 6908 5116 6916 5124
rect 7004 5116 7012 5124
rect 7308 5116 7316 5124
rect 7436 5116 7444 5124
rect 8204 5116 8212 5124
rect 8556 5336 8564 5344
rect 8652 5336 8660 5344
rect 9260 5896 9268 5904
rect 9244 5876 9252 5884
rect 9484 5876 9492 5884
rect 9580 5876 9588 5884
rect 9676 5876 9684 5884
rect 9004 5656 9012 5664
rect 9164 5856 9172 5864
rect 9180 5776 9188 5784
rect 9372 5716 9380 5724
rect 9372 5696 9380 5704
rect 9692 5856 9700 5864
rect 9580 5796 9588 5804
rect 9836 5776 9844 5784
rect 9484 5736 9492 5744
rect 9724 5736 9732 5744
rect 9884 6116 9892 6124
rect 9868 6096 9876 6104
rect 9884 6076 9892 6084
rect 9868 6056 9876 6064
rect 9900 5876 9908 5884
rect 10044 5816 10052 5824
rect 10044 5796 10052 5804
rect 9852 5716 9860 5724
rect 9884 5716 9892 5724
rect 9900 5716 9908 5724
rect 9452 5696 9460 5704
rect 9692 5696 9700 5704
rect 9692 5676 9700 5684
rect 10220 5676 10228 5684
rect 9420 5616 9428 5624
rect 9836 5536 9844 5544
rect 9404 5516 9412 5524
rect 9628 5516 9636 5524
rect 9020 5396 9028 5404
rect 9388 5476 9396 5484
rect 9196 5416 9204 5424
rect 9324 5396 9332 5404
rect 9196 5356 9204 5364
rect 10028 5496 10036 5504
rect 9852 5476 9860 5484
rect 10044 5396 10052 5404
rect 9644 5376 9652 5384
rect 9820 5376 9828 5384
rect 9468 5356 9476 5364
rect 9644 5356 9652 5364
rect 9868 5356 9876 5364
rect 10028 5356 10036 5364
rect 10044 5356 10052 5364
rect 10236 5356 10244 5364
rect 8988 5336 8996 5344
rect 9036 5336 9044 5344
rect 9084 5336 9092 5344
rect 9420 5336 9428 5344
rect 9772 5336 9780 5344
rect 8652 5296 8654 5304
rect 8654 5296 8660 5304
rect 8540 5256 8548 5264
rect 8524 5196 8532 5204
rect 9548 5316 9556 5324
rect 9548 5296 9556 5304
rect 9868 5296 9876 5304
rect 9180 5276 9188 5284
rect 9772 5276 9780 5284
rect 9068 5196 9076 5204
rect 9052 5156 9060 5164
rect 5852 5096 5860 5104
rect 5868 5096 5876 5104
rect 5884 5096 5892 5104
rect 6652 5096 6660 5104
rect 6188 5076 6196 5084
rect 6652 5076 6660 5084
rect 6844 5076 6852 5084
rect 6540 5056 6548 5064
rect 7004 5056 7012 5064
rect 7212 5056 7220 5064
rect 7356 5056 7364 5064
rect 6860 5036 6868 5044
rect 7132 5036 7140 5044
rect 5660 4996 5668 5004
rect 5596 4976 5604 4984
rect 5628 4976 5636 4984
rect 5836 4996 5844 5004
rect 6796 5016 6804 5024
rect 7068 5016 7076 5024
rect 6540 4996 6548 5004
rect 6396 4976 6404 4984
rect 6780 4976 6788 4984
rect 5692 4956 5700 4964
rect 5724 4956 5732 4964
rect 6108 4956 6116 4964
rect 6348 4936 6356 4944
rect 5596 4896 5604 4904
rect 5900 4896 5908 4904
rect 5692 4876 5700 4884
rect 6684 4916 6692 4924
rect 7228 4936 7236 4944
rect 7292 4936 7300 4944
rect 6972 4916 6980 4924
rect 6348 4896 6356 4904
rect 6508 4896 6516 4904
rect 6700 4896 6708 4904
rect 6332 4876 6340 4884
rect 6988 4876 6996 4884
rect 6508 4836 6516 4844
rect 6508 4736 6516 4744
rect 6588 4736 6596 4744
rect 5500 4716 5508 4724
rect 5500 4676 5508 4684
rect 5468 4636 5476 4644
rect 5596 4536 5604 4544
rect 5612 4456 5620 4464
rect 5452 4356 5460 4364
rect 5948 4716 5954 4724
rect 5954 4716 5956 4724
rect 6492 4716 6500 4724
rect 6956 4716 6964 4724
rect 5932 4676 5940 4684
rect 5964 4676 5972 4684
rect 6124 4676 6132 4684
rect 6604 4676 6612 4684
rect 5724 4656 5732 4664
rect 6284 4616 6292 4624
rect 6316 4616 6324 4624
rect 5948 4556 5956 4564
rect 6156 4556 6164 4564
rect 5836 4536 5844 4544
rect 6604 4536 6612 4544
rect 5916 4516 5924 4524
rect 6156 4516 6164 4524
rect 6332 4516 6340 4524
rect 6476 4516 6484 4524
rect 6588 4496 6596 4504
rect 6140 4476 6148 4484
rect 6492 4476 6500 4484
rect 6748 4476 6756 4484
rect 5836 4456 5844 4464
rect 6140 4456 6148 4464
rect 5644 4336 5652 4344
rect 6156 4336 6164 4344
rect 6620 4336 6628 4344
rect 7164 4896 7172 4904
rect 7500 5036 7508 5044
rect 7980 5096 7988 5104
rect 8748 5116 8756 5124
rect 8828 5116 8836 5124
rect 9036 5096 9044 5104
rect 8844 5076 8852 5084
rect 7868 5056 7876 5064
rect 7596 5036 7604 5044
rect 7516 4996 7524 5004
rect 7436 4916 7444 4924
rect 7452 4896 7460 4904
rect 7404 4876 7412 4884
rect 7580 4876 7588 4884
rect 7260 4736 7268 4744
rect 7612 4996 7620 5004
rect 7884 4956 7892 4964
rect 8076 4956 8084 4964
rect 8428 5056 8436 5064
rect 8460 5056 8468 5064
rect 8748 5056 8756 5064
rect 8972 5056 8980 5064
rect 8204 4976 8212 4984
rect 8220 4976 8228 4984
rect 7740 4936 7748 4944
rect 7788 4936 7796 4944
rect 7868 4936 7876 4944
rect 8124 4936 8132 4944
rect 8204 4936 8212 4944
rect 8348 4956 8356 4964
rect 8476 4976 8484 4984
rect 8764 4976 8772 4984
rect 8588 4956 8596 4964
rect 9692 5136 9700 5144
rect 10092 5296 10100 5304
rect 9484 5116 9492 5124
rect 9148 5076 9156 5084
rect 9388 5076 9396 5084
rect 9612 5076 9620 5084
rect 9708 5076 9716 5084
rect 9884 5076 9892 5084
rect 10028 5076 10036 5084
rect 9500 5056 9508 5064
rect 9148 4976 9156 4984
rect 9244 4956 9252 4964
rect 10172 4996 10180 5004
rect 8396 4936 8404 4944
rect 8428 4936 8436 4944
rect 8668 4936 8676 4944
rect 9036 4936 9044 4944
rect 9164 4936 9172 4944
rect 9404 4936 9412 4944
rect 9564 4936 9572 4944
rect 9596 4936 9604 4944
rect 9820 4936 9828 4944
rect 9900 4936 9908 4944
rect 8300 4916 8308 4924
rect 7644 4896 7652 4904
rect 7852 4736 7860 4744
rect 7372 4716 7380 4724
rect 7676 4716 7684 4724
rect 7036 4696 7044 4704
rect 7692 4696 7700 4704
rect 7260 4676 7268 4684
rect 7276 4596 7284 4604
rect 7388 4596 7396 4604
rect 7708 4636 7716 4644
rect 7836 4636 7844 4644
rect 7580 4596 7588 4604
rect 8668 4896 8676 4904
rect 8732 4756 8740 4764
rect 8252 4716 8260 4724
rect 8476 4716 8484 4724
rect 8556 4716 8564 4724
rect 8492 4696 8500 4704
rect 8252 4656 8260 4664
rect 8588 4656 8596 4664
rect 8284 4636 8292 4644
rect 8044 4596 8052 4604
rect 8572 4596 8580 4604
rect 8284 4576 8292 4584
rect 8780 4876 8788 4884
rect 9180 4916 9188 4924
rect 9388 4896 9396 4904
rect 10012 4896 10020 4904
rect 9612 4876 9620 4884
rect 8972 4776 8980 4784
rect 9148 4736 9156 4744
rect 9692 4756 9700 4764
rect 9580 4736 9588 4744
rect 10092 4736 10100 4744
rect 9340 4716 9348 4724
rect 8796 4696 8804 4704
rect 9692 4696 9700 4704
rect 9132 4676 9140 4684
rect 9228 4676 9236 4684
rect 9388 4676 9396 4684
rect 9580 4676 9588 4684
rect 9676 4676 9684 4684
rect 10252 4676 10260 4684
rect 9212 4656 9220 4664
rect 9916 4656 9924 4664
rect 8748 4636 8756 4644
rect 8892 4636 8900 4644
rect 8940 4636 8948 4644
rect 10204 4636 10212 4644
rect 8716 4576 8724 4584
rect 8316 4556 8324 4564
rect 8444 4556 8452 4564
rect 8572 4556 8580 4564
rect 8716 4556 8724 4564
rect 8028 4536 8036 4544
rect 6828 4516 6836 4524
rect 7148 4496 7156 4504
rect 6828 4456 6836 4464
rect 7052 4456 7060 4464
rect 6796 4356 6804 4364
rect 7036 4356 7044 4364
rect 4716 4316 4724 4324
rect 5100 4316 5108 4324
rect 5436 4316 5444 4324
rect 5612 4316 5620 4324
rect 6380 4316 6388 4324
rect 4860 4296 4868 4304
rect 5068 4296 5076 4304
rect 5212 4276 5220 4284
rect 4316 4236 4324 4244
rect 4540 4236 4548 4244
rect 4700 4236 4708 4244
rect 4780 4236 4788 4244
rect 3612 4136 3620 4144
rect 3852 4116 3860 4124
rect 3452 4096 3460 4104
rect 3596 4096 3604 4104
rect 3388 4056 3396 4064
rect 3452 4036 3460 4044
rect 3372 3936 3380 3944
rect 3612 3896 3620 3904
rect 3260 3876 3268 3884
rect 3372 3876 3380 3884
rect 3596 3876 3604 3884
rect 3644 3816 3652 3824
rect 3420 3776 3428 3784
rect 3836 4076 3844 4084
rect 3820 3896 3828 3904
rect 4060 4136 4068 4144
rect 4076 3976 4084 3984
rect 3932 3916 3940 3924
rect 3868 3896 3876 3904
rect 3948 3776 3956 3784
rect 3708 3756 3716 3764
rect 4044 3756 4052 3764
rect 3420 3736 3428 3744
rect 3628 3736 3636 3744
rect 3660 3736 3668 3744
rect 3404 3716 3412 3724
rect 4028 3696 4036 3704
rect 4060 3696 4068 3704
rect 4076 3696 4084 3704
rect 3692 3676 3700 3684
rect 3916 3676 3924 3684
rect 3724 3616 3732 3624
rect 3372 3516 3380 3524
rect 3804 3516 3812 3524
rect 3596 3496 3604 3504
rect 3372 3476 3380 3484
rect 3580 3456 3588 3464
rect 3628 3456 3636 3464
rect 3228 3436 3236 3444
rect 3596 3436 3604 3444
rect 4012 3436 4020 3444
rect 3452 3396 3460 3404
rect 3228 3296 3236 3304
rect 3404 3296 3412 3304
rect 2812 3276 2820 3284
rect 3212 3276 3220 3284
rect 3404 3256 3412 3264
rect 2524 3216 2532 3224
rect 2284 3156 2292 3164
rect 2492 3156 2500 3164
rect 3084 3136 3092 3144
rect 3644 3376 3652 3384
rect 3836 3356 3844 3364
rect 4364 4136 4372 4144
rect 4476 4136 4484 4144
rect 4668 4136 4676 4144
rect 4108 3736 4116 3744
rect 4140 4096 4148 4104
rect 4524 4116 4532 4124
rect 4732 4096 4740 4104
rect 4172 4056 4180 4064
rect 4332 4056 4340 4064
rect 4588 4056 4596 4064
rect 4380 3936 4388 3944
rect 4604 3896 4612 3904
rect 4620 3896 4628 3904
rect 4284 3876 4292 3884
rect 4396 3876 4404 3884
rect 4556 3856 4564 3864
rect 4140 3836 4148 3844
rect 4364 3796 4372 3804
rect 4156 3756 4164 3764
rect 4284 3756 4292 3764
rect 4492 3716 4500 3724
rect 4300 3696 4308 3704
rect 4508 3696 4516 3704
rect 4124 3576 4132 3584
rect 4476 3516 4484 3524
rect 4732 3756 4740 3764
rect 4764 3756 4772 3764
rect 4748 3676 4756 3684
rect 4572 3556 4580 3564
rect 4300 3496 4308 3504
rect 4508 3496 4516 3504
rect 4540 3496 4548 3504
rect 4092 3476 4100 3484
rect 4124 3456 4132 3464
rect 4236 3436 4244 3444
rect 4284 3436 4292 3444
rect 4156 3336 4164 3344
rect 4076 3316 4084 3324
rect 3612 3296 3620 3304
rect 4092 3296 4100 3304
rect 3612 3276 3620 3284
rect 4060 3276 4068 3284
rect 3612 3256 3620 3264
rect 3788 3256 3796 3264
rect 3148 3116 3156 3124
rect 3452 3116 3460 3124
rect 3532 3116 3540 3124
rect 3756 3116 3764 3124
rect 2412 3096 2420 3104
rect 2476 3096 2484 3104
rect 2844 3096 2852 3104
rect 2860 3096 2868 3104
rect 2460 3016 2468 3024
rect 2092 2956 2100 2964
rect 1980 2936 1988 2944
rect 1756 2916 1764 2924
rect 2028 2916 2036 2924
rect 2316 2916 2324 2924
rect 1836 2896 1844 2904
rect 1596 2876 1604 2884
rect 1836 2876 1844 2884
rect 1548 2856 1556 2864
rect 1292 2756 1300 2764
rect 1228 2736 1236 2744
rect 1084 2716 1092 2724
rect 1452 2716 1460 2724
rect 1148 2676 1156 2684
rect 1244 2676 1252 2684
rect 1356 2656 1364 2664
rect 1356 2636 1364 2644
rect 1356 2616 1364 2624
rect 1132 2596 1140 2604
rect 1340 2576 1348 2584
rect 1004 2556 1012 2564
rect 572 2536 580 2544
rect 748 2536 756 2544
rect 780 2536 788 2544
rect 1228 2536 1236 2544
rect 892 2496 900 2504
rect 700 2476 708 2484
rect 508 2376 516 2384
rect 492 2336 500 2344
rect 652 2336 660 2344
rect 492 2316 500 2324
rect 876 2296 884 2304
rect 652 2276 660 2284
rect 684 2276 692 2284
rect 876 2276 884 2284
rect 492 2256 500 2264
rect 684 2256 692 2264
rect 524 2156 532 2164
rect 652 2156 660 2164
rect 668 2116 676 2124
rect 508 2016 516 2024
rect 652 1876 660 1884
rect 636 1856 644 1864
rect 652 1756 660 1764
rect 524 1736 532 1744
rect 668 1716 676 1724
rect 540 1516 548 1524
rect 540 1476 548 1484
rect 652 1476 660 1484
rect 668 1416 676 1424
rect 540 1336 548 1344
rect 652 1296 660 1304
rect 652 1136 660 1144
rect 700 2176 708 2184
rect 988 2476 996 2484
rect 1212 2496 1220 2504
rect 1004 2316 1012 2324
rect 1308 2336 1316 2344
rect 1324 2316 1332 2324
rect 1100 2256 1108 2264
rect 1132 2256 1140 2264
rect 1292 2256 1300 2264
rect 1308 2256 1316 2264
rect 956 2176 964 2184
rect 1180 2176 1188 2184
rect 956 2156 964 2164
rect 972 2136 980 2144
rect 1324 2096 1332 2104
rect 1164 2076 1172 2084
rect 956 2056 964 2064
rect 956 1956 964 1964
rect 860 1936 868 1944
rect 764 1876 772 1884
rect 956 1876 964 1884
rect 716 1756 724 1764
rect 860 1856 868 1864
rect 1164 1856 1172 1864
rect 1308 1856 1316 1864
rect 1340 1836 1348 1844
rect 1116 1796 1124 1804
rect 1340 1796 1348 1804
rect 764 1736 772 1744
rect 1180 1736 1188 1744
rect 1212 1736 1220 1744
rect 748 1696 756 1704
rect 748 1516 756 1524
rect 1212 1676 1220 1684
rect 1116 1656 1124 1664
rect 940 1556 948 1564
rect 972 1556 980 1564
rect 1148 1496 1156 1504
rect 764 1476 772 1484
rect 876 1436 884 1444
rect 732 1356 740 1364
rect 988 1476 996 1484
rect 1324 1476 1332 1484
rect 1116 1416 1124 1424
rect 1996 2856 2004 2864
rect 1852 2796 1860 2804
rect 2092 2896 2100 2904
rect 2284 2856 2292 2864
rect 2332 2856 2340 2864
rect 2236 2816 2244 2824
rect 2252 2756 2260 2764
rect 2028 2716 2036 2724
rect 1660 2696 1668 2704
rect 2252 2696 2260 2704
rect 2012 2676 2020 2684
rect 1660 2656 1668 2664
rect 1692 2656 1700 2664
rect 2092 2656 2100 2664
rect 1660 2616 1668 2624
rect 1420 2576 1428 2584
rect 1804 2536 1812 2544
rect 1836 2536 1844 2544
rect 2028 2536 2036 2544
rect 1436 2496 1444 2504
rect 1820 2496 1828 2504
rect 2012 2396 2020 2404
rect 1596 2336 1604 2344
rect 1980 2316 1988 2324
rect 1756 2296 1764 2304
rect 1772 2296 1780 2304
rect 1548 2276 1556 2284
rect 1644 2256 1652 2264
rect 1628 2236 1634 2244
rect 1634 2236 1636 2244
rect 1836 2236 1844 2244
rect 1804 2196 1812 2204
rect 1388 2156 1396 2164
rect 1644 2156 1652 2164
rect 1772 2156 1780 2164
rect 1548 2076 1556 2084
rect 1804 1916 1812 1924
rect 1420 1856 1428 1864
rect 1612 1856 1620 1864
rect 1756 1856 1764 1864
rect 1772 1856 1780 1864
rect 1820 1856 1828 1864
rect 1580 1836 1588 1844
rect 1628 1816 1636 1824
rect 1644 1796 1652 1804
rect 1436 1756 1444 1764
rect 1788 1716 1796 1724
rect 1820 1716 1828 1724
rect 1628 1596 1636 1604
rect 1548 1516 1556 1524
rect 1612 1496 1620 1504
rect 1644 1476 1652 1484
rect 1580 1396 1588 1404
rect 1212 1356 1220 1364
rect 1676 1356 1684 1364
rect 732 1336 740 1344
rect 1196 1336 1204 1344
rect 876 1316 884 1324
rect 876 1296 884 1304
rect 1564 1296 1572 1304
rect 940 1276 948 1284
rect 892 1236 900 1244
rect 908 1136 916 1144
rect 972 1256 980 1264
rect 1660 1256 1668 1264
rect 1372 1176 1380 1184
rect 748 1116 756 1124
rect 940 1096 948 1104
rect 1116 1096 1124 1104
rect 1164 1096 1172 1104
rect 1196 1096 1204 1104
rect 1356 1096 1364 1104
rect 972 1076 980 1084
rect 764 1056 772 1064
rect 524 1036 532 1044
rect 908 1036 916 1044
rect 476 996 484 1004
rect 684 996 692 1004
rect 204 956 212 964
rect 652 956 660 964
rect 428 936 436 944
rect 508 916 516 924
rect 892 916 900 924
rect 428 896 436 904
rect 236 796 244 804
rect 428 736 436 744
rect 444 676 452 684
rect 92 656 100 664
rect 76 596 84 604
rect 204 556 212 564
rect 924 976 932 984
rect 1196 976 1204 984
rect 1324 936 1332 944
rect 1116 916 1124 924
rect 1116 896 1124 904
rect 1340 876 1348 884
rect 956 736 964 744
rect 892 716 900 724
rect 540 676 548 684
rect 972 696 980 704
rect 1100 676 1108 684
rect 1308 676 1316 684
rect 956 656 964 664
rect 652 556 660 564
rect 684 556 692 564
rect 316 516 324 524
rect 956 616 964 624
rect 1148 596 1156 604
rect 860 556 868 564
rect 1100 556 1108 564
rect 1132 556 1140 564
rect 892 536 900 544
rect 300 496 308 504
rect 620 496 628 504
rect 220 396 228 404
rect 1356 596 1364 604
rect 1324 556 1332 564
rect 1564 1156 1572 1164
rect 1388 1096 1396 1104
rect 2236 2536 2244 2544
rect 2092 2496 2100 2504
rect 2076 2396 2084 2404
rect 2204 2336 2212 2344
rect 2092 2276 2100 2284
rect 2172 2276 2180 2284
rect 2060 2236 2068 2244
rect 2316 2776 2324 2784
rect 2316 2756 2324 2764
rect 2524 3076 2532 3084
rect 2716 3076 2724 3084
rect 3052 3076 3060 3084
rect 3308 3076 3316 3084
rect 3340 3076 3348 3084
rect 3532 3076 3540 3084
rect 3756 3076 3764 3084
rect 2668 3056 2676 3064
rect 3180 3036 3188 3044
rect 2540 2996 2548 3004
rect 2684 2936 2692 2944
rect 2924 2996 2932 3004
rect 2716 2976 2724 2984
rect 2892 2936 2900 2944
rect 2892 2896 2900 2904
rect 3164 3016 3172 3024
rect 3116 2956 3124 2964
rect 2892 2816 2900 2824
rect 2940 2816 2948 2824
rect 2700 2756 2708 2764
rect 2476 2696 2484 2704
rect 2988 2776 2996 2784
rect 2924 2716 2932 2724
rect 2460 2676 2468 2684
rect 2492 2656 2500 2664
rect 2748 2656 2756 2664
rect 2892 2656 2900 2664
rect 2940 2656 2948 2664
rect 3100 2656 3108 2664
rect 3132 2656 3140 2664
rect 2364 2536 2372 2544
rect 2492 2536 2500 2544
rect 3132 2616 3140 2624
rect 3148 2596 3156 2604
rect 3324 3016 3332 3024
rect 3372 2996 3380 3004
rect 3836 3176 3844 3184
rect 4204 3136 4212 3144
rect 5276 4256 5284 4264
rect 5164 4176 5172 4184
rect 5052 4156 5060 4164
rect 5260 4156 5268 4164
rect 4924 4136 4932 4144
rect 4940 4136 4948 4144
rect 4972 4116 4980 4124
rect 5388 4276 5396 4284
rect 5756 4276 5764 4284
rect 5916 4256 5924 4264
rect 5660 4236 5668 4244
rect 5068 4136 5076 4144
rect 5308 4136 5316 4144
rect 5388 4116 5396 4124
rect 5628 4116 5636 4124
rect 5756 4216 5764 4224
rect 6380 4296 6388 4304
rect 7436 4516 7444 4524
rect 7900 4516 7908 4524
rect 8124 4516 8132 4524
rect 8476 4516 8484 4524
rect 7260 4496 7268 4504
rect 7468 4476 7476 4484
rect 7836 4356 7844 4364
rect 7884 4356 7892 4364
rect 7900 4356 7908 4364
rect 7212 4316 7220 4324
rect 7260 4316 7268 4324
rect 7324 4316 7332 4324
rect 7452 4316 7460 4324
rect 7708 4316 7716 4324
rect 7468 4296 7476 4304
rect 7548 4296 7556 4304
rect 6156 4276 6164 4284
rect 7660 4276 7668 4284
rect 7692 4276 7700 4284
rect 6188 4256 6196 4264
rect 6604 4256 6612 4264
rect 6780 4256 6788 4264
rect 6012 4236 6020 4244
rect 6348 4196 6356 4204
rect 6156 4176 6164 4184
rect 5964 4156 5972 4164
rect 5980 4156 5988 4164
rect 5756 4136 5764 4144
rect 5420 4096 5428 4104
rect 5740 4076 5748 4084
rect 5964 4076 5972 4084
rect 5292 3996 5300 4004
rect 5484 3996 5492 4004
rect 5068 3936 5076 3944
rect 4844 3916 4852 3924
rect 5068 3896 5076 3904
rect 4828 3876 4836 3884
rect 5516 3936 5524 3944
rect 5724 3936 5732 3944
rect 5868 3936 5876 3944
rect 6092 3936 6100 3944
rect 5484 3876 5492 3884
rect 5868 3876 5876 3884
rect 6204 4156 6212 4164
rect 6668 4216 6676 4224
rect 6588 4196 6596 4204
rect 6412 4136 6420 4144
rect 6460 4136 6468 4144
rect 6188 4096 6196 4104
rect 6188 4056 6196 4064
rect 6428 4056 6436 4064
rect 6812 4236 6820 4244
rect 6892 4236 6900 4244
rect 7196 4196 7204 4204
rect 7068 4156 7076 4164
rect 7116 4156 7124 4164
rect 7564 4216 7572 4224
rect 7388 4156 7396 4164
rect 7484 4156 7492 4164
rect 7244 4136 7252 4144
rect 6732 4096 6740 4104
rect 6844 4096 6852 4104
rect 6172 3936 6180 3944
rect 6636 3936 6644 3944
rect 6380 3916 6388 3924
rect 7372 4096 7380 4104
rect 6972 4056 6980 4064
rect 6748 3976 6756 3984
rect 6860 3976 6868 3984
rect 6988 3976 6996 3984
rect 7260 3916 7268 3924
rect 6828 3896 6836 3904
rect 7164 3896 7172 3904
rect 6188 3876 6196 3884
rect 6828 3876 6836 3884
rect 5260 3836 5268 3844
rect 4796 3776 4804 3784
rect 4956 3756 4964 3764
rect 5500 3856 5508 3864
rect 5708 3856 5716 3864
rect 6060 3856 6068 3864
rect 6156 3856 6164 3864
rect 5196 3756 5204 3764
rect 5420 3756 5428 3764
rect 5532 3736 5540 3744
rect 6636 3856 6644 3864
rect 6412 3776 6420 3784
rect 6588 3756 6596 3764
rect 7100 3836 7108 3844
rect 6828 3796 6836 3804
rect 6988 3776 6996 3784
rect 7020 3776 7028 3784
rect 6172 3736 6180 3744
rect 4988 3716 4996 3724
rect 5196 3716 5204 3724
rect 5420 3716 5428 3724
rect 5740 3696 5748 3704
rect 5532 3676 5540 3684
rect 6172 3716 6180 3724
rect 6588 3716 6596 3724
rect 6972 3716 6980 3724
rect 7468 4076 7476 4084
rect 7484 4076 7492 4084
rect 7404 4056 7412 4064
rect 7484 3916 7492 3924
rect 7388 3896 7396 3904
rect 7468 3876 7476 3884
rect 7612 3876 7620 3884
rect 7244 3856 7252 3864
rect 7196 3816 7204 3824
rect 7180 3776 7188 3784
rect 7100 3736 7108 3744
rect 6172 3676 6180 3684
rect 5756 3636 5764 3644
rect 4924 3536 4932 3544
rect 4780 3516 4788 3524
rect 4796 3496 4804 3504
rect 4460 3476 4468 3484
rect 4572 3456 4580 3464
rect 4620 3436 4628 3444
rect 4716 3436 4724 3444
rect 4332 3396 4340 3404
rect 4940 3356 4948 3364
rect 4316 3336 4324 3344
rect 4508 3336 4516 3344
rect 4620 3336 4628 3344
rect 6604 3676 6612 3684
rect 6396 3556 6404 3564
rect 6572 3556 6580 3564
rect 5148 3536 5156 3544
rect 5372 3536 5380 3544
rect 5804 3536 5812 3544
rect 5900 3536 5908 3544
rect 6124 3536 6132 3544
rect 5388 3516 5396 3524
rect 5324 3476 5332 3484
rect 5804 3476 5812 3484
rect 6124 3476 6132 3484
rect 5148 3456 5156 3464
rect 5468 3456 5476 3464
rect 5916 3456 5924 3464
rect 5660 3436 5668 3444
rect 5180 3316 5188 3324
rect 5724 3396 5732 3404
rect 6284 3396 6292 3404
rect 5612 3376 5620 3384
rect 5692 3376 5700 3384
rect 5724 3376 5732 3384
rect 5740 3376 5748 3384
rect 6060 3376 6068 3384
rect 6092 3376 6100 3384
rect 6172 3376 6180 3384
rect 5500 3356 5508 3364
rect 5516 3356 5524 3364
rect 5292 3336 5300 3344
rect 6540 3496 6548 3504
rect 6572 3476 6580 3484
rect 6940 3556 6948 3564
rect 6780 3496 6788 3504
rect 7164 3496 7172 3504
rect 7116 3476 7124 3484
rect 7068 3456 7076 3464
rect 6844 3436 6852 3444
rect 6764 3416 6772 3424
rect 6764 3396 6772 3404
rect 6636 3356 6644 3364
rect 7212 3776 7220 3784
rect 7468 3756 7476 3764
rect 7388 3736 7396 3744
rect 7500 3696 7508 3704
rect 7228 3516 7236 3524
rect 7244 3476 7252 3484
rect 7228 3456 7236 3464
rect 7324 3436 7332 3444
rect 7180 3376 7188 3384
rect 7580 3516 7588 3524
rect 7500 3476 7508 3484
rect 7404 3376 7412 3384
rect 7564 3456 7572 3464
rect 6204 3336 6212 3344
rect 6540 3336 6548 3344
rect 6924 3336 6932 3344
rect 7100 3336 7108 3344
rect 7308 3336 7316 3344
rect 7388 3336 7396 3344
rect 7436 3336 7444 3344
rect 7484 3336 7492 3344
rect 4524 3296 4532 3304
rect 4716 3296 4724 3304
rect 5004 3296 5012 3304
rect 5196 3296 5204 3304
rect 5948 3296 5956 3304
rect 6284 3296 6292 3304
rect 6540 3296 6548 3304
rect 5500 3276 5508 3284
rect 7276 3316 7284 3324
rect 6860 3296 6868 3304
rect 6620 3256 6628 3264
rect 6844 3256 6852 3264
rect 4620 3176 4628 3184
rect 4572 3136 4580 3144
rect 5772 3176 5780 3184
rect 5436 3156 5444 3164
rect 5132 3136 5138 3144
rect 5138 3136 5140 3144
rect 5356 3136 5364 3144
rect 5468 3136 5476 3144
rect 6156 3156 6164 3164
rect 6412 3156 6420 3164
rect 5884 3136 5892 3144
rect 6652 3136 6660 3144
rect 6860 3136 6868 3144
rect 5260 3116 5268 3124
rect 4284 3096 4292 3104
rect 4828 3096 4836 3104
rect 5052 3096 5060 3104
rect 5564 3096 5572 3104
rect 6428 3096 6436 3104
rect 4204 3076 4212 3084
rect 4572 3076 4580 3084
rect 4636 3076 4644 3084
rect 4748 3076 4756 3084
rect 4828 3076 4836 3084
rect 5564 3076 5572 3084
rect 5788 3076 5796 3084
rect 5996 3076 6004 3084
rect 6652 3076 6660 3084
rect 3868 3056 3876 3064
rect 3980 3056 3988 3064
rect 4428 3036 4436 3044
rect 4540 3036 4548 3044
rect 4476 3016 4484 3024
rect 4524 3016 4532 3024
rect 4236 2956 4244 2964
rect 4348 2936 4356 2944
rect 3420 2916 3428 2924
rect 3196 2896 3204 2904
rect 3596 2916 3604 2924
rect 3788 2916 3796 2924
rect 4652 3056 4660 3064
rect 4700 2996 4708 3004
rect 5036 3056 5044 3064
rect 5244 3056 5252 3064
rect 5372 3056 5380 3064
rect 5644 3056 5652 3064
rect 6204 3056 6212 3064
rect 6876 3056 6884 3064
rect 4924 3036 4932 3044
rect 4972 3036 4980 3044
rect 4988 3036 4996 3044
rect 4908 2956 4916 2964
rect 4572 2916 4580 2924
rect 3804 2896 3812 2904
rect 4236 2896 4244 2904
rect 4316 2896 4324 2904
rect 4924 2896 4932 2904
rect 3356 2856 3364 2864
rect 3580 2856 3588 2864
rect 3596 2796 3604 2804
rect 3596 2756 3604 2764
rect 3836 2756 3844 2764
rect 4540 2876 4548 2884
rect 4316 2776 4324 2784
rect 4092 2756 4100 2764
rect 4012 2736 4020 2744
rect 4668 2756 4676 2764
rect 4876 2756 4884 2764
rect 3228 2716 3236 2724
rect 3372 2716 3380 2724
rect 4012 2716 4020 2724
rect 4316 2716 4324 2724
rect 3212 2676 3220 2684
rect 2764 2556 2772 2564
rect 3020 2556 3028 2564
rect 2812 2536 2820 2544
rect 3644 2696 3652 2704
rect 4220 2696 4228 2704
rect 4492 2696 4500 2704
rect 3564 2656 3572 2664
rect 3996 2676 4004 2684
rect 4204 2676 4212 2684
rect 4300 2676 4308 2684
rect 3788 2656 3796 2664
rect 3868 2656 3876 2664
rect 3884 2636 3892 2644
rect 3436 2596 3444 2604
rect 3420 2556 3428 2564
rect 3612 2556 3620 2564
rect 3868 2616 3876 2624
rect 3660 2596 3668 2604
rect 3836 2556 3844 2564
rect 3036 2536 3044 2544
rect 3644 2536 3652 2544
rect 3372 2516 3380 2524
rect 4092 2556 4100 2564
rect 4300 2556 4308 2564
rect 4316 2556 4324 2564
rect 4092 2536 4100 2544
rect 4108 2536 4116 2544
rect 7228 3116 7236 3124
rect 7212 3096 7220 3104
rect 8428 4336 8436 4344
rect 8476 4336 8484 4344
rect 8188 4316 8196 4324
rect 7884 4296 7892 4304
rect 8092 4276 8100 4284
rect 7916 4256 7924 4264
rect 7948 4256 7956 4264
rect 7740 4216 7748 4224
rect 7836 4156 7844 4164
rect 8412 4296 8420 4304
rect 8604 4496 8612 4504
rect 8812 4496 8820 4504
rect 8540 4316 8548 4324
rect 8220 4276 8228 4284
rect 8332 4196 8340 4204
rect 8492 4196 8500 4204
rect 8524 4196 8532 4204
rect 8812 4356 8820 4364
rect 8620 4336 8628 4344
rect 8620 4316 8628 4324
rect 8636 4276 8644 4284
rect 8828 4336 8836 4344
rect 9228 4556 9236 4564
rect 9116 4536 9124 4544
rect 9212 4536 9220 4544
rect 9132 4476 9140 4484
rect 9180 4436 9188 4444
rect 9212 4336 9220 4344
rect 8924 4316 8932 4324
rect 8844 4296 8852 4304
rect 9132 4276 9140 4284
rect 9036 4236 9044 4244
rect 8604 4176 8612 4184
rect 8956 4156 8964 4164
rect 7964 4136 7972 4144
rect 8124 4136 8132 4144
rect 7676 4116 7684 4124
rect 7836 4116 7844 4124
rect 7932 4116 7940 4124
rect 8348 4116 8356 4124
rect 8732 4116 8740 4124
rect 8492 4096 8494 4104
rect 8494 4096 8500 4104
rect 8956 4096 8964 4104
rect 7836 4076 7844 4084
rect 8732 4076 8740 4084
rect 9148 4256 9156 4264
rect 9164 4256 9172 4264
rect 9356 4316 9364 4324
rect 10028 4596 10036 4604
rect 9548 4556 9556 4564
rect 9580 4556 9588 4564
rect 9404 4536 9412 4544
rect 9772 4536 9780 4544
rect 9788 4496 9796 4504
rect 9884 4456 9892 4464
rect 9548 4356 9556 4364
rect 9612 4336 9620 4344
rect 9852 4336 9860 4344
rect 9388 4296 9396 4304
rect 9372 4276 9380 4284
rect 9820 4276 9828 4284
rect 9132 4176 9140 4184
rect 9148 4176 9156 4184
rect 9036 4156 9044 4164
rect 9036 4116 9044 4124
rect 9132 4096 9140 4104
rect 8892 3956 8900 3964
rect 8988 3956 8996 3964
rect 9068 3956 9076 3964
rect 7900 3936 7908 3944
rect 8540 3936 8548 3944
rect 9932 4296 9940 4304
rect 9500 4176 9508 4184
rect 10060 4196 10068 4204
rect 9900 4136 9908 4144
rect 9276 4116 9284 4124
rect 9484 4116 9492 4124
rect 9708 4116 9716 4124
rect 9276 4096 9284 4104
rect 9580 4076 9588 4084
rect 9916 4076 9924 4084
rect 9260 4056 9268 4064
rect 9628 4016 9636 4024
rect 9436 3936 9444 3944
rect 9212 3916 9220 3924
rect 7692 3896 7700 3904
rect 9100 3896 9108 3904
rect 7916 3876 7924 3884
rect 8092 3876 8100 3884
rect 8460 3876 8468 3884
rect 8764 3876 8772 3884
rect 8780 3876 8788 3884
rect 7676 3856 7684 3864
rect 7820 3836 7828 3844
rect 8044 3856 8052 3864
rect 7676 3776 7684 3784
rect 7692 3756 7700 3764
rect 7868 3736 7876 3744
rect 7884 3676 7892 3684
rect 7676 3556 7684 3564
rect 7900 3516 7908 3524
rect 8300 3836 8308 3844
rect 8364 3816 8372 3824
rect 8476 3816 8484 3824
rect 8316 3776 8324 3784
rect 8172 3756 8180 3764
rect 8604 3756 8612 3764
rect 8732 3796 8740 3804
rect 8396 3736 8404 3744
rect 8700 3736 8708 3744
rect 8172 3696 8180 3704
rect 8140 3676 8148 3684
rect 8124 3616 8132 3624
rect 7916 3476 7924 3484
rect 7692 3456 7700 3464
rect 7708 3376 7716 3384
rect 7820 3376 7828 3384
rect 7308 3276 7316 3284
rect 7644 3276 7652 3284
rect 7276 3076 7284 3084
rect 7420 3076 7428 3084
rect 7356 3056 7364 3064
rect 7964 3316 7972 3324
rect 7948 3276 7956 3284
rect 7740 3236 7748 3244
rect 7884 3236 7892 3244
rect 7516 3076 7524 3084
rect 7676 3076 7684 3084
rect 6060 3036 6068 3044
rect 6348 3036 6356 3044
rect 6924 3036 6932 3044
rect 7068 3036 7076 3044
rect 5564 2956 5572 2964
rect 5132 2936 5140 2944
rect 5164 2936 5172 2944
rect 5356 2936 5364 2944
rect 5724 2936 5732 2944
rect 6012 2936 6020 2944
rect 5132 2836 5140 2844
rect 4972 2736 4980 2744
rect 4892 2696 4900 2704
rect 4972 2696 4980 2704
rect 4588 2676 4596 2684
rect 4508 2636 4516 2644
rect 4556 2636 4564 2644
rect 4492 2576 4500 2584
rect 4748 2616 4756 2624
rect 5356 2916 5364 2924
rect 6140 2976 6148 2984
rect 6252 2956 6260 2964
rect 6572 2956 6580 2964
rect 6092 2936 6100 2944
rect 6236 2936 6244 2944
rect 6572 2936 6580 2944
rect 6812 2936 6820 2944
rect 6908 2936 6916 2944
rect 6748 2916 6756 2924
rect 5580 2896 5588 2904
rect 6236 2896 6244 2904
rect 6332 2896 6340 2904
rect 6444 2896 6452 2904
rect 6540 2896 6548 2904
rect 7020 3016 7028 3024
rect 7004 2996 7012 3004
rect 7228 2996 7236 3004
rect 6972 2976 6980 2984
rect 7292 2976 7300 2984
rect 7004 2916 7012 2924
rect 7100 2896 7108 2904
rect 7196 2896 7204 2904
rect 5180 2736 5188 2744
rect 5532 2716 5540 2724
rect 5164 2696 5172 2704
rect 5516 2676 5524 2684
rect 5628 2676 5636 2684
rect 5196 2656 5204 2664
rect 5484 2656 5492 2664
rect 5612 2656 5620 2664
rect 5324 2636 5332 2644
rect 5372 2636 5380 2644
rect 5148 2596 5156 2604
rect 6060 2876 6068 2884
rect 6716 2776 6724 2784
rect 6636 2736 6644 2744
rect 7148 2796 7156 2804
rect 6188 2716 6196 2724
rect 6268 2716 6276 2724
rect 6492 2716 6500 2724
rect 6748 2716 6756 2724
rect 6892 2716 6900 2724
rect 6028 2696 6036 2704
rect 6620 2696 6628 2704
rect 6188 2676 6196 2684
rect 5836 2656 5844 2664
rect 6268 2656 6276 2664
rect 6556 2656 6564 2664
rect 5788 2616 5796 2624
rect 5900 2596 5908 2604
rect 4620 2556 4628 2564
rect 4764 2556 4772 2564
rect 5132 2556 5140 2564
rect 5980 2556 5988 2564
rect 6204 2556 6212 2564
rect 6940 2656 6948 2664
rect 6828 2596 6836 2604
rect 6620 2576 6628 2584
rect 6652 2576 6660 2584
rect 6780 2576 6788 2584
rect 4380 2536 4388 2544
rect 4476 2536 4484 2544
rect 4972 2536 4980 2544
rect 5324 2536 5332 2544
rect 5548 2536 5556 2544
rect 5980 2536 5988 2544
rect 6396 2536 6404 2544
rect 6476 2536 6484 2544
rect 6764 2536 6772 2544
rect 4540 2516 4548 2524
rect 5084 2516 5092 2524
rect 5756 2516 5764 2524
rect 6188 2516 6196 2524
rect 7596 2996 7604 3004
rect 7404 2976 7412 2984
rect 7564 2956 7572 2964
rect 7644 2896 7652 2904
rect 7708 3016 7716 3024
rect 7788 2996 7796 3004
rect 8092 3116 8100 3124
rect 8060 3076 8068 3084
rect 7916 3056 7924 3064
rect 7932 3036 7940 3044
rect 7868 2976 7876 2984
rect 7676 2956 7684 2964
rect 7692 2956 7700 2964
rect 7884 2896 7892 2904
rect 8012 2916 8020 2924
rect 7996 2876 8004 2884
rect 7564 2756 7572 2764
rect 7660 2756 7668 2764
rect 7788 2736 7796 2744
rect 8108 3076 8116 3084
rect 8092 3056 8100 3064
rect 8348 3576 8356 3584
rect 8380 3576 8388 3584
rect 8572 3576 8580 3584
rect 9452 3876 9460 3884
rect 9212 3856 9220 3864
rect 9132 3836 9140 3844
rect 8972 3796 8980 3804
rect 8988 3776 8996 3784
rect 9276 3756 9284 3764
rect 9356 3756 9364 3764
rect 9452 3756 9460 3764
rect 8844 3736 8852 3744
rect 9164 3736 9172 3744
rect 9500 3736 9508 3744
rect 8828 3716 8836 3724
rect 9020 3716 9028 3724
rect 9180 3716 9188 3724
rect 9260 3716 9268 3724
rect 9468 3716 9476 3724
rect 9020 3556 9028 3564
rect 9452 3516 9460 3524
rect 8492 3496 8500 3504
rect 9036 3496 9044 3504
rect 9228 3496 9236 3504
rect 9244 3496 9252 3504
rect 8348 3476 8356 3484
rect 8572 3476 8580 3484
rect 8812 3476 8820 3484
rect 8476 3456 8484 3464
rect 8572 3456 8580 3464
rect 9020 3456 9028 3464
rect 8588 3436 8596 3444
rect 8988 3436 8996 3444
rect 8268 3376 8276 3384
rect 8428 3356 8436 3364
rect 8188 3336 8196 3344
rect 8428 3316 8436 3324
rect 8188 3296 8196 3304
rect 8380 3296 8388 3304
rect 9468 3476 9476 3484
rect 9068 3436 9076 3444
rect 10268 4176 10276 4184
rect 9884 3956 9892 3964
rect 10076 3956 10084 3964
rect 9660 3916 9668 3924
rect 9852 3916 9860 3924
rect 9644 3896 9652 3904
rect 9692 3756 9700 3764
rect 10092 3876 10100 3884
rect 10092 3796 10100 3804
rect 9820 3736 9828 3744
rect 10012 3736 10020 3744
rect 9852 3716 9860 3724
rect 9676 3536 9684 3544
rect 9900 3536 9908 3544
rect 10092 3516 10100 3524
rect 9692 3476 9700 3484
rect 9916 3476 9924 3484
rect 10252 3476 10260 3484
rect 9644 3356 9652 3364
rect 9836 3356 9844 3364
rect 8716 3336 8724 3344
rect 8860 3336 8868 3344
rect 9164 3336 9172 3344
rect 9244 3336 9252 3344
rect 9388 3336 9396 3344
rect 9612 3336 9620 3344
rect 8652 3316 8660 3324
rect 10060 3356 10068 3364
rect 9916 3336 9924 3344
rect 10044 3336 10052 3344
rect 8652 3296 8660 3304
rect 9484 3296 9492 3304
rect 8988 3156 8996 3164
rect 8540 3136 8548 3144
rect 8284 3116 8292 3124
rect 8396 3076 8404 3084
rect 8140 2996 8148 3004
rect 8236 2996 8244 3004
rect 8300 2996 8308 3004
rect 8460 2996 8468 3004
rect 8076 2976 8084 2984
rect 8092 2916 8100 2924
rect 8332 2916 8340 2924
rect 8332 2896 8340 2904
rect 8380 2836 8388 2844
rect 8060 2716 8068 2724
rect 7164 2696 7172 2704
rect 8204 2696 8212 2704
rect 8108 2676 8116 2684
rect 8124 2676 8132 2684
rect 7468 2636 7476 2644
rect 7500 2636 7508 2644
rect 7132 2596 7140 2604
rect 7004 2576 7012 2584
rect 7420 2556 7428 2564
rect 6876 2536 6884 2544
rect 6956 2516 6964 2524
rect 2332 2496 2340 2504
rect 2492 2496 2500 2504
rect 2540 2496 2548 2504
rect 2796 2496 2804 2504
rect 2876 2496 2884 2504
rect 3644 2496 3652 2504
rect 4972 2496 4974 2504
rect 4974 2496 4980 2504
rect 5084 2496 5092 2504
rect 5980 2496 5988 2504
rect 6956 2496 6964 2504
rect 7180 2496 7188 2504
rect 2428 2316 2436 2324
rect 2476 2316 2484 2324
rect 2412 2256 2420 2264
rect 2252 2116 2260 2124
rect 2428 2136 2436 2144
rect 2844 2316 2852 2324
rect 2508 2296 2516 2304
rect 7420 2496 7428 2504
rect 3388 2476 3396 2484
rect 5532 2476 5540 2484
rect 7404 2476 7412 2484
rect 5308 2456 5316 2464
rect 3100 2436 3108 2444
rect 3724 2356 3732 2364
rect 4684 2356 4692 2364
rect 5148 2356 5156 2364
rect 2524 2276 2532 2284
rect 2940 2276 2948 2284
rect 3068 2276 3076 2284
rect 2668 2216 2676 2224
rect 1996 2096 2004 2104
rect 2316 2096 2324 2104
rect 2060 2076 2068 2084
rect 2012 1956 2014 1964
rect 2014 1956 2020 1964
rect 2236 1956 2244 1964
rect 1884 1936 1892 1944
rect 2684 2056 2692 2064
rect 2684 1956 2692 1964
rect 2332 1936 2340 1944
rect 2476 1936 2484 1944
rect 2268 1916 2276 1924
rect 2700 1936 2708 1944
rect 2476 1856 2484 1864
rect 2684 1856 2692 1864
rect 1884 1796 1892 1804
rect 1868 1736 1876 1744
rect 2012 1736 2020 1744
rect 2044 1736 2052 1744
rect 2460 1816 2468 1824
rect 2908 2156 2916 2164
rect 2908 2096 2916 2104
rect 2780 1916 2788 1924
rect 3020 2156 3028 2164
rect 3932 2336 3940 2344
rect 4028 2336 4036 2344
rect 4236 2336 4244 2344
rect 4396 2336 4404 2344
rect 3180 2316 3188 2324
rect 3484 2316 3492 2324
rect 3628 2276 3636 2284
rect 3788 2276 3796 2284
rect 4044 2276 4052 2284
rect 4076 2276 4084 2284
rect 4412 2276 4420 2284
rect 2988 2096 2996 2104
rect 2940 1876 2948 1884
rect 2972 1856 2980 1864
rect 2940 1816 2948 1824
rect 2476 1756 2484 1764
rect 2252 1736 2260 1744
rect 2092 1716 2100 1724
rect 2028 1676 2036 1684
rect 2700 1756 2708 1764
rect 2796 1756 2804 1764
rect 2796 1716 2804 1724
rect 2700 1696 2708 1704
rect 2940 1696 2948 1704
rect 1852 1616 1860 1624
rect 2092 1536 2100 1544
rect 2332 1536 2340 1544
rect 2540 1536 2548 1544
rect 2300 1476 2308 1484
rect 2332 1476 2340 1484
rect 2028 1336 2036 1344
rect 2252 1416 2260 1424
rect 2316 1376 2324 1384
rect 2716 1436 2724 1444
rect 2700 1396 2708 1404
rect 2924 1376 2932 1384
rect 2108 1356 2116 1364
rect 2444 1356 2452 1364
rect 3004 2076 3012 2084
rect 3164 2076 3172 2084
rect 3004 1916 3012 1924
rect 3308 2256 3316 2264
rect 3372 2256 3378 2264
rect 3378 2256 3380 2264
rect 3484 2256 3492 2264
rect 3404 2236 3412 2244
rect 3420 2236 3428 2244
rect 3564 2236 3572 2244
rect 3244 2076 3252 2084
rect 3388 2016 3396 2024
rect 3372 1956 3380 1964
rect 3212 1936 3220 1944
rect 3180 1896 3188 1904
rect 3196 1876 3204 1884
rect 3020 1856 3028 1864
rect 3180 1856 3188 1864
rect 3036 1756 3044 1764
rect 3020 1656 3028 1664
rect 3132 1476 3140 1484
rect 3164 1476 3172 1484
rect 3148 1456 3156 1464
rect 3372 1856 3380 1864
rect 3212 1756 3220 1764
rect 3932 2256 3940 2264
rect 3868 2216 3876 2224
rect 3596 2156 3604 2164
rect 3836 2136 3844 2144
rect 3820 1956 3828 1964
rect 3852 1956 3860 1964
rect 3628 1936 3636 1944
rect 3596 1876 3604 1884
rect 3404 1756 3412 1764
rect 3228 1716 3236 1724
rect 3388 1696 3396 1704
rect 3660 1776 3668 1784
rect 3484 1716 3492 1724
rect 3484 1696 3492 1704
rect 3836 1796 3844 1804
rect 3692 1716 3700 1724
rect 3692 1696 3700 1704
rect 3692 1676 3700 1684
rect 3676 1656 3684 1664
rect 4412 2236 4420 2244
rect 4188 2216 4196 2224
rect 4060 2176 4068 2184
rect 5132 2316 5140 2324
rect 4924 2296 4932 2304
rect 4940 2296 4948 2304
rect 5276 2336 5284 2344
rect 5516 2336 5524 2344
rect 5292 2316 5300 2324
rect 5356 2296 5364 2304
rect 4812 2276 4820 2284
rect 4748 2256 4756 2264
rect 4940 2256 4948 2264
rect 5228 2256 5236 2264
rect 4636 2236 4644 2244
rect 4572 2156 4580 2164
rect 3932 2136 3940 2144
rect 4060 2136 4068 2144
rect 4268 2136 4276 2144
rect 4316 2136 4324 2144
rect 4476 2136 4484 2144
rect 4492 2136 4500 2144
rect 4540 2136 4548 2144
rect 4492 2116 4500 2124
rect 3916 2096 3924 2104
rect 4508 2096 4516 2104
rect 4076 1956 4084 1964
rect 4284 1936 4292 1944
rect 4140 1836 4148 1844
rect 4492 1936 4500 1944
rect 4476 1876 4484 1884
rect 4508 1876 4516 1884
rect 4316 1856 4324 1864
rect 4492 1856 4500 1864
rect 4268 1816 4276 1824
rect 4092 1776 4100 1784
rect 3900 1756 3908 1764
rect 4252 1756 4260 1764
rect 4300 1756 4308 1764
rect 3900 1716 3908 1724
rect 3932 1536 3940 1544
rect 4076 1536 4084 1544
rect 3916 1516 3924 1524
rect 3372 1476 3380 1484
rect 3452 1476 3460 1484
rect 3532 1476 3540 1484
rect 3644 1476 3652 1484
rect 3820 1476 3828 1484
rect 4156 1476 4164 1484
rect 4300 1476 4308 1484
rect 3388 1456 3396 1464
rect 3468 1436 3476 1444
rect 3420 1396 3428 1404
rect 3468 1396 3476 1404
rect 3596 1456 3604 1464
rect 3628 1416 3636 1424
rect 3596 1376 3604 1384
rect 2092 1336 2100 1344
rect 2476 1336 2484 1344
rect 2780 1336 2788 1344
rect 2988 1336 2996 1344
rect 1836 1176 1844 1184
rect 1836 1156 1844 1164
rect 2012 1096 2020 1104
rect 1756 1076 1764 1084
rect 2012 1076 2020 1084
rect 1628 1016 1636 1024
rect 1772 996 1780 1004
rect 1404 976 1412 984
rect 1836 976 1844 984
rect 1532 956 1540 964
rect 1772 956 1780 964
rect 1868 956 1876 964
rect 1404 916 1412 924
rect 1628 916 1636 924
rect 1644 916 1652 924
rect 1548 896 1556 904
rect 1740 876 1748 884
rect 1596 836 1604 844
rect 1532 736 1540 744
rect 2444 1316 2452 1324
rect 2556 1316 2564 1324
rect 2108 1296 2116 1304
rect 2572 1296 2580 1304
rect 2764 1296 2772 1304
rect 3116 1296 3124 1304
rect 3148 1296 3156 1304
rect 2972 1276 2980 1284
rect 3420 1216 3428 1224
rect 2668 1156 2676 1164
rect 3164 1156 3172 1164
rect 3324 1156 3332 1164
rect 2876 1136 2884 1144
rect 3372 1136 3380 1144
rect 2092 1096 2100 1104
rect 2668 1096 2676 1104
rect 2892 1096 2900 1104
rect 3084 1096 3092 1104
rect 2444 1076 2452 1084
rect 2108 1056 2116 1064
rect 2252 1036 2260 1044
rect 2732 1036 2740 1044
rect 2076 1016 2084 1024
rect 2060 976 2068 984
rect 2060 956 2068 964
rect 1740 716 1748 724
rect 1964 716 1972 724
rect 2044 716 2052 724
rect 1740 696 1748 704
rect 1948 696 1956 704
rect 1532 676 1540 684
rect 2028 676 2036 684
rect 1868 636 1876 644
rect 1580 576 1588 584
rect 1564 556 1572 564
rect 1164 476 1172 484
rect 1804 516 1812 524
rect 1836 516 1844 524
rect 1788 476 1796 484
rect 1820 476 1828 484
rect 892 456 900 464
rect 1564 456 1572 464
rect 428 316 436 324
rect 876 316 884 324
rect 188 296 196 304
rect 1532 356 1540 364
rect 1068 336 1076 344
rect 2476 996 2484 1004
rect 2268 976 2276 984
rect 2284 956 2292 964
rect 3116 996 3124 1004
rect 2492 976 2500 984
rect 2924 976 2932 984
rect 2940 976 2948 984
rect 2524 956 2532 964
rect 2972 956 2980 964
rect 3196 956 3204 964
rect 2940 936 2948 944
rect 2652 916 2660 924
rect 2668 916 2676 924
rect 2748 916 2756 924
rect 2764 916 2772 924
rect 3084 896 3092 904
rect 2636 736 2644 744
rect 2892 856 2900 864
rect 3180 876 3188 884
rect 3100 816 3108 824
rect 3404 1116 3412 1124
rect 3564 1136 3572 1144
rect 3580 1056 3588 1064
rect 3532 996 3540 1004
rect 3404 936 3412 944
rect 3772 1316 3780 1324
rect 4236 1356 4244 1364
rect 3772 1196 3780 1204
rect 3852 1176 3860 1184
rect 4044 1176 4052 1184
rect 4012 1156 4020 1164
rect 3644 1076 3652 1084
rect 3628 1056 3636 1064
rect 3996 1056 4004 1064
rect 4044 1036 4052 1044
rect 3772 1016 3780 1024
rect 3612 996 3620 1004
rect 4076 1176 4084 1184
rect 4204 1136 4212 1144
rect 4284 1136 4292 1144
rect 4236 1116 4244 1124
rect 4188 1076 4196 1084
rect 4460 1736 4468 1744
rect 4476 1676 4484 1684
rect 4476 1456 4484 1464
rect 4460 1336 4468 1344
rect 4444 1156 4452 1164
rect 4300 1116 4308 1124
rect 4428 1036 4436 1044
rect 4524 1836 4532 1844
rect 4572 2076 4580 2084
rect 4732 1936 4740 1944
rect 5068 2236 5076 2244
rect 4972 2196 4980 2204
rect 4812 2136 4820 2144
rect 5052 2096 5060 2104
rect 5164 2096 5172 2104
rect 4812 1916 4820 1924
rect 5020 1916 5028 1924
rect 5420 2236 5428 2244
rect 5484 2196 5492 2204
rect 5804 2456 5812 2464
rect 5724 2236 5732 2244
rect 6108 2436 6116 2444
rect 7276 2376 7284 2384
rect 6028 2336 6036 2344
rect 7500 2616 7508 2624
rect 8236 2656 8244 2664
rect 7660 2596 7668 2604
rect 7932 2596 7940 2604
rect 7580 2556 7588 2564
rect 7852 2556 7860 2564
rect 7884 2556 7892 2564
rect 8076 2596 8084 2604
rect 8108 2596 8116 2604
rect 7644 2536 7652 2544
rect 7884 2536 7892 2544
rect 7980 2536 7988 2544
rect 8284 2536 8292 2544
rect 8284 2516 8292 2524
rect 7644 2496 7652 2504
rect 8076 2396 8084 2404
rect 8124 2396 8132 2404
rect 7788 2336 7796 2344
rect 7964 2336 7972 2344
rect 7980 2336 7988 2344
rect 6236 2316 6244 2324
rect 6684 2316 6692 2324
rect 6908 2316 6916 2324
rect 7324 2316 7332 2324
rect 7468 2316 7476 2324
rect 6252 2296 6260 2304
rect 6028 2256 6036 2264
rect 5964 2236 5972 2244
rect 6172 2236 6180 2244
rect 5788 2196 5796 2204
rect 5868 2196 5876 2204
rect 5532 2176 5540 2184
rect 5612 2156 5620 2164
rect 5724 2116 5732 2124
rect 7132 2296 7140 2304
rect 7564 2296 7572 2304
rect 8332 2316 8340 2324
rect 6700 2276 6708 2284
rect 6892 2276 6900 2284
rect 7660 2276 7668 2284
rect 7772 2276 7780 2284
rect 8012 2276 8020 2284
rect 8300 2276 8308 2284
rect 8316 2276 8324 2284
rect 6924 2256 6932 2264
rect 6972 2256 6980 2264
rect 7132 2256 7140 2264
rect 7180 2256 7188 2264
rect 6476 2196 6484 2204
rect 6524 2196 6532 2204
rect 6364 2156 6372 2164
rect 7068 2216 7076 2224
rect 7356 2196 7364 2204
rect 7404 2196 7412 2204
rect 7852 2256 7860 2264
rect 7708 2216 7716 2224
rect 7708 2196 7716 2204
rect 7276 2156 7284 2164
rect 8060 2236 8068 2244
rect 7932 2216 7940 2224
rect 7868 2156 7876 2164
rect 6380 2136 6388 2144
rect 7052 2136 7060 2144
rect 6588 2116 6596 2124
rect 7484 2116 7492 2124
rect 5740 2096 5748 2104
rect 5948 2096 5956 2104
rect 6156 2096 6164 2104
rect 6812 2096 6820 2104
rect 7036 2096 7044 2104
rect 7388 2096 7396 2104
rect 5388 2056 5396 2064
rect 4716 1856 4724 1864
rect 4700 1796 4708 1804
rect 4556 1756 4564 1764
rect 4540 1636 4548 1644
rect 4588 1516 4596 1524
rect 4556 1376 4564 1384
rect 5020 1876 5028 1884
rect 5180 1896 5188 1904
rect 5260 1876 5268 1884
rect 5468 1876 5476 1884
rect 4956 1776 4964 1784
rect 5036 1776 5044 1784
rect 4940 1756 4948 1764
rect 5148 1756 5156 1764
rect 4796 1736 4804 1744
rect 4988 1736 4996 1744
rect 4796 1716 4804 1724
rect 5484 1796 5492 1804
rect 5628 1796 5636 1804
rect 5260 1736 5268 1744
rect 5420 1716 5428 1724
rect 5372 1696 5380 1704
rect 4764 1636 4772 1644
rect 5212 1656 5220 1664
rect 4924 1576 4932 1584
rect 5164 1536 5172 1544
rect 4956 1516 4964 1524
rect 4780 1496 4788 1504
rect 4716 1416 4724 1424
rect 4748 1416 4756 1424
rect 4588 1356 4596 1364
rect 4668 1336 4676 1344
rect 4524 1316 4532 1324
rect 4700 1296 4708 1304
rect 4556 1156 4564 1164
rect 4540 1116 4548 1124
rect 4684 1096 4692 1104
rect 4636 1036 4644 1044
rect 4268 956 4276 964
rect 3740 936 3748 944
rect 3948 936 3956 944
rect 4060 936 4068 944
rect 4188 916 4196 924
rect 3964 896 3972 904
rect 3164 716 3172 724
rect 3388 716 3396 724
rect 3084 696 3092 704
rect 2636 676 2644 684
rect 2668 676 2676 684
rect 3084 676 3092 684
rect 3180 676 3188 684
rect 3388 676 3396 684
rect 3724 676 3732 684
rect 2396 656 2404 664
rect 2204 616 2212 624
rect 1884 556 1892 564
rect 2012 556 2014 564
rect 2014 556 2020 564
rect 2236 556 2244 564
rect 1868 476 1876 484
rect 2700 616 2708 624
rect 2460 596 2468 604
rect 2332 556 2340 564
rect 2556 556 2564 564
rect 2300 516 2308 524
rect 2332 496 2338 504
rect 2338 496 2340 504
rect 2444 436 2452 444
rect 2476 436 2484 444
rect 2188 356 2196 364
rect 2268 356 2276 364
rect 3308 616 3316 624
rect 2876 596 2884 604
rect 2748 576 2756 584
rect 3356 576 3364 584
rect 2956 556 2964 564
rect 3100 556 3108 564
rect 3564 556 3572 564
rect 3132 536 3140 544
rect 3196 536 3204 544
rect 3340 536 3348 544
rect 3420 536 3428 544
rect 3516 536 3524 544
rect 3580 516 3588 524
rect 3676 556 3684 564
rect 3756 556 3764 564
rect 4028 876 4036 884
rect 4188 876 4196 884
rect 4252 836 4260 844
rect 3820 736 3828 744
rect 4172 676 4180 684
rect 3820 656 3828 664
rect 3788 596 3796 604
rect 3820 576 3828 584
rect 4460 936 4468 944
rect 4652 936 4660 944
rect 4428 876 4436 884
rect 4700 796 4708 804
rect 4636 736 4644 744
rect 4492 696 4500 704
rect 4412 676 4420 684
rect 4444 556 4452 564
rect 3772 536 3780 544
rect 3964 536 3972 544
rect 4012 536 4020 544
rect 4204 536 4212 544
rect 4268 536 4276 544
rect 3820 516 3828 524
rect 2892 476 2900 484
rect 3308 396 3316 404
rect 3100 356 3108 364
rect 2844 336 2852 344
rect 1292 316 1300 324
rect 1836 316 1844 324
rect 2652 316 2660 324
rect 2716 316 2724 324
rect 1740 296 1748 304
rect 1836 296 1844 304
rect 2412 296 2420 304
rect 620 276 628 284
rect 1196 276 1204 284
rect 1276 276 1284 284
rect 1740 276 1748 284
rect 412 256 420 264
rect 988 256 996 264
rect 1068 256 1076 264
rect 268 236 276 244
rect 748 236 756 244
rect 300 196 308 204
rect 492 196 500 204
rect 92 156 100 164
rect 924 216 932 224
rect 764 176 772 184
rect 556 136 564 144
rect 700 136 708 144
rect 1148 216 1156 224
rect 1356 216 1364 224
rect 1452 196 1460 204
rect 1004 156 1012 164
rect 1356 156 1364 164
rect 1388 156 1396 164
rect 1004 116 1012 124
rect 3532 356 3540 364
rect 3772 336 3780 344
rect 4092 496 4100 504
rect 4636 676 4644 684
rect 4636 596 4644 604
rect 4764 1396 4772 1404
rect 4812 1376 4820 1384
rect 4908 1176 4916 1184
rect 4780 1096 4788 1104
rect 4796 1056 4804 1064
rect 4732 996 4740 1004
rect 4860 936 4868 944
rect 4732 716 4740 724
rect 4892 916 4900 924
rect 4940 1096 4948 1104
rect 4924 896 4932 904
rect 5004 1496 5012 1504
rect 5148 1416 5156 1424
rect 5020 1356 5028 1364
rect 5340 1456 5348 1464
rect 5228 1336 5236 1344
rect 5340 1296 5348 1304
rect 5212 1276 5220 1284
rect 5020 1156 5028 1164
rect 5164 1156 5172 1164
rect 5004 1096 5012 1104
rect 5356 1096 5364 1104
rect 5372 1076 5380 1084
rect 5340 1036 5348 1044
rect 5356 1016 5364 1024
rect 5564 1476 5572 1484
rect 6380 2076 6388 2084
rect 7260 2076 7268 2084
rect 6956 2016 6964 2024
rect 7484 2076 7492 2084
rect 7692 2076 7700 2084
rect 7468 1976 7476 1984
rect 6108 1936 6116 1944
rect 6796 1936 6804 1944
rect 5724 1916 5732 1924
rect 5916 1916 5924 1924
rect 6700 1916 6702 1924
rect 6702 1916 6708 1924
rect 6780 1916 6788 1924
rect 5932 1896 5940 1904
rect 6780 1896 6788 1904
rect 6812 1896 6820 1904
rect 5708 1876 5716 1884
rect 6300 1876 6308 1884
rect 6492 1876 6500 1884
rect 6684 1876 6692 1884
rect 5788 1856 5796 1864
rect 6044 1856 6052 1864
rect 5820 1816 5828 1824
rect 5900 1756 5908 1764
rect 5788 1736 5796 1744
rect 5868 1736 5876 1744
rect 5676 1656 5684 1664
rect 5788 1516 5796 1524
rect 5820 1476 5828 1484
rect 5788 1456 5796 1464
rect 5660 1416 5668 1424
rect 5452 1336 5460 1344
rect 5820 1336 5828 1344
rect 5452 1276 5460 1284
rect 5804 1256 5812 1264
rect 5676 1156 5684 1164
rect 5452 1116 5460 1124
rect 5468 1076 5476 1084
rect 5596 1036 5598 1044
rect 5598 1036 5604 1044
rect 5580 1016 5588 1024
rect 5020 976 5028 984
rect 5100 936 5108 944
rect 5212 936 5220 944
rect 5548 936 5556 944
rect 5100 856 5108 864
rect 5676 956 5684 964
rect 5884 1676 5892 1684
rect 6076 1836 6084 1844
rect 6124 1736 6132 1744
rect 6284 1736 6292 1744
rect 6236 1656 6244 1664
rect 5884 1496 5892 1504
rect 5900 1476 5908 1484
rect 6684 1856 6692 1864
rect 6684 1756 6692 1764
rect 6444 1736 6452 1744
rect 6684 1716 6692 1724
rect 6700 1696 6708 1704
rect 6780 1696 6788 1704
rect 6444 1656 6452 1664
rect 6508 1636 6516 1644
rect 6492 1516 6500 1524
rect 6460 1476 6468 1484
rect 6060 1456 6068 1464
rect 6300 1456 6308 1464
rect 5916 1336 5924 1344
rect 6060 1336 6068 1344
rect 5900 1256 5908 1264
rect 6268 1256 6276 1264
rect 6700 1536 6708 1544
rect 6924 1536 6932 1544
rect 6796 1516 6804 1524
rect 6796 1496 6804 1504
rect 6684 1456 6692 1464
rect 6716 1456 6724 1464
rect 7036 1856 7044 1864
rect 7660 1956 7668 1964
rect 7676 1896 7684 1904
rect 7340 1876 7348 1884
rect 7372 1876 7380 1884
rect 6988 1776 6996 1784
rect 7212 1776 7220 1784
rect 7020 1716 7028 1724
rect 7452 1736 7460 1744
rect 7452 1696 7460 1704
rect 7244 1536 7252 1544
rect 7804 1816 7812 1824
rect 7644 1796 7652 1804
rect 7676 1776 7684 1784
rect 7804 1736 7812 1744
rect 7804 1716 7812 1724
rect 7852 1716 7860 1724
rect 8172 2216 8180 2224
rect 8988 3116 8996 3124
rect 9052 3116 9060 3124
rect 9196 3116 9204 3124
rect 9452 3116 9460 3124
rect 9692 3116 9700 3124
rect 8732 3076 8740 3084
rect 8812 3036 8820 3044
rect 8940 3036 8948 3044
rect 8732 2976 8740 2984
rect 8908 2936 8916 2944
rect 8556 2916 8564 2924
rect 8540 2896 8548 2904
rect 8556 2896 8564 2904
rect 8940 2876 8948 2884
rect 8620 2856 8628 2864
rect 8524 2736 8532 2744
rect 8428 2696 8436 2704
rect 9244 3096 9252 3104
rect 9484 3096 9492 3104
rect 9660 3096 9668 3104
rect 9244 3076 9252 3084
rect 9484 3056 9492 3064
rect 9020 3036 9028 3044
rect 9580 2996 9588 3004
rect 9628 2996 9636 3004
rect 9228 2976 9236 2984
rect 9132 2956 9140 2964
rect 9372 2956 9380 2964
rect 9612 2976 9620 2984
rect 9372 2916 9380 2924
rect 10044 3076 10052 3084
rect 9836 2976 9844 2984
rect 9692 2936 9700 2944
rect 9900 2936 9908 2944
rect 9884 2916 9892 2924
rect 9916 2916 9924 2924
rect 9148 2896 9156 2904
rect 9180 2876 9188 2884
rect 9676 2876 9684 2884
rect 8764 2716 8772 2724
rect 8956 2716 8964 2724
rect 8572 2676 8580 2684
rect 8620 2676 8628 2684
rect 8764 2676 8772 2684
rect 8844 2676 8852 2684
rect 8444 2556 8452 2564
rect 8508 2556 8516 2564
rect 8588 2556 8596 2564
rect 8396 2536 8404 2544
rect 8412 2276 8420 2284
rect 8492 2276 8500 2284
rect 8396 2256 8404 2264
rect 8124 2136 8132 2144
rect 7916 2096 7924 2104
rect 8124 2096 8132 2104
rect 8284 2096 8292 2104
rect 8556 2176 8564 2184
rect 8860 2636 8868 2644
rect 8956 2636 8964 2644
rect 8780 2576 8788 2584
rect 8764 2516 8772 2524
rect 8748 2436 8756 2444
rect 8940 2556 8948 2564
rect 8812 2536 8820 2544
rect 9148 2596 9156 2604
rect 9052 2536 9060 2544
rect 9036 2516 9044 2524
rect 8956 2476 8964 2484
rect 8780 2436 8788 2444
rect 8620 2336 8628 2344
rect 9516 2796 9524 2804
rect 9500 2716 9508 2724
rect 9212 2656 9220 2664
rect 9196 2636 9204 2644
rect 9660 2736 9668 2744
rect 9516 2696 9524 2704
rect 9692 2696 9700 2704
rect 9724 2676 9732 2684
rect 9436 2656 9444 2664
rect 9628 2576 9636 2584
rect 9852 2576 9860 2584
rect 9228 2516 9236 2524
rect 9244 2516 9252 2524
rect 9596 2516 9604 2524
rect 9596 2476 9604 2484
rect 9276 2336 9284 2344
rect 8844 2316 8852 2324
rect 8956 2316 8964 2324
rect 9164 2316 9172 2324
rect 9468 2316 9476 2324
rect 9612 2316 9620 2324
rect 9180 2296 9188 2304
rect 8988 2276 8996 2284
rect 9260 2276 9268 2284
rect 9596 2276 9604 2284
rect 8604 2256 8612 2264
rect 8636 2176 8644 2184
rect 8588 2156 8596 2164
rect 8700 2156 8708 2164
rect 8924 2156 8932 2164
rect 8668 2136 8676 2144
rect 8364 2116 8372 2124
rect 9132 2156 9140 2164
rect 8764 2136 8772 2144
rect 8988 2136 8996 2144
rect 9036 2136 9044 2144
rect 9244 2136 9252 2144
rect 8364 2096 8372 2104
rect 8492 2016 8500 2024
rect 8332 1976 8340 1984
rect 8364 1956 8372 1964
rect 7884 1916 7892 1924
rect 8124 1916 8132 1924
rect 8348 1916 8356 1924
rect 8124 1896 8132 1904
rect 9452 2156 9460 2164
rect 9468 2156 9476 2164
rect 9180 2116 9188 2124
rect 9420 2116 9428 2124
rect 9164 2096 9172 2104
rect 9468 1976 9476 1984
rect 9244 1956 9252 1964
rect 8588 1936 8596 1944
rect 8796 1936 8804 1944
rect 9148 1936 9156 1944
rect 9900 2896 9908 2904
rect 9916 2796 9924 2804
rect 9948 2716 9956 2724
rect 10076 2716 10084 2724
rect 9948 2696 9956 2704
rect 10124 2676 10132 2684
rect 10076 2596 10084 2604
rect 9708 2536 9716 2544
rect 9692 2496 9700 2504
rect 9868 2476 9876 2484
rect 9820 2296 9828 2304
rect 9820 2276 9828 2284
rect 9900 2336 9908 2344
rect 9916 2236 9924 2244
rect 9884 2156 9892 2164
rect 10236 2196 10244 2204
rect 10060 2136 10068 2144
rect 10108 2136 10116 2144
rect 9884 2116 9892 2124
rect 9868 1936 9876 1944
rect 8796 1916 8804 1924
rect 8988 1916 8996 1924
rect 9660 1896 9668 1904
rect 7900 1876 7908 1884
rect 9244 1876 9252 1884
rect 9420 1876 9428 1884
rect 9564 1876 9572 1884
rect 8572 1856 8580 1864
rect 8044 1836 8052 1844
rect 8316 1836 8324 1844
rect 8380 1756 8388 1764
rect 8140 1736 8148 1744
rect 8268 1736 8276 1744
rect 7916 1716 7924 1724
rect 7452 1516 7460 1524
rect 7596 1516 7604 1524
rect 7468 1496 7476 1504
rect 7692 1496 7700 1504
rect 7020 1456 7028 1464
rect 7244 1456 7252 1464
rect 6940 1396 6948 1404
rect 6924 1376 6932 1384
rect 7004 1376 7012 1384
rect 6348 1316 6356 1324
rect 6572 1316 6580 1324
rect 6796 1316 6804 1324
rect 7372 1376 7380 1384
rect 7036 1316 7044 1324
rect 6348 1276 6356 1284
rect 6540 1276 6548 1284
rect 6556 1276 6564 1284
rect 6796 1276 6804 1284
rect 8156 1696 8164 1704
rect 8300 1676 8308 1684
rect 8060 1656 8068 1664
rect 8460 1536 8468 1544
rect 8812 1816 8820 1824
rect 8940 1816 8948 1824
rect 8748 1756 8756 1764
rect 9132 1816 9140 1824
rect 9676 1816 9684 1824
rect 9804 1816 9812 1824
rect 8588 1736 8596 1744
rect 8748 1656 8756 1664
rect 8236 1496 8244 1504
rect 8892 1496 8900 1504
rect 9020 1756 9028 1764
rect 9436 1756 9444 1764
rect 9884 1896 9892 1904
rect 10092 1876 10100 1884
rect 10252 1836 10260 1844
rect 10220 1796 10228 1804
rect 10060 1776 10068 1784
rect 8956 1736 8964 1744
rect 9436 1736 9444 1744
rect 9228 1696 9236 1704
rect 9324 1516 9332 1524
rect 9404 1516 9412 1524
rect 8972 1476 8980 1484
rect 8988 1476 8996 1484
rect 9404 1476 9412 1484
rect 9596 1476 9604 1484
rect 7868 1456 7876 1464
rect 7660 1376 7668 1384
rect 7868 1376 7876 1384
rect 8012 1376 8020 1384
rect 7596 1336 7604 1344
rect 7596 1316 7604 1324
rect 7692 1316 7700 1324
rect 7916 1316 7924 1324
rect 7900 1296 7908 1304
rect 7596 1276 7604 1284
rect 7404 1256 7412 1264
rect 6812 1196 6820 1204
rect 6380 1136 6388 1144
rect 6620 1136 6628 1144
rect 7484 1136 7492 1144
rect 5916 1116 5924 1124
rect 5932 1116 5940 1124
rect 5948 1116 5956 1124
rect 6156 1116 6164 1124
rect 7036 1116 7044 1124
rect 7708 1116 7714 1124
rect 7714 1116 7716 1124
rect 5900 1076 5908 1084
rect 6316 1096 6324 1104
rect 6524 1096 6532 1104
rect 6956 1096 6964 1104
rect 7708 1096 7716 1104
rect 6620 1076 6628 1084
rect 7068 1056 7076 1064
rect 7244 1056 7252 1064
rect 7388 1056 7396 1064
rect 7852 1056 7860 1064
rect 6956 1036 6964 1044
rect 7212 1036 7220 1044
rect 6748 976 6756 984
rect 7452 976 7460 984
rect 6092 956 6100 964
rect 6764 956 6772 964
rect 6892 956 6900 964
rect 7132 956 7140 964
rect 5884 936 5892 944
rect 6140 936 6148 944
rect 6540 936 6548 944
rect 6556 936 6564 944
rect 7244 936 7252 944
rect 5788 916 5796 924
rect 5868 916 5876 924
rect 5212 876 5220 884
rect 5180 816 5188 824
rect 5420 816 5428 824
rect 5340 776 5348 784
rect 5100 736 5108 744
rect 5788 876 5796 884
rect 5804 796 5812 804
rect 6124 896 6132 904
rect 6284 896 6292 904
rect 7452 916 7460 924
rect 7148 896 7156 904
rect 5884 876 5892 884
rect 6092 876 6100 884
rect 4892 696 4900 704
rect 4908 696 4916 704
rect 4716 596 4724 604
rect 5132 696 5140 704
rect 5548 696 5556 704
rect 6012 696 6020 704
rect 5468 676 5476 684
rect 5084 656 5092 664
rect 5100 656 5108 664
rect 5212 656 5220 664
rect 5628 656 5636 664
rect 5852 616 5860 624
rect 6092 656 6100 664
rect 6124 656 6132 664
rect 6284 636 6292 644
rect 6044 576 6052 584
rect 5452 556 5460 564
rect 4540 536 4548 544
rect 4940 536 4948 544
rect 5260 536 5268 544
rect 5580 536 5588 544
rect 6156 536 6164 544
rect 4476 516 4484 524
rect 4364 496 4372 504
rect 4124 476 4132 484
rect 3836 336 3844 344
rect 3500 296 3508 304
rect 2860 276 2868 284
rect 2956 276 2964 284
rect 3084 276 3092 284
rect 3116 276 3124 284
rect 3308 276 3316 284
rect 3532 276 3540 284
rect 1756 256 1764 264
rect 2652 256 2660 264
rect 1628 236 1636 244
rect 2044 236 2052 244
rect 2076 236 2084 244
rect 2380 236 2388 244
rect 2572 236 2580 244
rect 2716 236 2724 244
rect 2732 236 2740 244
rect 3308 236 3316 244
rect 1548 196 1556 204
rect 1852 196 1860 204
rect 1628 156 1636 164
rect 1820 156 1828 164
rect 2044 156 2052 164
rect 1532 136 1540 144
rect 1900 136 1908 144
rect 1980 136 1988 144
rect 2444 196 2452 204
rect 2348 176 2356 184
rect 2172 156 2180 164
rect 2156 136 2164 144
rect 1212 96 1220 104
rect 1468 96 1476 104
rect 3372 216 3380 224
rect 3820 276 3828 284
rect 3708 196 3716 204
rect 3804 196 3812 204
rect 2812 156 2820 164
rect 2956 156 2964 164
rect 3180 156 3188 164
rect 4156 316 4164 324
rect 3964 296 3972 304
rect 4380 436 4388 444
rect 4460 436 4468 444
rect 4556 516 4564 524
rect 4604 436 4612 444
rect 4940 436 4948 444
rect 4940 356 4948 364
rect 4716 336 4724 344
rect 4716 316 4724 324
rect 5148 516 5156 524
rect 5148 496 5156 504
rect 5244 476 5252 484
rect 5948 516 5956 524
rect 6172 516 6180 524
rect 5788 496 5796 504
rect 5676 476 5684 484
rect 5548 456 5556 464
rect 5612 456 5620 464
rect 5708 456 5716 464
rect 5772 436 5780 444
rect 5628 356 5636 364
rect 5388 316 5396 324
rect 5628 316 5636 324
rect 4604 296 4612 304
rect 4940 296 4948 304
rect 5132 296 5140 304
rect 5404 296 5412 304
rect 4412 276 4420 284
rect 4716 276 4724 284
rect 5036 276 5044 284
rect 5180 276 5188 284
rect 5420 276 5428 284
rect 4364 176 4372 184
rect 4188 156 4196 164
rect 3692 136 3700 144
rect 3868 136 3876 144
rect 4076 136 4084 144
rect 2732 116 2740 124
rect 3404 96 3412 104
rect 3596 96 3604 104
rect 3628 96 3636 104
rect 2684 16 2692 24
rect 4092 116 4100 124
rect 4188 96 4196 104
rect 3852 76 3860 84
rect 4076 76 4084 84
rect 4044 16 4052 24
rect 4076 16 4084 24
rect 5468 236 5476 244
rect 5868 476 5876 484
rect 7244 876 7252 884
rect 6716 756 6724 764
rect 6492 736 6500 744
rect 6716 716 6724 724
rect 6700 696 6708 704
rect 7580 776 7588 784
rect 7372 756 7380 764
rect 7388 756 7396 764
rect 7020 736 7028 744
rect 6476 676 6484 684
rect 6396 556 6404 564
rect 7036 696 7044 704
rect 7372 676 7380 684
rect 6956 616 6964 624
rect 7180 556 7188 564
rect 6572 536 6580 544
rect 6620 536 6628 544
rect 7068 536 7076 544
rect 7580 596 7588 604
rect 7500 556 7508 564
rect 7276 536 7284 544
rect 7388 536 7396 544
rect 6972 516 6980 524
rect 6972 496 6980 504
rect 7692 936 7700 944
rect 8076 1016 8084 1024
rect 8444 1396 8452 1404
rect 9308 1456 9316 1464
rect 9564 1456 9572 1464
rect 8780 1436 8788 1444
rect 9180 1436 9188 1444
rect 8524 1396 8532 1404
rect 8364 1356 8372 1364
rect 8364 1316 8372 1324
rect 8348 1276 8356 1284
rect 8124 1256 8132 1264
rect 8268 1256 8276 1264
rect 8684 1256 8692 1264
rect 8236 1156 8244 1164
rect 8492 1136 8500 1144
rect 8700 1136 8708 1144
rect 8460 1076 8468 1084
rect 8284 1036 8292 1044
rect 8508 1036 8516 1044
rect 8092 996 8100 1004
rect 8300 956 8308 964
rect 7916 936 7924 944
rect 8556 956 8564 964
rect 8236 896 8244 904
rect 8556 896 8564 904
rect 7836 836 7844 844
rect 8316 836 8324 844
rect 8476 836 8484 844
rect 7660 756 7668 764
rect 8028 716 8036 724
rect 8108 716 8116 724
rect 8700 716 8708 724
rect 8716 716 8724 724
rect 8028 696 8036 704
rect 8044 696 8052 704
rect 8476 696 8484 704
rect 7692 676 7700 684
rect 7820 676 7828 684
rect 8684 676 8692 684
rect 8236 636 8244 644
rect 8332 636 8340 644
rect 8316 596 8324 604
rect 7740 576 7748 584
rect 7804 576 7812 584
rect 8092 576 8100 584
rect 8284 556 8292 564
rect 7932 536 7940 544
rect 8300 536 8308 544
rect 8460 536 8468 544
rect 8428 496 8436 504
rect 8460 496 8468 504
rect 7052 476 7060 484
rect 8124 476 8132 484
rect 6332 436 6340 444
rect 7532 436 7540 444
rect 7644 436 7652 444
rect 6636 396 6644 404
rect 5868 336 5876 344
rect 6236 336 6244 344
rect 5852 316 5860 324
rect 6076 316 6084 324
rect 6284 316 6292 324
rect 6492 316 6500 324
rect 7052 376 7060 384
rect 6284 276 6292 284
rect 6524 276 6532 284
rect 6668 276 6676 284
rect 6844 276 6852 284
rect 6076 236 6084 244
rect 6860 236 6868 244
rect 7036 236 7044 244
rect 6028 216 6036 224
rect 4620 176 4628 184
rect 4636 136 4644 144
rect 5068 156 5076 164
rect 5100 156 5108 164
rect 5548 156 5556 164
rect 5788 156 5796 164
rect 4412 116 4420 124
rect 4604 116 4612 124
rect 4876 116 4884 124
rect 4412 96 4420 104
rect 4860 96 4868 104
rect 4684 16 4692 24
rect 5100 116 5108 124
rect 5340 116 5348 124
rect 6844 216 6852 224
rect 6636 156 6644 164
rect 6012 136 6020 144
rect 6780 136 6788 144
rect 5564 116 5572 124
rect 6028 116 6036 124
rect 6908 216 6916 224
rect 7196 336 7204 344
rect 7068 316 7076 324
rect 7196 316 7204 324
rect 7292 316 7300 324
rect 7484 296 7492 304
rect 7068 276 7076 284
rect 7276 276 7284 284
rect 7244 236 7252 244
rect 7228 176 7236 184
rect 7260 176 7268 184
rect 7948 356 7956 364
rect 7708 336 7716 344
rect 8172 336 8180 344
rect 8268 336 8276 344
rect 7708 296 7716 304
rect 7948 296 7956 304
rect 8172 276 8180 284
rect 8252 276 8260 284
rect 7740 236 7748 244
rect 8108 236 8116 244
rect 7852 176 7860 184
rect 8348 176 8356 184
rect 8492 416 8500 424
rect 8716 576 8724 584
rect 8716 476 8724 484
rect 9164 1416 9172 1424
rect 9596 1396 9604 1404
rect 9740 1536 9748 1544
rect 9868 1536 9876 1544
rect 10076 1696 10084 1704
rect 9756 1516 9764 1524
rect 10060 1516 10068 1524
rect 9772 1496 9780 1504
rect 9740 1476 9748 1484
rect 9980 1496 9988 1504
rect 9820 1456 9828 1464
rect 9852 1456 9860 1464
rect 9612 1376 9620 1384
rect 8828 1336 8836 1344
rect 9132 1336 9140 1344
rect 9180 1336 9188 1344
rect 9228 1336 9236 1344
rect 9692 1336 9700 1344
rect 9868 1336 9876 1344
rect 10012 1336 10020 1344
rect 8780 1296 8788 1304
rect 8796 1296 8804 1304
rect 8924 1136 8932 1144
rect 8924 1056 8932 1064
rect 8908 956 8916 964
rect 8908 896 8916 904
rect 8892 716 8900 724
rect 8924 696 8932 704
rect 9244 1316 9252 1324
rect 9404 1296 9412 1304
rect 9676 1276 9684 1284
rect 10028 1196 10036 1204
rect 10060 1196 10068 1204
rect 9244 1156 9252 1164
rect 9916 1136 9924 1144
rect 9820 1116 9828 1124
rect 9468 1096 9476 1104
rect 9916 1076 9924 1084
rect 9148 1056 9156 1064
rect 9388 1056 9396 1064
rect 9404 1056 9412 1064
rect 9820 1056 9828 1064
rect 9260 1016 9268 1024
rect 9420 996 9428 1004
rect 9132 956 9140 964
rect 9148 956 9156 964
rect 9244 956 9252 964
rect 9580 956 9588 964
rect 9164 916 9172 924
rect 9612 956 9620 964
rect 9596 916 9604 924
rect 9820 936 9828 944
rect 9868 916 9876 924
rect 9820 896 9828 904
rect 10108 896 10116 904
rect 9900 876 9908 884
rect 9644 736 9652 744
rect 9324 716 9332 724
rect 9532 716 9540 724
rect 9836 716 9844 724
rect 9884 716 9892 724
rect 9004 676 9012 684
rect 9164 676 9172 684
rect 9532 676 9540 684
rect 8780 636 8788 644
rect 8812 636 8820 644
rect 9036 596 9044 604
rect 9148 596 9156 604
rect 9660 656 9668 664
rect 9196 616 9204 624
rect 9180 576 9188 584
rect 9564 576 9572 584
rect 9804 556 9812 564
rect 9820 536 9828 544
rect 8780 516 8788 524
rect 9356 516 9364 524
rect 9804 496 9812 504
rect 8956 436 8964 444
rect 8732 376 8740 384
rect 8924 336 8932 344
rect 8940 336 8948 344
rect 9148 336 9156 344
rect 9500 336 9508 344
rect 8700 316 8708 324
rect 9724 316 9732 324
rect 8844 276 8852 284
rect 9820 296 9828 304
rect 9884 696 9892 704
rect 9852 576 9860 584
rect 9996 536 10004 544
rect 10092 736 10100 744
rect 10188 716 10196 724
rect 10092 536 10100 544
rect 10108 516 10116 524
rect 10044 316 10052 324
rect 8924 276 8932 284
rect 9308 276 9316 284
rect 9500 276 9508 284
rect 9740 276 9748 284
rect 10012 276 10020 284
rect 10140 276 10148 284
rect 8860 256 8868 264
rect 9820 256 9828 264
rect 8652 236 8660 244
rect 8748 236 8756 244
rect 8780 236 8788 244
rect 8972 236 8980 244
rect 10028 236 10036 244
rect 8492 196 8500 204
rect 8748 196 8756 204
rect 8524 156 8532 164
rect 8636 156 8644 164
rect 7356 136 7364 144
rect 7420 136 7428 144
rect 7692 136 7700 144
rect 8028 136 8036 144
rect 8140 136 8148 144
rect 8348 136 8356 144
rect 8428 136 8436 144
rect 7516 116 7524 124
rect 7676 116 7684 124
rect 8076 116 8084 124
rect 8124 116 8132 124
rect 8940 136 8948 144
rect 9532 216 9540 224
rect 9836 216 9844 224
rect 9596 196 9604 204
rect 9148 176 9156 184
rect 9244 176 9252 184
rect 9356 176 9364 184
rect 9436 176 9444 184
rect 9884 176 9892 184
rect 9036 156 9044 164
rect 9020 136 9028 144
rect 8588 116 8596 124
rect 9484 156 9492 164
rect 9692 136 9700 144
rect 10012 136 10020 144
rect 9676 116 9684 124
rect 5548 96 5556 104
rect 5788 96 5796 104
rect 6028 96 6034 104
rect 6034 96 6036 104
rect 8588 96 8596 104
rect 8748 96 8756 104
rect 9196 96 9204 104
rect 9468 96 9474 104
rect 9474 96 9476 104
rect 10012 96 10020 104
rect 6012 76 6020 84
rect 6236 76 6244 84
rect 5148 16 5156 24
rect 7356 16 7364 24
<< metal3 >>
rect 3588 7617 3612 7623
rect 5172 7617 5180 7623
rect 1780 7597 1820 7603
rect 6093 7564 6099 7576
rect 3364 7537 3388 7543
rect 3396 7537 4268 7543
rect 4612 7537 5020 7543
rect 5028 7537 6172 7543
rect 6180 7537 6188 7543
rect 9284 7537 9644 7543
rect 564 7517 572 7523
rect 1108 7517 1116 7523
rect 1444 7517 1452 7523
rect 2532 7517 2588 7523
rect 2724 7517 2732 7523
rect 3940 7517 4220 7523
rect 4356 7517 4812 7523
rect 5300 7517 5404 7523
rect 5412 7517 6380 7523
rect 6596 7517 6611 7523
rect 7060 7517 7756 7523
rect 317 7504 323 7516
rect 8413 7504 8419 7523
rect 8628 7517 8844 7523
rect 9252 7517 9820 7523
rect 9917 7504 9923 7523
rect 2804 7497 3484 7503
rect 3492 7497 3708 7503
rect 5844 7497 5852 7503
rect 5860 7497 7548 7503
rect 7556 7497 7676 7503
rect 8212 7497 8220 7503
rect 9492 7497 9500 7503
rect 9556 7497 9708 7503
rect 308 7477 316 7483
rect 532 7477 556 7483
rect 756 7477 1228 7483
rect 1700 7477 1708 7483
rect 2276 7477 2476 7483
rect 2500 7477 2524 7483
rect 3460 7477 3708 7483
rect 3716 7477 3916 7483
rect 4132 7477 4147 7483
rect 4276 7477 4380 7483
rect 4388 7477 4396 7483
rect 5316 7477 5356 7483
rect 5972 7477 6860 7483
rect 6868 7477 7004 7483
rect 7444 7477 7452 7483
rect 8445 7477 8460 7483
rect 8740 7477 8748 7483
rect 8852 7477 8860 7483
rect 9188 7477 9836 7483
rect 9933 7477 9948 7483
rect 7101 7464 7107 7476
rect 1220 7457 1836 7463
rect 2964 7457 3036 7463
rect 3860 7457 3948 7463
rect 3956 7457 4540 7463
rect 4548 7457 4604 7463
rect 4852 7457 6012 7463
rect 8212 7457 9180 7463
rect 9284 7457 9292 7463
rect 9316 7457 9500 7463
rect 1124 7437 2524 7443
rect 2532 7437 2732 7443
rect 3476 7437 3500 7443
rect 5844 7437 7036 7443
rect 8772 7437 9596 7443
rect 9604 7437 10060 7443
rect 292 7417 316 7423
rect 916 7417 940 7423
rect 4276 7417 4460 7423
rect 5508 7417 5580 7423
rect 580 7397 668 7403
rect 2724 7397 3116 7403
rect 5092 7397 5132 7403
rect 5364 7397 6028 7403
rect 6036 7397 7068 7403
rect 7076 7397 7884 7403
rect 7988 7397 8300 7403
rect 8324 7397 8732 7403
rect 68 7377 76 7383
rect 100 7377 508 7383
rect 877 7377 2236 7383
rect 877 7364 883 7377
rect 5668 7377 5836 7383
rect 5860 7377 6236 7383
rect 6244 7377 6492 7383
rect 6660 7377 7180 7383
rect 7540 7377 7548 7383
rect 7796 7377 7820 7383
rect 7844 7377 8060 7383
rect 10276 7377 10339 7383
rect 1092 7357 1340 7363
rect 1780 7357 2012 7363
rect 2436 7357 3644 7363
rect 3652 7357 3836 7363
rect 4212 7357 4732 7363
rect 5332 7357 5340 7363
rect 5348 7357 6140 7363
rect 6500 7357 8044 7363
rect 8052 7357 8268 7363
rect 8276 7357 8284 7363
rect 8356 7357 9580 7363
rect 308 7337 316 7343
rect 324 7337 428 7343
rect 644 7337 652 7343
rect 2756 7337 2764 7343
rect 3092 7337 3100 7343
rect 3380 7337 4204 7343
rect 4852 7337 4860 7343
rect 5188 7337 5548 7343
rect 5556 7337 5564 7343
rect 5796 7337 7452 7343
rect 7780 7337 7795 7343
rect 7892 7337 9708 7343
rect 1869 7324 1875 7336
rect 4653 7324 4659 7336
rect 196 7317 1852 7323
rect 2452 7317 3324 7323
rect 3332 7317 3340 7323
rect 3620 7317 3628 7323
rect 4100 7317 4204 7323
rect 5172 7317 5852 7323
rect 5876 7317 6124 7323
rect 6148 7317 7468 7323
rect 7476 7317 7484 7323
rect 8180 7317 8492 7323
rect 8564 7317 8572 7323
rect 8596 7317 9052 7323
rect 9620 7317 9916 7323
rect 10276 7317 10339 7323
rect 660 7297 1084 7303
rect 1316 7297 1324 7303
rect 1556 7297 1564 7303
rect 1860 7297 2492 7303
rect 2500 7297 3228 7303
rect 3236 7297 4444 7303
rect 4452 7297 4460 7303
rect 4660 7297 4844 7303
rect 4932 7297 5180 7303
rect 5780 7297 5788 7303
rect 5892 7297 5900 7303
rect 6132 7297 6172 7303
rect 6180 7297 6316 7303
rect 6356 7297 6364 7303
rect 6388 7297 6572 7303
rect 6820 7297 8044 7303
rect 8052 7297 8060 7303
rect 8484 7297 8492 7303
rect 8500 7297 9036 7303
rect 9620 7297 9644 7303
rect 9924 7297 9932 7303
rect 5581 7284 5587 7296
rect 276 7277 1244 7283
rect 1316 7277 1548 7283
rect 1556 7277 1580 7283
rect 1588 7277 1628 7283
rect 1988 7277 2012 7283
rect 2660 7277 2716 7283
rect 2756 7277 3516 7283
rect 3524 7277 3980 7283
rect 4228 7277 4972 7283
rect 5860 7277 5900 7283
rect 5908 7277 6588 7283
rect 6596 7277 6604 7283
rect 6964 7277 7468 7283
rect 7476 7277 7964 7283
rect 884 7257 892 7263
rect 3108 7257 3116 7263
rect 4404 7257 4604 7263
rect 4612 7257 4956 7263
rect 4964 7257 4988 7263
rect 1652 7197 1660 7203
rect 8100 7177 8268 7183
rect 3620 7157 5228 7163
rect 8276 7157 8412 7163
rect 772 7137 780 7143
rect 1108 7137 2732 7143
rect 4260 7137 4876 7143
rect 5220 7137 6572 7143
rect 7188 7137 7388 7143
rect 8020 7137 8636 7143
rect 269 7123 275 7136
rect 269 7117 284 7123
rect 436 7117 1628 7123
rect 1636 7117 1644 7123
rect 1652 7117 2556 7123
rect 2564 7117 2620 7123
rect 2628 7117 2636 7123
rect 2772 7117 2796 7123
rect 3700 7117 3708 7123
rect 3764 7117 3772 7123
rect 4548 7117 4556 7123
rect 4564 7117 4892 7123
rect 4980 7117 4988 7123
rect 5220 7117 5228 7123
rect 5780 7117 6012 7123
rect 6132 7117 6172 7123
rect 6932 7117 6940 7123
rect 6948 7117 7164 7123
rect 7460 7117 7484 7123
rect 7620 7117 7708 7123
rect 7956 7117 8828 7123
rect 8861 7117 8876 7123
rect 9060 7117 9212 7123
rect 9860 7117 9868 7123
rect 692 7097 764 7103
rect 948 7097 1068 7103
rect 1092 7097 1100 7103
rect 1124 7097 1132 7103
rect 1156 7097 1420 7103
rect 1444 7097 1532 7103
rect 1572 7097 2332 7103
rect 2340 7097 3372 7103
rect 3396 7097 3468 7103
rect 3876 7097 4540 7103
rect 4820 7097 4988 7103
rect 6340 7097 6588 7103
rect 7124 7097 7164 7103
rect 7172 7097 7948 7103
rect 8036 7097 8172 7103
rect 8404 7097 8604 7103
rect 8644 7097 9436 7103
rect 644 7077 652 7083
rect 660 7077 2108 7083
rect 2244 7077 2252 7083
rect 2340 7077 2348 7083
rect 3028 7077 3036 7083
rect 3092 7077 3100 7083
rect 3348 7077 4316 7083
rect 4484 7077 4876 7083
rect 4884 7077 5132 7083
rect 5236 7077 5244 7083
rect 5460 7077 5468 7083
rect 6020 7077 7100 7083
rect 7252 7077 7340 7083
rect 7556 7077 8636 7083
rect 8884 7077 8892 7083
rect 8948 7077 9436 7083
rect 212 7057 1308 7063
rect 1316 7057 1644 7063
rect 1652 7057 2444 7063
rect 2740 7057 3532 7063
rect 3540 7057 3692 7063
rect 3876 7057 4012 7063
rect 4100 7057 4115 7063
rect 4468 7057 5372 7063
rect 5380 7057 5388 7063
rect 5796 7057 5884 7063
rect 5892 7057 6124 7063
rect 6964 7057 7868 7063
rect 9428 7057 9628 7063
rect 788 7037 956 7043
rect 1124 7037 1244 7043
rect 1796 7037 1804 7043
rect 2116 7037 3116 7043
rect 3124 7037 3980 7043
rect 3988 7037 4732 7043
rect 4740 7037 4748 7043
rect 6788 7037 7500 7043
rect 9684 7037 9692 7043
rect 1876 7017 1884 7023
rect 2596 7017 3884 7023
rect 7380 7017 9132 7023
rect 2260 6997 2284 7003
rect 3028 6997 3340 7003
rect 5796 6997 6012 7003
rect 9652 6997 10236 7003
rect 221 6977 268 6983
rect 221 6963 227 6977
rect 660 6977 684 6983
rect 2468 6977 2924 6983
rect 4420 6977 4444 6983
rect 212 6957 227 6963
rect 548 6957 668 6963
rect 2100 6957 4204 6963
rect 4564 6957 4604 6963
rect 6612 6957 6780 6963
rect 7204 6957 7468 6963
rect 7684 6957 7692 6963
rect 7972 6957 9436 6963
rect 9444 6957 9452 6963
rect 9652 6957 9884 6963
rect 884 6937 892 6943
rect 980 6937 1324 6943
rect 1860 6937 1868 6943
rect 2644 6937 2652 6943
rect 3316 6937 4236 6943
rect 4324 6937 4332 6943
rect 4548 6937 4828 6943
rect 4996 6937 5068 6943
rect 5076 6937 5084 6943
rect 5412 6937 5420 6943
rect 5908 6937 5980 6943
rect 6228 6937 6268 6943
rect 6292 6937 6540 6943
rect 6548 6937 6668 6943
rect 7012 6937 7228 6943
rect 7236 6937 7244 6943
rect 7476 6937 7644 6943
rect 7652 6937 8012 6943
rect 8116 6937 8588 6943
rect 8804 6937 8819 6943
rect 2973 6924 2979 6936
rect 884 6917 2284 6923
rect 2356 6917 2732 6923
rect 2941 6917 2956 6923
rect 3508 6917 4076 6923
rect 4612 6917 4620 6923
rect 4980 6917 5052 6923
rect 5060 6917 5196 6923
rect 6276 6917 7004 6923
rect 7012 6917 7212 6923
rect 7220 6917 8396 6923
rect 8813 6923 8819 6937
rect 8836 6937 8908 6943
rect 8916 6937 9100 6943
rect 9524 6937 9532 6943
rect 9668 6937 9676 6943
rect 8813 6917 8860 6923
rect 9380 6917 10108 6923
rect 436 6897 444 6903
rect 1188 6897 1628 6903
rect 2436 6897 2748 6903
rect 3316 6897 3484 6903
rect 3764 6897 3788 6903
rect 3988 6897 3996 6903
rect 4004 6897 4028 6903
rect 4084 6897 4844 6903
rect 5188 6897 5996 6903
rect 6004 6897 6012 6903
rect 6212 6897 6227 6903
rect 6685 6897 6956 6903
rect 509 6884 515 6896
rect 973 6884 979 6896
rect 1181 6884 1187 6896
rect 2077 6884 2083 6896
rect 3309 6884 3315 6896
rect 4877 6884 4883 6896
rect 6317 6884 6323 6896
rect 6685 6884 6691 6897
rect 7412 6897 7564 6903
rect 7780 6897 7788 6903
rect 7828 6897 8012 6903
rect 8020 6897 8108 6903
rect 8116 6897 9372 6903
rect 9380 6897 9692 6903
rect 9700 6897 9724 6903
rect 2084 6877 2956 6883
rect 4228 6877 4876 6883
rect 6996 6877 9116 6883
rect 9332 6877 9340 6883
rect 9444 6877 9452 6883
rect 9508 6877 9660 6883
rect 2420 6857 3164 6863
rect 3540 6857 3548 6863
rect 3780 6857 3788 6863
rect 6308 6857 6364 6863
rect 8676 6857 8684 6863
rect 1332 6837 1340 6843
rect 4196 6837 4204 6843
rect 8349 6837 8508 6843
rect 4269 6824 4275 6836
rect 4701 6824 4707 6836
rect 4941 6824 4947 6836
rect 8349 6823 8355 6837
rect 8276 6817 8355 6823
rect 2580 6777 2636 6783
rect 1860 6757 1884 6763
rect 2932 6757 2940 6763
rect 5044 6757 5052 6763
rect 5764 6757 5772 6763
rect 1620 6737 1900 6743
rect 1908 6737 2364 6743
rect 2372 6737 2380 6743
rect 2676 6737 2684 6743
rect 2724 6737 3244 6743
rect 3988 6737 4044 6743
rect 4052 6737 4412 6743
rect 5092 6737 5260 6743
rect 5412 6737 6172 6743
rect 6180 6737 6732 6743
rect 9540 6737 9564 6743
rect 77 6724 83 6736
rect 7501 6724 7507 6736
rect 516 6717 1212 6723
rect 1636 6717 2716 6723
rect 3172 6717 3180 6723
rect 3476 6717 3484 6723
rect 3828 6717 3836 6723
rect 4244 6717 4508 6723
rect 4692 6717 4748 6723
rect 4756 6717 4771 6723
rect 5476 6717 6844 6723
rect 6852 6717 7100 6723
rect 7236 6717 7292 6723
rect 7300 6717 7308 6723
rect 7492 6717 7500 6723
rect 7716 6717 7740 6723
rect 8580 6717 8588 6723
rect 8916 6717 9068 6723
rect 9364 6717 9372 6723
rect 9572 6717 9660 6723
rect 9876 6717 10252 6723
rect 532 6697 972 6703
rect 1133 6697 1148 6703
rect 1668 6697 1932 6703
rect 2756 6697 4060 6703
rect 4068 6697 4588 6703
rect 5604 6697 5820 6703
rect 5860 6697 5868 6703
rect 5876 6697 6188 6703
rect 6196 6697 6332 6703
rect 6500 6697 9004 6703
rect 9012 6697 9900 6703
rect 564 6677 684 6683
rect 756 6677 764 6683
rect 1124 6677 1132 6683
rect 1252 6677 1308 6683
rect 1812 6677 2076 6683
rect 2292 6677 2364 6683
rect 2372 6677 2796 6683
rect 2836 6677 3132 6683
rect 3460 6677 3484 6683
rect 4052 6677 4060 6683
rect 4260 6677 4268 6683
rect 4484 6677 4492 6683
rect 5044 6677 5084 6683
rect 5092 6677 5228 6683
rect 5236 6677 5276 6683
rect 5540 6677 5564 6683
rect 5572 6677 5628 6683
rect 6068 6677 6076 6683
rect 6084 6677 7820 6683
rect 7940 6677 8092 6683
rect 8564 6677 8572 6683
rect 8884 6677 9020 6683
rect 9204 6677 9340 6683
rect 9668 6677 9836 6683
rect 8461 6664 8467 6676
rect 9021 6664 9027 6676
rect 100 6657 108 6663
rect 692 6657 2428 6663
rect 2980 6657 4588 6663
rect 5572 6657 5612 6663
rect 6036 6657 6156 6663
rect 6164 6657 6172 6663
rect 6276 6657 6284 6663
rect 6628 6657 7116 6663
rect 7284 6657 7292 6663
rect 7668 6657 7683 6663
rect 7700 6657 7724 6663
rect 7876 6657 7916 6663
rect 9060 6657 9676 6663
rect 1652 6637 1660 6643
rect 1764 6637 1852 6643
rect 2516 6637 2828 6643
rect 3492 6637 3676 6643
rect 4020 6637 4060 6643
rect 5220 6637 5324 6643
rect 5332 6637 5436 6643
rect 5444 6637 5788 6643
rect 6836 6637 6860 6643
rect 6980 6637 7068 6643
rect 8788 6637 9388 6643
rect 4349 6624 4355 6636
rect 116 6617 268 6623
rect 1396 6617 1436 6623
rect 2500 6617 2668 6623
rect 7796 6617 8060 6623
rect 9572 6617 9804 6623
rect 308 6597 668 6603
rect 756 6597 1116 6603
rect 2116 6597 2716 6603
rect 3108 6597 4044 6603
rect 4884 6597 5404 6603
rect 5636 6597 5772 6603
rect 6093 6603 6099 6616
rect 6093 6597 6300 6603
rect 6308 6597 6476 6603
rect 6484 6597 6492 6603
rect 7044 6597 7180 6603
rect 7524 6597 7836 6603
rect 8788 6597 8796 6603
rect 1092 6577 1100 6583
rect 1940 6577 1948 6583
rect 2068 6577 2220 6583
rect 2276 6577 2892 6583
rect 3556 6577 3612 6583
rect 3796 6577 3820 6583
rect 6756 6577 7164 6583
rect 7684 6577 7740 6583
rect 8772 6577 8908 6583
rect 212 6557 300 6563
rect 692 6557 972 6563
rect 980 6557 1324 6563
rect 1332 6557 2412 6563
rect 2644 6557 2844 6563
rect 2852 6557 4716 6563
rect 5700 6557 5708 6563
rect 6164 6557 6268 6563
rect 6276 6557 6364 6563
rect 6964 6557 7356 6563
rect 7860 6557 7948 6563
rect 7972 6557 9564 6563
rect 9844 6557 10124 6563
rect 4829 6544 4835 6556
rect 644 6537 1660 6543
rect 1796 6537 1852 6543
rect 2404 6537 2412 6543
rect 2420 6537 2620 6543
rect 2628 6537 2748 6543
rect 2804 6537 2812 6543
rect 3092 6537 3100 6543
rect 3252 6537 3260 6543
rect 3412 6537 3420 6543
rect 3588 6537 3740 6543
rect 4340 6537 4380 6543
rect 4484 6537 4828 6543
rect 5284 6537 5292 6543
rect 5572 6537 5884 6543
rect 6116 6537 6172 6543
rect 6916 6537 7020 6543
rect 7140 6537 7148 6543
rect 7556 6537 7596 6543
rect 7796 6537 7804 6543
rect 7860 6537 8044 6543
rect 8228 6537 8236 6543
rect 8260 6537 8268 6543
rect 8276 6537 9116 6543
rect 9188 6537 9212 6543
rect 3965 6524 3971 6536
rect 9677 6524 9683 6536
rect 10013 6524 10019 6536
rect 852 6517 876 6523
rect 1316 6517 1324 6523
rect 1380 6517 1516 6523
rect 1540 6517 1996 6523
rect 2004 6517 3180 6523
rect 3188 6517 3964 6523
rect 4932 6517 5868 6523
rect 5892 6517 6572 6523
rect 6580 6517 6588 6523
rect 7380 6517 7900 6523
rect 7908 6517 9132 6523
rect 84 6497 636 6503
rect 644 6497 668 6503
rect 964 6497 1628 6503
rect 1860 6497 1900 6503
rect 2084 6497 2108 6503
rect 2436 6497 2636 6503
rect 2660 6497 4172 6503
rect 4340 6497 4396 6503
rect 4404 6497 4444 6503
rect 4500 6497 4524 6503
rect 4532 6497 4556 6503
rect 4900 6497 5532 6503
rect 5764 6497 5779 6503
rect 6020 6497 6076 6503
rect 6100 6497 6332 6503
rect 6340 6497 6348 6503
rect 6580 6497 6604 6503
rect 7364 6497 7372 6503
rect 7444 6497 7852 6503
rect 7876 6497 8252 6503
rect 8356 6497 8364 6503
rect 8548 6497 8556 6503
rect 8772 6497 8796 6503
rect 9620 6497 9660 6503
rect 9908 6497 10044 6503
rect 1300 6477 2844 6483
rect 2852 6477 2860 6483
rect 3252 6477 3804 6483
rect 3812 6477 5084 6483
rect 7172 6477 7596 6483
rect 7604 6477 7612 6483
rect 7876 6477 8140 6483
rect 8260 6477 10012 6483
rect 3972 6457 3980 6463
rect 7492 6457 9820 6463
rect 6772 6437 7500 6443
rect 7508 6437 9436 6443
rect 8820 6377 8988 6383
rect 4532 6357 4908 6363
rect 6356 6357 6364 6363
rect 8484 6357 8572 6363
rect 8580 6357 9420 6363
rect 9796 6357 9868 6363
rect 1108 6337 1420 6343
rect 1428 6337 3180 6343
rect 3636 6337 3820 6343
rect 4052 6337 4060 6343
rect 4196 6337 4316 6343
rect 4324 6337 4492 6343
rect 4628 6337 4636 6343
rect 4996 6337 5020 6343
rect 5220 6337 5372 6343
rect 5524 6337 5532 6343
rect 5604 6337 6012 6343
rect 6372 6337 6588 6343
rect 6756 6337 6812 6343
rect 8260 6337 9148 6343
rect 100 6317 108 6323
rect 676 6317 684 6323
rect 900 6317 924 6323
rect 1348 6317 1532 6323
rect 1636 6317 2492 6323
rect 2500 6317 2780 6323
rect 2916 6317 2940 6323
rect 3236 6317 3244 6323
rect 3540 6317 3548 6323
rect 3780 6317 5020 6323
rect 5300 6317 5820 6323
rect 5828 6317 5836 6323
rect 5892 6317 5900 6323
rect 6132 6317 7036 6323
rect 8036 6317 8316 6323
rect 8484 6317 9356 6323
rect 9668 6317 10220 6323
rect 6125 6304 6131 6316
rect 308 6297 444 6303
rect 2468 6297 2492 6303
rect 2804 6297 4348 6303
rect 4516 6297 4684 6303
rect 4692 6297 4940 6303
rect 5028 6297 5452 6303
rect 5492 6297 5900 6303
rect 6596 6297 7276 6303
rect 7988 6297 8908 6303
rect 8916 6297 9404 6303
rect 9716 6297 10220 6303
rect 436 6277 652 6283
rect 660 6277 2556 6283
rect 2772 6277 2924 6283
rect 2932 6277 3020 6283
rect 3572 6277 4236 6283
rect 4660 6277 4684 6283
rect 4692 6277 5596 6283
rect 5876 6277 6476 6283
rect 6484 6277 6604 6283
rect 7012 6277 7027 6283
rect 7044 6277 7052 6283
rect 7060 6277 7084 6283
rect 7220 6277 7804 6283
rect 8020 6277 8035 6283
rect 8436 6277 8451 6283
rect 9028 6277 9164 6283
rect 9364 6277 9372 6283
rect 9476 6277 9596 6283
rect 9844 6277 10076 6283
rect 8909 6264 8915 6276
rect 468 6257 524 6263
rect 1124 6257 1427 6263
rect 228 6237 236 6243
rect 1421 6243 1427 6257
rect 1444 6257 1452 6263
rect 1620 6257 1660 6263
rect 1892 6257 2044 6263
rect 2692 6257 2700 6263
rect 3124 6257 3452 6263
rect 3812 6257 3820 6263
rect 4020 6257 4044 6263
rect 4244 6257 4476 6263
rect 4916 6257 4940 6263
rect 4964 6257 5180 6263
rect 5396 6257 5804 6263
rect 6084 6257 6108 6263
rect 6116 6257 6140 6263
rect 6244 6257 6252 6263
rect 6372 6257 6604 6263
rect 6788 6257 7372 6263
rect 8068 6257 8835 6263
rect 1421 6237 1564 6243
rect 1604 6237 1612 6243
rect 1908 6237 2508 6243
rect 4020 6237 4332 6243
rect 5812 6237 5916 6243
rect 8020 6237 8076 6243
rect 8548 6237 8556 6243
rect 8564 6237 8716 6243
rect 8772 6237 8812 6243
rect 8829 6243 8835 6257
rect 9828 6257 9836 6263
rect 8829 6237 9820 6243
rect 116 6217 236 6223
rect 660 6217 1996 6223
rect 4068 6217 4124 6223
rect 7252 6217 7452 6223
rect 7860 6217 9164 6223
rect 84 6197 92 6203
rect 1092 6197 1324 6203
rect 1476 6197 1548 6203
rect 2260 6197 2444 6203
rect 2724 6197 2908 6203
rect 4916 6197 4972 6203
rect 9652 6197 9676 6203
rect 9789 6203 9795 6216
rect 9789 6197 10028 6203
rect 852 6177 940 6183
rect 1140 6177 1164 6183
rect 1261 6177 1836 6183
rect 1261 6163 1267 6177
rect 2644 6177 3420 6183
rect 4708 6177 4812 6183
rect 5220 6177 5276 6183
rect 7364 6177 7404 6183
rect 7636 6177 7676 6183
rect 10020 6177 10044 6183
rect 884 6157 1267 6163
rect 1300 6157 2156 6163
rect 2212 6157 3587 6163
rect 877 6144 883 6156
rect 212 6137 476 6143
rect 500 6137 636 6143
rect 1604 6137 1628 6143
rect 1748 6137 1756 6143
rect 1780 6137 2460 6143
rect 2500 6137 2844 6143
rect 3581 6143 3587 6157
rect 3764 6157 4572 6163
rect 4580 6157 5100 6163
rect 5668 6157 5820 6163
rect 6004 6157 6028 6163
rect 6340 6157 6364 6163
rect 6868 6157 6924 6163
rect 7124 6157 8108 6163
rect 9524 6157 9532 6163
rect 3581 6137 3852 6143
rect 3860 6137 3948 6143
rect 3972 6137 3980 6143
rect 3988 6137 4316 6143
rect 4324 6137 4620 6143
rect 4788 6137 4796 6143
rect 5236 6137 5436 6143
rect 6068 6137 6236 6143
rect 6244 6137 6380 6143
rect 6564 6137 6796 6143
rect 7140 6137 7148 6143
rect 7428 6137 7852 6143
rect 8564 6137 8652 6143
rect 8996 6137 9004 6143
rect 9220 6137 9228 6143
rect 9348 6137 9756 6143
rect 10084 6137 10204 6143
rect 1092 6117 1132 6123
rect 1316 6117 2524 6123
rect 3604 6117 3980 6123
rect 3988 6117 3996 6123
rect 4004 6117 5676 6123
rect 5748 6117 6572 6123
rect 6612 6117 7148 6123
rect 7156 6117 7180 6123
rect 7588 6117 7644 6123
rect 7684 6117 7692 6123
rect 7885 6123 7891 6136
rect 8333 6124 8339 6136
rect 7700 6117 7891 6123
rect 8900 6117 9164 6123
rect 9172 6117 9884 6123
rect 9892 6117 9916 6123
rect 468 6097 524 6103
rect 660 6097 1180 6103
rect 1412 6097 1612 6103
rect 1636 6097 1644 6103
rect 1988 6097 1996 6103
rect 2308 6097 2332 6103
rect 2468 6097 2892 6103
rect 2980 6097 2988 6103
rect 653 6084 659 6096
rect 3101 6084 3107 6103
rect 3316 6097 3324 6103
rect 3556 6097 3772 6103
rect 3780 6097 4300 6103
rect 4308 6097 4508 6103
rect 4541 6097 4556 6103
rect 4756 6097 4764 6103
rect 5012 6097 5404 6103
rect 6020 6097 6156 6103
rect 6260 6097 7020 6103
rect 7220 6097 7235 6103
rect 7229 6084 7235 6097
rect 8676 6097 8892 6103
rect 9012 6097 9372 6103
rect 8013 6084 8019 6096
rect 884 6077 892 6083
rect 980 6077 1100 6083
rect 1108 6077 1308 6083
rect 1972 6077 2204 6083
rect 3572 6077 3740 6083
rect 3748 6077 4268 6083
rect 4276 6077 4492 6083
rect 4500 6077 4924 6083
rect 5588 6077 5836 6083
rect 5844 6077 6604 6083
rect 6692 6077 6924 6083
rect 9188 6077 9340 6083
rect 9876 6077 9884 6083
rect 2308 6057 2316 6063
rect 2932 6057 5004 6063
rect 5236 6057 5244 6063
rect 5636 6057 6332 6063
rect 6340 6057 6348 6063
rect 8116 6057 8124 6063
rect 2205 6044 2211 6056
rect 6781 6044 6787 6056
rect 564 6037 732 6043
rect 4100 6037 4108 6043
rect 5412 6037 5628 6043
rect 8996 5997 9004 6003
rect 5261 5984 5267 5996
rect 9268 5977 9388 5983
rect 452 5957 556 5963
rect 2948 5957 3612 5963
rect 644 5937 764 5943
rect 1124 5937 1580 5943
rect 1588 5937 2428 5943
rect 2532 5937 2988 5943
rect 4660 5937 5036 5943
rect 5428 5937 5724 5943
rect 5732 5937 6124 5943
rect 6468 5937 6476 5943
rect 7860 5937 7948 5943
rect 765 5924 771 5936
rect 9037 5924 9043 5936
rect 1652 5917 1948 5923
rect 1956 5917 2716 5923
rect 2724 5917 2732 5923
rect 3364 5917 4044 5923
rect 4820 5917 4940 5923
rect 4996 5917 5228 5923
rect 5508 5917 5516 5923
rect 5956 5917 6076 5923
rect 6084 5917 6108 5923
rect 6308 5917 6316 5923
rect 6324 5917 6492 5923
rect 6564 5917 7292 5923
rect 7300 5917 8524 5923
rect 8532 5917 8540 5923
rect 8580 5917 8604 5923
rect 8708 5917 8716 5923
rect 9604 5917 9692 5923
rect 4253 5904 4259 5916
rect 676 5897 716 5903
rect 724 5897 780 5903
rect 2020 5897 2028 5903
rect 2516 5897 2700 5903
rect 3364 5897 3580 5903
rect 5012 5897 5724 5903
rect 5732 5897 5788 5903
rect 6548 5897 7020 5903
rect 7028 5897 7948 5903
rect 7956 5897 7980 5903
rect 8052 5897 8156 5903
rect 8804 5897 9260 5903
rect 6541 5884 6547 5896
rect 212 5877 236 5883
rect 868 5877 876 5883
rect 1348 5877 3020 5883
rect 3188 5877 3324 5883
rect 3588 5877 3596 5883
rect 3796 5877 4236 5883
rect 4244 5877 4252 5883
rect 4484 5877 4732 5883
rect 5364 5877 5388 5883
rect 5412 5877 6316 5883
rect 6324 5877 6428 5883
rect 6756 5877 6771 5883
rect 6820 5877 6844 5883
rect 7156 5877 7308 5883
rect 7316 5877 8268 5883
rect 8292 5877 8940 5883
rect 8948 5877 8956 5883
rect 9252 5877 9484 5883
rect 9684 5877 9900 5883
rect 3021 5864 3027 5876
rect 228 5857 1388 5863
rect 1812 5857 2284 5863
rect 2500 5857 2524 5863
rect 3028 5857 3964 5863
rect 4692 5857 4700 5863
rect 5492 5857 5500 5863
rect 5508 5857 5580 5863
rect 6164 5857 6332 5863
rect 6468 5857 7084 5863
rect 7092 5857 7660 5863
rect 7700 5857 7788 5863
rect 7892 5857 8508 5863
rect 8516 5857 8524 5863
rect 9172 5857 9692 5863
rect 2292 5837 4284 5843
rect 5892 5837 7868 5843
rect 2356 5817 4492 5823
rect 6868 5817 6972 5823
rect 7428 5817 7516 5823
rect 7732 5817 7740 5823
rect 7940 5817 8012 5823
rect 3156 5797 3164 5803
rect 3604 5797 3660 5803
rect 4692 5797 4716 5803
rect 8132 5797 8364 5803
rect 8484 5797 8492 5803
rect 9588 5797 10044 5803
rect 2781 5784 2787 5796
rect 708 5777 972 5783
rect 1108 5777 1116 5783
rect 1684 5777 2716 5783
rect 3396 5777 3452 5783
rect 3844 5777 4924 5783
rect 6820 5777 6924 5783
rect 7188 5777 7196 5783
rect 8324 5777 8348 5783
rect 8820 5777 9180 5783
rect 9812 5777 9836 5783
rect 308 5757 316 5763
rect 1636 5757 1884 5763
rect 2356 5757 2364 5763
rect 2372 5757 2476 5763
rect 2756 5757 2908 5763
rect 3028 5757 3052 5763
rect 3188 5757 3580 5763
rect 3588 5757 4508 5763
rect 4516 5757 4908 5763
rect 5684 5757 5692 5763
rect 6356 5757 6492 5763
rect 6772 5757 7740 5763
rect 196 5737 1116 5743
rect 1364 5737 1420 5743
rect 1636 5737 1660 5743
rect 2532 5737 2956 5743
rect 2964 5737 3916 5743
rect 3924 5737 4108 5743
rect 4228 5737 4236 5743
rect 4372 5737 4796 5743
rect 4804 5737 4812 5743
rect 5236 5737 5244 5743
rect 5252 5737 5484 5743
rect 5524 5737 5580 5743
rect 5588 5737 5932 5743
rect 6372 5737 6604 5743
rect 6836 5737 6844 5743
rect 6932 5737 7500 5743
rect 7924 5737 8060 5743
rect 8148 5737 8163 5743
rect 9124 5737 9436 5743
rect 9444 5737 9484 5743
rect 9700 5737 9724 5743
rect 9901 5724 9907 5743
rect 500 5717 652 5723
rect 1204 5717 1212 5723
rect 1380 5717 3036 5723
rect 3060 5717 3180 5723
rect 3204 5717 3372 5723
rect 3652 5717 3788 5723
rect 4052 5717 4076 5723
rect 4084 5717 4572 5723
rect 4932 5717 5164 5723
rect 5348 5717 5452 5723
rect 5460 5717 5468 5723
rect 5924 5717 6364 5723
rect 6500 5717 7148 5723
rect 7156 5717 7276 5723
rect 7508 5717 9372 5723
rect 9380 5717 9852 5723
rect 205 5704 211 5716
rect 1085 5704 1091 5716
rect 9885 5704 9891 5716
rect 212 5697 1004 5703
rect 1364 5697 1900 5703
rect 2116 5697 2124 5703
rect 2340 5697 2348 5703
rect 2564 5697 3564 5703
rect 3588 5697 3596 5703
rect 3604 5697 4556 5703
rect 4564 5697 4572 5703
rect 4628 5697 5132 5703
rect 5364 5697 5388 5703
rect 5908 5697 6108 5703
rect 6132 5697 6492 5703
rect 6500 5697 6508 5703
rect 6820 5697 6828 5703
rect 6964 5697 7020 5703
rect 7284 5697 7292 5703
rect 7492 5697 7500 5703
rect 8676 5697 9372 5703
rect 9380 5697 9388 5703
rect 9460 5697 9468 5703
rect 9476 5697 9500 5703
rect 9700 5697 9708 5703
rect 8093 5684 8099 5696
rect 8509 5684 8515 5696
rect 420 5677 428 5683
rect 436 5677 508 5683
rect 516 5677 1804 5683
rect 1892 5677 2780 5683
rect 3892 5677 4332 5683
rect 4356 5677 4476 5683
rect 4676 5677 4780 5683
rect 4788 5677 4796 5683
rect 5277 5677 6588 5683
rect 660 5657 940 5663
rect 948 5657 1116 5663
rect 1428 5657 1468 5663
rect 1652 5657 1676 5663
rect 2580 5657 3004 5663
rect 3492 5657 3644 5663
rect 5277 5663 5283 5677
rect 6596 5677 7404 5683
rect 8820 5677 9692 5683
rect 9700 5677 10220 5683
rect 4340 5657 5283 5663
rect 5700 5657 5708 5663
rect 2516 5637 2572 5643
rect 2676 5637 2700 5643
rect 2756 5637 3900 5643
rect 3908 5637 4092 5643
rect 4925 5624 4931 5643
rect 2580 5617 3836 5623
rect 3796 5597 3804 5603
rect 3236 5577 4204 5583
rect 1220 5557 1676 5563
rect 1684 5557 2828 5563
rect 3396 5557 3420 5563
rect 7716 5557 8092 5563
rect 8100 5557 8700 5563
rect 68 5537 220 5543
rect 996 5537 1068 5543
rect 3172 5537 3180 5543
rect 3316 5537 3468 5543
rect 3476 5537 4716 5543
rect 5412 5537 5420 5543
rect 6052 5537 6060 5543
rect 6372 5537 6524 5543
rect 6532 5537 6588 5543
rect 6820 5537 6956 5543
rect 7108 5537 7500 5543
rect 7508 5537 8492 5543
rect 8724 5537 8732 5543
rect 5181 5524 5187 5536
rect 9837 5524 9843 5536
rect 212 5517 268 5523
rect 740 5517 995 5523
rect 989 5504 995 5517
rect 1588 5517 1596 5523
rect 2052 5517 2060 5523
rect 2148 5517 2156 5523
rect 2724 5517 2940 5523
rect 2948 5517 4332 5523
rect 4372 5517 4508 5523
rect 4596 5517 4812 5523
rect 5412 5517 6524 5523
rect 6836 5517 6844 5523
rect 6852 5517 7452 5523
rect 7460 5517 7932 5523
rect 8180 5517 8236 5523
rect 8244 5517 8268 5523
rect 8436 5517 9404 5523
rect 9636 5517 9740 5523
rect 7933 5504 7939 5516
rect 660 5497 668 5503
rect 692 5497 924 5503
rect 1476 5497 1836 5503
rect 2036 5497 2044 5503
rect 2500 5497 2508 5503
rect 2532 5497 3180 5503
rect 3252 5497 3916 5503
rect 3924 5497 3932 5503
rect 4276 5497 4284 5503
rect 4596 5497 4604 5503
rect 4612 5497 4668 5503
rect 4724 5497 5180 5503
rect 5188 5497 5228 5503
rect 5396 5497 5932 5503
rect 6436 5497 7052 5503
rect 7060 5497 7548 5503
rect 7716 5497 7724 5503
rect 7956 5497 7980 5503
rect 8516 5497 8956 5503
rect 8964 5497 8972 5503
rect 9076 5497 10028 5503
rect 452 5477 732 5483
rect 932 5477 1148 5483
rect 1348 5477 1356 5483
rect 1844 5477 3580 5483
rect 5460 5477 5500 5483
rect 5732 5477 5740 5483
rect 6068 5477 6156 5483
rect 6612 5477 6620 5483
rect 6740 5477 6755 5483
rect 6820 5477 6844 5483
rect 6964 5477 7004 5483
rect 7028 5477 7260 5483
rect 7300 5477 7324 5483
rect 7396 5477 7500 5483
rect 7668 5477 8588 5483
rect 8596 5477 8956 5483
rect 9396 5477 9404 5483
rect 9444 5477 9852 5483
rect 909 5464 915 5476
rect 6717 5464 6723 5476
rect 7389 5464 7395 5476
rect 1012 5457 2444 5463
rect 3156 5457 3484 5463
rect 3812 5457 3868 5463
rect 5268 5457 5276 5463
rect 5284 5457 5356 5463
rect 5716 5457 6332 5463
rect 7700 5457 7724 5463
rect 8580 5457 8604 5463
rect 8628 5457 8652 5463
rect 8660 5457 8764 5463
rect 8996 5457 9036 5463
rect 532 5437 700 5443
rect 2708 5437 2716 5443
rect 2724 5437 3676 5443
rect 3972 5437 3996 5443
rect 7268 5437 8956 5443
rect 1149 5424 1155 5436
rect 2708 5417 2748 5423
rect 3620 5417 3628 5423
rect 6356 5417 6364 5423
rect 916 5397 1612 5403
rect 2116 5397 3004 5403
rect 3700 5397 5100 5403
rect 5124 5397 5500 5403
rect 6084 5397 6595 5403
rect 1860 5377 2060 5383
rect 2228 5377 2508 5383
rect 2532 5377 2540 5383
rect 3412 5377 3900 5383
rect 4052 5377 4060 5383
rect 4932 5377 5356 5383
rect 6244 5377 6300 5383
rect 6589 5383 6595 5397
rect 6628 5397 7660 5403
rect 8068 5397 8140 5403
rect 8413 5403 8419 5416
rect 8413 5397 8460 5403
rect 8557 5397 8892 5403
rect 8557 5384 8563 5397
rect 8948 5397 9020 5403
rect 9197 5403 9203 5416
rect 9197 5397 9324 5403
rect 9828 5397 10044 5403
rect 6589 5377 6876 5383
rect 7156 5377 7180 5383
rect 7380 5377 8172 5383
rect 8756 5377 9644 5383
rect 212 5357 252 5363
rect 340 5357 524 5363
rect 1348 5357 1356 5363
rect 1812 5357 1836 5363
rect 2036 5357 3436 5363
rect 3613 5357 4220 5363
rect 308 5337 908 5343
rect 1140 5337 1244 5343
rect 1252 5337 1436 5343
rect 1588 5337 2108 5343
rect 2228 5337 2268 5343
rect 2276 5337 2380 5343
rect 2733 5337 2748 5343
rect 2836 5337 2844 5343
rect 2868 5337 2972 5343
rect 3613 5343 3619 5357
rect 4244 5357 4364 5363
rect 4564 5357 6012 5363
rect 6196 5357 6220 5363
rect 6228 5357 6716 5363
rect 6980 5357 7180 5363
rect 7188 5357 7228 5363
rect 7428 5357 7516 5363
rect 8292 5357 8732 5363
rect 8740 5357 8924 5363
rect 8980 5357 9196 5363
rect 9444 5357 9468 5363
rect 9652 5357 9868 5363
rect 9924 5357 10028 5363
rect 10052 5357 10236 5363
rect 2980 5337 3619 5343
rect 3636 5337 3644 5343
rect 4116 5337 4124 5343
rect 4244 5337 4252 5343
rect 4756 5337 4924 5343
rect 4948 5337 5228 5343
rect 5844 5337 6124 5343
rect 6388 5337 6716 5343
rect 7060 5337 7068 5343
rect 7076 5337 7500 5343
rect 8420 5337 8428 5343
rect 8468 5337 8556 5343
rect 8644 5337 8652 5343
rect 8660 5337 8988 5343
rect 9428 5337 9596 5343
rect 9604 5337 9772 5343
rect 9780 5337 10012 5343
rect 5229 5324 5235 5336
rect 660 5317 668 5323
rect 2308 5317 2828 5323
rect 2836 5317 3180 5323
rect 3636 5317 3868 5323
rect 3956 5317 4796 5323
rect 4804 5317 4860 5323
rect 6372 5317 6380 5323
rect 6724 5317 7628 5323
rect 7860 5317 7868 5323
rect 7876 5317 9548 5323
rect 10276 5317 10339 5323
rect 1581 5304 1587 5316
rect 6141 5304 6147 5316
rect 1380 5297 1404 5303
rect 1652 5297 3020 5303
rect 3412 5297 3420 5303
rect 4052 5297 4108 5303
rect 4420 5297 4572 5303
rect 5012 5297 5020 5303
rect 5252 5297 5340 5303
rect 5492 5297 5708 5303
rect 5732 5297 5916 5303
rect 6308 5297 6476 5303
rect 6484 5297 6508 5303
rect 6516 5297 6988 5303
rect 6996 5297 7388 5303
rect 7396 5297 7532 5303
rect 7684 5297 8652 5303
rect 8660 5297 8668 5303
rect 8964 5297 9340 5303
rect 9348 5297 9548 5303
rect 9780 5297 9868 5303
rect 9876 5297 9884 5303
rect 10084 5297 10092 5303
rect 4797 5284 4803 5296
rect 916 5277 1228 5283
rect 1588 5277 1756 5283
rect 2276 5277 2284 5283
rect 2548 5277 2732 5283
rect 3204 5277 3212 5283
rect 4820 5277 5244 5283
rect 6292 5277 6684 5283
rect 6692 5277 7148 5283
rect 7412 5277 7628 5283
rect 8052 5277 8204 5283
rect 8484 5277 8524 5283
rect 8532 5277 9180 5283
rect 9380 5277 9708 5283
rect 9716 5277 9772 5283
rect 516 5257 1100 5263
rect 1572 5257 2348 5263
rect 2820 5257 4220 5263
rect 4228 5257 5260 5263
rect 5348 5257 5692 5263
rect 6340 5257 7068 5263
rect 7076 5257 7964 5263
rect 7972 5257 8428 5263
rect 8548 5257 8556 5263
rect 900 5237 2476 5243
rect 3268 5237 3276 5243
rect 3700 5237 3884 5243
rect 6676 5237 7772 5243
rect 84 5217 92 5223
rect 5956 5217 6124 5223
rect 6516 5217 6524 5223
rect 7716 5217 9612 5223
rect 7620 5197 8524 5203
rect 8532 5197 9068 5203
rect 3540 5177 3564 5183
rect 7204 5177 7212 5183
rect 8196 5177 8460 5183
rect 900 5157 908 5163
rect 2724 5157 2796 5163
rect 3188 5157 3932 5163
rect 5636 5157 5932 5163
rect 6036 5157 7468 5163
rect 452 5137 524 5143
rect 676 5137 1580 5143
rect 2132 5137 2220 5143
rect 3220 5137 3804 5143
rect 5204 5137 5500 5143
rect 5508 5137 6492 5143
rect 6564 5137 6668 5143
rect 7268 5137 7868 5143
rect 7876 5137 9692 5143
rect -51 5083 -45 5123
rect 500 5117 956 5123
rect 964 5117 972 5123
rect 1220 5117 1228 5123
rect 1572 5117 1580 5123
rect 1844 5117 2476 5123
rect 2948 5117 2956 5123
rect 3396 5117 4252 5123
rect 4260 5117 4300 5123
rect 5460 5117 5724 5123
rect 6196 5117 6284 5123
rect 6916 5117 7004 5123
rect 7300 5117 7308 5123
rect 7348 5117 7404 5123
rect 7412 5117 7436 5123
rect 8196 5117 8204 5123
rect 8468 5117 8748 5123
rect 8820 5117 8828 5123
rect 9469 5117 9484 5123
rect 5869 5104 5875 5116
rect 6653 5104 6659 5116
rect 996 5097 1084 5103
rect 1892 5097 2124 5103
rect 2164 5097 3148 5103
rect 3156 5097 4108 5103
rect 4116 5097 4300 5103
rect 4308 5097 4588 5103
rect 4596 5097 4812 5103
rect 5508 5097 5852 5103
rect 5892 5097 5916 5103
rect 5924 5097 6108 5103
rect 6660 5097 7980 5103
rect 7988 5097 8044 5103
rect 8461 5097 9036 5103
rect -51 5077 252 5083
rect 452 5077 460 5083
rect 660 5077 1132 5083
rect 1220 5077 1228 5083
rect 1348 5077 1372 5083
rect 2020 5077 2508 5083
rect 2804 5077 3244 5083
rect 3604 5077 3612 5083
rect 3956 5077 4172 5083
rect 4404 5077 4572 5083
rect 5316 5077 5404 5083
rect 5492 5077 6172 5083
rect 6180 5077 6188 5083
rect 6660 5077 6668 5083
rect 8461 5083 8467 5097
rect 6852 5077 8467 5083
rect 8852 5077 9148 5083
rect 9396 5077 9612 5083
rect 9668 5077 9708 5083
rect 9892 5077 10028 5083
rect 100 5057 524 5063
rect 900 5057 940 5063
rect 1012 5057 1676 5063
rect 2484 5057 2572 5063
rect 3108 5057 3260 5063
rect 3460 5057 3724 5063
rect 4404 5057 4412 5063
rect 5204 5057 5452 5063
rect 5460 5057 6540 5063
rect 7220 5057 7356 5063
rect 7492 5057 7868 5063
rect 7876 5057 8428 5063
rect 8756 5057 8972 5063
rect 9508 5057 9628 5063
rect 516 5037 684 5043
rect 1524 5037 1532 5043
rect 2596 5037 4092 5043
rect 6868 5037 6892 5043
rect 7140 5037 7500 5043
rect 7604 5037 7612 5043
rect 3268 5017 3468 5023
rect 3876 5017 4060 5023
rect 6804 5017 7068 5023
rect 4372 4997 4396 5003
rect 5668 4997 5836 5003
rect 6548 4997 6956 5003
rect 7524 4997 7612 5003
rect 9940 4997 10172 5003
rect 2941 4984 2947 4996
rect -51 4977 12 4983
rect 221 4977 252 4983
rect 221 4963 227 4977
rect 909 4977 972 4983
rect 909 4964 915 4977
rect 3940 4977 3948 4983
rect 4836 4977 5596 4983
rect 5636 4977 6396 4983
rect 6404 4977 6780 4983
rect 8212 4977 8220 4983
rect 8228 4977 8476 4983
rect 8573 4977 8764 4983
rect 212 4957 227 4963
rect 1124 4957 1516 4963
rect 1572 4957 1580 4963
rect 1828 4957 1900 4963
rect 2452 4957 2796 4963
rect 3492 4957 3644 4963
rect 4084 4957 4284 4963
rect 4292 4957 4524 4963
rect 4532 4957 4540 4963
rect 5572 4957 5692 4963
rect 5732 4957 5740 4963
rect 6116 4957 6156 4963
rect 6180 4957 7884 4963
rect 7892 4957 7900 4963
rect 7917 4957 8076 4963
rect 4605 4944 4611 4956
rect 1236 4937 1372 4943
rect 1524 4937 2940 4943
rect 2996 4937 3820 4943
rect 3828 4937 4172 4943
rect 4596 4937 4604 4943
rect 4941 4937 4956 4943
rect 5188 4937 6348 4943
rect 6356 4937 6380 4943
rect 6388 4937 7036 4943
rect 7044 4937 7228 4943
rect 7236 4937 7244 4943
rect 7300 4937 7308 4943
rect 7748 4937 7763 4943
rect 676 4917 1196 4923
rect 1588 4917 1596 4923
rect 1684 4917 1836 4923
rect 1844 4917 2060 4923
rect 2484 4917 2572 4923
rect 2772 4917 3260 4923
rect 5188 4917 5852 4923
rect 6532 4917 6684 4923
rect 6980 4917 7436 4923
rect 7757 4923 7763 4937
rect 7780 4937 7788 4943
rect 7917 4943 7923 4957
rect 8573 4963 8579 4977
rect 8356 4957 8579 4963
rect 9252 4957 9820 4963
rect 9828 4957 10204 4963
rect 7876 4937 7923 4943
rect 8116 4937 8124 4943
rect 8148 4937 8204 4943
rect 8404 4937 8412 4943
rect 8436 4937 8668 4943
rect 9044 4937 9068 4943
rect 9172 4937 9404 4943
rect 9572 4937 9580 4943
rect 9604 4937 9619 4943
rect 9613 4924 9619 4937
rect 9764 4937 9820 4943
rect 9908 4937 9932 4943
rect 7757 4917 8300 4923
rect 8596 4917 9180 4923
rect 1108 4897 1116 4903
rect 1124 4897 1548 4903
rect 1572 4897 1660 4903
rect 1668 4897 1772 4903
rect 1908 4897 1916 4903
rect 3028 4897 3036 4903
rect 4084 4897 4092 4903
rect 4157 4897 4172 4903
rect 4468 4897 4956 4903
rect 4964 4897 4972 4903
rect 5604 4897 5900 4903
rect 6356 4897 6508 4903
rect 6708 4897 6844 4903
rect 7028 4897 7164 4903
rect 7444 4897 7452 4903
rect 7620 4897 7644 4903
rect 7668 4897 8668 4903
rect 9396 4897 9420 4903
rect 10020 4897 10028 4903
rect 2797 4884 2803 4896
rect 9613 4884 9619 4896
rect 1108 4877 1132 4883
rect 3636 4877 4140 4883
rect 4148 4877 4524 4883
rect 4532 4877 4604 4883
rect 4612 4877 4620 4883
rect 5700 4877 5740 4883
rect 6340 4877 6988 4883
rect 7412 4877 7580 4883
rect 7588 4877 8780 4883
rect 916 4857 1404 4863
rect 3236 4857 3500 4863
rect 3844 4857 3852 4863
rect 4356 4857 4492 4863
rect 4500 4857 4572 4863
rect 4148 4837 4796 4843
rect 6516 4837 6588 4843
rect 2116 4817 2140 4823
rect 8829 4777 8972 4783
rect 8829 4763 8835 4777
rect 8740 4757 8835 4763
rect 9700 4757 9724 4763
rect 452 4737 460 4743
rect 1892 4737 2556 4743
rect 2564 4737 3036 4743
rect 3044 4737 3596 4743
rect 3604 4737 3964 4743
rect 4564 4737 4940 4743
rect 5044 4737 5052 4743
rect 5268 4737 5820 4743
rect 5828 4737 6188 4743
rect 6516 4737 6572 4743
rect 7268 4737 7660 4743
rect 7828 4737 7852 4743
rect 7876 4737 9148 4743
rect 9396 4737 9580 4743
rect 9940 4737 10092 4743
rect 77 4724 83 4736
rect 1789 4724 1795 4736
rect 6589 4724 6595 4736
rect -51 4683 -45 4723
rect 260 4717 524 4723
rect 916 4717 924 4723
rect 948 4717 1212 4723
rect 1556 4717 1564 4723
rect 2020 4717 2044 4723
rect 2484 4717 2508 4723
rect 2532 4717 2556 4723
rect 2708 4717 2716 4723
rect 2996 4717 3820 4723
rect 3828 4717 3836 4723
rect 4484 4717 4492 4723
rect 4548 4717 4572 4723
rect 4580 4717 5196 4723
rect 5476 4717 5500 4723
rect 5956 4717 6300 4723
rect 6500 4717 6572 4723
rect 6948 4717 6956 4723
rect 7684 4717 7948 4723
rect 7972 4717 8252 4723
rect 8564 4717 8588 4723
rect 2804 4697 3564 4703
rect 5188 4697 5276 4703
rect 5284 4697 5580 4703
rect 6516 4697 7036 4703
rect 7940 4697 7964 4703
rect 7972 4697 8492 4703
rect 8500 4697 8636 4703
rect 8772 4697 8796 4703
rect 9684 4697 9692 4703
rect -51 4677 12 4683
rect 84 4677 92 4683
rect 100 4677 444 4683
rect 676 4677 700 4683
rect 1140 4677 1148 4683
rect 2372 4677 2460 4683
rect 2820 4677 2828 4683
rect 3380 4677 3404 4683
rect 4276 4677 4300 4683
rect 4932 4677 4956 4683
rect 5508 4677 5532 4683
rect 5540 4677 5932 4683
rect 5956 4677 5964 4683
rect 6132 4677 6588 4683
rect 6612 4677 6636 4683
rect 6644 4677 7260 4683
rect 7268 4677 8908 4683
rect 8916 4677 9132 4683
rect 9156 4677 9228 4683
rect 9236 4677 9388 4683
rect 9588 4677 9596 4683
rect 9684 4677 9708 4683
rect 10020 4677 10252 4683
rect 909 4664 915 4676
rect 3581 4664 3587 4676
rect 9917 4664 9923 4676
rect 1156 4657 1596 4663
rect 1796 4657 1811 4663
rect 20 4637 924 4643
rect 1188 4637 1420 4643
rect 676 4597 684 4603
rect 1380 4597 1404 4603
rect 1805 4603 1811 4657
rect 1908 4657 1916 4663
rect 2676 4657 2700 4663
rect 2708 4657 2956 4663
rect 3156 4657 3180 4663
rect 4468 4657 4476 4663
rect 7012 4657 8252 4663
rect 8260 4657 8508 4663
rect 8596 4657 8764 4663
rect 8916 4657 8940 4663
rect 9204 4657 9212 4663
rect 2525 4644 2531 4656
rect 2260 4637 2268 4643
rect 3476 4637 3612 4643
rect 3876 4637 4732 4643
rect 5476 4637 6124 4643
rect 7716 4637 7836 4643
rect 8260 4637 8284 4643
rect 8756 4637 8764 4643
rect 8900 4637 8940 4643
rect 2260 4617 2268 4623
rect 4308 4617 4572 4623
rect 6292 4617 6316 4623
rect 1805 4597 1836 4603
rect 1924 4597 2300 4603
rect 2509 4603 2515 4616
rect 2509 4597 3196 4603
rect 5172 4597 5244 4603
rect 7284 4597 7388 4603
rect 7396 4597 7580 4603
rect 8052 4597 8572 4603
rect 9892 4597 9900 4603
rect 9908 4597 10028 4603
rect -51 4577 12 4583
rect 1348 4577 1372 4583
rect 2068 4577 2108 4583
rect 2276 4577 2284 4583
rect 2292 4577 2460 4583
rect 3860 4577 3916 4583
rect 4068 4577 4140 4583
rect 4276 4577 4300 4583
rect 7764 4577 8284 4583
rect 212 4557 236 4563
rect 532 4557 908 4563
rect 1620 4557 2572 4563
rect 2948 4557 3100 4563
rect 3108 4557 3148 4563
rect 3812 4557 4156 4563
rect 4180 4557 4732 4563
rect 4740 4557 4828 4563
rect 5956 4557 5964 4563
rect 5972 4557 6108 4563
rect 6164 4557 7004 4563
rect 8324 4557 8444 4563
rect 8580 4557 8716 4563
rect 9556 4557 9580 4563
rect 244 4537 316 4543
rect 548 4537 556 4543
rect 996 4537 1100 4543
rect 1140 4537 1148 4543
rect 1604 4537 1612 4543
rect 1700 4537 1715 4543
rect 1940 4537 2412 4543
rect 2420 4537 2444 4543
rect 2468 4537 2492 4543
rect 2820 4537 2908 4543
rect 2916 4537 2956 4543
rect 3380 4537 3388 4543
rect 3588 4537 4348 4543
rect 4356 4537 4508 4543
rect 4660 4537 4732 4543
rect 5348 4537 5356 4543
rect 5604 4537 5740 4543
rect 5844 4537 6316 4543
rect 6324 4537 6604 4543
rect 6612 4537 6620 4543
rect 6628 4537 7484 4543
rect 8052 4537 9004 4543
rect 9012 4537 9020 4543
rect 9028 4537 9116 4543
rect 9220 4537 9404 4543
rect 9780 4537 9795 4543
rect 1252 4517 1436 4523
rect 1444 4517 2076 4523
rect 2084 4517 2988 4523
rect 3620 4517 3644 4523
rect 3844 4517 3868 4523
rect 3940 4517 4268 4523
rect 6340 4517 6476 4523
rect 6708 4517 6716 4523
rect 6724 4517 6828 4523
rect 7444 4517 7900 4523
rect 8132 4517 8156 4523
rect 8484 4517 8780 4523
rect 5917 4504 5923 4516
rect 308 4497 316 4503
rect 676 4497 684 4503
rect 1428 4497 1900 4503
rect 1908 4497 2956 4503
rect 3156 4497 3388 4503
rect 3860 4497 3868 4503
rect 4068 4497 4076 4503
rect 4756 4497 5020 4503
rect 5028 4497 5036 4503
rect 6500 4497 6588 4503
rect 7156 4497 7164 4503
rect 7268 4497 7276 4503
rect 8820 4497 8892 4503
rect 9668 4497 9692 4503
rect 9700 4497 9788 4503
rect 9133 4484 9139 4496
rect 1252 4477 1548 4483
rect 1556 4477 2460 4483
rect 2468 4477 2492 4483
rect 2772 4477 2780 4483
rect 2804 4477 3356 4483
rect 3364 4477 3388 4483
rect 3844 4477 4796 4483
rect 4804 4477 5372 4483
rect 6484 4477 6492 4483
rect 7188 4477 7468 4483
rect 500 4457 748 4463
rect 1604 4457 1612 4463
rect 2260 4457 2268 4463
rect 2804 4457 3004 4463
rect 5620 4457 5836 4463
rect 5844 4457 6140 4463
rect 6148 4457 6828 4463
rect 6836 4457 7052 4463
rect 3165 4444 3171 4456
rect 692 4437 892 4443
rect 2052 4437 2668 4443
rect 7252 4437 9164 4443
rect 9172 4437 9180 4443
rect 1165 4384 1171 4396
rect 1588 4377 1644 4383
rect 3204 4377 3884 4383
rect 2644 4357 3660 4363
rect 5396 4357 5452 4363
rect 7844 4357 7884 4363
rect 7908 4357 8812 4363
rect 8820 4357 9500 4363
rect 9508 4357 9548 4363
rect 212 4337 284 4343
rect 3572 4337 3612 4343
rect 4932 4337 5180 4343
rect 5652 4337 6156 4343
rect 6612 4337 6620 4343
rect 6628 4337 7852 4343
rect 8436 4337 8476 4343
rect 8628 4337 8828 4343
rect 9220 4337 9612 4343
rect 564 4317 572 4323
rect 909 4317 915 4336
rect 9853 4324 9859 4336
rect 948 4317 1004 4323
rect 1364 4317 1644 4323
rect 2260 4317 2268 4323
rect 2340 4317 2460 4323
rect 2468 4317 2796 4323
rect 3380 4317 3596 4323
rect 3620 4317 3756 4323
rect 3828 4317 4316 4323
rect 4324 4317 4332 4323
rect 4532 4317 4572 4323
rect 5092 4317 5100 4323
rect 5604 4317 5612 4323
rect 6372 4317 6380 4323
rect 6388 4317 7100 4323
rect 7220 4317 7260 4323
rect 7460 4317 7468 4323
rect 7716 4317 8188 4323
rect 8196 4317 8540 4323
rect 8612 4317 8620 4323
rect 7325 4304 7331 4316
rect 1428 4297 1436 4303
rect 1748 4297 2556 4303
rect 2692 4297 2700 4303
rect 3396 4297 3804 4303
rect 3812 4297 3820 4303
rect 4244 4297 4860 4303
rect 4868 4297 5068 4303
rect 6388 4297 7244 4303
rect 7252 4297 7292 4303
rect 7556 4297 7708 4303
rect 7892 4297 8412 4303
rect 8724 4297 8844 4303
rect 9396 4297 9932 4303
rect 3149 4284 3155 4296
rect 100 4277 220 4283
rect 548 4277 556 4283
rect 900 4277 908 4283
rect 1012 4277 1020 4283
rect 1796 4277 1820 4283
rect 2260 4277 2268 4283
rect 2484 4277 2716 4283
rect 4228 4277 4540 4283
rect 5220 4277 5388 4283
rect 5732 4277 5756 4283
rect 6164 4277 6268 4283
rect 6276 4277 7628 4283
rect 7652 4277 7660 4283
rect 7684 4277 7692 4283
rect 8036 4277 8092 4283
rect 8228 4277 8556 4283
rect 8644 4277 8732 4283
rect 9236 4277 9372 4283
rect 9828 4277 9843 4283
rect 3997 4264 4003 4276
rect 9165 4264 9171 4276
rect 676 4257 2012 4263
rect 3012 4257 3164 4263
rect 3172 4257 3404 4263
rect 3588 4257 3948 4263
rect 4084 4257 4684 4263
rect 5060 4257 5276 4263
rect 5924 4257 6188 4263
rect 6612 4257 6668 4263
rect 6788 4257 7164 4263
rect 7172 4257 7916 4263
rect 7956 4257 8300 4263
rect 9140 4257 9148 4263
rect -51 4237 12 4243
rect 772 4237 780 4243
rect 2596 4237 2956 4243
rect 3412 4237 3420 4243
rect 3796 4237 4316 4243
rect 4548 4237 4700 4243
rect 5668 4237 6012 4243
rect 6020 4237 6140 4243
rect 6356 4237 6812 4243
rect 6900 4237 8332 4243
rect 8612 4237 9036 4243
rect 1581 4224 1587 4236
rect 452 4217 924 4223
rect 1828 4217 2492 4223
rect 2532 4217 3660 4223
rect 6484 4217 6668 4223
rect 6676 4217 7340 4223
rect 7556 4217 7564 4223
rect 7604 4217 7740 4223
rect 916 4197 1612 4203
rect 2708 4197 2716 4203
rect 2740 4197 3420 4203
rect 6596 4197 7180 4203
rect 7268 4197 8332 4203
rect 8500 4197 8524 4203
rect 1604 4177 2092 4183
rect 2893 4177 2956 4183
rect 212 4157 236 4163
rect 1204 4157 1228 4163
rect 1812 4157 1836 4163
rect 2893 4163 2899 4177
rect 5156 4177 5164 4183
rect 6164 4177 8412 4183
rect 8420 4177 8604 4183
rect 10276 4177 10339 4183
rect 2708 4157 2899 4163
rect 2916 4157 3132 4163
rect 5060 4157 5260 4163
rect 5988 4157 6188 4163
rect 6212 4157 6828 4163
rect 7124 4157 7340 4163
rect 7396 4157 7404 4163
rect 7428 4157 7484 4163
rect 7844 4157 8236 4163
rect 8244 4157 8956 4163
rect 8964 4157 8972 4163
rect 9044 4157 9564 4163
rect 9572 4157 9916 4163
rect 2461 4144 2467 4156
rect 228 4137 316 4143
rect 772 4137 1116 4143
rect 1124 4137 1388 4143
rect 2020 4137 2028 4143
rect 2500 4137 2924 4143
rect 3620 4137 3628 4143
rect 4068 4137 4364 4143
rect 4660 4137 4668 4143
rect 4948 4137 4963 4143
rect 5076 4137 5308 4143
rect 5748 4137 5756 4143
rect 5764 4137 6188 4143
rect 6420 4137 6460 4143
rect 6756 4137 7244 4143
rect 7252 4137 7964 4143
rect 8132 4137 8716 4143
rect 9284 4137 9548 4143
rect 9908 4137 9923 4143
rect 1588 4117 1820 4123
rect 2804 4117 3148 4123
rect 3156 4117 3180 4123
rect 3380 4117 3852 4123
rect 4477 4123 4483 4136
rect 4477 4117 4524 4123
rect 4925 4123 4931 4136
rect 5389 4124 5395 4136
rect 8733 4124 8739 4136
rect 9277 4124 9283 4136
rect 9917 4124 9923 4137
rect 4925 4117 4972 4123
rect 5636 4117 6028 4123
rect 6036 4117 6700 4123
rect 6708 4117 7484 4123
rect 7684 4117 7708 4123
rect 7732 4117 7836 4123
rect 7876 4117 7932 4123
rect 8356 4117 8604 4123
rect 8900 4117 9036 4123
rect 9492 4117 9708 4123
rect 765 4104 771 4116
rect 324 4097 332 4103
rect 1108 4097 1116 4103
rect 1213 4097 1228 4103
rect 1428 4097 1580 4103
rect 2484 4097 3452 4103
rect 3604 4097 3612 4103
rect 4052 4097 4140 4103
rect 4148 4097 4188 4103
rect 4580 4097 4732 4103
rect 4740 4097 4748 4103
rect 5428 4097 5708 4103
rect 5716 4097 6076 4103
rect 6180 4097 6188 4103
rect 6740 4097 6748 4103
rect 6852 4097 6892 4103
rect 7636 4097 8492 4103
rect 8516 4097 8956 4103
rect 9140 4097 9276 4103
rect 9284 4097 9884 4103
rect 525 4084 531 4096
rect 660 4077 1196 4083
rect 1204 4077 2236 4083
rect 2244 4077 2540 4083
rect 2548 4077 2652 4083
rect 2708 4077 2732 4083
rect 2884 4077 3020 4083
rect 3028 4077 3836 4083
rect 5748 4077 5756 4083
rect 5972 4077 6172 4083
rect 6180 4077 6780 4083
rect 6788 4077 7468 4083
rect 7492 4077 7676 4083
rect 7716 4077 7836 4083
rect 7924 4077 8732 4083
rect 8740 4077 8812 4083
rect 9076 4077 9516 4083
rect 9572 4077 9580 4083
rect 1620 4057 2476 4063
rect 3396 4057 3404 4063
rect 4164 4057 4172 4063
rect 4340 4057 4588 4063
rect 5764 4057 6188 4063
rect 6196 4057 6428 4063
rect 6980 4057 7404 4063
rect 7412 4057 7548 4063
rect 3460 4037 5356 4043
rect 7380 4037 7692 4043
rect 9620 4017 9628 4023
rect 5300 3997 5484 4003
rect 4084 3977 5340 3983
rect 6756 3977 6860 3983
rect 6868 3977 6988 3983
rect 1181 3957 1772 3963
rect 1181 3943 1187 3957
rect 9892 3957 10076 3963
rect 484 3937 1187 3943
rect 1204 3937 1228 3943
rect 1236 3937 1884 3943
rect 2244 3937 2284 3943
rect 2740 3937 2908 3943
rect 4388 3937 5004 3943
rect 5076 3937 5132 3943
rect 5524 3937 5532 3943
rect 5540 3937 5548 3943
rect 5732 3937 5836 3943
rect 5876 3937 6012 3943
rect 6148 3937 6172 3943
rect 7908 3937 8524 3943
rect 8548 3937 8620 3943
rect 8868 3937 9436 3943
rect 3373 3924 3379 3936
rect 4381 3924 4387 3936
rect 1108 3917 2876 3923
rect 2916 3917 2924 3923
rect 3924 3917 3932 3923
rect 4852 3917 5516 3923
rect 5524 3917 6156 3923
rect 6388 3917 6396 3923
rect 7268 3917 7276 3923
rect 7492 3917 9132 3923
rect 9140 3917 9212 3923
rect 9220 3917 9228 3923
rect 9668 3917 9852 3923
rect 429 3904 435 3916
rect 6829 3904 6835 3916
rect 7389 3904 7395 3916
rect 1156 3897 1420 3903
rect 1556 3897 1612 3903
rect 1620 3897 1868 3903
rect 2468 3897 2588 3903
rect 2724 3897 3196 3903
rect 3204 3897 3612 3903
rect 3828 3897 3868 3903
rect 4068 3897 4604 3903
rect 4628 3897 4652 3903
rect 5076 3897 6620 3903
rect 7172 3897 7260 3903
rect 7668 3897 7692 3903
rect 8468 3897 9100 3903
rect 9108 3897 9116 3903
rect 9124 3897 9260 3903
rect 9652 3897 9660 3903
rect 205 3877 220 3883
rect 340 3877 1020 3883
rect 1124 3877 1196 3883
rect 1220 3877 1596 3883
rect 1604 3877 1740 3883
rect 1764 3877 1884 3883
rect 1892 3877 3020 3883
rect 3268 3877 3372 3883
rect 3604 3877 3916 3883
rect 4292 3877 4300 3883
rect 4404 3877 4828 3883
rect 4836 3877 4844 3883
rect 5492 3877 5628 3883
rect 5652 3877 5868 3883
rect 6020 3877 6188 3883
rect 6196 3877 6508 3883
rect 6516 3877 6652 3883
rect 6820 3877 6828 3883
rect 7140 3877 7260 3883
rect 7268 3877 7468 3883
rect 7620 3877 7708 3883
rect 7924 3877 8092 3883
rect 8452 3877 8460 3883
rect 8788 3877 9452 3883
rect 9460 3877 9852 3883
rect 10052 3877 10092 3883
rect 3133 3864 3139 3876
rect 292 3857 636 3863
rect 644 3857 652 3863
rect 1780 3857 1788 3863
rect 2484 3857 2716 3863
rect 2916 3857 2956 3863
rect 3172 3857 3628 3863
rect 3636 3857 4556 3863
rect 5508 3857 5532 3863
rect 5716 3857 6060 3863
rect 6068 3857 6092 3863
rect 6644 3857 6796 3863
rect 7252 3857 7660 3863
rect 7684 3857 8044 3863
rect 8308 3857 8732 3863
rect 8740 3857 9164 3863
rect 9172 3857 9212 3863
rect 260 3837 300 3843
rect 740 3837 1004 3843
rect 1028 3837 4140 3843
rect 5268 3837 5564 3843
rect 7828 3837 7836 3843
rect 8308 3837 9100 3843
rect 9124 3837 9132 3843
rect 244 3817 2092 3823
rect 2132 3817 2748 3823
rect 7204 3817 7843 3823
rect 244 3797 252 3803
rect 2020 3797 2044 3803
rect 2532 3797 2540 3803
rect 4308 3797 4364 3803
rect 6836 3797 7820 3803
rect 7837 3803 7843 3817
rect 8372 3817 8476 3823
rect 7837 3797 8732 3803
rect 8980 3797 9468 3803
rect 9924 3797 10092 3803
rect -51 3777 12 3783
rect 228 3777 1148 3783
rect 1860 3777 3420 3783
rect 3956 3777 3964 3783
rect 4749 3777 4796 3783
rect 292 3757 444 3763
rect 1684 3757 1804 3763
rect 2036 3757 2268 3763
rect 2420 3757 3708 3763
rect 3716 3757 4044 3763
rect 4164 3757 4284 3763
rect 4749 3763 4755 3777
rect 6420 3777 6428 3783
rect 7005 3777 7020 3783
rect 7188 3777 7212 3783
rect 7444 3777 7676 3783
rect 8772 3777 8988 3783
rect 4740 3757 4755 3763
rect 4772 3757 4956 3763
rect 5188 3757 5196 3763
rect 6868 3757 7468 3763
rect 7700 3757 8163 3763
rect 5421 3744 5427 3756
rect 676 3737 732 3743
rect 1348 3737 1356 3743
rect 1748 3737 2012 3743
rect 2260 3737 2524 3743
rect 2676 3737 2684 3743
rect 3172 3737 3180 3743
rect 3405 3737 3420 3743
rect 3636 3737 3660 3743
rect 4116 3737 5420 3743
rect 5540 3737 5548 3743
rect 6180 3737 6188 3743
rect 6196 3737 7052 3743
rect 7060 3737 7068 3743
rect 7348 3737 7388 3743
rect 7860 3737 7868 3743
rect 8157 3743 8163 3757
rect 8180 3757 8460 3763
rect 8484 3757 8604 3763
rect 9284 3757 9356 3763
rect 9460 3757 9692 3763
rect 8157 3737 8396 3743
rect 8852 3737 8908 3743
rect 9172 3737 9292 3743
rect 9508 3737 9612 3743
rect 9860 3737 10012 3743
rect 2589 3724 2595 3736
rect 2036 3717 2332 3723
rect 2468 3717 2476 3723
rect 3412 3717 3436 3723
rect 4308 3717 4492 3723
rect 4996 3717 5196 3723
rect 5204 3717 5420 3723
rect 6596 3717 6956 3723
rect 6980 3717 6988 3723
rect 7101 3723 7107 3736
rect 7101 3717 8828 3723
rect 9028 3717 9180 3723
rect 9188 3717 9260 3723
rect 9821 3723 9827 3736
rect 9821 3717 9852 3723
rect 6173 3704 6179 3716
rect 9469 3704 9475 3716
rect 916 3697 956 3703
rect 1588 3697 1596 3703
rect 2596 3697 2636 3703
rect 2788 3697 2940 3703
rect 3188 3697 3772 3703
rect 3780 3697 4028 3703
rect 4036 3697 4060 3703
rect 4308 3697 4316 3703
rect 4516 3697 4524 3703
rect 5748 3697 5756 3703
rect 7492 3697 7500 3703
rect 7700 3697 8172 3703
rect 1117 3684 1123 3696
rect 4749 3684 4755 3696
rect 5533 3684 5539 3696
rect 1348 3677 3180 3683
rect 3700 3677 3804 3683
rect 3812 3677 3916 3683
rect 6180 3677 6604 3683
rect 8148 3677 8236 3683
rect 68 3657 204 3663
rect 1140 3657 1756 3663
rect 2244 3657 2252 3663
rect 5764 3637 5900 3643
rect 3732 3617 3740 3623
rect 8132 3617 8140 3623
rect 2564 3597 2588 3603
rect 1844 3577 4124 3583
rect 8356 3577 8380 3583
rect 8388 3577 8572 3583
rect 1108 3557 1116 3563
rect 6404 3557 6572 3563
rect 6580 3557 6940 3563
rect 7684 3557 7708 3563
rect 340 3537 1340 3543
rect 4932 3537 5148 3543
rect 5380 3537 5788 3543
rect 6132 3537 6636 3543
rect 6644 3537 7612 3543
rect 7620 3537 7708 3543
rect 7956 3537 8348 3543
rect 8356 3537 9676 3543
rect 9684 3537 9708 3543
rect 5805 3524 5811 3536
rect 9901 3524 9907 3536
rect 100 3517 444 3523
rect 676 3517 1628 3523
rect 2477 3517 2492 3523
rect 2532 3517 3372 3523
rect 3380 3517 3388 3523
rect 4484 3517 4780 3523
rect 5156 3517 5388 3523
rect 5812 3517 6860 3523
rect 7236 3517 7580 3523
rect 7812 3517 7820 3523
rect 7828 3517 7900 3523
rect 8356 3517 9388 3523
rect 9396 3517 9452 3523
rect 10100 3517 10115 3523
rect 2029 3504 2035 3516
rect 68 3497 316 3503
rect 900 3497 908 3503
rect 964 3497 1196 3503
rect 1412 3497 1660 3503
rect 2036 3497 3356 3503
rect 3380 3497 3596 3503
rect 3604 3497 3996 3503
rect 4004 3497 4300 3503
rect 4308 3497 4508 3503
rect 4548 3497 4780 3503
rect 6548 3497 6572 3503
rect 6580 3497 6780 3503
rect 7172 3497 7372 3503
rect 7716 3497 8492 3503
rect 8500 3497 8508 3503
rect 9044 3497 9228 3503
rect 9252 3497 9324 3503
rect 4797 3484 4803 3496
rect 212 3477 236 3483
rect 900 3477 956 3483
rect 964 3477 2092 3483
rect 2228 3477 2252 3483
rect 2292 3477 2444 3483
rect 2692 3477 2716 3483
rect 2932 3477 2972 3483
rect 3156 3477 3164 3483
rect 3380 3477 3388 3483
rect 3588 3477 4092 3483
rect 4468 3477 4476 3483
rect 4484 3477 4556 3483
rect 5332 3477 5347 3483
rect 5796 3477 5804 3483
rect 5812 3477 6044 3483
rect 6132 3477 6140 3483
rect 6148 3477 6364 3483
rect 6436 3477 6572 3483
rect 7124 3477 7132 3483
rect 7236 3477 7244 3483
rect 7540 3477 7916 3483
rect 7924 3477 8300 3483
rect 8356 3477 8572 3483
rect 8820 3477 8908 3483
rect 8980 3477 9132 3483
rect 9140 3477 9468 3483
rect 9684 3477 9692 3483
rect 9924 3477 10252 3483
rect 445 3464 451 3476
rect 3581 3464 3587 3476
rect 548 3457 940 3463
rect 1188 3457 1452 3463
rect 1652 3457 1788 3463
rect 1812 3457 1820 3463
rect 2020 3457 3571 3463
rect 1780 3437 2044 3443
rect 2244 3437 2268 3443
rect 3156 3437 3228 3443
rect 3565 3443 3571 3457
rect 3613 3457 3628 3463
rect 3876 3457 4124 3463
rect 4132 3457 4284 3463
rect 4516 3457 4572 3463
rect 4589 3457 5148 3463
rect 3565 3437 3596 3443
rect 3604 3437 3996 3443
rect 4244 3437 4259 3443
rect 4589 3443 4595 3457
rect 5332 3457 5468 3463
rect 5844 3457 5916 3463
rect 7076 3457 7228 3463
rect 7364 3457 7564 3463
rect 8372 3457 8476 3463
rect 8580 3457 9020 3463
rect 4292 3437 4595 3443
rect 4612 3437 4620 3443
rect 4628 3437 4716 3443
rect 4996 3437 5660 3443
rect 6852 3437 6860 3443
rect 7332 3437 7388 3443
rect 7396 3437 8588 3443
rect 8884 3437 8988 3443
rect 8996 3437 9068 3443
rect 308 3417 332 3423
rect 2221 3423 2227 3436
rect 2221 3417 2572 3423
rect 2276 3397 3452 3403
rect 4324 3397 4332 3403
rect 5732 3397 6284 3403
rect 6628 3397 6764 3403
rect 2132 3377 2387 3383
rect 2381 3364 2387 3377
rect 2740 3377 3644 3383
rect 5700 3377 5724 3383
rect 5748 3377 5756 3383
rect 6100 3377 6108 3383
rect 6164 3377 6172 3383
rect 7716 3377 7820 3383
rect 8260 3377 8268 3383
rect 2148 3357 2156 3363
rect 2564 3357 2780 3363
rect 2804 3357 2828 3363
rect 2852 3357 2972 3363
rect 3188 3357 3196 3363
rect 3412 3357 3836 3363
rect 3844 3357 3852 3363
rect 4948 3357 4988 3363
rect 5524 3357 5548 3363
rect 5556 3357 6012 3363
rect 6020 3357 6636 3363
rect 7988 3357 8124 3363
rect 8132 3357 8428 3363
rect 8436 3357 9372 3363
rect 9540 3357 9644 3363
rect 9844 3357 10060 3363
rect 676 3337 684 3343
rect 916 3337 972 3343
rect 1012 3337 1132 3343
rect 1588 3337 1596 3343
rect 2116 3337 4156 3343
rect 4164 3337 4172 3343
rect 4516 3337 4524 3343
rect 5092 3337 5292 3343
rect 5300 3337 5388 3343
rect 5396 3337 6140 3343
rect 6148 3337 6188 3343
rect 6525 3337 6540 3343
rect 6916 3337 6924 3343
rect 7076 3337 7100 3343
rect 7316 3337 7388 3343
rect 7444 3337 7452 3343
rect 7492 3337 8172 3343
rect 8196 3337 8364 3343
rect 8701 3337 8716 3343
rect 212 3317 988 3323
rect 996 3317 1004 3323
rect 1588 3317 1708 3323
rect 1940 3317 3356 3323
rect 4084 3317 4604 3323
rect 5188 3317 5532 3323
rect 5540 3317 6268 3323
rect 6276 3317 7132 3323
rect 7652 3317 7964 3323
rect 8436 3317 8604 3323
rect 8701 3323 8707 3337
rect 8852 3337 8860 3343
rect 9172 3337 9244 3343
rect 9620 3337 9916 3343
rect 10036 3337 10044 3343
rect 8660 3317 8707 3323
rect 228 3297 236 3303
rect 452 3297 460 3303
rect 1444 3297 1692 3303
rect 1892 3297 1916 3303
rect 1924 3297 3100 3303
rect 3172 3297 3180 3303
rect 3236 3297 3404 3303
rect 3620 3297 4092 3303
rect 4100 3297 4316 3303
rect 4532 3297 4556 3303
rect 4724 3297 5004 3303
rect 5188 3297 5196 3303
rect 5412 3297 5948 3303
rect 5956 3297 6236 3303
rect 6292 3297 6307 3303
rect 6516 3297 6540 3303
rect 6548 3297 6716 3303
rect 6852 3297 6860 3303
rect 6868 3297 7276 3303
rect 7284 3297 7516 3303
rect 7956 3297 8188 3303
rect 8388 3297 8652 3303
rect 9492 3297 9532 3303
rect 7949 3284 7955 3296
rect 1604 3277 1612 3283
rect 2244 3277 2284 3283
rect 2820 3277 2844 3283
rect 3220 3277 3244 3283
rect 3252 3277 3612 3283
rect 3748 3277 3820 3283
rect 3828 3277 4060 3283
rect 5508 3277 6204 3283
rect 7316 3277 7644 3283
rect 1140 3257 1164 3263
rect 3412 3257 3612 3263
rect 3796 3257 3916 3263
rect 6852 3257 6876 3263
rect 6068 3237 7740 3243
rect 7748 3237 7884 3243
rect 2525 3203 2531 3216
rect 1604 3197 3052 3203
rect 1069 3177 3836 3183
rect 1069 3163 1075 3177
rect 5044 3177 5772 3183
rect 948 3157 1075 3163
rect 2292 3157 2380 3163
rect 2388 3157 2492 3163
rect 5444 3157 6156 3163
rect 6164 3157 6412 3163
rect 516 3137 876 3143
rect 1540 3137 2524 3143
rect 3092 3137 3868 3143
rect 4212 3137 4220 3143
rect 5124 3137 5132 3143
rect 5476 3137 5484 3143
rect 6644 3137 6652 3143
rect 6852 3137 6860 3143
rect 8548 3137 10076 3143
rect 5357 3124 5363 3136
rect 292 3117 652 3123
rect 1092 3117 1100 3123
rect 1204 3117 1212 3123
rect 1380 3117 1852 3123
rect 2084 3117 2460 3123
rect 2468 3117 2956 3123
rect 2980 3117 3148 3123
rect 3460 3117 3532 3123
rect 3620 3117 3756 3123
rect 3764 3117 3772 3123
rect 4068 3117 4492 3123
rect 4500 3117 4988 3123
rect 4996 3117 5244 3123
rect 5252 3117 5260 3123
rect 5396 3117 7228 3123
rect 7860 3117 8076 3123
rect 8084 3117 8092 3123
rect 8292 3117 8988 3123
rect 8996 3117 9052 3123
rect 9204 3117 9219 3123
rect 9300 3117 9452 3123
rect 9460 3117 9692 3123
rect 10276 3117 10339 3123
rect 692 3097 1532 3103
rect 2420 3097 2428 3103
rect 2484 3097 2844 3103
rect 2868 3097 2876 3103
rect 4292 3097 4828 3103
rect 5060 3097 5148 3103
rect 6180 3097 6428 3103
rect 6884 3097 7212 3103
rect 8596 3097 9244 3103
rect 9284 3097 9484 3103
rect 9492 3097 9660 3103
rect 4285 3084 4291 3096
rect 1092 3077 1244 3083
rect 1252 3077 2412 3083
rect 2532 3077 2716 3083
rect 2756 3077 3052 3083
rect 3316 3077 3340 3083
rect 3540 3077 3548 3083
rect 3741 3077 3756 3083
rect 4189 3077 4204 3083
rect 4580 3077 4588 3083
rect 4628 3077 4636 3083
rect 4836 3077 5180 3083
rect 5188 3077 5388 3083
rect 5444 3077 5564 3083
rect 5732 3077 5788 3083
rect 5956 3077 5996 3083
rect 6084 3077 6652 3083
rect 6660 3077 6892 3083
rect 7284 3077 7420 3083
rect 7524 3077 7548 3083
rect 7684 3077 8060 3083
rect 8077 3077 8108 3083
rect 724 3057 1164 3063
rect 1188 3057 1196 3063
rect 1220 3057 1388 3063
rect 1620 3057 1644 3063
rect 2052 3057 2076 3063
rect 2100 3057 2220 3063
rect 2548 3057 2668 3063
rect 3876 3057 3980 3063
rect 4164 3057 4556 3063
rect 4564 3057 4652 3063
rect 4948 3057 5036 3063
rect 5044 3057 5244 3063
rect 5652 3057 6204 3063
rect 6884 3057 6908 3063
rect 8077 3063 8083 3077
rect 8404 3077 8412 3083
rect 8740 3077 9100 3083
rect 9252 3077 9260 3083
rect 10036 3077 10044 3083
rect 7924 3057 8083 3063
rect 8100 3057 9484 3063
rect 9492 3057 10092 3063
rect 196 2997 204 3003
rect 525 3003 531 3056
rect 2164 3037 2220 3043
rect 2228 3037 2716 3043
rect 3188 3037 3212 3043
rect 4356 3037 4428 3043
rect 4916 3037 4924 3043
rect 4996 3037 5036 3043
rect 6068 3037 6092 3043
rect 6340 3037 6348 3043
rect 6932 3037 7068 3043
rect 7076 3037 7932 3043
rect 8116 3037 8812 3043
rect 8916 3037 8940 3043
rect 4477 3024 4483 3036
rect 2468 3017 2556 3023
rect 4532 3017 4940 3023
rect 6356 3017 7020 3023
rect 7229 3017 7708 3023
rect 516 2997 531 3003
rect 1268 2997 1324 3003
rect 1620 2997 1788 3003
rect 2548 2997 2732 3003
rect 2836 2997 2844 3003
rect 2852 2997 2924 3003
rect 3325 3003 3331 3016
rect 7229 3004 7235 3017
rect 3325 2997 3372 3003
rect 6996 2997 7004 3003
rect 7604 2997 7788 3003
rect 8148 2997 8236 3003
rect 8308 2997 8460 3003
rect 9588 2997 9628 3003
rect 4701 2984 4707 2996
rect 2660 2977 2716 2983
rect 3092 2977 4700 2983
rect 6980 2977 7292 2983
rect 7412 2977 7676 2983
rect 7860 2977 7868 2983
rect 8084 2977 8732 2983
rect 9236 2977 9308 2983
rect 9620 2977 9836 2983
rect 68 2957 92 2963
rect 125 2957 284 2963
rect 125 2943 131 2957
rect 644 2957 652 2963
rect 1636 2957 2092 2963
rect 2676 2957 3116 2963
rect 3124 2957 3244 2963
rect 5572 2957 6124 2963
rect 6141 2957 6252 2963
rect 84 2937 131 2943
rect 436 2937 444 2943
rect 676 2937 732 2943
rect 1988 2937 2243 2943
rect 1316 2917 1420 2923
rect 1764 2917 2028 2923
rect 2237 2923 2243 2937
rect 2660 2937 2684 2943
rect 2900 2937 3196 2943
rect 3572 2937 4348 2943
rect 5140 2937 5164 2943
rect 5332 2937 5356 2943
rect 6004 2937 6012 2943
rect 6141 2943 6147 2957
rect 6724 2957 7564 2963
rect 7636 2957 7676 2963
rect 7700 2957 8332 2963
rect 9133 2944 9139 2956
rect 9373 2944 9379 2956
rect 6100 2937 6147 2943
rect 6244 2937 6268 2943
rect 6580 2937 6588 2943
rect 6900 2937 6908 2943
rect 6916 2937 7052 2943
rect 7524 2937 8908 2943
rect 9700 2937 9708 2943
rect 9908 2937 9932 2943
rect 2237 2917 2316 2923
rect 2324 2917 2332 2923
rect 3428 2917 3596 2923
rect 3956 2917 4572 2923
rect 5364 2917 6604 2923
rect 6756 2917 7004 2923
rect 7316 2917 7948 2923
rect 7956 2917 8012 2923
rect 8036 2917 8092 2923
rect 8340 2917 8540 2923
rect 8548 2917 8556 2923
rect 9380 2917 9676 2923
rect 9684 2917 9884 2923
rect 9892 2917 9916 2923
rect 436 2897 668 2903
rect 740 2897 844 2903
rect 852 2897 972 2903
rect 1844 2897 2012 2903
rect 2100 2897 2860 2903
rect 2900 2897 2956 2903
rect 3108 2897 3196 2903
rect 3204 2897 3804 2903
rect 3812 2897 3820 2903
rect 4228 2897 4236 2903
rect 4324 2897 4348 2903
rect 4932 2897 4940 2903
rect 5588 2897 5772 2903
rect 6036 2897 6220 2903
rect 6228 2897 6236 2903
rect 6340 2897 6348 2903
rect 6452 2897 6540 2903
rect 7108 2897 7196 2903
rect 7252 2897 7468 2903
rect 7476 2897 7644 2903
rect 7876 2897 7884 2903
rect 8276 2897 8332 2903
rect 8340 2897 8348 2903
rect 8388 2897 8540 2903
rect 8548 2897 8556 2903
rect 9060 2897 9148 2903
rect 9156 2897 9228 2903
rect 9908 2897 9916 2903
rect 9677 2884 9683 2896
rect 660 2877 764 2883
rect 3748 2877 4540 2883
rect 4548 2877 4908 2883
rect 6068 2877 6172 2883
rect 7428 2877 7996 2883
rect 8948 2877 9180 2883
rect 2292 2857 2332 2863
rect 3588 2857 3603 2863
rect 276 2837 700 2843
rect 708 2837 1180 2843
rect 2900 2817 2940 2823
rect 3597 2804 3603 2857
rect 7892 2857 8620 2863
rect 4276 2837 5132 2843
rect 7508 2837 8380 2843
rect 1188 2797 1548 2803
rect 1556 2797 1852 2803
rect 6692 2797 7148 2803
rect 2324 2777 2332 2783
rect 2932 2777 2988 2783
rect 6724 2777 6732 2783
rect 948 2757 1260 2763
rect 1268 2757 1292 2763
rect 2260 2757 2316 2763
rect 2708 2757 2716 2763
rect 3604 2757 3836 2763
rect 3844 2757 4092 2763
rect 4660 2757 4668 2763
rect 6740 2757 7564 2763
rect 628 2737 1084 2743
rect 1092 2737 1228 2743
rect 1236 2737 3100 2743
rect 3108 2737 4012 2743
rect 4020 2737 4268 2743
rect 4276 2737 4972 2743
rect 6628 2737 6636 2743
rect 6644 2737 7596 2743
rect 7620 2737 7788 2743
rect 8532 2737 8540 2743
rect 8724 2737 9660 2743
rect 1092 2717 1452 2723
rect 2036 2717 2860 2723
rect 2909 2717 2924 2723
rect 3220 2717 3228 2723
rect 3380 2717 3788 2723
rect 3796 2717 4012 2723
rect 4020 2717 4028 2723
rect 4324 2717 4716 2723
rect 4724 2717 5532 2723
rect 6180 2717 6188 2723
rect 6276 2717 6332 2723
rect 6500 2717 6732 2723
rect 6820 2717 6892 2723
rect 8068 2717 8764 2723
rect 8932 2717 8956 2723
rect 9316 2717 9500 2723
rect 9956 2717 9964 2723
rect 9988 2717 10076 2723
rect 1661 2704 1667 2716
rect 2244 2697 2252 2703
rect 2484 2697 3596 2703
rect 3652 2697 4108 2703
rect 4132 2697 4220 2703
rect 4228 2697 4236 2703
rect 4244 2697 4284 2703
rect 4500 2697 4892 2703
rect 4964 2697 4972 2703
rect 5172 2697 6028 2703
rect 6612 2697 6620 2703
rect 6628 2697 7116 2703
rect 7172 2697 7196 2703
rect 7684 2697 8204 2703
rect 8436 2697 9516 2703
rect 9700 2697 9948 2703
rect 228 2677 243 2683
rect 237 2664 243 2677
rect 452 2677 700 2683
rect 916 2677 956 2683
rect 1140 2677 1148 2683
rect 1252 2677 1260 2683
rect 1652 2677 2012 2683
rect 2020 2677 2188 2683
rect 2260 2677 2460 2683
rect 2468 2677 2476 2683
rect 2484 2677 3212 2683
rect 3220 2677 3580 2683
rect 3604 2677 3996 2683
rect 4004 2677 4204 2683
rect 4308 2677 4323 2683
rect 4461 2677 4588 2683
rect 212 2657 220 2663
rect 676 2657 1356 2663
rect 1668 2657 1692 2663
rect 2004 2657 2092 2663
rect 2132 2657 2492 2663
rect 2756 2657 2892 2663
rect 2948 2657 3100 2663
rect 3572 2657 3788 2663
rect 3796 2657 3868 2663
rect 4461 2663 4467 2677
rect 4612 2677 5516 2683
rect 5620 2677 5628 2683
rect 5764 2677 5852 2683
rect 5860 2677 6188 2683
rect 6196 2677 7692 2683
rect 7860 2677 8108 2683
rect 8132 2677 8572 2683
rect 8628 2677 8716 2683
rect 8772 2677 8844 2683
rect 9012 2677 9724 2683
rect 9844 2677 10124 2683
rect 4116 2657 4467 2663
rect 4484 2657 5196 2663
rect 5492 2657 5612 2663
rect 5732 2657 5836 2663
rect 6164 2657 6268 2663
rect 6564 2657 6940 2663
rect 8244 2657 9212 2663
rect 9444 2657 9484 2663
rect 1364 2637 1788 2643
rect 1828 2637 3180 2643
rect 3188 2637 3356 2643
rect 3892 2637 4508 2643
rect 4564 2637 5324 2643
rect 5380 2637 5388 2643
rect 7460 2637 7468 2643
rect 7492 2637 7500 2643
rect 7668 2637 8860 2643
rect 228 2617 252 2623
rect 3140 2617 3868 2623
rect 3156 2597 3436 2603
rect 3588 2597 3660 2603
rect 4308 2597 5148 2603
rect 5789 2603 5795 2616
rect 5789 2597 5900 2603
rect 6644 2597 6828 2603
rect 7140 2597 7660 2603
rect 7924 2597 7932 2603
rect 8084 2597 8108 2603
rect 8452 2597 9148 2603
rect 9972 2597 10076 2603
rect 701 2584 707 2596
rect 1348 2577 1420 2583
rect 4468 2577 4492 2583
rect 6628 2577 6652 2583
rect 6788 2577 7004 2583
rect 7012 2577 8780 2583
rect 9636 2577 9852 2583
rect 1012 2557 1116 2563
rect 1124 2557 2748 2563
rect 2772 2557 3020 2563
rect 3028 2557 3420 2563
rect 3556 2557 3612 2563
rect 3844 2557 4092 2563
rect 4324 2557 4620 2563
rect 4756 2557 4764 2563
rect 6212 2557 7372 2563
rect 7380 2557 7420 2563
rect 7556 2557 7580 2563
rect 7860 2557 7884 2563
rect 8452 2557 8508 2563
rect 8548 2557 8588 2563
rect 8820 2557 8940 2563
rect 8948 2557 9148 2563
rect 6205 2544 6211 2556
rect 84 2537 92 2543
rect 436 2537 444 2543
rect 564 2537 572 2543
rect 756 2537 780 2543
rect 1236 2537 1244 2543
rect 1252 2537 1292 2543
rect 1796 2537 1804 2543
rect 1821 2537 1836 2543
rect 2004 2537 2028 2543
rect 2228 2537 2236 2543
rect 2356 2537 2364 2543
rect 2388 2537 2492 2543
rect 2804 2537 2812 2543
rect 3044 2537 3052 2543
rect 3076 2537 3644 2543
rect 4084 2537 4092 2543
rect 4116 2537 4380 2543
rect 4980 2537 4988 2543
rect 5012 2537 5324 2543
rect 5556 2537 5756 2543
rect 5972 2537 5980 2543
rect 6404 2537 6476 2543
rect 6756 2537 6764 2543
rect 7044 2537 7644 2543
rect 7892 2537 7980 2543
rect 8292 2537 8300 2543
rect 8404 2537 8476 2543
rect 8708 2537 8812 2543
rect 9252 2537 9676 2543
rect 9684 2537 9708 2543
rect 2260 2517 3372 2523
rect 4477 2523 4483 2536
rect 6957 2524 6963 2536
rect 4477 2517 4540 2523
rect 5092 2517 5596 2523
rect 5764 2517 5772 2523
rect 5780 2517 5916 2523
rect 8260 2517 8284 2523
rect 8772 2517 9020 2523
rect 9053 2523 9059 2536
rect 9245 2524 9251 2536
rect 9044 2517 9059 2523
rect 9220 2517 9228 2523
rect 9268 2517 9596 2523
rect 6189 2504 6195 2516
rect 452 2497 476 2503
rect 900 2497 1212 2503
rect 1220 2497 1228 2503
rect 1284 2497 1436 2503
rect 1812 2497 1820 2503
rect 2100 2497 2332 2503
rect 2548 2497 2796 2503
rect 2852 2497 2876 2503
rect 3636 2497 3644 2503
rect 4292 2497 4972 2503
rect 4980 2497 4988 2503
rect 5044 2497 5084 2503
rect 5972 2497 5980 2503
rect 6964 2497 6972 2503
rect 7172 2497 7180 2503
rect 7428 2497 7644 2503
rect 7652 2497 7676 2503
rect 7684 2497 9308 2503
rect 9316 2497 9692 2503
rect 212 2477 700 2483
rect 708 2477 796 2483
rect 916 2477 988 2483
rect 3396 2477 3420 2483
rect 5524 2477 5532 2483
rect 5540 2477 7148 2483
rect 7156 2477 7404 2483
rect 7412 2477 7420 2483
rect 8964 2477 9596 2483
rect 9620 2477 9868 2483
rect 5316 2457 5804 2463
rect 6100 2437 6108 2443
rect 6116 2437 6172 2443
rect 6180 2437 8748 2443
rect 8756 2437 8780 2443
rect 436 2397 460 2403
rect 2020 2397 2076 2403
rect 8084 2397 8124 2403
rect 468 2377 508 2383
rect 7188 2377 7276 2383
rect 3732 2357 3740 2363
rect 4692 2357 4707 2363
rect 5140 2357 5148 2363
rect 653 2344 659 2356
rect 244 2337 492 2343
rect 804 2337 1308 2343
rect 1604 2337 2172 2343
rect 2212 2337 3932 2343
rect 3940 2337 3948 2343
rect 4036 2337 4060 2343
rect 4244 2337 4396 2343
rect 5284 2337 5516 2343
rect 6036 2337 6620 2343
rect 7796 2337 7916 2343
rect 7956 2337 7964 2343
rect 7988 2337 8620 2343
rect 500 2317 652 2323
rect 660 2317 1004 2323
rect 1332 2317 1884 2323
rect 1908 2317 1980 2323
rect 1988 2317 2092 2323
rect 2436 2317 2460 2323
rect 2468 2317 2476 2323
rect 2852 2317 2860 2323
rect 3165 2317 3180 2323
rect 3492 2317 3500 2323
rect 3620 2317 5132 2323
rect 5156 2317 5292 2323
rect 6244 2317 6252 2323
rect 6260 2317 6684 2323
rect 6692 2317 6700 2323
rect 6740 2317 6908 2323
rect 7332 2317 7347 2323
rect 7908 2317 7916 2323
rect 7924 2317 8332 2323
rect 8852 2317 8956 2323
rect 8964 2317 9164 2323
rect 9277 2317 9283 2336
rect 9476 2317 9612 2323
rect 9901 2323 9907 2336
rect 9892 2317 9907 2323
rect 884 2297 1644 2303
rect 1780 2297 2028 2303
rect 2244 2297 2268 2303
rect 2276 2297 2508 2303
rect 2532 2297 4924 2303
rect 4948 2297 4956 2303
rect 5348 2297 5356 2303
rect 5428 2297 6236 2303
rect 6244 2297 6252 2303
rect 7140 2297 7164 2303
rect 7469 2303 7475 2316
rect 7469 2297 7564 2303
rect 7700 2297 8140 2303
rect 8148 2297 9180 2303
rect 9524 2297 9820 2303
rect 9828 2297 9836 2303
rect 660 2277 684 2283
rect 884 2277 1324 2283
rect 1556 2277 1564 2283
rect 1572 2277 1868 2283
rect 2180 2277 2188 2283
rect 2532 2277 2780 2283
rect 2804 2277 2940 2283
rect 3076 2277 3084 2283
rect 3220 2277 3484 2283
rect 3796 2277 4044 2283
rect 4372 2277 4412 2283
rect 4788 2277 4812 2283
rect 4916 2277 6700 2283
rect 6900 2277 6972 2283
rect 6980 2277 7308 2283
rect 7316 2277 7340 2283
rect 7668 2277 7772 2283
rect 8004 2277 8012 2283
rect 8324 2277 8412 2283
rect 8420 2277 8492 2283
rect 8996 2277 9148 2283
rect 9268 2277 9292 2283
rect 9492 2277 9596 2283
rect 9828 2277 9932 2283
rect 3485 2264 3491 2276
rect 500 2257 684 2263
rect 1108 2257 1132 2263
rect 1316 2257 1644 2263
rect 1652 2257 2108 2263
rect 2420 2257 3308 2263
rect 3364 2257 3372 2263
rect 3380 2257 3468 2263
rect 3940 2257 4748 2263
rect 6020 2257 6028 2263
rect 6036 2257 6140 2263
rect 6980 2257 7068 2263
rect 7092 2257 7132 2263
rect 7172 2257 7180 2263
rect 7860 2257 8396 2263
rect 8612 2257 9516 2263
rect 1620 2237 1628 2243
rect 1844 2237 2060 2243
rect 3581 2243 3587 2256
rect 3572 2237 3587 2243
rect 4420 2237 4636 2243
rect 4836 2237 5068 2243
rect 5428 2237 5724 2243
rect 5972 2237 6172 2243
rect 8068 2237 8156 2243
rect 8996 2237 9916 2243
rect 2660 2217 2668 2223
rect 3876 2217 4188 2223
rect 7940 2217 8172 2223
rect 1812 2197 1820 2203
rect 3140 2197 4972 2203
rect 5492 2197 5564 2203
rect 5796 2197 5868 2203
rect 6484 2197 6524 2203
rect 7364 2197 7404 2203
rect 7412 2197 7708 2203
rect 8420 2197 10236 2203
rect 708 2177 723 2183
rect 964 2177 972 2183
rect 1012 2177 1180 2183
rect 4013 2177 4060 2183
rect 308 2157 524 2163
rect 660 2157 956 2163
rect 964 2157 1388 2163
rect 1652 2157 1660 2163
rect 1684 2157 1772 2163
rect 2580 2157 2908 2163
rect 3012 2157 3020 2163
rect 4013 2163 4019 2177
rect 8564 2177 8636 2183
rect 3604 2157 4019 2163
rect 4036 2157 4572 2163
rect 4580 2157 4604 2163
rect 5620 2157 6092 2163
rect 6372 2157 7100 2163
rect 7124 2157 7132 2163
rect 7140 2157 7276 2163
rect 7876 2157 8588 2163
rect 8708 2157 8924 2163
rect 9012 2157 9132 2163
rect 9476 2157 9484 2163
rect 100 2137 220 2143
rect 228 2137 316 2143
rect 932 2137 972 2143
rect 980 2137 1004 2143
rect 1268 2137 2428 2143
rect 2436 2137 3532 2143
rect 3540 2137 3564 2143
rect 3828 2137 3836 2143
rect 3940 2137 4044 2143
rect 4068 2137 4268 2143
rect 4308 2137 4316 2143
rect 4324 2137 4476 2143
rect 4500 2137 4540 2143
rect 4548 2137 4556 2143
rect 4804 2137 4812 2143
rect 6388 2137 7020 2143
rect 7060 2137 7404 2143
rect 7972 2137 8124 2143
rect 8676 2137 8691 2143
rect 8772 2137 8988 2143
rect 9140 2137 9244 2143
rect 9252 2137 9804 2143
rect 10068 2137 10108 2143
rect 8365 2124 8371 2136
rect 676 2117 2252 2123
rect 2260 2117 4492 2123
rect 4500 2117 4508 2123
rect 5732 2117 5740 2123
rect 5748 2117 5852 2123
rect 5892 2117 6588 2123
rect 6884 2117 7484 2123
rect 9037 2123 9043 2136
rect 9037 2117 9180 2123
rect 9428 2117 9884 2123
rect 1332 2097 1548 2103
rect 2324 2097 2908 2103
rect 2996 2097 3916 2103
rect 3924 2097 4508 2103
rect 5060 2097 5164 2103
rect 5732 2097 5740 2103
rect 5956 2097 6156 2103
rect 6820 2097 6828 2103
rect 7044 2097 7244 2103
rect 7252 2097 7260 2103
rect 7396 2097 7548 2103
rect 7796 2097 7916 2103
rect 8132 2097 8284 2103
rect 8372 2097 8380 2103
rect 9156 2097 9164 2103
rect 2061 2084 2067 2096
rect 7693 2084 7699 2096
rect 1172 2077 1548 2083
rect 3172 2077 3244 2083
rect 4036 2077 4572 2083
rect 6388 2077 6396 2083
rect 6404 2077 7212 2083
rect 4948 2057 5388 2063
rect 2685 1964 2691 2056
rect 3396 2017 3404 2023
rect 8484 2017 8492 2023
rect 7476 1977 8332 1983
rect 964 1957 972 1963
rect 1012 1957 2012 1963
rect 2228 1957 2236 1963
rect 3380 1957 3404 1963
rect 3828 1957 3836 1963
rect 3844 1957 3852 1963
rect 7636 1957 7660 1963
rect 8356 1957 8364 1963
rect 9236 1957 9244 1963
rect 868 1937 988 1943
rect 996 1937 1827 1943
rect 292 1917 1628 1923
rect 1796 1917 1804 1923
rect 1821 1923 1827 1937
rect 1892 1937 1900 1943
rect 2132 1937 2332 1943
rect 2340 1937 2476 1943
rect 2708 1937 3148 1943
rect 3220 1937 3628 1943
rect 4740 1937 4828 1943
rect 6116 1937 6796 1943
rect 6820 1937 8588 1943
rect 8804 1937 8835 1943
rect 4285 1924 4291 1936
rect 4493 1924 4499 1936
rect 1821 1917 2252 1923
rect 2260 1917 2268 1923
rect 2452 1917 2780 1923
rect 2836 1917 3004 1923
rect 4820 1917 4844 1923
rect 4996 1917 5020 1923
rect 5700 1917 5724 1923
rect 5924 1917 5948 1923
rect 6228 1917 6684 1923
rect 6692 1917 6700 1923
rect 6788 1917 6796 1923
rect 6804 1917 7660 1923
rect 7828 1917 7884 1923
rect 7908 1917 8124 1923
rect 8132 1917 8348 1923
rect 8804 1917 8812 1923
rect 8829 1923 8835 1937
rect 9156 1937 9452 1943
rect 9460 1937 9868 1943
rect 8829 1917 8988 1923
rect 212 1897 524 1903
rect 532 1897 2668 1903
rect 3172 1897 3180 1903
rect 3188 1897 5180 1903
rect 660 1877 668 1883
rect 852 1877 860 1883
rect 964 1877 988 1883
rect 1204 1877 2940 1883
rect 2948 1877 3196 1883
rect 3604 1877 4348 1883
rect 4452 1877 4476 1883
rect 301 1864 307 1876
rect 637 1864 643 1876
rect 861 1864 867 1876
rect 4493 1864 4499 1897
rect 5940 1897 5980 1903
rect 6772 1897 6780 1903
rect 6820 1897 7372 1903
rect 7380 1897 7628 1903
rect 8132 1897 8812 1903
rect 9396 1897 9660 1903
rect 9892 1897 9900 1903
rect 7677 1884 7683 1896
rect 4516 1877 4812 1883
rect 4820 1877 5020 1883
rect 5268 1877 5324 1883
rect 5476 1877 5491 1883
rect 5716 1877 6300 1883
rect 6500 1877 6620 1883
rect 6692 1877 6716 1883
rect 7380 1877 7676 1883
rect 7892 1877 7900 1883
rect 7908 1877 8908 1883
rect 8916 1877 9244 1883
rect 9428 1877 9564 1883
rect 10109 1883 10115 1896
rect 10100 1877 10115 1883
rect 1172 1857 1308 1863
rect 1316 1857 1420 1863
rect 1620 1857 1756 1863
rect 1780 1857 1820 1863
rect 1844 1857 2476 1863
rect 2660 1857 2684 1863
rect 2980 1857 3020 1863
rect 3188 1857 3372 1863
rect 3924 1857 4316 1863
rect 4708 1857 4716 1863
rect 6052 1857 6684 1863
rect 6708 1857 7036 1863
rect 8036 1857 8556 1863
rect 8564 1857 8572 1863
rect 1348 1837 1580 1843
rect 4148 1837 4300 1843
rect 4308 1837 4332 1843
rect 4356 1837 4524 1843
rect 5956 1837 6076 1843
rect 7805 1824 7811 1843
rect 7972 1837 8044 1843
rect 8324 1837 8444 1843
rect 10260 1837 10339 1843
rect 244 1817 252 1823
rect 1636 1817 1996 1823
rect 2948 1817 3004 1823
rect 4276 1817 4284 1823
rect 5828 1817 6156 1823
rect 8820 1817 8940 1823
rect 8948 1817 9132 1823
rect 9684 1817 9804 1823
rect 996 1797 1116 1803
rect 1140 1797 1340 1803
rect 1364 1797 1644 1803
rect 1892 1797 1900 1803
rect 5492 1797 5628 1803
rect 7652 1797 7788 1803
rect 7796 1797 7804 1803
rect 9908 1797 10220 1803
rect 3668 1777 4092 1783
rect 4964 1777 5036 1783
rect 6996 1777 7212 1783
rect 7684 1777 7692 1783
rect 68 1757 92 1763
rect 436 1757 444 1763
rect 676 1757 716 1763
rect 724 1757 956 1763
rect 1444 1757 1612 1763
rect 2468 1757 2476 1763
rect 2804 1757 3036 1763
rect 3044 1757 3212 1763
rect 3412 1757 3900 1763
rect 4260 1757 4300 1763
rect 4948 1757 5148 1763
rect 5204 1757 5900 1763
rect 6692 1757 8364 1763
rect 8372 1757 8380 1763
rect 8388 1757 8540 1763
rect 8756 1757 9020 1763
rect 653 1744 659 1756
rect 2701 1744 2707 1756
rect 84 1737 524 1743
rect 772 1737 844 1743
rect 1188 1737 1212 1743
rect 1876 1737 2012 1743
rect 2020 1737 2044 1743
rect 2260 1737 2540 1743
rect 2900 1737 4044 1743
rect 4052 1737 4460 1743
rect 4557 1743 4563 1756
rect 4548 1737 4563 1743
rect 4756 1737 4796 1743
rect 4813 1737 4988 1743
rect 676 1717 748 1723
rect 756 1717 1260 1723
rect 1796 1717 1820 1723
rect 2036 1717 2092 1723
rect 2276 1717 2652 1723
rect 2660 1717 2796 1723
rect 2989 1717 3228 1723
rect 756 1697 1548 1703
rect 2532 1697 2700 1703
rect 2989 1703 2995 1717
rect 3476 1717 3484 1723
rect 3588 1717 3692 1723
rect 3908 1717 3916 1723
rect 4813 1723 4819 1737
rect 5268 1737 5788 1743
rect 5796 1737 5836 1743
rect 5876 1737 6124 1743
rect 6132 1737 6140 1743
rect 6292 1737 6444 1743
rect 7284 1737 7292 1743
rect 7300 1737 7452 1743
rect 7796 1737 7804 1743
rect 7812 1737 8140 1743
rect 8276 1737 8588 1743
rect 8596 1737 8956 1743
rect 9453 1743 9459 1756
rect 9444 1737 9459 1743
rect 7021 1724 7027 1736
rect 4804 1717 4819 1723
rect 5428 1717 5436 1723
rect 5444 1717 6684 1723
rect 7604 1717 7804 1723
rect 7837 1717 7852 1723
rect 7908 1717 7916 1723
rect 2948 1697 2995 1703
rect 3108 1697 3372 1703
rect 3380 1697 3388 1703
rect 3476 1697 3484 1703
rect 3700 1697 5148 1703
rect 6708 1697 6716 1703
rect 6788 1697 7164 1703
rect 7220 1697 7452 1703
rect 7460 1697 7468 1703
rect 7732 1697 8140 1703
rect 8148 1697 8156 1703
rect 9220 1697 9228 1703
rect 9940 1697 10076 1703
rect 2020 1677 2028 1683
rect 2036 1677 3043 1683
rect 436 1657 444 1663
rect 1124 1657 1580 1663
rect 3037 1663 3043 1677
rect 3364 1677 3692 1683
rect 3860 1677 4460 1683
rect 4468 1677 4476 1683
rect 5892 1677 5916 1683
rect 5924 1677 7244 1683
rect 7476 1677 8300 1683
rect 3037 1657 3676 1663
rect 5220 1657 5676 1663
rect 6244 1657 6444 1663
rect 8068 1657 8748 1663
rect 2452 1637 3676 1643
rect 3684 1637 4540 1643
rect 4772 1637 4780 1643
rect 6516 1637 7788 1643
rect 1844 1617 1852 1623
rect 1636 1597 1644 1603
rect 4932 1577 4940 1583
rect 212 1557 284 1563
rect 292 1557 428 1563
rect 948 1557 972 1563
rect 324 1537 428 1543
rect 436 1537 620 1543
rect 2084 1537 2092 1543
rect 2340 1537 2348 1543
rect 2532 1537 2540 1543
rect 3940 1537 4076 1543
rect 4516 1537 5164 1543
rect 6708 1537 6924 1543
rect 8468 1537 8524 1543
rect 9748 1537 9868 1543
rect 7245 1524 7251 1536
rect 228 1517 524 1523
rect 532 1517 540 1523
rect 756 1517 940 1523
rect 1556 1517 1772 1523
rect 1780 1517 3356 1523
rect 3924 1517 4508 1523
rect 4580 1517 4588 1523
rect 4964 1517 5532 1523
rect 5540 1517 5788 1523
rect 6468 1517 6492 1523
rect 6804 1517 7228 1523
rect 7460 1517 7475 1523
rect 9316 1517 9324 1523
rect 9412 1517 9436 1523
rect 9764 1517 10060 1523
rect 5885 1504 5891 1516
rect 8893 1504 8899 1516
rect 100 1497 1148 1503
rect 1620 1497 2700 1503
rect 2708 1497 3324 1503
rect 3588 1497 4780 1503
rect 5012 1497 5452 1503
rect 6804 1497 6812 1503
rect 7028 1497 7468 1503
rect 7700 1497 7964 1503
rect 8964 1497 9772 1503
rect 9796 1497 9980 1503
rect 8237 1484 8243 1496
rect 548 1477 556 1483
rect 644 1477 652 1483
rect 772 1477 876 1483
rect 980 1477 988 1483
rect 1332 1477 1436 1483
rect 1652 1477 1660 1483
rect 2308 1477 2332 1483
rect 2564 1477 2908 1483
rect 2916 1477 3020 1483
rect 3140 1477 3164 1483
rect 3380 1477 3452 1483
rect 3652 1477 3820 1483
rect 4148 1477 4156 1483
rect 4308 1477 4316 1483
rect 5572 1477 5724 1483
rect 5828 1477 5900 1483
rect 6052 1477 6460 1483
rect 6468 1477 7884 1483
rect 8996 1477 9004 1483
rect 9412 1477 9427 1483
rect 9604 1477 9740 1483
rect 5341 1464 5347 1476
rect 436 1457 2764 1463
rect 3396 1457 3596 1463
rect 3972 1457 4476 1463
rect 5796 1457 6060 1463
rect 6308 1457 6684 1463
rect 6692 1457 6700 1463
rect 6724 1457 6924 1463
rect 7252 1457 7292 1463
rect 7876 1457 8012 1463
rect 8052 1457 9308 1463
rect 9332 1457 9564 1463
rect 9828 1457 9852 1463
rect 852 1437 876 1443
rect 2356 1437 2716 1443
rect 8788 1437 8796 1443
rect 8980 1437 9180 1443
rect 676 1417 684 1423
rect 1108 1417 1116 1423
rect 2260 1417 2268 1423
rect 2285 1417 3628 1423
rect 2285 1403 2291 1417
rect 4724 1417 4748 1423
rect 5668 1417 7020 1423
rect 9172 1417 9212 1423
rect 1588 1397 2291 1403
rect 3428 1397 3468 1403
rect 4772 1397 4780 1403
rect 8452 1397 8524 1403
rect 9540 1397 9596 1403
rect 1757 1377 2316 1383
rect 740 1357 1212 1363
rect 1757 1363 1763 1377
rect 2324 1377 2572 1383
rect 2916 1377 2924 1383
rect 4548 1377 4556 1383
rect 6932 1377 7004 1383
rect 7380 1377 7388 1383
rect 7668 1377 7868 1383
rect 8964 1377 9612 1383
rect 1684 1357 1763 1363
rect 4244 1357 4316 1363
rect 5028 1357 5036 1363
rect 6708 1357 8364 1363
rect 68 1337 92 1343
rect 324 1337 428 1343
rect 548 1337 732 1343
rect 2020 1337 2028 1343
rect 2100 1337 2476 1343
rect 2484 1337 2780 1343
rect 2788 1337 2876 1343
rect 2884 1337 2988 1343
rect 4468 1337 4668 1343
rect 4676 1337 5228 1343
rect 5364 1337 5452 1343
rect 5812 1337 5820 1343
rect 5908 1337 5916 1343
rect 6068 1337 7404 1343
rect 7412 1337 7596 1343
rect 7604 1337 8476 1343
rect 8820 1337 8828 1343
rect 9188 1337 9228 1343
rect 9236 1337 9244 1343
rect 9492 1337 9692 1343
rect 9876 1337 10012 1343
rect 3773 1324 3779 1336
rect 852 1317 876 1323
rect 884 1317 2444 1323
rect 2548 1317 2556 1323
rect 4532 1317 5356 1323
rect 5492 1317 6348 1323
rect 6580 1317 6588 1323
rect 7044 1317 7132 1323
rect 7588 1317 7596 1323
rect 7620 1317 7692 1323
rect 7924 1317 7932 1323
rect 8372 1317 9244 1323
rect 9252 1317 9260 1323
rect 100 1297 108 1303
rect 292 1297 300 1303
rect 308 1297 652 1303
rect 884 1297 1308 1303
rect 1428 1297 1564 1303
rect 2116 1297 2124 1303
rect 2564 1297 2572 1303
rect 2772 1297 2860 1303
rect 3124 1297 3148 1303
rect 4580 1297 4684 1303
rect 4692 1297 4700 1303
rect 6276 1297 7900 1303
rect 7956 1297 8780 1303
rect 8804 1297 9132 1303
rect 9140 1297 9404 1303
rect 5213 1284 5219 1296
rect 948 1277 2972 1283
rect 5460 1277 5676 1283
rect 5684 1277 5884 1283
rect 5892 1277 6348 1283
rect 6452 1277 6540 1283
rect 6564 1277 6796 1283
rect 7604 1277 8348 1283
rect 8356 1277 8380 1283
rect 9028 1277 9676 1283
rect 980 1257 988 1263
rect 5812 1257 5820 1263
rect 5892 1257 5900 1263
rect 6260 1257 6268 1263
rect 7412 1257 8124 1263
rect 8276 1257 8684 1263
rect 564 1237 892 1243
rect 900 1237 972 1243
rect 6820 1197 6828 1203
rect 10036 1197 10060 1203
rect 1380 1177 1836 1183
rect 2724 1177 3852 1183
rect 4052 1177 4076 1183
rect 4916 1177 4924 1183
rect 2676 1157 2684 1163
rect 3332 1157 3644 1163
rect 4452 1157 4556 1163
rect 4564 1157 4652 1163
rect 4660 1157 5020 1163
rect 5028 1157 5164 1163
rect 8020 1157 8236 1163
rect 8909 1157 9244 1163
rect 1565 1144 1571 1156
rect 660 1137 908 1143
rect 1636 1137 2876 1143
rect 2884 1137 3372 1143
rect 3380 1137 3564 1143
rect 3572 1137 4204 1143
rect 4212 1137 4284 1143
rect 5828 1137 6380 1143
rect 6628 1137 6636 1143
rect 7492 1137 7804 1143
rect 8276 1137 8492 1143
rect 8909 1143 8915 1157
rect 8708 1137 8915 1143
rect 9140 1137 9916 1143
rect 244 1117 444 1123
rect 756 1117 860 1123
rect 868 1117 972 1123
rect 980 1117 3404 1123
rect 3412 1117 3484 1123
rect 3492 1117 3820 1123
rect 3828 1117 4236 1123
rect 4532 1117 4540 1123
rect 4548 1117 4588 1123
rect 5220 1117 5452 1123
rect 5460 1117 5484 1123
rect 5956 1117 6140 1123
rect 6148 1117 6156 1123
rect 6500 1117 7036 1123
rect 7716 1117 7724 1123
rect 8596 1117 9820 1123
rect 228 1097 236 1103
rect 948 1097 1116 1103
rect 1172 1097 1196 1103
rect 1348 1097 1356 1103
rect 1396 1097 2012 1103
rect 2084 1097 2092 1103
rect 2676 1097 2844 1103
rect 3092 1097 4492 1103
rect 4500 1097 4684 1103
rect 4788 1097 4940 1103
rect 4948 1097 5004 1103
rect 5348 1097 5356 1103
rect 5364 1097 6316 1103
rect 6324 1097 6396 1103
rect 6532 1097 6956 1103
rect 7268 1097 7708 1103
rect 7716 1097 7820 1103
rect 2893 1084 2899 1096
rect 9469 1084 9475 1096
rect 212 1077 236 1083
rect 980 1077 1644 1083
rect 1764 1077 1772 1083
rect 2004 1077 2012 1083
rect 2436 1077 2444 1083
rect 3556 1077 3644 1083
rect 3844 1077 4188 1083
rect 5364 1077 5372 1083
rect 5412 1077 5468 1083
rect 5860 1077 5900 1083
rect 5908 1077 6620 1083
rect 6628 1077 7900 1083
rect 8468 1077 8476 1083
rect 9828 1077 9916 1083
rect 765 1064 771 1076
rect 4797 1064 4803 1076
rect 868 1057 2108 1063
rect 2116 1057 3196 1063
rect 3588 1057 3596 1063
rect 3652 1057 3996 1063
rect 5044 1057 7068 1063
rect 7076 1057 7100 1063
rect 7252 1057 7388 1063
rect 7492 1057 7852 1063
rect 8356 1057 8812 1063
rect 8820 1057 8924 1063
rect 8932 1057 9148 1063
rect 9412 1057 9644 1063
rect 9700 1057 9820 1063
rect 9389 1044 9395 1056
rect 212 1037 524 1043
rect 916 1037 2252 1043
rect 2468 1037 2732 1043
rect 4052 1037 4428 1043
rect 4436 1037 4636 1043
rect 5332 1037 5340 1043
rect 5604 1037 5932 1043
rect 6964 1037 7212 1043
rect 8292 1037 8508 1043
rect 1620 1017 1628 1023
rect 2004 1017 2076 1023
rect 2692 1017 3772 1023
rect 3780 1017 3852 1023
rect 5364 1017 5580 1023
rect 8020 1017 8076 1023
rect 484 997 684 1003
rect 1780 997 2428 1003
rect 2484 997 3116 1003
rect 3540 997 3548 1003
rect 4740 997 4812 1003
rect 8100 997 8124 1003
rect 9261 1003 9267 1016
rect 9261 997 9420 1003
rect 3613 984 3619 996
rect 653 977 924 983
rect 653 964 659 977
rect 1076 977 1196 983
rect 1412 977 1836 983
rect 2068 977 2236 983
rect 2260 977 2268 983
rect 2500 977 2924 983
rect 2948 977 3612 983
rect 6756 977 7452 983
rect 7460 977 9155 983
rect 9149 964 9155 977
rect 1268 957 1532 963
rect 1780 957 1868 963
rect 2292 957 2524 963
rect 2532 957 2540 963
rect 2740 957 2972 963
rect 5636 957 5676 963
rect 6100 957 6684 963
rect 6772 957 6892 963
rect 7124 957 7132 963
rect 7140 957 8300 963
rect 8308 957 8348 963
rect 8564 957 8572 963
rect 9156 957 9244 963
rect 9588 957 9612 963
rect 3197 944 3203 956
rect 436 937 860 943
rect 1316 937 1324 943
rect 1332 937 2940 943
rect 3380 937 3404 943
rect 3748 937 3948 943
rect 3988 937 4060 943
rect 4468 937 4652 943
rect 4660 937 4860 943
rect 5108 937 5212 943
rect 5220 937 5548 943
rect 5892 937 5900 943
rect 6132 937 6140 943
rect 6356 937 6540 943
rect 6564 937 6579 943
rect 7140 937 7244 943
rect 7668 937 7692 943
rect 7924 937 7996 943
rect 8292 937 9820 943
rect 516 917 892 923
rect 1124 917 1404 923
rect 1652 917 1660 923
rect 1668 917 2652 923
rect 2772 917 3404 923
rect 4180 917 4188 923
rect 4196 917 4892 923
rect 5876 917 7452 923
rect 7460 917 8028 923
rect 8692 917 9164 923
rect 9172 917 9228 923
rect 9604 917 9868 923
rect 436 897 972 903
rect 1076 897 1116 903
rect 1556 897 3084 903
rect 3092 897 3100 903
rect 3956 897 3964 903
rect 4196 897 4924 903
rect 6132 897 6268 903
rect 6276 897 6284 903
rect 7156 897 7164 903
rect 7172 897 7932 903
rect 7988 897 8236 903
rect 8548 897 8556 903
rect 8868 897 8876 903
rect 8884 897 8908 903
rect 9316 897 9820 903
rect 9828 897 10108 903
rect 4189 884 4195 896
rect 1348 877 1724 883
rect 1748 877 3180 883
rect 3188 877 4028 883
rect 4436 877 4524 883
rect 5220 877 5228 883
rect 5780 877 5788 883
rect 5892 877 6092 883
rect 6100 877 6140 883
rect 7252 877 7260 883
rect 9828 877 9900 883
rect 2900 857 3628 863
rect 4964 857 5100 863
rect 5108 857 5804 863
rect 5812 857 6156 863
rect 564 837 1596 843
rect 1604 837 1676 843
rect 4260 837 4748 843
rect 5796 837 7836 843
rect 7844 837 8316 843
rect 8468 837 8476 843
rect 3101 824 3107 836
rect 4708 797 4716 803
rect 5780 797 5804 803
rect 237 784 243 796
rect 5236 777 5340 783
rect 5348 777 5596 783
rect 7588 777 7596 783
rect 6724 757 6732 763
rect 7556 757 7660 763
rect 420 737 428 743
rect 436 737 956 743
rect 2644 737 2716 743
rect 4644 737 4652 743
rect 5108 737 5340 743
rect 7012 737 7020 743
rect 7108 737 9500 743
rect 9508 737 9644 743
rect 1533 724 1539 736
rect 6493 724 6499 736
rect 10093 724 10099 736
rect 877 717 892 723
rect 1652 717 1740 723
rect 1956 717 1964 723
rect 2052 717 3164 723
rect 3172 717 3388 723
rect 3396 717 4732 723
rect 6724 717 8028 723
rect 8036 717 8044 723
rect 8100 717 8108 723
rect 8692 717 8700 723
rect 8724 717 8892 723
rect 9332 717 9436 723
rect 9540 717 9555 723
rect 9844 717 9884 723
rect 10180 717 10188 723
rect 1956 697 2028 703
rect 3092 697 4492 703
rect 4900 697 4908 703
rect 4916 697 5132 703
rect 5540 697 5548 703
rect 5556 697 5820 703
rect 5828 697 6012 703
rect 6692 697 6700 703
rect 7044 697 7916 703
rect 8484 697 8924 703
rect 973 684 979 696
rect 1741 684 1747 696
rect 9885 684 9891 696
rect 429 677 444 683
rect 548 677 556 683
rect 1108 677 1308 683
rect 1316 677 1324 683
rect 1540 677 1660 683
rect 2036 677 2044 683
rect 2628 677 2636 683
rect 2676 677 3084 683
rect 3188 677 3388 683
rect 3396 677 3404 683
rect 3732 677 4172 683
rect 4180 677 4412 683
rect 4420 677 4636 683
rect 5092 677 5212 683
rect 5460 677 5468 683
rect 5476 677 6476 683
rect 6484 677 7292 683
rect 7364 677 7372 683
rect 7700 677 7820 683
rect 7908 677 8684 683
rect 8692 677 9004 683
rect 9012 677 9020 683
rect 9172 677 9532 683
rect 5085 664 5091 676
rect 948 657 956 663
rect 964 657 1740 663
rect 2484 657 3820 663
rect 3828 657 3836 663
rect 5220 657 5228 663
rect 5236 657 5628 663
rect 6100 657 6124 663
rect 7236 657 9660 663
rect 6244 637 6284 643
rect 8244 637 8252 643
rect 8260 637 8332 643
rect 8788 637 8796 643
rect 2205 624 2211 636
rect 964 617 988 623
rect 2628 617 2700 623
rect 5860 617 5884 623
rect 7748 617 9196 623
rect 84 597 92 603
rect 1156 597 1356 603
rect 2404 597 2460 603
rect 3668 597 3788 603
rect 4644 597 4716 603
rect 7588 597 8316 603
rect 9044 597 9148 603
rect 1325 577 1580 583
rect 1325 564 1331 577
rect 2573 577 2748 583
rect 212 557 636 563
rect 660 557 684 563
rect 1108 557 1132 563
rect 1572 557 1612 563
rect 2020 557 2236 563
rect 2573 563 2579 577
rect 3364 577 3820 583
rect 4100 577 4684 583
rect 7748 577 7804 583
rect 8004 577 8012 583
rect 8020 577 8092 583
rect 8724 577 9180 583
rect 9572 577 9852 583
rect 6397 564 6403 576
rect 2564 557 2579 563
rect 2964 557 2979 563
rect 3108 557 3116 563
rect 3572 557 3660 563
rect 3764 557 3948 563
rect 3956 557 4444 563
rect 5460 557 5628 563
rect 7188 557 7500 563
rect 861 544 867 556
rect 1885 544 1891 556
rect 2333 544 2339 556
rect 3677 544 3683 556
rect 900 537 1068 543
rect 1076 537 1884 543
rect 2340 537 3132 543
rect 3181 537 3196 543
rect 3348 537 3420 543
rect 3972 537 4012 543
rect 4228 537 4268 543
rect 4548 537 4796 543
rect 4948 537 5228 543
rect 5236 537 5260 543
rect 5588 537 5596 543
rect 6580 537 6620 543
rect 6996 537 7068 543
rect 7284 537 7292 543
rect 7332 537 7388 543
rect 7684 537 7932 543
rect 8260 537 8300 543
rect 8477 543 8483 556
rect 9805 544 9811 556
rect 8468 537 8483 543
rect 9828 537 9996 543
rect 10100 537 10115 543
rect 308 517 316 523
rect 324 517 1004 523
rect 1844 517 2076 523
rect 2308 517 2412 523
rect 2420 517 2460 523
rect 3517 523 3523 536
rect 3517 517 3580 523
rect 3773 523 3779 536
rect 3773 517 3820 523
rect 4205 523 4211 536
rect 3828 517 4460 523
rect 4365 504 4371 517
rect 4484 517 4556 523
rect 5156 517 5948 523
rect 5956 517 6172 523
rect 6980 517 8780 523
rect 9364 517 9388 523
rect 10116 517 10172 523
rect 308 497 316 503
rect 324 497 620 503
rect 628 497 1948 503
rect 2340 497 2668 503
rect 4100 497 4300 503
rect 5124 497 5148 503
rect 5764 497 5788 503
rect 5796 497 6972 503
rect 6980 497 8428 503
rect 8932 497 9804 503
rect 957 477 1164 483
rect 957 463 963 477
rect 1540 477 1788 483
rect 1796 477 1820 483
rect 1876 477 2892 483
rect 3316 477 4124 483
rect 5252 477 5676 483
rect 5684 477 5868 483
rect 6964 477 7052 483
rect 8132 477 8716 483
rect 900 457 963 463
rect 1572 457 1580 463
rect 4708 457 5100 463
rect 5556 457 5612 463
rect 5620 457 5708 463
rect 5716 457 6044 463
rect 2212 437 2444 443
rect 2452 437 2476 443
rect 4388 437 4460 443
rect 4468 437 4604 443
rect 4612 437 4940 443
rect 5780 437 6332 443
rect 7540 437 7644 443
rect 7652 437 8956 443
rect 7444 417 8492 423
rect 3316 397 3324 403
rect 6596 397 6636 403
rect 7060 377 8732 383
rect 2196 357 2268 363
rect 3540 357 3980 363
rect 4948 357 4956 363
rect 7956 357 8012 363
rect 1956 337 2844 343
rect 3780 337 3836 343
rect 3844 337 4716 343
rect 5188 337 5868 343
rect 5876 337 5900 343
rect 7204 337 7708 343
rect 7796 337 8172 343
rect 8180 337 8252 343
rect 8948 337 9148 343
rect 1069 324 1075 336
rect 6237 324 6243 336
rect 8269 324 8275 336
rect 8925 324 8931 336
rect 9501 324 9507 336
rect 420 317 428 323
rect 868 317 876 323
rect 1300 317 1836 323
rect 2660 317 2716 323
rect 2740 317 4156 323
rect 4724 317 5356 323
rect 5364 317 5388 323
rect 5636 317 5852 323
rect 6084 317 6236 323
rect 6292 317 6492 323
rect 7076 317 7196 323
rect 7300 317 7308 323
rect 7684 317 8268 323
rect 8324 317 8700 323
rect 9732 317 9747 323
rect 9764 317 10044 323
rect 7485 304 7491 316
rect 196 297 652 303
rect 1732 297 1740 303
rect 2756 297 3500 303
rect 3508 297 3964 303
rect 4612 297 4940 303
rect 4948 297 5132 303
rect 5140 297 5148 303
rect 7716 297 7740 303
rect 7924 297 7948 303
rect 8276 297 9820 303
rect 5405 284 5411 296
rect 628 277 940 283
rect 1268 277 1276 283
rect 1748 277 2860 283
rect 3092 277 3116 283
rect 3316 277 3532 283
rect 3828 277 4412 283
rect 4708 277 4716 283
rect 5188 277 5196 283
rect 5428 277 6284 283
rect 6532 277 6668 283
rect 6852 277 7068 283
rect 7284 277 7292 283
rect 7300 277 8172 283
rect 8260 277 8268 283
rect 8292 277 8844 283
rect 8932 277 8947 283
rect 9316 277 9500 283
rect 9700 277 9708 283
rect 9716 277 9740 283
rect 10020 277 10140 283
rect 2957 264 2963 276
rect 420 257 764 263
rect 772 257 988 263
rect 1076 257 1084 263
rect 1092 257 1756 263
rect 1764 257 2476 263
rect 2557 257 2652 263
rect 148 237 268 243
rect 756 237 1420 243
rect 2052 237 2076 243
rect 2557 243 2563 257
rect 5204 257 8860 263
rect 8868 257 8876 263
rect 8884 257 9820 263
rect 2388 237 2563 243
rect 2580 237 2716 243
rect 2740 237 3308 243
rect 5476 237 6076 243
rect 6868 237 7036 243
rect 7252 237 7740 243
rect 8116 237 8652 243
rect 8788 237 8956 243
rect 8980 237 10028 243
rect 932 217 1148 223
rect 1828 217 3372 223
rect 6020 217 6028 223
rect 6852 217 6908 223
rect 8493 217 9532 223
rect 8493 204 8499 217
rect 308 197 492 203
rect 1460 197 1548 203
rect 1588 197 1852 203
rect 2052 197 2444 203
rect 3716 197 3804 203
rect 8756 197 9596 203
rect 772 177 860 183
rect 2356 177 3148 183
rect 4372 177 4396 183
rect 4628 177 5315 183
rect 100 157 140 163
rect 1396 157 1628 163
rect 2180 157 2812 163
rect 3188 157 3196 163
rect 4196 157 5068 163
rect 5076 157 5100 163
rect 5108 157 5116 163
rect 5309 163 5315 177
rect 7236 177 7260 183
rect 7860 177 8316 183
rect 8356 177 8988 183
rect 9156 177 9171 183
rect 9252 177 9356 183
rect 9444 177 9820 183
rect 9892 177 9964 183
rect 5309 157 5548 163
rect 5796 157 5964 163
rect 6644 157 8508 163
rect 8532 157 8636 163
rect 8916 157 9036 163
rect 9492 157 9756 163
rect 564 137 700 143
rect 708 137 1532 143
rect 1908 137 1980 143
rect 1988 137 2156 143
rect 3700 137 3868 143
rect 3876 137 3948 143
rect 4084 137 4092 143
rect 4644 137 4700 143
rect 6020 137 6028 143
rect 6788 137 7324 143
rect 7428 137 7436 143
rect 7700 137 8012 143
rect 8036 137 8067 143
rect 1012 117 2732 123
rect 4100 117 4412 123
rect 4420 117 4604 123
rect 4612 117 4652 123
rect 4884 117 5100 123
rect 5348 117 5564 123
rect 5572 117 6028 123
rect 7524 117 7676 123
rect 8061 123 8067 137
rect 8116 137 8131 143
rect 8125 124 8131 137
rect 8148 137 8348 143
rect 8436 137 8940 143
rect 8948 137 9020 143
rect 9028 137 9692 143
rect 9700 137 9708 143
rect 9876 137 10012 143
rect 8061 117 8076 123
rect 8516 117 8588 123
rect 9524 117 9676 123
rect 1220 97 1468 103
rect 3396 97 3404 103
rect 3604 97 3628 103
rect 3636 97 4172 103
rect 4180 97 4188 103
rect 4404 97 4412 103
rect 4420 97 4860 103
rect 5556 97 5788 103
rect 6036 97 7676 103
rect 8596 97 8748 103
rect 8756 97 9196 103
rect 9476 97 9852 103
rect 10020 97 10035 103
rect 3860 77 4076 83
rect 6020 77 6236 83
rect 2692 17 2700 23
rect 4052 17 4076 23
rect 4692 17 4700 23
<< m4contact >>
rect 5180 7616 5188 7624
rect 6092 7556 6100 7564
rect 4268 7536 4276 7544
rect 5020 7536 5028 7544
rect 6172 7536 6180 7544
rect 9644 7536 9652 7544
rect 316 7516 324 7524
rect 572 7516 580 7524
rect 1116 7516 1124 7524
rect 1436 7516 1444 7524
rect 2588 7516 2596 7524
rect 2732 7516 2740 7524
rect 4220 7516 4228 7524
rect 4812 7516 4820 7524
rect 5404 7516 5412 7524
rect 6588 7516 6596 7524
rect 9820 7516 9828 7524
rect 3484 7496 3492 7504
rect 5836 7496 5844 7504
rect 7676 7496 7684 7504
rect 8220 7496 8228 7504
rect 8412 7496 8420 7504
rect 9500 7496 9508 7504
rect 9548 7496 9556 7504
rect 9916 7496 9924 7504
rect 300 7476 308 7484
rect 1692 7476 1700 7484
rect 2476 7476 2484 7484
rect 4124 7476 4132 7484
rect 4268 7476 4276 7484
rect 4396 7476 4404 7484
rect 7004 7476 7012 7484
rect 7100 7476 7108 7484
rect 7452 7476 7460 7484
rect 8460 7476 8468 7484
rect 8748 7476 8756 7484
rect 8844 7476 8852 7484
rect 9836 7476 9844 7484
rect 9948 7476 9956 7484
rect 76 7456 84 7464
rect 92 7456 100 7464
rect 908 7456 916 7464
rect 2028 7456 2036 7464
rect 4540 7456 4548 7464
rect 6012 7456 6020 7464
rect 6188 7456 6196 7464
rect 9180 7456 9188 7464
rect 9276 7456 9284 7464
rect 9308 7456 9316 7464
rect 9708 7456 9716 7464
rect 3500 7436 3508 7444
rect 9596 7436 9604 7444
rect 316 7416 324 7424
rect 908 7416 916 7424
rect 6572 7416 6580 7424
rect 7468 7416 7476 7424
rect 9036 7416 9044 7424
rect 572 7396 580 7404
rect 3180 7396 3188 7404
rect 7884 7396 7892 7404
rect 8316 7396 8324 7404
rect 76 7376 84 7384
rect 92 7376 100 7384
rect 3740 7376 3748 7384
rect 6236 7376 6244 7384
rect 7244 7376 7252 7384
rect 7548 7376 7556 7384
rect 8140 7376 8148 7384
rect 9260 7376 9268 7384
rect 4092 7356 4100 7364
rect 5212 7356 5220 7364
rect 5340 7356 5348 7364
rect 8284 7356 8292 7364
rect 316 7336 324 7344
rect 636 7336 644 7344
rect 764 7336 772 7344
rect 1868 7336 1876 7344
rect 2764 7336 2772 7344
rect 3084 7336 3092 7344
rect 3228 7336 3236 7344
rect 3372 7336 3380 7344
rect 4652 7336 4660 7344
rect 4844 7336 4852 7344
rect 5180 7336 5188 7344
rect 5564 7336 5572 7344
rect 7452 7336 7460 7344
rect 7708 7336 7716 7344
rect 7772 7336 7780 7344
rect 7884 7336 7892 7344
rect 9708 7336 9716 7344
rect 2444 7316 2452 7324
rect 3340 7316 3348 7324
rect 3612 7316 3620 7324
rect 4092 7316 4100 7324
rect 4444 7316 4452 7324
rect 5868 7316 5876 7324
rect 7484 7316 7492 7324
rect 8172 7316 8180 7324
rect 8556 7316 8564 7324
rect 9052 7316 9060 7324
rect 9612 7316 9620 7324
rect 10268 7316 10276 7324
rect 1308 7296 1316 7304
rect 1564 7296 1572 7304
rect 2492 7296 2500 7304
rect 4460 7296 4468 7304
rect 4844 7296 4852 7304
rect 5180 7296 5188 7304
rect 5580 7296 5588 7304
rect 5772 7296 5780 7304
rect 5884 7296 5892 7304
rect 6172 7296 6180 7304
rect 6348 7296 6356 7304
rect 6380 7296 6388 7304
rect 8044 7296 8052 7304
rect 8476 7296 8484 7304
rect 9644 7296 9652 7304
rect 9916 7296 9924 7304
rect 1244 7276 1252 7284
rect 1548 7276 1556 7284
rect 2716 7276 2724 7284
rect 2748 7276 2756 7284
rect 3980 7276 3988 7284
rect 4220 7276 4228 7284
rect 4972 7276 4980 7284
rect 5900 7276 5908 7284
rect 6604 7276 6612 7284
rect 6956 7276 6964 7284
rect 7964 7276 7972 7284
rect 428 7256 436 7264
rect 892 7256 900 7264
rect 3116 7256 3124 7264
rect 3324 7256 3332 7264
rect 3532 7256 3540 7264
rect 4396 7256 4404 7264
rect 4604 7256 4612 7264
rect 4988 7256 4996 7264
rect 7372 7256 7380 7264
rect 8268 7256 8276 7264
rect 8828 7256 8836 7264
rect 9692 7256 9700 7264
rect 2236 7216 2244 7224
rect 7180 7216 7188 7224
rect 9420 7216 9428 7224
rect 9436 7216 9444 7224
rect 1660 7196 1668 7204
rect 2460 7176 2468 7184
rect 8268 7176 8276 7184
rect 5228 7156 5236 7164
rect 8172 7156 8180 7164
rect 8268 7156 8276 7164
rect 780 7136 788 7144
rect 2732 7136 2740 7144
rect 5212 7136 5220 7144
rect 7180 7136 7188 7144
rect 8012 7136 8020 7144
rect 9868 7136 9876 7144
rect 284 7116 292 7124
rect 1628 7116 1636 7124
rect 2620 7116 2628 7124
rect 2796 7116 2804 7124
rect 2908 7116 2916 7124
rect 3708 7116 3716 7124
rect 3756 7116 3764 7124
rect 4540 7116 4548 7124
rect 4988 7116 4996 7124
rect 5212 7116 5220 7124
rect 5772 7116 5780 7124
rect 6172 7116 6180 7124
rect 6924 7116 6932 7124
rect 7452 7116 7460 7124
rect 8828 7116 8836 7124
rect 8876 7116 8884 7124
rect 8972 7116 8980 7124
rect 8988 7116 8996 7124
rect 9628 7116 9636 7124
rect 9852 7116 9860 7124
rect 684 7096 692 7104
rect 1068 7096 1076 7104
rect 1100 7096 1108 7104
rect 1132 7096 1140 7104
rect 1532 7096 1540 7104
rect 1564 7096 1572 7104
rect 3372 7096 3380 7104
rect 3868 7096 3876 7104
rect 4812 7096 4820 7104
rect 7116 7096 7124 7104
rect 8028 7096 8036 7104
rect 8396 7096 8404 7104
rect 9852 7096 9860 7104
rect 636 7076 644 7084
rect 2108 7076 2116 7084
rect 2252 7076 2260 7084
rect 2348 7076 2356 7084
rect 2460 7076 2468 7084
rect 3020 7076 3028 7084
rect 3084 7076 3092 7084
rect 3340 7076 3348 7084
rect 4476 7076 4484 7084
rect 5228 7076 5236 7084
rect 5468 7076 5476 7084
rect 6012 7076 6020 7084
rect 7100 7076 7108 7084
rect 7340 7076 7348 7084
rect 7548 7076 7556 7084
rect 8876 7076 8884 7084
rect 204 7056 212 7064
rect 1308 7056 1316 7064
rect 2444 7056 2452 7064
rect 3532 7056 3540 7064
rect 3692 7056 3700 7064
rect 4092 7056 4100 7064
rect 5388 7056 5396 7064
rect 5788 7056 5796 7064
rect 5884 7056 5892 7064
rect 6780 7056 6788 7064
rect 9420 7056 9428 7064
rect 780 7036 788 7044
rect 1788 7036 1796 7044
rect 2108 7036 2116 7044
rect 3116 7036 3124 7044
rect 4732 7036 4740 7044
rect 5900 7036 5908 7044
rect 7500 7036 7508 7044
rect 9676 7036 9684 7044
rect 1884 7016 1892 7024
rect 2588 7016 2596 7024
rect 6796 7016 6804 7024
rect 7372 7016 7380 7024
rect 9468 7016 9476 7024
rect 2252 6996 2260 7004
rect 3020 6996 3028 7004
rect 6924 6996 6932 7004
rect 684 6976 692 6984
rect 2924 6976 2932 6984
rect 8556 6976 8564 6984
rect 9068 6976 9076 6984
rect 2092 6956 2100 6964
rect 4556 6956 4564 6964
rect 6604 6956 6612 6964
rect 7196 6956 7204 6964
rect 7692 6956 7700 6964
rect 9436 6956 9444 6964
rect 876 6936 884 6944
rect 1852 6936 1860 6944
rect 2636 6936 2644 6944
rect 2972 6936 2980 6944
rect 4332 6936 4340 6944
rect 4828 6936 4836 6944
rect 5084 6936 5092 6944
rect 5404 6936 5412 6944
rect 5900 6936 5908 6944
rect 6268 6936 6276 6944
rect 6540 6936 6548 6944
rect 7004 6936 7012 6944
rect 7228 6936 7236 6944
rect 7644 6936 7652 6944
rect 8012 6936 8020 6944
rect 8588 6936 8596 6944
rect 2284 6916 2292 6924
rect 2348 6916 2356 6924
rect 2956 6916 2964 6924
rect 3500 6916 3508 6924
rect 4604 6916 4612 6924
rect 4972 6916 4980 6924
rect 5052 6916 5060 6924
rect 7212 6916 7220 6924
rect 8396 6916 8404 6924
rect 8828 6936 8836 6944
rect 8908 6936 8916 6944
rect 9532 6936 9540 6944
rect 9660 6936 9668 6944
rect 9372 6916 9380 6924
rect 428 6896 436 6904
rect 508 6896 516 6904
rect 972 6896 980 6904
rect 1180 6896 1188 6904
rect 2076 6896 2084 6904
rect 2428 6896 2436 6904
rect 3308 6896 3316 6904
rect 3484 6896 3492 6904
rect 3996 6896 4004 6904
rect 4844 6896 4852 6904
rect 4876 6896 4884 6904
rect 6012 6896 6020 6904
rect 6204 6896 6212 6904
rect 6316 6896 6324 6904
rect 6956 6896 6964 6904
rect 7788 6896 7796 6904
rect 7820 6896 7828 6904
rect 9692 6896 9700 6904
rect 9724 6896 9732 6904
rect 4220 6876 4228 6884
rect 6684 6876 6692 6884
rect 9116 6876 9124 6884
rect 9324 6876 9332 6884
rect 9452 6876 9460 6884
rect 9500 6876 9508 6884
rect 1548 6856 1556 6864
rect 3548 6856 3556 6864
rect 3788 6856 3796 6864
rect 8684 6856 8692 6864
rect 1340 6836 1348 6844
rect 4204 6836 4212 6844
rect 4268 6836 4276 6844
rect 4700 6836 4708 6844
rect 4940 6836 4948 6844
rect 6988 6836 6996 6844
rect 76 6816 84 6824
rect 5596 6816 5604 6824
rect 972 6796 980 6804
rect 2636 6776 2644 6784
rect 316 6756 324 6764
rect 1884 6756 1892 6764
rect 2924 6756 2932 6764
rect 4268 6756 4276 6764
rect 5052 6756 5060 6764
rect 5756 6756 5764 6764
rect 2364 6736 2372 6744
rect 2668 6736 2676 6744
rect 3980 6736 3988 6744
rect 4412 6736 4420 6744
rect 5084 6736 5092 6744
rect 6732 6736 6740 6744
rect 6972 6736 6980 6744
rect 9532 6736 9540 6744
rect 76 6716 84 6724
rect 508 6716 516 6724
rect 1356 6716 1364 6724
rect 3180 6716 3188 6724
rect 3484 6716 3492 6724
rect 3596 6716 3604 6724
rect 3836 6716 3844 6724
rect 4748 6716 4756 6724
rect 5084 6716 5092 6724
rect 5468 6716 5476 6724
rect 7100 6716 7108 6724
rect 7228 6716 7236 6724
rect 7292 6716 7300 6724
rect 7484 6716 7492 6724
rect 7500 6716 7508 6724
rect 7740 6716 7748 6724
rect 8572 6716 8580 6724
rect 9068 6716 9076 6724
rect 9372 6716 9380 6724
rect 9564 6716 9572 6724
rect 972 6696 980 6704
rect 1148 6696 1156 6704
rect 1660 6696 1668 6704
rect 2268 6696 2276 6704
rect 5596 6696 5604 6704
rect 5852 6696 5860 6704
rect 6188 6696 6196 6704
rect 6492 6696 6500 6704
rect 9900 6696 9908 6704
rect 684 6676 692 6684
rect 748 6676 756 6684
rect 1132 6676 1140 6684
rect 1244 6676 1252 6684
rect 2284 6676 2292 6684
rect 2796 6676 2804 6684
rect 2828 6676 2836 6684
rect 4044 6676 4052 6684
rect 4252 6676 4260 6684
rect 4492 6676 4500 6684
rect 5084 6676 5092 6684
rect 5228 6676 5236 6684
rect 5564 6676 5572 6684
rect 6060 6676 6068 6684
rect 7820 6676 7828 6684
rect 8460 6676 8468 6684
rect 8556 6676 8564 6684
rect 8876 6676 8884 6684
rect 9020 6676 9028 6684
rect 9660 6676 9668 6684
rect 108 6656 116 6664
rect 684 6656 692 6664
rect 2700 6656 2708 6664
rect 2972 6656 2980 6664
rect 5836 6656 5844 6664
rect 6028 6656 6036 6664
rect 6156 6656 6164 6664
rect 6268 6656 6276 6664
rect 7116 6656 7124 6664
rect 7276 6656 7284 6664
rect 7660 6656 7668 6664
rect 7692 6656 7700 6664
rect 7868 6656 7876 6664
rect 9052 6656 9060 6664
rect 1548 6636 1556 6644
rect 1644 6636 1652 6644
rect 1852 6636 1860 6644
rect 2828 6636 2836 6644
rect 3484 6636 3492 6644
rect 4012 6636 4020 6644
rect 4348 6636 4356 6644
rect 5212 6636 5220 6644
rect 5788 6636 5796 6644
rect 6860 6636 6868 6644
rect 6972 6636 6980 6644
rect 8780 6636 8788 6644
rect 108 6616 116 6624
rect 2668 6616 2676 6624
rect 5180 6616 5188 6624
rect 7788 6616 7796 6624
rect 300 6596 308 6604
rect 748 6596 756 6604
rect 2108 6596 2116 6604
rect 3100 6596 3108 6604
rect 4252 6596 4260 6604
rect 4876 6596 4884 6604
rect 5772 6596 5780 6604
rect 6300 6596 6308 6604
rect 6492 6596 6500 6604
rect 6764 6596 6772 6604
rect 8796 6596 8804 6604
rect 220 6576 228 6584
rect 1084 6576 1092 6584
rect 1948 6576 1956 6584
rect 2220 6576 2228 6584
rect 2268 6576 2276 6584
rect 3548 6576 3556 6584
rect 3628 6576 3636 6584
rect 3788 6576 3796 6584
rect 7740 6576 7748 6584
rect 8764 6576 8772 6584
rect 300 6556 308 6564
rect 2412 6556 2420 6564
rect 2508 6556 2516 6564
rect 2636 6556 2644 6564
rect 4716 6556 4724 6564
rect 5708 6556 5716 6564
rect 6156 6556 6164 6564
rect 6364 6556 6372 6564
rect 6956 6556 6964 6564
rect 7948 6556 7956 6564
rect 7964 6556 7972 6564
rect 1660 6536 1668 6544
rect 1788 6536 1796 6544
rect 2396 6536 2404 6544
rect 2748 6536 2756 6544
rect 2812 6536 2820 6544
rect 3100 6536 3108 6544
rect 3260 6536 3268 6544
rect 3404 6536 3412 6544
rect 3964 6536 3972 6544
rect 4332 6536 4340 6544
rect 4828 6536 4836 6544
rect 5292 6536 5300 6544
rect 5420 6536 5428 6544
rect 6172 6536 6180 6544
rect 7148 6536 7156 6544
rect 7548 6536 7556 6544
rect 7788 6536 7796 6544
rect 7852 6536 7860 6544
rect 8092 6536 8100 6544
rect 8236 6536 8244 6544
rect 8268 6536 8276 6544
rect 9212 6536 9220 6544
rect 9676 6536 9684 6544
rect 10012 6536 10020 6544
rect 844 6516 852 6524
rect 1324 6516 1332 6524
rect 1996 6516 2004 6524
rect 4924 6516 4932 6524
rect 5868 6516 5876 6524
rect 6588 6516 6596 6524
rect 7372 6516 7380 6524
rect 7900 6516 7908 6524
rect 668 6496 676 6504
rect 1900 6496 1908 6504
rect 2108 6496 2116 6504
rect 2636 6496 2644 6504
rect 2652 6496 2660 6504
rect 4332 6496 4340 6504
rect 4444 6496 4452 6504
rect 4524 6496 4532 6504
rect 4556 6496 4564 6504
rect 5756 6496 5764 6504
rect 6012 6496 6020 6504
rect 6348 6496 6356 6504
rect 6604 6496 6612 6504
rect 7372 6496 7380 6504
rect 7852 6496 7860 6504
rect 7868 6496 7876 6504
rect 8348 6496 8356 6504
rect 8460 6496 8468 6504
rect 8540 6496 8548 6504
rect 8796 6496 8804 6504
rect 9660 6496 9668 6504
rect 9900 6496 9908 6504
rect 412 6476 420 6484
rect 2844 6476 2852 6484
rect 3244 6476 3252 6484
rect 3804 6476 3812 6484
rect 7612 6476 7620 6484
rect 8140 6476 8148 6484
rect 876 6456 884 6464
rect 2636 6456 2644 6464
rect 3980 6456 3988 6464
rect 7484 6456 7492 6464
rect 6764 6436 6772 6444
rect 2236 6416 2244 6424
rect 3148 6396 3156 6404
rect 8812 6376 8820 6384
rect 3116 6356 3124 6364
rect 6348 6356 6356 6364
rect 1100 6336 1108 6344
rect 1420 6336 1428 6344
rect 3180 6336 3188 6344
rect 3628 6336 3636 6344
rect 4060 6336 4068 6344
rect 4620 6336 4628 6344
rect 5020 6336 5028 6344
rect 5516 6336 5524 6344
rect 5596 6336 5604 6344
rect 6252 6336 6260 6344
rect 6364 6336 6372 6344
rect 108 6316 116 6324
rect 684 6316 692 6324
rect 2908 6316 2916 6324
rect 3244 6316 3252 6324
rect 3532 6316 3540 6324
rect 5020 6316 5028 6324
rect 5292 6316 5300 6324
rect 5836 6316 5844 6324
rect 5884 6316 5892 6324
rect 6124 6316 6132 6324
rect 8476 6316 8484 6324
rect 9660 6316 9668 6324
rect 300 6296 308 6304
rect 2236 6296 2244 6304
rect 2492 6296 2500 6304
rect 2796 6296 2804 6304
rect 4348 6296 4356 6304
rect 4940 6296 4948 6304
rect 5020 6296 5028 6304
rect 5900 6296 5908 6304
rect 6588 6296 6596 6304
rect 7276 6296 7284 6304
rect 7980 6296 7988 6304
rect 9404 6296 9412 6304
rect 9708 6296 9716 6304
rect 428 6276 436 6284
rect 2556 6276 2564 6284
rect 4652 6276 4660 6284
rect 5596 6276 5604 6284
rect 5868 6276 5876 6284
rect 6476 6276 6484 6284
rect 7004 6276 7012 6284
rect 7036 6276 7044 6284
rect 7084 6276 7092 6284
rect 8012 6276 8020 6284
rect 8428 6276 8436 6284
rect 8684 6276 8692 6284
rect 8908 6276 8916 6284
rect 9372 6276 9380 6284
rect 9836 6276 9844 6284
rect 92 6256 100 6264
rect 236 6236 244 6244
rect 1452 6256 1460 6264
rect 1612 6256 1620 6264
rect 2476 6256 2484 6264
rect 2684 6256 2692 6264
rect 3116 6256 3124 6264
rect 3820 6256 3828 6264
rect 4012 6256 4020 6264
rect 4236 6256 4244 6264
rect 4956 6256 4964 6264
rect 5372 6256 5380 6264
rect 5388 6256 5396 6264
rect 6108 6256 6116 6264
rect 6236 6256 6244 6264
rect 6604 6256 6612 6264
rect 7372 6256 7380 6264
rect 1596 6236 1604 6244
rect 1900 6236 1908 6244
rect 2860 6236 2868 6244
rect 4012 6236 4020 6244
rect 7340 6236 7348 6244
rect 8812 6236 8820 6244
rect 9836 6256 9844 6264
rect 108 6216 116 6224
rect 2332 6216 2340 6224
rect 4060 6216 4068 6224
rect 92 6196 100 6204
rect 1468 6196 1476 6204
rect 2684 6196 2692 6204
rect 2908 6196 2916 6204
rect 5372 6196 5380 6204
rect 9676 6196 9684 6204
rect 844 6176 852 6184
rect 1132 6176 1140 6184
rect 476 6156 484 6164
rect 2636 6176 2644 6184
rect 4012 6176 4020 6184
rect 4220 6176 4228 6184
rect 4812 6176 4820 6184
rect 5276 6176 5284 6184
rect 7180 6176 7188 6184
rect 7356 6176 7364 6184
rect 7628 6176 7636 6184
rect 2156 6156 2164 6164
rect 636 6136 644 6144
rect 876 6136 884 6144
rect 1628 6136 1636 6144
rect 1756 6136 1764 6144
rect 2460 6136 2468 6144
rect 2492 6136 2500 6144
rect 3564 6136 3572 6144
rect 5100 6156 5108 6164
rect 6364 6156 6372 6164
rect 6860 6156 6868 6164
rect 7116 6156 7124 6164
rect 9516 6156 9524 6164
rect 3948 6136 3956 6144
rect 3964 6136 3972 6144
rect 3980 6136 3988 6144
rect 4620 6136 4628 6144
rect 4780 6136 4788 6144
rect 6060 6136 6068 6144
rect 6380 6136 6388 6144
rect 6796 6136 6804 6144
rect 7132 6136 7140 6144
rect 7340 6136 7348 6144
rect 7852 6136 7860 6144
rect 8332 6136 8340 6144
rect 8652 6136 8660 6144
rect 9004 6136 9012 6144
rect 9228 6136 9236 6144
rect 9756 6136 9764 6144
rect 1084 6116 1092 6124
rect 1132 6116 1140 6124
rect 2524 6116 2532 6124
rect 3980 6116 3988 6124
rect 5740 6116 5748 6124
rect 6604 6116 6612 6124
rect 7180 6116 7188 6124
rect 7692 6116 7700 6124
rect 9164 6116 9172 6124
rect 9916 6116 9924 6124
rect 652 6096 660 6104
rect 1180 6096 1188 6104
rect 1612 6096 1620 6104
rect 1644 6096 1652 6104
rect 1996 6096 2004 6104
rect 2076 6096 2084 6104
rect 2332 6096 2340 6104
rect 2460 6096 2468 6104
rect 2972 6096 2980 6104
rect 3324 6096 3332 6104
rect 4556 6096 4564 6104
rect 4764 6096 4772 6104
rect 7020 6096 7028 6104
rect 8012 6096 8020 6104
rect 8668 6096 8676 6104
rect 9372 6096 9380 6104
rect 9868 6096 9876 6104
rect 892 6076 900 6084
rect 972 6076 980 6084
rect 2492 6076 2500 6084
rect 3100 6076 3108 6084
rect 3740 6076 3748 6084
rect 4924 6076 4932 6084
rect 6604 6076 6612 6084
rect 6684 6076 6692 6084
rect 7228 6076 7236 6084
rect 9868 6076 9876 6084
rect 1532 6056 1540 6064
rect 2300 6056 2308 6064
rect 5228 6056 5236 6064
rect 6348 6056 6356 6064
rect 6780 6056 6788 6064
rect 8124 6056 8132 6064
rect 9804 6056 9812 6064
rect 9868 6056 9876 6064
rect 556 6036 564 6044
rect 2204 6036 2212 6044
rect 4108 6036 4116 6044
rect 6796 6036 6804 6044
rect 2012 6016 2020 6024
rect 3580 6016 3588 6024
rect 6524 6016 6532 6024
rect 9004 5996 9012 6004
rect 5260 5976 5268 5984
rect 556 5956 564 5964
rect 2908 5956 2916 5964
rect 6044 5956 6052 5964
rect 8332 5956 8340 5964
rect 636 5936 644 5944
rect 1580 5936 1588 5944
rect 2428 5936 2436 5944
rect 2508 5936 2516 5944
rect 2524 5936 2532 5944
rect 3596 5936 3604 5944
rect 4652 5936 4660 5944
rect 5420 5936 5428 5944
rect 6124 5936 6132 5944
rect 6460 5936 6468 5944
rect 7820 5936 7828 5944
rect 764 5916 772 5924
rect 1644 5916 1652 5924
rect 1948 5916 1956 5924
rect 2716 5916 2724 5924
rect 4044 5916 4052 5924
rect 4252 5916 4260 5924
rect 4812 5916 4820 5924
rect 5228 5916 5236 5924
rect 5516 5916 5524 5924
rect 5948 5916 5956 5924
rect 6108 5916 6116 5924
rect 6300 5916 6308 5924
rect 6492 5916 6500 5924
rect 7292 5916 7300 5924
rect 8540 5916 8548 5924
rect 8572 5916 8580 5924
rect 8716 5916 8724 5924
rect 8732 5916 8740 5924
rect 9036 5916 9044 5924
rect 9580 5916 9588 5924
rect 1804 5896 1812 5904
rect 2012 5896 2020 5904
rect 2268 5896 2276 5904
rect 3580 5896 3588 5904
rect 3804 5896 3812 5904
rect 4028 5896 4036 5904
rect 5004 5896 5012 5904
rect 5788 5896 5796 5904
rect 6076 5896 6084 5904
rect 7948 5896 7956 5904
rect 7980 5896 7988 5904
rect 8044 5896 8052 5904
rect 236 5876 244 5884
rect 860 5876 868 5884
rect 3020 5876 3028 5884
rect 3324 5876 3332 5884
rect 3596 5876 3604 5884
rect 3788 5876 3796 5884
rect 4236 5876 4244 5884
rect 5356 5876 5364 5884
rect 5404 5876 5412 5884
rect 6428 5876 6436 5884
rect 6540 5876 6548 5884
rect 6748 5876 6756 5884
rect 6812 5876 6820 5884
rect 7148 5876 7156 5884
rect 8268 5876 8276 5884
rect 8284 5876 8292 5884
rect 8940 5876 8948 5884
rect 9580 5876 9588 5884
rect 3964 5856 3972 5864
rect 4684 5856 4692 5864
rect 5388 5856 5396 5864
rect 5484 5856 5492 5864
rect 5580 5856 5588 5864
rect 6156 5856 6164 5864
rect 6460 5856 6468 5864
rect 7660 5856 7668 5864
rect 7788 5856 7796 5864
rect 7884 5856 7892 5864
rect 8524 5856 8532 5864
rect 8604 5856 8612 5864
rect 7868 5836 7876 5844
rect 2332 5816 2340 5824
rect 2348 5816 2356 5824
rect 5932 5816 5940 5824
rect 7724 5816 7732 5824
rect 8012 5816 8020 5824
rect 10044 5816 10052 5824
rect 2268 5796 2276 5804
rect 3164 5796 3172 5804
rect 3436 5796 3444 5804
rect 3596 5796 3604 5804
rect 4684 5796 4692 5804
rect 8124 5796 8132 5804
rect 8476 5796 8484 5804
rect 1100 5776 1108 5784
rect 1676 5776 1684 5784
rect 2780 5776 2788 5784
rect 3836 5776 3844 5784
rect 6924 5776 6932 5784
rect 7196 5776 7204 5784
rect 8348 5776 8356 5784
rect 9804 5776 9812 5784
rect 316 5756 324 5764
rect 412 5756 420 5764
rect 1628 5756 1636 5764
rect 2364 5756 2372 5764
rect 2476 5756 2484 5764
rect 3052 5756 3060 5764
rect 3180 5756 3188 5764
rect 4508 5756 4516 5764
rect 5676 5756 5684 5764
rect 6348 5756 6356 5764
rect 6764 5756 6772 5764
rect 76 5736 84 5744
rect 1116 5736 1124 5744
rect 1356 5736 1364 5744
rect 3916 5736 3924 5744
rect 4220 5736 4228 5744
rect 4812 5736 4820 5744
rect 5228 5736 5236 5744
rect 5484 5736 5492 5744
rect 5516 5736 5524 5744
rect 5580 5736 5588 5744
rect 6364 5736 6372 5744
rect 6844 5736 6852 5744
rect 6924 5736 6932 5744
rect 8140 5736 8148 5744
rect 9116 5736 9124 5744
rect 9436 5736 9444 5744
rect 9692 5736 9700 5744
rect 652 5716 660 5724
rect 732 5716 740 5724
rect 1212 5716 1220 5724
rect 3036 5716 3044 5724
rect 3052 5716 3060 5724
rect 3196 5716 3204 5724
rect 3884 5716 3892 5724
rect 4044 5716 4052 5724
rect 4076 5716 4084 5724
rect 4924 5716 4932 5724
rect 5340 5716 5348 5724
rect 5452 5716 5460 5724
rect 6364 5716 6372 5724
rect 7148 5716 7156 5724
rect 7500 5716 7508 5724
rect 9852 5716 9860 5724
rect 9900 5716 9908 5724
rect 204 5696 212 5704
rect 1084 5696 1092 5704
rect 1356 5696 1364 5704
rect 2108 5696 2116 5704
rect 2332 5696 2340 5704
rect 3564 5696 3572 5704
rect 3580 5696 3588 5704
rect 4556 5696 4564 5704
rect 4620 5696 4628 5704
rect 5356 5696 5364 5704
rect 6124 5696 6132 5704
rect 6508 5696 6516 5704
rect 6812 5696 6820 5704
rect 6956 5696 6964 5704
rect 7292 5696 7300 5704
rect 7500 5696 7508 5704
rect 8092 5696 8100 5704
rect 8508 5696 8516 5704
rect 8668 5696 8676 5704
rect 9388 5696 9396 5704
rect 9468 5696 9476 5704
rect 9500 5696 9508 5704
rect 9708 5696 9716 5704
rect 9884 5696 9892 5704
rect 428 5676 436 5684
rect 508 5676 516 5684
rect 4476 5676 4484 5684
rect 4668 5676 4676 5684
rect 4796 5676 4804 5684
rect 652 5656 660 5664
rect 1468 5656 1476 5664
rect 1676 5656 1684 5664
rect 7404 5676 7412 5684
rect 8812 5676 8820 5684
rect 5708 5656 5716 5664
rect 7724 5656 7732 5664
rect 9004 5656 9012 5664
rect 2508 5636 2516 5644
rect 2668 5636 2676 5644
rect 2748 5636 2756 5644
rect 924 5616 932 5624
rect 2572 5616 2580 5624
rect 4924 5616 4932 5624
rect 8956 5616 8964 5624
rect 9420 5616 9428 5624
rect 3788 5596 3796 5604
rect 4204 5576 4212 5584
rect 1212 5556 1220 5564
rect 2828 5556 2836 5564
rect 3420 5556 3428 5564
rect 3916 5556 3924 5564
rect 4492 5556 4500 5564
rect 4828 5556 4836 5564
rect 7404 5556 7412 5564
rect 2748 5536 2756 5544
rect 3180 5536 3188 5544
rect 3308 5536 3316 5544
rect 4716 5536 4724 5544
rect 5420 5536 5428 5544
rect 6044 5536 6052 5544
rect 6588 5536 6596 5544
rect 6956 5536 6964 5544
rect 7020 5536 7028 5544
rect 7100 5536 7108 5544
rect 8716 5536 8724 5544
rect 732 5516 740 5524
rect 1596 5516 1604 5524
rect 2060 5516 2068 5524
rect 2156 5516 2164 5524
rect 2716 5516 2724 5524
rect 4332 5516 4340 5524
rect 4364 5516 4372 5524
rect 4588 5516 4596 5524
rect 5180 5516 5188 5524
rect 6524 5516 6532 5524
rect 6828 5516 6836 5524
rect 6844 5516 6852 5524
rect 7452 5516 7460 5524
rect 7932 5516 7940 5524
rect 8236 5516 8244 5524
rect 8268 5516 8276 5524
rect 8300 5516 8308 5524
rect 8428 5516 8436 5524
rect 9740 5516 9748 5524
rect 9836 5516 9844 5524
rect 652 5496 660 5504
rect 924 5496 932 5504
rect 1468 5496 1476 5504
rect 2044 5496 2052 5504
rect 2508 5496 2516 5504
rect 2524 5496 2532 5504
rect 3244 5496 3252 5504
rect 3932 5496 3940 5504
rect 4284 5496 4292 5504
rect 4604 5496 4612 5504
rect 4668 5496 4676 5504
rect 4716 5496 4724 5504
rect 5228 5496 5236 5504
rect 5932 5496 5940 5504
rect 6428 5496 6436 5504
rect 7548 5496 7556 5504
rect 7708 5496 7716 5504
rect 7948 5496 7956 5504
rect 7980 5496 7988 5504
rect 8508 5496 8516 5504
rect 8972 5496 8980 5504
rect 9068 5496 9076 5504
rect 732 5476 740 5484
rect 908 5476 916 5484
rect 1356 5476 1364 5484
rect 3580 5476 3588 5484
rect 3820 5476 3828 5484
rect 5452 5476 5460 5484
rect 5740 5476 5748 5484
rect 5836 5476 5844 5484
rect 6156 5476 6164 5484
rect 6604 5476 6612 5484
rect 6716 5476 6724 5484
rect 6732 5476 6740 5484
rect 6812 5476 6820 5484
rect 6956 5476 6964 5484
rect 7260 5476 7268 5484
rect 7292 5476 7300 5484
rect 7388 5476 7396 5484
rect 7660 5476 7668 5484
rect 8588 5476 8596 5484
rect 9404 5476 9412 5484
rect 9436 5476 9444 5484
rect 2444 5456 2452 5464
rect 3868 5456 3876 5464
rect 5356 5456 5364 5464
rect 7724 5456 7732 5464
rect 8172 5456 8180 5464
rect 8572 5456 8580 5464
rect 8620 5456 8628 5464
rect 8652 5456 8660 5464
rect 8988 5456 8996 5464
rect 9036 5456 9044 5464
rect 524 5436 532 5444
rect 1148 5436 1156 5444
rect 2220 5436 2228 5444
rect 2700 5436 2708 5444
rect 2716 5436 2724 5444
rect 3964 5436 3972 5444
rect 3996 5436 4004 5444
rect 5580 5436 5588 5444
rect 8956 5436 8964 5444
rect 1788 5416 1796 5424
rect 2700 5416 2708 5424
rect 3404 5416 3412 5424
rect 3628 5416 3636 5424
rect 6364 5416 6372 5424
rect 7196 5416 7204 5424
rect 7852 5416 7860 5424
rect 908 5396 916 5404
rect 2108 5396 2116 5404
rect 3692 5396 3700 5404
rect 5116 5396 5124 5404
rect 2220 5376 2228 5384
rect 2524 5376 2532 5384
rect 3404 5376 3412 5384
rect 4044 5376 4052 5384
rect 4924 5376 4932 5384
rect 5884 5376 5892 5384
rect 6572 5376 6580 5384
rect 7660 5396 7668 5404
rect 9820 5396 9828 5404
rect 7180 5376 7188 5384
rect 8172 5376 8180 5384
rect 8556 5376 8564 5384
rect 9820 5376 9828 5384
rect 316 5356 324 5364
rect 1148 5356 1156 5364
rect 1340 5356 1348 5364
rect 2028 5356 2036 5364
rect 1244 5336 1252 5344
rect 2108 5336 2116 5344
rect 2748 5336 2756 5344
rect 2828 5336 2836 5344
rect 2860 5336 2868 5344
rect 4236 5356 4244 5364
rect 4556 5356 4564 5364
rect 6124 5356 6132 5364
rect 6188 5356 6196 5364
rect 6220 5356 6228 5364
rect 6972 5356 6980 5364
rect 7228 5356 7236 5364
rect 7420 5356 7428 5364
rect 8924 5356 8932 5364
rect 8972 5356 8980 5364
rect 9436 5356 9444 5364
rect 9916 5356 9924 5364
rect 3644 5336 3652 5344
rect 4124 5336 4132 5344
rect 4204 5336 4212 5344
rect 4236 5336 4244 5344
rect 4924 5336 4932 5344
rect 4940 5336 4948 5344
rect 5228 5336 5236 5344
rect 5580 5336 5588 5344
rect 6380 5336 6388 5344
rect 6716 5336 6724 5344
rect 7052 5336 7060 5344
rect 7500 5336 7508 5344
rect 8428 5336 8436 5344
rect 8460 5336 8468 5344
rect 8636 5336 8644 5344
rect 9036 5336 9044 5344
rect 9084 5336 9092 5344
rect 9596 5336 9604 5344
rect 10012 5336 10020 5344
rect 652 5316 660 5324
rect 3420 5316 3428 5324
rect 3628 5316 3636 5324
rect 6364 5316 6372 5324
rect 6476 5316 6484 5324
rect 6700 5316 6708 5324
rect 7852 5316 7860 5324
rect 9548 5316 9556 5324
rect 10268 5316 10276 5324
rect 1404 5296 1412 5304
rect 1580 5296 1588 5304
rect 3420 5296 3428 5304
rect 4044 5296 4052 5304
rect 4796 5296 4804 5304
rect 5020 5296 5028 5304
rect 5244 5296 5252 5304
rect 5724 5296 5732 5304
rect 6140 5296 6148 5304
rect 6300 5296 6308 5304
rect 6508 5296 6516 5304
rect 6988 5296 6996 5304
rect 7388 5296 7396 5304
rect 7676 5296 7684 5304
rect 8668 5296 8676 5304
rect 8956 5296 8964 5304
rect 9340 5296 9348 5304
rect 9772 5296 9780 5304
rect 9884 5296 9892 5304
rect 10076 5296 10084 5304
rect 1756 5276 1764 5284
rect 2284 5276 2292 5284
rect 2540 5276 2548 5284
rect 3212 5276 3220 5284
rect 4812 5276 4820 5284
rect 6684 5276 6692 5284
rect 7404 5276 7412 5284
rect 8476 5276 8484 5284
rect 8524 5276 8532 5284
rect 9372 5276 9380 5284
rect 9708 5276 9716 5284
rect 1100 5256 1108 5264
rect 2812 5256 2820 5264
rect 4220 5256 4228 5264
rect 5260 5256 5268 5264
rect 5340 5256 5348 5264
rect 7964 5256 7972 5264
rect 8556 5256 8564 5264
rect 892 5236 900 5244
rect 2476 5236 2484 5244
rect 3260 5236 3268 5244
rect 3884 5236 3892 5244
rect 6668 5236 6676 5244
rect 92 5216 100 5224
rect 460 5216 468 5224
rect 1228 5216 1236 5224
rect 6124 5216 6132 5224
rect 6508 5216 6516 5224
rect 9612 5216 9620 5224
rect 3420 5196 3428 5204
rect 3644 5196 3652 5204
rect 4124 5196 4132 5204
rect 7612 5196 7620 5204
rect 3532 5176 3540 5184
rect 7196 5176 7204 5184
rect 8460 5176 8468 5184
rect 908 5156 916 5164
rect 2796 5156 2804 5164
rect 6028 5156 6036 5164
rect 7468 5156 7476 5164
rect 7964 5156 7972 5164
rect 9052 5156 9060 5164
rect 524 5136 532 5144
rect 1580 5136 1588 5144
rect 2220 5136 2228 5144
rect 3804 5136 3812 5144
rect 5500 5136 5508 5144
rect 6492 5136 6500 5144
rect 6668 5136 6676 5144
rect 7260 5136 7268 5144
rect 972 5116 980 5124
rect 1228 5116 1236 5124
rect 1580 5116 1588 5124
rect 2940 5116 2948 5124
rect 3388 5116 3396 5124
rect 4252 5116 4260 5124
rect 5868 5116 5876 5124
rect 6652 5116 6660 5124
rect 7292 5116 7300 5124
rect 7340 5116 7348 5124
rect 7404 5116 7412 5124
rect 8188 5116 8196 5124
rect 8460 5116 8468 5124
rect 8812 5116 8820 5124
rect 9484 5116 9492 5124
rect 1084 5096 1092 5104
rect 2156 5096 2164 5104
rect 4108 5096 4116 5104
rect 4588 5096 4596 5104
rect 4812 5096 4820 5104
rect 5916 5096 5924 5104
rect 6108 5096 6116 5104
rect 8044 5096 8052 5104
rect 444 5076 452 5084
rect 1132 5076 1140 5084
rect 1212 5076 1220 5084
rect 2668 5076 2676 5084
rect 3612 5076 3620 5084
rect 5404 5076 5412 5084
rect 5484 5076 5492 5084
rect 6172 5076 6180 5084
rect 6668 5076 6676 5084
rect 9660 5076 9668 5084
rect 940 5056 948 5064
rect 1004 5056 1012 5064
rect 2572 5056 2580 5064
rect 3100 5056 3108 5064
rect 4396 5056 4404 5064
rect 5452 5056 5460 5064
rect 7004 5056 7012 5064
rect 7484 5056 7492 5064
rect 8428 5056 8436 5064
rect 8460 5056 8468 5064
rect 9628 5056 9636 5064
rect 1532 5036 1540 5044
rect 2588 5036 2596 5044
rect 6892 5036 6900 5044
rect 7612 5036 7620 5044
rect 3260 5016 3268 5024
rect 3852 5016 3860 5024
rect 4060 5016 4068 5024
rect 4396 4996 4404 5004
rect 6956 4996 6964 5004
rect 9932 4996 9940 5004
rect 2668 4976 2676 4984
rect 2940 4976 2948 4984
rect 3948 4976 3956 4984
rect 1580 4956 1588 4964
rect 2444 4956 2452 4964
rect 3260 4956 3268 4964
rect 4284 4956 4292 4964
rect 4540 4956 4548 4964
rect 5564 4956 5572 4964
rect 5740 4956 5748 4964
rect 6156 4956 6164 4964
rect 6172 4956 6180 4964
rect 7900 4956 7908 4964
rect 2940 4936 2948 4944
rect 3820 4936 3828 4944
rect 4588 4936 4596 4944
rect 4604 4936 4612 4944
rect 4956 4936 4964 4944
rect 6380 4936 6388 4944
rect 7036 4936 7044 4944
rect 7244 4936 7252 4944
rect 7308 4936 7316 4944
rect 668 4916 676 4924
rect 1196 4916 1204 4924
rect 1580 4916 1588 4924
rect 1836 4916 1844 4924
rect 2572 4916 2580 4924
rect 2588 4916 2596 4924
rect 5852 4916 5860 4924
rect 6524 4916 6532 4924
rect 7772 4936 7780 4944
rect 9148 4976 9156 4984
rect 8588 4956 8596 4964
rect 9820 4956 9828 4964
rect 10204 4956 10212 4964
rect 8108 4936 8116 4944
rect 8140 4936 8148 4944
rect 8412 4936 8420 4944
rect 9068 4936 9076 4944
rect 9580 4936 9588 4944
rect 9756 4936 9764 4944
rect 9932 4936 9940 4944
rect 8588 4916 8596 4924
rect 9612 4916 9620 4924
rect 668 4896 676 4904
rect 1100 4896 1108 4904
rect 1548 4896 1556 4904
rect 1772 4896 1780 4904
rect 1916 4896 1924 4904
rect 2796 4896 2804 4904
rect 3036 4896 3044 4904
rect 4092 4896 4100 4904
rect 4172 4896 4180 4904
rect 4460 4896 4468 4904
rect 4972 4896 4980 4904
rect 6844 4896 6852 4904
rect 7020 4896 7028 4904
rect 7436 4896 7444 4904
rect 7612 4896 7620 4904
rect 7660 4896 7668 4904
rect 9420 4896 9428 4904
rect 9612 4896 9620 4904
rect 10028 4896 10036 4904
rect 1100 4876 1108 4884
rect 3628 4876 3636 4884
rect 4620 4876 4628 4884
rect 5740 4876 5748 4884
rect 908 4856 916 4864
rect 3852 4856 3860 4864
rect 4796 4836 4804 4844
rect 6588 4836 6596 4844
rect 2140 4816 2148 4824
rect 5260 4816 5268 4824
rect 236 4796 244 4804
rect 9724 4756 9732 4764
rect 460 4736 468 4744
rect 1548 4736 1556 4744
rect 1884 4736 1892 4744
rect 2556 4736 2564 4744
rect 3964 4736 3972 4744
rect 5052 4736 5060 4744
rect 5820 4736 5828 4744
rect 6188 4736 6196 4744
rect 6572 4736 6580 4744
rect 7660 4736 7668 4744
rect 7820 4736 7828 4744
rect 7868 4736 7876 4744
rect 9388 4736 9396 4744
rect 9932 4736 9940 4744
rect 76 4716 84 4724
rect 908 4716 916 4724
rect 1548 4716 1556 4724
rect 1788 4716 1796 4724
rect 2508 4716 2516 4724
rect 2556 4716 2564 4724
rect 2700 4716 2708 4724
rect 2988 4716 2996 4724
rect 3836 4716 3844 4724
rect 4476 4716 4484 4724
rect 5196 4716 5204 4724
rect 5468 4716 5476 4724
rect 6300 4716 6308 4724
rect 6572 4716 6580 4724
rect 6588 4716 6596 4724
rect 6940 4716 6948 4724
rect 7372 4716 7380 4724
rect 7948 4716 7956 4724
rect 7964 4716 7972 4724
rect 8476 4716 8484 4724
rect 8588 4716 8596 4724
rect 9340 4716 9348 4724
rect 3564 4696 3572 4704
rect 3596 4696 3604 4704
rect 5180 4696 5188 4704
rect 5580 4696 5588 4704
rect 6508 4696 6516 4704
rect 7692 4696 7700 4704
rect 7932 4696 7940 4704
rect 7964 4696 7972 4704
rect 8636 4696 8644 4704
rect 8764 4696 8772 4704
rect 9676 4696 9684 4704
rect 12 4676 20 4684
rect 76 4676 84 4684
rect 908 4676 916 4684
rect 1148 4676 1156 4684
rect 1916 4676 1924 4684
rect 2364 4676 2372 4684
rect 2812 4676 2820 4684
rect 3372 4676 3380 4684
rect 3580 4676 3588 4684
rect 5532 4676 5540 4684
rect 5948 4676 5956 4684
rect 6588 4676 6596 4684
rect 6636 4676 6644 4684
rect 8908 4676 8916 4684
rect 9148 4676 9156 4684
rect 9596 4676 9604 4684
rect 9708 4676 9716 4684
rect 9916 4676 9924 4684
rect 10012 4676 10020 4684
rect 12 4636 20 4644
rect 668 4596 676 4604
rect 1916 4656 1924 4664
rect 2668 4656 2676 4664
rect 4460 4656 4468 4664
rect 5164 4656 5172 4664
rect 5724 4656 5732 4664
rect 7004 4656 7012 4664
rect 8508 4656 8516 4664
rect 8764 4656 8772 4664
rect 8908 4656 8916 4664
rect 8940 4656 8948 4664
rect 9196 4656 9204 4664
rect 2268 4636 2276 4644
rect 2524 4636 2532 4644
rect 3612 4636 3620 4644
rect 6124 4636 6132 4644
rect 8252 4636 8260 4644
rect 8764 4636 8772 4644
rect 10204 4636 10212 4644
rect 2252 4616 2260 4624
rect 2284 4616 2292 4624
rect 5164 4596 5172 4604
rect 9884 4596 9892 4604
rect 9900 4596 9908 4604
rect 2060 4576 2068 4584
rect 2268 4576 2276 4584
rect 3852 4576 3860 4584
rect 7756 4576 7764 4584
rect 8716 4576 8724 4584
rect 908 4556 916 4564
rect 3100 4556 3108 4564
rect 4156 4556 4164 4564
rect 4172 4556 4180 4564
rect 4732 4556 4740 4564
rect 5964 4556 5972 4564
rect 6108 4556 6116 4564
rect 7004 4556 7012 4564
rect 9228 4556 9236 4564
rect 236 4536 244 4544
rect 540 4536 548 4544
rect 1100 4536 1108 4544
rect 1148 4536 1156 4544
rect 1596 4536 1604 4544
rect 1692 4536 1700 4544
rect 2412 4536 2420 4544
rect 2444 4536 2452 4544
rect 2908 4536 2916 4544
rect 3372 4536 3380 4544
rect 3580 4536 3588 4544
rect 4348 4536 4356 4544
rect 4652 4536 4660 4544
rect 4732 4536 4740 4544
rect 5356 4536 5364 4544
rect 5740 4536 5748 4544
rect 6316 4536 6324 4544
rect 6620 4536 6628 4544
rect 7484 4536 7492 4544
rect 8028 4536 8036 4544
rect 8044 4536 8052 4544
rect 9004 4536 9012 4544
rect 9020 4536 9028 4544
rect 9772 4536 9780 4544
rect 2988 4516 2996 4524
rect 3932 4516 3940 4524
rect 6156 4516 6164 4524
rect 6700 4516 6708 4524
rect 6716 4516 6724 4524
rect 8156 4516 8164 4524
rect 8780 4516 8788 4524
rect 316 4496 324 4504
rect 668 4496 676 4504
rect 1420 4496 1428 4504
rect 2956 4496 2964 4504
rect 3148 4496 3156 4504
rect 3852 4496 3860 4504
rect 4076 4496 4084 4504
rect 4236 4496 4244 4504
rect 4748 4496 4756 4504
rect 5020 4496 5028 4504
rect 5308 4496 5316 4504
rect 5916 4496 5924 4504
rect 6492 4496 6500 4504
rect 7164 4496 7172 4504
rect 7276 4496 7284 4504
rect 8604 4496 8612 4504
rect 8892 4496 8900 4504
rect 9132 4496 9140 4504
rect 9660 4496 9668 4504
rect 9692 4496 9700 4504
rect 1548 4476 1556 4484
rect 2492 4476 2500 4484
rect 2780 4476 2788 4484
rect 2796 4476 2804 4484
rect 3356 4476 3364 4484
rect 3388 4476 3396 4484
rect 3836 4476 3844 4484
rect 4796 4476 4804 4484
rect 6140 4476 6148 4484
rect 6476 4476 6484 4484
rect 6748 4476 6756 4484
rect 7180 4476 7188 4484
rect 1612 4456 1620 4464
rect 1692 4456 1700 4464
rect 2268 4456 2276 4464
rect 2796 4456 2804 4464
rect 9884 4456 9892 4464
rect 684 4436 692 4444
rect 892 4436 900 4444
rect 2668 4436 2676 4444
rect 3164 4436 3172 4444
rect 7244 4436 7252 4444
rect 9164 4436 9172 4444
rect 1164 4376 1172 4384
rect 1580 4376 1588 4384
rect 2636 4356 2644 4364
rect 6796 4356 6804 4364
rect 7036 4356 7044 4364
rect 9500 4356 9508 4364
rect 908 4336 916 4344
rect 2796 4336 2804 4344
rect 3564 4336 3572 4344
rect 4012 4336 4020 4344
rect 5180 4336 5188 4344
rect 5644 4336 5652 4344
rect 6604 4336 6612 4344
rect 7852 4336 7860 4344
rect 572 4316 580 4324
rect 1644 4316 1652 4324
rect 2252 4316 2260 4324
rect 2332 4316 2340 4324
rect 2796 4316 2804 4324
rect 3596 4316 3604 4324
rect 3756 4316 3764 4324
rect 4332 4316 4340 4324
rect 4572 4316 4580 4324
rect 4716 4316 4724 4324
rect 5084 4316 5092 4324
rect 5436 4316 5444 4324
rect 5596 4316 5604 4324
rect 6364 4316 6372 4324
rect 7100 4316 7108 4324
rect 7468 4316 7476 4324
rect 8604 4316 8612 4324
rect 8924 4316 8932 4324
rect 9356 4316 9364 4324
rect 9852 4316 9860 4324
rect 1420 4296 1428 4304
rect 1740 4296 1748 4304
rect 2684 4296 2692 4304
rect 3388 4296 3396 4304
rect 3820 4296 3828 4304
rect 7244 4296 7252 4304
rect 7292 4296 7300 4304
rect 7324 4296 7332 4304
rect 7468 4296 7476 4304
rect 7708 4296 7716 4304
rect 8716 4296 8724 4304
rect 540 4276 548 4284
rect 908 4276 916 4284
rect 1020 4276 1028 4284
rect 2252 4276 2260 4284
rect 3148 4276 3156 4284
rect 3996 4276 4004 4284
rect 5724 4276 5732 4284
rect 6268 4276 6276 4284
rect 7628 4276 7636 4284
rect 7644 4276 7652 4284
rect 7676 4276 7684 4284
rect 8028 4276 8036 4284
rect 8556 4276 8564 4284
rect 8732 4276 8740 4284
rect 9132 4276 9140 4284
rect 9164 4276 9172 4284
rect 9228 4276 9236 4284
rect 9820 4276 9828 4284
rect 2700 4256 2708 4264
rect 3948 4256 3956 4264
rect 4076 4256 4084 4264
rect 5052 4256 5060 4264
rect 6668 4256 6676 4264
rect 7164 4256 7172 4264
rect 8300 4256 8308 4264
rect 9132 4256 9140 4264
rect 764 4236 772 4244
rect 1580 4236 1588 4244
rect 2588 4236 2596 4244
rect 3228 4236 3236 4244
rect 3404 4236 3412 4244
rect 4780 4236 4788 4244
rect 6140 4236 6148 4244
rect 6348 4236 6356 4244
rect 8332 4236 8340 4244
rect 8604 4236 8612 4244
rect 444 4216 452 4224
rect 5756 4216 5764 4224
rect 6476 4216 6484 4224
rect 7340 4216 7348 4224
rect 7548 4216 7556 4224
rect 7596 4216 7604 4224
rect 908 4196 916 4204
rect 2700 4196 2708 4204
rect 2732 4196 2740 4204
rect 6348 4196 6356 4204
rect 7180 4196 7188 4204
rect 7196 4196 7204 4204
rect 7260 4196 7268 4204
rect 10060 4196 10068 4204
rect 5148 4176 5156 4184
rect 8412 4176 8420 4184
rect 9132 4176 9140 4184
rect 9148 4176 9156 4184
rect 9500 4176 9508 4184
rect 2908 4156 2916 4164
rect 5964 4156 5972 4164
rect 6188 4156 6196 4164
rect 6828 4156 6836 4164
rect 7068 4156 7076 4164
rect 7340 4156 7348 4164
rect 7404 4156 7412 4164
rect 7420 4156 7428 4164
rect 8236 4156 8244 4164
rect 8972 4156 8980 4164
rect 9564 4156 9572 4164
rect 9916 4156 9924 4164
rect 220 4136 228 4144
rect 2012 4136 2020 4144
rect 2460 4136 2468 4144
rect 2492 4136 2500 4144
rect 3628 4136 3636 4144
rect 4652 4136 4660 4144
rect 4940 4136 4948 4144
rect 5068 4136 5076 4144
rect 5388 4136 5396 4144
rect 5740 4136 5748 4144
rect 6188 4136 6196 4144
rect 6748 4136 6756 4144
rect 8716 4136 8724 4144
rect 8732 4136 8740 4144
rect 9276 4136 9284 4144
rect 9548 4136 9556 4144
rect 1580 4116 1588 4124
rect 2796 4116 2804 4124
rect 3180 4116 3188 4124
rect 3372 4116 3380 4124
rect 6028 4116 6036 4124
rect 6700 4116 6708 4124
rect 7484 4116 7492 4124
rect 7708 4116 7716 4124
rect 7724 4116 7732 4124
rect 7868 4116 7876 4124
rect 8604 4116 8612 4124
rect 8892 4116 8900 4124
rect 9916 4116 9924 4124
rect 332 4096 340 4104
rect 524 4096 532 4104
rect 764 4096 772 4104
rect 1100 4096 1108 4104
rect 1228 4096 1236 4104
rect 3612 4096 3620 4104
rect 4044 4096 4052 4104
rect 4188 4096 4196 4104
rect 4572 4096 4580 4104
rect 4748 4096 4756 4104
rect 5708 4096 5716 4104
rect 6076 4096 6084 4104
rect 6172 4096 6180 4104
rect 6748 4096 6756 4104
rect 6892 4096 6900 4104
rect 7372 4096 7380 4104
rect 7628 4096 7636 4104
rect 8508 4096 8516 4104
rect 9884 4096 9892 4104
rect 652 4076 660 4084
rect 1196 4076 1204 4084
rect 2732 4076 2740 4084
rect 2876 4076 2884 4084
rect 3020 4076 3028 4084
rect 5756 4076 5764 4084
rect 6172 4076 6180 4084
rect 6780 4076 6788 4084
rect 7676 4076 7684 4084
rect 7708 4076 7716 4084
rect 7916 4076 7924 4084
rect 8812 4076 8820 4084
rect 9068 4076 9076 4084
rect 9516 4076 9524 4084
rect 9564 4076 9572 4084
rect 9916 4076 9924 4084
rect 236 4056 244 4064
rect 1612 4056 1620 4064
rect 3404 4056 3412 4064
rect 4156 4056 4164 4064
rect 5756 4056 5764 4064
rect 7548 4056 7556 4064
rect 9260 4056 9268 4064
rect 5356 4036 5364 4044
rect 7372 4036 7380 4044
rect 7692 4036 7700 4044
rect 76 4016 84 4024
rect 9612 4016 9620 4024
rect 5340 3976 5348 3984
rect 476 3936 484 3944
rect 8892 3956 8900 3964
rect 8988 3956 8996 3964
rect 9068 3956 9076 3964
rect 1228 3936 1236 3944
rect 1884 3936 1892 3944
rect 2284 3936 2292 3944
rect 2908 3936 2916 3944
rect 5004 3936 5012 3944
rect 5068 3936 5076 3944
rect 5132 3936 5140 3944
rect 5532 3936 5540 3944
rect 5548 3936 5556 3944
rect 5836 3936 5844 3944
rect 6012 3936 6020 3944
rect 6092 3936 6100 3944
rect 6140 3936 6148 3944
rect 6636 3936 6644 3944
rect 8524 3936 8532 3944
rect 8620 3936 8628 3944
rect 8860 3936 8868 3944
rect 428 3916 436 3924
rect 2876 3916 2884 3924
rect 2924 3916 2932 3924
rect 3372 3916 3380 3924
rect 3916 3916 3924 3924
rect 4380 3916 4388 3924
rect 5516 3916 5524 3924
rect 6156 3916 6164 3924
rect 6396 3916 6404 3924
rect 6828 3916 6836 3924
rect 7276 3916 7284 3924
rect 7388 3916 7396 3924
rect 9132 3916 9140 3924
rect 9228 3916 9236 3924
rect 1148 3896 1156 3904
rect 1548 3896 1556 3904
rect 2588 3896 2596 3904
rect 2716 3896 2724 3904
rect 3196 3896 3204 3904
rect 4060 3896 4068 3904
rect 4652 3896 4660 3904
rect 6620 3896 6628 3904
rect 7260 3896 7268 3904
rect 7660 3896 7668 3904
rect 8460 3896 8468 3904
rect 9116 3896 9124 3904
rect 9260 3896 9268 3904
rect 9660 3896 9668 3904
rect 220 3876 228 3884
rect 236 3876 244 3884
rect 332 3876 340 3884
rect 1020 3876 1028 3884
rect 1196 3876 1204 3884
rect 1596 3876 1604 3884
rect 1740 3876 1748 3884
rect 1756 3876 1764 3884
rect 3132 3876 3140 3884
rect 3916 3876 3924 3884
rect 4300 3876 4308 3884
rect 4844 3876 4852 3884
rect 5628 3876 5636 3884
rect 5644 3876 5652 3884
rect 5868 3876 5876 3884
rect 6012 3876 6020 3884
rect 6508 3876 6516 3884
rect 6652 3876 6660 3884
rect 6812 3876 6820 3884
rect 7132 3876 7140 3884
rect 7260 3876 7268 3884
rect 7708 3876 7716 3884
rect 8444 3876 8452 3884
rect 8764 3876 8772 3884
rect 9852 3876 9860 3884
rect 10044 3876 10052 3884
rect 284 3856 292 3864
rect 636 3856 644 3864
rect 668 3856 676 3864
rect 1788 3856 1796 3864
rect 3164 3856 3172 3864
rect 3628 3856 3636 3864
rect 5532 3856 5540 3864
rect 6092 3856 6100 3864
rect 6156 3856 6164 3864
rect 6796 3856 6804 3864
rect 7660 3856 7668 3864
rect 8300 3856 8308 3864
rect 8732 3856 8740 3864
rect 9164 3856 9172 3864
rect 300 3836 308 3844
rect 1004 3836 1012 3844
rect 1020 3836 1028 3844
rect 5564 3836 5572 3844
rect 7100 3836 7108 3844
rect 7836 3836 7844 3844
rect 9100 3836 9108 3844
rect 9116 3836 9124 3844
rect 2124 3816 2132 3824
rect 3644 3816 3652 3824
rect 236 3796 244 3804
rect 2012 3796 2020 3804
rect 2524 3796 2532 3804
rect 4300 3796 4308 3804
rect 7820 3796 7828 3804
rect 9468 3796 9476 3804
rect 9916 3796 9924 3804
rect 220 3776 228 3784
rect 3964 3776 3972 3784
rect 1804 3756 1812 3764
rect 2012 3756 2020 3764
rect 2028 3756 2036 3764
rect 2412 3756 2420 3764
rect 4044 3756 4052 3764
rect 6428 3776 6436 3784
rect 6988 3776 6996 3784
rect 7020 3776 7028 3784
rect 7436 3776 7444 3784
rect 8316 3776 8324 3784
rect 8764 3776 8772 3784
rect 5180 3756 5188 3764
rect 6588 3756 6596 3764
rect 6860 3756 6868 3764
rect 1356 3736 1364 3744
rect 1740 3736 1748 3744
rect 2524 3736 2532 3744
rect 2588 3736 2596 3744
rect 2684 3736 2692 3744
rect 3164 3736 3172 3744
rect 3420 3736 3428 3744
rect 4108 3736 4116 3744
rect 5420 3736 5428 3744
rect 5548 3736 5556 3744
rect 6188 3736 6196 3744
rect 7052 3736 7060 3744
rect 7068 3736 7076 3744
rect 7340 3736 7348 3744
rect 7852 3736 7860 3744
rect 8460 3756 8468 3764
rect 8476 3756 8484 3764
rect 8700 3736 8708 3744
rect 8908 3736 8916 3744
rect 9292 3736 9300 3744
rect 9612 3736 9620 3744
rect 9852 3736 9860 3744
rect 2332 3716 2340 3724
rect 2460 3716 2468 3724
rect 3436 3716 3444 3724
rect 4300 3716 4308 3724
rect 6956 3716 6964 3724
rect 6988 3716 6996 3724
rect 1116 3696 1124 3704
rect 1596 3696 1604 3704
rect 2636 3696 2644 3704
rect 3180 3696 3188 3704
rect 3772 3696 3780 3704
rect 4076 3696 4084 3704
rect 4316 3696 4324 3704
rect 4524 3696 4532 3704
rect 4748 3696 4756 3704
rect 5532 3696 5540 3704
rect 5756 3696 5764 3704
rect 6172 3696 6180 3704
rect 7484 3696 7492 3704
rect 7692 3696 7700 3704
rect 9468 3696 9476 3704
rect 1340 3676 1348 3684
rect 3804 3676 3812 3684
rect 7884 3676 7892 3684
rect 8236 3676 8244 3684
rect 1132 3656 1140 3664
rect 1756 3656 1764 3664
rect 2236 3656 2244 3664
rect 5900 3636 5908 3644
rect 3740 3616 3748 3624
rect 8140 3616 8148 3624
rect 2588 3596 2596 3604
rect 1100 3556 1108 3564
rect 4572 3556 4580 3564
rect 7708 3556 7716 3564
rect 9020 3556 9028 3564
rect 332 3536 340 3544
rect 5788 3536 5796 3544
rect 5900 3536 5908 3544
rect 6124 3536 6132 3544
rect 6636 3536 6644 3544
rect 7612 3536 7620 3544
rect 7708 3536 7716 3544
rect 7948 3536 7956 3544
rect 8348 3536 8356 3544
rect 9708 3536 9716 3544
rect 92 3516 100 3524
rect 1628 3516 1636 3524
rect 2028 3516 2036 3524
rect 2492 3516 2500 3524
rect 2524 3516 2532 3524
rect 3388 3516 3396 3524
rect 3804 3516 3812 3524
rect 5148 3516 5156 3524
rect 5804 3516 5812 3524
rect 6860 3516 6868 3524
rect 7804 3516 7812 3524
rect 7820 3516 7828 3524
rect 8348 3516 8356 3524
rect 9388 3516 9396 3524
rect 9900 3516 9908 3524
rect 10092 3516 10100 3524
rect 316 3496 324 3504
rect 908 3496 916 3504
rect 1340 3496 1348 3504
rect 1404 3496 1412 3504
rect 3356 3496 3364 3504
rect 3372 3496 3380 3504
rect 3996 3496 4004 3504
rect 4780 3496 4788 3504
rect 6572 3496 6580 3504
rect 7372 3496 7380 3504
rect 7708 3496 7716 3504
rect 8508 3496 8516 3504
rect 9324 3496 9332 3504
rect 444 3476 452 3484
rect 892 3476 900 3484
rect 2220 3476 2228 3484
rect 2716 3476 2724 3484
rect 2972 3476 2980 3484
rect 3148 3476 3156 3484
rect 3388 3476 3396 3484
rect 3580 3476 3588 3484
rect 4476 3476 4484 3484
rect 4556 3476 4564 3484
rect 4796 3476 4804 3484
rect 5324 3476 5332 3484
rect 5788 3476 5796 3484
rect 6044 3476 6052 3484
rect 6140 3476 6148 3484
rect 6364 3476 6372 3484
rect 6428 3476 6436 3484
rect 7132 3476 7140 3484
rect 7228 3476 7236 3484
rect 7500 3476 7508 3484
rect 7532 3476 7540 3484
rect 8300 3476 8308 3484
rect 8908 3476 8916 3484
rect 8972 3476 8980 3484
rect 9132 3476 9140 3484
rect 9676 3476 9684 3484
rect 220 3456 228 3464
rect 1132 3456 1140 3464
rect 1788 3456 1796 3464
rect 1820 3456 1828 3464
rect 1772 3436 1780 3444
rect 2220 3436 2228 3444
rect 2236 3436 2244 3444
rect 3148 3436 3156 3444
rect 3628 3456 3636 3464
rect 3868 3456 3876 3464
rect 4284 3456 4292 3464
rect 4508 3456 4516 3464
rect 3996 3436 4004 3444
rect 4012 3436 4020 3444
rect 4236 3436 4244 3444
rect 5324 3456 5332 3464
rect 5836 3456 5844 3464
rect 7356 3456 7364 3464
rect 7692 3456 7700 3464
rect 8364 3456 8372 3464
rect 4604 3436 4612 3444
rect 4988 3436 4996 3444
rect 6860 3436 6868 3444
rect 7388 3436 7396 3444
rect 8876 3436 8884 3444
rect 9068 3436 9076 3444
rect 332 3416 340 3424
rect 3180 3416 3188 3424
rect 6764 3416 6772 3424
rect 4316 3396 4324 3404
rect 6620 3396 6628 3404
rect 2012 3376 2020 3384
rect 5612 3376 5620 3384
rect 5756 3376 5764 3384
rect 6060 3376 6068 3384
rect 6108 3376 6116 3384
rect 6156 3376 6164 3384
rect 7180 3376 7188 3384
rect 7404 3376 7412 3384
rect 8252 3376 8260 3384
rect 1244 3356 1252 3364
rect 2156 3356 2164 3364
rect 2828 3356 2836 3364
rect 2844 3356 2852 3364
rect 3180 3356 3188 3364
rect 3404 3356 3412 3364
rect 3852 3356 3860 3364
rect 4988 3356 4996 3364
rect 5500 3356 5508 3364
rect 5548 3356 5556 3364
rect 6012 3356 6020 3364
rect 7980 3356 7988 3364
rect 8124 3356 8132 3364
rect 9372 3356 9380 3364
rect 9532 3356 9540 3364
rect 684 3336 692 3344
rect 1132 3336 1140 3344
rect 1596 3336 1604 3344
rect 2108 3336 2116 3344
rect 4172 3336 4180 3344
rect 4316 3336 4324 3344
rect 4524 3336 4532 3344
rect 4620 3336 4628 3344
rect 5084 3336 5092 3344
rect 5388 3336 5396 3344
rect 6140 3336 6148 3344
rect 6188 3336 6196 3344
rect 6204 3336 6212 3344
rect 6540 3336 6548 3344
rect 6908 3336 6916 3344
rect 7068 3336 7076 3344
rect 7452 3336 7460 3344
rect 8172 3336 8180 3344
rect 8364 3336 8372 3344
rect 988 3316 996 3324
rect 1580 3316 1588 3324
rect 3356 3316 3364 3324
rect 4604 3316 4612 3324
rect 5532 3316 5540 3324
rect 6268 3316 6276 3324
rect 7132 3316 7140 3324
rect 7276 3316 7284 3324
rect 7644 3316 7652 3324
rect 7964 3316 7972 3324
rect 8604 3316 8612 3324
rect 8844 3336 8852 3344
rect 9388 3336 9396 3344
rect 10028 3336 10036 3344
rect 236 3296 244 3304
rect 460 3296 468 3304
rect 1884 3296 1892 3304
rect 3100 3296 3108 3304
rect 3180 3296 3188 3304
rect 4316 3296 4324 3304
rect 4556 3296 4564 3304
rect 5180 3296 5188 3304
rect 5404 3296 5412 3304
rect 6236 3296 6244 3304
rect 6284 3296 6292 3304
rect 6508 3296 6516 3304
rect 6716 3296 6724 3304
rect 6844 3296 6852 3304
rect 7276 3296 7284 3304
rect 7516 3296 7524 3304
rect 7948 3296 7956 3304
rect 9532 3296 9540 3304
rect 1612 3276 1620 3284
rect 2284 3276 2292 3284
rect 2380 3276 2388 3284
rect 2844 3276 2852 3284
rect 3244 3276 3252 3284
rect 3740 3276 3748 3284
rect 3820 3276 3828 3284
rect 4060 3276 4068 3284
rect 6204 3276 6212 3284
rect 1132 3256 1140 3264
rect 1244 3256 1252 3264
rect 3916 3256 3924 3264
rect 6620 3256 6628 3264
rect 6876 3256 6884 3264
rect 6060 3236 6068 3244
rect 1596 3196 1604 3204
rect 3052 3196 3060 3204
rect 4620 3176 4628 3184
rect 5036 3176 5044 3184
rect 2380 3156 2388 3164
rect 8988 3156 8996 3164
rect 2524 3136 2532 3144
rect 3868 3136 3876 3144
rect 4220 3136 4228 3144
rect 4572 3136 4580 3144
rect 5116 3136 5124 3144
rect 5484 3136 5492 3144
rect 5884 3136 5892 3144
rect 6636 3136 6644 3144
rect 6844 3136 6852 3144
rect 10076 3136 10084 3144
rect 652 3116 660 3124
rect 1084 3116 1092 3124
rect 1212 3116 1220 3124
rect 2460 3116 2468 3124
rect 2956 3116 2964 3124
rect 2972 3116 2980 3124
rect 3612 3116 3620 3124
rect 3772 3116 3780 3124
rect 4060 3116 4068 3124
rect 4492 3116 4500 3124
rect 4988 3116 4996 3124
rect 5244 3116 5252 3124
rect 5356 3116 5364 3124
rect 5388 3116 5396 3124
rect 7852 3116 7860 3124
rect 8076 3116 8084 3124
rect 9196 3116 9204 3124
rect 9292 3116 9300 3124
rect 10268 3116 10276 3124
rect 684 3096 692 3104
rect 2428 3096 2436 3104
rect 2876 3096 2884 3104
rect 5148 3096 5156 3104
rect 5564 3096 5572 3104
rect 6172 3096 6180 3104
rect 6876 3096 6884 3104
rect 8588 3096 8596 3104
rect 9244 3096 9252 3104
rect 9276 3096 9284 3104
rect 1244 3076 1252 3084
rect 2412 3076 2420 3084
rect 2748 3076 2756 3084
rect 3548 3076 3556 3084
rect 3756 3076 3764 3084
rect 4204 3076 4212 3084
rect 4284 3076 4292 3084
rect 4588 3076 4596 3084
rect 4620 3076 4628 3084
rect 4748 3076 4756 3084
rect 5180 3076 5188 3084
rect 5388 3076 5396 3084
rect 5436 3076 5444 3084
rect 5724 3076 5732 3084
rect 5948 3076 5956 3084
rect 6076 3076 6084 3084
rect 6892 3076 6900 3084
rect 7548 3076 7556 3084
rect 1164 3056 1172 3064
rect 1180 3056 1188 3064
rect 1212 3056 1220 3064
rect 1612 3056 1620 3064
rect 2076 3056 2084 3064
rect 2220 3056 2228 3064
rect 2540 3056 2548 3064
rect 4156 3056 4164 3064
rect 4556 3056 4564 3064
rect 4940 3056 4948 3064
rect 5372 3056 5380 3064
rect 6908 3056 6916 3064
rect 7356 3056 7364 3064
rect 8412 3076 8420 3084
rect 9100 3076 9108 3084
rect 9260 3076 9268 3084
rect 10028 3076 10036 3084
rect 10092 3056 10100 3064
rect 204 2996 212 3004
rect 2156 3036 2164 3044
rect 2716 3036 2724 3044
rect 3212 3036 3220 3044
rect 4348 3036 4356 3044
rect 4476 3036 4484 3044
rect 4540 3036 4548 3044
rect 4908 3036 4916 3044
rect 4972 3036 4980 3044
rect 5036 3036 5044 3044
rect 6092 3036 6100 3044
rect 6332 3036 6340 3044
rect 8108 3036 8116 3044
rect 8908 3036 8916 3044
rect 9020 3036 9028 3044
rect 2556 3016 2564 3024
rect 3164 3016 3172 3024
rect 4940 3016 4948 3024
rect 6348 3016 6356 3024
rect 1260 2996 1268 3004
rect 2732 2996 2740 3004
rect 2828 2996 2836 3004
rect 2844 2996 2852 3004
rect 6988 2996 6996 3004
rect 2652 2976 2660 2984
rect 3084 2976 3092 2984
rect 4700 2976 4708 2984
rect 6140 2976 6148 2984
rect 7676 2976 7684 2984
rect 7852 2976 7860 2984
rect 9308 2976 9316 2984
rect 9612 2976 9620 2984
rect 652 2956 660 2964
rect 1628 2956 1636 2964
rect 2668 2956 2676 2964
rect 3244 2956 3252 2964
rect 4236 2956 4244 2964
rect 4908 2956 4916 2964
rect 6124 2956 6132 2964
rect 300 2936 308 2944
rect 444 2936 452 2944
rect 668 2936 676 2944
rect 1420 2916 1428 2924
rect 2652 2936 2660 2944
rect 3196 2936 3204 2944
rect 3564 2936 3572 2944
rect 5324 2936 5332 2944
rect 5724 2936 5732 2944
rect 5996 2936 6004 2944
rect 6572 2956 6580 2964
rect 6716 2956 6724 2964
rect 7628 2956 7636 2964
rect 8332 2956 8340 2964
rect 6268 2936 6276 2944
rect 6588 2936 6596 2944
rect 6812 2936 6820 2944
rect 6892 2936 6900 2944
rect 7052 2936 7060 2944
rect 7516 2936 7524 2944
rect 9132 2936 9140 2944
rect 9372 2936 9380 2944
rect 9708 2936 9716 2944
rect 9932 2936 9940 2944
rect 2332 2916 2340 2924
rect 3788 2916 3796 2924
rect 3948 2916 3956 2924
rect 6604 2916 6612 2924
rect 7308 2916 7316 2924
rect 7948 2916 7956 2924
rect 8028 2916 8036 2924
rect 8540 2916 8548 2924
rect 8556 2916 8564 2924
rect 9676 2916 9684 2924
rect 428 2896 436 2904
rect 668 2896 676 2904
rect 844 2896 852 2904
rect 972 2896 980 2904
rect 2012 2896 2020 2904
rect 2860 2896 2868 2904
rect 2956 2896 2964 2904
rect 3100 2896 3108 2904
rect 3820 2896 3828 2904
rect 4220 2896 4228 2904
rect 4348 2896 4356 2904
rect 4940 2896 4948 2904
rect 5772 2896 5780 2904
rect 6028 2896 6036 2904
rect 6220 2896 6228 2904
rect 6348 2896 6356 2904
rect 7244 2896 7252 2904
rect 7468 2896 7476 2904
rect 7868 2896 7876 2904
rect 8268 2896 8276 2904
rect 8348 2896 8356 2904
rect 8380 2896 8388 2904
rect 9052 2896 9060 2904
rect 9228 2896 9236 2904
rect 9676 2896 9684 2904
rect 9916 2896 9924 2904
rect 764 2876 772 2884
rect 1596 2876 1604 2884
rect 1836 2876 1844 2884
rect 3740 2876 3748 2884
rect 4908 2876 4916 2884
rect 6172 2876 6180 2884
rect 7420 2876 7428 2884
rect 1548 2856 1556 2864
rect 1996 2856 2004 2864
rect 3356 2856 3364 2864
rect 1180 2836 1188 2844
rect 2236 2816 2244 2824
rect 7884 2856 7892 2864
rect 4268 2836 4276 2844
rect 7500 2836 7508 2844
rect 1548 2796 1556 2804
rect 6684 2796 6692 2804
rect 9516 2796 9524 2804
rect 9916 2796 9924 2804
rect 2332 2776 2340 2784
rect 2924 2776 2932 2784
rect 4316 2776 4324 2784
rect 6732 2776 6740 2784
rect 1260 2756 1268 2764
rect 2716 2756 2724 2764
rect 4652 2756 4660 2764
rect 4876 2756 4884 2764
rect 6732 2756 6740 2764
rect 7660 2756 7668 2764
rect 620 2736 628 2744
rect 1084 2736 1092 2744
rect 3100 2736 3108 2744
rect 4268 2736 4276 2744
rect 5180 2736 5188 2744
rect 6620 2736 6628 2744
rect 7596 2736 7604 2744
rect 7612 2736 7620 2744
rect 8540 2736 8548 2744
rect 8716 2736 8724 2744
rect 1660 2716 1668 2724
rect 2860 2716 2868 2724
rect 2924 2716 2932 2724
rect 3212 2716 3220 2724
rect 3788 2716 3796 2724
rect 4028 2716 4036 2724
rect 4716 2716 4724 2724
rect 6172 2716 6180 2724
rect 6332 2716 6340 2724
rect 6732 2716 6740 2724
rect 6748 2716 6756 2724
rect 6812 2716 6820 2724
rect 8924 2716 8932 2724
rect 9308 2716 9316 2724
rect 9964 2716 9972 2724
rect 9980 2716 9988 2724
rect 2236 2696 2244 2704
rect 3596 2696 3604 2704
rect 4108 2696 4116 2704
rect 4124 2696 4132 2704
rect 4236 2696 4244 2704
rect 4284 2696 4292 2704
rect 4956 2696 4964 2704
rect 6604 2696 6612 2704
rect 7116 2696 7124 2704
rect 7196 2696 7204 2704
rect 7676 2696 7684 2704
rect 220 2676 228 2684
rect 956 2676 964 2684
rect 1132 2676 1140 2684
rect 1260 2676 1268 2684
rect 1644 2676 1652 2684
rect 2188 2676 2196 2684
rect 2252 2676 2260 2684
rect 2476 2676 2484 2684
rect 3580 2676 3588 2684
rect 3596 2676 3604 2684
rect 4300 2676 4308 2684
rect 220 2656 228 2664
rect 1996 2656 2004 2664
rect 2124 2656 2132 2664
rect 3132 2656 3140 2664
rect 4108 2656 4116 2664
rect 4604 2676 4612 2684
rect 5612 2676 5620 2684
rect 5756 2676 5764 2684
rect 5852 2676 5860 2684
rect 7692 2676 7700 2684
rect 7852 2676 7860 2684
rect 8716 2676 8724 2684
rect 9004 2676 9012 2684
rect 9836 2676 9844 2684
rect 4476 2656 4484 2664
rect 5724 2656 5732 2664
rect 6156 2656 6164 2664
rect 9484 2656 9492 2664
rect 1788 2636 1796 2644
rect 1820 2636 1828 2644
rect 3180 2636 3188 2644
rect 3356 2636 3364 2644
rect 5388 2636 5396 2644
rect 7452 2636 7460 2644
rect 7484 2636 7492 2644
rect 7660 2636 7668 2644
rect 8956 2636 8964 2644
rect 9196 2636 9204 2644
rect 220 2616 228 2624
rect 1356 2616 1364 2624
rect 1660 2616 1668 2624
rect 4748 2616 4756 2624
rect 7500 2616 7508 2624
rect 1132 2596 1140 2604
rect 3580 2596 3588 2604
rect 4300 2596 4308 2604
rect 6636 2596 6644 2604
rect 7916 2596 7924 2604
rect 8444 2596 8452 2604
rect 9964 2596 9972 2604
rect 700 2576 708 2584
rect 4460 2576 4468 2584
rect 9628 2576 9636 2584
rect 1116 2556 1124 2564
rect 2748 2556 2756 2564
rect 3548 2556 3556 2564
rect 4300 2556 4308 2564
rect 4748 2556 4756 2564
rect 5132 2556 5140 2564
rect 5980 2556 5988 2564
rect 7372 2556 7380 2564
rect 7548 2556 7556 2564
rect 8540 2556 8548 2564
rect 8812 2556 8820 2564
rect 9148 2556 9156 2564
rect 76 2536 84 2544
rect 428 2536 436 2544
rect 556 2536 564 2544
rect 748 2536 756 2544
rect 1244 2536 1252 2544
rect 1292 2536 1300 2544
rect 1788 2536 1796 2544
rect 1836 2536 1844 2544
rect 1996 2536 2004 2544
rect 2220 2536 2228 2544
rect 2348 2536 2356 2544
rect 2380 2536 2388 2544
rect 2796 2536 2804 2544
rect 3052 2536 3060 2544
rect 3068 2536 3076 2544
rect 4076 2536 4084 2544
rect 4988 2536 4996 2544
rect 5004 2536 5012 2544
rect 5756 2536 5764 2544
rect 5964 2536 5972 2544
rect 6204 2536 6212 2544
rect 6748 2536 6756 2544
rect 6876 2536 6884 2544
rect 6956 2536 6964 2544
rect 7036 2536 7044 2544
rect 7644 2536 7652 2544
rect 8300 2536 8308 2544
rect 8476 2536 8484 2544
rect 8700 2536 8708 2544
rect 9244 2536 9252 2544
rect 9676 2536 9684 2544
rect 2252 2516 2260 2524
rect 5596 2516 5604 2524
rect 5772 2516 5780 2524
rect 5916 2516 5924 2524
rect 8252 2516 8260 2524
rect 9020 2516 9028 2524
rect 9212 2516 9220 2524
rect 9260 2516 9268 2524
rect 476 2496 484 2504
rect 1228 2496 1236 2504
rect 1276 2496 1284 2504
rect 1804 2496 1812 2504
rect 2492 2496 2500 2504
rect 2844 2496 2852 2504
rect 3628 2496 3636 2504
rect 4284 2496 4292 2504
rect 4988 2496 4996 2504
rect 5036 2496 5044 2504
rect 5084 2496 5092 2504
rect 5964 2496 5972 2504
rect 6188 2496 6196 2504
rect 6972 2496 6980 2504
rect 7164 2496 7172 2504
rect 7676 2496 7684 2504
rect 9308 2496 9316 2504
rect 204 2476 212 2484
rect 796 2476 804 2484
rect 908 2476 916 2484
rect 988 2476 996 2484
rect 3420 2476 3428 2484
rect 5516 2476 5524 2484
rect 7148 2476 7156 2484
rect 7420 2476 7428 2484
rect 9612 2476 9620 2484
rect 3100 2436 3108 2444
rect 6092 2436 6100 2444
rect 6172 2436 6180 2444
rect 428 2396 436 2404
rect 460 2376 468 2384
rect 7180 2376 7188 2384
rect 652 2356 660 2364
rect 3740 2356 3748 2364
rect 4684 2356 4692 2364
rect 5132 2356 5140 2364
rect 796 2336 804 2344
rect 2172 2336 2180 2344
rect 3948 2336 3956 2344
rect 4060 2336 4068 2344
rect 6620 2336 6628 2344
rect 7916 2336 7924 2344
rect 7948 2336 7956 2344
rect 9276 2336 9284 2344
rect 652 2316 660 2324
rect 1884 2316 1892 2324
rect 1900 2316 1908 2324
rect 2092 2316 2100 2324
rect 2460 2316 2468 2324
rect 2860 2316 2868 2324
rect 3180 2316 3188 2324
rect 3500 2316 3508 2324
rect 3612 2316 3620 2324
rect 5148 2316 5156 2324
rect 6252 2316 6260 2324
rect 6700 2316 6708 2324
rect 6732 2316 6740 2324
rect 7324 2316 7332 2324
rect 7900 2316 7908 2324
rect 7916 2316 7924 2324
rect 9884 2316 9892 2324
rect 1644 2296 1652 2304
rect 1756 2296 1764 2304
rect 1772 2296 1780 2304
rect 2028 2296 2036 2304
rect 2236 2296 2244 2304
rect 2268 2296 2276 2304
rect 2524 2296 2532 2304
rect 4924 2296 4932 2304
rect 4956 2296 4964 2304
rect 5340 2296 5348 2304
rect 5420 2296 5428 2304
rect 6236 2296 6244 2304
rect 7164 2296 7172 2304
rect 7692 2296 7700 2304
rect 8140 2296 8148 2304
rect 9516 2296 9524 2304
rect 9836 2296 9844 2304
rect 1324 2276 1332 2284
rect 1564 2276 1572 2284
rect 1868 2276 1876 2284
rect 2092 2276 2100 2284
rect 2188 2276 2196 2284
rect 2780 2276 2788 2284
rect 2796 2276 2804 2284
rect 3084 2276 3092 2284
rect 3212 2276 3220 2284
rect 3484 2276 3492 2284
rect 3628 2276 3636 2284
rect 4076 2276 4084 2284
rect 4364 2276 4372 2284
rect 4780 2276 4788 2284
rect 4908 2276 4916 2284
rect 6972 2276 6980 2284
rect 7308 2276 7316 2284
rect 7340 2276 7348 2284
rect 7996 2276 8004 2284
rect 8300 2276 8308 2284
rect 9148 2276 9156 2284
rect 9292 2276 9300 2284
rect 9484 2276 9492 2284
rect 9932 2276 9940 2284
rect 684 2256 692 2264
rect 1292 2256 1300 2264
rect 2108 2256 2116 2264
rect 3308 2256 3316 2264
rect 3356 2256 3364 2264
rect 3468 2256 3476 2264
rect 3580 2256 3588 2264
rect 4940 2256 4948 2264
rect 5228 2256 5236 2264
rect 6012 2256 6020 2264
rect 6140 2256 6148 2264
rect 6924 2256 6932 2264
rect 7068 2256 7076 2264
rect 7084 2256 7092 2264
rect 7164 2256 7172 2264
rect 9516 2256 9524 2264
rect 1612 2236 1620 2244
rect 3404 2236 3412 2244
rect 3420 2236 3428 2244
rect 4828 2236 4836 2244
rect 8156 2236 8164 2244
rect 8988 2236 8996 2244
rect 2652 2216 2660 2224
rect 7068 2216 7076 2224
rect 7708 2216 7716 2224
rect 1820 2196 1828 2204
rect 3132 2196 3140 2204
rect 5564 2196 5572 2204
rect 8412 2196 8420 2204
rect 700 2176 708 2184
rect 972 2176 980 2184
rect 1004 2176 1012 2184
rect 1660 2156 1668 2164
rect 1676 2156 1684 2164
rect 2572 2156 2580 2164
rect 3004 2156 3012 2164
rect 5532 2176 5540 2184
rect 4028 2156 4036 2164
rect 4604 2156 4612 2164
rect 6092 2156 6100 2164
rect 7100 2156 7108 2164
rect 7116 2156 7124 2164
rect 7132 2156 7140 2164
rect 9004 2156 9012 2164
rect 9452 2156 9460 2164
rect 9484 2156 9492 2164
rect 9884 2156 9892 2164
rect 220 2136 228 2144
rect 924 2136 932 2144
rect 1004 2136 1012 2144
rect 1260 2136 1268 2144
rect 3532 2136 3540 2144
rect 3564 2136 3572 2144
rect 3820 2136 3828 2144
rect 4044 2136 4052 2144
rect 4300 2136 4308 2144
rect 4556 2136 4564 2144
rect 4796 2136 4804 2144
rect 6380 2136 6388 2144
rect 7020 2136 7028 2144
rect 7052 2136 7060 2144
rect 7404 2136 7412 2144
rect 7964 2136 7972 2144
rect 8364 2136 8372 2144
rect 8668 2136 8676 2144
rect 9132 2136 9140 2144
rect 9804 2136 9812 2144
rect 668 2116 676 2124
rect 4508 2116 4516 2124
rect 5740 2116 5748 2124
rect 5852 2116 5860 2124
rect 5884 2116 5892 2124
rect 6876 2116 6884 2124
rect 1548 2096 1556 2104
rect 1996 2096 2004 2104
rect 2060 2096 2068 2104
rect 5724 2096 5732 2104
rect 6828 2096 6836 2104
rect 7244 2096 7252 2104
rect 7260 2096 7268 2104
rect 7548 2096 7556 2104
rect 7692 2096 7700 2104
rect 7788 2096 7796 2104
rect 8380 2096 8388 2104
rect 9148 2096 9156 2104
rect 3004 2076 3012 2084
rect 4028 2076 4036 2084
rect 6396 2076 6404 2084
rect 7212 2076 7220 2084
rect 7260 2076 7268 2084
rect 7484 2076 7492 2084
rect 956 2056 964 2064
rect 4940 2056 4948 2064
rect 220 2016 228 2024
rect 508 2016 516 2024
rect 3404 2016 3412 2024
rect 6956 2016 6964 2024
rect 8476 2016 8484 2024
rect 9468 1976 9476 1984
rect 972 1956 980 1964
rect 1004 1956 1012 1964
rect 2220 1956 2228 1964
rect 3404 1956 3412 1964
rect 3836 1956 3844 1964
rect 4076 1956 4084 1964
rect 7628 1956 7636 1964
rect 8348 1956 8356 1964
rect 9228 1956 9236 1964
rect 988 1936 996 1944
rect 1628 1916 1636 1924
rect 1788 1916 1796 1924
rect 1900 1936 1908 1944
rect 2124 1936 2132 1944
rect 3148 1936 3156 1944
rect 4828 1936 4836 1944
rect 6812 1936 6820 1944
rect 8588 1936 8596 1944
rect 2252 1916 2260 1924
rect 2444 1916 2452 1924
rect 2828 1916 2836 1924
rect 4284 1916 4292 1924
rect 4492 1916 4500 1924
rect 4844 1916 4852 1924
rect 4988 1916 4996 1924
rect 5692 1916 5700 1924
rect 5948 1916 5956 1924
rect 6220 1916 6228 1924
rect 6684 1916 6692 1924
rect 6796 1916 6804 1924
rect 7660 1916 7668 1924
rect 7820 1916 7828 1924
rect 7900 1916 7908 1924
rect 8812 1916 8820 1924
rect 9452 1936 9460 1944
rect 524 1896 532 1904
rect 2668 1896 2676 1904
rect 3164 1896 3172 1904
rect 300 1876 308 1884
rect 636 1876 644 1884
rect 668 1876 676 1884
rect 764 1876 772 1884
rect 844 1876 852 1884
rect 860 1876 868 1884
rect 988 1876 996 1884
rect 1196 1876 1204 1884
rect 4348 1876 4356 1884
rect 4444 1876 4452 1884
rect 5980 1896 5988 1904
rect 6764 1896 6772 1904
rect 7372 1896 7380 1904
rect 7628 1896 7636 1904
rect 8124 1896 8132 1904
rect 8812 1896 8820 1904
rect 9388 1896 9396 1904
rect 9900 1896 9908 1904
rect 10108 1896 10116 1904
rect 4812 1876 4820 1884
rect 5324 1876 5332 1884
rect 5468 1876 5476 1884
rect 6492 1876 6500 1884
rect 6620 1876 6628 1884
rect 6716 1876 6724 1884
rect 7340 1876 7348 1884
rect 7676 1876 7684 1884
rect 7884 1876 7892 1884
rect 8908 1876 8916 1884
rect 9244 1876 9252 1884
rect 1836 1856 1844 1864
rect 2652 1856 2660 1864
rect 3916 1856 3924 1864
rect 4700 1856 4708 1864
rect 5788 1856 5796 1864
rect 6700 1856 6708 1864
rect 7036 1856 7044 1864
rect 8028 1856 8036 1864
rect 8556 1856 8564 1864
rect 4300 1836 4308 1844
rect 4332 1836 4340 1844
rect 4348 1836 4356 1844
rect 5948 1836 5956 1844
rect 7964 1836 7972 1844
rect 8444 1836 8452 1844
rect 236 1816 244 1824
rect 428 1816 436 1824
rect 1996 1816 2004 1824
rect 2460 1816 2468 1824
rect 3004 1816 3012 1824
rect 4284 1816 4292 1824
rect 6156 1816 6164 1824
rect 7804 1816 7812 1824
rect 988 1796 996 1804
rect 1132 1796 1140 1804
rect 1356 1796 1364 1804
rect 1900 1796 1908 1804
rect 3836 1796 3844 1804
rect 4700 1796 4708 1804
rect 7788 1796 7796 1804
rect 7804 1796 7812 1804
rect 9900 1796 9908 1804
rect 7692 1776 7700 1784
rect 10060 1776 10068 1784
rect 428 1756 436 1764
rect 668 1756 676 1764
rect 956 1756 964 1764
rect 1612 1756 1620 1764
rect 2460 1756 2468 1764
rect 3404 1756 3412 1764
rect 5196 1756 5204 1764
rect 8364 1756 8372 1764
rect 8540 1756 8548 1764
rect 9436 1756 9444 1764
rect 9452 1756 9460 1764
rect 652 1736 660 1744
rect 844 1736 852 1744
rect 2540 1736 2548 1744
rect 2700 1736 2708 1744
rect 2892 1736 2900 1744
rect 4044 1736 4052 1744
rect 4540 1736 4548 1744
rect 4748 1736 4756 1744
rect 748 1716 756 1724
rect 1260 1716 1268 1724
rect 2028 1716 2036 1724
rect 2268 1716 2276 1724
rect 2652 1716 2660 1724
rect 1548 1696 1556 1704
rect 2524 1696 2532 1704
rect 3468 1716 3476 1724
rect 3580 1716 3588 1724
rect 3916 1716 3924 1724
rect 5836 1736 5844 1744
rect 6140 1736 6148 1744
rect 7020 1736 7028 1744
rect 7276 1736 7284 1744
rect 7292 1736 7300 1744
rect 7788 1736 7796 1744
rect 5436 1716 5444 1724
rect 7596 1716 7604 1724
rect 7852 1716 7860 1724
rect 7900 1716 7908 1724
rect 3100 1696 3108 1704
rect 3372 1696 3380 1704
rect 3468 1696 3476 1704
rect 5148 1696 5156 1704
rect 5372 1696 5380 1704
rect 6716 1696 6724 1704
rect 7164 1696 7172 1704
rect 7212 1696 7220 1704
rect 7468 1696 7476 1704
rect 7724 1696 7732 1704
rect 8140 1696 8148 1704
rect 9212 1696 9220 1704
rect 9932 1696 9940 1704
rect 1212 1676 1220 1684
rect 2012 1676 2020 1684
rect 428 1656 436 1664
rect 1580 1656 1588 1664
rect 3020 1656 3028 1664
rect 3356 1676 3364 1684
rect 3852 1676 3860 1684
rect 4460 1676 4468 1684
rect 5916 1676 5924 1684
rect 7244 1676 7252 1684
rect 7468 1676 7476 1684
rect 2444 1636 2452 1644
rect 3676 1636 3684 1644
rect 4780 1636 4788 1644
rect 7788 1636 7796 1644
rect 1836 1616 1844 1624
rect 1644 1596 1652 1604
rect 4940 1576 4948 1584
rect 428 1556 436 1564
rect 316 1536 324 1544
rect 620 1536 628 1544
rect 2076 1536 2084 1544
rect 2348 1536 2356 1544
rect 2524 1536 2532 1544
rect 3932 1536 3940 1544
rect 4508 1536 4516 1544
rect 8524 1536 8532 1544
rect 524 1516 532 1524
rect 940 1516 948 1524
rect 1772 1516 1780 1524
rect 3356 1516 3364 1524
rect 4508 1516 4516 1524
rect 4572 1516 4580 1524
rect 5532 1516 5540 1524
rect 5884 1516 5892 1524
rect 6460 1516 6468 1524
rect 7228 1516 7236 1524
rect 7244 1516 7252 1524
rect 7452 1516 7460 1524
rect 7596 1516 7604 1524
rect 8892 1516 8900 1524
rect 9308 1516 9316 1524
rect 9436 1516 9444 1524
rect 92 1496 100 1504
rect 2700 1496 2708 1504
rect 3324 1496 3332 1504
rect 3580 1496 3588 1504
rect 5452 1496 5460 1504
rect 6812 1496 6820 1504
rect 7020 1496 7028 1504
rect 7964 1496 7972 1504
rect 8956 1496 8964 1504
rect 9788 1496 9796 1504
rect 556 1476 564 1484
rect 636 1476 644 1484
rect 876 1476 884 1484
rect 972 1476 980 1484
rect 1436 1476 1444 1484
rect 1660 1476 1668 1484
rect 2556 1476 2564 1484
rect 2908 1476 2916 1484
rect 3020 1476 3028 1484
rect 3532 1476 3540 1484
rect 4140 1476 4148 1484
rect 4316 1476 4324 1484
rect 5340 1476 5348 1484
rect 5724 1476 5732 1484
rect 6044 1476 6052 1484
rect 7884 1476 7892 1484
rect 8236 1476 8244 1484
rect 8972 1476 8980 1484
rect 9004 1476 9012 1484
rect 9404 1476 9412 1484
rect 2764 1456 2772 1464
rect 3148 1456 3156 1464
rect 3964 1456 3972 1464
rect 4476 1456 4484 1464
rect 6700 1456 6708 1464
rect 6924 1456 6932 1464
rect 7020 1456 7028 1464
rect 7292 1456 7300 1464
rect 8012 1456 8020 1464
rect 8044 1456 8052 1464
rect 9308 1456 9316 1464
rect 9324 1456 9332 1464
rect 844 1436 852 1444
rect 2348 1436 2356 1444
rect 3468 1436 3476 1444
rect 8796 1436 8804 1444
rect 8972 1436 8980 1444
rect 684 1416 692 1424
rect 1100 1416 1108 1424
rect 2268 1416 2276 1424
rect 5148 1416 5156 1424
rect 7020 1416 7028 1424
rect 9212 1416 9220 1424
rect 2700 1396 2708 1404
rect 4780 1396 4788 1404
rect 6940 1396 6948 1404
rect 9532 1396 9540 1404
rect 2572 1376 2580 1384
rect 2908 1376 2916 1384
rect 3596 1376 3604 1384
rect 4540 1376 4548 1384
rect 4812 1376 4820 1384
rect 7388 1376 7396 1384
rect 8012 1376 8020 1384
rect 8956 1376 8964 1384
rect 2108 1356 2116 1364
rect 2444 1356 2452 1364
rect 4316 1356 4324 1364
rect 4588 1356 4596 1364
rect 5036 1356 5044 1364
rect 6700 1356 6708 1364
rect 428 1336 436 1344
rect 1196 1336 1204 1344
rect 2012 1336 2020 1344
rect 2876 1336 2884 1344
rect 3772 1336 3780 1344
rect 5356 1336 5364 1344
rect 5804 1336 5812 1344
rect 5900 1336 5908 1344
rect 7404 1336 7412 1344
rect 8476 1336 8484 1344
rect 8812 1336 8820 1344
rect 9132 1336 9140 1344
rect 9244 1336 9252 1344
rect 9484 1336 9492 1344
rect 844 1316 852 1324
rect 2540 1316 2548 1324
rect 5356 1316 5364 1324
rect 5484 1316 5492 1324
rect 6588 1316 6596 1324
rect 6796 1316 6804 1324
rect 7132 1316 7140 1324
rect 7580 1316 7588 1324
rect 7612 1316 7620 1324
rect 7932 1316 7940 1324
rect 9260 1316 9268 1324
rect 92 1296 100 1304
rect 284 1296 292 1304
rect 876 1296 884 1304
rect 1308 1296 1316 1304
rect 1420 1296 1428 1304
rect 2124 1296 2132 1304
rect 2556 1296 2564 1304
rect 2860 1296 2868 1304
rect 4572 1296 4580 1304
rect 4684 1296 4692 1304
rect 5212 1296 5220 1304
rect 5340 1296 5348 1304
rect 6268 1296 6276 1304
rect 7948 1296 7956 1304
rect 9132 1296 9140 1304
rect 5676 1276 5684 1284
rect 5884 1276 5892 1284
rect 6348 1276 6356 1284
rect 6444 1276 6452 1284
rect 8380 1276 8388 1284
rect 9020 1276 9028 1284
rect 988 1256 996 1264
rect 1660 1256 1668 1264
rect 5820 1256 5828 1264
rect 5884 1256 5892 1264
rect 6252 1256 6260 1264
rect 556 1236 564 1244
rect 972 1236 980 1244
rect 3420 1216 3428 1224
rect 76 1196 84 1204
rect 3772 1196 3780 1204
rect 6828 1196 6836 1204
rect 2716 1176 2724 1184
rect 4924 1176 4932 1184
rect 1836 1156 1844 1164
rect 2684 1156 2692 1164
rect 3164 1156 3172 1164
rect 3644 1156 3652 1164
rect 4012 1156 4020 1164
rect 4652 1156 4660 1164
rect 5676 1156 5684 1164
rect 8012 1156 8020 1164
rect 1564 1136 1572 1144
rect 1628 1136 1636 1144
rect 4284 1136 4292 1144
rect 5820 1136 5828 1144
rect 6636 1136 6644 1144
rect 7804 1136 7812 1144
rect 8268 1136 8276 1144
rect 8924 1136 8932 1144
rect 9132 1136 9140 1144
rect 860 1116 868 1124
rect 972 1116 980 1124
rect 3484 1116 3492 1124
rect 3820 1116 3828 1124
rect 4300 1116 4308 1124
rect 4524 1116 4532 1124
rect 4588 1116 4596 1124
rect 5212 1116 5220 1124
rect 5484 1116 5492 1124
rect 5916 1116 5924 1124
rect 5932 1116 5940 1124
rect 6140 1116 6148 1124
rect 6492 1116 6500 1124
rect 7724 1116 7732 1124
rect 8588 1116 8596 1124
rect 236 1096 244 1104
rect 1340 1096 1348 1104
rect 2076 1096 2084 1104
rect 2844 1096 2852 1104
rect 4492 1096 4500 1104
rect 5340 1096 5348 1104
rect 6396 1096 6404 1104
rect 7260 1096 7268 1104
rect 7820 1096 7828 1104
rect 764 1076 772 1084
rect 1644 1076 1652 1084
rect 1772 1076 1780 1084
rect 1996 1076 2004 1084
rect 2428 1076 2436 1084
rect 2892 1076 2900 1084
rect 3548 1076 3556 1084
rect 3836 1076 3844 1084
rect 4796 1076 4804 1084
rect 5356 1076 5364 1084
rect 5404 1076 5412 1084
rect 5852 1076 5860 1084
rect 7900 1076 7908 1084
rect 8476 1076 8484 1084
rect 9468 1076 9476 1084
rect 9820 1076 9828 1084
rect 860 1056 868 1064
rect 3196 1056 3204 1064
rect 3596 1056 3604 1064
rect 3628 1056 3636 1064
rect 3644 1056 3652 1064
rect 5036 1056 5044 1064
rect 7100 1056 7108 1064
rect 7484 1056 7492 1064
rect 8348 1056 8356 1064
rect 8812 1056 8820 1064
rect 9644 1056 9652 1064
rect 9692 1056 9700 1064
rect 204 1036 212 1044
rect 2460 1036 2468 1044
rect 5324 1036 5332 1044
rect 5932 1036 5940 1044
rect 9388 1036 9396 1044
rect 1612 1016 1620 1024
rect 1996 1016 2004 1024
rect 2684 1016 2692 1024
rect 3852 1016 3860 1024
rect 8012 1016 8020 1024
rect 2428 996 2436 1004
rect 3548 996 3556 1004
rect 4812 996 4820 1004
rect 8124 996 8132 1004
rect 1068 976 1076 984
rect 2236 976 2244 984
rect 2252 976 2260 984
rect 3612 976 3620 984
rect 5020 976 5028 984
rect 204 956 212 964
rect 1260 956 1268 964
rect 2060 956 2068 964
rect 2540 956 2548 964
rect 2732 956 2740 964
rect 4268 956 4276 964
rect 5628 956 5636 964
rect 6684 956 6692 964
rect 7116 956 7124 964
rect 8348 956 8356 964
rect 8572 956 8580 964
rect 8908 956 8916 964
rect 9132 956 9140 964
rect 860 936 868 944
rect 1308 936 1316 944
rect 3196 936 3204 944
rect 3372 936 3380 944
rect 3980 936 3988 944
rect 5900 936 5908 944
rect 6124 936 6132 944
rect 6348 936 6356 944
rect 6556 936 6564 944
rect 7132 936 7140 944
rect 7660 936 7668 944
rect 7996 936 8004 944
rect 8284 936 8292 944
rect 9820 936 9828 944
rect 1628 916 1636 924
rect 1660 916 1668 924
rect 2668 916 2676 924
rect 2748 916 2756 924
rect 2764 916 2772 924
rect 3404 916 3412 924
rect 4172 916 4180 924
rect 5788 916 5796 924
rect 8028 916 8036 924
rect 8684 916 8692 924
rect 9228 916 9236 924
rect 428 896 436 904
rect 972 896 980 904
rect 1068 896 1076 904
rect 1548 896 1556 904
rect 3100 896 3108 904
rect 3948 896 3956 904
rect 4188 896 4196 904
rect 6268 896 6276 904
rect 7164 896 7172 904
rect 7932 896 7940 904
rect 7980 896 7988 904
rect 8540 896 8548 904
rect 8860 896 8868 904
rect 8876 896 8884 904
rect 9308 896 9316 904
rect 1724 876 1732 884
rect 4028 876 4036 884
rect 4524 876 4532 884
rect 5228 876 5236 884
rect 5772 876 5780 884
rect 6140 876 6148 884
rect 7260 876 7268 884
rect 9820 876 9828 884
rect 3628 856 3636 864
rect 4956 856 4964 864
rect 5804 856 5812 864
rect 6156 856 6164 864
rect 556 836 564 844
rect 1676 836 1684 844
rect 3100 836 3108 844
rect 4748 836 4756 844
rect 5788 836 5796 844
rect 8460 836 8468 844
rect 5180 816 5188 824
rect 5420 816 5428 824
rect 4716 796 4724 804
rect 5772 796 5780 804
rect 236 776 244 784
rect 5228 776 5236 784
rect 5596 776 5604 784
rect 7596 776 7604 784
rect 6732 756 6740 764
rect 7372 756 7380 764
rect 7388 756 7396 764
rect 7548 756 7556 764
rect 412 736 420 744
rect 2716 736 2724 744
rect 3820 736 3828 744
rect 4652 736 4660 744
rect 5340 736 5348 744
rect 7004 736 7012 744
rect 7100 736 7108 744
rect 9500 736 9508 744
rect 892 716 900 724
rect 1532 716 1540 724
rect 1644 716 1652 724
rect 1948 716 1956 724
rect 6492 716 6500 724
rect 8044 716 8052 724
rect 8092 716 8100 724
rect 8684 716 8692 724
rect 9436 716 9444 724
rect 9532 716 9540 724
rect 10092 716 10100 724
rect 10172 716 10180 724
rect 2028 696 2036 704
rect 5532 696 5540 704
rect 5820 696 5828 704
rect 6684 696 6692 704
rect 7916 696 7924 704
rect 8028 696 8036 704
rect 8044 696 8052 704
rect 444 676 452 684
rect 556 676 564 684
rect 972 676 980 684
rect 1324 676 1332 684
rect 1660 676 1668 684
rect 1740 676 1748 684
rect 2044 676 2052 684
rect 2620 676 2628 684
rect 3084 676 3092 684
rect 3404 676 3412 684
rect 5084 676 5092 684
rect 5212 676 5220 684
rect 5452 676 5460 684
rect 7292 676 7300 684
rect 7356 676 7364 684
rect 7900 676 7908 684
rect 9020 676 9028 684
rect 9884 676 9892 684
rect 92 656 100 664
rect 940 656 948 664
rect 1740 656 1748 664
rect 2396 656 2404 664
rect 2476 656 2484 664
rect 3836 656 3844 664
rect 5100 656 5108 664
rect 5228 656 5236 664
rect 7228 656 7236 664
rect 1868 636 1876 644
rect 2204 636 2212 644
rect 6236 636 6244 644
rect 8252 636 8260 644
rect 8796 636 8804 644
rect 8812 636 8820 644
rect 988 616 996 624
rect 2620 616 2628 624
rect 3308 616 3316 624
rect 5884 616 5892 624
rect 6956 616 6964 624
rect 7740 616 7748 624
rect 92 596 100 604
rect 2396 596 2404 604
rect 2876 596 2884 604
rect 3660 596 3668 604
rect 636 556 644 564
rect 1612 556 1620 564
rect 4092 576 4100 584
rect 4684 576 4692 584
rect 6044 576 6052 584
rect 6396 576 6404 584
rect 7996 576 8004 584
rect 8012 576 8020 584
rect 2956 556 2964 564
rect 3116 556 3124 564
rect 3660 556 3668 564
rect 3948 556 3956 564
rect 5628 556 5636 564
rect 8284 556 8292 564
rect 8476 556 8484 564
rect 860 536 868 544
rect 1068 536 1076 544
rect 1884 536 1892 544
rect 2332 536 2340 544
rect 3132 536 3140 544
rect 3196 536 3204 544
rect 3676 536 3684 544
rect 4220 536 4228 544
rect 4796 536 4804 544
rect 5228 536 5236 544
rect 5596 536 5604 544
rect 6156 536 6164 544
rect 6988 536 6996 544
rect 7292 536 7300 544
rect 7324 536 7332 544
rect 7676 536 7684 544
rect 8252 536 8260 544
rect 8300 536 8308 544
rect 9804 536 9812 544
rect 10092 536 10100 544
rect 300 516 308 524
rect 1004 516 1012 524
rect 1804 516 1812 524
rect 2076 516 2084 524
rect 2412 516 2420 524
rect 2460 516 2468 524
rect 4460 516 4468 524
rect 9388 516 9396 524
rect 10172 516 10180 524
rect 316 496 324 504
rect 1948 496 1956 504
rect 2668 496 2676 504
rect 4300 496 4308 504
rect 5116 496 5124 504
rect 5756 496 5764 504
rect 8460 496 8468 504
rect 8924 496 8932 504
rect 1532 476 1540 484
rect 3308 476 3316 484
rect 6956 476 6964 484
rect 1580 456 1588 464
rect 4700 456 4708 464
rect 5100 456 5108 464
rect 6044 456 6052 464
rect 2204 436 2212 444
rect 7436 416 7444 424
rect 220 396 228 404
rect 3324 396 3332 404
rect 6588 396 6596 404
rect 1532 356 1540 364
rect 3100 356 3108 364
rect 3980 356 3988 364
rect 4956 356 4964 364
rect 5628 356 5636 364
rect 8012 356 8020 364
rect 1948 336 1956 344
rect 5180 336 5188 344
rect 5900 336 5908 344
rect 7788 336 7796 344
rect 8252 336 8260 344
rect 412 316 420 324
rect 860 316 868 324
rect 1068 316 1076 324
rect 2732 316 2740 324
rect 5356 316 5364 324
rect 6236 316 6244 324
rect 7308 316 7316 324
rect 7484 316 7492 324
rect 7676 316 7684 324
rect 8268 316 8276 324
rect 8316 316 8324 324
rect 8924 316 8932 324
rect 9500 316 9508 324
rect 9724 316 9732 324
rect 9756 316 9764 324
rect 652 296 660 304
rect 1724 296 1732 304
rect 1836 296 1844 304
rect 2412 296 2420 304
rect 2748 296 2756 304
rect 3964 296 3972 304
rect 5148 296 5156 304
rect 7740 296 7748 304
rect 7916 296 7924 304
rect 8268 296 8276 304
rect 940 276 948 284
rect 1196 276 1204 284
rect 1260 276 1268 284
rect 2860 276 2868 284
rect 4700 276 4708 284
rect 5036 276 5044 284
rect 5196 276 5204 284
rect 5404 276 5412 284
rect 7292 276 7300 284
rect 8268 276 8276 284
rect 8284 276 8292 284
rect 8924 276 8932 284
rect 9692 276 9700 284
rect 9708 276 9716 284
rect 764 256 772 264
rect 1084 256 1092 264
rect 2476 256 2484 264
rect 140 236 148 244
rect 1420 236 1428 244
rect 1628 236 1636 244
rect 2956 256 2964 264
rect 5196 256 5204 264
rect 8876 256 8884 264
rect 8748 236 8756 244
rect 8956 236 8964 244
rect 1356 216 1364 224
rect 1820 216 1828 224
rect 6012 216 6020 224
rect 6028 216 6036 224
rect 9836 216 9844 224
rect 1580 196 1588 204
rect 2044 196 2052 204
rect 860 176 868 184
rect 3148 176 3156 184
rect 4396 176 4404 184
rect 140 156 148 164
rect 1004 156 1012 164
rect 1356 156 1364 164
rect 1820 156 1828 164
rect 2044 156 2052 164
rect 2956 156 2964 164
rect 3196 156 3204 164
rect 4188 156 4196 164
rect 5116 156 5124 164
rect 8316 176 8324 184
rect 8988 176 8996 184
rect 9148 176 9156 184
rect 9820 176 9828 184
rect 9964 176 9972 184
rect 5964 156 5972 164
rect 8508 156 8516 164
rect 8908 156 8916 164
rect 9756 156 9764 164
rect 3948 136 3956 144
rect 4092 136 4100 144
rect 4700 136 4708 144
rect 6028 136 6036 144
rect 7324 136 7332 144
rect 7356 136 7364 144
rect 7436 136 7444 144
rect 8012 136 8020 144
rect 2732 116 2740 124
rect 4652 116 4660 124
rect 5100 116 5108 124
rect 8108 136 8116 144
rect 9708 136 9716 144
rect 9868 136 9876 144
rect 8508 116 8516 124
rect 9516 116 9524 124
rect 3388 96 3396 104
rect 4172 96 4180 104
rect 4396 96 4404 104
rect 4860 96 4868 104
rect 7676 96 7684 104
rect 9852 96 9860 104
rect 10012 96 10020 104
rect 2700 16 2708 24
rect 4700 16 4708 24
rect 5148 16 5156 24
rect 7356 16 7364 24
<< metal4 >>
rect 77 7384 83 7456
rect 93 7384 99 7456
rect 276 7117 284 7123
rect 77 6724 83 6816
rect 109 6624 115 6656
rect 93 6204 99 6256
rect 109 6224 115 6316
rect 77 4724 83 5736
rect 205 5704 211 7056
rect 301 6604 307 7476
rect 317 7424 323 7516
rect 573 7404 579 7516
rect 909 7424 915 7456
rect 317 6764 323 7336
rect 429 6944 435 7256
rect 637 7084 643 7336
rect 685 6984 691 7096
rect 13 4644 19 4676
rect 77 4024 83 4676
rect 93 3524 99 5216
rect 221 4144 227 6576
rect 301 6304 307 6556
rect 413 6484 419 6496
rect 237 5884 243 6236
rect 413 5764 419 6476
rect 429 6284 435 6896
rect 509 6724 515 6896
rect 317 5364 323 5756
rect 237 4544 243 4796
rect 237 3904 243 4056
rect 212 3877 220 3883
rect 221 3784 227 3856
rect 237 3804 243 3876
rect 77 1204 83 2536
rect 205 2484 211 2996
rect 221 2684 227 3456
rect 221 2624 227 2656
rect 221 2024 227 2136
rect 237 1824 243 3296
rect 93 1304 99 1496
rect 285 1304 291 3856
rect 301 3824 307 3836
rect 317 3504 323 4496
rect 333 3884 339 4096
rect 429 3924 435 5676
rect 445 4224 451 5076
rect 461 4744 467 5216
rect 477 3944 483 6156
rect 509 5684 515 6716
rect 685 6664 691 6676
rect 557 5964 563 6036
rect 637 5944 643 6136
rect 653 5724 659 6096
rect 653 5504 659 5656
rect 525 5144 531 5436
rect 669 4924 675 6496
rect 685 6324 691 6656
rect 749 6604 755 6676
rect 669 4604 675 4896
rect 541 4284 547 4536
rect 669 4504 675 4576
rect 685 4444 691 6316
rect 765 5924 771 7336
rect 781 7044 787 7136
rect 877 6664 883 6936
rect 893 6584 899 7256
rect 973 6904 979 6936
rect 973 6804 979 6896
rect 845 6184 851 6516
rect 861 5884 867 6576
rect 877 6144 883 6456
rect 893 6084 899 6116
rect 973 6084 979 6696
rect 1101 6344 1107 7096
rect 1117 6124 1123 7516
rect 1140 6697 1148 6703
rect 1133 6184 1139 6676
rect 733 5524 739 5716
rect 733 5484 739 5516
rect 893 5244 899 6076
rect 1085 5704 1091 6116
rect 1181 6104 1187 6896
rect 1245 6684 1251 7276
rect 1309 7064 1315 7296
rect 1437 6984 1443 7516
rect 1316 6517 1324 6523
rect 925 5524 931 5616
rect 909 5404 915 5476
rect 909 5164 915 5256
rect 909 4724 915 4856
rect 909 4564 915 4676
rect 333 3424 339 3536
rect 301 1884 307 2936
rect 429 2904 435 3916
rect 445 3384 451 3476
rect 429 2404 435 2536
rect 205 964 211 1036
rect 93 604 99 656
rect 221 404 227 1056
rect 237 1004 243 1096
rect 237 784 243 796
rect 301 524 307 1876
rect 429 1764 435 1816
rect 429 1564 435 1656
rect 317 504 323 1536
rect 429 904 435 1336
rect 413 324 419 736
rect 445 684 451 2936
rect 461 2384 467 3296
rect 477 2504 483 2536
rect 509 2024 515 3576
rect 525 1904 531 4096
rect 541 3584 547 4276
rect 573 3884 579 4316
rect 765 4104 771 4236
rect 637 3864 643 3896
rect 653 3124 659 4076
rect 653 2964 659 3116
rect 669 2944 675 3856
rect 893 3484 899 4436
rect 909 4324 915 4336
rect 909 4204 915 4276
rect 557 2544 563 2556
rect 525 1524 531 1716
rect 621 1544 627 2736
rect 653 2344 659 2356
rect 637 1484 643 1876
rect 653 1744 659 2316
rect 669 2124 675 2896
rect 685 2264 691 3096
rect 701 2584 707 2596
rect 708 2177 716 2183
rect 557 1244 563 1476
rect 557 684 563 836
rect 436 677 444 683
rect 653 304 659 1736
rect 669 1724 675 1756
rect 749 1724 755 2536
rect 765 1884 771 2876
rect 797 2344 803 2476
rect 845 1884 851 2896
rect 909 2484 915 3496
rect 925 2144 931 5496
rect 1101 5283 1107 5776
rect 1117 5744 1123 5756
rect 1085 5277 1107 5283
rect 941 1964 947 5056
rect 973 2904 979 5116
rect 1085 5104 1091 5277
rect 989 3324 995 4276
rect 1005 3844 1011 5056
rect 1101 4904 1107 5256
rect 1021 4264 1027 4276
rect 1021 3844 1027 3876
rect 1101 3564 1107 4076
rect 1117 3704 1123 5736
rect 1213 5564 1219 5716
rect 1149 5364 1155 5436
rect 1341 5364 1347 6836
rect 1357 5744 1363 6716
rect 1357 5484 1363 5696
rect 1229 5124 1235 5216
rect 1085 2744 1091 3116
rect 845 1444 851 1736
rect 685 1104 691 1416
rect 765 664 771 1076
rect 845 1043 851 1316
rect 861 1124 867 1876
rect 957 1764 963 2056
rect 973 1964 979 2176
rect 989 1944 995 2476
rect 1005 2144 1011 2176
rect 989 1804 995 1876
rect 877 1304 883 1476
rect 845 1037 867 1043
rect 861 944 867 1037
rect 765 264 771 656
rect 861 544 867 936
rect 884 717 892 723
rect 941 664 947 1516
rect 973 1244 979 1476
rect 1101 1424 1107 3296
rect 1117 2564 1123 3696
rect 1133 3664 1139 5076
rect 1213 5064 1219 5076
rect 1149 4644 1155 4676
rect 1149 3904 1155 4536
rect 1165 4384 1171 4396
rect 1197 4084 1203 4916
rect 1245 4784 1251 5336
rect 1213 4097 1228 4103
rect 1213 4084 1219 4097
rect 1133 3344 1139 3456
rect 1133 3264 1139 3336
rect 1149 3304 1155 3896
rect 1197 3884 1203 4076
rect 1213 3064 1219 3116
rect 1181 2844 1187 3056
rect 1133 2604 1139 2676
rect 1133 1804 1139 2576
rect 1229 2504 1235 3936
rect 1341 3504 1347 3676
rect 1245 3364 1251 3376
rect 1245 3104 1251 3256
rect 1245 2544 1251 3076
rect 1261 2684 1267 2756
rect 1357 2624 1363 3736
rect 1405 3504 1411 5296
rect 1421 4504 1427 6336
rect 1444 6257 1452 6263
rect 1469 6204 1475 6976
rect 1549 6864 1555 7276
rect 1565 7104 1571 7296
rect 1549 6644 1555 6856
rect 1597 6124 1603 6236
rect 1469 5504 1475 5656
rect 1533 5044 1539 6056
rect 1549 4904 1555 5236
rect 1549 4744 1555 4896
rect 1549 4484 1555 4716
rect 1421 2924 1427 4296
rect 1549 3904 1555 4436
rect 1549 2804 1555 2856
rect 1229 2484 1235 2496
rect 1197 1344 1203 1876
rect 1261 1724 1267 2136
rect 1213 1323 1219 1676
rect 1197 1317 1219 1323
rect 989 1264 995 1276
rect 973 904 979 1116
rect 1069 984 1075 1276
rect 1069 904 1075 976
rect 973 684 979 896
rect 141 164 147 236
rect 861 184 867 316
rect 941 284 947 656
rect 1005 164 1011 516
rect 1069 324 1075 536
rect 1085 264 1091 676
rect 1197 284 1203 1317
rect 1261 964 1267 1716
rect 1277 1044 1283 2496
rect 1293 2264 1299 2536
rect 1565 2284 1571 6116
rect 1613 6104 1619 6256
rect 1629 6144 1635 7116
rect 1661 6704 1667 7196
rect 1581 5304 1587 5936
rect 1629 5764 1635 6136
rect 1645 6104 1651 6636
rect 1661 6544 1667 6696
rect 1597 5484 1603 5516
rect 1581 5144 1587 5296
rect 1581 4964 1587 5116
rect 1581 4384 1587 4916
rect 1581 4124 1587 4236
rect 1597 3884 1603 4536
rect 1613 4064 1619 4456
rect 1597 3704 1603 3756
rect 1629 3524 1635 5756
rect 1645 4324 1651 5916
rect 1693 5784 1699 7476
rect 1869 7124 1875 7336
rect 1789 6544 1795 7036
rect 1853 6644 1859 6936
rect 1677 5664 1683 5776
rect 1700 4537 1708 4543
rect 1325 2264 1331 2276
rect 1549 1704 1555 2096
rect 1261 284 1267 956
rect 1309 944 1315 1296
rect 1348 1097 1356 1103
rect 1325 684 1331 1036
rect 1421 244 1427 1296
rect 1533 724 1539 1176
rect 1549 904 1555 1696
rect 1581 1664 1587 3316
rect 1597 3204 1603 3336
rect 1613 3183 1619 3276
rect 1597 3177 1619 3183
rect 1597 2884 1603 3177
rect 1629 2964 1635 3516
rect 1613 2164 1619 2236
rect 1613 1764 1619 2156
rect 1629 1924 1635 2956
rect 1645 2684 1651 4316
rect 1693 4264 1699 4456
rect 1741 4304 1747 5776
rect 1757 5284 1763 6136
rect 1741 3744 1747 3876
rect 1645 2304 1651 2676
rect 1661 2624 1667 2716
rect 1629 1144 1635 1916
rect 1645 1604 1651 2296
rect 1741 2264 1747 3736
rect 1757 2304 1763 3656
rect 1773 3444 1779 4896
rect 1789 4724 1795 5416
rect 1789 3844 1795 3856
rect 1805 3764 1811 5896
rect 1789 3464 1795 3476
rect 1789 2544 1795 2636
rect 1805 2523 1811 3756
rect 1821 2644 1827 3456
rect 1837 2884 1843 4916
rect 1869 4664 1875 7116
rect 1885 6764 1891 7016
rect 1901 6244 1907 6496
rect 1949 5924 1955 6576
rect 1997 6104 2003 6516
rect 2013 5904 2019 6016
rect 2029 5364 2035 7456
rect 2237 7124 2243 7216
rect 2109 7044 2115 7076
rect 2253 7004 2259 7076
rect 2077 6104 2083 6896
rect 2093 6504 2099 6956
rect 2349 6924 2355 7076
rect 2445 7064 2451 7316
rect 2461 7084 2467 7176
rect 2109 6504 2115 6596
rect 2269 6584 2275 6696
rect 2285 6684 2291 6916
rect 2045 5404 2051 5496
rect 1885 3944 1891 4736
rect 1917 4684 1923 4896
rect 1908 4657 1916 4663
rect 2061 4584 2067 5516
rect 2109 5404 2115 5696
rect 2157 5524 2163 6156
rect 2205 6044 2211 6063
rect 2013 3804 2019 4136
rect 2013 3444 2019 3756
rect 1828 2537 1836 2543
rect 1789 2517 1811 2523
rect 1757 2264 1763 2296
rect 1565 1104 1571 1136
rect 1613 564 1619 1016
rect 1629 924 1635 1136
rect 1645 1084 1651 1596
rect 1661 1484 1667 2156
rect 1773 1524 1779 2296
rect 1789 1924 1795 2517
rect 1805 2344 1811 2496
rect 1885 2324 1891 3296
rect 2013 2904 2019 3376
rect 1997 2664 2003 2856
rect 2004 2537 2012 2543
rect 1901 2324 1907 2336
rect 1812 2197 1820 2203
rect 1837 1864 1843 1876
rect 1645 724 1651 1076
rect 1661 943 1667 1256
rect 1661 937 1683 943
rect 1661 684 1667 916
rect 1677 844 1683 937
rect 1533 364 1539 476
rect 1357 164 1363 216
rect 1581 204 1587 456
rect 1725 304 1731 876
rect 1741 684 1747 1496
rect 1837 1164 1843 1616
rect 1773 1084 1779 1096
rect 1869 724 1875 2276
rect 1741 664 1747 676
rect 1869 644 1875 716
rect 1885 544 1891 2316
rect 2029 2304 2035 3516
rect 2109 3344 2115 5336
rect 2157 5104 2163 5516
rect 2221 5444 2227 6576
rect 2349 6524 2355 6916
rect 2237 6304 2243 6416
rect 2365 6243 2371 6736
rect 2413 6564 2419 6696
rect 2397 6364 2403 6536
rect 2349 6237 2371 6243
rect 2333 6104 2339 6216
rect 2269 5804 2275 5896
rect 2221 5144 2227 5376
rect 2276 5277 2284 5283
rect 2141 4244 2147 4816
rect 2253 4624 2259 4676
rect 2253 4324 2259 4616
rect 2269 4584 2275 4636
rect 2221 3444 2227 3476
rect 2237 3444 2243 3656
rect 2077 3064 2083 3076
rect 2093 2284 2099 2316
rect 2109 2264 2115 3336
rect 2157 3044 2163 3356
rect 2125 2664 2131 2676
rect 2173 2304 2179 2336
rect 2189 2284 2195 2676
rect 2221 2544 2227 3056
rect 2237 2704 2243 2816
rect 2253 2684 2259 4276
rect 1901 1804 1907 1936
rect 1997 1884 2003 2096
rect 1997 1824 2003 1876
rect 2013 1344 2019 1676
rect 1997 1024 2003 1076
rect 1805 524 1811 536
rect 1949 504 1955 716
rect 2029 704 2035 1716
rect 2061 964 2067 2096
rect 2084 1537 2092 1543
rect 2109 1364 2115 2076
rect 2221 1944 2227 1956
rect 2125 1304 2131 1936
rect 2045 664 2051 676
rect 2077 524 2083 1096
rect 2237 984 2243 2296
rect 2253 1924 2259 2516
rect 2269 2304 2275 4456
rect 2285 3944 2291 4616
rect 2301 3903 2307 6056
rect 2349 5824 2355 6237
rect 2429 5944 2435 6896
rect 2477 6264 2483 6336
rect 2493 6304 2499 7296
rect 2589 7024 2595 7516
rect 2733 7144 2739 7516
rect 2621 6784 2627 7116
rect 2637 6784 2643 6936
rect 2461 6104 2467 6136
rect 2333 5704 2339 5816
rect 2477 5764 2483 6256
rect 2493 6144 2499 6296
rect 2333 5244 2339 5696
rect 2285 3897 2307 3903
rect 2285 3284 2291 3897
rect 2333 3724 2339 4316
rect 2333 2784 2339 2916
rect 2349 2544 2355 4836
rect 2365 4684 2371 5756
rect 2445 4964 2451 5456
rect 2365 4644 2371 4676
rect 2445 4544 2451 4956
rect 2413 3764 2419 4536
rect 2461 4144 2467 4876
rect 2381 3164 2387 3276
rect 2413 3084 2419 3756
rect 2461 3504 2467 3716
rect 2477 3524 2483 5236
rect 2493 4484 2499 6076
rect 2509 5944 2515 6556
rect 2637 6504 2643 6556
rect 2653 6504 2659 6776
rect 2669 6624 2675 6736
rect 2637 6344 2643 6456
rect 2525 5944 2531 6116
rect 2509 5504 2515 5636
rect 2525 5484 2531 5496
rect 2525 5384 2531 5396
rect 2493 4124 2499 4136
rect 2525 3804 2531 4636
rect 2525 3524 2531 3736
rect 2484 3517 2492 3523
rect 2381 2544 2387 2556
rect 2461 2324 2467 3116
rect 2477 2084 2483 2676
rect 2493 2504 2499 3496
rect 2525 3144 2531 3516
rect 2525 2304 2531 3136
rect 2541 3064 2547 5276
rect 2557 4744 2563 6276
rect 2637 6184 2643 6336
rect 2685 6204 2691 6256
rect 2573 5064 2579 5616
rect 2669 5084 2675 5636
rect 2701 5444 2707 6656
rect 2749 6544 2755 7276
rect 2765 6924 2771 7336
rect 2788 7117 2796 7123
rect 2797 6304 2803 6676
rect 2829 6644 2835 6676
rect 2717 5524 2723 5916
rect 2813 5843 2819 6536
rect 2845 6144 2851 6476
rect 2861 6244 2867 6576
rect 2909 6344 2915 7116
rect 3085 7084 3091 7336
rect 3181 7324 3187 7396
rect 3229 7284 3235 7336
rect 3021 7004 3027 7076
rect 3117 7044 3123 7256
rect 2925 6764 2931 6976
rect 2948 6917 2956 6923
rect 2973 6664 2979 6936
rect 2909 6204 2915 6316
rect 2909 5964 2915 6196
rect 2973 6104 2979 6656
rect 3101 6544 3107 6596
rect 3117 6264 3123 6356
rect 3101 6084 3107 6103
rect 2797 5837 2819 5843
rect 2781 5784 2787 5803
rect 2749 5544 2755 5636
rect 2573 4924 2579 4956
rect 2589 4924 2595 5036
rect 2669 4964 2675 4976
rect 2701 4724 2707 5416
rect 2445 1884 2451 1916
rect 2269 1484 2275 1716
rect 2269 1424 2275 1476
rect 2253 984 2259 996
rect 1949 344 1955 496
rect 2205 444 2211 636
rect 2333 544 2339 1816
rect 2461 1764 2467 1816
rect 2349 1444 2355 1536
rect 2445 1364 2451 1636
rect 2429 1004 2435 1076
rect 2397 604 2403 656
rect 2461 524 2467 1036
rect 2477 664 2483 2056
rect 2525 1704 2531 2296
rect 2541 1744 2547 3056
rect 2557 3024 2563 4716
rect 2573 2164 2579 4696
rect 2669 4444 2675 4656
rect 2589 3904 2595 4236
rect 2589 3604 2595 3736
rect 2637 3704 2643 4356
rect 2685 4204 2691 4296
rect 2701 4204 2707 4256
rect 2717 3904 2723 5436
rect 2740 5337 2748 5343
rect 2797 5164 2803 5837
rect 2829 5344 2835 5556
rect 2797 4904 2803 4916
rect 2797 4484 2803 4896
rect 2813 4684 2819 5256
rect 2941 4984 2947 5116
rect 2772 4477 2780 4483
rect 2797 4344 2803 4456
rect 2797 4124 2803 4316
rect 2909 4164 2915 4536
rect 2653 2944 2659 2976
rect 2532 1537 2540 1543
rect 2541 964 2547 1316
rect 2557 1304 2563 1476
rect 2573 1384 2579 2156
rect 2653 1944 2659 2216
rect 2669 1904 2675 2956
rect 2653 1724 2659 1856
rect 2669 924 2675 1896
rect 2685 1164 2691 3736
rect 2708 3477 2716 3483
rect 2701 1744 2707 3096
rect 2717 2764 2723 3036
rect 2733 3004 2739 4076
rect 2877 3924 2883 4076
rect 2909 3944 2915 4156
rect 2733 2164 2739 2996
rect 2749 2564 2755 3076
rect 2829 3004 2835 3356
rect 2845 3284 2851 3356
rect 2877 3104 2883 3916
rect 2868 3097 2876 3103
rect 2701 1504 2707 1736
rect 2685 1024 2691 1156
rect 2413 304 2419 516
rect 1837 264 1843 296
rect 2477 264 2483 656
rect 2621 624 2627 676
rect 2669 504 2675 916
rect 1629 244 1635 256
rect 1821 164 1827 216
rect 2045 164 2051 196
rect 2701 24 2707 1396
rect 2717 744 2723 1176
rect 2733 964 2739 2076
rect 2733 324 2739 956
rect 2749 924 2755 2556
rect 2797 2284 2803 2536
rect 2845 2504 2851 2996
rect 2861 2904 2867 3096
rect 2925 2784 2931 3916
rect 2916 2717 2924 2723
rect 2861 2344 2867 2716
rect 2861 2324 2867 2336
rect 2781 2244 2787 2276
rect 2829 1924 2835 1936
rect 2941 1744 2947 4936
rect 2989 4524 2995 4716
rect 2957 3124 2963 4496
rect 3021 4084 3027 5876
rect 3037 5724 3043 5756
rect 3053 5724 3059 5756
rect 3037 4904 3043 5716
rect 3037 4884 3043 4896
rect 3101 4564 3107 5056
rect 3149 4504 3155 6396
rect 3181 6344 3187 6716
rect 3245 6484 3251 7136
rect 3325 7104 3331 7256
rect 3325 7064 3331 7096
rect 3341 7084 3347 7316
rect 3373 7104 3379 7336
rect 3165 5724 3171 5796
rect 3181 5764 3187 6336
rect 3245 6324 3251 6336
rect 3261 5843 3267 6536
rect 3245 5837 3267 5843
rect 3172 5537 3180 5543
rect 3245 5504 3251 5837
rect 3309 5544 3315 6896
rect 3325 5884 3331 6096
rect 3309 5444 3315 5536
rect 3149 4284 3155 4496
rect 3165 4444 3171 4463
rect 2973 3124 2979 3476
rect 2957 2904 2963 3116
rect 3053 2544 3059 3196
rect 3085 2284 3091 2976
rect 3101 2904 3107 3296
rect 3101 2444 3107 2736
rect 3133 2664 3139 3876
rect 3165 3744 3171 3856
rect 3149 3464 3155 3476
rect 3085 2264 3091 2276
rect 3012 2157 3020 2163
rect 3005 1824 3011 2076
rect 3149 1944 3155 3436
rect 3165 3024 3171 3716
rect 3181 3704 3187 4116
rect 3181 3364 3187 3416
rect 3181 2644 3187 3296
rect 3197 2944 3203 3896
rect 3213 3044 3219 5276
rect 3261 5244 3267 5256
rect 3261 4964 3267 5016
rect 3373 4724 3379 7096
rect 3405 6544 3411 6916
rect 3485 6904 3491 7496
rect 4132 7477 4140 7483
rect 3501 6924 3507 7436
rect 3620 7317 3628 7323
rect 3533 7064 3539 7256
rect 3485 6644 3491 6716
rect 3549 6584 3555 6856
rect 3405 5384 3411 5416
rect 3421 5404 3427 5556
rect 3421 5324 3427 5356
rect 3421 5204 3427 5296
rect 3229 4244 3235 4256
rect 3245 2964 3251 3276
rect 3172 2317 3180 2323
rect 2765 924 2771 1456
rect 2861 1304 2867 1376
rect 2733 124 2739 316
rect 2749 304 2755 916
rect 2861 284 2867 1296
rect 2877 604 2883 1336
rect 2893 1084 2899 1736
rect 3021 1484 3027 1656
rect 2909 1384 2915 1476
rect 3101 904 3107 1696
rect 3076 677 3084 683
rect 2964 557 2972 563
rect 3101 364 3107 836
rect 3133 544 3139 936
rect 2957 164 2963 256
rect 3149 184 3155 1456
rect 3165 1164 3171 1896
rect 3197 1064 3203 2936
rect 3213 2284 3219 2716
rect 3341 2304 3347 4716
rect 3373 4684 3379 4696
rect 3357 3504 3363 4476
rect 3373 4124 3379 4536
rect 3389 4484 3395 5116
rect 3373 3924 3379 4116
rect 3389 3524 3395 4296
rect 3405 4124 3411 4236
rect 3405 4064 3411 4096
rect 3412 3737 3420 3743
rect 3437 3724 3443 5796
rect 3533 5184 3539 6316
rect 3565 5704 3571 6136
rect 3581 5904 3587 6016
rect 3597 5944 3603 6716
rect 3629 6344 3635 6576
rect 3597 5804 3603 5876
rect 3581 5484 3587 5696
rect 3629 5324 3635 5416
rect 3693 5404 3699 7056
rect 3709 6664 3715 7116
rect 3741 6084 3747 7376
rect 4093 7324 4099 7356
rect 4221 7284 4227 7516
rect 4269 7484 4275 7536
rect 3757 6284 3763 7116
rect 3869 7104 3875 7276
rect 3789 6584 3795 6856
rect 3981 6744 3987 7276
rect 4100 7057 4108 7063
rect 4221 6904 4227 7276
rect 4397 7264 4403 7476
rect 3837 6704 3843 6716
rect 3805 5904 3811 6476
rect 3789 5604 3795 5876
rect 3645 5204 3651 5336
rect 3805 5144 3811 5896
rect 3837 5784 3843 6696
rect 3965 6244 3971 6536
rect 3981 6144 3987 6456
rect 3965 5864 3971 6136
rect 3821 5484 3827 5496
rect 3565 4344 3571 4696
rect 3581 4544 3587 4676
rect 3581 3643 3587 4536
rect 3597 4324 3603 4696
rect 3613 4644 3619 5076
rect 3565 3637 3587 3643
rect 3357 3324 3363 3476
rect 3357 3084 3363 3316
rect 3357 2664 3363 2856
rect 3357 2264 3363 2636
rect 3309 1684 3315 2256
rect 3373 1704 3379 3496
rect 3389 3484 3395 3496
rect 3357 1524 3363 1676
rect 3197 944 3203 1056
rect 3188 537 3196 543
rect 3309 484 3315 616
rect 3197 164 3203 476
rect 3325 404 3331 1496
rect 3389 664 3395 2656
rect 3405 2244 3411 3356
rect 3421 2244 3427 2456
rect 3501 2344 3507 2696
rect 3549 2564 3555 3076
rect 3565 2944 3571 3637
rect 3501 2324 3507 2336
rect 3405 1964 3411 2016
rect 3405 924 3411 1756
rect 3469 1724 3475 2256
rect 3421 1224 3427 1676
rect 3469 1444 3475 1696
rect 3421 1104 3427 1216
rect 3485 1124 3491 2276
rect 3533 1484 3539 2136
rect 3549 1084 3555 2556
rect 3565 2144 3571 2936
rect 3581 2904 3587 3476
rect 3581 2684 3587 2896
rect 3597 2704 3603 4316
rect 3757 4304 3763 4316
rect 3821 4304 3827 4936
rect 3853 4904 3859 5016
rect 3837 4484 3843 4716
rect 3853 4584 3859 4856
rect 3869 4484 3875 5456
rect 3885 5244 3891 5716
rect 3917 5564 3923 5736
rect 3933 4524 3939 5496
rect 3949 4984 3955 5496
rect 3997 5444 4003 6896
rect 4013 6264 4019 6276
rect 4013 6184 4019 6236
rect 4013 6104 4019 6176
rect 4029 5904 4035 6256
rect 4045 5924 4051 6676
rect 4205 6384 4211 6836
rect 4061 6284 4067 6336
rect 4045 5724 4051 5916
rect 3965 4744 3971 5436
rect 4045 5304 4051 5376
rect 4061 5024 4067 6216
rect 4221 6184 4227 6876
rect 4269 6764 4275 6836
rect 4253 6604 4259 6676
rect 4333 6544 4339 6936
rect 4413 6644 4419 6736
rect 3629 3864 3635 4136
rect 3620 3457 3628 3463
rect 3597 2684 3603 2696
rect 3581 2604 3587 2636
rect 3581 2244 3587 2256
rect 3581 1724 3587 2216
rect 3581 1504 3587 1716
rect 3549 1004 3555 1076
rect 3405 684 3411 916
rect 3581 684 3587 1496
rect 3597 1384 3603 2676
rect 3613 2324 3619 3116
rect 3613 984 3619 2316
rect 3629 2284 3635 2496
rect 3645 1164 3651 3816
rect 3741 3284 3747 3616
rect 3773 3124 3779 3696
rect 3805 3524 3811 3676
rect 3869 3464 3875 4476
rect 4013 4344 4019 4896
rect 4077 4504 4083 5716
rect 4093 4904 4099 5236
rect 4109 5104 4115 6036
rect 4237 5884 4243 6256
rect 4205 5344 4211 5576
rect 4125 5204 4131 5336
rect 4221 5264 4227 5736
rect 4164 4897 4172 4903
rect 4093 4884 4099 4896
rect 3917 3884 3923 3916
rect 3853 3364 3859 3456
rect 3748 3077 3756 3083
rect 3741 2364 3747 2876
rect 3789 2724 3795 2916
rect 3821 2904 3827 3276
rect 3869 3144 3875 3456
rect 3917 3264 3923 3876
rect 3965 3524 3971 3776
rect 3997 3504 4003 4276
rect 4045 3784 4051 4096
rect 4061 3904 4067 3936
rect 4013 3464 4019 3776
rect 4013 3444 4019 3456
rect 3949 2924 3955 3376
rect 3821 2324 3827 2576
rect 3949 2344 3955 2916
rect 3821 2144 3827 2316
rect 4029 2164 4035 2716
rect 4045 2144 4051 3756
rect 4061 3284 4067 3896
rect 4077 3704 4083 4256
rect 4109 3744 4115 4256
rect 4061 3124 4067 3276
rect 4157 3064 4163 4056
rect 4173 3344 4179 4556
rect 4237 4504 4243 5336
rect 4253 5124 4259 5916
rect 4333 5524 4339 6496
rect 4349 6304 4355 6636
rect 4445 6504 4451 7316
rect 4285 4964 4291 5496
rect 4189 4104 4195 4496
rect 4333 4324 4339 5516
rect 4349 4544 4355 6296
rect 4365 5504 4371 5516
rect 4381 3924 4387 5536
rect 4397 5004 4403 5056
rect 4461 4904 4467 7296
rect 4541 7124 4547 7456
rect 4477 6104 4483 7076
rect 4477 5684 4483 6096
rect 4493 5564 4499 6676
rect 4557 6504 4563 6956
rect 4605 6924 4611 7256
rect 4525 6444 4531 6496
rect 4493 5524 4499 5556
rect 4509 5044 4515 5756
rect 4477 4724 4483 5036
rect 4468 4657 4476 4663
rect 4301 3804 4307 3876
rect 4244 3437 4252 3443
rect 4212 3137 4220 3143
rect 4196 3077 4204 3083
rect 4237 2964 4243 3236
rect 4221 2884 4227 2896
rect 4237 2704 4243 2956
rect 4269 2844 4275 3436
rect 4285 3084 4291 3456
rect 4301 2784 4307 3716
rect 4525 3704 4531 6436
rect 4621 6144 4627 6336
rect 4653 6284 4659 7336
rect 4813 7104 4819 7516
rect 4845 7304 4851 7336
rect 4548 6097 4556 6103
rect 4685 5804 4691 5856
rect 4701 5764 4707 6836
rect 4557 5364 4563 5696
rect 4317 3404 4323 3696
rect 4317 3324 4323 3336
rect 4317 2784 4323 3296
rect 4477 3244 4483 3476
rect 4349 3044 4355 3076
rect 4349 2983 4355 3036
rect 4349 2977 4371 2983
rect 4340 2897 4348 2903
rect 4109 2664 4115 2696
rect 4061 2344 4067 2436
rect 4077 2284 4083 2536
rect 3837 1804 3843 1956
rect 3917 1864 3923 1876
rect 3917 1724 3923 1856
rect 3629 864 3635 1056
rect 3389 104 3395 656
rect 3661 564 3667 596
rect 3677 544 3683 1636
rect 3773 1204 3779 1336
rect 3821 744 3827 1116
rect 3837 664 3843 1076
rect 3853 1024 3859 1676
rect 3933 1544 3939 2056
rect 3949 564 3955 896
rect 3949 144 3955 556
rect 3965 304 3971 1456
rect 4013 1144 4019 1156
rect 3981 364 3987 936
rect 4029 884 4035 2076
rect 4045 1744 4051 2136
rect 4077 1964 4083 2116
rect 4141 1504 4147 1856
rect 4141 1484 4147 1496
rect 4269 964 4275 2736
rect 4285 2504 4291 2696
rect 4308 2677 4316 2683
rect 4301 2564 4307 2596
rect 4285 1924 4291 2496
rect 4365 2284 4371 2977
rect 4477 2744 4483 3036
rect 4301 2124 4307 2136
rect 4333 1844 4339 2136
rect 4349 1844 4355 1876
rect 4285 1144 4291 1816
rect 4301 1144 4307 1836
rect 4461 1684 4467 2576
rect 4477 1464 4483 2656
rect 4493 1924 4499 3116
rect 4509 2124 4515 3456
rect 4525 3124 4531 3336
rect 4541 3044 4547 4956
rect 4557 3484 4563 5356
rect 4589 5104 4595 5516
rect 4605 4944 4611 5496
rect 4573 3564 4579 4096
rect 4557 3104 4563 3296
rect 4573 3084 4579 3136
rect 4589 3084 4595 4936
rect 4621 4884 4627 5696
rect 4669 5504 4675 5676
rect 4717 5564 4723 6556
rect 4717 5504 4723 5536
rect 4733 4564 4739 7036
rect 4756 6717 4764 6723
rect 4829 6544 4835 6936
rect 4845 6904 4851 7296
rect 4973 6924 4979 7276
rect 4989 7124 4995 7256
rect 4845 6304 4851 6896
rect 4877 6604 4883 6896
rect 4765 6104 4771 6136
rect 4653 4544 4659 4556
rect 4653 3904 4659 4136
rect 4605 3444 4611 3516
rect 4557 2144 4563 3056
rect 4605 2704 4611 3316
rect 4621 3184 4627 3336
rect 4605 2164 4611 2676
rect 4621 2304 4627 3076
rect 4701 2984 4707 3756
rect 4653 2744 4659 2756
rect 4717 2724 4723 4316
rect 4733 3764 4739 4536
rect 4749 4104 4755 4496
rect 4781 4244 4787 5756
rect 4797 5684 4803 6296
rect 4813 5924 4819 6176
rect 4925 6084 4931 6516
rect 4941 6304 4947 6836
rect 5021 6344 5027 7536
rect 5181 7344 5187 7616
rect 6093 7524 6099 7556
rect 5181 7304 5187 7336
rect 5213 7144 5219 7356
rect 5053 6764 5059 6916
rect 5085 6744 5091 6936
rect 5085 6684 5091 6716
rect 5213 6644 5219 7116
rect 5229 7084 5235 7156
rect 5229 6684 5235 7076
rect 5181 6624 5187 6636
rect 5021 6304 5027 6316
rect 4813 5783 4819 5916
rect 4813 5777 4835 5783
rect 4797 4844 4803 5296
rect 4813 5284 4819 5736
rect 4829 5564 4835 5777
rect 4925 5724 4931 6076
rect 4925 5624 4931 5643
rect 4925 5344 4931 5376
rect 4941 5344 4947 6296
rect 4957 6264 4963 6276
rect 5005 5544 5011 5896
rect 5021 5304 5027 6296
rect 5101 5924 5107 6156
rect 5181 5524 5187 6616
rect 5293 6324 5299 6536
rect 5293 6304 5299 6316
rect 5229 5924 5235 6056
rect 5261 5984 5267 6116
rect 5229 5504 5235 5736
rect 4749 3084 4755 3696
rect 4781 3484 4787 3496
rect 4797 3484 4803 4476
rect 4692 2357 4700 2363
rect 4317 1364 4323 1376
rect 4093 144 4099 576
rect 4173 104 4179 916
rect 4189 164 4195 896
rect 4221 544 4227 556
rect 4301 504 4307 1116
rect 4493 1104 4499 1916
rect 4509 1544 4515 2116
rect 4701 1804 4707 1856
rect 4548 1737 4556 1743
rect 4509 1524 4515 1536
rect 4541 1384 4547 1736
rect 4573 1304 4579 1516
rect 4589 1124 4595 1356
rect 4525 884 4531 1116
rect 4653 744 4659 1156
rect 4685 1084 4691 1296
rect 4685 584 4691 1076
rect 4717 804 4723 2716
rect 4797 2643 4803 3476
rect 4813 3044 4819 5096
rect 4948 4937 4956 4943
rect 4845 3884 4851 4316
rect 4948 4137 4956 4143
rect 4797 2637 4819 2643
rect 4749 2564 4755 2616
rect 4749 844 4755 1736
rect 4781 1644 4787 2276
rect 4813 1884 4819 2637
rect 4829 1944 4835 2236
rect 4845 1924 4851 3036
rect 4909 2964 4915 3036
rect 4941 3024 4947 3056
rect 4973 3044 4979 4896
rect 5021 4504 5027 5296
rect 5053 4264 5059 4736
rect 5197 4704 5203 4716
rect 5165 4604 5171 4656
rect 5085 4324 5091 4476
rect 5181 4344 5187 4696
rect 5156 4177 5164 4183
rect 5069 3944 5075 4136
rect 4989 3364 4995 3436
rect 4877 2664 4883 2756
rect 4909 2284 4915 2876
rect 4845 1864 4851 1916
rect 4781 1404 4787 1616
rect 4797 544 4803 1076
rect 4813 1004 4819 1376
rect 4925 1184 4931 2296
rect 4941 2264 4947 2896
rect 4964 2697 4972 2703
rect 4957 2304 4963 2696
rect 4989 2544 4995 3116
rect 5005 2724 5011 3936
rect 5037 3044 5043 3176
rect 5005 2544 5011 2716
rect 5085 2504 5091 3336
rect 5117 3104 5123 3136
rect 5133 2804 5139 3936
rect 5149 3524 5155 3776
rect 5181 3764 5187 4336
rect 5181 3304 5187 3356
rect 4941 1584 4947 2056
rect 4989 1924 4995 2496
rect 5037 1364 5043 2496
rect 5133 2364 5139 2556
rect 5149 2324 5155 3096
rect 5181 3084 5187 3296
rect 5181 2744 5187 2876
rect 5149 1704 5155 2316
rect 5197 1764 5203 2796
rect 5229 2264 5235 5336
rect 5245 3124 5251 5296
rect 5261 5264 5267 5976
rect 5261 3444 5267 4816
rect 5277 4644 5283 6176
rect 5341 5724 5347 7356
rect 5389 7064 5395 7296
rect 5389 6264 5395 7056
rect 5405 6944 5411 7516
rect 5373 6204 5379 6256
rect 5364 5877 5372 5883
rect 5389 5864 5395 5916
rect 5405 5884 5411 6936
rect 5469 6724 5475 7076
rect 5565 6684 5571 7336
rect 5421 5944 5427 6536
rect 5517 5924 5523 6336
rect 5357 5464 5363 5696
rect 5309 4504 5315 4636
rect 5341 3984 5347 5256
rect 5405 5084 5411 5876
rect 5485 5744 5491 5856
rect 5517 5744 5523 5916
rect 5581 5864 5587 7296
rect 5773 7124 5779 7296
rect 5597 6704 5603 6816
rect 5757 6664 5763 6756
rect 5773 6604 5779 7116
rect 5789 6644 5795 7056
rect 5837 6664 5843 7496
rect 5773 6584 5779 6596
rect 5597 6284 5603 6336
rect 5597 5884 5603 6276
rect 5684 5757 5692 5763
rect 5357 4044 5363 4536
rect 5332 3477 5340 3483
rect 5325 2944 5331 3456
rect 5357 3124 5363 4036
rect 5389 3344 5395 4136
rect 5405 3304 5411 5076
rect 5421 3744 5427 5536
rect 5453 5484 5459 5716
rect 5453 5064 5459 5476
rect 5485 5084 5491 5736
rect 5581 5444 5587 5736
rect 5709 5703 5715 6556
rect 5764 6497 5772 6503
rect 5709 5697 5731 5703
rect 5709 5664 5715 5676
rect 5389 3084 5395 3116
rect 5437 3084 5443 4316
rect 5453 4124 5459 5056
rect 5476 4717 5484 4723
rect 5501 3364 5507 5136
rect 5533 3944 5539 4676
rect 5485 3124 5491 3136
rect 5325 1884 5331 2936
rect 5348 2297 5356 2303
rect 5149 1424 5155 1696
rect 5037 1064 5043 1356
rect 5021 904 5027 976
rect 4397 104 4403 176
rect 4653 124 4659 436
rect 4701 284 4707 456
rect 4701 144 4707 276
rect 4701 24 4707 136
rect 4861 104 4867 556
rect 4957 364 4963 856
rect 5037 284 5043 1056
rect 5085 444 5091 676
rect 5101 464 5107 656
rect 5101 124 5107 356
rect 5117 164 5123 496
rect 5181 364 5187 816
rect 5181 344 5187 356
rect 5149 24 5155 296
rect 5197 284 5203 1756
rect 5213 1124 5219 1296
rect 5213 684 5219 1116
rect 5325 1044 5331 1876
rect 5373 1704 5379 3056
rect 5389 2444 5395 2636
rect 5517 2484 5523 3916
rect 5533 3844 5539 3856
rect 5549 3744 5555 3936
rect 5565 3844 5571 4956
rect 5581 4704 5587 5336
rect 5597 4324 5603 4336
rect 5645 3884 5651 4336
rect 5709 4104 5715 5656
rect 5725 5304 5731 5697
rect 5741 5484 5747 6116
rect 5789 5904 5795 6636
rect 5837 5484 5843 6316
rect 5725 4684 5731 5296
rect 5741 4884 5747 4956
rect 5853 4924 5859 6696
rect 5869 6524 5875 7316
rect 5885 7064 5891 7296
rect 5901 7044 5907 7276
rect 6013 7084 6019 7456
rect 6173 7304 6179 7536
rect 9645 7524 9651 7536
rect 6596 7517 6604 7523
rect 8413 7504 8419 7523
rect 9917 7517 9932 7523
rect 9492 7497 9500 7503
rect 6173 7124 6179 7296
rect 6189 7284 6195 7456
rect 5869 6284 5875 6516
rect 5901 6304 5907 6936
rect 6013 6504 6019 6896
rect 6029 6644 6035 6656
rect 6061 6144 6067 6676
rect 6173 6664 6179 7116
rect 6189 6704 6195 7276
rect 6212 6897 6220 6903
rect 6157 6564 6163 6656
rect 6173 6544 6179 6656
rect 5933 5504 5939 5816
rect 6045 5563 6051 5956
rect 6077 5904 6083 6036
rect 6109 5924 6115 6256
rect 6125 5944 6131 6316
rect 6125 5704 6131 5936
rect 6029 5557 6051 5563
rect 5933 5464 5939 5496
rect 5869 5124 5875 5136
rect 5725 4284 5731 4656
rect 5725 4244 5731 4276
rect 5741 4144 5747 4536
rect 5821 4243 5827 4736
rect 5805 4237 5827 4243
rect 5533 3324 5539 3696
rect 5565 3444 5571 3836
rect 5341 1304 5347 1476
rect 5357 1324 5363 1336
rect 5229 784 5235 876
rect 5341 744 5347 1096
rect 5357 1084 5363 1316
rect 5229 544 5235 656
rect 5357 324 5363 1076
rect 5405 284 5411 1076
rect 5421 824 5427 2296
rect 5565 2204 5571 3096
rect 5613 2684 5619 3376
rect 5725 2664 5731 2936
rect 5437 1724 5443 2176
rect 5476 1877 5484 1883
rect 5533 1524 5539 2176
rect 5741 2124 5747 4136
rect 5757 4124 5763 4216
rect 5757 4084 5763 4096
rect 5757 3704 5763 4056
rect 5805 3524 5811 4237
rect 5869 4063 5875 5116
rect 5885 4124 5891 5376
rect 5917 4504 5923 5096
rect 5853 4057 5875 4063
rect 5837 3904 5843 3936
rect 5757 3364 5763 3376
rect 5757 2544 5763 2676
rect 5725 2104 5731 2116
rect 5757 2104 5763 2536
rect 5773 2524 5779 2896
rect 5700 1917 5708 1923
rect 5453 684 5459 1496
rect 5725 1484 5731 2096
rect 5789 1864 5795 3476
rect 5853 2684 5859 4057
rect 5933 3944 5939 5456
rect 5949 4704 5955 5316
rect 6029 5164 6035 5557
rect 6045 5444 6051 5536
rect 6125 5224 6131 5356
rect 6141 5304 6147 5556
rect 6157 5484 6163 5856
rect 6173 5764 6179 6536
rect 6237 6264 6243 7376
rect 6573 7344 6579 7416
rect 6269 6944 6275 6956
rect 6269 6664 6275 6936
rect 6221 5364 6227 5756
rect 6173 4964 6179 5076
rect 6157 4944 6163 4956
rect 6189 4744 6195 5356
rect 6253 4703 6259 6336
rect 6301 5924 6307 6596
rect 6301 4724 6307 5296
rect 6253 4697 6275 4703
rect 5949 4684 5955 4696
rect 5965 4164 5971 4556
rect 5869 3044 5875 3876
rect 5901 3544 5907 3636
rect 5885 3044 5891 3136
rect 5949 3084 5955 3096
rect 5965 2544 5971 4096
rect 6013 3884 6019 3936
rect 5885 2124 5891 2136
rect 5837 1724 5843 1736
rect 5485 1124 5491 1316
rect 5677 1164 5683 1276
rect 5805 1104 5811 1336
rect 5821 1144 5827 1256
rect 5533 564 5539 696
rect 5597 544 5603 776
rect 5629 564 5635 956
rect 5773 804 5779 876
rect 5789 844 5795 916
rect 5805 864 5811 1096
rect 5821 704 5827 1136
rect 5853 1084 5859 2116
rect 5885 1284 5891 1516
rect 5901 1344 5907 1716
rect 5917 1684 5923 2516
rect 5965 2484 5971 2496
rect 5949 1844 5955 1916
rect 5981 1904 5987 2556
rect 6013 2264 6019 3356
rect 6029 2904 6035 4116
rect 6045 3484 6051 3576
rect 6061 3244 6067 3376
rect 6077 3084 6083 4096
rect 6093 3924 6099 3936
rect 6093 3044 6099 3856
rect 6125 3544 6131 4636
rect 6141 4244 6147 4476
rect 6157 3924 6163 4516
rect 6269 4284 6275 4697
rect 6317 4544 6323 6896
rect 6349 6504 6355 7296
rect 6605 6964 6611 7276
rect 6493 6604 6499 6696
rect 6349 6364 6355 6496
rect 6365 6344 6371 6556
rect 6365 6164 6371 6336
rect 6349 5764 6355 6056
rect 6365 6044 6371 6156
rect 6365 5744 6371 6036
rect 6365 5724 6371 5736
rect 6365 5324 6371 5416
rect 6381 5344 6387 6136
rect 6429 5504 6435 5876
rect 6461 5864 6467 5936
rect 6461 5844 6467 5856
rect 6477 5324 6483 6276
rect 6365 5284 6371 5316
rect 6493 5144 6499 5916
rect 6509 5304 6515 5696
rect 6525 5524 6531 6016
rect 6541 5884 6547 6936
rect 6589 6304 6595 6516
rect 6605 6504 6611 6956
rect 6685 6884 6691 6903
rect 6605 6264 6611 6496
rect 6605 6124 6611 6256
rect 6349 4204 6355 4236
rect 6173 4104 6179 4116
rect 6109 3304 6115 3376
rect 6125 2964 6131 3536
rect 6141 3344 6147 3476
rect 6157 3384 6163 3856
rect 6173 3704 6179 4076
rect 6189 3744 6195 4136
rect 6365 3484 6371 4316
rect 6205 3344 6211 3356
rect 6141 2784 6147 2976
rect 6173 2744 6179 2876
rect 6093 2164 6099 2436
rect 5901 1324 5907 1336
rect 5885 624 5891 1256
rect 5917 1104 5923 1116
rect 5933 1044 5939 1116
rect 5629 364 5635 556
rect 5757 504 5763 576
rect 5901 344 5907 936
rect 6045 684 6051 1476
rect 6125 944 6131 1956
rect 6141 1744 6147 2256
rect 6157 1824 6163 2656
rect 6173 2444 6179 2716
rect 6189 2504 6195 3336
rect 6237 3304 6243 3316
rect 6205 2544 6211 3276
rect 6221 1924 6227 2896
rect 6237 2304 6243 3296
rect 6269 2944 6275 3316
rect 6292 3297 6300 3303
rect 6253 2324 6259 2516
rect 6269 1304 6275 2936
rect 6333 2724 6339 3036
rect 6349 2904 6355 3016
rect 6381 2144 6387 4936
rect 6493 4504 6499 5136
rect 6509 4704 6515 5216
rect 6525 4924 6531 5516
rect 6589 5484 6595 5536
rect 6605 5484 6611 6076
rect 6685 6064 6691 6076
rect 6733 5504 6739 6736
rect 6765 6444 6771 6596
rect 6781 6144 6787 7056
rect 6797 6183 6803 7016
rect 6925 7004 6931 7116
rect 7005 6944 7011 7476
rect 7101 7084 7107 7476
rect 7245 7364 7251 7376
rect 7453 7344 7459 7476
rect 7469 7404 7475 7416
rect 7181 7144 7187 7216
rect 7101 6983 7107 7076
rect 7085 6977 7107 6983
rect 6861 6644 6867 6696
rect 6797 6177 6819 6183
rect 6797 6144 6803 6156
rect 6781 6064 6787 6096
rect 6797 6044 6803 6136
rect 6813 5884 6819 6177
rect 6861 6164 6867 6636
rect 6957 6564 6963 6896
rect 6973 6644 6979 6736
rect 6989 6704 6995 6836
rect 7085 6284 7091 6977
rect 7012 6277 7020 6283
rect 6756 5877 6764 5883
rect 6765 5764 6771 5876
rect 6525 4564 6531 4916
rect 6573 4744 6579 5376
rect 6701 5324 6707 5496
rect 6813 5484 6819 5696
rect 6845 5524 6851 5736
rect 6740 5477 6748 5483
rect 6717 5344 6723 5476
rect 6669 5144 6675 5236
rect 6589 4724 6595 4836
rect 6477 4224 6483 4476
rect 6397 3904 6403 3916
rect 6429 3484 6435 3776
rect 6509 3304 6515 3876
rect 6573 3504 6579 4716
rect 6605 4164 6611 4336
rect 6532 3337 6540 3343
rect 6573 2744 6579 2956
rect 6589 2944 6595 3756
rect 6605 2924 6611 3956
rect 6621 3904 6627 4536
rect 6637 3964 6643 4676
rect 6637 3883 6643 3936
rect 6653 3884 6659 5116
rect 6669 5084 6675 5136
rect 6685 4644 6691 5276
rect 6717 4524 6723 5336
rect 6669 4264 6675 4336
rect 6701 4124 6707 4516
rect 6749 4244 6755 4476
rect 6749 4104 6755 4136
rect 6621 3877 6643 3883
rect 6621 3404 6627 3877
rect 6605 2704 6611 2916
rect 6621 2763 6627 3256
rect 6637 3144 6643 3536
rect 6685 2764 6691 2796
rect 6621 2757 6643 2763
rect 6621 2344 6627 2736
rect 6637 2604 6643 2757
rect 6397 1844 6403 2076
rect 6621 1884 6627 2336
rect 6701 2324 6707 3056
rect 6717 2964 6723 3296
rect 6468 1517 6476 1523
rect 6253 1264 6259 1276
rect 6141 884 6147 1116
rect 6269 904 6275 1296
rect 6349 944 6355 1276
rect 6493 1124 6499 1876
rect 6397 944 6403 1096
rect 5197 264 5203 276
rect 6013 224 6019 676
rect 6045 464 6051 576
rect 6157 544 6163 856
rect 6493 724 6499 1116
rect 6564 937 6572 943
rect 6237 324 6243 636
rect 6397 557 6403 576
rect 6589 404 6595 1316
rect 6637 1144 6643 1916
rect 6685 964 6691 1916
rect 6717 1884 6723 2956
rect 6733 2724 6739 2756
rect 6733 2324 6739 2556
rect 6749 2544 6755 2716
rect 6765 2564 6771 3416
rect 6701 1464 6707 1856
rect 6717 1704 6723 1716
rect 6701 1364 6707 1456
rect 6685 704 6691 956
rect 6733 764 6739 2116
rect 6765 1904 6771 2536
rect 6781 2244 6787 4076
rect 6797 3864 6803 4356
rect 6829 4164 6835 5516
rect 6861 5243 6867 6156
rect 6925 5744 6931 5776
rect 6845 5237 6867 5243
rect 6845 4904 6851 5237
rect 6925 5084 6931 5736
rect 6957 5544 6963 5696
rect 7021 5544 7027 6096
rect 6893 4664 6899 5036
rect 6941 4724 6947 5176
rect 6957 5004 6963 5476
rect 6973 5344 6979 5356
rect 6829 3784 6835 3916
rect 6845 3304 6851 3896
rect 6989 3784 6995 5296
rect 7005 4664 7011 5056
rect 7021 4904 7027 5536
rect 7037 4944 7043 6276
rect 7101 5544 7107 6716
rect 7117 6664 7123 7096
rect 7117 6164 7123 6576
rect 7005 4564 7011 4656
rect 7037 4344 7043 4356
rect 7012 3777 7020 3783
rect 6861 3524 6867 3756
rect 7053 3744 7059 5336
rect 7101 4324 7107 5536
rect 7117 5044 7123 6156
rect 7133 5863 7139 6136
rect 7149 5884 7155 6536
rect 7181 6164 7187 6176
rect 7133 5857 7155 5863
rect 7149 5724 7155 5857
rect 7181 5384 7187 6116
rect 7197 5744 7203 5776
rect 7197 5424 7203 5476
rect 7197 5184 7203 5416
rect 7069 4164 7075 4216
rect 7101 3844 7107 4316
rect 7165 4264 7171 4496
rect 7181 4204 7187 4476
rect 7197 4204 7203 4316
rect 7133 3884 7139 4196
rect 6957 3724 6963 3736
rect 6980 3717 6988 3723
rect 6861 3444 6867 3516
rect 7069 3344 7075 3736
rect 7213 3544 7219 6916
rect 7229 6724 7235 6936
rect 7229 6084 7235 6096
rect 7261 5484 7267 5496
rect 7229 3724 7235 5356
rect 7261 5144 7267 5276
rect 7245 4444 7251 4936
rect 7277 4504 7283 6296
rect 7293 5924 7299 6716
rect 7341 6244 7347 7076
rect 7373 7024 7379 7256
rect 7453 7124 7459 7336
rect 7373 6504 7379 6516
rect 7373 6264 7379 6496
rect 7293 5484 7299 5696
rect 7293 5144 7299 5476
rect 7341 5124 7347 6136
rect 7357 5844 7363 6176
rect 7405 5564 7411 5676
rect 7389 5304 7395 5476
rect 7405 5284 7411 5556
rect 7421 5364 7427 5676
rect 7453 5524 7459 7116
rect 7485 7104 7491 7316
rect 7549 7084 7555 7376
rect 7677 7324 7683 7496
rect 7885 7344 7891 7396
rect 7780 7337 7788 7343
rect 7501 6724 7507 7036
rect 7485 6464 7491 6716
rect 7549 6544 7555 7076
rect 7709 7044 7715 7336
rect 7501 5704 7507 5716
rect 7501 5344 7507 5696
rect 7549 5504 7555 6536
rect 7613 6484 7619 6756
rect 7629 6144 7635 6176
rect 7277 4484 7283 4496
rect 7293 4304 7299 5116
rect 7309 4904 7315 4936
rect 7373 4303 7379 4716
rect 7357 4297 7379 4303
rect 7133 3484 7139 3496
rect 7229 3484 7235 3716
rect 6852 3137 6860 3143
rect 6877 3104 6883 3256
rect 6893 2944 6899 3076
rect 6909 3064 6915 3336
rect 7133 3324 7139 3476
rect 6813 2724 6819 2936
rect 6797 1924 6803 2176
rect 6813 1944 6819 2236
rect 6877 2124 6883 2536
rect 6813 1504 6819 1936
rect 6797 1324 6803 1336
rect 6829 1204 6835 2096
rect 6925 1464 6931 2256
rect 6957 2024 6963 2536
rect 6973 2284 6979 2496
rect 6941 1404 6947 1476
rect 6957 484 6963 616
rect 6989 544 6995 2996
rect 7021 1744 7027 2136
rect 7037 1864 7043 2536
rect 7053 2144 7059 2936
rect 7069 2264 7075 2276
rect 7069 2144 7075 2216
rect 7021 1504 7027 1736
rect 7021 1464 7027 1496
rect 7085 1484 7091 2256
rect 7117 2164 7123 2696
rect 7021 1424 7027 1456
rect 7133 1324 7139 2156
rect 7101 744 7107 1056
rect 7117 964 7123 1256
rect 7133 944 7139 1316
rect 7149 1264 7155 2476
rect 7165 2304 7171 2496
rect 7181 2384 7187 3376
rect 7245 2904 7251 4296
rect 7261 3904 7267 4196
rect 7165 2264 7171 2296
rect 7197 1884 7203 2696
rect 7261 2104 7267 3876
rect 7277 3324 7283 3916
rect 7325 3444 7331 4296
rect 7341 4184 7347 4216
rect 7357 3464 7363 4297
rect 7373 4104 7379 4176
rect 7405 4164 7411 5116
rect 7373 3504 7379 4036
rect 7213 1704 7219 2076
rect 7165 904 7171 1696
rect 7245 1684 7251 2096
rect 7261 1924 7267 2076
rect 7277 1744 7283 3296
rect 7357 3064 7363 3436
rect 7309 2284 7315 2916
rect 7373 2564 7379 3496
rect 7389 3444 7395 3916
rect 7437 3784 7443 4896
rect 7469 4724 7475 5156
rect 7469 4324 7475 4716
rect 7485 4544 7491 5056
rect 7613 5044 7619 5196
rect 7469 4284 7475 4296
rect 7485 3704 7491 4116
rect 7549 4064 7555 4216
rect 7613 3544 7619 4816
rect 7629 4284 7635 5676
rect 7645 4284 7651 6936
rect 7693 6664 7699 6956
rect 7668 6657 7676 6663
rect 7741 6584 7747 6716
rect 7789 6624 7795 6896
rect 7821 6684 7827 6896
rect 7661 5484 7667 5856
rect 7661 4904 7667 5396
rect 7677 5304 7683 5456
rect 7693 5223 7699 6116
rect 7789 5864 7795 6536
rect 7853 6504 7859 6536
rect 7853 6144 7859 6156
rect 7821 5904 7827 5936
rect 7869 5844 7875 6496
rect 7885 5864 7891 7336
rect 7965 6564 7971 7276
rect 8013 6944 8019 7136
rect 8045 7104 8051 7296
rect 8141 7144 8147 7376
rect 8173 7164 8179 7316
rect 7949 6544 7955 6556
rect 7732 5817 7747 5823
rect 7709 5484 7715 5496
rect 7725 5464 7731 5656
rect 7853 5344 7859 5416
rect 7693 5217 7715 5223
rect 7661 4744 7667 4896
rect 7629 4104 7635 4276
rect 7661 4244 7667 4736
rect 7693 4684 7699 4696
rect 7709 4304 7715 5217
rect 7757 4937 7772 4943
rect 7757 4584 7763 4937
rect 7828 4737 7836 4743
rect 7853 4344 7859 5316
rect 7869 4744 7875 5836
rect 7901 5363 7907 6516
rect 7965 6244 7971 6556
rect 8093 6504 8099 6536
rect 7981 5904 7987 6296
rect 8020 6277 8028 6283
rect 7901 5357 7923 5363
rect 7501 3484 7507 3536
rect 7405 2884 7411 3376
rect 7421 2484 7427 2876
rect 7453 2644 7459 3336
rect 7533 3324 7539 3476
rect 7517 2944 7523 3296
rect 7540 3077 7548 3083
rect 7613 3064 7619 3536
rect 7629 3044 7635 4096
rect 7661 3864 7667 3896
rect 7597 2904 7603 3036
rect 7332 2317 7340 2323
rect 7341 1884 7347 2276
rect 7341 1844 7347 1876
rect 7245 1524 7251 1676
rect 7012 737 7020 743
rect 7229 664 7235 1516
rect 7293 1464 7299 1736
rect 7261 884 7267 1096
rect 7293 684 7299 1456
rect 7357 684 7363 1696
rect 7373 764 7379 1896
rect 7389 1364 7395 1376
rect 7405 1344 7411 2136
rect 7469 1704 7475 2896
rect 7501 2844 7507 2876
rect 7485 2104 7491 2636
rect 7501 2624 7507 2836
rect 7597 2744 7603 2896
rect 7549 2104 7555 2556
rect 7469 1524 7475 1676
rect 7460 1517 7468 1523
rect 7485 1064 7491 2076
rect 7597 1724 7603 2736
rect 7629 1964 7635 2956
rect 7645 2544 7651 3316
rect 7677 2984 7683 4076
rect 7693 3704 7699 4036
rect 7709 3884 7715 4076
rect 7709 3564 7715 3876
rect 7709 3504 7715 3536
rect 7725 3504 7731 4116
rect 7821 3524 7827 3796
rect 7661 2644 7667 2756
rect 7677 2704 7683 2976
rect 7693 2684 7699 3456
rect 7805 2523 7811 3516
rect 7837 3444 7843 3836
rect 7853 3744 7859 4336
rect 7853 3124 7859 3336
rect 7853 2684 7859 2976
rect 7869 2904 7875 2916
rect 7885 2864 7891 3676
rect 7805 2517 7827 2523
rect 7629 1904 7635 1956
rect 7597 784 7603 1516
rect 7613 1324 7619 1356
rect 7661 1344 7667 1916
rect 7677 1884 7683 2496
rect 7693 2304 7699 2476
rect 7661 944 7667 1336
rect 7373 704 7379 756
rect 7389 744 7395 756
rect 7549 744 7555 756
rect 7293 544 7299 676
rect 7677 544 7683 1836
rect 7693 1784 7699 2096
rect 7709 1844 7715 2216
rect 7789 1804 7795 2096
rect 7821 1924 7827 2517
rect 7901 2324 7907 4956
rect 7917 4084 7923 5357
rect 7933 4704 7939 5516
rect 7949 5504 7955 5896
rect 8013 5824 8019 6096
rect 8125 5804 8131 6056
rect 8148 5737 8156 5743
rect 8093 5524 8099 5696
rect 7965 5164 7971 5256
rect 7981 5044 7987 5496
rect 8173 5384 8179 5456
rect 8189 5124 8195 5456
rect 7949 4724 7955 5036
rect 7965 4724 7971 4736
rect 7949 4644 7955 4716
rect 7949 3544 7955 3816
rect 7965 3324 7971 4696
rect 8045 4544 8051 5096
rect 8029 4284 8035 4536
rect 7949 2924 7955 3296
rect 8077 3124 8083 4696
rect 8109 3044 8115 4936
rect 8141 3624 8147 4936
rect 8221 4644 8227 7496
rect 8445 7477 8460 7483
rect 8445 7464 8451 7477
rect 8269 7184 8275 7256
rect 8269 7164 8275 7176
rect 8269 5884 8275 6536
rect 8285 5884 8291 7356
rect 8564 7317 8572 7323
rect 8397 6924 8403 7096
rect 8461 6504 8467 6676
rect 8333 5964 8339 6136
rect 8269 5524 8275 5876
rect 8349 5784 8355 6496
rect 8436 6277 8451 6283
rect 8461 6263 8467 6456
rect 8477 6324 8483 7296
rect 8557 6684 8563 6976
rect 8445 6257 8467 6263
rect 7917 2344 7923 2596
rect 7956 2337 7964 2343
rect 7805 1824 7811 1843
rect 7725 1124 7731 1696
rect 7789 1644 7795 1736
rect 7805 1144 7811 1796
rect 7805 1044 7811 1136
rect 7821 1104 7827 1916
rect 7844 1717 7852 1723
rect 7885 1484 7891 1876
rect 7901 1724 7907 1916
rect 7821 644 7827 1096
rect 7901 1084 7907 1716
rect 7901 684 7907 1076
rect 7917 704 7923 2316
rect 7997 2264 8003 2276
rect 7965 1844 7971 2136
rect 8125 1904 8131 3356
rect 7965 1504 7971 1836
rect 8013 1464 8019 1476
rect 7933 904 7939 1316
rect 8013 1164 8019 1376
rect 8013 1024 8019 1116
rect 7981 904 7987 916
rect 7293 284 7299 536
rect 6029 144 6035 216
rect 7325 144 7331 536
rect 7437 144 7443 416
rect 7485 303 7491 316
rect 7485 297 7500 303
rect 7357 24 7363 136
rect 7677 104 7683 316
rect 7741 304 7747 616
rect 7789 344 7795 636
rect 7917 304 7923 696
rect 7997 584 8003 936
rect 8029 924 8035 1856
rect 8141 1704 8147 2296
rect 8157 2244 8163 4516
rect 8237 4164 8243 5516
rect 8253 4103 8259 4636
rect 8301 4264 8307 5516
rect 8429 5344 8435 5516
rect 8429 5064 8435 5336
rect 8445 5043 8451 6257
rect 8477 5804 8483 6316
rect 8573 5924 8579 6716
rect 8509 5504 8515 5696
rect 8461 5204 8467 5336
rect 8461 5124 8467 5176
rect 8461 5064 8467 5116
rect 8445 5037 8467 5043
rect 8461 4984 8467 5037
rect 8413 4284 8419 4936
rect 8237 4097 8259 4103
rect 8237 3684 8243 4097
rect 8301 3484 8307 3856
rect 8317 3764 8323 3776
rect 8253 2524 8259 3376
rect 8029 704 8035 916
rect 8045 724 8051 1456
rect 8093 724 8099 1696
rect 8237 1484 8243 1496
rect 8269 1144 8275 2896
rect 8301 2643 8307 3476
rect 8333 2964 8339 4236
rect 8356 3537 8364 3543
rect 8285 2637 8307 2643
rect 8045 684 8051 696
rect 8013 364 8019 576
rect 8125 544 8131 996
rect 8253 544 8259 636
rect 8253 284 8259 336
rect 8269 324 8275 1136
rect 8285 944 8291 2637
rect 8301 2284 8307 2536
rect 8333 2524 8339 2956
rect 8349 2904 8355 3516
rect 8365 3344 8371 3456
rect 8365 2144 8371 3336
rect 8413 3084 8419 4176
rect 8429 3843 8435 4976
rect 8477 4724 8483 5276
rect 8477 4704 8483 4716
rect 8509 4664 8515 5496
rect 8525 5284 8531 5856
rect 8445 3864 8451 3876
rect 8429 3837 8451 3843
rect 8349 1964 8355 1976
rect 8365 1764 8371 2136
rect 8381 2104 8387 2896
rect 8413 2204 8419 2976
rect 8445 2604 8451 3837
rect 8461 3764 8467 3896
rect 8509 3504 8515 4096
rect 8525 3944 8531 4336
rect 8541 2924 8547 5916
rect 8573 5464 8579 5496
rect 8589 5484 8595 6936
rect 8685 6284 8691 6856
rect 8557 5264 8563 5376
rect 8557 4284 8563 5256
rect 8589 4924 8595 4956
rect 8580 4717 8588 4723
rect 8605 4504 8611 5856
rect 8653 5464 8659 6136
rect 8669 5704 8675 6096
rect 8717 5704 8723 5916
rect 8541 2583 8547 2736
rect 8525 2577 8547 2583
rect 8381 1284 8387 2096
rect 8445 1844 8451 2176
rect 8477 2024 8483 2536
rect 8525 1544 8531 2577
rect 8557 1864 8563 2916
rect 8477 1084 8483 1336
rect 8349 964 8355 1056
rect 8285 564 8291 936
rect 8541 904 8547 1756
rect 8573 1324 8579 4256
rect 8605 4124 8611 4236
rect 8605 3324 8611 4116
rect 8621 3944 8627 5456
rect 8637 4704 8643 5336
rect 8669 5304 8675 5696
rect 8717 5484 8723 5536
rect 8717 4304 8723 4576
rect 8733 4284 8739 5916
rect 8733 3864 8739 4136
rect 8589 1944 8595 3096
rect 8701 2544 8707 3736
rect 8717 2684 8723 2736
rect 8676 2137 8684 2143
rect 8573 964 8579 1316
rect 8589 1124 8595 1936
rect 8269 304 8275 316
rect 8285 284 8291 556
rect 8269 264 8275 276
rect 8301 264 8307 536
rect 8461 504 8467 836
rect 8685 724 8691 916
rect 8477 544 8483 556
rect 8317 184 8323 316
rect 8749 244 8755 7476
rect 8829 7124 8835 7256
rect 8829 6944 8835 7116
rect 8765 4704 8771 6576
rect 8765 4664 8771 4696
rect 8765 4624 8771 4636
rect 8781 4524 8787 6636
rect 8797 6504 8803 6596
rect 8813 6244 8819 6376
rect 8845 5784 8851 7476
rect 9549 7464 9555 7496
rect 9709 7464 9715 7476
rect 9284 7457 9292 7463
rect 8861 7117 8876 7123
rect 8877 7084 8883 7096
rect 8877 6684 8883 7076
rect 8909 6284 8915 6936
rect 8973 6544 8979 7116
rect 8813 5124 8819 5676
rect 8893 4504 8899 5776
rect 8909 4684 8915 6276
rect 8941 4664 8947 5876
rect 8957 5524 8963 5616
rect 8957 5304 8963 5436
rect 8973 5364 8979 5496
rect 8989 5464 8995 7116
rect 9005 6004 9011 6136
rect 9005 5664 9011 5696
rect 8765 3884 8771 3896
rect 8765 3784 8771 3836
rect 8813 3043 8819 4076
rect 8861 3944 8867 4176
rect 8893 3964 8899 4116
rect 8797 3037 8819 3043
rect 8797 1444 8803 3037
rect 8813 1924 8819 2556
rect 8813 1363 8819 1896
rect 8797 1357 8819 1363
rect 8797 644 8803 1357
rect 8813 1064 8819 1336
rect 8861 904 8867 3936
rect 8877 3444 8883 3856
rect 8909 3744 8915 4656
rect 8925 4244 8931 4316
rect 8909 3484 8915 3736
rect 8909 3044 8915 3476
rect 8925 2244 8931 2716
rect 8957 2644 8963 5296
rect 9021 4544 9027 6676
rect 9037 6644 9043 7416
rect 9053 6664 9059 7316
rect 9069 6724 9075 6976
rect 9117 6644 9123 6876
rect 9037 5924 9043 6476
rect 9037 5384 9043 5456
rect 9037 5184 9043 5336
rect 9053 5164 9059 5516
rect 9069 5504 9075 6636
rect 9085 5344 9091 5356
rect 8973 3484 8979 4156
rect 8989 3164 8995 3956
rect 9005 2684 9011 4536
rect 9069 4084 9075 4936
rect 9021 3544 9027 3556
rect 9069 3444 9075 3956
rect 9117 3904 9123 5736
rect 9149 4684 9155 4976
rect 9133 4284 9139 4496
rect 9149 4244 9155 4676
rect 9165 4444 9171 6116
rect 9133 3924 9139 4176
rect 9117 3504 9123 3836
rect 9149 3524 9155 4176
rect 9165 3864 9171 4276
rect 9101 3084 9107 3096
rect 8893 1464 8899 1516
rect 8909 964 8915 1876
rect 8925 1144 8931 1856
rect 8957 1504 8963 2236
rect 8973 1444 8979 1476
rect 8813 644 8819 696
rect 8877 264 8883 896
rect 8909 164 8915 956
rect 8925 504 8931 1136
rect 8925 324 8931 496
rect 8932 277 8940 283
rect 8957 244 8963 1376
rect 8989 184 8995 2236
rect 9005 2164 9011 2676
rect 9021 2524 9027 3036
rect 9133 2944 9139 3476
rect 9005 1484 9011 2156
rect 9133 2144 9139 2936
rect 9149 2564 9155 2836
rect 9181 2484 9187 7456
rect 9309 7384 9315 7456
rect 9261 7364 9267 7376
rect 9421 7064 9427 7216
rect 9373 6924 9379 7036
rect 9437 6984 9443 7216
rect 9549 7044 9555 7456
rect 9604 7437 9612 7443
rect 9204 6537 9212 6543
rect 9204 4657 9212 4663
rect 9229 4564 9235 6136
rect 9325 5783 9331 6876
rect 9373 6724 9379 6916
rect 9373 6104 9379 6276
rect 9325 5777 9347 5783
rect 9341 5304 9347 5777
rect 9373 5284 9379 6096
rect 9204 3117 9212 3123
rect 9229 2924 9235 3916
rect 9245 3104 9251 4276
rect 9261 3924 9267 4056
rect 9261 3084 9267 3896
rect 9277 3104 9283 4136
rect 9341 3843 9347 4716
rect 9357 4244 9363 4316
rect 9373 4284 9379 5276
rect 9389 4744 9395 5696
rect 9405 5484 9411 6296
rect 9437 5744 9443 6956
rect 9453 6764 9459 6876
rect 9469 6644 9475 7016
rect 9501 5704 9507 6876
rect 9533 6744 9539 6936
rect 9565 6183 9571 6716
rect 9549 6177 9571 6183
rect 9524 6157 9532 6163
rect 9469 5684 9475 5696
rect 9421 4904 9427 5616
rect 9325 3837 9347 3843
rect 9293 3383 9299 3736
rect 9325 3504 9331 3837
rect 9389 3524 9395 4736
rect 9293 3377 9315 3383
rect 9293 3104 9299 3116
rect 9309 2984 9315 3377
rect 9197 2644 9203 2656
rect 9149 2284 9155 2476
rect 9149 2104 9155 2276
rect 9229 1964 9235 2896
rect 9309 2724 9315 2976
rect 9373 2944 9379 3356
rect 9245 1884 9251 2536
rect 9213 1424 9219 1696
rect 9133 1304 9139 1336
rect 9021 684 9027 1276
rect 9133 964 9139 1136
rect 9229 924 9235 1376
rect 9245 1344 9251 1356
rect 9261 1324 9267 2516
rect 9277 2317 9283 2336
rect 9284 2277 9292 2283
rect 9309 1844 9315 2496
rect 9389 1904 9395 3336
rect 9437 1783 9443 5356
rect 9549 5324 9555 6177
rect 9581 5884 9587 5916
rect 9476 5117 9484 5123
rect 9501 4184 9507 4356
rect 9549 4144 9555 5316
rect 9581 4944 9587 4956
rect 9597 4684 9603 5336
rect 9613 5224 9619 7316
rect 9629 5084 9635 7116
rect 9613 4924 9619 4936
rect 9565 4084 9571 4156
rect 9469 3704 9475 3796
rect 9517 2804 9523 4076
rect 9613 4024 9619 4896
rect 9533 3304 9539 3356
rect 9613 2984 9619 3736
rect 9485 2284 9491 2656
rect 9629 2584 9635 5056
rect 9517 2264 9523 2296
rect 9476 2157 9484 2163
rect 9453 1944 9459 2156
rect 9421 1777 9443 1783
rect 9309 1524 9315 1536
rect 9421 1503 9427 1777
rect 9437 1524 9443 1756
rect 9453 1744 9459 1756
rect 9421 1497 9443 1503
rect 9412 1477 9420 1483
rect 9309 904 9315 1456
rect 9389 524 9395 1036
rect 9437 724 9443 1497
rect 9469 1084 9475 1976
rect 9533 1404 9539 1776
rect 9645 1064 9651 7296
rect 9661 6684 9667 6936
rect 9661 6504 9667 6676
rect 9677 6564 9683 7036
rect 9693 6904 9699 7256
rect 9661 6324 9667 6496
rect 9661 5084 9667 6316
rect 9677 6204 9683 6536
rect 9709 6304 9715 7336
rect 9700 5737 9708 5743
rect 9709 5284 9715 5696
rect 9661 4504 9667 5076
rect 9725 4764 9731 6896
rect 9741 5524 9747 6556
rect 9757 5783 9763 6136
rect 9805 5784 9811 6056
rect 9757 5777 9779 5783
rect 9773 5304 9779 5777
rect 9821 5404 9827 7516
rect 9917 7504 9923 7517
rect 9940 7477 9948 7483
rect 9837 6284 9843 7476
rect 9853 7124 9859 7136
rect 9837 5524 9843 6256
rect 9853 6044 9859 7096
rect 9869 6104 9875 7136
rect 9901 6504 9907 6696
rect 9917 6644 9923 7296
rect 9876 6077 9884 6083
rect 9821 4964 9827 5376
rect 9757 4944 9763 4956
rect 9677 3484 9683 4696
rect 9700 4677 9708 4683
rect 9780 4537 9788 4543
rect 9677 2924 9683 3476
rect 9677 2544 9683 2896
rect 9693 1064 9699 4496
rect 9853 4324 9859 5716
rect 9828 4277 9836 4283
rect 9853 3884 9859 4316
rect 9709 2944 9715 3536
rect 9789 1504 9795 2576
rect 9837 2304 9843 2676
rect 9501 324 9507 736
rect 9540 717 9548 723
rect 9693 284 9699 1056
rect 9805 544 9811 2136
rect 9821 944 9827 1076
rect 9732 317 9740 323
rect 9156 177 9164 183
rect 8116 137 8124 143
rect 8509 124 8515 156
rect 9709 144 9715 276
rect 9757 164 9763 316
rect 9821 184 9827 876
rect 9837 224 9843 236
rect 9853 104 9859 3736
rect 9869 144 9875 6056
rect 9885 5704 9891 6036
rect 9901 5724 9907 5736
rect 9885 5684 9891 5696
rect 9917 5364 9923 6116
rect 9885 4604 9891 5296
rect 9933 5004 9939 6576
rect 10013 5344 10019 6536
rect 9933 4744 9939 4936
rect 10013 4684 10019 4856
rect 10029 4844 10035 4896
rect 9885 4104 9891 4456
rect 9901 3524 9907 4596
rect 9917 4164 9923 4676
rect 9917 4124 9923 4136
rect 9917 3804 9923 4076
rect 10045 3884 10051 5816
rect 10269 5324 10275 5376
rect 10077 5304 10083 5316
rect 9917 2904 9923 2916
rect 9917 2804 9923 2876
rect 9892 2317 9900 2323
rect 9933 2284 9939 2936
rect 9981 2724 9987 3376
rect 10029 3084 10035 3336
rect 9965 2604 9971 2716
rect 9885 684 9891 2156
rect 9901 1804 9907 1896
rect 9933 1704 9939 2276
rect 10061 1784 10067 4196
rect 10077 3144 10083 5296
rect 10205 4644 10211 4956
rect 10100 3517 10108 3523
rect 10093 724 10099 3056
rect 10109 1884 10115 1896
rect 10100 537 10108 543
rect 10173 524 10179 716
rect 9965 184 9971 276
rect 10020 97 10028 103
<< m5contact >>
rect 268 7116 276 7124
rect 428 6936 436 6944
rect 412 6496 420 6504
rect 236 3896 244 3904
rect 204 3876 212 3884
rect 220 3856 228 3864
rect 300 3816 308 3824
rect 652 5316 660 5324
rect 668 4576 676 4584
rect 876 6656 884 6664
rect 1068 7096 1076 7104
rect 972 6936 980 6944
rect 860 6576 868 6584
rect 892 6576 900 6584
rect 892 6116 900 6124
rect 1084 6576 1092 6584
rect 1132 7096 1140 7104
rect 1132 6696 1140 6704
rect 1116 6116 1124 6124
rect 1132 6116 1140 6124
rect 2476 7476 2484 7484
rect 1532 7096 1540 7104
rect 1436 6976 1444 6984
rect 1468 6976 1476 6984
rect 1308 6516 1316 6524
rect 924 5516 932 5524
rect 908 5256 916 5264
rect 508 3576 516 3584
rect 444 3376 452 3384
rect 220 1056 228 1064
rect 236 996 244 1004
rect 236 796 244 804
rect 476 2536 484 2544
rect 636 3896 644 3904
rect 572 3876 580 3884
rect 540 3576 548 3584
rect 908 4316 916 4324
rect 684 3336 692 3344
rect 556 2556 564 2564
rect 524 1716 532 1724
rect 652 2336 660 2344
rect 700 2596 708 2604
rect 716 2176 724 2184
rect 668 1876 676 1884
rect 428 676 436 684
rect 636 556 644 564
rect 1116 5756 1124 5764
rect 988 4276 996 4284
rect 1100 4876 1108 4884
rect 1100 4536 1108 4544
rect 1020 4256 1028 4264
rect 1100 4096 1108 4104
rect 1100 4076 1108 4084
rect 1100 3296 1108 3304
rect 956 2676 964 2684
rect 940 1956 948 1964
rect 668 1716 676 1724
rect 684 1096 692 1104
rect 1004 1956 1012 1964
rect 860 1056 868 1064
rect 764 656 772 664
rect 876 716 884 724
rect 1212 5056 1220 5064
rect 1148 4636 1156 4644
rect 1164 4396 1172 4404
rect 1244 4776 1252 4784
rect 1212 4076 1220 4084
rect 1148 3296 1156 3304
rect 1164 3056 1172 3064
rect 1132 2576 1140 2584
rect 1244 3376 1252 3384
rect 1244 3096 1252 3104
rect 1260 2996 1268 3004
rect 1436 6256 1444 6264
rect 1564 6116 1572 6124
rect 1596 6116 1604 6124
rect 1548 5236 1556 5244
rect 1548 4436 1556 4444
rect 1228 2476 1236 2484
rect 988 1276 996 1284
rect 1068 1276 1076 1284
rect 1084 676 1092 684
rect 988 616 996 624
rect 1596 5476 1604 5484
rect 1596 3756 1604 3764
rect 1868 7116 1876 7124
rect 1692 5776 1700 5784
rect 1740 5776 1748 5784
rect 1708 4536 1716 4544
rect 1324 2256 1332 2264
rect 1356 1796 1364 1804
rect 1436 1476 1444 1484
rect 1276 1036 1284 1044
rect 1356 1096 1364 1104
rect 1324 1036 1332 1044
rect 1532 1176 1540 1184
rect 1612 3056 1620 3064
rect 1612 2156 1620 2164
rect 1692 4256 1700 4264
rect 1756 3876 1764 3884
rect 1788 3836 1796 3844
rect 1788 3476 1796 3484
rect 2236 7116 2244 7124
rect 2092 6496 2100 6504
rect 2044 5396 2052 5404
rect 1868 4656 1876 4664
rect 1900 4656 1908 4664
rect 2204 6036 2212 6044
rect 2028 3756 2036 3764
rect 2012 3436 2020 3444
rect 1820 2536 1828 2544
rect 1740 2256 1748 2264
rect 1756 2256 1764 2264
rect 1676 2156 1684 2164
rect 1564 1096 1572 1104
rect 1804 2336 1812 2344
rect 2012 2536 2020 2544
rect 1900 2336 1908 2344
rect 1868 2276 1876 2284
rect 1804 2196 1812 2204
rect 1836 1876 1844 1884
rect 1740 1496 1748 1504
rect 1772 1096 1780 1104
rect 1868 716 1876 724
rect 2348 6516 2356 6524
rect 2412 6696 2420 6704
rect 2396 6356 2404 6364
rect 2268 5276 2276 5284
rect 2252 4676 2260 4684
rect 2140 4236 2148 4244
rect 2124 3816 2132 3824
rect 2076 3076 2084 3084
rect 2124 2676 2132 2684
rect 2172 2296 2180 2304
rect 1996 1876 2004 1884
rect 1804 536 1812 544
rect 2108 2076 2116 2084
rect 2092 1536 2100 1544
rect 2220 1936 2228 1944
rect 2044 656 2052 664
rect 2476 6336 2484 6344
rect 2716 7276 2724 7284
rect 2732 7136 2740 7144
rect 2620 6776 2628 6784
rect 2652 6776 2660 6784
rect 2332 5236 2340 5244
rect 2348 4836 2356 4844
rect 2364 4636 2372 4644
rect 2460 4876 2468 4884
rect 2700 6656 2708 6664
rect 2636 6336 2644 6344
rect 2524 5476 2532 5484
rect 2524 5396 2532 5404
rect 2508 4716 2516 4724
rect 2492 4116 2500 4124
rect 2476 3516 2484 3524
rect 2460 3496 2468 3504
rect 2492 3496 2500 3504
rect 2428 3096 2436 3104
rect 2380 2556 2388 2564
rect 2780 7116 2788 7124
rect 2764 6916 2772 6924
rect 2860 6576 2868 6584
rect 3180 7316 3188 7324
rect 3228 7276 3236 7284
rect 3244 7136 3252 7144
rect 2940 6916 2948 6924
rect 2908 6336 2916 6344
rect 2844 6136 2852 6144
rect 3100 6076 3108 6084
rect 2780 5776 2788 5784
rect 2572 4956 2580 4964
rect 2668 4956 2676 4964
rect 2476 2076 2484 2084
rect 2476 2056 2484 2064
rect 2444 1876 2452 1884
rect 2332 1816 2340 1824
rect 2268 1476 2276 1484
rect 2252 996 2260 1004
rect 2572 4696 2580 4704
rect 2684 4196 2692 4204
rect 2732 5336 2740 5344
rect 2860 5336 2868 5344
rect 2796 4916 2804 4924
rect 2764 4476 2772 4484
rect 2732 4196 2740 4204
rect 2540 1536 2548 1544
rect 2652 1936 2660 1944
rect 2700 3476 2708 3484
rect 2700 3096 2708 3104
rect 2860 3096 2868 3104
rect 2732 2156 2740 2164
rect 2732 2076 2740 2084
rect 1628 256 1636 264
rect 1836 256 1844 264
rect 2908 2716 2916 2724
rect 2860 2336 2868 2344
rect 2780 2236 2788 2244
rect 2828 1936 2836 1944
rect 3036 5756 3044 5764
rect 3036 4876 3044 4884
rect 3324 7096 3332 7104
rect 3324 7056 3332 7064
rect 3244 6336 3252 6344
rect 3164 5716 3172 5724
rect 3196 5716 3204 5724
rect 3164 5536 3172 5544
rect 3308 5436 3316 5444
rect 3164 4436 3172 4444
rect 3068 2536 3076 2544
rect 3164 3716 3172 3724
rect 3148 3456 3156 3464
rect 3084 2256 3092 2264
rect 3132 2196 3140 2204
rect 3020 2156 3028 2164
rect 3260 5256 3268 5264
rect 3404 6916 3412 6924
rect 4140 7476 4148 7484
rect 3628 7316 3636 7324
rect 3420 5396 3428 5404
rect 3420 5356 3428 5364
rect 3340 4716 3348 4724
rect 3372 4716 3380 4724
rect 3228 4256 3236 4264
rect 3164 2316 3172 2324
rect 2940 1736 2948 1744
rect 2860 1376 2868 1384
rect 2844 1096 2852 1104
rect 3132 936 3140 944
rect 3068 676 3076 684
rect 2972 556 2980 564
rect 3116 556 3124 564
rect 3372 4696 3380 4704
rect 3404 4116 3412 4124
rect 3404 4096 3412 4104
rect 3404 3736 3412 3744
rect 3708 6656 3716 6664
rect 3868 7276 3876 7284
rect 4108 7056 4116 7064
rect 4220 6896 4228 6904
rect 3836 6696 3844 6704
rect 3756 6276 3764 6284
rect 3820 6256 3828 6264
rect 3964 6236 3972 6244
rect 3948 6136 3956 6144
rect 3980 6116 3988 6124
rect 3820 5496 3828 5504
rect 3628 4876 3636 4884
rect 3388 3496 3396 3504
rect 3356 3476 3364 3484
rect 3356 3076 3364 3084
rect 3356 2656 3364 2664
rect 3340 2296 3348 2304
rect 3388 2656 3396 2664
rect 3308 1676 3316 1684
rect 3180 536 3188 544
rect 3196 476 3204 484
rect 3308 476 3316 484
rect 3372 936 3380 944
rect 3500 2696 3508 2704
rect 3420 2476 3428 2484
rect 3420 2456 3428 2464
rect 3500 2336 3508 2344
rect 3420 1676 3428 1684
rect 3420 1096 3428 1104
rect 3580 2896 3588 2904
rect 3852 4896 3860 4904
rect 3852 4496 3860 4504
rect 3948 5496 3956 5504
rect 4012 6636 4020 6644
rect 4012 6276 4020 6284
rect 4028 6256 4036 6264
rect 4012 6096 4020 6104
rect 4204 6376 4212 6384
rect 4060 6276 4068 6284
rect 4412 6636 4420 6644
rect 4012 4896 4020 4904
rect 3868 4476 3876 4484
rect 3756 4296 3764 4304
rect 3612 4096 3620 4104
rect 3612 3456 3620 3464
rect 3580 2636 3588 2644
rect 3580 2236 3588 2244
rect 3580 2216 3588 2224
rect 3596 1056 3604 1064
rect 4092 5236 4100 5244
rect 4236 5356 4244 5364
rect 4156 4896 4164 4904
rect 4092 4876 4100 4884
rect 4156 4556 4164 4564
rect 3948 4256 3956 4264
rect 3916 3916 3924 3924
rect 3852 3456 3860 3464
rect 3740 3076 3748 3084
rect 3964 3516 3972 3524
rect 4108 4256 4116 4264
rect 4060 3936 4068 3944
rect 4012 3776 4020 3784
rect 4044 3776 4052 3784
rect 4012 3456 4020 3464
rect 3996 3436 4004 3444
rect 3948 3376 3956 3384
rect 3820 2576 3828 2584
rect 3820 2316 3828 2324
rect 4188 4496 4196 4504
rect 4380 5536 4388 5544
rect 4364 5496 4372 5504
rect 4476 6096 4484 6104
rect 4524 6436 4532 6444
rect 4492 5516 4500 5524
rect 4476 5036 4484 5044
rect 4508 5036 4516 5044
rect 4476 4656 4484 4664
rect 4252 3436 4260 3444
rect 4268 3436 4276 3444
rect 4236 3236 4244 3244
rect 4204 3136 4212 3144
rect 4188 3076 4196 3084
rect 4220 2876 4228 2884
rect 4540 6096 4548 6104
rect 4652 5936 4660 5944
rect 4700 5756 4708 5764
rect 4316 3316 4324 3324
rect 4476 3236 4484 3244
rect 4348 3076 4356 3084
rect 4332 2896 4340 2904
rect 4300 2776 4308 2784
rect 4124 2696 4132 2704
rect 4060 2436 4068 2444
rect 3932 2056 3940 2064
rect 3916 1876 3924 1884
rect 3644 1056 3652 1064
rect 3580 676 3588 684
rect 3388 656 3396 664
rect 4012 1136 4020 1144
rect 4076 2116 4084 2124
rect 4140 1856 4148 1864
rect 4140 1496 4148 1504
rect 4316 2676 4324 2684
rect 4476 2736 4484 2744
rect 4332 2136 4340 2144
rect 4300 2116 4308 2124
rect 4444 1876 4452 1884
rect 4316 1476 4324 1484
rect 4524 3116 4532 3124
rect 4572 4316 4580 4324
rect 4556 3096 4564 3104
rect 4716 5556 4724 5564
rect 4764 6716 4772 6724
rect 4796 6296 4804 6304
rect 4844 6296 4852 6304
rect 4764 6136 4772 6144
rect 4780 6136 4788 6144
rect 4780 5756 4788 5764
rect 4652 4556 4660 4564
rect 4700 3756 4708 3764
rect 4604 3516 4612 3524
rect 4572 3076 4580 3084
rect 4604 2696 4612 2704
rect 4652 2736 4660 2744
rect 6092 7516 6100 7524
rect 5084 6736 5092 6744
rect 5180 6636 5188 6644
rect 4924 5616 4932 5624
rect 4956 6276 4964 6284
rect 5004 5536 5012 5544
rect 5100 5916 5108 5924
rect 5292 6296 5300 6304
rect 5260 6116 5268 6124
rect 5116 5396 5124 5404
rect 4812 5276 4820 5284
rect 4732 3756 4740 3764
rect 4780 3476 4788 3484
rect 4700 2356 4708 2364
rect 4620 2296 4628 2304
rect 4316 1376 4324 1384
rect 4300 1136 4308 1144
rect 4220 556 4228 564
rect 4556 1736 4564 1744
rect 4684 1076 4692 1084
rect 4940 4936 4948 4944
rect 4844 4316 4852 4324
rect 4956 4136 4964 4144
rect 4812 3036 4820 3044
rect 4844 3036 4852 3044
rect 4796 2136 4804 2144
rect 5196 4696 5204 4704
rect 5084 4476 5092 4484
rect 5164 4176 5172 4184
rect 4876 2656 4884 2664
rect 4844 1856 4852 1864
rect 4780 1616 4788 1624
rect 4972 2696 4980 2704
rect 5004 2716 5012 2724
rect 5116 3096 5124 3104
rect 5148 3776 5156 3784
rect 5180 3356 5188 3364
rect 5132 2796 5140 2804
rect 5180 2876 5188 2884
rect 5196 2796 5204 2804
rect 5388 7296 5396 7304
rect 5388 5916 5396 5924
rect 5372 5876 5380 5884
rect 5276 4636 5284 4644
rect 5308 4636 5316 4644
rect 5756 6656 5764 6664
rect 5772 6576 5780 6584
rect 5596 5876 5604 5884
rect 5692 5756 5700 5764
rect 5340 3476 5348 3484
rect 5260 3436 5268 3444
rect 5772 6496 5780 6504
rect 5740 6116 5748 6124
rect 5708 5676 5716 5684
rect 5580 5336 5588 5344
rect 5484 4716 5492 4724
rect 5452 4116 5460 4124
rect 5484 3116 5492 3124
rect 5356 2296 5364 2304
rect 5020 896 5028 904
rect 4860 556 4868 564
rect 4460 516 4468 524
rect 4652 436 4660 444
rect 5084 436 5092 444
rect 5100 356 5108 364
rect 5180 356 5188 364
rect 5532 3836 5540 3844
rect 5596 4336 5604 4344
rect 6604 7516 6612 7524
rect 9644 7516 9652 7524
rect 8412 7496 8420 7504
rect 9484 7496 9492 7504
rect 6188 7276 6196 7284
rect 5884 6316 5892 6324
rect 6028 6636 6036 6644
rect 6220 6896 6228 6904
rect 6172 6656 6180 6664
rect 6076 6036 6084 6044
rect 5948 5916 5956 5924
rect 5932 5456 5940 5464
rect 5868 5136 5876 5144
rect 5724 4676 5732 4684
rect 5724 4236 5732 4244
rect 5628 3876 5636 3884
rect 5564 3436 5572 3444
rect 5548 3356 5556 3364
rect 5388 2436 5396 2444
rect 5404 1076 5412 1084
rect 5724 3076 5732 3084
rect 5596 2516 5604 2524
rect 5436 2176 5444 2184
rect 5484 1876 5492 1884
rect 5756 4116 5764 4124
rect 5756 4096 5764 4104
rect 5788 3536 5796 3544
rect 5916 4496 5924 4504
rect 5884 4116 5892 4124
rect 5836 3896 5844 3904
rect 5756 3356 5764 3364
rect 5724 2116 5732 2124
rect 5756 2096 5764 2104
rect 5708 1916 5716 1924
rect 5836 3456 5844 3464
rect 5948 5316 5956 5324
rect 6140 5556 6148 5564
rect 6044 5436 6052 5444
rect 6572 7336 6580 7344
rect 6380 7296 6388 7304
rect 6268 6956 6276 6964
rect 6172 5756 6180 5764
rect 6220 5756 6228 5764
rect 6108 5096 6116 5104
rect 6156 4936 6164 4944
rect 5948 4696 5956 4704
rect 6108 4556 6116 4564
rect 5964 4096 5972 4104
rect 5932 3936 5940 3944
rect 5948 3096 5956 3104
rect 5868 3036 5876 3044
rect 5884 3036 5892 3044
rect 5996 2936 6004 2944
rect 5964 2536 5972 2544
rect 5884 2136 5892 2144
rect 5836 1716 5844 1724
rect 5804 1096 5812 1104
rect 5532 556 5540 564
rect 5900 1716 5908 1724
rect 5964 2476 5972 2484
rect 6044 3576 6052 3584
rect 6092 3916 6100 3924
rect 6140 3936 6148 3944
rect 6956 7276 6964 7284
rect 6364 6036 6372 6044
rect 6460 5836 6468 5844
rect 6364 5276 6372 5284
rect 6684 6876 6692 6884
rect 6188 4156 6196 4164
rect 6172 4116 6180 4124
rect 6108 3296 6116 3304
rect 6204 3356 6212 3364
rect 6172 3096 6180 3104
rect 6140 2776 6148 2784
rect 6172 2736 6180 2744
rect 6124 1956 6132 1964
rect 5900 1316 5908 1324
rect 5916 1096 5924 1104
rect 5756 576 5764 584
rect 6236 3316 6244 3324
rect 6300 3296 6308 3304
rect 6252 2516 6260 2524
rect 6684 6056 6692 6064
rect 7244 7356 7252 7364
rect 7468 7396 7476 7404
rect 6860 6696 6868 6704
rect 6796 6156 6804 6164
rect 6780 6136 6788 6144
rect 6780 6096 6788 6104
rect 6988 6696 6996 6704
rect 7020 6276 7028 6284
rect 6764 5876 6772 5884
rect 6700 5496 6708 5504
rect 6732 5496 6740 5504
rect 6588 5476 6596 5484
rect 6748 5476 6756 5484
rect 6700 5316 6708 5324
rect 6524 4556 6532 4564
rect 6396 3896 6404 3904
rect 6588 4676 6596 4684
rect 6604 4156 6612 4164
rect 6604 3956 6612 3964
rect 6524 3336 6532 3344
rect 6636 3956 6644 3964
rect 6620 3896 6628 3904
rect 6684 4636 6692 4644
rect 6668 4336 6676 4344
rect 6748 4236 6756 4244
rect 6572 2736 6580 2744
rect 6700 3056 6708 3064
rect 6684 2756 6692 2764
rect 6636 1916 6644 1924
rect 6396 1836 6404 1844
rect 6476 1516 6484 1524
rect 6252 1276 6260 1284
rect 6444 1276 6452 1284
rect 6396 936 6404 944
rect 6012 676 6020 684
rect 6044 676 6052 684
rect 6572 936 6580 944
rect 6396 576 6404 584
rect 6636 1136 6644 1144
rect 6732 2776 6740 2784
rect 6732 2556 6740 2564
rect 6764 2556 6772 2564
rect 6764 2536 6772 2544
rect 6732 2116 6740 2124
rect 6716 1716 6724 1724
rect 6940 5176 6948 5184
rect 6924 5076 6932 5084
rect 6972 5336 6980 5344
rect 6892 4656 6900 4664
rect 6892 4096 6900 4104
rect 6812 3876 6820 3884
rect 6844 3896 6852 3904
rect 6828 3776 6836 3784
rect 7196 6956 7204 6964
rect 7116 6576 7124 6584
rect 7036 4336 7044 4344
rect 7004 3776 7012 3784
rect 7180 6156 7188 6164
rect 7196 5736 7204 5744
rect 7196 5476 7204 5484
rect 7116 5036 7124 5044
rect 7068 4216 7076 4224
rect 7196 4316 7204 4324
rect 7132 4196 7140 4204
rect 6956 3736 6964 3744
rect 6972 3716 6980 3724
rect 7276 6656 7284 6664
rect 7228 6096 7236 6104
rect 7260 5496 7268 5504
rect 7260 5276 7268 5284
rect 7292 5136 7300 5144
rect 7356 5836 7364 5844
rect 7420 5676 7428 5684
rect 7484 7096 7492 7104
rect 7788 7336 7796 7344
rect 7676 7316 7684 7324
rect 7708 7036 7716 7044
rect 7612 6756 7620 6764
rect 7628 6136 7636 6144
rect 7628 5676 7636 5684
rect 7276 4476 7284 4484
rect 7308 4896 7316 4904
rect 7228 3716 7236 3724
rect 7212 3536 7220 3544
rect 7132 3496 7140 3504
rect 6860 3136 6868 3144
rect 6780 2236 6788 2244
rect 6812 2236 6820 2244
rect 6796 2176 6804 2184
rect 6796 1336 6804 1344
rect 6940 1476 6948 1484
rect 7068 2276 7076 2284
rect 7068 2136 7076 2144
rect 7100 2156 7108 2164
rect 7084 1476 7092 1484
rect 7116 1256 7124 1264
rect 7340 4176 7348 4184
rect 7340 4156 7348 4164
rect 7340 3736 7348 3744
rect 7372 4176 7380 4184
rect 7420 4156 7428 4164
rect 7324 3436 7332 3444
rect 7356 3436 7364 3444
rect 7196 1876 7204 1884
rect 7148 1256 7156 1264
rect 7260 1916 7268 1924
rect 7468 4716 7476 4724
rect 7612 4896 7620 4904
rect 7612 4816 7620 4824
rect 7468 4276 7476 4284
rect 7596 4216 7604 4224
rect 7676 6656 7684 6664
rect 7868 6656 7876 6664
rect 7676 5456 7684 5464
rect 7852 6156 7860 6164
rect 7820 5896 7828 5904
rect 8172 7316 8180 7324
rect 8140 7136 8148 7144
rect 8028 7096 8036 7104
rect 8044 7096 8052 7104
rect 7948 6536 7956 6544
rect 7724 5816 7732 5824
rect 7708 5476 7716 5484
rect 7724 5456 7732 5464
rect 7852 5336 7860 5344
rect 7692 4676 7700 4684
rect 7836 4736 7844 4744
rect 8092 6496 8100 6504
rect 8140 6476 8148 6484
rect 7964 6236 7972 6244
rect 8028 6276 8036 6284
rect 7676 4276 7684 4284
rect 7660 4236 7668 4244
rect 7708 4116 7716 4124
rect 7500 3536 7508 3544
rect 7404 2876 7412 2884
rect 7532 3316 7540 3324
rect 7532 3076 7540 3084
rect 7612 3056 7620 3064
rect 7596 3036 7604 3044
rect 7628 3036 7636 3044
rect 7596 2896 7604 2904
rect 7340 2316 7348 2324
rect 7340 1836 7348 1844
rect 7020 736 7028 744
rect 7356 1696 7364 1704
rect 7388 1356 7396 1364
rect 7500 2876 7508 2884
rect 7612 2736 7620 2744
rect 7484 2096 7492 2104
rect 7468 1696 7476 1704
rect 7468 1516 7476 1524
rect 7724 3496 7732 3504
rect 7868 4116 7876 4124
rect 7836 3436 7844 3444
rect 7852 3336 7860 3344
rect 7868 2916 7876 2924
rect 7580 1316 7588 1324
rect 7612 1356 7620 1364
rect 7692 2476 7700 2484
rect 7676 1836 7684 1844
rect 7660 1336 7668 1344
rect 7388 736 7396 744
rect 7548 736 7556 744
rect 7372 696 7380 704
rect 7356 676 7364 684
rect 7708 1836 7716 1844
rect 8044 5896 8052 5904
rect 8156 5736 8164 5744
rect 8092 5516 8100 5524
rect 8188 5456 8196 5464
rect 7948 5036 7956 5044
rect 7980 5036 7988 5044
rect 7964 4736 7972 4744
rect 7948 4636 7956 4644
rect 7948 3816 7956 3824
rect 8076 4696 8084 4704
rect 7980 3356 7988 3364
rect 8444 7456 8452 7464
rect 8316 7396 8324 7404
rect 8236 6536 8244 6544
rect 8572 7316 8580 7324
rect 8460 6456 8468 6464
rect 8428 6276 8436 6284
rect 8540 6496 8548 6504
rect 8220 4636 8228 4644
rect 8028 2916 8036 2924
rect 7964 2336 7972 2344
rect 7804 1816 7812 1824
rect 7836 1716 7844 1724
rect 7804 1036 7812 1044
rect 7996 2256 8004 2264
rect 8012 1476 8020 1484
rect 7932 1316 7940 1324
rect 7948 1296 7956 1304
rect 8012 1116 8020 1124
rect 7980 916 7988 924
rect 7788 636 7796 644
rect 7820 636 7828 644
rect 7308 316 7316 324
rect 5964 156 5972 164
rect 7500 296 7508 304
rect 8460 5196 8468 5204
rect 8428 4976 8436 4984
rect 8460 4976 8468 4984
rect 8412 4276 8420 4284
rect 8316 3756 8324 3764
rect 8172 3336 8180 3344
rect 8092 1696 8100 1704
rect 8236 1496 8244 1504
rect 8364 3536 8372 3544
rect 8044 676 8052 684
rect 8124 536 8132 544
rect 8332 2516 8340 2524
rect 8476 4696 8484 4704
rect 8524 4336 8532 4344
rect 8444 3856 8452 3864
rect 8412 2976 8420 2984
rect 8348 1976 8356 1984
rect 8476 3756 8484 3764
rect 8572 5496 8580 5504
rect 8572 4716 8580 4724
rect 8716 5696 8724 5704
rect 8604 4316 8612 4324
rect 8572 4256 8580 4264
rect 8444 2176 8452 2184
rect 8540 2556 8548 2564
rect 8716 5476 8724 5484
rect 8716 4136 8724 4144
rect 8684 2136 8692 2144
rect 8572 1316 8580 1324
rect 8252 276 8260 284
rect 8476 536 8484 544
rect 8268 256 8276 264
rect 8300 256 8308 264
rect 8764 4616 8772 4624
rect 9708 7476 9716 7484
rect 9292 7456 9300 7464
rect 9548 7456 9556 7464
rect 8876 7116 8884 7124
rect 8876 7096 8884 7104
rect 8972 6536 8980 6544
rect 8844 5776 8852 5784
rect 8892 5776 8900 5784
rect 8924 5356 8932 5364
rect 8956 5516 8964 5524
rect 9004 5696 9012 5704
rect 8860 4176 8868 4184
rect 8764 3896 8772 3904
rect 8764 3836 8772 3844
rect 8844 3336 8852 3344
rect 8876 3856 8884 3864
rect 8924 4236 8932 4244
rect 9036 6636 9044 6644
rect 9068 6636 9076 6644
rect 9116 6636 9124 6644
rect 9036 6476 9044 6484
rect 9052 5516 9060 5524
rect 9036 5376 9044 5384
rect 9036 5176 9044 5184
rect 9084 5356 9092 5364
rect 9020 3536 9028 3544
rect 9132 4256 9140 4264
rect 9148 4236 9156 4244
rect 9100 3836 9108 3844
rect 9148 3516 9156 3524
rect 9116 3496 9124 3504
rect 9100 3096 9108 3104
rect 8924 2236 8932 2244
rect 8956 2236 8964 2244
rect 8892 1456 8900 1464
rect 8924 1856 8932 1864
rect 8812 696 8820 704
rect 8924 316 8932 324
rect 8940 276 8948 284
rect 9052 2896 9060 2904
rect 9148 2836 9156 2844
rect 9308 7376 9316 7384
rect 9260 7356 9268 7364
rect 9372 7036 9380 7044
rect 9612 7436 9620 7444
rect 9548 7036 9556 7044
rect 9436 6976 9444 6984
rect 9196 6536 9204 6544
rect 9212 4656 9220 4664
rect 9228 4276 9236 4284
rect 9244 4276 9252 4284
rect 9212 3116 9220 3124
rect 9260 3916 9268 3924
rect 9452 6756 9460 6764
rect 9468 6636 9476 6644
rect 9532 6156 9540 6164
rect 9468 5676 9476 5684
rect 9436 5476 9444 5484
rect 9372 4276 9380 4284
rect 9356 4236 9364 4244
rect 9292 3096 9300 3104
rect 9228 2916 9236 2924
rect 9196 2656 9204 2664
rect 9212 2516 9220 2524
rect 9148 2476 9156 2484
rect 9180 2476 9188 2484
rect 9228 1376 9236 1384
rect 9132 1136 9140 1144
rect 9244 1356 9252 1364
rect 9276 2336 9284 2344
rect 9276 2276 9284 2284
rect 9308 1836 9316 1844
rect 9468 5116 9476 5124
rect 9580 4956 9588 4964
rect 9628 5076 9636 5084
rect 9612 4936 9620 4944
rect 9612 2476 9620 2484
rect 9468 2156 9476 2164
rect 9308 1536 9316 1544
rect 9452 1736 9460 1744
rect 9420 1476 9428 1484
rect 9324 1456 9332 1464
rect 9532 1776 9540 1784
rect 9484 1336 9492 1344
rect 9676 6556 9684 6564
rect 9708 5736 9716 5744
rect 9740 6556 9748 6564
rect 9932 7516 9940 7524
rect 9932 7476 9940 7484
rect 10268 7316 10276 7324
rect 9852 7136 9860 7144
rect 9916 6636 9924 6644
rect 9932 6576 9940 6584
rect 9884 6076 9892 6084
rect 9852 6036 9860 6044
rect 9756 4956 9764 4964
rect 9660 3896 9668 3904
rect 9692 4676 9700 4684
rect 9788 4536 9796 4544
rect 9836 4276 9844 4284
rect 9788 2576 9796 2584
rect 9548 716 9556 724
rect 9740 316 9748 324
rect 9164 176 9172 184
rect 8012 136 8020 144
rect 8124 136 8132 144
rect 9836 236 9844 244
rect 9516 116 9524 124
rect 9884 6036 9892 6044
rect 9900 5736 9908 5744
rect 9884 5676 9892 5684
rect 10012 4856 10020 4864
rect 10028 4836 10036 4844
rect 9916 4136 9924 4144
rect 10268 5376 10276 5384
rect 10076 5316 10084 5324
rect 9980 3376 9988 3384
rect 9916 2916 9924 2924
rect 9916 2876 9924 2884
rect 9900 2316 9908 2324
rect 10108 3516 10116 3524
rect 10268 3116 10276 3124
rect 10108 1876 10116 1884
rect 10108 536 10116 544
rect 9964 276 9972 284
rect 10028 96 10036 104
<< metal5 >>
rect 6100 7517 6604 7523
rect 9652 7517 9787 7523
rect 9925 7517 9932 7523
rect 8413 7504 8419 7515
rect 9492 7497 10011 7503
rect 2484 7477 4140 7483
rect 9157 7477 9708 7483
rect 9940 7477 9947 7483
rect 8445 7464 8451 7475
rect 9300 7457 9548 7463
rect 9605 7437 9612 7443
rect 7476 7397 8316 7403
rect 7252 7357 9260 7363
rect 6580 7337 7788 7343
rect 3188 7317 3628 7323
rect 7684 7317 8172 7323
rect 8580 7317 10268 7323
rect 5396 7297 6380 7303
rect 2724 7277 2843 7283
rect 2853 7277 3228 7283
rect 3236 7277 3868 7283
rect 6196 7277 6956 7283
rect 2740 7137 3244 7143
rect 8148 7137 9852 7143
rect 276 7117 1868 7123
rect 2244 7117 2780 7123
rect 8869 7117 8876 7123
rect 1076 7097 1132 7103
rect 1540 7097 2683 7103
rect 2693 7097 3324 7103
rect 7492 7097 8028 7103
rect 8052 7097 8876 7103
rect 3332 7057 4108 7063
rect 7716 7037 9372 7043
rect 9541 7037 9548 7043
rect 1444 6977 1468 6983
rect 6276 6957 7196 6963
rect 436 6937 972 6943
rect 2772 6917 2940 6923
rect 2948 6917 3404 6923
rect 6213 6897 6220 6903
rect 6685 6884 6691 6895
rect 2628 6777 2652 6783
rect 7620 6757 9452 6763
rect 4837 6737 5084 6743
rect 4485 6717 4764 6723
rect 1125 6697 1132 6703
rect 2420 6697 3836 6703
rect 6868 6697 6988 6703
rect 884 6657 2700 6663
rect 2708 6657 3708 6663
rect 5764 6657 5787 6663
rect 6180 6657 7276 6663
rect 7684 6657 7868 6663
rect 4005 6637 4012 6643
rect 5188 6637 5755 6643
rect 5765 6637 6028 6643
rect 9044 6637 9068 6643
rect 868 6577 892 6583
rect 1092 6577 1115 6583
rect 2853 6577 2860 6583
rect 5780 6577 7116 6583
rect 9917 6583 9923 6636
rect 9917 6577 9932 6583
rect 9684 6557 9740 6563
rect 7956 6537 8236 6543
rect 8980 6537 9196 6543
rect 1316 6517 1947 6523
rect 1957 6517 2348 6523
rect 420 6497 2092 6503
rect 5765 6497 5772 6503
rect 8100 6497 8540 6503
rect 8148 6477 9036 6483
rect 8453 6457 8460 6463
rect 4532 6437 6139 6443
rect 4197 6377 4204 6383
rect 2484 6337 2636 6343
rect 2916 6337 3244 6343
rect 5797 6317 5884 6323
rect 4804 6297 4844 6303
rect 4852 6297 5292 6303
rect 3764 6277 4012 6283
rect 4068 6277 4956 6283
rect 7028 6277 8028 6283
rect 8436 6277 8443 6283
rect 1444 6257 3355 6263
rect 3828 6257 3995 6263
rect 4005 6257 4028 6263
rect 7941 6237 7964 6243
rect 6804 6157 7180 6163
rect 7860 6157 9532 6163
rect 3956 6137 4764 6143
rect 4788 6137 4795 6143
rect 6788 6137 7628 6143
rect 900 6117 1116 6123
rect 1140 6117 1564 6123
rect 1572 6117 1596 6123
rect 3988 6117 3995 6123
rect 5268 6117 5740 6123
rect 3365 6097 4012 6103
rect 4484 6097 4540 6103
rect 6725 6097 6780 6103
rect 6788 6097 7228 6103
rect 3101 6084 3107 6095
rect 7621 6077 9884 6083
rect 6685 6064 6691 6075
rect 2205 6044 2211 6055
rect 6084 6037 6364 6043
rect 9860 6037 9884 6043
rect 4421 5937 4652 5943
rect 5108 5917 5388 5923
rect 5396 5917 5948 5923
rect 7828 5897 8044 5903
rect 5380 5877 5499 5883
rect 5509 5877 5596 5883
rect 6149 5877 6764 5883
rect 7732 5817 7739 5823
rect 2781 5784 2787 5795
rect 1700 5777 1740 5783
rect 8852 5777 8892 5783
rect 1124 5757 2395 5763
rect 3044 5757 4700 5763
rect 4708 5757 4780 5763
rect 4837 5757 5692 5763
rect 6180 5757 6220 5763
rect 7204 5737 8156 5743
rect 9716 5737 9723 5743
rect 9893 5737 9900 5743
rect 3172 5717 3196 5723
rect 8549 5697 8716 5703
rect 8724 5697 9004 5703
rect 5716 5677 6683 5683
rect 6693 5677 7420 5683
rect 7636 5677 9468 5683
rect 9765 5677 9884 5683
rect 4925 5624 4931 5635
rect 4709 5557 4716 5563
rect 3172 5537 4380 5543
rect 4388 5537 5004 5543
rect 4500 5517 5179 5523
rect 8100 5517 8956 5523
rect 8964 5517 9052 5523
rect 3828 5497 3948 5503
rect 3956 5497 4364 5503
rect 6708 5497 6732 5503
rect 7268 5497 8572 5503
rect 1604 5477 2524 5483
rect 6596 5477 6748 5483
rect 7204 5477 7708 5483
rect 8724 5477 9436 5483
rect 5940 5457 7676 5463
rect 7732 5457 8188 5463
rect 3301 5437 3308 5443
rect 2052 5397 2524 5403
rect 3428 5397 5116 5403
rect 9044 5377 10268 5383
rect 3428 5357 4236 5363
rect 8932 5357 9084 5363
rect 2740 5337 2860 5343
rect 5588 5337 6972 5343
rect 7860 5337 7867 5343
rect 660 5317 667 5323
rect 5956 5317 6700 5323
rect 9733 5317 10076 5323
rect 2276 5277 2395 5283
rect 4581 5277 4812 5283
rect 6373 5277 7260 5283
rect 916 5257 3260 5263
rect 1556 5237 2332 5243
rect 4100 5237 5083 5243
rect 8261 5197 8460 5203
rect 6948 5177 9036 5183
rect 5876 5137 6203 5143
rect 7300 5137 7323 5143
rect 9476 5117 9755 5123
rect 6116 5097 6459 5103
rect 6917 5077 6924 5083
rect 1220 5057 1531 5063
rect 4484 5037 4508 5043
rect 7124 5037 7131 5043
rect 7956 5037 7980 5043
rect 8436 4977 8460 4983
rect 2580 4957 2668 4963
rect 9588 4957 9756 4963
rect 4948 4937 5499 4943
rect 6164 4937 9612 4943
rect 2804 4917 2843 4923
rect 3860 4897 3867 4903
rect 4020 4897 4156 4903
rect 4164 4897 4219 4903
rect 7316 4897 7612 4903
rect 1108 4877 1115 4883
rect 2468 4877 3036 4883
rect 3589 4877 3628 4883
rect 3845 4877 4092 4883
rect 2356 4837 3291 4843
rect 10021 4837 10028 4843
rect 7844 4737 7964 4743
rect 2516 4717 3340 4723
rect 3348 4717 3372 4723
rect 5492 4717 5499 4723
rect 7476 4717 8572 4723
rect 2580 4697 3372 4703
rect 5204 4697 5948 4703
rect 8084 4697 8476 4703
rect 2213 4677 2252 4683
rect 6596 4677 7227 4683
rect 7237 4677 7692 4683
rect 9125 4677 9691 4683
rect 1876 4657 1900 4663
rect 1908 4657 2459 4663
rect 2469 4657 4475 4663
rect 6900 4657 9212 4663
rect 2341 4637 2364 4643
rect 5284 4637 5308 4643
rect 7956 4637 7963 4643
rect 8765 4624 8771 4635
rect 4164 4557 4652 4563
rect 6116 4557 6524 4563
rect 1108 4537 1708 4543
rect 9701 4537 9788 4543
rect 3860 4497 3867 4503
rect 5924 4497 6779 4503
rect 2772 4477 3868 4483
rect 4485 4477 4699 4483
rect 5093 4477 6011 4483
rect 6021 4477 7276 4483
rect 3165 4444 3171 4455
rect 1541 4437 1548 4443
rect 1157 4397 1164 4403
rect 5604 4337 5723 4343
rect 6676 4337 6907 4343
rect 6917 4337 7036 4343
rect 8532 4337 8539 4343
rect 916 4317 923 4323
rect 4580 4317 4827 4323
rect 4837 4317 4844 4323
rect 7204 4317 8604 4323
rect 3764 4297 3931 4303
rect 996 4277 2779 4283
rect 7476 4277 7676 4283
rect 8420 4277 9228 4283
rect 9252 4277 9372 4283
rect 9701 4277 9836 4283
rect 1700 4257 3228 4263
rect 3956 4257 4108 4263
rect 8580 4257 9115 4263
rect 9140 4257 9147 4263
rect 5732 4237 5979 4243
rect 7668 4237 7675 4243
rect 9364 4237 9371 4243
rect 7076 4217 7596 4223
rect 2692 4197 2732 4203
rect 5157 4177 5164 4183
rect 7348 4177 7372 4183
rect 6196 4157 6604 4163
rect 7348 4157 7420 4163
rect 4901 4137 4923 4143
rect 4933 4137 4956 4143
rect 8724 4137 9916 4143
rect 1125 4117 1139 4123
rect 1108 4097 1115 4103
rect 1133 4083 1139 4117
rect 2405 4117 2492 4123
rect 3397 4117 3404 4123
rect 5445 4117 5452 4123
rect 5892 4117 6172 4123
rect 6180 4117 6203 4123
rect 7716 4117 7868 4123
rect 3412 4097 3547 4103
rect 3557 4097 3612 4103
rect 5764 4097 5964 4103
rect 5972 4097 6363 4103
rect 6900 4097 7355 4103
rect 1213 4084 1219 4095
rect 1108 4077 1139 4083
rect 6612 3957 6636 3963
rect 3973 3937 4060 3943
rect 5940 3937 6140 3943
rect 3924 3917 3995 3923
rect 6100 3917 6715 3923
rect 9268 3917 9275 3923
rect 644 3897 1947 3903
rect 212 3877 219 3883
rect 237 3863 243 3896
rect 5844 3897 6396 3903
rect 6628 3897 6844 3903
rect 8772 3897 9660 3903
rect 580 3877 1756 3883
rect 5636 3877 6812 3883
rect 228 3857 243 3863
rect 8452 3857 8876 3863
rect 1789 3844 1795 3855
rect 5533 3844 5539 3855
rect 9108 3837 9307 3843
rect 308 3817 2124 3823
rect 7941 3817 7948 3823
rect 4020 3777 4044 3783
rect 6836 3777 7004 3783
rect 1604 3757 2028 3763
rect 4708 3757 4732 3763
rect 8324 3757 8476 3763
rect 3412 3737 3419 3743
rect 6964 3737 7340 3743
rect 6980 3717 7228 3723
rect 516 3577 540 3583
rect 5796 3537 6715 3543
rect 6725 3537 7212 3543
rect 7508 3537 7739 3543
rect 8357 3537 8364 3543
rect 9028 3537 9147 3543
rect 2484 3517 3835 3523
rect 3972 3517 4604 3523
rect 9317 3517 10108 3523
rect 2468 3497 2492 3503
rect 7140 3497 7724 3503
rect 3389 3485 3395 3496
rect 1796 3477 2700 3483
rect 4788 3477 5340 3483
rect 3156 3457 3612 3463
rect 3860 3457 4012 3463
rect 4581 3457 5836 3463
rect 4004 3437 4252 3443
rect 4260 3437 4268 3443
rect 5268 3437 5275 3443
rect 7332 3437 7356 3443
rect 3941 3377 3948 3383
rect 9957 3377 9980 3383
rect 5541 3357 5548 3363
rect 5573 3357 5756 3363
rect 6212 3357 6779 3363
rect 7973 3357 7980 3363
rect 677 3337 684 3343
rect 6149 3337 6524 3343
rect 6532 3337 7852 3343
rect 8180 3337 8844 3343
rect 6244 3317 7532 3323
rect 1108 3297 1148 3303
rect 6116 3297 6300 3303
rect 4244 3237 4476 3243
rect 4212 3137 4571 3143
rect 6757 3137 6860 3143
rect 4532 3117 5484 3123
rect 9220 3117 10268 3123
rect 2436 3097 2683 3103
rect 2693 3097 2700 3103
rect 2868 3097 2875 3103
rect 4564 3097 5116 3103
rect 5285 3097 5948 3103
rect 5989 3097 6172 3103
rect 9108 3097 9292 3103
rect 2084 3077 2395 3083
rect 3364 3077 3740 3083
rect 3748 3077 3931 3083
rect 4196 3077 4348 3083
rect 4580 3077 5724 3083
rect 5765 3077 7532 3083
rect 1172 3057 1612 3063
rect 6693 3057 6700 3063
rect 4820 3037 4844 3043
rect 5861 3037 5868 3043
rect 7604 3037 7628 3043
rect 1221 2997 1260 3003
rect 6004 2937 6011 2943
rect 7876 2917 8028 2923
rect 9236 2917 9916 2923
rect 3588 2897 4332 2903
rect 7604 2897 9052 2903
rect 2917 2877 4220 2883
rect 4228 2877 5180 2883
rect 7412 2877 7500 2883
rect 5140 2797 5196 2803
rect 4293 2777 4300 2783
rect 6148 2777 6211 2783
rect 6205 2763 6211 2777
rect 6701 2777 6732 2783
rect 6205 2757 6684 2763
rect 4484 2737 4652 2743
rect 6701 2743 6707 2777
rect 6580 2737 6707 2743
rect 7365 2737 7612 2743
rect 2916 2717 5004 2723
rect 3508 2697 4124 2703
rect 4612 2697 4972 2703
rect 964 2677 2124 2683
rect 2885 2677 4316 2683
rect 3396 2657 4876 2663
rect 4884 2657 4891 2663
rect 8933 2657 9196 2663
rect 3557 2637 3580 2643
rect 677 2597 700 2603
rect 1125 2577 1132 2583
rect 3828 2577 3835 2583
rect 564 2557 2380 2563
rect 6740 2557 6764 2563
rect 7845 2557 8540 2563
rect 484 2537 1820 2543
rect 2020 2537 3068 2543
rect 5972 2537 6764 2543
rect 5604 2517 6252 2523
rect 8340 2517 9212 2523
rect 9220 2517 9243 2523
rect 1236 2477 1531 2483
rect 3397 2477 3420 2483
rect 5972 2477 7692 2483
rect 9156 2477 9180 2483
rect 9188 2477 9612 2483
rect 9620 2477 9723 2483
rect 3365 2437 4060 2443
rect 4068 2437 5388 2443
rect 1253 2357 4700 2363
rect 660 2337 667 2343
rect 1812 2337 1900 2343
rect 2868 2337 3500 2343
rect 7877 2337 7964 2343
rect 9277 2325 9283 2336
rect 3172 2317 3820 2323
rect 7333 2317 7340 2323
rect 9605 2317 9900 2323
rect 2180 2297 3340 2303
rect 3348 2297 4620 2303
rect 4628 2297 5356 2303
rect 1876 2277 2907 2283
rect 7076 2277 9276 2283
rect 1332 2257 1723 2263
rect 1733 2257 1740 2263
rect 1764 2257 3084 2263
rect 2788 2237 3580 2243
rect 6788 2237 6812 2243
rect 8932 2237 8956 2243
rect 1797 2197 1804 2203
rect 3109 2197 3132 2203
rect 677 2177 716 2183
rect 6789 2177 6796 2183
rect 1620 2157 1676 2163
rect 2740 2157 3020 2163
rect 7108 2157 9468 2163
rect 4340 2137 4796 2143
rect 7076 2137 8684 2143
rect 4084 2117 4300 2123
rect 5732 2117 6203 2123
rect 6213 2117 6732 2123
rect 2116 2077 2476 2083
rect 2484 2077 2732 2083
rect 2469 2057 2476 2063
rect 8349 1965 8355 1976
rect 948 1957 1004 1963
rect 6132 1957 6139 1963
rect 1733 1937 2220 1943
rect 2660 1937 2828 1943
rect 5716 1917 5851 1923
rect 5861 1917 6636 1923
rect 6644 1917 7260 1923
rect 676 1877 1836 1883
rect 2004 1877 2444 1883
rect 3397 1877 3916 1883
rect 4452 1877 4475 1883
rect 4485 1877 5484 1883
rect 7204 1877 10108 1883
rect 4148 1857 4844 1863
rect 8357 1857 8924 1863
rect 7301 1837 7340 1843
rect 7684 1837 7708 1843
rect 7805 1824 7811 1835
rect 453 1797 1356 1803
rect 2948 1737 4556 1743
rect 9381 1737 9452 1743
rect 532 1717 668 1723
rect 5844 1717 5900 1723
rect 6717 1705 6723 1716
rect 7813 1717 7836 1723
rect 6725 1697 7356 1703
rect 7476 1697 8092 1703
rect 3316 1677 3420 1683
rect 4788 1617 4795 1623
rect 2021 1537 2092 1543
rect 2149 1537 2540 1543
rect 6484 1517 7227 1523
rect 7237 1517 7468 1523
rect 1748 1497 4140 1503
rect 8244 1497 8251 1503
rect 1444 1477 2268 1483
rect 4293 1477 4316 1483
rect 6948 1477 7084 1483
rect 8020 1477 9420 1483
rect 8900 1457 9324 1463
rect 2868 1377 2875 1383
rect 9236 1377 9243 1383
rect 4317 1365 4323 1376
rect 7396 1357 7612 1363
rect 7685 1357 9244 1363
rect 6804 1337 7603 1343
rect 5908 1317 7580 1323
rect 7597 1323 7603 1337
rect 7668 1337 9484 1343
rect 7597 1317 7907 1323
rect 7901 1303 7907 1317
rect 7940 1317 8572 1323
rect 7901 1297 7948 1303
rect 996 1277 1068 1283
rect 6260 1277 6444 1283
rect 7124 1257 7148 1263
rect 4020 1137 4300 1143
rect 6644 1137 9115 1143
rect 9125 1137 9132 1143
rect 8005 1117 8012 1123
rect 692 1097 1356 1103
rect 1572 1097 1772 1103
rect 2852 1097 3420 1103
rect 5812 1097 5916 1103
rect 4692 1077 5404 1083
rect 228 1057 860 1063
rect 3604 1057 3644 1063
rect 1284 1037 1324 1043
rect 244 997 2252 1003
rect 3140 937 3372 943
rect 6404 937 6572 943
rect 7813 917 7980 923
rect 229 797 236 803
rect 6181 737 7020 743
rect 7396 737 7548 743
rect 884 717 1868 723
rect 9445 717 9548 723
rect 7380 697 8812 703
rect 436 677 1084 683
rect 3076 677 3580 683
rect 6020 677 6044 683
rect 7364 677 8044 683
rect 772 657 2044 663
rect 2052 657 3388 663
rect 7796 637 7820 643
rect 996 617 1019 623
rect 6397 565 6403 576
rect 644 557 2972 563
rect 3124 557 4220 563
rect 4868 557 5532 563
rect 1812 537 3180 543
rect 8132 537 8476 543
rect 9477 537 10108 543
rect 4468 517 5019 523
rect 3204 477 3308 483
rect 4660 437 5084 443
rect 5108 357 5180 363
rect 7316 317 8924 323
rect 9733 317 9740 323
rect 7493 297 7500 303
rect 8260 277 8940 283
rect 9972 277 10011 283
rect 1636 257 1836 263
rect 8276 257 8300 263
rect 9844 237 9883 243
rect 8229 177 9164 183
rect 5972 157 7291 163
rect 8020 137 8124 143
rect 7621 117 9516 123
rect 9637 97 10028 103
<< m6contact >>
rect 8411 7515 8421 7525
rect 9787 7515 9797 7525
rect 9915 7515 9925 7525
rect 10011 7495 10021 7505
rect 8443 7475 8453 7485
rect 9147 7475 9157 7485
rect 9947 7475 9957 7485
rect 9595 7435 9605 7445
rect 9307 7384 9317 7385
rect 9307 7376 9308 7384
rect 9308 7376 9316 7384
rect 9316 7376 9317 7384
rect 9307 7375 9317 7376
rect 2843 7275 2853 7285
rect 8859 7115 8869 7125
rect 2683 7095 2693 7105
rect 9531 7035 9541 7045
rect 9435 6984 9445 6985
rect 9435 6976 9436 6984
rect 9436 6976 9444 6984
rect 9444 6976 9445 6984
rect 9435 6975 9445 6976
rect 4219 6904 4229 6905
rect 4219 6896 4220 6904
rect 4220 6896 4228 6904
rect 4228 6896 4229 6904
rect 4219 6895 4229 6896
rect 6203 6895 6213 6905
rect 6683 6895 6693 6905
rect 4827 6735 4837 6745
rect 4475 6715 4485 6725
rect 1115 6695 1125 6705
rect 5787 6655 5797 6665
rect 3995 6635 4005 6645
rect 4411 6644 4421 6645
rect 4411 6636 4412 6644
rect 4412 6636 4420 6644
rect 4420 6636 4421 6644
rect 4411 6635 4421 6636
rect 5755 6635 5765 6645
rect 9115 6644 9125 6645
rect 9115 6636 9116 6644
rect 9116 6636 9124 6644
rect 9124 6636 9125 6644
rect 9115 6635 9125 6636
rect 9467 6644 9477 6645
rect 9467 6636 9468 6644
rect 9468 6636 9476 6644
rect 9476 6636 9477 6644
rect 9467 6635 9477 6636
rect 1115 6575 1125 6585
rect 2843 6575 2853 6585
rect 1947 6515 1957 6525
rect 5755 6495 5765 6505
rect 8443 6455 8453 6465
rect 6139 6435 6149 6445
rect 4187 6375 4197 6385
rect 2395 6364 2405 6365
rect 2395 6356 2396 6364
rect 2396 6356 2404 6364
rect 2404 6356 2405 6364
rect 2395 6355 2405 6356
rect 5787 6315 5797 6325
rect 8443 6275 8453 6285
rect 3355 6255 3365 6265
rect 3995 6255 4005 6265
rect 3963 6244 3973 6245
rect 3963 6236 3964 6244
rect 3964 6236 3972 6244
rect 3972 6236 3973 6244
rect 3963 6235 3973 6236
rect 7931 6235 7941 6245
rect 2843 6144 2853 6145
rect 2843 6136 2844 6144
rect 2844 6136 2852 6144
rect 2852 6136 2853 6144
rect 2843 6135 2853 6136
rect 4795 6135 4805 6145
rect 3995 6115 4005 6125
rect 3099 6095 3109 6105
rect 3355 6095 3365 6105
rect 6715 6095 6725 6105
rect 6683 6075 6693 6085
rect 7611 6075 7621 6085
rect 2203 6055 2213 6065
rect 4411 5935 4421 5945
rect 5499 5875 5509 5885
rect 6139 5875 6149 5885
rect 6459 5844 6469 5845
rect 6459 5836 6460 5844
rect 6460 5836 6468 5844
rect 6468 5836 6469 5844
rect 6459 5835 6469 5836
rect 7355 5844 7365 5845
rect 7355 5836 7356 5844
rect 7356 5836 7364 5844
rect 7364 5836 7365 5844
rect 7355 5835 7365 5836
rect 7739 5815 7749 5825
rect 2779 5795 2789 5805
rect 2395 5755 2405 5765
rect 4827 5755 4837 5765
rect 9723 5735 9733 5745
rect 9883 5735 9893 5745
rect 8539 5695 8549 5705
rect 6683 5675 6693 5685
rect 9755 5675 9765 5685
rect 4923 5635 4933 5645
rect 4699 5555 4709 5565
rect 6139 5564 6149 5565
rect 6139 5556 6140 5564
rect 6140 5556 6148 5564
rect 6148 5556 6149 5564
rect 6139 5555 6149 5556
rect 923 5524 933 5525
rect 923 5516 924 5524
rect 924 5516 932 5524
rect 932 5516 933 5524
rect 923 5515 933 5516
rect 5179 5515 5189 5525
rect 3291 5435 3301 5445
rect 6043 5444 6053 5445
rect 6043 5436 6044 5444
rect 6044 5436 6052 5444
rect 6052 5436 6053 5444
rect 6043 5435 6053 5436
rect 7867 5335 7877 5345
rect 667 5315 677 5325
rect 9723 5315 9733 5325
rect 2395 5275 2405 5285
rect 4571 5275 4581 5285
rect 6363 5284 6373 5285
rect 6363 5276 6364 5284
rect 6364 5276 6372 5284
rect 6372 5276 6373 5284
rect 6363 5275 6373 5276
rect 5083 5235 5093 5245
rect 8251 5195 8261 5205
rect 6203 5135 6213 5145
rect 7323 5135 7333 5145
rect 9755 5115 9765 5125
rect 6459 5095 6469 5105
rect 6907 5075 6917 5085
rect 9627 5084 9637 5085
rect 9627 5076 9628 5084
rect 9628 5076 9636 5084
rect 9636 5076 9637 5084
rect 9627 5075 9637 5076
rect 1531 5055 1541 5065
rect 7131 5035 7141 5045
rect 5499 4935 5509 4945
rect 2843 4915 2853 4925
rect 3867 4895 3877 4905
rect 4219 4895 4229 4905
rect 1115 4875 1125 4885
rect 3579 4875 3589 4885
rect 3835 4875 3845 4885
rect 10011 4864 10021 4865
rect 10011 4856 10012 4864
rect 10012 4856 10020 4864
rect 10020 4856 10021 4864
rect 10011 4855 10021 4856
rect 3291 4835 3301 4845
rect 10011 4835 10021 4845
rect 7611 4824 7621 4825
rect 7611 4816 7612 4824
rect 7612 4816 7620 4824
rect 7620 4816 7621 4824
rect 7611 4815 7621 4816
rect 1243 4784 1253 4785
rect 1243 4776 1244 4784
rect 1244 4776 1252 4784
rect 1252 4776 1253 4784
rect 1243 4775 1253 4776
rect 5499 4715 5509 4725
rect 2203 4675 2213 4685
rect 5723 4684 5733 4685
rect 5723 4676 5724 4684
rect 5724 4676 5732 4684
rect 5732 4676 5733 4684
rect 5723 4675 5733 4676
rect 7227 4675 7237 4685
rect 9115 4675 9125 4685
rect 9691 4684 9701 4685
rect 9691 4676 9692 4684
rect 9692 4676 9700 4684
rect 9700 4676 9701 4684
rect 9691 4675 9701 4676
rect 2459 4655 2469 4665
rect 4475 4664 4485 4665
rect 4475 4656 4476 4664
rect 4476 4656 4484 4664
rect 4484 4656 4485 4664
rect 4475 4655 4485 4656
rect 1147 4644 1157 4645
rect 1147 4636 1148 4644
rect 1148 4636 1156 4644
rect 1156 4636 1157 4644
rect 1147 4635 1157 4636
rect 2331 4635 2341 4645
rect 6683 4644 6693 4645
rect 6683 4636 6684 4644
rect 6684 4636 6692 4644
rect 6692 4636 6693 4644
rect 6683 4635 6693 4636
rect 7963 4635 7973 4645
rect 8219 4644 8229 4645
rect 8219 4636 8220 4644
rect 8220 4636 8228 4644
rect 8228 4636 8229 4644
rect 8219 4635 8229 4636
rect 8763 4635 8773 4645
rect 667 4584 677 4585
rect 667 4576 668 4584
rect 668 4576 676 4584
rect 676 4576 677 4584
rect 667 4575 677 4576
rect 9691 4535 9701 4545
rect 3867 4495 3877 4505
rect 4187 4504 4197 4505
rect 4187 4496 4188 4504
rect 4188 4496 4196 4504
rect 4196 4496 4197 4504
rect 4187 4495 4197 4496
rect 6779 4495 6789 4505
rect 4475 4475 4485 4485
rect 4699 4475 4709 4485
rect 5083 4484 5093 4485
rect 5083 4476 5084 4484
rect 5084 4476 5092 4484
rect 5092 4476 5093 4484
rect 5083 4475 5093 4476
rect 6011 4475 6021 4485
rect 3163 4455 3173 4465
rect 1531 4435 1541 4445
rect 1147 4395 1157 4405
rect 5723 4335 5733 4345
rect 6907 4335 6917 4345
rect 8539 4335 8549 4345
rect 923 4315 933 4325
rect 4827 4315 4837 4325
rect 3931 4295 3941 4305
rect 2779 4275 2789 4285
rect 9691 4275 9701 4285
rect 1019 4264 1029 4265
rect 1019 4256 1020 4264
rect 1020 4256 1028 4264
rect 1028 4256 1029 4264
rect 1019 4255 1029 4256
rect 9115 4255 9125 4265
rect 9147 4255 9157 4265
rect 2139 4244 2149 4245
rect 2139 4236 2140 4244
rect 2140 4236 2148 4244
rect 2148 4236 2149 4244
rect 2139 4235 2149 4236
rect 5979 4235 5989 4245
rect 6747 4244 6757 4245
rect 6747 4236 6748 4244
rect 6748 4236 6756 4244
rect 6756 4236 6757 4244
rect 6747 4235 6757 4236
rect 7675 4235 7685 4245
rect 8923 4244 8933 4245
rect 8923 4236 8924 4244
rect 8924 4236 8932 4244
rect 8932 4236 8933 4244
rect 8923 4235 8933 4236
rect 9147 4244 9157 4245
rect 9147 4236 9148 4244
rect 9148 4236 9156 4244
rect 9156 4236 9157 4244
rect 9147 4235 9157 4236
rect 9371 4235 9381 4245
rect 7131 4204 7141 4205
rect 7131 4196 7132 4204
rect 7132 4196 7140 4204
rect 7140 4196 7141 4204
rect 7131 4195 7141 4196
rect 5147 4175 5157 4185
rect 8859 4184 8869 4185
rect 8859 4176 8860 4184
rect 8860 4176 8868 4184
rect 8868 4176 8869 4184
rect 8859 4175 8869 4176
rect 4891 4135 4901 4145
rect 4923 4135 4933 4145
rect 1115 4115 1125 4125
rect 1115 4095 1125 4105
rect 2395 4115 2405 4125
rect 3387 4115 3397 4125
rect 5435 4115 5445 4125
rect 5755 4124 5765 4125
rect 5755 4116 5756 4124
rect 5756 4116 5764 4124
rect 5764 4116 5765 4124
rect 5755 4115 5765 4116
rect 6203 4115 6213 4125
rect 1211 4095 1221 4105
rect 3547 4095 3557 4105
rect 6363 4095 6373 4105
rect 7355 4095 7365 4105
rect 3963 3935 3973 3945
rect 3995 3915 4005 3925
rect 6715 3915 6725 3925
rect 9275 3915 9285 3925
rect 219 3875 229 3885
rect 1947 3895 1957 3905
rect 1787 3855 1797 3865
rect 5531 3855 5541 3865
rect 8763 3844 8773 3845
rect 8763 3836 8764 3844
rect 8764 3836 8772 3844
rect 8772 3836 8773 3844
rect 8763 3835 8773 3836
rect 9307 3835 9317 3845
rect 7931 3815 7941 3825
rect 5147 3784 5157 3785
rect 5147 3776 5148 3784
rect 5148 3776 5156 3784
rect 5156 3776 5157 3784
rect 5147 3775 5157 3776
rect 3419 3735 3429 3745
rect 3163 3724 3173 3725
rect 3163 3716 3164 3724
rect 3164 3716 3172 3724
rect 3172 3716 3173 3724
rect 3163 3715 3173 3716
rect 6043 3584 6053 3585
rect 6043 3576 6044 3584
rect 6044 3576 6052 3584
rect 6052 3576 6053 3584
rect 6043 3575 6053 3576
rect 6715 3535 6725 3545
rect 7739 3535 7749 3545
rect 8347 3535 8357 3545
rect 9147 3535 9157 3545
rect 3835 3515 3845 3525
rect 9147 3524 9157 3525
rect 9147 3516 9148 3524
rect 9148 3516 9156 3524
rect 9156 3516 9157 3524
rect 9147 3515 9157 3516
rect 9307 3515 9317 3525
rect 9115 3504 9125 3505
rect 9115 3496 9116 3504
rect 9116 3496 9124 3504
rect 9124 3496 9125 3504
rect 9115 3495 9125 3496
rect 3355 3484 3365 3485
rect 3355 3476 3356 3484
rect 3356 3476 3364 3484
rect 3364 3476 3365 3484
rect 3355 3475 3365 3476
rect 3387 3475 3397 3485
rect 4571 3455 4581 3465
rect 2011 3444 2021 3445
rect 2011 3436 2012 3444
rect 2012 3436 2020 3444
rect 2020 3436 2021 3444
rect 2011 3435 2021 3436
rect 5275 3435 5285 3445
rect 5563 3444 5573 3445
rect 7835 3444 7845 3445
rect 5563 3436 5564 3444
rect 5564 3436 5572 3444
rect 5572 3436 5573 3444
rect 7835 3436 7836 3444
rect 7836 3436 7844 3444
rect 7844 3436 7845 3444
rect 5563 3435 5573 3436
rect 7835 3435 7845 3436
rect 443 3384 453 3385
rect 443 3376 444 3384
rect 444 3376 452 3384
rect 452 3376 453 3384
rect 443 3375 453 3376
rect 1243 3384 1253 3385
rect 1243 3376 1244 3384
rect 1244 3376 1252 3384
rect 1252 3376 1253 3384
rect 1243 3375 1253 3376
rect 3931 3375 3941 3385
rect 9947 3375 9957 3385
rect 5179 3364 5189 3365
rect 5179 3356 5180 3364
rect 5180 3356 5188 3364
rect 5188 3356 5189 3364
rect 5179 3355 5189 3356
rect 5531 3355 5541 3365
rect 5563 3355 5573 3365
rect 6779 3355 6789 3365
rect 7963 3355 7973 3365
rect 667 3335 677 3345
rect 6139 3335 6149 3345
rect 4315 3324 4325 3325
rect 4315 3316 4316 3324
rect 4316 3316 4324 3324
rect 4324 3316 4325 3324
rect 4315 3315 4325 3316
rect 4571 3135 4581 3145
rect 6747 3135 6757 3145
rect 1243 3104 1253 3105
rect 1243 3096 1244 3104
rect 1244 3096 1252 3104
rect 1252 3096 1253 3104
rect 1243 3095 1253 3096
rect 2683 3095 2693 3105
rect 2875 3095 2885 3105
rect 5275 3095 5285 3105
rect 5979 3095 5989 3105
rect 2395 3075 2405 3085
rect 3931 3075 3941 3085
rect 5755 3075 5765 3085
rect 6683 3055 6693 3065
rect 7611 3064 7621 3065
rect 7611 3056 7612 3064
rect 7612 3056 7620 3064
rect 7620 3056 7621 3064
rect 7611 3055 7621 3056
rect 5851 3035 5861 3045
rect 5883 3044 5893 3045
rect 5883 3036 5884 3044
rect 5884 3036 5892 3044
rect 5892 3036 5893 3044
rect 5883 3035 5893 3036
rect 1211 2995 1221 3005
rect 8411 2984 8421 2985
rect 8411 2976 8412 2984
rect 8412 2976 8420 2984
rect 8420 2976 8421 2984
rect 8411 2975 8421 2976
rect 6011 2935 6021 2945
rect 2907 2875 2917 2885
rect 9915 2884 9925 2885
rect 9915 2876 9916 2884
rect 9916 2876 9924 2884
rect 9924 2876 9925 2884
rect 9915 2875 9925 2876
rect 9147 2844 9157 2845
rect 9147 2836 9148 2844
rect 9148 2836 9156 2844
rect 9156 2836 9157 2844
rect 9147 2835 9157 2836
rect 4283 2775 4293 2785
rect 6171 2744 6181 2745
rect 6171 2736 6172 2744
rect 6172 2736 6180 2744
rect 6180 2736 6181 2744
rect 6171 2735 6181 2736
rect 7355 2735 7365 2745
rect 2875 2675 2885 2685
rect 3355 2664 3365 2665
rect 3355 2656 3356 2664
rect 3356 2656 3364 2664
rect 3364 2656 3365 2664
rect 3355 2655 3365 2656
rect 4891 2655 4901 2665
rect 8923 2655 8933 2665
rect 3547 2635 3557 2645
rect 667 2595 677 2605
rect 1115 2575 1125 2585
rect 3835 2575 3845 2585
rect 9787 2584 9797 2585
rect 9787 2576 9788 2584
rect 9788 2576 9796 2584
rect 9796 2576 9797 2584
rect 9787 2575 9797 2576
rect 7835 2555 7845 2565
rect 9243 2515 9253 2525
rect 1531 2475 1541 2485
rect 3387 2475 3397 2485
rect 9723 2475 9733 2485
rect 3419 2464 3429 2465
rect 3419 2456 3420 2464
rect 3420 2456 3428 2464
rect 3428 2456 3429 2464
rect 3419 2455 3429 2456
rect 3355 2435 3365 2445
rect 1243 2355 1253 2365
rect 667 2335 677 2345
rect 7867 2335 7877 2345
rect 7323 2315 7333 2325
rect 9275 2315 9285 2325
rect 9595 2315 9605 2325
rect 2907 2275 2917 2285
rect 1723 2255 1733 2265
rect 7995 2264 8005 2265
rect 7995 2256 7996 2264
rect 7996 2256 8004 2264
rect 8004 2256 8005 2264
rect 7995 2255 8005 2256
rect 3579 2224 3589 2225
rect 3579 2216 3580 2224
rect 3580 2216 3588 2224
rect 3588 2216 3589 2224
rect 3579 2215 3589 2216
rect 1787 2195 1797 2205
rect 3099 2195 3109 2205
rect 667 2175 677 2185
rect 5435 2184 5445 2185
rect 5435 2176 5436 2184
rect 5436 2176 5444 2184
rect 5444 2176 5445 2184
rect 5435 2175 5445 2176
rect 6779 2175 6789 2185
rect 8443 2184 8453 2185
rect 8443 2176 8444 2184
rect 8444 2176 8452 2184
rect 8452 2176 8453 2184
rect 8443 2175 8453 2176
rect 5883 2144 5893 2145
rect 5883 2136 5884 2144
rect 5884 2136 5892 2144
rect 5892 2136 5893 2144
rect 5883 2135 5893 2136
rect 6203 2115 6213 2125
rect 5755 2104 5765 2105
rect 5755 2096 5756 2104
rect 5756 2096 5764 2104
rect 5764 2096 5765 2104
rect 5755 2095 5765 2096
rect 7483 2104 7493 2105
rect 7483 2096 7484 2104
rect 7484 2096 7492 2104
rect 7492 2096 7493 2104
rect 7483 2095 7493 2096
rect 2459 2055 2469 2065
rect 3931 2064 3941 2065
rect 3931 2056 3932 2064
rect 3932 2056 3940 2064
rect 3940 2056 3941 2064
rect 3931 2055 3941 2056
rect 6139 1955 6149 1965
rect 8347 1955 8357 1965
rect 1723 1935 1733 1945
rect 5851 1915 5861 1925
rect 3387 1875 3397 1885
rect 4475 1875 4485 1885
rect 8347 1855 8357 1865
rect 6395 1844 6405 1845
rect 6395 1836 6396 1844
rect 6396 1836 6404 1844
rect 6404 1836 6405 1844
rect 6395 1835 6405 1836
rect 7291 1835 7301 1845
rect 7803 1835 7813 1845
rect 9307 1844 9317 1845
rect 9307 1836 9308 1844
rect 9308 1836 9316 1844
rect 9316 1836 9317 1844
rect 9307 1835 9317 1836
rect 2331 1824 2341 1825
rect 2331 1816 2332 1824
rect 2332 1816 2340 1824
rect 2340 1816 2341 1824
rect 2331 1815 2341 1816
rect 443 1795 453 1805
rect 9531 1784 9541 1785
rect 9531 1776 9532 1784
rect 9532 1776 9540 1784
rect 9540 1776 9541 1784
rect 9531 1775 9541 1776
rect 9371 1735 9381 1745
rect 7803 1715 7813 1725
rect 6715 1695 6725 1705
rect 4795 1615 4805 1625
rect 2011 1535 2021 1545
rect 2139 1535 2149 1545
rect 9307 1544 9317 1545
rect 9307 1536 9308 1544
rect 9308 1536 9316 1544
rect 9316 1536 9317 1544
rect 9307 1535 9317 1536
rect 7227 1515 7237 1525
rect 8251 1495 8261 1505
rect 4283 1475 4293 1485
rect 2875 1375 2885 1385
rect 9243 1375 9253 1385
rect 4315 1355 4325 1365
rect 7675 1355 7685 1365
rect 1531 1184 1541 1185
rect 1531 1176 1532 1184
rect 1532 1176 1540 1184
rect 1540 1176 1541 1184
rect 1531 1175 1541 1176
rect 9115 1135 9125 1145
rect 7995 1115 8005 1125
rect 7803 1044 7813 1045
rect 7803 1036 7804 1044
rect 7804 1036 7812 1044
rect 7812 1036 7813 1044
rect 7803 1035 7813 1036
rect 7803 915 7813 925
rect 5019 904 5029 905
rect 5019 896 5020 904
rect 5020 896 5028 904
rect 5028 896 5029 904
rect 5019 895 5029 896
rect 219 795 229 805
rect 6171 735 6181 745
rect 9435 715 9445 725
rect 1019 615 1029 625
rect 5755 584 5765 585
rect 5755 576 5756 584
rect 5756 576 5764 584
rect 5764 576 5765 584
rect 5755 575 5765 576
rect 6395 555 6405 565
rect 9467 535 9477 545
rect 5019 515 5029 525
rect 9723 315 9733 325
rect 7483 295 7493 305
rect 10011 275 10021 285
rect 9883 235 9893 245
rect 8219 175 8229 185
rect 7291 155 7301 165
rect 7611 115 7621 125
rect 9627 95 9637 105
<< metal6 >>
rect 1115 6585 1125 6695
rect 667 4585 677 5315
rect 923 4325 933 5515
rect 219 805 229 3875
rect 443 1805 453 3375
rect 667 2605 677 3335
rect 667 2185 677 2335
rect 1019 625 1029 4255
rect 1115 4125 1125 4875
rect 1147 4405 1157 4635
rect 1115 2585 1125 4095
rect 1211 3005 1221 4095
rect 1243 3385 1253 4775
rect 1531 4445 1541 5055
rect 1947 3905 1957 6515
rect 2203 4685 2213 6055
rect 2395 5765 2405 6355
rect 1243 2365 1253 3095
rect 1531 1185 1541 2475
rect 1723 1945 1733 2255
rect 1787 2205 1797 3855
rect 2011 1545 2021 3435
rect 2139 1545 2149 4235
rect 2331 1825 2341 4635
rect 2395 4125 2405 5275
rect 2395 3085 2405 4115
rect 2459 2065 2469 4655
rect 2683 3105 2693 7095
rect 2843 6585 2853 7275
rect 3995 6265 4005 6635
rect 2779 4285 2789 5795
rect 2843 4925 2853 6135
rect 3355 6105 3365 6255
rect 2875 2685 2885 3095
rect 2875 1385 2885 2675
rect 2907 2285 2917 2875
rect 3099 2205 3109 6095
rect 3291 4845 3301 5435
rect 3163 3725 3173 4455
rect 3355 3485 3365 6095
rect 3387 3485 3397 4115
rect 3355 2445 3365 2655
rect 3387 1885 3397 2475
rect 3419 2465 3429 3735
rect 3547 2645 3557 4095
rect 3579 2225 3589 4875
rect 3835 3525 3845 4875
rect 3867 4505 3877 4895
rect 3835 2585 3845 3515
rect 3931 3385 3941 4295
rect 3963 3945 3973 6235
rect 3995 3925 4005 6115
rect 4187 4505 4197 6375
rect 4219 4905 4229 6895
rect 4411 5945 4421 6635
rect 4475 4665 4485 6715
rect 3931 2065 3941 3075
rect 4283 1485 4293 2775
rect 4315 1365 4325 3315
rect 4475 1885 4485 4475
rect 4571 3465 4581 5275
rect 4699 4485 4709 5555
rect 4571 3145 4581 3455
rect 4795 1625 4805 6135
rect 4827 5765 4837 6735
rect 5755 6505 5765 6635
rect 5787 6325 5797 6655
rect 6139 5885 6149 6435
rect 4827 4325 4837 5755
rect 4923 4145 4933 5635
rect 5083 4485 5093 5235
rect 4891 2665 4901 4135
rect 5147 3785 5157 4175
rect 5179 3365 5189 5515
rect 5499 4945 5509 5875
rect 6139 5565 6149 5875
rect 5499 4725 5509 4935
rect 5723 4345 5733 4675
rect 5275 3105 5285 3435
rect 5435 2185 5445 4115
rect 5531 3365 5541 3855
rect 5563 3365 5573 3435
rect 5755 3085 5765 4115
rect 5979 3105 5989 4235
rect 5019 525 5029 895
rect 5755 585 5765 2095
rect 5851 1925 5861 3035
rect 5883 2145 5893 3035
rect 6011 2945 6021 4475
rect 6043 3585 6053 5435
rect 6203 5145 6213 6895
rect 6683 6085 6693 6895
rect 6139 1965 6149 3335
rect 6171 745 6181 2735
rect 6203 2125 6213 4115
rect 6363 4105 6373 5275
rect 6459 5105 6469 5835
rect 6683 5685 6693 6075
rect 6683 3065 6693 4635
rect 6715 3925 6725 6095
rect 6395 565 6405 1835
rect 6715 1705 6725 3535
rect 6747 3145 6757 4235
rect 6779 3365 6789 4495
rect 6907 4345 6917 5075
rect 7131 4205 7141 5035
rect 6779 2185 6789 3355
rect 7227 1525 7237 4675
rect 7323 2325 7333 5135
rect 7355 4105 7365 5835
rect 7611 4825 7621 6075
rect 7355 2745 7365 4095
rect 7291 165 7301 1835
rect 7483 305 7493 2095
rect 7611 125 7621 3055
rect 7675 1365 7685 4235
rect 7739 3545 7749 5815
rect 7835 2565 7845 3435
rect 7867 2345 7877 5335
rect 7931 3825 7941 6235
rect 7963 3365 7973 4635
rect 7803 1725 7813 1835
rect 7995 1125 8005 2255
rect 7803 925 7813 1035
rect 8219 185 8229 4635
rect 8251 1505 8261 5195
rect 8347 1965 8357 3535
rect 8411 2985 8421 7515
rect 8443 6465 8453 7475
rect 8443 2185 8453 6275
rect 8539 4345 8549 5695
rect 8763 3845 8773 4635
rect 8859 4185 8869 7115
rect 9115 4685 9125 6635
rect 9115 4265 9125 4675
rect 9147 4265 9157 7475
rect 8923 2665 8933 4235
rect 9147 3545 9157 4235
rect 8347 1865 8357 1955
rect 9115 1145 9125 3495
rect 9147 2845 9157 3515
rect 9243 1385 9253 2515
rect 9275 2325 9285 3915
rect 9307 3845 9317 7375
rect 9307 3525 9317 3835
rect 9307 1545 9317 1835
rect 9371 1745 9381 4235
rect 9435 725 9445 6975
rect 9467 545 9477 6635
rect 9531 1785 9541 7035
rect 9595 2325 9605 7435
rect 9723 5325 9733 5735
rect 9755 5125 9765 5675
rect 9627 105 9637 5075
rect 9691 4545 9701 4675
rect 9691 4285 9701 4535
rect 9787 2585 9797 7515
rect 9723 325 9733 2475
rect 9883 245 9893 5735
rect 9915 2885 9925 7515
rect 9947 3385 9957 7475
rect 10011 4865 10021 7495
rect 10011 285 10021 4835
use FILL  FILL_38_12
timestamp 1612251222
transform 1 0 10246 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_11
timestamp 1612251222
transform 1 0 10230 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_10
timestamp 1612251222
transform 1 0 10214 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_9
timestamp 1612251222
transform 1 0 10198 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_8
timestamp 1612251222
transform 1 0 10182 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_7
timestamp 1612251222
transform 1 0 10166 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_6
timestamp 1612251222
transform 1 0 10150 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_5
timestamp 1612251222
transform 1 0 10134 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_4
timestamp 1612251222
transform 1 0 10118 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_3
timestamp 1612251222
transform 1 0 10102 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_2
timestamp 1612251222
transform 1 0 10086 0 1 7410
box -4 -6 20 206
use FILL  FILL_38_1
timestamp 1612251222
transform 1 0 10070 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_192
timestamp 1612251222
transform 1 0 9904 0 1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_192
timestamp 1612251222
transform 1 0 9888 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_192
timestamp 1612251222
transform 1 0 9872 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_192
timestamp 1612251222
transform 1 0 9856 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_567
timestamp 1612251222
transform 1 0 9690 0 1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_567
timestamp 1612251222
transform 1 0 9674 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_567
timestamp 1612251222
transform 1 0 9658 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_567
timestamp 1612251222
transform 1 0 9642 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_566
timestamp 1612251222
transform 1 0 9476 0 1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_566
timestamp 1612251222
transform 1 0 9460 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_566
timestamp 1612251222
transform 1 0 9444 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_566
timestamp 1612251222
transform 1 0 9428 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_854
timestamp 1612251222
transform 1 0 9262 0 1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_854
timestamp 1612251222
transform 1 0 9246 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_854
timestamp 1612251222
transform 1 0 9230 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_854
timestamp 1612251222
transform 1 0 9214 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_776
timestamp 1612251222
transform -1 0 9214 0 1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_776
timestamp 1612251222
transform -1 0 9048 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_776
timestamp 1612251222
transform -1 0 9032 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_776
timestamp 1612251222
transform -1 0 9016 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_223
timestamp 1612251222
transform 1 0 8834 0 1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_223
timestamp 1612251222
transform 1 0 8818 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_223
timestamp 1612251222
transform 1 0 8802 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_223
timestamp 1612251222
transform 1 0 8786 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_221
timestamp 1612251222
transform -1 0 8786 0 1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_221
timestamp 1612251222
transform -1 0 8620 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_221
timestamp 1612251222
transform -1 0 8604 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_221
timestamp 1612251222
transform -1 0 8588 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_742
timestamp 1612251222
transform 1 0 8406 0 1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_742
timestamp 1612251222
transform 1 0 8390 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_742
timestamp 1612251222
transform 1 0 8374 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_742
timestamp 1612251222
transform 1 0 8358 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_331
timestamp 1612251222
transform 1 0 8192 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_331
timestamp 1612251222
transform 1 0 8176 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_331
timestamp 1612251222
transform 1 0 8160 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_331
timestamp 1612251222
transform 1 0 8144 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_331
timestamp 1612251222
transform 1 0 8128 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_838
timestamp 1612251222
transform 1 0 7962 0 1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_838
timestamp 1612251222
transform 1 0 7946 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_838
timestamp 1612251222
transform 1 0 7930 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_838
timestamp 1612251222
transform 1 0 7914 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_837
timestamp 1612251222
transform 1 0 7748 0 1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_837
timestamp 1612251222
transform 1 0 7732 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_837
timestamp 1612251222
transform 1 0 7716 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_837
timestamp 1612251222
transform 1 0 7700 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_419
timestamp 1612251222
transform 1 0 7534 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_419
timestamp 1612251222
transform 1 0 7518 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_419
timestamp 1612251222
transform 1 0 7502 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_419
timestamp 1612251222
transform 1 0 7486 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_419
timestamp 1612251222
transform 1 0 7470 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_295
timestamp 1612251222
transform -1 0 7470 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_295
timestamp 1612251222
transform -1 0 7304 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_295
timestamp 1612251222
transform -1 0 7288 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_295
timestamp 1612251222
transform -1 0 7272 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_295
timestamp 1612251222
transform -1 0 7256 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_505
timestamp 1612251222
transform 1 0 7074 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_505
timestamp 1612251222
transform 1 0 7058 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_505
timestamp 1612251222
transform 1 0 7042 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_505
timestamp 1612251222
transform 1 0 7026 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_505
timestamp 1612251222
transform 1 0 7010 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_825
timestamp 1612251222
transform 1 0 6844 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_825
timestamp 1612251222
transform 1 0 6828 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_825
timestamp 1612251222
transform 1 0 6812 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_825
timestamp 1612251222
transform 1 0 6796 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_825
timestamp 1612251222
transform 1 0 6780 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_347
timestamp 1612251222
transform 1 0 6614 0 1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_347
timestamp 1612251222
transform 1 0 6598 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_347
timestamp 1612251222
transform 1 0 6582 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_347
timestamp 1612251222
transform 1 0 6566 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_69
timestamp 1612251222
transform 1 0 6400 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_69
timestamp 1612251222
transform 1 0 6384 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_69
timestamp 1612251222
transform 1 0 6368 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_69
timestamp 1612251222
transform 1 0 6352 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_69
timestamp 1612251222
transform 1 0 6336 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_68
timestamp 1612251222
transform 1 0 6170 0 1 7410
box -4 -6 170 206
use FILL  FILL2_POR2X1_68
timestamp 1612251222
transform 1 0 6154 0 1 7410
box -4 -6 20 206
use FILL  FILL1_POR2X1_68
timestamp 1612251222
transform 1 0 6138 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_68
timestamp 1612251222
transform 1 0 6122 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_68
timestamp 1612251222
transform 1 0 6106 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_297
timestamp 1612251222
transform 1 0 5940 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_297
timestamp 1612251222
transform 1 0 5924 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_297
timestamp 1612251222
transform 1 0 5908 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_297
timestamp 1612251222
transform 1 0 5892 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_297
timestamp 1612251222
transform 1 0 5876 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_296
timestamp 1612251222
transform -1 0 5876 0 1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_296
timestamp 1612251222
transform -1 0 5710 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_296
timestamp 1612251222
transform -1 0 5694 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_296
timestamp 1612251222
transform -1 0 5678 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_401
timestamp 1612251222
transform 1 0 5496 0 1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_401
timestamp 1612251222
transform 1 0 5480 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_401
timestamp 1612251222
transform 1 0 5464 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_401
timestamp 1612251222
transform 1 0 5448 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_396
timestamp 1612251222
transform 1 0 5282 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_396
timestamp 1612251222
transform 1 0 5266 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_396
timestamp 1612251222
transform 1 0 5250 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_396
timestamp 1612251222
transform 1 0 5234 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_396
timestamp 1612251222
transform 1 0 5218 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_33
timestamp 1612251222
transform 1 0 5052 0 1 7410
box -4 -6 170 206
use FILL  FILL2_POR2X1_33
timestamp 1612251222
transform 1 0 5036 0 1 7410
box -4 -6 20 206
use FILL  FILL1_POR2X1_33
timestamp 1612251222
transform 1 0 5020 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_33
timestamp 1612251222
transform 1 0 5004 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_33
timestamp 1612251222
transform 1 0 4988 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_20
timestamp 1612251222
transform 1 0 4822 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_20
timestamp 1612251222
transform 1 0 4806 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_20
timestamp 1612251222
transform 1 0 4790 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_20
timestamp 1612251222
transform 1 0 4774 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_20
timestamp 1612251222
transform 1 0 4758 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_19
timestamp 1612251222
transform 1 0 4592 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_19
timestamp 1612251222
transform 1 0 4576 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_19
timestamp 1612251222
transform 1 0 4560 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_19
timestamp 1612251222
transform 1 0 4544 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_19
timestamp 1612251222
transform 1 0 4528 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_5
timestamp 1612251222
transform 1 0 4362 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_5
timestamp 1612251222
transform 1 0 4346 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_5
timestamp 1612251222
transform 1 0 4330 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_5
timestamp 1612251222
transform 1 0 4314 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_5
timestamp 1612251222
transform 1 0 4298 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_612
timestamp 1612251222
transform -1 0 4298 0 1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_612
timestamp 1612251222
transform -1 0 4132 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_612
timestamp 1612251222
transform -1 0 4116 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_612
timestamp 1612251222
transform -1 0 4100 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_414
timestamp 1612251222
transform 1 0 3918 0 1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_414
timestamp 1612251222
transform 1 0 3902 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_414
timestamp 1612251222
transform 1 0 3886 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_414
timestamp 1612251222
transform 1 0 3870 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_4
timestamp 1612251222
transform 1 0 3704 0 1 7410
box -4 -6 170 206
use FILL  FILL2_POR2X1_4
timestamp 1612251222
transform 1 0 3688 0 1 7410
box -4 -6 20 206
use FILL  FILL1_POR2X1_4
timestamp 1612251222
transform 1 0 3672 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_4
timestamp 1612251222
transform 1 0 3656 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_4
timestamp 1612251222
transform 1 0 3640 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_5
timestamp 1612251222
transform -1 0 3640 0 1 7410
box -4 -6 170 206
use FILL  FILL2_POR2X1_5
timestamp 1612251222
transform -1 0 3474 0 1 7410
box -4 -6 20 206
use FILL  FILL1_POR2X1_5
timestamp 1612251222
transform -1 0 3458 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_5
timestamp 1612251222
transform -1 0 3442 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_5
timestamp 1612251222
transform -1 0 3426 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_37
timestamp 1612251222
transform -1 0 3410 0 1 7410
box -4 -6 170 206
use FILL  FILL2_POR2X1_37
timestamp 1612251222
transform -1 0 3244 0 1 7410
box -4 -6 20 206
use FILL  FILL1_POR2X1_37
timestamp 1612251222
transform -1 0 3228 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_37
timestamp 1612251222
transform -1 0 3212 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_37
timestamp 1612251222
transform -1 0 3196 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_461
timestamp 1612251222
transform 1 0 3014 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_461
timestamp 1612251222
transform 1 0 2998 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_461
timestamp 1612251222
transform 1 0 2982 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_461
timestamp 1612251222
transform 1 0 2966 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_461
timestamp 1612251222
transform 1 0 2950 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_413
timestamp 1612251222
transform 1 0 2784 0 1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_413
timestamp 1612251222
transform 1 0 2768 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_413
timestamp 1612251222
transform 1 0 2752 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_413
timestamp 1612251222
transform 1 0 2736 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_607
timestamp 1612251222
transform -1 0 2736 0 1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_607
timestamp 1612251222
transform -1 0 2570 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_607
timestamp 1612251222
transform -1 0 2554 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_607
timestamp 1612251222
transform -1 0 2538 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_646
timestamp 1612251222
transform -1 0 2522 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_646
timestamp 1612251222
transform -1 0 2356 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_646
timestamp 1612251222
transform -1 0 2340 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_646
timestamp 1612251222
transform -1 0 2324 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_646
timestamp 1612251222
transform -1 0 2308 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_647
timestamp 1612251222
transform -1 0 2292 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_647
timestamp 1612251222
transform -1 0 2126 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_647
timestamp 1612251222
transform -1 0 2110 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_647
timestamp 1612251222
transform -1 0 2094 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_647
timestamp 1612251222
transform -1 0 2078 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_656
timestamp 1612251222
transform -1 0 2062 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_656
timestamp 1612251222
transform -1 0 1896 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_656
timestamp 1612251222
transform -1 0 1880 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_656
timestamp 1612251222
transform -1 0 1864 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_656
timestamp 1612251222
transform -1 0 1848 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_663
timestamp 1612251222
transform 1 0 1666 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_663
timestamp 1612251222
transform 1 0 1650 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_663
timestamp 1612251222
transform 1 0 1634 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_663
timestamp 1612251222
transform 1 0 1618 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_663
timestamp 1612251222
transform 1 0 1602 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_662
timestamp 1612251222
transform 1 0 1436 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_662
timestamp 1612251222
transform 1 0 1420 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_662
timestamp 1612251222
transform 1 0 1404 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_662
timestamp 1612251222
transform 1 0 1388 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_662
timestamp 1612251222
transform 1 0 1372 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_660
timestamp 1612251222
transform 1 0 1206 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_660
timestamp 1612251222
transform 1 0 1190 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_660
timestamp 1612251222
transform 1 0 1174 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_660
timestamp 1612251222
transform 1 0 1158 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_660
timestamp 1612251222
transform 1 0 1142 0 1 7410
box -4 -6 20 206
use POR2X1  POR2X1_690
timestamp 1612251222
transform -1 0 1142 0 1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_690
timestamp 1612251222
transform -1 0 976 0 1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_690
timestamp 1612251222
transform -1 0 960 0 1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_690
timestamp 1612251222
transform -1 0 944 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_691
timestamp 1612251222
transform -1 0 928 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_691
timestamp 1612251222
transform -1 0 762 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_691
timestamp 1612251222
transform -1 0 746 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_691
timestamp 1612251222
transform -1 0 730 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_691
timestamp 1612251222
transform -1 0 714 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_655
timestamp 1612251222
transform 1 0 532 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_655
timestamp 1612251222
transform 1 0 516 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_655
timestamp 1612251222
transform 1 0 500 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_655
timestamp 1612251222
transform 1 0 484 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_655
timestamp 1612251222
transform 1 0 468 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_648
timestamp 1612251222
transform 1 0 302 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_648
timestamp 1612251222
transform 1 0 286 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_648
timestamp 1612251222
transform 1 0 270 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_648
timestamp 1612251222
transform 1 0 254 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_648
timestamp 1612251222
transform 1 0 238 0 1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_602
timestamp 1612251222
transform 1 0 72 0 1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_602
timestamp 1612251222
transform 1 0 56 0 1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_602
timestamp 1612251222
transform 1 0 40 0 1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_602
timestamp 1612251222
transform 1 0 24 0 1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_602
timestamp 1612251222
transform 1 0 8 0 1 7410
box -4 -6 20 206
use FILL  FILL_37_12
timestamp 1612251222
transform -1 0 10262 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_11
timestamp 1612251222
transform -1 0 10246 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_10
timestamp 1612251222
transform -1 0 10230 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_9
timestamp 1612251222
transform -1 0 10214 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_8
timestamp 1612251222
transform -1 0 10198 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_7
timestamp 1612251222
transform -1 0 10182 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_6
timestamp 1612251222
transform -1 0 10166 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_5
timestamp 1612251222
transform -1 0 10150 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_4
timestamp 1612251222
transform -1 0 10134 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_3
timestamp 1612251222
transform -1 0 10118 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_2
timestamp 1612251222
transform -1 0 10102 0 -1 7410
box -4 -6 20 206
use FILL  FILL_37_1
timestamp 1612251222
transform -1 0 10086 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_580
timestamp 1612251222
transform 1 0 9904 0 -1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_580
timestamp 1612251222
transform 1 0 9888 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_580
timestamp 1612251222
transform 1 0 9872 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_580
timestamp 1612251222
transform 1 0 9856 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_171
timestamp 1612251222
transform 1 0 9690 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_171
timestamp 1612251222
transform 1 0 9674 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_171
timestamp 1612251222
transform 1 0 9658 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_171
timestamp 1612251222
transform 1 0 9642 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_171
timestamp 1612251222
transform 1 0 9626 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_355
timestamp 1612251222
transform -1 0 9626 0 -1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_355
timestamp 1612251222
transform -1 0 9460 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_355
timestamp 1612251222
transform -1 0 9444 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_355
timestamp 1612251222
transform -1 0 9428 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_507
timestamp 1612251222
transform 1 0 9246 0 -1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_507
timestamp 1612251222
transform 1 0 9230 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_507
timestamp 1612251222
transform 1 0 9214 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_507
timestamp 1612251222
transform 1 0 9198 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_504
timestamp 1612251222
transform 1 0 9032 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_504
timestamp 1612251222
transform 1 0 9016 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_504
timestamp 1612251222
transform 1 0 9000 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_504
timestamp 1612251222
transform 1 0 8984 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_504
timestamp 1612251222
transform 1 0 8968 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_481
timestamp 1612251222
transform 1 0 8802 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_481
timestamp 1612251222
transform 1 0 8786 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_481
timestamp 1612251222
transform 1 0 8770 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_481
timestamp 1612251222
transform 1 0 8754 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_481
timestamp 1612251222
transform 1 0 8738 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_294
timestamp 1612251222
transform 1 0 8572 0 -1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_294
timestamp 1612251222
transform 1 0 8556 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_294
timestamp 1612251222
transform 1 0 8540 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_294
timestamp 1612251222
transform 1 0 8524 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_827
timestamp 1612251222
transform -1 0 8524 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_827
timestamp 1612251222
transform -1 0 8358 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_827
timestamp 1612251222
transform -1 0 8342 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_827
timestamp 1612251222
transform -1 0 8326 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_827
timestamp 1612251222
transform -1 0 8310 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_67
timestamp 1612251222
transform -1 0 8294 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_67
timestamp 1612251222
transform -1 0 8128 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_67
timestamp 1612251222
transform -1 0 8112 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_67
timestamp 1612251222
transform -1 0 8096 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_67
timestamp 1612251222
transform -1 0 8080 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_826
timestamp 1612251222
transform -1 0 8064 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_826
timestamp 1612251222
transform -1 0 7898 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_826
timestamp 1612251222
transform -1 0 7882 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_826
timestamp 1612251222
transform -1 0 7866 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_826
timestamp 1612251222
transform -1 0 7850 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_202
timestamp 1612251222
transform -1 0 7834 0 -1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_202
timestamp 1612251222
transform -1 0 7668 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_202
timestamp 1612251222
transform -1 0 7652 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_202
timestamp 1612251222
transform -1 0 7636 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_58
timestamp 1612251222
transform 1 0 7454 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_58
timestamp 1612251222
transform 1 0 7438 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_58
timestamp 1612251222
transform 1 0 7422 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_58
timestamp 1612251222
transform 1 0 7406 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_58
timestamp 1612251222
transform 1 0 7390 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_346
timestamp 1612251222
transform -1 0 7390 0 -1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_346
timestamp 1612251222
transform -1 0 7224 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_346
timestamp 1612251222
transform -1 0 7208 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_346
timestamp 1612251222
transform -1 0 7192 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_402
timestamp 1612251222
transform 1 0 7010 0 -1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_402
timestamp 1612251222
transform 1 0 6994 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_402
timestamp 1612251222
transform 1 0 6978 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_402
timestamp 1612251222
transform 1 0 6962 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_96
timestamp 1612251222
transform 1 0 6796 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_96
timestamp 1612251222
transform 1 0 6780 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_96
timestamp 1612251222
transform 1 0 6764 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_96
timestamp 1612251222
transform 1 0 6748 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_96
timestamp 1612251222
transform 1 0 6732 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_94
timestamp 1612251222
transform 1 0 6566 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_94
timestamp 1612251222
transform 1 0 6550 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_94
timestamp 1612251222
transform 1 0 6534 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_94
timestamp 1612251222
transform 1 0 6518 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_94
timestamp 1612251222
transform 1 0 6502 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_55
timestamp 1612251222
transform 1 0 6336 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_55
timestamp 1612251222
transform 1 0 6320 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_55
timestamp 1612251222
transform 1 0 6304 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_55
timestamp 1612251222
transform 1 0 6288 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_55
timestamp 1612251222
transform 1 0 6272 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_293
timestamp 1612251222
transform 1 0 6106 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_293
timestamp 1612251222
transform 1 0 6090 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_293
timestamp 1612251222
transform 1 0 6074 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_293
timestamp 1612251222
transform 1 0 6058 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_293
timestamp 1612251222
transform 1 0 6042 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_23
timestamp 1612251222
transform 1 0 5876 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_23
timestamp 1612251222
transform 1 0 5860 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_23
timestamp 1612251222
transform 1 0 5844 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_23
timestamp 1612251222
transform 1 0 5828 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_23
timestamp 1612251222
transform 1 0 5812 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_395
timestamp 1612251222
transform -1 0 5812 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_395
timestamp 1612251222
transform -1 0 5646 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_395
timestamp 1612251222
transform -1 0 5630 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_395
timestamp 1612251222
transform -1 0 5614 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_395
timestamp 1612251222
transform -1 0 5598 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_54
timestamp 1612251222
transform -1 0 5582 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_POR2X1_54
timestamp 1612251222
transform -1 0 5416 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_POR2X1_54
timestamp 1612251222
transform -1 0 5400 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_54
timestamp 1612251222
transform -1 0 5384 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_54
timestamp 1612251222
transform -1 0 5368 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_24
timestamp 1612251222
transform -1 0 5352 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_24
timestamp 1612251222
transform -1 0 5186 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_24
timestamp 1612251222
transform -1 0 5170 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_24
timestamp 1612251222
transform -1 0 5154 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_24
timestamp 1612251222
transform -1 0 5138 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_14
timestamp 1612251222
transform 1 0 4956 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_14
timestamp 1612251222
transform 1 0 4940 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_14
timestamp 1612251222
transform 1 0 4924 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_14
timestamp 1612251222
transform 1 0 4908 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_14
timestamp 1612251222
transform 1 0 4892 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_293
timestamp 1612251222
transform -1 0 4892 0 -1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_293
timestamp 1612251222
transform -1 0 4726 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_293
timestamp 1612251222
transform -1 0 4710 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_293
timestamp 1612251222
transform -1 0 4694 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_611
timestamp 1612251222
transform -1 0 4678 0 -1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_611
timestamp 1612251222
transform -1 0 4512 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_611
timestamp 1612251222
transform -1 0 4496 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_611
timestamp 1612251222
transform -1 0 4480 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_610
timestamp 1612251222
transform -1 0 4464 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_610
timestamp 1612251222
transform -1 0 4298 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_610
timestamp 1612251222
transform -1 0 4282 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_610
timestamp 1612251222
transform -1 0 4266 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_610
timestamp 1612251222
transform -1 0 4250 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_415
timestamp 1612251222
transform -1 0 4234 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_415
timestamp 1612251222
transform -1 0 4068 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_415
timestamp 1612251222
transform -1 0 4052 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_415
timestamp 1612251222
transform -1 0 4036 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_415
timestamp 1612251222
transform -1 0 4020 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_416
timestamp 1612251222
transform -1 0 4004 0 -1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_416
timestamp 1612251222
transform -1 0 3838 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_416
timestamp 1612251222
transform -1 0 3822 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_416
timestamp 1612251222
transform -1 0 3806 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_462
timestamp 1612251222
transform 1 0 3624 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_462
timestamp 1612251222
transform 1 0 3608 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_462
timestamp 1612251222
transform 1 0 3592 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_462
timestamp 1612251222
transform 1 0 3576 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_462
timestamp 1612251222
transform 1 0 3560 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_232
timestamp 1612251222
transform -1 0 3560 0 -1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_232
timestamp 1612251222
transform -1 0 3394 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_232
timestamp 1612251222
transform -1 0 3378 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_232
timestamp 1612251222
transform -1 0 3362 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_606
timestamp 1612251222
transform -1 0 3346 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_606
timestamp 1612251222
transform -1 0 3180 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_606
timestamp 1612251222
transform -1 0 3164 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_606
timestamp 1612251222
transform -1 0 3148 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_606
timestamp 1612251222
transform -1 0 3132 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_411
timestamp 1612251222
transform -1 0 3116 0 -1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_411
timestamp 1612251222
transform -1 0 2950 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_411
timestamp 1612251222
transform -1 0 2934 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_411
timestamp 1612251222
transform -1 0 2918 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_634
timestamp 1612251222
transform 1 0 2736 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_634
timestamp 1612251222
transform 1 0 2720 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_634
timestamp 1612251222
transform 1 0 2704 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_634
timestamp 1612251222
transform 1 0 2688 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_634
timestamp 1612251222
transform 1 0 2672 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_412
timestamp 1612251222
transform -1 0 2672 0 -1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_412
timestamp 1612251222
transform -1 0 2506 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_412
timestamp 1612251222
transform -1 0 2490 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_412
timestamp 1612251222
transform -1 0 2474 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_642
timestamp 1612251222
transform -1 0 2458 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_642
timestamp 1612251222
transform -1 0 2292 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_642
timestamp 1612251222
transform -1 0 2276 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_642
timestamp 1612251222
transform -1 0 2260 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_642
timestamp 1612251222
transform -1 0 2244 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_400
timestamp 1612251222
transform 1 0 2062 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_400
timestamp 1612251222
transform 1 0 2046 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_400
timestamp 1612251222
transform 1 0 2030 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_400
timestamp 1612251222
transform 1 0 2014 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_400
timestamp 1612251222
transform 1 0 1998 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_394
timestamp 1612251222
transform 1 0 1832 0 -1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_394
timestamp 1612251222
transform 1 0 1816 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_394
timestamp 1612251222
transform 1 0 1800 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_394
timestamp 1612251222
transform 1 0 1784 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_393
timestamp 1612251222
transform 1 0 1618 0 -1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_393
timestamp 1612251222
transform 1 0 1602 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_393
timestamp 1612251222
transform 1 0 1586 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_393
timestamp 1612251222
transform 1 0 1570 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_688
timestamp 1612251222
transform -1 0 1570 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_688
timestamp 1612251222
transform -1 0 1404 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_688
timestamp 1612251222
transform -1 0 1388 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_688
timestamp 1612251222
transform -1 0 1372 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_688
timestamp 1612251222
transform -1 0 1356 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_590
timestamp 1612251222
transform -1 0 1340 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_590
timestamp 1612251222
transform -1 0 1174 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_590
timestamp 1612251222
transform -1 0 1158 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_590
timestamp 1612251222
transform -1 0 1142 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_590
timestamp 1612251222
transform -1 0 1126 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_689
timestamp 1612251222
transform -1 0 1110 0 -1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_689
timestamp 1612251222
transform -1 0 944 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_689
timestamp 1612251222
transform -1 0 928 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_689
timestamp 1612251222
transform -1 0 912 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_649
timestamp 1612251222
transform -1 0 896 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_649
timestamp 1612251222
transform -1 0 730 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_649
timestamp 1612251222
transform -1 0 714 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_649
timestamp 1612251222
transform -1 0 698 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_649
timestamp 1612251222
transform -1 0 682 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_600
timestamp 1612251222
transform -1 0 666 0 -1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_600
timestamp 1612251222
transform -1 0 500 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_600
timestamp 1612251222
transform -1 0 484 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_600
timestamp 1612251222
transform -1 0 468 0 -1 7410
box -4 -6 20 206
use PAND2X1  PAND2X1_645
timestamp 1612251222
transform -1 0 452 0 -1 7410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_645
timestamp 1612251222
transform -1 0 286 0 -1 7410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_645
timestamp 1612251222
transform -1 0 270 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_645
timestamp 1612251222
transform -1 0 254 0 -1 7410
box -4 -6 20 206
use FILL  FILL_PAND2X1_645
timestamp 1612251222
transform -1 0 238 0 -1 7410
box -4 -6 20 206
use POR2X1  POR2X1_601
timestamp 1612251222
transform -1 0 222 0 -1 7410
box -4 -6 170 206
use FILL  FILL1_POR2X1_601
timestamp 1612251222
transform -1 0 56 0 -1 7410
box -4 -6 20 206
use FILL  FILL0_POR2X1_601
timestamp 1612251222
transform -1 0 40 0 -1 7410
box -4 -6 20 206
use FILL  FILL_POR2X1_601
timestamp 1612251222
transform -1 0 24 0 -1 7410
box -4 -6 20 206
use FILL  FILL_36_10
timestamp 1612251222
transform 1 0 10246 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_9
timestamp 1612251222
transform 1 0 10230 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_8
timestamp 1612251222
transform 1 0 10214 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_7
timestamp 1612251222
transform 1 0 10198 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_6
timestamp 1612251222
transform 1 0 10182 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_5
timestamp 1612251222
transform 1 0 10166 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_4
timestamp 1612251222
transform 1 0 10150 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_3
timestamp 1612251222
transform 1 0 10134 0 1 7010
box -4 -6 20 206
use FILL  FILL_35_1
timestamp 1612251222
transform -1 0 10268 0 -1 7010
box -4 -6 20 206
use FILL  FILL_36_2
timestamp 1612251222
transform 1 0 10118 0 1 7010
box -4 -6 20 206
use FILL  FILL_36_1
timestamp 1612251222
transform 1 0 10102 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_506
timestamp 1612251222
transform 1 0 10086 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_506
timestamp 1612251222
transform 1 0 10070 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_506
timestamp 1612251222
transform 1 0 10054 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_506
timestamp 1612251222
transform 1 0 10038 0 -1 7010
box -4 -6 20 206
use POR2X1  POR2X1_839
timestamp 1612251222
transform -1 0 10102 0 1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_839
timestamp 1612251222
transform -1 0 9936 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_839
timestamp 1612251222
transform -1 0 9920 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_839
timestamp 1612251222
transform -1 0 9904 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_836
timestamp 1612251222
transform 1 0 9872 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_836
timestamp 1612251222
transform 1 0 9856 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_836
timestamp 1612251222
transform 1 0 9840 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_836
timestamp 1612251222
transform 1 0 9824 0 -1 7010
box -4 -6 20 206
use POR2X1  POR2X1_852
timestamp 1612251222
transform -1 0 9888 0 1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_852
timestamp 1612251222
transform -1 0 9722 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_852
timestamp 1612251222
transform -1 0 9706 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_852
timestamp 1612251222
transform -1 0 9690 0 1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_823
timestamp 1612251222
transform 1 0 9658 0 -1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_823
timestamp 1612251222
transform 1 0 9642 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_823
timestamp 1612251222
transform 1 0 9626 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_823
timestamp 1612251222
transform 1 0 9610 0 -1 7010
box -4 -6 20 206
use POR2X1  POR2X1_508
timestamp 1612251222
transform -1 0 9674 0 1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_508
timestamp 1612251222
transform -1 0 9508 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_508
timestamp 1612251222
transform -1 0 9492 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_508
timestamp 1612251222
transform -1 0 9476 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_823
timestamp 1612251222
transform 1 0 9594 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_627
timestamp 1612251222
transform -1 0 9460 0 1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_627
timestamp 1612251222
transform -1 0 9294 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_627
timestamp 1612251222
transform -1 0 9278 0 1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_824
timestamp 1612251222
transform 1 0 9428 0 -1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_824
timestamp 1612251222
transform 1 0 9412 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_824
timestamp 1612251222
transform 1 0 9396 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_824
timestamp 1612251222
transform 1 0 9380 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_824
timestamp 1612251222
transform 1 0 9364 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_627
timestamp 1612251222
transform -1 0 9262 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_627
timestamp 1612251222
transform -1 0 9246 0 1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_292
timestamp 1612251222
transform -1 0 9364 0 -1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_292
timestamp 1612251222
transform -1 0 9198 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_292
timestamp 1612251222
transform -1 0 9182 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_292
timestamp 1612251222
transform -1 0 9166 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_292
timestamp 1612251222
transform -1 0 9150 0 -1 7010
box -4 -6 20 206
use POR2X1  POR2X1_629
timestamp 1612251222
transform -1 0 9230 0 1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_629
timestamp 1612251222
transform -1 0 9064 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_629
timestamp 1612251222
transform -1 0 9048 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_629
timestamp 1612251222
transform -1 0 9032 0 1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_16
timestamp 1612251222
transform -1 0 9134 0 -1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_16
timestamp 1612251222
transform -1 0 8968 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_16
timestamp 1612251222
transform -1 0 8952 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_16
timestamp 1612251222
transform -1 0 8936 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_626
timestamp 1612251222
transform 1 0 8850 0 1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_626
timestamp 1612251222
transform 1 0 8834 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_626
timestamp 1612251222
transform 1 0 8818 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_626
timestamp 1612251222
transform 1 0 8802 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_626
timestamp 1612251222
transform 1 0 8786 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_16
timestamp 1612251222
transform -1 0 8920 0 -1 7010
box -4 -6 20 206
use POR2X1  POR2X1_194
timestamp 1612251222
transform -1 0 8904 0 -1 7010
box -4 -6 170 206
use PAND2X1  PAND2X1_39
timestamp 1612251222
transform 1 0 8620 0 1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_39
timestamp 1612251222
transform 1 0 8604 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_39
timestamp 1612251222
transform 1 0 8588 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_39
timestamp 1612251222
transform 1 0 8572 0 1 7010
box -4 -6 20 206
use FILL  FILL1_POR2X1_194
timestamp 1612251222
transform -1 0 8738 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_194
timestamp 1612251222
transform -1 0 8722 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_194
timestamp 1612251222
transform -1 0 8706 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_39
timestamp 1612251222
transform 1 0 8556 0 1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_625
timestamp 1612251222
transform 1 0 8390 0 1 7010
box -4 -6 170 206
use POR2X1  POR2X1_200
timestamp 1612251222
transform -1 0 8690 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_200
timestamp 1612251222
transform -1 0 8524 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_200
timestamp 1612251222
transform -1 0 8508 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_200
timestamp 1612251222
transform -1 0 8492 0 -1 7010
box -4 -6 20 206
use FILL  FILL2_PAND2X1_625
timestamp 1612251222
transform 1 0 8374 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_625
timestamp 1612251222
transform 1 0 8358 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_625
timestamp 1612251222
transform 1 0 8342 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_625
timestamp 1612251222
transform 1 0 8326 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_195
timestamp 1612251222
transform 1 0 8310 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_195
timestamp 1612251222
transform 1 0 8294 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_195
timestamp 1612251222
transform 1 0 8278 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_195
timestamp 1612251222
transform 1 0 8262 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_43
timestamp 1612251222
transform 1 0 8160 0 1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_43
timestamp 1612251222
transform 1 0 8144 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_43
timestamp 1612251222
transform 1 0 8128 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_43
timestamp 1612251222
transform 1 0 8112 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_43
timestamp 1612251222
transform 1 0 8096 0 1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_41
timestamp 1612251222
transform 1 0 8096 0 -1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_41
timestamp 1612251222
transform 1 0 8080 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_41
timestamp 1612251222
transform 1 0 8064 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_41
timestamp 1612251222
transform 1 0 8048 0 -1 7010
box -4 -6 20 206
use POR2X1  POR2X1_66
timestamp 1612251222
transform 1 0 7930 0 1 7010
box -4 -6 170 206
use FILL  FILL2_POR2X1_66
timestamp 1612251222
transform 1 0 7914 0 1 7010
box -4 -6 20 206
use FILL  FILL1_POR2X1_66
timestamp 1612251222
transform 1 0 7898 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_66
timestamp 1612251222
transform 1 0 7882 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_66
timestamp 1612251222
transform 1 0 7866 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_41
timestamp 1612251222
transform 1 0 8032 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_393
timestamp 1612251222
transform -1 0 8032 0 -1 7010
box -4 -6 170 206
use POR2X1  POR2X1_61
timestamp 1612251222
transform 1 0 7700 0 1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_393
timestamp 1612251222
transform -1 0 7866 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_393
timestamp 1612251222
transform -1 0 7850 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_393
timestamp 1612251222
transform -1 0 7834 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_393
timestamp 1612251222
transform -1 0 7818 0 -1 7010
box -4 -6 20 206
use FILL  FILL2_POR2X1_61
timestamp 1612251222
transform 1 0 7684 0 1 7010
box -4 -6 20 206
use FILL  FILL1_POR2X1_61
timestamp 1612251222
transform 1 0 7668 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_61
timestamp 1612251222
transform 1 0 7652 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_61
timestamp 1612251222
transform 1 0 7636 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_400
timestamp 1612251222
transform -1 0 7802 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_400
timestamp 1612251222
transform -1 0 7636 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_400
timestamp 1612251222
transform -1 0 7620 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_400
timestamp 1612251222
transform -1 0 7604 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_60
timestamp 1612251222
transform 1 0 7470 0 1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_60
timestamp 1612251222
transform 1 0 7454 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_60
timestamp 1612251222
transform 1 0 7438 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_60
timestamp 1612251222
transform 1 0 7422 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_60
timestamp 1612251222
transform 1 0 7406 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_403
timestamp 1612251222
transform -1 0 7588 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_403
timestamp 1612251222
transform -1 0 7422 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_403
timestamp 1612251222
transform -1 0 7406 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_403
timestamp 1612251222
transform -1 0 7390 0 -1 7010
box -4 -6 20 206
use POR2X1  POR2X1_404
timestamp 1612251222
transform -1 0 7406 0 1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_404
timestamp 1612251222
transform -1 0 7240 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_404
timestamp 1612251222
transform -1 0 7224 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_404
timestamp 1612251222
transform -1 0 7208 0 1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_399
timestamp 1612251222
transform 1 0 7208 0 -1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_399
timestamp 1612251222
transform 1 0 7192 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_399
timestamp 1612251222
transform 1 0 7176 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_397
timestamp 1612251222
transform -1 0 7192 0 1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_397
timestamp 1612251222
transform -1 0 7026 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_397
timestamp 1612251222
transform -1 0 7010 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_399
timestamp 1612251222
transform 1 0 7160 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_399
timestamp 1612251222
transform 1 0 7144 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_397
timestamp 1612251222
transform -1 0 6994 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_397
timestamp 1612251222
transform -1 0 6978 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_398
timestamp 1612251222
transform 1 0 6978 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_398
timestamp 1612251222
transform 1 0 6962 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_398
timestamp 1612251222
transform 1 0 6946 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_398
timestamp 1612251222
transform 1 0 6930 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_82
timestamp 1612251222
transform 1 0 6764 0 -1 7010
box -4 -6 170 206
use PAND2X1  PAND2X1_83
timestamp 1612251222
transform -1 0 6962 0 1 7010
box -4 -6 170 206
use FILL  FILL1_PAND2X1_82
timestamp 1612251222
transform 1 0 6732 0 -1 7010
box -4 -6 20 206
use FILL  FILL2_PAND2X1_82
timestamp 1612251222
transform 1 0 6748 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_83
timestamp 1612251222
transform -1 0 6748 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_83
timestamp 1612251222
transform -1 0 6764 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_83
timestamp 1612251222
transform -1 0 6780 0 1 7010
box -4 -6 20 206
use FILL  FILL2_PAND2X1_83
timestamp 1612251222
transform -1 0 6796 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_82
timestamp 1612251222
transform 1 0 6700 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_82
timestamp 1612251222
transform 1 0 6716 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_27
timestamp 1612251222
transform -1 0 6700 0 -1 7010
box -4 -6 170 206
use POR2X1  POR2X1_35
timestamp 1612251222
transform 1 0 6566 0 1 7010
box -4 -6 170 206
use FILL  FILL_PAND2X1_27
timestamp 1612251222
transform -1 0 6486 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_27
timestamp 1612251222
transform -1 0 6502 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_27
timestamp 1612251222
transform -1 0 6518 0 -1 7010
box -4 -6 20 206
use FILL  FILL2_PAND2X1_27
timestamp 1612251222
transform -1 0 6534 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_35
timestamp 1612251222
transform 1 0 6502 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_35
timestamp 1612251222
transform 1 0 6518 0 1 7010
box -4 -6 20 206
use FILL  FILL1_POR2X1_35
timestamp 1612251222
transform 1 0 6534 0 1 7010
box -4 -6 20 206
use FILL  FILL2_POR2X1_35
timestamp 1612251222
transform 1 0 6550 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_34
timestamp 1612251222
transform -1 0 6502 0 1 7010
box -4 -6 170 206
use FILL  FILL2_POR2X1_34
timestamp 1612251222
transform -1 0 6336 0 1 7010
box -4 -6 20 206
use FILL  FILL1_POR2X1_34
timestamp 1612251222
transform -1 0 6320 0 1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_32
timestamp 1612251222
transform 1 0 6304 0 -1 7010
box -4 -6 170 206
use FILL  FILL0_POR2X1_34
timestamp 1612251222
transform -1 0 6304 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_34
timestamp 1612251222
transform -1 0 6288 0 1 7010
box -4 -6 20 206
use FILL  FILL2_PAND2X1_32
timestamp 1612251222
transform 1 0 6288 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_32
timestamp 1612251222
transform 1 0 6272 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_32
timestamp 1612251222
transform 1 0 6256 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_32
timestamp 1612251222
transform 1 0 6240 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_617
timestamp 1612251222
transform -1 0 6240 0 -1 7010
box -4 -6 170 206
use PAND2X1  PAND2X1_6
timestamp 1612251222
transform 1 0 6106 0 1 7010
box -4 -6 170 206
use FILL  FILL1_PAND2X1_617
timestamp 1612251222
transform -1 0 6058 0 -1 7010
box -4 -6 20 206
use FILL  FILL2_PAND2X1_617
timestamp 1612251222
transform -1 0 6074 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_6
timestamp 1612251222
transform 1 0 6042 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_6
timestamp 1612251222
transform 1 0 6058 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_6
timestamp 1612251222
transform 1 0 6074 0 1 7010
box -4 -6 20 206
use FILL  FILL2_PAND2X1_6
timestamp 1612251222
transform 1 0 6090 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_617
timestamp 1612251222
transform -1 0 6026 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_617
timestamp 1612251222
transform -1 0 6042 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_49
timestamp 1612251222
transform -1 0 6010 0 -1 7010
box -4 -6 170 206
use PAND2X1  PAND2X1_616
timestamp 1612251222
transform -1 0 6042 0 1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_616
timestamp 1612251222
transform -1 0 5876 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_49
timestamp 1612251222
transform -1 0 5796 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_49
timestamp 1612251222
transform -1 0 5812 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_49
timestamp 1612251222
transform -1 0 5828 0 -1 7010
box -4 -6 20 206
use FILL  FILL2_PAND2X1_49
timestamp 1612251222
transform -1 0 5844 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_616
timestamp 1612251222
transform -1 0 5828 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_616
timestamp 1612251222
transform -1 0 5844 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_616
timestamp 1612251222
transform -1 0 5860 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_621
timestamp 1612251222
transform -1 0 5812 0 1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_621
timestamp 1612251222
transform -1 0 5646 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_621
timestamp 1612251222
transform -1 0 5630 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_621
timestamp 1612251222
transform -1 0 5614 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_622
timestamp 1612251222
transform 1 0 5614 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_622
timestamp 1612251222
transform 1 0 5598 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_672
timestamp 1612251222
transform 1 0 5432 0 1 7010
box -4 -6 170 206
use FILL  FILL0_POR2X1_622
timestamp 1612251222
transform 1 0 5582 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_622
timestamp 1612251222
transform 1 0 5566 0 -1 7010
box -4 -6 20 206
use FILL  FILL2_PAND2X1_672
timestamp 1612251222
transform 1 0 5416 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_672
timestamp 1612251222
transform 1 0 5400 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_672
timestamp 1612251222
transform 1 0 5384 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_672
timestamp 1612251222
transform 1 0 5368 0 1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_619
timestamp 1612251222
transform 1 0 5400 0 -1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_619
timestamp 1612251222
transform 1 0 5384 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_619
timestamp 1612251222
transform 1 0 5368 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_619
timestamp 1612251222
transform 1 0 5352 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_619
timestamp 1612251222
transform 1 0 5336 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_618
timestamp 1612251222
transform 1 0 5170 0 -1 7010
box -4 -6 170 206
use PAND2X1  PAND2X1_671
timestamp 1612251222
transform 1 0 5202 0 1 7010
box -4 -6 170 206
use FILL  FILL1_PAND2X1_671
timestamp 1612251222
transform 1 0 5170 0 1 7010
box -4 -6 20 206
use FILL  FILL2_PAND2X1_671
timestamp 1612251222
transform 1 0 5186 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_618
timestamp 1612251222
transform 1 0 5106 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_618
timestamp 1612251222
transform 1 0 5122 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_618
timestamp 1612251222
transform 1 0 5138 0 -1 7010
box -4 -6 20 206
use FILL  FILL2_PAND2X1_618
timestamp 1612251222
transform 1 0 5154 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_671
timestamp 1612251222
transform 1 0 5138 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_671
timestamp 1612251222
transform 1 0 5154 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_8
timestamp 1612251222
transform 1 0 4972 0 1 7010
box -4 -6 170 206
use FILL  FILL2_POR2X1_8
timestamp 1612251222
transform 1 0 4956 0 1 7010
box -4 -6 20 206
use FILL  FILL1_POR2X1_8
timestamp 1612251222
transform 1 0 4940 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_8
timestamp 1612251222
transform 1 0 4924 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_8
timestamp 1612251222
transform 1 0 4908 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_14
timestamp 1612251222
transform -1 0 5106 0 -1 7010
box -4 -6 170 206
use FILL  FILL2_POR2X1_14
timestamp 1612251222
transform -1 0 4940 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_POR2X1_14
timestamp 1612251222
transform -1 0 4924 0 -1 7010
box -4 -6 20 206
use POR2X1  POR2X1_104
timestamp 1612251222
transform -1 0 4908 0 1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_104
timestamp 1612251222
transform -1 0 4742 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_14
timestamp 1612251222
transform -1 0 4908 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_14
timestamp 1612251222
transform -1 0 4892 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_104
timestamp 1612251222
transform -1 0 4726 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_104
timestamp 1612251222
transform -1 0 4710 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_38
timestamp 1612251222
transform -1 0 4876 0 -1 7010
box -4 -6 170 206
use FILL  FILL2_POR2X1_38
timestamp 1612251222
transform -1 0 4710 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_POR2X1_38
timestamp 1612251222
transform -1 0 4694 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_38
timestamp 1612251222
transform -1 0 4678 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_38
timestamp 1612251222
transform -1 0 4662 0 -1 7010
box -4 -6 20 206
use POR2X1  POR2X1_126
timestamp 1612251222
transform 1 0 4528 0 1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_126
timestamp 1612251222
transform 1 0 4512 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_126
timestamp 1612251222
transform 1 0 4496 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_126
timestamp 1612251222
transform 1 0 4480 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_671
timestamp 1612251222
transform -1 0 4646 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_671
timestamp 1612251222
transform -1 0 4480 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_671
timestamp 1612251222
transform -1 0 4464 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_671
timestamp 1612251222
transform -1 0 4448 0 -1 7010
box -4 -6 20 206
use POR2X1  POR2X1_102
timestamp 1612251222
transform -1 0 4480 0 1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_102
timestamp 1612251222
transform -1 0 4314 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_102
timestamp 1612251222
transform -1 0 4298 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_102
timestamp 1612251222
transform -1 0 4282 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_672
timestamp 1612251222
transform -1 0 4432 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_672
timestamp 1612251222
transform -1 0 4266 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_672
timestamp 1612251222
transform -1 0 4250 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_672
timestamp 1612251222
transform -1 0 4234 0 -1 7010
box -4 -6 20 206
use POR2X1  POR2X1_119
timestamp 1612251222
transform -1 0 4266 0 1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_119
timestamp 1612251222
transform -1 0 4100 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_119
timestamp 1612251222
transform -1 0 4084 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_119
timestamp 1612251222
transform -1 0 4068 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_236
timestamp 1612251222
transform 1 0 4052 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_236
timestamp 1612251222
transform 1 0 4036 0 -1 7010
box -4 -6 20 206
use POR2X1  POR2X1_609
timestamp 1612251222
transform -1 0 4052 0 1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_609
timestamp 1612251222
transform -1 0 3886 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_609
timestamp 1612251222
transform -1 0 3870 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_236
timestamp 1612251222
transform 1 0 4020 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_236
timestamp 1612251222
transform 1 0 4004 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_609
timestamp 1612251222
transform -1 0 3854 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_395
timestamp 1612251222
transform -1 0 4004 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_395
timestamp 1612251222
transform -1 0 3838 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_395
timestamp 1612251222
transform -1 0 3822 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_395
timestamp 1612251222
transform -1 0 3806 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_401
timestamp 1612251222
transform -1 0 3790 0 -1 7010
box -4 -6 170 206
use PAND2X1  PAND2X1_608
timestamp 1612251222
transform 1 0 3672 0 1 7010
box -4 -6 170 206
use FILL  FILL1_PAND2X1_401
timestamp 1612251222
transform -1 0 3608 0 -1 7010
box -4 -6 20 206
use FILL  FILL2_PAND2X1_401
timestamp 1612251222
transform -1 0 3624 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_608
timestamp 1612251222
transform 1 0 3608 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_608
timestamp 1612251222
transform 1 0 3624 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_608
timestamp 1612251222
transform 1 0 3640 0 1 7010
box -4 -6 20 206
use FILL  FILL2_PAND2X1_608
timestamp 1612251222
transform 1 0 3656 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_401
timestamp 1612251222
transform -1 0 3576 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_401
timestamp 1612251222
transform -1 0 3592 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_402
timestamp 1612251222
transform -1 0 3560 0 -1 7010
box -4 -6 170 206
use PAND2X1  PAND2X1_240
timestamp 1612251222
transform 1 0 3442 0 1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_240
timestamp 1612251222
transform 1 0 3426 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_402
timestamp 1612251222
transform -1 0 3346 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_402
timestamp 1612251222
transform -1 0 3362 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_402
timestamp 1612251222
transform -1 0 3378 0 -1 7010
box -4 -6 20 206
use FILL  FILL2_PAND2X1_402
timestamp 1612251222
transform -1 0 3394 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_240
timestamp 1612251222
transform 1 0 3378 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_240
timestamp 1612251222
transform 1 0 3394 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_240
timestamp 1612251222
transform 1 0 3410 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_234
timestamp 1612251222
transform 1 0 3212 0 1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_234
timestamp 1612251222
transform 1 0 3196 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_234
timestamp 1612251222
transform 1 0 3180 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_234
timestamp 1612251222
transform 1 0 3164 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_233
timestamp 1612251222
transform -1 0 3330 0 -1 7010
box -4 -6 170 206
use PAND2X1  PAND2X1_404
timestamp 1612251222
transform 1 0 2998 0 1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_404
timestamp 1612251222
transform 1 0 2982 0 1 7010
box -4 -6 20 206
use FILL  FILL1_POR2X1_233
timestamp 1612251222
transform -1 0 3164 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_233
timestamp 1612251222
transform -1 0 3148 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_233
timestamp 1612251222
transform -1 0 3132 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_404
timestamp 1612251222
transform 1 0 2966 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_404
timestamp 1612251222
transform 1 0 2950 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_404
timestamp 1612251222
transform 1 0 2934 0 1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_410
timestamp 1612251222
transform 1 0 2950 0 -1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_410
timestamp 1612251222
transform 1 0 2934 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_410
timestamp 1612251222
transform 1 0 2918 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_410
timestamp 1612251222
transform 1 0 2902 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_410
timestamp 1612251222
transform 1 0 2886 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_403
timestamp 1612251222
transform 1 0 2768 0 1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_403
timestamp 1612251222
transform 1 0 2752 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_403
timestamp 1612251222
transform 1 0 2736 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_403
timestamp 1612251222
transform 1 0 2720 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_403
timestamp 1612251222
transform 1 0 2704 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_290
timestamp 1612251222
transform 1 0 2720 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_290
timestamp 1612251222
transform 1 0 2704 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_290
timestamp 1612251222
transform 1 0 2688 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_290
timestamp 1612251222
transform 1 0 2672 0 -1 7010
box -4 -6 20 206
use POR2X1  POR2X1_399
timestamp 1612251222
transform 1 0 2538 0 1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_399
timestamp 1612251222
transform 1 0 2522 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_399
timestamp 1612251222
transform 1 0 2506 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_399
timestamp 1612251222
transform 1 0 2490 0 1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_520
timestamp 1612251222
transform -1 0 2672 0 -1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_520
timestamp 1612251222
transform -1 0 2506 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_520
timestamp 1612251222
transform -1 0 2490 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_520
timestamp 1612251222
transform -1 0 2474 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_398
timestamp 1612251222
transform 1 0 2324 0 1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_398
timestamp 1612251222
transform 1 0 2308 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_398
timestamp 1612251222
transform 1 0 2292 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_520
timestamp 1612251222
transform -1 0 2458 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_398
timestamp 1612251222
transform 1 0 2276 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_398
timestamp 1612251222
transform 1 0 2260 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_824
timestamp 1612251222
transform -1 0 2442 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_824
timestamp 1612251222
transform -1 0 2276 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_824
timestamp 1612251222
transform -1 0 2260 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_824
timestamp 1612251222
transform -1 0 2244 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_836
timestamp 1612251222
transform -1 0 2260 0 1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_836
timestamp 1612251222
transform -1 0 2094 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_836
timestamp 1612251222
transform -1 0 2078 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_836
timestamp 1612251222
transform -1 0 2062 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_836
timestamp 1612251222
transform -1 0 2046 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_823
timestamp 1612251222
transform 1 0 2062 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_823
timestamp 1612251222
transform 1 0 2046 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_823
timestamp 1612251222
transform 1 0 2030 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_823
timestamp 1612251222
transform 1 0 2014 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_835
timestamp 1612251222
transform 1 0 1848 0 -1 7010
box -4 -6 170 206
use PAND2X1  PAND2X1_839
timestamp 1612251222
transform -1 0 2030 0 1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_839
timestamp 1612251222
transform -1 0 1864 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_835
timestamp 1612251222
transform 1 0 1784 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_835
timestamp 1612251222
transform 1 0 1800 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_835
timestamp 1612251222
transform 1 0 1816 0 -1 7010
box -4 -6 20 206
use FILL  FILL2_PAND2X1_835
timestamp 1612251222
transform 1 0 1832 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_839
timestamp 1612251222
transform -1 0 1816 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_839
timestamp 1612251222
transform -1 0 1832 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_839
timestamp 1612251222
transform -1 0 1848 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_122
timestamp 1612251222
transform 1 0 1634 0 1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_122
timestamp 1612251222
transform 1 0 1618 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_122
timestamp 1612251222
transform 1 0 1602 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_122
timestamp 1612251222
transform 1 0 1586 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_822
timestamp 1612251222
transform 1 0 1618 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_822
timestamp 1612251222
transform 1 0 1602 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_822
timestamp 1612251222
transform 1 0 1586 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_121
timestamp 1612251222
transform 1 0 1420 0 1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_121
timestamp 1612251222
transform 1 0 1404 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_822
timestamp 1612251222
transform 1 0 1570 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_120
timestamp 1612251222
transform -1 0 1570 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_PAND2X1_121
timestamp 1612251222
transform 1 0 1388 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_121
timestamp 1612251222
transform 1 0 1372 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_121
timestamp 1612251222
transform 1 0 1356 0 1 7010
box -4 -6 20 206
use FILL  FILL2_PAND2X1_120
timestamp 1612251222
transform -1 0 1404 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_120
timestamp 1612251222
transform -1 0 1388 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_120
timestamp 1612251222
transform -1 0 1372 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_120
timestamp 1612251222
transform -1 0 1356 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_722
timestamp 1612251222
transform 1 0 1190 0 1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_722
timestamp 1612251222
transform 1 0 1174 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_722
timestamp 1612251222
transform 1 0 1158 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_722
timestamp 1612251222
transform 1 0 1142 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_722
timestamp 1612251222
transform 1 0 1126 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_591
timestamp 1612251222
transform 1 0 1174 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_591
timestamp 1612251222
transform 1 0 1158 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_591
timestamp 1612251222
transform 1 0 1142 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_591
timestamp 1612251222
transform 1 0 1126 0 -1 7010
box -4 -6 20 206
use POR2X1  POR2X1_666
timestamp 1612251222
transform -1 0 1126 0 1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_666
timestamp 1612251222
transform -1 0 960 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_666
timestamp 1612251222
transform -1 0 944 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_666
timestamp 1612251222
transform -1 0 928 0 1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_718
timestamp 1612251222
transform 1 0 960 0 -1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_718
timestamp 1612251222
transform 1 0 944 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_718
timestamp 1612251222
transform 1 0 928 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_718
timestamp 1612251222
transform 1 0 912 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_718
timestamp 1612251222
transform 1 0 896 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_719
timestamp 1612251222
transform 1 0 746 0 1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_719
timestamp 1612251222
transform 1 0 730 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_719
timestamp 1612251222
transform 1 0 714 0 1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_664
timestamp 1612251222
transform -1 0 896 0 -1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_664
timestamp 1612251222
transform -1 0 730 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_719
timestamp 1612251222
transform 1 0 698 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_719
timestamp 1612251222
transform 1 0 682 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_664
timestamp 1612251222
transform -1 0 714 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_664
timestamp 1612251222
transform -1 0 698 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_664
timestamp 1612251222
transform -1 0 682 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_756
timestamp 1612251222
transform -1 0 682 0 1 7010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_756
timestamp 1612251222
transform -1 0 516 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_756
timestamp 1612251222
transform -1 0 500 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_756
timestamp 1612251222
transform -1 0 484 0 1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_756
timestamp 1612251222
transform -1 0 468 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_665
timestamp 1612251222
transform 1 0 500 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_665
timestamp 1612251222
transform 1 0 484 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_665
timestamp 1612251222
transform 1 0 468 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_665
timestamp 1612251222
transform 1 0 452 0 -1 7010
box -4 -6 20 206
use POR2X1  POR2X1_757
timestamp 1612251222
transform -1 0 452 0 1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_757
timestamp 1612251222
transform -1 0 286 0 1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_757
timestamp 1612251222
transform -1 0 270 0 1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_757
timestamp 1612251222
transform -1 0 254 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_755
timestamp 1612251222
transform -1 0 452 0 -1 7010
box -4 -6 170 206
use FILL  FILL1_POR2X1_755
timestamp 1612251222
transform -1 0 286 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_POR2X1_755
timestamp 1612251222
transform -1 0 270 0 -1 7010
box -4 -6 20 206
use FILL  FILL_POR2X1_755
timestamp 1612251222
transform -1 0 254 0 -1 7010
box -4 -6 20 206
use PAND2X1  PAND2X1_791
timestamp 1612251222
transform -1 0 238 0 -1 7010
box -4 -6 170 206
use PAND2X1  PAND2X1_532
timestamp 1612251222
transform -1 0 238 0 1 7010
box -4 -6 170 206
use FILL  FILL_PAND2X1_791
timestamp 1612251222
transform -1 0 24 0 -1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_791
timestamp 1612251222
transform -1 0 40 0 -1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_791
timestamp 1612251222
transform -1 0 56 0 -1 7010
box -4 -6 20 206
use FILL  FILL2_PAND2X1_791
timestamp 1612251222
transform -1 0 72 0 -1 7010
box -4 -6 20 206
use FILL  FILL_PAND2X1_532
timestamp 1612251222
transform -1 0 24 0 1 7010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_532
timestamp 1612251222
transform -1 0 40 0 1 7010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_532
timestamp 1612251222
transform -1 0 56 0 1 7010
box -4 -6 20 206
use FILL  FILL2_PAND2X1_532
timestamp 1612251222
transform -1 0 72 0 1 7010
box -4 -6 20 206
use POR2X1  POR2X1_835
timestamp 1612251222
transform -1 0 10268 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_835
timestamp 1612251222
transform -1 0 10102 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_835
timestamp 1612251222
transform -1 0 10086 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_835
timestamp 1612251222
transform -1 0 10070 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_239
timestamp 1612251222
transform 1 0 9888 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_239
timestamp 1612251222
transform 1 0 9872 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_239
timestamp 1612251222
transform 1 0 9856 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_239
timestamp 1612251222
transform 1 0 9840 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_239
timestamp 1612251222
transform 1 0 9824 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_821
timestamp 1612251222
transform 1 0 9658 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_821
timestamp 1612251222
transform 1 0 9642 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_821
timestamp 1612251222
transform 1 0 9626 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_821
timestamp 1612251222
transform 1 0 9610 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_821
timestamp 1612251222
transform 1 0 9594 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_510
timestamp 1612251222
transform -1 0 9594 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_510
timestamp 1612251222
transform -1 0 9428 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_510
timestamp 1612251222
transform -1 0 9412 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_510
timestamp 1612251222
transform -1 0 9396 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_447
timestamp 1612251222
transform -1 0 9380 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_447
timestamp 1612251222
transform -1 0 9214 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_447
timestamp 1612251222
transform -1 0 9198 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_447
timestamp 1612251222
transform -1 0 9182 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_420
timestamp 1612251222
transform 1 0 9000 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_420
timestamp 1612251222
transform 1 0 8984 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_420
timestamp 1612251222
transform 1 0 8968 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_420
timestamp 1612251222
transform 1 0 8952 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_420
timestamp 1612251222
transform 1 0 8936 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_630
timestamp 1612251222
transform -1 0 8936 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_630
timestamp 1612251222
transform -1 0 8770 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_630
timestamp 1612251222
transform -1 0 8754 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_630
timestamp 1612251222
transform -1 0 8738 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_631
timestamp 1612251222
transform 1 0 8556 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_631
timestamp 1612251222
transform 1 0 8540 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_631
timestamp 1612251222
transform 1 0 8524 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_631
timestamp 1612251222
transform 1 0 8508 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_199
timestamp 1612251222
transform -1 0 8508 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_199
timestamp 1612251222
transform -1 0 8342 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_199
timestamp 1612251222
transform -1 0 8326 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_199
timestamp 1612251222
transform -1 0 8310 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_207
timestamp 1612251222
transform -1 0 8294 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_207
timestamp 1612251222
transform -1 0 8128 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_207
timestamp 1612251222
transform -1 0 8112 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_207
timestamp 1612251222
transform -1 0 8096 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_214
timestamp 1612251222
transform 1 0 7914 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_214
timestamp 1612251222
transform 1 0 7898 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_214
timestamp 1612251222
transform 1 0 7882 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_214
timestamp 1612251222
transform 1 0 7866 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_206
timestamp 1612251222
transform 1 0 7700 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_206
timestamp 1612251222
transform 1 0 7684 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_206
timestamp 1612251222
transform 1 0 7668 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_206
timestamp 1612251222
transform 1 0 7652 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_208
timestamp 1612251222
transform 1 0 7486 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_208
timestamp 1612251222
transform 1 0 7470 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_208
timestamp 1612251222
transform 1 0 7454 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_208
timestamp 1612251222
transform 1 0 7438 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_57
timestamp 1612251222
transform 1 0 7272 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_57
timestamp 1612251222
transform 1 0 7256 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_57
timestamp 1612251222
transform 1 0 7240 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_57
timestamp 1612251222
transform 1 0 7224 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_57
timestamp 1612251222
transform 1 0 7208 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_98
timestamp 1612251222
transform 1 0 7042 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_98
timestamp 1612251222
transform 1 0 7026 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_98
timestamp 1612251222
transform 1 0 7010 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_98
timestamp 1612251222
transform 1 0 6994 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_232
timestamp 1612251222
transform 1 0 6828 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_232
timestamp 1612251222
transform 1 0 6812 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_232
timestamp 1612251222
transform 1 0 6796 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_232
timestamp 1612251222
transform 1 0 6780 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_232
timestamp 1612251222
transform 1 0 6764 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_88
timestamp 1612251222
transform 1 0 6598 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_88
timestamp 1612251222
transform 1 0 6582 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_88
timestamp 1612251222
transform 1 0 6566 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_88
timestamp 1612251222
transform 1 0 6550 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_88
timestamp 1612251222
transform 1 0 6534 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_87
timestamp 1612251222
transform 1 0 6368 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_87
timestamp 1612251222
transform 1 0 6352 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_87
timestamp 1612251222
transform 1 0 6336 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_87
timestamp 1612251222
transform 1 0 6320 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_29
timestamp 1612251222
transform 1 0 6154 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_29
timestamp 1612251222
transform 1 0 6138 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_29
timestamp 1612251222
transform 1 0 6122 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_29
timestamp 1612251222
transform 1 0 6106 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_29
timestamp 1612251222
transform 1 0 6090 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_670
timestamp 1612251222
transform -1 0 6090 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_670
timestamp 1612251222
transform -1 0 5924 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_670
timestamp 1612251222
transform -1 0 5908 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_670
timestamp 1612251222
transform -1 0 5892 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_670
timestamp 1612251222
transform -1 0 5876 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_673
timestamp 1612251222
transform -1 0 5860 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_673
timestamp 1612251222
transform -1 0 5694 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_673
timestamp 1612251222
transform -1 0 5678 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_673
timestamp 1612251222
transform -1 0 5662 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_4
timestamp 1612251222
transform -1 0 5646 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_4
timestamp 1612251222
transform -1 0 5480 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_4
timestamp 1612251222
transform -1 0 5464 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_4
timestamp 1612251222
transform -1 0 5448 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_4
timestamp 1612251222
transform -1 0 5432 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_37
timestamp 1612251222
transform 1 0 5250 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_37
timestamp 1612251222
transform 1 0 5234 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_37
timestamp 1612251222
transform 1 0 5218 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_37
timestamp 1612251222
transform 1 0 5202 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_37
timestamp 1612251222
transform 1 0 5186 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_8
timestamp 1612251222
transform 1 0 5020 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_8
timestamp 1612251222
transform 1 0 5004 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_8
timestamp 1612251222
transform 1 0 4988 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_8
timestamp 1612251222
transform 1 0 4972 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_8
timestamp 1612251222
transform 1 0 4956 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_380
timestamp 1612251222
transform 1 0 4790 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_380
timestamp 1612251222
transform 1 0 4774 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_380
timestamp 1612251222
transform 1 0 4758 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_380
timestamp 1612251222
transform 1 0 4742 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_379
timestamp 1612251222
transform 1 0 4576 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_379
timestamp 1612251222
transform 1 0 4560 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_379
timestamp 1612251222
transform 1 0 4544 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_379
timestamp 1612251222
transform 1 0 4528 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_379
timestamp 1612251222
transform 1 0 4512 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_77
timestamp 1612251222
transform -1 0 4512 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_77
timestamp 1612251222
transform -1 0 4346 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_77
timestamp 1612251222
transform -1 0 4330 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_77
timestamp 1612251222
transform -1 0 4314 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_673
timestamp 1612251222
transform -1 0 4298 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_673
timestamp 1612251222
transform -1 0 4132 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_673
timestamp 1612251222
transform -1 0 4116 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_673
timestamp 1612251222
transform -1 0 4100 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_673
timestamp 1612251222
transform -1 0 4084 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_668
timestamp 1612251222
transform -1 0 4068 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_668
timestamp 1612251222
transform -1 0 3902 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_668
timestamp 1612251222
transform -1 0 3886 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_668
timestamp 1612251222
transform -1 0 3870 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_668
timestamp 1612251222
transform -1 0 3854 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_669
timestamp 1612251222
transform -1 0 3838 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_669
timestamp 1612251222
transform -1 0 3672 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_669
timestamp 1612251222
transform -1 0 3656 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_669
timestamp 1612251222
transform -1 0 3640 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_720
timestamp 1612251222
transform 1 0 3458 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_720
timestamp 1612251222
transform 1 0 3442 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_720
timestamp 1612251222
transform 1 0 3426 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_720
timestamp 1612251222
transform 1 0 3410 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_720
timestamp 1612251222
transform 1 0 3394 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_667
timestamp 1612251222
transform 1 0 3228 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_667
timestamp 1612251222
transform 1 0 3212 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_667
timestamp 1612251222
transform 1 0 3196 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_667
timestamp 1612251222
transform 1 0 3180 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_517
timestamp 1612251222
transform -1 0 3180 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_517
timestamp 1612251222
transform -1 0 3014 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_517
timestamp 1612251222
transform -1 0 2998 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_517
timestamp 1612251222
transform -1 0 2982 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_559
timestamp 1612251222
transform -1 0 2966 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_559
timestamp 1612251222
transform -1 0 2800 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_559
timestamp 1612251222
transform -1 0 2784 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_559
timestamp 1612251222
transform -1 0 2768 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_559
timestamp 1612251222
transform -1 0 2752 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_518
timestamp 1612251222
transform -1 0 2736 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_518
timestamp 1612251222
transform -1 0 2570 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_518
timestamp 1612251222
transform -1 0 2554 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_518
timestamp 1612251222
transform -1 0 2538 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_264
timestamp 1612251222
transform 1 0 2356 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_264
timestamp 1612251222
transform 1 0 2340 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_264
timestamp 1612251222
transform 1 0 2324 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_264
timestamp 1612251222
transform 1 0 2308 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_264
timestamp 1612251222
transform 1 0 2292 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_838
timestamp 1612251222
transform -1 0 2292 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_838
timestamp 1612251222
transform -1 0 2126 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_838
timestamp 1612251222
transform -1 0 2110 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_838
timestamp 1612251222
transform -1 0 2094 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_838
timestamp 1612251222
transform -1 0 2078 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_41
timestamp 1612251222
transform 1 0 1896 0 1 6610
box -4 -6 170 206
use FILL  FILL2_POR2X1_41
timestamp 1612251222
transform 1 0 1880 0 1 6610
box -4 -6 20 206
use FILL  FILL1_POR2X1_41
timestamp 1612251222
transform 1 0 1864 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_41
timestamp 1612251222
transform 1 0 1848 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_41
timestamp 1612251222
transform 1 0 1832 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_852
timestamp 1612251222
transform -1 0 1832 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_852
timestamp 1612251222
transform -1 0 1666 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_852
timestamp 1612251222
transform -1 0 1650 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_852
timestamp 1612251222
transform -1 0 1634 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_852
timestamp 1612251222
transform -1 0 1618 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_194
timestamp 1612251222
transform 1 0 1436 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_194
timestamp 1612251222
transform 1 0 1420 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_194
timestamp 1612251222
transform 1 0 1404 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_194
timestamp 1612251222
transform 1 0 1388 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_194
timestamp 1612251222
transform 1 0 1372 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_16
timestamp 1612251222
transform 1 0 1206 0 1 6610
box -4 -6 170 206
use FILL  FILL2_POR2X1_16
timestamp 1612251222
transform 1 0 1190 0 1 6610
box -4 -6 20 206
use FILL  FILL1_POR2X1_16
timestamp 1612251222
transform 1 0 1174 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_16
timestamp 1612251222
transform 1 0 1158 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_16
timestamp 1612251222
transform 1 0 1142 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_605
timestamp 1612251222
transform -1 0 1142 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_605
timestamp 1612251222
transform -1 0 976 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_605
timestamp 1612251222
transform -1 0 960 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_605
timestamp 1612251222
transform -1 0 944 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_605
timestamp 1612251222
transform -1 0 928 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_686
timestamp 1612251222
transform 1 0 746 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_686
timestamp 1612251222
transform 1 0 730 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_686
timestamp 1612251222
transform 1 0 714 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_686
timestamp 1612251222
transform 1 0 698 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_686
timestamp 1612251222
transform 1 0 682 0 1 6610
box -4 -6 20 206
use POR2X1  POR2X1_684
timestamp 1612251222
transform 1 0 516 0 1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_684
timestamp 1612251222
transform 1 0 500 0 1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_684
timestamp 1612251222
transform 1 0 484 0 1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_684
timestamp 1612251222
transform 1 0 468 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_788
timestamp 1612251222
transform 1 0 302 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_788
timestamp 1612251222
transform 1 0 286 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_788
timestamp 1612251222
transform 1 0 270 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_788
timestamp 1612251222
transform 1 0 254 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_788
timestamp 1612251222
transform 1 0 238 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_792
timestamp 1612251222
transform 1 0 72 0 1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_792
timestamp 1612251222
transform 1 0 56 0 1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_792
timestamp 1612251222
transform 1 0 40 0 1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_792
timestamp 1612251222
transform 1 0 24 0 1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_792
timestamp 1612251222
transform 1 0 8 0 1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_822
timestamp 1612251222
transform 1 0 10102 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_822
timestamp 1612251222
transform 1 0 10086 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_822
timestamp 1612251222
transform 1 0 10070 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_822
timestamp 1612251222
transform 1 0 10054 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_822
timestamp 1612251222
transform 1 0 10038 0 -1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_224
timestamp 1612251222
transform -1 0 10038 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_224
timestamp 1612251222
transform -1 0 9872 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_224
timestamp 1612251222
transform -1 0 9856 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_224
timestamp 1612251222
transform -1 0 9840 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_224
timestamp 1612251222
transform -1 0 9824 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_509
timestamp 1612251222
transform 1 0 9642 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_509
timestamp 1612251222
transform 1 0 9626 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_509
timestamp 1612251222
transform 1 0 9610 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_509
timestamp 1612251222
transform 1 0 9594 0 -1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_52
timestamp 1612251222
transform -1 0 9594 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_52
timestamp 1612251222
transform -1 0 9428 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_52
timestamp 1612251222
transform -1 0 9412 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_52
timestamp 1612251222
transform -1 0 9396 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_52
timestamp 1612251222
transform -1 0 9380 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_555
timestamp 1612251222
transform 1 0 9198 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_555
timestamp 1612251222
transform 1 0 9182 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_555
timestamp 1612251222
transform 1 0 9166 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_555
timestamp 1612251222
transform 1 0 9150 0 -1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_628
timestamp 1612251222
transform -1 0 9150 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_628
timestamp 1612251222
transform -1 0 8984 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_628
timestamp 1612251222
transform -1 0 8968 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_628
timestamp 1612251222
transform -1 0 8952 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_628
timestamp 1612251222
transform -1 0 8936 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_632
timestamp 1612251222
transform 1 0 8754 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_632
timestamp 1612251222
transform 1 0 8738 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_632
timestamp 1612251222
transform 1 0 8722 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_632
timestamp 1612251222
transform 1 0 8706 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_219
timestamp 1612251222
transform 1 0 8540 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_219
timestamp 1612251222
transform 1 0 8524 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_219
timestamp 1612251222
transform 1 0 8508 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_219
timestamp 1612251222
transform 1 0 8492 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_215
timestamp 1612251222
transform 1 0 8326 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_215
timestamp 1612251222
transform 1 0 8310 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_215
timestamp 1612251222
transform 1 0 8294 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_215
timestamp 1612251222
transform 1 0 8278 0 -1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_394
timestamp 1612251222
transform -1 0 8278 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_394
timestamp 1612251222
transform -1 0 8112 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_394
timestamp 1612251222
transform -1 0 8096 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_394
timestamp 1612251222
transform -1 0 8080 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_394
timestamp 1612251222
transform -1 0 8064 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_198
timestamp 1612251222
transform -1 0 8048 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_198
timestamp 1612251222
transform -1 0 7882 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_198
timestamp 1612251222
transform -1 0 7866 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_198
timestamp 1612251222
transform -1 0 7850 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_201
timestamp 1612251222
transform -1 0 7834 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_201
timestamp 1612251222
transform -1 0 7668 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_201
timestamp 1612251222
transform -1 0 7652 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_201
timestamp 1612251222
transform -1 0 7636 0 -1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_291
timestamp 1612251222
transform -1 0 7620 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_291
timestamp 1612251222
transform -1 0 7454 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_291
timestamp 1612251222
transform -1 0 7438 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_291
timestamp 1612251222
transform -1 0 7422 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_291
timestamp 1612251222
transform -1 0 7406 0 -1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_93
timestamp 1612251222
transform -1 0 7390 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_93
timestamp 1612251222
transform -1 0 7224 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_93
timestamp 1612251222
transform -1 0 7208 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_93
timestamp 1612251222
transform -1 0 7192 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_93
timestamp 1612251222
transform -1 0 7176 0 -1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_234
timestamp 1612251222
transform -1 0 7160 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_234
timestamp 1612251222
transform -1 0 6994 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_234
timestamp 1612251222
transform -1 0 6978 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_234
timestamp 1612251222
transform -1 0 6962 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_234
timestamp 1612251222
transform -1 0 6946 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_240
timestamp 1612251222
transform -1 0 6930 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_240
timestamp 1612251222
transform -1 0 6764 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_240
timestamp 1612251222
transform -1 0 6748 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_240
timestamp 1612251222
transform -1 0 6732 0 -1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_233
timestamp 1612251222
transform 1 0 6550 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_233
timestamp 1612251222
transform 1 0 6534 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_233
timestamp 1612251222
transform 1 0 6518 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_233
timestamp 1612251222
transform 1 0 6502 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_233
timestamp 1612251222
transform 1 0 6486 0 -1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_102
timestamp 1612251222
transform 1 0 6320 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_102
timestamp 1612251222
transform 1 0 6304 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_102
timestamp 1612251222
transform 1 0 6288 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_102
timestamp 1612251222
transform 1 0 6272 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_102
timestamp 1612251222
transform 1 0 6256 0 -1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_236
timestamp 1612251222
transform 1 0 6090 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_236
timestamp 1612251222
transform 1 0 6074 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_236
timestamp 1612251222
transform 1 0 6058 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_236
timestamp 1612251222
transform 1 0 6042 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_236
timestamp 1612251222
transform 1 0 6026 0 -1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_54
timestamp 1612251222
transform 1 0 5860 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_54
timestamp 1612251222
transform 1 0 5844 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_54
timestamp 1612251222
transform 1 0 5828 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_54
timestamp 1612251222
transform 1 0 5812 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_54
timestamp 1612251222
transform 1 0 5796 0 -1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_104
timestamp 1612251222
transform -1 0 5796 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_104
timestamp 1612251222
transform -1 0 5630 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_104
timestamp 1612251222
transform -1 0 5614 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_104
timestamp 1612251222
transform -1 0 5598 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_104
timestamp 1612251222
transform -1 0 5582 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_28
timestamp 1612251222
transform -1 0 5566 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_POR2X1_28
timestamp 1612251222
transform -1 0 5400 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_POR2X1_28
timestamp 1612251222
transform -1 0 5384 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_28
timestamp 1612251222
transform -1 0 5368 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_28
timestamp 1612251222
transform -1 0 5352 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_19
timestamp 1612251222
transform -1 0 5336 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_POR2X1_19
timestamp 1612251222
transform -1 0 5170 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_POR2X1_19
timestamp 1612251222
transform -1 0 5154 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_19
timestamp 1612251222
transform -1 0 5138 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_19
timestamp 1612251222
transform -1 0 5122 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_20
timestamp 1612251222
transform -1 0 5106 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_POR2X1_20
timestamp 1612251222
transform -1 0 4940 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_POR2X1_20
timestamp 1612251222
transform -1 0 4924 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_20
timestamp 1612251222
transform -1 0 4908 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_20
timestamp 1612251222
transform -1 0 4892 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_42
timestamp 1612251222
transform -1 0 4876 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_POR2X1_42
timestamp 1612251222
transform -1 0 4710 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_POR2X1_42
timestamp 1612251222
transform -1 0 4694 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_42
timestamp 1612251222
transform -1 0 4678 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_42
timestamp 1612251222
transform -1 0 4662 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_23
timestamp 1612251222
transform 1 0 4480 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_POR2X1_23
timestamp 1612251222
transform 1 0 4464 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_POR2X1_23
timestamp 1612251222
transform 1 0 4448 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_23
timestamp 1612251222
transform 1 0 4432 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_23
timestamp 1612251222
transform 1 0 4416 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_670
timestamp 1612251222
transform -1 0 4416 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_670
timestamp 1612251222
transform -1 0 4250 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_670
timestamp 1612251222
transform -1 0 4234 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_670
timestamp 1612251222
transform -1 0 4218 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_825
timestamp 1612251222
transform -1 0 4202 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_825
timestamp 1612251222
transform -1 0 4036 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_825
timestamp 1612251222
transform -1 0 4020 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_825
timestamp 1612251222
transform -1 0 4004 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_396
timestamp 1612251222
transform -1 0 3988 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_396
timestamp 1612251222
transform -1 0 3822 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_396
timestamp 1612251222
transform -1 0 3806 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_396
timestamp 1612251222
transform -1 0 3790 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_397
timestamp 1612251222
transform -1 0 3774 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_397
timestamp 1612251222
transform -1 0 3608 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_397
timestamp 1612251222
transform -1 0 3592 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_397
timestamp 1612251222
transform -1 0 3576 0 -1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_334
timestamp 1612251222
transform 1 0 3394 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_334
timestamp 1612251222
transform 1 0 3378 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_334
timestamp 1612251222
transform 1 0 3362 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_334
timestamp 1612251222
transform 1 0 3346 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_334
timestamp 1612251222
transform 1 0 3330 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_291
timestamp 1612251222
transform 1 0 3164 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_291
timestamp 1612251222
transform 1 0 3148 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_291
timestamp 1612251222
transform 1 0 3132 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_291
timestamp 1612251222
transform 1 0 3116 0 -1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_837
timestamp 1612251222
transform -1 0 3116 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_837
timestamp 1612251222
transform -1 0 2950 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_837
timestamp 1612251222
transform -1 0 2934 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_837
timestamp 1612251222
transform -1 0 2918 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_837
timestamp 1612251222
transform -1 0 2902 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_43
timestamp 1612251222
transform -1 0 2886 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_POR2X1_43
timestamp 1612251222
transform -1 0 2720 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_POR2X1_43
timestamp 1612251222
transform -1 0 2704 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_43
timestamp 1612251222
transform -1 0 2688 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_43
timestamp 1612251222
transform -1 0 2672 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_519
timestamp 1612251222
transform -1 0 2656 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_519
timestamp 1612251222
transform -1 0 2490 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_519
timestamp 1612251222
transform -1 0 2474 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_519
timestamp 1612251222
transform -1 0 2458 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_827
timestamp 1612251222
transform -1 0 2442 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_827
timestamp 1612251222
transform -1 0 2276 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_827
timestamp 1612251222
transform -1 0 2260 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_827
timestamp 1612251222
transform -1 0 2244 0 -1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_195
timestamp 1612251222
transform 1 0 2062 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_195
timestamp 1612251222
transform 1 0 2046 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_195
timestamp 1612251222
transform 1 0 2030 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_195
timestamp 1612251222
transform 1 0 2014 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_195
timestamp 1612251222
transform 1 0 1998 0 -1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_124
timestamp 1612251222
transform 1 0 1832 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_124
timestamp 1612251222
transform 1 0 1816 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_124
timestamp 1612251222
transform 1 0 1800 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_124
timestamp 1612251222
transform 1 0 1784 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_124
timestamp 1612251222
transform 1 0 1768 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_821
timestamp 1612251222
transform 1 0 1602 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_821
timestamp 1612251222
transform 1 0 1586 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_821
timestamp 1612251222
transform 1 0 1570 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_821
timestamp 1612251222
transform 1 0 1554 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_39
timestamp 1612251222
transform -1 0 1554 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_POR2X1_39
timestamp 1612251222
transform -1 0 1388 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_POR2X1_39
timestamp 1612251222
transform -1 0 1372 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_39
timestamp 1612251222
transform -1 0 1356 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_39
timestamp 1612251222
transform -1 0 1340 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_683
timestamp 1612251222
transform -1 0 1324 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_683
timestamp 1612251222
transform -1 0 1158 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_683
timestamp 1612251222
transform -1 0 1142 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_683
timestamp 1612251222
transform -1 0 1126 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_604
timestamp 1612251222
transform 1 0 944 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_604
timestamp 1612251222
transform 1 0 928 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_604
timestamp 1612251222
transform 1 0 912 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_604
timestamp 1612251222
transform 1 0 896 0 -1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_644
timestamp 1612251222
transform -1 0 896 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_644
timestamp 1612251222
transform -1 0 730 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_644
timestamp 1612251222
transform -1 0 714 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_644
timestamp 1612251222
transform -1 0 698 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_644
timestamp 1612251222
transform -1 0 682 0 -1 6610
box -4 -6 20 206
use PAND2X1  PAND2X1_758
timestamp 1612251222
transform -1 0 666 0 -1 6610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_758
timestamp 1612251222
transform -1 0 500 0 -1 6610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_758
timestamp 1612251222
transform -1 0 484 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_758
timestamp 1612251222
transform -1 0 468 0 -1 6610
box -4 -6 20 206
use FILL  FILL_PAND2X1_758
timestamp 1612251222
transform -1 0 452 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_759
timestamp 1612251222
transform -1 0 436 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_759
timestamp 1612251222
transform -1 0 270 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_759
timestamp 1612251222
transform -1 0 254 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_759
timestamp 1612251222
transform -1 0 238 0 -1 6610
box -4 -6 20 206
use POR2X1  POR2X1_533
timestamp 1612251222
transform 1 0 56 0 -1 6610
box -4 -6 170 206
use FILL  FILL1_POR2X1_533
timestamp 1612251222
transform 1 0 40 0 -1 6610
box -4 -6 20 206
use FILL  FILL0_POR2X1_533
timestamp 1612251222
transform 1 0 24 0 -1 6610
box -4 -6 20 206
use FILL  FILL_POR2X1_533
timestamp 1612251222
transform 1 0 8 0 -1 6610
box -4 -6 20 206
use FILL  FILL_32_1
timestamp 1612251222
transform 1 0 10252 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_238
timestamp 1612251222
transform -1 0 10252 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_238
timestamp 1612251222
transform -1 0 10086 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_238
timestamp 1612251222
transform -1 0 10070 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_238
timestamp 1612251222
transform -1 0 10054 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_238
timestamp 1612251222
transform -1 0 10038 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_242
timestamp 1612251222
transform -1 0 10022 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_242
timestamp 1612251222
transform -1 0 9856 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_242
timestamp 1612251222
transform -1 0 9840 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_242
timestamp 1612251222
transform -1 0 9824 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_227
timestamp 1612251222
transform -1 0 9808 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_227
timestamp 1612251222
transform -1 0 9642 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_227
timestamp 1612251222
transform -1 0 9626 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_227
timestamp 1612251222
transform -1 0 9610 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_340
timestamp 1612251222
transform 1 0 9428 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_340
timestamp 1612251222
transform 1 0 9412 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_340
timestamp 1612251222
transform 1 0 9396 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_340
timestamp 1612251222
transform 1 0 9380 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_258
timestamp 1612251222
transform -1 0 9380 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_258
timestamp 1612251222
transform -1 0 9214 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_258
timestamp 1612251222
transform -1 0 9198 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_258
timestamp 1612251222
transform -1 0 9182 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_258
timestamp 1612251222
transform -1 0 9166 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_259
timestamp 1612251222
transform 1 0 8984 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_259
timestamp 1612251222
transform 1 0 8968 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_259
timestamp 1612251222
transform 1 0 8952 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_259
timestamp 1612251222
transform 1 0 8936 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_7
timestamp 1612251222
transform -1 0 8936 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_7
timestamp 1612251222
transform -1 0 8770 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_7
timestamp 1612251222
transform -1 0 8754 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_7
timestamp 1612251222
transform -1 0 8738 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_7
timestamp 1612251222
transform -1 0 8722 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_228
timestamp 1612251222
transform 1 0 8540 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_228
timestamp 1612251222
transform 1 0 8524 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_228
timestamp 1612251222
transform 1 0 8508 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_228
timestamp 1612251222
transform 1 0 8492 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_197
timestamp 1612251222
transform -1 0 8492 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_197
timestamp 1612251222
transform -1 0 8326 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_197
timestamp 1612251222
transform -1 0 8310 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_197
timestamp 1612251222
transform -1 0 8294 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_345
timestamp 1612251222
transform -1 0 8278 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_345
timestamp 1612251222
transform -1 0 8112 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_345
timestamp 1612251222
transform -1 0 8096 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_345
timestamp 1612251222
transform -1 0 8080 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_244
timestamp 1612251222
transform -1 0 8064 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_244
timestamp 1612251222
transform -1 0 7898 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_244
timestamp 1612251222
transform -1 0 7882 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_244
timestamp 1612251222
transform -1 0 7866 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_99
timestamp 1612251222
transform -1 0 7850 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_99
timestamp 1612251222
transform -1 0 7684 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_99
timestamp 1612251222
transform -1 0 7668 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_99
timestamp 1612251222
transform -1 0 7652 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_100
timestamp 1612251222
transform 1 0 7470 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_100
timestamp 1612251222
transform 1 0 7454 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_100
timestamp 1612251222
transform 1 0 7438 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_100
timestamp 1612251222
transform 1 0 7422 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_86
timestamp 1612251222
transform 1 0 7256 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_86
timestamp 1612251222
transform 1 0 7240 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_86
timestamp 1612251222
transform 1 0 7224 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_86
timestamp 1612251222
transform 1 0 7208 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_86
timestamp 1612251222
transform 1 0 7192 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_85
timestamp 1612251222
transform 1 0 7026 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_85
timestamp 1612251222
transform 1 0 7010 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_85
timestamp 1612251222
transform 1 0 6994 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_85
timestamp 1612251222
transform 1 0 6978 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_85
timestamp 1612251222
transform 1 0 6962 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_243
timestamp 1612251222
transform 1 0 6796 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_243
timestamp 1612251222
transform 1 0 6780 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_243
timestamp 1612251222
transform 1 0 6764 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_243
timestamp 1612251222
transform 1 0 6748 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_92
timestamp 1612251222
transform 1 0 6582 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_92
timestamp 1612251222
transform 1 0 6566 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_92
timestamp 1612251222
transform 1 0 6550 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_92
timestamp 1612251222
transform 1 0 6534 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_92
timestamp 1612251222
transform 1 0 6518 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_77
timestamp 1612251222
transform 1 0 6352 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_77
timestamp 1612251222
transform 1 0 6336 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_77
timestamp 1612251222
transform 1 0 6320 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_77
timestamp 1612251222
transform 1 0 6304 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_77
timestamp 1612251222
transform 1 0 6288 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_38
timestamp 1612251222
transform 1 0 6122 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_38
timestamp 1612251222
transform 1 0 6106 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_38
timestamp 1612251222
transform 1 0 6090 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_38
timestamp 1612251222
transform 1 0 6074 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_38
timestamp 1612251222
transform 1 0 6058 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_624
timestamp 1612251222
transform 1 0 5892 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_624
timestamp 1612251222
transform 1 0 5876 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_624
timestamp 1612251222
transform 1 0 5860 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_624
timestamp 1612251222
transform 1 0 5844 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_55
timestamp 1612251222
transform -1 0 5844 0 1 6210
box -4 -6 170 206
use FILL  FILL2_POR2X1_55
timestamp 1612251222
transform -1 0 5678 0 1 6210
box -4 -6 20 206
use FILL  FILL1_POR2X1_55
timestamp 1612251222
transform -1 0 5662 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_55
timestamp 1612251222
transform -1 0 5646 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_55
timestamp 1612251222
transform -1 0 5630 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_377
timestamp 1612251222
transform 1 0 5448 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_377
timestamp 1612251222
transform 1 0 5432 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_377
timestamp 1612251222
transform 1 0 5416 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_377
timestamp 1612251222
transform 1 0 5400 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_463
timestamp 1612251222
transform -1 0 5400 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_463
timestamp 1612251222
transform -1 0 5234 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_463
timestamp 1612251222
transform -1 0 5218 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_463
timestamp 1612251222
transform -1 0 5202 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_463
timestamp 1612251222
transform -1 0 5186 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_460
timestamp 1612251222
transform 1 0 5004 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_460
timestamp 1612251222
transform 1 0 4988 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_460
timestamp 1612251222
transform 1 0 4972 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_460
timestamp 1612251222
transform 1 0 4956 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_460
timestamp 1612251222
transform 1 0 4940 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_33
timestamp 1612251222
transform -1 0 4940 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_33
timestamp 1612251222
transform -1 0 4774 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_33
timestamp 1612251222
transform -1 0 4758 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_33
timestamp 1612251222
transform -1 0 4742 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_33
timestamp 1612251222
transform -1 0 4726 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_94
timestamp 1612251222
transform -1 0 4710 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_94
timestamp 1612251222
transform -1 0 4544 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_94
timestamp 1612251222
transform -1 0 4528 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_94
timestamp 1612251222
transform -1 0 4512 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_153
timestamp 1612251222
transform -1 0 4496 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_153
timestamp 1612251222
transform -1 0 4330 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_153
timestamp 1612251222
transform -1 0 4314 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_153
timestamp 1612251222
transform -1 0 4298 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_96
timestamp 1612251222
transform -1 0 4282 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_96
timestamp 1612251222
transform -1 0 4116 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_96
timestamp 1612251222
transform -1 0 4100 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_96
timestamp 1612251222
transform -1 0 4084 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_472
timestamp 1612251222
transform -1 0 4068 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_472
timestamp 1612251222
transform -1 0 3902 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_472
timestamp 1612251222
transform -1 0 3886 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_472
timestamp 1612251222
transform -1 0 3870 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_472
timestamp 1612251222
transform -1 0 3854 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_721
timestamp 1612251222
transform -1 0 3838 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_721
timestamp 1612251222
transform -1 0 3672 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_721
timestamp 1612251222
transform -1 0 3656 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_721
timestamp 1612251222
transform -1 0 3640 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_721
timestamp 1612251222
transform -1 0 3624 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_826
timestamp 1612251222
transform -1 0 3608 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_826
timestamp 1612251222
transform -1 0 3442 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_826
timestamp 1612251222
transform -1 0 3426 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_826
timestamp 1612251222
transform -1 0 3410 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_640
timestamp 1612251222
transform 1 0 3228 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_640
timestamp 1612251222
transform 1 0 3212 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_640
timestamp 1612251222
transform 1 0 3196 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_640
timestamp 1612251222
transform 1 0 3180 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_640
timestamp 1612251222
transform 1 0 3164 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_633
timestamp 1612251222
transform 1 0 2998 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_633
timestamp 1612251222
transform 1 0 2982 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_633
timestamp 1612251222
transform 1 0 2966 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_633
timestamp 1612251222
transform 1 0 2950 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_633
timestamp 1612251222
transform 1 0 2934 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_118
timestamp 1612251222
transform 1 0 2768 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_118
timestamp 1612251222
transform 1 0 2752 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_118
timestamp 1612251222
transform 1 0 2736 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_118
timestamp 1612251222
transform 1 0 2720 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_123
timestamp 1612251222
transform -1 0 2720 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_123
timestamp 1612251222
transform -1 0 2554 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_123
timestamp 1612251222
transform -1 0 2538 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_123
timestamp 1612251222
transform -1 0 2522 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_123
timestamp 1612251222
transform -1 0 2506 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_48
timestamp 1612251222
transform -1 0 2490 0 1 6210
box -4 -6 170 206
use FILL  FILL2_POR2X1_48
timestamp 1612251222
transform -1 0 2324 0 1 6210
box -4 -6 20 206
use FILL  FILL1_POR2X1_48
timestamp 1612251222
transform -1 0 2308 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_48
timestamp 1612251222
transform -1 0 2292 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_48
timestamp 1612251222
transform -1 0 2276 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_199
timestamp 1612251222
transform -1 0 2260 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_199
timestamp 1612251222
transform -1 0 2094 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_199
timestamp 1612251222
transform -1 0 2078 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_199
timestamp 1612251222
transform -1 0 2062 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_199
timestamp 1612251222
transform -1 0 2046 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_207
timestamp 1612251222
transform 1 0 1864 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_207
timestamp 1612251222
transform 1 0 1848 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_207
timestamp 1612251222
transform 1 0 1832 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_207
timestamp 1612251222
transform 1 0 1816 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_207
timestamp 1612251222
transform 1 0 1800 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_200
timestamp 1612251222
transform 1 0 1634 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_200
timestamp 1612251222
transform 1 0 1618 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_200
timestamp 1612251222
transform 1 0 1602 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_200
timestamp 1612251222
transform 1 0 1586 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_200
timestamp 1612251222
transform 1 0 1570 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_681
timestamp 1612251222
transform 1 0 1404 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_681
timestamp 1612251222
transform 1 0 1388 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_681
timestamp 1612251222
transform 1 0 1372 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_681
timestamp 1612251222
transform 1 0 1356 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_682
timestamp 1612251222
transform -1 0 1356 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_682
timestamp 1612251222
transform -1 0 1190 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_682
timestamp 1612251222
transform -1 0 1174 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_682
timestamp 1612251222
transform -1 0 1158 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_685
timestamp 1612251222
transform -1 0 1142 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_685
timestamp 1612251222
transform -1 0 976 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_685
timestamp 1612251222
transform -1 0 960 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_685
timestamp 1612251222
transform -1 0 944 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_685
timestamp 1612251222
transform -1 0 928 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_687
timestamp 1612251222
transform -1 0 912 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_687
timestamp 1612251222
transform -1 0 746 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_687
timestamp 1612251222
transform -1 0 730 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_687
timestamp 1612251222
transform -1 0 714 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_687
timestamp 1612251222
transform -1 0 698 0 1 6210
box -4 -6 20 206
use POR2X1  POR2X1_534
timestamp 1612251222
transform -1 0 682 0 1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_534
timestamp 1612251222
transform -1 0 516 0 1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_534
timestamp 1612251222
transform -1 0 500 0 1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_534
timestamp 1612251222
transform -1 0 484 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_535
timestamp 1612251222
transform -1 0 468 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_535
timestamp 1612251222
transform -1 0 302 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_535
timestamp 1612251222
transform -1 0 286 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_535
timestamp 1612251222
transform -1 0 270 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_535
timestamp 1612251222
transform -1 0 254 0 1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_856
timestamp 1612251222
transform 1 0 72 0 1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_856
timestamp 1612251222
transform 1 0 56 0 1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_856
timestamp 1612251222
transform 1 0 40 0 1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_856
timestamp 1612251222
transform 1 0 24 0 1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_856
timestamp 1612251222
transform 1 0 8 0 1 6210
box -4 -6 20 206
use FILL  FILL_31_1
timestamp 1612251222
transform -1 0 10268 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_241
timestamp 1612251222
transform -1 0 10252 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_241
timestamp 1612251222
transform -1 0 10086 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_241
timestamp 1612251222
transform -1 0 10070 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_241
timestamp 1612251222
transform -1 0 10054 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_226
timestamp 1612251222
transform 1 0 9872 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_226
timestamp 1612251222
transform 1 0 9856 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_226
timestamp 1612251222
transform 1 0 9840 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_226
timestamp 1612251222
transform 1 0 9824 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_226
timestamp 1612251222
transform 1 0 9808 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_503
timestamp 1612251222
transform -1 0 9808 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_503
timestamp 1612251222
transform -1 0 9642 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_503
timestamp 1612251222
transform -1 0 9626 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_503
timestamp 1612251222
transform -1 0 9610 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_503
timestamp 1612251222
transform -1 0 9594 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_338
timestamp 1612251222
transform -1 0 9578 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_338
timestamp 1612251222
transform -1 0 9412 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_338
timestamp 1612251222
transform -1 0 9396 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_338
timestamp 1612251222
transform -1 0 9380 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_97
timestamp 1612251222
transform -1 0 9364 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_97
timestamp 1612251222
transform -1 0 9198 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_97
timestamp 1612251222
transform -1 0 9182 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_97
timestamp 1612251222
transform -1 0 9166 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_89
timestamp 1612251222
transform 1 0 8984 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_89
timestamp 1612251222
transform 1 0 8968 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_89
timestamp 1612251222
transform 1 0 8952 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_89
timestamp 1612251222
transform 1 0 8936 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_89
timestamp 1612251222
transform 1 0 8920 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_257
timestamp 1612251222
transform -1 0 8920 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_257
timestamp 1612251222
transform -1 0 8754 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_257
timestamp 1612251222
transform -1 0 8738 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_257
timestamp 1612251222
transform -1 0 8722 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_257
timestamp 1612251222
transform -1 0 8706 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_193
timestamp 1612251222
transform 1 0 8524 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_193
timestamp 1612251222
transform 1 0 8508 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_193
timestamp 1612251222
transform 1 0 8492 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_193
timestamp 1612251222
transform 1 0 8476 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_196
timestamp 1612251222
transform 1 0 8310 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_196
timestamp 1612251222
transform 1 0 8294 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_196
timestamp 1612251222
transform 1 0 8278 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_196
timestamp 1612251222
transform 1 0 8262 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_261
timestamp 1612251222
transform 1 0 8096 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_261
timestamp 1612251222
transform 1 0 8080 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_261
timestamp 1612251222
transform 1 0 8064 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_261
timestamp 1612251222
transform 1 0 8048 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_261
timestamp 1612251222
transform 1 0 8032 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_348
timestamp 1612251222
transform -1 0 8032 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_348
timestamp 1612251222
transform -1 0 7866 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_348
timestamp 1612251222
transform -1 0 7850 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_348
timestamp 1612251222
transform -1 0 7834 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_360
timestamp 1612251222
transform 1 0 7652 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_360
timestamp 1612251222
transform 1 0 7636 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_360
timestamp 1612251222
transform 1 0 7620 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_360
timestamp 1612251222
transform 1 0 7604 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_101
timestamp 1612251222
transform -1 0 7604 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_101
timestamp 1612251222
transform -1 0 7438 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_101
timestamp 1612251222
transform -1 0 7422 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_101
timestamp 1612251222
transform -1 0 7406 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_334
timestamp 1612251222
transform 1 0 7224 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_334
timestamp 1612251222
transform 1 0 7208 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_334
timestamp 1612251222
transform 1 0 7192 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_334
timestamp 1612251222
transform 1 0 7176 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_15
timestamp 1612251222
transform -1 0 7176 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_15
timestamp 1612251222
transform -1 0 7010 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_15
timestamp 1612251222
transform -1 0 6994 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_15
timestamp 1612251222
transform -1 0 6978 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_15
timestamp 1612251222
transform -1 0 6962 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_290
timestamp 1612251222
transform -1 0 6946 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_290
timestamp 1612251222
transform -1 0 6780 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_290
timestamp 1612251222
transform -1 0 6764 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_290
timestamp 1612251222
transform -1 0 6748 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_290
timestamp 1612251222
transform -1 0 6732 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_235
timestamp 1612251222
transform 1 0 6550 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_235
timestamp 1612251222
transform 1 0 6534 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_235
timestamp 1612251222
transform 1 0 6518 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_235
timestamp 1612251222
transform 1 0 6502 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_235
timestamp 1612251222
transform 1 0 6486 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_10
timestamp 1612251222
transform 1 0 6320 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_10
timestamp 1612251222
transform 1 0 6304 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_10
timestamp 1612251222
transform 1 0 6288 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_10
timestamp 1612251222
transform 1 0 6272 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_10
timestamp 1612251222
transform 1 0 6256 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_613
timestamp 1612251222
transform -1 0 6256 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_613
timestamp 1612251222
transform -1 0 6090 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_613
timestamp 1612251222
transform -1 0 6074 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_613
timestamp 1612251222
transform -1 0 6058 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_613
timestamp 1612251222
transform -1 0 6042 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_620
timestamp 1612251222
transform -1 0 6026 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_620
timestamp 1612251222
transform -1 0 5860 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_620
timestamp 1612251222
transform -1 0 5844 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_620
timestamp 1612251222
transform -1 0 5828 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_623
timestamp 1612251222
transform 1 0 5646 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_623
timestamp 1612251222
transform 1 0 5630 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_623
timestamp 1612251222
transform 1 0 5614 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_623
timestamp 1612251222
transform 1 0 5598 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_378
timestamp 1612251222
transform -1 0 5598 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_378
timestamp 1612251222
transform -1 0 5432 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_378
timestamp 1612251222
transform -1 0 5416 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_378
timestamp 1612251222
transform -1 0 5400 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_459
timestamp 1612251222
transform 1 0 5218 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_459
timestamp 1612251222
transform 1 0 5202 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_459
timestamp 1612251222
transform 1 0 5186 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_459
timestamp 1612251222
transform 1 0 5170 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_459
timestamp 1612251222
transform 1 0 5154 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_159
timestamp 1612251222
transform 1 0 4988 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_159
timestamp 1612251222
transform 1 0 4972 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_159
timestamp 1612251222
transform 1 0 4956 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_159
timestamp 1612251222
transform 1 0 4940 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_159
timestamp 1612251222
transform 1 0 4924 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_409
timestamp 1612251222
transform 1 0 4758 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_409
timestamp 1612251222
transform 1 0 4742 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_409
timestamp 1612251222
transform 1 0 4726 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_409
timestamp 1612251222
transform 1 0 4710 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_29
timestamp 1612251222
transform 1 0 4544 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_POR2X1_29
timestamp 1612251222
transform 1 0 4528 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_POR2X1_29
timestamp 1612251222
transform 1 0 4512 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_29
timestamp 1612251222
transform 1 0 4496 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_29
timestamp 1612251222
transform 1 0 4480 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_24
timestamp 1612251222
transform 1 0 4314 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_POR2X1_24
timestamp 1612251222
transform 1 0 4298 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_POR2X1_24
timestamp 1612251222
transform 1 0 4282 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_24
timestamp 1612251222
transform 1 0 4266 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_24
timestamp 1612251222
transform 1 0 4250 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_49
timestamp 1612251222
transform -1 0 4250 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_POR2X1_49
timestamp 1612251222
transform -1 0 4084 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_POR2X1_49
timestamp 1612251222
transform -1 0 4068 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_49
timestamp 1612251222
transform -1 0 4052 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_49
timestamp 1612251222
transform -1 0 4036 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_407
timestamp 1612251222
transform -1 0 4020 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_407
timestamp 1612251222
transform -1 0 3854 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_407
timestamp 1612251222
transform -1 0 3838 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_407
timestamp 1612251222
transform -1 0 3822 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_407
timestamp 1612251222
transform -1 0 3806 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_82
timestamp 1612251222
transform -1 0 3790 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_82
timestamp 1612251222
transform -1 0 3624 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_82
timestamp 1612251222
transform -1 0 3608 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_82
timestamp 1612251222
transform -1 0 3592 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_46
timestamp 1612251222
transform -1 0 3576 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_POR2X1_46
timestamp 1612251222
transform -1 0 3410 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_POR2X1_46
timestamp 1612251222
transform -1 0 3394 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_46
timestamp 1612251222
transform -1 0 3378 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_46
timestamp 1612251222
transform -1 0 3362 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_650
timestamp 1612251222
transform -1 0 3346 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_650
timestamp 1612251222
transform -1 0 3180 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_650
timestamp 1612251222
transform -1 0 3164 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_650
timestamp 1612251222
transform -1 0 3148 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_650
timestamp 1612251222
transform -1 0 3132 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_654
timestamp 1612251222
transform -1 0 3116 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_654
timestamp 1612251222
transform -1 0 2950 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_654
timestamp 1612251222
transform -1 0 2934 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_654
timestamp 1612251222
transform -1 0 2918 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_654
timestamp 1612251222
transform -1 0 2902 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_277
timestamp 1612251222
transform -1 0 2886 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_277
timestamp 1612251222
transform -1 0 2720 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_277
timestamp 1612251222
transform -1 0 2704 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_277
timestamp 1612251222
transform -1 0 2688 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_117
timestamp 1612251222
transform 1 0 2506 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_117
timestamp 1612251222
transform 1 0 2490 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_117
timestamp 1612251222
transform 1 0 2474 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_117
timestamp 1612251222
transform 1 0 2458 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_196
timestamp 1612251222
transform 1 0 2292 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_196
timestamp 1612251222
transform 1 0 2276 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_196
timestamp 1612251222
transform 1 0 2260 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_196
timestamp 1612251222
transform 1 0 2244 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_196
timestamp 1612251222
transform 1 0 2228 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_828
timestamp 1612251222
transform -1 0 2228 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_828
timestamp 1612251222
transform -1 0 2062 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_828
timestamp 1612251222
transform -1 0 2046 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_828
timestamp 1612251222
transform -1 0 2030 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_828
timestamp 1612251222
transform -1 0 2014 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_599
timestamp 1612251222
transform -1 0 1998 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_599
timestamp 1612251222
transform -1 0 1832 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_599
timestamp 1612251222
transform -1 0 1816 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_599
timestamp 1612251222
transform -1 0 1800 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_661
timestamp 1612251222
transform -1 0 1784 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_661
timestamp 1612251222
transform -1 0 1618 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_661
timestamp 1612251222
transform -1 0 1602 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_661
timestamp 1612251222
transform -1 0 1586 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_661
timestamp 1612251222
transform -1 0 1570 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_596
timestamp 1612251222
transform -1 0 1554 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_596
timestamp 1612251222
transform -1 0 1388 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_596
timestamp 1612251222
transform -1 0 1372 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_596
timestamp 1612251222
transform -1 0 1356 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_596
timestamp 1612251222
transform -1 0 1340 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_603
timestamp 1612251222
transform -1 0 1324 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_603
timestamp 1612251222
transform -1 0 1158 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_603
timestamp 1612251222
transform -1 0 1142 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_603
timestamp 1612251222
transform -1 0 1126 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_597
timestamp 1612251222
transform -1 0 1110 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_597
timestamp 1612251222
transform -1 0 944 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_597
timestamp 1612251222
transform -1 0 928 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_597
timestamp 1612251222
transform -1 0 912 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_761
timestamp 1612251222
transform -1 0 896 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_761
timestamp 1612251222
transform -1 0 730 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_761
timestamp 1612251222
transform -1 0 714 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_761
timestamp 1612251222
transform -1 0 698 0 -1 6210
box -4 -6 20 206
use POR2X1  POR2X1_829
timestamp 1612251222
transform -1 0 682 0 -1 6210
box -4 -6 170 206
use FILL  FILL1_POR2X1_829
timestamp 1612251222
transform -1 0 516 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_POR2X1_829
timestamp 1612251222
transform -1 0 500 0 -1 6210
box -4 -6 20 206
use FILL  FILL_POR2X1_829
timestamp 1612251222
transform -1 0 484 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_855
timestamp 1612251222
transform -1 0 468 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_855
timestamp 1612251222
transform -1 0 302 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_855
timestamp 1612251222
transform -1 0 286 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_855
timestamp 1612251222
transform -1 0 270 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_855
timestamp 1612251222
transform -1 0 254 0 -1 6210
box -4 -6 20 206
use PAND2X1  PAND2X1_854
timestamp 1612251222
transform -1 0 238 0 -1 6210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_854
timestamp 1612251222
transform -1 0 72 0 -1 6210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_854
timestamp 1612251222
transform -1 0 56 0 -1 6210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_854
timestamp 1612251222
transform -1 0 40 0 -1 6210
box -4 -6 20 206
use FILL  FILL_PAND2X1_854
timestamp 1612251222
transform -1 0 24 0 -1 6210
box -4 -6 20 206
use FILL  FILL_30_13
timestamp 1612251222
transform 1 0 10246 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_12
timestamp 1612251222
transform 1 0 10230 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_11
timestamp 1612251222
transform 1 0 10214 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_10
timestamp 1612251222
transform 1 0 10198 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_9
timestamp 1612251222
transform 1 0 10182 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_8
timestamp 1612251222
transform 1 0 10166 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_7
timestamp 1612251222
transform 1 0 10150 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_6
timestamp 1612251222
transform 1 0 10134 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_5
timestamp 1612251222
transform 1 0 10118 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_4
timestamp 1612251222
transform 1 0 10102 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_3
timestamp 1612251222
transform 1 0 10086 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_2
timestamp 1612251222
transform 1 0 10070 0 1 5810
box -4 -6 20 206
use FILL  FILL_30_1
timestamp 1612251222
transform 1 0 10054 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_358
timestamp 1612251222
transform 1 0 9888 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_358
timestamp 1612251222
transform 1 0 9872 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_358
timestamp 1612251222
transform 1 0 9856 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_358
timestamp 1612251222
transform 1 0 9840 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_350
timestamp 1612251222
transform 1 0 9674 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_350
timestamp 1612251222
transform 1 0 9658 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_350
timestamp 1612251222
transform 1 0 9642 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_350
timestamp 1612251222
transform 1 0 9626 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_351
timestamp 1612251222
transform 1 0 9460 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_351
timestamp 1612251222
transform 1 0 9444 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_351
timestamp 1612251222
transform 1 0 9428 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_351
timestamp 1612251222
transform 1 0 9412 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_562
timestamp 1612251222
transform 1 0 9246 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_562
timestamp 1612251222
transform 1 0 9230 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_562
timestamp 1612251222
transform 1 0 9214 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_562
timestamp 1612251222
transform 1 0 9198 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_339
timestamp 1612251222
transform 1 0 9032 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_339
timestamp 1612251222
transform 1 0 9016 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_339
timestamp 1612251222
transform 1 0 9000 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_339
timestamp 1612251222
transform 1 0 8984 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_252
timestamp 1612251222
transform -1 0 8984 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_252
timestamp 1612251222
transform -1 0 8818 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_252
timestamp 1612251222
transform -1 0 8802 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_252
timestamp 1612251222
transform -1 0 8786 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_252
timestamp 1612251222
transform -1 0 8770 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_556
timestamp 1612251222
transform 1 0 8588 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_556
timestamp 1612251222
transform 1 0 8572 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_556
timestamp 1612251222
transform 1 0 8556 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_556
timestamp 1612251222
transform 1 0 8540 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_45
timestamp 1612251222
transform -1 0 8540 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_45
timestamp 1612251222
transform -1 0 8374 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_45
timestamp 1612251222
transform -1 0 8358 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_45
timestamp 1612251222
transform -1 0 8342 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_45
timestamp 1612251222
transform -1 0 8326 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_363
timestamp 1612251222
transform 1 0 8144 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_363
timestamp 1612251222
transform 1 0 8128 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_363
timestamp 1612251222
transform 1 0 8112 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_363
timestamp 1612251222
transform 1 0 8096 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_359
timestamp 1612251222
transform 1 0 7930 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_359
timestamp 1612251222
transform 1 0 7914 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_359
timestamp 1612251222
transform 1 0 7898 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_359
timestamp 1612251222
transform 1 0 7882 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_349
timestamp 1612251222
transform 1 0 7716 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_349
timestamp 1612251222
transform 1 0 7700 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_349
timestamp 1612251222
transform 1 0 7684 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_349
timestamp 1612251222
transform 1 0 7668 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_342
timestamp 1612251222
transform 1 0 7502 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_342
timestamp 1612251222
transform 1 0 7486 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_342
timestamp 1612251222
transform 1 0 7470 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_342
timestamp 1612251222
transform 1 0 7454 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_248
timestamp 1612251222
transform 1 0 7288 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_248
timestamp 1612251222
transform 1 0 7272 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_248
timestamp 1612251222
transform 1 0 7256 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_248
timestamp 1612251222
transform 1 0 7240 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_248
timestamp 1612251222
transform 1 0 7224 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_247
timestamp 1612251222
transform 1 0 7058 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_247
timestamp 1612251222
transform 1 0 7042 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_247
timestamp 1612251222
transform 1 0 7026 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_247
timestamp 1612251222
transform 1 0 7010 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_84
timestamp 1612251222
transform 1 0 6844 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_84
timestamp 1612251222
transform 1 0 6828 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_84
timestamp 1612251222
transform 1 0 6812 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_84
timestamp 1612251222
transform 1 0 6796 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_490
timestamp 1612251222
transform -1 0 6796 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_490
timestamp 1612251222
transform -1 0 6630 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_490
timestamp 1612251222
transform -1 0 6614 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_490
timestamp 1612251222
transform -1 0 6598 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_490
timestamp 1612251222
transform -1 0 6582 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_528
timestamp 1612251222
transform -1 0 6566 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_528
timestamp 1612251222
transform -1 0 6400 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_528
timestamp 1612251222
transform -1 0 6384 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_528
timestamp 1612251222
transform -1 0 6368 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_528
timestamp 1612251222
transform -1 0 6352 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_530
timestamp 1612251222
transform -1 0 6336 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_530
timestamp 1612251222
transform -1 0 6170 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_530
timestamp 1612251222
transform -1 0 6154 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_530
timestamp 1612251222
transform -1 0 6138 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_530
timestamp 1612251222
transform -1 0 6122 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_133
timestamp 1612251222
transform -1 0 6106 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_133
timestamp 1612251222
transform -1 0 5940 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_133
timestamp 1612251222
transform -1 0 5924 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_133
timestamp 1612251222
transform -1 0 5908 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_133
timestamp 1612251222
transform -1 0 5892 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_126
timestamp 1612251222
transform 1 0 5710 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_126
timestamp 1612251222
transform 1 0 5694 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_126
timestamp 1612251222
transform 1 0 5678 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_126
timestamp 1612251222
transform 1 0 5662 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_126
timestamp 1612251222
transform 1 0 5646 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_9
timestamp 1612251222
transform 1 0 5480 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_9
timestamp 1612251222
transform 1 0 5464 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_9
timestamp 1612251222
transform 1 0 5448 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_9
timestamp 1612251222
transform 1 0 5432 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_9
timestamp 1612251222
transform 1 0 5416 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_62
timestamp 1612251222
transform -1 0 5416 0 1 5810
box -4 -6 170 206
use FILL  FILL2_POR2X1_62
timestamp 1612251222
transform -1 0 5250 0 1 5810
box -4 -6 20 206
use FILL  FILL1_POR2X1_62
timestamp 1612251222
transform -1 0 5234 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_62
timestamp 1612251222
transform -1 0 5218 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_62
timestamp 1612251222
transform -1 0 5202 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_375
timestamp 1612251222
transform 1 0 5020 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_375
timestamp 1612251222
transform 1 0 5004 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_375
timestamp 1612251222
transform 1 0 4988 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_375
timestamp 1612251222
transform 1 0 4972 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_375
timestamp 1612251222
transform 1 0 4956 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_32
timestamp 1612251222
transform -1 0 4956 0 1 5810
box -4 -6 170 206
use FILL  FILL2_POR2X1_32
timestamp 1612251222
transform -1 0 4790 0 1 5810
box -4 -6 20 206
use FILL  FILL1_POR2X1_32
timestamp 1612251222
transform -1 0 4774 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_32
timestamp 1612251222
transform -1 0 4758 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_32
timestamp 1612251222
transform -1 0 4742 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_34
timestamp 1612251222
transform -1 0 4726 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_34
timestamp 1612251222
transform -1 0 4560 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_34
timestamp 1612251222
transform -1 0 4544 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_34
timestamp 1612251222
transform -1 0 4528 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_34
timestamp 1612251222
transform -1 0 4512 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_35
timestamp 1612251222
transform -1 0 4496 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_35
timestamp 1612251222
transform -1 0 4330 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_35
timestamp 1612251222
transform -1 0 4314 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_35
timestamp 1612251222
transform -1 0 4298 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_35
timestamp 1612251222
transform -1 0 4282 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_263
timestamp 1612251222
transform -1 0 4266 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_263
timestamp 1612251222
transform -1 0 4100 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_263
timestamp 1612251222
transform -1 0 4084 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_263
timestamp 1612251222
transform -1 0 4068 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_845
timestamp 1612251222
transform -1 0 4052 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_845
timestamp 1612251222
transform -1 0 3886 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_845
timestamp 1612251222
transform -1 0 3870 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_845
timestamp 1612251222
transform -1 0 3854 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_845
timestamp 1612251222
transform -1 0 3838 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_85
timestamp 1612251222
transform -1 0 3822 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_85
timestamp 1612251222
transform -1 0 3656 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_85
timestamp 1612251222
transform -1 0 3640 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_85
timestamp 1612251222
transform -1 0 3624 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_243
timestamp 1612251222
transform -1 0 3608 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_243
timestamp 1612251222
transform -1 0 3442 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_243
timestamp 1612251222
transform -1 0 3426 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_243
timestamp 1612251222
transform -1 0 3410 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_243
timestamp 1612251222
transform -1 0 3394 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_83
timestamp 1612251222
transform -1 0 3378 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_83
timestamp 1612251222
transform -1 0 3212 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_83
timestamp 1612251222
transform -1 0 3196 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_83
timestamp 1612251222
transform -1 0 3180 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_229
timestamp 1612251222
transform 1 0 2998 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_229
timestamp 1612251222
transform 1 0 2982 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_229
timestamp 1612251222
transform 1 0 2966 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_229
timestamp 1612251222
transform 1 0 2950 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_278
timestamp 1612251222
transform -1 0 2950 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_278
timestamp 1612251222
transform -1 0 2784 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_278
timestamp 1612251222
transform -1 0 2768 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_278
timestamp 1612251222
transform -1 0 2752 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_265
timestamp 1612251222
transform -1 0 2736 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_265
timestamp 1612251222
transform -1 0 2570 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_265
timestamp 1612251222
transform -1 0 2554 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_265
timestamp 1612251222
transform -1 0 2538 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_327
timestamp 1612251222
transform -1 0 2522 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_327
timestamp 1612251222
transform -1 0 2356 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_327
timestamp 1612251222
transform -1 0 2340 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_327
timestamp 1612251222
transform -1 0 2324 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_327
timestamp 1612251222
transform -1 0 2308 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_208
timestamp 1612251222
transform -1 0 2292 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_208
timestamp 1612251222
transform -1 0 2126 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_208
timestamp 1612251222
transform -1 0 2110 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_208
timestamp 1612251222
transform -1 0 2094 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_208
timestamp 1612251222
transform -1 0 2078 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_214
timestamp 1612251222
transform -1 0 2062 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_214
timestamp 1612251222
transform -1 0 1896 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_214
timestamp 1612251222
transform -1 0 1880 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_214
timestamp 1612251222
transform -1 0 1864 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_214
timestamp 1612251222
transform -1 0 1848 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_853
timestamp 1612251222
transform -1 0 1832 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_853
timestamp 1612251222
transform -1 0 1666 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_853
timestamp 1612251222
transform -1 0 1650 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_853
timestamp 1612251222
transform -1 0 1634 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_853
timestamp 1612251222
transform -1 0 1618 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_857
timestamp 1612251222
transform -1 0 1602 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_857
timestamp 1612251222
transform -1 0 1436 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_857
timestamp 1612251222
transform -1 0 1420 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_857
timestamp 1612251222
transform -1 0 1404 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_857
timestamp 1612251222
transform -1 0 1388 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_249
timestamp 1612251222
transform -1 0 1372 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_249
timestamp 1612251222
transform -1 0 1206 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_249
timestamp 1612251222
transform -1 0 1190 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_249
timestamp 1612251222
transform -1 0 1174 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_249
timestamp 1612251222
transform -1 0 1158 0 1 5810
box -4 -6 20 206
use POR2X1  POR2X1_595
timestamp 1612251222
transform -1 0 1142 0 1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_595
timestamp 1612251222
transform -1 0 976 0 1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_595
timestamp 1612251222
transform -1 0 960 0 1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_595
timestamp 1612251222
transform -1 0 944 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_729
timestamp 1612251222
transform 1 0 762 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_729
timestamp 1612251222
transform 1 0 746 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_729
timestamp 1612251222
transform 1 0 730 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_729
timestamp 1612251222
transform 1 0 714 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_729
timestamp 1612251222
transform 1 0 698 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_800
timestamp 1612251222
transform -1 0 698 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_800
timestamp 1612251222
transform -1 0 532 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_800
timestamp 1612251222
transform -1 0 516 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_800
timestamp 1612251222
transform -1 0 500 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_800
timestamp 1612251222
transform -1 0 484 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_801
timestamp 1612251222
transform -1 0 468 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_801
timestamp 1612251222
transform -1 0 302 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_801
timestamp 1612251222
transform -1 0 286 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_801
timestamp 1612251222
transform -1 0 270 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_801
timestamp 1612251222
transform -1 0 254 0 1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_863
timestamp 1612251222
transform -1 0 238 0 1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_863
timestamp 1612251222
transform -1 0 72 0 1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_863
timestamp 1612251222
transform -1 0 56 0 1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_863
timestamp 1612251222
transform -1 0 40 0 1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_863
timestamp 1612251222
transform -1 0 24 0 1 5810
box -4 -6 20 206
use FILL  FILL_29_13
timestamp 1612251222
transform -1 0 10262 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_12
timestamp 1612251222
transform -1 0 10246 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_11
timestamp 1612251222
transform -1 0 10230 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_10
timestamp 1612251222
transform -1 0 10214 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_9
timestamp 1612251222
transform -1 0 10198 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_8
timestamp 1612251222
transform -1 0 10182 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_7
timestamp 1612251222
transform -1 0 10166 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_6
timestamp 1612251222
transform -1 0 10150 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_5
timestamp 1612251222
transform -1 0 10134 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_4
timestamp 1612251222
transform -1 0 10118 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_3
timestamp 1612251222
transform -1 0 10102 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_2
timestamp 1612251222
transform -1 0 10086 0 -1 5810
box -4 -6 20 206
use FILL  FILL_29_1
timestamp 1612251222
transform -1 0 10070 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_333
timestamp 1612251222
transform 1 0 9888 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_333
timestamp 1612251222
transform 1 0 9872 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_333
timestamp 1612251222
transform 1 0 9856 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_333
timestamp 1612251222
transform 1 0 9840 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_502
timestamp 1612251222
transform 1 0 9674 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_502
timestamp 1612251222
transform 1 0 9658 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_502
timestamp 1612251222
transform 1 0 9642 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_502
timestamp 1612251222
transform 1 0 9626 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_237
timestamp 1612251222
transform 1 0 9460 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_237
timestamp 1612251222
transform 1 0 9444 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_237
timestamp 1612251222
transform 1 0 9428 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_237
timestamp 1612251222
transform 1 0 9412 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_237
timestamp 1612251222
transform 1 0 9396 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_253
timestamp 1612251222
transform -1 0 9396 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_253
timestamp 1612251222
transform -1 0 9230 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_253
timestamp 1612251222
transform -1 0 9214 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_253
timestamp 1612251222
transform -1 0 9198 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_253
timestamp 1612251222
transform -1 0 9182 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_341
timestamp 1612251222
transform 1 0 9000 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_341
timestamp 1612251222
transform 1 0 8984 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_341
timestamp 1612251222
transform 1 0 8968 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_341
timestamp 1612251222
transform 1 0 8952 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_254
timestamp 1612251222
transform 1 0 8786 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_254
timestamp 1612251222
transform 1 0 8770 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_254
timestamp 1612251222
transform 1 0 8754 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_254
timestamp 1612251222
transform 1 0 8738 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_483
timestamp 1612251222
transform -1 0 8738 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_483
timestamp 1612251222
transform -1 0 8572 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_483
timestamp 1612251222
transform -1 0 8556 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_483
timestamp 1612251222
transform -1 0 8540 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_260
timestamp 1612251222
transform -1 0 8524 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_260
timestamp 1612251222
transform -1 0 8358 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_260
timestamp 1612251222
transform -1 0 8342 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_260
timestamp 1612251222
transform -1 0 8326 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_205
timestamp 1612251222
transform 1 0 8144 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_205
timestamp 1612251222
transform 1 0 8128 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_205
timestamp 1612251222
transform 1 0 8112 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_205
timestamp 1612251222
transform 1 0 8096 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_344
timestamp 1612251222
transform -1 0 8096 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_344
timestamp 1612251222
transform -1 0 7930 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_344
timestamp 1612251222
transform -1 0 7914 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_344
timestamp 1612251222
transform -1 0 7898 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_256
timestamp 1612251222
transform 1 0 7716 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_256
timestamp 1612251222
transform 1 0 7700 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_256
timestamp 1612251222
transform 1 0 7684 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_256
timestamp 1612251222
transform 1 0 7668 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_256
timestamp 1612251222
transform 1 0 7652 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_65
timestamp 1612251222
transform 1 0 7486 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_65
timestamp 1612251222
transform 1 0 7470 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_65
timestamp 1612251222
transform 1 0 7454 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_65
timestamp 1612251222
transform 1 0 7438 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_65
timestamp 1612251222
transform 1 0 7422 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_246
timestamp 1612251222
transform 1 0 7256 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_246
timestamp 1612251222
transform 1 0 7240 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_246
timestamp 1612251222
transform 1 0 7224 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_246
timestamp 1612251222
transform 1 0 7208 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_246
timestamp 1612251222
transform 1 0 7192 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_204
timestamp 1612251222
transform 1 0 7026 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_204
timestamp 1612251222
transform 1 0 7010 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_204
timestamp 1612251222
transform 1 0 6994 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_204
timestamp 1612251222
transform 1 0 6978 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_81
timestamp 1612251222
transform 1 0 6812 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_81
timestamp 1612251222
transform 1 0 6796 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_81
timestamp 1612251222
transform 1 0 6780 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_81
timestamp 1612251222
transform 1 0 6764 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_81
timestamp 1612251222
transform 1 0 6748 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_63
timestamp 1612251222
transform 1 0 6582 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_63
timestamp 1612251222
transform 1 0 6566 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_63
timestamp 1612251222
transform 1 0 6550 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_63
timestamp 1612251222
transform 1 0 6534 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_63
timestamp 1612251222
transform 1 0 6518 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_73
timestamp 1612251222
transform -1 0 6518 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_73
timestamp 1612251222
transform -1 0 6352 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_73
timestamp 1612251222
transform -1 0 6336 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_73
timestamp 1612251222
transform -1 0 6320 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_73
timestamp 1612251222
transform -1 0 6304 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_548
timestamp 1612251222
transform 1 0 6122 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_548
timestamp 1612251222
transform 1 0 6106 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_548
timestamp 1612251222
transform 1 0 6090 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_548
timestamp 1612251222
transform 1 0 6074 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_143
timestamp 1612251222
transform 1 0 5908 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_143
timestamp 1612251222
transform 1 0 5892 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_143
timestamp 1612251222
transform 1 0 5876 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_143
timestamp 1612251222
transform 1 0 5860 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_143
timestamp 1612251222
transform 1 0 5844 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_529
timestamp 1612251222
transform 1 0 5678 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_529
timestamp 1612251222
transform 1 0 5662 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_529
timestamp 1612251222
transform 1 0 5646 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_529
timestamp 1612251222
transform 1 0 5630 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_529
timestamp 1612251222
transform 1 0 5614 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_615
timestamp 1612251222
transform 1 0 5448 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_615
timestamp 1612251222
transform 1 0 5432 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_615
timestamp 1612251222
transform 1 0 5416 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_615
timestamp 1612251222
transform 1 0 5400 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_615
timestamp 1612251222
transform 1 0 5384 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_28
timestamp 1612251222
transform 1 0 5218 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_28
timestamp 1612251222
transform 1 0 5202 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_28
timestamp 1612251222
transform 1 0 5186 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_28
timestamp 1612251222
transform 1 0 5170 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_28
timestamp 1612251222
transform 1 0 5154 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_376
timestamp 1612251222
transform -1 0 5154 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_376
timestamp 1612251222
transform -1 0 4988 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_376
timestamp 1612251222
transform -1 0 4972 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_376
timestamp 1612251222
transform -1 0 4956 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_159
timestamp 1612251222
transform 1 0 4774 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_159
timestamp 1612251222
transform 1 0 4758 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_159
timestamp 1612251222
transform 1 0 4742 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_159
timestamp 1612251222
transform 1 0 4726 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_27
timestamp 1612251222
transform 1 0 4560 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_POR2X1_27
timestamp 1612251222
transform 1 0 4544 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_POR2X1_27
timestamp 1612251222
transform 1 0 4528 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_27
timestamp 1612251222
transform 1 0 4512 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_27
timestamp 1612251222
transform 1 0 4496 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_10
timestamp 1612251222
transform 1 0 4330 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_POR2X1_10
timestamp 1612251222
transform 1 0 4314 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_POR2X1_10
timestamp 1612251222
transform 1 0 4298 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_10
timestamp 1612251222
transform 1 0 4282 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_10
timestamp 1612251222
transform 1 0 4266 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_63
timestamp 1612251222
transform -1 0 4266 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_POR2X1_63
timestamp 1612251222
transform -1 0 4100 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_POR2X1_63
timestamp 1612251222
transform -1 0 4084 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_63
timestamp 1612251222
transform -1 0 4068 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_63
timestamp 1612251222
transform -1 0 4052 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_813
timestamp 1612251222
transform 1 0 3870 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_813
timestamp 1612251222
transform 1 0 3854 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_813
timestamp 1612251222
transform 1 0 3838 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_813
timestamp 1612251222
transform 1 0 3822 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_235
timestamp 1612251222
transform -1 0 3822 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_235
timestamp 1612251222
transform -1 0 3656 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_235
timestamp 1612251222
transform -1 0 3640 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_235
timestamp 1612251222
transform -1 0 3624 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_230
timestamp 1612251222
transform -1 0 3608 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_230
timestamp 1612251222
transform -1 0 3442 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_230
timestamp 1612251222
transform -1 0 3426 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_230
timestamp 1612251222
transform -1 0 3410 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_231
timestamp 1612251222
transform -1 0 3394 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_231
timestamp 1612251222
transform -1 0 3228 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_231
timestamp 1612251222
transform -1 0 3212 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_231
timestamp 1612251222
transform -1 0 3196 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_231
timestamp 1612251222
transform -1 0 3180 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_641
timestamp 1612251222
transform 1 0 2998 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_641
timestamp 1612251222
transform 1 0 2982 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_641
timestamp 1612251222
transform 1 0 2966 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_641
timestamp 1612251222
transform 1 0 2950 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_641
timestamp 1612251222
transform 1 0 2934 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_734
timestamp 1612251222
transform -1 0 2934 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_734
timestamp 1612251222
transform -1 0 2768 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_734
timestamp 1612251222
transform -1 0 2752 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_734
timestamp 1612251222
transform -1 0 2736 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_734
timestamp 1612251222
transform -1 0 2720 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_406
timestamp 1612251222
transform 1 0 2538 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_406
timestamp 1612251222
transform 1 0 2522 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_406
timestamp 1612251222
transform 1 0 2506 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_406
timestamp 1612251222
transform 1 0 2490 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_405
timestamp 1612251222
transform 1 0 2324 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_405
timestamp 1612251222
transform 1 0 2308 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_405
timestamp 1612251222
transform 1 0 2292 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_405
timestamp 1612251222
transform 1 0 2276 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_405
timestamp 1612251222
transform 1 0 2260 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_198
timestamp 1612251222
transform 1 0 2094 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_198
timestamp 1612251222
transform 1 0 2078 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_198
timestamp 1612251222
transform 1 0 2062 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_198
timestamp 1612251222
transform 1 0 2046 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_198
timestamp 1612251222
transform 1 0 2030 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_57
timestamp 1612251222
transform 1 0 1864 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_POR2X1_57
timestamp 1612251222
transform 1 0 1848 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_POR2X1_57
timestamp 1612251222
transform 1 0 1832 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_57
timestamp 1612251222
transform 1 0 1816 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_57
timestamp 1612251222
transform 1 0 1800 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_737
timestamp 1612251222
transform 1 0 1634 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_737
timestamp 1612251222
transform 1 0 1618 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_737
timestamp 1612251222
transform 1 0 1602 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_737
timestamp 1612251222
transform 1 0 1586 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_737
timestamp 1612251222
transform 1 0 1570 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_733
timestamp 1612251222
transform 1 0 1404 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_733
timestamp 1612251222
transform 1 0 1388 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_733
timestamp 1612251222
transform 1 0 1372 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_733
timestamp 1612251222
transform 1 0 1356 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_733
timestamp 1612251222
transform 1 0 1340 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_193
timestamp 1612251222
transform 1 0 1174 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_193
timestamp 1612251222
transform 1 0 1158 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_193
timestamp 1612251222
transform 1 0 1142 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_193
timestamp 1612251222
transform 1 0 1126 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_193
timestamp 1612251222
transform 1 0 1110 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_13
timestamp 1612251222
transform -1 0 1110 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_POR2X1_13
timestamp 1612251222
transform -1 0 944 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_POR2X1_13
timestamp 1612251222
transform -1 0 928 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_13
timestamp 1612251222
transform -1 0 912 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_13
timestamp 1612251222
transform -1 0 896 0 -1 5810
box -4 -6 20 206
use PAND2X1  PAND2X1_643
timestamp 1612251222
transform 1 0 714 0 -1 5810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_643
timestamp 1612251222
transform 1 0 698 0 -1 5810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_643
timestamp 1612251222
transform 1 0 682 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_643
timestamp 1612251222
transform 1 0 666 0 -1 5810
box -4 -6 20 206
use FILL  FILL_PAND2X1_643
timestamp 1612251222
transform 1 0 650 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_760
timestamp 1612251222
transform 1 0 484 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_760
timestamp 1612251222
transform 1 0 468 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_760
timestamp 1612251222
transform 1 0 452 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_760
timestamp 1612251222
transform 1 0 436 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_281
timestamp 1612251222
transform -1 0 436 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_281
timestamp 1612251222
transform -1 0 270 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_281
timestamp 1612251222
transform -1 0 254 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_281
timestamp 1612251222
transform -1 0 238 0 -1 5810
box -4 -6 20 206
use POR2X1  POR2X1_282
timestamp 1612251222
transform -1 0 222 0 -1 5810
box -4 -6 170 206
use FILL  FILL1_POR2X1_282
timestamp 1612251222
transform -1 0 56 0 -1 5810
box -4 -6 20 206
use FILL  FILL0_POR2X1_282
timestamp 1612251222
transform -1 0 40 0 -1 5810
box -4 -6 20 206
use FILL  FILL_POR2X1_282
timestamp 1612251222
transform -1 0 24 0 -1 5810
box -4 -6 20 206
use FILL  FILL_28_12
timestamp 1612251222
transform 1 0 10246 0 1 5410
box -4 -6 20 206
use FILL  FILL_28_11
timestamp 1612251222
transform 1 0 10230 0 1 5410
box -4 -6 20 206
use FILL  FILL_28_10
timestamp 1612251222
transform 1 0 10214 0 1 5410
box -4 -6 20 206
use FILL  FILL_28_9
timestamp 1612251222
transform 1 0 10198 0 1 5410
box -4 -6 20 206
use FILL  FILL_28_8
timestamp 1612251222
transform 1 0 10182 0 1 5410
box -4 -6 20 206
use FILL  FILL_28_7
timestamp 1612251222
transform 1 0 10166 0 1 5410
box -4 -6 20 206
use FILL  FILL_28_6
timestamp 1612251222
transform 1 0 10150 0 1 5410
box -4 -6 20 206
use FILL  FILL_28_5
timestamp 1612251222
transform 1 0 10134 0 1 5410
box -4 -6 20 206
use FILL  FILL_28_4
timestamp 1612251222
transform 1 0 10118 0 1 5410
box -4 -6 20 206
use FILL  FILL_28_3
timestamp 1612251222
transform 1 0 10102 0 1 5410
box -4 -6 20 206
use FILL  FILL_28_2
timestamp 1612251222
transform 1 0 10086 0 1 5410
box -4 -6 20 206
use FILL  FILL_28_1
timestamp 1612251222
transform 1 0 10070 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_785
timestamp 1612251222
transform -1 0 10070 0 1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_785
timestamp 1612251222
transform -1 0 9904 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_785
timestamp 1612251222
transform -1 0 9888 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_785
timestamp 1612251222
transform -1 0 9872 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_853
timestamp 1612251222
transform -1 0 9856 0 1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_853
timestamp 1612251222
transform -1 0 9690 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_853
timestamp 1612251222
transform -1 0 9674 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_853
timestamp 1612251222
transform -1 0 9658 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_857
timestamp 1612251222
transform -1 0 9642 0 1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_857
timestamp 1612251222
transform -1 0 9476 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_857
timestamp 1612251222
transform -1 0 9460 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_857
timestamp 1612251222
transform -1 0 9444 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_230
timestamp 1612251222
transform -1 0 9428 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_230
timestamp 1612251222
transform -1 0 9262 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_230
timestamp 1612251222
transform -1 0 9246 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_230
timestamp 1612251222
transform -1 0 9230 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_230
timestamp 1612251222
transform -1 0 9214 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_231
timestamp 1612251222
transform -1 0 9198 0 1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_231
timestamp 1612251222
transform -1 0 9032 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_231
timestamp 1612251222
transform -1 0 9016 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_231
timestamp 1612251222
transform -1 0 9000 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_13
timestamp 1612251222
transform -1 0 8984 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_13
timestamp 1612251222
transform -1 0 8818 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_13
timestamp 1612251222
transform -1 0 8802 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_13
timestamp 1612251222
transform -1 0 8786 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_13
timestamp 1612251222
transform -1 0 8770 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_795
timestamp 1612251222
transform -1 0 8754 0 1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_795
timestamp 1612251222
transform -1 0 8588 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_795
timestamp 1612251222
transform -1 0 8572 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_795
timestamp 1612251222
transform -1 0 8556 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_702
timestamp 1612251222
transform 1 0 8374 0 1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_702
timestamp 1612251222
transform 1 0 8358 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_702
timestamp 1612251222
transform 1 0 8342 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_702
timestamp 1612251222
transform 1 0 8326 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_48
timestamp 1612251222
transform 1 0 8160 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_48
timestamp 1612251222
transform 1 0 8144 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_48
timestamp 1612251222
transform 1 0 8128 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_48
timestamp 1612251222
transform 1 0 8112 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_48
timestamp 1612251222
transform 1 0 8096 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_482
timestamp 1612251222
transform 1 0 7930 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_482
timestamp 1612251222
transform 1 0 7914 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_482
timestamp 1612251222
transform 1 0 7898 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_482
timestamp 1612251222
transform 1 0 7882 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_482
timestamp 1612251222
transform 1 0 7866 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_833
timestamp 1612251222
transform 1 0 7700 0 1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_833
timestamp 1612251222
transform 1 0 7684 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_833
timestamp 1612251222
transform 1 0 7668 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_833
timestamp 1612251222
transform 1 0 7652 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_255
timestamp 1612251222
transform 1 0 7486 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_255
timestamp 1612251222
transform 1 0 7470 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_255
timestamp 1612251222
transform 1 0 7454 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_255
timestamp 1612251222
transform 1 0 7438 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_255
timestamp 1612251222
transform 1 0 7422 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_150
timestamp 1612251222
transform -1 0 7422 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_150
timestamp 1612251222
transform -1 0 7256 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_150
timestamp 1612251222
transform -1 0 7240 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_150
timestamp 1612251222
transform -1 0 7224 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_150
timestamp 1612251222
transform -1 0 7208 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_495
timestamp 1612251222
transform 1 0 7026 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_495
timestamp 1612251222
transform 1 0 7010 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_495
timestamp 1612251222
transform 1 0 6994 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_495
timestamp 1612251222
transform 1 0 6978 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_495
timestamp 1612251222
transform 1 0 6962 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_786
timestamp 1612251222
transform 1 0 6796 0 1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_786
timestamp 1612251222
transform 1 0 6780 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_786
timestamp 1612251222
transform 1 0 6764 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_786
timestamp 1612251222
transform 1 0 6748 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_262
timestamp 1612251222
transform -1 0 6748 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_262
timestamp 1612251222
transform -1 0 6582 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_262
timestamp 1612251222
transform -1 0 6566 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_262
timestamp 1612251222
transform -1 0 6550 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_262
timestamp 1612251222
transform -1 0 6534 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_266
timestamp 1612251222
transform 1 0 6352 0 1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_266
timestamp 1612251222
transform 1 0 6336 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_266
timestamp 1612251222
transform 1 0 6320 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_266
timestamp 1612251222
transform 1 0 6304 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_549
timestamp 1612251222
transform -1 0 6304 0 1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_549
timestamp 1612251222
transform -1 0 6138 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_549
timestamp 1612251222
transform -1 0 6122 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_549
timestamp 1612251222
transform -1 0 6106 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_547
timestamp 1612251222
transform -1 0 6090 0 1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_547
timestamp 1612251222
transform -1 0 5924 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_547
timestamp 1612251222
transform -1 0 5908 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_547
timestamp 1612251222
transform -1 0 5892 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_813
timestamp 1612251222
transform 1 0 5710 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_813
timestamp 1612251222
transform 1 0 5694 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_813
timestamp 1612251222
transform 1 0 5678 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_813
timestamp 1612251222
transform 1 0 5662 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_813
timestamp 1612251222
transform 1 0 5646 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_263
timestamp 1612251222
transform 1 0 5480 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_263
timestamp 1612251222
transform 1 0 5464 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_263
timestamp 1612251222
transform 1 0 5448 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_263
timestamp 1612251222
transform 1 0 5432 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_263
timestamp 1612251222
transform 1 0 5416 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_614
timestamp 1612251222
transform -1 0 5416 0 1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_614
timestamp 1612251222
transform -1 0 5250 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_614
timestamp 1612251222
transform -1 0 5234 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_614
timestamp 1612251222
transform -1 0 5218 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_749
timestamp 1612251222
transform -1 0 5202 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_749
timestamp 1612251222
transform -1 0 5036 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_749
timestamp 1612251222
transform -1 0 5020 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_749
timestamp 1612251222
transform -1 0 5004 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_749
timestamp 1612251222
transform -1 0 4988 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_87
timestamp 1612251222
transform 1 0 4806 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_87
timestamp 1612251222
transform 1 0 4790 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_87
timestamp 1612251222
transform 1 0 4774 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_87
timestamp 1612251222
transform 1 0 4758 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_87
timestamp 1612251222
transform 1 0 4742 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_68
timestamp 1612251222
transform 1 0 4576 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_68
timestamp 1612251222
transform 1 0 4560 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_68
timestamp 1612251222
transform 1 0 4544 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_68
timestamp 1612251222
transform 1 0 4528 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_68
timestamp 1612251222
transform 1 0 4512 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_62
timestamp 1612251222
transform -1 0 4512 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_62
timestamp 1612251222
transform -1 0 4346 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_62
timestamp 1612251222
transform -1 0 4330 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_62
timestamp 1612251222
transform -1 0 4314 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_62
timestamp 1612251222
transform -1 0 4298 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_143
timestamp 1612251222
transform -1 0 4282 0 1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_143
timestamp 1612251222
transform -1 0 4116 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_143
timestamp 1612251222
transform -1 0 4100 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_143
timestamp 1612251222
transform -1 0 4084 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_65
timestamp 1612251222
transform 1 0 3902 0 1 5410
box -4 -6 170 206
use FILL  FILL2_POR2X1_65
timestamp 1612251222
transform 1 0 3886 0 1 5410
box -4 -6 20 206
use FILL  FILL1_POR2X1_65
timestamp 1612251222
transform 1 0 3870 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_65
timestamp 1612251222
transform 1 0 3854 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_65
timestamp 1612251222
transform 1 0 3838 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_73
timestamp 1612251222
transform -1 0 3838 0 1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_73
timestamp 1612251222
transform -1 0 3672 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_73
timestamp 1612251222
transform -1 0 3656 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_73
timestamp 1612251222
transform -1 0 3640 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_86
timestamp 1612251222
transform 1 0 3458 0 1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_86
timestamp 1612251222
transform 1 0 3442 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_86
timestamp 1612251222
transform 1 0 3426 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_86
timestamp 1612251222
transform 1 0 3410 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_206
timestamp 1612251222
transform -1 0 3410 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_206
timestamp 1612251222
transform -1 0 3244 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_206
timestamp 1612251222
transform -1 0 3228 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_206
timestamp 1612251222
transform -1 0 3212 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_206
timestamp 1612251222
transform -1 0 3196 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_490
timestamp 1612251222
transform -1 0 3180 0 1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_490
timestamp 1612251222
transform -1 0 3014 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_490
timestamp 1612251222
transform -1 0 2998 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_490
timestamp 1612251222
transform -1 0 2982 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_262
timestamp 1612251222
transform -1 0 2966 0 1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_262
timestamp 1612251222
transform -1 0 2800 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_262
timestamp 1612251222
transform -1 0 2784 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_262
timestamp 1612251222
transform -1 0 2768 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_266
timestamp 1612251222
transform -1 0 2752 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_266
timestamp 1612251222
transform -1 0 2586 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_266
timestamp 1612251222
transform -1 0 2570 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_266
timestamp 1612251222
transform -1 0 2554 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_266
timestamp 1612251222
transform -1 0 2538 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_267
timestamp 1612251222
transform -1 0 2522 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_267
timestamp 1612251222
transform -1 0 2356 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_267
timestamp 1612251222
transform -1 0 2340 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_267
timestamp 1612251222
transform -1 0 2324 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_267
timestamp 1612251222
transform -1 0 2308 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_52
timestamp 1612251222
transform 1 0 2126 0 1 5410
box -4 -6 170 206
use FILL  FILL2_POR2X1_52
timestamp 1612251222
transform 1 0 2110 0 1 5410
box -4 -6 20 206
use FILL  FILL1_POR2X1_52
timestamp 1612251222
transform 1 0 2094 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_52
timestamp 1612251222
transform 1 0 2078 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_52
timestamp 1612251222
transform 1 0 2062 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_723
timestamp 1612251222
transform -1 0 2062 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_723
timestamp 1612251222
transform -1 0 1896 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_723
timestamp 1612251222
transform -1 0 1880 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_723
timestamp 1612251222
transform -1 0 1864 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_723
timestamp 1612251222
transform -1 0 1848 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_7
timestamp 1612251222
transform -1 0 1832 0 1 5410
box -4 -6 170 206
use FILL  FILL2_POR2X1_7
timestamp 1612251222
transform -1 0 1666 0 1 5410
box -4 -6 20 206
use FILL  FILL1_POR2X1_7
timestamp 1612251222
transform -1 0 1650 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_7
timestamp 1612251222
transform -1 0 1634 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_7
timestamp 1612251222
transform -1 0 1618 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_215
timestamp 1612251222
transform -1 0 1602 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_215
timestamp 1612251222
transform -1 0 1436 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_215
timestamp 1612251222
transform -1 0 1420 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_215
timestamp 1612251222
transform -1 0 1404 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_215
timestamp 1612251222
transform -1 0 1388 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_219
timestamp 1612251222
transform -1 0 1372 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_219
timestamp 1612251222
transform -1 0 1206 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_219
timestamp 1612251222
transform -1 0 1190 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_219
timestamp 1612251222
transform -1 0 1174 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_219
timestamp 1612251222
transform -1 0 1158 0 1 5410
box -4 -6 20 206
use POR2X1  POR2X1_536
timestamp 1612251222
transform 1 0 976 0 1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_536
timestamp 1612251222
transform 1 0 960 0 1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_536
timestamp 1612251222
transform 1 0 944 0 1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_536
timestamp 1612251222
transform 1 0 928 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_222
timestamp 1612251222
transform -1 0 928 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_222
timestamp 1612251222
transform -1 0 762 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_222
timestamp 1612251222
transform -1 0 746 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_222
timestamp 1612251222
transform -1 0 730 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_222
timestamp 1612251222
transform -1 0 714 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_538
timestamp 1612251222
transform -1 0 698 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_538
timestamp 1612251222
transform -1 0 532 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_538
timestamp 1612251222
transform -1 0 516 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_538
timestamp 1612251222
transform -1 0 500 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_538
timestamp 1612251222
transform -1 0 484 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_539
timestamp 1612251222
transform -1 0 468 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_539
timestamp 1612251222
transform -1 0 302 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_539
timestamp 1612251222
transform -1 0 286 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_539
timestamp 1612251222
transform -1 0 270 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_539
timestamp 1612251222
transform -1 0 254 0 1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_285
timestamp 1612251222
transform -1 0 238 0 1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_285
timestamp 1612251222
transform -1 0 72 0 1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_285
timestamp 1612251222
transform -1 0 56 0 1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_285
timestamp 1612251222
transform -1 0 40 0 1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_285
timestamp 1612251222
transform -1 0 24 0 1 5410
box -4 -6 20 206
use FILL  FILL_27_1
timestamp 1612251222
transform -1 0 10262 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_164
timestamp 1612251222
transform 1 0 10080 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_164
timestamp 1612251222
transform 1 0 10064 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_164
timestamp 1612251222
transform 1 0 10048 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_164
timestamp 1612251222
transform 1 0 10032 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_164
timestamp 1612251222
transform 1 0 10016 0 -1 5410
box -4 -6 20 206
use POR2X1  POR2X1_775
timestamp 1612251222
transform 1 0 9850 0 -1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_775
timestamp 1612251222
transform 1 0 9834 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_775
timestamp 1612251222
transform 1 0 9818 0 -1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_775
timestamp 1612251222
transform 1 0 9802 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_109
timestamp 1612251222
transform -1 0 9802 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_109
timestamp 1612251222
transform -1 0 9636 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_109
timestamp 1612251222
transform -1 0 9620 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_109
timestamp 1612251222
transform -1 0 9604 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_109
timestamp 1612251222
transform -1 0 9588 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_173
timestamp 1612251222
transform -1 0 9572 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_173
timestamp 1612251222
transform -1 0 9406 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_173
timestamp 1612251222
transform -1 0 9390 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_173
timestamp 1612251222
transform -1 0 9374 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_173
timestamp 1612251222
transform -1 0 9358 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_229
timestamp 1612251222
transform 1 0 9176 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_229
timestamp 1612251222
transform 1 0 9160 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_229
timestamp 1612251222
transform 1 0 9144 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_229
timestamp 1612251222
transform 1 0 9128 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_229
timestamp 1612251222
transform 1 0 9112 0 -1 5410
box -4 -6 20 206
use POR2X1  POR2X1_332
timestamp 1612251222
transform -1 0 9112 0 -1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_332
timestamp 1612251222
transform -1 0 8946 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_332
timestamp 1612251222
transform -1 0 8930 0 -1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_332
timestamp 1612251222
transform -1 0 8914 0 -1 5410
box -4 -6 20 206
use POR2X1  POR2X1_112
timestamp 1612251222
transform 1 0 8732 0 -1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_112
timestamp 1612251222
transform 1 0 8716 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_112
timestamp 1612251222
transform 1 0 8700 0 -1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_112
timestamp 1612251222
transform 1 0 8684 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_135
timestamp 1612251222
transform -1 0 8684 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_135
timestamp 1612251222
transform -1 0 8518 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_135
timestamp 1612251222
transform -1 0 8502 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_135
timestamp 1612251222
transform -1 0 8486 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_135
timestamp 1612251222
transform -1 0 8470 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_111
timestamp 1612251222
transform -1 0 8454 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_111
timestamp 1612251222
transform -1 0 8288 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_111
timestamp 1612251222
transform -1 0 8272 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_111
timestamp 1612251222
transform -1 0 8256 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_111
timestamp 1612251222
transform -1 0 8240 0 -1 5410
box -4 -6 20 206
use POR2X1  POR2X1_203
timestamp 1612251222
transform -1 0 8224 0 -1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_203
timestamp 1612251222
transform -1 0 8058 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_203
timestamp 1612251222
transform -1 0 8042 0 -1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_203
timestamp 1612251222
transform -1 0 8026 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_72
timestamp 1612251222
transform 1 0 7844 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_72
timestamp 1612251222
transform 1 0 7828 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_72
timestamp 1612251222
transform 1 0 7812 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_72
timestamp 1612251222
transform 1 0 7796 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_72
timestamp 1612251222
transform 1 0 7780 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_71
timestamp 1612251222
transform 1 0 7614 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_71
timestamp 1612251222
transform 1 0 7598 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_71
timestamp 1612251222
transform 1 0 7582 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_71
timestamp 1612251222
transform 1 0 7566 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_71
timestamp 1612251222
transform 1 0 7550 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_245
timestamp 1612251222
transform -1 0 7550 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_245
timestamp 1612251222
transform -1 0 7384 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_245
timestamp 1612251222
transform -1 0 7368 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_245
timestamp 1612251222
transform -1 0 7352 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_245
timestamp 1612251222
transform -1 0 7336 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_46
timestamp 1612251222
transform 1 0 7154 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_46
timestamp 1612251222
transform 1 0 7138 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_46
timestamp 1612251222
transform 1 0 7122 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_46
timestamp 1612251222
transform 1 0 7106 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_46
timestamp 1612251222
transform 1 0 7090 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_527
timestamp 1612251222
transform -1 0 7090 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_527
timestamp 1612251222
transform -1 0 6924 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_527
timestamp 1612251222
transform -1 0 6908 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_527
timestamp 1612251222
transform -1 0 6892 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_527
timestamp 1612251222
transform -1 0 6876 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_80
timestamp 1612251222
transform 1 0 6694 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_80
timestamp 1612251222
transform 1 0 6678 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_80
timestamp 1612251222
transform 1 0 6662 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_80
timestamp 1612251222
transform 1 0 6646 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_80
timestamp 1612251222
transform 1 0 6630 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_42
timestamp 1612251222
transform 1 0 6464 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_42
timestamp 1612251222
transform 1 0 6448 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_42
timestamp 1612251222
transform 1 0 6432 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_42
timestamp 1612251222
transform 1 0 6416 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_42
timestamp 1612251222
transform 1 0 6400 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_531
timestamp 1612251222
transform -1 0 6400 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_531
timestamp 1612251222
transform -1 0 6234 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_531
timestamp 1612251222
transform -1 0 6218 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_531
timestamp 1612251222
transform -1 0 6202 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_531
timestamp 1612251222
transform -1 0 6186 0 -1 5410
box -4 -6 20 206
use POR2X1  POR2X1_6
timestamp 1612251222
transform -1 0 6170 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_POR2X1_6
timestamp 1612251222
transform -1 0 6004 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_POR2X1_6
timestamp 1612251222
transform -1 0 5988 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_6
timestamp 1612251222
transform -1 0 5972 0 -1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_6
timestamp 1612251222
transform -1 0 5956 0 -1 5410
box -4 -6 20 206
use POR2X1  POR2X1_845
timestamp 1612251222
transform -1 0 5940 0 -1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_845
timestamp 1612251222
transform -1 0 5774 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_845
timestamp 1612251222
transform -1 0 5758 0 -1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_845
timestamp 1612251222
transform -1 0 5742 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_202
timestamp 1612251222
transform -1 0 5726 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_202
timestamp 1612251222
transform -1 0 5560 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_202
timestamp 1612251222
transform -1 0 5544 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_202
timestamp 1612251222
transform -1 0 5528 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_202
timestamp 1612251222
transform -1 0 5512 0 -1 5410
box -4 -6 20 206
use POR2X1  POR2X1_69
timestamp 1612251222
transform 1 0 5330 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_POR2X1_69
timestamp 1612251222
transform 1 0 5314 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_POR2X1_69
timestamp 1612251222
transform 1 0 5298 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_69
timestamp 1612251222
transform 1 0 5282 0 -1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_69
timestamp 1612251222
transform 1 0 5266 0 -1 5410
box -4 -6 20 206
use POR2X1  POR2X1_15
timestamp 1612251222
transform -1 0 5266 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_POR2X1_15
timestamp 1612251222
transform -1 0 5100 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_POR2X1_15
timestamp 1612251222
transform -1 0 5084 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_15
timestamp 1612251222
transform -1 0 5068 0 -1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_15
timestamp 1612251222
transform -1 0 5052 0 -1 5410
box -4 -6 20 206
use POR2X1  POR2X1_88
timestamp 1612251222
transform -1 0 5036 0 -1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_88
timestamp 1612251222
transform -1 0 4870 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_88
timestamp 1612251222
transform -1 0 4854 0 -1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_88
timestamp 1612251222
transform -1 0 4838 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_340
timestamp 1612251222
transform -1 0 4822 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_340
timestamp 1612251222
transform -1 0 4656 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_340
timestamp 1612251222
transform -1 0 4640 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_340
timestamp 1612251222
transform -1 0 4624 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_340
timestamp 1612251222
transform -1 0 4608 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_350
timestamp 1612251222
transform -1 0 4592 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_350
timestamp 1612251222
transform -1 0 4426 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_350
timestamp 1612251222
transform -1 0 4410 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_350
timestamp 1612251222
transform -1 0 4394 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_350
timestamp 1612251222
transform -1 0 4378 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_341
timestamp 1612251222
transform 1 0 4196 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_341
timestamp 1612251222
transform 1 0 4180 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_341
timestamp 1612251222
transform 1 0 4164 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_341
timestamp 1612251222
transform 1 0 4148 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_341
timestamp 1612251222
transform 1 0 4132 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_201
timestamp 1612251222
transform -1 0 4132 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_201
timestamp 1612251222
transform -1 0 3966 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_201
timestamp 1612251222
transform -1 0 3950 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_201
timestamp 1612251222
transform -1 0 3934 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_201
timestamp 1612251222
transform -1 0 3918 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_100
timestamp 1612251222
transform -1 0 3902 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_100
timestamp 1612251222
transform -1 0 3736 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_100
timestamp 1612251222
transform -1 0 3720 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_100
timestamp 1612251222
transform -1 0 3704 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_100
timestamp 1612251222
transform -1 0 3688 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_101
timestamp 1612251222
transform -1 0 3672 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_101
timestamp 1612251222
transform -1 0 3506 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_101
timestamp 1612251222
transform -1 0 3490 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_101
timestamp 1612251222
transform -1 0 3474 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_101
timestamp 1612251222
transform -1 0 3458 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_358
timestamp 1612251222
transform -1 0 3442 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_358
timestamp 1612251222
transform -1 0 3276 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_358
timestamp 1612251222
transform -1 0 3260 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_358
timestamp 1612251222
transform -1 0 3244 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_358
timestamp 1612251222
transform -1 0 3228 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_197
timestamp 1612251222
transform -1 0 3212 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_197
timestamp 1612251222
transform -1 0 3046 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_197
timestamp 1612251222
transform -1 0 3030 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_197
timestamp 1612251222
transform -1 0 3014 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_197
timestamp 1612251222
transform -1 0 2998 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_228
timestamp 1612251222
transform 1 0 2816 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_228
timestamp 1612251222
transform 1 0 2800 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_228
timestamp 1612251222
transform 1 0 2784 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_228
timestamp 1612251222
transform 1 0 2768 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_228
timestamp 1612251222
transform 1 0 2752 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_716
timestamp 1612251222
transform -1 0 2752 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_716
timestamp 1612251222
transform -1 0 2586 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_716
timestamp 1612251222
transform -1 0 2570 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_716
timestamp 1612251222
transform -1 0 2554 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_716
timestamp 1612251222
transform -1 0 2538 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_572
timestamp 1612251222
transform 1 0 2356 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_572
timestamp 1612251222
transform 1 0 2340 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_572
timestamp 1612251222
transform 1 0 2324 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_572
timestamp 1612251222
transform 1 0 2308 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_572
timestamp 1612251222
transform 1 0 2292 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_217
timestamp 1612251222
transform -1 0 2292 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_217
timestamp 1612251222
transform -1 0 2126 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_217
timestamp 1612251222
transform -1 0 2110 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_217
timestamp 1612251222
transform -1 0 2094 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_217
timestamp 1612251222
transform -1 0 2078 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_216
timestamp 1612251222
transform -1 0 2062 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_216
timestamp 1612251222
transform -1 0 1896 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_216
timestamp 1612251222
transform -1 0 1880 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_216
timestamp 1612251222
transform -1 0 1864 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_216
timestamp 1612251222
transform -1 0 1848 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_218
timestamp 1612251222
transform -1 0 1832 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_218
timestamp 1612251222
transform -1 0 1666 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_218
timestamp 1612251222
transform -1 0 1650 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_218
timestamp 1612251222
transform -1 0 1634 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_218
timestamp 1612251222
transform -1 0 1618 0 -1 5410
box -4 -6 20 206
use POR2X1  POR2X1_385
timestamp 1612251222
transform -1 0 1602 0 -1 5410
box -4 -6 170 206
use FILL  FILL1_POR2X1_385
timestamp 1612251222
transform -1 0 1436 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_POR2X1_385
timestamp 1612251222
transform -1 0 1420 0 -1 5410
box -4 -6 20 206
use FILL  FILL_POR2X1_385
timestamp 1612251222
transform -1 0 1404 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_593
timestamp 1612251222
transform -1 0 1388 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_593
timestamp 1612251222
transform -1 0 1222 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_593
timestamp 1612251222
transform -1 0 1206 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_593
timestamp 1612251222
transform -1 0 1190 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_593
timestamp 1612251222
transform -1 0 1174 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_537
timestamp 1612251222
transform -1 0 1158 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_537
timestamp 1612251222
transform -1 0 992 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_537
timestamp 1612251222
transform -1 0 976 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_537
timestamp 1612251222
transform -1 0 960 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_537
timestamp 1612251222
transform -1 0 944 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_799
timestamp 1612251222
transform -1 0 928 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_799
timestamp 1612251222
transform -1 0 762 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_799
timestamp 1612251222
transform -1 0 746 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_799
timestamp 1612251222
transform -1 0 730 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_799
timestamp 1612251222
transform -1 0 714 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_802
timestamp 1612251222
transform -1 0 698 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_802
timestamp 1612251222
transform -1 0 532 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_802
timestamp 1612251222
transform -1 0 516 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_802
timestamp 1612251222
transform -1 0 500 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_802
timestamp 1612251222
transform -1 0 484 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_809
timestamp 1612251222
transform 1 0 302 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_809
timestamp 1612251222
transform 1 0 286 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_809
timestamp 1612251222
transform 1 0 270 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_809
timestamp 1612251222
transform 1 0 254 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_809
timestamp 1612251222
transform 1 0 238 0 -1 5410
box -4 -6 20 206
use PAND2X1  PAND2X1_567
timestamp 1612251222
transform -1 0 238 0 -1 5410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_567
timestamp 1612251222
transform -1 0 72 0 -1 5410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_567
timestamp 1612251222
transform -1 0 56 0 -1 5410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_567
timestamp 1612251222
transform -1 0 40 0 -1 5410
box -4 -6 20 206
use FILL  FILL_PAND2X1_567
timestamp 1612251222
transform -1 0 24 0 -1 5410
box -4 -6 20 206
use FILL  FILL_26_12
timestamp 1612251222
transform 1 0 10246 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_11
timestamp 1612251222
transform 1 0 10230 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_10
timestamp 1612251222
transform 1 0 10214 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_9
timestamp 1612251222
transform 1 0 10198 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_8
timestamp 1612251222
transform 1 0 10182 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_7
timestamp 1612251222
transform 1 0 10166 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_6
timestamp 1612251222
transform 1 0 10150 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_5
timestamp 1612251222
transform 1 0 10134 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_4
timestamp 1612251222
transform 1 0 10118 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_3
timestamp 1612251222
transform 1 0 10102 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_2
timestamp 1612251222
transform 1 0 10086 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_1
timestamp 1612251222
transform 1 0 10070 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_168
timestamp 1612251222
transform -1 0 10070 0 1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_168
timestamp 1612251222
transform -1 0 9904 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_168
timestamp 1612251222
transform -1 0 9888 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_168
timestamp 1612251222
transform -1 0 9872 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_165
timestamp 1612251222
transform 1 0 9690 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_165
timestamp 1612251222
transform 1 0 9674 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_165
timestamp 1612251222
transform 1 0 9658 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_165
timestamp 1612251222
transform 1 0 9642 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_165
timestamp 1612251222
transform 1 0 9626 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_174
timestamp 1612251222
transform 1 0 9460 0 1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_174
timestamp 1612251222
transform 1 0 9444 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_174
timestamp 1612251222
transform 1 0 9428 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_174
timestamp 1612251222
transform 1 0 9412 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_175
timestamp 1612251222
transform -1 0 9412 0 1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_175
timestamp 1612251222
transform -1 0 9246 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_175
timestamp 1612251222
transform -1 0 9230 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_175
timestamp 1612251222
transform -1 0 9214 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_456
timestamp 1612251222
transform 1 0 9032 0 1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_456
timestamp 1612251222
transform 1 0 9016 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_456
timestamp 1612251222
transform 1 0 9000 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_456
timestamp 1612251222
transform 1 0 8984 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_445
timestamp 1612251222
transform 1 0 8818 0 1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_445
timestamp 1612251222
transform 1 0 8802 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_445
timestamp 1612251222
transform 1 0 8786 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_445
timestamp 1612251222
transform 1 0 8770 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_455
timestamp 1612251222
transform -1 0 8770 0 1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_455
timestamp 1612251222
transform -1 0 8604 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_455
timestamp 1612251222
transform -1 0 8588 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_455
timestamp 1612251222
transform -1 0 8572 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_715
timestamp 1612251222
transform -1 0 8556 0 1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_715
timestamp 1612251222
transform -1 0 8390 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_715
timestamp 1612251222
transform -1 0 8374 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_715
timestamp 1612251222
transform -1 0 8358 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_541
timestamp 1612251222
transform 1 0 8176 0 1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_541
timestamp 1612251222
transform 1 0 8160 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_541
timestamp 1612251222
transform 1 0 8144 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_541
timestamp 1612251222
transform 1 0 8128 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_323
timestamp 1612251222
transform 1 0 7962 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_323
timestamp 1612251222
transform 1 0 7946 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_323
timestamp 1612251222
transform 1 0 7930 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_323
timestamp 1612251222
transform 1 0 7914 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_323
timestamp 1612251222
transform 1 0 7898 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_74
timestamp 1612251222
transform -1 0 7898 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_74
timestamp 1612251222
transform -1 0 7732 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_74
timestamp 1612251222
transform -1 0 7716 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_74
timestamp 1612251222
transform -1 0 7700 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_74
timestamp 1612251222
transform -1 0 7684 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_579
timestamp 1612251222
transform 1 0 7502 0 1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_579
timestamp 1612251222
transform 1 0 7486 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_579
timestamp 1612251222
transform 1 0 7470 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_579
timestamp 1612251222
transform 1 0 7454 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_573
timestamp 1612251222
transform -1 0 7454 0 1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_573
timestamp 1612251222
transform -1 0 7288 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_573
timestamp 1612251222
transform -1 0 7272 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_573
timestamp 1612251222
transform -1 0 7256 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_499
timestamp 1612251222
transform -1 0 7240 0 1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_499
timestamp 1612251222
transform -1 0 7074 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_499
timestamp 1612251222
transform -1 0 7058 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_499
timestamp 1612251222
transform -1 0 7042 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_316
timestamp 1612251222
transform -1 0 7026 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_316
timestamp 1612251222
transform -1 0 6860 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_316
timestamp 1612251222
transform -1 0 6844 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_316
timestamp 1612251222
transform -1 0 6828 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_316
timestamp 1612251222
transform -1 0 6812 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_184
timestamp 1612251222
transform 1 0 6630 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_184
timestamp 1612251222
transform 1 0 6614 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_184
timestamp 1612251222
transform 1 0 6598 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_184
timestamp 1612251222
transform 1 0 6582 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_184
timestamp 1612251222
transform 1 0 6566 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_497
timestamp 1612251222
transform -1 0 6566 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_497
timestamp 1612251222
transform -1 0 6400 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_497
timestamp 1612251222
transform -1 0 6384 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_497
timestamp 1612251222
transform -1 0 6368 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_497
timestamp 1612251222
transform -1 0 6352 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_110
timestamp 1612251222
transform 1 0 6170 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_110
timestamp 1612251222
transform 1 0 6154 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_110
timestamp 1612251222
transform 1 0 6138 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_110
timestamp 1612251222
transform 1 0 6122 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_110
timestamp 1612251222
transform 1 0 6106 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_565
timestamp 1612251222
transform 1 0 5940 0 1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_565
timestamp 1612251222
transform 1 0 5924 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_565
timestamp 1612251222
transform 1 0 5908 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_565
timestamp 1612251222
transform 1 0 5892 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_525
timestamp 1612251222
transform -1 0 5892 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_525
timestamp 1612251222
transform -1 0 5726 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_525
timestamp 1612251222
transform -1 0 5710 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_525
timestamp 1612251222
transform -1 0 5694 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_525
timestamp 1612251222
transform -1 0 5678 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_550
timestamp 1612251222
transform -1 0 5662 0 1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_550
timestamp 1612251222
transform -1 0 5496 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_550
timestamp 1612251222
transform -1 0 5480 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_550
timestamp 1612251222
transform -1 0 5464 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_754
timestamp 1612251222
transform 1 0 5282 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_754
timestamp 1612251222
transform 1 0 5266 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_754
timestamp 1612251222
transform 1 0 5250 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_754
timestamp 1612251222
transform 1 0 5234 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_754
timestamp 1612251222
transform 1 0 5218 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_522
timestamp 1612251222
transform -1 0 5218 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_522
timestamp 1612251222
transform -1 0 5052 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_522
timestamp 1612251222
transform -1 0 5036 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_522
timestamp 1612251222
transform -1 0 5020 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_522
timestamp 1612251222
transform -1 0 5004 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_523
timestamp 1612251222
transform -1 0 4988 0 1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_523
timestamp 1612251222
transform -1 0 4822 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_523
timestamp 1612251222
transform -1 0 4806 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_523
timestamp 1612251222
transform -1 0 4790 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_820
timestamp 1612251222
transform -1 0 4774 0 1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_820
timestamp 1612251222
transform -1 0 4608 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_820
timestamp 1612251222
transform -1 0 4592 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_820
timestamp 1612251222
transform -1 0 4576 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_847
timestamp 1612251222
transform 1 0 4394 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_847
timestamp 1612251222
transform 1 0 4378 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_847
timestamp 1612251222
transform 1 0 4362 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_847
timestamp 1612251222
transform 1 0 4346 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_847
timestamp 1612251222
transform 1 0 4330 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_58
timestamp 1612251222
transform -1 0 4330 0 1 5010
box -4 -6 170 206
use FILL  FILL2_POR2X1_58
timestamp 1612251222
transform -1 0 4164 0 1 5010
box -4 -6 20 206
use FILL  FILL1_POR2X1_58
timestamp 1612251222
transform -1 0 4148 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_58
timestamp 1612251222
transform -1 0 4132 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_58
timestamp 1612251222
transform -1 0 4116 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_61
timestamp 1612251222
transform 1 0 3934 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_61
timestamp 1612251222
transform 1 0 3918 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_61
timestamp 1612251222
transform 1 0 3902 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_61
timestamp 1612251222
transform 1 0 3886 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_61
timestamp 1612251222
transform 1 0 3870 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_849
timestamp 1612251222
transform 1 0 3704 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_849
timestamp 1612251222
transform 1 0 3688 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_849
timestamp 1612251222
transform 1 0 3672 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_849
timestamp 1612251222
transform 1 0 3656 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_849
timestamp 1612251222
transform 1 0 3640 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_338
timestamp 1612251222
transform -1 0 3640 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_338
timestamp 1612251222
transform -1 0 3474 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_338
timestamp 1612251222
transform -1 0 3458 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_338
timestamp 1612251222
transform -1 0 3442 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_338
timestamp 1612251222
transform -1 0 3426 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_844
timestamp 1612251222
transform 1 0 3244 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_844
timestamp 1612251222
transform 1 0 3228 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_844
timestamp 1612251222
transform 1 0 3212 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_844
timestamp 1612251222
transform 1 0 3196 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_844
timestamp 1612251222
transform 1 0 3180 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_521
timestamp 1612251222
transform -1 0 3180 0 1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_521
timestamp 1612251222
transform -1 0 3014 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_521
timestamp 1612251222
transform -1 0 2998 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_521
timestamp 1612251222
transform -1 0 2982 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_523
timestamp 1612251222
transform -1 0 2966 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_523
timestamp 1612251222
transform -1 0 2800 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_523
timestamp 1612251222
transform -1 0 2784 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_523
timestamp 1612251222
transform -1 0 2768 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_523
timestamp 1612251222
transform -1 0 2752 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_560
timestamp 1612251222
transform -1 0 2736 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_560
timestamp 1612251222
transform -1 0 2570 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_560
timestamp 1612251222
transform -1 0 2554 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_560
timestamp 1612251222
transform -1 0 2538 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_560
timestamp 1612251222
transform -1 0 2522 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_476
timestamp 1612251222
transform -1 0 2506 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_476
timestamp 1612251222
transform -1 0 2340 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_476
timestamp 1612251222
transform -1 0 2324 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_476
timestamp 1612251222
transform -1 0 2308 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_476
timestamp 1612251222
transform -1 0 2292 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_576
timestamp 1612251222
transform 1 0 2110 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_576
timestamp 1612251222
transform 1 0 2094 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_576
timestamp 1612251222
transform 1 0 2078 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_576
timestamp 1612251222
transform 1 0 2062 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_576
timestamp 1612251222
transform 1 0 2046 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_571
timestamp 1612251222
transform -1 0 2046 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_571
timestamp 1612251222
transform -1 0 1880 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_571
timestamp 1612251222
transform -1 0 1864 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_571
timestamp 1612251222
transform -1 0 1848 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_571
timestamp 1612251222
transform -1 0 1832 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_557
timestamp 1612251222
transform 1 0 1650 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_557
timestamp 1612251222
transform 1 0 1634 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_557
timestamp 1612251222
transform 1 0 1618 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_557
timestamp 1612251222
transform 1 0 1602 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_557
timestamp 1612251222
transform 1 0 1586 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_653
timestamp 1612251222
transform 1 0 1420 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_653
timestamp 1612251222
transform 1 0 1404 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_653
timestamp 1612251222
transform 1 0 1388 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_653
timestamp 1612251222
transform 1 0 1372 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_653
timestamp 1612251222
transform 1 0 1356 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_652
timestamp 1612251222
transform 1 0 1190 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_652
timestamp 1612251222
transform 1 0 1174 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_652
timestamp 1612251222
transform 1 0 1158 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_652
timestamp 1612251222
transform 1 0 1142 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_652
timestamp 1612251222
transform 1 0 1126 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_250
timestamp 1612251222
transform 1 0 960 0 1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_250
timestamp 1612251222
transform 1 0 944 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_250
timestamp 1612251222
transform 1 0 928 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_250
timestamp 1612251222
transform 1 0 912 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_364
timestamp 1612251222
transform -1 0 912 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_364
timestamp 1612251222
transform -1 0 746 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_364
timestamp 1612251222
transform -1 0 730 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_364
timestamp 1612251222
transform -1 0 714 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_364
timestamp 1612251222
transform -1 0 698 0 1 5010
box -4 -6 20 206
use POR2X1  POR2X1_283
timestamp 1612251222
transform -1 0 682 0 1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_283
timestamp 1612251222
transform -1 0 516 0 1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_283
timestamp 1612251222
transform -1 0 500 0 1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_283
timestamp 1612251222
transform -1 0 484 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_223
timestamp 1612251222
transform -1 0 468 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_223
timestamp 1612251222
transform -1 0 302 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_223
timestamp 1612251222
transform -1 0 286 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_223
timestamp 1612251222
transform -1 0 270 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_223
timestamp 1612251222
transform -1 0 254 0 1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_286
timestamp 1612251222
transform 1 0 72 0 1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_286
timestamp 1612251222
transform 1 0 56 0 1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_286
timestamp 1612251222
transform 1 0 40 0 1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_286
timestamp 1612251222
transform 1 0 24 0 1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_286
timestamp 1612251222
transform 1 0 8 0 1 5010
box -4 -6 20 206
use FILL  FILL_25_5
timestamp 1612251222
transform -1 0 10268 0 -1 5010
box -4 -6 20 206
use FILL  FILL_25_4
timestamp 1612251222
transform -1 0 10252 0 -1 5010
box -4 -6 20 206
use FILL  FILL_25_3
timestamp 1612251222
transform -1 0 10236 0 -1 5010
box -4 -6 20 206
use FILL  FILL_25_2
timestamp 1612251222
transform -1 0 10220 0 -1 5010
box -4 -6 20 206
use FILL  FILL_25_1
timestamp 1612251222
transform -1 0 10204 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_578
timestamp 1612251222
transform 1 0 10022 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_578
timestamp 1612251222
transform 1 0 10006 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_578
timestamp 1612251222
transform 1 0 9990 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_578
timestamp 1612251222
transform 1 0 9974 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_577
timestamp 1612251222
transform 1 0 9808 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_577
timestamp 1612251222
transform 1 0 9792 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_577
timestamp 1612251222
transform 1 0 9776 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_577
timestamp 1612251222
transform 1 0 9760 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_569
timestamp 1612251222
transform 1 0 9594 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_569
timestamp 1612251222
transform 1 0 9578 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_569
timestamp 1612251222
transform 1 0 9562 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_569
timestamp 1612251222
transform 1 0 9546 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_570
timestamp 1612251222
transform 1 0 9380 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_570
timestamp 1612251222
transform 1 0 9364 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_570
timestamp 1612251222
transform 1 0 9348 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_570
timestamp 1612251222
transform 1 0 9332 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_465
timestamp 1612251222
transform 1 0 9166 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_465
timestamp 1612251222
transform 1 0 9150 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_465
timestamp 1612251222
transform 1 0 9134 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_465
timestamp 1612251222
transform 1 0 9118 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_563
timestamp 1612251222
transform 1 0 8952 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_563
timestamp 1612251222
transform 1 0 8936 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_563
timestamp 1612251222
transform 1 0 8920 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_563
timestamp 1612251222
transform 1 0 8904 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_553
timestamp 1612251222
transform 1 0 8738 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_553
timestamp 1612251222
transform 1 0 8722 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_553
timestamp 1612251222
transform 1 0 8706 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_553
timestamp 1612251222
transform 1 0 8690 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_272
timestamp 1612251222
transform -1 0 8690 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_272
timestamp 1612251222
transform -1 0 8524 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_272
timestamp 1612251222
transform -1 0 8508 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_272
timestamp 1612251222
transform -1 0 8492 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_272
timestamp 1612251222
transform -1 0 8476 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_76
timestamp 1612251222
transform 1 0 8294 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_76
timestamp 1612251222
transform 1 0 8278 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_76
timestamp 1612251222
transform 1 0 8262 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_76
timestamp 1612251222
transform 1 0 8246 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_274
timestamp 1612251222
transform -1 0 8246 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_274
timestamp 1612251222
transform -1 0 8080 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_274
timestamp 1612251222
transform -1 0 8064 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_274
timestamp 1612251222
transform -1 0 8048 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_275
timestamp 1612251222
transform 1 0 7866 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_275
timestamp 1612251222
transform 1 0 7850 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_275
timestamp 1612251222
transform 1 0 7834 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_275
timestamp 1612251222
transform 1 0 7818 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_275
timestamp 1612251222
transform 1 0 7802 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_575
timestamp 1612251222
transform -1 0 7802 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_575
timestamp 1612251222
transform -1 0 7636 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_575
timestamp 1612251222
transform -1 0 7620 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_575
timestamp 1612251222
transform -1 0 7604 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_501
timestamp 1612251222
transform 1 0 7422 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_501
timestamp 1612251222
transform 1 0 7406 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_501
timestamp 1612251222
transform 1 0 7390 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_501
timestamp 1612251222
transform 1 0 7374 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_496
timestamp 1612251222
transform 1 0 7208 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_496
timestamp 1612251222
transform 1 0 7192 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_496
timestamp 1612251222
transform 1 0 7176 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_496
timestamp 1612251222
transform 1 0 7160 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_496
timestamp 1612251222
transform 1 0 7144 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_576
timestamp 1612251222
transform 1 0 6978 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_576
timestamp 1612251222
transform 1 0 6962 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_576
timestamp 1612251222
transform 1 0 6946 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_576
timestamp 1612251222
transform 1 0 6930 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_500
timestamp 1612251222
transform 1 0 6764 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_500
timestamp 1612251222
transform 1 0 6748 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_500
timestamp 1612251222
transform 1 0 6732 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_500
timestamp 1612251222
transform 1 0 6716 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_78
timestamp 1612251222
transform -1 0 6716 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_78
timestamp 1612251222
transform -1 0 6550 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_78
timestamp 1612251222
transform -1 0 6534 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_78
timestamp 1612251222
transform -1 0 6518 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_79
timestamp 1612251222
transform 1 0 6336 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_79
timestamp 1612251222
transform 1 0 6320 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_79
timestamp 1612251222
transform 1 0 6304 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_79
timestamp 1612251222
transform 1 0 6288 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_79
timestamp 1612251222
transform 1 0 6272 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_571
timestamp 1612251222
transform 1 0 6106 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_571
timestamp 1612251222
transform 1 0 6090 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_571
timestamp 1612251222
transform 1 0 6074 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_571
timestamp 1612251222
transform 1 0 6058 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_560
timestamp 1612251222
transform 1 0 5892 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_560
timestamp 1612251222
transform 1 0 5876 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_560
timestamp 1612251222
transform 1 0 5860 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_560
timestamp 1612251222
transform 1 0 5844 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_546
timestamp 1612251222
transform 1 0 5678 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_546
timestamp 1612251222
transform 1 0 5662 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_546
timestamp 1612251222
transform 1 0 5646 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_546
timestamp 1612251222
transform 1 0 5630 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_844
timestamp 1612251222
transform -1 0 5630 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_844
timestamp 1612251222
transform -1 0 5464 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_844
timestamp 1612251222
transform -1 0 5448 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_844
timestamp 1612251222
transform -1 0 5432 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_849
timestamp 1612251222
transform -1 0 5416 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_849
timestamp 1612251222
transform -1 0 5250 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_849
timestamp 1612251222
transform -1 0 5234 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_849
timestamp 1612251222
transform -1 0 5218 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_521
timestamp 1612251222
transform -1 0 5202 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_521
timestamp 1612251222
transform -1 0 5036 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_521
timestamp 1612251222
transform -1 0 5020 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_521
timestamp 1612251222
transform -1 0 5004 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_521
timestamp 1612251222
transform -1 0 4988 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_819
timestamp 1612251222
transform -1 0 4972 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_819
timestamp 1612251222
transform -1 0 4806 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_819
timestamp 1612251222
transform -1 0 4790 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_819
timestamp 1612251222
transform -1 0 4774 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_818
timestamp 1612251222
transform 1 0 4592 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_818
timestamp 1612251222
transform 1 0 4576 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_818
timestamp 1612251222
transform 1 0 4560 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_818
timestamp 1612251222
transform 1 0 4544 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_818
timestamp 1612251222
transform 1 0 4528 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_817
timestamp 1612251222
transform -1 0 4528 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_817
timestamp 1612251222
transform -1 0 4362 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_817
timestamp 1612251222
transform -1 0 4346 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_817
timestamp 1612251222
transform -1 0 4330 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_381
timestamp 1612251222
transform 1 0 4148 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_381
timestamp 1612251222
transform 1 0 4132 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_381
timestamp 1612251222
transform 1 0 4116 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_381
timestamp 1612251222
transform 1 0 4100 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_9
timestamp 1612251222
transform -1 0 4100 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_POR2X1_9
timestamp 1612251222
transform -1 0 3934 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_POR2X1_9
timestamp 1612251222
transform -1 0 3918 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_9
timestamp 1612251222
transform -1 0 3902 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_9
timestamp 1612251222
transform -1 0 3886 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_98
timestamp 1612251222
transform -1 0 3870 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_98
timestamp 1612251222
transform -1 0 3704 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_98
timestamp 1612251222
transform -1 0 3688 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_98
timestamp 1612251222
transform -1 0 3672 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_98
timestamp 1612251222
transform -1 0 3656 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_99
timestamp 1612251222
transform 1 0 3474 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_99
timestamp 1612251222
transform 1 0 3458 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_99
timestamp 1612251222
transform 1 0 3442 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_99
timestamp 1612251222
transform 1 0 3426 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_99
timestamp 1612251222
transform 1 0 3410 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_351
timestamp 1612251222
transform 1 0 3244 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_351
timestamp 1612251222
transform 1 0 3228 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_351
timestamp 1612251222
transform 1 0 3212 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_351
timestamp 1612251222
transform 1 0 3196 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_351
timestamp 1612251222
transform 1 0 3180 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_60
timestamp 1612251222
transform 1 0 3014 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_POR2X1_60
timestamp 1612251222
transform 1 0 2998 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_POR2X1_60
timestamp 1612251222
transform 1 0 2982 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_60
timestamp 1612251222
transform 1 0 2966 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_60
timestamp 1612251222
transform 1 0 2950 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_522
timestamp 1612251222
transform 1 0 2784 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_522
timestamp 1612251222
transform 1 0 2768 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_522
timestamp 1612251222
transform 1 0 2752 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_522
timestamp 1612251222
transform 1 0 2736 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_339
timestamp 1612251222
transform 1 0 2570 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_339
timestamp 1612251222
transform 1 0 2554 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_339
timestamp 1612251222
transform 1 0 2538 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_339
timestamp 1612251222
transform 1 0 2522 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_339
timestamp 1612251222
transform 1 0 2506 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_475
timestamp 1612251222
transform -1 0 2506 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_475
timestamp 1612251222
transform -1 0 2340 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_475
timestamp 1612251222
transform -1 0 2324 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_475
timestamp 1612251222
transform -1 0 2308 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_475
timestamp 1612251222
transform -1 0 2292 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_479
timestamp 1612251222
transform -1 0 2276 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_479
timestamp 1612251222
transform -1 0 2110 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_479
timestamp 1612251222
transform -1 0 2094 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_479
timestamp 1612251222
transform -1 0 2078 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_479
timestamp 1612251222
transform -1 0 2062 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_561
timestamp 1612251222
transform 1 0 1880 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_561
timestamp 1612251222
transform 1 0 1864 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_561
timestamp 1612251222
transform 1 0 1848 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_561
timestamp 1612251222
transform 1 0 1832 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_561
timestamp 1612251222
transform 1 0 1816 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_473
timestamp 1612251222
transform 1 0 1650 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_473
timestamp 1612251222
transform 1 0 1634 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_473
timestamp 1612251222
transform 1 0 1618 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_473
timestamp 1612251222
transform 1 0 1602 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_473
timestamp 1612251222
transform 1 0 1586 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_361
timestamp 1612251222
transform -1 0 1586 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_361
timestamp 1612251222
transform -1 0 1420 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_361
timestamp 1612251222
transform -1 0 1404 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_361
timestamp 1612251222
transform -1 0 1388 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_361
timestamp 1612251222
transform -1 0 1372 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_594
timestamp 1612251222
transform 1 0 1190 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_594
timestamp 1612251222
transform 1 0 1174 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_594
timestamp 1612251222
transform 1 0 1158 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_594
timestamp 1612251222
transform 1 0 1142 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_329
timestamp 1612251222
transform -1 0 1142 0 -1 5010
box -4 -6 170 206
use FILL  FILL1_POR2X1_329
timestamp 1612251222
transform -1 0 976 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_POR2X1_329
timestamp 1612251222
transform -1 0 960 0 -1 5010
box -4 -6 20 206
use FILL  FILL_POR2X1_329
timestamp 1612251222
transform -1 0 944 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_355
timestamp 1612251222
transform -1 0 928 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_355
timestamp 1612251222
transform -1 0 762 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_355
timestamp 1612251222
transform -1 0 746 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_355
timestamp 1612251222
transform -1 0 730 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_355
timestamp 1612251222
transform -1 0 714 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_356
timestamp 1612251222
transform -1 0 698 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_356
timestamp 1612251222
transform -1 0 532 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_356
timestamp 1612251222
transform -1 0 516 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_356
timestamp 1612251222
transform -1 0 500 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_356
timestamp 1612251222
transform -1 0 484 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_365
timestamp 1612251222
transform -1 0 468 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_365
timestamp 1612251222
transform -1 0 302 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_365
timestamp 1612251222
transform -1 0 286 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_365
timestamp 1612251222
transform -1 0 270 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_365
timestamp 1612251222
transform -1 0 254 0 -1 5010
box -4 -6 20 206
use PAND2X1  PAND2X1_367
timestamp 1612251222
transform -1 0 238 0 -1 5010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_367
timestamp 1612251222
transform -1 0 72 0 -1 5010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_367
timestamp 1612251222
transform -1 0 56 0 -1 5010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_367
timestamp 1612251222
transform -1 0 40 0 -1 5010
box -4 -6 20 206
use FILL  FILL_PAND2X1_367
timestamp 1612251222
transform -1 0 24 0 -1 5010
box -4 -6 20 206
use POR2X1  POR2X1_170
timestamp 1612251222
transform 1 0 10102 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_170
timestamp 1612251222
transform 1 0 10086 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_170
timestamp 1612251222
transform 1 0 10070 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_170
timestamp 1612251222
transform 1 0 10054 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_169
timestamp 1612251222
transform 1 0 9888 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_169
timestamp 1612251222
transform 1 0 9872 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_169
timestamp 1612251222
transform 1 0 9856 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_169
timestamp 1612251222
transform 1 0 9840 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_166
timestamp 1612251222
transform 1 0 9674 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_166
timestamp 1612251222
transform 1 0 9658 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_166
timestamp 1612251222
transform 1 0 9642 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_166
timestamp 1612251222
transform 1 0 9626 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_166
timestamp 1612251222
transform 1 0 9610 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_315
timestamp 1612251222
transform -1 0 9610 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_315
timestamp 1612251222
transform -1 0 9444 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_315
timestamp 1612251222
transform -1 0 9428 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_315
timestamp 1612251222
transform -1 0 9412 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_315
timestamp 1612251222
transform -1 0 9396 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_318
timestamp 1612251222
transform 1 0 9214 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_318
timestamp 1612251222
transform 1 0 9198 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_318
timestamp 1612251222
transform 1 0 9182 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_318
timestamp 1612251222
transform 1 0 9166 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_127
timestamp 1612251222
transform -1 0 9166 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_127
timestamp 1612251222
transform -1 0 9000 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_127
timestamp 1612251222
transform -1 0 8984 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_127
timestamp 1612251222
transform -1 0 8968 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_127
timestamp 1612251222
transform -1 0 8952 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_735
timestamp 1612251222
transform 1 0 8770 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_735
timestamp 1612251222
transform 1 0 8754 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_735
timestamp 1612251222
transform 1 0 8738 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_735
timestamp 1612251222
transform 1 0 8722 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_658
timestamp 1612251222
transform 1 0 8556 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_658
timestamp 1612251222
transform 1 0 8540 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_658
timestamp 1612251222
transform 1 0 8524 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_658
timestamp 1612251222
transform 1 0 8508 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_75
timestamp 1612251222
transform -1 0 8508 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_75
timestamp 1612251222
transform -1 0 8342 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_75
timestamp 1612251222
transform -1 0 8326 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_75
timestamp 1612251222
transform -1 0 8310 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_75
timestamp 1612251222
transform -1 0 8294 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_131
timestamp 1612251222
transform -1 0 8278 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_131
timestamp 1612251222
transform -1 0 8112 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_131
timestamp 1612251222
transform -1 0 8096 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_131
timestamp 1612251222
transform -1 0 8080 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_131
timestamp 1612251222
transform -1 0 8064 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_140
timestamp 1612251222
transform -1 0 8048 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_140
timestamp 1612251222
transform -1 0 7882 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_140
timestamp 1612251222
transform -1 0 7866 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_140
timestamp 1612251222
transform -1 0 7850 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_130
timestamp 1612251222
transform 1 0 7668 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_130
timestamp 1612251222
transform 1 0 7652 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_130
timestamp 1612251222
transform 1 0 7636 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_130
timestamp 1612251222
transform 1 0 7620 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_138
timestamp 1612251222
transform -1 0 7620 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_138
timestamp 1612251222
transform -1 0 7454 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_138
timestamp 1612251222
transform -1 0 7438 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_138
timestamp 1612251222
transform -1 0 7422 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_136
timestamp 1612251222
transform 1 0 7240 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_136
timestamp 1612251222
transform 1 0 7224 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_136
timestamp 1612251222
transform 1 0 7208 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_136
timestamp 1612251222
transform 1 0 7192 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_136
timestamp 1612251222
transform 1 0 7176 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_267
timestamp 1612251222
transform 1 0 7010 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_267
timestamp 1612251222
transform 1 0 6994 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_267
timestamp 1612251222
transform 1 0 6978 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_267
timestamp 1612251222
transform 1 0 6962 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_641
timestamp 1612251222
transform -1 0 6962 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_641
timestamp 1612251222
transform -1 0 6796 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_641
timestamp 1612251222
transform -1 0 6780 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_641
timestamp 1612251222
transform -1 0 6764 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_767
timestamp 1612251222
transform 1 0 6582 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_767
timestamp 1612251222
transform 1 0 6566 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_767
timestamp 1612251222
transform 1 0 6550 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_767
timestamp 1612251222
transform 1 0 6534 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_767
timestamp 1612251222
transform 1 0 6518 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_557
timestamp 1612251222
transform -1 0 6518 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_557
timestamp 1612251222
transform -1 0 6352 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_557
timestamp 1612251222
transform -1 0 6336 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_557
timestamp 1612251222
transform -1 0 6320 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_561
timestamp 1612251222
transform -1 0 6304 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_561
timestamp 1612251222
transform -1 0 6138 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_561
timestamp 1612251222
transform -1 0 6122 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_561
timestamp 1612251222
transform -1 0 6106 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_129
timestamp 1612251222
transform 1 0 5924 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_129
timestamp 1612251222
transform 1 0 5908 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_129
timestamp 1612251222
transform 1 0 5892 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_129
timestamp 1612251222
transform 1 0 5876 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_129
timestamp 1612251222
transform 1 0 5860 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_559
timestamp 1612251222
transform 1 0 5694 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_559
timestamp 1612251222
transform 1 0 5678 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_559
timestamp 1612251222
transform 1 0 5662 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_559
timestamp 1612251222
transform 1 0 5646 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_90
timestamp 1612251222
transform 1 0 5480 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_90
timestamp 1612251222
transform 1 0 5464 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_90
timestamp 1612251222
transform 1 0 5448 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_90
timestamp 1612251222
transform 1 0 5432 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_90
timestamp 1612251222
transform 1 0 5416 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_225
timestamp 1612251222
transform 1 0 5250 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_225
timestamp 1612251222
transform 1 0 5234 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_225
timestamp 1612251222
transform 1 0 5218 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_225
timestamp 1612251222
transform 1 0 5202 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_225
timestamp 1612251222
transform 1 0 5186 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_846
timestamp 1612251222
transform -1 0 5186 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_846
timestamp 1612251222
transform -1 0 5020 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_846
timestamp 1612251222
transform -1 0 5004 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_846
timestamp 1612251222
transform -1 0 4988 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_846
timestamp 1612251222
transform -1 0 4972 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_848
timestamp 1612251222
transform -1 0 4956 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_848
timestamp 1612251222
transform -1 0 4790 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_848
timestamp 1612251222
transform -1 0 4774 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_848
timestamp 1612251222
transform -1 0 4758 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_848
timestamp 1612251222
transform -1 0 4742 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_382
timestamp 1612251222
transform 1 0 4560 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_382
timestamp 1612251222
transform 1 0 4544 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_382
timestamp 1612251222
transform 1 0 4528 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_382
timestamp 1612251222
transform 1 0 4512 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_224
timestamp 1612251222
transform -1 0 4512 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_224
timestamp 1612251222
transform -1 0 4346 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_224
timestamp 1612251222
transform -1 0 4330 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_224
timestamp 1612251222
transform -1 0 4314 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_227
timestamp 1612251222
transform -1 0 4298 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_227
timestamp 1612251222
transform -1 0 4132 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_227
timestamp 1612251222
transform -1 0 4116 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_227
timestamp 1612251222
transform -1 0 4100 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_227
timestamp 1612251222
transform -1 0 4084 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_509
timestamp 1612251222
transform -1 0 4068 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_509
timestamp 1612251222
transform -1 0 3902 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_509
timestamp 1612251222
transform -1 0 3886 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_509
timestamp 1612251222
transform -1 0 3870 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_509
timestamp 1612251222
transform -1 0 3854 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_289
timestamp 1612251222
transform -1 0 3838 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_289
timestamp 1612251222
transform -1 0 3672 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_289
timestamp 1612251222
transform -1 0 3656 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_289
timestamp 1612251222
transform -1 0 3640 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_89
timestamp 1612251222
transform -1 0 3624 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_89
timestamp 1612251222
transform -1 0 3458 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_89
timestamp 1612251222
transform -1 0 3442 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_89
timestamp 1612251222
transform -1 0 3426 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_97
timestamp 1612251222
transform -1 0 3410 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_97
timestamp 1612251222
transform -1 0 3244 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_97
timestamp 1612251222
transform -1 0 3228 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_97
timestamp 1612251222
transform -1 0 3212 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_97
timestamp 1612251222
transform -1 0 3196 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_84
timestamp 1612251222
transform -1 0 3180 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_84
timestamp 1612251222
transform -1 0 3014 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_84
timestamp 1612251222
transform -1 0 2998 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_84
timestamp 1612251222
transform -1 0 2982 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_84
timestamp 1612251222
transform -1 0 2966 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_71
timestamp 1612251222
transform 1 0 2784 0 1 4610
box -4 -6 170 206
use FILL  FILL2_POR2X1_71
timestamp 1612251222
transform 1 0 2768 0 1 4610
box -4 -6 20 206
use FILL  FILL1_POR2X1_71
timestamp 1612251222
transform 1 0 2752 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_71
timestamp 1612251222
transform 1 0 2736 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_71
timestamp 1612251222
transform 1 0 2720 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_786
timestamp 1612251222
transform -1 0 2720 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_786
timestamp 1612251222
transform -1 0 2554 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_786
timestamp 1612251222
transform -1 0 2538 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_786
timestamp 1612251222
transform -1 0 2522 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_786
timestamp 1612251222
transform -1 0 2506 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_598
timestamp 1612251222
transform -1 0 2490 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_598
timestamp 1612251222
transform -1 0 2324 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_598
timestamp 1612251222
transform -1 0 2308 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_598
timestamp 1612251222
transform -1 0 2292 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_598
timestamp 1612251222
transform -1 0 2276 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_493
timestamp 1612251222
transform 1 0 2094 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_493
timestamp 1612251222
transform 1 0 2078 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_493
timestamp 1612251222
transform 1 0 2062 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_493
timestamp 1612251222
transform 1 0 2046 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_493
timestamp 1612251222
transform 1 0 2030 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_492
timestamp 1612251222
transform 1 0 1864 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_492
timestamp 1612251222
transform 1 0 1848 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_492
timestamp 1612251222
transform 1 0 1832 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_492
timestamp 1612251222
transform 1 0 1816 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_741
timestamp 1612251222
transform -1 0 1816 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_741
timestamp 1612251222
transform -1 0 1650 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_741
timestamp 1612251222
transform -1 0 1634 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_741
timestamp 1612251222
transform -1 0 1618 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_741
timestamp 1612251222
transform -1 0 1602 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_674
timestamp 1612251222
transform -1 0 1586 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_674
timestamp 1612251222
transform -1 0 1420 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_674
timestamp 1612251222
transform -1 0 1404 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_674
timestamp 1612251222
transform -1 0 1388 0 1 4610
box -4 -6 20 206
use POR2X1  POR2X1_331
timestamp 1612251222
transform -1 0 1372 0 1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_331
timestamp 1612251222
transform -1 0 1206 0 1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_331
timestamp 1612251222
transform -1 0 1190 0 1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_331
timestamp 1612251222
transform -1 0 1174 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_742
timestamp 1612251222
transform -1 0 1158 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_742
timestamp 1612251222
transform -1 0 992 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_742
timestamp 1612251222
transform -1 0 976 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_742
timestamp 1612251222
transform -1 0 960 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_742
timestamp 1612251222
transform -1 0 944 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_362
timestamp 1612251222
transform -1 0 928 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_362
timestamp 1612251222
transform -1 0 762 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_362
timestamp 1612251222
transform -1 0 746 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_362
timestamp 1612251222
transform -1 0 730 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_362
timestamp 1612251222
transform -1 0 714 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_366
timestamp 1612251222
transform -1 0 698 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_366
timestamp 1612251222
transform -1 0 532 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_366
timestamp 1612251222
transform -1 0 516 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_366
timestamp 1612251222
transform -1 0 500 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_366
timestamp 1612251222
transform -1 0 484 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_810
timestamp 1612251222
transform -1 0 468 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_810
timestamp 1612251222
transform -1 0 302 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_810
timestamp 1612251222
transform -1 0 286 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_810
timestamp 1612251222
transform -1 0 270 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_810
timestamp 1612251222
transform -1 0 254 0 1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_864
timestamp 1612251222
transform 1 0 72 0 1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_864
timestamp 1612251222
transform 1 0 56 0 1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_864
timestamp 1612251222
transform 1 0 40 0 1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_864
timestamp 1612251222
transform 1 0 24 0 1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_864
timestamp 1612251222
transform 1 0 8 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_1
timestamp 1612251222
transform -1 0 10268 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_211
timestamp 1612251222
transform -1 0 10252 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_211
timestamp 1612251222
transform -1 0 10086 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_211
timestamp 1612251222
transform -1 0 10070 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_211
timestamp 1612251222
transform -1 0 10054 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_91
timestamp 1612251222
transform 1 0 9872 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_91
timestamp 1612251222
transform 1 0 9856 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_91
timestamp 1612251222
transform 1 0 9840 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_91
timestamp 1612251222
transform 1 0 9824 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_91
timestamp 1612251222
transform 1 0 9808 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_418
timestamp 1612251222
transform -1 0 9808 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_418
timestamp 1612251222
transform -1 0 9642 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_418
timestamp 1612251222
transform -1 0 9626 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_418
timestamp 1612251222
transform -1 0 9610 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_418
timestamp 1612251222
transform -1 0 9594 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_446
timestamp 1612251222
transform -1 0 9578 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_446
timestamp 1612251222
transform -1 0 9412 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_446
timestamp 1612251222
transform -1 0 9396 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_446
timestamp 1612251222
transform -1 0 9380 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_454
timestamp 1612251222
transform 1 0 9198 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_454
timestamp 1612251222
transform 1 0 9182 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_454
timestamp 1612251222
transform 1 0 9166 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_454
timestamp 1612251222
transform 1 0 9150 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_125
timestamp 1612251222
transform -1 0 9150 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_125
timestamp 1612251222
transform -1 0 8984 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_125
timestamp 1612251222
transform -1 0 8968 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_125
timestamp 1612251222
transform -1 0 8952 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_125
timestamp 1612251222
transform -1 0 8936 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_128
timestamp 1612251222
transform -1 0 8920 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_128
timestamp 1612251222
transform -1 0 8754 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_128
timestamp 1612251222
transform -1 0 8738 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_128
timestamp 1612251222
transform -1 0 8722 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_554
timestamp 1612251222
transform 1 0 8540 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_554
timestamp 1612251222
transform 1 0 8524 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_554
timestamp 1612251222
transform 1 0 8508 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_554
timestamp 1612251222
transform 1 0 8492 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_574
timestamp 1612251222
transform -1 0 8492 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_574
timestamp 1612251222
transform -1 0 8326 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_574
timestamp 1612251222
transform -1 0 8310 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_574
timestamp 1612251222
transform -1 0 8294 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_516
timestamp 1612251222
transform 1 0 8112 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_516
timestamp 1612251222
transform 1 0 8096 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_516
timestamp 1612251222
transform 1 0 8080 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_516
timestamp 1612251222
transform 1 0 8064 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_516
timestamp 1612251222
transform 1 0 8048 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_515
timestamp 1612251222
transform 1 0 7882 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_515
timestamp 1612251222
transform 1 0 7866 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_515
timestamp 1612251222
transform 1 0 7850 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_515
timestamp 1612251222
transform 1 0 7834 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_141
timestamp 1612251222
transform 1 0 7668 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_141
timestamp 1612251222
transform 1 0 7652 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_141
timestamp 1612251222
transform 1 0 7636 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_141
timestamp 1612251222
transform 1 0 7620 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_139
timestamp 1612251222
transform 1 0 7454 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_139
timestamp 1612251222
transform 1 0 7438 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_139
timestamp 1612251222
transform 1 0 7422 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_139
timestamp 1612251222
transform 1 0 7406 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_514
timestamp 1612251222
transform 1 0 7240 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_514
timestamp 1612251222
transform 1 0 7224 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_514
timestamp 1612251222
transform 1 0 7208 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_514
timestamp 1612251222
transform 1 0 7192 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_572
timestamp 1612251222
transform -1 0 7192 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_572
timestamp 1612251222
transform -1 0 7026 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_572
timestamp 1612251222
transform -1 0 7010 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_572
timestamp 1612251222
transform -1 0 6994 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_265
timestamp 1612251222
transform 1 0 6812 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_265
timestamp 1612251222
transform 1 0 6796 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_265
timestamp 1612251222
transform 1 0 6780 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_265
timestamp 1612251222
transform 1 0 6764 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_265
timestamp 1612251222
transform 1 0 6748 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_491
timestamp 1612251222
transform 1 0 6582 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_491
timestamp 1612251222
transform 1 0 6566 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_491
timestamp 1612251222
transform 1 0 6550 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_491
timestamp 1612251222
transform 1 0 6534 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_491
timestamp 1612251222
transform 1 0 6518 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_558
timestamp 1612251222
transform -1 0 6518 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_558
timestamp 1612251222
transform -1 0 6352 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_558
timestamp 1612251222
transform -1 0 6336 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_558
timestamp 1612251222
transform -1 0 6320 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_494
timestamp 1612251222
transform 1 0 6138 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_494
timestamp 1612251222
transform 1 0 6122 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_494
timestamp 1612251222
transform 1 0 6106 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_494
timestamp 1612251222
transform 1 0 6090 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_494
timestamp 1612251222
transform 1 0 6074 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_264
timestamp 1612251222
transform 1 0 5908 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_264
timestamp 1612251222
transform 1 0 5892 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_264
timestamp 1612251222
transform 1 0 5876 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_264
timestamp 1612251222
transform 1 0 5860 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_517
timestamp 1612251222
transform -1 0 5860 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_517
timestamp 1612251222
transform -1 0 5694 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_517
timestamp 1612251222
transform -1 0 5678 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_517
timestamp 1612251222
transform -1 0 5662 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_517
timestamp 1612251222
transform -1 0 5646 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_667
timestamp 1612251222
transform -1 0 5630 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_667
timestamp 1612251222
transform -1 0 5464 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_667
timestamp 1612251222
transform -1 0 5448 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_667
timestamp 1612251222
transform -1 0 5432 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_667
timestamp 1612251222
transform -1 0 5416 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_816
timestamp 1612251222
transform -1 0 5400 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_816
timestamp 1612251222
transform -1 0 5234 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_816
timestamp 1612251222
transform -1 0 5218 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_816
timestamp 1612251222
transform -1 0 5202 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_815
timestamp 1612251222
transform 1 0 5020 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_815
timestamp 1612251222
transform 1 0 5004 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_815
timestamp 1612251222
transform 1 0 4988 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_815
timestamp 1612251222
transform 1 0 4972 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_814
timestamp 1612251222
transform 1 0 4806 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_814
timestamp 1612251222
transform 1 0 4790 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_814
timestamp 1612251222
transform 1 0 4774 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_814
timestamp 1612251222
transform 1 0 4758 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_814
timestamp 1612251222
transform 1 0 4742 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_226
timestamp 1612251222
transform -1 0 4742 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_226
timestamp 1612251222
transform -1 0 4576 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_226
timestamp 1612251222
transform -1 0 4560 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_226
timestamp 1612251222
transform -1 0 4544 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_502
timestamp 1612251222
transform -1 0 4528 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_502
timestamp 1612251222
transform -1 0 4362 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_502
timestamp 1612251222
transform -1 0 4346 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_502
timestamp 1612251222
transform -1 0 4330 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_502
timestamp 1612251222
transform -1 0 4314 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_503
timestamp 1612251222
transform -1 0 4298 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_503
timestamp 1612251222
transform -1 0 4132 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_503
timestamp 1612251222
transform -1 0 4116 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_503
timestamp 1612251222
transform -1 0 4100 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_93
timestamp 1612251222
transform -1 0 4084 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_93
timestamp 1612251222
transform -1 0 3918 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_93
timestamp 1612251222
transform -1 0 3902 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_93
timestamp 1612251222
transform -1 0 3886 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_859
timestamp 1612251222
transform -1 0 3870 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_859
timestamp 1612251222
transform -1 0 3704 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_859
timestamp 1612251222
transform -1 0 3688 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_859
timestamp 1612251222
transform -1 0 3672 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_859
timestamp 1612251222
transform -1 0 3656 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_333
timestamp 1612251222
transform -1 0 3640 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_333
timestamp 1612251222
transform -1 0 3474 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_333
timestamp 1612251222
transform -1 0 3458 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_333
timestamp 1612251222
transform -1 0 3442 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_333
timestamp 1612251222
transform -1 0 3426 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_474
timestamp 1612251222
transform -1 0 3410 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_474
timestamp 1612251222
transform -1 0 3244 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_474
timestamp 1612251222
transform -1 0 3228 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_474
timestamp 1612251222
transform -1 0 3212 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_474
timestamp 1612251222
transform -1 0 3196 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_500
timestamp 1612251222
transform -1 0 3180 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_500
timestamp 1612251222
transform -1 0 3014 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_500
timestamp 1612251222
transform -1 0 2998 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_500
timestamp 1612251222
transform -1 0 2982 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_500
timestamp 1612251222
transform -1 0 2966 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_497
timestamp 1612251222
transform 1 0 2784 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_497
timestamp 1612251222
transform 1 0 2768 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_497
timestamp 1612251222
transform 1 0 2752 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_497
timestamp 1612251222
transform 1 0 2736 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_150
timestamp 1612251222
transform -1 0 2736 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_150
timestamp 1612251222
transform -1 0 2570 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_150
timestamp 1612251222
transform -1 0 2554 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_150
timestamp 1612251222
transform -1 0 2538 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_558
timestamp 1612251222
transform -1 0 2522 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_558
timestamp 1612251222
transform -1 0 2356 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_558
timestamp 1612251222
transform -1 0 2340 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_558
timestamp 1612251222
transform -1 0 2324 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_558
timestamp 1612251222
transform -1 0 2308 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_717
timestamp 1612251222
transform -1 0 2292 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_717
timestamp 1612251222
transform -1 0 2126 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_717
timestamp 1612251222
transform -1 0 2110 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_717
timestamp 1612251222
transform -1 0 2094 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_717
timestamp 1612251222
transform -1 0 2078 0 -1 4610
box -4 -6 20 206
use POR2X1  POR2X1_491
timestamp 1612251222
transform 1 0 1896 0 -1 4610
box -4 -6 170 206
use FILL  FILL1_POR2X1_491
timestamp 1612251222
transform 1 0 1880 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_POR2X1_491
timestamp 1612251222
transform 1 0 1864 0 -1 4610
box -4 -6 20 206
use FILL  FILL_POR2X1_491
timestamp 1612251222
transform 1 0 1848 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_736
timestamp 1612251222
transform 1 0 1682 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_736
timestamp 1612251222
transform 1 0 1666 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_736
timestamp 1612251222
transform 1 0 1650 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_736
timestamp 1612251222
transform 1 0 1634 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_736
timestamp 1612251222
transform 1 0 1618 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_186
timestamp 1612251222
transform -1 0 1618 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_186
timestamp 1612251222
transform -1 0 1452 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_186
timestamp 1612251222
transform -1 0 1436 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_186
timestamp 1612251222
transform -1 0 1420 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_186
timestamp 1612251222
transform -1 0 1404 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_330
timestamp 1612251222
transform 1 0 1222 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_330
timestamp 1612251222
transform 1 0 1206 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_330
timestamp 1612251222
transform 1 0 1190 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_330
timestamp 1612251222
transform 1 0 1174 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_330
timestamp 1612251222
transform 1 0 1158 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_675
timestamp 1612251222
transform -1 0 1158 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_675
timestamp 1612251222
transform -1 0 992 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_675
timestamp 1612251222
transform -1 0 976 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_675
timestamp 1612251222
transform -1 0 960 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_675
timestamp 1612251222
transform -1 0 944 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_806
timestamp 1612251222
transform -1 0 928 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_806
timestamp 1612251222
transform -1 0 762 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_806
timestamp 1612251222
transform -1 0 746 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_806
timestamp 1612251222
transform -1 0 730 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_806
timestamp 1612251222
transform -1 0 714 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_354
timestamp 1612251222
transform 1 0 532 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_354
timestamp 1612251222
transform 1 0 516 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_354
timestamp 1612251222
transform 1 0 500 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_354
timestamp 1612251222
transform 1 0 484 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_354
timestamp 1612251222
transform 1 0 468 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_288
timestamp 1612251222
transform 1 0 302 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_288
timestamp 1612251222
transform 1 0 286 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_288
timestamp 1612251222
transform 1 0 270 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_288
timestamp 1612251222
transform 1 0 254 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_288
timestamp 1612251222
transform 1 0 238 0 -1 4610
box -4 -6 20 206
use PAND2X1  PAND2X1_866
timestamp 1612251222
transform -1 0 238 0 -1 4610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_866
timestamp 1612251222
transform -1 0 72 0 -1 4610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_866
timestamp 1612251222
transform -1 0 56 0 -1 4610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_866
timestamp 1612251222
transform -1 0 40 0 -1 4610
box -4 -6 20 206
use FILL  FILL_PAND2X1_866
timestamp 1612251222
transform -1 0 24 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_12
timestamp 1612251222
transform 1 0 10252 0 1 4210
box -4 -6 20 206
use FILL  FILL_22_11
timestamp 1612251222
transform 1 0 10236 0 1 4210
box -4 -6 20 206
use FILL  FILL_22_10
timestamp 1612251222
transform 1 0 10220 0 1 4210
box -4 -6 20 206
use FILL  FILL_22_9
timestamp 1612251222
transform 1 0 10204 0 1 4210
box -4 -6 20 206
use FILL  FILL_22_8
timestamp 1612251222
transform 1 0 10188 0 1 4210
box -4 -6 20 206
use FILL  FILL_22_7
timestamp 1612251222
transform 1 0 10172 0 1 4210
box -4 -6 20 206
use FILL  FILL_22_6
timestamp 1612251222
transform 1 0 10156 0 1 4210
box -4 -6 20 206
use FILL  FILL_22_5
timestamp 1612251222
transform 1 0 10140 0 1 4210
box -4 -6 20 206
use FILL  FILL_22_4
timestamp 1612251222
transform 1 0 10124 0 1 4210
box -4 -6 20 206
use FILL  FILL_22_3
timestamp 1612251222
transform 1 0 10108 0 1 4210
box -4 -6 20 206
use FILL  FILL_22_2
timestamp 1612251222
transform 1 0 10092 0 1 4210
box -4 -6 20 206
use FILL  FILL_22_1
timestamp 1612251222
transform 1 0 10076 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_319
timestamp 1612251222
transform 1 0 9910 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_319
timestamp 1612251222
transform 1 0 9894 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_319
timestamp 1612251222
transform 1 0 9878 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_319
timestamp 1612251222
transform 1 0 9862 0 1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_314
timestamp 1612251222
transform -1 0 9862 0 1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_314
timestamp 1612251222
transform -1 0 9696 0 1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_314
timestamp 1612251222
transform -1 0 9680 0 1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_314
timestamp 1612251222
transform -1 0 9664 0 1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_314
timestamp 1612251222
transform -1 0 9648 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_714
timestamp 1612251222
transform -1 0 9632 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_714
timestamp 1612251222
transform -1 0 9466 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_714
timestamp 1612251222
transform -1 0 9450 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_714
timestamp 1612251222
transform -1 0 9434 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_724
timestamp 1612251222
transform -1 0 9418 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_724
timestamp 1612251222
transform -1 0 9252 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_724
timestamp 1612251222
transform -1 0 9236 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_724
timestamp 1612251222
transform -1 0 9220 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_270
timestamp 1612251222
transform -1 0 9204 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_270
timestamp 1612251222
transform -1 0 9038 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_270
timestamp 1612251222
transform -1 0 9022 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_270
timestamp 1612251222
transform -1 0 9006 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_659
timestamp 1612251222
transform 1 0 8824 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_659
timestamp 1612251222
transform 1 0 8808 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_659
timestamp 1612251222
transform 1 0 8792 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_659
timestamp 1612251222
transform 1 0 8776 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_222
timestamp 1612251222
transform 1 0 8610 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_222
timestamp 1612251222
transform 1 0 8594 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_222
timestamp 1612251222
transform 1 0 8578 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_222
timestamp 1612251222
transform 1 0 8562 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_657
timestamp 1612251222
transform 1 0 8396 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_657
timestamp 1612251222
transform 1 0 8380 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_657
timestamp 1612251222
transform 1 0 8364 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_657
timestamp 1612251222
transform 1 0 8348 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_115
timestamp 1612251222
transform 1 0 8182 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_115
timestamp 1612251222
transform 1 0 8166 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_115
timestamp 1612251222
transform 1 0 8150 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_115
timestamp 1612251222
transform 1 0 8134 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_276
timestamp 1612251222
transform -1 0 8134 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_276
timestamp 1612251222
transform -1 0 7968 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_276
timestamp 1612251222
transform -1 0 7952 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_276
timestamp 1612251222
transform -1 0 7936 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_217
timestamp 1612251222
transform -1 0 7920 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_217
timestamp 1612251222
transform -1 0 7754 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_217
timestamp 1612251222
transform -1 0 7738 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_217
timestamp 1612251222
transform -1 0 7722 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_860
timestamp 1612251222
transform 1 0 7540 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_860
timestamp 1612251222
transform 1 0 7524 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_860
timestamp 1612251222
transform 1 0 7508 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_860
timestamp 1612251222
transform 1 0 7492 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_861
timestamp 1612251222
transform -1 0 7492 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_861
timestamp 1612251222
transform -1 0 7326 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_861
timestamp 1612251222
transform -1 0 7310 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_861
timestamp 1612251222
transform -1 0 7294 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_361
timestamp 1612251222
transform -1 0 7278 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_361
timestamp 1612251222
transform -1 0 7112 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_361
timestamp 1612251222
transform -1 0 7096 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_361
timestamp 1612251222
transform -1 0 7080 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_327
timestamp 1612251222
transform -1 0 7064 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_327
timestamp 1612251222
transform -1 0 6898 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_327
timestamp 1612251222
transform -1 0 6882 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_327
timestamp 1612251222
transform -1 0 6866 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_493
timestamp 1612251222
transform -1 0 6850 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_493
timestamp 1612251222
transform -1 0 6684 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_493
timestamp 1612251222
transform -1 0 6668 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_493
timestamp 1612251222
transform -1 0 6652 0 1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_117
timestamp 1612251222
transform -1 0 6636 0 1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_117
timestamp 1612251222
transform -1 0 6470 0 1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_117
timestamp 1612251222
transform -1 0 6454 0 1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_117
timestamp 1612251222
transform -1 0 6438 0 1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_117
timestamp 1612251222
transform -1 0 6422 0 1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_519
timestamp 1612251222
transform -1 0 6406 0 1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_519
timestamp 1612251222
transform -1 0 6240 0 1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_519
timestamp 1612251222
transform -1 0 6224 0 1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_519
timestamp 1612251222
transform -1 0 6208 0 1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_519
timestamp 1612251222
transform -1 0 6192 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_383
timestamp 1612251222
transform -1 0 6176 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_383
timestamp 1612251222
transform -1 0 6010 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_383
timestamp 1612251222
transform -1 0 5994 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_383
timestamp 1612251222
transform -1 0 5978 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_520
timestamp 1612251222
transform -1 0 5962 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_520
timestamp 1612251222
transform -1 0 5796 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_520
timestamp 1612251222
transform -1 0 5780 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_520
timestamp 1612251222
transform -1 0 5764 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_721
timestamp 1612251222
transform 1 0 5582 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_721
timestamp 1612251222
transform 1 0 5566 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_721
timestamp 1612251222
transform 1 0 5550 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_721
timestamp 1612251222
transform 1 0 5534 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_720
timestamp 1612251222
transform 1 0 5368 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_720
timestamp 1612251222
transform 1 0 5352 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_720
timestamp 1612251222
transform 1 0 5336 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_720
timestamp 1612251222
transform 1 0 5320 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_750
timestamp 1612251222
transform -1 0 5320 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_750
timestamp 1612251222
transform -1 0 5154 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_750
timestamp 1612251222
transform -1 0 5138 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_750
timestamp 1612251222
transform -1 0 5122 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_749
timestamp 1612251222
transform -1 0 5106 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_749
timestamp 1612251222
transform -1 0 4940 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_749
timestamp 1612251222
transform -1 0 4924 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_749
timestamp 1612251222
transform -1 0 4908 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_92
timestamp 1612251222
transform -1 0 4892 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_92
timestamp 1612251222
transform -1 0 4726 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_92
timestamp 1612251222
transform -1 0 4710 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_92
timestamp 1612251222
transform -1 0 4694 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_618
timestamp 1612251222
transform 1 0 4512 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_618
timestamp 1612251222
transform 1 0 4496 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_618
timestamp 1612251222
transform 1 0 4480 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_618
timestamp 1612251222
transform 1 0 4464 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_384
timestamp 1612251222
transform 1 0 4298 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_384
timestamp 1612251222
transform 1 0 4282 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_384
timestamp 1612251222
transform 1 0 4266 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_384
timestamp 1612251222
transform 1 0 4250 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_133
timestamp 1612251222
transform -1 0 4250 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_133
timestamp 1612251222
transform -1 0 4084 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_133
timestamp 1612251222
transform -1 0 4068 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_133
timestamp 1612251222
transform -1 0 4052 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_529
timestamp 1612251222
transform -1 0 4036 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_529
timestamp 1612251222
transform -1 0 3870 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_529
timestamp 1612251222
transform -1 0 3854 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_529
timestamp 1612251222
transform -1 0 3838 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_494
timestamp 1612251222
transform -1 0 3822 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_494
timestamp 1612251222
transform -1 0 3656 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_494
timestamp 1612251222
transform -1 0 3640 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_494
timestamp 1612251222
transform -1 0 3624 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_80
timestamp 1612251222
transform -1 0 3608 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_80
timestamp 1612251222
transform -1 0 3442 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_80
timestamp 1612251222
transform -1 0 3426 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_80
timestamp 1612251222
transform -1 0 3410 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_81
timestamp 1612251222
transform -1 0 3394 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_81
timestamp 1612251222
transform -1 0 3228 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_81
timestamp 1612251222
transform -1 0 3212 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_81
timestamp 1612251222
transform -1 0 3196 0 1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_573
timestamp 1612251222
transform -1 0 3180 0 1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_573
timestamp 1612251222
transform -1 0 3014 0 1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_573
timestamp 1612251222
transform -1 0 2998 0 1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_573
timestamp 1612251222
transform -1 0 2982 0 1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_573
timestamp 1612251222
transform -1 0 2966 0 1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_501
timestamp 1612251222
transform 1 0 2784 0 1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_501
timestamp 1612251222
transform 1 0 2768 0 1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_501
timestamp 1612251222
transform 1 0 2752 0 1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_501
timestamp 1612251222
transform 1 0 2736 0 1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_501
timestamp 1612251222
transform 1 0 2720 0 1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_659
timestamp 1612251222
transform -1 0 2720 0 1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_659
timestamp 1612251222
transform -1 0 2554 0 1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_659
timestamp 1612251222
transform -1 0 2538 0 1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_659
timestamp 1612251222
transform -1 0 2522 0 1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_659
timestamp 1612251222
transform -1 0 2506 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_498
timestamp 1612251222
transform 1 0 2324 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_498
timestamp 1612251222
transform 1 0 2308 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_498
timestamp 1612251222
transform 1 0 2292 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_498
timestamp 1612251222
transform 1 0 2276 0 1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_676
timestamp 1612251222
transform -1 0 2276 0 1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_676
timestamp 1612251222
transform -1 0 2110 0 1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_676
timestamp 1612251222
transform -1 0 2094 0 1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_676
timestamp 1612251222
transform -1 0 2078 0 1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_676
timestamp 1612251222
transform -1 0 2062 0 1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_204
timestamp 1612251222
transform -1 0 2046 0 1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_204
timestamp 1612251222
transform -1 0 1880 0 1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_204
timestamp 1612251222
transform -1 0 1864 0 1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_204
timestamp 1612251222
transform -1 0 1848 0 1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_204
timestamp 1612251222
transform -1 0 1832 0 1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_205
timestamp 1612251222
transform -1 0 1816 0 1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_205
timestamp 1612251222
transform -1 0 1650 0 1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_205
timestamp 1612251222
transform -1 0 1634 0 1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_205
timestamp 1612251222
transform -1 0 1618 0 1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_205
timestamp 1612251222
transform -1 0 1602 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_680
timestamp 1612251222
transform 1 0 1420 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_680
timestamp 1612251222
transform 1 0 1404 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_680
timestamp 1612251222
transform 1 0 1388 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_680
timestamp 1612251222
transform 1 0 1372 0 1 4210
box -4 -6 20 206
use POR2X1  POR2X1_187
timestamp 1612251222
transform -1 0 1372 0 1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_187
timestamp 1612251222
transform -1 0 1206 0 1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_187
timestamp 1612251222
transform -1 0 1190 0 1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_187
timestamp 1612251222
transform -1 0 1174 0 1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_740
timestamp 1612251222
transform 1 0 992 0 1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_740
timestamp 1612251222
transform 1 0 976 0 1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_740
timestamp 1612251222
transform 1 0 960 0 1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_740
timestamp 1612251222
transform 1 0 944 0 1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_740
timestamp 1612251222
transform 1 0 928 0 1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_730
timestamp 1612251222
transform -1 0 928 0 1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_730
timestamp 1612251222
transform -1 0 762 0 1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_730
timestamp 1612251222
transform -1 0 746 0 1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_730
timestamp 1612251222
transform -1 0 730 0 1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_730
timestamp 1612251222
transform -1 0 714 0 1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_798
timestamp 1612251222
transform 1 0 532 0 1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_798
timestamp 1612251222
transform 1 0 516 0 1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_798
timestamp 1612251222
transform 1 0 500 0 1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_798
timestamp 1612251222
transform 1 0 484 0 1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_798
timestamp 1612251222
transform 1 0 468 0 1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_807
timestamp 1612251222
transform -1 0 468 0 1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_807
timestamp 1612251222
transform -1 0 302 0 1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_807
timestamp 1612251222
transform -1 0 286 0 1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_807
timestamp 1612251222
transform -1 0 270 0 1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_807
timestamp 1612251222
transform -1 0 254 0 1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_812
timestamp 1612251222
transform -1 0 238 0 1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_812
timestamp 1612251222
transform -1 0 72 0 1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_812
timestamp 1612251222
transform -1 0 56 0 1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_812
timestamp 1612251222
transform -1 0 40 0 1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_812
timestamp 1612251222
transform -1 0 24 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_12
timestamp 1612251222
transform -1 0 10262 0 -1 4210
box -4 -6 20 206
use FILL  FILL_21_11
timestamp 1612251222
transform -1 0 10246 0 -1 4210
box -4 -6 20 206
use FILL  FILL_21_10
timestamp 1612251222
transform -1 0 10230 0 -1 4210
box -4 -6 20 206
use FILL  FILL_21_9
timestamp 1612251222
transform -1 0 10214 0 -1 4210
box -4 -6 20 206
use FILL  FILL_21_8
timestamp 1612251222
transform -1 0 10198 0 -1 4210
box -4 -6 20 206
use FILL  FILL_21_7
timestamp 1612251222
transform -1 0 10182 0 -1 4210
box -4 -6 20 206
use FILL  FILL_21_6
timestamp 1612251222
transform -1 0 10166 0 -1 4210
box -4 -6 20 206
use FILL  FILL_21_5
timestamp 1612251222
transform -1 0 10150 0 -1 4210
box -4 -6 20 206
use FILL  FILL_21_4
timestamp 1612251222
transform -1 0 10134 0 -1 4210
box -4 -6 20 206
use FILL  FILL_21_3
timestamp 1612251222
transform -1 0 10118 0 -1 4210
box -4 -6 20 206
use FILL  FILL_21_2
timestamp 1612251222
transform -1 0 10102 0 -1 4210
box -4 -6 20 206
use FILL  FILL_21_1
timestamp 1612251222
transform -1 0 10086 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_367
timestamp 1612251222
transform 1 0 9904 0 -1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_367
timestamp 1612251222
transform 1 0 9888 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_367
timestamp 1612251222
transform 1 0 9872 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_367
timestamp 1612251222
transform 1 0 9856 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_317
timestamp 1612251222
transform 1 0 9690 0 -1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_317
timestamp 1612251222
transform 1 0 9674 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_317
timestamp 1612251222
transform 1 0 9658 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_317
timestamp 1612251222
transform 1 0 9642 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_704
timestamp 1612251222
transform 1 0 9476 0 -1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_704
timestamp 1612251222
transform 1 0 9460 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_704
timestamp 1612251222
transform 1 0 9444 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_704
timestamp 1612251222
transform 1 0 9428 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_313
timestamp 1612251222
transform 1 0 9262 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_313
timestamp 1612251222
transform 1 0 9246 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_313
timestamp 1612251222
transform 1 0 9230 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_313
timestamp 1612251222
transform 1 0 9214 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_313
timestamp 1612251222
transform 1 0 9198 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_703
timestamp 1612251222
transform 1 0 9032 0 -1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_703
timestamp 1612251222
transform 1 0 9016 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_703
timestamp 1612251222
transform 1 0 9000 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_703
timestamp 1612251222
transform 1 0 8984 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_417
timestamp 1612251222
transform -1 0 8984 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_417
timestamp 1612251222
transform -1 0 8818 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_417
timestamp 1612251222
transform -1 0 8802 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_417
timestamp 1612251222
transform -1 0 8786 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_417
timestamp 1612251222
transform -1 0 8770 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_268
timestamp 1612251222
transform -1 0 8754 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_268
timestamp 1612251222
transform -1 0 8588 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_268
timestamp 1612251222
transform -1 0 8572 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_268
timestamp 1612251222
transform -1 0 8556 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_268
timestamp 1612251222
transform -1 0 8540 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_269
timestamp 1612251222
transform -1 0 8524 0 -1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_269
timestamp 1612251222
transform -1 0 8358 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_269
timestamp 1612251222
transform -1 0 8342 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_269
timestamp 1612251222
transform -1 0 8326 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_271
timestamp 1612251222
transform -1 0 8310 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_271
timestamp 1612251222
transform -1 0 8144 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_271
timestamp 1612251222
transform -1 0 8128 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_271
timestamp 1612251222
transform -1 0 8112 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_271
timestamp 1612251222
transform -1 0 8096 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_366
timestamp 1612251222
transform 1 0 7914 0 -1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_366
timestamp 1612251222
transform 1 0 7898 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_366
timestamp 1612251222
transform 1 0 7882 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_366
timestamp 1612251222
transform 1 0 7866 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_106
timestamp 1612251222
transform -1 0 7866 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_106
timestamp 1612251222
transform -1 0 7700 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_106
timestamp 1612251222
transform -1 0 7684 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_106
timestamp 1612251222
transform -1 0 7668 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_106
timestamp 1612251222
transform -1 0 7652 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_362
timestamp 1612251222
transform 1 0 7470 0 -1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_362
timestamp 1612251222
transform 1 0 7454 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_362
timestamp 1612251222
transform 1 0 7438 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_362
timestamp 1612251222
transform 1 0 7422 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_474
timestamp 1612251222
transform -1 0 7422 0 -1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_474
timestamp 1612251222
transform -1 0 7256 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_474
timestamp 1612251222
transform -1 0 7240 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_474
timestamp 1612251222
transform -1 0 7224 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_218
timestamp 1612251222
transform 1 0 7042 0 -1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_218
timestamp 1612251222
transform 1 0 7026 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_218
timestamp 1612251222
transform 1 0 7010 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_218
timestamp 1612251222
transform 1 0 6994 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_216
timestamp 1612251222
transform 1 0 6828 0 -1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_216
timestamp 1612251222
transform 1 0 6812 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_216
timestamp 1612251222
transform 1 0 6796 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_216
timestamp 1612251222
transform 1 0 6780 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_124
timestamp 1612251222
transform 1 0 6614 0 -1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_124
timestamp 1612251222
transform 1 0 6598 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_124
timestamp 1612251222
transform 1 0 6582 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_124
timestamp 1612251222
transform 1 0 6566 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_123
timestamp 1612251222
transform 1 0 6400 0 -1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_123
timestamp 1612251222
transform 1 0 6384 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_123
timestamp 1612251222
transform 1 0 6368 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_123
timestamp 1612251222
transform 1 0 6352 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_492
timestamp 1612251222
transform 1 0 6186 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_492
timestamp 1612251222
transform 1 0 6170 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_492
timestamp 1612251222
transform 1 0 6154 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_492
timestamp 1612251222
transform 1 0 6138 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_492
timestamp 1612251222
transform 1 0 6122 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_118
timestamp 1612251222
transform 1 0 5956 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_118
timestamp 1612251222
transform 1 0 5940 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_118
timestamp 1612251222
transform 1 0 5924 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_118
timestamp 1612251222
transform 1 0 5908 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_118
timestamp 1612251222
transform 1 0 5892 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_518
timestamp 1612251222
transform 1 0 5726 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_518
timestamp 1612251222
transform 1 0 5710 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_518
timestamp 1612251222
transform 1 0 5694 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_518
timestamp 1612251222
transform 1 0 5678 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_518
timestamp 1612251222
transform 1 0 5662 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_384
timestamp 1612251222
transform -1 0 5662 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_384
timestamp 1612251222
transform -1 0 5496 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_384
timestamp 1612251222
transform -1 0 5480 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_384
timestamp 1612251222
transform -1 0 5464 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_384
timestamp 1612251222
transform -1 0 5448 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_668
timestamp 1612251222
transform -1 0 5432 0 -1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_668
timestamp 1612251222
transform -1 0 5266 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_668
timestamp 1612251222
transform -1 0 5250 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_668
timestamp 1612251222
transform -1 0 5234 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_669
timestamp 1612251222
transform 1 0 5052 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_669
timestamp 1612251222
transform 1 0 5036 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_669
timestamp 1612251222
transform 1 0 5020 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_669
timestamp 1612251222
transform 1 0 5004 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_669
timestamp 1612251222
transform 1 0 4988 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_750
timestamp 1612251222
transform -1 0 4988 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_750
timestamp 1612251222
transform -1 0 4822 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_750
timestamp 1612251222
transform -1 0 4806 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_750
timestamp 1612251222
transform -1 0 4790 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_750
timestamp 1612251222
transform -1 0 4774 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_751
timestamp 1612251222
transform -1 0 4758 0 -1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_751
timestamp 1612251222
transform -1 0 4592 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_751
timestamp 1612251222
transform -1 0 4576 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_751
timestamp 1612251222
transform -1 0 4560 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_391
timestamp 1612251222
transform -1 0 4544 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_391
timestamp 1612251222
transform -1 0 4378 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_391
timestamp 1612251222
transform -1 0 4362 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_391
timestamp 1612251222
transform -1 0 4346 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_391
timestamp 1612251222
transform -1 0 4330 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_383
timestamp 1612251222
transform 1 0 4148 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_383
timestamp 1612251222
transform 1 0 4132 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_383
timestamp 1612251222
transform 1 0 4116 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_383
timestamp 1612251222
transform 1 0 4100 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_383
timestamp 1612251222
transform 1 0 4084 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_392
timestamp 1612251222
transform -1 0 4084 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_392
timestamp 1612251222
transform -1 0 3918 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_392
timestamp 1612251222
transform -1 0 3902 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_392
timestamp 1612251222
transform -1 0 3886 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_392
timestamp 1612251222
transform -1 0 3870 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_171
timestamp 1612251222
transform -1 0 3854 0 -1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_171
timestamp 1612251222
transform -1 0 3688 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_171
timestamp 1612251222
transform -1 0 3672 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_171
timestamp 1612251222
transform -1 0 3656 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_658
timestamp 1612251222
transform -1 0 3640 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_658
timestamp 1612251222
transform -1 0 3474 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_658
timestamp 1612251222
transform -1 0 3458 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_658
timestamp 1612251222
transform -1 0 3442 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_658
timestamp 1612251222
transform -1 0 3426 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_735
timestamp 1612251222
transform -1 0 3410 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_735
timestamp 1612251222
transform -1 0 3244 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_735
timestamp 1612251222
transform -1 0 3228 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_735
timestamp 1612251222
transform -1 0 3212 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_735
timestamp 1612251222
transform -1 0 3196 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_72
timestamp 1612251222
transform -1 0 3180 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_POR2X1_72
timestamp 1612251222
transform -1 0 3014 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_POR2X1_72
timestamp 1612251222
transform -1 0 2998 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_72
timestamp 1612251222
transform -1 0 2982 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_72
timestamp 1612251222
transform -1 0 2966 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_657
timestamp 1612251222
transform -1 0 2950 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_657
timestamp 1612251222
transform -1 0 2784 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_657
timestamp 1612251222
transform -1 0 2768 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_657
timestamp 1612251222
transform -1 0 2752 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_657
timestamp 1612251222
transform -1 0 2736 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_203
timestamp 1612251222
transform -1 0 2720 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_203
timestamp 1612251222
transform -1 0 2554 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_203
timestamp 1612251222
transform -1 0 2538 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_203
timestamp 1612251222
transform -1 0 2522 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_203
timestamp 1612251222
transform -1 0 2506 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_188
timestamp 1612251222
transform -1 0 2490 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_188
timestamp 1612251222
transform -1 0 2324 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_188
timestamp 1612251222
transform -1 0 2308 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_188
timestamp 1612251222
transform -1 0 2292 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_188
timestamp 1612251222
transform -1 0 2276 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_189
timestamp 1612251222
transform -1 0 2260 0 -1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_189
timestamp 1612251222
transform -1 0 2094 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_189
timestamp 1612251222
transform -1 0 2078 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_189
timestamp 1612251222
transform -1 0 2062 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_679
timestamp 1612251222
transform -1 0 2046 0 -1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_679
timestamp 1612251222
transform -1 0 1880 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_679
timestamp 1612251222
transform -1 0 1864 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_679
timestamp 1612251222
transform -1 0 1848 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_728
timestamp 1612251222
transform -1 0 1832 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_728
timestamp 1612251222
transform -1 0 1666 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_728
timestamp 1612251222
transform -1 0 1650 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_728
timestamp 1612251222
transform -1 0 1634 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_728
timestamp 1612251222
transform -1 0 1618 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_192
timestamp 1612251222
transform -1 0 1602 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_192
timestamp 1612251222
transform -1 0 1436 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_192
timestamp 1612251222
transform -1 0 1420 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_192
timestamp 1612251222
transform -1 0 1404 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_192
timestamp 1612251222
transform -1 0 1388 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_191
timestamp 1612251222
transform 1 0 1206 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_191
timestamp 1612251222
transform 1 0 1190 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_191
timestamp 1612251222
transform 1 0 1174 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_191
timestamp 1612251222
transform 1 0 1158 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_191
timestamp 1612251222
transform 1 0 1142 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_221
timestamp 1612251222
transform -1 0 1142 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_221
timestamp 1612251222
transform -1 0 976 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_221
timestamp 1612251222
transform -1 0 960 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_221
timestamp 1612251222
transform -1 0 944 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_221
timestamp 1612251222
transform -1 0 928 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_739
timestamp 1612251222
transform 1 0 746 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_739
timestamp 1612251222
transform 1 0 730 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_739
timestamp 1612251222
transform 1 0 714 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_739
timestamp 1612251222
transform 1 0 698 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_739
timestamp 1612251222
transform 1 0 682 0 -1 4210
box -4 -6 20 206
use POR2X1  POR2X1_79
timestamp 1612251222
transform 1 0 516 0 -1 4210
box -4 -6 170 206
use FILL  FILL1_POR2X1_79
timestamp 1612251222
transform 1 0 500 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_POR2X1_79
timestamp 1612251222
transform 1 0 484 0 -1 4210
box -4 -6 20 206
use FILL  FILL_POR2X1_79
timestamp 1612251222
transform 1 0 468 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_805
timestamp 1612251222
transform 1 0 302 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_805
timestamp 1612251222
transform 1 0 286 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_805
timestamp 1612251222
transform 1 0 270 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_805
timestamp 1612251222
transform 1 0 254 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_805
timestamp 1612251222
transform 1 0 238 0 -1 4210
box -4 -6 20 206
use PAND2X1  PAND2X1_811
timestamp 1612251222
transform -1 0 238 0 -1 4210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_811
timestamp 1612251222
transform -1 0 72 0 -1 4210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_811
timestamp 1612251222
transform -1 0 56 0 -1 4210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_811
timestamp 1612251222
transform -1 0 40 0 -1 4210
box -4 -6 20 206
use FILL  FILL_PAND2X1_811
timestamp 1612251222
transform -1 0 24 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_2
timestamp 1612251222
transform 1 0 10252 0 1 3810
box -4 -6 20 206
use FILL  FILL_20_1
timestamp 1612251222
transform 1 0 10236 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_364
timestamp 1612251222
transform 1 0 10070 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_364
timestamp 1612251222
transform 1 0 10054 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_364
timestamp 1612251222
transform 1 0 10038 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_364
timestamp 1612251222
transform 1 0 10022 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_212
timestamp 1612251222
transform 1 0 9856 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_212
timestamp 1612251222
transform 1 0 9840 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_212
timestamp 1612251222
transform 1 0 9824 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_212
timestamp 1612251222
transform 1 0 9808 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_352
timestamp 1612251222
transform 1 0 9642 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_352
timestamp 1612251222
transform 1 0 9626 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_352
timestamp 1612251222
transform 1 0 9610 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_352
timestamp 1612251222
transform 1 0 9594 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_167
timestamp 1612251222
transform 1 0 9428 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_167
timestamp 1612251222
transform 1 0 9412 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_167
timestamp 1612251222
transform 1 0 9396 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_167
timestamp 1612251222
transform 1 0 9380 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_167
timestamp 1612251222
transform 1 0 9364 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_179
timestamp 1612251222
transform 1 0 9198 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_179
timestamp 1612251222
transform 1 0 9182 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_179
timestamp 1612251222
transform 1 0 9166 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_179
timestamp 1612251222
transform 1 0 9150 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_179
timestamp 1612251222
transform 1 0 9134 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_176
timestamp 1612251222
transform -1 0 9134 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_176
timestamp 1612251222
transform -1 0 8968 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_176
timestamp 1612251222
transform -1 0 8952 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_176
timestamp 1612251222
transform -1 0 8936 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_176
timestamp 1612251222
transform -1 0 8920 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_388
timestamp 1612251222
transform -1 0 8904 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_388
timestamp 1612251222
transform -1 0 8738 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_388
timestamp 1612251222
transform -1 0 8722 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_388
timestamp 1612251222
transform -1 0 8706 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_538
timestamp 1612251222
transform 1 0 8524 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_538
timestamp 1612251222
transform 1 0 8508 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_538
timestamp 1612251222
transform 1 0 8492 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_538
timestamp 1612251222
transform 1 0 8476 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_336
timestamp 1612251222
transform -1 0 8476 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_336
timestamp 1612251222
transform -1 0 8310 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_336
timestamp 1612251222
transform -1 0 8294 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_336
timestamp 1612251222
transform -1 0 8278 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_303
timestamp 1612251222
transform 1 0 8096 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_303
timestamp 1612251222
transform 1 0 8080 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_303
timestamp 1612251222
transform 1 0 8064 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_303
timestamp 1612251222
transform 1 0 8048 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_716
timestamp 1612251222
transform 1 0 7882 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_716
timestamp 1612251222
transform 1 0 7866 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_716
timestamp 1612251222
transform 1 0 7850 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_716
timestamp 1612251222
transform 1 0 7834 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_723
timestamp 1612251222
transform 1 0 7668 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_723
timestamp 1612251222
transform 1 0 7652 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_723
timestamp 1612251222
transform 1 0 7636 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_723
timestamp 1612251222
transform 1 0 7620 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_105
timestamp 1612251222
transform 1 0 7454 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_105
timestamp 1612251222
transform 1 0 7438 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_105
timestamp 1612251222
transform 1 0 7422 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_105
timestamp 1612251222
transform 1 0 7406 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_717
timestamp 1612251222
transform -1 0 7406 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_717
timestamp 1612251222
transform -1 0 7240 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_717
timestamp 1612251222
transform -1 0 7224 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_717
timestamp 1612251222
transform -1 0 7208 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_116
timestamp 1612251222
transform -1 0 7192 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_116
timestamp 1612251222
transform -1 0 7026 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_116
timestamp 1612251222
transform -1 0 7010 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_116
timestamp 1612251222
transform -1 0 6994 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_392
timestamp 1612251222
transform 1 0 6812 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_392
timestamp 1612251222
transform 1 0 6796 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_392
timestamp 1612251222
transform 1 0 6780 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_392
timestamp 1612251222
transform 1 0 6764 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_473
timestamp 1612251222
transform -1 0 6764 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_473
timestamp 1612251222
transform -1 0 6598 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_473
timestamp 1612251222
transform -1 0 6582 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_473
timestamp 1612251222
transform -1 0 6566 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_137
timestamp 1612251222
transform 1 0 6384 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_137
timestamp 1612251222
transform 1 0 6368 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_137
timestamp 1612251222
transform 1 0 6352 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_137
timestamp 1612251222
transform 1 0 6336 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_134
timestamp 1612251222
transform 1 0 6170 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_134
timestamp 1612251222
transform 1 0 6154 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_134
timestamp 1612251222
transform 1 0 6138 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_134
timestamp 1612251222
transform 1 0 6122 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_134
timestamp 1612251222
transform 1 0 6106 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_634
timestamp 1612251222
transform -1 0 6106 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_634
timestamp 1612251222
transform -1 0 5940 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_634
timestamp 1612251222
transform -1 0 5924 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_634
timestamp 1612251222
transform -1 0 5908 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_132
timestamp 1612251222
transform -1 0 5892 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_132
timestamp 1612251222
transform -1 0 5726 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_132
timestamp 1612251222
transform -1 0 5710 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_132
timestamp 1612251222
transform -1 0 5694 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_132
timestamp 1612251222
transform -1 0 5678 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_412
timestamp 1612251222
transform 1 0 5496 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_412
timestamp 1612251222
transform 1 0 5480 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_412
timestamp 1612251222
transform 1 0 5464 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_412
timestamp 1612251222
transform 1 0 5448 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_412
timestamp 1612251222
transform 1 0 5432 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_391
timestamp 1612251222
transform 1 0 5266 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_391
timestamp 1612251222
transform 1 0 5250 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_391
timestamp 1612251222
transform 1 0 5234 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_391
timestamp 1612251222
transform 1 0 5218 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_526
timestamp 1612251222
transform 1 0 5052 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_526
timestamp 1612251222
transform 1 0 5036 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_526
timestamp 1612251222
transform 1 0 5020 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_526
timestamp 1612251222
transform 1 0 5004 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_526
timestamp 1612251222
transform 1 0 4988 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_381
timestamp 1612251222
transform 1 0 4822 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_381
timestamp 1612251222
transform 1 0 4806 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_381
timestamp 1612251222
transform 1 0 4790 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_381
timestamp 1612251222
transform 1 0 4774 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_381
timestamp 1612251222
transform 1 0 4758 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_619
timestamp 1612251222
transform 1 0 4592 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_619
timestamp 1612251222
transform 1 0 4576 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_619
timestamp 1612251222
transform 1 0 4560 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_619
timestamp 1612251222
transform 1 0 4544 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_414
timestamp 1612251222
transform 1 0 4378 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_414
timestamp 1612251222
transform 1 0 4362 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_414
timestamp 1612251222
transform 1 0 4346 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_414
timestamp 1612251222
transform 1 0 4330 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_414
timestamp 1612251222
transform 1 0 4314 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_789
timestamp 1612251222
transform -1 0 4314 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_789
timestamp 1612251222
transform -1 0 4148 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_789
timestamp 1612251222
transform -1 0 4132 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_789
timestamp 1612251222
transform -1 0 4116 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_789
timestamp 1612251222
transform -1 0 4100 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_67
timestamp 1612251222
transform 1 0 3918 0 1 3810
box -4 -6 170 206
use FILL  FILL2_POR2X1_67
timestamp 1612251222
transform 1 0 3902 0 1 3810
box -4 -6 20 206
use FILL  FILL1_POR2X1_67
timestamp 1612251222
transform 1 0 3886 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_67
timestamp 1612251222
transform 1 0 3870 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_67
timestamp 1612251222
transform 1 0 3854 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_548
timestamp 1612251222
transform -1 0 3854 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_548
timestamp 1612251222
transform -1 0 3688 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_548
timestamp 1612251222
transform -1 0 3672 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_548
timestamp 1612251222
transform -1 0 3656 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_548
timestamp 1612251222
transform -1 0 3640 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_185
timestamp 1612251222
transform -1 0 3624 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_185
timestamp 1612251222
transform -1 0 3458 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_185
timestamp 1612251222
transform -1 0 3442 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_185
timestamp 1612251222
transform -1 0 3426 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_185
timestamp 1612251222
transform -1 0 3410 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_860
timestamp 1612251222
transform -1 0 3394 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_860
timestamp 1612251222
transform -1 0 3228 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_860
timestamp 1612251222
transform -1 0 3212 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_860
timestamp 1612251222
transform -1 0 3196 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_860
timestamp 1612251222
transform -1 0 3180 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_510
timestamp 1612251222
transform -1 0 3164 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_510
timestamp 1612251222
transform -1 0 2998 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_510
timestamp 1612251222
transform -1 0 2982 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_510
timestamp 1612251222
transform -1 0 2966 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_510
timestamp 1612251222
transform -1 0 2950 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_574
timestamp 1612251222
transform -1 0 2934 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_574
timestamp 1612251222
transform -1 0 2768 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_574
timestamp 1612251222
transform -1 0 2752 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_574
timestamp 1612251222
transform -1 0 2736 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_574
timestamp 1612251222
transform -1 0 2720 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_184
timestamp 1612251222
transform -1 0 2704 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_184
timestamp 1612251222
transform -1 0 2538 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_184
timestamp 1612251222
transform -1 0 2522 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_184
timestamp 1612251222
transform -1 0 2506 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_575
timestamp 1612251222
transform -1 0 2490 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_575
timestamp 1612251222
transform -1 0 2324 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_575
timestamp 1612251222
transform -1 0 2308 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_575
timestamp 1612251222
transform -1 0 2292 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_575
timestamp 1612251222
transform -1 0 2276 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_579
timestamp 1612251222
transform -1 0 2260 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_579
timestamp 1612251222
transform -1 0 2094 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_579
timestamp 1612251222
transform -1 0 2078 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_579
timestamp 1612251222
transform -1 0 2062 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_579
timestamp 1612251222
transform -1 0 2046 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_468
timestamp 1612251222
transform 1 0 1864 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_468
timestamp 1612251222
transform 1 0 1848 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_468
timestamp 1612251222
transform 1 0 1832 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_468
timestamp 1612251222
transform 1 0 1816 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_468
timestamp 1612251222
transform 1 0 1800 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_794
timestamp 1612251222
transform -1 0 1800 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_794
timestamp 1612251222
transform -1 0 1634 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_794
timestamp 1612251222
transform -1 0 1618 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_794
timestamp 1612251222
transform -1 0 1602 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_794
timestamp 1612251222
transform -1 0 1586 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_440
timestamp 1612251222
transform 1 0 1404 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_440
timestamp 1612251222
transform 1 0 1388 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_440
timestamp 1612251222
transform 1 0 1372 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_440
timestamp 1612251222
transform 1 0 1356 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_440
timestamp 1612251222
transform 1 0 1340 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_437
timestamp 1612251222
transform 1 0 1174 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_437
timestamp 1612251222
transform 1 0 1158 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_437
timestamp 1612251222
transform 1 0 1142 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_437
timestamp 1612251222
transform 1 0 1126 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_487
timestamp 1612251222
transform -1 0 1126 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_487
timestamp 1612251222
transform -1 0 960 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_487
timestamp 1612251222
transform -1 0 944 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_487
timestamp 1612251222
transform -1 0 928 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_489
timestamp 1612251222
transform -1 0 912 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_489
timestamp 1612251222
transform -1 0 746 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_489
timestamp 1612251222
transform -1 0 730 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_489
timestamp 1612251222
transform -1 0 714 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_489
timestamp 1612251222
transform -1 0 698 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_78
timestamp 1612251222
transform -1 0 682 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_78
timestamp 1612251222
transform -1 0 516 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_78
timestamp 1612251222
transform -1 0 500 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_78
timestamp 1612251222
transform -1 0 484 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_78
timestamp 1612251222
transform -1 0 468 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_767
timestamp 1612251222
transform -1 0 452 0 1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_767
timestamp 1612251222
transform -1 0 286 0 1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_767
timestamp 1612251222
transform -1 0 270 0 1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_767
timestamp 1612251222
transform -1 0 254 0 1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_774
timestamp 1612251222
transform -1 0 238 0 1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_774
timestamp 1612251222
transform -1 0 72 0 1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_774
timestamp 1612251222
transform -1 0 56 0 1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_774
timestamp 1612251222
transform -1 0 40 0 1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_774
timestamp 1612251222
transform -1 0 24 0 1 3810
box -4 -6 20 206
use POR2X1  POR2X1_365
timestamp 1612251222
transform -1 0 10268 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_365
timestamp 1612251222
transform -1 0 10102 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_365
timestamp 1612251222
transform -1 0 10086 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_365
timestamp 1612251222
transform -1 0 10070 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_353
timestamp 1612251222
transform 1 0 10102 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_353
timestamp 1612251222
transform 1 0 10086 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_353
timestamp 1612251222
transform 1 0 10070 0 1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_353
timestamp 1612251222
transform 1 0 10054 0 1 3410
box -4 -6 20 206
use POR2X1  POR2X1_357
timestamp 1612251222
transform 1 0 9888 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_357
timestamp 1612251222
transform 1 0 9872 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_357
timestamp 1612251222
transform 1 0 9856 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_357
timestamp 1612251222
transform 1 0 9840 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_443
timestamp 1612251222
transform 1 0 9888 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_443
timestamp 1612251222
transform 1 0 9872 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_443
timestamp 1612251222
transform 1 0 9856 0 1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_443
timestamp 1612251222
transform 1 0 9840 0 1 3410
box -4 -6 20 206
use POR2X1  POR2X1_182
timestamp 1612251222
transform 1 0 9674 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_182
timestamp 1612251222
transform 1 0 9658 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_182
timestamp 1612251222
transform 1 0 9642 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_182
timestamp 1612251222
transform 1 0 9626 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_441
timestamp 1612251222
transform 1 0 9674 0 1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_441
timestamp 1612251222
transform 1 0 9658 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_441
timestamp 1612251222
transform 1 0 9642 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_441
timestamp 1612251222
transform 1 0 9626 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_441
timestamp 1612251222
transform 1 0 9610 0 1 3410
box -4 -6 20 206
use POR2X1  POR2X1_180
timestamp 1612251222
transform 1 0 9460 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_180
timestamp 1612251222
transform 1 0 9444 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_524
timestamp 1612251222
transform 1 0 9444 0 1 3410
box -4 -6 170 206
use FILL  FILL0_POR2X1_180
timestamp 1612251222
transform 1 0 9428 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_180
timestamp 1612251222
transform 1 0 9412 0 -1 3810
box -4 -6 20 206
use FILL  FILL2_PAND2X1_524
timestamp 1612251222
transform 1 0 9428 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_524
timestamp 1612251222
transform 1 0 9412 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_524
timestamp 1612251222
transform 1 0 9396 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_524
timestamp 1612251222
transform 1 0 9380 0 1 3410
box -4 -6 20 206
use POR2X1  POR2X1_181
timestamp 1612251222
transform 1 0 9246 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_181
timestamp 1612251222
transform 1 0 9230 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_181
timestamp 1612251222
transform 1 0 9214 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_181
timestamp 1612251222
transform 1 0 9198 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_471
timestamp 1612251222
transform 1 0 9214 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_471
timestamp 1612251222
transform 1 0 9198 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_471
timestamp 1612251222
transform 1 0 9182 0 1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_471
timestamp 1612251222
transform 1 0 9166 0 1 3410
box -4 -6 20 206
use POR2X1  POR2X1_540
timestamp 1612251222
transform -1 0 9198 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_540
timestamp 1612251222
transform -1 0 9032 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_540
timestamp 1612251222
transform -1 0 9016 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_540
timestamp 1612251222
transform -1 0 9000 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_543
timestamp 1612251222
transform 1 0 9000 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_543
timestamp 1612251222
transform 1 0 8984 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_543
timestamp 1612251222
transform 1 0 8968 0 1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_543
timestamp 1612251222
transform 1 0 8952 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_178
timestamp 1612251222
transform 1 0 8818 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_178
timestamp 1612251222
transform 1 0 8802 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_178
timestamp 1612251222
transform 1 0 8786 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_178
timestamp 1612251222
transform 1 0 8770 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_178
timestamp 1612251222
transform 1 0 8754 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_312
timestamp 1612251222
transform 1 0 8786 0 1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_312
timestamp 1612251222
transform 1 0 8770 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_312
timestamp 1612251222
transform 1 0 8754 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_312
timestamp 1612251222
transform 1 0 8738 0 1 3410
box -4 -6 20 206
use POR2X1  POR2X1_337
timestamp 1612251222
transform 1 0 8588 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_337
timestamp 1612251222
transform 1 0 8572 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_312
timestamp 1612251222
transform 1 0 8722 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_337
timestamp 1612251222
transform 1 0 8556 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_337
timestamp 1612251222
transform 1 0 8540 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_370
timestamp 1612251222
transform 1 0 8556 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_370
timestamp 1612251222
transform 1 0 8540 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_370
timestamp 1612251222
transform 1 0 8524 0 1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_370
timestamp 1612251222
transform 1 0 8508 0 1 3410
box -4 -6 20 206
use POR2X1  POR2X1_335
timestamp 1612251222
transform 1 0 8374 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_335
timestamp 1612251222
transform 1 0 8358 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_335
timestamp 1612251222
transform 1 0 8342 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_335
timestamp 1612251222
transform 1 0 8326 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_309
timestamp 1612251222
transform -1 0 8508 0 1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_309
timestamp 1612251222
transform -1 0 8342 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_309
timestamp 1612251222
transform -1 0 8326 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_309
timestamp 1612251222
transform -1 0 8310 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_309
timestamp 1612251222
transform -1 0 8294 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_311
timestamp 1612251222
transform 1 0 8160 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_311
timestamp 1612251222
transform 1 0 8144 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_311
timestamp 1612251222
transform 1 0 8128 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_311
timestamp 1612251222
transform 1 0 8112 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_311
timestamp 1612251222
transform 1 0 8096 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_831
timestamp 1612251222
transform 1 0 8112 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_831
timestamp 1612251222
transform 1 0 8096 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_831
timestamp 1612251222
transform 1 0 8080 0 1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_831
timestamp 1612251222
transform 1 0 8064 0 1 3410
box -4 -6 20 206
use POR2X1  POR2X1_301
timestamp 1612251222
transform -1 0 8096 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_301
timestamp 1612251222
transform -1 0 7930 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_301
timestamp 1612251222
transform -1 0 7914 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_301
timestamp 1612251222
transform -1 0 7898 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_273
timestamp 1612251222
transform 1 0 7898 0 1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_273
timestamp 1612251222
transform 1 0 7882 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_273
timestamp 1612251222
transform 1 0 7866 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_498
timestamp 1612251222
transform -1 0 7882 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_498
timestamp 1612251222
transform -1 0 7716 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_273
timestamp 1612251222
transform 1 0 7850 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_273
timestamp 1612251222
transform 1 0 7834 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_498
timestamp 1612251222
transform -1 0 7700 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_498
timestamp 1612251222
transform -1 0 7684 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_498
timestamp 1612251222
transform -1 0 7668 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_251
timestamp 1612251222
transform 1 0 7668 0 1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_251
timestamp 1612251222
transform 1 0 7652 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_251
timestamp 1612251222
transform 1 0 7636 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_251
timestamp 1612251222
transform 1 0 7620 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_251
timestamp 1612251222
transform 1 0 7604 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_310
timestamp 1612251222
transform 1 0 7486 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_310
timestamp 1612251222
transform 1 0 7470 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_310
timestamp 1612251222
transform 1 0 7454 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_310
timestamp 1612251222
transform 1 0 7438 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_310
timestamp 1612251222
transform 1 0 7422 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_778
timestamp 1612251222
transform -1 0 7604 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_778
timestamp 1612251222
transform -1 0 7438 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_778
timestamp 1612251222
transform -1 0 7422 0 1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_778
timestamp 1612251222
transform -1 0 7406 0 1 3410
box -4 -6 20 206
use POR2X1  POR2X1_114
timestamp 1612251222
transform -1 0 7422 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_114
timestamp 1612251222
transform -1 0 7256 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_114
timestamp 1612251222
transform -1 0 7240 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_114
timestamp 1612251222
transform -1 0 7224 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_372
timestamp 1612251222
transform 1 0 7224 0 1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_372
timestamp 1612251222
transform 1 0 7208 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_372
timestamp 1612251222
transform 1 0 7192 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_372
timestamp 1612251222
transform 1 0 7176 0 1 3410
box -4 -6 20 206
use POR2X1  POR2X1_390
timestamp 1612251222
transform -1 0 7208 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_390
timestamp 1612251222
transform -1 0 7042 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_390
timestamp 1612251222
transform -1 0 7026 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_390
timestamp 1612251222
transform -1 0 7010 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_372
timestamp 1612251222
transform 1 0 7160 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_103
timestamp 1612251222
transform -1 0 7160 0 1 3410
box -4 -6 170 206
use PAND2X1  PAND2X1_153
timestamp 1612251222
transform -1 0 6994 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_103
timestamp 1612251222
transform -1 0 6994 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_103
timestamp 1612251222
transform -1 0 6978 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_103
timestamp 1612251222
transform -1 0 6962 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_103
timestamp 1612251222
transform -1 0 6946 0 1 3410
box -4 -6 20 206
use FILL  FILL2_PAND2X1_153
timestamp 1612251222
transform -1 0 6828 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_153
timestamp 1612251222
transform -1 0 6812 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_153
timestamp 1612251222
transform -1 0 6796 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_153
timestamp 1612251222
transform -1 0 6780 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_772
timestamp 1612251222
transform 1 0 6764 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_772
timestamp 1612251222
transform 1 0 6748 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_772
timestamp 1612251222
transform 1 0 6732 0 1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_772
timestamp 1612251222
transform 1 0 6716 0 1 3410
box -4 -6 20 206
use POR2X1  POR2X1_650
timestamp 1612251222
transform 1 0 6598 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_650
timestamp 1612251222
transform 1 0 6582 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_650
timestamp 1612251222
transform 1 0 6566 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_650
timestamp 1612251222
transform 1 0 6550 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_768
timestamp 1612251222
transform 1 0 6550 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_768
timestamp 1612251222
transform 1 0 6534 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_768
timestamp 1612251222
transform 1 0 6518 0 1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_768
timestamp 1612251222
transform 1 0 6502 0 1 3410
box -4 -6 20 206
use POR2X1  POR2X1_113
timestamp 1612251222
transform 1 0 6384 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_113
timestamp 1612251222
transform 1 0 6368 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_113
timestamp 1612251222
transform 1 0 6352 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_113
timestamp 1612251222
transform 1 0 6336 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_489
timestamp 1612251222
transform 1 0 6336 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_489
timestamp 1612251222
transform 1 0 6320 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_489
timestamp 1612251222
transform 1 0 6304 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_107
timestamp 1612251222
transform 1 0 6170 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_107
timestamp 1612251222
transform 1 0 6154 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_107
timestamp 1612251222
transform 1 0 6138 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_107
timestamp 1612251222
transform 1 0 6122 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_489
timestamp 1612251222
transform 1 0 6288 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_488
timestamp 1612251222
transform 1 0 6122 0 1 3410
box -4 -6 170 206
use FILL  FILL_PAND2X1_107
timestamp 1612251222
transform 1 0 6106 0 -1 3810
box -4 -6 20 206
use FILL  FILL2_PAND2X1_488
timestamp 1612251222
transform 1 0 6106 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_488
timestamp 1612251222
transform 1 0 6090 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_488
timestamp 1612251222
transform 1 0 6074 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_488
timestamp 1612251222
transform 1 0 6058 0 1 3410
box -4 -6 20 206
use POR2X1  POR2X1_640
timestamp 1612251222
transform 1 0 5940 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_640
timestamp 1612251222
transform 1 0 5924 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_640
timestamp 1612251222
transform 1 0 5908 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_640
timestamp 1612251222
transform 1 0 5892 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_278
timestamp 1612251222
transform 1 0 5892 0 1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_278
timestamp 1612251222
transform 1 0 5876 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_278
timestamp 1612251222
transform 1 0 5860 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_278
timestamp 1612251222
transform 1 0 5844 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_278
timestamp 1612251222
transform 1 0 5828 0 1 3410
box -4 -6 20 206
use POR2X1  POR2X1_633
timestamp 1612251222
transform 1 0 5726 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_633
timestamp 1612251222
transform 1 0 5710 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_633
timestamp 1612251222
transform 1 0 5694 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_633
timestamp 1612251222
transform 1 0 5678 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_818
timestamp 1612251222
transform -1 0 5828 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_818
timestamp 1612251222
transform -1 0 5662 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_818
timestamp 1612251222
transform -1 0 5646 0 1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_818
timestamp 1612251222
transform -1 0 5630 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_277
timestamp 1612251222
transform 1 0 5512 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_277
timestamp 1612251222
transform 1 0 5496 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_277
timestamp 1612251222
transform 1 0 5480 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_277
timestamp 1612251222
transform 1 0 5464 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_277
timestamp 1612251222
transform 1 0 5448 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_751
timestamp 1612251222
transform 1 0 5448 0 1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_751
timestamp 1612251222
transform 1 0 5432 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_382
timestamp 1612251222
transform -1 0 5448 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_382
timestamp 1612251222
transform -1 0 5282 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_382
timestamp 1612251222
transform -1 0 5266 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_751
timestamp 1612251222
transform 1 0 5416 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_751
timestamp 1612251222
transform 1 0 5400 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_751
timestamp 1612251222
transform 1 0 5384 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_382
timestamp 1612251222
transform -1 0 5250 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_382
timestamp 1612251222
transform -1 0 5234 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_415
timestamp 1612251222
transform -1 0 5384 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_415
timestamp 1612251222
transform -1 0 5218 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_415
timestamp 1612251222
transform -1 0 5202 0 1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_415
timestamp 1612251222
transform -1 0 5186 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_621
timestamp 1612251222
transform -1 0 5170 0 1 3410
box -4 -6 170 206
use PAND2X1  PAND2X1_817
timestamp 1612251222
transform -1 0 5218 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_621
timestamp 1612251222
transform -1 0 5004 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_817
timestamp 1612251222
transform -1 0 5004 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_817
timestamp 1612251222
transform -1 0 5020 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_817
timestamp 1612251222
transform -1 0 5036 0 -1 3810
box -4 -6 20 206
use FILL  FILL2_PAND2X1_817
timestamp 1612251222
transform -1 0 5052 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_621
timestamp 1612251222
transform -1 0 4956 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_621
timestamp 1612251222
transform -1 0 4972 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_621
timestamp 1612251222
transform -1 0 4988 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_622
timestamp 1612251222
transform -1 0 4988 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_622
timestamp 1612251222
transform -1 0 4822 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_622
timestamp 1612251222
transform -1 0 4806 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_622
timestamp 1612251222
transform -1 0 4790 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_622
timestamp 1612251222
transform -1 0 4774 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_617
timestamp 1612251222
transform 1 0 4774 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_617
timestamp 1612251222
transform 1 0 4758 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_617
timestamp 1612251222
transform 1 0 4742 0 1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_617
timestamp 1612251222
transform 1 0 4726 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_624
timestamp 1612251222
transform -1 0 4758 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_624
timestamp 1612251222
transform -1 0 4592 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_624
timestamp 1612251222
transform -1 0 4576 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_66
timestamp 1612251222
transform 1 0 4560 0 1 3410
box -4 -6 170 206
use FILL  FILL0_PAND2X1_624
timestamp 1612251222
transform -1 0 4560 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_624
timestamp 1612251222
transform -1 0 4544 0 -1 3810
box -4 -6 20 206
use FILL  FILL2_PAND2X1_66
timestamp 1612251222
transform 1 0 4544 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_66
timestamp 1612251222
transform 1 0 4528 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_66
timestamp 1612251222
transform 1 0 4512 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_66
timestamp 1612251222
transform 1 0 4496 0 1 3410
box -4 -6 20 206
use POR2X1  POR2X1_748
timestamp 1612251222
transform -1 0 4528 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_748
timestamp 1612251222
transform -1 0 4362 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_748
timestamp 1612251222
transform -1 0 4346 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_748
timestamp 1612251222
transform -1 0 4330 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_154
timestamp 1612251222
transform -1 0 4496 0 1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_154
timestamp 1612251222
transform -1 0 4330 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_154
timestamp 1612251222
transform -1 0 4314 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_154
timestamp 1612251222
transform -1 0 4298 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_154
timestamp 1612251222
transform -1 0 4282 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_793
timestamp 1612251222
transform -1 0 4314 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_793
timestamp 1612251222
transform -1 0 4148 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_793
timestamp 1612251222
transform -1 0 4132 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_793
timestamp 1612251222
transform -1 0 4116 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_793
timestamp 1612251222
transform -1 0 4100 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_129
timestamp 1612251222
transform 1 0 4100 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_129
timestamp 1612251222
transform 1 0 4084 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_129
timestamp 1612251222
transform 1 0 4068 0 1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_129
timestamp 1612251222
transform 1 0 4052 0 1 3410
box -4 -6 20 206
use POR2X1  POR2X1_172
timestamp 1612251222
transform -1 0 4084 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_172
timestamp 1612251222
transform -1 0 3918 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_172
timestamp 1612251222
transform -1 0 3902 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_172
timestamp 1612251222
transform -1 0 3886 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_431
timestamp 1612251222
transform -1 0 4052 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_431
timestamp 1612251222
transform -1 0 3886 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_431
timestamp 1612251222
transform -1 0 3870 0 1 3410
box -4 -6 20 206
use POR2X1  POR2X1_530
timestamp 1612251222
transform 1 0 3704 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_530
timestamp 1612251222
transform 1 0 3688 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_431
timestamp 1612251222
transform -1 0 3854 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_530
timestamp 1612251222
transform 1 0 3672 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_530
timestamp 1612251222
transform 1 0 3656 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_434
timestamp 1612251222
transform -1 0 3838 0 1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_434
timestamp 1612251222
transform -1 0 3672 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_434
timestamp 1612251222
transform -1 0 3656 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_434
timestamp 1612251222
transform -1 0 3640 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_434
timestamp 1612251222
transform -1 0 3624 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_174
timestamp 1612251222
transform -1 0 3656 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_174
timestamp 1612251222
transform -1 0 3490 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_174
timestamp 1612251222
transform -1 0 3474 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_174
timestamp 1612251222
transform -1 0 3458 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_174
timestamp 1612251222
transform -1 0 3442 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_677
timestamp 1612251222
transform -1 0 3608 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_677
timestamp 1612251222
transform -1 0 3442 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_677
timestamp 1612251222
transform -1 0 3426 0 1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_677
timestamp 1612251222
transform -1 0 3410 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_244
timestamp 1612251222
transform -1 0 3426 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_244
timestamp 1612251222
transform -1 0 3260 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_244
timestamp 1612251222
transform -1 0 3244 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_244
timestamp 1612251222
transform -1 0 3228 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_244
timestamp 1612251222
transform -1 0 3212 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_316
timestamp 1612251222
transform -1 0 3394 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_316
timestamp 1612251222
transform -1 0 3228 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_316
timestamp 1612251222
transform -1 0 3212 0 1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_316
timestamp 1612251222
transform -1 0 3196 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_861
timestamp 1612251222
transform -1 0 3196 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_861
timestamp 1612251222
transform -1 0 3030 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_861
timestamp 1612251222
transform -1 0 3014 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_861
timestamp 1612251222
transform -1 0 2998 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_436
timestamp 1612251222
transform -1 0 3180 0 1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_436
timestamp 1612251222
transform -1 0 3014 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_436
timestamp 1612251222
transform -1 0 2998 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_861
timestamp 1612251222
transform -1 0 2982 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_865
timestamp 1612251222
transform -1 0 2966 0 -1 3810
box -4 -6 170 206
use FILL  FILL0_PAND2X1_436
timestamp 1612251222
transform -1 0 2982 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_436
timestamp 1612251222
transform -1 0 2966 0 1 3410
box -4 -6 20 206
use FILL  FILL2_PAND2X1_865
timestamp 1612251222
transform -1 0 2800 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_865
timestamp 1612251222
transform -1 0 2784 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_865
timestamp 1612251222
transform -1 0 2768 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_865
timestamp 1612251222
transform -1 0 2752 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_851
timestamp 1612251222
transform -1 0 2950 0 1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_851
timestamp 1612251222
transform -1 0 2784 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_851
timestamp 1612251222
transform -1 0 2768 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_851
timestamp 1612251222
transform -1 0 2752 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_851
timestamp 1612251222
transform -1 0 2736 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_858
timestamp 1612251222
transform -1 0 2720 0 1 3410
box -4 -6 170 206
use PAND2X1  PAND2X1_862
timestamp 1612251222
transform 1 0 2570 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_862
timestamp 1612251222
transform 1 0 2554 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_858
timestamp 1612251222
transform -1 0 2506 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_858
timestamp 1612251222
transform -1 0 2522 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_858
timestamp 1612251222
transform -1 0 2538 0 1 3410
box -4 -6 20 206
use FILL  FILL2_PAND2X1_858
timestamp 1612251222
transform -1 0 2554 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_862
timestamp 1612251222
transform 1 0 2506 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_862
timestamp 1612251222
transform 1 0 2522 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_862
timestamp 1612251222
transform 1 0 2538 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_795
timestamp 1612251222
transform -1 0 2506 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_795
timestamp 1612251222
transform -1 0 2340 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_795
timestamp 1612251222
transform -1 0 2324 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_795
timestamp 1612251222
transform -1 0 2308 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_275
timestamp 1612251222
transform -1 0 2490 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_275
timestamp 1612251222
transform -1 0 2324 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_275
timestamp 1612251222
transform -1 0 2308 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_795
timestamp 1612251222
transform -1 0 2292 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_678
timestamp 1612251222
transform -1 0 2276 0 -1 3810
box -4 -6 170 206
use FILL  FILL_POR2X1_275
timestamp 1612251222
transform -1 0 2292 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_276
timestamp 1612251222
transform -1 0 2276 0 1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_678
timestamp 1612251222
transform -1 0 2110 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_678
timestamp 1612251222
transform -1 0 2094 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_678
timestamp 1612251222
transform -1 0 2078 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_678
timestamp 1612251222
transform -1 0 2062 0 -1 3810
box -4 -6 20 206
use FILL  FILL2_PAND2X1_276
timestamp 1612251222
transform -1 0 2110 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_276
timestamp 1612251222
transform -1 0 2094 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_276
timestamp 1612251222
transform -1 0 2078 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_276
timestamp 1612251222
transform -1 0 2062 0 1 3410
box -4 -6 20 206
use POR2X1  POR2X1_173
timestamp 1612251222
transform -1 0 2046 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_173
timestamp 1612251222
transform -1 0 1880 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_173
timestamp 1612251222
transform -1 0 1864 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_173
timestamp 1612251222
transform -1 0 1848 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_589
timestamp 1612251222
transform -1 0 2046 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_589
timestamp 1612251222
transform -1 0 1880 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_589
timestamp 1612251222
transform -1 0 1864 0 1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_589
timestamp 1612251222
transform -1 0 1848 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_592
timestamp 1612251222
transform -1 0 1832 0 1 3410
box -4 -6 170 206
use PAND2X1  PAND2X1_175
timestamp 1612251222
transform -1 0 1832 0 -1 3810
box -4 -6 170 206
use FILL  FILL_PAND2X1_592
timestamp 1612251222
transform -1 0 1618 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_592
timestamp 1612251222
transform -1 0 1634 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_592
timestamp 1612251222
transform -1 0 1650 0 1 3410
box -4 -6 20 206
use FILL  FILL2_PAND2X1_592
timestamp 1612251222
transform -1 0 1666 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_175
timestamp 1612251222
transform -1 0 1618 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_175
timestamp 1612251222
transform -1 0 1634 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_175
timestamp 1612251222
transform -1 0 1650 0 -1 3810
box -4 -6 20 206
use FILL  FILL2_PAND2X1_175
timestamp 1612251222
transform -1 0 1666 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_804
timestamp 1612251222
transform -1 0 1602 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_804
timestamp 1612251222
transform -1 0 1436 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_804
timestamp 1612251222
transform -1 0 1420 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_850
timestamp 1612251222
transform 1 0 1436 0 1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_850
timestamp 1612251222
transform 1 0 1420 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_850
timestamp 1612251222
transform 1 0 1404 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_804
timestamp 1612251222
transform -1 0 1404 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_804
timestamp 1612251222
transform -1 0 1388 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_850
timestamp 1612251222
transform 1 0 1388 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_850
timestamp 1612251222
transform 1 0 1372 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_360
timestamp 1612251222
transform -1 0 1372 0 1 3410
box -4 -6 170 206
use PAND2X1  PAND2X1_808
timestamp 1612251222
transform -1 0 1372 0 -1 3810
box -4 -6 170 206
use FILL  FILL0_PAND2X1_360
timestamp 1612251222
transform -1 0 1174 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_360
timestamp 1612251222
transform -1 0 1190 0 1 3410
box -4 -6 20 206
use FILL  FILL2_PAND2X1_360
timestamp 1612251222
transform -1 0 1206 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_808
timestamp 1612251222
transform -1 0 1174 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_808
timestamp 1612251222
transform -1 0 1190 0 -1 3810
box -4 -6 20 206
use FILL  FILL2_PAND2X1_808
timestamp 1612251222
transform -1 0 1206 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_360
timestamp 1612251222
transform -1 0 1158 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_808
timestamp 1612251222
transform -1 0 1158 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_488
timestamp 1612251222
transform -1 0 1142 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_POR2X1_488
timestamp 1612251222
transform -1 0 976 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_POR2X1_488
timestamp 1612251222
transform -1 0 960 0 -1 3810
box -4 -6 20 206
use FILL  FILL_POR2X1_488
timestamp 1612251222
transform -1 0 944 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_343
timestamp 1612251222
transform -1 0 1142 0 1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_343
timestamp 1612251222
transform -1 0 976 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_343
timestamp 1612251222
transform -1 0 960 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_343
timestamp 1612251222
transform -1 0 944 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_343
timestamp 1612251222
transform -1 0 928 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_363
timestamp 1612251222
transform -1 0 928 0 -1 3810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_363
timestamp 1612251222
transform -1 0 762 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_363
timestamp 1612251222
transform -1 0 746 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_363
timestamp 1612251222
transform -1 0 730 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_296
timestamp 1612251222
transform -1 0 912 0 1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_296
timestamp 1612251222
transform -1 0 746 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_296
timestamp 1612251222
transform -1 0 730 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_363
timestamp 1612251222
transform -1 0 714 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_772
timestamp 1612251222
transform -1 0 698 0 -1 3810
box -4 -6 170 206
use FILL  FILL0_PAND2X1_296
timestamp 1612251222
transform -1 0 714 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_296
timestamp 1612251222
transform -1 0 698 0 1 3410
box -4 -6 20 206
use FILL  FILL2_PAND2X1_772
timestamp 1612251222
transform -1 0 532 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_772
timestamp 1612251222
transform -1 0 516 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_772
timestamp 1612251222
transform -1 0 500 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_772
timestamp 1612251222
transform -1 0 484 0 -1 3810
box -4 -6 20 206
use POR2X1  POR2X1_297
timestamp 1612251222
transform -1 0 682 0 1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_297
timestamp 1612251222
transform -1 0 516 0 1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_297
timestamp 1612251222
transform -1 0 500 0 1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_297
timestamp 1612251222
transform -1 0 484 0 1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_568
timestamp 1612251222
transform -1 0 468 0 1 3410
box -4 -6 170 206
use PAND2X1  PAND2X1_773
timestamp 1612251222
transform -1 0 468 0 -1 3810
box -4 -6 170 206
use FILL  FILL1_PAND2X1_568
timestamp 1612251222
transform -1 0 286 0 1 3410
box -4 -6 20 206
use FILL  FILL2_PAND2X1_568
timestamp 1612251222
transform -1 0 302 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_773
timestamp 1612251222
transform -1 0 286 0 -1 3810
box -4 -6 20 206
use FILL  FILL2_PAND2X1_773
timestamp 1612251222
transform -1 0 302 0 -1 3810
box -4 -6 20 206
use FILL  FILL_PAND2X1_568
timestamp 1612251222
transform -1 0 254 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_568
timestamp 1612251222
transform -1 0 270 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_773
timestamp 1612251222
transform -1 0 254 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_773
timestamp 1612251222
transform -1 0 270 0 -1 3810
box -4 -6 20 206
use PAND2X1  PAND2X1_578
timestamp 1612251222
transform -1 0 238 0 1 3410
box -4 -6 170 206
use PAND2X1  PAND2X1_580
timestamp 1612251222
transform -1 0 238 0 -1 3810
box -4 -6 170 206
use FILL  FILL_PAND2X1_578
timestamp 1612251222
transform -1 0 24 0 1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_578
timestamp 1612251222
transform -1 0 40 0 1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_578
timestamp 1612251222
transform -1 0 56 0 1 3410
box -4 -6 20 206
use FILL  FILL2_PAND2X1_578
timestamp 1612251222
transform -1 0 72 0 1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_580
timestamp 1612251222
transform -1 0 24 0 -1 3810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_580
timestamp 1612251222
transform -1 0 40 0 -1 3810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_580
timestamp 1612251222
transform -1 0 56 0 -1 3810
box -4 -6 20 206
use FILL  FILL2_PAND2X1_580
timestamp 1612251222
transform -1 0 72 0 -1 3810
box -4 -6 20 206
use FILL  FILL_17_12
timestamp 1612251222
transform -1 0 10262 0 -1 3410
box -4 -6 20 206
use FILL  FILL_17_11
timestamp 1612251222
transform -1 0 10246 0 -1 3410
box -4 -6 20 206
use FILL  FILL_17_10
timestamp 1612251222
transform -1 0 10230 0 -1 3410
box -4 -6 20 206
use FILL  FILL_17_9
timestamp 1612251222
transform -1 0 10214 0 -1 3410
box -4 -6 20 206
use FILL  FILL_17_8
timestamp 1612251222
transform -1 0 10198 0 -1 3410
box -4 -6 20 206
use FILL  FILL_17_7
timestamp 1612251222
transform -1 0 10182 0 -1 3410
box -4 -6 20 206
use FILL  FILL_17_6
timestamp 1612251222
transform -1 0 10166 0 -1 3410
box -4 -6 20 206
use FILL  FILL_17_5
timestamp 1612251222
transform -1 0 10150 0 -1 3410
box -4 -6 20 206
use FILL  FILL_17_4
timestamp 1612251222
transform -1 0 10134 0 -1 3410
box -4 -6 20 206
use FILL  FILL_17_3
timestamp 1612251222
transform -1 0 10118 0 -1 3410
box -4 -6 20 206
use FILL  FILL_17_2
timestamp 1612251222
transform -1 0 10102 0 -1 3410
box -4 -6 20 206
use FILL  FILL_17_1
timestamp 1612251222
transform -1 0 10086 0 -1 3410
box -4 -6 20 206
use POR2X1  POR2X1_545
timestamp 1612251222
transform 1 0 9904 0 -1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_545
timestamp 1612251222
transform 1 0 9888 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_545
timestamp 1612251222
transform 1 0 9872 0 -1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_545
timestamp 1612251222
transform 1 0 9856 0 -1 3410
box -4 -6 20 206
use POR2X1  POR2X1_551
timestamp 1612251222
transform -1 0 9856 0 -1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_551
timestamp 1612251222
transform -1 0 9690 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_551
timestamp 1612251222
transform -1 0 9674 0 -1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_551
timestamp 1612251222
transform -1 0 9658 0 -1 3410
box -4 -6 20 206
use POR2X1  POR2X1_564
timestamp 1612251222
transform 1 0 9476 0 -1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_564
timestamp 1612251222
transform 1 0 9460 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_564
timestamp 1612251222
transform 1 0 9444 0 -1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_564
timestamp 1612251222
transform 1 0 9428 0 -1 3410
box -4 -6 20 206
use POR2X1  POR2X1_552
timestamp 1612251222
transform 1 0 9262 0 -1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_552
timestamp 1612251222
transform 1 0 9246 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_552
timestamp 1612251222
transform 1 0 9230 0 -1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_552
timestamp 1612251222
transform 1 0 9214 0 -1 3410
box -4 -6 20 206
use POR2X1  POR2X1_542
timestamp 1612251222
transform 1 0 9048 0 -1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_542
timestamp 1612251222
transform 1 0 9032 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_542
timestamp 1612251222
transform 1 0 9016 0 -1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_542
timestamp 1612251222
transform 1 0 9000 0 -1 3410
box -4 -6 20 206
use POR2X1  POR2X1_464
timestamp 1612251222
transform 1 0 8834 0 -1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_464
timestamp 1612251222
transform 1 0 8818 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_464
timestamp 1612251222
transform 1 0 8802 0 -1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_464
timestamp 1612251222
transform 1 0 8786 0 -1 3410
box -4 -6 20 206
use POR2X1  POR2X1_457
timestamp 1612251222
transform 1 0 8620 0 -1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_457
timestamp 1612251222
transform 1 0 8604 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_457
timestamp 1612251222
transform 1 0 8588 0 -1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_457
timestamp 1612251222
transform 1 0 8572 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_368
timestamp 1612251222
transform 1 0 8406 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_368
timestamp 1612251222
transform 1 0 8390 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_368
timestamp 1612251222
transform 1 0 8374 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_368
timestamp 1612251222
transform 1 0 8358 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_368
timestamp 1612251222
transform 1 0 8342 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_369
timestamp 1612251222
transform 1 0 8176 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_369
timestamp 1612251222
transform 1 0 8160 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_369
timestamp 1612251222
transform 1 0 8144 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_369
timestamp 1612251222
transform 1 0 8128 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_369
timestamp 1612251222
transform 1 0 8112 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_300
timestamp 1612251222
transform 1 0 7946 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_300
timestamp 1612251222
transform 1 0 7930 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_300
timestamp 1612251222
transform 1 0 7914 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_300
timestamp 1612251222
transform 1 0 7898 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_300
timestamp 1612251222
transform 1 0 7882 0 -1 3410
box -4 -6 20 206
use POR2X1  POR2X1_843
timestamp 1612251222
transform 1 0 7716 0 -1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_843
timestamp 1612251222
transform 1 0 7700 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_843
timestamp 1612251222
transform 1 0 7684 0 -1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_843
timestamp 1612251222
transform 1 0 7668 0 -1 3410
box -4 -6 20 206
use POR2X1  POR2X1_343
timestamp 1612251222
transform -1 0 7668 0 -1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_343
timestamp 1612251222
transform -1 0 7502 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_343
timestamp 1612251222
transform -1 0 7486 0 -1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_343
timestamp 1612251222
transform -1 0 7470 0 -1 3410
box -4 -6 20 206
use POR2X1  POR2X1_458
timestamp 1612251222
transform 1 0 7288 0 -1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_458
timestamp 1612251222
transform 1 0 7272 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_458
timestamp 1612251222
transform 1 0 7256 0 -1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_458
timestamp 1612251222
transform 1 0 7240 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_250
timestamp 1612251222
transform 1 0 7074 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_250
timestamp 1612251222
transform 1 0 7058 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_250
timestamp 1612251222
transform 1 0 7042 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_250
timestamp 1612251222
transform 1 0 7026 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_250
timestamp 1612251222
transform 1 0 7010 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_371
timestamp 1612251222
transform 1 0 6844 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_371
timestamp 1612251222
transform 1 0 6828 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_371
timestamp 1612251222
transform 1 0 6812 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_371
timestamp 1612251222
transform 1 0 6796 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_371
timestamp 1612251222
transform 1 0 6780 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_122
timestamp 1612251222
transform 1 0 6614 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_122
timestamp 1612251222
transform 1 0 6598 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_122
timestamp 1612251222
transform 1 0 6582 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_122
timestamp 1612251222
transform 1 0 6566 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_122
timestamp 1612251222
transform 1 0 6550 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_487
timestamp 1612251222
transform -1 0 6550 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_487
timestamp 1612251222
transform -1 0 6384 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_487
timestamp 1612251222
transform -1 0 6368 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_487
timestamp 1612251222
transform -1 0 6352 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_487
timestamp 1612251222
transform -1 0 6336 0 -1 3410
box -4 -6 20 206
use POR2X1  POR2X1_486
timestamp 1612251222
transform -1 0 6320 0 -1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_486
timestamp 1612251222
transform -1 0 6154 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_486
timestamp 1612251222
transform -1 0 6138 0 -1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_486
timestamp 1612251222
transform -1 0 6122 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_484
timestamp 1612251222
transform 1 0 5940 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_484
timestamp 1612251222
transform 1 0 5924 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_484
timestamp 1612251222
transform 1 0 5908 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_484
timestamp 1612251222
transform 1 0 5892 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_484
timestamp 1612251222
transform 1 0 5876 0 -1 3410
box -4 -6 20 206
use POR2X1  POR2X1_705
timestamp 1612251222
transform 1 0 5710 0 -1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_705
timestamp 1612251222
transform 1 0 5694 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_705
timestamp 1612251222
transform 1 0 5678 0 -1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_705
timestamp 1612251222
transform 1 0 5662 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_485
timestamp 1612251222
transform 1 0 5496 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_485
timestamp 1612251222
transform 1 0 5480 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_485
timestamp 1612251222
transform 1 0 5464 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_485
timestamp 1612251222
transform 1 0 5448 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_485
timestamp 1612251222
transform 1 0 5432 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_416
timestamp 1612251222
transform 1 0 5266 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_416
timestamp 1612251222
transform 1 0 5250 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_416
timestamp 1612251222
transform 1 0 5234 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_416
timestamp 1612251222
transform 1 0 5218 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_416
timestamp 1612251222
transform 1 0 5202 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_819
timestamp 1612251222
transform -1 0 5202 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_819
timestamp 1612251222
transform -1 0 5036 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_819
timestamp 1612251222
transform -1 0 5020 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_819
timestamp 1612251222
transform -1 0 5004 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_819
timestamp 1612251222
transform -1 0 4988 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_820
timestamp 1612251222
transform -1 0 4972 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_820
timestamp 1612251222
transform -1 0 4806 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_820
timestamp 1612251222
transform -1 0 4790 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_820
timestamp 1612251222
transform -1 0 4774 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_820
timestamp 1612251222
transform -1 0 4758 0 -1 3410
box -4 -6 20 206
use POR2X1  POR2X1_847
timestamp 1612251222
transform -1 0 4742 0 -1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_847
timestamp 1612251222
transform -1 0 4576 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_847
timestamp 1612251222
transform -1 0 4560 0 -1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_847
timestamp 1612251222
transform -1 0 4544 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_790
timestamp 1612251222
transform -1 0 4528 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_790
timestamp 1612251222
transform -1 0 4362 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_790
timestamp 1612251222
transform -1 0 4346 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_790
timestamp 1612251222
transform -1 0 4330 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_790
timestamp 1612251222
transform -1 0 4314 0 -1 3410
box -4 -6 20 206
use POR2X1  POR2X1_616
timestamp 1612251222
transform 1 0 4132 0 -1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_616
timestamp 1612251222
transform 1 0 4116 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_616
timestamp 1612251222
transform 1 0 4100 0 -1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_616
timestamp 1612251222
transform 1 0 4084 0 -1 3410
box -4 -6 20 206
use POR2X1  POR2X1_268
timestamp 1612251222
transform -1 0 4084 0 -1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_268
timestamp 1612251222
transform -1 0 3918 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_268
timestamp 1612251222
transform -1 0 3902 0 -1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_268
timestamp 1612251222
transform -1 0 3886 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_269
timestamp 1612251222
transform -1 0 3870 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_269
timestamp 1612251222
transform -1 0 3704 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_269
timestamp 1612251222
transform -1 0 3688 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_269
timestamp 1612251222
transform -1 0 3672 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_269
timestamp 1612251222
transform -1 0 3656 0 -1 3410
box -4 -6 20 206
use POR2X1  POR2X1_432
timestamp 1612251222
transform -1 0 3640 0 -1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_432
timestamp 1612251222
transform -1 0 3474 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_432
timestamp 1612251222
transform -1 0 3458 0 -1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_432
timestamp 1612251222
transform -1 0 3442 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_435
timestamp 1612251222
transform -1 0 3426 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_435
timestamp 1612251222
transform -1 0 3260 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_435
timestamp 1612251222
transform -1 0 3244 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_435
timestamp 1612251222
transform -1 0 3228 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_435
timestamp 1612251222
transform -1 0 3212 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_832
timestamp 1612251222
transform -1 0 3196 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_832
timestamp 1612251222
transform -1 0 3030 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_832
timestamp 1612251222
transform -1 0 3014 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_832
timestamp 1612251222
transform -1 0 2998 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_832
timestamp 1612251222
transform -1 0 2982 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_841
timestamp 1612251222
transform 1 0 2800 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_841
timestamp 1612251222
transform 1 0 2784 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_841
timestamp 1612251222
transform 1 0 2768 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_841
timestamp 1612251222
transform 1 0 2752 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_841
timestamp 1612251222
transform 1 0 2736 0 -1 3410
box -4 -6 20 206
use POR2X1  POR2X1_271
timestamp 1612251222
transform -1 0 2736 0 -1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_271
timestamp 1612251222
transform -1 0 2570 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_271
timestamp 1612251222
transform -1 0 2554 0 -1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_271
timestamp 1612251222
transform -1 0 2538 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_831
timestamp 1612251222
transform 1 0 2356 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_831
timestamp 1612251222
transform 1 0 2340 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_831
timestamp 1612251222
transform 1 0 2324 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_831
timestamp 1612251222
transform 1 0 2308 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_831
timestamp 1612251222
transform 1 0 2292 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_274
timestamp 1612251222
transform 1 0 2126 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_274
timestamp 1612251222
transform 1 0 2110 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_274
timestamp 1612251222
transform 1 0 2094 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_274
timestamp 1612251222
transform 1 0 2078 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_274
timestamp 1612251222
transform 1 0 2062 0 -1 3410
box -4 -6 20 206
use POR2X1  POR2X1_273
timestamp 1612251222
transform 1 0 1896 0 -1 3410
box -4 -6 170 206
use FILL  FILL1_POR2X1_273
timestamp 1612251222
transform 1 0 1880 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_POR2X1_273
timestamp 1612251222
transform 1 0 1864 0 -1 3410
box -4 -6 20 206
use FILL  FILL_POR2X1_273
timestamp 1612251222
transform 1 0 1848 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_390
timestamp 1612251222
transform 1 0 1682 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_390
timestamp 1612251222
transform 1 0 1666 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_390
timestamp 1612251222
transform 1 0 1650 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_390
timestamp 1612251222
transform 1 0 1634 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_390
timestamp 1612251222
transform 1 0 1618 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_842
timestamp 1612251222
transform -1 0 1618 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_842
timestamp 1612251222
transform -1 0 1452 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_842
timestamp 1612251222
transform -1 0 1436 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_842
timestamp 1612251222
transform -1 0 1420 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_842
timestamp 1612251222
transform -1 0 1404 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_389
timestamp 1612251222
transform 1 0 1222 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_389
timestamp 1612251222
transform 1 0 1206 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_389
timestamp 1612251222
transform 1 0 1190 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_389
timestamp 1612251222
transform 1 0 1174 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_389
timestamp 1612251222
transform 1 0 1158 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_843
timestamp 1612251222
transform 1 0 992 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_843
timestamp 1612251222
transform 1 0 976 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_843
timestamp 1612251222
transform 1 0 960 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_843
timestamp 1612251222
transform 1 0 944 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_843
timestamp 1612251222
transform 1 0 928 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_349
timestamp 1612251222
transform -1 0 928 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_349
timestamp 1612251222
transform -1 0 762 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_349
timestamp 1612251222
transform -1 0 746 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_349
timestamp 1612251222
transform -1 0 730 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_349
timestamp 1612251222
transform -1 0 714 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_359
timestamp 1612251222
transform -1 0 698 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_359
timestamp 1612251222
transform -1 0 532 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_359
timestamp 1612251222
transform -1 0 516 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_359
timestamp 1612251222
transform -1 0 500 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_359
timestamp 1612251222
transform -1 0 484 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_347
timestamp 1612251222
transform -1 0 468 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_347
timestamp 1612251222
transform -1 0 302 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_347
timestamp 1612251222
transform -1 0 286 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_347
timestamp 1612251222
transform -1 0 270 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_347
timestamp 1612251222
transform -1 0 254 0 -1 3410
box -4 -6 20 206
use PAND2X1  PAND2X1_287
timestamp 1612251222
transform -1 0 238 0 -1 3410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_287
timestamp 1612251222
transform -1 0 72 0 -1 3410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_287
timestamp 1612251222
transform -1 0 56 0 -1 3410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_287
timestamp 1612251222
transform -1 0 40 0 -1 3410
box -4 -6 20 206
use FILL  FILL_PAND2X1_287
timestamp 1612251222
transform -1 0 24 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_13
timestamp 1612251222
transform 1 0 10252 0 1 3010
box -4 -6 20 206
use FILL  FILL_16_12
timestamp 1612251222
transform 1 0 10236 0 1 3010
box -4 -6 20 206
use FILL  FILL_16_11
timestamp 1612251222
transform 1 0 10220 0 1 3010
box -4 -6 20 206
use FILL  FILL_16_10
timestamp 1612251222
transform 1 0 10204 0 1 3010
box -4 -6 20 206
use FILL  FILL_16_9
timestamp 1612251222
transform 1 0 10188 0 1 3010
box -4 -6 20 206
use FILL  FILL_16_8
timestamp 1612251222
transform 1 0 10172 0 1 3010
box -4 -6 20 206
use FILL  FILL_16_7
timestamp 1612251222
transform 1 0 10156 0 1 3010
box -4 -6 20 206
use FILL  FILL_16_6
timestamp 1612251222
transform 1 0 10140 0 1 3010
box -4 -6 20 206
use FILL  FILL_16_5
timestamp 1612251222
transform 1 0 10124 0 1 3010
box -4 -6 20 206
use FILL  FILL_16_4
timestamp 1612251222
transform 1 0 10108 0 1 3010
box -4 -6 20 206
use FILL  FILL_16_3
timestamp 1612251222
transform 1 0 10092 0 1 3010
box -4 -6 20 206
use FILL  FILL_16_2
timestamp 1612251222
transform 1 0 10076 0 1 3010
box -4 -6 20 206
use FILL  FILL_16_1
timestamp 1612251222
transform 1 0 10060 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_444
timestamp 1612251222
transform -1 0 10060 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_444
timestamp 1612251222
transform -1 0 9894 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_444
timestamp 1612251222
transform -1 0 9878 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_444
timestamp 1612251222
transform -1 0 9862 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_544
timestamp 1612251222
transform 1 0 9680 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_544
timestamp 1612251222
transform 1 0 9664 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_544
timestamp 1612251222
transform 1 0 9648 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_544
timestamp 1612251222
transform 1 0 9632 0 1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_438
timestamp 1612251222
transform 1 0 9466 0 1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_438
timestamp 1612251222
transform 1 0 9450 0 1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_438
timestamp 1612251222
transform 1 0 9434 0 1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_438
timestamp 1612251222
transform 1 0 9418 0 1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_438
timestamp 1612251222
transform 1 0 9402 0 1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_373
timestamp 1612251222
transform 1 0 9236 0 1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_373
timestamp 1612251222
transform 1 0 9220 0 1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_373
timestamp 1612251222
transform 1 0 9204 0 1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_373
timestamp 1612251222
transform 1 0 9188 0 1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_373
timestamp 1612251222
transform 1 0 9172 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_663
timestamp 1612251222
transform 1 0 9006 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_663
timestamp 1612251222
transform 1 0 8990 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_663
timestamp 1612251222
transform 1 0 8974 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_663
timestamp 1612251222
transform 1 0 8958 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_325
timestamp 1612251222
transform 1 0 8792 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_325
timestamp 1612251222
transform 1 0 8776 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_325
timestamp 1612251222
transform 1 0 8760 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_325
timestamp 1612251222
transform 1 0 8744 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_374
timestamp 1612251222
transform -1 0 8744 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_374
timestamp 1612251222
transform -1 0 8578 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_374
timestamp 1612251222
transform -1 0 8562 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_374
timestamp 1612251222
transform -1 0 8546 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_787
timestamp 1612251222
transform 1 0 8364 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_787
timestamp 1612251222
transform 1 0 8348 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_787
timestamp 1612251222
transform 1 0 8332 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_787
timestamp 1612251222
transform 1 0 8316 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_284
timestamp 1612251222
transform -1 0 8316 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_284
timestamp 1612251222
transform -1 0 8150 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_284
timestamp 1612251222
transform -1 0 8134 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_284
timestamp 1612251222
transform -1 0 8118 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_249
timestamp 1612251222
transform -1 0 8102 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_249
timestamp 1612251222
transform -1 0 7936 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_249
timestamp 1612251222
transform -1 0 7920 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_249
timestamp 1612251222
transform -1 0 7904 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_287
timestamp 1612251222
transform -1 0 7888 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_287
timestamp 1612251222
transform -1 0 7722 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_287
timestamp 1612251222
transform -1 0 7706 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_287
timestamp 1612251222
transform -1 0 7690 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_734
timestamp 1612251222
transform 1 0 7508 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_734
timestamp 1612251222
transform 1 0 7492 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_734
timestamp 1612251222
transform 1 0 7476 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_734
timestamp 1612251222
transform 1 0 7460 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_475
timestamp 1612251222
transform -1 0 7460 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_475
timestamp 1612251222
transform -1 0 7294 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_475
timestamp 1612251222
transform -1 0 7278 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_475
timestamp 1612251222
transform -1 0 7262 0 1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_611
timestamp 1612251222
transform -1 0 7246 0 1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_611
timestamp 1612251222
transform -1 0 7080 0 1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_611
timestamp 1612251222
transform -1 0 7064 0 1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_611
timestamp 1612251222
transform -1 0 7048 0 1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_611
timestamp 1612251222
transform -1 0 7032 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_773
timestamp 1612251222
transform 1 0 6850 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_773
timestamp 1612251222
transform 1 0 6834 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_773
timestamp 1612251222
transform 1 0 6818 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_773
timestamp 1612251222
transform 1 0 6802 0 1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_283
timestamp 1612251222
transform 1 0 6636 0 1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_283
timestamp 1612251222
transform 1 0 6620 0 1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_283
timestamp 1612251222
transform 1 0 6604 0 1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_283
timestamp 1612251222
transform 1 0 6588 0 1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_283
timestamp 1612251222
transform 1 0 6572 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_642
timestamp 1612251222
transform 1 0 6406 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_642
timestamp 1612251222
transform 1 0 6390 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_642
timestamp 1612251222
transform 1 0 6374 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_642
timestamp 1612251222
transform 1 0 6358 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_462
timestamp 1612251222
transform 1 0 6192 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_462
timestamp 1612251222
transform 1 0 6176 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_462
timestamp 1612251222
transform 1 0 6160 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_462
timestamp 1612251222
transform 1 0 6144 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_859
timestamp 1612251222
transform 1 0 5978 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_859
timestamp 1612251222
transform 1 0 5962 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_859
timestamp 1612251222
transform 1 0 5946 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_859
timestamp 1612251222
transform 1 0 5930 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_848
timestamp 1612251222
transform 1 0 5764 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_848
timestamp 1612251222
transform 1 0 5748 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_848
timestamp 1612251222
transform 1 0 5732 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_848
timestamp 1612251222
transform 1 0 5716 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_790
timestamp 1612251222
transform 1 0 5550 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_790
timestamp 1612251222
transform 1 0 5534 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_790
timestamp 1612251222
transform 1 0 5518 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_790
timestamp 1612251222
transform 1 0 5502 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_753
timestamp 1612251222
transform 1 0 5336 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_753
timestamp 1612251222
transform 1 0 5320 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_753
timestamp 1612251222
transform 1 0 5304 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_753
timestamp 1612251222
transform 1 0 5288 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_754
timestamp 1612251222
transform -1 0 5288 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_754
timestamp 1612251222
transform -1 0 5122 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_754
timestamp 1612251222
transform -1 0 5106 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_754
timestamp 1612251222
transform -1 0 5090 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_615
timestamp 1612251222
transform -1 0 5074 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_615
timestamp 1612251222
transform -1 0 4908 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_615
timestamp 1612251222
transform -1 0 4892 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_615
timestamp 1612251222
transform -1 0 4876 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_90
timestamp 1612251222
transform -1 0 4860 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_90
timestamp 1612251222
transform -1 0 4694 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_90
timestamp 1612251222
transform -1 0 4678 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_90
timestamp 1612251222
transform -1 0 4662 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_625
timestamp 1612251222
transform -1 0 4646 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_625
timestamp 1612251222
transform -1 0 4480 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_625
timestamp 1612251222
transform -1 0 4464 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_625
timestamp 1612251222
transform -1 0 4448 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_245
timestamp 1612251222
transform 1 0 4266 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_245
timestamp 1612251222
transform 1 0 4250 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_245
timestamp 1612251222
transform 1 0 4234 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_245
timestamp 1612251222
transform 1 0 4218 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_246
timestamp 1612251222
transform -1 0 4218 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_246
timestamp 1612251222
transform -1 0 4052 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_246
timestamp 1612251222
transform -1 0 4036 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_246
timestamp 1612251222
transform -1 0 4020 0 1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_342
timestamp 1612251222
transform -1 0 4004 0 1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_342
timestamp 1612251222
transform -1 0 3838 0 1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_342
timestamp 1612251222
transform -1 0 3822 0 1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_342
timestamp 1612251222
transform -1 0 3806 0 1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_342
timestamp 1612251222
transform -1 0 3790 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_433
timestamp 1612251222
transform -1 0 3774 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_433
timestamp 1612251222
transform -1 0 3608 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_433
timestamp 1612251222
transform -1 0 3592 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_433
timestamp 1612251222
transform -1 0 3576 0 1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_834
timestamp 1612251222
transform -1 0 3560 0 1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_834
timestamp 1612251222
transform -1 0 3394 0 1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_834
timestamp 1612251222
transform -1 0 3378 0 1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_834
timestamp 1612251222
transform -1 0 3362 0 1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_834
timestamp 1612251222
transform -1 0 3346 0 1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_840
timestamp 1612251222
transform -1 0 3330 0 1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_840
timestamp 1612251222
transform -1 0 3164 0 1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_840
timestamp 1612251222
transform -1 0 3148 0 1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_840
timestamp 1612251222
transform -1 0 3132 0 1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_840
timestamp 1612251222
transform -1 0 3116 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_255
timestamp 1612251222
transform -1 0 3100 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_255
timestamp 1612251222
transform -1 0 2934 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_255
timestamp 1612251222
transform -1 0 2918 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_255
timestamp 1612251222
transform -1 0 2902 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_75
timestamp 1612251222
transform -1 0 2886 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_75
timestamp 1612251222
transform -1 0 2720 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_75
timestamp 1612251222
transform -1 0 2704 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_75
timestamp 1612251222
transform -1 0 2688 0 1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_301
timestamp 1612251222
transform 1 0 2506 0 1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_301
timestamp 1612251222
transform 1 0 2490 0 1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_301
timestamp 1612251222
transform 1 0 2474 0 1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_301
timestamp 1612251222
transform 1 0 2458 0 1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_301
timestamp 1612251222
transform 1 0 2442 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_300
timestamp 1612251222
transform -1 0 2442 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_300
timestamp 1612251222
transform -1 0 2276 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_300
timestamp 1612251222
transform -1 0 2260 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_300
timestamp 1612251222
transform -1 0 2244 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_272
timestamp 1612251222
transform 1 0 2062 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_272
timestamp 1612251222
transform 1 0 2046 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_272
timestamp 1612251222
transform 1 0 2030 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_272
timestamp 1612251222
transform 1 0 2014 0 1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_141
timestamp 1612251222
transform 1 0 1848 0 1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_141
timestamp 1612251222
transform 1 0 1832 0 1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_141
timestamp 1612251222
transform 1 0 1816 0 1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_141
timestamp 1612251222
transform 1 0 1800 0 1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_141
timestamp 1612251222
transform 1 0 1784 0 1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_139
timestamp 1612251222
transform 1 0 1618 0 1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_139
timestamp 1612251222
transform 1 0 1602 0 1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_139
timestamp 1612251222
transform 1 0 1586 0 1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_139
timestamp 1612251222
transform 1 0 1570 0 1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_139
timestamp 1612251222
transform 1 0 1554 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_131
timestamp 1612251222
transform -1 0 1554 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_131
timestamp 1612251222
transform -1 0 1388 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_131
timestamp 1612251222
transform -1 0 1372 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_131
timestamp 1612251222
transform -1 0 1356 0 1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_140
timestamp 1612251222
transform 1 0 1174 0 1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_140
timestamp 1612251222
transform 1 0 1158 0 1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_140
timestamp 1612251222
transform 1 0 1142 0 1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_140
timestamp 1612251222
transform 1 0 1126 0 1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_140
timestamp 1612251222
transform 1 0 1110 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_103
timestamp 1612251222
transform -1 0 1110 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_103
timestamp 1612251222
transform -1 0 944 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_103
timestamp 1612251222
transform -1 0 928 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_103
timestamp 1612251222
transform -1 0 912 0 1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_768
timestamp 1612251222
transform -1 0 896 0 1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_768
timestamp 1612251222
transform -1 0 730 0 1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_768
timestamp 1612251222
transform -1 0 714 0 1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_768
timestamp 1612251222
transform -1 0 698 0 1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_768
timestamp 1612251222
transform -1 0 682 0 1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_137
timestamp 1612251222
transform 1 0 500 0 1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_137
timestamp 1612251222
transform 1 0 484 0 1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_137
timestamp 1612251222
transform 1 0 468 0 1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_137
timestamp 1612251222
transform 1 0 452 0 1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_137
timestamp 1612251222
transform 1 0 436 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_134
timestamp 1612251222
transform 1 0 270 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_134
timestamp 1612251222
transform 1 0 254 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_134
timestamp 1612251222
transform 1 0 238 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_134
timestamp 1612251222
transform 1 0 222 0 1 3010
box -4 -6 20 206
use POR2X1  POR2X1_125
timestamp 1612251222
transform -1 0 222 0 1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_125
timestamp 1612251222
transform -1 0 56 0 1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_125
timestamp 1612251222
transform -1 0 40 0 1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_125
timestamp 1612251222
transform -1 0 24 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_12
timestamp 1612251222
transform -1 0 10262 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_11
timestamp 1612251222
transform -1 0 10246 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_10
timestamp 1612251222
transform -1 0 10230 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_9
timestamp 1612251222
transform -1 0 10214 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_8
timestamp 1612251222
transform -1 0 10198 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_7
timestamp 1612251222
transform -1 0 10182 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_6
timestamp 1612251222
transform -1 0 10166 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_5
timestamp 1612251222
transform -1 0 10150 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_4
timestamp 1612251222
transform -1 0 10134 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_3
timestamp 1612251222
transform -1 0 10118 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_2
timestamp 1612251222
transform -1 0 10102 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_1
timestamp 1612251222
transform -1 0 10086 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_442
timestamp 1612251222
transform 1 0 9904 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_442
timestamp 1612251222
transform 1 0 9888 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_442
timestamp 1612251222
transform 1 0 9872 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_442
timestamp 1612251222
transform 1 0 9856 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_442
timestamp 1612251222
transform 1 0 9840 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_177
timestamp 1612251222
transform 1 0 9674 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_177
timestamp 1612251222
transform 1 0 9658 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_177
timestamp 1612251222
transform 1 0 9642 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_177
timestamp 1612251222
transform 1 0 9626 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_177
timestamp 1612251222
transform 1 0 9610 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_439
timestamp 1612251222
transform -1 0 9610 0 -1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_439
timestamp 1612251222
transform -1 0 9444 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_439
timestamp 1612251222
transform -1 0 9428 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_439
timestamp 1612251222
transform -1 0 9412 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_183
timestamp 1612251222
transform -1 0 9396 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_183
timestamp 1612251222
transform -1 0 9230 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_183
timestamp 1612251222
transform -1 0 9214 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_183
timestamp 1612251222
transform -1 0 9198 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_183
timestamp 1612251222
transform -1 0 9182 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_280
timestamp 1612251222
transform -1 0 9166 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_280
timestamp 1612251222
transform -1 0 9000 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_280
timestamp 1612251222
transform -1 0 8984 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_280
timestamp 1612251222
transform -1 0 8968 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_280
timestamp 1612251222
transform -1 0 8952 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_298
timestamp 1612251222
transform -1 0 8936 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_298
timestamp 1612251222
transform -1 0 8770 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_298
timestamp 1612251222
transform -1 0 8754 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_298
timestamp 1612251222
transform -1 0 8738 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_298
timestamp 1612251222
transform -1 0 8722 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_322
timestamp 1612251222
transform 1 0 8540 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_322
timestamp 1612251222
transform 1 0 8524 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_322
timestamp 1612251222
transform 1 0 8508 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_322
timestamp 1612251222
transform 1 0 8492 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_322
timestamp 1612251222
transform 1 0 8476 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_279
timestamp 1612251222
transform 1 0 8310 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_279
timestamp 1612251222
transform 1 0 8294 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_279
timestamp 1612251222
transform 1 0 8278 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_279
timestamp 1612251222
transform 1 0 8262 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_279
timestamp 1612251222
transform 1 0 8246 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_302
timestamp 1612251222
transform 1 0 8080 0 -1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_302
timestamp 1612251222
transform 1 0 8064 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_302
timestamp 1612251222
transform 1 0 8048 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_302
timestamp 1612251222
transform 1 0 8032 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_299
timestamp 1612251222
transform -1 0 8032 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_299
timestamp 1612251222
transform -1 0 7866 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_299
timestamp 1612251222
transform -1 0 7850 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_299
timestamp 1612251222
transform -1 0 7834 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_299
timestamp 1612251222
transform -1 0 7818 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_405
timestamp 1612251222
transform 1 0 7636 0 -1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_405
timestamp 1612251222
transform 1 0 7620 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_405
timestamp 1612251222
transform 1 0 7604 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_405
timestamp 1612251222
transform 1 0 7588 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_406
timestamp 1612251222
transform -1 0 7588 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_406
timestamp 1612251222
transform -1 0 7422 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_406
timestamp 1612251222
transform -1 0 7406 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_406
timestamp 1612251222
transform -1 0 7390 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_406
timestamp 1612251222
transform -1 0 7374 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_288
timestamp 1612251222
transform 1 0 7192 0 -1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_288
timestamp 1612251222
transform 1 0 7176 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_288
timestamp 1612251222
transform 1 0 7160 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_288
timestamp 1612251222
transform 1 0 7144 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_479
timestamp 1612251222
transform 1 0 6978 0 -1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_479
timestamp 1612251222
transform 1 0 6962 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_479
timestamp 1612251222
transform 1 0 6946 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_479
timestamp 1612251222
transform 1 0 6930 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_595
timestamp 1612251222
transform -1 0 6930 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_595
timestamp 1612251222
transform -1 0 6764 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_595
timestamp 1612251222
transform -1 0 6748 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_595
timestamp 1612251222
transform -1 0 6732 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_595
timestamp 1612251222
transform -1 0 6716 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_476
timestamp 1612251222
transform 1 0 6534 0 -1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_476
timestamp 1612251222
transform 1 0 6518 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_476
timestamp 1612251222
transform 1 0 6502 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_476
timestamp 1612251222
transform 1 0 6486 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_612
timestamp 1612251222
transform 1 0 6320 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_612
timestamp 1612251222
transform 1 0 6304 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_612
timestamp 1612251222
transform 1 0 6288 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_612
timestamp 1612251222
transform 1 0 6272 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_612
timestamp 1612251222
transform 1 0 6256 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_610
timestamp 1612251222
transform -1 0 6256 0 -1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_610
timestamp 1612251222
transform -1 0 6090 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_610
timestamp 1612251222
transform -1 0 6074 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_610
timestamp 1612251222
transform -1 0 6058 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_413
timestamp 1612251222
transform -1 0 6042 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_413
timestamp 1612251222
transform -1 0 5876 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_413
timestamp 1612251222
transform -1 0 5860 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_413
timestamp 1612251222
transform -1 0 5844 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_413
timestamp 1612251222
transform -1 0 5828 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_461
timestamp 1612251222
transform -1 0 5812 0 -1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_461
timestamp 1612251222
transform -1 0 5646 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_461
timestamp 1612251222
transform -1 0 5630 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_461
timestamp 1612251222
transform -1 0 5614 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_814
timestamp 1612251222
transform -1 0 5598 0 -1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_814
timestamp 1612251222
transform -1 0 5432 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_814
timestamp 1612251222
transform -1 0 5416 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_814
timestamp 1612251222
transform -1 0 5400 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_815
timestamp 1612251222
transform -1 0 5384 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_815
timestamp 1612251222
transform -1 0 5218 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_815
timestamp 1612251222
transform -1 0 5202 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_815
timestamp 1612251222
transform -1 0 5186 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_815
timestamp 1612251222
transform -1 0 5170 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_846
timestamp 1612251222
transform -1 0 5154 0 -1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_846
timestamp 1612251222
transform -1 0 4988 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_846
timestamp 1612251222
transform -1 0 4972 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_846
timestamp 1612251222
transform -1 0 4956 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_623
timestamp 1612251222
transform -1 0 4940 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_623
timestamp 1612251222
transform -1 0 4774 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_623
timestamp 1612251222
transform -1 0 4758 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_623
timestamp 1612251222
transform -1 0 4742 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_623
timestamp 1612251222
transform -1 0 4726 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_225
timestamp 1612251222
transform 1 0 4544 0 -1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_225
timestamp 1612251222
transform 1 0 4528 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_225
timestamp 1612251222
transform 1 0 4512 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_225
timestamp 1612251222
transform 1 0 4496 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_614
timestamp 1612251222
transform 1 0 4330 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_614
timestamp 1612251222
transform 1 0 4314 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_614
timestamp 1612251222
transform 1 0 4298 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_614
timestamp 1612251222
transform 1 0 4282 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_614
timestamp 1612251222
transform 1 0 4266 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_247
timestamp 1612251222
transform -1 0 4266 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_247
timestamp 1612251222
transform -1 0 4100 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_247
timestamp 1612251222
transform -1 0 4084 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_247
timestamp 1612251222
transform -1 0 4068 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_247
timestamp 1612251222
transform -1 0 4052 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_248
timestamp 1612251222
transform -1 0 4036 0 -1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_248
timestamp 1612251222
transform -1 0 3870 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_248
timestamp 1612251222
transform -1 0 3854 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_248
timestamp 1612251222
transform -1 0 3838 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_495
timestamp 1612251222
transform -1 0 3822 0 -1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_495
timestamp 1612251222
transform -1 0 3656 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_495
timestamp 1612251222
transform -1 0 3640 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_495
timestamp 1612251222
transform -1 0 3624 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_833
timestamp 1612251222
transform -1 0 3608 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_833
timestamp 1612251222
transform -1 0 3442 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_833
timestamp 1612251222
transform -1 0 3426 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_833
timestamp 1612251222
transform -1 0 3410 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_833
timestamp 1612251222
transform -1 0 3394 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_499
timestamp 1612251222
transform -1 0 3378 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_499
timestamp 1612251222
transform -1 0 3212 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_499
timestamp 1612251222
transform -1 0 3196 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_499
timestamp 1612251222
transform -1 0 3180 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_499
timestamp 1612251222
transform -1 0 3164 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_270
timestamp 1612251222
transform -1 0 3148 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_270
timestamp 1612251222
transform -1 0 2982 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_270
timestamp 1612251222
transform -1 0 2966 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_270
timestamp 1612251222
transform -1 0 2950 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_270
timestamp 1612251222
transform -1 0 2934 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_74
timestamp 1612251222
transform -1 0 2918 0 -1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_74
timestamp 1612251222
transform -1 0 2752 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_74
timestamp 1612251222
transform -1 0 2736 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_74
timestamp 1612251222
transform -1 0 2720 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_76
timestamp 1612251222
transform -1 0 2704 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_76
timestamp 1612251222
transform -1 0 2538 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_76
timestamp 1612251222
transform -1 0 2522 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_76
timestamp 1612251222
transform -1 0 2506 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_76
timestamp 1612251222
transform -1 0 2490 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_332
timestamp 1612251222
transform 1 0 2308 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_332
timestamp 1612251222
transform 1 0 2292 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_332
timestamp 1612251222
transform 1 0 2276 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_332
timestamp 1612251222
transform 1 0 2260 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_332
timestamp 1612251222
transform 1 0 2244 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_45
timestamp 1612251222
transform 1 0 2078 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_POR2X1_45
timestamp 1612251222
transform 1 0 2062 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_POR2X1_45
timestamp 1612251222
transform 1 0 2046 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_45
timestamp 1612251222
transform 1 0 2030 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_45
timestamp 1612251222
transform 1 0 2014 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_138
timestamp 1612251222
transform -1 0 2014 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_138
timestamp 1612251222
transform -1 0 1848 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_138
timestamp 1612251222
transform -1 0 1832 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_138
timestamp 1612251222
transform -1 0 1816 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_138
timestamp 1612251222
transform -1 0 1800 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_130
timestamp 1612251222
transform -1 0 1784 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_130
timestamp 1612251222
transform -1 0 1618 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_130
timestamp 1612251222
transform -1 0 1602 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_130
timestamp 1612251222
transform -1 0 1586 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_130
timestamp 1612251222
transform -1 0 1570 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_190
timestamp 1612251222
transform -1 0 1554 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_190
timestamp 1612251222
transform -1 0 1388 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_190
timestamp 1612251222
transform -1 0 1372 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_190
timestamp 1612251222
transform -1 0 1356 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_190
timestamp 1612251222
transform -1 0 1340 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_251
timestamp 1612251222
transform -1 0 1324 0 -1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_251
timestamp 1612251222
transform -1 0 1158 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_251
timestamp 1612251222
transform -1 0 1142 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_251
timestamp 1612251222
transform -1 0 1126 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_113
timestamp 1612251222
transform 1 0 944 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_113
timestamp 1612251222
transform 1 0 928 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_113
timestamp 1612251222
transform 1 0 912 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_113
timestamp 1612251222
transform 1 0 896 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_113
timestamp 1612251222
transform 1 0 880 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_107
timestamp 1612251222
transform 1 0 714 0 -1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_107
timestamp 1612251222
transform 1 0 698 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_107
timestamp 1612251222
transform 1 0 682 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_107
timestamp 1612251222
transform 1 0 666 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_132
timestamp 1612251222
transform -1 0 666 0 -1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_132
timestamp 1612251222
transform -1 0 500 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_132
timestamp 1612251222
transform -1 0 484 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_132
timestamp 1612251222
transform -1 0 468 0 -1 3010
box -4 -6 20 206
use POR2X1  POR2X1_127
timestamp 1612251222
transform -1 0 452 0 -1 3010
box -4 -6 170 206
use FILL  FILL1_POR2X1_127
timestamp 1612251222
transform -1 0 286 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_POR2X1_127
timestamp 1612251222
transform -1 0 270 0 -1 3010
box -4 -6 20 206
use FILL  FILL_POR2X1_127
timestamp 1612251222
transform -1 0 254 0 -1 3010
box -4 -6 20 206
use PAND2X1  PAND2X1_128
timestamp 1612251222
transform 1 0 72 0 -1 3010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_128
timestamp 1612251222
transform 1 0 56 0 -1 3010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_128
timestamp 1612251222
transform 1 0 40 0 -1 3010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_128
timestamp 1612251222
transform 1 0 24 0 -1 3010
box -4 -6 20 206
use FILL  FILL_PAND2X1_128
timestamp 1612251222
transform 1 0 8 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_11
timestamp 1612251222
transform 1 0 10252 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_10
timestamp 1612251222
transform 1 0 10236 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_9
timestamp 1612251222
transform 1 0 10220 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_8
timestamp 1612251222
transform 1 0 10204 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_7
timestamp 1612251222
transform 1 0 10188 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_6
timestamp 1612251222
transform 1 0 10172 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_5
timestamp 1612251222
transform 1 0 10156 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_4
timestamp 1612251222
transform 1 0 10140 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_3
timestamp 1612251222
transform 1 0 10124 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_2
timestamp 1612251222
transform 1 0 10108 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_1
timestamp 1612251222
transform 1 0 10092 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_191
timestamp 1612251222
transform 1 0 9926 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_191
timestamp 1612251222
transform 1 0 9910 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_191
timestamp 1612251222
transform 1 0 9894 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_191
timestamp 1612251222
transform 1 0 9878 0 1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_189
timestamp 1612251222
transform 1 0 9712 0 1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_189
timestamp 1612251222
transform 1 0 9696 0 1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_189
timestamp 1612251222
transform 1 0 9680 0 1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_189
timestamp 1612251222
transform 1 0 9664 0 1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_189
timestamp 1612251222
transform 1 0 9648 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_190
timestamp 1612251222
transform 1 0 9482 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_190
timestamp 1612251222
transform 1 0 9466 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_190
timestamp 1612251222
transform 1 0 9450 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_190
timestamp 1612251222
transform 1 0 9434 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_675
timestamp 1612251222
transform -1 0 9434 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_675
timestamp 1612251222
transform -1 0 9268 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_675
timestamp 1612251222
transform -1 0 9252 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_675
timestamp 1612251222
transform -1 0 9236 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_736
timestamp 1612251222
transform -1 0 9220 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_736
timestamp 1612251222
transform -1 0 9054 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_736
timestamp 1612251222
transform -1 0 9038 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_736
timestamp 1612251222
transform -1 0 9022 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_737
timestamp 1612251222
transform 1 0 8840 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_737
timestamp 1612251222
transform 1 0 8824 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_737
timestamp 1612251222
transform 1 0 8808 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_737
timestamp 1612251222
transform 1 0 8792 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_188
timestamp 1612251222
transform -1 0 8792 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_188
timestamp 1612251222
transform -1 0 8626 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_188
timestamp 1612251222
transform -1 0 8610 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_188
timestamp 1612251222
transform -1 0 8594 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_842
timestamp 1612251222
transform 1 0 8412 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_842
timestamp 1612251222
transform 1 0 8396 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_842
timestamp 1612251222
transform 1 0 8380 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_842
timestamp 1612251222
transform 1 0 8364 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_806
timestamp 1612251222
transform 1 0 8198 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_806
timestamp 1612251222
transform 1 0 8182 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_806
timestamp 1612251222
transform 1 0 8166 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_806
timestamp 1612251222
transform 1 0 8150 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_850
timestamp 1612251222
transform -1 0 8150 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_850
timestamp 1612251222
transform -1 0 7984 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_850
timestamp 1612251222
transform -1 0 7968 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_850
timestamp 1612251222
transform -1 0 7952 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_656
timestamp 1612251222
transform 1 0 7770 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_656
timestamp 1612251222
transform 1 0 7754 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_656
timestamp 1612251222
transform 1 0 7738 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_656
timestamp 1612251222
transform 1 0 7722 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_647
timestamp 1612251222
transform 1 0 7556 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_647
timestamp 1612251222
transform 1 0 7540 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_647
timestamp 1612251222
transform 1 0 7524 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_647
timestamp 1612251222
transform 1 0 7508 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_865
timestamp 1612251222
transform 1 0 7342 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_865
timestamp 1612251222
transform 1 0 7326 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_865
timestamp 1612251222
transform 1 0 7310 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_865
timestamp 1612251222
transform 1 0 7294 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_862
timestamp 1612251222
transform 1 0 7128 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_862
timestamp 1612251222
transform 1 0 7112 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_862
timestamp 1612251222
transform 1 0 7096 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_862
timestamp 1612251222
transform 1 0 7080 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_286
timestamp 1612251222
transform 1 0 6914 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_286
timestamp 1612251222
transform 1 0 6898 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_286
timestamp 1612251222
transform 1 0 6882 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_286
timestamp 1612251222
transform 1 0 6866 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_649
timestamp 1612251222
transform 1 0 6700 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_649
timestamp 1612251222
transform 1 0 6684 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_649
timestamp 1612251222
transform 1 0 6668 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_649
timestamp 1612251222
transform 1 0 6652 0 1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_281
timestamp 1612251222
transform -1 0 6652 0 1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_281
timestamp 1612251222
transform -1 0 6486 0 1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_281
timestamp 1612251222
transform -1 0 6470 0 1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_281
timestamp 1612251222
transform -1 0 6454 0 1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_281
timestamp 1612251222
transform -1 0 6438 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_472
timestamp 1612251222
transform 1 0 6256 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_472
timestamp 1612251222
transform 1 0 6240 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_472
timestamp 1612251222
transform 1 0 6224 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_472
timestamp 1612251222
transform 1 0 6208 0 1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_816
timestamp 1612251222
transform -1 0 6208 0 1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_816
timestamp 1612251222
transform -1 0 6042 0 1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_816
timestamp 1612251222
transform -1 0 6026 0 1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_816
timestamp 1612251222
transform -1 0 6010 0 1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_816
timestamp 1612251222
transform -1 0 5994 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_793
timestamp 1612251222
transform 1 0 5812 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_793
timestamp 1612251222
transform 1 0 5796 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_793
timestamp 1612251222
transform 1 0 5780 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_793
timestamp 1612251222
transform 1 0 5764 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_789
timestamp 1612251222
transform 1 0 5598 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_789
timestamp 1612251222
transform 1 0 5582 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_789
timestamp 1612251222
transform 1 0 5566 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_789
timestamp 1612251222
transform 1 0 5550 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_496
timestamp 1612251222
transform -1 0 5550 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_496
timestamp 1612251222
transform -1 0 5384 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_496
timestamp 1612251222
transform -1 0 5368 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_496
timestamp 1612251222
transform -1 0 5352 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_504
timestamp 1612251222
transform 1 0 5170 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_504
timestamp 1612251222
transform 1 0 5154 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_504
timestamp 1612251222
transform 1 0 5138 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_504
timestamp 1612251222
transform 1 0 5122 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_628
timestamp 1612251222
transform 1 0 4956 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_628
timestamp 1612251222
transform 1 0 4940 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_628
timestamp 1612251222
transform 1 0 4924 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_628
timestamp 1612251222
transform 1 0 4908 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_626
timestamp 1612251222
transform -1 0 4908 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_626
timestamp 1612251222
transform -1 0 4742 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_626
timestamp 1612251222
transform -1 0 4726 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_626
timestamp 1612251222
transform -1 0 4710 0 1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_631
timestamp 1612251222
transform -1 0 4694 0 1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_631
timestamp 1612251222
transform -1 0 4528 0 1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_631
timestamp 1612251222
transform -1 0 4512 0 1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_631
timestamp 1612251222
transform -1 0 4496 0 1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_631
timestamp 1612251222
transform -1 0 4480 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_505
timestamp 1612251222
transform 1 0 4298 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_505
timestamp 1612251222
transform 1 0 4282 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_505
timestamp 1612251222
transform 1 0 4266 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_505
timestamp 1612251222
transform 1 0 4250 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_482
timestamp 1612251222
transform -1 0 4250 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_482
timestamp 1612251222
transform -1 0 4084 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_482
timestamp 1612251222
transform -1 0 4068 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_482
timestamp 1612251222
transform -1 0 4052 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_252
timestamp 1612251222
transform -1 0 4036 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_252
timestamp 1612251222
transform -1 0 3870 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_252
timestamp 1612251222
transform -1 0 3854 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_252
timestamp 1612251222
transform -1 0 3838 0 1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_483
timestamp 1612251222
transform -1 0 3822 0 1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_483
timestamp 1612251222
transform -1 0 3656 0 1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_483
timestamp 1612251222
transform -1 0 3640 0 1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_483
timestamp 1612251222
transform -1 0 3624 0 1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_483
timestamp 1612251222
transform -1 0 3608 0 1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_254
timestamp 1612251222
transform -1 0 3592 0 1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_254
timestamp 1612251222
transform -1 0 3426 0 1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_254
timestamp 1612251222
transform -1 0 3410 0 1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_254
timestamp 1612251222
transform -1 0 3394 0 1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_254
timestamp 1612251222
transform -1 0 3378 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_253
timestamp 1612251222
transform 1 0 3196 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_253
timestamp 1612251222
transform 1 0 3180 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_253
timestamp 1612251222
transform 1 0 3164 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_253
timestamp 1612251222
transform 1 0 3148 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_516
timestamp 1612251222
transform -1 0 3148 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_516
timestamp 1612251222
transform -1 0 2982 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_516
timestamp 1612251222
transform -1 0 2966 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_516
timestamp 1612251222
transform -1 0 2950 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_256
timestamp 1612251222
transform -1 0 2934 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_256
timestamp 1612251222
transform -1 0 2768 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_256
timestamp 1612251222
transform -1 0 2752 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_256
timestamp 1612251222
transform -1 0 2736 0 1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_541
timestamp 1612251222
transform -1 0 2720 0 1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_541
timestamp 1612251222
transform -1 0 2554 0 1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_541
timestamp 1612251222
transform -1 0 2538 0 1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_541
timestamp 1612251222
transform -1 0 2522 0 1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_541
timestamp 1612251222
transform -1 0 2506 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_135
timestamp 1612251222
transform -1 0 2490 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_135
timestamp 1612251222
transform -1 0 2324 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_135
timestamp 1612251222
transform -1 0 2308 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_135
timestamp 1612251222
transform -1 0 2292 0 1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_702
timestamp 1612251222
transform -1 0 2276 0 1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_702
timestamp 1612251222
transform -1 0 2110 0 1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_702
timestamp 1612251222
transform -1 0 2094 0 1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_702
timestamp 1612251222
transform -1 0 2078 0 1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_702
timestamp 1612251222
transform -1 0 2062 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_183
timestamp 1612251222
transform -1 0 2046 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_183
timestamp 1612251222
transform -1 0 1880 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_183
timestamp 1612251222
transform -1 0 1864 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_183
timestamp 1612251222
transform -1 0 1848 0 1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_116
timestamp 1612251222
transform 1 0 1666 0 1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_116
timestamp 1612251222
transform 1 0 1650 0 1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_116
timestamp 1612251222
transform 1 0 1634 0 1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_116
timestamp 1612251222
transform 1 0 1618 0 1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_116
timestamp 1612251222
transform 1 0 1602 0 1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_114
timestamp 1612251222
transform 1 0 1436 0 1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_114
timestamp 1612251222
transform 1 0 1420 0 1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_114
timestamp 1612251222
transform 1 0 1404 0 1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_114
timestamp 1612251222
transform 1 0 1388 0 1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_114
timestamp 1612251222
transform 1 0 1372 0 1 2610
box -4 -6 20 206
use POR2X1  POR2X1_106
timestamp 1612251222
transform 1 0 1206 0 1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_106
timestamp 1612251222
transform 1 0 1190 0 1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_106
timestamp 1612251222
transform 1 0 1174 0 1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_106
timestamp 1612251222
transform 1 0 1158 0 1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_540
timestamp 1612251222
transform -1 0 1158 0 1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_540
timestamp 1612251222
transform -1 0 992 0 1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_540
timestamp 1612251222
transform -1 0 976 0 1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_540
timestamp 1612251222
transform -1 0 960 0 1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_540
timestamp 1612251222
transform -1 0 944 0 1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_553
timestamp 1612251222
transform -1 0 928 0 1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_553
timestamp 1612251222
transform -1 0 762 0 1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_553
timestamp 1612251222
transform -1 0 746 0 1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_553
timestamp 1612251222
transform -1 0 730 0 1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_553
timestamp 1612251222
transform -1 0 714 0 1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_554
timestamp 1612251222
transform -1 0 698 0 1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_554
timestamp 1612251222
transform -1 0 532 0 1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_554
timestamp 1612251222
transform -1 0 516 0 1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_554
timestamp 1612251222
transform -1 0 500 0 1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_554
timestamp 1612251222
transform -1 0 484 0 1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_563
timestamp 1612251222
transform -1 0 468 0 1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_563
timestamp 1612251222
transform -1 0 302 0 1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_563
timestamp 1612251222
transform -1 0 286 0 1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_563
timestamp 1612251222
transform -1 0 270 0 1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_563
timestamp 1612251222
transform -1 0 254 0 1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_570
timestamp 1612251222
transform -1 0 238 0 1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_570
timestamp 1612251222
transform -1 0 72 0 1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_570
timestamp 1612251222
transform -1 0 56 0 1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_570
timestamp 1612251222
transform -1 0 40 0 1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_570
timestamp 1612251222
transform -1 0 24 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_11
timestamp 1612251222
transform -1 0 10262 0 -1 2610
box -4 -6 20 206
use FILL  FILL_13_10
timestamp 1612251222
transform -1 0 10246 0 -1 2610
box -4 -6 20 206
use FILL  FILL_13_9
timestamp 1612251222
transform -1 0 10230 0 -1 2610
box -4 -6 20 206
use FILL  FILL_13_8
timestamp 1612251222
transform -1 0 10214 0 -1 2610
box -4 -6 20 206
use FILL  FILL_13_7
timestamp 1612251222
transform -1 0 10198 0 -1 2610
box -4 -6 20 206
use FILL  FILL_13_6
timestamp 1612251222
transform -1 0 10182 0 -1 2610
box -4 -6 20 206
use FILL  FILL_13_5
timestamp 1612251222
transform -1 0 10166 0 -1 2610
box -4 -6 20 206
use FILL  FILL_13_4
timestamp 1612251222
transform -1 0 10150 0 -1 2610
box -4 -6 20 206
use FILL  FILL_13_3
timestamp 1612251222
transform -1 0 10134 0 -1 2610
box -4 -6 20 206
use FILL  FILL_13_2
timestamp 1612251222
transform -1 0 10118 0 -1 2610
box -4 -6 20 206
use FILL  FILL_13_1
timestamp 1612251222
transform -1 0 10102 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_187
timestamp 1612251222
transform 1 0 9920 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_187
timestamp 1612251222
transform 1 0 9904 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_187
timestamp 1612251222
transform 1 0 9888 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_187
timestamp 1612251222
transform 1 0 9872 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_187
timestamp 1612251222
transform 1 0 9856 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_172
timestamp 1612251222
transform 1 0 9690 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_172
timestamp 1612251222
transform 1 0 9674 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_172
timestamp 1612251222
transform 1 0 9658 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_172
timestamp 1612251222
transform 1 0 9642 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_172
timestamp 1612251222
transform 1 0 9626 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_437
timestamp 1612251222
transform -1 0 9626 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_437
timestamp 1612251222
transform -1 0 9460 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_437
timestamp 1612251222
transform -1 0 9444 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_437
timestamp 1612251222
transform -1 0 9428 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_437
timestamp 1612251222
transform -1 0 9412 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_674
timestamp 1612251222
transform 1 0 9230 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_674
timestamp 1612251222
transform 1 0 9214 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_674
timestamp 1612251222
transform 1 0 9198 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_674
timestamp 1612251222
transform 1 0 9182 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_674
timestamp 1612251222
transform 1 0 9166 0 -1 2610
box -4 -6 20 206
use POR2X1  POR2X1_741
timestamp 1612251222
transform 1 0 9000 0 -1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_741
timestamp 1612251222
transform 1 0 8984 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_741
timestamp 1612251222
transform 1 0 8968 0 -1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_741
timestamp 1612251222
transform 1 0 8952 0 -1 2610
box -4 -6 20 206
use POR2X1  POR2X1_539
timestamp 1612251222
transform 1 0 8786 0 -1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_539
timestamp 1612251222
transform 1 0 8770 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_539
timestamp 1612251222
transform 1 0 8754 0 -1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_539
timestamp 1612251222
transform 1 0 8738 0 -1 2610
box -4 -6 20 206
use POR2X1  POR2X1_733
timestamp 1612251222
transform 1 0 8572 0 -1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_733
timestamp 1612251222
transform 1 0 8556 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_733
timestamp 1612251222
transform 1 0 8540 0 -1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_733
timestamp 1612251222
transform 1 0 8524 0 -1 2610
box -4 -6 20 206
use POR2X1  POR2X1_830
timestamp 1612251222
transform 1 0 8358 0 -1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_830
timestamp 1612251222
transform 1 0 8342 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_830
timestamp 1612251222
transform 1 0 8326 0 -1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_830
timestamp 1612251222
transform 1 0 8310 0 -1 2610
box -4 -6 20 206
use POR2X1  POR2X1_841
timestamp 1612251222
transform -1 0 8310 0 -1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_841
timestamp 1612251222
transform -1 0 8144 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_841
timestamp 1612251222
transform -1 0 8128 0 -1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_841
timestamp 1612251222
transform -1 0 8112 0 -1 2610
box -4 -6 20 206
use POR2X1  POR2X1_851
timestamp 1612251222
transform -1 0 8096 0 -1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_851
timestamp 1612251222
transform -1 0 7930 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_851
timestamp 1612251222
transform -1 0 7914 0 -1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_851
timestamp 1612251222
transform -1 0 7898 0 -1 2610
box -4 -6 20 206
use POR2X1  POR2X1_858
timestamp 1612251222
transform -1 0 7882 0 -1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_858
timestamp 1612251222
transform -1 0 7716 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_858
timestamp 1612251222
transform -1 0 7700 0 -1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_858
timestamp 1612251222
transform -1 0 7684 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_108
timestamp 1612251222
transform -1 0 7668 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_108
timestamp 1612251222
transform -1 0 7502 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_108
timestamp 1612251222
transform -1 0 7486 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_108
timestamp 1612251222
transform -1 0 7470 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_108
timestamp 1612251222
transform -1 0 7454 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_536
timestamp 1612251222
transform -1 0 7438 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_536
timestamp 1612251222
transform -1 0 7272 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_536
timestamp 1612251222
transform -1 0 7256 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_536
timestamp 1612251222
transform -1 0 7240 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_536
timestamp 1612251222
transform -1 0 7224 0 -1 2610
box -4 -6 20 206
use POR2X1  POR2X1_537
timestamp 1612251222
transform -1 0 7208 0 -1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_537
timestamp 1612251222
transform -1 0 7042 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_537
timestamp 1612251222
transform -1 0 7026 0 -1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_537
timestamp 1612251222
transform -1 0 7010 0 -1 2610
box -4 -6 20 206
use POR2X1  POR2X1_121
timestamp 1612251222
transform -1 0 6994 0 -1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_121
timestamp 1612251222
transform -1 0 6828 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_121
timestamp 1612251222
transform -1 0 6812 0 -1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_121
timestamp 1612251222
transform -1 0 6796 0 -1 2610
box -4 -6 20 206
use POR2X1  POR2X1_643
timestamp 1612251222
transform -1 0 6780 0 -1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_643
timestamp 1612251222
transform -1 0 6614 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_643
timestamp 1612251222
transform -1 0 6598 0 -1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_643
timestamp 1612251222
transform -1 0 6582 0 -1 2610
box -4 -6 20 206
use POR2X1  POR2X1_285
timestamp 1612251222
transform 1 0 6400 0 -1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_285
timestamp 1612251222
transform 1 0 6384 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_285
timestamp 1612251222
transform 1 0 6368 0 -1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_285
timestamp 1612251222
transform 1 0 6352 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_282
timestamp 1612251222
transform 1 0 6186 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_282
timestamp 1612251222
transform 1 0 6170 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_282
timestamp 1612251222
transform 1 0 6154 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_282
timestamp 1612251222
transform 1 0 6138 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_282
timestamp 1612251222
transform 1 0 6122 0 -1 2610
box -4 -6 20 206
use POR2X1  POR2X1_185
timestamp 1612251222
transform 1 0 5956 0 -1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_185
timestamp 1612251222
transform 1 0 5940 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_185
timestamp 1612251222
transform 1 0 5924 0 -1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_185
timestamp 1612251222
transform 1 0 5908 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_411
timestamp 1612251222
transform 1 0 5742 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_411
timestamp 1612251222
transform 1 0 5726 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_411
timestamp 1612251222
transform 1 0 5710 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_411
timestamp 1612251222
transform 1 0 5694 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_411
timestamp 1612251222
transform 1 0 5678 0 -1 2610
box -4 -6 20 206
use POR2X1  POR2X1_410
timestamp 1612251222
transform 1 0 5512 0 -1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_410
timestamp 1612251222
transform 1 0 5496 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_410
timestamp 1612251222
transform 1 0 5480 0 -1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_410
timestamp 1612251222
transform 1 0 5464 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_748
timestamp 1612251222
transform 1 0 5298 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_748
timestamp 1612251222
transform 1 0 5282 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_748
timestamp 1612251222
transform 1 0 5266 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_748
timestamp 1612251222
transform 1 0 5250 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_748
timestamp 1612251222
transform 1 0 5234 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_699
timestamp 1612251222
transform 1 0 5068 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_699
timestamp 1612251222
transform 1 0 5052 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_699
timestamp 1612251222
transform 1 0 5036 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_699
timestamp 1612251222
transform 1 0 5020 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_699
timestamp 1612251222
transform 1 0 5004 0 -1 2610
box -4 -6 20 206
use POR2X1  POR2X1_627
timestamp 1612251222
transform -1 0 5004 0 -1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_627
timestamp 1612251222
transform -1 0 4838 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_627
timestamp 1612251222
transform -1 0 4822 0 -1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_627
timestamp 1612251222
transform -1 0 4806 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_629
timestamp 1612251222
transform -1 0 4790 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_629
timestamp 1612251222
transform -1 0 4624 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_629
timestamp 1612251222
transform -1 0 4608 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_629
timestamp 1612251222
transform -1 0 4592 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_629
timestamp 1612251222
transform -1 0 4576 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_507
timestamp 1612251222
transform -1 0 4560 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_507
timestamp 1612251222
transform -1 0 4394 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_507
timestamp 1612251222
transform -1 0 4378 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_507
timestamp 1612251222
transform -1 0 4362 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_507
timestamp 1612251222
transform -1 0 4346 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_630
timestamp 1612251222
transform -1 0 4330 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_630
timestamp 1612251222
transform -1 0 4164 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_630
timestamp 1612251222
transform -1 0 4148 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_630
timestamp 1612251222
transform -1 0 4132 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_630
timestamp 1612251222
transform -1 0 4116 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_508
timestamp 1612251222
transform -1 0 4100 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_508
timestamp 1612251222
transform -1 0 3934 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_508
timestamp 1612251222
transform -1 0 3918 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_508
timestamp 1612251222
transform -1 0 3902 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_508
timestamp 1612251222
transform -1 0 3886 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_632
timestamp 1612251222
transform -1 0 3870 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_632
timestamp 1612251222
transform -1 0 3704 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_632
timestamp 1612251222
transform -1 0 3688 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_632
timestamp 1612251222
transform -1 0 3672 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_632
timestamp 1612251222
transform -1 0 3656 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_513
timestamp 1612251222
transform -1 0 3640 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_513
timestamp 1612251222
transform -1 0 3474 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_513
timestamp 1612251222
transform -1 0 3458 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_513
timestamp 1612251222
transform -1 0 3442 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_513
timestamp 1612251222
transform -1 0 3426 0 -1 2610
box -4 -6 20 206
use POR2X1  POR2X1_56
timestamp 1612251222
transform -1 0 3410 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_POR2X1_56
timestamp 1612251222
transform -1 0 3244 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_POR2X1_56
timestamp 1612251222
transform -1 0 3228 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_56
timestamp 1612251222
transform -1 0 3212 0 -1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_56
timestamp 1612251222
transform -1 0 3196 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_456
timestamp 1612251222
transform 1 0 3014 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_456
timestamp 1612251222
transform 1 0 2998 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_456
timestamp 1612251222
transform 1 0 2982 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_456
timestamp 1612251222
transform 1 0 2966 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_456
timestamp 1612251222
transform 1 0 2950 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_515
timestamp 1612251222
transform 1 0 2784 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_515
timestamp 1612251222
transform 1 0 2768 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_515
timestamp 1612251222
transform 1 0 2752 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_515
timestamp 1612251222
transform 1 0 2736 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_515
timestamp 1612251222
transform 1 0 2720 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_344
timestamp 1612251222
transform -1 0 2720 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_344
timestamp 1612251222
transform -1 0 2554 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_344
timestamp 1612251222
transform -1 0 2538 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_344
timestamp 1612251222
transform -1 0 2522 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_344
timestamp 1612251222
transform -1 0 2506 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_514
timestamp 1612251222
transform 1 0 2324 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_514
timestamp 1612251222
transform 1 0 2308 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_514
timestamp 1612251222
transform 1 0 2292 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_514
timestamp 1612251222
transform 1 0 2276 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_514
timestamp 1612251222
transform 1 0 2260 0 -1 2610
box -4 -6 20 206
use POR2X1  POR2X1_136
timestamp 1612251222
transform -1 0 2260 0 -1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_136
timestamp 1612251222
transform -1 0 2094 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_136
timestamp 1612251222
transform -1 0 2078 0 -1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_136
timestamp 1612251222
transform -1 0 2062 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_556
timestamp 1612251222
transform -1 0 2046 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_556
timestamp 1612251222
transform -1 0 1880 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_556
timestamp 1612251222
transform -1 0 1864 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_556
timestamp 1612251222
transform -1 0 1848 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_556
timestamp 1612251222
transform -1 0 1832 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_115
timestamp 1612251222
transform -1 0 1816 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_115
timestamp 1612251222
transform -1 0 1650 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_115
timestamp 1612251222
transform -1 0 1634 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_115
timestamp 1612251222
transform -1 0 1618 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_115
timestamp 1612251222
transform -1 0 1602 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_830
timestamp 1612251222
transform 1 0 1420 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_830
timestamp 1612251222
transform 1 0 1404 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_830
timestamp 1612251222
transform 1 0 1388 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_830
timestamp 1612251222
transform 1 0 1372 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_830
timestamp 1612251222
transform 1 0 1356 0 -1 2610
box -4 -6 20 206
use POR2X1  POR2X1_108
timestamp 1612251222
transform 1 0 1190 0 -1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_108
timestamp 1612251222
transform 1 0 1174 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_108
timestamp 1612251222
transform 1 0 1158 0 -1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_108
timestamp 1612251222
transform 1 0 1142 0 -1 2610
box -4 -6 20 206
use POR2X1  POR2X1_178
timestamp 1612251222
transform 1 0 976 0 -1 2610
box -4 -6 170 206
use FILL  FILL1_POR2X1_178
timestamp 1612251222
transform 1 0 960 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_POR2X1_178
timestamp 1612251222
transform 1 0 944 0 -1 2610
box -4 -6 20 206
use FILL  FILL_POR2X1_178
timestamp 1612251222
transform 1 0 928 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_105
timestamp 1612251222
transform 1 0 762 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_105
timestamp 1612251222
transform 1 0 746 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_105
timestamp 1612251222
transform 1 0 730 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_105
timestamp 1612251222
transform 1 0 714 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_105
timestamp 1612251222
transform 1 0 698 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_348
timestamp 1612251222
transform 1 0 532 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_348
timestamp 1612251222
transform 1 0 516 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_348
timestamp 1612251222
transform 1 0 500 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_348
timestamp 1612251222
transform 1 0 484 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_348
timestamp 1612251222
transform 1 0 468 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_562
timestamp 1612251222
transform -1 0 468 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_562
timestamp 1612251222
transform -1 0 302 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_562
timestamp 1612251222
transform -1 0 286 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_562
timestamp 1612251222
transform -1 0 270 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_562
timestamp 1612251222
transform -1 0 254 0 -1 2610
box -4 -6 20 206
use PAND2X1  PAND2X1_577
timestamp 1612251222
transform 1 0 72 0 -1 2610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_577
timestamp 1612251222
transform 1 0 56 0 -1 2610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_577
timestamp 1612251222
transform 1 0 40 0 -1 2610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_577
timestamp 1612251222
transform 1 0 24 0 -1 2610
box -4 -6 20 206
use FILL  FILL_PAND2X1_577
timestamp 1612251222
transform 1 0 8 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_13
timestamp 1612251222
transform 1 0 10252 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_12
timestamp 1612251222
transform 1 0 10236 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_11
timestamp 1612251222
transform 1 0 10220 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_10
timestamp 1612251222
transform 1 0 10204 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_9
timestamp 1612251222
transform 1 0 10188 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_8
timestamp 1612251222
transform 1 0 10172 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_7
timestamp 1612251222
transform 1 0 10156 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_6
timestamp 1612251222
transform 1 0 10140 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_5
timestamp 1612251222
transform 1 0 10124 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_4
timestamp 1612251222
transform 1 0 10108 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_3
timestamp 1612251222
transform 1 0 10092 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_2
timestamp 1612251222
transform 1 0 10076 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_1
timestamp 1612251222
transform 1 0 10060 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_739
timestamp 1612251222
transform 1 0 9894 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_739
timestamp 1612251222
transform 1 0 9878 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_739
timestamp 1612251222
transform 1 0 9862 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_739
timestamp 1612251222
transform 1 0 9846 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_727
timestamp 1612251222
transform -1 0 9846 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_727
timestamp 1612251222
transform -1 0 9680 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_727
timestamp 1612251222
transform -1 0 9664 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_727
timestamp 1612251222
transform -1 0 9648 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_440
timestamp 1612251222
transform -1 0 9632 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_440
timestamp 1612251222
transform -1 0 9466 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_440
timestamp 1612251222
transform -1 0 9450 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_440
timestamp 1612251222
transform -1 0 9434 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_732
timestamp 1612251222
transform 1 0 9252 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_732
timestamp 1612251222
transform 1 0 9236 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_732
timestamp 1612251222
transform 1 0 9220 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_732
timestamp 1612251222
transform 1 0 9204 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_151
timestamp 1612251222
transform -1 0 9204 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_151
timestamp 1612251222
transform -1 0 9038 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_151
timestamp 1612251222
transform -1 0 9022 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_151
timestamp 1612251222
transform -1 0 9006 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_186
timestamp 1612251222
transform 1 0 8824 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_186
timestamp 1612251222
transform 1 0 8808 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_186
timestamp 1612251222
transform 1 0 8792 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_186
timestamp 1612251222
transform 1 0 8776 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_662
timestamp 1612251222
transform 1 0 8610 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_662
timestamp 1612251222
transform 1 0 8594 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_662
timestamp 1612251222
transform 1 0 8578 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_662
timestamp 1612251222
transform 1 0 8562 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_308
timestamp 1612251222
transform 1 0 8396 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_308
timestamp 1612251222
transform 1 0 8380 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_308
timestamp 1612251222
transform 1 0 8364 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_308
timestamp 1612251222
transform 1 0 8348 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_512
timestamp 1612251222
transform -1 0 8348 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_512
timestamp 1612251222
transform -1 0 8182 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_512
timestamp 1612251222
transform -1 0 8166 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_512
timestamp 1612251222
transform -1 0 8150 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_840
timestamp 1612251222
transform 1 0 7968 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_840
timestamp 1612251222
transform 1 0 7952 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_840
timestamp 1612251222
transform 1 0 7936 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_840
timestamp 1612251222
transform 1 0 7920 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_660
timestamp 1612251222
transform 1 0 7754 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_660
timestamp 1612251222
transform 1 0 7738 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_660
timestamp 1612251222
transform 1 0 7722 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_660
timestamp 1612251222
transform 1 0 7706 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_784
timestamp 1612251222
transform 1 0 7540 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_784
timestamp 1612251222
transform 1 0 7524 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_784
timestamp 1612251222
transform 1 0 7508 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_784
timestamp 1612251222
transform 1 0 7492 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_777
timestamp 1612251222
transform 1 0 7326 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_777
timestamp 1612251222
transform 1 0 7310 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_777
timestamp 1612251222
transform 1 0 7294 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_777
timestamp 1612251222
transform 1 0 7278 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_389
timestamp 1612251222
transform 1 0 7112 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_389
timestamp 1612251222
transform 1 0 7096 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_389
timestamp 1612251222
transform 1 0 7080 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_389
timestamp 1612251222
transform 1 0 7064 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_654
timestamp 1612251222
transform 1 0 6898 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_654
timestamp 1612251222
transform 1 0 6882 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_654
timestamp 1612251222
transform 1 0 6866 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_654
timestamp 1612251222
transform 1 0 6850 0 1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_119
timestamp 1612251222
transform 1 0 6684 0 1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_119
timestamp 1612251222
transform 1 0 6668 0 1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_119
timestamp 1612251222
transform 1 0 6652 0 1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_119
timestamp 1612251222
transform 1 0 6636 0 1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_119
timestamp 1612251222
transform 1 0 6620 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_706
timestamp 1612251222
transform 1 0 6454 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_706
timestamp 1612251222
transform 1 0 6438 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_706
timestamp 1612251222
transform 1 0 6422 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_706
timestamp 1612251222
transform 1 0 6406 0 1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_693
timestamp 1612251222
transform 1 0 6240 0 1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_693
timestamp 1612251222
transform 1 0 6224 0 1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_693
timestamp 1612251222
transform 1 0 6208 0 1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_693
timestamp 1612251222
transform 1 0 6192 0 1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_693
timestamp 1612251222
transform 1 0 6176 0 1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_701
timestamp 1612251222
transform 1 0 6010 0 1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_701
timestamp 1612251222
transform 1 0 5994 0 1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_701
timestamp 1612251222
transform 1 0 5978 0 1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_701
timestamp 1612251222
transform 1 0 5962 0 1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_701
timestamp 1612251222
transform 1 0 5946 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_709
timestamp 1612251222
transform 1 0 5780 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_709
timestamp 1612251222
transform 1 0 5764 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_709
timestamp 1612251222
transform 1 0 5748 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_709
timestamp 1612251222
transform 1 0 5732 0 1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_637
timestamp 1612251222
transform 1 0 5566 0 1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_637
timestamp 1612251222
transform 1 0 5550 0 1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_637
timestamp 1612251222
transform 1 0 5534 0 1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_637
timestamp 1612251222
transform 1 0 5518 0 1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_637
timestamp 1612251222
transform 1 0 5502 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_585
timestamp 1612251222
transform 1 0 5336 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_585
timestamp 1612251222
transform 1 0 5320 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_585
timestamp 1612251222
transform 1 0 5304 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_585
timestamp 1612251222
transform 1 0 5288 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_586
timestamp 1612251222
transform 1 0 5122 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_586
timestamp 1612251222
transform 1 0 5106 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_586
timestamp 1612251222
transform 1 0 5090 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_586
timestamp 1612251222
transform 1 0 5074 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_422
timestamp 1612251222
transform 1 0 4908 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_422
timestamp 1612251222
transform 1 0 4892 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_422
timestamp 1612251222
transform 1 0 4876 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_422
timestamp 1612251222
transform 1 0 4860 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_387
timestamp 1612251222
transform -1 0 4860 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_387
timestamp 1612251222
transform -1 0 4694 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_387
timestamp 1612251222
transform -1 0 4678 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_387
timestamp 1612251222
transform -1 0 4662 0 1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_777
timestamp 1612251222
transform 1 0 4480 0 1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_777
timestamp 1612251222
transform 1 0 4464 0 1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_777
timestamp 1612251222
transform 1 0 4448 0 1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_777
timestamp 1612251222
transform 1 0 4432 0 1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_777
timestamp 1612251222
transform 1 0 4416 0 1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_784
timestamp 1612251222
transform -1 0 4416 0 1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_784
timestamp 1612251222
transform -1 0 4250 0 1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_784
timestamp 1612251222
transform -1 0 4234 0 1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_784
timestamp 1612251222
transform -1 0 4218 0 1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_784
timestamp 1612251222
transform -1 0 4202 0 1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_778
timestamp 1612251222
transform 1 0 4020 0 1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_778
timestamp 1612251222
transform 1 0 4004 0 1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_778
timestamp 1612251222
transform 1 0 3988 0 1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_778
timestamp 1612251222
transform 1 0 3972 0 1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_778
timestamp 1612251222
transform 1 0 3956 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_371
timestamp 1612251222
transform -1 0 3956 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_371
timestamp 1612251222
transform -1 0 3790 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_371
timestamp 1612251222
transform -1 0 3774 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_371
timestamp 1612251222
transform -1 0 3758 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_372
timestamp 1612251222
transform -1 0 3742 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_372
timestamp 1612251222
transform -1 0 3576 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_372
timestamp 1612251222
transform -1 0 3560 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_372
timestamp 1612251222
transform -1 0 3544 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_423
timestamp 1612251222
transform -1 0 3528 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_423
timestamp 1612251222
transform -1 0 3362 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_423
timestamp 1612251222
transform -1 0 3346 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_423
timestamp 1612251222
transform -1 0 3330 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_110
timestamp 1612251222
transform 1 0 3148 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_110
timestamp 1612251222
transform 1 0 3132 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_110
timestamp 1612251222
transform 1 0 3116 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_110
timestamp 1612251222
transform 1 0 3100 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_417
timestamp 1612251222
transform -1 0 3100 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_417
timestamp 1612251222
transform -1 0 2934 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_417
timestamp 1612251222
transform -1 0 2918 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_417
timestamp 1612251222
transform -1 0 2902 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_368
timestamp 1612251222
transform -1 0 2886 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_368
timestamp 1612251222
transform -1 0 2720 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_368
timestamp 1612251222
transform -1 0 2704 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_368
timestamp 1612251222
transform -1 0 2688 0 1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_458
timestamp 1612251222
transform 1 0 2506 0 1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_458
timestamp 1612251222
transform 1 0 2490 0 1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_458
timestamp 1612251222
transform 1 0 2474 0 1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_458
timestamp 1612251222
transform 1 0 2458 0 1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_458
timestamp 1612251222
transform 1 0 2442 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_111
timestamp 1612251222
transform -1 0 2442 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_111
timestamp 1612251222
transform -1 0 2276 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_111
timestamp 1612251222
transform -1 0 2260 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_111
timestamp 1612251222
transform -1 0 2244 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_310
timestamp 1612251222
transform -1 0 2228 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_310
timestamp 1612251222
transform -1 0 2062 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_310
timestamp 1612251222
transform -1 0 2046 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_310
timestamp 1612251222
transform -1 0 2030 0 1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_715
timestamp 1612251222
transform -1 0 2014 0 1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_715
timestamp 1612251222
transform -1 0 1848 0 1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_715
timestamp 1612251222
transform -1 0 1832 0 1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_715
timestamp 1612251222
transform -1 0 1816 0 1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_715
timestamp 1612251222
transform -1 0 1800 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_309
timestamp 1612251222
transform -1 0 1784 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_309
timestamp 1612251222
transform -1 0 1618 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_309
timestamp 1612251222
transform -1 0 1602 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_309
timestamp 1612251222
transform -1 0 1586 0 1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_294
timestamp 1612251222
transform -1 0 1570 0 1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_294
timestamp 1612251222
transform -1 0 1404 0 1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_294
timestamp 1612251222
transform -1 0 1388 0 1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_294
timestamp 1612251222
transform -1 0 1372 0 1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_294
timestamp 1612251222
transform -1 0 1356 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_179
timestamp 1612251222
transform -1 0 1340 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_179
timestamp 1612251222
transform -1 0 1174 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_179
timestamp 1612251222
transform -1 0 1158 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_179
timestamp 1612251222
transform -1 0 1142 0 1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_181
timestamp 1612251222
transform -1 0 1126 0 1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_181
timestamp 1612251222
transform -1 0 960 0 1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_181
timestamp 1612251222
transform -1 0 944 0 1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_181
timestamp 1612251222
transform -1 0 928 0 1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_181
timestamp 1612251222
transform -1 0 912 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_292
timestamp 1612251222
transform -1 0 896 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_292
timestamp 1612251222
transform -1 0 730 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_292
timestamp 1612251222
transform -1 0 714 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_292
timestamp 1612251222
transform -1 0 698 0 1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_346
timestamp 1612251222
transform -1 0 682 0 1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_346
timestamp 1612251222
transform -1 0 516 0 1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_346
timestamp 1612251222
transform -1 0 500 0 1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_346
timestamp 1612251222
transform -1 0 484 0 1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_346
timestamp 1612251222
transform -1 0 468 0 1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_260
timestamp 1612251222
transform -1 0 452 0 1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_260
timestamp 1612251222
transform -1 0 286 0 1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_260
timestamp 1612251222
transform -1 0 270 0 1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_260
timestamp 1612251222
transform -1 0 254 0 1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_260
timestamp 1612251222
transform -1 0 238 0 1 2210
box -4 -6 20 206
use POR2X1  POR2X1_261
timestamp 1612251222
transform -1 0 222 0 1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_261
timestamp 1612251222
transform -1 0 56 0 1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_261
timestamp 1612251222
transform -1 0 40 0 1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_261
timestamp 1612251222
transform -1 0 24 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_1
timestamp 1612251222
transform -1 0 10268 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_740
timestamp 1612251222
transform 1 0 10086 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_740
timestamp 1612251222
transform 1 0 10070 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_740
timestamp 1612251222
transform 1 0 10054 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_740
timestamp 1612251222
transform 1 0 10038 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_738
timestamp 1612251222
transform 1 0 9872 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_738
timestamp 1612251222
transform 1 0 9856 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_738
timestamp 1612251222
transform 1 0 9840 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_738
timestamp 1612251222
transform 1 0 9824 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_731
timestamp 1612251222
transform 1 0 9658 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_731
timestamp 1612251222
transform 1 0 9642 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_731
timestamp 1612251222
transform 1 0 9626 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_731
timestamp 1612251222
transform 1 0 9610 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_726
timestamp 1612251222
transform 1 0 9444 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_726
timestamp 1612251222
transform 1 0 9428 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_726
timestamp 1612251222
transform 1 0 9412 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_726
timestamp 1612251222
transform 1 0 9396 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_152
timestamp 1612251222
transform 1 0 9230 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_152
timestamp 1612251222
transform 1 0 9214 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_152
timestamp 1612251222
transform 1 0 9198 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_152
timestamp 1612251222
transform 1 0 9182 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_152
timestamp 1612251222
transform 1 0 9166 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_594
timestamp 1612251222
transform -1 0 9166 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_594
timestamp 1612251222
transform -1 0 9000 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_594
timestamp 1612251222
transform -1 0 8984 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_594
timestamp 1612251222
transform -1 0 8968 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_594
timestamp 1612251222
transform -1 0 8952 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_653
timestamp 1612251222
transform 1 0 8770 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_653
timestamp 1612251222
transform 1 0 8754 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_653
timestamp 1612251222
transform 1 0 8738 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_653
timestamp 1612251222
transform 1 0 8722 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_661
timestamp 1612251222
transform -1 0 8722 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_661
timestamp 1612251222
transform -1 0 8556 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_661
timestamp 1612251222
transform -1 0 8540 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_661
timestamp 1612251222
transform -1 0 8524 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_306
timestamp 1612251222
transform 1 0 8342 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_306
timestamp 1612251222
transform 1 0 8326 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_306
timestamp 1612251222
transform 1 0 8310 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_306
timestamp 1612251222
transform 1 0 8294 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_306
timestamp 1612251222
transform 1 0 8278 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_832
timestamp 1612251222
transform 1 0 8112 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_832
timestamp 1612251222
transform 1 0 8096 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_832
timestamp 1612251222
transform 1 0 8080 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_832
timestamp 1612251222
transform 1 0 8064 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_513
timestamp 1612251222
transform 1 0 7898 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_513
timestamp 1612251222
transform 1 0 7882 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_513
timestamp 1612251222
transform 1 0 7866 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_513
timestamp 1612251222
transform 1 0 7850 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_307
timestamp 1612251222
transform 1 0 7684 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_307
timestamp 1612251222
transform 1 0 7668 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_307
timestamp 1612251222
transform 1 0 7652 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_307
timestamp 1612251222
transform 1 0 7636 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_655
timestamp 1612251222
transform 1 0 7470 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_655
timestamp 1612251222
transform 1 0 7454 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_655
timestamp 1612251222
transform 1 0 7438 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_655
timestamp 1612251222
transform 1 0 7422 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_305
timestamp 1612251222
transform 1 0 7256 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_305
timestamp 1612251222
transform 1 0 7240 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_305
timestamp 1612251222
transform 1 0 7224 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_305
timestamp 1612251222
transform 1 0 7208 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_305
timestamp 1612251222
transform 1 0 7192 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_385
timestamp 1612251222
transform 1 0 7026 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_385
timestamp 1612251222
transform 1 0 7010 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_385
timestamp 1612251222
transform 1 0 6994 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_385
timestamp 1612251222
transform 1 0 6978 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_385
timestamp 1612251222
transform 1 0 6962 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_725
timestamp 1612251222
transform 1 0 6796 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_725
timestamp 1612251222
transform 1 0 6780 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_725
timestamp 1612251222
transform 1 0 6764 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_725
timestamp 1612251222
transform 1 0 6748 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_713
timestamp 1612251222
transform 1 0 6582 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_713
timestamp 1612251222
transform 1 0 6566 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_713
timestamp 1612251222
transform 1 0 6550 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_713
timestamp 1612251222
transform 1 0 6534 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_692
timestamp 1612251222
transform 1 0 6368 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_692
timestamp 1612251222
transform 1 0 6352 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_692
timestamp 1612251222
transform 1 0 6336 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_692
timestamp 1612251222
transform 1 0 6320 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_692
timestamp 1612251222
transform 1 0 6304 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_711
timestamp 1612251222
transform 1 0 6138 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_711
timestamp 1612251222
transform 1 0 6122 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_711
timestamp 1612251222
transform 1 0 6106 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_711
timestamp 1612251222
transform 1 0 6090 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_710
timestamp 1612251222
transform 1 0 5924 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_710
timestamp 1612251222
transform 1 0 5908 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_710
timestamp 1612251222
transform 1 0 5892 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_710
timestamp 1612251222
transform 1 0 5876 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_698
timestamp 1612251222
transform 1 0 5710 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_698
timestamp 1612251222
transform 1 0 5694 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_698
timestamp 1612251222
transform 1 0 5678 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_698
timestamp 1612251222
transform 1 0 5662 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_698
timestamp 1612251222
transform 1 0 5646 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_753
timestamp 1612251222
transform -1 0 5646 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_753
timestamp 1612251222
transform -1 0 5480 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_753
timestamp 1612251222
transform -1 0 5464 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_753
timestamp 1612251222
transform -1 0 5448 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_753
timestamp 1612251222
transform -1 0 5432 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_638
timestamp 1612251222
transform -1 0 5416 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_638
timestamp 1612251222
transform -1 0 5250 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_638
timestamp 1612251222
transform -1 0 5234 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_638
timestamp 1612251222
transform -1 0 5218 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_638
timestamp 1612251222
transform -1 0 5202 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_651
timestamp 1612251222
transform -1 0 5186 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_651
timestamp 1612251222
transform -1 0 5020 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_651
timestamp 1612251222
transform -1 0 5004 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_651
timestamp 1612251222
transform -1 0 4988 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_651
timestamp 1612251222
transform -1 0 4972 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_620
timestamp 1612251222
transform 1 0 4790 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_620
timestamp 1612251222
transform 1 0 4774 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_620
timestamp 1612251222
transform 1 0 4758 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_620
timestamp 1612251222
transform 1 0 4742 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_620
timestamp 1612251222
transform 1 0 4726 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_613
timestamp 1612251222
transform 1 0 4560 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_613
timestamp 1612251222
transform 1 0 4544 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_613
timestamp 1612251222
transform 1 0 4528 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_613
timestamp 1612251222
transform 1 0 4512 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_305
timestamp 1612251222
transform -1 0 4512 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_305
timestamp 1612251222
transform -1 0 4346 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_305
timestamp 1612251222
transform -1 0 4330 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_305
timestamp 1612251222
transform -1 0 4314 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_506
timestamp 1612251222
transform -1 0 4298 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_506
timestamp 1612251222
transform -1 0 4132 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_506
timestamp 1612251222
transform -1 0 4116 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_506
timestamp 1612251222
transform -1 0 4100 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_506
timestamp 1612251222
transform -1 0 4084 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_239
timestamp 1612251222
transform 1 0 3902 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_239
timestamp 1612251222
transform 1 0 3886 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_239
timestamp 1612251222
transform 1 0 3870 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_239
timestamp 1612251222
transform 1 0 3854 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_512
timestamp 1612251222
transform -1 0 3854 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_512
timestamp 1612251222
transform -1 0 3688 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_512
timestamp 1612251222
transform -1 0 3672 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_512
timestamp 1612251222
transform -1 0 3656 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_512
timestamp 1612251222
transform -1 0 3640 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_242
timestamp 1612251222
transform -1 0 3624 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_242
timestamp 1612251222
transform -1 0 3458 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_242
timestamp 1612251222
transform -1 0 3442 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_242
timestamp 1612251222
transform -1 0 3426 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_242
timestamp 1612251222
transform -1 0 3410 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_465
timestamp 1612251222
transform 1 0 3228 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_465
timestamp 1612251222
transform 1 0 3212 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_465
timestamp 1612251222
transform 1 0 3196 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_465
timestamp 1612251222
transform 1 0 3180 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_465
timestamp 1612251222
transform 1 0 3164 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_455
timestamp 1612251222
transform 1 0 2998 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_455
timestamp 1612251222
transform 1 0 2982 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_455
timestamp 1612251222
transform 1 0 2966 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_455
timestamp 1612251222
transform 1 0 2950 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_455
timestamp 1612251222
transform 1 0 2934 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_775
timestamp 1612251222
transform -1 0 2934 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_775
timestamp 1612251222
transform -1 0 2768 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_775
timestamp 1612251222
transform -1 0 2752 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_775
timestamp 1612251222
transform -1 0 2736 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_775
timestamp 1612251222
transform -1 0 2720 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_785
timestamp 1612251222
transform -1 0 2704 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_785
timestamp 1612251222
transform -1 0 2538 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_785
timestamp 1612251222
transform -1 0 2522 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_785
timestamp 1612251222
transform -1 0 2506 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_785
timestamp 1612251222
transform -1 0 2490 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_109
timestamp 1612251222
transform -1 0 2474 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_109
timestamp 1612251222
transform -1 0 2308 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_109
timestamp 1612251222
transform -1 0 2292 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_109
timestamp 1612251222
transform -1 0 2276 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_112
timestamp 1612251222
transform -1 0 2260 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_112
timestamp 1612251222
transform -1 0 2094 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_112
timestamp 1612251222
transform -1 0 2078 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_112
timestamp 1612251222
transform -1 0 2062 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_112
timestamp 1612251222
transform -1 0 2046 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_787
timestamp 1612251222
transform -1 0 2030 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_787
timestamp 1612251222
transform -1 0 1864 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_787
timestamp 1612251222
transform -1 0 1848 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_787
timestamp 1612251222
transform -1 0 1832 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_787
timestamp 1612251222
transform -1 0 1816 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_335
timestamp 1612251222
transform -1 0 1800 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_335
timestamp 1612251222
transform -1 0 1634 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_335
timestamp 1612251222
transform -1 0 1618 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_335
timestamp 1612251222
transform -1 0 1602 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_335
timestamp 1612251222
transform -1 0 1586 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_337
timestamp 1612251222
transform -1 0 1570 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_337
timestamp 1612251222
transform -1 0 1404 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_337
timestamp 1612251222
transform -1 0 1388 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_337
timestamp 1612251222
transform -1 0 1372 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_337
timestamp 1612251222
transform -1 0 1356 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_311
timestamp 1612251222
transform -1 0 1340 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_311
timestamp 1612251222
transform -1 0 1174 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_311
timestamp 1612251222
transform -1 0 1158 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_311
timestamp 1612251222
transform -1 0 1142 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_336
timestamp 1612251222
transform 1 0 960 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_336
timestamp 1612251222
transform 1 0 944 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_336
timestamp 1612251222
transform 1 0 928 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_336
timestamp 1612251222
transform 1 0 912 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_336
timestamp 1612251222
transform 1 0 896 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_295
timestamp 1612251222
transform -1 0 896 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_295
timestamp 1612251222
transform -1 0 730 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_295
timestamp 1612251222
transform -1 0 714 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_295
timestamp 1612251222
transform -1 0 698 0 -1 2210
box -4 -6 20 206
use POR2X1  POR2X1_481
timestamp 1612251222
transform -1 0 682 0 -1 2210
box -4 -6 170 206
use FILL  FILL1_POR2X1_481
timestamp 1612251222
transform -1 0 516 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_POR2X1_481
timestamp 1612251222
transform -1 0 500 0 -1 2210
box -4 -6 20 206
use FILL  FILL_POR2X1_481
timestamp 1612251222
transform -1 0 484 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_555
timestamp 1612251222
transform 1 0 302 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_555
timestamp 1612251222
transform 1 0 286 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_555
timestamp 1612251222
transform 1 0 270 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_555
timestamp 1612251222
transform 1 0 254 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_555
timestamp 1612251222
transform 1 0 238 0 -1 2210
box -4 -6 20 206
use PAND2X1  PAND2X1_345
timestamp 1612251222
transform 1 0 72 0 -1 2210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_345
timestamp 1612251222
transform 1 0 56 0 -1 2210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_345
timestamp 1612251222
transform 1 0 40 0 -1 2210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_345
timestamp 1612251222
transform 1 0 24 0 -1 2210
box -4 -6 20 206
use FILL  FILL_PAND2X1_345
timestamp 1612251222
transform 1 0 8 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_1
timestamp 1612251222
transform 1 0 10252 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_480
timestamp 1612251222
transform 1 0 10086 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_480
timestamp 1612251222
transform 1 0 10070 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_480
timestamp 1612251222
transform 1 0 10054 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_480
timestamp 1612251222
transform 1 0 10038 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_478
timestamp 1612251222
transform 1 0 9872 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_478
timestamp 1612251222
transform 1 0 9856 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_478
timestamp 1612251222
transform 1 0 9840 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_478
timestamp 1612251222
transform 1 0 9824 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_477
timestamp 1612251222
transform 1 0 9658 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_477
timestamp 1612251222
transform 1 0 9642 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_477
timestamp 1612251222
transform 1 0 9626 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_477
timestamp 1612251222
transform 1 0 9610 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_434
timestamp 1612251222
transform -1 0 9610 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_434
timestamp 1612251222
transform -1 0 9444 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_434
timestamp 1612251222
transform -1 0 9428 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_434
timestamp 1612251222
transform -1 0 9412 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_431
timestamp 1612251222
transform 1 0 9230 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_431
timestamp 1612251222
transform 1 0 9214 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_431
timestamp 1612251222
transform 1 0 9198 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_431
timestamp 1612251222
transform 1 0 9182 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_431
timestamp 1612251222
transform 1 0 9166 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_652
timestamp 1612251222
transform -1 0 9166 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_652
timestamp 1612251222
transform -1 0 9000 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_652
timestamp 1612251222
transform -1 0 8984 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_652
timestamp 1612251222
transform -1 0 8968 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_799
timestamp 1612251222
transform 1 0 8786 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_799
timestamp 1612251222
transform 1 0 8770 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_799
timestamp 1612251222
transform 1 0 8754 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_799
timestamp 1612251222
transform 1 0 8738 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_424
timestamp 1612251222
transform 1 0 8572 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_424
timestamp 1612251222
transform 1 0 8556 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_424
timestamp 1612251222
transform 1 0 8540 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_424
timestamp 1612251222
transform 1 0 8524 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_424
timestamp 1612251222
transform 1 0 8508 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_142
timestamp 1612251222
transform 1 0 8342 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_142
timestamp 1612251222
transform 1 0 8326 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_142
timestamp 1612251222
transform 1 0 8310 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_142
timestamp 1612251222
transform 1 0 8294 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_142
timestamp 1612251222
transform 1 0 8278 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_423
timestamp 1612251222
transform 1 0 8112 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_423
timestamp 1612251222
transform 1 0 8096 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_423
timestamp 1612251222
transform 1 0 8080 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_423
timestamp 1612251222
transform 1 0 8064 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_423
timestamp 1612251222
transform 1 0 8048 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_433
timestamp 1612251222
transform 1 0 7882 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_433
timestamp 1612251222
transform 1 0 7866 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_433
timestamp 1612251222
transform 1 0 7850 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_433
timestamp 1612251222
transform 1 0 7834 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_433
timestamp 1612251222
transform 1 0 7818 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_590
timestamp 1612251222
transform 1 0 7652 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_590
timestamp 1612251222
transform 1 0 7636 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_590
timestamp 1612251222
transform 1 0 7620 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_590
timestamp 1612251222
transform 1 0 7604 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_807
timestamp 1612251222
transform 1 0 7438 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_807
timestamp 1612251222
transform 1 0 7422 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_807
timestamp 1612251222
transform 1 0 7406 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_807
timestamp 1612251222
transform 1 0 7390 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_646
timestamp 1612251222
transform 1 0 7224 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_646
timestamp 1612251222
transform 1 0 7208 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_646
timestamp 1612251222
transform 1 0 7192 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_646
timestamp 1612251222
transform 1 0 7176 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_609
timestamp 1612251222
transform 1 0 7010 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_609
timestamp 1612251222
transform 1 0 6994 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_609
timestamp 1612251222
transform 1 0 6978 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_609
timestamp 1612251222
transform 1 0 6962 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_609
timestamp 1612251222
transform 1 0 6946 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_120
timestamp 1612251222
transform 1 0 6780 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_120
timestamp 1612251222
transform 1 0 6764 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_120
timestamp 1612251222
transform 1 0 6748 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_120
timestamp 1612251222
transform 1 0 6732 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_758
timestamp 1612251222
transform -1 0 6732 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_758
timestamp 1612251222
transform -1 0 6566 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_758
timestamp 1612251222
transform -1 0 6550 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_758
timestamp 1612251222
transform -1 0 6534 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_759
timestamp 1612251222
transform -1 0 6518 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_759
timestamp 1612251222
transform -1 0 6352 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_759
timestamp 1612251222
transform -1 0 6336 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_759
timestamp 1612251222
transform -1 0 6320 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_759
timestamp 1612251222
transform -1 0 6304 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_792
timestamp 1612251222
transform -1 0 6288 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_792
timestamp 1612251222
transform -1 0 6122 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_792
timestamp 1612251222
transform -1 0 6106 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_792
timestamp 1612251222
transform -1 0 6090 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_805
timestamp 1612251222
transform 1 0 5908 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_805
timestamp 1612251222
transform 1 0 5892 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_805
timestamp 1612251222
transform 1 0 5876 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_805
timestamp 1612251222
transform 1 0 5860 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_700
timestamp 1612251222
transform 1 0 5694 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_700
timestamp 1612251222
transform 1 0 5678 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_700
timestamp 1612251222
transform 1 0 5662 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_700
timestamp 1612251222
transform 1 0 5646 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_700
timestamp 1612251222
transform 1 0 5630 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_378
timestamp 1612251222
transform 1 0 5464 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_378
timestamp 1612251222
transform 1 0 5448 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_378
timestamp 1612251222
transform 1 0 5432 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_378
timestamp 1612251222
transform 1 0 5416 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_378
timestamp 1612251222
transform 1 0 5400 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_377
timestamp 1612251222
transform 1 0 5234 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_377
timestamp 1612251222
transform 1 0 5218 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_377
timestamp 1612251222
transform 1 0 5202 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_377
timestamp 1612251222
transform 1 0 5186 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_377
timestamp 1612251222
transform 1 0 5170 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_584
timestamp 1612251222
transform 1 0 5004 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_584
timestamp 1612251222
transform 1 0 4988 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_584
timestamp 1612251222
transform 1 0 4972 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_584
timestamp 1612251222
transform 1 0 4956 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_583
timestamp 1612251222
transform 1 0 4790 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_583
timestamp 1612251222
transform 1 0 4774 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_583
timestamp 1612251222
transform 1 0 4758 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_583
timestamp 1612251222
transform 1 0 4742 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_448
timestamp 1612251222
transform -1 0 4742 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_448
timestamp 1612251222
transform -1 0 4576 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_448
timestamp 1612251222
transform -1 0 4560 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_448
timestamp 1612251222
transform -1 0 4544 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_448
timestamp 1612251222
transform -1 0 4528 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_419
timestamp 1612251222
transform -1 0 4512 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_419
timestamp 1612251222
transform -1 0 4346 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_419
timestamp 1612251222
transform -1 0 4330 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_419
timestamp 1612251222
transform -1 0 4314 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_528
timestamp 1612251222
transform -1 0 4298 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_528
timestamp 1612251222
transform -1 0 4132 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_528
timestamp 1612251222
transform -1 0 4116 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_528
timestamp 1612251222
transform -1 0 4100 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_307
timestamp 1612251222
transform -1 0 4084 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_307
timestamp 1612251222
transform -1 0 3918 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_307
timestamp 1612251222
transform -1 0 3902 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_307
timestamp 1612251222
transform -1 0 3886 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_307
timestamp 1612251222
transform -1 0 3870 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_308
timestamp 1612251222
transform -1 0 3854 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_308
timestamp 1612251222
transform -1 0 3688 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_308
timestamp 1612251222
transform -1 0 3672 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_308
timestamp 1612251222
transform -1 0 3656 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_308
timestamp 1612251222
transform -1 0 3640 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_453
timestamp 1612251222
transform -1 0 3624 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_453
timestamp 1612251222
transform -1 0 3458 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_453
timestamp 1612251222
transform -1 0 3442 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_453
timestamp 1612251222
transform -1 0 3426 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_453
timestamp 1612251222
transform -1 0 3410 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_471
timestamp 1612251222
transform -1 0 3394 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_471
timestamp 1612251222
transform -1 0 3228 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_471
timestamp 1612251222
transform -1 0 3212 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_471
timestamp 1612251222
transform -1 0 3196 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_471
timestamp 1612251222
transform -1 0 3180 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_464
timestamp 1612251222
transform 1 0 2998 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_464
timestamp 1612251222
transform 1 0 2982 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_464
timestamp 1612251222
transform 1 0 2966 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_464
timestamp 1612251222
transform 1 0 2950 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_464
timestamp 1612251222
transform 1 0 2934 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_457
timestamp 1612251222
transform 1 0 2768 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_457
timestamp 1612251222
transform 1 0 2752 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_457
timestamp 1612251222
transform 1 0 2736 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_457
timestamp 1612251222
transform 1 0 2720 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_457
timestamp 1612251222
transform 1 0 2704 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_318
timestamp 1612251222
transform -1 0 2704 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_318
timestamp 1612251222
transform -1 0 2538 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_318
timestamp 1612251222
transform -1 0 2522 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_318
timestamp 1612251222
transform -1 0 2506 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_318
timestamp 1612251222
transform -1 0 2490 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_298
timestamp 1612251222
transform 1 0 2308 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_298
timestamp 1612251222
transform 1 0 2292 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_298
timestamp 1612251222
transform 1 0 2276 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_298
timestamp 1612251222
transform 1 0 2260 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_151
timestamp 1612251222
transform -1 0 2260 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_151
timestamp 1612251222
transform -1 0 2094 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_151
timestamp 1612251222
transform -1 0 2078 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_151
timestamp 1612251222
transform -1 0 2062 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_151
timestamp 1612251222
transform -1 0 2046 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_357
timestamp 1612251222
transform 1 0 1864 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_357
timestamp 1612251222
transform 1 0 1848 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_357
timestamp 1612251222
transform 1 0 1832 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_357
timestamp 1612251222
transform 1 0 1816 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_357
timestamp 1612251222
transform 1 0 1800 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_211
timestamp 1612251222
transform -1 0 1800 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_211
timestamp 1612251222
transform -1 0 1634 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_211
timestamp 1612251222
transform -1 0 1618 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_211
timestamp 1612251222
transform -1 0 1602 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_211
timestamp 1612251222
transform -1 0 1586 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_352
timestamp 1612251222
transform 1 0 1404 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_352
timestamp 1612251222
transform 1 0 1388 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_352
timestamp 1612251222
transform 1 0 1372 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_352
timestamp 1612251222
transform 1 0 1356 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_352
timestamp 1612251222
transform 1 0 1340 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_212
timestamp 1612251222
transform -1 0 1340 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_212
timestamp 1612251222
transform -1 0 1174 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_212
timestamp 1612251222
transform -1 0 1158 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_212
timestamp 1612251222
transform -1 0 1142 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_212
timestamp 1612251222
transform -1 0 1126 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_182
timestamp 1612251222
transform 1 0 944 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_182
timestamp 1612251222
transform 1 0 928 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_182
timestamp 1612251222
transform 1 0 912 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_182
timestamp 1612251222
transform 1 0 896 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_182
timestamp 1612251222
transform 1 0 880 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_312
timestamp 1612251222
transform -1 0 880 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_312
timestamp 1612251222
transform -1 0 714 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_312
timestamp 1612251222
transform -1 0 698 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_312
timestamp 1612251222
transform -1 0 682 0 1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_319
timestamp 1612251222
transform -1 0 666 0 1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_319
timestamp 1612251222
transform -1 0 500 0 1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_319
timestamp 1612251222
transform -1 0 484 0 1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_319
timestamp 1612251222
transform -1 0 468 0 1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_319
timestamp 1612251222
transform -1 0 452 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_279
timestamp 1612251222
transform 1 0 270 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_279
timestamp 1612251222
transform 1 0 254 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_279
timestamp 1612251222
transform 1 0 238 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_279
timestamp 1612251222
transform 1 0 222 0 1 1810
box -4 -6 20 206
use POR2X1  POR2X1_257
timestamp 1612251222
transform -1 0 222 0 1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_257
timestamp 1612251222
transform -1 0 56 0 1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_257
timestamp 1612251222
transform -1 0 40 0 1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_257
timestamp 1612251222
transform -1 0 24 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_2
timestamp 1612251222
transform -1 0 10268 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_1
timestamp 1612251222
transform -1 0 10252 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_469
timestamp 1612251222
transform 1 0 10070 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_469
timestamp 1612251222
transform 1 0 10054 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_469
timestamp 1612251222
transform 1 0 10038 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_469
timestamp 1612251222
transform 1 0 10022 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_468
timestamp 1612251222
transform 1 0 9856 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_468
timestamp 1612251222
transform 1 0 9840 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_468
timestamp 1612251222
transform 1 0 9824 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_468
timestamp 1612251222
transform 1 0 9808 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_470
timestamp 1612251222
transform 1 0 9642 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_470
timestamp 1612251222
transform 1 0 9626 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_470
timestamp 1612251222
transform 1 0 9610 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_470
timestamp 1612251222
transform 1 0 9594 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_466
timestamp 1612251222
transform 1 0 9428 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_466
timestamp 1612251222
transform 1 0 9412 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_466
timestamp 1612251222
transform 1 0 9396 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_466
timestamp 1612251222
transform 1 0 9380 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_453
timestamp 1612251222
transform 1 0 9214 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_453
timestamp 1612251222
transform 1 0 9198 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_453
timestamp 1612251222
transform 1 0 9182 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_453
timestamp 1612251222
transform 1 0 9166 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_449
timestamp 1612251222
transform 1 0 9000 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_449
timestamp 1612251222
transform 1 0 8984 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_449
timestamp 1612251222
transform 1 0 8968 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_449
timestamp 1612251222
transform 1 0 8952 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_593
timestamp 1612251222
transform 1 0 8786 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_593
timestamp 1612251222
transform 1 0 8770 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_593
timestamp 1612251222
transform 1 0 8754 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_593
timestamp 1612251222
transform 1 0 8738 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_592
timestamp 1612251222
transform 1 0 8572 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_592
timestamp 1612251222
transform 1 0 8556 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_592
timestamp 1612251222
transform 1 0 8540 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_592
timestamp 1612251222
transform 1 0 8524 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_589
timestamp 1612251222
transform 1 0 8358 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_589
timestamp 1612251222
transform 1 0 8342 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_589
timestamp 1612251222
transform 1 0 8326 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_589
timestamp 1612251222
transform 1 0 8310 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_589
timestamp 1612251222
transform 1 0 8294 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_56
timestamp 1612251222
transform 1 0 8128 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_56
timestamp 1612251222
transform 1 0 8112 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_56
timestamp 1612251222
transform 1 0 8096 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_56
timestamp 1612251222
transform 1 0 8080 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_56
timestamp 1612251222
transform 1 0 8064 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_591
timestamp 1612251222
transform 1 0 7898 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_591
timestamp 1612251222
transform 1 0 7882 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_591
timestamp 1612251222
transform 1 0 7866 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_591
timestamp 1612251222
transform 1 0 7850 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_591
timestamp 1612251222
transform 1 0 7834 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_304
timestamp 1612251222
transform -1 0 7834 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_304
timestamp 1612251222
transform -1 0 7668 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_304
timestamp 1612251222
transform -1 0 7652 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_304
timestamp 1612251222
transform -1 0 7636 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_304
timestamp 1612251222
transform -1 0 7620 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_511
timestamp 1612251222
transform 1 0 7438 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_511
timestamp 1612251222
transform 1 0 7422 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_511
timestamp 1612251222
transform 1 0 7406 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_511
timestamp 1612251222
transform 1 0 7390 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_511
timestamp 1612251222
transform 1 0 7374 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_606
timestamp 1612251222
transform -1 0 7374 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_606
timestamp 1612251222
transform -1 0 7208 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_606
timestamp 1612251222
transform -1 0 7192 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_606
timestamp 1612251222
transform -1 0 7176 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_607
timestamp 1612251222
transform 1 0 6994 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_607
timestamp 1612251222
transform 1 0 6978 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_607
timestamp 1612251222
transform 1 0 6962 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_607
timestamp 1612251222
transform 1 0 6946 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_607
timestamp 1612251222
transform 1 0 6930 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_608
timestamp 1612251222
transform 1 0 6764 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_608
timestamp 1612251222
transform 1 0 6748 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_608
timestamp 1612251222
transform 1 0 6732 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_608
timestamp 1612251222
transform 1 0 6716 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_585
timestamp 1612251222
transform -1 0 6716 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_585
timestamp 1612251222
transform -1 0 6550 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_585
timestamp 1612251222
transform -1 0 6534 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_585
timestamp 1612251222
transform -1 0 6518 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_585
timestamp 1612251222
transform -1 0 6502 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_791
timestamp 1612251222
transform -1 0 6486 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_791
timestamp 1612251222
transform -1 0 6320 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_791
timestamp 1612251222
transform -1 0 6304 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_791
timestamp 1612251222
transform -1 0 6288 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_757
timestamp 1612251222
transform 1 0 6106 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_757
timestamp 1612251222
transform 1 0 6090 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_757
timestamp 1612251222
transform 1 0 6074 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_757
timestamp 1612251222
transform 1 0 6058 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_757
timestamp 1612251222
transform 1 0 6042 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_756
timestamp 1612251222
transform 1 0 5876 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_756
timestamp 1612251222
transform 1 0 5860 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_756
timestamp 1612251222
transform 1 0 5844 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_756
timestamp 1612251222
transform 1 0 5828 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_463
timestamp 1612251222
transform 1 0 5662 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_463
timestamp 1612251222
transform 1 0 5646 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_463
timestamp 1612251222
transform 1 0 5630 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_463
timestamp 1612251222
transform 1 0 5614 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_459
timestamp 1612251222
transform 1 0 5448 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_459
timestamp 1612251222
transform 1 0 5432 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_459
timestamp 1612251222
transform 1 0 5416 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_459
timestamp 1612251222
transform 1 0 5400 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_376
timestamp 1612251222
transform 1 0 5234 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_376
timestamp 1612251222
transform 1 0 5218 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_376
timestamp 1612251222
transform 1 0 5202 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_376
timestamp 1612251222
transform 1 0 5186 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_376
timestamp 1612251222
transform 1 0 5170 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_636
timestamp 1612251222
transform -1 0 5170 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_636
timestamp 1612251222
transform -1 0 5004 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_636
timestamp 1612251222
transform -1 0 4988 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_636
timestamp 1612251222
transform -1 0 4972 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_636
timestamp 1612251222
transform -1 0 4956 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_639
timestamp 1612251222
transform 1 0 4774 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_639
timestamp 1612251222
transform 1 0 4758 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_639
timestamp 1612251222
transform 1 0 4742 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_639
timestamp 1612251222
transform 1 0 4726 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_639
timestamp 1612251222
transform 1 0 4710 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_421
timestamp 1612251222
transform 1 0 4544 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_421
timestamp 1612251222
transform 1 0 4528 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_421
timestamp 1612251222
transform 1 0 4512 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_421
timestamp 1612251222
transform 1 0 4496 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_420
timestamp 1612251222
transform -1 0 4496 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_420
timestamp 1612251222
transform -1 0 4330 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_420
timestamp 1612251222
transform -1 0 4314 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_420
timestamp 1612251222
transform -1 0 4298 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_447
timestamp 1612251222
transform -1 0 4282 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_447
timestamp 1612251222
transform -1 0 4116 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_447
timestamp 1612251222
transform -1 0 4100 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_447
timestamp 1612251222
transform -1 0 4084 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_447
timestamp 1612251222
transform -1 0 4068 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_304
timestamp 1612251222
transform 1 0 3886 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_304
timestamp 1612251222
transform 1 0 3870 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_304
timestamp 1612251222
transform 1 0 3854 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_304
timestamp 1612251222
transform 1 0 3838 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_306
timestamp 1612251222
transform 1 0 3672 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_306
timestamp 1612251222
transform 1 0 3656 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_306
timestamp 1612251222
transform 1 0 3640 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_306
timestamp 1612251222
transform 1 0 3624 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_449
timestamp 1612251222
transform 1 0 3458 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_449
timestamp 1612251222
transform 1 0 3442 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_449
timestamp 1612251222
transform 1 0 3426 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_449
timestamp 1612251222
transform 1 0 3410 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_449
timestamp 1612251222
transform 1 0 3394 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_237
timestamp 1612251222
transform -1 0 3394 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_237
timestamp 1612251222
transform -1 0 3228 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_237
timestamp 1612251222
transform -1 0 3212 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_237
timestamp 1612251222
transform -1 0 3196 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_241
timestamp 1612251222
transform 1 0 3014 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_241
timestamp 1612251222
transform 1 0 2998 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_241
timestamp 1612251222
transform 1 0 2982 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_241
timestamp 1612251222
transform 1 0 2966 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_241
timestamp 1612251222
transform 1 0 2950 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_445
timestamp 1612251222
transform 1 0 2784 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_445
timestamp 1612251222
transform 1 0 2768 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_445
timestamp 1612251222
transform 1 0 2752 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_445
timestamp 1612251222
transform 1 0 2736 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_445
timestamp 1612251222
transform 1 0 2720 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_299
timestamp 1612251222
transform -1 0 2720 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_299
timestamp 1612251222
transform -1 0 2554 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_299
timestamp 1612251222
transform -1 0 2538 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_299
timestamp 1612251222
transform -1 0 2522 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_302
timestamp 1612251222
transform -1 0 2506 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_302
timestamp 1612251222
transform -1 0 2340 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_302
timestamp 1612251222
transform -1 0 2324 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_302
timestamp 1612251222
transform -1 0 2308 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_302
timestamp 1612251222
transform -1 0 2292 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_303
timestamp 1612251222
transform -1 0 2276 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_303
timestamp 1612251222
transform -1 0 2110 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_303
timestamp 1612251222
transform -1 0 2094 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_303
timestamp 1612251222
transform -1 0 2078 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_303
timestamp 1612251222
transform -1 0 2062 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_353
timestamp 1612251222
transform -1 0 2046 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_353
timestamp 1612251222
transform -1 0 1880 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_353
timestamp 1612251222
transform -1 0 1864 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_353
timestamp 1612251222
transform -1 0 1848 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_353
timestamp 1612251222
transform -1 0 1832 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_566
timestamp 1612251222
transform -1 0 1816 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_566
timestamp 1612251222
transform -1 0 1650 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_566
timestamp 1612251222
transform -1 0 1634 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_566
timestamp 1612251222
transform -1 0 1618 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_566
timestamp 1612251222
transform -1 0 1602 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_370
timestamp 1612251222
transform 1 0 1420 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_370
timestamp 1612251222
transform 1 0 1404 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_370
timestamp 1612251222
transform 1 0 1388 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_370
timestamp 1612251222
transform 1 0 1372 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_370
timestamp 1612251222
transform 1 0 1356 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_220
timestamp 1612251222
transform 1 0 1190 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_220
timestamp 1612251222
transform 1 0 1174 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_220
timestamp 1612251222
transform 1 0 1158 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_220
timestamp 1612251222
transform 1 0 1142 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_220
timestamp 1612251222
transform 1 0 1126 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_180
timestamp 1612251222
transform 1 0 960 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_180
timestamp 1612251222
transform 1 0 944 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_180
timestamp 1612251222
transform 1 0 928 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_180
timestamp 1612251222
transform 1 0 912 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_180
timestamp 1612251222
transform 1 0 896 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_176
timestamp 1612251222
transform 1 0 730 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_176
timestamp 1612251222
transform 1 0 714 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_176
timestamp 1612251222
transform 1 0 698 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_176
timestamp 1612251222
transform 1 0 682 0 -1 1810
box -4 -6 20 206
use POR2X1  POR2X1_258
timestamp 1612251222
transform -1 0 682 0 -1 1810
box -4 -6 170 206
use FILL  FILL1_POR2X1_258
timestamp 1612251222
transform -1 0 516 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_POR2X1_258
timestamp 1612251222
transform -1 0 500 0 -1 1810
box -4 -6 20 206
use FILL  FILL_POR2X1_258
timestamp 1612251222
transform -1 0 484 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_284
timestamp 1612251222
transform -1 0 468 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_284
timestamp 1612251222
transform -1 0 302 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_284
timestamp 1612251222
transform -1 0 286 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_284
timestamp 1612251222
transform -1 0 270 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_284
timestamp 1612251222
transform -1 0 254 0 -1 1810
box -4 -6 20 206
use PAND2X1  PAND2X1_259
timestamp 1612251222
transform 1 0 72 0 -1 1810
box -4 -6 170 206
use FILL  FILL2_PAND2X1_259
timestamp 1612251222
transform 1 0 56 0 -1 1810
box -4 -6 20 206
use FILL  FILL1_PAND2X1_259
timestamp 1612251222
transform 1 0 40 0 -1 1810
box -4 -6 20 206
use FILL  FILL0_PAND2X1_259
timestamp 1612251222
transform 1 0 24 0 -1 1810
box -4 -6 20 206
use FILL  FILL_PAND2X1_259
timestamp 1612251222
transform 1 0 8 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_4
timestamp 1612251222
transform 1 0 10252 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_3
timestamp 1612251222
transform 1 0 10236 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_2
timestamp 1612251222
transform 1 0 10220 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_1
timestamp 1612251222
transform 1 0 10204 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_354
timestamp 1612251222
transform 1 0 10038 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_354
timestamp 1612251222
transform 1 0 10022 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_354
timestamp 1612251222
transform 1 0 10006 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_354
timestamp 1612251222
transform 1 0 9990 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_326
timestamp 1612251222
transform 1 0 9824 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_326
timestamp 1612251222
transform 1 0 9808 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_326
timestamp 1612251222
transform 1 0 9792 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_326
timestamp 1612251222
transform 1 0 9776 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_798
timestamp 1612251222
transform -1 0 9776 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_798
timestamp 1612251222
transform -1 0 9610 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_798
timestamp 1612251222
transform -1 0 9594 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_798
timestamp 1612251222
transform -1 0 9578 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_436
timestamp 1612251222
transform 1 0 9396 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_436
timestamp 1612251222
transform 1 0 9380 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_436
timestamp 1612251222
transform 1 0 9364 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_436
timestamp 1612251222
transform 1 0 9348 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_532
timestamp 1612251222
transform -1 0 9348 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_532
timestamp 1612251222
transform -1 0 9182 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_532
timestamp 1612251222
transform -1 0 9166 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_532
timestamp 1612251222
transform -1 0 9150 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_533
timestamp 1612251222
transform 1 0 8968 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_533
timestamp 1612251222
transform 1 0 8952 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_533
timestamp 1612251222
transform 1 0 8936 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_533
timestamp 1612251222
transform 1 0 8920 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_533
timestamp 1612251222
transform 1 0 8904 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_802
timestamp 1612251222
transform -1 0 8904 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_802
timestamp 1612251222
transform -1 0 8738 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_802
timestamp 1612251222
transform -1 0 8722 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_802
timestamp 1612251222
transform -1 0 8706 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_147
timestamp 1612251222
transform 1 0 8524 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_147
timestamp 1612251222
transform 1 0 8508 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_147
timestamp 1612251222
transform 1 0 8492 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_147
timestamp 1612251222
transform 1 0 8476 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_794
timestamp 1612251222
transform -1 0 8476 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_794
timestamp 1612251222
transform -1 0 8310 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_794
timestamp 1612251222
transform -1 0 8294 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_794
timestamp 1612251222
transform -1 0 8278 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_804
timestamp 1612251222
transform -1 0 8262 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_804
timestamp 1612251222
transform -1 0 8096 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_804
timestamp 1612251222
transform -1 0 8080 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_804
timestamp 1612251222
transform -1 0 8064 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_718
timestamp 1612251222
transform -1 0 8048 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_718
timestamp 1612251222
transform -1 0 7882 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_718
timestamp 1612251222
transform -1 0 7866 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_718
timestamp 1612251222
transform -1 0 7850 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_435
timestamp 1612251222
transform 1 0 7668 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_435
timestamp 1612251222
transform 1 0 7652 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_435
timestamp 1612251222
transform 1 0 7636 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_435
timestamp 1612251222
transform 1 0 7620 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_432
timestamp 1612251222
transform 1 0 7454 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_432
timestamp 1612251222
transform 1 0 7438 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_432
timestamp 1612251222
transform 1 0 7422 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_432
timestamp 1612251222
transform 1 0 7406 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_432
timestamp 1612251222
transform 1 0 7390 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_600
timestamp 1612251222
transform 1 0 7224 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_600
timestamp 1612251222
transform 1 0 7208 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_600
timestamp 1612251222
transform 1 0 7192 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_600
timestamp 1612251222
transform 1 0 7176 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_600
timestamp 1612251222
transform 1 0 7160 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_666
timestamp 1612251222
transform 1 0 6994 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_666
timestamp 1612251222
transform 1 0 6978 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_666
timestamp 1612251222
transform 1 0 6962 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_666
timestamp 1612251222
transform 1 0 6946 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_666
timestamp 1612251222
transform 1 0 6930 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_664
timestamp 1612251222
transform 1 0 6764 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_664
timestamp 1612251222
transform 1 0 6748 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_664
timestamp 1612251222
transform 1 0 6732 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_664
timestamp 1612251222
transform 1 0 6716 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_755
timestamp 1612251222
transform -1 0 6716 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_755
timestamp 1612251222
transform -1 0 6550 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_755
timestamp 1612251222
transform -1 0 6534 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_755
timestamp 1612251222
transform -1 0 6518 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_755
timestamp 1612251222
transform -1 0 6502 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_586
timestamp 1612251222
transform -1 0 6486 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_586
timestamp 1612251222
transform -1 0 6320 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_586
timestamp 1612251222
transform -1 0 6304 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_586
timestamp 1612251222
transform -1 0 6288 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_586
timestamp 1612251222
transform -1 0 6272 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_637
timestamp 1612251222
transform -1 0 6256 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_637
timestamp 1612251222
transform -1 0 6090 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_637
timestamp 1612251222
transform -1 0 6074 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_637
timestamp 1612251222
transform -1 0 6058 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_95
timestamp 1612251222
transform 1 0 5876 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_95
timestamp 1612251222
transform 1 0 5860 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_95
timestamp 1612251222
transform 1 0 5844 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_95
timestamp 1612251222
transform 1 0 5828 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_95
timestamp 1612251222
transform 1 0 5812 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_379
timestamp 1612251222
transform -1 0 5812 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_379
timestamp 1612251222
transform -1 0 5646 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_379
timestamp 1612251222
transform -1 0 5630 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_379
timestamp 1612251222
transform -1 0 5614 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_380
timestamp 1612251222
transform -1 0 5598 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_380
timestamp 1612251222
transform -1 0 5432 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_380
timestamp 1612251222
transform -1 0 5416 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_380
timestamp 1612251222
transform -1 0 5400 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_380
timestamp 1612251222
transform -1 0 5384 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_460
timestamp 1612251222
transform -1 0 5368 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_460
timestamp 1612251222
transform -1 0 5202 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_460
timestamp 1612251222
transform -1 0 5186 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_460
timestamp 1612251222
transform -1 0 5170 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_375
timestamp 1612251222
transform 1 0 4988 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_375
timestamp 1612251222
transform 1 0 4972 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_375
timestamp 1612251222
transform 1 0 4956 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_375
timestamp 1612251222
transform 1 0 4940 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_588
timestamp 1612251222
transform 1 0 4774 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_588
timestamp 1612251222
transform 1 0 4758 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_588
timestamp 1612251222
transform 1 0 4742 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_588
timestamp 1612251222
transform 1 0 4726 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_386
timestamp 1612251222
transform 1 0 4560 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_386
timestamp 1612251222
transform 1 0 4544 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_386
timestamp 1612251222
transform 1 0 4528 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_386
timestamp 1612251222
transform 1 0 4512 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_699
timestamp 1612251222
transform -1 0 4512 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_699
timestamp 1612251222
transform -1 0 4346 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_699
timestamp 1612251222
transform -1 0 4330 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_699
timestamp 1612251222
transform -1 0 4314 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_155
timestamp 1612251222
transform 1 0 4132 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_155
timestamp 1612251222
transform 1 0 4116 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_155
timestamp 1612251222
transform 1 0 4100 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_155
timestamp 1612251222
transform 1 0 4084 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_155
timestamp 1612251222
transform 1 0 4068 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_743
timestamp 1612251222
transform 1 0 3902 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_743
timestamp 1612251222
transform 1 0 3886 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_743
timestamp 1612251222
transform 1 0 3870 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_743
timestamp 1612251222
transform 1 0 3854 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_796
timestamp 1612251222
transform -1 0 3854 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_796
timestamp 1612251222
transform -1 0 3688 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_796
timestamp 1612251222
transform -1 0 3672 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_796
timestamp 1612251222
transform -1 0 3656 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_796
timestamp 1612251222
transform -1 0 3640 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_454
timestamp 1612251222
transform -1 0 3624 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_454
timestamp 1612251222
transform -1 0 3458 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_454
timestamp 1612251222
transform -1 0 3442 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_454
timestamp 1612251222
transform -1 0 3426 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_454
timestamp 1612251222
transform -1 0 3410 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_466
timestamp 1612251222
transform -1 0 3394 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_466
timestamp 1612251222
transform -1 0 3228 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_466
timestamp 1612251222
transform -1 0 3212 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_466
timestamp 1612251222
transform -1 0 3196 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_466
timestamp 1612251222
transform -1 0 3180 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_470
timestamp 1612251222
transform -1 0 3164 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_470
timestamp 1612251222
transform -1 0 2998 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_470
timestamp 1612251222
transform -1 0 2982 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_470
timestamp 1612251222
transform -1 0 2966 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_470
timestamp 1612251222
transform -1 0 2950 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_477
timestamp 1612251222
transform -1 0 2934 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_477
timestamp 1612251222
transform -1 0 2768 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_477
timestamp 1612251222
transform -1 0 2752 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_477
timestamp 1612251222
transform -1 0 2736 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_477
timestamp 1612251222
transform -1 0 2720 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_480
timestamp 1612251222
transform 1 0 2538 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_480
timestamp 1612251222
transform 1 0 2522 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_480
timestamp 1612251222
transform 1 0 2506 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_480
timestamp 1612251222
transform 1 0 2490 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_480
timestamp 1612251222
transform 1 0 2474 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_478
timestamp 1612251222
transform 1 0 2308 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_478
timestamp 1612251222
transform 1 0 2292 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_478
timestamp 1612251222
transform 1 0 2276 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_478
timestamp 1612251222
transform 1 0 2260 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_478
timestamp 1612251222
transform 1 0 2244 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_469
timestamp 1612251222
transform 1 0 2078 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_469
timestamp 1612251222
transform 1 0 2062 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_469
timestamp 1612251222
transform 1 0 2046 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_469
timestamp 1612251222
transform 1 0 2030 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_469
timestamp 1612251222
transform 1 0 2014 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_444
timestamp 1612251222
transform 1 0 1848 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_444
timestamp 1612251222
transform 1 0 1832 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_444
timestamp 1612251222
transform 1 0 1816 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_444
timestamp 1612251222
transform 1 0 1800 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_444
timestamp 1612251222
transform 1 0 1784 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_442
timestamp 1612251222
transform 1 0 1618 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_442
timestamp 1612251222
transform 1 0 1602 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_442
timestamp 1612251222
transform 1 0 1586 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_442
timestamp 1612251222
transform 1 0 1570 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_369
timestamp 1612251222
transform -1 0 1570 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_369
timestamp 1612251222
transform -1 0 1404 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_369
timestamp 1612251222
transform -1 0 1388 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_369
timestamp 1612251222
transform -1 0 1372 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_543
timestamp 1612251222
transform -1 0 1356 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_543
timestamp 1612251222
transform -1 0 1190 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_543
timestamp 1612251222
transform -1 0 1174 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_543
timestamp 1612251222
transform -1 0 1158 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_543
timestamp 1612251222
transform -1 0 1142 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_388
timestamp 1612251222
transform 1 0 960 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_388
timestamp 1612251222
transform 1 0 944 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_388
timestamp 1612251222
transform 1 0 928 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_388
timestamp 1612251222
transform 1 0 912 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_388
timestamp 1612251222
transform 1 0 896 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_177
timestamp 1612251222
transform 1 0 730 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_177
timestamp 1612251222
transform 1 0 714 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_177
timestamp 1612251222
transform 1 0 698 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_177
timestamp 1612251222
transform 1 0 682 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_703
timestamp 1612251222
transform 1 0 516 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_703
timestamp 1612251222
transform 1 0 500 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_703
timestamp 1612251222
transform 1 0 484 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_703
timestamp 1612251222
transform 1 0 468 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_703
timestamp 1612251222
transform 1 0 452 0 1 1410
box -4 -6 20 206
use POR2X1  POR2X1_280
timestamp 1612251222
transform -1 0 452 0 1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_280
timestamp 1612251222
transform -1 0 286 0 1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_280
timestamp 1612251222
transform -1 0 270 0 1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_280
timestamp 1612251222
transform -1 0 254 0 1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_542
timestamp 1612251222
transform -1 0 238 0 1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_542
timestamp 1612251222
transform -1 0 72 0 1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_542
timestamp 1612251222
transform -1 0 56 0 1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_542
timestamp 1612251222
transform -1 0 40 0 1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_542
timestamp 1612251222
transform -1 0 24 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_13
timestamp 1612251222
transform -1 0 10262 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_12
timestamp 1612251222
transform -1 0 10246 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_11
timestamp 1612251222
transform -1 0 10230 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_10
timestamp 1612251222
transform -1 0 10214 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_9
timestamp 1612251222
transform -1 0 10198 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_8
timestamp 1612251222
transform -1 0 10182 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_7
timestamp 1612251222
transform -1 0 10166 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_6
timestamp 1612251222
transform -1 0 10150 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_5
timestamp 1612251222
transform -1 0 10134 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_4
timestamp 1612251222
transform -1 0 10118 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_3
timestamp 1612251222
transform -1 0 10102 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_2
timestamp 1612251222
transform -1 0 10086 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_1
timestamp 1612251222
transform -1 0 10070 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_324
timestamp 1612251222
transform -1 0 10054 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_324
timestamp 1612251222
transform -1 0 9888 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_324
timestamp 1612251222
transform -1 0 9872 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_324
timestamp 1612251222
transform -1 0 9856 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_321
timestamp 1612251222
transform 1 0 9674 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_321
timestamp 1612251222
transform 1 0 9658 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_321
timestamp 1612251222
transform 1 0 9642 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_321
timestamp 1612251222
transform 1 0 9626 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_321
timestamp 1612251222
transform 1 0 9610 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_535
timestamp 1612251222
transform 1 0 9444 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_535
timestamp 1612251222
transform 1 0 9428 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_535
timestamp 1612251222
transform 1 0 9412 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_535
timestamp 1612251222
transform 1 0 9396 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_534
timestamp 1612251222
transform 1 0 9230 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_534
timestamp 1612251222
transform 1 0 9214 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_534
timestamp 1612251222
transform 1 0 9198 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_534
timestamp 1612251222
transform 1 0 9182 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_534
timestamp 1612251222
transform 1 0 9166 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_448
timestamp 1612251222
transform 1 0 9000 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_448
timestamp 1612251222
transform 1 0 8984 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_448
timestamp 1612251222
transform 1 0 8968 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_448
timestamp 1612251222
transform 1 0 8952 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_422
timestamp 1612251222
transform 1 0 8786 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_422
timestamp 1612251222
transform 1 0 8770 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_422
timestamp 1612251222
transform 1 0 8754 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_422
timestamp 1612251222
transform 1 0 8738 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_422
timestamp 1612251222
transform 1 0 8722 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_788
timestamp 1612251222
transform -1 0 8722 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_788
timestamp 1612251222
transform -1 0 8556 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_788
timestamp 1612251222
transform -1 0 8540 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_788
timestamp 1612251222
transform -1 0 8524 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_144
timestamp 1612251222
transform 1 0 8342 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_144
timestamp 1612251222
transform 1 0 8326 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_144
timestamp 1612251222
transform 1 0 8310 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_144
timestamp 1612251222
transform 1 0 8294 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_144
timestamp 1612251222
transform 1 0 8278 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_602
timestamp 1612251222
transform 1 0 8112 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_602
timestamp 1612251222
transform 1 0 8096 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_602
timestamp 1612251222
transform 1 0 8080 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_602
timestamp 1612251222
transform 1 0 8064 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_601
timestamp 1612251222
transform 1 0 7898 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_601
timestamp 1612251222
transform 1 0 7882 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_601
timestamp 1612251222
transform 1 0 7866 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_601
timestamp 1612251222
transform 1 0 7850 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_601
timestamp 1612251222
transform 1 0 7834 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_722
timestamp 1612251222
transform 1 0 7668 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_722
timestamp 1612251222
transform 1 0 7652 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_722
timestamp 1612251222
transform 1 0 7636 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_722
timestamp 1612251222
transform 1 0 7620 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_696
timestamp 1612251222
transform -1 0 7620 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_696
timestamp 1612251222
transform -1 0 7454 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_696
timestamp 1612251222
transform -1 0 7438 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_696
timestamp 1612251222
transform -1 0 7422 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_696
timestamp 1612251222
transform -1 0 7406 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_719
timestamp 1612251222
transform 1 0 7224 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_719
timestamp 1612251222
transform 1 0 7208 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_719
timestamp 1612251222
transform 1 0 7192 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_719
timestamp 1612251222
transform 1 0 7176 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_665
timestamp 1612251222
transform 1 0 7010 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_665
timestamp 1612251222
transform 1 0 6994 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_665
timestamp 1612251222
transform 1 0 6978 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_665
timestamp 1612251222
transform 1 0 6962 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_665
timestamp 1612251222
transform 1 0 6946 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_387
timestamp 1612251222
transform 1 0 6780 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_387
timestamp 1612251222
transform 1 0 6764 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_387
timestamp 1612251222
transform 1 0 6748 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_387
timestamp 1612251222
transform 1 0 6732 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_387
timestamp 1612251222
transform 1 0 6716 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_651
timestamp 1612251222
transform 1 0 6550 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_651
timestamp 1612251222
transform 1 0 6534 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_651
timestamp 1612251222
transform 1 0 6518 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_651
timestamp 1612251222
transform 1 0 6502 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_53
timestamp 1612251222
transform 1 0 6336 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_53
timestamp 1612251222
transform 1 0 6320 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_53
timestamp 1612251222
transform 1 0 6304 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_53
timestamp 1612251222
transform 1 0 6288 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_53
timestamp 1612251222
transform 1 0 6272 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_638
timestamp 1612251222
transform 1 0 6106 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_638
timestamp 1612251222
transform 1 0 6090 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_638
timestamp 1612251222
transform 1 0 6074 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_638
timestamp 1612251222
transform 1 0 6058 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_588
timestamp 1612251222
transform 1 0 5892 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_588
timestamp 1612251222
transform 1 0 5876 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_588
timestamp 1612251222
transform 1 0 5860 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_588
timestamp 1612251222
transform 1 0 5844 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_588
timestamp 1612251222
transform 1 0 5828 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_18
timestamp 1612251222
transform -1 0 5828 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_18
timestamp 1612251222
transform -1 0 5662 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_18
timestamp 1612251222
transform -1 0 5646 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_18
timestamp 1612251222
transform -1 0 5630 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_18
timestamp 1612251222
transform -1 0 5614 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_752
timestamp 1612251222
transform 1 0 5432 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_752
timestamp 1612251222
transform 1 0 5416 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_752
timestamp 1612251222
transform 1 0 5400 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_752
timestamp 1612251222
transform 1 0 5384 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_752
timestamp 1612251222
transform 1 0 5368 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_752
timestamp 1612251222
transform 1 0 5202 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_752
timestamp 1612251222
transform 1 0 5186 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_752
timestamp 1612251222
transform 1 0 5170 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_752
timestamp 1612251222
transform 1 0 5154 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_22
timestamp 1612251222
transform 1 0 4988 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_POR2X1_22
timestamp 1612251222
transform 1 0 4972 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_POR2X1_22
timestamp 1612251222
transform 1 0 4956 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_22
timestamp 1612251222
transform 1 0 4940 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_22
timestamp 1612251222
transform 1 0 4924 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_408
timestamp 1612251222
transform -1 0 4924 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_408
timestamp 1612251222
transform -1 0 4758 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_408
timestamp 1612251222
transform -1 0 4742 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_408
timestamp 1612251222
transform -1 0 4726 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_328
timestamp 1612251222
transform -1 0 4710 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_328
timestamp 1612251222
transform -1 0 4544 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_328
timestamp 1612251222
transform -1 0 4528 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_328
timestamp 1612251222
transform -1 0 4512 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_53
timestamp 1612251222
transform -1 0 4496 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_POR2X1_53
timestamp 1612251222
transform -1 0 4330 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_POR2X1_53
timestamp 1612251222
transform -1 0 4314 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_53
timestamp 1612251222
transform -1 0 4298 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_53
timestamp 1612251222
transform -1 0 4282 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_156
timestamp 1612251222
transform -1 0 4266 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_156
timestamp 1612251222
transform -1 0 4100 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_156
timestamp 1612251222
transform -1 0 4084 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_156
timestamp 1612251222
transform -1 0 4068 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_156
timestamp 1612251222
transform -1 0 4052 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_780
timestamp 1612251222
transform -1 0 4036 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_780
timestamp 1612251222
transform -1 0 3870 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_780
timestamp 1612251222
transform -1 0 3854 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_780
timestamp 1612251222
transform -1 0 3838 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_780
timestamp 1612251222
transform -1 0 3822 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_783
timestamp 1612251222
transform -1 0 3806 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_783
timestamp 1612251222
transform -1 0 3640 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_783
timestamp 1612251222
transform -1 0 3624 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_783
timestamp 1612251222
transform -1 0 3608 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_783
timestamp 1612251222
transform -1 0 3592 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_424
timestamp 1612251222
transform -1 0 3576 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_424
timestamp 1612251222
transform -1 0 3410 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_424
timestamp 1612251222
transform -1 0 3394 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_424
timestamp 1612251222
transform -1 0 3378 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_446
timestamp 1612251222
transform 1 0 3196 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_446
timestamp 1612251222
transform 1 0 3180 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_446
timestamp 1612251222
transform 1 0 3164 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_446
timestamp 1612251222
transform 1 0 3148 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_446
timestamp 1612251222
transform 1 0 3132 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_418
timestamp 1612251222
transform 1 0 2966 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_418
timestamp 1612251222
transform 1 0 2950 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_418
timestamp 1612251222
transform 1 0 2934 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_418
timestamp 1612251222
transform 1 0 2918 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_238
timestamp 1612251222
transform 1 0 2752 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_238
timestamp 1612251222
transform 1 0 2736 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_238
timestamp 1612251222
transform 1 0 2720 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_238
timestamp 1612251222
transform 1 0 2704 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_776
timestamp 1612251222
transform 1 0 2538 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_776
timestamp 1612251222
transform 1 0 2522 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_776
timestamp 1612251222
transform 1 0 2506 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_776
timestamp 1612251222
transform 1 0 2490 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_776
timestamp 1612251222
transform 1 0 2474 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_91
timestamp 1612251222
transform -1 0 2474 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_91
timestamp 1612251222
transform -1 0 2308 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_91
timestamp 1612251222
transform -1 0 2292 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_91
timestamp 1612251222
transform -1 0 2276 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_315
timestamp 1612251222
transform 1 0 2094 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_315
timestamp 1612251222
transform 1 0 2078 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_315
timestamp 1612251222
transform 1 0 2062 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_315
timestamp 1612251222
transform 1 0 2046 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_727
timestamp 1612251222
transform -1 0 2046 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_727
timestamp 1612251222
transform -1 0 1880 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_727
timestamp 1612251222
transform -1 0 1864 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_727
timestamp 1612251222
transform -1 0 1848 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_727
timestamp 1612251222
transform -1 0 1832 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_443
timestamp 1612251222
transform 1 0 1650 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_443
timestamp 1612251222
transform 1 0 1634 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_443
timestamp 1612251222
transform 1 0 1618 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_443
timestamp 1612251222
transform 1 0 1602 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_443
timestamp 1612251222
transform 1 0 1586 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_803
timestamp 1612251222
transform -1 0 1586 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_803
timestamp 1612251222
transform -1 0 1420 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_803
timestamp 1612251222
transform -1 0 1404 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_803
timestamp 1612251222
transform -1 0 1388 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_803
timestamp 1612251222
transform -1 0 1372 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_704
timestamp 1612251222
transform 1 0 1190 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_704
timestamp 1612251222
transform 1 0 1174 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_704
timestamp 1612251222
transform 1 0 1158 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_704
timestamp 1612251222
transform 1 0 1142 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_704
timestamp 1612251222
transform 1 0 1126 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_439
timestamp 1612251222
transform 1 0 960 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_439
timestamp 1612251222
transform 1 0 944 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_439
timestamp 1612251222
transform 1 0 928 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_439
timestamp 1612251222
transform 1 0 912 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_439
timestamp 1612251222
transform 1 0 896 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_313
timestamp 1612251222
transform -1 0 896 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_313
timestamp 1612251222
transform -1 0 730 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_313
timestamp 1612251222
transform -1 0 714 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_313
timestamp 1612251222
transform -1 0 698 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_317
timestamp 1612251222
transform 1 0 516 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_317
timestamp 1612251222
transform 1 0 500 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_317
timestamp 1612251222
transform 1 0 484 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_317
timestamp 1612251222
transform 1 0 468 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_317
timestamp 1612251222
transform 1 0 452 0 -1 1410
box -4 -6 20 206
use POR2X1  POR2X1_314
timestamp 1612251222
transform 1 0 286 0 -1 1410
box -4 -6 170 206
use FILL  FILL1_POR2X1_314
timestamp 1612251222
transform 1 0 270 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_POR2X1_314
timestamp 1612251222
transform 1 0 254 0 -1 1410
box -4 -6 20 206
use FILL  FILL_POR2X1_314
timestamp 1612251222
transform 1 0 238 0 -1 1410
box -4 -6 20 206
use PAND2X1  PAND2X1_552
timestamp 1612251222
transform 1 0 72 0 -1 1410
box -4 -6 170 206
use FILL  FILL2_PAND2X1_552
timestamp 1612251222
transform 1 0 56 0 -1 1410
box -4 -6 20 206
use FILL  FILL1_PAND2X1_552
timestamp 1612251222
transform 1 0 40 0 -1 1410
box -4 -6 20 206
use FILL  FILL0_PAND2X1_552
timestamp 1612251222
transform 1 0 24 0 -1 1410
box -4 -6 20 206
use FILL  FILL_PAND2X1_552
timestamp 1612251222
transform 1 0 8 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_12
timestamp 1612251222
transform 1 0 10246 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_11
timestamp 1612251222
transform 1 0 10230 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_10
timestamp 1612251222
transform 1 0 10214 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_9
timestamp 1612251222
transform 1 0 10198 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_8
timestamp 1612251222
transform 1 0 10182 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_7
timestamp 1612251222
transform 1 0 10166 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_6
timestamp 1612251222
transform 1 0 10150 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_5
timestamp 1612251222
transform 1 0 10134 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_4
timestamp 1612251222
transform 1 0 10118 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_3
timestamp 1612251222
transform 1 0 10102 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_2
timestamp 1612251222
transform 1 0 10086 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_1
timestamp 1612251222
transform 1 0 10070 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_320
timestamp 1612251222
transform 1 0 9904 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_320
timestamp 1612251222
transform 1 0 9888 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_320
timestamp 1612251222
transform 1 0 9872 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_320
timestamp 1612251222
transform 1 0 9856 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_320
timestamp 1612251222
transform 1 0 9840 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_145
timestamp 1612251222
transform -1 0 9840 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_145
timestamp 1612251222
transform -1 0 9674 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_145
timestamp 1612251222
transform -1 0 9658 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_145
timestamp 1612251222
transform -1 0 9642 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_145
timestamp 1612251222
transform -1 0 9626 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_209
timestamp 1612251222
transform 1 0 9444 0 1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_209
timestamp 1612251222
transform 1 0 9428 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_209
timestamp 1612251222
transform 1 0 9412 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_209
timestamp 1612251222
transform 1 0 9396 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_149
timestamp 1612251222
transform 1 0 9230 0 1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_149
timestamp 1612251222
transform 1 0 9214 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_149
timestamp 1612251222
transform 1 0 9198 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_149
timestamp 1612251222
transform 1 0 9182 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_684
timestamp 1612251222
transform -1 0 9182 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_684
timestamp 1612251222
transform -1 0 9016 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_684
timestamp 1612251222
transform -1 0 9000 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_684
timestamp 1612251222
transform -1 0 8984 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_684
timestamp 1612251222
transform -1 0 8968 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_603
timestamp 1612251222
transform -1 0 8952 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_603
timestamp 1612251222
transform -1 0 8786 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_603
timestamp 1612251222
transform -1 0 8770 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_603
timestamp 1612251222
transform -1 0 8754 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_603
timestamp 1612251222
transform -1 0 8738 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_605
timestamp 1612251222
transform -1 0 8722 0 1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_605
timestamp 1612251222
transform -1 0 8556 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_605
timestamp 1612251222
transform -1 0 8540 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_605
timestamp 1612251222
transform -1 0 8524 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_677
timestamp 1612251222
transform -1 0 8508 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_677
timestamp 1612251222
transform -1 0 8342 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_677
timestamp 1612251222
transform -1 0 8326 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_677
timestamp 1612251222
transform -1 0 8310 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_677
timestamp 1612251222
transform -1 0 8294 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_645
timestamp 1612251222
transform -1 0 8278 0 1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_645
timestamp 1612251222
transform -1 0 8112 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_645
timestamp 1612251222
transform -1 0 8096 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_645
timestamp 1612251222
transform -1 0 8080 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_648
timestamp 1612251222
transform -1 0 8064 0 1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_648
timestamp 1612251222
transform -1 0 7898 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_648
timestamp 1612251222
transform -1 0 7882 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_648
timestamp 1612251222
transform -1 0 7866 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_407
timestamp 1612251222
transform 1 0 7684 0 1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_407
timestamp 1612251222
transform 1 0 7668 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_407
timestamp 1612251222
transform 1 0 7652 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_407
timestamp 1612251222
transform 1 0 7636 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_779
timestamp 1612251222
transform 1 0 7470 0 1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_779
timestamp 1612251222
transform 1 0 7454 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_779
timestamp 1612251222
transform 1 0 7438 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_779
timestamp 1612251222
transform 1 0 7422 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_708
timestamp 1612251222
transform -1 0 7422 0 1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_708
timestamp 1612251222
transform -1 0 7256 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_708
timestamp 1612251222
transform -1 0 7240 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_708
timestamp 1612251222
transform -1 0 7224 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_697
timestamp 1612251222
transform 1 0 7042 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_697
timestamp 1612251222
transform 1 0 7026 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_697
timestamp 1612251222
transform 1 0 7010 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_697
timestamp 1612251222
transform 1 0 6994 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_697
timestamp 1612251222
transform 1 0 6978 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_712
timestamp 1612251222
transform -1 0 6978 0 1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_712
timestamp 1612251222
transform -1 0 6812 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_712
timestamp 1612251222
transform -1 0 6796 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_712
timestamp 1612251222
transform -1 0 6780 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_766
timestamp 1612251222
transform 1 0 6598 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_766
timestamp 1612251222
transform 1 0 6582 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_766
timestamp 1612251222
transform 1 0 6566 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_766
timestamp 1612251222
transform 1 0 6550 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_766
timestamp 1612251222
transform 1 0 6534 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_386
timestamp 1612251222
transform 1 0 6368 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_386
timestamp 1612251222
transform 1 0 6352 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_386
timestamp 1612251222
transform 1 0 6336 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_386
timestamp 1612251222
transform 1 0 6320 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_386
timestamp 1612251222
transform 1 0 6304 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_59
timestamp 1612251222
transform 1 0 6138 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_59
timestamp 1612251222
transform 1 0 6122 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_59
timestamp 1612251222
transform 1 0 6106 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_59
timestamp 1612251222
transform 1 0 6090 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_59
timestamp 1612251222
transform 1 0 6074 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_26
timestamp 1612251222
transform 1 0 5908 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_26
timestamp 1612251222
transform 1 0 5892 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_26
timestamp 1612251222
transform 1 0 5876 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_26
timestamp 1612251222
transform 1 0 5860 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_26
timestamp 1612251222
transform 1 0 5844 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_64
timestamp 1612251222
transform 1 0 5678 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_64
timestamp 1612251222
transform 1 0 5662 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_64
timestamp 1612251222
transform 1 0 5646 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_64
timestamp 1612251222
transform 1 0 5630 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_64
timestamp 1612251222
transform 1 0 5614 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_21
timestamp 1612251222
transform 1 0 5448 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_21
timestamp 1612251222
transform 1 0 5432 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_21
timestamp 1612251222
transform 1 0 5416 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_21
timestamp 1612251222
transform 1 0 5400 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_21
timestamp 1612251222
transform 1 0 5384 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_21
timestamp 1612251222
transform -1 0 5384 0 1 1010
box -4 -6 170 206
use FILL  FILL2_POR2X1_21
timestamp 1612251222
transform -1 0 5218 0 1 1010
box -4 -6 20 206
use FILL  FILL1_POR2X1_21
timestamp 1612251222
transform -1 0 5202 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_21
timestamp 1612251222
transform -1 0 5186 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_21
timestamp 1612251222
transform -1 0 5170 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_3
timestamp 1612251222
transform 1 0 4988 0 1 1010
box -4 -6 170 206
use FILL  FILL2_POR2X1_3
timestamp 1612251222
transform 1 0 4972 0 1 1010
box -4 -6 20 206
use FILL  FILL1_POR2X1_3
timestamp 1612251222
transform 1 0 4956 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_3
timestamp 1612251222
transform 1 0 4940 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_3
timestamp 1612251222
transform 1 0 4924 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_12
timestamp 1612251222
transform 1 0 4758 0 1 1010
box -4 -6 170 206
use FILL  FILL2_POR2X1_12
timestamp 1612251222
transform 1 0 4742 0 1 1010
box -4 -6 20 206
use FILL  FILL1_POR2X1_12
timestamp 1612251222
transform 1 0 4726 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_12
timestamp 1612251222
transform 1 0 4710 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_12
timestamp 1612251222
transform 1 0 4694 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_36
timestamp 1612251222
transform 1 0 4528 0 1 1010
box -4 -6 170 206
use FILL  FILL2_POR2X1_36
timestamp 1612251222
transform 1 0 4512 0 1 1010
box -4 -6 20 206
use FILL  FILL1_POR2X1_36
timestamp 1612251222
transform 1 0 4496 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_36
timestamp 1612251222
transform 1 0 4480 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_36
timestamp 1612251222
transform 1 0 4464 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_64
timestamp 1612251222
transform -1 0 4464 0 1 1010
box -4 -6 170 206
use FILL  FILL2_POR2X1_64
timestamp 1612251222
transform -1 0 4298 0 1 1010
box -4 -6 20 206
use FILL  FILL1_POR2X1_64
timestamp 1612251222
transform -1 0 4282 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_64
timestamp 1612251222
transform -1 0 4266 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_64
timestamp 1612251222
transform -1 0 4250 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_744
timestamp 1612251222
transform -1 0 4234 0 1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_744
timestamp 1612251222
transform -1 0 4068 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_744
timestamp 1612251222
transform -1 0 4052 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_744
timestamp 1612251222
transform -1 0 4036 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_547
timestamp 1612251222
transform -1 0 4020 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_547
timestamp 1612251222
transform -1 0 3854 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_547
timestamp 1612251222
transform -1 0 3838 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_547
timestamp 1612251222
transform -1 0 3822 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_547
timestamp 1612251222
transform -1 0 3806 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_779
timestamp 1612251222
transform 1 0 3624 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_779
timestamp 1612251222
transform 1 0 3608 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_779
timestamp 1612251222
transform 1 0 3592 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_779
timestamp 1612251222
transform 1 0 3576 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_779
timestamp 1612251222
transform 1 0 3560 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_527
timestamp 1612251222
transform 1 0 3394 0 1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_527
timestamp 1612251222
transform 1 0 3378 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_527
timestamp 1612251222
transform 1 0 3362 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_527
timestamp 1612251222
transform 1 0 3346 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_549
timestamp 1612251222
transform -1 0 3346 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_549
timestamp 1612251222
transform -1 0 3180 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_549
timestamp 1612251222
transform -1 0 3164 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_549
timestamp 1612251222
transform -1 0 3148 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_549
timestamp 1612251222
transform -1 0 3132 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_693
timestamp 1612251222
transform -1 0 3116 0 1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_693
timestamp 1612251222
transform -1 0 2950 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_693
timestamp 1612251222
transform -1 0 2934 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_693
timestamp 1612251222
transform -1 0 2918 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_485
timestamp 1612251222
transform -1 0 2902 0 1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_485
timestamp 1612251222
transform -1 0 2736 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_485
timestamp 1612251222
transform -1 0 2720 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_485
timestamp 1612251222
transform -1 0 2704 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_323
timestamp 1612251222
transform -1 0 2688 0 1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_323
timestamp 1612251222
transform -1 0 2522 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_323
timestamp 1612251222
transform -1 0 2506 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_323
timestamp 1612251222
transform -1 0 2490 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_325
timestamp 1612251222
transform -1 0 2474 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_325
timestamp 1612251222
transform -1 0 2308 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_325
timestamp 1612251222
transform -1 0 2292 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_325
timestamp 1612251222
transform -1 0 2276 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_325
timestamp 1612251222
transform -1 0 2260 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_165
timestamp 1612251222
transform 1 0 2078 0 1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_165
timestamp 1612251222
transform 1 0 2062 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_165
timestamp 1612251222
transform 1 0 2046 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_165
timestamp 1612251222
transform 1 0 2030 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_170
timestamp 1612251222
transform -1 0 2030 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_170
timestamp 1612251222
transform -1 0 1864 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_170
timestamp 1612251222
transform -1 0 1848 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_170
timestamp 1612251222
transform -1 0 1832 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_170
timestamp 1612251222
transform -1 0 1816 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_724
timestamp 1612251222
transform -1 0 1800 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_724
timestamp 1612251222
transform -1 0 1634 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_724
timestamp 1612251222
transform -1 0 1618 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_724
timestamp 1612251222
transform -1 0 1602 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_724
timestamp 1612251222
transform -1 0 1586 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_714
timestamp 1612251222
transform 1 0 1404 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_714
timestamp 1612251222
transform 1 0 1388 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_714
timestamp 1612251222
transform 1 0 1372 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_714
timestamp 1612251222
transform 1 0 1356 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_714
timestamp 1612251222
transform 1 0 1340 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_169
timestamp 1612251222
transform 1 0 1174 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_169
timestamp 1612251222
transform 1 0 1158 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_169
timestamp 1612251222
transform 1 0 1142 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_169
timestamp 1612251222
transform 1 0 1126 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_169
timestamp 1612251222
transform 1 0 1110 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_166
timestamp 1612251222
transform 1 0 944 0 1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_166
timestamp 1612251222
transform 1 0 928 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_166
timestamp 1612251222
transform 1 0 912 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_166
timestamp 1612251222
transform 1 0 896 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_167
timestamp 1612251222
transform 1 0 730 0 1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_167
timestamp 1612251222
transform 1 0 714 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_167
timestamp 1612251222
transform 1 0 698 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_167
timestamp 1612251222
transform 1 0 682 0 1 1010
box -4 -6 20 206
use POR2X1  POR2X1_765
timestamp 1612251222
transform -1 0 682 0 1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_765
timestamp 1612251222
transform -1 0 516 0 1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_765
timestamp 1612251222
transform -1 0 500 0 1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_765
timestamp 1612251222
transform -1 0 484 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_564
timestamp 1612251222
transform -1 0 468 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_564
timestamp 1612251222
transform -1 0 302 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_564
timestamp 1612251222
transform -1 0 286 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_564
timestamp 1612251222
transform -1 0 270 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_564
timestamp 1612251222
transform -1 0 254 0 1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_569
timestamp 1612251222
transform -1 0 238 0 1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_569
timestamp 1612251222
transform -1 0 72 0 1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_569
timestamp 1612251222
transform -1 0 56 0 1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_569
timestamp 1612251222
transform -1 0 40 0 1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_569
timestamp 1612251222
transform -1 0 24 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_13
timestamp 1612251222
transform -1 0 10262 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_12
timestamp 1612251222
transform -1 0 10246 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_11
timestamp 1612251222
transform -1 0 10230 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_10
timestamp 1612251222
transform -1 0 10214 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_9
timestamp 1612251222
transform -1 0 10198 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_8
timestamp 1612251222
transform -1 0 10182 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_7
timestamp 1612251222
transform -1 0 10166 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_6
timestamp 1612251222
transform -1 0 10150 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_5
timestamp 1612251222
transform -1 0 10134 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_4
timestamp 1612251222
transform -1 0 10118 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_3
timestamp 1612251222
transform -1 0 10102 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_2
timestamp 1612251222
transform -1 0 10086 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_1
timestamp 1612251222
transform -1 0 10070 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_213
timestamp 1612251222
transform 1 0 9888 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_213
timestamp 1612251222
transform 1 0 9872 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_213
timestamp 1612251222
transform 1 0 9856 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_213
timestamp 1612251222
transform 1 0 9840 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_146
timestamp 1612251222
transform -1 0 9840 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_146
timestamp 1612251222
transform -1 0 9674 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_146
timestamp 1612251222
transform -1 0 9658 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_146
timestamp 1612251222
transform -1 0 9642 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_146
timestamp 1612251222
transform -1 0 9626 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_148
timestamp 1612251222
transform -1 0 9610 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_148
timestamp 1612251222
transform -1 0 9444 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_148
timestamp 1612251222
transform -1 0 9428 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_148
timestamp 1612251222
transform -1 0 9412 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_329
timestamp 1612251222
transform 1 0 9230 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_329
timestamp 1612251222
transform 1 0 9214 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_329
timestamp 1612251222
transform 1 0 9198 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_329
timestamp 1612251222
transform 1 0 9182 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_329
timestamp 1612251222
transform 1 0 9166 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_421
timestamp 1612251222
transform -1 0 9166 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_421
timestamp 1612251222
transform -1 0 9000 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_421
timestamp 1612251222
transform -1 0 8984 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_421
timestamp 1612251222
transform -1 0 8968 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_421
timestamp 1612251222
transform -1 0 8952 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_604
timestamp 1612251222
transform -1 0 8936 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_604
timestamp 1612251222
transform -1 0 8770 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_604
timestamp 1612251222
transform -1 0 8754 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_604
timestamp 1612251222
transform -1 0 8738 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_604
timestamp 1612251222
transform -1 0 8722 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_683
timestamp 1612251222
transform 1 0 8540 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_683
timestamp 1612251222
transform 1 0 8524 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_683
timestamp 1612251222
transform 1 0 8508 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_683
timestamp 1612251222
transform 1 0 8492 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_683
timestamp 1612251222
transform 1 0 8476 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_678
timestamp 1612251222
transform 1 0 8310 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_678
timestamp 1612251222
transform 1 0 8294 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_678
timestamp 1612251222
transform 1 0 8278 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_678
timestamp 1612251222
transform 1 0 8262 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_834
timestamp 1612251222
transform -1 0 8262 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_834
timestamp 1612251222
transform -1 0 8096 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_834
timestamp 1612251222
transform -1 0 8080 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_834
timestamp 1612251222
transform -1 0 8064 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_644
timestamp 1612251222
transform 1 0 7882 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_644
timestamp 1612251222
transform 1 0 7866 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_644
timestamp 1612251222
transform 1 0 7850 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_644
timestamp 1612251222
transform 1 0 7834 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_597
timestamp 1612251222
transform 1 0 7668 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_597
timestamp 1612251222
transform 1 0 7652 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_597
timestamp 1612251222
transform 1 0 7636 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_597
timestamp 1612251222
transform 1 0 7620 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_597
timestamp 1612251222
transform 1 0 7604 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_596
timestamp 1612251222
transform 1 0 7438 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_596
timestamp 1612251222
transform 1 0 7422 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_596
timestamp 1612251222
transform 1 0 7406 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_596
timestamp 1612251222
transform 1 0 7390 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_743
timestamp 1612251222
transform 1 0 7224 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_743
timestamp 1612251222
transform 1 0 7208 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_743
timestamp 1612251222
transform 1 0 7192 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_743
timestamp 1612251222
transform 1 0 7176 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_743
timestamp 1612251222
transform 1 0 7160 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_765
timestamp 1612251222
transform -1 0 7160 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_765
timestamp 1612251222
transform -1 0 6994 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_765
timestamp 1612251222
transform -1 0 6978 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_765
timestamp 1612251222
transform -1 0 6962 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_765
timestamp 1612251222
transform -1 0 6946 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_770
timestamp 1612251222
transform -1 0 6930 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_770
timestamp 1612251222
transform -1 0 6764 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_770
timestamp 1612251222
transform -1 0 6748 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_770
timestamp 1612251222
transform -1 0 6732 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_328
timestamp 1612251222
transform 1 0 6550 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_328
timestamp 1612251222
transform 1 0 6534 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_328
timestamp 1612251222
transform 1 0 6518 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_328
timestamp 1612251222
transform 1 0 6502 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_328
timestamp 1612251222
transform 1 0 6486 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_707
timestamp 1612251222
transform 1 0 6320 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_707
timestamp 1612251222
transform 1 0 6304 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_707
timestamp 1612251222
transform 1 0 6288 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_707
timestamp 1612251222
transform 1 0 6272 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_695
timestamp 1612251222
transform 1 0 6106 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_695
timestamp 1612251222
transform 1 0 6090 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_695
timestamp 1612251222
transform 1 0 6074 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_695
timestamp 1612251222
transform 1 0 6058 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_695
timestamp 1612251222
transform 1 0 6042 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_40
timestamp 1612251222
transform 1 0 5876 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_40
timestamp 1612251222
transform 1 0 5860 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_40
timestamp 1612251222
transform 1 0 5844 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_40
timestamp 1612251222
transform 1 0 5828 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_40
timestamp 1612251222
transform 1 0 5812 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_409
timestamp 1612251222
transform -1 0 5812 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_409
timestamp 1612251222
transform -1 0 5646 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_409
timestamp 1612251222
transform -1 0 5630 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_409
timestamp 1612251222
transform -1 0 5614 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_409
timestamp 1612251222
transform -1 0 5598 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_22
timestamp 1612251222
transform -1 0 5582 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_22
timestamp 1612251222
transform -1 0 5416 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_22
timestamp 1612251222
transform -1 0 5400 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_22
timestamp 1612251222
transform -1 0 5384 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_22
timestamp 1612251222
transform -1 0 5368 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_3
timestamp 1612251222
transform 1 0 5186 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_3
timestamp 1612251222
transform 1 0 5170 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_3
timestamp 1612251222
transform 1 0 5154 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_3
timestamp 1612251222
transform 1 0 5138 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_3
timestamp 1612251222
transform 1 0 5122 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_12
timestamp 1612251222
transform -1 0 5122 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_12
timestamp 1612251222
transform -1 0 4956 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_12
timestamp 1612251222
transform -1 0 4940 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_12
timestamp 1612251222
transform -1 0 4924 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_12
timestamp 1612251222
transform -1 0 4908 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_587
timestamp 1612251222
transform -1 0 4892 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_587
timestamp 1612251222
transform -1 0 4726 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_587
timestamp 1612251222
transform -1 0 4710 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_587
timestamp 1612251222
transform -1 0 4694 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_51
timestamp 1612251222
transform -1 0 4678 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_POR2X1_51
timestamp 1612251222
transform -1 0 4512 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_POR2X1_51
timestamp 1612251222
transform -1 0 4496 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_51
timestamp 1612251222
transform -1 0 4480 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_51
timestamp 1612251222
transform -1 0 4464 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_44
timestamp 1612251222
transform -1 0 4448 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_POR2X1_44
timestamp 1612251222
transform -1 0 4282 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_POR2X1_44
timestamp 1612251222
transform -1 0 4266 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_44
timestamp 1612251222
transform -1 0 4250 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_44
timestamp 1612251222
transform -1 0 4234 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_50
timestamp 1612251222
transform -1 0 4218 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_POR2X1_50
timestamp 1612251222
transform -1 0 4052 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_POR2X1_50
timestamp 1612251222
transform -1 0 4036 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_50
timestamp 1612251222
transform -1 0 4020 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_50
timestamp 1612251222
transform -1 0 4004 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_95
timestamp 1612251222
transform -1 0 3988 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_95
timestamp 1612251222
transform -1 0 3822 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_95
timestamp 1612251222
transform -1 0 3806 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_95
timestamp 1612251222
transform -1 0 3790 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_70
timestamp 1612251222
transform -1 0 3774 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_POR2X1_70
timestamp 1612251222
transform -1 0 3608 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_POR2X1_70
timestamp 1612251222
transform -1 0 3592 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_70
timestamp 1612251222
transform -1 0 3576 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_70
timestamp 1612251222
transform -1 0 3560 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_511
timestamp 1612251222
transform 1 0 3378 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_511
timestamp 1612251222
transform 1 0 3362 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_511
timestamp 1612251222
transform 1 0 3346 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_511
timestamp 1612251222
transform 1 0 3330 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_531
timestamp 1612251222
transform 1 0 3164 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_531
timestamp 1612251222
transform 1 0 3148 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_531
timestamp 1612251222
transform 1 0 3132 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_531
timestamp 1612251222
transform 1 0 3116 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_427
timestamp 1612251222
transform 1 0 2950 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_427
timestamp 1612251222
transform 1 0 2934 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_427
timestamp 1612251222
transform 1 0 2918 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_427
timestamp 1612251222
transform 1 0 2902 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_697
timestamp 1612251222
transform 1 0 2736 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_697
timestamp 1612251222
transform 1 0 2720 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_697
timestamp 1612251222
transform 1 0 2704 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_697
timestamp 1612251222
transform 1 0 2688 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_164
timestamp 1612251222
transform -1 0 2688 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_164
timestamp 1612251222
transform -1 0 2522 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_164
timestamp 1612251222
transform -1 0 2506 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_164
timestamp 1612251222
transform -1 0 2490 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_565
timestamp 1612251222
transform -1 0 2474 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_565
timestamp 1612251222
transform -1 0 2308 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_565
timestamp 1612251222
transform -1 0 2292 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_565
timestamp 1612251222
transform -1 0 2276 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_565
timestamp 1612251222
transform -1 0 2260 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_168
timestamp 1612251222
transform -1 0 2244 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_168
timestamp 1612251222
transform -1 0 2078 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_168
timestamp 1612251222
transform -1 0 2062 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_168
timestamp 1612251222
transform -1 0 2046 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_168
timestamp 1612251222
transform -1 0 2030 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_374
timestamp 1612251222
transform 1 0 1848 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_374
timestamp 1612251222
transform 1 0 1832 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_374
timestamp 1612251222
transform 1 0 1816 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_374
timestamp 1612251222
transform 1 0 1800 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_374
timestamp 1612251222
transform 1 0 1784 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_322
timestamp 1612251222
transform 1 0 1618 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_322
timestamp 1612251222
transform 1 0 1602 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_322
timestamp 1612251222
transform 1 0 1586 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_322
timestamp 1612251222
transform 1 0 1570 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_373
timestamp 1612251222
transform -1 0 1570 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_373
timestamp 1612251222
transform -1 0 1404 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_373
timestamp 1612251222
transform -1 0 1388 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_373
timestamp 1612251222
transform -1 0 1372 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_438
timestamp 1612251222
transform -1 0 1356 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_438
timestamp 1612251222
transform -1 0 1190 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_438
timestamp 1612251222
transform -1 0 1174 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_438
timestamp 1612251222
transform -1 0 1158 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_544
timestamp 1612251222
transform -1 0 1142 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_544
timestamp 1612251222
transform -1 0 976 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_544
timestamp 1612251222
transform -1 0 960 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_544
timestamp 1612251222
transform -1 0 944 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_544
timestamp 1612251222
transform -1 0 928 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_326
timestamp 1612251222
transform -1 0 912 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_326
timestamp 1612251222
transform -1 0 746 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_326
timestamp 1612251222
transform -1 0 730 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_326
timestamp 1612251222
transform -1 0 714 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_326
timestamp 1612251222
transform -1 0 698 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_551
timestamp 1612251222
transform -1 0 682 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_551
timestamp 1612251222
transform -1 0 516 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_551
timestamp 1612251222
transform -1 0 500 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_551
timestamp 1612251222
transform -1 0 484 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_551
timestamp 1612251222
transform -1 0 468 0 -1 1010
box -4 -6 20 206
use POR2X1  POR2X1_766
timestamp 1612251222
transform -1 0 452 0 -1 1010
box -4 -6 170 206
use FILL  FILL1_POR2X1_766
timestamp 1612251222
transform -1 0 286 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_POR2X1_766
timestamp 1612251222
transform -1 0 270 0 -1 1010
box -4 -6 20 206
use FILL  FILL_POR2X1_766
timestamp 1612251222
transform -1 0 254 0 -1 1010
box -4 -6 20 206
use PAND2X1  PAND2X1_770
timestamp 1612251222
transform -1 0 238 0 -1 1010
box -4 -6 170 206
use FILL  FILL2_PAND2X1_770
timestamp 1612251222
transform -1 0 72 0 -1 1010
box -4 -6 20 206
use FILL  FILL1_PAND2X1_770
timestamp 1612251222
transform -1 0 56 0 -1 1010
box -4 -6 20 206
use FILL  FILL0_PAND2X1_770
timestamp 1612251222
transform -1 0 40 0 -1 1010
box -4 -6 20 206
use FILL  FILL_PAND2X1_770
timestamp 1612251222
transform -1 0 24 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1
timestamp 1612251222
transform 1 0 10252 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_160
timestamp 1612251222
transform 1 0 10086 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_160
timestamp 1612251222
transform 1 0 10070 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_160
timestamp 1612251222
transform 1 0 10054 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_160
timestamp 1612251222
transform 1 0 10038 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_745
timestamp 1612251222
transform 1 0 9872 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_745
timestamp 1612251222
transform 1 0 9856 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_745
timestamp 1612251222
transform 1 0 9840 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_745
timestamp 1612251222
transform 1 0 9824 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_745
timestamp 1612251222
transform 1 0 9808 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_746
timestamp 1612251222
transform 1 0 9642 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_746
timestamp 1612251222
transform 1 0 9626 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_746
timestamp 1612251222
transform 1 0 9610 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_746
timestamp 1612251222
transform 1 0 9594 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_746
timestamp 1612251222
transform 1 0 9578 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_856
timestamp 1612251222
transform -1 0 9578 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_856
timestamp 1612251222
transform -1 0 9412 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_856
timestamp 1612251222
transform -1 0 9396 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_856
timestamp 1612251222
transform -1 0 9380 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_863
timestamp 1612251222
transform -1 0 9364 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_863
timestamp 1612251222
transform -1 0 9198 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_863
timestamp 1612251222
transform -1 0 9182 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_863
timestamp 1612251222
transform -1 0 9166 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_829
timestamp 1612251222
transform 1 0 8984 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_829
timestamp 1612251222
transform 1 0 8968 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_829
timestamp 1612251222
transform 1 0 8952 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_829
timestamp 1612251222
transform 1 0 8936 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_829
timestamp 1612251222
transform 1 0 8920 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_686
timestamp 1612251222
transform -1 0 8920 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_686
timestamp 1612251222
transform -1 0 8754 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_686
timestamp 1612251222
transform -1 0 8738 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_686
timestamp 1612251222
transform -1 0 8722 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_760
timestamp 1612251222
transform -1 0 8706 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_760
timestamp 1612251222
transform -1 0 8540 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_760
timestamp 1612251222
transform -1 0 8524 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_760
timestamp 1612251222
transform -1 0 8508 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_760
timestamp 1612251222
transform -1 0 8492 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_828
timestamp 1612251222
transform 1 0 8310 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_828
timestamp 1612251222
transform 1 0 8294 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_828
timestamp 1612251222
transform 1 0 8278 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_828
timestamp 1612251222
transform 1 0 8262 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_598
timestamp 1612251222
transform 1 0 8096 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_598
timestamp 1612251222
transform 1 0 8080 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_598
timestamp 1612251222
transform 1 0 8064 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_598
timestamp 1612251222
transform 1 0 8048 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_744
timestamp 1612251222
transform -1 0 8048 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_744
timestamp 1612251222
transform -1 0 7882 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_744
timestamp 1612251222
transform -1 0 7866 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_744
timestamp 1612251222
transform -1 0 7850 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_744
timestamp 1612251222
transform -1 0 7834 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_780
timestamp 1612251222
transform 1 0 7652 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_780
timestamp 1612251222
transform 1 0 7636 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_780
timestamp 1612251222
transform 1 0 7620 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_780
timestamp 1612251222
transform 1 0 7604 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_811
timestamp 1612251222
transform -1 0 7604 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_811
timestamp 1612251222
transform -1 0 7438 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_811
timestamp 1612251222
transform -1 0 7422 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_811
timestamp 1612251222
transform -1 0 7406 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_688
timestamp 1612251222
transform -1 0 7390 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_688
timestamp 1612251222
transform -1 0 7224 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_688
timestamp 1612251222
transform -1 0 7208 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_688
timestamp 1612251222
transform -1 0 7192 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_690
timestamp 1612251222
transform 1 0 7010 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_690
timestamp 1612251222
transform 1 0 6994 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_690
timestamp 1612251222
transform 1 0 6978 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_690
timestamp 1612251222
transform 1 0 6962 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_690
timestamp 1612251222
transform 1 0 6946 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_771
timestamp 1612251222
transform 1 0 6780 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_771
timestamp 1612251222
transform 1 0 6764 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_771
timestamp 1612251222
transform 1 0 6748 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_771
timestamp 1612251222
transform 1 0 6732 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_764
timestamp 1612251222
transform -1 0 6732 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_764
timestamp 1612251222
transform -1 0 6566 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_764
timestamp 1612251222
transform -1 0 6550 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_764
timestamp 1612251222
transform -1 0 6534 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_764
timestamp 1612251222
transform -1 0 6518 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_428
timestamp 1612251222
transform -1 0 6502 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_428
timestamp 1612251222
transform -1 0 6336 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_428
timestamp 1612251222
transform -1 0 6320 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_428
timestamp 1612251222
transform -1 0 6304 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_428
timestamp 1612251222
transform -1 0 6288 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_47
timestamp 1612251222
transform 1 0 6106 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_47
timestamp 1612251222
transform 1 0 6090 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_47
timestamp 1612251222
transform 1 0 6074 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_47
timestamp 1612251222
transform 1 0 6058 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_47
timestamp 1612251222
transform 1 0 6042 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_44
timestamp 1612251222
transform -1 0 6042 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_44
timestamp 1612251222
transform -1 0 5876 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_44
timestamp 1612251222
transform -1 0 5860 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_44
timestamp 1612251222
transform -1 0 5844 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_44
timestamp 1612251222
transform -1 0 5828 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_408
timestamp 1612251222
transform 1 0 5646 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_408
timestamp 1612251222
transform 1 0 5630 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_408
timestamp 1612251222
transform 1 0 5614 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_408
timestamp 1612251222
transform 1 0 5598 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_408
timestamp 1612251222
transform 1 0 5582 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_36
timestamp 1612251222
transform -1 0 5582 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_36
timestamp 1612251222
transform -1 0 5416 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_36
timestamp 1612251222
transform -1 0 5400 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_36
timestamp 1612251222
transform -1 0 5384 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_36
timestamp 1612251222
transform -1 0 5368 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_1
timestamp 1612251222
transform 1 0 5186 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_1
timestamp 1612251222
transform 1 0 5170 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_1
timestamp 1612251222
transform 1 0 5154 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_1
timestamp 1612251222
transform 1 0 5138 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_1
timestamp 1612251222
transform 1 0 5122 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_30
timestamp 1612251222
transform -1 0 5122 0 1 610
box -4 -6 170 206
use FILL  FILL2_POR2X1_30
timestamp 1612251222
transform -1 0 4956 0 1 610
box -4 -6 20 206
use FILL  FILL1_POR2X1_30
timestamp 1612251222
transform -1 0 4940 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_30
timestamp 1612251222
transform -1 0 4924 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_30
timestamp 1612251222
transform -1 0 4908 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_31
timestamp 1612251222
transform -1 0 4892 0 1 610
box -4 -6 170 206
use FILL  FILL2_POR2X1_31
timestamp 1612251222
transform -1 0 4726 0 1 610
box -4 -6 20 206
use FILL  FILL1_POR2X1_31
timestamp 1612251222
transform -1 0 4710 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_31
timestamp 1612251222
transform -1 0 4694 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_31
timestamp 1612251222
transform -1 0 4678 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_26
timestamp 1612251222
transform -1 0 4662 0 1 610
box -4 -6 170 206
use FILL  FILL2_POR2X1_26
timestamp 1612251222
transform -1 0 4496 0 1 610
box -4 -6 20 206
use FILL  FILL1_POR2X1_26
timestamp 1612251222
transform -1 0 4480 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_26
timestamp 1612251222
transform -1 0 4464 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_26
timestamp 1612251222
transform -1 0 4448 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_47
timestamp 1612251222
transform -1 0 4432 0 1 610
box -4 -6 170 206
use FILL  FILL2_POR2X1_47
timestamp 1612251222
transform -1 0 4266 0 1 610
box -4 -6 20 206
use FILL  FILL1_POR2X1_47
timestamp 1612251222
transform -1 0 4250 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_47
timestamp 1612251222
transform -1 0 4234 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_47
timestamp 1612251222
transform -1 0 4218 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_40
timestamp 1612251222
transform -1 0 4202 0 1 610
box -4 -6 170 206
use FILL  FILL2_POR2X1_40
timestamp 1612251222
transform -1 0 4036 0 1 610
box -4 -6 20 206
use FILL  FILL1_POR2X1_40
timestamp 1612251222
transform -1 0 4020 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_40
timestamp 1612251222
transform -1 0 4004 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_40
timestamp 1612251222
transform -1 0 3988 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_698
timestamp 1612251222
transform 1 0 3806 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_698
timestamp 1612251222
transform 1 0 3790 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_698
timestamp 1612251222
transform 1 0 3774 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_698
timestamp 1612251222
transform 1 0 3758 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_59
timestamp 1612251222
transform -1 0 3758 0 1 610
box -4 -6 170 206
use FILL  FILL2_POR2X1_59
timestamp 1612251222
transform -1 0 3592 0 1 610
box -4 -6 20 206
use FILL  FILL1_POR2X1_59
timestamp 1612251222
transform -1 0 3576 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_59
timestamp 1612251222
transform -1 0 3560 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_59
timestamp 1612251222
transform -1 0 3544 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_701
timestamp 1612251222
transform 1 0 3362 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_701
timestamp 1612251222
transform 1 0 3346 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_701
timestamp 1612251222
transform 1 0 3330 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_701
timestamp 1612251222
transform 1 0 3314 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_428
timestamp 1612251222
transform 1 0 3148 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_428
timestamp 1612251222
transform 1 0 3132 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_428
timestamp 1612251222
transform 1 0 3116 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_428
timestamp 1612251222
transform 1 0 3100 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_696
timestamp 1612251222
transform -1 0 3100 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_696
timestamp 1612251222
transform -1 0 2934 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_696
timestamp 1612251222
transform -1 0 2918 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_696
timestamp 1612251222
transform -1 0 2902 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_708
timestamp 1612251222
transform -1 0 2886 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_708
timestamp 1612251222
transform -1 0 2720 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_708
timestamp 1612251222
transform -1 0 2704 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_708
timestamp 1612251222
transform -1 0 2688 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_708
timestamp 1612251222
transform -1 0 2672 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_550
timestamp 1612251222
transform -1 0 2656 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_550
timestamp 1612251222
transform -1 0 2490 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_550
timestamp 1612251222
transform -1 0 2474 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_550
timestamp 1612251222
transform -1 0 2458 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_550
timestamp 1612251222
transform -1 0 2442 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_706
timestamp 1612251222
transform -1 0 2426 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_706
timestamp 1612251222
transform -1 0 2260 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_706
timestamp 1612251222
transform -1 0 2244 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_706
timestamp 1612251222
transform -1 0 2228 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_706
timestamp 1612251222
transform -1 0 2212 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_526
timestamp 1612251222
transform 1 0 2030 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_526
timestamp 1612251222
transform 1 0 2014 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_526
timestamp 1612251222
transform 1 0 1998 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_526
timestamp 1612251222
transform 1 0 1982 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_152
timestamp 1612251222
transform -1 0 1982 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_152
timestamp 1612251222
transform -1 0 1816 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_152
timestamp 1612251222
transform -1 0 1800 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_152
timestamp 1612251222
transform -1 0 1784 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_441
timestamp 1612251222
transform -1 0 1768 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_441
timestamp 1612251222
transform -1 0 1602 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_441
timestamp 1612251222
transform -1 0 1586 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_441
timestamp 1612251222
transform -1 0 1570 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_144
timestamp 1612251222
transform -1 0 1554 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_144
timestamp 1612251222
transform -1 0 1388 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_144
timestamp 1612251222
transform -1 0 1372 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_144
timestamp 1612251222
transform -1 0 1356 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_147
timestamp 1612251222
transform -1 0 1340 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_147
timestamp 1612251222
transform -1 0 1174 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_147
timestamp 1612251222
transform -1 0 1158 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_147
timestamp 1612251222
transform -1 0 1142 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_147
timestamp 1612251222
transform -1 0 1126 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_142
timestamp 1612251222
transform 1 0 944 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_142
timestamp 1612251222
transform 1 0 928 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_142
timestamp 1612251222
transform 1 0 912 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_142
timestamp 1612251222
transform 1 0 896 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_321
timestamp 1612251222
transform -1 0 896 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_321
timestamp 1612251222
transform -1 0 730 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_321
timestamp 1612251222
transform -1 0 714 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_321
timestamp 1612251222
transform -1 0 698 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_545
timestamp 1612251222
transform 1 0 516 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_545
timestamp 1612251222
transform 1 0 500 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_545
timestamp 1612251222
transform 1 0 484 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_545
timestamp 1612251222
transform 1 0 468 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_545
timestamp 1612251222
transform 1 0 452 0 1 610
box -4 -6 20 206
use POR2X1  POR2X1_764
timestamp 1612251222
transform -1 0 452 0 1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_764
timestamp 1612251222
transform -1 0 286 0 1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_764
timestamp 1612251222
transform -1 0 270 0 1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_764
timestamp 1612251222
transform -1 0 254 0 1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_771
timestamp 1612251222
transform 1 0 72 0 1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_771
timestamp 1612251222
transform 1 0 56 0 1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_771
timestamp 1612251222
transform 1 0 40 0 1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_771
timestamp 1612251222
transform 1 0 24 0 1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_771
timestamp 1612251222
transform 1 0 8 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1
timestamp 1612251222
transform -1 0 10268 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_356
timestamp 1612251222
transform 1 0 10086 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_356
timestamp 1612251222
transform 1 0 10070 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_356
timestamp 1612251222
transform 1 0 10054 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_356
timestamp 1612251222
transform 1 0 10038 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_781
timestamp 1612251222
transform -1 0 10038 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_781
timestamp 1612251222
transform -1 0 9872 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_781
timestamp 1612251222
transform -1 0 9856 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_781
timestamp 1612251222
transform -1 0 9840 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_747
timestamp 1612251222
transform -1 0 9824 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_747
timestamp 1612251222
transform -1 0 9658 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_747
timestamp 1612251222
transform -1 0 9642 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_747
timestamp 1612251222
transform -1 0 9626 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_747
timestamp 1612251222
transform -1 0 9610 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_782
timestamp 1612251222
transform -1 0 9594 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_782
timestamp 1612251222
transform -1 0 9428 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_782
timestamp 1612251222
transform -1 0 9412 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_782
timestamp 1612251222
transform -1 0 9396 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_797
timestamp 1612251222
transform -1 0 9380 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_797
timestamp 1612251222
transform -1 0 9214 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_797
timestamp 1612251222
transform -1 0 9198 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_797
timestamp 1612251222
transform -1 0 9182 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_855
timestamp 1612251222
transform 1 0 9000 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_855
timestamp 1612251222
transform 1 0 8984 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_855
timestamp 1612251222
transform 1 0 8968 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_855
timestamp 1612251222
transform 1 0 8952 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_154
timestamp 1612251222
transform 1 0 8786 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_154
timestamp 1612251222
transform 1 0 8770 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_154
timestamp 1612251222
transform 1 0 8754 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_154
timestamp 1612251222
transform 1 0 8738 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_803
timestamp 1612251222
transform -1 0 8738 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_803
timestamp 1612251222
transform -1 0 8572 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_803
timestamp 1612251222
transform -1 0 8556 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_803
timestamp 1612251222
transform -1 0 8540 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_808
timestamp 1612251222
transform -1 0 8524 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_808
timestamp 1612251222
transform -1 0 8358 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_808
timestamp 1612251222
transform -1 0 8342 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_808
timestamp 1612251222
transform -1 0 8326 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_599
timestamp 1612251222
transform -1 0 8310 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_599
timestamp 1612251222
transform -1 0 8144 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_599
timestamp 1612251222
transform -1 0 8128 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_599
timestamp 1612251222
transform -1 0 8112 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_599
timestamp 1612251222
transform -1 0 8096 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_796
timestamp 1612251222
transform 1 0 7914 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_796
timestamp 1612251222
transform 1 0 7898 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_796
timestamp 1612251222
transform 1 0 7882 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_796
timestamp 1612251222
transform 1 0 7866 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_783
timestamp 1612251222
transform 1 0 7700 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_783
timestamp 1612251222
transform 1 0 7684 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_783
timestamp 1612251222
transform 1 0 7668 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_783
timestamp 1612251222
transform 1 0 7652 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_691
timestamp 1612251222
transform 1 0 7486 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_691
timestamp 1612251222
transform 1 0 7470 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_691
timestamp 1612251222
transform 1 0 7454 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_691
timestamp 1612251222
transform 1 0 7438 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_689
timestamp 1612251222
transform 1 0 7272 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_689
timestamp 1612251222
transform 1 0 7256 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_689
timestamp 1612251222
transform 1 0 7240 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_689
timestamp 1612251222
transform 1 0 7224 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_689
timestamp 1612251222
transform 1 0 7208 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_774
timestamp 1612251222
transform 1 0 7042 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_774
timestamp 1612251222
transform 1 0 7026 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_774
timestamp 1612251222
transform 1 0 7010 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_774
timestamp 1612251222
transform 1 0 6994 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_584
timestamp 1612251222
transform -1 0 6994 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_584
timestamp 1612251222
transform -1 0 6828 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_584
timestamp 1612251222
transform -1 0 6812 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_584
timestamp 1612251222
transform -1 0 6796 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_584
timestamp 1612251222
transform -1 0 6780 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_769
timestamp 1612251222
transform 1 0 6598 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_769
timestamp 1612251222
transform 1 0 6582 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_769
timestamp 1612251222
transform 1 0 6566 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_769
timestamp 1612251222
transform 1 0 6550 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_763
timestamp 1612251222
transform 1 0 6384 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_763
timestamp 1612251222
transform 1 0 6368 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_763
timestamp 1612251222
transform 1 0 6352 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_763
timestamp 1612251222
transform 1 0 6336 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_763
timestamp 1612251222
transform 1 0 6320 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_762
timestamp 1612251222
transform 1 0 6154 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_762
timestamp 1612251222
transform 1 0 6138 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_762
timestamp 1612251222
transform 1 0 6122 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_762
timestamp 1612251222
transform 1 0 6106 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_762
timestamp 1612251222
transform 1 0 6090 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_25
timestamp 1612251222
transform 1 0 5924 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_25
timestamp 1612251222
transform 1 0 5908 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_25
timestamp 1612251222
transform 1 0 5892 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_25
timestamp 1612251222
transform 1 0 5876 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_25
timestamp 1612251222
transform 1 0 5860 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_587
timestamp 1612251222
transform 1 0 5694 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_587
timestamp 1612251222
transform 1 0 5678 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_587
timestamp 1612251222
transform 1 0 5662 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_587
timestamp 1612251222
transform 1 0 5646 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_587
timestamp 1612251222
transform 1 0 5630 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_31
timestamp 1612251222
transform -1 0 5630 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_31
timestamp 1612251222
transform -1 0 5464 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_31
timestamp 1612251222
transform -1 0 5448 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_31
timestamp 1612251222
transform -1 0 5432 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_31
timestamp 1612251222
transform -1 0 5416 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_50
timestamp 1612251222
transform 1 0 5234 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_50
timestamp 1612251222
transform 1 0 5218 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_50
timestamp 1612251222
transform 1 0 5202 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_50
timestamp 1612251222
transform 1 0 5186 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_50
timestamp 1612251222
transform 1 0 5170 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_1
timestamp 1612251222
transform -1 0 5170 0 -1 610
box -4 -6 170 206
use FILL  FILL2_POR2X1_1
timestamp 1612251222
transform -1 0 5004 0 -1 610
box -4 -6 20 206
use FILL  FILL1_POR2X1_1
timestamp 1612251222
transform -1 0 4988 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_1
timestamp 1612251222
transform -1 0 4972 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_1
timestamp 1612251222
transform -1 0 4956 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_25
timestamp 1612251222
transform -1 0 4940 0 -1 610
box -4 -6 170 206
use FILL  FILL2_POR2X1_25
timestamp 1612251222
transform -1 0 4774 0 -1 610
box -4 -6 20 206
use FILL  FILL1_POR2X1_25
timestamp 1612251222
transform -1 0 4758 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_25
timestamp 1612251222
transform -1 0 4742 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_25
timestamp 1612251222
transform -1 0 4726 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_18
timestamp 1612251222
transform 1 0 4544 0 -1 610
box -4 -6 170 206
use FILL  FILL2_POR2X1_18
timestamp 1612251222
transform 1 0 4528 0 -1 610
box -4 -6 20 206
use FILL  FILL1_POR2X1_18
timestamp 1612251222
transform 1 0 4512 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_18
timestamp 1612251222
transform 1 0 4496 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_18
timestamp 1612251222
transform 1 0 4480 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_762
timestamp 1612251222
transform -1 0 4480 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_762
timestamp 1612251222
transform -1 0 4314 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_762
timestamp 1612251222
transform -1 0 4298 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_762
timestamp 1612251222
transform -1 0 4282 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_635
timestamp 1612251222
transform 1 0 4100 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_635
timestamp 1612251222
transform 1 0 4084 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_635
timestamp 1612251222
transform 1 0 4068 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_635
timestamp 1612251222
transform 1 0 4052 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_635
timestamp 1612251222
transform 1 0 4036 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_709
timestamp 1612251222
transform -1 0 4036 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_709
timestamp 1612251222
transform -1 0 3870 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_709
timestamp 1612251222
transform -1 0 3854 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_709
timestamp 1612251222
transform -1 0 3838 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_709
timestamp 1612251222
transform -1 0 3822 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_700
timestamp 1612251222
transform 1 0 3640 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_700
timestamp 1612251222
transform 1 0 3624 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_700
timestamp 1612251222
transform 1 0 3608 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_700
timestamp 1612251222
transform 1 0 3592 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_710
timestamp 1612251222
transform -1 0 3592 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_710
timestamp 1612251222
transform -1 0 3426 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_710
timestamp 1612251222
transform -1 0 3410 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_710
timestamp 1612251222
transform -1 0 3394 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_710
timestamp 1612251222
transform -1 0 3378 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_711
timestamp 1612251222
transform -1 0 3362 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_711
timestamp 1612251222
transform -1 0 3196 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_711
timestamp 1612251222
transform -1 0 3180 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_711
timestamp 1612251222
transform -1 0 3164 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_711
timestamp 1612251222
transform -1 0 3148 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_763
timestamp 1612251222
transform -1 0 3132 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_763
timestamp 1612251222
transform -1 0 2966 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_763
timestamp 1612251222
transform -1 0 2950 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_763
timestamp 1612251222
transform -1 0 2934 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_525
timestamp 1612251222
transform -1 0 2918 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_525
timestamp 1612251222
transform -1 0 2752 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_525
timestamp 1612251222
transform -1 0 2736 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_525
timestamp 1612251222
transform -1 0 2720 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_546
timestamp 1612251222
transform 1 0 2538 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_546
timestamp 1612251222
transform 1 0 2522 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_546
timestamp 1612251222
transform 1 0 2506 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_546
timestamp 1612251222
transform 1 0 2490 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_546
timestamp 1612251222
transform 1 0 2474 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_692
timestamp 1612251222
transform 1 0 2308 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_692
timestamp 1612251222
transform 1 0 2292 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_692
timestamp 1612251222
transform 1 0 2276 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_692
timestamp 1612251222
transform 1 0 2260 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_486
timestamp 1612251222
transform -1 0 2260 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_486
timestamp 1612251222
transform -1 0 2094 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_486
timestamp 1612251222
transform -1 0 2078 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_486
timestamp 1612251222
transform -1 0 2062 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_486
timestamp 1612251222
transform -1 0 2046 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_484
timestamp 1612251222
transform 1 0 1864 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_484
timestamp 1612251222
transform 1 0 1848 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_484
timestamp 1612251222
transform 1 0 1832 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_484
timestamp 1612251222
transform 1 0 1816 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_726
timestamp 1612251222
transform -1 0 1816 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_726
timestamp 1612251222
transform -1 0 1650 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_726
timestamp 1612251222
transform -1 0 1634 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_726
timestamp 1612251222
transform -1 0 1618 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_726
timestamp 1612251222
transform -1 0 1602 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_732
timestamp 1612251222
transform -1 0 1586 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_732
timestamp 1612251222
transform -1 0 1420 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_732
timestamp 1612251222
transform -1 0 1404 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_732
timestamp 1612251222
transform -1 0 1388 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_732
timestamp 1612251222
transform -1 0 1372 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_731
timestamp 1612251222
transform -1 0 1356 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_731
timestamp 1612251222
transform -1 0 1190 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_731
timestamp 1612251222
transform -1 0 1174 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_731
timestamp 1612251222
transform -1 0 1158 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_731
timestamp 1612251222
transform -1 0 1142 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_738
timestamp 1612251222
transform -1 0 1126 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_738
timestamp 1612251222
transform -1 0 960 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_738
timestamp 1612251222
transform -1 0 944 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_738
timestamp 1612251222
transform -1 0 928 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_738
timestamp 1612251222
transform -1 0 912 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_320
timestamp 1612251222
transform -1 0 896 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_320
timestamp 1612251222
transform -1 0 730 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_320
timestamp 1612251222
transform -1 0 714 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_320
timestamp 1612251222
transform -1 0 698 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_324
timestamp 1612251222
transform -1 0 682 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_324
timestamp 1612251222
transform -1 0 516 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_324
timestamp 1612251222
transform -1 0 500 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_324
timestamp 1612251222
transform -1 0 484 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_324
timestamp 1612251222
transform -1 0 468 0 -1 610
box -4 -6 20 206
use POR2X1  POR2X1_524
timestamp 1612251222
transform 1 0 286 0 -1 610
box -4 -6 170 206
use FILL  FILL1_POR2X1_524
timestamp 1612251222
transform 1 0 270 0 -1 610
box -4 -6 20 206
use FILL  FILL0_POR2X1_524
timestamp 1612251222
transform 1 0 254 0 -1 610
box -4 -6 20 206
use FILL  FILL_POR2X1_524
timestamp 1612251222
transform 1 0 238 0 -1 610
box -4 -6 20 206
use PAND2X1  PAND2X1_769
timestamp 1612251222
transform -1 0 238 0 -1 610
box -4 -6 170 206
use FILL  FILL2_PAND2X1_769
timestamp 1612251222
transform -1 0 72 0 -1 610
box -4 -6 20 206
use FILL  FILL1_PAND2X1_769
timestamp 1612251222
transform -1 0 56 0 -1 610
box -4 -6 20 206
use FILL  FILL0_PAND2X1_769
timestamp 1612251222
transform -1 0 40 0 -1 610
box -4 -6 20 206
use FILL  FILL_PAND2X1_769
timestamp 1612251222
transform -1 0 24 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_5
timestamp 1612251222
transform 1 0 10252 0 1 210
box -4 -6 20 206
use FILL  FILL_1_12
timestamp 1612251222
transform -1 0 10246 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_13
timestamp 1612251222
transform -1 0 10262 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_4
timestamp 1612251222
transform 1 0 10236 0 1 210
box -4 -6 20 206
use FILL  FILL_1_11
timestamp 1612251222
transform -1 0 10230 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_2
timestamp 1612251222
transform 1 0 10204 0 1 210
box -4 -6 20 206
use FILL  FILL_2_3
timestamp 1612251222
transform 1 0 10220 0 1 210
box -4 -6 20 206
use FILL  FILL_1_9
timestamp 1612251222
transform -1 0 10198 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_10
timestamp 1612251222
transform -1 0 10214 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_1
timestamp 1612251222
transform 1 0 10188 0 1 210
box -4 -6 20 206
use FILL  FILL_1_8
timestamp 1612251222
transform -1 0 10182 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_6
timestamp 1612251222
transform -1 0 10150 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_7
timestamp 1612251222
transform -1 0 10166 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_162
timestamp 1612251222
transform -1 0 10188 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_162
timestamp 1612251222
transform -1 0 10022 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_162
timestamp 1612251222
transform -1 0 10006 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_162
timestamp 1612251222
transform -1 0 9990 0 1 210
box -4 -6 20 206
use FILL  FILL_1_5
timestamp 1612251222
transform -1 0 10134 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_4
timestamp 1612251222
transform -1 0 10118 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_3
timestamp 1612251222
transform -1 0 10102 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_2
timestamp 1612251222
transform -1 0 10086 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_1
timestamp 1612251222
transform -1 0 10070 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_161
timestamp 1612251222
transform 1 0 9808 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_161
timestamp 1612251222
transform 1 0 9792 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_568
timestamp 1612251222
transform -1 0 10054 0 -1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_568
timestamp 1612251222
transform -1 0 9888 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_568
timestamp 1612251222
transform -1 0 9872 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_568
timestamp 1612251222
transform -1 0 9856 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_161
timestamp 1612251222
transform 1 0 9776 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_161
timestamp 1612251222
transform 1 0 9760 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_289
timestamp 1612251222
transform 1 0 9674 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_289
timestamp 1612251222
transform 1 0 9658 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_289
timestamp 1612251222
transform 1 0 9642 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_289
timestamp 1612251222
transform 1 0 9626 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_289
timestamp 1612251222
transform 1 0 9610 0 -1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_680
timestamp 1612251222
transform -1 0 9760 0 1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_680
timestamp 1612251222
transform -1 0 9594 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_680
timestamp 1612251222
transform -1 0 9578 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_680
timestamp 1612251222
transform -1 0 9562 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_680
timestamp 1612251222
transform -1 0 9546 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_220
timestamp 1612251222
transform 1 0 9444 0 -1 210
box -4 -6 170 206
use PAND2X1  PAND2X1_158
timestamp 1612251222
transform -1 0 9530 0 1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_158
timestamp 1612251222
transform -1 0 9364 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_158
timestamp 1612251222
transform -1 0 9348 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_158
timestamp 1612251222
transform -1 0 9332 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_158
timestamp 1612251222
transform -1 0 9316 0 1 210
box -4 -6 20 206
use FILL  FILL1_POR2X1_220
timestamp 1612251222
transform 1 0 9428 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_220
timestamp 1612251222
transform 1 0 9412 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_220
timestamp 1612251222
transform 1 0 9396 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_156
timestamp 1612251222
transform 1 0 9134 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_156
timestamp 1612251222
transform 1 0 9118 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_156
timestamp 1612251222
transform 1 0 9102 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_156
timestamp 1612251222
transform 1 0 9086 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_210
timestamp 1612251222
transform 1 0 9230 0 -1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_210
timestamp 1612251222
transform 1 0 9214 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_210
timestamp 1612251222
transform 1 0 9198 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_210
timestamp 1612251222
transform 1 0 9182 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_155
timestamp 1612251222
transform 1 0 8920 0 1 210
box -4 -6 170 206
use POR2X1  POR2X1_330
timestamp 1612251222
transform 1 0 9016 0 -1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_330
timestamp 1612251222
transform 1 0 9000 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_330
timestamp 1612251222
transform 1 0 8984 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_330
timestamp 1612251222
transform 1 0 8968 0 -1 210
box -4 -6 20 206
use FILL  FILL1_POR2X1_155
timestamp 1612251222
transform 1 0 8904 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_155
timestamp 1612251222
transform 1 0 8888 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_155
timestamp 1612251222
transform 1 0 8872 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_163
timestamp 1612251222
transform -1 0 8968 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_163
timestamp 1612251222
transform -1 0 8802 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_163
timestamp 1612251222
transform -1 0 8786 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_163
timestamp 1612251222
transform -1 0 8770 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_163
timestamp 1612251222
transform -1 0 8754 0 -1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_682
timestamp 1612251222
transform -1 0 8872 0 1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_682
timestamp 1612251222
transform -1 0 8706 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_682
timestamp 1612251222
transform -1 0 8690 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_682
timestamp 1612251222
transform -1 0 8674 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_682
timestamp 1612251222
transform -1 0 8658 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_467
timestamp 1612251222
transform 1 0 8572 0 -1 210
box -4 -6 170 206
use PAND2X1  PAND2X1_679
timestamp 1612251222
transform 1 0 8476 0 1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_679
timestamp 1612251222
transform 1 0 8460 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_679
timestamp 1612251222
transform 1 0 8444 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_679
timestamp 1612251222
transform 1 0 8428 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_679
timestamp 1612251222
transform 1 0 8412 0 1 210
box -4 -6 20 206
use FILL  FILL1_POR2X1_467
timestamp 1612251222
transform 1 0 8556 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_467
timestamp 1612251222
transform 1 0 8540 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_467
timestamp 1612251222
transform 1 0 8524 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_676
timestamp 1612251222
transform 1 0 8246 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_676
timestamp 1612251222
transform 1 0 8230 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_676
timestamp 1612251222
transform 1 0 8214 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_728
timestamp 1612251222
transform -1 0 8524 0 -1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_728
timestamp 1612251222
transform -1 0 8358 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_728
timestamp 1612251222
transform -1 0 8342 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_728
timestamp 1612251222
transform -1 0 8326 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_676
timestamp 1612251222
transform 1 0 8198 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_730
timestamp 1612251222
transform 1 0 8144 0 -1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_730
timestamp 1612251222
transform 1 0 8128 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_730
timestamp 1612251222
transform 1 0 8112 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_730
timestamp 1612251222
transform 1 0 8096 0 -1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_681
timestamp 1612251222
transform -1 0 8198 0 1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_681
timestamp 1612251222
transform -1 0 8032 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_681
timestamp 1612251222
transform -1 0 8016 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_681
timestamp 1612251222
transform -1 0 8000 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_681
timestamp 1612251222
transform -1 0 7984 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_685
timestamp 1612251222
transform -1 0 8096 0 -1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_685
timestamp 1612251222
transform -1 0 7930 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_685
timestamp 1612251222
transform -1 0 7914 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_685
timestamp 1612251222
transform -1 0 7898 0 -1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_761
timestamp 1612251222
transform -1 0 7968 0 1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_761
timestamp 1612251222
transform -1 0 7802 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_761
timestamp 1612251222
transform -1 0 7786 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_761
timestamp 1612251222
transform -1 0 7770 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_761
timestamp 1612251222
transform -1 0 7754 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_687
timestamp 1612251222
transform -1 0 7882 0 -1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_687
timestamp 1612251222
transform -1 0 7716 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_864
timestamp 1612251222
transform -1 0 7738 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_864
timestamp 1612251222
transform -1 0 7572 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_864
timestamp 1612251222
transform -1 0 7556 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_864
timestamp 1612251222
transform -1 0 7540 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_687
timestamp 1612251222
transform -1 0 7700 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_687
timestamp 1612251222
transform -1 0 7684 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_866
timestamp 1612251222
transform -1 0 7524 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_866
timestamp 1612251222
transform -1 0 7358 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_729
timestamp 1612251222
transform 1 0 7502 0 -1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_729
timestamp 1612251222
transform 1 0 7486 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_729
timestamp 1612251222
transform 1 0 7470 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_729
timestamp 1612251222
transform 1 0 7454 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_866
timestamp 1612251222
transform -1 0 7342 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_866
timestamp 1612251222
transform -1 0 7326 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_800
timestamp 1612251222
transform -1 0 7454 0 -1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_800
timestamp 1612251222
transform -1 0 7288 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_800
timestamp 1612251222
transform -1 0 7272 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_800
timestamp 1612251222
transform -1 0 7256 0 -1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_583
timestamp 1612251222
transform -1 0 7310 0 1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_583
timestamp 1612251222
transform -1 0 7144 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_583
timestamp 1612251222
transform -1 0 7128 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_583
timestamp 1612251222
transform -1 0 7112 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_583
timestamp 1612251222
transform -1 0 7096 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_801
timestamp 1612251222
transform -1 0 7240 0 -1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_801
timestamp 1612251222
transform -1 0 7074 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_801
timestamp 1612251222
transform -1 0 7058 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_801
timestamp 1612251222
transform -1 0 7042 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_810
timestamp 1612251222
transform -1 0 7080 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_810
timestamp 1612251222
transform -1 0 6914 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_810
timestamp 1612251222
transform -1 0 6898 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_810
timestamp 1612251222
transform -1 0 6882 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_809
timestamp 1612251222
transform -1 0 7026 0 -1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_809
timestamp 1612251222
transform -1 0 6860 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_809
timestamp 1612251222
transform -1 0 6844 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_636
timestamp 1612251222
transform -1 0 6866 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_636
timestamp 1612251222
transform -1 0 6700 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_636
timestamp 1612251222
transform -1 0 6684 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_636
timestamp 1612251222
transform -1 0 6668 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_809
timestamp 1612251222
transform -1 0 6828 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_812
timestamp 1612251222
transform -1 0 6812 0 -1 210
box -4 -6 170 206
use POR2X1  POR2X1_639
timestamp 1612251222
transform 1 0 6486 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_639
timestamp 1612251222
transform 1 0 6470 0 1 210
box -4 -6 20 206
use FILL  FILL1_POR2X1_812
timestamp 1612251222
transform -1 0 6646 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_812
timestamp 1612251222
transform -1 0 6630 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_812
timestamp 1612251222
transform -1 0 6614 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_639
timestamp 1612251222
transform 1 0 6454 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_639
timestamp 1612251222
transform 1 0 6438 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_452
timestamp 1612251222
transform 1 0 6432 0 -1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_452
timestamp 1612251222
transform 1 0 6416 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_452
timestamp 1612251222
transform 1 0 6400 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_452
timestamp 1612251222
transform 1 0 6384 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_451
timestamp 1612251222
transform 1 0 6272 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_451
timestamp 1612251222
transform 1 0 6256 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_451
timestamp 1612251222
transform 1 0 6240 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_451
timestamp 1612251222
transform 1 0 6224 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_450
timestamp 1612251222
transform 1 0 6218 0 -1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_450
timestamp 1612251222
transform 1 0 6202 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_450
timestamp 1612251222
transform 1 0 6186 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_450
timestamp 1612251222
transform 1 0 6170 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_635
timestamp 1612251222
transform 1 0 6058 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_635
timestamp 1612251222
transform 1 0 6042 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_635
timestamp 1612251222
transform 1 0 6026 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_635
timestamp 1612251222
transform 1 0 6010 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_427
timestamp 1612251222
transform 1 0 6004 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_427
timestamp 1612251222
transform 1 0 5988 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_427
timestamp 1612251222
transform 1 0 5972 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_427
timestamp 1612251222
transform 1 0 5956 0 -1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_70
timestamp 1612251222
transform 1 0 5844 0 1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_70
timestamp 1612251222
transform 1 0 5828 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_70
timestamp 1612251222
transform 1 0 5812 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_70
timestamp 1612251222
transform 1 0 5796 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_70
timestamp 1612251222
transform 1 0 5780 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_427
timestamp 1612251222
transform 1 0 5940 0 -1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_426
timestamp 1612251222
transform 1 0 5774 0 -1 210
box -4 -6 170 206
use PAND2X1  PAND2X1_51
timestamp 1612251222
transform 1 0 5614 0 1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_51
timestamp 1612251222
transform 1 0 5598 0 1 210
box -4 -6 20 206
use FILL  FILL2_PAND2X1_426
timestamp 1612251222
transform 1 0 5758 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_426
timestamp 1612251222
transform 1 0 5742 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_426
timestamp 1612251222
transform 1 0 5726 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_426
timestamp 1612251222
transform 1 0 5710 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_51
timestamp 1612251222
transform 1 0 5582 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_51
timestamp 1612251222
transform 1 0 5566 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_51
timestamp 1612251222
transform 1 0 5550 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_694
timestamp 1612251222
transform 1 0 5544 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_694
timestamp 1612251222
transform 1 0 5528 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_694
timestamp 1612251222
transform 1 0 5512 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_694
timestamp 1612251222
transform 1 0 5496 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_694
timestamp 1612251222
transform 1 0 5480 0 -1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_582
timestamp 1612251222
transform 1 0 5314 0 -1 210
box -4 -6 170 206
use PAND2X1  PAND2X1_30
timestamp 1612251222
transform 1 0 5384 0 1 210
box -4 -6 170 206
use FILL  FILL0_PAND2X1_30
timestamp 1612251222
transform 1 0 5336 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_30
timestamp 1612251222
transform 1 0 5352 0 1 210
box -4 -6 20 206
use FILL  FILL2_PAND2X1_30
timestamp 1612251222
transform 1 0 5368 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_582
timestamp 1612251222
transform 1 0 5250 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_582
timestamp 1612251222
transform 1 0 5266 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_582
timestamp 1612251222
transform 1 0 5282 0 -1 210
box -4 -6 20 206
use FILL  FILL2_PAND2X1_582
timestamp 1612251222
transform 1 0 5298 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_30
timestamp 1612251222
transform 1 0 5320 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_430
timestamp 1612251222
transform 1 0 5154 0 1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_430
timestamp 1612251222
transform 1 0 5138 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_430
timestamp 1612251222
transform 1 0 5122 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_430
timestamp 1612251222
transform 1 0 5106 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_430
timestamp 1612251222
transform 1 0 5090 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_581
timestamp 1612251222
transform 1 0 5084 0 -1 210
box -4 -6 170 206
use PAND2X1  PAND2X1_429
timestamp 1612251222
transform 1 0 4924 0 1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_429
timestamp 1612251222
transform 1 0 4908 0 1 210
box -4 -6 20 206
use FILL  FILL2_PAND2X1_581
timestamp 1612251222
transform 1 0 5068 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_581
timestamp 1612251222
transform 1 0 5052 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_581
timestamp 1612251222
transform 1 0 5036 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_581
timestamp 1612251222
transform 1 0 5020 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_429
timestamp 1612251222
transform 1 0 4892 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_429
timestamp 1612251222
transform 1 0 4876 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_429
timestamp 1612251222
transform 1 0 4860 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_157
timestamp 1612251222
transform 1 0 4854 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_157
timestamp 1612251222
transform 1 0 4838 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_157
timestamp 1612251222
transform 1 0 4822 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_157
timestamp 1612251222
transform 1 0 4806 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_157
timestamp 1612251222
transform 1 0 4790 0 -1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_2
timestamp 1612251222
transform 1 0 4624 0 -1 210
box -4 -6 170 206
use PAND2X1  PAND2X1_11
timestamp 1612251222
transform 1 0 4694 0 1 210
box -4 -6 170 206
use FILL  FILL0_PAND2X1_11
timestamp 1612251222
transform 1 0 4646 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_11
timestamp 1612251222
transform 1 0 4662 0 1 210
box -4 -6 20 206
use FILL  FILL2_PAND2X1_11
timestamp 1612251222
transform 1 0 4678 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_2
timestamp 1612251222
transform 1 0 4560 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_2
timestamp 1612251222
transform 1 0 4576 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_2
timestamp 1612251222
transform 1 0 4592 0 -1 210
box -4 -6 20 206
use FILL  FILL2_PAND2X1_2
timestamp 1612251222
transform 1 0 4608 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_11
timestamp 1612251222
transform 1 0 4630 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_17
timestamp 1612251222
transform -1 0 4630 0 1 210
box -4 -6 170 206
use FILL  FILL2_POR2X1_17
timestamp 1612251222
transform -1 0 4464 0 1 210
box -4 -6 20 206
use FILL  FILL1_POR2X1_17
timestamp 1612251222
transform -1 0 4448 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_17
timestamp 1612251222
transform -1 0 4432 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_17
timestamp 1612251222
transform -1 0 4416 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_425
timestamp 1612251222
transform 1 0 4394 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_425
timestamp 1612251222
transform 1 0 4378 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_581
timestamp 1612251222
transform -1 0 4400 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_581
timestamp 1612251222
transform -1 0 4234 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_581
timestamp 1612251222
transform -1 0 4218 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_425
timestamp 1612251222
transform 1 0 4362 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_425
timestamp 1612251222
transform 1 0 4346 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_425
timestamp 1612251222
transform 1 0 4330 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_581
timestamp 1612251222
transform -1 0 4202 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_17
timestamp 1612251222
transform 1 0 4164 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_17
timestamp 1612251222
transform 1 0 4148 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_17
timestamp 1612251222
transform 1 0 4132 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_17
timestamp 1612251222
transform 1 0 4116 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_17
timestamp 1612251222
transform 1 0 4100 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_582
timestamp 1612251222
transform -1 0 4186 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_582
timestamp 1612251222
transform -1 0 4020 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_582
timestamp 1612251222
transform -1 0 4004 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_582
timestamp 1612251222
transform -1 0 3988 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_11
timestamp 1612251222
transform -1 0 4100 0 -1 210
box -4 -6 170 206
use FILL  FILL2_POR2X1_11
timestamp 1612251222
transform -1 0 3934 0 -1 210
box -4 -6 20 206
use FILL  FILL1_POR2X1_11
timestamp 1612251222
transform -1 0 3918 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_11
timestamp 1612251222
transform -1 0 3902 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_11
timestamp 1612251222
transform -1 0 3886 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_157
timestamp 1612251222
transform 1 0 3806 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_157
timestamp 1612251222
transform 1 0 3790 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_157
timestamp 1612251222
transform 1 0 3774 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_157
timestamp 1612251222
transform 1 0 3758 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_2
timestamp 1612251222
transform -1 0 3870 0 -1 210
box -4 -6 170 206
use FILL  FILL2_POR2X1_2
timestamp 1612251222
transform -1 0 3704 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_425
timestamp 1612251222
transform -1 0 3758 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_425
timestamp 1612251222
transform -1 0 3592 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_425
timestamp 1612251222
transform -1 0 3576 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_425
timestamp 1612251222
transform -1 0 3560 0 1 210
box -4 -6 20 206
use FILL  FILL1_POR2X1_2
timestamp 1612251222
transform -1 0 3688 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_2
timestamp 1612251222
transform -1 0 3672 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_2
timestamp 1612251222
transform -1 0 3656 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_158
timestamp 1612251222
transform -1 0 3544 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_158
timestamp 1612251222
transform -1 0 3378 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_158
timestamp 1612251222
transform -1 0 3362 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_158
timestamp 1612251222
transform -1 0 3346 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_429
timestamp 1612251222
transform -1 0 3640 0 -1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_429
timestamp 1612251222
transform -1 0 3474 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_429
timestamp 1612251222
transform -1 0 3458 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_429
timestamp 1612251222
transform -1 0 3442 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_426
timestamp 1612251222
transform -1 0 3330 0 1 210
box -4 -6 170 206
use POR2X1  POR2X1_430
timestamp 1612251222
transform -1 0 3426 0 -1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_430
timestamp 1612251222
transform -1 0 3260 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_430
timestamp 1612251222
transform -1 0 3244 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_430
timestamp 1612251222
transform -1 0 3228 0 -1 210
box -4 -6 20 206
use FILL  FILL1_POR2X1_426
timestamp 1612251222
transform -1 0 3164 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_426
timestamp 1612251222
transform -1 0 3148 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_426
timestamp 1612251222
transform -1 0 3132 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_451
timestamp 1612251222
transform -1 0 3212 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_451
timestamp 1612251222
transform -1 0 3046 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_451
timestamp 1612251222
transform -1 0 3030 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_451
timestamp 1612251222
transform -1 0 3014 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_451
timestamp 1612251222
transform -1 0 2998 0 -1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_450
timestamp 1612251222
transform -1 0 3116 0 1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_450
timestamp 1612251222
transform -1 0 2950 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_450
timestamp 1612251222
transform -1 0 2934 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_450
timestamp 1612251222
transform -1 0 2918 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_450
timestamp 1612251222
transform -1 0 2902 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_452
timestamp 1612251222
transform -1 0 2982 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_452
timestamp 1612251222
transform -1 0 2816 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_695
timestamp 1612251222
transform -1 0 2886 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_695
timestamp 1612251222
transform -1 0 2720 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_695
timestamp 1612251222
transform -1 0 2704 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_695
timestamp 1612251222
transform -1 0 2688 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_452
timestamp 1612251222
transform -1 0 2800 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_452
timestamp 1612251222
transform -1 0 2784 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_452
timestamp 1612251222
transform -1 0 2768 0 -1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_712
timestamp 1612251222
transform -1 0 2672 0 1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_712
timestamp 1612251222
transform -1 0 2506 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_712
timestamp 1612251222
transform -1 0 2490 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_712
timestamp 1612251222
transform -1 0 2474 0 1 210
box -4 -6 20 206
use POR2X1  POR2X1_694
timestamp 1612251222
transform -1 0 2752 0 -1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_694
timestamp 1612251222
transform -1 0 2586 0 -1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_694
timestamp 1612251222
transform -1 0 2570 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_694
timestamp 1612251222
transform -1 0 2554 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_712
timestamp 1612251222
transform -1 0 2458 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_707
timestamp 1612251222
transform -1 0 2538 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_707
timestamp 1612251222
transform -1 0 2372 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_707
timestamp 1612251222
transform -1 0 2356 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_707
timestamp 1612251222
transform -1 0 2340 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_707
timestamp 1612251222
transform -1 0 2324 0 -1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_705
timestamp 1612251222
transform -1 0 2442 0 1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_705
timestamp 1612251222
transform -1 0 2276 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_705
timestamp 1612251222
transform -1 0 2260 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_705
timestamp 1612251222
transform -1 0 2244 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_705
timestamp 1612251222
transform -1 0 2228 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_467
timestamp 1612251222
transform 1 0 2142 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_467
timestamp 1612251222
transform 1 0 2126 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_467
timestamp 1612251222
transform 1 0 2110 0 -1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_713
timestamp 1612251222
transform -1 0 2212 0 1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_713
timestamp 1612251222
transform -1 0 2046 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_713
timestamp 1612251222
transform -1 0 2030 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_713
timestamp 1612251222
transform -1 0 2014 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_713
timestamp 1612251222
transform -1 0 1998 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_467
timestamp 1612251222
transform 1 0 2094 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_467
timestamp 1612251222
transform 1 0 2078 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_163
timestamp 1612251222
transform 1 0 1816 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_163
timestamp 1612251222
transform 1 0 1800 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_163
timestamp 1612251222
transform 1 0 1784 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_163
timestamp 1612251222
transform 1 0 1768 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_725
timestamp 1612251222
transform -1 0 2078 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_725
timestamp 1612251222
transform -1 0 1912 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_725
timestamp 1612251222
transform -1 0 1896 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_725
timestamp 1612251222
transform -1 0 1880 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_725
timestamp 1612251222
transform -1 0 1864 0 -1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_160
timestamp 1612251222
transform -1 0 1768 0 1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_160
timestamp 1612251222
transform -1 0 1602 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_210
timestamp 1612251222
transform -1 0 1848 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_210
timestamp 1612251222
transform -1 0 1682 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_210
timestamp 1612251222
transform -1 0 1666 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_210
timestamp 1612251222
transform -1 0 1650 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_210
timestamp 1612251222
transform -1 0 1634 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_160
timestamp 1612251222
transform -1 0 1586 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_160
timestamp 1612251222
transform -1 0 1570 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_160
timestamp 1612251222
transform -1 0 1554 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_162
timestamp 1612251222
transform 1 0 1452 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_162
timestamp 1612251222
transform 1 0 1436 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_162
timestamp 1612251222
transform 1 0 1420 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_162
timestamp 1612251222
transform 1 0 1404 0 -1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_209
timestamp 1612251222
transform -1 0 1538 0 1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_209
timestamp 1612251222
transform -1 0 1372 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_209
timestamp 1612251222
transform -1 0 1356 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_209
timestamp 1612251222
transform -1 0 1340 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_209
timestamp 1612251222
transform -1 0 1324 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_162
timestamp 1612251222
transform 1 0 1388 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_145
timestamp 1612251222
transform -1 0 1308 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_145
timestamp 1612251222
transform -1 0 1142 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_145
timestamp 1612251222
transform -1 0 1126 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_145
timestamp 1612251222
transform -1 0 1110 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_213
timestamp 1612251222
transform -1 0 1388 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_213
timestamp 1612251222
transform -1 0 1222 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_213
timestamp 1612251222
transform -1 0 1206 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_213
timestamp 1612251222
transform -1 0 1190 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_213
timestamp 1612251222
transform -1 0 1174 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_146
timestamp 1612251222
transform -1 0 1094 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_146
timestamp 1612251222
transform -1 0 928 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_146
timestamp 1612251222
transform -1 0 912 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_161
timestamp 1612251222
transform 1 0 992 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_161
timestamp 1612251222
transform 1 0 976 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_161
timestamp 1612251222
transform 1 0 960 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_161
timestamp 1612251222
transform 1 0 944 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_161
timestamp 1612251222
transform 1 0 928 0 -1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_146
timestamp 1612251222
transform -1 0 896 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_149
timestamp 1612251222
transform -1 0 880 0 1 210
box -4 -6 170 206
use PAND2X1  PAND2X1_148
timestamp 1612251222
transform -1 0 928 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_148
timestamp 1612251222
transform -1 0 762 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_148
timestamp 1612251222
transform -1 0 746 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_148
timestamp 1612251222
transform -1 0 730 0 -1 210
box -4 -6 20 206
use FILL  FILL2_PAND2X1_149
timestamp 1612251222
transform -1 0 714 0 1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_149
timestamp 1612251222
transform -1 0 698 0 1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_149
timestamp 1612251222
transform -1 0 682 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_149
timestamp 1612251222
transform -1 0 666 0 1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_148
timestamp 1612251222
transform -1 0 714 0 -1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_797
timestamp 1612251222
transform 1 0 532 0 -1 210
box -4 -6 170 206
use POR2X1  POR2X1_747
timestamp 1612251222
transform -1 0 650 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_747
timestamp 1612251222
transform -1 0 484 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_747
timestamp 1612251222
transform -1 0 468 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_747
timestamp 1612251222
transform -1 0 452 0 1 210
box -4 -6 20 206
use FILL  FILL2_PAND2X1_797
timestamp 1612251222
transform 1 0 516 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_797
timestamp 1612251222
transform 1 0 500 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_797
timestamp 1612251222
transform 1 0 484 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_797
timestamp 1612251222
transform 1 0 468 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_745
timestamp 1612251222
transform -1 0 436 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_745
timestamp 1612251222
transform -1 0 270 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_745
timestamp 1612251222
transform -1 0 254 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_745
timestamp 1612251222
transform -1 0 238 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_782
timestamp 1612251222
transform 1 0 302 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_782
timestamp 1612251222
transform 1 0 286 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_782
timestamp 1612251222
transform 1 0 270 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_782
timestamp 1612251222
transform 1 0 254 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_782
timestamp 1612251222
transform 1 0 238 0 -1 210
box -4 -6 20 206
use POR2X1  POR2X1_746
timestamp 1612251222
transform -1 0 222 0 1 210
box -4 -6 170 206
use FILL  FILL1_POR2X1_746
timestamp 1612251222
transform -1 0 56 0 1 210
box -4 -6 20 206
use FILL  FILL0_POR2X1_746
timestamp 1612251222
transform -1 0 40 0 1 210
box -4 -6 20 206
use FILL  FILL_POR2X1_746
timestamp 1612251222
transform -1 0 24 0 1 210
box -4 -6 20 206
use PAND2X1  PAND2X1_781
timestamp 1612251222
transform 1 0 72 0 -1 210
box -4 -6 170 206
use FILL  FILL2_PAND2X1_781
timestamp 1612251222
transform 1 0 56 0 -1 210
box -4 -6 20 206
use FILL  FILL1_PAND2X1_781
timestamp 1612251222
transform 1 0 40 0 -1 210
box -4 -6 20 206
use FILL  FILL0_PAND2X1_781
timestamp 1612251222
transform 1 0 24 0 -1 210
box -4 -6 20 206
use FILL  FILL_PAND2X1_781
timestamp 1612251222
transform 1 0 8 0 -1 210
box -4 -6 20 206
<< labels >>
rlabel metal2 s 1104 7680 1104 7680 6 INPUT_0
port 0 nsew
rlabel metal2 s 2784 7680 2784 7680 6 D_INPUT_0
port 1 nsew
rlabel metal2 s 3728 7680 3728 7680 6 INPUT_1
port 2 nsew
rlabel metal2 s 5168 7680 5168 7680 6 D_INPUT_1
port 3 nsew
rlabel metal2 s 3584 7680 3584 7680 6 INPUT_2
port 4 nsew
rlabel metal2 s 3360 7680 3360 7680 6 D_INPUT_2
port 5 nsew
rlabel metal2 s 4352 7680 4352 7680 6 INPUT_3
port 6 nsew
rlabel metal2 s 3920 7680 3920 7680 6 D_INPUT_3
port 7 nsew
rlabel metal2 s 4048 -40 4048 -40 8 INPUT_4
port 8 nsew
rlabel metal2 s 4672 -40 4672 -40 8 D_INPUT_4
port 9 nsew
rlabel metal2 s 3824 -40 3824 -40 8 INPUT_5
port 10 nsew
rlabel metal2 s 4608 -40 4608 -40 8 D_INPUT_5
port 11 nsew
rlabel metal2 s 5104 -40 5104 -40 8 INPUT_6
port 12 nsew
rlabel metal2 s 4384 -40 4384 -40 8 D_INPUT_6
port 13 nsew
rlabel metal2 s 3600 -40 3600 -40 8 INPUT_7
port 14 nsew
rlabel metal2 s 5136 -40 5136 -40 8 D_INPUT_7
port 15 nsew
rlabel metal3 s 10336 5320 10336 5320 6 D_GATE_222
port 16 nsew
rlabel metal3 s 10336 4180 10336 4180 6 D_GATE_366
port 17 nsew
rlabel metal3 s 10336 1840 10336 1840 6 D_GATE_479
port 18 nsew
rlabel metal3 s 10336 7380 10336 7380 6 D_GATE_579
port 19 nsew
rlabel metal3 s 10336 3120 10336 3120 6 D_GATE_662
port 20 nsew
rlabel metal3 s 10336 7320 10336 7320 6 D_GATE_741
port 21 nsew
rlabel metal2 s 6672 -40 6672 -40 8 D_GATE_811
port 22 nsew
rlabel metal2 s 7344 -40 7344 -40 8 D_GATE_865
port 23 nsew
rlabel metal3 s -48 5120 -48 5120 4 GATE_222
port 24 nsew
rlabel metal3 s -48 4980 -48 4980 4 GATE_366
port 25 nsew
rlabel metal2 s 2656 -40 2656 -40 8 GATE_479
port 26 nsew
rlabel metal3 s -48 3780 -48 3780 4 GATE_579
port 27 nsew
rlabel metal2 s 1776 7680 1776 7680 6 GATE_662
port 28 nsew
rlabel metal3 s -48 4720 -48 4720 4 GATE_741
port 29 nsew
rlabel metal3 s -48 4240 -48 4240 4 GATE_811
port 30 nsew
rlabel metal3 s -48 4580 -48 4580 4 GATE_865
port 31 nsew
rlabel metal3 s -48 4800 -48 4800 4 gate
port 32 nsew
rlabel metal2 s 6560 7680 6560 7680 6 type:
port 33 nsew
rlabel metal3 s -48 6500 -48 6500 4 AND;
port 34 nsew
rlabel metal3 s 10336 340 10336 340 6 name:
port 35 nsew
rlabel metal2 s 7568 7680 7568 7680 6 GATE_0_I0
port 36 nsew
rlabel space -51 -43 10339 7683 1 vdd
rlabel space -51 -43 10339 7683 1 gnd
<< end >>
