*** TEST 004 partitioning ***
*
* ngSPICE test for PLS experiments
*
* AES SBOX PLS test init file generator - protected dualRail SBOX area illuminated
*
* Author: Jan Belohoubek, 08/2020
* jan.belohoubek@fit.cvut.cz
*
* https://users.fit.cvut.cz/~belohja4/
*
*
* **************************************

.include ../../models.lib
.include ../../tsmc180nmcmos.lib
.include pDualRail.spice

* **************************************
* --- Test ---
* **************************************

* --- Settings
.param showPlots = 0
.param writeFile = 1
.param run_inputSet = 0

* redefine defaults ...
.include test00X_settings.inc

.csparam showPlots = {showPlots}
.csparam writeFile = {writeFile}
.csparam run_inputSet = {run_inputSet}

.global showPlots writeFile run_inputSet

* --- End of Settins

Vtrig LaserTrig 0 0 PWL(0ns 0V 20ns 0V 21ns SUPP)

.param beamDistanceTop = 0
.param beamDistanceBot = 0

.global LaserTrig beamDistanceTop beamDistanceBot

* --- inputs
Vvin0 INPUT_0 0 0 PWL(0ns 0V 5ns  0V 7ns  0V)
Vvin1 INPUT_1 0 0 PWL(0ns 0V 6ns  0V 8ns  0V)
Vvin2 INPUT_2 0 0 PWL(0ns 0V 7ns  0V 9ns  0V)
Vvin3 INPUT_3 0 0 PWL(0ns 0V 8ns  0V 10ns 0V)
Vvin4 INPUT_4 0 0 PWL(0ns 0V 9ns  0V 11ns 0V)
Vvin5 INPUT_5 0 0 PWL(0ns 0V 10ns 0V 12ns 0V)
Vvin6 INPUT_6 0 0 PWL(0ns 0V 11ns 0V 13ns 0V)
Vvin7 INPUT_7 0 0 PWL(0ns 0V 12ns 0V 14ns 0V)

Vvin0D D_INPUT_0 0 0 PWL(0ns 0V 5ns  0V 7ns  0V)
Vvin1D D_INPUT_1 0 0 PWL(0ns 0V 6ns  0V 8ns  0V)
Vvin2D D_INPUT_2 0 0 PWL(0ns 0V 7ns  0V 9ns  0V)
Vvin3D D_INPUT_3 0 0 PWL(0ns 0V 8ns  0V 10ns 0V)
Vvin4D D_INPUT_4 0 0 PWL(0ns 0V 9ns  0V 11ns 0V)
Vvin5D D_INPUT_5 0 0 PWL(0ns 0V 10ns 0V 12ns 0V)
Vvin6D D_INPUT_6 0 0 PWL(0ns 0V 11ns 0V 13ns 0V)
Vvin7D D_INPUT_7 0 0 PWL(0ns 0V 12ns 0V 14ns 0V)


* --- outputs
C0 VSS GATE_222 10fF
C1 VSS GATE_366 10fF
C2 VSS GATE_479 10fF
C3 VSS GATE_579 10fF
C4 VSS GATE_662 10fF
C5 VSS GATE_741 10fF
C6 VSS GATE_811 10fF
C7 VSS GATE_865 10fF

C0d VSS D_GATE_222 10fF
C1d VSS D_GATE_366 10fF
C2d VSS D_GATE_479 10fF
C3d VSS D_GATE_579 10fF
C4d VSS D_GATE_662 10fF
C5d VSS D_GATE_741 10fF
C6d VSS D_GATE_811 10fF
C7d VSS D_GATE_865 10fF

* --- circuit layout model

Xsbox1 
+ PAND2X1_812/A PAND2X1_366/A PAND2X1_479/B POR2X1_660/A POR2X1_216/Y POR2X1_351/B POR2X1_852/A POR2X1_243/Y POR2X1_472/Y PAND2X1_739/B PAND2X1_863/A PAND2X1_550/Y PAND2X1_724/B PAND2X1_339/Y PAND2X1_721/B POR2X1_362/B POR2X1_858/B PAND2X1_359/B PAND2X1_477/B PAND2X1_362/A PAND2X1_773/B PAND2X1_351/A PAND2X1_714/Y PAND2X1_466/B PAND2X1_350/A PAND2X1_862/B PAND2X1_656/B POR2X1_206/A POR2X1_857/B POR2X1_207/B POR2X1_466/A POR2X1_856/B POR2X1_568/A POR2X1_139/Y PAND2X1_649/A PAND2X1_560/B PAND2X1_207/A PAND2X1_783/Y PAND2X1_840/Y POR2X1_632/Y POR2X1_392/B POR2X1_566/A POR2X1_452/Y POR2X1_723/B POR2X1_552/Y PAND2X1_717/Y PAND2X1_211/A PAND2X1_785/Y PAND2X1_209/A PAND2X1_353/Y PAND2X1_731/B 
+ PAND2X1_725/A PAND2X1_651/Y PAND2X1_472/B PAND2X1_841/Y POR2X1_734/A POR2X1_569/A POR2X1_860/A PAND2X1_658/A POR2X1_640/Y POR2X1_553/Y POR2X1_796/A PAND2X1_725/B PAND2X1_726/B PAND2X1_390/Y PAND2X1_365/A PAND2X1_644/Y PAND2X1_675/A PAND2X1_551/A PAND2X1_645/B PAND2X1_573/B PAND2X1_736/A PAND2X1_123/Y PAND2X1_835/Y PAND2X1_182/A PAND2X1_175/B PAND2X1_781/Y PAND2X1_641/Y PAND2X1_443/Y PAND2X1_545/Y PAND2X1_169/Y PAND2X1_191/Y PAND2X1_555/A PAND2X1_213/B PAND2X1_508/B PAND2X1_719/Y PAND2X1_200/B POR2X1_805/A PAND2X1_467/B POR2X1_730/B POR2X1_149/A POR2X1_467/Y POR2X1_210/Y POR2X1_244/B POR2X1_343/Y POR2X1_444/A POR2X1_785/B POR2X1_559/Y POR2X1_558/B POR2X1_572/B POR2X1_791/Y POR2X1_449/Y 
+ POR2X1_360/A POR2X1_556/A POR2X1_713/B POR2X1_768/Y POR2X1_213/B POR2X1_726/Y POR2X1_403/A POR2X1_554/Y POR2X1_639/Y POR2X1_324/Y POR2X1_644/Y POR2X1_200/A POR2X1_840/B POR2X1_500/A POR2X1_205/A POR2X1_646/Y POR2X1_722/A POR2X1_540/Y POR2X1_181/Y POR2X1_782/A POR2X1_555/B POR2X1_649/B PAND2X1_241/Y PAND2X1_349/B PAND2X1_730/A PAND2X1_341/A PAND2X1_148/Y PAND2X1_467/Y PAND2X1_546/Y PAND2X1_794/B PAND2X1_653/Y PAND2X1_479/A PAND2X1_737/B PAND2X1_192/Y PAND2X1_324/Y PAND2X1_718/Y PAND2X1_714/A PAND2X1_388/Y PAND2X1_830/Y POR2X1_574/Y POR2X1_863/B POR2X1_730/Y POR2X1_550/Y POR2X1_339/Y POR2X1_724/A POR2X1_561/Y PAND2X1_345/Y PAND2X1_444/Y PAND2X1_140/A POR2X1_359/B PAND2X1_553/A 
+ PAND2X1_190/Y PAND2X1_193/Y PAND2X1_639/B PAND2X1_449/Y PAND2X1_793/Y PAND2X1_575/B POR2X1_805/B POR2X1_710/Y POR2X1_542/Y POR2X1_797/A POR2X1_523/Y POR2X1_639/A POR2X1_228/Y POR2X1_551/A POR2X1_728/B PAND2X1_852/B PAND2X1_244/B PAND2X1_476/A POR2X1_812/B POR2X1_362/Y POR2X1_476/Y PAND2X1_660/B PAND2X1_218/A POR2X1_712/Y POR2X1_651/Y POR2X1_717/Y POR2X1_795/B POR2X1_566/B POR2X1_149/Y POR2X1_353/Y POR2X1_731/A POR2X1_851/A POR2X1_783/Y POR2X1_477/A POR2X1_840/Y POR2X1_794/B POR2X1_773/A POR2X1_724/B POR2X1_350/B PAND2X1_555/Y PAND2X1_658/B POR2X1_679/Y PAND2X1_137/Y PAND2X1_768/Y PAND2X1_403/B PAND2X1_805/A PAND2X1_474/A PAND2X1_723/A PAND2X1_303/Y PAND2X1_564/B PAND2X1_787/Y 
+ POR2X1_862/A POR2X1_550/B POR2X1_720/Y POR2X1_508/A POR2X1_349/Y POR2X1_788/A PAND2X1_850/Y PAND2X1_242/Y POR2X1_647/Y PAND2X1_620/Y PAND2X1_206/B PAND2X1_182/B PAND2X1_552/A PAND2X1_336/Y PAND2X1_785/A PAND2X1_771/B PAND2X1_139/Y PAND2X1_857/A POR2X1_463/Y PAND2X1_854/Y PAND2X1_568/B POR2X1_348/A POR2X1_623/A POR2X1_341/A PAND2X1_561/Y POR2X1_402/A POR2X1_241/Y POR2X1_715/A PAND2X1_348/Y PAND2X1_466/A PAND2X1_795/B PAND2X1_206/A PAND2X1_734/B POR2X1_208/Y POR2X1_337/Y PAND2X1_842/Y PAND2X1_205/A PAND2X1_214/B PAND2X1_796/B PAND2X1_352/B POR2X1_713/Y POR2X1_711/Y POR2X1_624/Y PAND2X1_650/A PAND2X1_563/A PAND2X1_853/B PAND2X1_346/Y PAND2X1_569/B POR2X1_356/Y POR2X1_453/Y POR2X1_140/B 
+ POR2X1_192/Y POR2X1_137/Y POR2X1_850/B POR2X1_190/Y POR2X1_788/Y POR2X1_661/B POR2X1_479/B POR2X1_737/A POR2X1_141/A POR2X1_771/A POR2X1_193/Y POR2X1_718/A POR2X1_558/Y POR2X1_440/Y POR2X1_61/Y POR2X1_347/A POR2X1_84/Y POR2X1_830/Y PAND2X1_844/B PAND2X1_623/Y PAND2X1_501/B PAND2X1_61/Y PAND2X1_402/B PAND2X1_840/A PAND2X1_499/Y PAND2X1_556/B PAND2X1_643/Y PAND2X1_84/Y POR2X1_562/B POR2X1_439/Y POR2X1_180/Y POR2X1_853/A POR2X1_175/A POR2X1_544/Y POR2X1_203/Y POR2X1_573/A POR2X1_675/Y POR2X1_123/Y POR2X1_835/Y POR2X1_169/Y POR2X1_191/Y POR2X1_650/A POR2X1_786/Y POR2X1_444/Y POR2X1_390/B POR2X1_703/Y POR2X1_337/A POR2X1_722/B POR2X1_201/Y POR2X1_623/Y POR2X1_500/Y 
+ POR2X1_643/Y PAND2X1_341/B PAND2X1_558/Y PAND2X1_140/Y PAND2X1_792/B PAND2X1_711/B PAND2X1_647/B PAND2X1_652/A PAND2X1_493/Y PAND2X1_715/B PAND2X1_205/B PAND2X1_602/Y PAND2X1_713/A PAND2X1_347/Y PAND2X1_124/Y PAND2X1_782/Y PAND2X1_563/B PAND2X1_213/A PAND2X1_731/A PAND2X1_639/Y POR2X1_802/B POR2X1_802/A PAND2X1_802/B PAND2X1_798/Y POR2X1_567/A PAND2X1_539/Y PAND2X1_810/A POR2X1_510/Y PAND2X1_657/B POR2X1_774/Y POR2X1_35/Y PAND2X1_35/Y PAND2X1_455/Y PAND2X1_404/Y POR2X1_465/B POR2X1_404/Y PAND2X1_267/Y PAND2X1_631/A PAND2X1_798/B POR2X1_652/A POR2X1_631/B POR2X1_468/B POR2X1_319/Y PAND2X1_593/Y POR2X1_267/Y PAND2X1_354/A 
+ VSS VDD 
+ GATE_222 GATE_366 GATE_479 GATE_579 GATE_662 GATE_741 GATE_811 GATE_865 D_GATE_222 D_GATE_366 D_GATE_479 D_GATE_579 D_GATE_662 D_GATE_741 D_GATE_811 D_GATE_865 
+ AES_SBOX_3

.include outputs_2.plw

* **************************************
* --- Simulation Settings ---
* **************************************

.param SIM_LEN = 35ns
.csparam SIM_LEN = {SIM_LEN}

.tran 0.1ns 'SIM_LEN'
.param SIMSTEP = 'SIM_LEN/0.1ns'
.csparam SIMSTEP = {SIMSTEP}

* **************************************
* --- Simulation Control ---
* **************************************

.control
    .include ../inputsD.inc

    run
    
    if ('writeFile' > 0)   
      wrdata ivdd_3.out i(vvdd)
      wrdata ivss_3.out i(vvss)
      *snsave sim_3.snap
    end
    
    set wr_vecnames
    set wr_singlescale
    wrdata outputs_3.out V("GATE_222") V("GATE_366") V("GATE_479") V("GATE_579") V("GATE_662") V("GATE_741") V("GATE_811") V("GATE_865") V("D_GATE_222") V("D_GATE_366") V("D_GATE_479") V("D_GATE_579") V("D_GATE_662") V("D_GATE_741") V("D_GATE_811") V("D_GATE_865") 
    
    if ('showPlots' < 1)
        quit
    end
       
.endc

.end
