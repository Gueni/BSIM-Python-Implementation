* SPICE3 subcircuits originally created by qflow ...

.include tsmc180nmcmos.lib

VVDD VDDR 0 1.8V
R_VDD VDDR VDD 0.001
VVSS VSS 0 0V

.global VDD VSS 

.subckt MODEL_INV1X1 Y VSS A VDD
M1000 Y A VDD VDD TSMC180nmP w=2u l=0.2u
+  ad=1p pd=5u as=1p ps=5u
M1001 Y A VSS VSS TSMC180nmN w=1u l=0.2u
+  ad=0.5p pd=3u as=0.5p ps=3u
C0 Y A 0.08fF
C1 Y VDD 0.39fF
C2 A VDD 0.20fF
C3 VSS Y 0.16fF
C4 VSS A 0.05fF
C5 VSS VSS 0.12fF
C6 Y VSS 0.14fF
C7 A VSS 0.31fF
C8 VDD VSS 1.52fF
.ends

.subckt MODEL_NOR2X1 Y VSS A B a_36_216# VDD
M1000 a_36_216# A VDD VDD TSMC180nmP w=4u l=0.2u
+  ad=1.2p pd=8.6u as=2p ps=9u
M1001 Y B a_36_216# VDD TSMC180nmP w=4u l=0.2u
+  ad=2p pd=9u as=0p ps=0u
M1002 Y A VSS VSS TSMC180nmN w=1u l=0.2u
+  ad=0.6p pd=3.2u as=1p ps=6u
M1003 VSS B Y VSS TSMC180nmN w=1u l=0.2u
+  ad=0p pd=0u as=0p ps=0u
C0 B A 0.18fF
C1 B VDD 0.12fF
C2 A VDD 0.07fF
C3 VSS Y 0.26fF
C4 Y a_36_216# 0.01fF
C5 Y B 0.12fF
C6 VSS A 0.05fF
C7 Y A 0.07fF
C8 Y VDD 0.17fF
C9 VSS VSS 0.18fF
C10 Y VSS 0.12fF
C11 B VSS 0.28fF
C12 A VSS 0.31fF
C13 VDD VSS 1.73fF
.ends

.subckt MODEL_NAND2X1 Y VSS A B a_36_24# VDD
M1000 Y A VDD VDD TSMC180nmP w=2u l=0.2u
+  ad=1.2p pd=5.2u as=2p ps=10u
M1001 VDD B Y VDD TSMC180nmP w=2u l=0.2u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_36_24# A VSS VSS TSMC180nmN w=2u l=0.2u
+  ad=0.6p pd=4.6u as=1p ps=5u
M1003 Y B a_36_24# VSS TSMC180nmN w=2u l=0.2u
+  ad=1p pd=5u as=0p ps=0u
C0 Y VDD 0.57fF
C1 B A 0.22fF
C2 B VDD 0.27fF
C3 A VDD 0.20fF
C4 a_36_24# Y 0.01fF
C5 VSS Y 0.09fF
C6 Y B 0.10fF
C7 VSS A 0.05fF
C8 Y A 0.08fF
C9 VSS VSS 0.17fF
C10 Y VSS 0.11fF
C11 B VSS 0.19fF
C12 A VSS 0.25fF
C13 VDD VSS 1.73fF
.ends

.subckt MODEL_NAND2X1_SC1 Y VSS A B a_36_24# VDD
M1000 Y A VDD VDD TSMC180nmP w=2u l=0.2u
+  ad=1.2p pd=5.2u as=2p ps=10u
M1001 VDD B Y VDD TSMC180nmP w=2u l=0.2u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_36_24# A VSS VSS TSMC180nmN w=2u l=0.2u
+  ad=0.6p pd=4.6u as=1p ps=5u
M1003 Y B a_36_24# VSS TSMC180nmN w=2u l=0.2u
+  ad=1p pd=5u as=0p ps=0u
C0 Y VDD 0.57fF
C1 B A 0.22fF
C2 B VDD 0.27fF
C3 A VDD 0.20fF
C4 a_36_24# Y 0.01fF
C5 VSS Y 0.09fF
C6 Y B 0.10fF
C7 VSS A 0.05fF
C8 Y A 0.08fF
C9 VSS VSS 0.17fF
C10 Y VSS 0.11fF
C11 B VSS 0.19fF
C12 A VSS 0.25fF
C13 VDD VSS 1.73fF

R_FAULT Y VDD 1

.ends


* Simulation

.options TEMP = 25°C
.options TNOM = 25°C
.ic 
.tran 5e-12s 5e-08s 0s uic

* Place circuit netlist generated by TSaCt2 here!


