magic
tech scmos
timestamp 1612034806
<< nwell >>
rect -15 48 100 105
<< ntransistor >>
rect 13 7 15 11
rect 21 7 23 11
rect 29 7 31 11
rect 34 7 36 11
rect 42 7 44 27
rect 58 7 60 11
rect 74 7 76 42
rect 82 7 84 27
<< ptransistor >>
rect 8 89 10 93
rect 13 89 15 93
rect 21 89 23 93
rect 26 89 28 93
rect 34 77 36 93
rect 42 77 44 93
rect 58 54 60 93
rect 74 89 76 93
rect 82 54 84 93
<< ndiffusion >>
rect 12 7 13 11
rect 15 7 16 11
rect 20 7 21 11
rect 23 7 24 11
rect 28 7 29 11
rect 31 7 34 11
rect 36 7 37 11
rect 41 7 42 27
rect 44 7 45 27
rect 57 7 58 11
rect 60 7 61 11
rect 73 7 74 42
rect 76 7 77 42
rect 81 7 82 27
rect 84 7 85 27
<< pdiffusion >>
rect 7 89 8 93
rect 10 89 13 93
rect 15 89 16 93
rect 20 89 21 93
rect 23 89 26 93
rect 28 89 29 93
rect 33 77 34 93
rect 36 77 37 93
rect 41 77 42 93
rect 44 77 45 93
rect 57 54 58 93
rect 60 54 61 93
rect 73 89 74 93
rect 76 89 77 93
rect 81 54 82 93
rect 84 54 85 93
<< ndcontact >>
rect 8 7 12 11
rect 16 7 20 11
rect 24 7 28 11
rect 37 7 41 27
rect 45 7 49 27
rect 53 7 57 11
rect 61 7 65 11
rect 69 7 73 42
rect 77 7 81 42
rect 85 7 89 27
<< pdcontact >>
rect 3 89 7 93
rect 16 89 20 93
rect 29 77 33 93
rect 37 77 41 93
rect 45 77 49 93
rect 53 54 57 93
rect 61 54 65 93
rect 69 89 73 93
rect 77 54 81 93
rect 85 54 89 93
<< psubstratepcontact >>
rect -1 -2 3 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect -1 98 3 102
rect 37 98 41 102
<< polysilicon >>
rect 8 93 10 95
rect 13 93 15 95
rect 21 93 23 95
rect 26 93 28 95
rect 34 93 36 95
rect 42 93 44 95
rect 58 93 60 95
rect 74 93 76 95
rect 82 93 84 95
rect 8 53 10 89
rect 13 41 15 89
rect 21 53 23 89
rect 18 49 19 53
rect 13 11 15 37
rect 21 11 23 49
rect 26 41 28 89
rect 34 57 36 77
rect 42 50 44 77
rect 58 50 60 54
rect 34 48 60 50
rect 34 27 36 48
rect 58 44 59 48
rect 42 41 51 43
rect 42 27 44 41
rect 29 25 36 27
rect 29 11 31 25
rect 34 11 36 25
rect 58 11 60 44
rect 74 42 76 89
rect 82 49 84 54
rect 83 45 84 49
rect 82 27 84 45
rect 13 5 15 7
rect 21 5 23 7
rect 29 5 31 7
rect 34 5 36 7
rect 42 5 44 7
rect 58 5 60 7
rect 74 2 76 7
rect 82 5 84 7
<< polycontact >>
rect 6 49 10 53
rect 19 49 23 53
rect 13 37 17 41
rect 34 53 38 57
rect 26 37 30 41
rect 59 44 63 48
rect 51 39 55 43
rect 79 45 83 49
rect 73 -2 77 2
<< metal1 >>
rect -1 102 94 103
rect 3 98 37 102
rect 41 98 94 102
rect -1 97 94 98
rect 37 93 41 97
rect 61 93 65 97
rect 77 93 81 97
rect 3 88 7 89
rect 16 64 20 89
rect 45 64 49 77
rect 16 60 49 64
rect 8 53 12 57
rect 10 49 19 53
rect 27 49 31 60
rect 52 57 53 93
rect 38 54 53 57
rect 38 53 56 54
rect 27 45 34 49
rect 17 37 26 41
rect 13 33 20 37
rect 34 27 38 45
rect 52 43 56 53
rect 69 48 73 89
rect 89 54 90 93
rect 63 44 73 48
rect 78 45 79 49
rect 55 39 56 43
rect 8 23 37 27
rect 8 11 12 23
rect 24 11 28 23
rect 52 11 56 39
rect 69 42 73 44
rect 52 7 53 11
rect 86 27 90 54
rect 89 7 90 27
rect 16 3 20 7
rect 45 3 49 7
rect 61 3 65 7
rect 77 3 81 7
rect -1 2 94 3
rect 3 -2 26 2
rect 30 -2 73 2
rect 77 -2 94 2
rect -1 -3 94 -2
<< m2contact >>
rect 3 89 7 93
rect 29 89 33 93
rect 34 45 38 49
rect 79 45 83 49
<< metal2 >>
rect 7 89 29 93
rect 38 45 79 49
<< metal4 >>
rect 61 -1 67 3
<< labels >>
rlabel space -8 -3 99 105 1 vdd
rlabel space -8 -3 99 105 1 gnd
rlabel ptransistor 58 82 58 82 1 D$
rlabel ptransistor 60 82 60 82 1 S$
rlabel metal1 54 26 54 26 1 CTRL2
rlabel ntransistor 58 9 58 9 1 D$
rlabel ntransistor 60 9 60 9 1 S$
rlabel ntransistor 82 17 82 17 1 S$
rlabel ntransistor 84 17 84 17 1 D$
rlabel ptransistor 82 92 82 92 1 S$
rlabel ptransistor 84 92 84 92 1 D$
rlabel metal1 90 62 90 66 1 Y
port 5 n signal output
rlabel ptransistor 76 92 76 92 1 S$
rlabel ptransistor 74 92 74 92 1 D$
rlabel ntransistor 74 16 74 16 1 D$
rlabel ntransistor 76 16 76 16 1 S$
rlabel metal1 71 70 71 70 1 CTRL
rlabel metal1 8 53 8 57 1 B
port 3 n signal input
rlabel metal1 29 62 29 62 1 O
rlabel metal1 9 0 9 0 1 GND!
port 2 n power bidirectional
rlabel metal1 16 100 16 100 1 VDD!
port 1 n power bidirectional
rlabel metal1 13 33 13 37 1 A
port 4 n signal input
rlabel ptransistor 23 90 23 90 1 S$
rlabel ptransistor 21 90 21 90 1 D$
rlabel ptransistor 15 90 15 90 1 D$
rlabel ptransistor 13 90 13 90 1 S$
rlabel ptransistor 10 90 10 90 1 D$
rlabel ptransistor 8 90 8 90 1 S$
rlabel ptransistor 26 90 26 90 1 D$
rlabel ptransistor 28 90 28 90 1 S$
rlabel ptransistor 44 78 44 78 1 D$
rlabel ptransistor 42 78 42 78 1 S$
rlabel ptransistor 36 78 36 78 1 S$
rlabel ptransistor 34 78 34 78 1 D$
rlabel space -15 -3 100 105 1 vdd
rlabel space -15 -3 100 105 1 gnd
rlabel ntransistor 42 10 42 10 1 D$
rlabel ntransistor 44 9 44 9 1 S$
rlabel ntransistor 34 10 34 10 1 S$
rlabel ntransistor 36 9 36 9 1 D$
rlabel ntransistor 29 10 29 10 1 S$
rlabel ntransistor 31 9 31 9 1 D$
rlabel ntransistor 21 10 21 10 1 S$
rlabel ntransistor 23 9 23 9 1 D$
rlabel ntransistor 13 10 13 10 1 D$
rlabel ntransistor 15 9 15 9 1 S$
<< end >>
