magic
tech scmos
timestamp 1597936220
<< nwell >>
rect 0 50 104 107
<< ntransistor >>
rect 25 10 27 20
rect 30 10 32 20
rect 35 10 37 20
rect 43 10 45 20
rect 48 10 50 20
rect 53 10 55 20
rect 83 9 85 29
rect 91 9 93 29
<< ptransistor >>
rect 11 76 13 96
rect 27 72 29 96
rect 35 72 37 96
rect 43 72 45 96
rect 51 72 53 96
rect 67 76 69 96
rect 83 92 85 96
rect 91 56 93 96
<< ndiffusion >>
rect 24 10 25 20
rect 27 10 30 20
rect 32 10 35 20
rect 37 10 38 20
rect 42 10 43 20
rect 45 10 48 20
rect 50 10 53 20
rect 55 10 56 20
rect 82 9 83 29
rect 85 9 86 29
rect 90 9 91 29
rect 93 9 94 29
<< pdiffusion >>
rect 10 80 11 96
rect 6 76 11 80
rect 13 92 18 96
rect 13 76 14 92
rect 26 72 27 96
rect 29 92 35 96
rect 29 72 30 92
rect 34 72 35 92
rect 37 80 38 96
rect 42 80 43 96
rect 37 76 43 80
rect 37 72 38 76
rect 42 72 43 76
rect 45 92 51 96
rect 45 72 46 92
rect 50 72 51 92
rect 53 72 54 96
rect 62 92 67 96
rect 66 76 67 92
rect 69 80 70 96
rect 82 92 83 96
rect 85 92 86 96
rect 69 76 74 80
rect 90 56 91 96
rect 93 56 94 96
<< ndcontact >>
rect 20 10 24 20
rect 38 10 42 20
rect 56 10 60 20
rect 78 9 82 29
rect 86 9 90 29
rect 94 9 98 29
<< pdcontact >>
rect 6 80 10 96
rect 14 76 18 92
rect 22 72 26 96
rect 30 72 34 92
rect 38 80 42 96
rect 38 72 42 76
rect 46 72 50 92
rect 54 72 58 96
rect 62 76 66 92
rect 70 80 74 96
rect 78 92 82 96
rect 86 56 90 96
rect 94 56 98 96
<< psubstratepcontact >>
rect 7 1 11 5
rect 16 1 21 5
rect 28 1 32 5
rect 51 1 55 5
rect 62 1 66 5
rect 72 1 76 5
rect 94 1 98 5
<< nsubstratencontact >>
rect 3 100 7 104
rect 22 100 26 104
rect 38 100 42 104
rect 54 100 58 104
rect 70 100 74 104
rect 86 100 90 104
rect 97 100 101 104
<< polysilicon >>
rect 11 96 13 98
rect 27 96 29 98
rect 35 96 37 98
rect 43 96 45 98
rect 51 96 53 98
rect 67 96 69 98
rect 83 96 85 98
rect 91 96 93 98
rect 11 73 13 76
rect 10 69 13 73
rect 67 73 69 76
rect 27 69 29 72
rect 35 68 37 72
rect 33 65 37 68
rect 43 68 45 72
rect 51 69 53 72
rect 67 69 70 73
rect 43 65 47 68
rect 33 50 35 65
rect 32 46 35 50
rect 25 20 27 39
rect 30 20 32 46
rect 39 33 41 54
rect 45 43 47 65
rect 45 39 46 43
rect 35 31 45 33
rect 35 20 37 31
rect 43 20 45 31
rect 48 20 50 39
rect 53 20 55 46
rect 83 29 85 92
rect 91 40 93 56
rect 92 36 93 40
rect 91 29 93 36
rect 25 7 27 10
rect 30 7 32 10
rect 35 7 37 10
rect 43 7 45 10
rect 48 7 50 10
rect 53 7 55 10
rect 83 5 85 9
rect 91 7 93 9
<< polycontact >>
rect 6 69 10 73
rect 26 65 30 69
rect 70 69 74 73
rect 50 65 54 69
rect 38 54 42 58
rect 28 46 32 50
rect 23 39 27 43
rect 51 46 55 50
rect 46 39 50 43
rect 88 36 92 40
rect 82 1 86 5
<< metal1 >>
rect 2 104 102 105
rect 2 100 3 104
rect 7 100 22 104
rect 26 100 38 104
rect 42 100 54 104
rect 58 100 70 104
rect 74 100 86 104
rect 90 100 97 104
rect 101 100 102 104
rect 2 99 102 100
rect 22 96 26 99
rect 54 96 58 99
rect 86 96 90 99
rect 6 58 10 69
rect 70 58 74 69
rect 78 58 82 92
rect 6 54 38 58
rect 42 54 82 58
rect 98 56 99 59
rect 32 46 51 50
rect 27 39 46 43
rect 78 29 82 54
rect 87 36 88 40
rect 95 29 99 56
rect 18 23 62 27
rect 20 20 24 23
rect 56 20 60 23
rect 38 6 42 10
rect 98 26 99 29
rect 86 6 90 9
rect 6 5 99 6
rect 6 1 7 5
rect 11 1 16 5
rect 21 1 28 5
rect 32 1 38 5
rect 42 1 51 5
rect 55 1 62 5
rect 66 1 72 5
rect 76 1 82 5
rect 86 1 94 5
rect 98 1 99 5
rect 6 0 99 1
<< m2contact >>
rect 6 76 10 80
rect 14 92 18 96
rect 30 92 34 96
rect 38 76 42 80
rect 46 92 50 96
rect 62 92 66 96
rect 70 76 74 80
rect 26 61 30 65
rect 50 61 54 65
rect 88 36 92 40
rect 14 23 18 27
rect 62 23 66 27
rect 38 1 42 5
<< metal2 >>
rect 18 92 30 96
rect 34 92 46 96
rect 50 92 62 96
rect 10 76 38 80
rect 42 76 70 80
rect 14 27 18 76
rect 30 61 50 65
rect 38 5 42 61
rect 62 40 66 76
rect 62 36 88 40
rect 62 27 66 36
rect 38 0 42 1
<< labels >>
rlabel metal1 72 56 72 56 1 CTRL
rlabel metal1 46 3 46 3 1 GND!
port 5 n ground bidirectional
rlabel metal1 34 102 34 102 1 VDD!
port 4 n power bidirectional
rlabel pdcontact 64 86 64 86 1 VVDD
rlabel ndiffusion 33 18 33 18 1 VGND1
rlabel ndiffusion 46 18 46 18 1 VGND2
rlabel ntransistor 83 19 83 19 1 D$
rlabel ntransistor 85 19 85 19 1 S$
rlabel ptransistor 85 94 85 94 1 S$
rlabel ptransistor 83 94 83 94 1 D$
rlabel polycontact 23 39 23 43 1 A
port 2 n signal input
rlabel polycontact 28 46 28 50 1 B
port 1 n signal input
rlabel ntransistor 45 15 45 15 1 D$
rlabel ntransistor 50 15 50 15 1 D$
rlabel ntransistor 55 15 55 15 1 D$
rlabel ntransistor 35 15 35 15 1 D$
rlabel ntransistor 30 15 30 15 1 D$
rlabel ntransistor 25 15 25 15 1 D$
rlabel ntransistor 53 15 53 15 1 S$
rlabel ntransistor 48 15 48 15 1 S$
rlabel ntransistor 43 15 43 15 1 S$
rlabel ntransistor 37 15 37 15 1 S$
rlabel ntransistor 32 15 32 15 1 S$
rlabel ntransistor 27 15 27 15 1 S$
rlabel ntransistor 93 19 93 19 1 D$
rlabel ntransistor 91 19 91 19 1 S$
rlabel ptransistor 93 94 93 94 1 D$
rlabel ptransistor 91 94 91 94 1 S$
rlabel ptransistor 69 87 69 87 1 D$
rlabel ptransistor 51 87 51 87 1 D$
rlabel ptransistor 29 87 29 87 1 D$
rlabel ptransistor 43 87 43 87 1 D$
rlabel ptransistor 37 87 37 87 1 D$
rlabel ptransistor 11 88 11 88 1 D$
rlabel ptransistor 67 87 67 87 1 S$
rlabel ptransistor 53 87 53 87 1 S$
rlabel ptransistor 45 87 45 87 1 S$
rlabel ptransistor 35 87 35 87 1 S$
rlabel ptransistor 27 87 27 87 1 S$
rlabel ptransistor 13 88 13 88 1 S$
rlabel space 0 0 104 107 1 vdd
rlabel space 0 0 104 107 1 gnd
rlabel metal2 63 77 63 77 1 O
rlabel metal2 64 34 64 34 1 O
rlabel metal1 99 40 99 44 1 Y
port 3 n signal output
<< end >>
