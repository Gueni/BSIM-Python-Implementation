* SPICE3 file created from dualRail.ext - technology: scmos

.subckt POR2X1 VDD GND B A Y m4_208_n4# O CTRL2 a_16_28# CTRL a_76_344# a_56_344#
X0 a_16_28# A GND GND NMOS_MAGIC ad=0.44p pd=3.8u as=3.39p ps=17u w=0.4u l=0.2u
**devattr s=S d=D
X1 O CTRL VDD VDD PMOS_MAGIC ad=1.72p pd=7.8u as=5.94p ps=27.8u w=3.3u l=0.2u
**devattr s=S d=D
X2 CTRL GND GND GND NMOS_MAGIC ad=1.75p pd=8u as=0p ps=0u w=3.5u l=0.2u
**devattr s=S d=D
X3 a_56_344# B VDD VDD PMOS_MAGIC ad=0.21p pd=2u as=0p ps=0u w=0.7u l=0.2u
**devattr s=S d=D
X4 Y O GND GND NMOS_MAGIC ad=1p pd=5u as=0p ps=0u w=2u l=0.2u
**devattr s=S d=D
X5 Y O VDD VDD PMOS_MAGIC ad=1.95p pd=8.8u as=0p ps=0u w=3.9u l=0.2u
**devattr s=S d=D
X6 CTRL2 CTRL GND GND NMOS_MAGIC ad=0.2p pd=1.8u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X7 O CTRL2 a_76_344# VDD PMOS_MAGIC ad=0p pd=0u as=0.42p ps=2.6u w=0.7u l=0.2u
**devattr s=S d=D
X8 CTRL GND VDD VDD PMOS_MAGIC ad=0.2p pd=1.8u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X9 O CTRL a_16_28# GND NMOS_MAGIC ad=1.04p pd=5.2u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X10 a_76_344# A a_56_344# VDD PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=0.7u l=0.2u
**devattr s=S d=D
X11 a_16_28# B GND GND NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X12 CTRL2 CTRL VDD VDD PMOS_MAGIC ad=1.95p pd=8.8u as=0p ps=0u w=3.9u l=0.2u
**devattr s=S d=D
X13 O CTRL2 GND GND NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=2u l=0.2u
**devattr s=S d=D
C0 O A 0.13fF
C1 a_16_28# B 0.02fF
C2 O Y 0.05fF
C3 O a_76_344# 0.07fF
C4 a_16_28# A 0.10fF
C5 VDD B 0.36fF
C6 O a_16_28# 0.21fF
C7 CTRL2 VDD 1.37fF
C8 CTRL VDD 1.32fF
C9 VDD A 0.28fF
C10 O VDD 0.59fF
C11 B A 0.47fF
C12 VDD Y 0.54fF
C13 O B 0.08fF
C14 CTRL2 CTRL 0.32fF
C15 CTRL2 A 0.13fF
C16 a_76_344# VDD 0.05fF
C17 CTRL2 O 0.27fF
C18 CTRL A 0.16fF
C19 CTRL O 0.15fF
C20 Y 0 0.50fF
C21 A 0 0.35fF
C22 B 0 0.27fF
C23 VDD 0 4.59fF
C24 GND 0 -0.16fF
C25 m4_208_n4# 0 0.01fF
C26 a_16_28# 0 0.33fF
C27 a_76_344# 0 0.00fF
C28 O 0 0.33fF
C29 CTRL 0 0.70fF
C30 CTRL2 0 0.39fF
.ends

.subckt PAND2X1 VDD GND B A Y a_16_344# m4_208_n4# O a_56_28# CTRL2 CTRL a_76_28#
X0 a_56_28# A a_76_28# GND NMOS_MAGIC ad=0.15p pd=1.6u as=0.3p ps=2.2u w=0.5u l=0.2u
**devattr s=S d=D
X1 CTRL GND GND GND NMOS_MAGIC ad=1.75p pd=8u as=3.22p ps=15.2u w=3.5u l=0.2u
**devattr s=S d=D
X2 O B a_16_344# VDD PMOS_MAGIC ad=1.72p pd=8.8u as=0.77p ps=5u w=0.7u l=0.2u
**devattr s=S d=D
X3 Y O GND GND NMOS_MAGIC ad=1.1p pd=5.4u as=0p ps=0u w=2.2u l=0.2u
**devattr s=S d=D
X4 Y O VDD VDD PMOS_MAGIC ad=1.95p pd=8.8u as=5.31p ps=24.2u w=3.9u l=0.2u
**devattr s=S d=D
X5 CTRL2 CTRL GND GND NMOS_MAGIC ad=0.2p pd=1.8u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X6 a_16_344# CTRL2 VDD VDD PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=0.7u l=0.2u
**devattr s=S d=D
X7 CTRL GND VDD VDD PMOS_MAGIC ad=0.2p pd=1.8u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X8 a_76_28# CTRL GND GND NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=0.5u l=0.2u
**devattr s=S d=D
X9 O A a_16_344# VDD PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=0.7u l=0.2u
**devattr s=S d=D
X10 O B a_56_28# GND NMOS_MAGIC ad=1.25p pd=7u as=0p ps=0u w=0.5u l=0.2u
**devattr s=S d=D
X11 CTRL2 CTRL VDD VDD PMOS_MAGIC ad=1.95p pd=8.8u as=0p ps=0u w=3.9u l=0.2u
**devattr s=S d=D
X12 O CTRL VDD VDD PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=2.6u l=0.2u
**devattr s=S d=D
X13 O CTRL2 GND GND NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=2u l=0.2u
**devattr s=S d=D
C0 O A 0.17fF
C1 a_76_28# B 0.01fF
C2 O Y 0.05fF
C3 a_16_344# A 0.01fF
C4 O a_16_344# 0.17fF
C5 a_76_28# A 0.01fF
C6 VDD B 0.36fF
C7 O a_76_28# 0.05fF
C8 CTRL2 VDD 0.86fF
C9 a_56_28# a_76_28# 0.00fF
C10 CTRL VDD 1.37fF
C11 VDD A 0.28fF
C12 O VDD 0.78fF
C13 B A 0.49fF
C14 VDD Y 0.54fF
C15 a_16_344# VDD 0.19fF
C16 O B 0.13fF
C17 CTRL2 CTRL 0.34fF
C18 CTRL2 A 0.13fF
C19 a_16_344# B 0.01fF
C20 CTRL2 O 1.20fF
C21 CTRL A 0.16fF
C22 CTRL O 0.19fF
C23 Y 0 0.50fF
C24 A 0 0.34fF
C25 B 0 0.27fF
C26 VDD 0 4.59fF
C27 GND 0 -0.15fF
C28 m4_208_n4# 0 0.01fF
C29 a_76_28# 0 0.02fF
C30 a_16_344# 0 -0.00fF
C31 O 0 0.47fF
C32 CTRL 0 0.70fF
C33 CTRL2 0 0.39fF
.ends

.subckt dualRail INPUT_0 D_INPUT_0 INPUT_1 D_INPUT_1 INPUT_2 D_INPUT_2 INPUT_3 D_INPUT_3
+ INPUT_4 D_INPUT_4 INPUT_5 D_INPUT_5 INPUT_6 D_INPUT_6 INPUT_7 D_INPUT_7 D_GATE_222
+ D_GATE_366 D_GATE_479 D_GATE_579 D_GATE_662 D_GATE_741 D_GATE_811 D_GATE_865 GATE_222
+ GATE_366 GATE_479 GATE_579 GATE_662 GATE_741 GATE_811 GATE_865 gate type: AND; name:
+ GATE_0_I0
XPOR2X1_717 VDD GND POR2X1_717/B POR2X1_558/B POR2X1_717/Y POR2X1_717/m4_208_n4# POR2X1_717/O
+ POR2X1_717/CTRL2 POR2X1_717/a_16_28# POR2X1_717/CTRL POR2X1_717/a_76_344# POR2X1_717/a_56_344#
+ POR2X1
XPOR2X1_706 VDD GND POR2X1_706/B POR2X1_706/A POR2X1_713/A POR2X1_706/m4_208_n4# POR2X1_706/O
+ POR2X1_706/CTRL2 POR2X1_706/a_16_28# POR2X1_706/CTRL POR2X1_706/a_76_344# POR2X1_706/a_56_344#
+ POR2X1
XPOR2X1_728 VDD GND POR2X1_728/B POR2X1_728/A POR2X1_730/B POR2X1_728/m4_208_n4# POR2X1_728/O
+ POR2X1_728/CTRL2 POR2X1_728/a_16_28# POR2X1_728/CTRL POR2X1_728/a_76_344# POR2X1_728/a_56_344#
+ POR2X1
XPOR2X1_739 VDD GND POR2X1_192/Y POR2X1_730/Y POR2X1_740/A POR2X1_739/m4_208_n4# POR2X1_739/O
+ POR2X1_739/CTRL2 POR2X1_739/a_16_28# POR2X1_739/CTRL POR2X1_739/a_76_344# POR2X1_739/a_56_344#
+ POR2X1
XPOR2X1_514 VDD GND INPUT_0 POR2X1_138/A POR2X1_514/Y POR2X1_514/m4_208_n4# POR2X1_514/O
+ POR2X1_514/CTRL2 POR2X1_514/a_16_28# POR2X1_514/CTRL POR2X1_514/a_76_344# POR2X1_514/a_56_344#
+ POR2X1
XPOR2X1_503 VDD GND POR2X1_65/A POR2X1_503/A POR2X1_503/Y POR2X1_503/m4_208_n4# POR2X1_503/O
+ POR2X1_503/CTRL2 POR2X1_503/a_16_28# POR2X1_503/CTRL POR2X1_503/a_76_344# POR2X1_503/a_56_344#
+ POR2X1
XPOR2X1_525 VDD GND POR2X1_41/B POR2X1_52/A POR2X1_525/Y POR2X1_525/m4_208_n4# POR2X1_525/O
+ POR2X1_525/CTRL2 POR2X1_525/a_16_28# POR2X1_525/CTRL POR2X1_525/a_76_344# POR2X1_525/a_56_344#
+ POR2X1
XPOR2X1_547 VDD GND POR2X1_547/B POR2X1_620/B POR2X1_550/A POR2X1_547/m4_208_n4# POR2X1_547/O
+ POR2X1_547/CTRL2 POR2X1_547/a_16_28# POR2X1_547/CTRL POR2X1_547/a_76_344# POR2X1_547/a_56_344#
+ POR2X1
XPOR2X1_536 VDD GND POR2X1_13/A POR2X1_102/Y POR2X1_536/Y POR2X1_536/m4_208_n4# POR2X1_536/O
+ POR2X1_536/CTRL2 POR2X1_536/a_16_28# POR2X1_536/CTRL POR2X1_536/a_76_344# POR2X1_536/a_56_344#
+ POR2X1
XPOR2X1_569 VDD GND POR2X1_564/Y POR2X1_569/A POR2X1_569/Y POR2X1_569/m4_208_n4# POR2X1_569/O
+ POR2X1_569/CTRL2 POR2X1_569/a_16_28# POR2X1_569/CTRL POR2X1_569/a_76_344# POR2X1_569/a_56_344#
+ POR2X1
XPOR2X1_558 VDD GND POR2X1_558/B POR2X1_558/A POR2X1_558/Y POR2X1_558/m4_208_n4# POR2X1_558/O
+ POR2X1_558/CTRL2 POR2X1_558/a_16_28# POR2X1_558/CTRL POR2X1_558/a_76_344# POR2X1_558/a_56_344#
+ POR2X1
XPOR2X1_300 VDD GND POR2X1_60/A POR2X1_119/Y POR2X1_300/Y POR2X1_300/m4_208_n4# POR2X1_300/O
+ POR2X1_300/CTRL2 POR2X1_300/a_16_28# POR2X1_300/CTRL POR2X1_300/a_76_344# POR2X1_300/a_56_344#
+ POR2X1
XPOR2X1_333 VDD GND POR2X1_174/B POR2X1_333/A POR2X1_333/Y POR2X1_333/m4_208_n4# POR2X1_333/O
+ POR2X1_333/CTRL2 POR2X1_333/a_16_28# POR2X1_333/CTRL POR2X1_333/a_76_344# POR2X1_333/a_56_344#
+ POR2X1
XPOR2X1_344 VDD GND POR2X1_254/Y POR2X1_344/A POR2X1_344/Y POR2X1_344/m4_208_n4# POR2X1_344/O
+ POR2X1_344/CTRL2 POR2X1_344/a_16_28# POR2X1_344/CTRL POR2X1_344/a_76_344# POR2X1_344/a_56_344#
+ POR2X1
XPOR2X1_322 VDD GND POR2X1_57/A POR2X1_376/B POR2X1_322/Y POR2X1_322/m4_208_n4# POR2X1_322/O
+ POR2X1_322/CTRL2 POR2X1_322/a_16_28# POR2X1_322/CTRL POR2X1_322/a_76_344# POR2X1_322/a_56_344#
+ POR2X1
XPOR2X1_311 VDD GND POR2X1_83/B POR2X1_102/Y POR2X1_311/Y POR2X1_311/m4_208_n4# POR2X1_311/O
+ POR2X1_311/CTRL2 POR2X1_311/a_16_28# POR2X1_311/CTRL POR2X1_311/a_76_344# POR2X1_311/a_56_344#
+ POR2X1
XPOR2X1_355 VDD GND POR2X1_355/B POR2X1_355/A POR2X1_356/A POR2X1_355/m4_208_n4# POR2X1_355/O
+ POR2X1_355/CTRL2 POR2X1_355/a_16_28# POR2X1_355/CTRL POR2X1_355/a_76_344# POR2X1_355/a_56_344#
+ POR2X1
XPOR2X1_377 VDD GND POR2X1_7/B PAND2X1_94/A POR2X1_378/A POR2X1_377/m4_208_n4# POR2X1_377/O
+ POR2X1_377/CTRL2 POR2X1_377/a_16_28# POR2X1_377/CTRL POR2X1_377/a_76_344# POR2X1_377/a_56_344#
+ POR2X1
XPOR2X1_366 VDD GND POR2X1_362/Y POR2X1_366/A POR2X1_366/Y POR2X1_366/m4_208_n4# POR2X1_366/O
+ POR2X1_366/CTRL2 POR2X1_366/a_16_28# POR2X1_366/CTRL POR2X1_366/a_76_344# POR2X1_366/a_56_344#
+ POR2X1
XPOR2X1_399 VDD GND POR2X1_57/A POR2X1_399/A POR2X1_399/Y POR2X1_399/m4_208_n4# POR2X1_399/O
+ POR2X1_399/CTRL2 POR2X1_399/a_16_28# POR2X1_399/CTRL POR2X1_399/a_76_344# POR2X1_399/a_56_344#
+ POR2X1
XPOR2X1_388 VDD GND POR2X1_169/A POR2X1_180/B POR2X1_390/B POR2X1_388/m4_208_n4# POR2X1_388/O
+ POR2X1_388/CTRL2 POR2X1_388/a_16_28# POR2X1_388/CTRL POR2X1_388/a_76_344# POR2X1_388/a_56_344#
+ POR2X1
XPAND2X1_307 VDD GND POR2X1_305/Y POR2X1_304/Y PAND2X1_308/B PAND2X1_307/a_16_344#
+ PAND2X1_307/m4_208_n4# PAND2X1_307/O PAND2X1_307/a_56_28# PAND2X1_307/CTRL2 PAND2X1_307/CTRL
+ PAND2X1_307/a_76_28# PAND2X1
XPAND2X1_318 VDD GND POR2X1_316/Y POR2X1_315/Y PAND2X1_319/B PAND2X1_318/a_16_344#
+ PAND2X1_318/m4_208_n4# PAND2X1_318/O PAND2X1_318/a_56_28# PAND2X1_318/CTRL2 PAND2X1_318/CTRL
+ PAND2X1_318/a_76_28# PAND2X1
XPAND2X1_329 VDD GND POR2X1_596/A POR2X1_327/Y POR2X1_355/B PAND2X1_329/a_16_344#
+ POR2X1_149/m4_208_n4# PAND2X1_329/O PAND2X1_329/a_56_28# PAND2X1_329/CTRL2 PAND2X1_329/CTRL
+ PAND2X1_329/a_76_28# PAND2X1
XPAND2X1_841 VDD GND PAND2X1_841/B PAND2X1_831/Y PAND2X1_841/Y PAND2X1_841/a_16_344#
+ PAND2X1_841/m4_208_n4# PAND2X1_841/O PAND2X1_841/a_56_28# PAND2X1_841/CTRL2 PAND2X1_841/CTRL
+ PAND2X1_841/a_76_28# PAND2X1
XPAND2X1_830 VDD GND POR2X1_142/Y POR2X1_108/Y PAND2X1_830/Y PAND2X1_830/a_16_344#
+ PAND2X1_830/m4_208_n4# PAND2X1_830/O PAND2X1_830/a_56_28# PAND2X1_830/CTRL2 PAND2X1_830/CTRL
+ PAND2X1_830/a_76_28# PAND2X1
XPAND2X1_863 VDD GND PAND2X1_863/B PAND2X1_863/A PAND2X1_864/B PAND2X1_863/a_16_344#
+ PAND2X1_863/m4_208_n4# PAND2X1_863/O PAND2X1_863/a_56_28# PAND2X1_863/CTRL2 PAND2X1_863/CTRL
+ PAND2X1_863/a_76_28# PAND2X1
XPAND2X1_852 VDD GND PAND2X1_852/B PAND2X1_852/A PAND2X1_857/A PAND2X1_852/a_16_344#
+ POR2X1_821/m4_208_n4# PAND2X1_852/O PAND2X1_852/a_56_28# PAND2X1_852/CTRL2 PAND2X1_852/CTRL
+ PAND2X1_852/a_76_28# PAND2X1
XPOR2X1_130 VDD GND PAND2X1_6/Y POR2X1_130/A POR2X1_130/Y POR2X1_141/m4_208_n4# POR2X1_130/O
+ POR2X1_130/CTRL2 POR2X1_130/a_16_28# POR2X1_130/CTRL POR2X1_130/a_76_344# POR2X1_130/a_56_344#
+ POR2X1
XPOR2X1_141 VDD GND POR2X1_139/Y POR2X1_141/A POR2X1_141/Y POR2X1_141/m4_208_n4# POR2X1_141/O
+ POR2X1_141/CTRL2 POR2X1_141/a_16_28# POR2X1_141/CTRL POR2X1_141/a_76_344# POR2X1_141/a_56_344#
+ POR2X1
XPOR2X1_152 VDD GND POR2X1_48/A POR2X1_152/A POR2X1_152/Y POR2X1_152/m4_208_n4# POR2X1_152/O
+ POR2X1_152/CTRL2 POR2X1_152/a_16_28# POR2X1_152/CTRL POR2X1_152/a_76_344# POR2X1_152/a_56_344#
+ POR2X1
XPOR2X1_174 VDD GND POR2X1_174/B POR2X1_174/A POR2X1_175/A POR2X1_174/m4_208_n4# POR2X1_174/O
+ POR2X1_174/CTRL2 POR2X1_174/a_16_28# POR2X1_174/CTRL POR2X1_174/a_76_344# POR2X1_174/a_56_344#
+ POR2X1
XPOR2X1_163 VDD GND POR2X1_52/A POR2X1_163/A POR2X1_163/Y POR2X1_163/m4_208_n4# POR2X1_163/O
+ POR2X1_163/CTRL2 POR2X1_163/a_16_28# POR2X1_163/CTRL POR2X1_163/a_76_344# POR2X1_163/a_56_344#
+ POR2X1
XPOR2X1_185 VDD GND PAND2X1_55/Y PAND2X1_73/Y POR2X1_188/A POR2X1_185/m4_208_n4# POR2X1_185/O
+ POR2X1_185/CTRL2 POR2X1_185/a_16_28# POR2X1_185/CTRL POR2X1_185/a_76_344# POR2X1_185/a_56_344#
+ POR2X1
XPOR2X1_196 VDD GND POR2X1_702/B PAND2X1_48/Y POR2X1_196/Y POR2X1_196/m4_208_n4# POR2X1_196/O
+ POR2X1_196/CTRL2 POR2X1_196/a_16_28# POR2X1_196/CTRL POR2X1_196/a_76_344# POR2X1_196/a_56_344#
+ POR2X1
XPAND2X1_115 VDD GND PAND2X1_115/B POR2X1_106/Y PAND2X1_115/Y PAND2X1_115/a_16_344#
+ PAND2X1_115/m4_208_n4# PAND2X1_115/O PAND2X1_115/a_56_28# PAND2X1_115/CTRL2 PAND2X1_115/CTRL
+ PAND2X1_115/a_76_28# PAND2X1
XPAND2X1_126 VDD GND PAND2X1_90/A PAND2X1_6/A POR2X1_532/A PAND2X1_126/a_16_344# PAND2X1_126/m4_208_n4#
+ PAND2X1_126/O PAND2X1_126/a_56_28# PAND2X1_126/CTRL2 PAND2X1_126/CTRL PAND2X1_126/a_76_28#
+ PAND2X1
XPAND2X1_104 VDD GND PAND2X1_8/Y PAND2X1_6/A POR2X1_814/B PAND2X1_104/a_16_344# PAND2X1_104/m4_208_n4#
+ PAND2X1_104/O PAND2X1_104/a_56_28# PAND2X1_104/CTRL2 PAND2X1_104/CTRL PAND2X1_104/a_76_28#
+ PAND2X1
XPAND2X1_137 VDD GND POR2X1_134/Y POR2X1_132/Y PAND2X1_137/Y PAND2X1_137/a_16_344#
+ PAND2X1_137/m4_208_n4# PAND2X1_137/O PAND2X1_137/a_56_28# PAND2X1_137/CTRL2 PAND2X1_137/CTRL
+ PAND2X1_137/a_76_28# PAND2X1
XPAND2X1_148 VDD GND POR2X1_146/Y POR2X1_145/Y PAND2X1_148/Y PAND2X1_148/a_16_344#
+ PAND2X1_148/m4_208_n4# PAND2X1_148/O PAND2X1_148/a_56_28# PAND2X1_148/CTRL2 PAND2X1_148/CTRL
+ PAND2X1_148/a_76_28# PAND2X1
XPAND2X1_159 VDD GND PAND2X1_9/Y POR2X1_68/B POR2X1_750/B PAND2X1_159/a_16_344# PAND2X1_159/m4_208_n4#
+ PAND2X1_159/O PAND2X1_159/a_56_28# PAND2X1_159/CTRL2 PAND2X1_159/CTRL PAND2X1_159/a_76_28#
+ PAND2X1
XPOR2X1_70 VDD GND POR2X1_3/A POR2X1_51/A POR2X1_72/B POR2X1_70/m4_208_n4# POR2X1_70/O
+ POR2X1_70/CTRL2 POR2X1_70/a_16_28# POR2X1_70/CTRL POR2X1_70/a_76_344# POR2X1_70/a_56_344#
+ POR2X1
XPOR2X1_92 VDD GND D_INPUT_1 POR2X1_8/Y POR2X1_93/A POR2X1_92/m4_208_n4# POR2X1_92/O
+ POR2X1_92/CTRL2 POR2X1_92/a_16_28# POR2X1_92/CTRL POR2X1_92/a_76_344# POR2X1_92/a_56_344#
+ POR2X1
XPOR2X1_81 VDD GND POR2X1_60/A POR2X1_81/A POR2X1_81/Y POR2X1_81/m4_208_n4# POR2X1_81/O
+ POR2X1_81/CTRL2 POR2X1_81/a_16_28# POR2X1_81/CTRL POR2X1_81/a_76_344# POR2X1_81/a_56_344#
+ POR2X1
XPAND2X1_682 VDD GND POR2X1_750/B PAND2X1_69/A POR2X1_685/A PAND2X1_682/a_16_344#
+ PAND2X1_682/m4_208_n4# PAND2X1_682/O PAND2X1_682/a_56_28# PAND2X1_682/CTRL2 PAND2X1_682/CTRL
+ PAND2X1_682/a_76_28# PAND2X1
XPAND2X1_671 VDD GND PAND2X1_6/A INPUT_2 PAND2X1_671/Y PAND2X1_671/a_16_344# PAND2X1_671/m4_208_n4#
+ PAND2X1_671/O PAND2X1_671/a_56_28# PAND2X1_671/CTRL2 PAND2X1_671/CTRL PAND2X1_671/a_76_28#
+ PAND2X1
XPAND2X1_660 VDD GND PAND2X1_660/B PAND2X1_655/Y PAND2X1_660/Y PAND2X1_660/a_16_344#
+ PAND2X1_660/m4_208_n4# PAND2X1_660/O PAND2X1_660/a_56_28# PAND2X1_660/CTRL2 PAND2X1_660/CTRL
+ PAND2X1_660/a_76_28# PAND2X1
XPAND2X1_693 VDD GND PAND2X1_69/A PAND2X1_94/A POR2X1_706/A PAND2X1_693/a_16_344#
+ PAND2X1_693/m4_208_n4# PAND2X1_693/O PAND2X1_693/a_56_28# PAND2X1_693/CTRL2 PAND2X1_693/CTRL
+ PAND2X1_693/a_76_28# PAND2X1
XPAND2X1_3 VDD GND PAND2X1_3/B PAND2X1_3/A POR2X1_66/B PAND2X1_3/a_16_344# PAND2X1_3/m4_208_n4#
+ PAND2X1_3/O PAND2X1_3/a_56_28# PAND2X1_3/CTRL2 PAND2X1_3/CTRL PAND2X1_3/a_76_28#
+ PAND2X1
XPAND2X1_490 VDD GND PAND2X1_85/Y POR2X1_4/Y POR2X1_557/A PAND2X1_490/a_16_344# PAND2X1_63/m4_208_n4#
+ PAND2X1_490/O PAND2X1_490/a_56_28# PAND2X1_490/CTRL2 PAND2X1_490/CTRL PAND2X1_490/a_76_28#
+ PAND2X1
XPOR2X1_707 VDD GND POR2X1_707/B POR2X1_707/A POR2X1_707/Y POR2X1_707/m4_208_n4# POR2X1_707/O
+ POR2X1_707/CTRL2 POR2X1_707/a_16_28# POR2X1_707/CTRL POR2X1_707/a_76_344# POR2X1_707/a_56_344#
+ POR2X1
XPOR2X1_718 VDD GND POR2X1_593/B POR2X1_718/A POR2X1_722/B POR2X1_718/m4_208_n4# POR2X1_718/O
+ POR2X1_718/CTRL2 POR2X1_718/a_16_28# POR2X1_718/CTRL POR2X1_718/a_76_344# POR2X1_718/a_56_344#
+ POR2X1
XPOR2X1_729 VDD GND POR2X1_687/Y POR2X1_855/B POR2X1_729/Y POR2X1_729/m4_208_n4# POR2X1_729/O
+ POR2X1_729/CTRL2 POR2X1_729/a_16_28# POR2X1_729/CTRL POR2X1_729/a_76_344# POR2X1_729/a_56_344#
+ POR2X1
XPOR2X1_515 VDD GND POR2X1_446/B POR2X1_514/Y POR2X1_515/Y POR2X1_515/m4_208_n4# POR2X1_515/O
+ POR2X1_515/CTRL2 POR2X1_515/a_16_28# POR2X1_515/CTRL POR2X1_515/a_76_344# POR2X1_515/a_56_344#
+ POR2X1
XPOR2X1_526 VDD GND POR2X1_32/A POR2X1_669/B POR2X1_526/Y POR2X1_526/m4_208_n4# POR2X1_526/O
+ POR2X1_526/CTRL2 POR2X1_526/a_16_28# POR2X1_526/CTRL POR2X1_526/a_76_344# POR2X1_526/a_56_344#
+ POR2X1
XPOR2X1_504 VDD GND POR2X1_41/B POR2X1_416/B POR2X1_504/Y POR2X1_504/m4_208_n4# POR2X1_504/O
+ POR2X1_504/CTRL2 POR2X1_504/a_16_28# POR2X1_504/CTRL POR2X1_504/a_76_344# POR2X1_504/a_56_344#
+ POR2X1
XPOR2X1_548 VDD GND POR2X1_548/B POR2X1_548/A POR2X1_549/A POR2X1_548/m4_208_n4# POR2X1_548/O
+ POR2X1_548/CTRL2 POR2X1_548/a_16_28# POR2X1_548/CTRL POR2X1_548/a_76_344# POR2X1_548/a_56_344#
+ POR2X1
XPOR2X1_559 VDD GND POR2X1_559/B POR2X1_559/A POR2X1_559/Y POR2X1_559/m4_208_n4# POR2X1_559/O
+ POR2X1_559/CTRL2 POR2X1_559/a_16_28# POR2X1_559/CTRL POR2X1_559/a_76_344# POR2X1_559/a_56_344#
+ POR2X1
XPOR2X1_537 VDD GND POR2X1_537/B POR2X1_537/A POR2X1_537/Y POR2X1_537/m4_208_n4# POR2X1_537/O
+ POR2X1_537/CTRL2 POR2X1_537/a_16_28# POR2X1_537/CTRL POR2X1_537/a_76_344# POR2X1_537/a_56_344#
+ POR2X1
XPOR2X1_301 VDD GND POR2X1_76/A POR2X1_301/A POR2X1_303/B POR2X1_301/m4_208_n4# POR2X1_301/O
+ POR2X1_301/CTRL2 POR2X1_301/a_16_28# POR2X1_301/CTRL POR2X1_301/a_76_344# POR2X1_301/a_56_344#
+ POR2X1
XPOR2X1_334 VDD GND POR2X1_334/B POR2X1_334/A POR2X1_334/Y POR2X1_334/m4_208_n4# POR2X1_334/O
+ POR2X1_334/CTRL2 POR2X1_334/a_16_28# POR2X1_334/CTRL POR2X1_334/a_76_344# POR2X1_334/a_56_344#
+ POR2X1
XPOR2X1_323 VDD GND POR2X1_96/A POR2X1_110/Y POR2X1_323/Y POR2X1_164/m4_208_n4# POR2X1_323/O
+ POR2X1_323/CTRL2 POR2X1_323/a_16_28# POR2X1_323/CTRL POR2X1_323/a_76_344# POR2X1_323/a_56_344#
+ POR2X1
XPOR2X1_312 VDD GND POR2X1_55/Y POR2X1_65/A POR2X1_312/Y POR2X1_312/m4_208_n4# POR2X1_312/O
+ POR2X1_312/CTRL2 POR2X1_312/a_16_28# POR2X1_312/CTRL POR2X1_312/a_76_344# POR2X1_312/a_56_344#
+ POR2X1
XPOR2X1_345 VDD GND POR2X1_555/B POR2X1_345/A POR2X1_348/A POR2X1_345/m4_208_n4# POR2X1_345/O
+ POR2X1_345/CTRL2 POR2X1_345/a_16_28# POR2X1_345/CTRL POR2X1_345/a_76_344# POR2X1_345/a_56_344#
+ POR2X1
XPOR2X1_367 VDD GND POR2X1_365/Y POR2X1_366/Y D_GATE_366 POR2X1_367/m4_208_n4# POR2X1_367/O
+ POR2X1_367/CTRL2 POR2X1_367/a_16_28# POR2X1_367/CTRL POR2X1_367/a_76_344# POR2X1_367/a_56_344#
+ POR2X1
XPOR2X1_356 VDD GND POR2X1_356/B POR2X1_356/A POR2X1_356/Y POR2X1_356/m4_208_n4# POR2X1_356/O
+ POR2X1_356/CTRL2 POR2X1_356/a_16_28# POR2X1_356/CTRL POR2X1_356/a_76_344# POR2X1_356/a_56_344#
+ POR2X1
XPOR2X1_378 VDD GND POR2X1_296/B POR2X1_378/A POR2X1_378/Y POR2X1_378/m4_208_n4# POR2X1_378/O
+ POR2X1_378/CTRL2 POR2X1_378/a_16_28# POR2X1_378/CTRL POR2X1_378/a_76_344# POR2X1_378/a_56_344#
+ POR2X1
XPOR2X1_389 VDD GND POR2X1_537/B POR2X1_389/A POR2X1_389/Y POR2X1_389/m4_208_n4# POR2X1_389/O
+ POR2X1_389/CTRL2 POR2X1_389/a_16_28# POR2X1_389/CTRL POR2X1_389/a_76_344# POR2X1_389/a_56_344#
+ POR2X1
XPAND2X1_308 VDD GND PAND2X1_308/B POR2X1_306/Y PAND2X1_308/Y PAND2X1_308/a_16_344#
+ PAND2X1_308/m4_208_n4# PAND2X1_308/O PAND2X1_308/a_56_28# PAND2X1_308/CTRL2 PAND2X1_308/CTRL
+ PAND2X1_308/a_76_28# PAND2X1
XPAND2X1_319 VDD GND PAND2X1_319/B PAND2X1_317/Y PAND2X1_354/A PAND2X1_319/a_16_344#
+ PAND2X1_319/m4_208_n4# PAND2X1_319/O PAND2X1_319/a_56_28# PAND2X1_319/CTRL2 PAND2X1_319/CTRL
+ PAND2X1_319/a_76_28# PAND2X1
XPAND2X1_820 VDD GND PAND2X1_820/B POR2X1_818/Y POR2X1_847/A PAND2X1_820/a_16_344#
+ PAND2X1_820/m4_208_n4# PAND2X1_820/O PAND2X1_820/a_56_28# PAND2X1_820/CTRL2 PAND2X1_820/CTRL
+ PAND2X1_820/a_76_28# PAND2X1
XPAND2X1_831 VDD GND POR2X1_300/Y POR2X1_273/Y PAND2X1_831/Y PAND2X1_831/a_16_344#
+ PAND2X1_831/m4_208_n4# PAND2X1_831/O PAND2X1_831/a_56_28# PAND2X1_831/CTRL2 PAND2X1_831/CTRL
+ PAND2X1_831/a_76_28# PAND2X1
XPAND2X1_853 VDD GND PAND2X1_853/B PAND2X1_35/Y PAND2X1_857/B PAND2X1_853/a_16_344#
+ PAND2X1_853/m4_208_n4# PAND2X1_853/O PAND2X1_853/a_56_28# PAND2X1_853/CTRL2 PAND2X1_853/CTRL
+ PAND2X1_853/a_76_28# PAND2X1
XPAND2X1_864 VDD GND PAND2X1_864/B PAND2X1_810/A PAND2X1_866/A PAND2X1_864/a_16_344#
+ PAND2X1_864/m4_208_n4# PAND2X1_864/O PAND2X1_864/a_56_28# PAND2X1_864/CTRL2 PAND2X1_864/CTRL
+ PAND2X1_864/a_76_28# PAND2X1
XPAND2X1_842 VDD GND PAND2X1_830/Y POR2X1_184/Y PAND2X1_842/Y PAND2X1_842/a_16_344#
+ PAND2X1_842/m4_208_n4# PAND2X1_842/O PAND2X1_842/a_56_28# PAND2X1_842/CTRL2 PAND2X1_842/CTRL
+ PAND2X1_842/a_76_28# PAND2X1
XPOR2X1_142 VDD GND POR2X1_49/Y POR2X1_65/A POR2X1_142/Y POR2X1_142/m4_208_n4# POR2X1_142/O
+ POR2X1_142/CTRL2 POR2X1_142/a_16_28# POR2X1_142/CTRL POR2X1_142/a_76_344# POR2X1_142/a_56_344#
+ POR2X1
XPOR2X1_120 VDD GND POR2X1_294/B PAND2X1_39/B POR2X1_121/A POR2X1_120/m4_208_n4# POR2X1_120/O
+ POR2X1_120/CTRL2 POR2X1_120/a_16_28# POR2X1_120/CTRL POR2X1_120/a_76_344# POR2X1_120/a_56_344#
+ POR2X1
XPOR2X1_131 VDD GND POR2X1_13/A POR2X1_131/A POR2X1_131/Y POR2X1_131/m4_208_n4# POR2X1_131/O
+ POR2X1_131/CTRL2 POR2X1_131/a_16_28# POR2X1_131/CTRL POR2X1_131/a_76_344# POR2X1_131/a_56_344#
+ POR2X1
XPOR2X1_153 VDD GND INPUT_1 POR2X1_37/Y POR2X1_153/Y POR2X1_153/m4_208_n4# POR2X1_153/O
+ POR2X1_153/CTRL2 POR2X1_153/a_16_28# POR2X1_153/CTRL POR2X1_153/a_76_344# POR2X1_153/a_56_344#
+ POR2X1
XPOR2X1_175 VDD GND POR2X1_175/B POR2X1_175/A POR2X1_853/A POR2X1_175/m4_208_n4# POR2X1_175/O
+ POR2X1_175/CTRL2 POR2X1_175/a_16_28# POR2X1_175/CTRL POR2X1_175/a_76_344# POR2X1_175/a_56_344#
+ POR2X1
XPOR2X1_164 VDD GND POR2X1_20/B POR2X1_376/B POR2X1_164/Y POR2X1_164/m4_208_n4# POR2X1_164/O
+ POR2X1_164/CTRL2 POR2X1_164/a_16_28# POR2X1_164/CTRL POR2X1_164/a_76_344# POR2X1_164/a_56_344#
+ POR2X1
XPOR2X1_186 VDD GND POR2X1_186/B POR2X1_188/A POR2X1_186/Y POR2X1_186/m4_208_n4# POR2X1_186/O
+ POR2X1_186/CTRL2 POR2X1_186/a_16_28# POR2X1_186/CTRL POR2X1_186/a_76_344# POR2X1_186/a_56_344#
+ POR2X1
XPOR2X1_197 VDD GND PAND2X1_52/Y PAND2X1_56/Y POR2X1_197/Y POR2X1_197/m4_208_n4# POR2X1_197/O
+ POR2X1_197/CTRL2 POR2X1_197/a_16_28# POR2X1_197/CTRL POR2X1_197/a_76_344# POR2X1_197/a_56_344#
+ POR2X1
XPAND2X1_127 VDD GND POR2X1_532/A POR2X1_66/B POR2X1_128/A PAND2X1_127/a_16_344# PAND2X1_127/m4_208_n4#
+ PAND2X1_127/O PAND2X1_127/a_56_28# PAND2X1_127/CTRL2 PAND2X1_127/CTRL PAND2X1_127/a_76_28#
+ PAND2X1
XPAND2X1_116 VDD GND PAND2X1_115/Y PAND2X1_114/Y PAND2X1_216/B PAND2X1_116/a_16_344#
+ PAND2X1_116/m4_208_n4# PAND2X1_116/O PAND2X1_116/a_56_28# PAND2X1_116/CTRL2 PAND2X1_116/CTRL
+ PAND2X1_116/a_76_28# PAND2X1
XPAND2X1_105 VDD GND POR2X1_411/B POR2X1_77/Y POR2X1_251/A PAND2X1_105/a_16_344# PAND2X1_105/m4_208_n4#
+ PAND2X1_105/O PAND2X1_105/a_56_28# PAND2X1_105/CTRL2 PAND2X1_105/CTRL PAND2X1_105/a_76_28#
+ PAND2X1
XPAND2X1_138 VDD GND POR2X1_136/Y POR2X1_135/Y PAND2X1_139/B PAND2X1_138/a_16_344#
+ PAND2X1_138/m4_208_n4# PAND2X1_138/O PAND2X1_138/a_56_28# PAND2X1_138/CTRL2 PAND2X1_138/CTRL
+ PAND2X1_138/a_76_28# PAND2X1
XPAND2X1_149 VDD GND PAND2X1_148/Y PAND2X1_149/A PAND2X1_209/A PAND2X1_149/a_16_344#
+ PAND2X1_149/m4_208_n4# PAND2X1_149/O PAND2X1_149/a_56_28# PAND2X1_149/CTRL2 PAND2X1_149/CTRL
+ PAND2X1_149/a_76_28# PAND2X1
XPOR2X1_60 VDD GND POR2X1_38/Y POR2X1_60/A POR2X1_60/Y POR2X1_60/m4_208_n4# POR2X1_60/O
+ POR2X1_60/CTRL2 POR2X1_60/a_16_28# POR2X1_60/CTRL POR2X1_60/a_76_344# POR2X1_60/a_56_344#
+ POR2X1
XPOR2X1_71 VDD GND POR2X1_5/Y POR2X1_62/Y POR2X1_71/Y POR2X1_71/m4_208_n4# POR2X1_71/O
+ POR2X1_71/CTRL2 POR2X1_71/a_16_28# POR2X1_71/CTRL POR2X1_71/a_76_344# POR2X1_71/a_56_344#
+ POR2X1
XPOR2X1_82 VDD GND POR2X1_14/Y POR2X1_29/A POR2X1_83/A POR2X1_82/m4_208_n4# POR2X1_82/O
+ POR2X1_82/CTRL2 POR2X1_82/a_16_28# POR2X1_82/CTRL POR2X1_82/a_76_344# POR2X1_82/a_56_344#
+ POR2X1
XPOR2X1_93 VDD GND POR2X1_83/B POR2X1_93/A POR2X1_93/Y POR2X1_93/m4_208_n4# POR2X1_93/O
+ POR2X1_93/CTRL2 POR2X1_93/a_16_28# POR2X1_93/CTRL POR2X1_93/a_76_344# POR2X1_93/a_56_344#
+ POR2X1
XPAND2X1_683 VDD GND PAND2X1_58/A POR2X1_78/B POR2X1_686/B PAND2X1_683/a_16_344# PAND2X1_683/m4_208_n4#
+ PAND2X1_683/O PAND2X1_683/a_56_28# PAND2X1_683/CTRL2 PAND2X1_683/CTRL PAND2X1_683/a_76_28#
+ PAND2X1
XPAND2X1_661 VDD GND PAND2X1_661/B PAND2X1_653/Y PAND2X1_661/Y PAND2X1_661/a_16_344#
+ PAND2X1_661/m4_208_n4# PAND2X1_661/O PAND2X1_661/a_56_28# PAND2X1_661/CTRL2 PAND2X1_661/CTRL
+ PAND2X1_661/a_76_28# PAND2X1
XPAND2X1_650 VDD GND PAND2X1_641/Y PAND2X1_650/A PAND2X1_654/A PAND2X1_650/a_16_344#
+ PAND2X1_650/m4_208_n4# PAND2X1_650/O PAND2X1_650/a_56_28# PAND2X1_650/CTRL2 PAND2X1_650/CTRL
+ PAND2X1_650/a_76_28# PAND2X1
XPAND2X1_672 VDD GND PAND2X1_671/Y POR2X1_260/A POR2X1_673/A PAND2X1_672/a_16_344#
+ PAND2X1_672/m4_208_n4# PAND2X1_672/O PAND2X1_672/a_56_28# PAND2X1_672/CTRL2 PAND2X1_672/CTRL
+ PAND2X1_672/a_76_28# PAND2X1
XPAND2X1_694 VDD GND PAND2X1_425/Y POR2X1_614/A POR2X1_707/B PAND2X1_694/a_16_344#
+ PAND2X1_694/m4_208_n4# PAND2X1_694/O PAND2X1_694/a_56_28# PAND2X1_694/CTRL2 PAND2X1_694/CTRL
+ PAND2X1_694/a_76_28# PAND2X1
XPAND2X1_4 VDD GND D_INPUT_1 INPUT_0 PAND2X1_6/A PAND2X1_4/a_16_344# PAND2X1_4/m4_208_n4#
+ PAND2X1_4/O PAND2X1_4/a_56_28# PAND2X1_4/CTRL2 PAND2X1_4/CTRL PAND2X1_4/a_76_28#
+ PAND2X1
XPAND2X1_491 VDD GND POR2X1_590/A PAND2X1_32/B POR2X1_493/B PAND2X1_491/a_16_344#
+ PAND2X1_491/m4_208_n4# PAND2X1_491/O PAND2X1_491/a_56_28# PAND2X1_491/CTRL2 PAND2X1_491/CTRL
+ PAND2X1_491/a_76_28# PAND2X1
XPAND2X1_480 VDD GND PAND2X1_480/B PAND2X1_478/Y GATE_479 PAND2X1_480/a_16_344# PAND2X1_776/m4_208_n4#
+ PAND2X1_480/O PAND2X1_480/a_56_28# PAND2X1_480/CTRL2 PAND2X1_480/CTRL PAND2X1_480/a_76_28#
+ PAND2X1
XPOR2X1_708 VDD GND POR2X1_708/B POR2X1_779/A POR2X1_712/A POR2X1_708/m4_208_n4# POR2X1_708/O
+ POR2X1_708/CTRL2 POR2X1_708/a_16_28# POR2X1_708/CTRL POR2X1_708/a_76_344# POR2X1_708/a_56_344#
+ POR2X1
XPOR2X1_719 VDD GND POR2X1_719/B POR2X1_719/A POR2X1_722/A POR2X1_719/m4_208_n4# POR2X1_719/O
+ POR2X1_719/CTRL2 POR2X1_719/a_16_28# POR2X1_719/CTRL POR2X1_719/a_76_344# POR2X1_719/a_56_344#
+ POR2X1
XPOR2X1_516 VDD GND POR2X1_516/B POR2X1_516/A POR2X1_516/Y POR2X1_516/m4_208_n4# POR2X1_516/O
+ POR2X1_516/CTRL2 POR2X1_516/a_16_28# POR2X1_516/CTRL POR2X1_516/a_76_344# POR2X1_516/a_56_344#
+ POR2X1
XPOR2X1_505 VDD GND POR2X1_20/B POR2X1_23/Y POR2X1_505/Y POR2X1_505/m4_208_n4# POR2X1_505/O
+ POR2X1_505/CTRL2 POR2X1_505/a_16_28# POR2X1_505/CTRL POR2X1_505/a_76_344# POR2X1_505/a_56_344#
+ POR2X1
XPOR2X1_549 VDD GND POR2X1_549/B POR2X1_549/A POR2X1_565/B POR2X1_549/m4_208_n4# POR2X1_549/O
+ POR2X1_549/CTRL2 POR2X1_549/a_16_28# POR2X1_549/CTRL POR2X1_549/a_76_344# POR2X1_549/a_56_344#
+ POR2X1
XPOR2X1_538 VDD GND POR2X1_193/A POR2X1_538/A POR2X1_539/A POR2X1_538/m4_208_n4# POR2X1_538/O
+ POR2X1_538/CTRL2 POR2X1_538/a_16_28# POR2X1_538/CTRL POR2X1_538/a_76_344# POR2X1_538/a_56_344#
+ POR2X1
XPOR2X1_527 VDD GND POR2X1_65/A POR2X1_110/Y POR2X1_527/Y POR2X1_527/m4_208_n4# POR2X1_527/O
+ POR2X1_527/CTRL2 POR2X1_527/a_16_28# POR2X1_527/CTRL POR2X1_527/a_76_344# POR2X1_527/a_56_344#
+ POR2X1
XPOR2X1_335 VDD GND POR2X1_335/B POR2X1_335/A POR2X1_335/Y POR2X1_335/m4_208_n4# POR2X1_335/O
+ POR2X1_335/CTRL2 POR2X1_335/a_16_28# POR2X1_335/CTRL POR2X1_335/a_76_344# POR2X1_335/a_56_344#
+ POR2X1
XPOR2X1_313 VDD GND POR2X1_72/B POR2X1_90/Y POR2X1_313/Y POR2X1_313/m4_208_n4# POR2X1_313/O
+ POR2X1_313/CTRL2 POR2X1_313/a_16_28# POR2X1_313/CTRL POR2X1_313/a_76_344# POR2X1_313/a_56_344#
+ POR2X1
XPOR2X1_324 VDD GND POR2X1_324/B POR2X1_324/A POR2X1_324/Y POR2X1_324/m4_208_n4# POR2X1_324/O
+ POR2X1_324/CTRL2 POR2X1_324/a_16_28# POR2X1_324/CTRL POR2X1_324/a_76_344# POR2X1_324/a_56_344#
+ POR2X1
XPOR2X1_302 VDD GND POR2X1_302/B POR2X1_302/A POR2X1_302/Y POR2X1_302/m4_208_n4# POR2X1_302/O
+ POR2X1_302/CTRL2 POR2X1_302/a_16_28# POR2X1_302/CTRL POR2X1_302/a_76_344# POR2X1_302/a_56_344#
+ POR2X1
XPOR2X1_346 VDD GND POR2X1_346/B POR2X1_346/A POR2X1_347/A POR2X1_346/m4_208_n4# POR2X1_346/O
+ POR2X1_346/CTRL2 POR2X1_346/a_16_28# POR2X1_346/CTRL POR2X1_346/a_76_344# POR2X1_346/a_56_344#
+ POR2X1
XPOR2X1_357 VDD GND POR2X1_357/B POR2X1_353/Y POR2X1_357/Y POR2X1_357/m4_208_n4# POR2X1_357/O
+ POR2X1_357/CTRL2 POR2X1_357/a_16_28# POR2X1_357/CTRL POR2X1_357/a_76_344# POR2X1_357/a_56_344#
+ POR2X1
XPOR2X1_368 VDD GND POR2X1_7/A POR2X1_271/A POR2X1_368/Y POR2X1_368/m4_208_n4# POR2X1_368/O
+ POR2X1_368/CTRL2 POR2X1_368/a_16_28# POR2X1_368/CTRL POR2X1_368/a_76_344# POR2X1_368/a_56_344#
+ POR2X1
XPOR2X1_379 VDD GND POR2X1_260/B POR2X1_66/A POR2X1_379/Y POR2X1_379/m4_208_n4# POR2X1_379/O
+ POR2X1_379/CTRL2 POR2X1_379/a_16_28# POR2X1_379/CTRL POR2X1_379/a_76_344# POR2X1_379/a_56_344#
+ POR2X1
XPAND2X1_309 VDD GND POR2X1_814/A PAND2X1_58/A POR2X1_335/B PAND2X1_309/a_16_344#
+ PAND2X1_309/m4_208_n4# PAND2X1_309/O PAND2X1_309/a_56_28# PAND2X1_309/CTRL2 PAND2X1_309/CTRL
+ PAND2X1_309/a_76_28# PAND2X1
XPAND2X1_810 VDD GND PAND2X1_810/B PAND2X1_810/A PAND2X1_812/A PAND2X1_810/a_16_344#
+ PAND2X1_810/m4_208_n4# PAND2X1_810/O PAND2X1_810/a_56_28# PAND2X1_810/CTRL2 PAND2X1_810/CTRL
+ PAND2X1_810/a_76_28# PAND2X1
XPAND2X1_832 VDD GND POR2X1_433/Y POR2X1_423/Y PAND2X1_841/B PAND2X1_832/a_16_344#
+ PAND2X1_832/m4_208_n4# PAND2X1_832/O PAND2X1_832/a_56_28# PAND2X1_832/CTRL2 PAND2X1_832/CTRL
+ PAND2X1_832/a_76_28# PAND2X1
XPAND2X1_821 VDD GND PAND2X1_72/A POR2X1_294/B POR2X1_835/B PAND2X1_821/a_16_344#
+ PAND2X1_821/m4_208_n4# PAND2X1_821/O PAND2X1_821/a_56_28# PAND2X1_821/CTRL2 PAND2X1_821/CTRL
+ PAND2X1_821/a_76_28# PAND2X1
XPAND2X1_865 VDD GND PAND2X1_862/Y PAND2X1_865/A PAND2X1_865/Y PAND2X1_865/a_16_344#
+ PAND2X1_865/m4_208_n4# PAND2X1_865/O PAND2X1_865/a_56_28# PAND2X1_865/CTRL2 PAND2X1_865/CTRL
+ PAND2X1_865/a_76_28# PAND2X1
XPAND2X1_843 VDD GND POR2X1_278/Y POR2X1_251/Y PAND2X1_843/Y PAND2X1_843/a_16_344#
+ PAND2X1_843/m4_208_n4# PAND2X1_843/O PAND2X1_843/a_56_28# PAND2X1_843/CTRL2 PAND2X1_843/CTRL
+ PAND2X1_843/a_76_28# PAND2X1
XPAND2X1_854 VDD GND PAND2X1_535/Y PAND2X1_854/A PAND2X1_854/Y PAND2X1_854/a_16_344#
+ PAND2X1_854/m4_208_n4# PAND2X1_854/O PAND2X1_854/a_56_28# PAND2X1_854/CTRL2 PAND2X1_854/CTRL
+ PAND2X1_854/a_76_28# PAND2X1
XPOR2X1_110 VDD GND INPUT_0 POR2X1_14/Y POR2X1_110/Y POR2X1_110/m4_208_n4# POR2X1_110/O
+ POR2X1_110/CTRL2 POR2X1_110/a_16_28# POR2X1_110/CTRL POR2X1_110/a_76_344# POR2X1_110/a_56_344#
+ POR2X1
XPOR2X1_143 VDD GND INPUT_1 POR2X1_8/Y POR2X1_376/B POR2X1_143/m4_208_n4# POR2X1_143/O
+ POR2X1_143/CTRL2 POR2X1_143/a_16_28# POR2X1_143/CTRL POR2X1_143/a_76_344# POR2X1_143/a_56_344#
+ POR2X1
XPOR2X1_121 VDD GND POR2X1_121/B POR2X1_121/A POR2X1_121/Y POR2X1_121/m4_208_n4# POR2X1_121/O
+ POR2X1_121/CTRL2 POR2X1_121/a_16_28# POR2X1_121/CTRL POR2X1_121/a_76_344# POR2X1_121/a_56_344#
+ POR2X1
XPOR2X1_132 VDD GND POR2X1_90/Y POR2X1_96/A POR2X1_132/Y POR2X1_132/m4_208_n4# POR2X1_132/O
+ POR2X1_132/CTRL2 POR2X1_132/a_16_28# POR2X1_132/CTRL POR2X1_132/a_76_344# POR2X1_132/a_56_344#
+ POR2X1
XPOR2X1_154 VDD GND PAND2X1_6/Y PAND2X1_39/B POR2X1_156/B POR2X1_154/m4_208_n4# POR2X1_154/O
+ POR2X1_154/CTRL2 POR2X1_154/a_16_28# POR2X1_154/CTRL POR2X1_154/a_76_344# POR2X1_154/a_56_344#
+ POR2X1
XPOR2X1_165 VDD GND POR2X1_52/A POR2X1_73/Y POR2X1_165/Y POR2X1_165/m4_208_n4# POR2X1_165/O
+ POR2X1_165/CTRL2 POR2X1_165/a_16_28# POR2X1_165/CTRL POR2X1_165/a_76_344# POR2X1_165/a_56_344#
+ POR2X1
XPOR2X1_176 VDD GND POR2X1_83/B POR2X1_90/Y POR2X1_176/Y POR2X1_176/m4_208_n4# POR2X1_176/O
+ POR2X1_176/CTRL2 POR2X1_176/a_16_28# POR2X1_176/CTRL POR2X1_176/a_76_344# POR2X1_176/a_56_344#
+ POR2X1
XPOR2X1_198 VDD GND POR2X1_198/B POR2X1_197/Y POR2X1_208/A POR2X1_198/m4_208_n4# POR2X1_198/O
+ POR2X1_198/CTRL2 POR2X1_198/a_16_28# POR2X1_198/CTRL POR2X1_198/a_76_344# POR2X1_198/a_56_344#
+ POR2X1
XPOR2X1_187 VDD GND POR2X1_40/Y POR2X1_594/A POR2X1_187/Y POR2X1_187/m4_208_n4# POR2X1_187/O
+ POR2X1_187/CTRL2 POR2X1_187/a_16_28# POR2X1_187/CTRL POR2X1_187/a_76_344# POR2X1_187/a_56_344#
+ POR2X1
XPAND2X1_117 VDD GND PAND2X1_72/A PAND2X1_63/Y POR2X1_123/B PAND2X1_117/a_16_344#
+ PAND2X1_117/m4_208_n4# PAND2X1_117/O PAND2X1_117/a_56_28# PAND2X1_117/CTRL2 PAND2X1_117/CTRL
+ PAND2X1_117/a_76_28# PAND2X1
XPAND2X1_106 VDD GND POR2X1_105/Y PAND2X1_48/B POR2X1_554/B PAND2X1_106/a_16_344#
+ PAND2X1_106/m4_208_n4# PAND2X1_106/O PAND2X1_106/a_56_28# PAND2X1_106/CTRL2 PAND2X1_106/CTRL
+ PAND2X1_106/a_76_28# PAND2X1
XPAND2X1_139 VDD GND PAND2X1_139/B PAND2X1_137/Y PAND2X1_139/Y PAND2X1_139/a_16_344#
+ PAND2X1_139/m4_208_n4# PAND2X1_139/O PAND2X1_139/a_56_28# PAND2X1_139/CTRL2 PAND2X1_139/CTRL
+ PAND2X1_139/a_76_28# PAND2X1
XPAND2X1_128 VDD GND POR2X1_127/Y POR2X1_125/Y PAND2X1_140/A PAND2X1_128/a_16_344#
+ PAND2X1_128/m4_208_n4# PAND2X1_128/O PAND2X1_128/a_56_28# PAND2X1_128/CTRL2 PAND2X1_128/CTRL
+ PAND2X1_128/a_76_28# PAND2X1
XPOR2X1_61 VDD GND POR2X1_61/B POR2X1_61/A POR2X1_61/Y POR2X1_61/m4_208_n4# POR2X1_61/O
+ POR2X1_61/CTRL2 POR2X1_61/a_16_28# POR2X1_61/CTRL POR2X1_61/a_76_344# POR2X1_61/a_56_344#
+ POR2X1
XPOR2X1_50 VDD GND INPUT_6 INPUT_7 POR2X1_51/A POR2X1_50/m4_208_n4# POR2X1_50/O POR2X1_50/CTRL2
+ POR2X1_50/a_16_28# POR2X1_50/CTRL POR2X1_50/a_76_344# POR2X1_50/a_56_344# POR2X1
XPOR2X1_94 VDD GND POR2X1_14/Y POR2X1_94/A POR2X1_96/B POR2X1_94/m4_208_n4# POR2X1_94/O
+ POR2X1_94/CTRL2 POR2X1_94/a_16_28# POR2X1_94/CTRL POR2X1_94/a_76_344# POR2X1_94/a_56_344#
+ POR2X1
XPOR2X1_83 VDD GND POR2X1_83/B POR2X1_83/A POR2X1_83/Y POR2X1_83/m4_208_n4# POR2X1_83/O
+ POR2X1_83/CTRL2 POR2X1_83/a_16_28# POR2X1_83/CTRL POR2X1_83/a_76_344# POR2X1_83/a_56_344#
+ POR2X1
XPOR2X1_72 VDD GND POR2X1_72/B POR2X1_71/Y POR2X1_72/Y POR2X1_72/m4_208_n4# POR2X1_72/O
+ POR2X1_72/CTRL2 POR2X1_72/a_16_28# POR2X1_72/CTRL POR2X1_72/a_76_344# POR2X1_72/a_56_344#
+ POR2X1
XPAND2X1_640 VDD GND PAND2X1_640/B PAND2X1_633/Y PAND2X1_650/A PAND2X1_640/a_16_344#
+ PAND2X1_640/m4_208_n4# PAND2X1_640/O PAND2X1_640/a_56_28# PAND2X1_640/CTRL2 PAND2X1_640/CTRL
+ PAND2X1_640/a_76_28# PAND2X1
XPAND2X1_651 VDD GND PAND2X1_639/Y PAND2X1_651/A PAND2X1_651/Y PAND2X1_651/a_16_344#
+ PAND2X1_651/m4_208_n4# PAND2X1_651/O PAND2X1_651/a_56_28# PAND2X1_651/CTRL2 PAND2X1_651/CTRL
+ PAND2X1_651/a_76_28# PAND2X1
XPAND2X1_673 VDD GND POR2X1_672/Y POR2X1_670/Y PAND2X1_673/Y PAND2X1_673/a_16_344#
+ PAND2X1_673/m4_208_n4# PAND2X1_673/O PAND2X1_673/a_56_28# PAND2X1_673/CTRL2 PAND2X1_673/CTRL
+ PAND2X1_673/a_76_28# PAND2X1
XPAND2X1_662 VDD GND PAND2X1_661/Y PAND2X1_660/Y PAND2X1_662/Y PAND2X1_662/a_16_344#
+ PAND2X1_662/m4_208_n4# PAND2X1_662/O PAND2X1_662/a_56_28# PAND2X1_662/CTRL2 PAND2X1_662/CTRL
+ PAND2X1_662/a_76_28# PAND2X1
XPAND2X1_684 VDD GND POR2X1_296/B POR2X1_260/B POR2X1_686/A PAND2X1_684/a_16_344#
+ PAND2X1_684/m4_208_n4# PAND2X1_684/O PAND2X1_684/a_56_28# PAND2X1_684/CTRL2 PAND2X1_684/CTRL
+ PAND2X1_684/a_76_28# PAND2X1
XPAND2X1_695 VDD GND PAND2X1_48/B PAND2X1_23/Y POR2X1_707/A PAND2X1_695/a_16_344#
+ PAND2X1_695/m4_208_n4# PAND2X1_695/O PAND2X1_695/a_56_28# PAND2X1_695/CTRL2 PAND2X1_695/CTRL
+ PAND2X1_695/a_76_28# PAND2X1
XPAND2X1_5 VDD GND INPUT_3 D_INPUT_2 POR2X1_68/B PAND2X1_5/a_16_344# PAND2X1_5/m4_208_n4#
+ PAND2X1_5/O PAND2X1_5/a_56_28# PAND2X1_5/CTRL2 PAND2X1_5/CTRL PAND2X1_5/a_76_28#
+ PAND2X1
XPAND2X1_470 VDD GND PAND2X1_467/Y PAND2X1_470/A PAND2X1_477/A PAND2X1_470/a_16_344#
+ PAND2X1_470/m4_208_n4# PAND2X1_470/O PAND2X1_470/a_56_28# PAND2X1_470/CTRL2 PAND2X1_470/CTRL
+ PAND2X1_470/a_76_28# PAND2X1
XPAND2X1_481 VDD GND POR2X1_294/Y POR2X1_66/B POR2X1_555/A PAND2X1_481/a_16_344# PAND2X1_481/m4_208_n4#
+ PAND2X1_481/O PAND2X1_481/a_56_28# PAND2X1_481/CTRL2 PAND2X1_481/CTRL PAND2X1_481/a_76_28#
+ PAND2X1
XPAND2X1_492 VDD GND POR2X1_532/A PAND2X1_60/B POR2X1_493/A PAND2X1_492/a_16_344#
+ PAND2X1_492/m4_208_n4# PAND2X1_492/O PAND2X1_492/a_56_28# PAND2X1_492/CTRL2 PAND2X1_492/CTRL
+ PAND2X1_492/a_76_28# PAND2X1
XPOR2X1_709 VDD GND POR2X1_709/B POR2X1_709/A POR2X1_711/B POR2X1_709/m4_208_n4# POR2X1_709/O
+ POR2X1_709/CTRL2 POR2X1_709/a_16_28# POR2X1_709/CTRL POR2X1_709/a_76_344# POR2X1_709/a_56_344#
+ POR2X1
XPOR2X1_506 VDD GND POR2X1_506/B POR2X1_447/B POR2X1_508/B POR2X1_506/m4_208_n4# POR2X1_506/O
+ POR2X1_506/CTRL2 POR2X1_506/a_16_28# POR2X1_506/CTRL POR2X1_506/a_76_344# POR2X1_506/a_56_344#
+ POR2X1
XPOR2X1_517 VDD GND POR2X1_32/A POR2X1_667/A POR2X1_517/Y POR2X1_517/m4_208_n4# POR2X1_517/O
+ POR2X1_517/CTRL2 POR2X1_517/a_16_28# POR2X1_517/CTRL POR2X1_517/a_76_344# POR2X1_517/a_56_344#
+ POR2X1
XPOR2X1_528 VDD GND POR2X1_7/A POR2X1_57/A POR2X1_528/Y POR2X1_528/m4_208_n4# POR2X1_528/O
+ POR2X1_528/CTRL2 POR2X1_528/a_16_28# POR2X1_528/CTRL POR2X1_528/a_76_344# POR2X1_528/a_56_344#
+ POR2X1
XPOR2X1_539 VDD GND POR2X1_537/Y POR2X1_539/A POR2X1_567/A POR2X1_539/m4_208_n4# POR2X1_539/O
+ POR2X1_539/CTRL2 POR2X1_539/a_16_28# POR2X1_539/CTRL POR2X1_539/a_76_344# POR2X1_539/a_56_344#
+ POR2X1
XPOR2X1_303 VDD GND POR2X1_303/B POR2X1_302/Y POR2X1_566/A POR2X1_303/m4_208_n4# POR2X1_303/O
+ POR2X1_303/CTRL2 POR2X1_303/a_16_28# POR2X1_303/CTRL POR2X1_303/a_76_344# POR2X1_303/a_56_344#
+ POR2X1
XPOR2X1_314 VDD GND POR2X1_16/A POR2X1_65/A POR2X1_314/Y POR2X1_314/m4_208_n4# POR2X1_314/O
+ POR2X1_314/CTRL2 POR2X1_314/a_16_28# POR2X1_314/CTRL POR2X1_314/a_76_344# POR2X1_314/a_56_344#
+ POR2X1
XPOR2X1_325 VDD GND POR2X1_325/B POR2X1_325/A POR2X1_326/A POR2X1_325/m4_208_n4# POR2X1_325/O
+ POR2X1_325/CTRL2 POR2X1_325/a_16_28# POR2X1_325/CTRL POR2X1_325/a_76_344# POR2X1_325/a_56_344#
+ POR2X1
XPOR2X1_347 VDD GND POR2X1_347/B POR2X1_347/A POR2X1_360/A POR2X1_347/m4_208_n4# POR2X1_347/O
+ POR2X1_347/CTRL2 POR2X1_347/a_16_28# POR2X1_347/CTRL POR2X1_347/a_76_344# POR2X1_347/a_56_344#
+ POR2X1
XPOR2X1_358 VDD GND POR2X1_350/Y POR2X1_351/Y POR2X1_364/A POR2X1_333/m4_208_n4# POR2X1_358/O
+ POR2X1_358/CTRL2 POR2X1_358/a_16_28# POR2X1_358/CTRL POR2X1_358/a_76_344# POR2X1_358/a_56_344#
+ POR2X1
XPOR2X1_336 VDD GND POR2X1_538/A POR2X1_703/A POR2X1_337/A POR2X1_336/m4_208_n4# POR2X1_336/O
+ POR2X1_336/CTRL2 POR2X1_336/a_16_28# POR2X1_336/CTRL POR2X1_336/a_76_344# POR2X1_336/a_56_344#
+ POR2X1
XPOR2X1_369 VDD GND POR2X1_43/B POR2X1_119/Y POR2X1_369/Y POR2X1_369/m4_208_n4# POR2X1_369/O
+ POR2X1_369/CTRL2 POR2X1_369/a_16_28# POR2X1_369/CTRL POR2X1_369/a_76_344# POR2X1_369/a_56_344#
+ POR2X1
XPAND2X1_800 VDD GND POR2X1_760/Y PAND2X1_687/Y PAND2X1_801/B PAND2X1_800/a_16_344#
+ POR2X1_760/m4_208_n4# PAND2X1_800/O PAND2X1_800/a_56_28# PAND2X1_800/CTRL2 PAND2X1_800/CTRL
+ PAND2X1_800/a_76_28# PAND2X1
XPAND2X1_811 VDD GND PAND2X1_808/Y PAND2X1_811/A PAND2X1_811/Y PAND2X1_811/a_16_344#
+ PAND2X1_811/m4_208_n4# PAND2X1_811/O PAND2X1_811/a_56_28# PAND2X1_811/CTRL2 PAND2X1_811/CTRL
+ PAND2X1_811/a_76_28# PAND2X1
XPAND2X1_822 VDD GND POR2X1_590/A PAND2X1_65/B POR2X1_835/A PAND2X1_822/a_16_344#
+ PAND2X1_822/m4_208_n4# PAND2X1_822/O PAND2X1_822/a_56_28# PAND2X1_822/CTRL2 PAND2X1_822/CTRL
+ PAND2X1_822/a_76_28# PAND2X1
XPAND2X1_844 VDD GND PAND2X1_844/B POR2X1_497/Y PAND2X1_844/Y PAND2X1_844/a_16_344#
+ PAND2X1_351/m4_208_n4# PAND2X1_844/O PAND2X1_844/a_56_28# PAND2X1_844/CTRL2 PAND2X1_844/CTRL
+ PAND2X1_844/a_76_28# PAND2X1
XPAND2X1_833 VDD GND POR2X1_495/Y POR2X1_482/Y PAND2X1_840/A PAND2X1_833/a_16_344#
+ PAND2X1_833/m4_208_n4# PAND2X1_833/O PAND2X1_833/a_56_28# PAND2X1_833/CTRL2 PAND2X1_833/CTRL
+ PAND2X1_833/a_76_28# PAND2X1
XPAND2X1_855 VDD GND POR2X1_829/Y PAND2X1_691/Y PAND2X1_856/B PAND2X1_855/a_16_344#
+ PAND2X1_855/m4_208_n4# PAND2X1_855/O PAND2X1_855/a_56_28# PAND2X1_855/CTRL2 PAND2X1_855/CTRL
+ PAND2X1_855/a_76_28# PAND2X1
XPAND2X1_866 VDD GND PAND2X1_865/Y PAND2X1_866/A GATE_865 PAND2X1_866/a_16_344# PAND2X1_866/m4_208_n4#
+ PAND2X1_866/O PAND2X1_866/a_56_28# PAND2X1_866/CTRL2 PAND2X1_866/CTRL PAND2X1_866/a_76_28#
+ PAND2X1
XPOR2X1_100 VDD GND PAND2X1_86/Y PAND2X1_88/Y POR2X1_101/A POR2X1_100/m4_208_n4# POR2X1_100/O
+ POR2X1_100/CTRL2 POR2X1_100/a_16_28# POR2X1_100/CTRL POR2X1_100/a_76_344# POR2X1_100/a_56_344#
+ POR2X1
XPOR2X1_122 VDD GND POR2X1_57/A POR2X1_122/A POR2X1_122/Y POR2X1_122/m4_208_n4# POR2X1_122/O
+ POR2X1_122/CTRL2 POR2X1_122/a_16_28# POR2X1_122/CTRL POR2X1_122/a_76_344# POR2X1_122/a_56_344#
+ POR2X1
XPOR2X1_133 VDD GND POR2X1_8/Y POR2X1_38/B POR2X1_257/A POR2X1_133/m4_208_n4# POR2X1_133/O
+ POR2X1_133/CTRL2 POR2X1_133/a_16_28# POR2X1_133/CTRL POR2X1_133/a_76_344# POR2X1_133/a_56_344#
+ POR2X1
XPOR2X1_111 VDD GND POR2X1_32/A POR2X1_110/Y POR2X1_111/Y POR2X1_111/m4_208_n4# POR2X1_111/O
+ POR2X1_111/CTRL2 POR2X1_111/a_16_28# POR2X1_111/CTRL POR2X1_111/a_76_344# POR2X1_111/a_56_344#
+ POR2X1
XPOR2X1_144 VDD GND POR2X1_60/A POR2X1_376/B POR2X1_144/Y POR2X1_144/m4_208_n4# POR2X1_144/O
+ POR2X1_144/CTRL2 POR2X1_144/a_16_28# POR2X1_144/CTRL POR2X1_144/a_76_344# POR2X1_144/a_56_344#
+ POR2X1
XPOR2X1_155 VDD GND POR2X1_68/A POR2X1_407/A POR2X1_155/Y POR2X1_155/m4_208_n4# POR2X1_155/O
+ POR2X1_155/CTRL2 POR2X1_155/a_16_28# POR2X1_155/CTRL POR2X1_155/a_76_344# POR2X1_155/a_56_344#
+ POR2X1
XPOR2X1_166 VDD GND POR2X1_16/A POR2X1_40/Y POR2X1_166/Y POR2X1_166/m4_208_n4# POR2X1_166/O
+ POR2X1_166/CTRL2 POR2X1_166/a_16_28# POR2X1_166/CTRL POR2X1_166/a_76_344# POR2X1_166/a_56_344#
+ POR2X1
XPOR2X1_177 VDD GND POR2X1_49/Y POR2X1_72/B POR2X1_177/Y POR2X1_177/m4_208_n4# POR2X1_177/O
+ POR2X1_177/CTRL2 POR2X1_177/a_16_28# POR2X1_177/CTRL POR2X1_177/a_76_344# POR2X1_177/a_56_344#
+ POR2X1
XPOR2X1_199 VDD GND POR2X1_199/B POR2X1_196/Y POR2X1_207/B POR2X1_199/m4_208_n4# POR2X1_199/O
+ POR2X1_199/CTRL2 POR2X1_199/a_16_28# POR2X1_199/CTRL POR2X1_199/a_76_344# POR2X1_199/a_56_344#
+ POR2X1
XPOR2X1_188 VDD GND PAND2X1_39/B POR2X1_188/A POR2X1_188/Y POR2X1_733/m4_208_n4# POR2X1_188/O
+ POR2X1_188/CTRL2 POR2X1_188/a_16_28# POR2X1_188/CTRL POR2X1_188/a_76_344# POR2X1_188/a_56_344#
+ POR2X1
XPAND2X1_118 VDD GND POR2X1_78/A PAND2X1_72/A POR2X1_123/A PAND2X1_118/a_16_344# POR2X1_383/m4_208_n4#
+ PAND2X1_118/O PAND2X1_118/a_56_28# PAND2X1_118/CTRL2 PAND2X1_118/CTRL PAND2X1_118/a_76_28#
+ PAND2X1
XPAND2X1_107 VDD GND POR2X1_78/A PAND2X1_65/B POR2X1_113/A PAND2X1_107/a_16_344# PAND2X1_107/m4_208_n4#
+ PAND2X1_107/O PAND2X1_107/a_56_28# PAND2X1_107/CTRL2 PAND2X1_107/CTRL PAND2X1_107/a_76_28#
+ PAND2X1
XPAND2X1_129 VDD GND PAND2X1_90/A POR2X1_38/B POR2X1_130/A PAND2X1_129/a_16_344# PAND2X1_129/m4_208_n4#
+ PAND2X1_129/O PAND2X1_129/a_56_28# PAND2X1_129/CTRL2 PAND2X1_129/CTRL PAND2X1_129/a_76_28#
+ PAND2X1
XPOR2X1_62 VDD GND PAND2X1_9/Y POR2X1_94/A POR2X1_62/Y POR2X1_62/m4_208_n4# POR2X1_62/O
+ POR2X1_62/CTRL2 POR2X1_62/a_16_28# POR2X1_62/CTRL POR2X1_62/a_76_344# POR2X1_62/a_56_344#
+ POR2X1
XPOR2X1_40 VDD GND POR2X1_3/A POR2X1_25/Y POR2X1_40/Y POR2X1_40/m4_208_n4# POR2X1_40/O
+ POR2X1_40/CTRL2 POR2X1_40/a_16_28# POR2X1_40/CTRL POR2X1_40/a_76_344# POR2X1_40/a_56_344#
+ POR2X1
XPOR2X1_51 VDD GND POR2X1_51/B POR2X1_51/A POR2X1_52/A POR2X1_51/m4_208_n4# POR2X1_51/O
+ POR2X1_51/CTRL2 POR2X1_51/a_16_28# POR2X1_51/CTRL POR2X1_51/a_76_344# POR2X1_51/a_56_344#
+ POR2X1
XPOR2X1_84 VDD GND POR2X1_84/B POR2X1_84/A POR2X1_84/Y POR2X1_84/m4_208_n4# POR2X1_84/O
+ POR2X1_84/CTRL2 POR2X1_84/a_16_28# POR2X1_84/CTRL POR2X1_84/a_76_344# POR2X1_84/a_56_344#
+ POR2X1
XPOR2X1_73 VDD GND POR2X1_9/Y POR2X1_37/Y POR2X1_73/Y POR2X1_73/m4_208_n4# POR2X1_73/O
+ POR2X1_73/CTRL2 POR2X1_73/a_16_28# POR2X1_73/CTRL POR2X1_73/a_76_344# POR2X1_73/a_56_344#
+ POR2X1
XPOR2X1_95 VDD GND POR2X1_12/A POR2X1_51/A POR2X1_96/A POR2X1_95/m4_208_n4# POR2X1_95/O
+ POR2X1_95/CTRL2 POR2X1_95/a_16_28# POR2X1_95/CTRL POR2X1_95/a_76_344# POR2X1_95/a_56_344#
+ POR2X1
XPAND2X1_630 VDD GND PAND2X1_630/B POR2X1_628/Y PAND2X1_632/A PAND2X1_630/a_16_344#
+ PAND2X1_630/m4_208_n4# PAND2X1_630/O PAND2X1_630/a_56_28# PAND2X1_630/CTRL2 PAND2X1_630/CTRL
+ PAND2X1_630/a_76_28# PAND2X1
XPAND2X1_641 VDD GND POR2X1_265/Y PAND2X1_341/B PAND2X1_641/Y PAND2X1_641/a_16_344#
+ POR2X1_229/m4_208_n4# PAND2X1_641/O PAND2X1_641/a_56_28# PAND2X1_641/CTRL2 PAND2X1_641/CTRL
+ PAND2X1_641/a_76_28# PAND2X1
XPAND2X1_652 VDD GND PAND2X1_593/Y PAND2X1_652/A PAND2X1_652/Y PAND2X1_652/a_16_344#
+ POR2X1_594/m4_208_n4# PAND2X1_652/O PAND2X1_652/a_56_28# PAND2X1_652/CTRL2 PAND2X1_652/CTRL
+ PAND2X1_652/a_76_28# PAND2X1
XPAND2X1_674 VDD GND POR2X1_327/Y PAND2X1_72/A POR2X1_675/A PAND2X1_674/a_16_344#
+ PAND2X1_674/m4_208_n4# PAND2X1_674/O PAND2X1_674/a_56_28# PAND2X1_674/CTRL2 PAND2X1_674/CTRL
+ PAND2X1_674/a_76_28# PAND2X1
XPAND2X1_663 VDD GND PAND2X1_662/Y PAND2X1_659/Y GATE_662 PAND2X1_663/a_16_344# PAND2X1_663/m4_208_n4#
+ PAND2X1_663/O PAND2X1_663/a_56_28# PAND2X1_663/CTRL2 PAND2X1_663/CTRL PAND2X1_663/a_76_28#
+ PAND2X1
XPAND2X1_696 VDD GND POR2X1_502/A POR2X1_66/A POR2X1_708/B PAND2X1_696/a_16_344# PAND2X1_696/m4_208_n4#
+ PAND2X1_696/O PAND2X1_696/a_56_28# PAND2X1_696/CTRL2 PAND2X1_696/CTRL PAND2X1_696/a_76_28#
+ PAND2X1
XPAND2X1_685 VDD GND POR2X1_682/Y POR2X1_681/Y PAND2X1_687/A PAND2X1_685/a_16_344#
+ PAND2X1_685/m4_208_n4# PAND2X1_685/O PAND2X1_685/a_56_28# PAND2X1_685/CTRL2 PAND2X1_685/CTRL
+ PAND2X1_685/a_76_28# PAND2X1
XPAND2X1_6 VDD GND POR2X1_68/B PAND2X1_6/A PAND2X1_6/Y PAND2X1_6/a_16_344# PAND2X1_6/m4_208_n4#
+ PAND2X1_6/O PAND2X1_6/a_56_28# PAND2X1_6/CTRL2 PAND2X1_6/CTRL PAND2X1_6/a_76_28#
+ PAND2X1
XPAND2X1_482 VDD GND PAND2X1_60/B PAND2X1_6/Y POR2X1_483/A PAND2X1_482/a_16_344# PAND2X1_482/m4_208_n4#
+ PAND2X1_482/O PAND2X1_482/a_56_28# PAND2X1_482/CTRL2 PAND2X1_482/CTRL PAND2X1_482/a_76_28#
+ PAND2X1
XPAND2X1_471 VDD GND PAND2X1_471/B PAND2X1_464/Y PAND2X1_477/B PAND2X1_471/a_16_344#
+ POR2X1_237/m4_208_n4# PAND2X1_471/O PAND2X1_471/a_56_28# PAND2X1_471/CTRL2 PAND2X1_471/CTRL
+ PAND2X1_471/a_76_28# PAND2X1
XPAND2X1_460 VDD GND POR2X1_409/Y POR2X1_380/Y PAND2X1_460/Y PAND2X1_460/a_16_344#
+ PAND2X1_460/m4_208_n4# PAND2X1_460/O PAND2X1_460/a_56_28# PAND2X1_460/CTRL2 PAND2X1_460/CTRL
+ PAND2X1_460/a_76_28# PAND2X1
XPAND2X1_493 VDD GND POR2X1_492/Y POR2X1_491/Y PAND2X1_493/Y PAND2X1_493/a_16_344#
+ PAND2X1_493/m4_208_n4# PAND2X1_493/O PAND2X1_493/a_56_28# PAND2X1_493/CTRL2 PAND2X1_493/CTRL
+ PAND2X1_493/a_76_28# PAND2X1
XPAND2X1_290 VDD GND POR2X1_66/A POR2X1_78/B POR2X1_334/B PAND2X1_290/a_16_344# PAND2X1_290/m4_208_n4#
+ PAND2X1_290/O PAND2X1_290/a_56_28# PAND2X1_290/CTRL2 PAND2X1_290/CTRL PAND2X1_290/a_76_28#
+ PAND2X1
XPOR2X1_507 VDD GND POR2X1_507/B POR2X1_507/A POR2X1_508/A POR2X1_507/m4_208_n4# POR2X1_507/O
+ POR2X1_507/CTRL2 POR2X1_507/a_16_28# POR2X1_507/CTRL POR2X1_507/a_76_344# POR2X1_507/a_56_344#
+ POR2X1
XPOR2X1_518 VDD GND POR2X1_65/A POR2X1_73/Y POR2X1_518/Y POR2X1_518/m4_208_n4# POR2X1_518/O
+ POR2X1_518/CTRL2 POR2X1_518/a_16_28# POR2X1_518/CTRL POR2X1_518/a_76_344# POR2X1_518/a_56_344#
+ POR2X1
XPOR2X1_529 VDD GND D_INPUT_3 POR2X1_83/B POR2X1_529/Y POR2X1_529/m4_208_n4# POR2X1_529/O
+ POR2X1_529/CTRL2 POR2X1_529/a_16_28# POR2X1_529/CTRL POR2X1_529/a_76_344# POR2X1_529/a_56_344#
+ POR2X1
XPOR2X1_315 VDD GND POR2X1_32/A POR2X1_257/A POR2X1_315/Y POR2X1_315/m4_208_n4# POR2X1_315/O
+ POR2X1_315/CTRL2 POR2X1_315/a_16_28# POR2X1_315/CTRL POR2X1_315/a_76_344# POR2X1_315/a_56_344#
+ POR2X1
XPOR2X1_326 VDD GND POR2X1_324/Y POR2X1_326/A POR2X1_854/B POR2X1_324/m4_208_n4# POR2X1_326/O
+ POR2X1_326/CTRL2 POR2X1_326/a_16_28# POR2X1_326/CTRL POR2X1_326/a_76_344# POR2X1_326/a_56_344#
+ POR2X1
XPOR2X1_304 VDD GND POR2X1_56/B POR2X1_236/Y POR2X1_304/Y POR2X1_304/m4_208_n4# POR2X1_304/O
+ POR2X1_304/CTRL2 POR2X1_304/a_16_28# POR2X1_304/CTRL POR2X1_304/a_76_344# POR2X1_304/a_56_344#
+ POR2X1
XPOR2X1_348 VDD GND POR2X1_344/Y POR2X1_348/A POR2X1_359/B POR2X1_348/m4_208_n4# POR2X1_348/O
+ POR2X1_348/CTRL2 POR2X1_348/a_16_28# POR2X1_348/CTRL POR2X1_348/a_76_344# POR2X1_348/a_56_344#
+ POR2X1
XPOR2X1_359 VDD GND POR2X1_359/B POR2X1_349/Y POR2X1_359/Y POR2X1_359/m4_208_n4# POR2X1_359/O
+ POR2X1_359/CTRL2 POR2X1_359/a_16_28# POR2X1_359/CTRL POR2X1_359/a_76_344# POR2X1_359/a_56_344#
+ POR2X1
XPOR2X1_337 VDD GND POR2X1_335/Y POR2X1_337/A POR2X1_337/Y POR2X1_337/m4_208_n4# POR2X1_337/O
+ POR2X1_337/CTRL2 POR2X1_337/a_16_28# POR2X1_337/CTRL POR2X1_337/a_76_344# POR2X1_337/a_56_344#
+ POR2X1
XPOR2X1_860 VDD GND POR2X1_244/Y POR2X1_860/A POR2X1_861/A POR2X1_860/m4_208_n4# POR2X1_860/O
+ POR2X1_860/CTRL2 POR2X1_860/a_16_28# POR2X1_860/CTRL POR2X1_860/a_76_344# POR2X1_860/a_56_344#
+ POR2X1
XPAND2X1_801 VDD GND PAND2X1_801/B POR2X1_761/Y PAND2X1_809/A PAND2X1_801/a_16_344#
+ PAND2X1_801/m4_208_n4# PAND2X1_801/O PAND2X1_801/a_56_28# PAND2X1_801/CTRL2 PAND2X1_801/CTRL
+ PAND2X1_801/a_76_28# PAND2X1
XPAND2X1_812 VDD GND PAND2X1_811/Y PAND2X1_812/A GATE_811 PAND2X1_812/a_16_344# PAND2X1_811/m4_208_n4#
+ PAND2X1_812/O PAND2X1_812/a_56_28# PAND2X1_812/CTRL2 PAND2X1_812/CTRL PAND2X1_812/a_76_28#
+ PAND2X1
XPAND2X1_823 VDD GND POR2X1_383/A PAND2X1_52/B POR2X1_836/B PAND2X1_823/a_16_344#
+ POR2X1_852/m4_208_n4# PAND2X1_823/O PAND2X1_823/a_56_28# PAND2X1_823/CTRL2 PAND2X1_823/CTRL
+ PAND2X1_823/a_76_28# PAND2X1
XPAND2X1_834 VDD GND POR2X1_677/Y POR2X1_511/Y PAND2X1_840/B PAND2X1_834/a_16_344#
+ PAND2X1_834/m4_208_n4# PAND2X1_834/O PAND2X1_834/a_56_28# PAND2X1_834/CTRL2 PAND2X1_834/CTRL
+ PAND2X1_834/a_76_28# PAND2X1
XPAND2X1_845 VDD GND POR2X1_813/Y PAND2X1_673/Y PAND2X1_849/B PAND2X1_845/a_16_344#
+ PAND2X1_845/m4_208_n4# PAND2X1_845/O PAND2X1_845/a_56_28# PAND2X1_845/CTRL2 PAND2X1_845/CTRL
+ PAND2X1_845/a_76_28# PAND2X1
XPAND2X1_856 VDD GND PAND2X1_856/B PAND2X1_854/Y PAND2X1_863/A PAND2X1_856/a_16_344#
+ PAND2X1_856/m4_208_n4# PAND2X1_856/O PAND2X1_856/a_56_28# PAND2X1_856/CTRL2 PAND2X1_856/CTRL
+ PAND2X1_856/a_76_28# PAND2X1
XPOR2X1_101 VDD GND POR2X1_99/Y POR2X1_101/A POR2X1_101/Y POR2X1_101/m4_208_n4# POR2X1_101/O
+ POR2X1_101/CTRL2 POR2X1_101/a_16_28# POR2X1_101/CTRL POR2X1_101/a_76_344# POR2X1_101/a_56_344#
+ POR2X1
XPOR2X1_112 VDD GND POR2X1_775/A POR2X1_332/B POR2X1_112/Y POR2X1_112/m4_208_n4# POR2X1_112/O
+ POR2X1_112/CTRL2 POR2X1_112/a_16_28# POR2X1_112/CTRL POR2X1_112/a_76_344# POR2X1_112/a_56_344#
+ POR2X1
XPOR2X1_123 VDD GND POR2X1_123/B POR2X1_123/A POR2X1_123/Y POR2X1_123/m4_208_n4# POR2X1_123/O
+ POR2X1_123/CTRL2 POR2X1_123/a_16_28# POR2X1_123/CTRL POR2X1_123/a_76_344# POR2X1_123/a_56_344#
+ POR2X1
XPOR2X1_134 VDD GND POR2X1_96/A POR2X1_257/A POR2X1_134/Y POR2X1_134/m4_208_n4# POR2X1_134/O
+ POR2X1_134/CTRL2 POR2X1_134/a_16_28# POR2X1_134/CTRL POR2X1_134/a_76_344# POR2X1_134/a_56_344#
+ POR2X1
XPOR2X1_156 VDD GND POR2X1_156/B POR2X1_155/Y POR2X1_156/Y POR2X1_156/m4_208_n4# POR2X1_156/O
+ POR2X1_156/CTRL2 POR2X1_156/a_16_28# POR2X1_156/CTRL POR2X1_156/a_76_344# POR2X1_156/a_56_344#
+ POR2X1
XPOR2X1_145 VDD GND POR2X1_52/A POR2X1_77/Y POR2X1_145/Y POR2X1_145/m4_208_n4# POR2X1_145/O
+ POR2X1_145/CTRL2 POR2X1_145/a_16_28# POR2X1_145/CTRL POR2X1_145/a_76_344# POR2X1_145/a_56_344#
+ POR2X1
XPOR2X1_167 VDD GND POR2X1_65/A POR2X1_669/B POR2X1_167/Y POR2X1_167/m4_208_n4# POR2X1_167/O
+ POR2X1_167/CTRL2 POR2X1_167/a_16_28# POR2X1_167/CTRL POR2X1_167/a_76_344# POR2X1_167/a_56_344#
+ POR2X1
XPOR2X1_189 VDD GND POR2X1_96/A POR2X1_498/A POR2X1_189/Y POR2X1_189/m4_208_n4# POR2X1_189/O
+ POR2X1_189/CTRL2 POR2X1_189/a_16_28# POR2X1_189/CTRL POR2X1_189/a_76_344# POR2X1_189/a_56_344#
+ POR2X1
XPOR2X1_178 VDD GND POR2X1_55/Y POR2X1_416/B POR2X1_178/Y POR2X1_178/m4_208_n4# POR2X1_178/O
+ POR2X1_178/CTRL2 POR2X1_178/a_16_28# POR2X1_178/CTRL POR2X1_178/a_76_344# POR2X1_178/a_56_344#
+ POR2X1
XPAND2X1_108 VDD GND POR2X1_590/A PAND2X1_60/B POR2X1_114/B PAND2X1_108/a_16_344#
+ PAND2X1_108/m4_208_n4# PAND2X1_108/O PAND2X1_108/a_56_28# PAND2X1_108/CTRL2 PAND2X1_108/CTRL
+ PAND2X1_108/a_76_28# PAND2X1
XPAND2X1_119 VDD GND PAND2X1_94/A INPUT_1 POR2X1_121/B PAND2X1_119/a_16_344# PAND2X1_119/m4_208_n4#
+ PAND2X1_119/O PAND2X1_119/a_56_28# PAND2X1_119/CTRL2 PAND2X1_119/CTRL PAND2X1_119/a_76_28#
+ PAND2X1
XPOR2X1_41 VDD GND POR2X1_41/B POR2X1_40/Y POR2X1_41/Y POR2X1_41/m4_208_n4# POR2X1_41/O
+ POR2X1_41/CTRL2 POR2X1_41/a_16_28# POR2X1_41/CTRL POR2X1_41/a_76_344# POR2X1_41/a_56_344#
+ POR2X1
XPOR2X1_52 VDD GND POR2X1_49/Y POR2X1_52/A POR2X1_52/Y POR2X1_52/m4_208_n4# POR2X1_52/O
+ POR2X1_52/CTRL2 POR2X1_52/a_16_28# POR2X1_52/CTRL POR2X1_52/a_76_344# POR2X1_52/a_56_344#
+ POR2X1
XPOR2X1_30 VDD GND D_INPUT_4 D_INPUT_5 POR2X1_51/B POR2X1_30/m4_208_n4# POR2X1_30/O
+ POR2X1_30/CTRL2 POR2X1_30/a_16_28# POR2X1_30/CTRL POR2X1_30/a_76_344# POR2X1_30/a_56_344#
+ POR2X1
XPOR2X1_96 VDD GND POR2X1_96/B POR2X1_96/A POR2X1_96/Y POR2X1_96/m4_208_n4# POR2X1_96/O
+ POR2X1_96/CTRL2 POR2X1_96/a_16_28# POR2X1_96/CTRL POR2X1_96/a_76_344# POR2X1_96/a_56_344#
+ POR2X1
XPOR2X1_85 VDD GND POR2X1_20/B POR2X1_37/Y POR2X1_85/Y POR2X1_85/m4_208_n4# POR2X1_85/O
+ POR2X1_85/CTRL2 POR2X1_85/a_16_28# POR2X1_85/CTRL POR2X1_85/a_76_344# POR2X1_85/a_56_344#
+ POR2X1
XPOR2X1_63 VDD GND POR2X1_8/Y POR2X1_62/Y POR2X1_63/Y POR2X1_63/m4_208_n4# POR2X1_63/O
+ POR2X1_63/CTRL2 POR2X1_63/a_16_28# POR2X1_63/CTRL POR2X1_63/a_76_344# POR2X1_63/a_56_344#
+ POR2X1
XPOR2X1_74 VDD GND POR2X1_32/A POR2X1_73/Y POR2X1_74/Y POR2X1_74/m4_208_n4# POR2X1_74/O
+ POR2X1_74/CTRL2 POR2X1_74/a_16_28# POR2X1_74/CTRL POR2X1_74/a_76_344# POR2X1_74/a_56_344#
+ POR2X1
XPOR2X1_690 VDD GND INPUT_0 POR2X1_413/A POR2X1_690/Y POR2X1_690/m4_208_n4# POR2X1_690/O
+ POR2X1_690/CTRL2 POR2X1_690/a_16_28# POR2X1_690/CTRL POR2X1_690/a_76_344# POR2X1_690/a_56_344#
+ POR2X1
XPAND2X1_631 VDD GND POR2X1_625/Y PAND2X1_631/A PAND2X1_632/B PAND2X1_631/a_16_344#
+ PAND2X1_631/m4_208_n4# PAND2X1_631/O PAND2X1_631/a_56_28# PAND2X1_631/CTRL2 PAND2X1_631/CTRL
+ PAND2X1_631/a_76_28# PAND2X1
XPAND2X1_620 VDD GND POR2X1_613/Y POR2X1_528/Y PAND2X1_620/Y PAND2X1_620/a_16_344#
+ PAND2X1_620/m4_208_n4# PAND2X1_620/O PAND2X1_620/a_56_28# PAND2X1_620/CTRL2 PAND2X1_620/CTRL
+ PAND2X1_620/a_76_28# PAND2X1
XPAND2X1_653 VDD GND PAND2X1_652/Y POR2X1_594/Y PAND2X1_653/Y PAND2X1_653/a_16_344#
+ PAND2X1_653/m4_208_n4# PAND2X1_653/O PAND2X1_653/a_56_28# PAND2X1_653/CTRL2 PAND2X1_653/CTRL
+ PAND2X1_653/a_76_28# PAND2X1
XPAND2X1_664 VDD GND POR2X1_77/Y POR2X1_73/Y POR2X1_665/A PAND2X1_664/a_16_344# PAND2X1_664/m4_208_n4#
+ PAND2X1_664/O PAND2X1_664/a_56_28# PAND2X1_664/CTRL2 PAND2X1_664/CTRL PAND2X1_664/a_76_28#
+ PAND2X1
XPAND2X1_642 VDD GND PAND2X1_642/B POR2X1_416/Y PAND2X1_649/A PAND2X1_642/a_16_344#
+ PAND2X1_642/m4_208_n4# PAND2X1_642/O PAND2X1_642/a_56_28# PAND2X1_642/CTRL2 PAND2X1_642/CTRL
+ PAND2X1_642/a_76_28# PAND2X1
XPAND2X1_675 VDD GND POR2X1_674/Y PAND2X1_675/A PAND2X1_736/A PAND2X1_675/a_16_344#
+ PAND2X1_675/m4_208_n4# PAND2X1_675/O PAND2X1_675/a_56_28# PAND2X1_675/CTRL2 PAND2X1_675/CTRL
+ PAND2X1_675/a_76_28# PAND2X1
XPAND2X1_697 VDD GND POR2X1_383/A POR2X1_260/A POR2X1_779/A PAND2X1_697/a_16_344#
+ PAND2X1_697/m4_208_n4# PAND2X1_697/O PAND2X1_697/a_56_28# PAND2X1_697/CTRL2 PAND2X1_697/CTRL
+ PAND2X1_697/a_76_28# PAND2X1
XPAND2X1_686 VDD GND POR2X1_684/Y POR2X1_683/Y PAND2X1_687/B PAND2X1_686/a_16_344#
+ PAND2X1_686/m4_208_n4# PAND2X1_686/O PAND2X1_686/a_56_28# PAND2X1_686/CTRL2 PAND2X1_686/CTRL
+ PAND2X1_686/a_76_28# PAND2X1
XPAND2X1_7 VDD GND PAND2X1_6/Y POR2X1_66/B PAND2X1_7/Y PAND2X1_7/a_16_344# PAND2X1_7/m4_208_n4#
+ PAND2X1_7/O PAND2X1_7/a_56_28# PAND2X1_7/CTRL2 PAND2X1_7/CTRL PAND2X1_7/a_76_28#
+ PAND2X1
XPAND2X1_450 VDD GND POR2X1_427/Y POR2X1_426/Y PAND2X1_452/A PAND2X1_450/a_16_344#
+ PAND2X1_450/m4_208_n4# PAND2X1_450/O PAND2X1_450/a_56_28# PAND2X1_450/CTRL2 PAND2X1_450/CTRL
+ PAND2X1_450/a_76_28# PAND2X1
XPAND2X1_472 VDD GND PAND2X1_472/B PAND2X1_472/A PAND2X1_476/A PAND2X1_472/a_16_344#
+ PAND2X1_472/m4_208_n4# PAND2X1_472/O PAND2X1_472/a_56_28# PAND2X1_472/CTRL2 PAND2X1_472/CTRL
+ PAND2X1_472/a_76_28# PAND2X1
XPAND2X1_461 VDD GND POR2X1_413/Y POR2X1_411/Y PAND2X1_462/B PAND2X1_461/a_16_344#
+ PAND2X1_461/m4_208_n4# PAND2X1_461/O PAND2X1_461/a_56_28# PAND2X1_461/CTRL2 PAND2X1_461/CTRL
+ PAND2X1_461/a_76_28# PAND2X1
XPAND2X1_494 VDD GND POR2X1_383/Y POR2X1_260/B POR2X1_558/A PAND2X1_494/a_16_344#
+ PAND2X1_494/m4_208_n4# PAND2X1_494/O PAND2X1_494/a_56_28# PAND2X1_494/CTRL2 PAND2X1_494/CTRL
+ PAND2X1_494/a_76_28# PAND2X1
XPAND2X1_483 VDD GND POR2X1_482/Y POR2X1_252/Y PAND2X1_631/A PAND2X1_483/a_16_344#
+ PAND2X1_483/m4_208_n4# PAND2X1_483/O PAND2X1_483/a_56_28# PAND2X1_483/CTRL2 PAND2X1_483/CTRL
+ PAND2X1_483/a_76_28# PAND2X1
XPAND2X1_280 VDD GND POR2X1_383/A PAND2X1_48/B POR2X1_542/B PAND2X1_280/a_16_344#
+ PAND2X1_280/m4_208_n4# PAND2X1_280/O PAND2X1_280/a_56_28# PAND2X1_280/CTRL2 PAND2X1_280/CTRL
+ PAND2X1_280/a_76_28# PAND2X1
XPAND2X1_291 VDD GND PAND2X1_824/B PAND2X1_69/A POR2X1_334/A PAND2X1_291/a_16_344#
+ PAND2X1_291/m4_208_n4# PAND2X1_291/O PAND2X1_291/a_56_28# PAND2X1_291/CTRL2 PAND2X1_291/CTRL
+ PAND2X1_291/a_76_28# PAND2X1
XPOR2X1_508 VDD GND POR2X1_508/B POR2X1_508/A POR2X1_510/B POR2X1_508/m4_208_n4# POR2X1_508/O
+ POR2X1_508/CTRL2 POR2X1_508/a_16_28# POR2X1_508/CTRL POR2X1_508/a_76_344# POR2X1_508/a_56_344#
+ POR2X1
XPOR2X1_519 VDD GND POR2X1_46/Y POR2X1_416/B POR2X1_519/Y POR2X1_519/m4_208_n4# POR2X1_519/O
+ POR2X1_519/CTRL2 POR2X1_519/a_16_28# POR2X1_519/CTRL POR2X1_519/a_76_344# POR2X1_519/a_56_344#
+ POR2X1
XPOR2X1_316 VDD GND POR2X1_13/A POR2X1_81/A POR2X1_316/Y POR2X1_316/m4_208_n4# POR2X1_316/O
+ POR2X1_316/CTRL2 POR2X1_316/a_16_28# POR2X1_316/CTRL POR2X1_316/a_76_344# POR2X1_316/a_56_344#
+ POR2X1
XPOR2X1_305 VDD GND POR2X1_7/B POR2X1_90/Y POR2X1_305/Y POR2X1_305/m4_208_n4# POR2X1_305/O
+ POR2X1_305/CTRL2 POR2X1_305/a_16_28# POR2X1_305/CTRL POR2X1_305/a_76_344# POR2X1_305/a_56_344#
+ POR2X1
XPOR2X1_338 VDD GND POR2X1_333/Y POR2X1_334/Y POR2X1_351/B POR2X1_338/m4_208_n4# POR2X1_338/O
+ POR2X1_338/CTRL2 POR2X1_338/a_16_28# POR2X1_338/CTRL POR2X1_338/a_76_344# POR2X1_338/a_56_344#
+ POR2X1
XPOR2X1_349 VDD GND POR2X1_342/Y POR2X1_343/Y POR2X1_349/Y POR2X1_349/m4_208_n4# POR2X1_349/O
+ POR2X1_349/CTRL2 POR2X1_349/a_16_28# POR2X1_349/CTRL POR2X1_349/a_76_344# POR2X1_349/a_56_344#
+ POR2X1
XPOR2X1_327 VDD GND PAND2X1_63/Y POR2X1_264/Y POR2X1_327/Y POR2X1_327/m4_208_n4# POR2X1_327/O
+ POR2X1_327/CTRL2 POR2X1_327/a_16_28# POR2X1_327/CTRL POR2X1_327/a_76_344# POR2X1_327/a_56_344#
+ POR2X1
XPOR2X1_861 VDD GND POR2X1_624/Y POR2X1_861/A POR2X1_865/B POR2X1_861/m4_208_n4# POR2X1_861/O
+ POR2X1_861/CTRL2 POR2X1_861/a_16_28# POR2X1_861/CTRL POR2X1_861/a_76_344# POR2X1_861/a_56_344#
+ POR2X1
XPOR2X1_850 VDD GND POR2X1_850/B POR2X1_850/A POR2X1_858/B POR2X1_850/m4_208_n4# POR2X1_850/O
+ POR2X1_850/CTRL2 POR2X1_850/a_16_28# POR2X1_850/CTRL POR2X1_850/a_76_344# POR2X1_850/a_56_344#
+ POR2X1
XPAND2X1_813 VDD GND POR2X1_266/A POR2X1_62/Y POR2X1_845/A PAND2X1_813/a_16_344# POR2X1_845/m4_208_n4#
+ PAND2X1_813/O PAND2X1_813/a_56_28# PAND2X1_813/CTRL2 PAND2X1_813/CTRL PAND2X1_813/a_76_28#
+ PAND2X1
XPAND2X1_802 VDD GND PAND2X1_802/B PAND2X1_798/Y PAND2X1_809/B PAND2X1_802/a_16_344#
+ PAND2X1_802/m4_208_n4# PAND2X1_802/O PAND2X1_802/a_56_28# PAND2X1_802/CTRL2 PAND2X1_802/CTRL
+ PAND2X1_802/a_76_28# PAND2X1
XPAND2X1_846 VDD GND POR2X1_816/Y POR2X1_815/Y PAND2X1_848/A PAND2X1_846/a_16_344#
+ PAND2X1_846/m4_208_n4# PAND2X1_846/O PAND2X1_846/a_56_28# PAND2X1_846/CTRL2 PAND2X1_846/CTRL
+ PAND2X1_846/a_76_28# PAND2X1
XPAND2X1_835 VDD GND POR2X1_822/Y POR2X1_821/Y PAND2X1_835/Y PAND2X1_835/a_16_344#
+ PAND2X1_835/m4_208_n4# PAND2X1_835/O PAND2X1_835/a_56_28# PAND2X1_835/CTRL2 PAND2X1_835/CTRL
+ PAND2X1_835/a_76_28# PAND2X1
XPAND2X1_824 VDD GND PAND2X1_824/B POR2X1_66/A POR2X1_836/A PAND2X1_824/a_16_344#
+ PAND2X1_824/m4_208_n4# PAND2X1_824/O PAND2X1_824/a_56_28# PAND2X1_824/CTRL2 PAND2X1_824/CTRL
+ PAND2X1_824/a_76_28# PAND2X1
XPAND2X1_857 VDD GND PAND2X1_857/B PAND2X1_857/A PAND2X1_863/B PAND2X1_857/a_16_344#
+ PAND2X1_857/m4_208_n4# PAND2X1_857/O PAND2X1_857/a_56_28# PAND2X1_857/CTRL2 PAND2X1_857/CTRL
+ PAND2X1_857/a_76_28# PAND2X1
XPOR2X1_102 VDD GND POR2X1_8/Y POR2X1_54/Y POR2X1_102/Y POR2X1_102/m4_208_n4# POR2X1_102/O
+ POR2X1_102/CTRL2 POR2X1_102/a_16_28# POR2X1_102/CTRL POR2X1_102/a_76_344# POR2X1_102/a_56_344#
+ POR2X1
XPOR2X1_124 VDD GND POR2X1_124/B POR2X1_123/Y POR2X1_572/B POR2X1_124/m4_208_n4# POR2X1_124/O
+ POR2X1_124/CTRL2 POR2X1_124/a_16_28# POR2X1_124/CTRL POR2X1_124/a_76_344# POR2X1_124/a_56_344#
+ POR2X1
XPOR2X1_113 VDD GND POR2X1_113/B POR2X1_113/A POR2X1_113/Y POR2X1_113/m4_208_n4# POR2X1_113/O
+ POR2X1_113/CTRL2 POR2X1_113/a_16_28# POR2X1_113/CTRL POR2X1_113/a_76_344# POR2X1_113/a_56_344#
+ POR2X1
XPOR2X1_168 VDD GND POR2X1_776/B POR2X1_168/A POR2X1_170/B POR2X1_168/m4_208_n4# POR2X1_168/O
+ POR2X1_168/CTRL2 POR2X1_168/a_16_28# POR2X1_168/CTRL POR2X1_168/a_76_344# POR2X1_168/a_56_344#
+ POR2X1
XPOR2X1_157 VDD GND POR2X1_3/A POR2X1_36/B POR2X1_416/B POR2X1_157/m4_208_n4# POR2X1_157/O
+ POR2X1_157/CTRL2 POR2X1_157/a_16_28# POR2X1_157/CTRL POR2X1_157/a_76_344# POR2X1_157/a_56_344#
+ POR2X1
XPOR2X1_146 VDD GND POR2X1_39/B POR2X1_394/A POR2X1_146/Y POR2X1_146/m4_208_n4# POR2X1_146/O
+ POR2X1_146/CTRL2 POR2X1_146/a_16_28# POR2X1_146/CTRL POR2X1_146/a_76_344# POR2X1_146/a_56_344#
+ POR2X1
XPOR2X1_135 VDD GND POR2X1_60/A POR2X1_257/A POR2X1_135/Y POR2X1_135/m4_208_n4# POR2X1_135/O
+ POR2X1_135/CTRL2 POR2X1_135/a_16_28# POR2X1_135/CTRL POR2X1_135/a_76_344# POR2X1_135/a_56_344#
+ POR2X1
XPOR2X1_179 VDD GND POR2X1_39/B POR2X1_411/B POR2X1_179/Y POR2X1_311/m4_208_n4# POR2X1_179/O
+ POR2X1_179/CTRL2 POR2X1_179/a_16_28# POR2X1_179/CTRL POR2X1_179/a_76_344# POR2X1_179/a_56_344#
+ POR2X1
XPAND2X1_109 VDD GND POR2X1_78/A PAND2X1_32/B POR2X1_775/A PAND2X1_109/a_16_344# PAND2X1_109/m4_208_n4#
+ PAND2X1_109/O PAND2X1_109/a_56_28# PAND2X1_109/CTRL2 PAND2X1_109/CTRL PAND2X1_109/a_76_28#
+ PAND2X1
XPOR2X1_20 VDD GND POR2X1_20/B POR2X1_20/A POR2X1_20/Y POR2X1_20/m4_208_n4# POR2X1_20/O
+ POR2X1_20/CTRL2 POR2X1_20/a_16_28# POR2X1_20/CTRL POR2X1_20/a_76_344# POR2X1_20/a_56_344#
+ POR2X1
XPOR2X1_42 VDD GND D_INPUT_1 POR2X1_37/Y POR2X1_42/Y POR2X1_42/m4_208_n4# POR2X1_42/O
+ POR2X1_42/CTRL2 POR2X1_42/a_16_28# POR2X1_42/CTRL POR2X1_42/a_76_344# POR2X1_42/a_56_344#
+ POR2X1
XPOR2X1_31 VDD GND POR2X1_3/B POR2X1_51/B POR2X1_32/A POR2X1_31/m4_208_n4# POR2X1_31/O
+ POR2X1_31/CTRL2 POR2X1_31/a_16_28# POR2X1_31/CTRL POR2X1_31/a_76_344# POR2X1_31/a_56_344#
+ POR2X1
XPOR2X1_53 VDD GND INPUT_5 POR2X1_51/A POR2X1_56/B POR2X1_53/m4_208_n4# POR2X1_53/O
+ POR2X1_53/CTRL2 POR2X1_53/a_16_28# POR2X1_53/CTRL POR2X1_53/a_76_344# POR2X1_53/a_56_344#
+ POR2X1
XPOR2X1_86 VDD GND D_INPUT_0 POR2X1_85/Y POR2X1_86/Y POR2X1_86/m4_208_n4# POR2X1_86/O
+ POR2X1_86/CTRL2 POR2X1_86/a_16_28# POR2X1_86/CTRL POR2X1_86/a_76_344# POR2X1_86/a_56_344#
+ POR2X1
XPOR2X1_64 VDD GND POR2X1_22/A POR2X1_51/A POR2X1_65/A POR2X1_64/m4_208_n4# POR2X1_64/O
+ POR2X1_64/CTRL2 POR2X1_64/a_16_28# POR2X1_64/CTRL POR2X1_64/a_76_344# POR2X1_64/a_56_344#
+ POR2X1
XPOR2X1_75 VDD GND POR2X1_23/Y POR2X1_60/A POR2X1_75/Y POR2X1_75/m4_208_n4# POR2X1_75/O
+ POR2X1_75/CTRL2 POR2X1_75/a_16_28# POR2X1_75/CTRL POR2X1_75/a_76_344# POR2X1_75/a_56_344#
+ POR2X1
XPOR2X1_97 VDD GND POR2X1_97/B POR2X1_97/A POR2X1_99/B POR2X1_97/m4_208_n4# POR2X1_97/O
+ POR2X1_97/CTRL2 POR2X1_97/a_16_28# POR2X1_97/CTRL POR2X1_97/a_76_344# POR2X1_97/a_56_344#
+ POR2X1
XPOR2X1_680 VDD GND POR2X1_52/A POR2X1_594/A POR2X1_680/Y POR2X1_680/m4_208_n4# POR2X1_680/O
+ POR2X1_680/CTRL2 POR2X1_680/a_16_28# POR2X1_680/CTRL POR2X1_680/a_76_344# POR2X1_680/a_56_344#
+ POR2X1
XPOR2X1_691 VDD GND POR2X1_691/B POR2X1_691/A POR2X1_855/B POR2X1_691/m4_208_n4# POR2X1_691/O
+ POR2X1_691/CTRL2 POR2X1_691/a_16_28# POR2X1_691/CTRL POR2X1_691/a_76_344# POR2X1_691/a_56_344#
+ POR2X1
XPAND2X1_621 VDD GND POR2X1_617/Y POR2X1_616/Y PAND2X1_621/Y PAND2X1_621/a_16_344#
+ PAND2X1_621/m4_208_n4# PAND2X1_621/O PAND2X1_621/a_56_28# PAND2X1_621/CTRL2 PAND2X1_621/CTRL
+ PAND2X1_621/a_76_28# PAND2X1
XPAND2X1_610 VDD GND POR2X1_48/A POR2X1_40/Y POR2X1_612/B PAND2X1_610/a_16_344# PAND2X1_610/m4_208_n4#
+ PAND2X1_610/O PAND2X1_610/a_56_28# PAND2X1_610/CTRL2 PAND2X1_610/CTRL PAND2X1_610/a_76_28#
+ PAND2X1
XPAND2X1_643 VDD GND POR2X1_595/Y PAND2X1_643/A PAND2X1_643/Y PAND2X1_643/a_16_344#
+ PAND2X1_643/m4_208_n4# PAND2X1_643/O PAND2X1_643/a_56_28# PAND2X1_643/CTRL2 PAND2X1_643/CTRL
+ PAND2X1_643/a_76_28# PAND2X1
XPAND2X1_632 VDD GND PAND2X1_632/B PAND2X1_632/A PAND2X1_658/B PAND2X1_632/a_16_344#
+ PAND2X1_632/m4_208_n4# PAND2X1_632/O PAND2X1_632/a_56_28# PAND2X1_632/CTRL2 PAND2X1_632/CTRL
+ PAND2X1_632/a_76_28# PAND2X1
XPAND2X1_665 VDD GND POR2X1_664/Y POR2X1_66/B POR2X1_719/B PAND2X1_665/a_16_344# PAND2X1_665/m4_208_n4#
+ PAND2X1_665/O PAND2X1_665/a_56_28# PAND2X1_665/CTRL2 PAND2X1_665/CTRL PAND2X1_665/a_76_28#
+ PAND2X1
XPAND2X1_654 VDD GND PAND2X1_651/Y PAND2X1_654/A PAND2X1_661/B PAND2X1_654/a_16_344#
+ PAND2X1_654/m4_208_n4# PAND2X1_654/O PAND2X1_654/a_56_28# PAND2X1_654/CTRL2 PAND2X1_654/CTRL
+ PAND2X1_654/a_76_28# PAND2X1
XPAND2X1_676 VDD GND POR2X1_599/A POR2X1_257/A POR2X1_679/B PAND2X1_676/a_16_344#
+ PAND2X1_676/m4_208_n4# PAND2X1_676/O PAND2X1_676/a_56_28# PAND2X1_676/CTRL2 PAND2X1_676/CTRL
+ PAND2X1_676/a_76_28# PAND2X1
XPAND2X1_698 VDD GND POR2X1_532/A PAND2X1_65/B POR2X1_709/B PAND2X1_698/a_16_344#
+ PAND2X1_698/m4_208_n4# PAND2X1_698/O PAND2X1_698/a_56_28# PAND2X1_698/CTRL2 PAND2X1_698/CTRL
+ PAND2X1_698/a_76_28# PAND2X1
XPAND2X1_687 VDD GND PAND2X1_687/B PAND2X1_687/A PAND2X1_687/Y PAND2X1_687/a_16_344#
+ PAND2X1_687/m4_208_n4# PAND2X1_687/O PAND2X1_687/a_56_28# PAND2X1_687/CTRL2 PAND2X1_687/CTRL
+ PAND2X1_687/a_76_28# PAND2X1
XPAND2X1_8 VDD GND D_INPUT_3 INPUT_2 PAND2X1_8/Y PAND2X1_8/a_16_344# PAND2X1_8/m4_208_n4#
+ PAND2X1_8/O PAND2X1_8/a_56_28# PAND2X1_8/CTRL2 PAND2X1_8/CTRL PAND2X1_8/a_76_28#
+ PAND2X1
XPAND2X1_440 VDD GND PAND2X1_675/A POR2X1_437/Y PAND2X1_652/A PAND2X1_440/a_16_344#
+ PAND2X1_440/m4_208_n4# PAND2X1_440/O PAND2X1_440/a_56_28# PAND2X1_440/CTRL2 PAND2X1_440/CTRL
+ PAND2X1_440/a_76_28# PAND2X1
XPAND2X1_473 VDD GND PAND2X1_473/B PAND2X1_216/B PAND2X1_473/Y PAND2X1_473/a_16_344#
+ PAND2X1_473/m4_208_n4# PAND2X1_473/O PAND2X1_473/a_56_28# PAND2X1_473/CTRL2 PAND2X1_473/CTRL
+ PAND2X1_473/a_76_28# PAND2X1
XPAND2X1_451 VDD GND POR2X1_430/Y POR2X1_428/Y PAND2X1_452/B PAND2X1_451/a_16_344#
+ PAND2X1_451/m4_208_n4# PAND2X1_451/O PAND2X1_451/a_56_28# PAND2X1_451/CTRL2 PAND2X1_451/CTRL
+ PAND2X1_451/a_76_28# PAND2X1
XPAND2X1_462 VDD GND PAND2X1_462/B POR2X1_416/Y PAND2X1_472/A PAND2X1_462/a_16_344#
+ PAND2X1_462/m4_208_n4# PAND2X1_462/O PAND2X1_462/a_56_28# PAND2X1_462/CTRL2 PAND2X1_462/CTRL
+ PAND2X1_462/a_76_28# PAND2X1
XPAND2X1_495 VDD GND PAND2X1_55/Y PAND2X1_69/A POR2X1_833/A PAND2X1_495/a_16_344#
+ PAND2X1_495/m4_208_n4# PAND2X1_495/O PAND2X1_495/a_56_28# PAND2X1_495/CTRL2 PAND2X1_495/CTRL
+ PAND2X1_495/a_76_28# PAND2X1
XPAND2X1_484 VDD GND PAND2X1_69/A POR2X1_294/B POR2X1_486/B PAND2X1_484/a_16_344#
+ PAND2X1_484/m4_208_n4# PAND2X1_484/O PAND2X1_484/a_56_28# PAND2X1_484/CTRL2 PAND2X1_484/CTRL
+ PAND2X1_484/a_76_28# PAND2X1
XPAND2X1_270 VDD GND POR2X1_39/B POR2X1_20/B POR2X1_271/A PAND2X1_270/a_16_344# PAND2X1_270/m4_208_n4#
+ PAND2X1_270/O PAND2X1_270/a_56_28# PAND2X1_270/CTRL2 PAND2X1_270/CTRL PAND2X1_270/a_76_28#
+ PAND2X1
XPAND2X1_281 VDD GND POR2X1_383/A POR2X1_66/B POR2X1_285/B PAND2X1_281/a_16_344# PAND2X1_281/m4_208_n4#
+ PAND2X1_281/O PAND2X1_281/a_56_28# PAND2X1_281/CTRL2 PAND2X1_281/CTRL PAND2X1_281/a_76_28#
+ PAND2X1
XPAND2X1_292 VDD GND POR2X1_186/B PAND2X1_41/B POR2X1_346/B PAND2X1_292/a_16_344#
+ PAND2X1_292/m4_208_n4# PAND2X1_292/O PAND2X1_292/a_56_28# PAND2X1_292/CTRL2 PAND2X1_292/CTRL
+ PAND2X1_292/a_76_28# PAND2X1
XPOR2X1_509 VDD GND POR2X1_509/B POR2X1_509/A POR2X1_510/A POR2X1_509/m4_208_n4# POR2X1_509/O
+ POR2X1_509/CTRL2 POR2X1_509/a_16_28# POR2X1_509/CTRL POR2X1_509/a_76_344# POR2X1_509/a_56_344#
+ POR2X1
XPOR2X1_317 VDD GND POR2X1_317/B POR2X1_317/A POR2X1_317/Y POR2X1_317/m4_208_n4# POR2X1_317/O
+ POR2X1_317/CTRL2 POR2X1_317/a_16_28# POR2X1_317/CTRL POR2X1_317/a_76_344# POR2X1_317/a_56_344#
+ POR2X1
XPOR2X1_306 VDD GND POR2X1_43/B POR2X1_376/B POR2X1_306/Y POR2X1_306/m4_208_n4# POR2X1_306/O
+ POR2X1_306/CTRL2 POR2X1_306/a_16_28# POR2X1_306/CTRL POR2X1_306/a_76_344# POR2X1_306/a_56_344#
+ POR2X1
XPOR2X1_339 VDD GND POR2X1_61/Y POR2X1_332/Y POR2X1_339/Y POR2X1_339/m4_208_n4# POR2X1_339/O
+ POR2X1_339/CTRL2 POR2X1_339/a_16_28# POR2X1_339/CTRL POR2X1_339/a_76_344# POR2X1_339/a_56_344#
+ POR2X1
XPOR2X1_328 VDD GND INPUT_4 POR2X1_51/A POR2X1_329/A POR2X1_328/m4_208_n4# POR2X1_328/O
+ POR2X1_328/CTRL2 POR2X1_328/a_16_28# POR2X1_328/CTRL POR2X1_328/a_76_344# POR2X1_328/a_56_344#
+ POR2X1
XPOR2X1_840 VDD GND POR2X1_840/B POR2X1_834/Y POR2X1_840/Y POR2X1_840/m4_208_n4# POR2X1_840/O
+ POR2X1_840/CTRL2 POR2X1_840/a_16_28# POR2X1_840/CTRL POR2X1_840/a_76_344# POR2X1_840/a_56_344#
+ POR2X1
XPOR2X1_851 VDD GND POR2X1_840/Y POR2X1_851/A POR2X1_858/A POR2X1_851/m4_208_n4# POR2X1_851/O
+ POR2X1_851/CTRL2 POR2X1_851/a_16_28# POR2X1_851/CTRL POR2X1_851/a_76_344# POR2X1_851/a_56_344#
+ POR2X1
XPOR2X1_862 VDD GND POR2X1_862/B POR2X1_862/A POR2X1_862/Y POR2X1_862/m4_208_n4# POR2X1_862/O
+ POR2X1_862/CTRL2 POR2X1_862/a_16_28# POR2X1_862/CTRL POR2X1_862/a_76_344# POR2X1_862/a_56_344#
+ POR2X1
XPAND2X1_814 VDD GND POR2X1_283/A POR2X1_411/B POR2X1_815/A PAND2X1_814/a_16_344#
+ PAND2X1_814/m4_208_n4# PAND2X1_814/O PAND2X1_814/a_56_28# PAND2X1_814/CTRL2 PAND2X1_814/CTRL
+ PAND2X1_814/a_76_28# PAND2X1
XPAND2X1_803 VDD GND PAND2X1_797/Y PAND2X1_803/A PAND2X1_803/Y PAND2X1_803/a_16_344#
+ PAND2X1_803/m4_208_n4# PAND2X1_803/O PAND2X1_803/a_56_28# PAND2X1_803/CTRL2 PAND2X1_803/CTRL
+ PAND2X1_803/a_76_28# PAND2X1
XPAND2X1_847 VDD GND POR2X1_820/Y POR2X1_817/Y PAND2X1_848/B PAND2X1_847/a_16_344#
+ PAND2X1_847/m4_208_n4# PAND2X1_847/O PAND2X1_847/a_56_28# PAND2X1_847/CTRL2 PAND2X1_847/CTRL
+ PAND2X1_847/a_76_28# PAND2X1
XPAND2X1_836 VDD GND POR2X1_824/Y POR2X1_823/Y PAND2X1_839/B PAND2X1_836/a_16_344#
+ PAND2X1_836/m4_208_n4# PAND2X1_836/O PAND2X1_836/a_56_28# PAND2X1_836/CTRL2 PAND2X1_836/CTRL
+ PAND2X1_836/a_76_28# PAND2X1
XPAND2X1_825 VDD GND PAND2X1_94/Y PAND2X1_57/B POR2X1_837/B PAND2X1_825/a_16_344#
+ PAND2X1_825/m4_208_n4# PAND2X1_825/O PAND2X1_825/a_56_28# PAND2X1_825/CTRL2 PAND2X1_825/CTRL
+ PAND2X1_825/a_76_28# PAND2X1
XPAND2X1_858 VDD GND PAND2X1_858/B PAND2X1_850/Y PAND2X1_858/Y PAND2X1_858/a_16_344#
+ PAND2X1_858/m4_208_n4# PAND2X1_858/O PAND2X1_858/a_56_28# PAND2X1_858/CTRL2 PAND2X1_858/CTRL
+ PAND2X1_858/a_76_28# PAND2X1
XPOR2X1_114 VDD GND POR2X1_114/B POR2X1_113/Y POR2X1_114/Y POR2X1_114/m4_208_n4# POR2X1_114/O
+ POR2X1_114/CTRL2 POR2X1_114/a_16_28# POR2X1_114/CTRL POR2X1_114/a_76_344# POR2X1_114/a_56_344#
+ POR2X1
XPOR2X1_125 VDD GND POR2X1_96/A POR2X1_411/B POR2X1_125/Y POR2X1_125/m4_208_n4# POR2X1_125/O
+ POR2X1_125/CTRL2 POR2X1_125/a_16_28# POR2X1_125/CTRL POR2X1_125/a_76_344# POR2X1_125/a_56_344#
+ POR2X1
XPOR2X1_103 VDD GND POR2X1_48/A POR2X1_102/Y POR2X1_103/Y POR2X1_103/m4_208_n4# POR2X1_103/O
+ POR2X1_103/CTRL2 POR2X1_103/a_16_28# POR2X1_103/CTRL POR2X1_103/a_76_344# POR2X1_103/a_56_344#
+ POR2X1
XPOR2X1_158 VDD GND POR2X1_158/B POR2X1_416/B POR2X1_158/Y POR2X1_158/m4_208_n4# POR2X1_158/O
+ POR2X1_158/CTRL2 POR2X1_158/a_16_28# POR2X1_158/CTRL POR2X1_158/a_76_344# POR2X1_158/a_56_344#
+ POR2X1
XPOR2X1_147 VDD GND POR2X1_830/A POR2X1_147/A POR2X1_149/B POR2X1_147/m4_208_n4# POR2X1_147/O
+ POR2X1_147/CTRL2 POR2X1_147/a_16_28# POR2X1_147/CTRL POR2X1_147/a_76_344# POR2X1_147/a_56_344#
+ POR2X1
XPOR2X1_136 VDD GND POR2X1_7/B POR2X1_42/Y POR2X1_136/Y POR2X1_136/m4_208_n4# POR2X1_136/O
+ POR2X1_136/CTRL2 POR2X1_136/a_16_28# POR2X1_136/CTRL POR2X1_136/a_76_344# POR2X1_136/a_56_344#
+ POR2X1
XPOR2X1_169 VDD GND POR2X1_169/B POR2X1_169/A POR2X1_169/Y POR2X1_169/m4_208_n4# POR2X1_169/O
+ POR2X1_169/CTRL2 POR2X1_169/a_16_28# POR2X1_169/CTRL POR2X1_169/a_76_344# POR2X1_169/a_56_344#
+ POR2X1
XPOR2X1_10 VDD GND POR2X1_8/Y POR2X1_9/Y POR2X1_41/B POR2X1_10/m4_208_n4# POR2X1_10/O
+ POR2X1_10/CTRL2 POR2X1_10/a_16_28# POR2X1_10/CTRL POR2X1_10/a_76_344# POR2X1_10/a_56_344#
+ POR2X1
XPAND2X1_90 VDD GND POR2X1_94/A PAND2X1_90/A PAND2X1_90/Y PAND2X1_90/a_16_344# PAND2X1_90/m4_208_n4#
+ PAND2X1_90/O PAND2X1_90/a_56_28# PAND2X1_90/CTRL2 PAND2X1_90/CTRL PAND2X1_90/a_76_28#
+ PAND2X1
XPOR2X1_43 VDD GND POR2X1_43/B POR2X1_42/Y POR2X1_43/Y POR2X1_43/m4_208_n4# POR2X1_43/O
+ POR2X1_43/CTRL2 POR2X1_43/a_16_28# POR2X1_43/CTRL POR2X1_43/a_76_344# POR2X1_43/a_56_344#
+ POR2X1
XPOR2X1_32 VDD GND POR2X1_29/Y POR2X1_32/A POR2X1_32/Y POR2X1_32/m4_208_n4# POR2X1_32/O
+ POR2X1_32/CTRL2 POR2X1_32/a_16_28# POR2X1_32/CTRL POR2X1_32/a_76_344# POR2X1_32/a_56_344#
+ POR2X1
XPOR2X1_21 VDD GND D_INPUT_4 INPUT_5 POR2X1_22/A POR2X1_21/m4_208_n4# POR2X1_21/O
+ POR2X1_21/CTRL2 POR2X1_21/a_16_28# POR2X1_21/CTRL POR2X1_21/a_76_344# POR2X1_21/a_56_344#
+ POR2X1
XPOR2X1_54 VDD GND D_INPUT_0 D_INPUT_1 POR2X1_54/Y POR2X1_54/m4_208_n4# POR2X1_54/O
+ POR2X1_54/CTRL2 POR2X1_54/a_16_28# POR2X1_54/CTRL POR2X1_54/a_76_344# POR2X1_54/a_56_344#
+ POR2X1
XPOR2X1_87 VDD GND POR2X1_87/B POR2X1_68/A POR2X1_87/Y POR2X1_87/m4_208_n4# POR2X1_87/O
+ POR2X1_87/CTRL2 POR2X1_87/a_16_28# POR2X1_87/CTRL POR2X1_87/a_76_344# POR2X1_87/a_56_344#
+ POR2X1
XPOR2X1_65 VDD GND POR2X1_63/Y POR2X1_65/A POR2X1_65/Y POR2X1_65/m4_208_n4# POR2X1_65/O
+ POR2X1_65/CTRL2 POR2X1_65/a_16_28# POR2X1_65/CTRL POR2X1_65/a_76_344# POR2X1_65/a_56_344#
+ POR2X1
XPOR2X1_76 VDD GND POR2X1_76/B POR2X1_76/A POR2X1_76/Y POR2X1_76/m4_208_n4# POR2X1_76/O
+ POR2X1_76/CTRL2 POR2X1_76/a_16_28# POR2X1_76/CTRL POR2X1_76/a_76_344# POR2X1_76/a_56_344#
+ POR2X1
XPOR2X1_98 VDD GND POR2X1_98/B POR2X1_98/A POR2X1_99/A POR2X1_98/m4_208_n4# POR2X1_98/O
+ POR2X1_98/CTRL2 POR2X1_98/a_16_28# POR2X1_98/CTRL POR2X1_98/a_76_344# POR2X1_98/a_56_344#
+ POR2X1
XPOR2X1_670 VDD GND POR2X1_40/Y POR2X1_102/Y POR2X1_670/Y POR2X1_670/m4_208_n4# POR2X1_670/O
+ POR2X1_670/CTRL2 POR2X1_670/a_16_28# POR2X1_670/CTRL POR2X1_670/a_76_344# POR2X1_670/a_56_344#
+ POR2X1
XPOR2X1_681 VDD GND POR2X1_32/A POR2X1_153/Y POR2X1_681/Y POR2X1_681/m4_208_n4# POR2X1_681/O
+ POR2X1_681/CTRL2 POR2X1_681/a_16_28# POR2X1_681/CTRL POR2X1_681/a_76_344# POR2X1_681/a_56_344#
+ POR2X1
XPOR2X1_692 VDD GND POR2X1_20/B POR2X1_46/Y POR2X1_692/Y POR2X1_692/m4_208_n4# POR2X1_692/O
+ POR2X1_692/CTRL2 POR2X1_692/a_16_28# POR2X1_692/CTRL POR2X1_692/a_76_344# POR2X1_692/a_56_344#
+ POR2X1
XPAND2X1_622 VDD GND PAND2X1_621/Y POR2X1_619/Y PAND2X1_624/A PAND2X1_622/a_16_344#
+ PAND2X1_622/m4_208_n4# PAND2X1_622/O PAND2X1_622/a_56_28# PAND2X1_622/CTRL2 PAND2X1_622/CTRL
+ PAND2X1_622/a_76_28# PAND2X1
XPAND2X1_611 VDD GND POR2X1_54/Y POR2X1_68/B PAND2X1_612/B PAND2X1_611/a_16_344# PAND2X1_611/m4_208_n4#
+ PAND2X1_611/O PAND2X1_611/a_56_28# PAND2X1_611/CTRL2 PAND2X1_611/CTRL PAND2X1_611/a_76_28#
+ PAND2X1
XPAND2X1_600 VDD GND POR2X1_814/B PAND2X1_32/B POR2X1_602/B PAND2X1_600/a_16_344#
+ POR2X1_719/m4_208_n4# PAND2X1_600/O PAND2X1_600/a_56_28# PAND2X1_600/CTRL2 PAND2X1_600/CTRL
+ PAND2X1_600/a_76_28# PAND2X1
XPAND2X1_633 VDD GND POR2X1_278/A POR2X1_118/Y PAND2X1_633/Y PAND2X1_633/a_16_344#
+ PAND2X1_633/m4_208_n4# PAND2X1_633/O PAND2X1_633/a_56_28# PAND2X1_633/CTRL2 PAND2X1_633/CTRL
+ PAND2X1_633/a_76_28# PAND2X1
XPAND2X1_644 VDD GND POR2X1_761/A POR2X1_597/Y PAND2X1_644/Y PAND2X1_644/a_16_344#
+ PAND2X1_644/m4_208_n4# PAND2X1_644/O PAND2X1_644/a_56_28# PAND2X1_644/CTRL2 PAND2X1_644/CTRL
+ PAND2X1_644/a_76_28# PAND2X1
XPAND2X1_655 VDD GND PAND2X1_655/B PAND2X1_648/Y PAND2X1_655/Y PAND2X1_655/a_16_344#
+ PAND2X1_655/m4_208_n4# PAND2X1_655/O PAND2X1_655/a_56_28# PAND2X1_655/CTRL2 PAND2X1_655/CTRL
+ PAND2X1_655/a_76_28# PAND2X1
XPAND2X1_666 VDD GND POR2X1_121/A PAND2X1_20/A POR2X1_719/A PAND2X1_666/a_16_344#
+ PAND2X1_666/m4_208_n4# PAND2X1_666/O PAND2X1_666/a_56_28# PAND2X1_666/CTRL2 PAND2X1_666/CTRL
+ PAND2X1_666/a_76_28# PAND2X1
XPAND2X1_677 VDD GND POR2X1_614/A POR2X1_66/A POR2X1_678/A PAND2X1_677/a_16_344# PAND2X1_677/m4_208_n4#
+ PAND2X1_677/O PAND2X1_677/a_56_28# PAND2X1_677/CTRL2 PAND2X1_677/CTRL PAND2X1_677/a_76_28#
+ PAND2X1
XPAND2X1_688 VDD GND POR2X1_293/Y POR2X1_38/Y POR2X1_689/A PAND2X1_688/a_16_344# PAND2X1_688/m4_208_n4#
+ PAND2X1_688/O PAND2X1_688/a_56_28# PAND2X1_688/CTRL2 PAND2X1_688/CTRL PAND2X1_688/a_76_28#
+ PAND2X1
XPAND2X1_699 VDD GND POR2X1_260/A PAND2X1_94/A POR2X1_709/A PAND2X1_699/a_16_344#
+ PAND2X1_699/m4_208_n4# PAND2X1_699/O PAND2X1_699/a_56_28# PAND2X1_699/CTRL2 PAND2X1_699/CTRL
+ PAND2X1_699/a_76_28# PAND2X1
XPAND2X1_9 VDD GND D_INPUT_1 D_INPUT_0 PAND2X1_9/Y PAND2X1_9/a_16_344# PAND2X1_9/m4_208_n4#
+ PAND2X1_9/O PAND2X1_9/a_56_28# PAND2X1_9/CTRL2 PAND2X1_9/CTRL PAND2X1_9/a_76_28#
+ PAND2X1
XPAND2X1_430 VDD GND PAND2X1_429/Y POR2X1_750/B POR2X1_451/A PAND2X1_430/a_16_344#
+ PAND2X1_430/m4_208_n4# PAND2X1_430/O PAND2X1_430/a_56_28# PAND2X1_430/CTRL2 PAND2X1_430/CTRL
+ PAND2X1_430/a_76_28# PAND2X1
XPAND2X1_441 VDD GND POR2X1_68/A PAND2X1_41/B POR2X1_443/A PAND2X1_441/a_16_344# PAND2X1_441/m4_208_n4#
+ PAND2X1_441/O PAND2X1_441/a_56_28# PAND2X1_441/CTRL2 PAND2X1_441/CTRL PAND2X1_441/a_76_28#
+ PAND2X1
XPAND2X1_452 VDD GND PAND2X1_452/B PAND2X1_452/A PAND2X1_467/B PAND2X1_452/a_16_344#
+ PAND2X1_452/m4_208_n4# PAND2X1_452/O PAND2X1_452/a_56_28# PAND2X1_452/CTRL2 PAND2X1_452/CTRL
+ PAND2X1_452/a_76_28# PAND2X1
XPAND2X1_463 VDD GND PAND2X1_460/Y PAND2X1_459/Y PAND2X1_472/B PAND2X1_463/a_16_344#
+ PAND2X1_463/m4_208_n4# PAND2X1_463/O PAND2X1_463/a_56_28# PAND2X1_463/CTRL2 PAND2X1_463/CTRL
+ PAND2X1_463/a_76_28# PAND2X1
XPAND2X1_496 VDD GND PAND2X1_55/Y PAND2X1_20/A POR2X1_499/A PAND2X1_496/a_16_344#
+ PAND2X1_496/m4_208_n4# PAND2X1_496/O PAND2X1_496/a_56_28# PAND2X1_496/CTRL2 PAND2X1_496/CTRL
+ PAND2X1_496/a_76_28# PAND2X1
XPAND2X1_474 VDD GND PAND2X1_404/Y PAND2X1_474/A PAND2X1_474/Y PAND2X1_474/a_16_344#
+ PAND2X1_97/m4_208_n4# PAND2X1_474/O PAND2X1_474/a_56_28# PAND2X1_474/CTRL2 PAND2X1_474/CTRL
+ PAND2X1_474/a_76_28# PAND2X1
XPAND2X1_485 VDD GND POR2X1_590/A PAND2X1_57/B POR2X1_705/B PAND2X1_485/a_16_344#
+ PAND2X1_485/m4_208_n4# PAND2X1_485/O PAND2X1_485/a_56_28# PAND2X1_485/CTRL2 PAND2X1_485/CTRL
+ PAND2X1_485/a_76_28# PAND2X1
XPAND2X1_271 VDD GND POR2X1_270/Y POR2X1_269/Y POR2X1_276/B PAND2X1_271/a_16_344#
+ PAND2X1_271/m4_208_n4# PAND2X1_271/O PAND2X1_271/a_56_28# PAND2X1_271/CTRL2 PAND2X1_271/CTRL
+ PAND2X1_271/a_76_28# PAND2X1
XPAND2X1_282 VDD GND POR2X1_260/A POR2X1_590/A POR2X1_285/A PAND2X1_282/a_16_344#
+ PAND2X1_282/m4_208_n4# PAND2X1_282/O PAND2X1_282/a_56_28# PAND2X1_282/CTRL2 PAND2X1_282/CTRL
+ PAND2X1_282/a_76_28# PAND2X1
XPAND2X1_260 VDD GND POR2X1_416/B POR2X1_13/A POR2X1_261/A PAND2X1_260/a_16_344# PAND2X1_260/m4_208_n4#
+ PAND2X1_260/O PAND2X1_260/a_56_28# PAND2X1_260/CTRL2 PAND2X1_260/CTRL PAND2X1_260/a_76_28#
+ PAND2X1
XPAND2X1_293 VDD GND POR2X1_68/B INPUT_1 POR2X1_294/A PAND2X1_293/a_16_344# PAND2X1_293/m4_208_n4#
+ PAND2X1_293/O PAND2X1_293/a_56_28# PAND2X1_293/CTRL2 PAND2X1_293/CTRL PAND2X1_293/a_76_28#
+ PAND2X1
XPOR2X1_307 VDD GND POR2X1_307/B POR2X1_307/A POR2X1_307/Y POR2X1_307/m4_208_n4# POR2X1_307/O
+ POR2X1_307/CTRL2 POR2X1_307/a_16_28# POR2X1_307/CTRL POR2X1_307/a_76_344# POR2X1_307/a_56_344#
+ POR2X1
XPOR2X1_329 VDD GND POR2X1_760/A POR2X1_329/A POR2X1_329/Y POR2X1_329/m4_208_n4# POR2X1_329/O
+ POR2X1_329/CTRL2 POR2X1_329/a_16_28# POR2X1_329/CTRL POR2X1_329/a_76_344# POR2X1_329/a_56_344#
+ POR2X1
XPOR2X1_318 VDD GND POR2X1_445/A POR2X1_318/A POR2X1_319/A POR2X1_318/m4_208_n4# POR2X1_318/O
+ POR2X1_318/CTRL2 POR2X1_318/a_16_28# POR2X1_318/CTRL POR2X1_318/a_76_344# POR2X1_318/a_56_344#
+ POR2X1
XPOR2X1_830 VDD GND POR2X1_114/B POR2X1_830/A POR2X1_830/Y POR2X1_830/m4_208_n4# POR2X1_830/O
+ POR2X1_830/CTRL2 POR2X1_830/a_16_28# POR2X1_830/CTRL POR2X1_830/a_76_344# POR2X1_830/a_56_344#
+ POR2X1
XPOR2X1_852 VDD GND POR2X1_852/B POR2X1_852/A POR2X1_857/B POR2X1_852/m4_208_n4# POR2X1_852/O
+ POR2X1_852/CTRL2 POR2X1_852/a_16_28# POR2X1_852/CTRL POR2X1_852/a_76_344# POR2X1_852/a_56_344#
+ POR2X1
XPOR2X1_863 VDD GND POR2X1_863/B POR2X1_863/A POR2X1_864/A POR2X1_863/m4_208_n4# POR2X1_863/O
+ POR2X1_863/CTRL2 POR2X1_863/a_16_28# POR2X1_863/CTRL POR2X1_863/a_76_344# POR2X1_863/a_56_344#
+ POR2X1
XPOR2X1_841 VDD GND POR2X1_841/B POR2X1_832/Y POR2X1_851/A POR2X1_841/m4_208_n4# POR2X1_841/O
+ POR2X1_841/CTRL2 POR2X1_841/a_16_28# POR2X1_841/CTRL POR2X1_841/a_76_344# POR2X1_841/a_56_344#
+ POR2X1
XPAND2X1_804 VDD GND PAND2X1_804/B PAND2X1_804/A PAND2X1_808/B PAND2X1_804/a_16_344#
+ PAND2X1_804/m4_208_n4# PAND2X1_804/O PAND2X1_804/a_56_28# PAND2X1_804/CTRL2 PAND2X1_804/CTRL
+ PAND2X1_804/a_76_28# PAND2X1
XPAND2X1_815 VDD GND POR2X1_814/Y POR2X1_66/B POR2X1_846/B PAND2X1_815/a_16_344# PAND2X1_815/m4_208_n4#
+ PAND2X1_815/O PAND2X1_815/a_56_28# PAND2X1_815/CTRL2 PAND2X1_815/CTRL PAND2X1_815/a_76_28#
+ PAND2X1
XPAND2X1_837 VDD GND POR2X1_826/Y POR2X1_825/Y PAND2X1_838/B PAND2X1_837/a_16_344#
+ PAND2X1_837/m4_208_n4# PAND2X1_837/O PAND2X1_837/a_56_28# PAND2X1_837/CTRL2 PAND2X1_837/CTRL
+ PAND2X1_837/a_76_28# PAND2X1
XPAND2X1_826 VDD GND PAND2X1_96/B PAND2X1_55/Y POR2X1_837/A PAND2X1_826/a_16_344#
+ PAND2X1_826/m4_208_n4# PAND2X1_826/O PAND2X1_826/a_56_28# PAND2X1_826/CTRL2 PAND2X1_826/CTRL
+ PAND2X1_826/a_76_28# PAND2X1
XPAND2X1_848 VDD GND PAND2X1_848/B PAND2X1_848/A PAND2X1_859/A PAND2X1_848/a_16_344#
+ PAND2X1_848/m4_208_n4# PAND2X1_848/O PAND2X1_848/a_56_28# PAND2X1_848/CTRL2 PAND2X1_848/CTRL
+ PAND2X1_848/a_76_28# PAND2X1
XPAND2X1_859 VDD GND PAND2X1_859/B PAND2X1_859/A PAND2X1_862/B PAND2X1_859/a_16_344#
+ PAND2X1_859/m4_208_n4# PAND2X1_859/O PAND2X1_859/a_56_28# PAND2X1_859/CTRL2 PAND2X1_859/CTRL
+ PAND2X1_859/a_76_28# PAND2X1
XPOR2X1_104 VDD GND POR2X1_4/Y POR2X1_8/Y POR2X1_411/B POR2X1_104/m4_208_n4# POR2X1_104/O
+ POR2X1_104/CTRL2 POR2X1_104/a_16_28# POR2X1_104/CTRL POR2X1_104/a_76_344# POR2X1_104/a_56_344#
+ POR2X1
XPOR2X1_115 VDD GND POR2X1_554/B POR2X1_112/Y POR2X1_116/A POR2X1_115/m4_208_n4# POR2X1_115/O
+ POR2X1_115/CTRL2 POR2X1_115/a_16_28# POR2X1_115/CTRL POR2X1_115/a_76_344# POR2X1_115/a_56_344#
+ POR2X1
XPOR2X1_126 VDD GND POR2X1_4/Y POR2X1_37/Y POR2X1_394/A POR2X1_126/m4_208_n4# POR2X1_126/O
+ POR2X1_126/CTRL2 POR2X1_126/a_16_28# POR2X1_126/CTRL POR2X1_126/a_76_344# POR2X1_126/a_56_344#
+ POR2X1
XPOR2X1_159 VDD GND POR2X1_5/Y POR2X1_9/Y POR2X1_669/B POR2X1_159/m4_208_n4# POR2X1_159/O
+ POR2X1_159/CTRL2 POR2X1_159/a_16_28# POR2X1_159/CTRL POR2X1_159/a_76_344# POR2X1_159/a_56_344#
+ POR2X1
XPOR2X1_137 VDD GND POR2X1_137/B POR2X1_768/A POR2X1_137/Y POR2X1_113/m4_208_n4# POR2X1_137/O
+ POR2X1_137/CTRL2 POR2X1_137/a_16_28# POR2X1_137/CTRL POR2X1_137/a_76_344# POR2X1_137/a_56_344#
+ POR2X1
XPOR2X1_148 VDD GND POR2X1_148/B POR2X1_148/A POR2X1_149/A POR2X1_148/m4_208_n4# POR2X1_148/O
+ POR2X1_148/CTRL2 POR2X1_148/a_16_28# POR2X1_148/CTRL POR2X1_148/a_76_344# POR2X1_148/a_56_344#
+ POR2X1
XPAND2X1_80 VDD GND POR2X1_38/B POR2X1_68/B PAND2X1_81/B PAND2X1_80/a_16_344# PAND2X1_80/m4_208_n4#
+ PAND2X1_80/O PAND2X1_80/a_56_28# PAND2X1_80/CTRL2 PAND2X1_80/CTRL PAND2X1_80/a_76_28#
+ PAND2X1
XPOR2X1_11 VDD GND INPUT_4 D_INPUT_5 POR2X1_12/A POR2X1_11/m4_208_n4# POR2X1_11/O
+ POR2X1_11/CTRL2 POR2X1_11/a_16_28# POR2X1_11/CTRL POR2X1_11/a_76_344# POR2X1_11/a_56_344#
+ POR2X1
XPAND2X1_91 VDD GND PAND2X1_90/Y PAND2X1_52/B POR2X1_97/A PAND2X1_91/a_16_344# PAND2X1_91/m4_208_n4#
+ PAND2X1_91/O PAND2X1_91/a_56_28# PAND2X1_91/CTRL2 PAND2X1_91/CTRL PAND2X1_91/a_76_28#
+ PAND2X1
XPOR2X1_33 VDD GND POR2X1_33/B POR2X1_33/A POR2X1_35/B POR2X1_33/m4_208_n4# POR2X1_33/O
+ POR2X1_33/CTRL2 POR2X1_33/a_16_28# POR2X1_33/CTRL POR2X1_33/a_76_344# POR2X1_33/a_56_344#
+ POR2X1
XPOR2X1_44 VDD GND POR2X1_36/B POR2X1_51/B POR2X1_57/A POR2X1_44/m4_208_n4# POR2X1_44/O
+ POR2X1_44/CTRL2 POR2X1_44/a_16_28# POR2X1_44/CTRL POR2X1_44/a_76_344# POR2X1_44/a_56_344#
+ POR2X1
XPOR2X1_22 VDD GND POR2X1_3/B POR2X1_22/A POR2X1_43/B POR2X1_22/m4_208_n4# POR2X1_22/O
+ POR2X1_22/CTRL2 POR2X1_22/a_16_28# POR2X1_22/CTRL POR2X1_22/a_76_344# POR2X1_22/a_56_344#
+ POR2X1
XPOR2X1_66 VDD GND POR2X1_66/B POR2X1_66/A POR2X1_66/Y POR2X1_66/m4_208_n4# POR2X1_66/O
+ POR2X1_66/CTRL2 POR2X1_66/a_16_28# POR2X1_66/CTRL POR2X1_66/a_76_344# POR2X1_66/a_56_344#
+ POR2X1
XPOR2X1_77 VDD GND POR2X1_14/Y POR2X1_54/Y POR2X1_77/Y POR2X1_77/m4_208_n4# POR2X1_77/O
+ POR2X1_77/CTRL2 POR2X1_77/a_16_28# POR2X1_77/CTRL POR2X1_77/a_76_344# POR2X1_77/a_56_344#
+ POR2X1
XPOR2X1_55 VDD GND POR2X1_5/Y POR2X1_54/Y POR2X1_55/Y POR2X1_55/m4_208_n4# POR2X1_55/O
+ POR2X1_55/CTRL2 POR2X1_55/a_16_28# POR2X1_55/CTRL POR2X1_55/a_76_344# POR2X1_55/a_56_344#
+ POR2X1
XPOR2X1_671 VDD GND D_INPUT_2 POR2X1_4/Y POR2X1_672/A POR2X1_671/m4_208_n4# POR2X1_671/O
+ POR2X1_671/CTRL2 POR2X1_671/a_16_28# POR2X1_671/CTRL POR2X1_671/a_76_344# POR2X1_671/a_56_344#
+ POR2X1
XPOR2X1_99 VDD GND POR2X1_99/B POR2X1_99/A POR2X1_99/Y POR2X1_99/m4_208_n4# POR2X1_99/O
+ POR2X1_99/CTRL2 POR2X1_99/a_16_28# POR2X1_99/CTRL POR2X1_99/a_76_344# POR2X1_99/a_56_344#
+ POR2X1
XPOR2X1_88 VDD GND POR2X1_7/B POR2X1_88/A POR2X1_88/Y POR2X1_88/m4_208_n4# POR2X1_88/O
+ POR2X1_88/CTRL2 POR2X1_88/a_16_28# POR2X1_88/CTRL POR2X1_88/a_76_344# POR2X1_88/a_56_344#
+ POR2X1
XPOR2X1_660 VDD GND POR2X1_655/Y POR2X1_660/A POR2X1_660/Y POR2X1_660/m4_208_n4# POR2X1_660/O
+ POR2X1_660/CTRL2 POR2X1_660/a_16_28# POR2X1_660/CTRL POR2X1_660/a_76_344# POR2X1_660/a_56_344#
+ POR2X1
XPOR2X1_682 VDD GND POR2X1_39/B POR2X1_669/B POR2X1_682/Y POR2X1_682/m4_208_n4# POR2X1_682/O
+ POR2X1_682/CTRL2 POR2X1_682/a_16_28# POR2X1_682/CTRL POR2X1_682/a_76_344# POR2X1_682/a_56_344#
+ POR2X1
XPOR2X1_693 VDD GND POR2X1_14/Y POR2X1_39/B POR2X1_693/Y POR2X1_693/m4_208_n4# POR2X1_693/O
+ POR2X1_693/CTRL2 POR2X1_693/a_16_28# POR2X1_693/CTRL POR2X1_693/a_76_344# POR2X1_693/a_56_344#
+ POR2X1
XPAND2X1_612 VDD GND PAND2X1_612/B POR2X1_610/Y POR2X1_647/B PAND2X1_612/a_16_344#
+ PAND2X1_612/m4_208_n4# PAND2X1_612/O PAND2X1_612/a_56_28# PAND2X1_612/CTRL2 PAND2X1_612/CTRL
+ PAND2X1_612/a_76_28# PAND2X1
XPAND2X1_601 VDD GND PAND2X1_48/B POR2X1_78/B POR2X1_602/A PAND2X1_601/a_16_344# PAND2X1_601/m4_208_n4#
+ PAND2X1_601/O PAND2X1_601/a_56_28# PAND2X1_601/CTRL2 PAND2X1_601/CTRL PAND2X1_601/a_76_28#
+ PAND2X1
XPAND2X1_623 VDD GND PAND2X1_620/Y POR2X1_615/Y PAND2X1_623/Y PAND2X1_623/a_16_344#
+ PAND2X1_623/m4_208_n4# PAND2X1_623/O PAND2X1_623/a_56_28# PAND2X1_623/CTRL2 PAND2X1_623/CTRL
+ PAND2X1_623/a_76_28# PAND2X1
XPAND2X1_645 VDD GND PAND2X1_645/B PAND2X1_602/Y PAND2X1_645/Y PAND2X1_645/a_16_344#
+ PAND2X1_645/m4_208_n4# PAND2X1_645/O PAND2X1_645/a_56_28# PAND2X1_645/CTRL2 PAND2X1_645/CTRL
+ PAND2X1_645/a_76_28# PAND2X1
XPAND2X1_634 VDD GND POR2X1_413/A POR2X1_290/Y PAND2X1_640/B PAND2X1_634/a_16_344#
+ PAND2X1_634/m4_208_n4# PAND2X1_634/O PAND2X1_634/a_56_28# PAND2X1_634/CTRL2 PAND2X1_634/CTRL
+ PAND2X1_634/a_76_28# PAND2X1
XPAND2X1_656 VDD GND PAND2X1_656/B PAND2X1_656/A PAND2X1_660/B PAND2X1_656/a_16_344#
+ POR2X1_394/m4_208_n4# PAND2X1_656/O PAND2X1_656/a_56_28# PAND2X1_656/CTRL2 PAND2X1_656/CTRL
+ PAND2X1_656/a_76_28# PAND2X1
XPAND2X1_667 VDD GND POR2X1_264/Y PAND2X1_65/B POR2X1_720/B PAND2X1_667/a_16_344#
+ PAND2X1_667/m4_208_n4# PAND2X1_667/O PAND2X1_667/a_56_28# PAND2X1_667/CTRL2 PAND2X1_667/CTRL
+ PAND2X1_667/a_76_28# PAND2X1
XPAND2X1_678 VDD GND POR2X1_677/Y POR2X1_13/A POR2X1_679/A PAND2X1_678/a_16_344# PAND2X1_678/m4_208_n4#
+ PAND2X1_678/O PAND2X1_678/a_56_28# PAND2X1_678/CTRL2 PAND2X1_678/CTRL PAND2X1_678/a_76_28#
+ PAND2X1
XPAND2X1_689 VDD GND POR2X1_688/Y PAND2X1_32/B POR2X1_691/B PAND2X1_689/a_16_344#
+ PAND2X1_689/m4_208_n4# PAND2X1_689/O PAND2X1_689/a_56_28# PAND2X1_689/CTRL2 PAND2X1_689/CTRL
+ PAND2X1_689/a_76_28# PAND2X1
XPOR2X1_490 VDD GND PAND2X1_6/A POR2X1_85/Y POR2X1_490/Y POR2X1_490/m4_208_n4# POR2X1_490/O
+ POR2X1_490/CTRL2 POR2X1_490/a_16_28# POR2X1_490/CTRL POR2X1_490/a_76_344# POR2X1_490/a_56_344#
+ POR2X1
XPAND2X1_431 VDD GND POR2X1_383/A PAND2X1_72/A POR2X1_434/A PAND2X1_431/a_16_344#
+ PAND2X1_431/m4_208_n4# PAND2X1_431/O PAND2X1_431/a_56_28# PAND2X1_431/CTRL2 PAND2X1_431/CTRL
+ PAND2X1_431/a_76_28# PAND2X1
XPAND2X1_420 VDD GND POR2X1_590/A PAND2X1_96/B POR2X1_447/A PAND2X1_420/a_16_344#
+ PAND2X1_420/m4_208_n4# PAND2X1_420/O PAND2X1_420/a_56_28# PAND2X1_420/CTRL2 PAND2X1_420/CTRL
+ PAND2X1_420/a_76_28# PAND2X1
XPAND2X1_442 VDD GND POR2X1_814/B PAND2X1_41/B POR2X1_444/B PAND2X1_442/a_16_344#
+ PAND2X1_442/m4_208_n4# PAND2X1_442/O PAND2X1_442/a_56_28# PAND2X1_442/CTRL2 PAND2X1_442/CTRL
+ PAND2X1_442/a_76_28# PAND2X1
XPAND2X1_453 VDD GND PAND2X1_449/Y PAND2X1_453/A PAND2X1_466/A PAND2X1_453/a_16_344#
+ PAND2X1_453/m4_208_n4# PAND2X1_453/O PAND2X1_453/a_56_28# PAND2X1_453/CTRL2 PAND2X1_453/CTRL
+ PAND2X1_453/a_76_28# PAND2X1
XPAND2X1_464 VDD GND PAND2X1_464/B PAND2X1_457/Y PAND2X1_464/Y PAND2X1_464/a_16_344#
+ PAND2X1_464/m4_208_n4# PAND2X1_464/O PAND2X1_464/a_56_28# PAND2X1_464/CTRL2 PAND2X1_464/CTRL
+ PAND2X1_464/a_76_28# PAND2X1
XPAND2X1_497 VDD GND PAND2X1_71/Y PAND2X1_58/A POR2X1_844/B PAND2X1_497/a_16_344#
+ PAND2X1_79/m4_208_n4# PAND2X1_497/O PAND2X1_497/a_56_28# PAND2X1_497/CTRL2 PAND2X1_497/CTRL
+ PAND2X1_497/a_76_28# PAND2X1
XPAND2X1_475 VDD GND PAND2X1_474/Y POR2X1_406/Y PAND2X1_479/A PAND2X1_475/a_16_344#
+ PAND2X1_475/m4_208_n4# PAND2X1_475/O PAND2X1_475/a_56_28# PAND2X1_475/CTRL2 PAND2X1_475/CTRL
+ PAND2X1_475/a_76_28# PAND2X1
XPAND2X1_486 VDD GND POR2X1_485/Y POR2X1_484/Y PAND2X1_556/B PAND2X1_486/a_16_344#
+ POR2X1_526/m4_208_n4# PAND2X1_486/O PAND2X1_486/a_56_28# PAND2X1_486/CTRL2 PAND2X1_486/CTRL
+ PAND2X1_486/a_76_28# PAND2X1
XPAND2X1_272 VDD GND POR2X1_296/B PAND2X1_32/B POR2X1_274/B PAND2X1_272/a_16_344#
+ PAND2X1_272/m4_208_n4# PAND2X1_272/O PAND2X1_272/a_56_28# PAND2X1_272/CTRL2 PAND2X1_272/CTRL
+ PAND2X1_272/a_76_28# PAND2X1
XPAND2X1_250 VDD GND POR2X1_249/Y PAND2X1_65/B POR2X1_343/B PAND2X1_250/a_16_344#
+ PAND2X1_250/m4_208_n4# PAND2X1_250/O PAND2X1_250/a_56_28# PAND2X1_250/CTRL2 PAND2X1_250/CTRL
+ PAND2X1_250/a_76_28# PAND2X1
XPAND2X1_261 VDD GND POR2X1_260/Y POR2X1_814/B POR2X1_345/A PAND2X1_261/a_16_344#
+ PAND2X1_261/m4_208_n4# PAND2X1_261/O PAND2X1_261/a_56_28# PAND2X1_261/CTRL2 PAND2X1_261/CTRL
+ PAND2X1_261/a_76_28# PAND2X1
XPAND2X1_283 VDD GND POR2X1_814/A POR2X1_66/A POR2X1_286/B PAND2X1_283/a_16_344# PAND2X1_283/m4_208_n4#
+ PAND2X1_283/O PAND2X1_283/a_56_28# PAND2X1_283/CTRL2 PAND2X1_283/CTRL PAND2X1_283/a_76_28#
+ PAND2X1
XPAND2X1_294 VDD GND POR2X1_293/Y POR2X1_41/B POR2X1_481/A PAND2X1_294/a_16_344# PAND2X1_337/m4_208_n4#
+ PAND2X1_294/O PAND2X1_294/a_56_28# PAND2X1_294/CTRL2 PAND2X1_294/CTRL PAND2X1_294/a_76_28#
+ PAND2X1
XPOR2X1_308 VDD GND POR2X1_308/B POR2X1_307/Y POR2X1_353/A POR2X1_308/m4_208_n4# POR2X1_308/O
+ POR2X1_308/CTRL2 POR2X1_308/a_16_28# POR2X1_308/CTRL POR2X1_308/a_76_344# POR2X1_308/a_56_344#
+ POR2X1
XPOR2X1_319 VDD GND POR2X1_317/Y POR2X1_319/A POR2X1_319/Y POR2X1_367/m4_208_n4# POR2X1_319/O
+ POR2X1_319/CTRL2 POR2X1_319/a_16_28# POR2X1_319/CTRL POR2X1_319/a_76_344# POR2X1_319/a_56_344#
+ POR2X1
XPOR2X1_820 VDD GND POR2X1_820/B POR2X1_820/A POR2X1_820/Y POR2X1_820/m4_208_n4# POR2X1_820/O
+ POR2X1_820/CTRL2 POR2X1_820/a_16_28# POR2X1_820/CTRL POR2X1_820/a_76_344# POR2X1_820/a_56_344#
+ POR2X1
XPOR2X1_853 VDD GND POR2X1_35/Y POR2X1_853/A POR2X1_857/A POR2X1_853/m4_208_n4# POR2X1_853/O
+ POR2X1_853/CTRL2 POR2X1_853/a_16_28# POR2X1_853/CTRL POR2X1_853/a_76_344# POR2X1_853/a_56_344#
+ POR2X1
XPOR2X1_831 VDD GND POR2X1_274/A POR2X1_301/A POR2X1_841/B POR2X1_831/m4_208_n4# POR2X1_831/O
+ POR2X1_831/CTRL2 POR2X1_831/a_16_28# POR2X1_831/CTRL POR2X1_831/a_76_344# POR2X1_831/a_56_344#
+ POR2X1
XPOR2X1_842 VDD GND POR2X1_456/B POR2X1_830/Y POR2X1_850/B POR2X1_842/m4_208_n4# POR2X1_842/O
+ POR2X1_842/CTRL2 POR2X1_842/a_16_28# POR2X1_842/CTRL POR2X1_842/a_76_344# POR2X1_842/a_56_344#
+ POR2X1
XPOR2X1_864 VDD GND POR2X1_774/Y POR2X1_864/A POR2X1_866/B POR2X1_864/m4_208_n4# POR2X1_864/O
+ POR2X1_864/CTRL2 POR2X1_864/a_16_28# POR2X1_864/CTRL POR2X1_864/a_76_344# POR2X1_864/a_56_344#
+ POR2X1
XPAND2X1_805 VDD GND PAND2X1_793/Y PAND2X1_805/A PAND2X1_805/Y PAND2X1_805/a_16_344#
+ PAND2X1_805/m4_208_n4# PAND2X1_805/O PAND2X1_805/a_56_28# PAND2X1_805/CTRL2 PAND2X1_805/CTRL
+ PAND2X1_805/a_76_28# PAND2X1
XPAND2X1_816 VDD GND POR2X1_188/A PAND2X1_52/B POR2X1_846/A PAND2X1_816/a_16_344#
+ PAND2X1_816/m4_208_n4# PAND2X1_816/O PAND2X1_816/a_56_28# PAND2X1_816/CTRL2 PAND2X1_816/CTRL
+ PAND2X1_816/a_76_28# PAND2X1
XPAND2X1_838 VDD GND PAND2X1_838/B POR2X1_827/Y PAND2X1_852/A PAND2X1_838/a_16_344#
+ PAND2X1_195/m4_208_n4# PAND2X1_838/O PAND2X1_838/a_56_28# PAND2X1_838/CTRL2 PAND2X1_838/CTRL
+ PAND2X1_838/a_76_28# PAND2X1
XPAND2X1_827 VDD GND POR2X1_260/A POR2X1_296/B POR2X1_838/B PAND2X1_827/a_16_344#
+ PAND2X1_827/m4_208_n4# PAND2X1_827/O PAND2X1_827/a_56_28# PAND2X1_827/CTRL2 PAND2X1_827/CTRL
+ PAND2X1_827/a_76_28# PAND2X1
XPAND2X1_849 VDD GND PAND2X1_849/B PAND2X1_844/Y PAND2X1_859/B PAND2X1_849/a_16_344#
+ PAND2X1_849/m4_208_n4# PAND2X1_849/O PAND2X1_849/a_56_28# PAND2X1_849/CTRL2 PAND2X1_849/CTRL
+ PAND2X1_849/a_76_28# PAND2X1
XPOR2X1_105 VDD GND POR2X1_78/A POR2X1_814/B POR2X1_105/Y POR2X1_105/m4_208_n4# POR2X1_105/O
+ POR2X1_105/CTRL2 POR2X1_105/a_16_28# POR2X1_105/CTRL POR2X1_105/a_76_344# POR2X1_105/a_56_344#
+ POR2X1
XPOR2X1_116 VDD GND POR2X1_114/Y POR2X1_116/A POR2X1_116/Y POR2X1_116/m4_208_n4# POR2X1_116/O
+ POR2X1_116/CTRL2 POR2X1_116/a_16_28# POR2X1_116/CTRL POR2X1_116/a_76_344# POR2X1_116/a_56_344#
+ POR2X1
XPOR2X1_138 VDD GND POR2X1_702/A POR2X1_138/A POR2X1_139/A POR2X1_138/m4_208_n4# POR2X1_138/O
+ POR2X1_138/CTRL2 POR2X1_138/a_16_28# POR2X1_138/CTRL POR2X1_138/a_76_344# POR2X1_138/a_56_344#
+ POR2X1
XPOR2X1_149 VDD GND POR2X1_149/B POR2X1_149/A POR2X1_149/Y POR2X1_149/m4_208_n4# POR2X1_149/O
+ POR2X1_149/CTRL2 POR2X1_149/a_16_28# POR2X1_149/CTRL POR2X1_149/a_76_344# POR2X1_149/a_56_344#
+ POR2X1
XPOR2X1_127 VDD GND POR2X1_7/B POR2X1_394/A POR2X1_127/Y POR2X1_127/m4_208_n4# POR2X1_127/O
+ POR2X1_127/CTRL2 POR2X1_127/a_16_28# POR2X1_127/CTRL POR2X1_127/a_76_344# POR2X1_127/a_56_344#
+ POR2X1
XPAND2X1_70 VDD GND PAND2X1_95/B PAND2X1_3/B PAND2X1_72/A PAND2X1_70/a_16_344# PAND2X1_70/m4_208_n4#
+ PAND2X1_70/O PAND2X1_70/a_56_28# PAND2X1_70/CTRL2 PAND2X1_70/CTRL PAND2X1_70/a_76_28#
+ PAND2X1
XPAND2X1_81 VDD GND PAND2X1_81/B PAND2X1_60/B POR2X1_84/B PAND2X1_81/a_16_344# PAND2X1_81/m4_208_n4#
+ PAND2X1_81/O PAND2X1_81/a_56_28# PAND2X1_81/CTRL2 PAND2X1_81/CTRL PAND2X1_81/a_76_28#
+ PAND2X1
XPOR2X1_34 VDD GND POR2X1_34/B POR2X1_34/A POR2X1_34/Y POR2X1_34/m4_208_n4# POR2X1_34/O
+ POR2X1_34/CTRL2 POR2X1_34/a_16_28# POR2X1_34/CTRL POR2X1_34/a_76_344# POR2X1_34/a_56_344#
+ POR2X1
XPOR2X1_23 VDD GND POR2X1_4/Y POR2X1_14/Y POR2X1_23/Y POR2X1_23/m4_208_n4# POR2X1_23/O
+ POR2X1_23/CTRL2 POR2X1_23/a_16_28# POR2X1_23/CTRL POR2X1_23/a_76_344# POR2X1_23/a_56_344#
+ POR2X1
XPOR2X1_12 VDD GND POR2X1_3/B POR2X1_12/A POR2X1_13/A POR2X1_12/m4_208_n4# POR2X1_12/O
+ POR2X1_12/CTRL2 POR2X1_12/a_16_28# POR2X1_12/CTRL POR2X1_12/a_76_344# POR2X1_12/a_56_344#
+ POR2X1
XPAND2X1_92 VDD GND PAND2X1_8/Y INPUT_1 PAND2X1_93/B PAND2X1_92/a_16_344# PAND2X1_92/m4_208_n4#
+ PAND2X1_92/O PAND2X1_92/a_56_28# PAND2X1_92/CTRL2 PAND2X1_92/CTRL PAND2X1_92/a_76_28#
+ PAND2X1
XPOR2X1_78 VDD GND POR2X1_78/B POR2X1_78/A POR2X1_78/Y POR2X1_78/m4_208_n4# POR2X1_78/O
+ POR2X1_78/CTRL2 POR2X1_78/a_16_28# POR2X1_78/CTRL POR2X1_78/a_76_344# POR2X1_78/a_56_344#
+ POR2X1
XPOR2X1_67 VDD GND POR2X1_55/Y POR2X1_67/A POR2X1_67/Y POR2X1_67/m4_208_n4# POR2X1_67/O
+ POR2X1_67/CTRL2 POR2X1_67/a_16_28# POR2X1_67/CTRL POR2X1_67/a_76_344# POR2X1_67/a_56_344#
+ POR2X1
XPOR2X1_56 VDD GND POR2X1_56/B POR2X1_55/Y POR2X1_56/Y POR2X1_56/m4_208_n4# POR2X1_56/O
+ POR2X1_56/CTRL2 POR2X1_56/a_16_28# POR2X1_56/CTRL POR2X1_56/a_76_344# POR2X1_56/a_56_344#
+ POR2X1
XPOR2X1_45 VDD GND POR2X1_23/Y POR2X1_57/A POR2X1_45/Y POR2X1_45/m4_208_n4# POR2X1_45/O
+ POR2X1_45/CTRL2 POR2X1_45/a_16_28# POR2X1_45/CTRL POR2X1_45/a_76_344# POR2X1_45/a_56_344#
+ POR2X1
XPOR2X1_672 VDD GND POR2X1_416/B POR2X1_672/A POR2X1_672/Y POR2X1_672/m4_208_n4# POR2X1_672/O
+ POR2X1_672/CTRL2 POR2X1_672/a_16_28# POR2X1_672/CTRL POR2X1_672/a_76_344# POR2X1_672/a_56_344#
+ POR2X1
XPOR2X1_89 VDD GND POR2X1_60/A POR2X1_77/Y POR2X1_89/Y POR2X1_89/m4_208_n4# POR2X1_89/O
+ POR2X1_89/CTRL2 POR2X1_89/a_16_28# POR2X1_89/CTRL POR2X1_89/a_76_344# POR2X1_89/a_56_344#
+ POR2X1
XPOR2X1_650 VDD GND POR2X1_640/Y POR2X1_650/A POR2X1_654/B POR2X1_650/m4_208_n4# POR2X1_650/O
+ POR2X1_650/CTRL2 POR2X1_650/a_16_28# POR2X1_650/CTRL POR2X1_650/a_76_344# POR2X1_650/a_56_344#
+ POR2X1
XPOR2X1_661 VDD GND POR2X1_661/B POR2X1_661/A POR2X1_661/Y POR2X1_661/m4_208_n4# POR2X1_661/O
+ POR2X1_661/CTRL2 POR2X1_661/a_16_28# POR2X1_661/CTRL POR2X1_661/a_76_344# POR2X1_661/a_56_344#
+ POR2X1
XPOR2X1_683 VDD GND POR2X1_16/A POR2X1_43/B POR2X1_683/Y POR2X1_683/m4_208_n4# POR2X1_683/O
+ POR2X1_683/CTRL2 POR2X1_683/a_16_28# POR2X1_683/CTRL POR2X1_683/a_76_344# POR2X1_683/a_56_344#
+ POR2X1
XPOR2X1_694 VDD GND POR2X1_257/A POR2X1_425/Y POR2X1_694/Y POR2X1_694/m4_208_n4# POR2X1_694/O
+ POR2X1_694/CTRL2 POR2X1_694/a_16_28# POR2X1_694/CTRL POR2X1_694/a_76_344# POR2X1_694/a_56_344#
+ POR2X1
XPAND2X1_613 VDD GND PAND2X1_55/Y PAND2X1_41/B POR2X1_620/A PAND2X1_613/a_16_344#
+ PAND2X1_613/m4_208_n4# PAND2X1_613/O PAND2X1_613/a_56_28# PAND2X1_613/CTRL2 PAND2X1_613/CTRL
+ PAND2X1_613/a_76_28# PAND2X1
XPAND2X1_602 VDD GND POR2X1_601/Y POR2X1_600/Y PAND2X1_602/Y PAND2X1_602/a_16_344#
+ PAND2X1_602/m4_208_n4# PAND2X1_602/O PAND2X1_602/a_56_28# PAND2X1_602/CTRL2 PAND2X1_602/CTRL
+ PAND2X1_602/a_76_28# PAND2X1
XPAND2X1_624 VDD GND PAND2X1_623/Y PAND2X1_624/A PAND2X1_658/A PAND2X1_624/a_16_344#
+ PAND2X1_624/m4_208_n4# PAND2X1_624/O PAND2X1_624/a_56_28# PAND2X1_624/CTRL2 PAND2X1_624/CTRL
+ PAND2X1_624/a_76_28# PAND2X1
XPAND2X1_635 VDD GND POR2X1_582/Y POR2X1_428/Y PAND2X1_635/Y PAND2X1_635/a_16_344#
+ PAND2X1_635/m4_208_n4# PAND2X1_635/O PAND2X1_635/a_56_28# PAND2X1_635/CTRL2 PAND2X1_635/CTRL
+ PAND2X1_635/a_76_28# PAND2X1
XPAND2X1_646 VDD GND POR2X1_609/Y POR2X1_607/Y PAND2X1_647/B PAND2X1_646/a_16_344#
+ PAND2X1_646/m4_208_n4# PAND2X1_646/O PAND2X1_646/a_56_28# PAND2X1_646/CTRL2 PAND2X1_646/CTRL
+ PAND2X1_646/a_76_28# PAND2X1
XPAND2X1_657 VDD GND PAND2X1_657/B PAND2X1_217/B PAND2X1_659/A PAND2X1_657/a_16_344#
+ PAND2X1_657/m4_208_n4# PAND2X1_657/O PAND2X1_657/a_56_28# PAND2X1_657/CTRL2 PAND2X1_657/CTRL
+ PAND2X1_657/a_76_28# PAND2X1
XPAND2X1_679 VDD GND POR2X1_678/Y POR2X1_676/Y POR2X1_728/B PAND2X1_679/a_16_344#
+ PAND2X1_679/m4_208_n4# PAND2X1_679/O PAND2X1_679/a_56_28# PAND2X1_679/CTRL2 PAND2X1_679/CTRL
+ PAND2X1_679/a_76_28# PAND2X1
XPAND2X1_668 VDD GND POR2X1_416/B POR2X1_83/B POR2X1_669/A PAND2X1_668/a_16_344# PAND2X1_668/m4_208_n4#
+ PAND2X1_668/O PAND2X1_668/a_56_28# PAND2X1_668/CTRL2 PAND2X1_668/CTRL PAND2X1_668/a_76_28#
+ PAND2X1
XPOR2X1_480 VDD GND POR2X1_478/Y POR2X1_480/A D_GATE_479 POR2X1_480/m4_208_n4# POR2X1_480/O
+ POR2X1_480/CTRL2 POR2X1_480/a_16_28# POR2X1_480/CTRL POR2X1_480/a_76_344# POR2X1_480/a_56_344#
+ POR2X1
XPOR2X1_491 VDD GND POR2X1_32/A POR2X1_102/Y POR2X1_491/Y POR2X1_491/m4_208_n4# POR2X1_491/O
+ POR2X1_491/CTRL2 POR2X1_491/a_16_28# POR2X1_491/CTRL POR2X1_491/a_76_344# POR2X1_491/a_56_344#
+ POR2X1
XPAND2X1_421 VDD GND POR2X1_596/A PAND2X1_90/Y POR2X1_448/B PAND2X1_421/a_16_344#
+ PAND2X1_421/m4_208_n4# PAND2X1_421/O PAND2X1_421/a_56_28# PAND2X1_421/CTRL2 PAND2X1_421/CTRL
+ PAND2X1_421/a_76_28# PAND2X1
XPAND2X1_410 VDD GND POR2X1_52/A POR2X1_13/A POR2X1_411/A PAND2X1_410/a_16_344# PAND2X1_410/m4_208_n4#
+ PAND2X1_410/O PAND2X1_410/a_56_28# PAND2X1_410/CTRL2 PAND2X1_410/CTRL PAND2X1_410/a_76_28#
+ PAND2X1
XPAND2X1_432 VDD GND POR2X1_130/A PAND2X1_20/A POR2X1_435/B PAND2X1_432/a_16_344#
+ PAND2X1_432/m4_208_n4# PAND2X1_432/O PAND2X1_432/a_56_28# PAND2X1_432/CTRL2 PAND2X1_432/CTRL
+ PAND2X1_432/a_76_28# PAND2X1
XPAND2X1_454 VDD GND PAND2X1_454/B PAND2X1_446/Y PAND2X1_466/B PAND2X1_454/a_16_344#
+ PAND2X1_454/m4_208_n4# PAND2X1_454/O PAND2X1_454/a_56_28# PAND2X1_454/CTRL2 PAND2X1_454/CTRL
+ PAND2X1_454/a_76_28# PAND2X1
XPAND2X1_443 VDD GND POR2X1_441/Y POR2X1_91/Y PAND2X1_443/Y PAND2X1_443/a_16_344#
+ PAND2X1_443/m4_208_n4# PAND2X1_443/O PAND2X1_443/a_56_28# PAND2X1_443/CTRL2 PAND2X1_443/CTRL
+ PAND2X1_443/a_76_28# PAND2X1
XPAND2X1_476 VDD GND PAND2X1_473/Y PAND2X1_476/A PAND2X1_479/B PAND2X1_476/a_16_344#
+ PAND2X1_475/m4_208_n4# PAND2X1_476/O PAND2X1_476/a_56_28# PAND2X1_476/CTRL2 PAND2X1_476/CTRL
+ PAND2X1_476/a_76_28# PAND2X1
XPAND2X1_498 VDD GND POR2X1_188/Y PAND2X1_72/A POR2X1_501/B PAND2X1_498/a_16_344#
+ POR2X1_723/m4_208_n4# PAND2X1_498/O PAND2X1_498/a_56_28# PAND2X1_498/CTRL2 PAND2X1_498/CTRL
+ PAND2X1_498/a_76_28# PAND2X1
XPAND2X1_487 VDD GND PAND2X1_96/B PAND2X1_23/Y POR2X1_489/B PAND2X1_487/a_16_344#
+ POR2X1_489/m4_208_n4# PAND2X1_487/O PAND2X1_487/a_56_28# PAND2X1_487/CTRL2 PAND2X1_487/CTRL
+ PAND2X1_487/a_76_28# PAND2X1
XPAND2X1_465 VDD GND PAND2X1_465/B PAND2X1_455/Y PAND2X1_471/B PAND2X1_465/a_16_344#
+ PAND2X1_465/m4_208_n4# PAND2X1_465/O PAND2X1_465/a_56_28# PAND2X1_465/CTRL2 PAND2X1_465/CTRL
+ PAND2X1_465/a_76_28# PAND2X1
XPAND2X1_262 VDD GND PAND2X1_63/Y PAND2X1_41/B POR2X1_786/A PAND2X1_262/a_16_344#
+ PAND2X1_262/m4_208_n4# PAND2X1_262/O PAND2X1_262/a_56_28# PAND2X1_262/CTRL2 PAND2X1_262/CTRL
+ PAND2X1_262/a_76_28# PAND2X1
XPAND2X1_273 VDD GND POR2X1_407/A PAND2X1_69/A POR2X1_274/A PAND2X1_273/a_16_344#
+ PAND2X1_273/m4_208_n4# PAND2X1_273/O PAND2X1_273/a_56_28# PAND2X1_273/CTRL2 PAND2X1_273/CTRL
+ PAND2X1_273/a_76_28# PAND2X1
XPAND2X1_251 VDD GND POR2X1_105/Y PAND2X1_52/B POR2X1_343/A PAND2X1_251/a_16_344#
+ PAND2X1_251/m4_208_n4# PAND2X1_251/O PAND2X1_251/a_56_28# PAND2X1_251/CTRL2 PAND2X1_251/CTRL
+ PAND2X1_251/a_76_28# PAND2X1
XPAND2X1_240 VDD GND POR2X1_234/Y POR2X1_232/Y PAND2X1_243/B PAND2X1_240/a_16_344#
+ PAND2X1_240/m4_208_n4# PAND2X1_240/O PAND2X1_240/a_56_28# PAND2X1_240/CTRL2 PAND2X1_240/CTRL
+ PAND2X1_240/a_76_28# PAND2X1
XPAND2X1_284 VDD GND POR2X1_280/Y POR2X1_279/Y PAND2X1_284/Y PAND2X1_284/a_16_344#
+ PAND2X1_284/m4_208_n4# PAND2X1_284/O PAND2X1_284/a_56_28# PAND2X1_284/CTRL2 PAND2X1_284/CTRL
+ PAND2X1_284/a_76_28# PAND2X1
XPAND2X1_295 VDD GND POR2X1_294/Y PAND2X1_60/B POR2X1_346/A PAND2X1_295/a_16_344#
+ PAND2X1_295/m4_208_n4# PAND2X1_295/O PAND2X1_295/a_56_28# PAND2X1_295/CTRL2 PAND2X1_295/CTRL
+ PAND2X1_295/a_76_28# PAND2X1
XPOR2X1_309 VDD GND POR2X1_43/B POR2X1_283/A POR2X1_309/Y POR2X1_309/m4_208_n4# POR2X1_309/O
+ POR2X1_309/CTRL2 POR2X1_309/a_16_28# POR2X1_309/CTRL POR2X1_309/a_76_344# POR2X1_309/a_56_344#
+ POR2X1
XPOR2X1_821 VDD GND POR2X1_41/B POR2X1_72/B POR2X1_821/Y POR2X1_821/m4_208_n4# POR2X1_821/O
+ POR2X1_821/CTRL2 POR2X1_821/a_16_28# POR2X1_821/CTRL POR2X1_821/a_76_344# POR2X1_821/a_56_344#
+ POR2X1
XPOR2X1_810 VDD GND POR2X1_774/Y POR2X1_809/Y POR2X1_812/B POR2X1_810/m4_208_n4# POR2X1_810/O
+ POR2X1_810/CTRL2 POR2X1_810/a_16_28# POR2X1_810/CTRL POR2X1_810/a_76_344# POR2X1_810/a_56_344#
+ POR2X1
XPOR2X1_854 VDD GND POR2X1_854/B POR2X1_567/B POR2X1_856/B POR2X1_854/m4_208_n4# POR2X1_854/O
+ POR2X1_854/CTRL2 POR2X1_854/a_16_28# POR2X1_854/CTRL POR2X1_854/a_76_344# POR2X1_854/a_56_344#
+ POR2X1
XPOR2X1_843 VDD GND POR2X1_343/A POR2X1_287/B POR2X1_850/A POR2X1_843/m4_208_n4# POR2X1_843/O
+ POR2X1_843/CTRL2 POR2X1_843/a_16_28# POR2X1_843/CTRL POR2X1_843/a_76_344# POR2X1_843/a_56_344#
+ POR2X1
XPOR2X1_832 VDD GND POR2X1_832/B POR2X1_832/A POR2X1_832/Y POR2X1_832/m4_208_n4# POR2X1_832/O
+ POR2X1_832/CTRL2 POR2X1_832/a_16_28# POR2X1_832/CTRL POR2X1_832/a_76_344# POR2X1_832/a_56_344#
+ POR2X1
XPOR2X1_865 VDD GND POR2X1_865/B POR2X1_862/Y POR2X1_866/A POR2X1_865/m4_208_n4# POR2X1_865/O
+ POR2X1_865/CTRL2 POR2X1_865/a_16_28# POR2X1_865/CTRL POR2X1_865/a_76_344# POR2X1_865/a_56_344#
+ POR2X1
XPAND2X1_806 VDD GND PAND2X1_736/A PAND2X1_362/A PAND2X1_807/B PAND2X1_806/a_16_344#
+ PAND2X1_806/m4_208_n4# PAND2X1_806/O PAND2X1_806/a_56_28# PAND2X1_806/CTRL2 PAND2X1_806/CTRL
+ PAND2X1_806/a_76_28# PAND2X1
XPAND2X1_817 VDD GND PAND2X1_381/Y D_INPUT_1 POR2X1_847/B PAND2X1_817/a_16_344# PAND2X1_817/m4_208_n4#
+ PAND2X1_817/O PAND2X1_817/a_56_28# PAND2X1_817/CTRL2 PAND2X1_817/CTRL PAND2X1_817/a_76_28#
+ PAND2X1
XPAND2X1_828 VDD GND POR2X1_599/A POR2X1_409/B POR2X1_829/A PAND2X1_828/a_16_344#
+ PAND2X1_828/m4_208_n4# PAND2X1_828/O PAND2X1_828/a_56_28# PAND2X1_828/CTRL2 PAND2X1_828/CTRL
+ PAND2X1_828/a_76_28# PAND2X1
XPAND2X1_839 VDD GND PAND2X1_839/B PAND2X1_835/Y PAND2X1_852/B PAND2X1_839/a_16_344#
+ PAND2X1_839/m4_208_n4# PAND2X1_839/O PAND2X1_839/a_56_28# PAND2X1_839/CTRL2 PAND2X1_839/CTRL
+ PAND2X1_839/a_76_28# PAND2X1
XPOR2X1_106 VDD GND POR2X1_48/A POR2X1_251/A POR2X1_106/Y POR2X1_106/m4_208_n4# POR2X1_106/O
+ POR2X1_106/CTRL2 POR2X1_106/a_16_28# POR2X1_106/CTRL POR2X1_106/a_76_344# POR2X1_106/a_56_344#
+ POR2X1
XPOR2X1_117 VDD GND POR2X1_63/Y POR2X1_72/B POR2X1_117/Y POR2X1_117/m4_208_n4# POR2X1_117/O
+ POR2X1_117/CTRL2 POR2X1_117/a_16_28# POR2X1_117/CTRL POR2X1_117/a_76_344# POR2X1_117/a_56_344#
+ POR2X1
XPOR2X1_128 VDD GND POR2X1_128/B POR2X1_128/A POR2X1_140/B POR2X1_128/m4_208_n4# POR2X1_128/O
+ POR2X1_128/CTRL2 POR2X1_128/a_16_28# POR2X1_128/CTRL POR2X1_128/a_76_344# POR2X1_128/a_56_344#
+ POR2X1
XPOR2X1_139 VDD GND POR2X1_137/Y POR2X1_139/A POR2X1_139/Y POR2X1_139/m4_208_n4# POR2X1_139/O
+ POR2X1_139/CTRL2 POR2X1_139/a_16_28# POR2X1_139/CTRL POR2X1_139/a_76_344# POR2X1_139/a_56_344#
+ POR2X1
XPAND2X1_71 VDD GND PAND2X1_63/B POR2X1_68/B PAND2X1_71/Y PAND2X1_71/a_16_344# PAND2X1_71/m4_208_n4#
+ PAND2X1_71/O PAND2X1_71/a_56_28# PAND2X1_71/CTRL2 PAND2X1_71/CTRL PAND2X1_71/a_76_28#
+ PAND2X1
XPAND2X1_60 VDD GND PAND2X1_60/B PAND2X1_39/B POR2X1_61/A PAND2X1_60/a_16_344# PAND2X1_60/m4_208_n4#
+ PAND2X1_60/O PAND2X1_60/a_56_28# PAND2X1_60/CTRL2 PAND2X1_60/CTRL PAND2X1_60/a_76_28#
+ PAND2X1
XPOR2X1_35 VDD GND POR2X1_35/B POR2X1_34/Y POR2X1_35/Y POR2X1_35/m4_208_n4# POR2X1_35/O
+ POR2X1_35/CTRL2 POR2X1_35/a_16_28# POR2X1_35/CTRL POR2X1_35/a_76_344# POR2X1_35/a_56_344#
+ POR2X1
XPOR2X1_24 VDD GND POR2X1_43/B POR2X1_23/Y POR2X1_24/Y POR2X1_24/m4_208_n4# POR2X1_24/O
+ POR2X1_24/CTRL2 POR2X1_24/a_16_28# POR2X1_24/CTRL POR2X1_24/a_76_344# POR2X1_24/a_56_344#
+ POR2X1
XPOR2X1_13 VDD GND POR2X1_41/B POR2X1_13/A POR2X1_13/Y POR2X1_13/m4_208_n4# POR2X1_13/O
+ POR2X1_13/CTRL2 POR2X1_13/a_16_28# POR2X1_13/CTRL POR2X1_13/a_76_344# POR2X1_13/a_56_344#
+ POR2X1
XPAND2X1_93 VDD GND PAND2X1_93/B POR2X1_66/A POR2X1_98/B PAND2X1_93/a_16_344# PAND2X1_93/m4_208_n4#
+ PAND2X1_93/O PAND2X1_93/a_56_28# PAND2X1_93/CTRL2 PAND2X1_93/CTRL PAND2X1_93/a_76_28#
+ PAND2X1
XPAND2X1_82 VDD GND POR2X1_38/B PAND2X1_94/A PAND2X1_82/Y PAND2X1_82/a_16_344# PAND2X1_82/m4_208_n4#
+ PAND2X1_82/O PAND2X1_82/a_56_28# PAND2X1_82/CTRL2 PAND2X1_82/CTRL PAND2X1_82/a_76_28#
+ PAND2X1
XPOR2X1_68 VDD GND POR2X1_68/B POR2X1_68/A POR2X1_68/Y POR2X1_68/m4_208_n4# POR2X1_68/O
+ POR2X1_68/CTRL2 POR2X1_68/a_16_28# POR2X1_68/CTRL POR2X1_68/a_76_344# POR2X1_68/a_56_344#
+ POR2X1
XPOR2X1_46 VDD GND INPUT_1 POR2X1_14/Y POR2X1_46/Y POR2X1_46/m4_208_n4# POR2X1_46/O
+ POR2X1_46/CTRL2 POR2X1_46/a_16_28# POR2X1_46/CTRL POR2X1_46/a_76_344# POR2X1_46/a_56_344#
+ POR2X1
XPOR2X1_57 VDD GND POR2X1_5/Y POR2X1_57/A POR2X1_57/Y POR2X1_57/m4_208_n4# POR2X1_57/O
+ POR2X1_57/CTRL2 POR2X1_57/a_16_28# POR2X1_57/CTRL POR2X1_57/a_76_344# POR2X1_57/a_56_344#
+ POR2X1
XPOR2X1_79 VDD GND POR2X1_20/B POR2X1_79/A POR2X1_79/Y POR2X1_79/m4_208_n4# POR2X1_79/O
+ POR2X1_79/CTRL2 POR2X1_79/a_16_28# POR2X1_79/CTRL POR2X1_79/a_76_344# POR2X1_79/a_56_344#
+ POR2X1
XPOR2X1_640 VDD GND POR2X1_633/Y POR2X1_640/A POR2X1_640/Y POR2X1_640/m4_208_n4# POR2X1_640/O
+ POR2X1_640/CTRL2 POR2X1_640/a_16_28# POR2X1_640/CTRL POR2X1_640/a_76_344# POR2X1_640/a_56_344#
+ POR2X1
XPOR2X1_651 VDD GND POR2X1_638/Y POR2X1_639/Y POR2X1_651/Y POR2X1_651/m4_208_n4# POR2X1_651/O
+ POR2X1_651/CTRL2 POR2X1_651/a_16_28# POR2X1_651/CTRL POR2X1_651/a_76_344# POR2X1_651/a_56_344#
+ POR2X1
XPOR2X1_662 VDD GND POR2X1_660/Y POR2X1_661/Y POR2X1_662/Y POR2X1_662/m4_208_n4# POR2X1_662/O
+ POR2X1_662/CTRL2 POR2X1_662/a_16_28# POR2X1_662/CTRL POR2X1_662/a_76_344# POR2X1_662/a_56_344#
+ POR2X1
XPOR2X1_673 VDD GND POR2X1_673/B POR2X1_673/A POR2X1_673/Y POR2X1_673/m4_208_n4# POR2X1_673/O
+ POR2X1_673/CTRL2 POR2X1_673/a_16_28# POR2X1_673/CTRL POR2X1_673/a_76_344# POR2X1_673/a_56_344#
+ POR2X1
XPOR2X1_684 VDD GND POR2X1_13/A POR2X1_42/Y POR2X1_684/Y POR2X1_684/m4_208_n4# POR2X1_684/O
+ POR2X1_684/CTRL2 POR2X1_684/a_16_28# POR2X1_684/CTRL POR2X1_684/a_76_344# POR2X1_684/a_56_344#
+ POR2X1
XPOR2X1_695 VDD GND POR2X1_23/Y POR2X1_48/A POR2X1_695/Y POR2X1_695/m4_208_n4# POR2X1_695/O
+ POR2X1_695/CTRL2 POR2X1_695/a_16_28# POR2X1_695/CTRL POR2X1_695/a_76_344# POR2X1_695/a_56_344#
+ POR2X1
XPAND2X1_603 VDD GND POR2X1_68/A POR2X1_260/B POR2X1_605/B PAND2X1_603/a_16_344# PAND2X1_603/m4_208_n4#
+ PAND2X1_603/O PAND2X1_603/a_56_28# PAND2X1_603/CTRL2 PAND2X1_603/CTRL PAND2X1_603/a_76_28#
+ PAND2X1
XPAND2X1_614 VDD GND POR2X1_257/A POR2X1_77/Y POR2X1_754/A PAND2X1_614/a_16_344# PAND2X1_614/m4_208_n4#
+ PAND2X1_614/O PAND2X1_614/a_56_28# PAND2X1_614/CTRL2 PAND2X1_614/CTRL PAND2X1_614/a_76_28#
+ PAND2X1
XPAND2X1_636 VDD GND POR2X1_584/Y POR2X1_583/Y PAND2X1_639/B PAND2X1_636/a_16_344#
+ PAND2X1_636/m4_208_n4# PAND2X1_636/O PAND2X1_636/a_56_28# PAND2X1_636/CTRL2 PAND2X1_636/CTRL
+ PAND2X1_636/a_76_28# PAND2X1
XPAND2X1_625 VDD GND POR2X1_294/A POR2X1_66/Y POR2X1_631/A PAND2X1_625/a_16_344# PAND2X1_625/m4_208_n4#
+ PAND2X1_625/O PAND2X1_625/a_56_28# PAND2X1_625/CTRL2 PAND2X1_625/CTRL PAND2X1_625/a_76_28#
+ PAND2X1
XPAND2X1_647 VDD GND PAND2X1_647/B POR2X1_612/Y PAND2X1_656/B PAND2X1_647/a_16_344#
+ PAND2X1_400/m4_208_n4# PAND2X1_647/O PAND2X1_647/a_56_28# PAND2X1_647/CTRL2 PAND2X1_647/CTRL
+ PAND2X1_647/a_76_28# PAND2X1
XPAND2X1_669 VDD GND POR2X1_668/Y POR2X1_750/B POR2X1_720/A PAND2X1_669/a_16_344#
+ PAND2X1_669/m4_208_n4# PAND2X1_669/O PAND2X1_669/a_56_28# PAND2X1_669/CTRL2 PAND2X1_669/CTRL
+ PAND2X1_669/a_76_28# PAND2X1
XPAND2X1_658 VDD GND PAND2X1_658/B PAND2X1_658/A PAND2X1_659/B PAND2X1_658/a_16_344#
+ PAND2X1_658/m4_208_n4# PAND2X1_658/O PAND2X1_658/a_56_28# PAND2X1_658/CTRL2 PAND2X1_658/CTRL
+ PAND2X1_658/a_76_28# PAND2X1
XPOR2X1_470 VDD GND POR2X1_466/Y POR2X1_467/Y POR2X1_477/B POR2X1_470/m4_208_n4# POR2X1_470/O
+ POR2X1_470/CTRL2 POR2X1_470/a_16_28# POR2X1_470/CTRL POR2X1_470/a_76_344# POR2X1_470/a_56_344#
+ POR2X1
XPOR2X1_492 VDD GND POR2X1_60/A POR2X1_394/A POR2X1_492/Y POR2X1_492/m4_208_n4# POR2X1_492/O
+ POR2X1_492/CTRL2 POR2X1_492/a_16_28# POR2X1_492/CTRL POR2X1_492/a_76_344# POR2X1_492/a_56_344#
+ POR2X1
XPOR2X1_481 VDD GND POR2X1_7/B POR2X1_481/A POR2X1_481/Y POR2X1_481/m4_208_n4# POR2X1_481/O
+ POR2X1_481/CTRL2 POR2X1_481/a_16_28# POR2X1_481/CTRL POR2X1_481/a_76_344# POR2X1_481/a_56_344#
+ POR2X1
XPAND2X1_411 VDD GND POR2X1_410/Y POR2X1_814/B POR2X1_461/B PAND2X1_411/a_16_344#
+ PAND2X1_411/m4_208_n4# PAND2X1_411/O PAND2X1_411/a_56_28# PAND2X1_411/CTRL2 PAND2X1_411/CTRL
+ PAND2X1_411/a_76_28# PAND2X1
XPAND2X1_422 VDD GND PAND2X1_93/B POR2X1_260/B POR2X1_448/A PAND2X1_422/a_16_344#
+ PAND2X1_422/m4_208_n4# PAND2X1_422/O PAND2X1_422/a_56_28# PAND2X1_422/CTRL2 PAND2X1_422/CTRL
+ PAND2X1_422/a_76_28# PAND2X1
XPAND2X1_400 VDD GND POR2X1_394/Y POR2X1_393/Y PAND2X1_403/B PAND2X1_400/a_16_344#
+ PAND2X1_400/m4_208_n4# PAND2X1_400/O PAND2X1_400/a_56_28# PAND2X1_400/CTRL2 PAND2X1_400/CTRL
+ PAND2X1_400/a_76_28# PAND2X1
XPAND2X1_455 VDD GND PAND2X1_445/Y PAND2X1_76/Y PAND2X1_455/Y PAND2X1_455/a_16_344#
+ PAND2X1_455/m4_208_n4# PAND2X1_455/O PAND2X1_455/a_56_28# PAND2X1_455/CTRL2 PAND2X1_455/CTRL
+ PAND2X1_455/a_76_28# PAND2X1
XPAND2X1_433 VDD GND POR2X1_407/A PAND2X1_72/A POR2X1_832/A PAND2X1_433/a_16_344#
+ PAND2X1_433/m4_208_n4# PAND2X1_433/O PAND2X1_433/a_56_28# PAND2X1_433/CTRL2 PAND2X1_433/CTRL
+ PAND2X1_433/a_76_28# PAND2X1
XPAND2X1_444 VDD GND PAND2X1_443/Y POR2X1_442/Y PAND2X1_444/Y PAND2X1_444/a_16_344#
+ PAND2X1_444/m4_208_n4# PAND2X1_444/O PAND2X1_444/a_56_28# PAND2X1_444/CTRL2 PAND2X1_444/CTRL
+ PAND2X1_444/a_76_28# PAND2X1
XPAND2X1_488 VDD GND POR2X1_814/A POR2X1_260/A POR2X1_489/A PAND2X1_488/a_16_344#
+ PAND2X1_488/m4_208_n4# PAND2X1_488/O PAND2X1_488/a_56_28# PAND2X1_488/CTRL2 PAND2X1_488/CTRL
+ PAND2X1_488/a_76_28# PAND2X1
XPAND2X1_466 VDD GND PAND2X1_466/B PAND2X1_466/A PAND2X1_470/A PAND2X1_466/a_16_344#
+ PAND2X1_466/m4_208_n4# PAND2X1_466/O PAND2X1_466/a_56_28# PAND2X1_466/CTRL2 PAND2X1_466/CTRL
+ PAND2X1_466/a_76_28# PAND2X1
XPAND2X1_477 VDD GND PAND2X1_477/B PAND2X1_477/A PAND2X1_478/B PAND2X1_477/a_16_344#
+ PAND2X1_477/m4_208_n4# PAND2X1_477/O PAND2X1_477/a_56_28# PAND2X1_477/CTRL2 PAND2X1_477/CTRL
+ PAND2X1_477/a_76_28# PAND2X1
XPAND2X1_499 VDD GND POR2X1_496/Y POR2X1_495/Y PAND2X1_499/Y PAND2X1_499/a_16_344#
+ PAND2X1_499/m4_208_n4# PAND2X1_499/O PAND2X1_499/a_56_28# PAND2X1_499/CTRL2 PAND2X1_499/CTRL
+ PAND2X1_499/a_76_28# PAND2X1
XPAND2X1_230 VDD GND PAND2X1_32/B PAND2X1_6/Y POR2X1_231/A PAND2X1_230/a_16_344# PAND2X1_230/m4_208_n4#
+ PAND2X1_230/O PAND2X1_230/a_56_28# PAND2X1_230/CTRL2 PAND2X1_230/CTRL PAND2X1_230/a_76_28#
+ PAND2X1
XPAND2X1_263 VDD GND PAND2X1_90/A PAND2X1_58/A POR2X1_266/A PAND2X1_263/a_16_344#
+ PAND2X1_263/m4_208_n4# PAND2X1_263/O PAND2X1_263/a_56_28# PAND2X1_263/CTRL2 PAND2X1_263/CTRL
+ PAND2X1_263/a_76_28# PAND2X1
XPAND2X1_241 VDD GND POR2X1_238/Y POR2X1_237/Y PAND2X1_241/Y PAND2X1_241/a_16_344#
+ PAND2X1_241/m4_208_n4# PAND2X1_241/O PAND2X1_241/a_56_28# PAND2X1_241/CTRL2 PAND2X1_241/CTRL
+ PAND2X1_241/a_76_28# PAND2X1
XPAND2X1_252 VDD GND PAND2X1_60/B PAND2X1_55/Y POR2X1_483/B PAND2X1_252/a_16_344#
+ PAND2X1_252/m4_208_n4# PAND2X1_252/O PAND2X1_252/a_56_28# PAND2X1_252/CTRL2 PAND2X1_252/CTRL
+ PAND2X1_252/a_76_28# PAND2X1
XPAND2X1_285 VDD GND POR2X1_282/Y POR2X1_281/Y PAND2X1_286/B PAND2X1_285/a_16_344#
+ PAND2X1_567/m4_208_n4# PAND2X1_285/O PAND2X1_285/a_56_28# PAND2X1_285/CTRL2 PAND2X1_285/CTRL
+ PAND2X1_285/a_76_28# PAND2X1
XPAND2X1_296 VDD GND POR2X1_55/Y POR2X1_42/Y POR2X1_297/A PAND2X1_296/a_16_344# PAND2X1_296/m4_208_n4#
+ PAND2X1_296/O PAND2X1_296/a_56_28# PAND2X1_296/CTRL2 PAND2X1_296/CTRL PAND2X1_296/a_76_28#
+ PAND2X1
XPAND2X1_274 VDD GND POR2X1_273/Y POR2X1_272/Y POR2X1_275/A PAND2X1_274/a_16_344#
+ PAND2X1_274/m4_208_n4# PAND2X1_274/O PAND2X1_274/a_56_28# PAND2X1_274/CTRL2 PAND2X1_274/CTRL
+ PAND2X1_274/a_76_28# PAND2X1
XPOR2X1_811 VDD GND POR2X1_811/B POR2X1_811/A POR2X1_812/A POR2X1_811/m4_208_n4# POR2X1_811/O
+ POR2X1_811/CTRL2 POR2X1_811/a_16_28# POR2X1_811/CTRL POR2X1_811/a_76_344# POR2X1_811/a_56_344#
+ POR2X1
XPOR2X1_800 VDD GND POR2X1_687/Y POR2X1_800/A POR2X1_801/A POR2X1_800/m4_208_n4# POR2X1_800/O
+ POR2X1_800/CTRL2 POR2X1_800/a_16_28# POR2X1_800/CTRL POR2X1_800/a_76_344# POR2X1_800/a_56_344#
+ POR2X1
XPOR2X1_822 VDD GND POR2X1_65/A POR2X1_102/Y POR2X1_822/Y POR2X1_822/m4_208_n4# POR2X1_822/O
+ POR2X1_822/CTRL2 POR2X1_822/a_16_28# POR2X1_822/CTRL POR2X1_822/a_76_344# POR2X1_822/a_56_344#
+ POR2X1
XPOR2X1_833 VDD GND POR2X1_483/A POR2X1_833/A POR2X1_840/B POR2X1_833/m4_208_n4# POR2X1_833/O
+ POR2X1_833/CTRL2 POR2X1_833/a_16_28# POR2X1_833/CTRL POR2X1_833/a_76_344# POR2X1_833/a_56_344#
+ POR2X1
XPOR2X1_844 VDD GND POR2X1_844/B POR2X1_523/Y POR2X1_849/B POR2X1_844/m4_208_n4# POR2X1_844/O
+ POR2X1_844/CTRL2 POR2X1_844/a_16_28# POR2X1_844/CTRL POR2X1_844/a_76_344# POR2X1_844/a_56_344#
+ POR2X1
XPOR2X1_855 VDD GND POR2X1_855/B POR2X1_855/A POR2X1_855/Y POR2X1_855/m4_208_n4# POR2X1_855/O
+ POR2X1_855/CTRL2 POR2X1_855/a_16_28# POR2X1_855/CTRL POR2X1_855/a_76_344# POR2X1_855/a_56_344#
+ POR2X1
XPOR2X1_866 VDD GND POR2X1_866/B POR2X1_866/A D_GATE_865 POR2X1_866/m4_208_n4# POR2X1_866/O
+ POR2X1_866/CTRL2 POR2X1_866/a_16_28# POR2X1_866/CTRL POR2X1_866/a_76_344# POR2X1_866/a_56_344#
+ POR2X1
XPAND2X1_818 VDD GND POR2X1_376/B POR2X1_5/Y POR2X1_820/B PAND2X1_818/a_16_344# PAND2X1_818/m4_208_n4#
+ PAND2X1_818/O PAND2X1_818/a_56_28# PAND2X1_818/CTRL2 PAND2X1_818/CTRL PAND2X1_818/a_76_28#
+ PAND2X1
XPAND2X1_807 VDD GND PAND2X1_807/B PAND2X1_805/Y PAND2X1_811/A PAND2X1_807/a_16_344#
+ PAND2X1_807/m4_208_n4# PAND2X1_807/O PAND2X1_807/a_56_28# PAND2X1_807/CTRL2 PAND2X1_807/CTRL
+ PAND2X1_807/a_76_28# PAND2X1
XPAND2X1_829 VDD GND POR2X1_828/Y PAND2X1_65/B POR2X1_855/A PAND2X1_829/a_16_344#
+ PAND2X1_829/m4_208_n4# PAND2X1_829/O PAND2X1_829/a_56_28# PAND2X1_829/CTRL2 PAND2X1_829/CTRL
+ PAND2X1_829/a_76_28# PAND2X1
XPOR2X1_107 VDD GND POR2X1_65/A POR2X1_77/Y POR2X1_107/Y POR2X1_107/m4_208_n4# POR2X1_107/O
+ POR2X1_107/CTRL2 POR2X1_107/a_16_28# POR2X1_107/CTRL POR2X1_107/a_76_344# POR2X1_107/a_56_344#
+ POR2X1
XPOR2X1_118 VDD GND POR2X1_72/B POR2X1_77/Y POR2X1_118/Y POR2X1_118/m4_208_n4# POR2X1_118/O
+ POR2X1_118/CTRL2 POR2X1_118/a_16_28# POR2X1_118/CTRL POR2X1_118/a_76_344# POR2X1_118/a_56_344#
+ POR2X1
XPOR2X1_129 VDD GND POR2X1_29/A POR2X1_37/Y POR2X1_129/Y POR2X1_129/m4_208_n4# POR2X1_129/O
+ POR2X1_129/CTRL2 POR2X1_129/a_16_28# POR2X1_129/CTRL POR2X1_129/a_76_344# POR2X1_129/a_56_344#
+ POR2X1
XPAND2X1_61 VDD GND POR2X1_60/Y POR2X1_58/Y PAND2X1_61/Y PAND2X1_61/a_16_344# PAND2X1_61/m4_208_n4#
+ PAND2X1_61/O PAND2X1_61/a_56_28# PAND2X1_61/CTRL2 PAND2X1_61/CTRL PAND2X1_61/a_76_28#
+ PAND2X1
XPAND2X1_50 VDD GND D_INPUT_7 D_INPUT_6 PAND2X1_95/B PAND2X1_50/a_16_344# PAND2X1_50/m4_208_n4#
+ PAND2X1_50/O PAND2X1_50/a_56_28# PAND2X1_50/CTRL2 PAND2X1_50/CTRL PAND2X1_50/a_76_28#
+ PAND2X1
XPAND2X1_72 VDD GND PAND2X1_71/Y PAND2X1_72/A PAND2X1_72/Y PAND2X1_72/a_16_344# PAND2X1_72/m4_208_n4#
+ PAND2X1_72/O PAND2X1_72/a_56_28# PAND2X1_72/CTRL2 PAND2X1_72/CTRL PAND2X1_72/a_76_28#
+ PAND2X1
XPOR2X1_14 VDD GND INPUT_2 INPUT_3 POR2X1_14/Y POR2X1_14/m4_208_n4# POR2X1_14/O POR2X1_14/CTRL2
+ POR2X1_14/a_16_28# POR2X1_14/CTRL POR2X1_14/a_76_344# POR2X1_14/a_56_344# POR2X1
XPOR2X1_25 VDD GND D_INPUT_6 INPUT_7 POR2X1_25/Y POR2X1_25/m4_208_n4# POR2X1_25/O
+ POR2X1_25/CTRL2 POR2X1_25/a_16_28# POR2X1_25/CTRL POR2X1_25/a_76_344# POR2X1_25/a_56_344#
+ POR2X1
XPAND2X1_83 VDD GND PAND2X1_82/Y POR2X1_66/A POR2X1_84/A PAND2X1_83/a_16_344# PAND2X1_83/m4_208_n4#
+ PAND2X1_83/O PAND2X1_83/a_56_28# PAND2X1_83/CTRL2 PAND2X1_83/CTRL PAND2X1_83/a_76_28#
+ PAND2X1
XPAND2X1_94 VDD GND POR2X1_54/Y PAND2X1_94/A PAND2X1_94/Y PAND2X1_94/a_16_344# PAND2X1_94/m4_208_n4#
+ PAND2X1_94/O PAND2X1_94/a_56_28# PAND2X1_94/CTRL2 PAND2X1_94/CTRL PAND2X1_94/a_76_28#
+ PAND2X1
XPOR2X1_69 VDD GND POR2X1_39/B POR2X1_69/A POR2X1_69/Y POR2X1_69/m4_208_n4# POR2X1_69/O
+ POR2X1_69/CTRL2 POR2X1_69/a_16_28# POR2X1_69/CTRL POR2X1_69/a_76_344# POR2X1_69/a_56_344#
+ POR2X1
XPOR2X1_58 VDD GND POR2X1_43/B POR2X1_49/Y POR2X1_58/Y POR2X1_58/m4_208_n4# POR2X1_58/O
+ POR2X1_58/CTRL2 POR2X1_58/a_16_28# POR2X1_58/CTRL POR2X1_58/a_76_344# POR2X1_58/a_56_344#
+ POR2X1
XPOR2X1_47 VDD GND POR2X1_25/Y POR2X1_51/B POR2X1_48/A POR2X1_47/m4_208_n4# POR2X1_47/O
+ POR2X1_47/CTRL2 POR2X1_47/a_16_28# POR2X1_47/CTRL POR2X1_47/a_76_344# POR2X1_47/a_56_344#
+ POR2X1
XPOR2X1_36 VDD GND POR2X1_36/B POR2X1_22/A POR2X1_39/B POR2X1_36/m4_208_n4# POR2X1_36/O
+ POR2X1_36/CTRL2 POR2X1_36/a_16_28# POR2X1_36/CTRL POR2X1_36/a_76_344# POR2X1_36/a_56_344#
+ POR2X1
XPOR2X1_630 VDD GND POR2X1_630/B POR2X1_630/A POR2X1_632/B POR2X1_630/m4_208_n4# POR2X1_630/O
+ POR2X1_630/CTRL2 POR2X1_630/a_16_28# POR2X1_630/CTRL POR2X1_630/a_76_344# POR2X1_630/a_56_344#
+ POR2X1
XPOR2X1_641 VDD GND POR2X1_341/A POR2X1_267/B POR2X1_650/A POR2X1_641/m4_208_n4# POR2X1_641/O
+ POR2X1_641/CTRL2 POR2X1_641/a_16_28# POR2X1_641/CTRL POR2X1_641/a_76_344# POR2X1_641/a_56_344#
+ POR2X1
XPOR2X1_663 VDD GND POR2X1_663/B POR2X1_662/Y D_GATE_662 POR2X1_663/m4_208_n4# POR2X1_663/O
+ POR2X1_663/CTRL2 POR2X1_663/a_16_28# POR2X1_663/CTRL POR2X1_663/a_76_344# POR2X1_663/a_56_344#
+ POR2X1
XPOR2X1_652 VDD GND POR2X1_440/Y POR2X1_652/A POR2X1_652/Y POR2X1_652/m4_208_n4# POR2X1_652/O
+ POR2X1_652/CTRL2 POR2X1_652/a_16_28# POR2X1_652/CTRL POR2X1_652/a_76_344# POR2X1_652/a_56_344#
+ POR2X1
XPOR2X1_674 VDD GND POR2X1_72/B POR2X1_760/A POR2X1_674/Y POR2X1_674/m4_208_n4# POR2X1_674/O
+ POR2X1_674/CTRL2 POR2X1_674/a_16_28# POR2X1_674/CTRL POR2X1_674/a_76_344# POR2X1_674/a_56_344#
+ POR2X1
XPOR2X1_696 VDD GND POR2X1_83/B POR2X1_376/B POR2X1_696/Y POR2X1_696/m4_208_n4# POR2X1_696/O
+ POR2X1_696/CTRL2 POR2X1_696/a_16_28# POR2X1_696/CTRL POR2X1_696/a_76_344# POR2X1_696/a_56_344#
+ POR2X1
XPOR2X1_685 VDD GND POR2X1_685/B POR2X1_685/A POR2X1_687/B POR2X1_685/m4_208_n4# POR2X1_685/O
+ POR2X1_685/CTRL2 POR2X1_685/a_16_28# POR2X1_685/CTRL POR2X1_685/a_76_344# POR2X1_685/a_56_344#
+ POR2X1
XPAND2X1_604 VDD GND POR2X1_750/B PAND2X1_72/A POR2X1_605/A PAND2X1_604/a_16_344#
+ PAND2X1_604/m4_208_n4# PAND2X1_604/O PAND2X1_604/a_56_28# PAND2X1_604/CTRL2 PAND2X1_604/CTRL
+ PAND2X1_604/a_76_28# PAND2X1
XPAND2X1_615 VDD GND POR2X1_614/Y PAND2X1_58/A POR2X1_623/B PAND2X1_615/a_16_344#
+ PAND2X1_615/m4_208_n4# PAND2X1_615/O PAND2X1_615/a_56_28# PAND2X1_615/CTRL2 PAND2X1_615/CTRL
+ PAND2X1_615/a_76_28# PAND2X1
XPAND2X1_637 VDD GND POR2X1_586/Y POR2X1_585/Y PAND2X1_638/B PAND2X1_637/a_16_344#
+ PAND2X1_637/m4_208_n4# PAND2X1_637/O PAND2X1_637/a_56_28# PAND2X1_637/CTRL2 PAND2X1_637/CTRL
+ PAND2X1_637/a_76_28# PAND2X1
XPAND2X1_626 VDD GND POR2X1_750/B PAND2X1_96/B POR2X1_629/B PAND2X1_626/a_16_344#
+ PAND2X1_626/m4_208_n4# PAND2X1_626/O PAND2X1_626/a_56_28# PAND2X1_626/CTRL2 PAND2X1_626/CTRL
+ PAND2X1_626/a_76_28# PAND2X1
XPAND2X1_659 VDD GND PAND2X1_659/B PAND2X1_659/A PAND2X1_659/Y PAND2X1_659/a_16_344#
+ PAND2X1_203/m4_208_n4# PAND2X1_659/O PAND2X1_659/a_56_28# PAND2X1_659/CTRL2 PAND2X1_659/CTRL
+ PAND2X1_659/a_76_28# PAND2X1
XPAND2X1_648 VDD GND PAND2X1_645/Y PAND2X1_644/Y PAND2X1_648/Y PAND2X1_648/a_16_344#
+ PAND2X1_648/m4_208_n4# PAND2X1_648/O PAND2X1_648/a_56_28# PAND2X1_648/CTRL2 PAND2X1_648/CTRL
+ PAND2X1_648/a_76_28# PAND2X1
XPOR2X1_471 VDD GND POR2X1_464/Y POR2X1_471/A POR2X1_477/A POR2X1_471/m4_208_n4# POR2X1_471/O
+ POR2X1_471/CTRL2 POR2X1_471/a_16_28# POR2X1_471/CTRL POR2X1_471/a_76_344# POR2X1_471/a_56_344#
+ POR2X1
XPOR2X1_460 VDD GND POR2X1_460/B POR2X1_460/A POR2X1_460/Y POR2X1_460/m4_208_n4# POR2X1_460/O
+ POR2X1_460/CTRL2 POR2X1_460/a_16_28# POR2X1_460/CTRL POR2X1_460/a_76_344# POR2X1_460/a_56_344#
+ POR2X1
XPOR2X1_493 VDD GND POR2X1_493/B POR2X1_493/A POR2X1_558/B POR2X1_493/m4_208_n4# POR2X1_493/O
+ POR2X1_493/CTRL2 POR2X1_493/a_16_28# POR2X1_493/CTRL POR2X1_493/a_76_344# POR2X1_493/a_56_344#
+ POR2X1
XPOR2X1_482 VDD GND POR2X1_7/A POR2X1_60/A POR2X1_482/Y POR2X1_482/m4_208_n4# POR2X1_482/O
+ POR2X1_482/CTRL2 POR2X1_482/a_16_28# POR2X1_482/CTRL POR2X1_482/a_76_344# POR2X1_482/a_56_344#
+ POR2X1
XPAND2X1_412 VDD GND PAND2X1_57/B PAND2X1_90/A POR2X1_634/A PAND2X1_412/a_16_344#
+ PAND2X1_412/m4_208_n4# PAND2X1_412/O PAND2X1_412/a_56_28# PAND2X1_412/CTRL2 PAND2X1_412/CTRL
+ PAND2X1_412/a_76_28# PAND2X1
XPAND2X1_401 VDD GND POR2X1_396/Y POR2X1_395/Y PAND2X1_402/B PAND2X1_401/a_16_344#
+ PAND2X1_401/m4_208_n4# PAND2X1_401/O PAND2X1_401/a_56_28# PAND2X1_401/CTRL2 PAND2X1_401/CTRL
+ PAND2X1_401/a_76_28# PAND2X1
XPAND2X1_434 VDD GND POR2X1_431/Y POR2X1_172/Y PAND2X1_436/A PAND2X1_434/a_16_344#
+ PAND2X1_434/m4_208_n4# PAND2X1_434/O PAND2X1_434/a_56_28# PAND2X1_434/CTRL2 PAND2X1_434/CTRL
+ PAND2X1_434/a_76_28# PAND2X1
XPAND2X1_423 VDD GND PAND2X1_65/B PAND2X1_6/Y POR2X1_832/B PAND2X1_423/a_16_344# PAND2X1_423/m4_208_n4#
+ PAND2X1_423/O PAND2X1_423/a_56_28# PAND2X1_423/CTRL2 PAND2X1_423/CTRL PAND2X1_423/a_76_28#
+ PAND2X1
XPAND2X1_445 VDD GND POR2X1_315/Y POR2X1_237/Y PAND2X1_445/Y PAND2X1_445/a_16_344#
+ PAND2X1_445/m4_208_n4# PAND2X1_445/O PAND2X1_445/a_56_28# PAND2X1_445/CTRL2 PAND2X1_445/CTRL
+ PAND2X1_445/a_76_28# PAND2X1
XPAND2X1_489 VDD GND POR2X1_488/Y POR2X1_487/Y PAND2X1_557/A PAND2X1_489/a_16_344#
+ PAND2X1_489/m4_208_n4# PAND2X1_489/O PAND2X1_489/a_56_28# PAND2X1_489/CTRL2 PAND2X1_489/CTRL
+ PAND2X1_489/a_76_28# PAND2X1
XPAND2X1_456 VDD GND PAND2X1_254/Y POR2X1_184/Y PAND2X1_465/B PAND2X1_456/a_16_344#
+ PAND2X1_456/m4_208_n4# PAND2X1_456/O PAND2X1_456/a_56_28# PAND2X1_456/CTRL2 PAND2X1_456/CTRL
+ PAND2X1_456/a_76_28# PAND2X1
XPAND2X1_478 VDD GND PAND2X1_478/B PAND2X1_469/Y PAND2X1_478/Y PAND2X1_478/a_16_344#
+ PAND2X1_478/m4_208_n4# PAND2X1_478/O PAND2X1_478/a_56_28# PAND2X1_478/CTRL2 PAND2X1_478/CTRL
+ PAND2X1_478/a_76_28# PAND2X1
XPAND2X1_467 VDD GND PAND2X1_467/B POR2X1_163/Y PAND2X1_467/Y PAND2X1_467/a_16_344#
+ PAND2X1_467/m4_208_n4# PAND2X1_467/O PAND2X1_467/a_56_28# PAND2X1_467/CTRL2 PAND2X1_467/CTRL
+ PAND2X1_467/a_76_28# PAND2X1
XPOR2X1_290 VDD GND POR2X1_16/A POR2X1_83/B POR2X1_290/Y POR2X1_290/m4_208_n4# POR2X1_290/O
+ POR2X1_290/CTRL2 POR2X1_290/a_16_28# POR2X1_290/CTRL POR2X1_290/a_76_344# POR2X1_290/a_56_344#
+ POR2X1
XPAND2X1_220 VDD GND PAND2X1_213/Y PAND2X1_220/A PAND2X1_220/Y PAND2X1_220/a_16_344#
+ PAND2X1_220/m4_208_n4# PAND2X1_220/O PAND2X1_220/a_56_28# PAND2X1_220/CTRL2 PAND2X1_220/CTRL
+ PAND2X1_220/a_76_28# PAND2X1
XPAND2X1_253 VDD GND POR2X1_614/A PAND2X1_65/B POR2X1_254/A PAND2X1_253/a_16_344#
+ PAND2X1_253/m4_208_n4# PAND2X1_253/O PAND2X1_253/a_56_28# PAND2X1_253/CTRL2 PAND2X1_253/CTRL
+ PAND2X1_253/a_76_28# PAND2X1
XPAND2X1_231 VDD GND POR2X1_230/Y POR2X1_229/Y PAND2X1_341/B PAND2X1_231/a_16_344#
+ PAND2X1_231/m4_208_n4# PAND2X1_231/O PAND2X1_231/a_56_28# PAND2X1_231/CTRL2 PAND2X1_231/CTRL
+ PAND2X1_231/a_76_28# PAND2X1
XPAND2X1_242 VDD GND PAND2X1_241/Y POR2X1_239/Y PAND2X1_242/Y PAND2X1_242/a_16_344#
+ PAND2X1_242/m4_208_n4# PAND2X1_242/O PAND2X1_242/a_56_28# PAND2X1_242/CTRL2 PAND2X1_242/CTRL
+ PAND2X1_242/a_76_28# PAND2X1
XPAND2X1_264 VDD GND POR2X1_77/Y POR2X1_41/B POR2X1_667/A PAND2X1_264/a_16_344# PAND2X1_264/m4_208_n4#
+ PAND2X1_264/O PAND2X1_264/a_56_28# PAND2X1_264/CTRL2 PAND2X1_264/CTRL PAND2X1_264/a_76_28#
+ PAND2X1
XPAND2X1_286 VDD GND PAND2X1_286/B POR2X1_283/Y PAND2X1_288/A PAND2X1_286/a_16_344#
+ PAND2X1_286/m4_208_n4# PAND2X1_286/O PAND2X1_286/a_56_28# PAND2X1_286/CTRL2 PAND2X1_286/CTRL
+ PAND2X1_286/a_76_28# PAND2X1
XPAND2X1_275 VDD GND POR2X1_274/Y D_INPUT_0 POR2X1_276/A PAND2X1_275/a_16_344# PAND2X1_275/m4_208_n4#
+ PAND2X1_275/O PAND2X1_275/a_56_28# PAND2X1_275/CTRL2 PAND2X1_275/CTRL PAND2X1_275/a_76_28#
+ PAND2X1
XPAND2X1_297 VDD GND POR2X1_296/Y PAND2X1_57/B POR2X1_347/B PAND2X1_297/a_16_344#
+ PAND2X1_297/m4_208_n4# PAND2X1_297/O PAND2X1_297/a_56_28# PAND2X1_297/CTRL2 PAND2X1_297/CTRL
+ PAND2X1_297/a_76_28# PAND2X1
XPOR2X1_801 VDD GND POR2X1_801/B POR2X1_801/A POR2X1_809/B POR2X1_801/m4_208_n4# POR2X1_801/O
+ POR2X1_801/CTRL2 POR2X1_801/a_16_28# POR2X1_801/CTRL POR2X1_801/a_76_344# POR2X1_801/a_56_344#
+ POR2X1
XPOR2X1_812 VDD GND POR2X1_812/B POR2X1_812/A D_GATE_811 POR2X1_812/m4_208_n4# POR2X1_812/O
+ POR2X1_812/CTRL2 POR2X1_812/a_16_28# POR2X1_812/CTRL POR2X1_812/a_76_344# POR2X1_812/a_56_344#
+ POR2X1
XPOR2X1_823 VDD GND POR2X1_52/A POR2X1_236/Y POR2X1_823/Y POR2X1_823/m4_208_n4# POR2X1_823/O
+ POR2X1_823/CTRL2 POR2X1_823/a_16_28# POR2X1_823/CTRL POR2X1_823/a_76_344# POR2X1_823/a_56_344#
+ POR2X1
XPOR2X1_845 VDD GND POR2X1_673/Y POR2X1_845/A POR2X1_849/A POR2X1_845/m4_208_n4# POR2X1_845/O
+ POR2X1_845/CTRL2 POR2X1_845/a_16_28# POR2X1_845/CTRL POR2X1_845/a_76_344# POR2X1_845/a_56_344#
+ POR2X1
XPOR2X1_834 VDD GND POR2X1_513/B POR2X1_678/A POR2X1_834/Y POR2X1_834/m4_208_n4# POR2X1_834/O
+ POR2X1_834/CTRL2 POR2X1_834/a_16_28# POR2X1_834/CTRL POR2X1_834/a_76_344# POR2X1_834/a_56_344#
+ POR2X1
XPOR2X1_856 VDD GND POR2X1_856/B POR2X1_855/Y POR2X1_863/B POR2X1_856/m4_208_n4# POR2X1_856/O
+ POR2X1_856/CTRL2 POR2X1_856/a_16_28# POR2X1_856/CTRL POR2X1_856/a_76_344# POR2X1_856/a_56_344#
+ POR2X1
XPAND2X1_808 VDD GND PAND2X1_808/B PAND2X1_803/Y PAND2X1_808/Y PAND2X1_808/a_16_344#
+ PAND2X1_808/m4_208_n4# PAND2X1_808/O PAND2X1_808/a_56_28# PAND2X1_808/CTRL2 PAND2X1_808/CTRL
+ PAND2X1_808/a_76_28# PAND2X1
XPAND2X1_819 VDD GND POR2X1_54/Y PAND2X1_48/B PAND2X1_820/B PAND2X1_819/a_16_344#
+ PAND2X1_819/m4_208_n4# PAND2X1_819/O PAND2X1_819/a_56_28# PAND2X1_819/CTRL2 PAND2X1_819/CTRL
+ PAND2X1_819/a_76_28# PAND2X1
XPOR2X1_119 VDD GND D_INPUT_1 POR2X1_14/Y POR2X1_119/Y POR2X1_236/m4_208_n4# POR2X1_119/O
+ POR2X1_119/CTRL2 POR2X1_119/a_16_28# POR2X1_119/CTRL POR2X1_119/a_76_344# POR2X1_119/a_56_344#
+ POR2X1
XPOR2X1_108 VDD GND POR2X1_60/A POR2X1_102/Y POR2X1_108/Y POR2X1_108/m4_208_n4# POR2X1_108/O
+ POR2X1_108/CTRL2 POR2X1_108/a_16_28# POR2X1_108/CTRL POR2X1_108/a_76_344# POR2X1_108/a_56_344#
+ POR2X1
XPAND2X1_62 VDD GND POR2X1_54/Y POR2X1_9/Y PAND2X1_63/B PAND2X1_62/a_16_344# PAND2X1_62/m4_208_n4#
+ PAND2X1_62/O PAND2X1_62/a_56_28# PAND2X1_62/CTRL2 PAND2X1_62/CTRL PAND2X1_62/a_76_28#
+ PAND2X1
XPAND2X1_40 VDD GND PAND2X1_59/B PAND2X1_3/B PAND2X1_41/B PAND2X1_40/a_16_344# PAND2X1_40/m4_208_n4#
+ PAND2X1_40/O PAND2X1_40/a_56_28# PAND2X1_40/CTRL2 PAND2X1_40/CTRL PAND2X1_40/a_76_28#
+ PAND2X1
XPAND2X1_51 VDD GND PAND2X1_95/B PAND2X1_47/B PAND2X1_52/B PAND2X1_51/a_16_344# PAND2X1_51/m4_208_n4#
+ PAND2X1_51/O PAND2X1_51/a_56_28# PAND2X1_51/CTRL2 PAND2X1_51/CTRL PAND2X1_51/a_76_28#
+ PAND2X1
XPAND2X1_73 VDD GND PAND2X1_90/A PAND2X1_9/Y PAND2X1_73/Y PAND2X1_73/a_16_344# PAND2X1_73/m4_208_n4#
+ PAND2X1_73/O PAND2X1_73/a_56_28# PAND2X1_73/CTRL2 PAND2X1_73/CTRL PAND2X1_73/a_76_28#
+ PAND2X1
XPAND2X1_84 VDD GND POR2X1_83/Y POR2X1_81/Y PAND2X1_84/Y PAND2X1_84/a_16_344# PAND2X1_84/m4_208_n4#
+ PAND2X1_84/O PAND2X1_84/a_56_28# PAND2X1_84/CTRL2 PAND2X1_84/CTRL PAND2X1_84/a_76_28#
+ PAND2X1
XPAND2X1_95 VDD GND PAND2X1_95/B PAND2X1_11/Y PAND2X1_96/B PAND2X1_95/a_16_344# PAND2X1_95/m4_208_n4#
+ PAND2X1_95/O PAND2X1_95/a_56_28# PAND2X1_95/CTRL2 PAND2X1_95/CTRL PAND2X1_95/a_76_28#
+ PAND2X1
XPOR2X1_15 VDD GND POR2X1_9/Y POR2X1_14/Y POR2X1_16/A POR2X1_15/m4_208_n4# POR2X1_15/O
+ POR2X1_15/CTRL2 POR2X1_15/a_16_28# POR2X1_15/CTRL POR2X1_15/a_76_344# POR2X1_15/a_56_344#
+ POR2X1
XPOR2X1_26 VDD GND POR2X1_22/A POR2X1_25/Y POR2X1_83/B POR2X1_26/m4_208_n4# POR2X1_26/O
+ POR2X1_26/CTRL2 POR2X1_26/a_16_28# POR2X1_26/CTRL POR2X1_26/a_76_344# POR2X1_26/a_56_344#
+ POR2X1
XPOR2X1_37 VDD GND D_INPUT_2 D_INPUT_3 POR2X1_37/Y POR2X1_37/m4_208_n4# POR2X1_37/O
+ POR2X1_37/CTRL2 POR2X1_37/a_16_28# POR2X1_37/CTRL POR2X1_37/a_76_344# POR2X1_37/a_56_344#
+ POR2X1
XPOR2X1_48 VDD GND POR2X1_46/Y POR2X1_48/A POR2X1_48/Y POR2X1_48/m4_208_n4# POR2X1_48/O
+ POR2X1_48/CTRL2 POR2X1_48/a_16_28# POR2X1_48/CTRL POR2X1_48/a_76_344# POR2X1_48/a_56_344#
+ POR2X1
XPOR2X1_620 VDD GND POR2X1_620/B POR2X1_620/A POR2X1_623/A POR2X1_620/m4_208_n4# POR2X1_620/O
+ POR2X1_620/CTRL2 POR2X1_620/a_16_28# POR2X1_620/CTRL POR2X1_620/a_76_344# POR2X1_620/a_56_344#
+ POR2X1
XPOR2X1_59 VDD GND POR2X1_12/A POR2X1_25/Y POR2X1_60/A POR2X1_59/m4_208_n4# POR2X1_59/O
+ POR2X1_59/CTRL2 POR2X1_59/a_16_28# POR2X1_59/CTRL POR2X1_59/a_76_344# POR2X1_59/a_56_344#
+ POR2X1
XPOR2X1_631 VDD GND POR2X1_631/B POR2X1_631/A POR2X1_632/A POR2X1_631/m4_208_n4# POR2X1_631/O
+ POR2X1_631/CTRL2 POR2X1_631/a_16_28# POR2X1_631/CTRL POR2X1_631/a_76_344# POR2X1_631/a_56_344#
+ POR2X1
XPOR2X1_653 VDD GND POR2X1_653/B POR2X1_652/Y POR2X1_661/B POR2X1_653/m4_208_n4# POR2X1_653/O
+ POR2X1_653/CTRL2 POR2X1_653/a_16_28# POR2X1_653/CTRL POR2X1_653/a_76_344# POR2X1_653/a_56_344#
+ POR2X1
XPOR2X1_642 VDD GND POR2X1_462/B POR2X1_559/A POR2X1_649/B POR2X1_642/m4_208_n4# POR2X1_642/O
+ POR2X1_642/CTRL2 POR2X1_642/a_16_28# POR2X1_642/CTRL POR2X1_642/a_76_344# POR2X1_642/a_56_344#
+ POR2X1
XPOR2X1_686 VDD GND POR2X1_686/B POR2X1_686/A POR2X1_687/A POR2X1_686/m4_208_n4# POR2X1_686/O
+ POR2X1_686/CTRL2 POR2X1_686/a_16_28# POR2X1_686/CTRL POR2X1_686/a_76_344# POR2X1_686/a_56_344#
+ POR2X1
XPOR2X1_664 VDD GND PAND2X1_73/Y POR2X1_78/A POR2X1_664/Y POR2X1_664/m4_208_n4# POR2X1_664/O
+ POR2X1_664/CTRL2 POR2X1_664/a_16_28# POR2X1_664/CTRL POR2X1_664/a_76_344# POR2X1_664/a_56_344#
+ POR2X1
XPOR2X1_675 VDD GND POR2X1_439/Y POR2X1_675/A POR2X1_675/Y POR2X1_675/m4_208_n4# POR2X1_675/O
+ POR2X1_675/CTRL2 POR2X1_675/a_16_28# POR2X1_675/CTRL POR2X1_675/a_76_344# POR2X1_675/a_56_344#
+ POR2X1
XPOR2X1_697 VDD GND POR2X1_416/B POR2X1_236/Y POR2X1_697/Y POR2X1_697/m4_208_n4# POR2X1_697/O
+ POR2X1_697/CTRL2 POR2X1_697/a_16_28# POR2X1_697/CTRL POR2X1_697/a_76_344# POR2X1_697/a_56_344#
+ POR2X1
XPAND2X1_638 VDD GND PAND2X1_638/B POR2X1_588/Y PAND2X1_651/A PAND2X1_638/a_16_344#
+ PAND2X1_638/m4_208_n4# PAND2X1_638/O PAND2X1_638/a_56_28# PAND2X1_638/CTRL2 PAND2X1_638/CTRL
+ PAND2X1_638/a_76_28# PAND2X1
XPAND2X1_605 VDD GND POR2X1_604/Y POR2X1_603/Y PAND2X1_645/B PAND2X1_605/a_16_344#
+ PAND2X1_605/m4_208_n4# PAND2X1_605/O PAND2X1_605/a_56_28# PAND2X1_605/CTRL2 PAND2X1_605/CTRL
+ PAND2X1_605/a_76_28# PAND2X1
XPAND2X1_616 VDD GND POR2X1_814/B PAND2X1_20/A POR2X1_621/B PAND2X1_616/a_16_344#
+ PAND2X1_616/m4_208_n4# PAND2X1_616/O PAND2X1_616/a_56_28# PAND2X1_616/CTRL2 PAND2X1_616/CTRL
+ PAND2X1_616/a_76_28# PAND2X1
XPAND2X1_627 VDD GND PAND2X1_69/A PAND2X1_6/Y POR2X1_629/A PAND2X1_627/a_16_344# PAND2X1_627/m4_208_n4#
+ PAND2X1_627/O PAND2X1_627/a_56_28# PAND2X1_627/CTRL2 PAND2X1_627/CTRL PAND2X1_627/a_76_28#
+ PAND2X1
XPAND2X1_649 VDD GND PAND2X1_643/Y PAND2X1_649/A PAND2X1_655/B PAND2X1_649/a_16_344#
+ PAND2X1_649/m4_208_n4# PAND2X1_649/O PAND2X1_649/a_56_28# PAND2X1_649/CTRL2 PAND2X1_649/CTRL
+ PAND2X1_649/a_76_28# PAND2X1
XPOR2X1_450 VDD GND POR2X1_450/B POR2X1_450/A POR2X1_450/Y POR2X1_450/m4_208_n4# POR2X1_450/O
+ POR2X1_450/CTRL2 POR2X1_450/a_16_28# POR2X1_450/CTRL POR2X1_450/a_76_344# POR2X1_450/a_56_344#
+ POR2X1
XPOR2X1_461 VDD GND POR2X1_461/B POR2X1_461/A POR2X1_461/Y POR2X1_461/m4_208_n4# POR2X1_461/O
+ POR2X1_461/CTRL2 POR2X1_461/a_16_28# POR2X1_461/CTRL POR2X1_461/a_76_344# POR2X1_461/a_56_344#
+ POR2X1
XPOR2X1_483 VDD GND POR2X1_483/B POR2X1_483/A POR2X1_631/B POR2X1_483/m4_208_n4# POR2X1_483/O
+ POR2X1_483/CTRL2 POR2X1_483/a_16_28# POR2X1_483/CTRL POR2X1_483/a_76_344# POR2X1_483/a_56_344#
+ POR2X1
XPOR2X1_494 VDD GND POR2X1_13/A POR2X1_384/A POR2X1_494/Y POR2X1_494/m4_208_n4# POR2X1_494/O
+ POR2X1_494/CTRL2 POR2X1_494/a_16_28# POR2X1_494/CTRL POR2X1_494/a_76_344# POR2X1_494/a_56_344#
+ POR2X1
XPOR2X1_472 VDD GND POR2X1_472/B POR2X1_463/Y POR2X1_472/Y POR2X1_472/m4_208_n4# POR2X1_472/O
+ POR2X1_472/CTRL2 POR2X1_472/a_16_28# POR2X1_472/CTRL POR2X1_472/a_76_344# POR2X1_472/a_56_344#
+ POR2X1
XPAND2X1_413 VDD GND POR2X1_634/A INPUT_0 POR2X1_461/A PAND2X1_413/a_16_344# PAND2X1_413/m4_208_n4#
+ PAND2X1_413/O PAND2X1_413/a_56_28# PAND2X1_413/CTRL2 PAND2X1_413/CTRL PAND2X1_413/a_76_28#
+ PAND2X1
XPAND2X1_402 VDD GND PAND2X1_402/B POR2X1_397/Y PAND2X1_404/A PAND2X1_402/a_16_344#
+ PAND2X1_402/m4_208_n4# PAND2X1_402/O PAND2X1_402/a_56_28# PAND2X1_402/CTRL2 PAND2X1_402/CTRL
+ PAND2X1_402/a_76_28# PAND2X1
XPAND2X1_435 VDD GND POR2X1_433/Y POR2X1_432/Y PAND2X1_435/Y PAND2X1_435/a_16_344#
+ PAND2X1_435/m4_208_n4# PAND2X1_435/O PAND2X1_435/a_56_28# PAND2X1_435/CTRL2 PAND2X1_435/CTRL
+ PAND2X1_435/a_76_28# PAND2X1
XPAND2X1_424 VDD GND POR2X1_78/A PAND2X1_57/B POR2X1_449/A PAND2X1_424/a_16_344# POR2X1_592/m4_208_n4#
+ PAND2X1_424/O PAND2X1_424/a_56_28# PAND2X1_424/CTRL2 PAND2X1_424/CTRL PAND2X1_424/a_76_28#
+ PAND2X1
XPAND2X1_446 VDD GND POR2X1_418/Y POR2X1_417/Y PAND2X1_446/Y PAND2X1_446/a_16_344#
+ PAND2X1_446/m4_208_n4# PAND2X1_446/O PAND2X1_446/a_56_28# PAND2X1_446/CTRL2 PAND2X1_446/CTRL
+ PAND2X1_446/a_76_28# PAND2X1
XPAND2X1_479 VDD GND PAND2X1_479/B PAND2X1_479/A PAND2X1_480/B PAND2X1_479/a_16_344#
+ PAND2X1_479/m4_208_n4# PAND2X1_479/O PAND2X1_479/a_56_28# PAND2X1_479/CTRL2 PAND2X1_479/CTRL
+ PAND2X1_479/a_76_28# PAND2X1
XPAND2X1_468 VDD GND PAND2X1_652/A PAND2X1_798/B PAND2X1_469/B PAND2X1_468/a_16_344#
+ PAND2X1_468/m4_208_n4# PAND2X1_468/O PAND2X1_468/a_56_28# PAND2X1_468/CTRL2 PAND2X1_468/CTRL
+ PAND2X1_468/a_76_28# PAND2X1
XPAND2X1_457 VDD GND PAND2X1_787/A POR2X1_368/Y PAND2X1_457/Y PAND2X1_457/a_16_344#
+ PAND2X1_457/m4_208_n4# PAND2X1_457/O PAND2X1_457/a_56_28# PAND2X1_457/CTRL2 PAND2X1_457/CTRL
+ PAND2X1_457/a_76_28# PAND2X1
XPOR2X1_280 VDD GND POR2X1_48/A POR2X1_236/Y POR2X1_280/Y POR2X1_280/m4_208_n4# POR2X1_280/O
+ POR2X1_280/CTRL2 POR2X1_280/a_16_28# POR2X1_280/CTRL POR2X1_280/a_76_344# POR2X1_280/a_56_344#
+ POR2X1
XPOR2X1_291 VDD GND POR2X1_39/B POR2X1_234/A POR2X1_291/Y POR2X1_291/m4_208_n4# POR2X1_291/O
+ POR2X1_291/CTRL2 POR2X1_291/a_16_28# POR2X1_291/CTRL POR2X1_291/a_76_344# POR2X1_291/a_56_344#
+ POR2X1
XPAND2X1_221 VDD GND PAND2X1_220/Y PAND2X1_192/Y PAND2X1_221/Y PAND2X1_221/a_16_344#
+ PAND2X1_221/m4_208_n4# PAND2X1_221/O PAND2X1_221/a_56_28# PAND2X1_221/CTRL2 PAND2X1_221/CTRL
+ PAND2X1_221/a_76_28# PAND2X1
XPAND2X1_210 VDD GND POR2X1_163/Y POR2X1_158/Y PAND2X1_213/B PAND2X1_210/a_16_344#
+ PAND2X1_210/m4_208_n4# PAND2X1_210/O PAND2X1_210/a_56_28# PAND2X1_210/CTRL2 PAND2X1_210/CTRL
+ PAND2X1_210/a_76_28# PAND2X1
XPAND2X1_254 VDD GND POR2X1_253/Y POR2X1_252/Y PAND2X1_254/Y PAND2X1_254/a_16_344#
+ PAND2X1_254/m4_208_n4# PAND2X1_254/O PAND2X1_254/a_56_28# PAND2X1_254/CTRL2 PAND2X1_254/CTRL
+ PAND2X1_254/a_76_28# PAND2X1
XPAND2X1_243 VDD GND PAND2X1_243/B POR2X1_235/Y PAND2X1_244/B PAND2X1_243/a_16_344#
+ POR2X1_230/m4_208_n4# PAND2X1_243/O PAND2X1_243/a_56_28# PAND2X1_243/CTRL2 PAND2X1_243/CTRL
+ PAND2X1_243/a_76_28# PAND2X1
XPAND2X1_232 VDD GND POR2X1_260/A POR2X1_78/B POR2X1_240/B PAND2X1_232/a_16_344# PAND2X1_232/m4_208_n4#
+ PAND2X1_232/O PAND2X1_232/a_56_28# PAND2X1_232/CTRL2 PAND2X1_232/CTRL PAND2X1_232/a_76_28#
+ PAND2X1
XPAND2X1_265 VDD GND POR2X1_264/Y PAND2X1_41/B POR2X1_267/B PAND2X1_265/a_16_344#
+ PAND2X1_265/m4_208_n4# PAND2X1_265/O PAND2X1_265/a_56_28# PAND2X1_265/CTRL2 PAND2X1_265/CTRL
+ PAND2X1_265/a_76_28# PAND2X1
XPAND2X1_276 VDD GND POR2X1_275/Y POR2X1_271/Y PAND2X1_473/B PAND2X1_276/a_16_344#
+ PAND2X1_276/m4_208_n4# PAND2X1_276/O PAND2X1_276/a_56_28# PAND2X1_276/CTRL2 PAND2X1_276/CTRL
+ PAND2X1_276/a_76_28# PAND2X1
XPAND2X1_287 VDD GND PAND2X1_284/Y POR2X1_278/Y PAND2X1_287/Y PAND2X1_287/a_16_344#
+ PAND2X1_287/m4_208_n4# PAND2X1_287/O PAND2X1_287/a_56_28# PAND2X1_287/CTRL2 PAND2X1_287/CTRL
+ PAND2X1_287/a_76_28# PAND2X1
XPAND2X1_298 VDD GND PAND2X1_55/Y PAND2X1_32/B POR2X1_302/B PAND2X1_298/a_16_344#
+ PAND2X1_298/m4_208_n4# PAND2X1_298/O PAND2X1_298/a_56_28# PAND2X1_298/CTRL2 PAND2X1_298/CTRL
+ PAND2X1_298/a_76_28# PAND2X1
XPOR2X1_802 VDD GND POR2X1_802/B POR2X1_802/A POR2X1_809/A POR2X1_802/m4_208_n4# POR2X1_802/O
+ POR2X1_802/CTRL2 POR2X1_802/a_16_28# POR2X1_802/CTRL POR2X1_802/a_76_344# POR2X1_802/a_56_344#
+ POR2X1
XPOR2X1_824 VDD GND POR2X1_83/B POR2X1_234/A POR2X1_824/Y POR2X1_824/m4_208_n4# POR2X1_824/O
+ POR2X1_824/CTRL2 POR2X1_824/a_16_28# POR2X1_824/CTRL POR2X1_824/a_76_344# POR2X1_824/a_56_344#
+ POR2X1
XPOR2X1_835 VDD GND POR2X1_835/B POR2X1_835/A POR2X1_835/Y POR2X1_835/m4_208_n4# POR2X1_835/O
+ POR2X1_835/CTRL2 POR2X1_835/a_16_28# POR2X1_835/CTRL POR2X1_835/a_76_344# POR2X1_835/a_56_344#
+ POR2X1
XPOR2X1_813 VDD GND PAND2X1_63/B POR2X1_263/Y POR2X1_813/Y POR2X1_813/m4_208_n4# POR2X1_813/O
+ POR2X1_813/CTRL2 POR2X1_813/a_16_28# POR2X1_813/CTRL POR2X1_813/a_76_344# POR2X1_813/a_56_344#
+ POR2X1
XPOR2X1_857 VDD GND POR2X1_857/B POR2X1_857/A POR2X1_863/A POR2X1_857/m4_208_n4# POR2X1_857/O
+ POR2X1_857/CTRL2 POR2X1_857/a_16_28# POR2X1_857/CTRL POR2X1_857/a_76_344# POR2X1_857/a_56_344#
+ POR2X1
XPOR2X1_846 VDD GND POR2X1_846/B POR2X1_846/A POR2X1_846/Y POR2X1_846/m4_208_n4# POR2X1_846/O
+ POR2X1_846/CTRL2 POR2X1_846/a_16_28# POR2X1_846/CTRL POR2X1_846/a_76_344# POR2X1_846/a_56_344#
+ POR2X1
XPAND2X1_809 VDD GND PAND2X1_809/B PAND2X1_809/A PAND2X1_810/B PAND2X1_809/a_16_344#
+ PAND2X1_809/m4_208_n4# PAND2X1_809/O PAND2X1_809/a_56_28# PAND2X1_809/CTRL2 PAND2X1_809/CTRL
+ PAND2X1_809/a_76_28# PAND2X1
XPOR2X1_109 VDD GND POR2X1_32/A POR2X1_77/Y POR2X1_109/Y POR2X1_109/m4_208_n4# POR2X1_109/O
+ POR2X1_109/CTRL2 POR2X1_109/a_16_28# POR2X1_109/CTRL POR2X1_109/a_76_344# POR2X1_109/a_56_344#
+ POR2X1
XPAND2X1_30 VDD GND INPUT_5 INPUT_4 PAND2X1_47/B PAND2X1_30/a_16_344# PAND2X1_30/m4_208_n4#
+ PAND2X1_30/O PAND2X1_30/a_56_28# PAND2X1_30/CTRL2 PAND2X1_30/CTRL PAND2X1_30/a_76_28#
+ PAND2X1
XPAND2X1_52 VDD GND PAND2X1_52/B POR2X1_68/A PAND2X1_52/Y PAND2X1_52/a_16_344# PAND2X1_52/m4_208_n4#
+ PAND2X1_52/O PAND2X1_52/a_56_28# PAND2X1_52/CTRL2 PAND2X1_52/CTRL PAND2X1_52/a_76_28#
+ PAND2X1
XPAND2X1_41 VDD GND PAND2X1_41/B POR2X1_294/B PAND2X1_41/Y PAND2X1_41/a_16_344# PAND2X1_41/m4_208_n4#
+ PAND2X1_41/O PAND2X1_41/a_56_28# PAND2X1_41/CTRL2 PAND2X1_41/CTRL PAND2X1_41/a_76_28#
+ PAND2X1
XPAND2X1_63 VDD GND PAND2X1_63/B PAND2X1_8/Y PAND2X1_63/Y PAND2X1_63/a_16_344# PAND2X1_63/m4_208_n4#
+ PAND2X1_63/O PAND2X1_63/a_56_28# PAND2X1_63/CTRL2 PAND2X1_63/CTRL PAND2X1_63/a_76_28#
+ PAND2X1
XPAND2X1_74 VDD GND PAND2X1_73/Y PAND2X1_32/B POR2X1_76/B PAND2X1_74/a_16_344# PAND2X1_74/m4_208_n4#
+ PAND2X1_74/O PAND2X1_74/a_56_28# PAND2X1_74/CTRL2 PAND2X1_74/CTRL PAND2X1_74/a_76_28#
+ PAND2X1
XPOR2X1_16 VDD GND POR2X1_7/B POR2X1_16/A POR2X1_16/Y POR2X1_16/m4_208_n4# POR2X1_16/O
+ POR2X1_16/CTRL2 POR2X1_16/a_16_28# POR2X1_16/CTRL POR2X1_16/a_76_344# POR2X1_16/a_56_344#
+ POR2X1
XPAND2X1_85 VDD GND PAND2X1_90/A PAND2X1_20/A PAND2X1_85/Y PAND2X1_85/a_16_344# PAND2X1_85/m4_208_n4#
+ PAND2X1_85/O PAND2X1_85/a_56_28# PAND2X1_85/CTRL2 PAND2X1_85/CTRL PAND2X1_85/a_76_28#
+ PAND2X1
XPOR2X1_38 VDD GND POR2X1_38/B POR2X1_37/Y POR2X1_38/Y POR2X1_38/m4_208_n4# POR2X1_38/O
+ POR2X1_38/CTRL2 POR2X1_38/a_16_28# POR2X1_38/CTRL POR2X1_38/a_76_344# POR2X1_38/a_56_344#
+ POR2X1
XPOR2X1_49 VDD GND POR2X1_14/Y POR2X1_38/B POR2X1_49/Y POR2X1_49/m4_208_n4# POR2X1_49/O
+ POR2X1_49/CTRL2 POR2X1_49/a_16_28# POR2X1_49/CTRL POR2X1_49/a_76_344# POR2X1_49/a_56_344#
+ POR2X1
XPOR2X1_27 VDD GND POR2X1_7/A POR2X1_83/B POR2X1_27/Y POR2X1_27/m4_208_n4# POR2X1_27/O
+ POR2X1_27/CTRL2 POR2X1_27/a_16_28# POR2X1_27/CTRL POR2X1_27/a_76_344# POR2X1_27/a_56_344#
+ POR2X1
XPOR2X1_610 VDD GND PAND2X1_41/B PAND2X1_48/B POR2X1_610/Y POR2X1_610/m4_208_n4# POR2X1_610/O
+ POR2X1_610/CTRL2 POR2X1_610/a_16_28# POR2X1_610/CTRL POR2X1_610/a_76_344# POR2X1_610/a_56_344#
+ POR2X1
XPAND2X1_96 VDD GND PAND2X1_96/B PAND2X1_94/Y POR2X1_98/A PAND2X1_96/a_16_344# PAND2X1_96/m4_208_n4#
+ PAND2X1_96/O PAND2X1_96/a_56_28# PAND2X1_96/CTRL2 PAND2X1_96/CTRL PAND2X1_96/a_76_28#
+ PAND2X1
XPOR2X1_621 VDD GND POR2X1_621/B POR2X1_621/A POR2X1_622/A POR2X1_621/m4_208_n4# POR2X1_621/O
+ POR2X1_621/CTRL2 POR2X1_621/a_16_28# POR2X1_621/CTRL POR2X1_621/a_76_344# POR2X1_621/a_56_344#
+ POR2X1
XPOR2X1_632 VDD GND POR2X1_632/B POR2X1_632/A POR2X1_632/Y POR2X1_632/m4_208_n4# POR2X1_632/O
+ POR2X1_632/CTRL2 POR2X1_632/a_16_28# POR2X1_632/CTRL POR2X1_632/a_76_344# POR2X1_632/a_56_344#
+ POR2X1
XPOR2X1_654 VDD GND POR2X1_654/B POR2X1_651/Y POR2X1_661/A POR2X1_654/m4_208_n4# POR2X1_654/O
+ POR2X1_654/CTRL2 POR2X1_654/a_16_28# POR2X1_654/CTRL POR2X1_654/a_76_344# POR2X1_654/a_56_344#
+ POR2X1
XPOR2X1_643 VDD GND POR2X1_537/Y POR2X1_643/A POR2X1_643/Y POR2X1_643/m4_208_n4# POR2X1_643/O
+ POR2X1_643/CTRL2 POR2X1_643/a_16_28# POR2X1_643/CTRL POR2X1_643/a_76_344# POR2X1_643/a_56_344#
+ POR2X1
XPOR2X1_665 VDD GND POR2X1_7/B POR2X1_665/A POR2X1_665/Y POR2X1_665/m4_208_n4# POR2X1_665/O
+ POR2X1_665/CTRL2 POR2X1_665/a_16_28# POR2X1_665/CTRL POR2X1_665/a_76_344# POR2X1_665/a_56_344#
+ POR2X1
XPOR2X1_676 VDD GND POR2X1_614/A POR2X1_828/A POR2X1_676/Y POR2X1_676/m4_208_n4# POR2X1_676/O
+ POR2X1_676/CTRL2 POR2X1_676/a_16_28# POR2X1_676/CTRL POR2X1_676/a_76_344# POR2X1_676/a_56_344#
+ POR2X1
XPOR2X1_687 VDD GND POR2X1_687/B POR2X1_687/A POR2X1_687/Y POR2X1_687/m4_208_n4# POR2X1_687/O
+ POR2X1_687/CTRL2 POR2X1_687/a_16_28# POR2X1_687/CTRL POR2X1_687/a_76_344# POR2X1_687/a_56_344#
+ POR2X1
XPOR2X1_698 VDD GND POR2X1_65/A POR2X1_394/A POR2X1_698/Y POR2X1_698/m4_208_n4# POR2X1_698/O
+ POR2X1_698/CTRL2 POR2X1_698/a_16_28# POR2X1_698/CTRL POR2X1_698/a_76_344# POR2X1_698/a_56_344#
+ POR2X1
XPAND2X1_628 VDD GND PAND2X1_93/B PAND2X1_48/B POR2X1_630/B PAND2X1_628/a_16_344#
+ PAND2X1_628/m4_208_n4# PAND2X1_628/O PAND2X1_628/a_56_28# PAND2X1_628/CTRL2 PAND2X1_628/CTRL
+ PAND2X1_628/a_76_28# PAND2X1
XPAND2X1_617 VDD GND PAND2X1_52/B PAND2X1_39/B POR2X1_621/A PAND2X1_617/a_16_344#
+ PAND2X1_617/m4_208_n4# PAND2X1_617/O PAND2X1_617/a_56_28# PAND2X1_617/CTRL2 PAND2X1_617/CTRL
+ PAND2X1_617/a_76_28# PAND2X1
XPAND2X1_606 VDD GND POR2X1_119/Y POR2X1_102/Y POR2X1_607/A PAND2X1_606/a_16_344#
+ PAND2X1_606/m4_208_n4# PAND2X1_606/O PAND2X1_606/a_56_28# PAND2X1_606/CTRL2 PAND2X1_606/CTRL
+ PAND2X1_606/a_76_28# PAND2X1
XPAND2X1_639 VDD GND PAND2X1_639/B PAND2X1_635/Y PAND2X1_639/Y PAND2X1_639/a_16_344#
+ PAND2X1_639/m4_208_n4# PAND2X1_639/O PAND2X1_639/a_56_28# PAND2X1_639/CTRL2 PAND2X1_639/CTRL
+ PAND2X1_639/a_76_28# PAND2X1
XPOR2X1_451 VDD GND POR2X1_635/B POR2X1_451/A POR2X1_452/A POR2X1_451/m4_208_n4# POR2X1_451/O
+ POR2X1_451/CTRL2 POR2X1_451/a_16_28# POR2X1_451/CTRL POR2X1_451/a_76_344# POR2X1_451/a_56_344#
+ POR2X1
XPOR2X1_440 VDD GND POR2X1_440/B POR2X1_439/Y POR2X1_440/Y POR2X1_440/m4_208_n4# POR2X1_440/O
+ POR2X1_440/CTRL2 POR2X1_440/a_16_28# POR2X1_440/CTRL POR2X1_440/a_76_344# POR2X1_440/a_56_344#
+ POR2X1
XPOR2X1_462 VDD GND POR2X1_462/B POR2X1_461/Y POR2X1_472/B POR2X1_462/m4_208_n4# POR2X1_462/O
+ POR2X1_462/CTRL2 POR2X1_462/a_16_28# POR2X1_462/CTRL POR2X1_462/a_76_344# POR2X1_462/a_56_344#
+ POR2X1
XPOR2X1_473 VDD GND POR2X1_116/Y POR2X1_276/Y POR2X1_476/A POR2X1_473/m4_208_n4# POR2X1_473/O
+ POR2X1_473/CTRL2 POR2X1_473/a_16_28# POR2X1_473/CTRL POR2X1_473/a_76_344# POR2X1_473/a_56_344#
+ POR2X1
XPOR2X1_484 VDD GND POR2X1_41/B POR2X1_39/B POR2X1_484/Y POR2X1_484/m4_208_n4# POR2X1_484/O
+ POR2X1_484/CTRL2 POR2X1_484/a_16_28# POR2X1_484/CTRL POR2X1_484/a_76_344# POR2X1_484/a_56_344#
+ POR2X1
XPOR2X1_495 VDD GND POR2X1_39/B POR2X1_55/Y POR2X1_495/Y POR2X1_495/m4_208_n4# POR2X1_495/O
+ POR2X1_495/CTRL2 POR2X1_495/a_16_28# POR2X1_495/CTRL POR2X1_495/a_76_344# POR2X1_495/a_56_344#
+ POR2X1
XPAND2X1_403 VDD GND PAND2X1_403/B POR2X1_399/Y PAND2X1_403/Y PAND2X1_403/a_16_344#
+ PAND2X1_403/m4_208_n4# PAND2X1_403/O PAND2X1_403/a_56_28# PAND2X1_403/CTRL2 PAND2X1_403/CTRL
+ PAND2X1_403/a_76_28# PAND2X1
XPAND2X1_414 VDD GND PAND2X1_6/A INPUT_3 POR2X1_415/A PAND2X1_414/a_16_344# PAND2X1_414/m4_208_n4#
+ PAND2X1_414/O PAND2X1_414/a_56_28# PAND2X1_414/CTRL2 PAND2X1_414/CTRL PAND2X1_414/a_76_28#
+ PAND2X1
XPAND2X1_436 VDD GND PAND2X1_435/Y PAND2X1_436/A PAND2X1_798/B PAND2X1_436/a_16_344#
+ PAND2X1_436/m4_208_n4# PAND2X1_436/O PAND2X1_436/a_56_28# PAND2X1_436/CTRL2 PAND2X1_436/CTRL
+ PAND2X1_436/a_76_28# PAND2X1
XPAND2X1_425 VDD GND PAND2X1_18/B D_INPUT_5 PAND2X1_425/Y PAND2X1_425/a_16_344# PAND2X1_425/m4_208_n4#
+ PAND2X1_425/O PAND2X1_425/a_56_28# PAND2X1_425/CTRL2 PAND2X1_425/CTRL PAND2X1_425/a_76_28#
+ PAND2X1
XPAND2X1_458 VDD GND PAND2X1_717/A POR2X1_372/Y PAND2X1_464/B PAND2X1_458/a_16_344#
+ PAND2X1_458/m4_208_n4# PAND2X1_458/O PAND2X1_458/a_56_28# PAND2X1_458/CTRL2 PAND2X1_458/CTRL
+ PAND2X1_458/a_76_28# PAND2X1
XPAND2X1_447 VDD GND POR2X1_420/Y POR2X1_419/Y PAND2X1_454/B PAND2X1_447/a_16_344#
+ PAND2X1_447/m4_208_n4# PAND2X1_447/O PAND2X1_447/a_56_28# PAND2X1_447/CTRL2 PAND2X1_447/CTRL
+ PAND2X1_447/a_76_28# PAND2X1
XPAND2X1_469 VDD GND PAND2X1_469/B PAND2X1_444/Y PAND2X1_469/Y PAND2X1_469/a_16_344#
+ PAND2X1_469/m4_208_n4# PAND2X1_469/O PAND2X1_469/a_56_28# PAND2X1_469/CTRL2 PAND2X1_469/CTRL
+ PAND2X1_469/a_76_28# PAND2X1
XPOR2X1_270 VDD GND PAND2X1_20/A PAND2X1_69/A POR2X1_270/Y POR2X1_270/m4_208_n4# POR2X1_270/O
+ POR2X1_270/CTRL2 POR2X1_270/a_16_28# POR2X1_270/CTRL POR2X1_270/a_76_344# POR2X1_270/a_56_344#
+ POR2X1
XPOR2X1_281 VDD GND POR2X1_7/B POR2X1_236/Y POR2X1_281/Y POR2X1_281/m4_208_n4# POR2X1_281/O
+ POR2X1_281/CTRL2 POR2X1_281/a_16_28# POR2X1_281/CTRL POR2X1_281/a_76_344# POR2X1_281/a_56_344#
+ POR2X1
XPOR2X1_292 VDD GND POR2X1_40/Y POR2X1_150/Y POR2X1_292/Y POR2X1_295/m4_208_n4# POR2X1_292/O
+ POR2X1_292/CTRL2 POR2X1_292/a_16_28# POR2X1_292/CTRL POR2X1_292/a_76_344# POR2X1_292/a_56_344#
+ POR2X1
XPAND2X1_211 VDD GND PAND2X1_853/B PAND2X1_211/A PAND2X1_212/B PAND2X1_211/a_16_344#
+ PAND2X1_211/m4_208_n4# PAND2X1_211/O PAND2X1_211/a_56_28# PAND2X1_211/CTRL2 PAND2X1_211/CTRL
+ PAND2X1_211/a_76_28# PAND2X1
XPAND2X1_200 VDD GND PAND2X1_200/B PAND2X1_193/Y PAND2X1_200/Y PAND2X1_200/a_16_344#
+ PAND2X1_200/m4_208_n4# PAND2X1_200/O PAND2X1_200/a_56_28# PAND2X1_200/CTRL2 PAND2X1_200/CTRL
+ PAND2X1_200/a_76_28# PAND2X1
XPAND2X1_255 VDD GND POR2X1_260/A PAND2X1_90/A POR2X1_541/B PAND2X1_255/a_16_344#
+ PAND2X1_255/m4_208_n4# PAND2X1_255/O PAND2X1_255/a_56_28# PAND2X1_255/CTRL2 PAND2X1_255/CTRL
+ PAND2X1_255/a_76_28# PAND2X1
XPAND2X1_222 VDD GND PAND2X1_222/B PAND2X1_222/A PAND2X1_223/B PAND2X1_222/a_16_344#
+ PAND2X1_799/m4_208_n4# PAND2X1_222/O PAND2X1_222/a_56_28# PAND2X1_222/CTRL2 PAND2X1_222/CTRL
+ PAND2X1_222/a_76_28# PAND2X1
XPAND2X1_244 VDD GND PAND2X1_244/B PAND2X1_242/Y PAND2X1_860/A PAND2X1_244/a_16_344#
+ PAND2X1_244/m4_208_n4# PAND2X1_244/O PAND2X1_244/a_56_28# PAND2X1_244/CTRL2 PAND2X1_244/CTRL
+ PAND2X1_244/a_76_28# PAND2X1
XPAND2X1_233 VDD GND PAND2X1_94/A INPUT_0 PAND2X1_824/B PAND2X1_233/a_16_344# PAND2X1_233/m4_208_n4#
+ PAND2X1_233/O PAND2X1_233/a_56_28# PAND2X1_233/CTRL2 PAND2X1_233/CTRL PAND2X1_233/a_76_28#
+ PAND2X1
XPAND2X1_266 VDD GND POR2X1_263/Y POR2X1_262/Y PAND2X1_267/B PAND2X1_266/a_16_344#
+ PAND2X1_716/m4_208_n4# PAND2X1_266/O PAND2X1_266/a_56_28# PAND2X1_266/CTRL2 PAND2X1_266/CTRL
+ PAND2X1_266/a_76_28# PAND2X1
XPAND2X1_288 VDD GND PAND2X1_287/Y PAND2X1_288/A PAND2X1_362/A PAND2X1_288/a_16_344#
+ PAND2X1_288/m4_208_n4# PAND2X1_288/O PAND2X1_288/a_56_28# PAND2X1_288/CTRL2 PAND2X1_288/CTRL
+ PAND2X1_288/a_76_28# PAND2X1
XPAND2X1_277 VDD GND PAND2X1_48/B PAND2X1_90/A POR2X1_633/A PAND2X1_277/a_16_344#
+ PAND2X1_277/m4_208_n4# PAND2X1_277/O PAND2X1_277/a_56_28# PAND2X1_277/CTRL2 PAND2X1_277/CTRL
+ PAND2X1_277/a_76_28# PAND2X1
XPAND2X1_299 VDD GND POR2X1_121/B POR2X1_260/B POR2X1_302/A PAND2X1_299/a_16_344#
+ PAND2X1_299/m4_208_n4# PAND2X1_299/O PAND2X1_299/a_56_28# PAND2X1_299/CTRL2 PAND2X1_299/CTRL
+ PAND2X1_299/a_76_28# PAND2X1
XPOR2X1_803 VDD GND POR2X1_796/Y POR2X1_803/A POR2X1_808/B POR2X1_803/m4_208_n4# POR2X1_803/O
+ POR2X1_803/CTRL2 POR2X1_803/a_16_28# POR2X1_803/CTRL POR2X1_803/a_76_344# POR2X1_803/a_56_344#
+ POR2X1
XPOR2X1_836 VDD GND POR2X1_836/B POR2X1_836/A POR2X1_836/Y POR2X1_836/m4_208_n4# POR2X1_836/O
+ POR2X1_836/CTRL2 POR2X1_836/a_16_28# POR2X1_836/CTRL POR2X1_836/a_76_344# POR2X1_836/a_56_344#
+ POR2X1
XPOR2X1_825 VDD GND POR2X1_57/A POR2X1_96/B POR2X1_825/Y POR2X1_825/m4_208_n4# POR2X1_825/O
+ POR2X1_825/CTRL2 POR2X1_825/a_16_28# POR2X1_825/CTRL POR2X1_825/a_76_344# POR2X1_825/a_56_344#
+ POR2X1
XPOR2X1_814 VDD GND POR2X1_814/B POR2X1_814/A POR2X1_814/Y POR2X1_814/m4_208_n4# POR2X1_814/O
+ POR2X1_814/CTRL2 POR2X1_814/a_16_28# POR2X1_814/CTRL POR2X1_814/a_76_344# POR2X1_814/a_56_344#
+ POR2X1
XPOR2X1_847 VDD GND POR2X1_847/B POR2X1_847/A POR2X1_848/A POR2X1_847/m4_208_n4# POR2X1_847/O
+ POR2X1_847/CTRL2 POR2X1_847/a_16_28# POR2X1_847/CTRL POR2X1_847/a_76_344# POR2X1_847/a_56_344#
+ POR2X1
XPOR2X1_858 VDD GND POR2X1_858/B POR2X1_858/A POR2X1_862/B POR2X1_858/m4_208_n4# POR2X1_858/O
+ POR2X1_858/CTRL2 POR2X1_858/a_16_28# POR2X1_858/CTRL POR2X1_858/a_76_344# POR2X1_858/a_56_344#
+ POR2X1
XPAND2X1_42 VDD GND PAND2X1_90/A INPUT_1 POR2X1_296/B PAND2X1_42/a_16_344# PAND2X1_42/m4_208_n4#
+ PAND2X1_42/O PAND2X1_42/a_56_28# PAND2X1_42/CTRL2 PAND2X1_42/CTRL PAND2X1_42/a_76_28#
+ PAND2X1
XPAND2X1_53 VDD GND PAND2X1_95/B D_INPUT_5 PAND2X1_56/A PAND2X1_53/a_16_344# PAND2X1_53/m4_208_n4#
+ PAND2X1_53/O PAND2X1_53/a_56_28# PAND2X1_53/CTRL2 PAND2X1_53/CTRL PAND2X1_53/a_76_28#
+ PAND2X1
XPAND2X1_31 VDD GND PAND2X1_47/B PAND2X1_3/A PAND2X1_32/B PAND2X1_31/a_16_344# PAND2X1_31/m4_208_n4#
+ PAND2X1_31/O PAND2X1_31/a_56_28# PAND2X1_31/CTRL2 PAND2X1_31/CTRL PAND2X1_31/a_76_28#
+ PAND2X1
XPAND2X1_20 VDD GND PAND2X1_19/Y PAND2X1_20/A POR2X1_33/B PAND2X1_20/a_16_344# PAND2X1_20/m4_208_n4#
+ PAND2X1_20/O PAND2X1_20/a_56_28# PAND2X1_20/CTRL2 PAND2X1_20/CTRL PAND2X1_20/a_76_28#
+ PAND2X1
XPAND2X1_75 VDD GND PAND2X1_60/B PAND2X1_23/Y POR2X1_76/A PAND2X1_75/a_16_344# PAND2X1_75/m4_208_n4#
+ PAND2X1_75/O PAND2X1_75/a_56_28# PAND2X1_75/CTRL2 PAND2X1_75/CTRL PAND2X1_75/a_76_28#
+ PAND2X1
XPAND2X1_64 VDD GND PAND2X1_95/B PAND2X1_26/A PAND2X1_65/B PAND2X1_64/a_16_344# PAND2X1_64/m4_208_n4#
+ PAND2X1_64/O PAND2X1_64/a_56_28# PAND2X1_64/CTRL2 PAND2X1_64/CTRL PAND2X1_64/a_76_28#
+ PAND2X1
XPOR2X1_17 VDD GND D_INPUT_6 D_INPUT_7 POR2X1_36/B POR2X1_17/m4_208_n4# POR2X1_17/O
+ POR2X1_17/CTRL2 POR2X1_17/a_16_28# POR2X1_17/CTRL POR2X1_17/a_76_344# POR2X1_17/a_56_344#
+ POR2X1
XPAND2X1_86 VDD GND PAND2X1_85/Y INPUT_0 PAND2X1_86/Y PAND2X1_86/a_16_344# PAND2X1_86/m4_208_n4#
+ PAND2X1_86/O PAND2X1_86/a_56_28# PAND2X1_86/CTRL2 PAND2X1_86/CTRL PAND2X1_86/a_76_28#
+ PAND2X1
XPAND2X1_97 VDD GND POR2X1_91/Y POR2X1_89/Y PAND2X1_97/Y PAND2X1_97/a_16_344# PAND2X1_97/m4_208_n4#
+ PAND2X1_97/O PAND2X1_97/a_56_28# PAND2X1_97/CTRL2 PAND2X1_97/CTRL PAND2X1_97/a_76_28#
+ PAND2X1
XPOR2X1_611 VDD GND POR2X1_5/Y POR2X1_94/A POR2X1_612/A POR2X1_611/m4_208_n4# POR2X1_611/O
+ POR2X1_611/CTRL2 POR2X1_611/a_16_28# POR2X1_611/CTRL POR2X1_611/a_76_344# POR2X1_611/a_56_344#
+ POR2X1
XPOR2X1_600 VDD GND POR2X1_32/A POR2X1_411/B POR2X1_600/Y POR2X1_600/m4_208_n4# POR2X1_600/O
+ POR2X1_600/CTRL2 POR2X1_600/a_16_28# POR2X1_600/CTRL POR2X1_600/a_76_344# POR2X1_600/a_56_344#
+ POR2X1
XPOR2X1_28 VDD GND INPUT_0 D_INPUT_1 POR2X1_38/B POR2X1_28/m4_208_n4# POR2X1_28/O
+ POR2X1_28/CTRL2 POR2X1_28/a_16_28# POR2X1_28/CTRL POR2X1_28/a_76_344# POR2X1_28/a_56_344#
+ POR2X1
XPOR2X1_39 VDD GND POR2X1_39/B POR2X1_38/Y POR2X1_39/Y POR2X1_39/m4_208_n4# POR2X1_39/O
+ POR2X1_39/CTRL2 POR2X1_39/a_16_28# POR2X1_39/CTRL POR2X1_39/a_76_344# POR2X1_39/a_56_344#
+ POR2X1
XPOR2X1_622 VDD GND POR2X1_622/B POR2X1_622/A POR2X1_624/B POR2X1_622/m4_208_n4# POR2X1_622/O
+ POR2X1_622/CTRL2 POR2X1_622/a_16_28# POR2X1_622/CTRL POR2X1_622/a_76_344# POR2X1_622/a_56_344#
+ POR2X1
XPOR2X1_633 VDD GND POR2X1_123/A POR2X1_633/A POR2X1_633/Y POR2X1_633/m4_208_n4# POR2X1_633/O
+ POR2X1_633/CTRL2 POR2X1_633/a_16_28# POR2X1_633/CTRL POR2X1_633/a_76_344# POR2X1_633/a_56_344#
+ POR2X1
XPOR2X1_644 VDD GND POR2X1_644/B POR2X1_644/A POR2X1_644/Y POR2X1_644/m4_208_n4# POR2X1_644/O
+ POR2X1_644/CTRL2 POR2X1_644/a_16_28# POR2X1_644/CTRL POR2X1_644/a_76_344# POR2X1_644/a_56_344#
+ POR2X1
XPOR2X1_666 VDD GND POR2X1_20/B POR2X1_666/A POR2X1_666/Y POR2X1_666/m4_208_n4# POR2X1_666/O
+ POR2X1_666/CTRL2 POR2X1_666/a_16_28# POR2X1_666/CTRL POR2X1_666/a_76_344# POR2X1_666/a_56_344#
+ POR2X1
XPOR2X1_677 VDD GND POR2X1_83/B POR2X1_257/A POR2X1_677/Y POR2X1_677/m4_208_n4# POR2X1_677/O
+ POR2X1_677/CTRL2 POR2X1_677/a_16_28# POR2X1_677/CTRL POR2X1_677/a_76_344# POR2X1_677/a_56_344#
+ POR2X1
XPOR2X1_655 VDD GND POR2X1_648/Y POR2X1_655/A POR2X1_655/Y POR2X1_655/m4_208_n4# POR2X1_655/O
+ POR2X1_655/CTRL2 POR2X1_655/a_16_28# POR2X1_655/CTRL POR2X1_655/a_76_344# POR2X1_655/a_56_344#
+ POR2X1
XPOR2X1_688 VDD GND PAND2X1_39/B POR2X1_294/A POR2X1_688/Y POR2X1_688/m4_208_n4# POR2X1_688/O
+ POR2X1_688/CTRL2 POR2X1_688/a_16_28# POR2X1_688/CTRL POR2X1_688/a_76_344# POR2X1_688/a_56_344#
+ POR2X1
XPOR2X1_699 VDD GND POR2X1_14/Y POR2X1_416/B POR2X1_748/A POR2X1_699/m4_208_n4# POR2X1_699/O
+ POR2X1_699/CTRL2 POR2X1_699/a_16_28# POR2X1_699/CTRL POR2X1_699/a_76_344# POR2X1_699/a_56_344#
+ POR2X1
XPAND2X1_629 VDD GND POR2X1_627/Y POR2X1_626/Y PAND2X1_630/B PAND2X1_629/a_16_344#
+ PAND2X1_629/m4_208_n4# PAND2X1_629/O PAND2X1_629/a_56_28# PAND2X1_629/CTRL2 PAND2X1_629/CTRL
+ PAND2X1_629/a_76_28# PAND2X1
XPAND2X1_607 VDD GND POR2X1_606/Y PAND2X1_20/A POR2X1_646/B PAND2X1_607/a_16_344#
+ PAND2X1_607/m4_208_n4# PAND2X1_607/O PAND2X1_607/a_56_28# PAND2X1_607/CTRL2 PAND2X1_607/CTRL
+ PAND2X1_607/a_76_28# PAND2X1
XPAND2X1_618 VDD GND POR2X1_29/A D_INPUT_3 PAND2X1_618/Y PAND2X1_618/a_16_344# PAND2X1_618/m4_208_n4#
+ PAND2X1_618/O PAND2X1_618/a_56_28# PAND2X1_618/CTRL2 PAND2X1_618/CTRL PAND2X1_618/a_76_28#
+ PAND2X1
XPOR2X1_441 VDD GND POR2X1_40/Y POR2X1_49/Y POR2X1_441/Y POR2X1_441/m4_208_n4# POR2X1_441/O
+ POR2X1_441/CTRL2 POR2X1_441/a_16_28# POR2X1_441/CTRL POR2X1_441/a_76_344# POR2X1_441/a_56_344#
+ POR2X1
XPOR2X1_452 VDD GND POR2X1_450/Y POR2X1_452/A POR2X1_452/Y POR2X1_452/m4_208_n4# POR2X1_452/O
+ POR2X1_452/CTRL2 POR2X1_452/a_16_28# POR2X1_452/CTRL POR2X1_452/a_76_344# POR2X1_452/a_56_344#
+ POR2X1
XPOR2X1_430 VDD GND POR2X1_669/B POR2X1_430/A POR2X1_430/Y POR2X1_430/m4_208_n4# POR2X1_430/O
+ POR2X1_430/CTRL2 POR2X1_430/a_16_28# POR2X1_430/CTRL POR2X1_430/a_76_344# POR2X1_430/a_56_344#
+ POR2X1
XPOR2X1_474 VDD GND POR2X1_860/A POR2X1_404/Y POR2X1_475/A POR2X1_474/m4_208_n4# POR2X1_474/O
+ POR2X1_474/CTRL2 POR2X1_474/a_16_28# POR2X1_474/CTRL POR2X1_474/a_76_344# POR2X1_474/a_56_344#
+ POR2X1
XPOR2X1_485 VDD GND POR2X1_57/A POR2X1_102/Y POR2X1_485/Y POR2X1_485/m4_208_n4# POR2X1_485/O
+ POR2X1_485/CTRL2 POR2X1_485/a_16_28# POR2X1_485/CTRL POR2X1_485/a_76_344# POR2X1_485/a_56_344#
+ POR2X1
XPOR2X1_463 VDD GND POR2X1_459/Y POR2X1_460/Y POR2X1_463/Y POR2X1_463/m4_208_n4# POR2X1_463/O
+ POR2X1_463/CTRL2 POR2X1_463/a_16_28# POR2X1_463/CTRL POR2X1_463/a_76_344# POR2X1_463/a_56_344#
+ POR2X1
XPOR2X1_496 VDD GND POR2X1_20/B POR2X1_55/Y POR2X1_496/Y POR2X1_496/m4_208_n4# POR2X1_496/O
+ POR2X1_496/CTRL2 POR2X1_496/a_16_28# POR2X1_496/CTRL POR2X1_496/a_76_344# POR2X1_496/a_56_344#
+ POR2X1
XPAND2X1_404 VDD GND PAND2X1_403/Y PAND2X1_404/A PAND2X1_404/Y PAND2X1_404/a_16_344#
+ PAND2X1_404/m4_208_n4# PAND2X1_404/O PAND2X1_404/a_56_28# PAND2X1_404/CTRL2 PAND2X1_404/CTRL
+ PAND2X1_404/a_76_28# PAND2X1
XPAND2X1_437 VDD GND POR2X1_186/B PAND2X1_60/B POR2X1_440/B PAND2X1_437/a_16_344#
+ PAND2X1_437/m4_208_n4# PAND2X1_437/O PAND2X1_437/a_56_28# PAND2X1_437/CTRL2 PAND2X1_437/CTRL
+ PAND2X1_437/a_76_28# PAND2X1
XPAND2X1_426 VDD GND PAND2X1_425/Y POR2X1_121/B POR2X1_450/B PAND2X1_426/a_16_344#
+ PAND2X1_426/m4_208_n4# PAND2X1_426/O PAND2X1_426/a_56_28# PAND2X1_426/CTRL2 PAND2X1_426/CTRL
+ PAND2X1_426/a_76_28# PAND2X1
XPAND2X1_415 VDD GND POR2X1_414/Y POR2X1_293/Y POR2X1_416/A PAND2X1_415/a_16_344#
+ PAND2X1_415/m4_208_n4# PAND2X1_415/O PAND2X1_415/a_56_28# PAND2X1_415/CTRL2 PAND2X1_415/CTRL
+ PAND2X1_415/a_76_28# PAND2X1
XPAND2X1_448 VDD GND POR2X1_422/Y POR2X1_421/Y PAND2X1_453/A PAND2X1_448/a_16_344#
+ PAND2X1_448/m4_208_n4# PAND2X1_448/O PAND2X1_448/a_56_28# PAND2X1_448/CTRL2 PAND2X1_448/CTRL
+ PAND2X1_448/a_76_28# PAND2X1
XPAND2X1_459 VDD GND POR2X1_378/Y POR2X1_376/Y PAND2X1_459/Y PAND2X1_459/a_16_344#
+ PAND2X1_459/m4_208_n4# PAND2X1_459/O PAND2X1_459/a_56_28# PAND2X1_459/CTRL2 PAND2X1_459/CTRL
+ PAND2X1_459/a_76_28# PAND2X1
XPOR2X1_260 VDD GND POR2X1_260/B POR2X1_260/A POR2X1_260/Y POR2X1_260/m4_208_n4# POR2X1_260/O
+ POR2X1_260/CTRL2 POR2X1_260/a_16_28# POR2X1_260/CTRL POR2X1_260/a_76_344# POR2X1_260/a_56_344#
+ POR2X1
XPOR2X1_271 VDD GND POR2X1_271/B POR2X1_271/A POR2X1_271/Y POR2X1_271/m4_208_n4# POR2X1_271/O
+ POR2X1_271/CTRL2 POR2X1_271/a_16_28# POR2X1_271/CTRL POR2X1_271/a_76_344# POR2X1_271/a_56_344#
+ POR2X1
XPOR2X1_293 VDD GND D_INPUT_1 POR2X1_5/Y POR2X1_293/Y POR2X1_293/m4_208_n4# POR2X1_293/O
+ POR2X1_293/CTRL2 POR2X1_293/a_16_28# POR2X1_293/CTRL POR2X1_293/a_76_344# POR2X1_293/a_56_344#
+ POR2X1
XPOR2X1_282 VDD GND POR2X1_102/Y POR2X1_416/B POR2X1_282/Y POR2X1_282/m4_208_n4# POR2X1_282/O
+ POR2X1_282/CTRL2 POR2X1_282/a_16_28# POR2X1_282/CTRL POR2X1_282/a_76_344# POR2X1_282/a_56_344#
+ POR2X1
XPAND2X1_201 VDD GND POR2X1_65/Y PAND2X1_61/Y PAND2X1_206/A PAND2X1_201/a_16_344#
+ POR2X1_65/m4_208_n4# PAND2X1_201/O PAND2X1_201/a_56_28# PAND2X1_201/CTRL2 PAND2X1_201/CTRL
+ PAND2X1_201/a_76_28# PAND2X1
XPAND2X1_212 VDD GND PAND2X1_212/B PAND2X1_352/A PAND2X1_220/A PAND2X1_212/a_16_344#
+ PAND2X1_212/m4_208_n4# PAND2X1_212/O PAND2X1_212/a_56_28# PAND2X1_212/CTRL2 PAND2X1_212/CTRL
+ PAND2X1_212/a_76_28# PAND2X1
XPAND2X1_245 VDD GND PAND2X1_90/A POR2X1_66/A POR2X1_777/B PAND2X1_245/a_16_344# PAND2X1_245/m4_208_n4#
+ PAND2X1_245/O PAND2X1_245/a_56_28# PAND2X1_245/CTRL2 PAND2X1_245/CTRL PAND2X1_245/a_76_28#
+ PAND2X1
XPAND2X1_223 VDD GND PAND2X1_223/B PAND2X1_221/Y GATE_222 PAND2X1_223/a_16_344# PAND2X1_365/m4_208_n4#
+ PAND2X1_223/O PAND2X1_223/a_56_28# PAND2X1_223/CTRL2 PAND2X1_223/CTRL PAND2X1_223/a_76_28#
+ PAND2X1
XPAND2X1_234 VDD GND PAND2X1_824/B PAND2X1_48/B POR2X1_240/A PAND2X1_234/a_16_344#
+ PAND2X1_234/m4_208_n4# PAND2X1_234/O PAND2X1_234/a_56_28# PAND2X1_234/CTRL2 PAND2X1_234/CTRL
+ PAND2X1_234/a_76_28# PAND2X1
XPAND2X1_256 VDD GND POR2X1_541/B POR2X1_4/Y POR2X1_344/A PAND2X1_256/a_16_344# POR2X1_349/m4_208_n4#
+ PAND2X1_256/O PAND2X1_256/a_56_28# PAND2X1_256/CTRL2 PAND2X1_256/CTRL PAND2X1_256/a_76_28#
+ PAND2X1
XPAND2X1_267 VDD GND PAND2X1_267/B POR2X1_265/Y PAND2X1_267/Y PAND2X1_267/a_16_344#
+ PAND2X1_267/m4_208_n4# PAND2X1_267/O PAND2X1_267/a_56_28# PAND2X1_267/CTRL2 PAND2X1_267/CTRL
+ PAND2X1_267/a_76_28# PAND2X1
XPAND2X1_278 VDD GND POR2X1_633/A POR2X1_9/Y POR2X1_287/B PAND2X1_278/a_16_344# PAND2X1_278/m4_208_n4#
+ PAND2X1_278/O PAND2X1_278/a_56_28# PAND2X1_278/CTRL2 PAND2X1_278/CTRL PAND2X1_278/a_76_28#
+ PAND2X1
XPAND2X1_289 VDD GND POR2X1_814/A PAND2X1_52/B POR2X1_333/A PAND2X1_289/a_16_344#
+ PAND2X1_289/m4_208_n4# PAND2X1_289/O PAND2X1_289/a_56_28# PAND2X1_289/CTRL2 PAND2X1_289/CTRL
+ PAND2X1_289/a_76_28# PAND2X1
XPAND2X1_790 VDD GND POR2X1_754/Y POR2X1_753/Y PAND2X1_790/Y PAND2X1_790/a_16_344#
+ PAND2X1_790/m4_208_n4# PAND2X1_790/O PAND2X1_790/a_56_28# PAND2X1_790/CTRL2 PAND2X1_790/CTRL
+ PAND2X1_790/a_76_28# PAND2X1
XPOR2X1_826 VDD GND POR2X1_55/Y POR2X1_96/A POR2X1_826/Y POR2X1_826/m4_208_n4# POR2X1_826/O
+ POR2X1_826/CTRL2 POR2X1_826/a_16_28# POR2X1_826/CTRL POR2X1_826/a_76_344# POR2X1_826/a_56_344#
+ POR2X1
XPOR2X1_815 VDD GND POR2X1_7/B POR2X1_815/A POR2X1_815/Y POR2X1_815/m4_208_n4# POR2X1_815/O
+ POR2X1_815/CTRL2 POR2X1_815/a_16_28# POR2X1_815/CTRL POR2X1_815/a_76_344# POR2X1_815/a_56_344#
+ POR2X1
XPOR2X1_804 VDD GND POR2X1_804/B POR2X1_804/A POR2X1_808/A POR2X1_804/m4_208_n4# POR2X1_804/O
+ POR2X1_804/CTRL2 POR2X1_804/a_16_28# POR2X1_804/CTRL POR2X1_804/a_76_344# POR2X1_804/a_56_344#
+ POR2X1
XPOR2X1_837 VDD GND POR2X1_837/B POR2X1_837/A POR2X1_837/Y POR2X1_837/m4_208_n4# POR2X1_837/O
+ POR2X1_837/CTRL2 POR2X1_837/a_16_28# POR2X1_837/CTRL POR2X1_837/a_76_344# POR2X1_837/a_56_344#
+ POR2X1
XPOR2X1_848 VDD GND POR2X1_846/Y POR2X1_848/A POR2X1_848/Y POR2X1_848/m4_208_n4# POR2X1_848/O
+ POR2X1_848/CTRL2 POR2X1_848/a_16_28# POR2X1_848/CTRL POR2X1_848/a_76_344# POR2X1_848/a_56_344#
+ POR2X1
XPOR2X1_859 VDD GND POR2X1_848/Y POR2X1_859/A POR2X1_862/A POR2X1_859/m4_208_n4# POR2X1_859/O
+ POR2X1_859/CTRL2 POR2X1_859/a_16_28# POR2X1_859/CTRL POR2X1_859/a_76_344# POR2X1_859/a_56_344#
+ POR2X1
XPAND2X1_10 VDD GND PAND2X1_9/Y PAND2X1_8/Y POR2X1_294/B PAND2X1_10/a_16_344# PAND2X1_10/m4_208_n4#
+ PAND2X1_10/O PAND2X1_10/a_56_28# PAND2X1_10/CTRL2 PAND2X1_10/CTRL PAND2X1_10/a_76_28#
+ PAND2X1
XPAND2X1_21 VDD GND D_INPUT_5 INPUT_4 PAND2X1_26/A PAND2X1_21/a_16_344# PAND2X1_21/m4_208_n4#
+ PAND2X1_21/O PAND2X1_21/a_56_28# PAND2X1_21/CTRL2 PAND2X1_21/CTRL PAND2X1_21/a_76_28#
+ PAND2X1
XPAND2X1_32 VDD GND PAND2X1_32/B POR2X1_87/B POR2X1_34/A PAND2X1_32/a_16_344# PAND2X1_32/m4_208_n4#
+ PAND2X1_32/O PAND2X1_32/a_56_28# PAND2X1_32/CTRL2 PAND2X1_32/CTRL PAND2X1_32/a_76_28#
+ PAND2X1
XPAND2X1_43 VDD GND POR2X1_296/B PAND2X1_58/A POR2X1_195/A PAND2X1_43/a_16_344# PAND2X1_43/m4_208_n4#
+ PAND2X1_43/O PAND2X1_43/a_56_28# PAND2X1_43/CTRL2 PAND2X1_43/CTRL PAND2X1_43/a_76_28#
+ PAND2X1
XPAND2X1_65 VDD GND PAND2X1_65/B PAND2X1_63/Y PAND2X1_65/Y PAND2X1_65/a_16_344# PAND2X1_65/m4_208_n4#
+ PAND2X1_65/O PAND2X1_65/a_56_28# PAND2X1_65/CTRL2 PAND2X1_65/CTRL PAND2X1_65/a_76_28#
+ PAND2X1
XPAND2X1_76 VDD GND POR2X1_75/Y POR2X1_74/Y PAND2X1_76/Y PAND2X1_76/a_16_344# PAND2X1_76/m4_208_n4#
+ PAND2X1_76/O PAND2X1_76/a_56_28# PAND2X1_76/CTRL2 PAND2X1_76/CTRL PAND2X1_76/a_76_28#
+ PAND2X1
XPAND2X1_54 VDD GND INPUT_1 INPUT_0 POR2X1_94/A PAND2X1_54/a_16_344# PAND2X1_54/m4_208_n4#
+ PAND2X1_54/O PAND2X1_54/a_56_28# PAND2X1_54/CTRL2 PAND2X1_54/CTRL PAND2X1_54/a_76_28#
+ PAND2X1
XPAND2X1_87 VDD GND POR2X1_49/Y POR2X1_29/Y POR2X1_88/A PAND2X1_87/a_16_344# POR2X1_88/m4_208_n4#
+ PAND2X1_87/O PAND2X1_87/a_56_28# PAND2X1_87/CTRL2 PAND2X1_87/CTRL PAND2X1_87/a_76_28#
+ PAND2X1
XPAND2X1_98 VDD GND POR2X1_96/Y POR2X1_93/Y PAND2X1_99/B PAND2X1_98/a_16_344# PAND2X1_98/m4_208_n4#
+ PAND2X1_98/O PAND2X1_98/a_56_28# PAND2X1_98/CTRL2 PAND2X1_98/CTRL PAND2X1_98/a_76_28#
+ PAND2X1
XPOR2X1_601 VDD GND POR2X1_16/A POR2X1_48/A POR2X1_601/Y POR2X1_601/m4_208_n4# POR2X1_601/O
+ POR2X1_601/CTRL2 POR2X1_601/a_16_28# POR2X1_601/CTRL POR2X1_601/a_76_344# POR2X1_601/a_56_344#
+ POR2X1
XPOR2X1_29 VDD GND POR2X1_8/Y POR2X1_29/A POR2X1_29/Y POR2X1_29/m4_208_n4# POR2X1_29/O
+ POR2X1_29/CTRL2 POR2X1_29/a_16_28# POR2X1_29/CTRL POR2X1_29/a_76_344# POR2X1_29/a_56_344#
+ POR2X1
XPOR2X1_18 VDD GND POR2X1_12/A POR2X1_36/B POR2X1_20/B POR2X1_18/m4_208_n4# POR2X1_18/O
+ POR2X1_18/CTRL2 POR2X1_18/a_16_28# POR2X1_18/CTRL POR2X1_18/a_76_344# POR2X1_18/a_56_344#
+ POR2X1
XPOR2X1_612 VDD GND POR2X1_612/B POR2X1_612/A POR2X1_612/Y POR2X1_612/m4_208_n4# POR2X1_612/O
+ POR2X1_612/CTRL2 POR2X1_612/a_16_28# POR2X1_612/CTRL POR2X1_612/a_76_344# POR2X1_612/a_56_344#
+ POR2X1
XPOR2X1_623 VDD GND POR2X1_623/B POR2X1_623/A POR2X1_623/Y POR2X1_623/m4_208_n4# POR2X1_623/O
+ POR2X1_623/CTRL2 POR2X1_623/a_16_28# POR2X1_623/CTRL POR2X1_623/a_76_344# POR2X1_623/a_56_344#
+ POR2X1
XPOR2X1_634 VDD GND POR2X1_334/B POR2X1_634/A POR2X1_640/A POR2X1_634/m4_208_n4# POR2X1_634/O
+ POR2X1_634/CTRL2 POR2X1_634/a_16_28# POR2X1_634/CTRL POR2X1_634/a_76_344# POR2X1_634/a_56_344#
+ POR2X1
XPOR2X1_645 VDD GND POR2X1_788/A POR2X1_718/A POR2X1_648/A POR2X1_645/m4_208_n4# POR2X1_645/O
+ POR2X1_645/CTRL2 POR2X1_645/a_16_28# POR2X1_645/CTRL POR2X1_645/a_76_344# POR2X1_645/a_56_344#
+ POR2X1
XPOR2X1_667 VDD GND POR2X1_65/A POR2X1_667/A POR2X1_667/Y POR2X1_667/m4_208_n4# POR2X1_667/O
+ POR2X1_667/CTRL2 POR2X1_667/a_16_28# POR2X1_667/CTRL POR2X1_667/a_76_344# POR2X1_667/a_56_344#
+ POR2X1
XPOR2X1_678 VDD GND POR2X1_260/B POR2X1_678/A POR2X1_678/Y POR2X1_678/m4_208_n4# POR2X1_678/O
+ POR2X1_678/CTRL2 POR2X1_678/a_16_28# POR2X1_678/CTRL POR2X1_678/a_76_344# POR2X1_678/a_56_344#
+ POR2X1
XPOR2X1_656 VDD GND POR2X1_101/Y POR2X1_647/Y POR2X1_660/A POR2X1_656/m4_208_n4# POR2X1_656/O
+ POR2X1_656/CTRL2 POR2X1_656/a_16_28# POR2X1_656/CTRL POR2X1_656/a_76_344# POR2X1_656/a_56_344#
+ POR2X1
XPOR2X1_689 VDD GND POR2X1_32/A POR2X1_689/A POR2X1_689/Y POR2X1_689/m4_208_n4# POR2X1_689/O
+ POR2X1_689/CTRL2 POR2X1_689/a_16_28# POR2X1_689/CTRL POR2X1_689/a_76_344# POR2X1_689/a_56_344#
+ POR2X1
XPAND2X1_608 VDD GND POR2X1_73/Y POR2X1_16/A POR2X1_609/A PAND2X1_608/a_16_344# PAND2X1_608/m4_208_n4#
+ PAND2X1_608/O PAND2X1_608/a_56_28# PAND2X1_608/CTRL2 PAND2X1_608/CTRL PAND2X1_608/a_76_28#
+ PAND2X1
XPAND2X1_619 VDD GND PAND2X1_618/Y PAND2X1_69/A POR2X1_622/B PAND2X1_619/a_16_344#
+ PAND2X1_619/m4_208_n4# PAND2X1_619/O PAND2X1_619/a_56_28# PAND2X1_619/CTRL2 PAND2X1_619/CTRL
+ PAND2X1_619/a_76_28# PAND2X1
XPOR2X1_431 VDD GND POR2X1_72/B POR2X1_236/Y POR2X1_431/Y POR2X1_431/m4_208_n4# POR2X1_431/O
+ POR2X1_431/CTRL2 POR2X1_431/a_16_28# POR2X1_431/CTRL POR2X1_431/a_76_344# POR2X1_431/a_56_344#
+ POR2X1
XPOR2X1_442 VDD GND POR2X1_40/Y POR2X1_411/B POR2X1_442/Y POR2X1_442/m4_208_n4# POR2X1_442/O
+ POR2X1_442/CTRL2 POR2X1_442/a_16_28# POR2X1_442/CTRL POR2X1_442/a_76_344# POR2X1_442/a_56_344#
+ POR2X1
XPOR2X1_420 VDD GND POR2X1_96/A POR2X1_102/Y POR2X1_420/Y POR2X1_420/m4_208_n4# POR2X1_420/O
+ POR2X1_420/CTRL2 POR2X1_420/a_16_28# POR2X1_420/CTRL POR2X1_420/a_76_344# POR2X1_420/a_56_344#
+ POR2X1
XPOR2X1_453 VDD GND POR2X1_448/Y POR2X1_449/Y POR2X1_453/Y POR2X1_453/m4_208_n4# POR2X1_453/O
+ POR2X1_453/CTRL2 POR2X1_453/a_16_28# POR2X1_453/CTRL POR2X1_453/a_76_344# POR2X1_453/a_56_344#
+ POR2X1
XPOR2X1_464 VDD GND POR2X1_457/Y POR2X1_458/Y POR2X1_464/Y POR2X1_464/m4_208_n4# POR2X1_464/O
+ POR2X1_464/CTRL2 POR2X1_464/a_16_28# POR2X1_464/CTRL POR2X1_464/a_76_344# POR2X1_464/a_56_344#
+ POR2X1
XPOR2X1_486 VDD GND POR2X1_486/B POR2X1_705/B POR2X1_556/A POR2X1_486/m4_208_n4# POR2X1_486/O
+ POR2X1_486/CTRL2 POR2X1_486/a_16_28# POR2X1_486/CTRL POR2X1_486/a_76_344# POR2X1_486/a_56_344#
+ POR2X1
XPOR2X1_475 VDD GND POR2X1_734/B POR2X1_475/A POR2X1_479/B POR2X1_475/m4_208_n4# POR2X1_475/O
+ POR2X1_475/CTRL2 POR2X1_475/a_16_28# POR2X1_475/CTRL POR2X1_475/a_76_344# POR2X1_475/a_56_344#
+ POR2X1
XPOR2X1_497 VDD GND POR2X1_43/B POR2X1_71/Y POR2X1_497/Y POR2X1_71/m4_208_n4# POR2X1_497/O
+ POR2X1_497/CTRL2 POR2X1_497/a_16_28# POR2X1_497/CTRL POR2X1_497/a_76_344# POR2X1_497/a_56_344#
+ POR2X1
XPAND2X1_405 VDD GND POR2X1_760/A POR2X1_46/Y POR2X1_406/A PAND2X1_405/a_16_344# PAND2X1_405/m4_208_n4#
+ PAND2X1_405/O PAND2X1_405/a_56_28# PAND2X1_405/CTRL2 PAND2X1_405/CTRL PAND2X1_405/a_76_28#
+ PAND2X1
XPAND2X1_416 VDD GND POR2X1_415/Y POR2X1_260/A POR2X1_462/B PAND2X1_416/a_16_344#
+ PAND2X1_416/m4_208_n4# PAND2X1_416/O PAND2X1_416/a_56_28# PAND2X1_416/CTRL2 PAND2X1_416/CTRL
+ PAND2X1_416/a_76_28# PAND2X1
XPAND2X1_427 VDD GND POR2X1_614/A PAND2X1_72/A POR2X1_450/A PAND2X1_427/a_16_344#
+ PAND2X1_427/m4_208_n4# PAND2X1_427/O PAND2X1_427/a_56_28# PAND2X1_427/CTRL2 PAND2X1_427/CTRL
+ PAND2X1_427/a_76_28# PAND2X1
XPAND2X1_438 VDD GND PAND2X1_72/A PAND2X1_23/Y POR2X1_544/A PAND2X1_438/a_16_344#
+ PAND2X1_438/m4_208_n4# PAND2X1_438/O PAND2X1_438/a_56_28# PAND2X1_438/CTRL2 PAND2X1_438/CTRL
+ PAND2X1_438/a_76_28# PAND2X1
XPAND2X1_449 VDD GND POR2X1_424/Y POR2X1_423/Y PAND2X1_449/Y PAND2X1_449/a_16_344#
+ PAND2X1_449/m4_208_n4# PAND2X1_449/O PAND2X1_449/a_56_28# PAND2X1_449/CTRL2 PAND2X1_449/CTRL
+ PAND2X1_449/a_76_28# PAND2X1
XPOR2X1_250 VDD GND POR2X1_65/A POR2X1_250/A POR2X1_250/Y POR2X1_250/m4_208_n4# POR2X1_250/O
+ POR2X1_250/CTRL2 POR2X1_250/a_16_28# POR2X1_250/CTRL POR2X1_250/a_76_344# POR2X1_250/a_56_344#
+ POR2X1
XPOR2X1_261 VDD GND POR2X1_411/B POR2X1_261/A POR2X1_261/Y POR2X1_261/m4_208_n4# POR2X1_261/O
+ POR2X1_261/CTRL2 POR2X1_261/a_16_28# POR2X1_261/CTRL POR2X1_261/a_76_344# POR2X1_261/a_56_344#
+ POR2X1
XPOR2X1_294 VDD GND POR2X1_294/B POR2X1_294/A POR2X1_294/Y POR2X1_294/m4_208_n4# POR2X1_294/O
+ POR2X1_294/CTRL2 POR2X1_294/a_16_28# POR2X1_294/CTRL POR2X1_294/a_76_344# POR2X1_294/a_56_344#
+ POR2X1
XPOR2X1_283 VDD GND POR2X1_83/B POR2X1_283/A POR2X1_283/Y POR2X1_283/m4_208_n4# POR2X1_283/O
+ POR2X1_283/CTRL2 POR2X1_283/a_16_28# POR2X1_283/CTRL POR2X1_283/a_76_344# POR2X1_283/a_56_344#
+ POR2X1
XPOR2X1_272 VDD GND POR2X1_32/A POR2X1_42/Y POR2X1_272/Y POR2X1_272/m4_208_n4# POR2X1_272/O
+ POR2X1_272/CTRL2 POR2X1_272/a_16_28# POR2X1_272/CTRL POR2X1_272/a_76_344# POR2X1_272/a_56_344#
+ POR2X1
XPAND2X1_202 VDD GND POR2X1_69/Y POR2X1_67/Y PAND2X1_206/B PAND2X1_202/a_16_344# PAND2X1_202/m4_208_n4#
+ PAND2X1_202/O PAND2X1_202/a_56_28# PAND2X1_202/CTRL2 PAND2X1_202/CTRL PAND2X1_202/a_76_28#
+ PAND2X1
XPAND2X1_246 VDD GND POR2X1_777/B PAND2X1_9/Y POR2X1_342/B PAND2X1_246/a_16_344# PAND2X1_246/m4_208_n4#
+ PAND2X1_246/O PAND2X1_246/a_56_28# PAND2X1_246/CTRL2 PAND2X1_246/CTRL PAND2X1_246/a_76_28#
+ PAND2X1
XPAND2X1_213 VDD GND PAND2X1_213/B PAND2X1_213/A PAND2X1_213/Y PAND2X1_213/a_16_344#
+ PAND2X1_213/m4_208_n4# PAND2X1_213/O PAND2X1_213/a_56_28# PAND2X1_213/CTRL2 PAND2X1_213/CTRL
+ PAND2X1_213/a_76_28# PAND2X1
XPAND2X1_235 VDD GND PAND2X1_85/Y POR2X1_62/Y POR2X1_243/B PAND2X1_235/a_16_344# PAND2X1_235/m4_208_n4#
+ PAND2X1_235/O PAND2X1_235/a_56_28# PAND2X1_235/CTRL2 PAND2X1_235/CTRL PAND2X1_235/a_76_28#
+ PAND2X1
XPAND2X1_224 VDD GND POR2X1_532/A PAND2X1_32/B POR2X1_227/B PAND2X1_224/a_16_344#
+ PAND2X1_224/m4_208_n4# PAND2X1_224/O PAND2X1_224/a_56_28# PAND2X1_224/CTRL2 PAND2X1_224/CTRL
+ PAND2X1_224/a_76_28# PAND2X1
XPAND2X1_268 VDD GND PAND2X1_93/B PAND2X1_69/A POR2X1_269/A PAND2X1_268/a_16_344#
+ PAND2X1_268/m4_208_n4# PAND2X1_268/O PAND2X1_268/a_56_28# PAND2X1_268/CTRL2 PAND2X1_268/CTRL
+ PAND2X1_268/a_76_28# PAND2X1
XPAND2X1_279 VDD GND POR2X1_614/A PAND2X1_57/B POR2X1_284/B PAND2X1_279/a_16_344#
+ PAND2X1_279/m4_208_n4# PAND2X1_279/O PAND2X1_279/a_56_28# PAND2X1_279/CTRL2 PAND2X1_279/CTRL
+ PAND2X1_279/a_76_28# PAND2X1
XPAND2X1_257 VDD GND POR2X1_614/A PAND2X1_20/A POR2X1_259/B PAND2X1_257/a_16_344#
+ PAND2X1_257/m4_208_n4# PAND2X1_257/O PAND2X1_257/a_56_28# PAND2X1_257/CTRL2 PAND2X1_257/CTRL
+ PAND2X1_257/a_76_28# PAND2X1
XPAND2X1_780 VDD GND POR2X1_744/Y POR2X1_743/Y PAND2X1_783/B PAND2X1_780/a_16_344#
+ PAND2X1_780/m4_208_n4# PAND2X1_780/O PAND2X1_780/a_56_28# PAND2X1_780/CTRL2 PAND2X1_780/CTRL
+ PAND2X1_780/a_76_28# PAND2X1
XPAND2X1_791 VDD GND POR2X1_757/Y POR2X1_755/Y PAND2X1_792/B PAND2X1_791/a_16_344#
+ PAND2X1_791/m4_208_n4# PAND2X1_791/O PAND2X1_791/a_56_28# PAND2X1_791/CTRL2 PAND2X1_791/CTRL
+ PAND2X1_791/a_76_28# PAND2X1
XPOR2X1_827 VDD GND POR2X1_42/Y POR2X1_416/B POR2X1_827/Y POR2X1_827/m4_208_n4# POR2X1_827/O
+ POR2X1_827/CTRL2 POR2X1_827/a_16_28# POR2X1_827/CTRL POR2X1_827/a_76_344# POR2X1_827/a_56_344#
+ POR2X1
XPOR2X1_816 VDD GND POR2X1_52/A POR2X1_816/A POR2X1_816/Y POR2X1_816/m4_208_n4# POR2X1_816/O
+ POR2X1_816/CTRL2 POR2X1_816/a_16_28# POR2X1_816/CTRL POR2X1_816/a_76_344# POR2X1_816/a_56_344#
+ POR2X1
XPOR2X1_805 VDD GND POR2X1_805/B POR2X1_805/A POR2X1_805/Y POR2X1_805/m4_208_n4# POR2X1_805/O
+ POR2X1_805/CTRL2 POR2X1_805/a_16_28# POR2X1_805/CTRL POR2X1_805/a_76_344# POR2X1_805/a_56_344#
+ POR2X1
XPOR2X1_838 VDD GND POR2X1_838/B POR2X1_837/Y POR2X1_852/B POR2X1_838/m4_208_n4# POR2X1_838/O
+ POR2X1_838/CTRL2 POR2X1_838/a_16_28# POR2X1_838/CTRL POR2X1_838/a_76_344# POR2X1_838/a_56_344#
+ POR2X1
XPOR2X1_849 VDD GND POR2X1_849/B POR2X1_849/A POR2X1_859/A POR2X1_849/m4_208_n4# POR2X1_849/O
+ POR2X1_849/CTRL2 POR2X1_849/a_16_28# POR2X1_849/CTRL POR2X1_849/a_76_344# POR2X1_849/a_56_344#
+ POR2X1
XPAND2X1_22 VDD GND PAND2X1_26/A PAND2X1_3/A PAND2X1_58/A PAND2X1_22/a_16_344# PAND2X1_22/m4_208_n4#
+ PAND2X1_22/O PAND2X1_22/a_56_28# PAND2X1_22/CTRL2 PAND2X1_22/CTRL PAND2X1_22/a_76_28#
+ PAND2X1
XPAND2X1_44 VDD GND PAND2X1_47/B PAND2X1_18/B PAND2X1_57/B PAND2X1_44/a_16_344# PAND2X1_44/m4_208_n4#
+ PAND2X1_44/O PAND2X1_44/a_56_28# PAND2X1_44/CTRL2 PAND2X1_44/CTRL PAND2X1_44/a_76_28#
+ PAND2X1
XPAND2X1_11 VDD GND INPUT_5 D_INPUT_4 PAND2X1_11/Y PAND2X1_11/a_16_344# PAND2X1_11/m4_208_n4#
+ PAND2X1_11/O PAND2X1_11/a_56_28# PAND2X1_11/CTRL2 PAND2X1_11/CTRL PAND2X1_11/a_76_28#
+ PAND2X1
XPAND2X1_33 VDD GND POR2X1_24/Y POR2X1_20/Y PAND2X1_35/A PAND2X1_33/a_16_344# PAND2X1_33/m4_208_n4#
+ PAND2X1_33/O PAND2X1_33/a_56_28# PAND2X1_33/CTRL2 PAND2X1_33/CTRL PAND2X1_33/a_76_28#
+ PAND2X1
XPAND2X1_66 VDD GND POR2X1_83/B POR2X1_7/B POR2X1_67/A PAND2X1_66/a_16_344# PAND2X1_66/m4_208_n4#
+ PAND2X1_66/O PAND2X1_66/a_56_28# PAND2X1_66/CTRL2 PAND2X1_66/CTRL PAND2X1_66/a_76_28#
+ PAND2X1
XPAND2X1_77 VDD GND POR2X1_94/A PAND2X1_94/A POR2X1_78/A PAND2X1_77/a_16_344# PAND2X1_77/m4_208_n4#
+ PAND2X1_77/O PAND2X1_77/a_56_28# PAND2X1_77/CTRL2 PAND2X1_77/CTRL PAND2X1_77/a_76_28#
+ PAND2X1
XPAND2X1_55 VDD GND POR2X1_94/A POR2X1_68/B PAND2X1_55/Y PAND2X1_55/a_16_344# PAND2X1_55/m4_208_n4#
+ PAND2X1_55/O PAND2X1_55/a_56_28# PAND2X1_55/CTRL2 PAND2X1_55/CTRL PAND2X1_55/a_76_28#
+ PAND2X1
XPAND2X1_99 VDD GND PAND2X1_99/B PAND2X1_97/Y PAND2X1_99/Y PAND2X1_99/a_16_344# PAND2X1_99/m4_208_n4#
+ PAND2X1_99/O PAND2X1_99/a_56_28# PAND2X1_99/CTRL2 PAND2X1_99/CTRL PAND2X1_99/a_76_28#
+ PAND2X1
XPOR2X1_19 VDD GND PAND2X1_6/A POR2X1_5/Y POR2X1_20/A POR2X1_19/m4_208_n4# POR2X1_19/O
+ POR2X1_19/CTRL2 POR2X1_19/a_16_28# POR2X1_19/CTRL POR2X1_19/a_76_344# POR2X1_19/a_56_344#
+ POR2X1
XPOR2X1_602 VDD GND POR2X1_602/B POR2X1_602/A POR2X1_788/A POR2X1_602/m4_208_n4# POR2X1_602/O
+ POR2X1_602/CTRL2 POR2X1_602/a_16_28# POR2X1_602/CTRL POR2X1_602/a_76_344# POR2X1_602/a_56_344#
+ POR2X1
XPAND2X1_88 VDD GND POR2X1_87/Y POR2X1_66/B PAND2X1_88/Y PAND2X1_88/a_16_344# PAND2X1_88/m4_208_n4#
+ PAND2X1_88/O PAND2X1_88/a_56_28# PAND2X1_88/CTRL2 PAND2X1_88/CTRL PAND2X1_88/a_76_28#
+ PAND2X1
XPOR2X1_624 VDD GND POR2X1_624/B POR2X1_623/Y POR2X1_624/Y POR2X1_624/m4_208_n4# POR2X1_624/O
+ POR2X1_624/CTRL2 POR2X1_624/a_16_28# POR2X1_624/CTRL POR2X1_624/a_76_344# POR2X1_624/a_56_344#
+ POR2X1
XPOR2X1_635 VDD GND POR2X1_635/B POR2X1_635/A POR2X1_635/Y POR2X1_635/m4_208_n4# POR2X1_635/O
+ POR2X1_635/CTRL2 POR2X1_635/a_16_28# POR2X1_635/CTRL POR2X1_635/a_76_344# POR2X1_635/a_56_344#
+ POR2X1
XPOR2X1_613 VDD GND POR2X1_40/Y POR2X1_55/Y POR2X1_613/Y POR2X1_613/m4_208_n4# POR2X1_613/O
+ POR2X1_613/CTRL2 POR2X1_613/a_16_28# POR2X1_613/CTRL POR2X1_613/a_76_344# POR2X1_613/a_56_344#
+ POR2X1
XPOR2X1_657 VDD GND POR2X1_141/Y POR2X1_510/Y POR2X1_657/Y POR2X1_657/m4_208_n4# POR2X1_657/O
+ POR2X1_657/CTRL2 POR2X1_657/a_16_28# POR2X1_657/CTRL POR2X1_657/a_76_344# POR2X1_657/a_56_344#
+ POR2X1
XPOR2X1_668 VDD GND POR2X1_66/A POR2X1_260/A POR2X1_668/Y POR2X1_668/m4_208_n4# POR2X1_668/O
+ POR2X1_668/CTRL2 POR2X1_668/a_16_28# POR2X1_668/CTRL POR2X1_668/a_76_344# POR2X1_668/a_56_344#
+ POR2X1
XPOR2X1_646 VDD GND POR2X1_646/B POR2X1_646/A POR2X1_646/Y POR2X1_646/m4_208_n4# POR2X1_646/O
+ POR2X1_646/CTRL2 POR2X1_646/a_16_28# POR2X1_646/CTRL POR2X1_646/a_76_344# POR2X1_646/a_56_344#
+ POR2X1
XPOR2X1_679 VDD GND POR2X1_679/B POR2X1_679/A POR2X1_679/Y POR2X1_679/m4_208_n4# POR2X1_679/O
+ POR2X1_679/CTRL2 POR2X1_679/a_16_28# POR2X1_679/CTRL POR2X1_679/a_76_344# POR2X1_679/a_56_344#
+ POR2X1
XPAND2X1_609 VDD GND POR2X1_608/Y PAND2X1_60/B POR2X1_646/A PAND2X1_609/a_16_344#
+ PAND2X1_609/m4_208_n4# PAND2X1_609/O PAND2X1_609/a_56_28# PAND2X1_609/CTRL2 PAND2X1_609/CTRL
+ PAND2X1_609/a_76_28# PAND2X1
XPOR2X1_410 VDD GND POR2X1_260/B PAND2X1_52/B POR2X1_410/Y POR2X1_410/m4_208_n4# POR2X1_410/O
+ POR2X1_410/CTRL2 POR2X1_410/a_16_28# POR2X1_410/CTRL POR2X1_410/a_76_344# POR2X1_410/a_56_344#
+ POR2X1
XPOR2X1_443 VDD GND POR2X1_97/A POR2X1_443/A POR2X1_444/A POR2X1_443/m4_208_n4# POR2X1_443/O
+ POR2X1_443/CTRL2 POR2X1_443/a_16_28# POR2X1_443/CTRL POR2X1_443/a_76_344# POR2X1_443/a_56_344#
+ POR2X1
XPOR2X1_432 VDD GND POR2X1_20/B POR2X1_129/Y POR2X1_432/Y POR2X1_432/m4_208_n4# POR2X1_432/O
+ POR2X1_432/CTRL2 POR2X1_432/a_16_28# POR2X1_432/CTRL POR2X1_432/a_76_344# POR2X1_432/a_56_344#
+ POR2X1
XPOR2X1_421 VDD GND POR2X1_90/Y POR2X1_329/A POR2X1_421/Y POR2X1_421/m4_208_n4# POR2X1_421/O
+ POR2X1_421/CTRL2 POR2X1_421/a_16_28# POR2X1_421/CTRL POR2X1_421/a_76_344# POR2X1_421/a_56_344#
+ POR2X1
XPOR2X1_465 VDD GND POR2X1_465/B POR2X1_465/A POR2X1_471/A POR2X1_465/m4_208_n4# POR2X1_465/O
+ POR2X1_465/CTRL2 POR2X1_465/a_16_28# POR2X1_465/CTRL POR2X1_465/a_76_344# POR2X1_465/a_56_344#
+ POR2X1
XPOR2X1_454 VDD GND POR2X1_454/B POR2X1_454/A POR2X1_466/A POR2X1_454/m4_208_n4# POR2X1_454/O
+ POR2X1_454/CTRL2 POR2X1_454/a_16_28# POR2X1_454/CTRL POR2X1_454/a_76_344# POR2X1_454/a_56_344#
+ POR2X1
XPOR2X1_487 VDD GND POR2X1_23/Y POR2X1_96/A POR2X1_487/Y POR2X1_487/m4_208_n4# POR2X1_487/O
+ POR2X1_487/CTRL2 POR2X1_487/a_16_28# POR2X1_487/CTRL POR2X1_487/a_76_344# POR2X1_487/a_56_344#
+ POR2X1
XPOR2X1_476 VDD GND POR2X1_472/Y POR2X1_476/A POR2X1_476/Y POR2X1_476/m4_208_n4# POR2X1_476/O
+ POR2X1_476/CTRL2 POR2X1_476/a_16_28# POR2X1_476/CTRL POR2X1_476/a_76_344# POR2X1_476/a_56_344#
+ POR2X1
XPOR2X1_498 VDD GND POR2X1_72/B POR2X1_498/A POR2X1_498/Y POR2X1_498/m4_208_n4# POR2X1_498/O
+ POR2X1_498/CTRL2 POR2X1_498/a_16_28# POR2X1_498/CTRL POR2X1_498/a_76_344# POR2X1_498/a_56_344#
+ POR2X1
XPAND2X1_417 VDD GND POR2X1_814/A PAND2X1_48/B POR2X1_446/B PAND2X1_417/a_16_344#
+ PAND2X1_417/m4_208_n4# PAND2X1_417/O PAND2X1_417/a_56_28# PAND2X1_417/CTRL2 PAND2X1_417/CTRL
+ PAND2X1_417/a_76_28# PAND2X1
XPAND2X1_406 VDD GND POR2X1_405/Y PAND2X1_96/B POR2X1_734/B PAND2X1_406/a_16_344#
+ PAND2X1_406/m4_208_n4# PAND2X1_406/O PAND2X1_406/a_56_28# PAND2X1_406/CTRL2 PAND2X1_406/CTRL
+ PAND2X1_406/a_76_28# PAND2X1
XPAND2X1_428 VDD GND POR2X1_383/A PAND2X1_32/B POR2X1_635/B PAND2X1_428/a_16_344#
+ PAND2X1_428/m4_208_n4# PAND2X1_428/O PAND2X1_428/a_56_28# PAND2X1_428/CTRL2 PAND2X1_428/CTRL
+ PAND2X1_428/a_76_28# PAND2X1
XPAND2X1_439 VDD GND POR2X1_438/Y POR2X1_177/Y PAND2X1_675/A PAND2X1_439/a_16_344#
+ PAND2X1_439/m4_208_n4# PAND2X1_439/O PAND2X1_439/a_56_28# PAND2X1_439/CTRL2 PAND2X1_439/CTRL
+ PAND2X1_439/a_76_28# PAND2X1
XPOR2X1_240 VDD GND POR2X1_240/B POR2X1_240/A POR2X1_243/A POR2X1_240/m4_208_n4# POR2X1_240/O
+ POR2X1_240/CTRL2 POR2X1_240/a_16_28# POR2X1_240/CTRL POR2X1_240/a_76_344# POR2X1_240/a_56_344#
+ POR2X1
XPOR2X1_251 VDD GND POR2X1_52/A POR2X1_251/A POR2X1_251/Y POR2X1_251/m4_208_n4# POR2X1_251/O
+ POR2X1_251/CTRL2 POR2X1_251/a_16_28# POR2X1_251/CTRL POR2X1_251/a_76_344# POR2X1_251/a_56_344#
+ POR2X1
XPOR2X1_262 VDD GND POR2X1_40/Y POR2X1_63/Y POR2X1_262/Y POR2X1_262/m4_208_n4# POR2X1_262/O
+ POR2X1_262/CTRL2 POR2X1_262/a_16_28# POR2X1_262/CTRL POR2X1_262/a_76_344# POR2X1_262/a_56_344#
+ POR2X1
XPOR2X1_273 VDD GND POR2X1_39/B POR2X1_153/Y POR2X1_273/Y POR2X1_273/m4_208_n4# POR2X1_273/O
+ POR2X1_273/CTRL2 POR2X1_273/a_16_28# POR2X1_273/CTRL POR2X1_273/a_76_344# POR2X1_273/a_56_344#
+ POR2X1
XPOR2X1_295 VDD GND POR2X1_60/A POR2X1_481/A POR2X1_295/Y POR2X1_295/m4_208_n4# POR2X1_295/O
+ POR2X1_295/CTRL2 POR2X1_295/a_16_28# POR2X1_295/CTRL POR2X1_295/a_76_344# POR2X1_295/a_56_344#
+ POR2X1
XPOR2X1_284 VDD GND POR2X1_284/B POR2X1_542/B POR2X1_287/A POR2X1_284/m4_208_n4# POR2X1_284/O
+ POR2X1_284/CTRL2 POR2X1_284/a_16_28# POR2X1_284/CTRL POR2X1_284/a_76_344# POR2X1_284/a_56_344#
+ POR2X1
XPAND2X1_203 VDD GND PAND2X1_76/Y POR2X1_72/Y PAND2X1_205/A PAND2X1_203/a_16_344#
+ PAND2X1_203/m4_208_n4# PAND2X1_203/O PAND2X1_203/a_56_28# PAND2X1_203/CTRL2 PAND2X1_203/CTRL
+ PAND2X1_203/a_76_28# PAND2X1
XPAND2X1_214 VDD GND PAND2X1_214/B PAND2X1_214/A PAND2X1_219/A PAND2X1_214/a_16_344#
+ PAND2X1_214/m4_208_n4# PAND2X1_214/O PAND2X1_214/a_56_28# PAND2X1_214/CTRL2 PAND2X1_214/CTRL
+ PAND2X1_214/a_76_28# PAND2X1
XPAND2X1_225 VDD GND POR2X1_68/B D_INPUT_1 POR2X1_814/A PAND2X1_225/a_16_344# PAND2X1_225/m4_208_n4#
+ PAND2X1_225/O PAND2X1_225/a_56_28# PAND2X1_225/CTRL2 PAND2X1_225/CTRL PAND2X1_225/a_76_28#
+ PAND2X1
XPAND2X1_236 VDD GND POR2X1_29/A POR2X1_68/B POR2X1_383/A PAND2X1_236/a_16_344# PAND2X1_236/m4_208_n4#
+ PAND2X1_236/O PAND2X1_236/a_56_28# PAND2X1_236/CTRL2 PAND2X1_236/CTRL PAND2X1_236/a_76_28#
+ PAND2X1
XPAND2X1_269 VDD GND POR2X1_268/Y POR2X1_236/Y POR2X1_271/B PAND2X1_269/a_16_344#
+ PAND2X1_269/m4_208_n4# PAND2X1_269/O PAND2X1_269/a_56_28# PAND2X1_269/CTRL2 PAND2X1_269/CTRL
+ PAND2X1_269/a_76_28# PAND2X1
XPAND2X1_247 VDD GND POR2X1_41/B POR2X1_7/A POR2X1_248/A PAND2X1_247/a_16_344# PAND2X1_247/m4_208_n4#
+ PAND2X1_247/O PAND2X1_247/a_56_28# PAND2X1_247/CTRL2 PAND2X1_247/CTRL PAND2X1_247/a_76_28#
+ PAND2X1
XPAND2X1_258 VDD GND POR2X1_260/A POR2X1_78/A POR2X1_259/A PAND2X1_258/a_16_344# PAND2X1_258/m4_208_n4#
+ PAND2X1_258/O PAND2X1_258/a_56_28# PAND2X1_258/CTRL2 PAND2X1_258/CTRL PAND2X1_258/a_76_28#
+ PAND2X1
XPAND2X1_770 VDD GND POR2X1_766/Y POR2X1_765/Y PAND2X1_771/B PAND2X1_770/a_16_344#
+ PAND2X1_770/m4_208_n4# PAND2X1_770/O PAND2X1_770/a_56_28# PAND2X1_770/CTRL2 PAND2X1_770/CTRL
+ PAND2X1_770/a_76_28# PAND2X1
XPAND2X1_781 VDD GND POR2X1_746/Y POR2X1_745/Y PAND2X1_781/Y PAND2X1_781/a_16_344#
+ PAND2X1_781/m4_208_n4# PAND2X1_781/O PAND2X1_781/a_56_28# PAND2X1_781/CTRL2 PAND2X1_781/CTRL
+ PAND2X1_781/a_76_28# PAND2X1
XPAND2X1_792 VDD GND PAND2X1_792/B POR2X1_759/Y PAND2X1_805/A PAND2X1_792/a_16_344#
+ PAND2X1_792/m4_208_n4# PAND2X1_792/O PAND2X1_792/a_56_28# PAND2X1_792/CTRL2 PAND2X1_792/CTRL
+ PAND2X1_792/a_76_28# PAND2X1
XPOR2X1_817 VDD GND INPUT_1 POR2X1_817/A POR2X1_817/Y POR2X1_817/m4_208_n4# POR2X1_817/O
+ POR2X1_817/CTRL2 POR2X1_817/a_16_28# POR2X1_817/CTRL POR2X1_817/a_76_344# POR2X1_817/a_56_344#
+ POR2X1
XPOR2X1_806 VDD GND POR2X1_362/B POR2X1_675/Y POR2X1_807/A POR2X1_806/m4_208_n4# POR2X1_806/O
+ POR2X1_806/CTRL2 POR2X1_806/a_16_28# POR2X1_806/CTRL POR2X1_806/a_76_344# POR2X1_806/a_56_344#
+ POR2X1
XPOR2X1_839 VDD GND POR2X1_835/Y POR2X1_836/Y POR2X1_852/A POR2X1_836/m4_208_n4# POR2X1_839/O
+ POR2X1_839/CTRL2 POR2X1_839/a_16_28# POR2X1_839/CTRL POR2X1_839/a_76_344# POR2X1_839/a_56_344#
+ POR2X1
XPOR2X1_828 VDD GND POR2X1_407/Y POR2X1_828/A POR2X1_828/Y POR2X1_808/m4_208_n4# POR2X1_828/O
+ POR2X1_828/CTRL2 POR2X1_828/a_16_28# POR2X1_828/CTRL POR2X1_828/a_76_344# POR2X1_828/a_56_344#
+ POR2X1
XPAND2X1_12 VDD GND PAND2X1_11/Y PAND2X1_3/A POR2X1_260/B PAND2X1_12/a_16_344# PAND2X1_12/m4_208_n4#
+ PAND2X1_12/O PAND2X1_12/a_56_28# PAND2X1_12/CTRL2 PAND2X1_12/CTRL PAND2X1_12/a_76_28#
+ PAND2X1
XPAND2X1_34 VDD GND POR2X1_32/Y POR2X1_27/Y PAND2X1_35/B PAND2X1_34/a_16_344# PAND2X1_34/m4_208_n4#
+ PAND2X1_34/O PAND2X1_34/a_56_28# PAND2X1_34/CTRL2 PAND2X1_34/CTRL PAND2X1_34/a_76_28#
+ PAND2X1
XPAND2X1_23 VDD GND PAND2X1_94/A PAND2X1_6/A PAND2X1_23/Y PAND2X1_23/a_16_344# PAND2X1_23/m4_208_n4#
+ PAND2X1_23/O PAND2X1_23/a_56_28# PAND2X1_23/CTRL2 PAND2X1_23/CTRL PAND2X1_23/a_76_28#
+ PAND2X1
XPAND2X1_56 VDD GND PAND2X1_55/Y PAND2X1_56/A PAND2X1_56/Y PAND2X1_56/a_16_344# PAND2X1_56/m4_208_n4#
+ PAND2X1_56/O PAND2X1_56/a_56_28# PAND2X1_56/CTRL2 PAND2X1_56/CTRL PAND2X1_56/a_76_28#
+ PAND2X1
XPAND2X1_45 VDD GND PAND2X1_57/B PAND2X1_23/Y POR2X1_702/B PAND2X1_45/a_16_344# PAND2X1_45/m4_208_n4#
+ PAND2X1_45/O PAND2X1_45/a_56_28# PAND2X1_45/CTRL2 PAND2X1_45/CTRL PAND2X1_45/a_76_28#
+ PAND2X1
XPAND2X1_67 VDD GND POR2X1_66/Y PAND2X1_55/Y POR2X1_202/B PAND2X1_67/a_16_344# PAND2X1_67/m4_208_n4#
+ PAND2X1_67/O PAND2X1_67/a_56_28# PAND2X1_67/CTRL2 PAND2X1_67/CTRL PAND2X1_67/a_76_28#
+ PAND2X1
XPAND2X1_78 VDD GND POR2X1_77/Y POR2X1_16/A POR2X1_79/A PAND2X1_78/a_16_344# PAND2X1_78/m4_208_n4#
+ PAND2X1_78/O PAND2X1_78/a_56_28# PAND2X1_78/CTRL2 PAND2X1_78/CTRL PAND2X1_78/a_76_28#
+ PAND2X1
XPAND2X1_89 VDD GND POR2X1_78/A PAND2X1_60/B POR2X1_97/B PAND2X1_89/a_16_344# PAND2X1_89/m4_208_n4#
+ PAND2X1_89/O PAND2X1_89/a_56_28# PAND2X1_89/CTRL2 PAND2X1_89/CTRL PAND2X1_89/a_76_28#
+ PAND2X1
XPOR2X1_603 VDD GND POR2X1_13/A POR2X1_49/Y POR2X1_603/Y POR2X1_603/m4_208_n4# POR2X1_603/O
+ POR2X1_603/CTRL2 POR2X1_603/a_16_28# POR2X1_603/CTRL POR2X1_603/a_76_344# POR2X1_603/a_56_344#
+ POR2X1
XPOR2X1_614 VDD GND POR2X1_78/A POR2X1_614/A POR2X1_614/Y POR2X1_614/m4_208_n4# POR2X1_614/O
+ POR2X1_614/CTRL2 POR2X1_614/a_16_28# POR2X1_614/CTRL POR2X1_614/a_76_344# POR2X1_614/a_56_344#
+ POR2X1
XPOR2X1_636 VDD GND POR2X1_636/B POR2X1_636/A POR2X1_639/A POR2X1_636/m4_208_n4# POR2X1_636/O
+ POR2X1_636/CTRL2 POR2X1_636/a_16_28# POR2X1_636/CTRL POR2X1_636/a_76_344# POR2X1_636/a_56_344#
+ POR2X1
XPOR2X1_625 VDD GND POR2X1_67/A POR2X1_293/Y POR2X1_625/Y POR2X1_625/m4_208_n4# POR2X1_625/O
+ POR2X1_625/CTRL2 POR2X1_625/a_16_28# POR2X1_625/CTRL POR2X1_625/a_76_344# POR2X1_625/a_56_344#
+ POR2X1
XPOR2X1_669 VDD GND POR2X1_669/B POR2X1_669/A POR2X1_669/Y POR2X1_669/m4_208_n4# POR2X1_669/O
+ POR2X1_669/CTRL2 POR2X1_669/a_16_28# POR2X1_669/CTRL POR2X1_669/a_76_344# POR2X1_669/a_56_344#
+ POR2X1
XPOR2X1_658 VDD GND POR2X1_624/Y POR2X1_632/Y POR2X1_659/A POR2X1_658/m4_208_n4# POR2X1_658/O
+ POR2X1_658/CTRL2 POR2X1_658/a_16_28# POR2X1_658/CTRL POR2X1_658/a_76_344# POR2X1_658/a_56_344#
+ POR2X1
XPOR2X1_647 VDD GND POR2X1_647/B POR2X1_646/Y POR2X1_647/Y POR2X1_647/m4_208_n4# POR2X1_647/O
+ POR2X1_647/CTRL2 POR2X1_647/a_16_28# POR2X1_647/CTRL POR2X1_647/a_76_344# POR2X1_647/a_56_344#
+ POR2X1
XPOR2X1_400 VDD GND POR2X1_400/B POR2X1_400/A POR2X1_403/A POR2X1_400/m4_208_n4# POR2X1_400/O
+ POR2X1_400/CTRL2 POR2X1_400/a_16_28# POR2X1_400/CTRL POR2X1_400/a_76_344# POR2X1_400/a_56_344#
+ POR2X1
XPOR2X1_411 VDD GND POR2X1_411/B POR2X1_411/A POR2X1_411/Y POR2X1_411/m4_208_n4# POR2X1_411/O
+ POR2X1_411/CTRL2 POR2X1_411/a_16_28# POR2X1_411/CTRL POR2X1_411/a_76_344# POR2X1_411/a_56_344#
+ POR2X1
XPOR2X1_444 VDD GND POR2X1_444/B POR2X1_444/A POR2X1_444/Y POR2X1_444/m4_208_n4# POR2X1_444/O
+ POR2X1_444/CTRL2 POR2X1_444/a_16_28# POR2X1_444/CTRL POR2X1_444/a_76_344# POR2X1_444/a_56_344#
+ POR2X1
XPOR2X1_422 VDD GND POR2X1_13/A POR2X1_93/A POR2X1_422/Y POR2X1_422/m4_208_n4# POR2X1_422/O
+ POR2X1_422/CTRL2 POR2X1_422/a_16_28# POR2X1_422/CTRL POR2X1_422/a_76_344# POR2X1_422/a_56_344#
+ POR2X1
XPOR2X1_433 VDD GND POR2X1_72/B POR2X1_153/Y POR2X1_433/Y POR2X1_433/m4_208_n4# POR2X1_433/O
+ POR2X1_433/CTRL2 POR2X1_433/a_16_28# POR2X1_433/CTRL POR2X1_433/a_76_344# POR2X1_433/a_56_344#
+ POR2X1
XPOR2X1_455 VDD GND POR2X1_76/Y POR2X1_455/A POR2X1_465/B POR2X1_455/m4_208_n4# POR2X1_455/O
+ POR2X1_455/CTRL2 POR2X1_455/a_16_28# POR2X1_455/CTRL POR2X1_455/a_76_344# POR2X1_455/a_56_344#
+ POR2X1
XPOR2X1_466 VDD GND POR2X1_453/Y POR2X1_466/A POR2X1_466/Y POR2X1_466/m4_208_n4# POR2X1_466/O
+ POR2X1_466/CTRL2 POR2X1_466/a_16_28# POR2X1_466/CTRL POR2X1_466/a_76_344# POR2X1_466/a_56_344#
+ POR2X1
XPOR2X1_477 VDD GND POR2X1_477/B POR2X1_477/A POR2X1_477/Y POR2X1_477/m4_208_n4# POR2X1_477/O
+ POR2X1_477/CTRL2 POR2X1_477/a_16_28# POR2X1_477/CTRL POR2X1_477/a_76_344# POR2X1_477/a_56_344#
+ POR2X1
XPOR2X1_499 VDD GND POR2X1_833/A POR2X1_499/A POR2X1_500/A POR2X1_499/m4_208_n4# POR2X1_499/O
+ POR2X1_499/CTRL2 POR2X1_499/a_16_28# POR2X1_499/CTRL POR2X1_499/a_76_344# POR2X1_499/a_56_344#
+ POR2X1
XPOR2X1_488 VDD GND POR2X1_416/B POR2X1_283/A POR2X1_488/Y POR2X1_488/m4_208_n4# POR2X1_488/O
+ POR2X1_488/CTRL2 POR2X1_488/a_16_28# POR2X1_488/CTRL POR2X1_488/a_76_344# POR2X1_488/a_56_344#
+ POR2X1
XPAND2X1_418 VDD GND PAND2X1_52/B POR2X1_78/B POR2X1_446/A PAND2X1_418/a_16_344# PAND2X1_418/m4_208_n4#
+ PAND2X1_418/O PAND2X1_418/a_56_28# PAND2X1_418/CTRL2 PAND2X1_418/CTRL PAND2X1_418/a_76_28#
+ PAND2X1
XPAND2X1_407 VDD GND POR2X1_153/Y POR2X1_55/Y POR2X1_409/B PAND2X1_407/a_16_344# PAND2X1_407/m4_208_n4#
+ PAND2X1_407/O PAND2X1_407/a_56_28# PAND2X1_407/CTRL2 PAND2X1_407/CTRL PAND2X1_407/a_76_28#
+ PAND2X1
XPAND2X1_429 VDD GND PAND2X1_11/Y D_INPUT_7 PAND2X1_429/Y PAND2X1_429/a_16_344# PAND2X1_429/m4_208_n4#
+ PAND2X1_429/O PAND2X1_429/a_56_28# PAND2X1_429/CTRL2 PAND2X1_429/CTRL PAND2X1_429/a_76_28#
+ PAND2X1
XPOR2X1_241 VDD GND POR2X1_241/B POR2X1_776/A POR2X1_241/Y POR2X1_241/m4_208_n4# POR2X1_241/O
+ POR2X1_241/CTRL2 POR2X1_241/a_16_28# POR2X1_241/CTRL POR2X1_241/a_76_344# POR2X1_241/a_56_344#
+ POR2X1
XPOR2X1_230 VDD GND POR2X1_7/A POR2X1_32/A POR2X1_230/Y POR2X1_230/m4_208_n4# POR2X1_230/O
+ POR2X1_230/CTRL2 POR2X1_230/a_16_28# POR2X1_230/CTRL POR2X1_230/a_76_344# POR2X1_230/a_56_344#
+ POR2X1
XPOR2X1_252 VDD GND POR2X1_55/Y POR2X1_60/A POR2X1_252/Y POR2X1_252/m4_208_n4# POR2X1_252/O
+ POR2X1_252/CTRL2 POR2X1_252/a_16_28# POR2X1_252/CTRL POR2X1_252/a_76_344# POR2X1_252/a_56_344#
+ POR2X1
XPOR2X1_263 VDD GND POR2X1_43/B POR2X1_37/Y POR2X1_263/Y POR2X1_63/m4_208_n4# POR2X1_263/O
+ POR2X1_263/CTRL2 POR2X1_263/a_16_28# POR2X1_263/CTRL POR2X1_263/a_76_344# POR2X1_263/a_56_344#
+ POR2X1
XPOR2X1_274 VDD GND POR2X1_274/B POR2X1_274/A POR2X1_274/Y POR2X1_274/m4_208_n4# POR2X1_274/O
+ POR2X1_274/CTRL2 POR2X1_274/a_16_28# POR2X1_274/CTRL POR2X1_274/a_76_344# POR2X1_274/a_56_344#
+ POR2X1
XPOR2X1_285 VDD GND POR2X1_285/B POR2X1_285/A POR2X1_285/Y POR2X1_285/m4_208_n4# POR2X1_285/O
+ POR2X1_285/CTRL2 POR2X1_285/a_16_28# POR2X1_285/CTRL POR2X1_285/a_76_344# POR2X1_285/a_56_344#
+ POR2X1
XPOR2X1_296 VDD GND POR2X1_296/B PAND2X1_55/Y POR2X1_296/Y POR2X1_296/m4_208_n4# POR2X1_296/O
+ POR2X1_296/CTRL2 POR2X1_296/a_16_28# POR2X1_296/CTRL POR2X1_296/a_76_344# POR2X1_296/a_56_344#
+ POR2X1
XPAND2X1_237 VDD GND POR2X1_383/A POR2X1_66/A POR2X1_241/B PAND2X1_237/a_16_344# POR2X1_351/m4_208_n4#
+ PAND2X1_237/O PAND2X1_237/a_56_28# PAND2X1_237/CTRL2 PAND2X1_237/CTRL PAND2X1_237/a_76_28#
+ PAND2X1
XPAND2X1_215 VDD GND PAND2X1_215/B PAND2X1_205/Y PAND2X1_219/B PAND2X1_215/a_16_344#
+ POR2X1_385/m4_208_n4# PAND2X1_215/O PAND2X1_215/a_56_28# PAND2X1_215/CTRL2 PAND2X1_215/CTRL
+ PAND2X1_215/a_76_28# PAND2X1
XPAND2X1_204 VDD GND PAND2X1_84/Y POR2X1_79/Y PAND2X1_205/B PAND2X1_204/a_16_344#
+ POR2X1_679/m4_208_n4# PAND2X1_204/O PAND2X1_204/a_56_28# PAND2X1_204/CTRL2 PAND2X1_204/CTRL
+ PAND2X1_204/a_76_28# PAND2X1
XPAND2X1_226 VDD GND POR2X1_814/A PAND2X1_20/A POR2X1_227/A PAND2X1_226/a_16_344#
+ PAND2X1_226/m4_208_n4# PAND2X1_226/O PAND2X1_226/a_56_28# PAND2X1_226/CTRL2 PAND2X1_226/CTRL
+ PAND2X1_226/a_76_28# PAND2X1
XPAND2X1_259 VDD GND POR2X1_258/Y POR2X1_257/Y PAND2X1_555/A PAND2X1_259/a_16_344#
+ PAND2X1_259/m4_208_n4# PAND2X1_259/O PAND2X1_259/a_56_28# PAND2X1_259/CTRL2 PAND2X1_259/CTRL
+ PAND2X1_259/a_76_28# PAND2X1
XPAND2X1_248 VDD GND POR2X1_247/Y PAND2X1_48/B POR2X1_342/A PAND2X1_248/a_16_344#
+ PAND2X1_248/m4_208_n4# PAND2X1_248/O PAND2X1_248/a_56_28# PAND2X1_248/CTRL2 PAND2X1_248/CTRL
+ PAND2X1_248/a_76_28# PAND2X1
XPAND2X1_760 VDD GND POR2X1_327/Y PAND2X1_65/B POR2X1_800/A PAND2X1_760/a_16_344#
+ PAND2X1_760/m4_208_n4# PAND2X1_760/O PAND2X1_760/a_56_28# PAND2X1_760/CTRL2 PAND2X1_760/CTRL
+ PAND2X1_760/a_76_28# PAND2X1
XPAND2X1_771 VDD GND PAND2X1_771/B PAND2X1_769/Y PAND2X1_771/Y PAND2X1_771/a_16_344#
+ PAND2X1_771/m4_208_n4# PAND2X1_771/O PAND2X1_771/a_56_28# PAND2X1_771/CTRL2 PAND2X1_771/CTRL
+ PAND2X1_771/a_76_28# PAND2X1
XPAND2X1_782 VDD GND PAND2X1_781/Y POR2X1_747/Y PAND2X1_782/Y PAND2X1_782/a_16_344#
+ PAND2X1_782/m4_208_n4# PAND2X1_782/O PAND2X1_782/a_56_28# PAND2X1_782/CTRL2 PAND2X1_782/CTRL
+ PAND2X1_782/a_76_28# PAND2X1
XPAND2X1_793 VDD GND PAND2X1_790/Y PAND2X1_793/A PAND2X1_793/Y PAND2X1_793/a_16_344#
+ PAND2X1_793/m4_208_n4# PAND2X1_793/O PAND2X1_793/a_56_28# PAND2X1_793/CTRL2 PAND2X1_793/CTRL
+ PAND2X1_793/a_76_28# PAND2X1
XPAND2X1_590 VDD GND POR2X1_102/Y POR2X1_38/Y POR2X1_591/A PAND2X1_590/a_16_344# PAND2X1_590/m4_208_n4#
+ PAND2X1_590/O PAND2X1_590/a_56_28# PAND2X1_590/CTRL2 PAND2X1_590/CTRL PAND2X1_590/a_76_28#
+ PAND2X1
XPOR2X1_818 VDD GND POR2X1_68/B POR2X1_502/A POR2X1_818/Y POR2X1_818/m4_208_n4# POR2X1_818/O
+ POR2X1_818/CTRL2 POR2X1_818/a_16_28# POR2X1_818/CTRL POR2X1_818/a_76_344# POR2X1_818/a_56_344#
+ POR2X1
XPOR2X1_807 VDD GND POR2X1_805/Y POR2X1_807/A POR2X1_811/B POR2X1_807/m4_208_n4# POR2X1_807/O
+ POR2X1_807/CTRL2 POR2X1_807/a_16_28# POR2X1_807/CTRL POR2X1_807/a_76_344# POR2X1_807/a_56_344#
+ POR2X1
XPOR2X1_829 VDD GND POR2X1_65/A POR2X1_829/A POR2X1_829/Y POR2X1_829/m4_208_n4# POR2X1_829/O
+ POR2X1_829/CTRL2 POR2X1_829/a_16_28# POR2X1_829/CTRL POR2X1_829/a_76_344# POR2X1_829/a_56_344#
+ POR2X1
XPAND2X1_13 VDD GND POR2X1_260/B POR2X1_294/B POR2X1_193/A PAND2X1_13/a_16_344# PAND2X1_13/m4_208_n4#
+ PAND2X1_13/O PAND2X1_13/a_56_28# PAND2X1_13/CTRL2 PAND2X1_13/CTRL PAND2X1_13/a_76_28#
+ PAND2X1
XPAND2X1_35 VDD GND PAND2X1_35/B PAND2X1_35/A PAND2X1_35/Y PAND2X1_35/a_16_344# PAND2X1_35/m4_208_n4#
+ PAND2X1_35/O PAND2X1_35/a_56_28# PAND2X1_35/CTRL2 PAND2X1_35/CTRL PAND2X1_35/a_76_28#
+ PAND2X1
XPAND2X1_24 VDD GND PAND2X1_23/Y PAND2X1_58/A POR2X1_33/A PAND2X1_24/a_16_344# PAND2X1_24/m4_208_n4#
+ PAND2X1_24/O PAND2X1_24/a_56_28# PAND2X1_24/CTRL2 PAND2X1_24/CTRL PAND2X1_24/a_76_28#
+ PAND2X1
XPAND2X1_68 VDD GND POR2X1_49/Y POR2X1_5/Y POR2X1_69/A PAND2X1_68/a_16_344# PAND2X1_68/m4_208_n4#
+ PAND2X1_68/O PAND2X1_68/a_56_28# PAND2X1_68/CTRL2 PAND2X1_68/CTRL PAND2X1_68/a_76_28#
+ PAND2X1
XPAND2X1_46 VDD GND PAND2X1_94/A D_INPUT_1 PAND2X1_48/A PAND2X1_46/a_16_344# PAND2X1_46/m4_208_n4#
+ PAND2X1_46/O PAND2X1_46/a_56_28# PAND2X1_46/CTRL2 PAND2X1_46/CTRL PAND2X1_46/a_76_28#
+ PAND2X1
XPAND2X1_57 VDD GND PAND2X1_57/B POR2X1_68/B POR2X1_198/B PAND2X1_57/a_16_344# PAND2X1_57/m4_208_n4#
+ PAND2X1_57/O PAND2X1_57/a_56_28# PAND2X1_57/CTRL2 PAND2X1_57/CTRL PAND2X1_57/a_76_28#
+ PAND2X1
XPAND2X1_79 VDD GND POR2X1_78/Y PAND2X1_20/A PAND2X1_79/Y PAND2X1_79/a_16_344# PAND2X1_79/m4_208_n4#
+ PAND2X1_79/O PAND2X1_79/a_56_28# PAND2X1_79/CTRL2 PAND2X1_79/CTRL PAND2X1_79/a_76_28#
+ PAND2X1
XPOR2X1_604 VDD GND POR2X1_72/B POR2X1_669/B POR2X1_604/Y POR2X1_604/m4_208_n4# POR2X1_604/O
+ POR2X1_604/CTRL2 POR2X1_604/a_16_28# POR2X1_604/CTRL POR2X1_604/a_76_344# POR2X1_604/a_56_344#
+ POR2X1
XPOR2X1_626 VDD GND POR2X1_96/A POR2X1_669/B POR2X1_626/Y POR2X1_626/m4_208_n4# POR2X1_626/O
+ POR2X1_626/CTRL2 POR2X1_626/a_16_28# POR2X1_626/CTRL POR2X1_626/a_76_344# POR2X1_626/a_56_344#
+ POR2X1
XPOR2X1_615 VDD GND POR2X1_43/B POR2X1_754/A POR2X1_615/Y POR2X1_615/m4_208_n4# POR2X1_615/O
+ POR2X1_615/CTRL2 POR2X1_615/a_16_28# POR2X1_615/CTRL POR2X1_615/a_76_344# POR2X1_615/a_56_344#
+ POR2X1
XPOR2X1_659 VDD GND POR2X1_657/Y POR2X1_659/A POR2X1_663/B POR2X1_659/m4_208_n4# POR2X1_659/O
+ POR2X1_659/CTRL2 POR2X1_659/a_16_28# POR2X1_659/CTRL POR2X1_659/a_76_344# POR2X1_659/a_56_344#
+ POR2X1
XPOR2X1_648 VDD GND POR2X1_644/Y POR2X1_648/A POR2X1_648/Y POR2X1_648/m4_208_n4# POR2X1_648/O
+ POR2X1_648/CTRL2 POR2X1_648/a_16_28# POR2X1_648/CTRL POR2X1_648/a_76_344# POR2X1_648/a_56_344#
+ POR2X1
XPOR2X1_637 VDD GND POR2X1_637/B POR2X1_637/A POR2X1_638/A POR2X1_637/m4_208_n4# POR2X1_637/O
+ POR2X1_637/CTRL2 POR2X1_637/a_16_28# POR2X1_637/CTRL POR2X1_637/a_76_344# POR2X1_637/a_56_344#
+ POR2X1
XPOR2X1_401 VDD GND POR2X1_401/B POR2X1_401/A POR2X1_402/A POR2X1_401/m4_208_n4# POR2X1_401/O
+ POR2X1_401/CTRL2 POR2X1_401/a_16_28# POR2X1_401/CTRL POR2X1_401/a_76_344# POR2X1_401/a_56_344#
+ POR2X1
XPOR2X1_412 VDD GND POR2X1_37/Y POR2X1_57/A POR2X1_413/A POR2X1_412/m4_208_n4# POR2X1_412/O
+ POR2X1_412/CTRL2 POR2X1_412/a_16_28# POR2X1_412/CTRL POR2X1_412/a_76_344# POR2X1_412/a_56_344#
+ POR2X1
XPOR2X1_434 VDD GND POR2X1_174/A POR2X1_434/A POR2X1_436/B POR2X1_434/m4_208_n4# POR2X1_434/O
+ POR2X1_434/CTRL2 POR2X1_434/a_16_28# POR2X1_434/CTRL POR2X1_434/a_76_344# POR2X1_434/a_56_344#
+ POR2X1
XPOR2X1_423 VDD GND POR2X1_7/A POR2X1_65/A POR2X1_423/Y POR2X1_423/m4_208_n4# POR2X1_423/O
+ POR2X1_423/CTRL2 POR2X1_423/a_16_28# POR2X1_423/CTRL POR2X1_423/a_76_344# POR2X1_423/a_56_344#
+ POR2X1
XPOR2X1_456 VDD GND POR2X1_456/B POR2X1_254/Y POR2X1_465/A POR2X1_456/m4_208_n4# POR2X1_456/O
+ POR2X1_456/CTRL2 POR2X1_456/a_16_28# POR2X1_456/CTRL POR2X1_456/a_76_344# POR2X1_456/a_56_344#
+ POR2X1
XPOR2X1_445 VDD GND POR2X1_241/B POR2X1_445/A POR2X1_455/A POR2X1_445/m4_208_n4# POR2X1_445/O
+ POR2X1_445/CTRL2 POR2X1_445/a_16_28# POR2X1_445/CTRL POR2X1_445/a_76_344# POR2X1_445/a_56_344#
+ POR2X1
XPOR2X1_467 VDD GND POR2X1_210/A POR2X1_452/Y POR2X1_467/Y POR2X1_467/m4_208_n4# POR2X1_467/O
+ POR2X1_467/CTRL2 POR2X1_467/a_16_28# POR2X1_467/CTRL POR2X1_467/a_76_344# POR2X1_467/a_56_344#
+ POR2X1
XPOR2X1_478 VDD GND POR2X1_478/B POR2X1_477/Y POR2X1_478/Y POR2X1_478/m4_208_n4# POR2X1_478/O
+ POR2X1_478/CTRL2 POR2X1_478/a_16_28# POR2X1_478/CTRL POR2X1_478/a_76_344# POR2X1_478/a_56_344#
+ POR2X1
XPOR2X1_489 VDD GND POR2X1_489/B POR2X1_489/A POR2X1_557/B POR2X1_489/m4_208_n4# POR2X1_489/O
+ POR2X1_489/CTRL2 POR2X1_489/a_16_28# POR2X1_489/CTRL POR2X1_489/a_76_344# POR2X1_489/a_56_344#
+ POR2X1
XPAND2X1_408 VDD GND PAND2X1_26/A D_INPUT_6 PAND2X1_408/Y PAND2X1_408/a_16_344# PAND2X1_408/m4_208_n4#
+ PAND2X1_408/O PAND2X1_408/a_56_28# PAND2X1_408/CTRL2 PAND2X1_408/CTRL PAND2X1_408/a_76_28#
+ PAND2X1
XPAND2X1_419 VDD GND POR2X1_296/B PAND2X1_69/A POR2X1_447/B PAND2X1_419/a_16_344#
+ PAND2X1_419/m4_208_n4# PAND2X1_419/O PAND2X1_419/a_56_28# PAND2X1_419/CTRL2 PAND2X1_419/CTRL
+ PAND2X1_419/a_76_28# PAND2X1
XPOR2X1_242 VDD GND POR2X1_506/B POR2X1_241/Y POR2X1_244/B POR2X1_242/m4_208_n4# POR2X1_242/O
+ POR2X1_242/CTRL2 POR2X1_242/a_16_28# POR2X1_242/CTRL POR2X1_242/a_76_344# POR2X1_242/a_56_344#
+ POR2X1
XPOR2X1_231 VDD GND POR2X1_231/B POR2X1_231/A POR2X1_341/A POR2X1_231/m4_208_n4# POR2X1_231/O
+ POR2X1_231/CTRL2 POR2X1_231/a_16_28# POR2X1_231/CTRL POR2X1_231/a_76_344# POR2X1_231/a_56_344#
+ POR2X1
XPOR2X1_220 VDD GND POR2X1_220/B POR2X1_220/A POR2X1_220/Y POR2X1_220/m4_208_n4# POR2X1_220/O
+ POR2X1_220/CTRL2 POR2X1_220/a_16_28# POR2X1_220/CTRL POR2X1_220/a_76_344# POR2X1_220/a_56_344#
+ POR2X1
XPOR2X1_264 VDD GND POR2X1_294/B POR2X1_78/A POR2X1_264/Y POR2X1_264/m4_208_n4# POR2X1_264/O
+ POR2X1_264/CTRL2 POR2X1_264/a_16_28# POR2X1_264/CTRL POR2X1_264/a_76_344# POR2X1_264/a_56_344#
+ POR2X1
XPOR2X1_275 VDD GND INPUT_0 POR2X1_275/A POR2X1_275/Y POR2X1_275/m4_208_n4# POR2X1_275/O
+ POR2X1_275/CTRL2 POR2X1_275/a_16_28# POR2X1_275/CTRL POR2X1_275/a_76_344# POR2X1_275/a_56_344#
+ POR2X1
XPOR2X1_253 VDD GND POR2X1_65/A POR2X1_257/A POR2X1_253/Y POR2X1_56/m4_208_n4# POR2X1_253/O
+ POR2X1_253/CTRL2 POR2X1_253/a_16_28# POR2X1_253/CTRL POR2X1_253/a_76_344# POR2X1_253/a_56_344#
+ POR2X1
XPOR2X1_286 VDD GND POR2X1_286/B POR2X1_285/Y POR2X1_286/Y POR2X1_286/m4_208_n4# POR2X1_286/O
+ POR2X1_286/CTRL2 POR2X1_286/a_16_28# POR2X1_286/CTRL POR2X1_286/a_76_344# POR2X1_286/a_56_344#
+ POR2X1
XPOR2X1_297 VDD GND POR2X1_57/A POR2X1_297/A POR2X1_297/Y POR2X1_297/m4_208_n4# POR2X1_297/O
+ POR2X1_297/CTRL2 POR2X1_297/a_16_28# POR2X1_297/CTRL POR2X1_297/a_76_344# POR2X1_297/a_56_344#
+ POR2X1
XPAND2X1_216 VDD GND PAND2X1_216/B PAND2X1_656/A PAND2X1_218/A PAND2X1_216/a_16_344#
+ PAND2X1_216/m4_208_n4# PAND2X1_216/O PAND2X1_216/a_56_28# PAND2X1_216/CTRL2 PAND2X1_216/CTRL
+ PAND2X1_216/a_76_28# PAND2X1
XPAND2X1_227 VDD GND POR2X1_226/Y POR2X1_224/Y PAND2X1_340/B PAND2X1_227/a_16_344#
+ POR2X1_503/m4_208_n4# PAND2X1_227/O PAND2X1_227/a_56_28# PAND2X1_227/CTRL2 PAND2X1_227/CTRL
+ PAND2X1_227/a_76_28# PAND2X1
XPAND2X1_205 VDD GND PAND2X1_205/B PAND2X1_205/A PAND2X1_205/Y PAND2X1_205/a_16_344#
+ PAND2X1_205/m4_208_n4# PAND2X1_205/O PAND2X1_205/a_56_28# PAND2X1_205/CTRL2 PAND2X1_205/CTRL
+ PAND2X1_205/a_76_28# PAND2X1
XPAND2X1_249 VDD GND POR2X1_38/Y POR2X1_23/Y POR2X1_250/A PAND2X1_249/a_16_344# PAND2X1_249/m4_208_n4#
+ PAND2X1_249/O PAND2X1_249/a_56_28# PAND2X1_249/CTRL2 PAND2X1_249/CTRL PAND2X1_249/a_76_28#
+ PAND2X1
XPAND2X1_238 VDD GND PAND2X1_52/B PAND2X1_23/Y POR2X1_776/A PAND2X1_238/a_16_344#
+ POR2X1_241/m4_208_n4# PAND2X1_238/O PAND2X1_238/a_56_28# PAND2X1_238/CTRL2 PAND2X1_238/CTRL
+ PAND2X1_238/a_76_28# PAND2X1
XPAND2X1_750 VDD GND POR2X1_749/Y POR2X1_669/B POR2X1_751/A PAND2X1_750/a_16_344#
+ PAND2X1_750/m4_208_n4# PAND2X1_750/O PAND2X1_750/a_56_28# PAND2X1_750/CTRL2 PAND2X1_750/CTRL
+ PAND2X1_750/a_76_28# PAND2X1
XPAND2X1_772 VDD GND PAND2X1_768/Y PAND2X1_557/A PAND2X1_773/B PAND2X1_772/a_16_344#
+ PAND2X1_772/m4_208_n4# PAND2X1_772/O PAND2X1_772/a_56_28# PAND2X1_772/CTRL2 PAND2X1_772/CTRL
+ PAND2X1_772/a_76_28# PAND2X1
XPAND2X1_783 VDD GND PAND2X1_783/B PAND2X1_779/Y PAND2X1_783/Y PAND2X1_783/a_16_344#
+ PAND2X1_783/m4_208_n4# PAND2X1_783/O PAND2X1_783/a_56_28# PAND2X1_783/CTRL2 PAND2X1_783/CTRL
+ PAND2X1_783/a_76_28# PAND2X1
XPAND2X1_761 VDD GND POR2X1_644/A D_INPUT_0 POR2X1_801/B PAND2X1_761/a_16_344# PAND2X1_761/m4_208_n4#
+ PAND2X1_761/O PAND2X1_761/a_56_28# PAND2X1_761/CTRL2 PAND2X1_761/CTRL PAND2X1_761/a_76_28#
+ PAND2X1
XPAND2X1_794 VDD GND PAND2X1_794/B PAND2X1_787/Y PAND2X1_804/A PAND2X1_794/a_16_344#
+ PAND2X1_794/m4_208_n4# PAND2X1_794/O PAND2X1_794/a_56_28# PAND2X1_794/CTRL2 PAND2X1_794/CTRL
+ PAND2X1_794/a_76_28# PAND2X1
XPAND2X1_580 VDD GND PAND2X1_580/B PAND2X1_578/Y GATE_579 PAND2X1_580/a_16_344# PAND2X1_580/m4_208_n4#
+ PAND2X1_580/O PAND2X1_580/a_56_28# PAND2X1_580/CTRL2 PAND2X1_580/CTRL PAND2X1_580/a_76_28#
+ PAND2X1
XPAND2X1_591 VDD GND POR2X1_590/Y PAND2X1_65/B POR2X1_593/B PAND2X1_591/a_16_344#
+ PAND2X1_591/m4_208_n4# PAND2X1_591/O PAND2X1_591/a_56_28# PAND2X1_591/CTRL2 PAND2X1_591/CTRL
+ PAND2X1_591/a_76_28# PAND2X1
XPOR2X1_808 VDD GND POR2X1_808/B POR2X1_808/A POR2X1_811/A POR2X1_808/m4_208_n4# POR2X1_808/O
+ POR2X1_808/CTRL2 POR2X1_808/a_16_28# POR2X1_808/CTRL POR2X1_808/a_76_344# POR2X1_808/a_56_344#
+ POR2X1
XPOR2X1_819 VDD GND POR2X1_48/A POR2X1_94/A POR2X1_820/A POR2X1_819/m4_208_n4# POR2X1_819/O
+ POR2X1_819/CTRL2 POR2X1_819/a_16_28# POR2X1_819/CTRL POR2X1_819/a_76_344# POR2X1_819/a_56_344#
+ POR2X1
XPAND2X1_25 VDD GND D_INPUT_7 INPUT_6 PAND2X1_59/B PAND2X1_25/a_16_344# PAND2X1_25/m4_208_n4#
+ PAND2X1_25/O PAND2X1_25/a_56_28# PAND2X1_25/CTRL2 PAND2X1_25/CTRL PAND2X1_25/a_76_28#
+ PAND2X1
XPAND2X1_14 VDD GND D_INPUT_3 D_INPUT_2 PAND2X1_94/A PAND2X1_14/a_16_344# PAND2X1_14/m4_208_n4#
+ PAND2X1_14/O PAND2X1_14/a_56_28# PAND2X1_14/CTRL2 PAND2X1_14/CTRL PAND2X1_14/a_76_28#
+ PAND2X1
XPAND2X1_47 VDD GND PAND2X1_47/B PAND2X1_59/B PAND2X1_48/B PAND2X1_47/a_16_344# PAND2X1_47/m4_208_n4#
+ PAND2X1_47/O PAND2X1_47/a_56_28# PAND2X1_47/CTRL2 PAND2X1_47/CTRL PAND2X1_47/a_76_28#
+ PAND2X1
XPAND2X1_36 VDD GND PAND2X1_26/A PAND2X1_18/B PAND2X1_69/A PAND2X1_36/a_16_344# PAND2X1_36/m4_208_n4#
+ PAND2X1_36/O PAND2X1_36/a_56_28# PAND2X1_36/CTRL2 PAND2X1_36/CTRL PAND2X1_36/a_76_28#
+ PAND2X1
XPAND2X1_58 VDD GND POR2X1_68/A PAND2X1_58/A POR2X1_61/B PAND2X1_58/a_16_344# PAND2X1_58/m4_208_n4#
+ PAND2X1_58/O PAND2X1_58/a_56_28# PAND2X1_58/CTRL2 PAND2X1_58/CTRL PAND2X1_58/a_76_28#
+ PAND2X1
XPAND2X1_69 VDD GND POR2X1_68/Y PAND2X1_69/A POR2X1_202/A PAND2X1_69/a_16_344# PAND2X1_69/m4_208_n4#
+ PAND2X1_69/O PAND2X1_69/a_56_28# PAND2X1_69/CTRL2 PAND2X1_69/CTRL PAND2X1_69/a_76_28#
+ PAND2X1
XPOR2X1_616 VDD GND POR2X1_20/B POR2X1_411/B POR2X1_616/Y POR2X1_616/m4_208_n4# POR2X1_616/O
+ POR2X1_616/CTRL2 POR2X1_616/a_16_28# POR2X1_616/CTRL POR2X1_616/a_76_344# POR2X1_616/a_56_344#
+ POR2X1
XPOR2X1_605 VDD GND POR2X1_605/B POR2X1_605/A POR2X1_718/A POR2X1_605/m4_208_n4# POR2X1_605/O
+ POR2X1_605/CTRL2 POR2X1_605/a_16_28# POR2X1_605/CTRL POR2X1_605/a_76_344# POR2X1_605/a_56_344#
+ POR2X1
XPOR2X1_627 VDD GND POR2X1_7/A POR2X1_39/B POR2X1_627/Y POR2X1_627/m4_208_n4# POR2X1_627/O
+ POR2X1_627/CTRL2 POR2X1_627/a_16_28# POR2X1_627/CTRL POR2X1_627/a_76_344# POR2X1_627/a_56_344#
+ POR2X1
XPOR2X1_638 VDD GND POR2X1_638/B POR2X1_638/A POR2X1_638/Y POR2X1_638/m4_208_n4# POR2X1_638/O
+ POR2X1_638/CTRL2 POR2X1_638/a_16_28# POR2X1_638/CTRL POR2X1_638/a_76_344# POR2X1_638/a_56_344#
+ POR2X1
XPOR2X1_649 VDD GND POR2X1_649/B POR2X1_643/Y POR2X1_655/A POR2X1_649/m4_208_n4# POR2X1_649/O
+ POR2X1_649/CTRL2 POR2X1_649/a_16_28# POR2X1_649/CTRL POR2X1_649/a_76_344# POR2X1_649/a_56_344#
+ POR2X1
XPOR2X1_413 VDD GND D_INPUT_0 POR2X1_413/A POR2X1_413/Y POR2X1_413/m4_208_n4# POR2X1_413/O
+ POR2X1_413/CTRL2 POR2X1_413/a_16_28# POR2X1_413/CTRL POR2X1_413/a_76_344# POR2X1_413/a_56_344#
+ POR2X1
XPOR2X1_402 VDD GND POR2X1_402/B POR2X1_402/A POR2X1_404/B POR2X1_402/m4_208_n4# POR2X1_402/O
+ POR2X1_402/CTRL2 POR2X1_402/a_16_28# POR2X1_402/CTRL POR2X1_402/a_76_344# POR2X1_402/a_56_344#
+ POR2X1
XPOR2X1_424 VDD GND POR2X1_57/A POR2X1_77/Y POR2X1_424/Y POR2X1_424/m4_208_n4# POR2X1_424/O
+ POR2X1_424/CTRL2 POR2X1_424/a_16_28# POR2X1_424/CTRL POR2X1_424/a_76_344# POR2X1_424/a_56_344#
+ POR2X1
XPOR2X1_435 VDD GND POR2X1_435/B POR2X1_832/A POR2X1_435/Y POR2X1_722/m4_208_n4# POR2X1_435/O
+ POR2X1_435/CTRL2 POR2X1_435/a_16_28# POR2X1_435/CTRL POR2X1_435/a_76_344# POR2X1_435/a_56_344#
+ POR2X1
XPOR2X1_446 VDD GND POR2X1_446/B POR2X1_446/A POR2X1_454/B POR2X1_446/m4_208_n4# POR2X1_446/O
+ POR2X1_446/CTRL2 POR2X1_446/a_16_28# POR2X1_446/CTRL POR2X1_446/a_76_344# POR2X1_446/a_56_344#
+ POR2X1
XPOR2X1_457 VDD GND POR2X1_457/B POR2X1_370/Y POR2X1_457/Y POR2X1_457/m4_208_n4# POR2X1_457/O
+ POR2X1_457/CTRL2 POR2X1_457/a_16_28# POR2X1_457/CTRL POR2X1_457/a_76_344# POR2X1_457/a_56_344#
+ POR2X1
XPOR2X1_468 VDD GND POR2X1_468/B POR2X1_440/Y POR2X1_468/Y POR2X1_468/m4_208_n4# POR2X1_468/O
+ POR2X1_468/CTRL2 POR2X1_468/a_16_28# POR2X1_468/CTRL POR2X1_468/a_76_344# POR2X1_468/a_56_344#
+ POR2X1
XPOR2X1_479 VDD GND POR2X1_479/B POR2X1_476/Y POR2X1_480/A POR2X1_479/m4_208_n4# POR2X1_479/O
+ POR2X1_479/CTRL2 POR2X1_479/a_16_28# POR2X1_479/CTRL POR2X1_479/a_76_344# POR2X1_479/a_56_344#
+ POR2X1
XPAND2X1_409 VDD GND PAND2X1_408/Y POR2X1_407/Y POR2X1_460/A PAND2X1_409/a_16_344#
+ PAND2X1_409/m4_208_n4# PAND2X1_409/O PAND2X1_409/a_56_28# PAND2X1_409/CTRL2 PAND2X1_409/CTRL
+ PAND2X1_409/a_76_28# PAND2X1
XPOR2X1_210 VDD GND POR2X1_210/B POR2X1_210/A POR2X1_210/Y POR2X1_210/m4_208_n4# POR2X1_210/O
+ POR2X1_210/CTRL2 POR2X1_210/a_16_28# POR2X1_210/CTRL POR2X1_210/a_76_344# POR2X1_210/a_56_344#
+ POR2X1
XPOR2X1_221 VDD GND POR2X1_192/Y POR2X1_220/Y POR2X1_221/Y POR2X1_294/m4_208_n4# POR2X1_221/O
+ POR2X1_221/CTRL2 POR2X1_221/a_16_28# POR2X1_221/CTRL POR2X1_221/a_76_344# POR2X1_221/a_56_344#
+ POR2X1
XPOR2X1_232 VDD GND POR2X1_16/A POR2X1_416/B POR2X1_232/Y POR2X1_232/m4_208_n4# POR2X1_232/O
+ POR2X1_232/CTRL2 POR2X1_232/a_16_28# POR2X1_232/CTRL POR2X1_232/a_76_344# POR2X1_232/a_56_344#
+ POR2X1
XPOR2X1_243 VDD GND POR2X1_243/B POR2X1_243/A POR2X1_243/Y POR2X1_243/m4_208_n4# POR2X1_243/O
+ POR2X1_243/CTRL2 POR2X1_243/a_16_28# POR2X1_243/CTRL POR2X1_243/a_76_344# POR2X1_243/a_56_344#
+ POR2X1
XPOR2X1_265 VDD GND POR2X1_40/Y POR2X1_667/A POR2X1_265/Y POR2X1_265/m4_208_n4# POR2X1_265/O
+ POR2X1_265/CTRL2 POR2X1_265/a_16_28# POR2X1_265/CTRL POR2X1_265/a_76_344# POR2X1_265/a_56_344#
+ POR2X1
XPOR2X1_254 VDD GND POR2X1_483/B POR2X1_254/A POR2X1_254/Y POR2X1_254/m4_208_n4# POR2X1_254/O
+ POR2X1_254/CTRL2 POR2X1_254/a_16_28# POR2X1_254/CTRL POR2X1_254/a_76_344# POR2X1_254/a_56_344#
+ POR2X1
XPOR2X1_276 VDD GND POR2X1_276/B POR2X1_276/A POR2X1_276/Y POR2X1_366/m4_208_n4# POR2X1_276/O
+ POR2X1_276/CTRL2 POR2X1_276/a_16_28# POR2X1_276/CTRL POR2X1_276/a_76_344# POR2X1_276/a_56_344#
+ POR2X1
XPOR2X1_298 VDD GND POR2X1_32/A POR2X1_55/Y POR2X1_298/Y POR2X1_298/m4_208_n4# POR2X1_298/O
+ POR2X1_298/CTRL2 POR2X1_298/a_16_28# POR2X1_298/CTRL POR2X1_298/a_76_344# POR2X1_298/a_56_344#
+ POR2X1
XPOR2X1_287 VDD GND POR2X1_287/B POR2X1_287/A POR2X1_288/A POR2X1_287/m4_208_n4# POR2X1_287/O
+ POR2X1_287/CTRL2 POR2X1_287/a_16_28# POR2X1_287/CTRL POR2X1_287/a_76_344# POR2X1_287/a_56_344#
+ POR2X1
XPAND2X1_206 VDD GND PAND2X1_206/B PAND2X1_206/A PAND2X1_215/B PAND2X1_206/a_16_344#
+ PAND2X1_206/m4_208_n4# PAND2X1_206/O PAND2X1_206/a_56_28# PAND2X1_206/CTRL2 PAND2X1_206/CTRL
+ PAND2X1_206/a_76_28# PAND2X1
XPAND2X1_228 VDD GND POR2X1_52/Y POR2X1_7/Y PAND2X1_341/A PAND2X1_228/a_16_344# PAND2X1_228/m4_208_n4#
+ PAND2X1_228/O PAND2X1_228/a_56_28# PAND2X1_228/CTRL2 PAND2X1_228/CTRL PAND2X1_228/a_76_28#
+ PAND2X1
XPAND2X1_217 VDD GND PAND2X1_217/B PAND2X1_124/Y PAND2X1_218/B PAND2X1_217/a_16_344#
+ PAND2X1_217/m4_208_n4# PAND2X1_217/O PAND2X1_217/a_56_28# PAND2X1_217/CTRL2 PAND2X1_217/CTRL
+ PAND2X1_217/a_76_28# PAND2X1
XPAND2X1_239 VDD GND POR2X1_590/A PAND2X1_52/B POR2X1_506/B PAND2X1_239/a_16_344#
+ PAND2X1_239/m4_208_n4# PAND2X1_239/O PAND2X1_239/a_56_28# PAND2X1_239/CTRL2 PAND2X1_239/CTRL
+ PAND2X1_239/a_76_28# PAND2X1
XPAND2X1_740 VDD GND PAND2X1_739/Y PAND2X1_738/Y PAND2X1_740/Y PAND2X1_740/a_16_344#
+ PAND2X1_740/m4_208_n4# PAND2X1_740/O PAND2X1_740/a_56_28# PAND2X1_740/CTRL2 PAND2X1_740/CTRL
+ PAND2X1_740/a_76_28# PAND2X1
XPAND2X1_751 VDD GND POR2X1_750/Y POR2X1_66/B POR2X1_789/A PAND2X1_751/a_16_344# PAND2X1_751/m4_208_n4#
+ PAND2X1_751/O PAND2X1_751/a_56_28# PAND2X1_751/CTRL2 PAND2X1_751/CTRL PAND2X1_751/a_76_28#
+ PAND2X1
XPAND2X1_773 VDD GND PAND2X1_773/B POR2X1_767/Y PAND2X1_773/Y PAND2X1_773/a_16_344#
+ PAND2X1_773/m4_208_n4# PAND2X1_773/O PAND2X1_773/a_56_28# PAND2X1_773/CTRL2 PAND2X1_773/CTRL
+ PAND2X1_773/a_76_28# PAND2X1
XPAND2X1_762 VDD GND PAND2X1_11/Y INPUT_6 PAND2X1_762/Y PAND2X1_762/a_16_344# PAND2X1_762/m4_208_n4#
+ PAND2X1_762/O PAND2X1_762/a_56_28# PAND2X1_762/CTRL2 PAND2X1_762/CTRL PAND2X1_762/a_76_28#
+ PAND2X1
XPAND2X1_795 VDD GND PAND2X1_795/B PAND2X1_785/Y PAND2X1_804/B PAND2X1_795/a_16_344#
+ PAND2X1_795/m4_208_n4# PAND2X1_795/O PAND2X1_795/a_56_28# PAND2X1_795/CTRL2 PAND2X1_795/CTRL
+ PAND2X1_795/a_76_28# PAND2X1
XPAND2X1_784 VDD GND PAND2X1_778/Y PAND2X1_784/A PAND2X1_796/B PAND2X1_784/a_16_344#
+ PAND2X1_784/m4_208_n4# PAND2X1_784/O PAND2X1_784/a_56_28# PAND2X1_784/CTRL2 PAND2X1_784/CTRL
+ PAND2X1_784/a_76_28# PAND2X1
XPAND2X1_592 VDD GND POR2X1_589/Y POR2X1_423/Y PAND2X1_592/Y PAND2X1_592/a_16_344#
+ PAND2X1_592/m4_208_n4# PAND2X1_592/O PAND2X1_592/a_56_28# PAND2X1_592/CTRL2 PAND2X1_592/CTRL
+ PAND2X1_592/a_76_28# PAND2X1
XPAND2X1_570 VDD GND PAND2X1_570/B PAND2X1_562/Y PAND2X1_577/B PAND2X1_570/a_16_344#
+ PAND2X1_570/m4_208_n4# PAND2X1_570/O PAND2X1_570/a_56_28# PAND2X1_570/CTRL2 PAND2X1_570/CTRL
+ PAND2X1_570/a_76_28# PAND2X1
XPAND2X1_581 VDD GND PAND2X1_3/B INPUT_6 PAND2X1_581/Y PAND2X1_581/a_16_344# PAND2X1_581/m4_208_n4#
+ PAND2X1_581/O PAND2X1_581/a_56_28# PAND2X1_581/CTRL2 PAND2X1_581/CTRL PAND2X1_581/a_76_28#
+ PAND2X1
XPOR2X1_809 VDD GND POR2X1_809/B POR2X1_809/A POR2X1_809/Y POR2X1_809/m4_208_n4# POR2X1_809/O
+ POR2X1_809/CTRL2 POR2X1_809/a_16_28# POR2X1_809/CTRL POR2X1_809/a_76_344# POR2X1_809/a_56_344#
+ POR2X1
XPAND2X1_26 VDD GND PAND2X1_59/B PAND2X1_26/A POR2X1_66/A PAND2X1_26/a_16_344# PAND2X1_26/m4_208_n4#
+ PAND2X1_26/O PAND2X1_26/a_56_28# PAND2X1_26/CTRL2 PAND2X1_26/CTRL PAND2X1_26/a_76_28#
+ PAND2X1
XPAND2X1_15 VDD GND PAND2X1_94/A PAND2X1_9/Y POR2X1_78/B PAND2X1_15/a_16_344# PAND2X1_15/m4_208_n4#
+ PAND2X1_15/O PAND2X1_15/a_56_28# PAND2X1_15/CTRL2 PAND2X1_15/CTRL PAND2X1_15/a_76_28#
+ PAND2X1
XPAND2X1_48 VDD GND PAND2X1_48/B PAND2X1_48/A PAND2X1_48/Y PAND2X1_48/a_16_344# PAND2X1_48/m4_208_n4#
+ PAND2X1_48/O PAND2X1_48/a_56_28# PAND2X1_48/CTRL2 PAND2X1_48/CTRL PAND2X1_48/a_76_28#
+ PAND2X1
XPAND2X1_59 VDD GND PAND2X1_59/B PAND2X1_11/Y PAND2X1_60/B PAND2X1_59/a_16_344# PAND2X1_59/m4_208_n4#
+ PAND2X1_59/O PAND2X1_59/a_56_28# PAND2X1_59/CTRL2 PAND2X1_59/CTRL PAND2X1_59/a_76_28#
+ PAND2X1
XPAND2X1_37 VDD GND INPUT_3 INPUT_2 PAND2X1_90/A PAND2X1_37/a_16_344# PAND2X1_37/m4_208_n4#
+ PAND2X1_37/O PAND2X1_37/a_56_28# PAND2X1_37/CTRL2 PAND2X1_37/CTRL PAND2X1_37/a_76_28#
+ PAND2X1
XPOR2X1_617 VDD GND POR2X1_38/Y POR2X1_52/A POR2X1_617/Y POR2X1_617/m4_208_n4# POR2X1_617/O
+ POR2X1_617/CTRL2 POR2X1_617/a_16_28# POR2X1_617/CTRL POR2X1_617/a_76_344# POR2X1_617/a_56_344#
+ POR2X1
XPOR2X1_606 VDD GND POR2X1_590/A POR2X1_121/B POR2X1_606/Y POR2X1_606/m4_208_n4# POR2X1_606/O
+ POR2X1_606/CTRL2 POR2X1_606/a_16_28# POR2X1_606/CTRL POR2X1_606/a_76_344# POR2X1_606/a_56_344#
+ POR2X1
XPOR2X1_639 VDD GND POR2X1_635/Y POR2X1_639/A POR2X1_639/Y POR2X1_639/m4_208_n4# POR2X1_639/O
+ POR2X1_639/CTRL2 POR2X1_639/a_16_28# POR2X1_639/CTRL POR2X1_639/a_76_344# POR2X1_639/a_56_344#
+ POR2X1
XPOR2X1_628 VDD GND POR2X1_48/A POR2X1_93/A POR2X1_628/Y POR2X1_628/m4_208_n4# POR2X1_628/O
+ POR2X1_628/CTRL2 POR2X1_628/a_16_28# POR2X1_628/CTRL POR2X1_628/a_76_344# POR2X1_628/a_56_344#
+ POR2X1
XPOR2X1_414 VDD GND D_INPUT_3 POR2X1_4/Y POR2X1_414/Y POR2X1_414/m4_208_n4# POR2X1_414/O
+ POR2X1_414/CTRL2 POR2X1_414/a_16_28# POR2X1_414/CTRL POR2X1_414/a_76_344# POR2X1_414/a_56_344#
+ POR2X1
XPOR2X1_403 VDD GND POR2X1_403/B POR2X1_403/A POR2X1_403/Y POR2X1_403/m4_208_n4# POR2X1_403/O
+ POR2X1_403/CTRL2 POR2X1_403/a_16_28# POR2X1_403/CTRL POR2X1_403/a_76_344# POR2X1_403/a_56_344#
+ POR2X1
XPOR2X1_425 VDD GND INPUT_5 POR2X1_36/B POR2X1_425/Y POR2X1_425/m4_208_n4# POR2X1_425/O
+ POR2X1_425/CTRL2 POR2X1_425/a_16_28# POR2X1_425/CTRL POR2X1_425/a_76_344# POR2X1_425/a_56_344#
+ POR2X1
XPOR2X1_447 VDD GND POR2X1_447/B POR2X1_447/A POR2X1_454/A POR2X1_447/m4_208_n4# POR2X1_447/O
+ POR2X1_447/CTRL2 POR2X1_447/a_16_28# POR2X1_447/CTRL POR2X1_447/a_76_344# POR2X1_447/a_56_344#
+ POR2X1
XPOR2X1_458 VDD GND POR2X1_458/B POR2X1_717/B POR2X1_458/Y POR2X1_458/m4_208_n4# POR2X1_458/O
+ POR2X1_458/CTRL2 POR2X1_458/a_16_28# POR2X1_458/CTRL POR2X1_458/a_76_344# POR2X1_458/a_56_344#
+ POR2X1
XPOR2X1_436 VDD GND POR2X1_436/B POR2X1_435/Y POR2X1_468/B POR2X1_436/m4_208_n4# POR2X1_436/O
+ POR2X1_436/CTRL2 POR2X1_436/a_16_28# POR2X1_436/CTRL POR2X1_436/a_76_344# POR2X1_436/a_56_344#
+ POR2X1
XPOR2X1_469 VDD GND POR2X1_444/Y POR2X1_468/Y POR2X1_478/B POR2X1_469/m4_208_n4# POR2X1_469/O
+ POR2X1_469/CTRL2 POR2X1_469/a_16_28# POR2X1_469/CTRL POR2X1_469/a_76_344# POR2X1_469/a_56_344#
+ POR2X1
XPOR2X1_200 VDD GND POR2X1_193/Y POR2X1_200/A POR2X1_207/A POR2X1_200/m4_208_n4# POR2X1_200/O
+ POR2X1_200/CTRL2 POR2X1_200/a_16_28# POR2X1_200/CTRL POR2X1_200/a_76_344# POR2X1_200/a_56_344#
+ POR2X1
XPOR2X1_233 VDD GND D_INPUT_0 POR2X1_14/Y POR2X1_234/A POR2X1_233/m4_208_n4# POR2X1_233/O
+ POR2X1_233/CTRL2 POR2X1_233/a_16_28# POR2X1_233/CTRL POR2X1_233/a_76_344# POR2X1_233/a_56_344#
+ POR2X1
XPOR2X1_211 VDD GND POR2X1_566/B POR2X1_853/A POR2X1_212/A POR2X1_211/m4_208_n4# POR2X1_211/O
+ POR2X1_211/CTRL2 POR2X1_211/a_16_28# POR2X1_211/CTRL POR2X1_211/a_76_344# POR2X1_211/a_56_344#
+ POR2X1
XPOR2X1_222 VDD GND POR2X1_218/Y POR2X1_222/A POR2X1_222/Y POR2X1_222/m4_208_n4# POR2X1_222/O
+ POR2X1_222/CTRL2 POR2X1_222/a_16_28# POR2X1_222/CTRL POR2X1_222/a_76_344# POR2X1_222/a_56_344#
+ POR2X1
XPOR2X1_244 VDD GND POR2X1_244/B POR2X1_243/Y POR2X1_244/Y POR2X1_244/m4_208_n4# POR2X1_244/O
+ POR2X1_244/CTRL2 POR2X1_244/a_16_28# POR2X1_244/CTRL POR2X1_244/a_76_344# POR2X1_244/a_56_344#
+ POR2X1
XPOR2X1_277 VDD GND POR2X1_37/Y POR2X1_48/A POR2X1_278/A POR2X1_277/m4_208_n4# POR2X1_277/O
+ POR2X1_277/CTRL2 POR2X1_277/a_16_28# POR2X1_277/CTRL POR2X1_277/a_76_344# POR2X1_277/a_56_344#
+ POR2X1
XPOR2X1_266 VDD GND POR2X1_786/A POR2X1_266/A POR2X1_267/A POR2X1_266/m4_208_n4# POR2X1_266/O
+ POR2X1_266/CTRL2 POR2X1_266/a_16_28# POR2X1_266/CTRL POR2X1_266/a_76_344# POR2X1_266/a_56_344#
+ POR2X1
XPOR2X1_255 VDD GND POR2X1_37/Y POR2X1_416/B POR2X1_255/Y POR2X1_255/m4_208_n4# POR2X1_255/O
+ POR2X1_255/CTRL2 POR2X1_255/a_16_28# POR2X1_255/CTRL POR2X1_255/a_76_344# POR2X1_255/a_56_344#
+ POR2X1
XPOR2X1_299 VDD GND POR2X1_13/A POR2X1_119/Y POR2X1_299/Y POR2X1_299/m4_208_n4# POR2X1_299/O
+ POR2X1_299/CTRL2 POR2X1_299/a_16_28# POR2X1_299/CTRL POR2X1_299/a_76_344# POR2X1_299/a_56_344#
+ POR2X1
XPOR2X1_288 VDD GND POR2X1_286/Y POR2X1_288/A POR2X1_362/B POR2X1_288/m4_208_n4# POR2X1_288/O
+ POR2X1_288/CTRL2 POR2X1_288/a_16_28# POR2X1_288/CTRL POR2X1_288/a_76_344# POR2X1_288/a_56_344#
+ POR2X1
XPAND2X1_218 VDD GND PAND2X1_218/B PAND2X1_218/A PAND2X1_222/A PAND2X1_218/a_16_344#
+ POR2X1_7/m4_208_n4# PAND2X1_218/O PAND2X1_218/a_56_28# PAND2X1_218/CTRL2 PAND2X1_218/CTRL
+ PAND2X1_218/a_76_28# PAND2X1
XPAND2X1_207 VDD GND PAND2X1_200/Y PAND2X1_207/A PAND2X1_214/A PAND2X1_207/a_16_344#
+ PAND2X1_207/m4_208_n4# PAND2X1_207/O PAND2X1_207/a_56_28# PAND2X1_207/CTRL2 PAND2X1_207/CTRL
+ PAND2X1_207/a_76_28# PAND2X1
XPAND2X1_229 VDD GND PAND2X1_23/Y POR2X1_260/B POR2X1_231/B PAND2X1_229/a_16_344#
+ PAND2X1_229/m4_208_n4# PAND2X1_229/O PAND2X1_229/a_56_28# PAND2X1_229/CTRL2 PAND2X1_229/CTRL
+ PAND2X1_229/a_76_28# PAND2X1
XPAND2X1_741 VDD GND PAND2X1_741/B PAND2X1_736/Y PAND2X1_742/B PAND2X1_741/a_16_344#
+ PAND2X1_741/m4_208_n4# PAND2X1_741/O PAND2X1_741/a_56_28# PAND2X1_741/CTRL2 PAND2X1_741/CTRL
+ PAND2X1_741/a_76_28# PAND2X1
XPAND2X1_730 VDD GND PAND2X1_730/B PAND2X1_730/A PAND2X1_739/B PAND2X1_730/a_16_344#
+ PAND2X1_730/m4_208_n4# PAND2X1_730/O PAND2X1_730/a_56_28# PAND2X1_730/CTRL2 PAND2X1_730/CTRL
+ PAND2X1_730/a_76_28# PAND2X1
XPAND2X1_774 VDD GND PAND2X1_773/Y PAND2X1_771/Y PAND2X1_810/A PAND2X1_774/a_16_344#
+ PAND2X1_580/m4_208_n4# PAND2X1_774/O PAND2X1_774/a_56_28# PAND2X1_774/CTRL2 PAND2X1_774/CTRL
+ PAND2X1_774/a_76_28# PAND2X1
XPAND2X1_752 VDD GND PAND2X1_95/B INPUT_5 PAND2X1_752/Y PAND2X1_752/a_16_344# PAND2X1_752/m4_208_n4#
+ PAND2X1_752/O PAND2X1_752/a_56_28# PAND2X1_752/CTRL2 PAND2X1_752/CTRL PAND2X1_752/a_76_28#
+ PAND2X1
XPAND2X1_763 VDD GND PAND2X1_762/Y PAND2X1_48/A POR2X1_769/B PAND2X1_763/a_16_344#
+ PAND2X1_763/m4_208_n4# PAND2X1_763/O PAND2X1_763/a_56_28# PAND2X1_763/CTRL2 PAND2X1_763/CTRL
+ PAND2X1_763/a_76_28# PAND2X1
XPAND2X1_785 VDD GND PAND2X1_776/Y PAND2X1_785/A PAND2X1_785/Y PAND2X1_785/a_16_344#
+ PAND2X1_785/m4_208_n4# PAND2X1_785/O PAND2X1_785/a_56_28# PAND2X1_785/CTRL2 PAND2X1_785/CTRL
+ PAND2X1_785/a_76_28# PAND2X1
XPAND2X1_796 VDD GND PAND2X1_796/B PAND2X1_783/Y PAND2X1_803/A PAND2X1_796/a_16_344#
+ PAND2X1_796/m4_208_n4# PAND2X1_796/O PAND2X1_796/a_56_28# PAND2X1_796/CTRL2 PAND2X1_796/CTRL
+ PAND2X1_796/a_76_28# PAND2X1
XPAND2X1_560 VDD GND PAND2X1_560/B PAND2X1_844/B PAND2X1_571/A PAND2X1_560/a_16_344#
+ PAND2X1_560/m4_208_n4# PAND2X1_560/O PAND2X1_560/a_56_28# PAND2X1_560/CTRL2 PAND2X1_560/CTRL
+ PAND2X1_560/a_76_28# PAND2X1
XPAND2X1_571 VDD GND PAND2X1_561/Y PAND2X1_571/A PAND2X1_571/Y PAND2X1_571/a_16_344#
+ PAND2X1_571/m4_208_n4# PAND2X1_571/O PAND2X1_571/a_56_28# PAND2X1_571/CTRL2 PAND2X1_571/CTRL
+ PAND2X1_571/a_76_28# PAND2X1
XPAND2X1_582 VDD GND PAND2X1_581/Y POR2X1_614/A POR2X1_635/A PAND2X1_582/a_16_344#
+ PAND2X1_582/m4_208_n4# PAND2X1_582/O PAND2X1_582/a_56_28# PAND2X1_582/CTRL2 PAND2X1_582/CTRL
+ PAND2X1_582/a_76_28# PAND2X1
XPAND2X1_593 VDD GND PAND2X1_592/Y POR2X1_591/Y PAND2X1_593/Y PAND2X1_593/a_16_344#
+ PAND2X1_593/m4_208_n4# PAND2X1_593/O PAND2X1_593/a_56_28# PAND2X1_593/CTRL2 PAND2X1_593/CTRL
+ PAND2X1_593/a_76_28# PAND2X1
XPAND2X1_390 VDD GND PAND2X1_389/Y PAND2X1_388/Y PAND2X1_390/Y PAND2X1_390/a_16_344#
+ PAND2X1_390/m4_208_n4# PAND2X1_390/O PAND2X1_390/a_56_28# PAND2X1_390/CTRL2 PAND2X1_390/CTRL
+ PAND2X1_390/a_76_28# PAND2X1
XPAND2X1_16 VDD GND POR2X1_78/B POR2X1_66/B POR2X1_194/B PAND2X1_16/a_16_344# PAND2X1_16/m4_208_n4#
+ PAND2X1_16/O PAND2X1_16/a_56_28# PAND2X1_16/CTRL2 PAND2X1_16/CTRL PAND2X1_16/a_76_28#
+ PAND2X1
XPAND2X1_38 VDD GND PAND2X1_90/A POR2X1_29/A PAND2X1_39/B PAND2X1_38/a_16_344# PAND2X1_38/m4_208_n4#
+ PAND2X1_38/O PAND2X1_38/a_56_28# PAND2X1_38/CTRL2 PAND2X1_38/CTRL PAND2X1_38/a_76_28#
+ PAND2X1
XPAND2X1_49 VDD GND POR2X1_29/A PAND2X1_94/A POR2X1_68/A PAND2X1_49/a_16_344# PAND2X1_49/m4_208_n4#
+ PAND2X1_49/O PAND2X1_49/a_56_28# PAND2X1_49/CTRL2 PAND2X1_49/CTRL PAND2X1_49/a_76_28#
+ PAND2X1
XPAND2X1_27 VDD GND POR2X1_66/A PAND2X1_6/Y POR2X1_34/B PAND2X1_27/a_16_344# PAND2X1_27/m4_208_n4#
+ PAND2X1_27/O PAND2X1_27/a_56_28# PAND2X1_27/CTRL2 PAND2X1_27/CTRL PAND2X1_27/a_76_28#
+ PAND2X1
XPOR2X1_607 VDD GND POR2X1_20/B POR2X1_607/A POR2X1_607/Y POR2X1_607/m4_208_n4# POR2X1_607/O
+ POR2X1_607/CTRL2 POR2X1_607/a_16_28# POR2X1_607/CTRL POR2X1_607/a_76_344# POR2X1_607/a_56_344#
+ POR2X1
XPOR2X1_618 VDD GND INPUT_3 POR2X1_38/B POR2X1_619/A POR2X1_618/m4_208_n4# POR2X1_618/O
+ POR2X1_618/CTRL2 POR2X1_618/a_16_28# POR2X1_618/CTRL POR2X1_618/a_76_344# POR2X1_618/a_56_344#
+ POR2X1
XPOR2X1_629 VDD GND POR2X1_629/B POR2X1_629/A POR2X1_630/A POR2X1_629/m4_208_n4# POR2X1_629/O
+ POR2X1_629/CTRL2 POR2X1_629/a_16_28# POR2X1_629/CTRL POR2X1_629/a_76_344# POR2X1_629/a_56_344#
+ POR2X1
XPOR2X1_404 VDD GND POR2X1_404/B POR2X1_403/Y POR2X1_404/Y POR2X1_404/m4_208_n4# POR2X1_404/O
+ POR2X1_404/CTRL2 POR2X1_404/a_16_28# POR2X1_404/CTRL POR2X1_404/a_76_344# POR2X1_404/a_56_344#
+ POR2X1
XPOR2X1_415 VDD GND POR2X1_294/A POR2X1_415/A POR2X1_415/Y POR2X1_415/m4_208_n4# POR2X1_415/O
+ POR2X1_415/CTRL2 POR2X1_415/a_16_28# POR2X1_415/CTRL POR2X1_415/a_76_344# POR2X1_415/a_56_344#
+ POR2X1
XPOR2X1_426 VDD GND POR2X1_119/Y POR2X1_425/Y POR2X1_426/Y POR2X1_426/m4_208_n4# POR2X1_426/O
+ POR2X1_426/CTRL2 POR2X1_426/a_16_28# POR2X1_426/CTRL POR2X1_426/a_76_344# POR2X1_426/a_56_344#
+ POR2X1
XPOR2X1_437 VDD GND POR2X1_60/A POR2X1_150/Y POR2X1_437/Y POR2X1_437/m4_208_n4# POR2X1_437/O
+ POR2X1_437/CTRL2 POR2X1_437/a_16_28# POR2X1_437/CTRL POR2X1_437/a_76_344# POR2X1_437/a_56_344#
+ POR2X1
XPOR2X1_448 VDD GND POR2X1_448/B POR2X1_448/A POR2X1_448/Y POR2X1_448/m4_208_n4# POR2X1_448/O
+ POR2X1_448/CTRL2 POR2X1_448/a_16_28# POR2X1_448/CTRL POR2X1_448/a_76_344# POR2X1_448/a_56_344#
+ POR2X1
XPOR2X1_459 VDD GND POR2X1_459/B POR2X1_459/A POR2X1_459/Y POR2X1_459/m4_208_n4# POR2X1_459/O
+ POR2X1_459/CTRL2 POR2X1_459/a_16_28# POR2X1_459/CTRL POR2X1_459/a_76_344# POR2X1_459/a_56_344#
+ POR2X1
XPOR2X1_201 VDD GND POR2X1_61/Y PAND2X1_65/Y POR2X1_201/Y POR2X1_201/m4_208_n4# POR2X1_201/O
+ POR2X1_201/CTRL2 POR2X1_201/a_16_28# POR2X1_201/CTRL POR2X1_201/a_76_344# POR2X1_201/a_56_344#
+ POR2X1
XPOR2X1_223 VDD GND POR2X1_221/Y POR2X1_222/Y D_GATE_222 POR2X1_223/m4_208_n4# POR2X1_223/O
+ POR2X1_223/CTRL2 POR2X1_223/a_16_28# POR2X1_223/CTRL POR2X1_223/a_76_344# POR2X1_223/a_56_344#
+ POR2X1
XPOR2X1_234 VDD GND POR2X1_48/A POR2X1_234/A POR2X1_234/Y POR2X1_234/m4_208_n4# POR2X1_234/O
+ POR2X1_234/CTRL2 POR2X1_234/a_16_28# POR2X1_234/CTRL POR2X1_234/a_76_344# POR2X1_234/a_56_344#
+ POR2X1
XPOR2X1_212 VDD GND POR2X1_212/B POR2X1_212/A POR2X1_220/B POR2X1_212/m4_208_n4# POR2X1_212/O
+ POR2X1_212/CTRL2 POR2X1_212/a_16_28# POR2X1_212/CTRL POR2X1_212/a_76_344# POR2X1_212/a_56_344#
+ POR2X1
XPOR2X1_267 VDD GND POR2X1_267/B POR2X1_267/A POR2X1_267/Y POR2X1_267/m4_208_n4# POR2X1_267/O
+ POR2X1_267/CTRL2 POR2X1_267/a_16_28# POR2X1_267/CTRL POR2X1_267/a_76_344# POR2X1_267/a_56_344#
+ POR2X1
XPOR2X1_256 VDD GND PAND2X1_6/A POR2X1_255/Y POR2X1_256/Y POR2X1_256/m4_208_n4# POR2X1_256/O
+ POR2X1_256/CTRL2 POR2X1_256/a_16_28# POR2X1_256/CTRL POR2X1_256/a_76_344# POR2X1_256/a_56_344#
+ POR2X1
XPOR2X1_245 VDD GND POR2X1_83/B POR2X1_37/Y POR2X1_245/Y POR2X1_245/m4_208_n4# POR2X1_245/O
+ POR2X1_245/CTRL2 POR2X1_245/a_16_28# POR2X1_245/CTRL POR2X1_245/a_76_344# POR2X1_245/a_56_344#
+ POR2X1
XPOR2X1_278 VDD GND PAND2X1_9/Y POR2X1_278/A POR2X1_278/Y POR2X1_278/m4_208_n4# POR2X1_278/O
+ POR2X1_278/CTRL2 POR2X1_278/a_16_28# POR2X1_278/CTRL POR2X1_278/a_76_344# POR2X1_278/a_56_344#
+ POR2X1
XPOR2X1_289 VDD GND POR2X1_52/A POR2X1_283/A POR2X1_289/Y POR2X1_289/m4_208_n4# POR2X1_289/O
+ POR2X1_289/CTRL2 POR2X1_289/a_16_28# POR2X1_289/CTRL POR2X1_289/a_76_344# POR2X1_289/a_56_344#
+ POR2X1
XPAND2X1_208 VDD GND PAND2X1_198/Y PAND2X1_35/Y PAND2X1_214/B PAND2X1_208/a_16_344#
+ PAND2X1_208/m4_208_n4# PAND2X1_208/O PAND2X1_208/a_56_28# PAND2X1_208/CTRL2 PAND2X1_208/CTRL
+ PAND2X1_208/a_76_28# PAND2X1
XPAND2X1_219 VDD GND PAND2X1_219/B PAND2X1_219/A PAND2X1_222/B PAND2X1_219/a_16_344#
+ PAND2X1_219/m4_208_n4# PAND2X1_219/O PAND2X1_219/a_56_28# PAND2X1_219/CTRL2 PAND2X1_219/CTRL
+ PAND2X1_219/a_76_28# PAND2X1
XPOR2X1_790 VDD GND POR2X1_790/B POR2X1_790/A POR2X1_793/A POR2X1_790/m4_208_n4# POR2X1_790/O
+ POR2X1_790/CTRL2 POR2X1_790/a_16_28# POR2X1_790/CTRL POR2X1_790/a_76_344# POR2X1_790/a_56_344#
+ POR2X1
XPAND2X1_731 VDD GND PAND2X1_731/B PAND2X1_731/A PAND2X1_738/A PAND2X1_731/a_16_344#
+ PAND2X1_731/m4_208_n4# PAND2X1_731/O PAND2X1_731/a_56_28# PAND2X1_731/CTRL2 PAND2X1_731/CTRL
+ PAND2X1_731/a_76_28# PAND2X1
XPAND2X1_720 VDD GND POR2X1_669/Y POR2X1_667/Y PAND2X1_721/B PAND2X1_720/a_16_344#
+ PAND2X1_720/m4_208_n4# PAND2X1_720/O PAND2X1_720/a_56_28# PAND2X1_720/CTRL2 PAND2X1_720/CTRL
+ PAND2X1_720/a_76_28# PAND2X1
XPAND2X1_742 VDD GND PAND2X1_742/B PAND2X1_740/Y GATE_741 PAND2X1_742/a_16_344# PAND2X1_675/m4_208_n4#
+ PAND2X1_742/O PAND2X1_742/a_56_28# PAND2X1_742/CTRL2 PAND2X1_742/CTRL PAND2X1_742/a_76_28#
+ PAND2X1
XPAND2X1_753 VDD GND PAND2X1_752/Y POR2X1_188/A POR2X1_790/B PAND2X1_753/a_16_344#
+ PAND2X1_753/m4_208_n4# PAND2X1_753/O PAND2X1_753/a_56_28# PAND2X1_753/CTRL2 PAND2X1_753/CTRL
+ PAND2X1_753/a_76_28# PAND2X1
XPAND2X1_764 VDD GND POR2X1_532/A PAND2X1_41/B POR2X1_769/A PAND2X1_764/a_16_344#
+ PAND2X1_764/m4_208_n4# PAND2X1_764/O PAND2X1_764/a_56_28# PAND2X1_764/CTRL2 PAND2X1_764/CTRL
+ PAND2X1_764/a_76_28# PAND2X1
XPAND2X1_786 VDD GND POR2X1_262/Y PAND2X1_84/Y PAND2X1_795/B PAND2X1_786/a_16_344#
+ PAND2X1_786/m4_208_n4# PAND2X1_786/O PAND2X1_786/a_56_28# PAND2X1_786/CTRL2 PAND2X1_786/CTRL
+ PAND2X1_786/a_76_28# PAND2X1
XPAND2X1_775 VDD GND POR2X1_109/Y POR2X1_91/Y PAND2X1_785/A PAND2X1_775/a_16_344#
+ PAND2X1_775/m4_208_n4# PAND2X1_775/O PAND2X1_775/a_56_28# PAND2X1_775/CTRL2 PAND2X1_775/CTRL
+ PAND2X1_775/a_76_28# PAND2X1
XPAND2X1_797 VDD GND PAND2X1_782/Y PAND2X1_209/A PAND2X1_797/Y PAND2X1_797/a_16_344#
+ PAND2X1_797/m4_208_n4# PAND2X1_797/O PAND2X1_797/a_56_28# PAND2X1_797/CTRL2 PAND2X1_797/CTRL
+ PAND2X1_797/a_76_28# PAND2X1
XPAND2X1_572 VDD GND PAND2X1_267/Y PAND2X1_124/Y PAND2X1_576/B PAND2X1_572/a_16_344#
+ PAND2X1_572/m4_208_n4# PAND2X1_572/O PAND2X1_572/a_56_28# PAND2X1_572/CTRL2 PAND2X1_572/CTRL
+ PAND2X1_572/a_76_28# PAND2X1
XPAND2X1_561 VDD GND PAND2X1_558/Y PAND2X1_561/A PAND2X1_561/Y PAND2X1_561/a_16_344#
+ PAND2X1_561/m4_208_n4# PAND2X1_561/O PAND2X1_561/a_56_28# PAND2X1_561/CTRL2 PAND2X1_561/CTRL
+ PAND2X1_561/a_76_28# PAND2X1
XPAND2X1_550 VDD GND PAND2X1_550/B PAND2X1_546/Y PAND2X1_550/Y PAND2X1_550/a_16_344#
+ PAND2X1_550/m4_208_n4# PAND2X1_550/O PAND2X1_550/a_56_28# PAND2X1_550/CTRL2 PAND2X1_550/CTRL
+ PAND2X1_550/a_76_28# PAND2X1
XPAND2X1_583 VDD GND POR2X1_68/A PAND2X1_32/B POR2X1_636/B PAND2X1_583/a_16_344# PAND2X1_583/m4_208_n4#
+ PAND2X1_583/O PAND2X1_583/a_56_28# PAND2X1_583/CTRL2 PAND2X1_583/CTRL PAND2X1_583/a_76_28#
+ PAND2X1
XPAND2X1_594 VDD GND POR2X1_186/Y PAND2X1_96/B POR2X1_653/B PAND2X1_594/a_16_344#
+ PAND2X1_594/m4_208_n4# PAND2X1_594/O PAND2X1_594/a_56_28# PAND2X1_594/CTRL2 PAND2X1_594/CTRL
+ PAND2X1_594/a_76_28# PAND2X1
XPAND2X1_391 VDD GND POR2X1_384/Y POR2X1_382/Y PAND2X1_392/B PAND2X1_391/a_16_344#
+ PAND2X1_391/m4_208_n4# PAND2X1_391/O PAND2X1_391/a_56_28# PAND2X1_391/CTRL2 PAND2X1_391/CTRL
+ PAND2X1_391/a_76_28# PAND2X1
XPAND2X1_380 VDD GND POR2X1_379/Y POR2X1_532/A POR2X1_460/B PAND2X1_380/a_16_344#
+ PAND2X1_380/m4_208_n4# PAND2X1_380/O PAND2X1_380/a_56_28# PAND2X1_380/CTRL2 PAND2X1_380/CTRL
+ PAND2X1_380/a_76_28# PAND2X1
XPAND2X1_17 VDD GND INPUT_7 INPUT_6 PAND2X1_18/B PAND2X1_17/a_16_344# PAND2X1_17/m4_208_n4#
+ PAND2X1_17/O PAND2X1_17/a_56_28# PAND2X1_17/CTRL2 PAND2X1_17/CTRL PAND2X1_17/a_76_28#
+ PAND2X1
XPAND2X1_28 VDD GND INPUT_1 D_INPUT_0 POR2X1_29/A PAND2X1_28/a_16_344# PAND2X1_28/m4_208_n4#
+ PAND2X1_28/O PAND2X1_28/a_56_28# PAND2X1_28/CTRL2 PAND2X1_28/CTRL PAND2X1_28/a_76_28#
+ PAND2X1
XPAND2X1_39 VDD GND PAND2X1_39/B PAND2X1_69/A POR2X1_194/A PAND2X1_39/a_16_344# PAND2X1_39/m4_208_n4#
+ PAND2X1_39/O PAND2X1_39/a_56_28# PAND2X1_39/CTRL2 PAND2X1_39/CTRL PAND2X1_39/a_76_28#
+ PAND2X1
XPOR2X1_608 VDD GND POR2X1_78/B PAND2X1_73/Y POR2X1_608/Y POR2X1_608/m4_208_n4# POR2X1_608/O
+ POR2X1_608/CTRL2 POR2X1_608/a_16_28# POR2X1_608/CTRL POR2X1_608/a_76_344# POR2X1_608/a_56_344#
+ POR2X1
XPOR2X1_619 VDD GND POR2X1_39/B POR2X1_619/A POR2X1_619/Y POR2X1_619/m4_208_n4# POR2X1_619/O
+ POR2X1_619/CTRL2 POR2X1_619/a_16_28# POR2X1_619/CTRL POR2X1_619/a_76_344# POR2X1_619/a_56_344#
+ POR2X1
XPOR2X1_416 VDD GND POR2X1_416/B POR2X1_416/A POR2X1_416/Y POR2X1_416/m4_208_n4# POR2X1_416/O
+ POR2X1_416/CTRL2 POR2X1_416/a_16_28# POR2X1_416/CTRL POR2X1_416/a_76_344# POR2X1_416/a_56_344#
+ POR2X1
XPOR2X1_405 VDD GND PAND2X1_48/A POR2X1_327/Y POR2X1_405/Y POR2X1_405/m4_208_n4# POR2X1_405/O
+ POR2X1_405/CTRL2 POR2X1_405/a_16_28# POR2X1_405/CTRL POR2X1_405/a_76_344# POR2X1_405/a_56_344#
+ POR2X1
XPOR2X1_438 VDD GND POR2X1_23/Y POR2X1_72/B POR2X1_438/Y POR2X1_438/m4_208_n4# POR2X1_438/O
+ POR2X1_438/CTRL2 POR2X1_438/a_16_28# POR2X1_438/CTRL POR2X1_438/a_76_344# POR2X1_438/a_56_344#
+ POR2X1
XPOR2X1_427 VDD GND POR2X1_72/B POR2X1_257/A POR2X1_427/Y POR2X1_427/m4_208_n4# POR2X1_427/O
+ POR2X1_427/CTRL2 POR2X1_427/a_16_28# POR2X1_427/CTRL POR2X1_427/a_76_344# POR2X1_427/a_56_344#
+ POR2X1
XPOR2X1_449 VDD GND POR2X1_832/B POR2X1_449/A POR2X1_449/Y POR2X1_449/m4_208_n4# POR2X1_449/O
+ POR2X1_449/CTRL2 POR2X1_449/a_16_28# POR2X1_449/CTRL POR2X1_449/a_76_344# POR2X1_449/a_56_344#
+ POR2X1
XPOR2X1_202 VDD GND POR2X1_202/B POR2X1_202/A POR2X1_206/A POR2X1_202/m4_208_n4# POR2X1_202/O
+ POR2X1_202/CTRL2 POR2X1_202/a_16_28# POR2X1_202/CTRL POR2X1_202/a_76_344# POR2X1_202/a_56_344#
+ POR2X1
XPOR2X1_224 VDD GND POR2X1_32/A POR2X1_394/A POR2X1_224/Y POR2X1_224/m4_208_n4# POR2X1_224/O
+ POR2X1_224/CTRL2 POR2X1_224/a_16_28# POR2X1_224/CTRL POR2X1_224/a_76_344# POR2X1_224/a_56_344#
+ POR2X1
XPOR2X1_213 VDD GND POR2X1_213/B POR2X1_210/Y POR2X1_220/A POR2X1_213/m4_208_n4# POR2X1_213/O
+ POR2X1_213/CTRL2 POR2X1_213/a_16_28# POR2X1_213/CTRL POR2X1_213/a_76_344# POR2X1_213/a_56_344#
+ POR2X1
XPOR2X1_235 VDD GND PAND2X1_63/B POR2X1_85/Y POR2X1_235/Y POR2X1_85/m4_208_n4# POR2X1_235/O
+ POR2X1_235/CTRL2 POR2X1_235/a_16_28# POR2X1_235/CTRL POR2X1_235/a_76_344# POR2X1_235/a_56_344#
+ POR2X1
XPOR2X1_268 VDD GND POR2X1_39/B POR2X1_93/A POR2X1_268/Y POR2X1_268/m4_208_n4# POR2X1_268/O
+ POR2X1_268/CTRL2 POR2X1_268/a_16_28# POR2X1_268/CTRL POR2X1_268/a_76_344# POR2X1_268/a_56_344#
+ POR2X1
XPOR2X1_257 VDD GND POR2X1_20/B POR2X1_257/A POR2X1_257/Y POR2X1_257/m4_208_n4# POR2X1_257/O
+ POR2X1_257/CTRL2 POR2X1_257/a_16_28# POR2X1_257/CTRL POR2X1_257/a_76_344# POR2X1_257/a_56_344#
+ POR2X1
XPOR2X1_246 VDD GND POR2X1_9/Y POR2X1_245/Y POR2X1_246/Y POR2X1_246/m4_208_n4# POR2X1_246/O
+ POR2X1_246/CTRL2 POR2X1_246/a_16_28# POR2X1_246/CTRL POR2X1_246/a_76_344# POR2X1_246/a_56_344#
+ POR2X1
XPOR2X1_279 VDD GND POR2X1_57/A POR2X1_257/A POR2X1_279/Y POR2X1_279/m4_208_n4# POR2X1_279/O
+ POR2X1_279/CTRL2 POR2X1_279/a_16_28# POR2X1_279/CTRL POR2X1_279/a_76_344# POR2X1_279/a_56_344#
+ POR2X1
XPAND2X1_209 VDD GND POR2X1_152/Y PAND2X1_209/A PAND2X1_213/A PAND2X1_209/a_16_344#
+ PAND2X1_209/m4_208_n4# PAND2X1_209/O PAND2X1_209/a_56_28# PAND2X1_209/CTRL2 PAND2X1_209/CTRL
+ PAND2X1_209/a_76_28# PAND2X1
XPOR2X1_780 VDD GND POR2X1_780/B POR2X1_780/A POR2X1_783/A POR2X1_780/m4_208_n4# POR2X1_780/O
+ POR2X1_780/CTRL2 POR2X1_780/a_16_28# POR2X1_780/CTRL POR2X1_780/a_76_344# POR2X1_780/a_56_344#
+ POR2X1
XPOR2X1_791 VDD GND POR2X1_791/B POR2X1_791/A POR2X1_791/Y POR2X1_791/m4_208_n4# POR2X1_791/O
+ POR2X1_791/CTRL2 POR2X1_791/a_16_28# POR2X1_791/CTRL POR2X1_791/a_76_344# POR2X1_791/a_56_344#
+ POR2X1
XPAND2X1_710 VDD GND POR2X1_701/Y POR2X1_700/Y PAND2X1_711/B PAND2X1_710/a_16_344#
+ POR2X1_701/m4_208_n4# PAND2X1_710/O PAND2X1_710/a_56_28# PAND2X1_710/CTRL2 PAND2X1_710/CTRL
+ PAND2X1_710/a_76_28# PAND2X1
XPAND2X1_732 VDD GND PAND2X1_725/Y PAND2X1_732/A PAND2X1_738/B PAND2X1_732/a_16_344#
+ PAND2X1_732/m4_208_n4# PAND2X1_732/O PAND2X1_732/a_56_28# PAND2X1_732/CTRL2 PAND2X1_732/CTRL
+ PAND2X1_732/a_76_28# PAND2X1
XPAND2X1_721 VDD GND PAND2X1_721/B PAND2X1_673/Y PAND2X1_734/B PAND2X1_721/a_16_344#
+ PAND2X1_721/m4_208_n4# PAND2X1_721/O PAND2X1_721/a_56_28# PAND2X1_721/CTRL2 PAND2X1_721/CTRL
+ PAND2X1_721/a_76_28# PAND2X1
XPAND2X1_754 VDD GND POR2X1_614/Y PAND2X1_69/A POR2X1_790/A PAND2X1_754/a_16_344#
+ PAND2X1_754/m4_208_n4# PAND2X1_754/O PAND2X1_754/a_56_28# PAND2X1_754/CTRL2 PAND2X1_754/CTRL
+ PAND2X1_754/a_76_28# PAND2X1
XPAND2X1_743 VDD GND POR2X1_407/A POR2X1_66/B POR2X1_780/B PAND2X1_743/a_16_344# PAND2X1_743/m4_208_n4#
+ PAND2X1_743/O PAND2X1_743/a_56_28# PAND2X1_743/CTRL2 PAND2X1_743/CTRL PAND2X1_743/a_76_28#
+ PAND2X1
XPAND2X1_765 VDD GND POR2X1_78/B POR2X1_260/B POR2X1_770/B PAND2X1_765/a_16_344# PAND2X1_765/m4_208_n4#
+ PAND2X1_765/O PAND2X1_765/a_56_28# PAND2X1_765/CTRL2 PAND2X1_765/CTRL PAND2X1_765/a_76_28#
+ PAND2X1
XPAND2X1_798 VDD GND PAND2X1_798/B PAND2X1_354/A PAND2X1_798/Y PAND2X1_798/a_16_344#
+ PAND2X1_798/m4_208_n4# PAND2X1_798/O PAND2X1_798/a_56_28# PAND2X1_798/CTRL2 PAND2X1_798/CTRL
+ PAND2X1_798/a_76_28# PAND2X1
XPAND2X1_787 VDD GND PAND2X1_556/B PAND2X1_787/A PAND2X1_787/Y PAND2X1_787/a_16_344#
+ PAND2X1_787/m4_208_n4# PAND2X1_787/O PAND2X1_787/a_56_28# PAND2X1_787/CTRL2 PAND2X1_787/CTRL
+ PAND2X1_787/a_76_28# PAND2X1
XPAND2X1_776 VDD GND POR2X1_238/Y POR2X1_164/Y PAND2X1_776/Y PAND2X1_776/a_16_344#
+ PAND2X1_776/m4_208_n4# PAND2X1_776/O PAND2X1_776/a_56_28# PAND2X1_776/CTRL2 PAND2X1_776/CTRL
+ PAND2X1_776/a_76_28# PAND2X1
XPAND2X1_540 VDD GND POR2X1_183/Y POR2X1_178/Y PAND2X1_553/A PAND2X1_540/a_16_344#
+ PAND2X1_540/m4_208_n4# PAND2X1_540/O PAND2X1_540/a_56_28# PAND2X1_540/CTRL2 PAND2X1_540/CTRL
+ PAND2X1_540/a_76_28# PAND2X1
XPAND2X1_573 VDD GND PAND2X1_573/B PAND2X1_404/Y PAND2X1_575/A PAND2X1_573/a_16_344#
+ POR2X1_72/m4_208_n4# PAND2X1_573/O PAND2X1_573/a_56_28# PAND2X1_573/CTRL2 PAND2X1_573/CTRL
+ PAND2X1_573/a_76_28# PAND2X1
XPAND2X1_562 VDD GND PAND2X1_562/B PAND2X1_555/Y PAND2X1_562/Y PAND2X1_562/a_16_344#
+ PAND2X1_562/m4_208_n4# PAND2X1_562/O PAND2X1_562/a_56_28# PAND2X1_562/CTRL2 PAND2X1_562/CTRL
+ PAND2X1_562/a_76_28# PAND2X1
XPAND2X1_551 VDD GND PAND2X1_545/Y PAND2X1_551/A PAND2X1_551/Y PAND2X1_551/a_16_344#
+ POR2X1_765/m4_208_n4# PAND2X1_551/O PAND2X1_551/a_56_28# PAND2X1_551/CTRL2 PAND2X1_551/CTRL
+ PAND2X1_551/a_76_28# PAND2X1
XPAND2X1_595 VDD GND POR2X1_249/Y POR2X1_66/A POR2X1_643/A PAND2X1_595/a_16_344# PAND2X1_595/m4_208_n4#
+ PAND2X1_595/O PAND2X1_595/a_56_28# PAND2X1_595/CTRL2 PAND2X1_595/CTRL PAND2X1_595/a_76_28#
+ PAND2X1
XPAND2X1_584 VDD GND PAND2X1_52/B PAND2X1_6/Y POR2X1_636/A PAND2X1_584/a_16_344# POR2X1_771/m4_208_n4#
+ PAND2X1_584/O PAND2X1_584/a_56_28# PAND2X1_584/CTRL2 PAND2X1_584/CTRL PAND2X1_584/a_76_28#
+ PAND2X1
XPAND2X1_381 VDD GND POR2X1_260/B INPUT_3 PAND2X1_381/Y PAND2X1_381/a_16_344# PAND2X1_381/m4_208_n4#
+ PAND2X1_381/O PAND2X1_381/a_56_28# PAND2X1_381/CTRL2 PAND2X1_381/CTRL PAND2X1_381/a_76_28#
+ PAND2X1
XPAND2X1_370 VDD GND POR2X1_369/Y POR2X1_309/Y PAND2X1_787/A PAND2X1_370/a_16_344#
+ PAND2X1_370/m4_208_n4# PAND2X1_370/O PAND2X1_370/a_56_28# PAND2X1_370/CTRL2 PAND2X1_370/CTRL
+ PAND2X1_370/a_76_28# PAND2X1
XPAND2X1_392 VDD GND PAND2X1_392/B PAND2X1_390/Y PAND2X1_474/A PAND2X1_392/a_16_344#
+ PAND2X1_392/m4_208_n4# PAND2X1_392/O PAND2X1_392/a_56_28# PAND2X1_392/CTRL2 PAND2X1_392/CTRL
+ PAND2X1_392/a_76_28# PAND2X1
XPAND2X1_18 VDD GND PAND2X1_18/B PAND2X1_11/Y PAND2X1_20/A PAND2X1_18/a_16_344# PAND2X1_18/m4_208_n4#
+ PAND2X1_18/O PAND2X1_18/a_56_28# PAND2X1_18/CTRL2 PAND2X1_18/CTRL PAND2X1_18/a_76_28#
+ PAND2X1
XPAND2X1_29 VDD GND POR2X1_38/B PAND2X1_8/Y POR2X1_87/B PAND2X1_29/a_16_344# PAND2X1_29/m4_208_n4#
+ PAND2X1_29/O PAND2X1_29/a_56_28# PAND2X1_29/CTRL2 PAND2X1_29/CTRL PAND2X1_29/a_76_28#
+ PAND2X1
XPOR2X1_609 VDD GND POR2X1_60/A POR2X1_609/A POR2X1_609/Y POR2X1_609/m4_208_n4# POR2X1_609/O
+ POR2X1_609/CTRL2 POR2X1_609/a_16_28# POR2X1_609/CTRL POR2X1_609/a_76_344# POR2X1_609/a_56_344#
+ POR2X1
XPOR2X1_406 VDD GND POR2X1_96/A POR2X1_406/A POR2X1_406/Y POR2X1_406/m4_208_n4# POR2X1_406/O
+ POR2X1_406/CTRL2 POR2X1_406/a_16_28# POR2X1_406/CTRL POR2X1_406/a_76_344# POR2X1_406/a_56_344#
+ POR2X1
XPOR2X1_417 VDD GND POR2X1_48/A POR2X1_283/A POR2X1_417/Y POR2X1_417/m4_208_n4# POR2X1_417/O
+ POR2X1_417/CTRL2 POR2X1_417/a_16_28# POR2X1_417/CTRL POR2X1_417/a_76_344# POR2X1_417/a_56_344#
+ POR2X1
XPOR2X1_428 VDD GND POR2X1_32/A POR2X1_236/Y POR2X1_428/Y POR2X1_428/m4_208_n4# POR2X1_428/O
+ POR2X1_428/CTRL2 POR2X1_428/a_16_28# POR2X1_428/CTRL POR2X1_428/a_76_344# POR2X1_428/a_56_344#
+ POR2X1
XPOR2X1_439 VDD GND POR2X1_180/A POR2X1_544/A POR2X1_439/Y POR2X1_439/m4_208_n4# POR2X1_439/O
+ POR2X1_439/CTRL2 POR2X1_439/a_16_28# POR2X1_439/CTRL POR2X1_439/a_76_344# POR2X1_439/a_56_344#
+ POR2X1
XPOR2X1_214 VDD GND POR2X1_214/B POR2X1_208/Y POR2X1_219/B POR2X1_214/m4_208_n4# POR2X1_214/O
+ POR2X1_214/CTRL2 POR2X1_214/a_16_28# POR2X1_214/CTRL POR2X1_214/a_76_344# POR2X1_214/a_56_344#
+ POR2X1
XPOR2X1_203 VDD GND PAND2X1_72/Y POR2X1_76/Y POR2X1_203/Y POR2X1_203/m4_208_n4# POR2X1_203/O
+ POR2X1_203/CTRL2 POR2X1_203/a_16_28# POR2X1_203/CTRL POR2X1_203/a_76_344# POR2X1_203/a_56_344#
+ POR2X1
XPOR2X1_225 VDD GND INPUT_1 POR2X1_5/Y POR2X1_283/A POR2X1_225/m4_208_n4# POR2X1_225/O
+ POR2X1_225/CTRL2 POR2X1_225/a_16_28# POR2X1_225/CTRL POR2X1_225/a_76_344# POR2X1_225/a_56_344#
+ POR2X1
XPOR2X1_236 VDD GND POR2X1_5/Y POR2X1_38/B POR2X1_236/Y POR2X1_236/m4_208_n4# POR2X1_236/O
+ POR2X1_236/CTRL2 POR2X1_236/a_16_28# POR2X1_236/CTRL POR2X1_236/a_76_344# POR2X1_236/a_56_344#
+ POR2X1
XPOR2X1_247 VDD GND PAND2X1_6/Y POR2X1_294/B POR2X1_247/Y POR2X1_247/m4_208_n4# POR2X1_247/O
+ POR2X1_247/CTRL2 POR2X1_247/a_16_28# POR2X1_247/CTRL POR2X1_247/a_76_344# POR2X1_247/a_56_344#
+ POR2X1
XPOR2X1_258 VDD GND POR2X1_77/Y POR2X1_416/B POR2X1_258/Y POR2X1_258/m4_208_n4# POR2X1_258/O
+ POR2X1_258/CTRL2 POR2X1_258/a_16_28# POR2X1_258/CTRL POR2X1_258/a_76_344# POR2X1_258/a_56_344#
+ POR2X1
XPOR2X1_269 VDD GND POR2X1_383/A POR2X1_269/A POR2X1_269/Y POR2X1_269/m4_208_n4# POR2X1_269/O
+ POR2X1_269/CTRL2 POR2X1_269/a_16_28# POR2X1_269/CTRL POR2X1_269/a_76_344# POR2X1_269/a_56_344#
+ POR2X1
XPOR2X1_781 VDD GND POR2X1_781/B POR2X1_781/A POR2X1_782/A POR2X1_781/m4_208_n4# POR2X1_781/O
+ POR2X1_781/CTRL2 POR2X1_781/a_16_28# POR2X1_781/CTRL POR2X1_781/a_76_344# POR2X1_781/a_56_344#
+ POR2X1
XPOR2X1_770 VDD GND POR2X1_770/B POR2X1_770/A POR2X1_771/A POR2X1_770/m4_208_n4# POR2X1_770/O
+ POR2X1_770/CTRL2 POR2X1_770/a_16_28# POR2X1_770/CTRL POR2X1_770/a_76_344# POR2X1_770/a_56_344#
+ POR2X1
XPOR2X1_792 VDD GND POR2X1_792/B POR2X1_791/Y POR2X1_805/B POR2X1_792/m4_208_n4# POR2X1_792/O
+ POR2X1_792/CTRL2 POR2X1_792/a_16_28# POR2X1_792/CTRL POR2X1_792/a_76_344# POR2X1_792/a_56_344#
+ POR2X1
XPAND2X1_700 VDD GND PAND2X1_90/Y PAND2X1_60/B POR2X1_710/B PAND2X1_700/a_16_344#
+ PAND2X1_700/m4_208_n4# PAND2X1_700/O PAND2X1_700/a_56_28# PAND2X1_700/CTRL2 PAND2X1_700/CTRL
+ PAND2X1_700/a_76_28# PAND2X1
XPAND2X1_711 VDD GND PAND2X1_711/B PAND2X1_711/A PAND2X1_726/B PAND2X1_711/a_16_344#
+ POR2X1_428/m4_208_n4# PAND2X1_711/O PAND2X1_711/a_56_28# PAND2X1_711/CTRL2 PAND2X1_711/CTRL
+ PAND2X1_711/a_76_28# PAND2X1
XPAND2X1_722 VDD GND PAND2X1_719/Y PAND2X1_718/Y PAND2X1_733/A PAND2X1_722/a_16_344#
+ PAND2X1_722/m4_208_n4# PAND2X1_722/O PAND2X1_722/a_56_28# PAND2X1_722/CTRL2 PAND2X1_722/CTRL
+ PAND2X1_722/a_76_28# PAND2X1
XPAND2X1_733 VDD GND PAND2X1_723/Y PAND2X1_733/A PAND2X1_733/Y PAND2X1_733/a_16_344#
+ PAND2X1_733/m4_208_n4# PAND2X1_733/O PAND2X1_733/a_56_28# PAND2X1_733/CTRL2 PAND2X1_733/CTRL
+ PAND2X1_733/a_76_28# PAND2X1
XPAND2X1_755 VDD GND POR2X1_664/Y PAND2X1_60/B POR2X1_791/B PAND2X1_755/a_16_344#
+ PAND2X1_755/m4_208_n4# PAND2X1_755/O PAND2X1_755/a_56_28# PAND2X1_755/CTRL2 PAND2X1_755/CTRL
+ PAND2X1_755/a_76_28# PAND2X1
XPAND2X1_744 VDD GND POR2X1_532/A PAND2X1_57/B POR2X1_780/A PAND2X1_744/a_16_344#
+ PAND2X1_744/m4_208_n4# PAND2X1_744/O PAND2X1_744/a_56_28# PAND2X1_744/CTRL2 PAND2X1_744/CTRL
+ PAND2X1_744/a_76_28# PAND2X1
XPAND2X1_799 VDD GND PAND2X1_593/Y PAND2X1_539/Y PAND2X1_802/B PAND2X1_799/a_16_344#
+ PAND2X1_799/m4_208_n4# PAND2X1_799/O PAND2X1_799/a_56_28# PAND2X1_799/CTRL2 PAND2X1_799/CTRL
+ PAND2X1_799/a_76_28# PAND2X1
XPAND2X1_777 VDD GND POR2X1_305/Y POR2X1_245/Y PAND2X1_784/A PAND2X1_777/a_16_344#
+ PAND2X1_777/m4_208_n4# PAND2X1_777/O PAND2X1_777/a_56_28# PAND2X1_777/CTRL2 PAND2X1_777/CTRL
+ PAND2X1_777/a_76_28# PAND2X1
XPAND2X1_766 VDD GND PAND2X1_90/Y PAND2X1_65/B POR2X1_770/A PAND2X1_766/a_16_344#
+ PAND2X1_766/m4_208_n4# PAND2X1_766/O PAND2X1_766/a_56_28# PAND2X1_766/CTRL2 PAND2X1_766/CTRL
+ PAND2X1_766/a_76_28# PAND2X1
XPAND2X1_788 VDD GND PAND2X1_602/Y POR2X1_533/Y PAND2X1_794/B PAND2X1_788/a_16_344#
+ PAND2X1_788/m4_208_n4# PAND2X1_788/O PAND2X1_788/a_56_28# PAND2X1_788/CTRL2 PAND2X1_788/CTRL
+ PAND2X1_788/a_76_28# PAND2X1
XPAND2X1_530 VDD GND POR2X1_590/A PAND2X1_69/A POR2X1_548/A PAND2X1_530/a_16_344#
+ POR2X1_548/m4_208_n4# PAND2X1_530/O PAND2X1_530/a_56_28# PAND2X1_530/CTRL2 PAND2X1_530/CTRL
+ PAND2X1_530/a_76_28# PAND2X1
XPAND2X1_574 VDD GND POR2X1_516/Y PAND2X1_657/B PAND2X1_575/B PAND2X1_574/a_16_344#
+ PAND2X1_574/m4_208_n4# PAND2X1_574/O PAND2X1_574/a_56_28# PAND2X1_574/CTRL2 PAND2X1_574/CTRL
+ PAND2X1_574/a_76_28# PAND2X1
XPAND2X1_541 VDD GND POR2X1_272/Y POR2X1_255/Y PAND2X1_553/B PAND2X1_541/a_16_344#
+ PAND2X1_344/m4_208_n4# PAND2X1_541/O PAND2X1_541/a_56_28# PAND2X1_541/CTRL2 PAND2X1_541/CTRL
+ PAND2X1_541/a_76_28# PAND2X1
XPAND2X1_563 VDD GND PAND2X1_563/B PAND2X1_563/A PAND2X1_570/B PAND2X1_563/a_16_344#
+ PAND2X1_562/m4_208_n4# PAND2X1_563/O PAND2X1_563/a_56_28# PAND2X1_563/CTRL2 PAND2X1_563/CTRL
+ PAND2X1_563/a_76_28# PAND2X1
XPAND2X1_552 VDD GND PAND2X1_552/B PAND2X1_552/A PAND2X1_564/B PAND2X1_552/a_16_344#
+ PAND2X1_552/m4_208_n4# PAND2X1_552/O PAND2X1_552/a_56_28# PAND2X1_552/CTRL2 PAND2X1_552/CTRL
+ PAND2X1_552/a_76_28# PAND2X1
XPAND2X1_585 VDD GND POR2X1_294/A PAND2X1_58/A POR2X1_637/B PAND2X1_585/a_16_344#
+ PAND2X1_585/m4_208_n4# PAND2X1_585/O PAND2X1_585/a_56_28# PAND2X1_585/CTRL2 PAND2X1_585/CTRL
+ PAND2X1_585/a_76_28# PAND2X1
XPAND2X1_596 VDD GND POR2X1_329/A POR2X1_57/A POR2X1_597/A PAND2X1_596/a_16_344# PAND2X1_596/m4_208_n4#
+ PAND2X1_596/O PAND2X1_596/a_56_28# PAND2X1_596/CTRL2 PAND2X1_596/CTRL PAND2X1_596/a_76_28#
+ PAND2X1
XPAND2X1_382 VDD GND PAND2X1_381/Y POR2X1_29/A POR2X1_391/B PAND2X1_382/a_16_344#
+ PAND2X1_382/m4_208_n4# PAND2X1_382/O PAND2X1_382/a_56_28# PAND2X1_382/CTRL2 PAND2X1_382/CTRL
+ PAND2X1_382/a_76_28# PAND2X1
XPAND2X1_360 VDD GND PAND2X1_347/Y PAND2X1_860/A PAND2X1_360/Y PAND2X1_360/a_16_344#
+ PAND2X1_360/m4_208_n4# PAND2X1_360/O PAND2X1_360/a_56_28# PAND2X1_360/CTRL2 PAND2X1_360/CTRL
+ PAND2X1_360/a_76_28# PAND2X1
XPAND2X1_371 VDD GND PAND2X1_32/B POR2X1_68/B POR2X1_778/B PAND2X1_371/a_16_344# PAND2X1_371/m4_208_n4#
+ PAND2X1_371/O PAND2X1_371/a_56_28# PAND2X1_371/CTRL2 PAND2X1_371/CTRL PAND2X1_371/a_76_28#
+ PAND2X1
XPAND2X1_393 VDD GND PAND2X1_41/B PAND2X1_39/B POR2X1_400/B PAND2X1_393/a_16_344#
+ PAND2X1_393/m4_208_n4# PAND2X1_393/O PAND2X1_393/a_56_28# PAND2X1_393/CTRL2 PAND2X1_393/CTRL
+ PAND2X1_393/a_76_28# PAND2X1
XPAND2X1_19 VDD GND POR2X1_68/B POR2X1_4/Y PAND2X1_19/Y PAND2X1_19/a_16_344# PAND2X1_19/m4_208_n4#
+ PAND2X1_19/O PAND2X1_19/a_56_28# PAND2X1_19/CTRL2 PAND2X1_19/CTRL PAND2X1_19/a_76_28#
+ PAND2X1
XPAND2X1_190 VDD GND POR2X1_184/Y POR2X1_183/Y PAND2X1_190/Y PAND2X1_190/a_16_344#
+ POR2X1_131/m4_208_n4# PAND2X1_190/O PAND2X1_190/a_56_28# PAND2X1_190/CTRL2 PAND2X1_190/CTRL
+ PAND2X1_190/a_76_28# PAND2X1
XPOR2X1_407 VDD GND PAND2X1_55/Y POR2X1_407/A POR2X1_407/Y POR2X1_407/m4_208_n4# POR2X1_407/O
+ POR2X1_407/CTRL2 POR2X1_407/a_16_28# POR2X1_407/CTRL POR2X1_407/a_76_344# POR2X1_407/a_56_344#
+ POR2X1
XPOR2X1_429 VDD GND INPUT_7 POR2X1_12/A POR2X1_430/A POR2X1_429/m4_208_n4# POR2X1_429/O
+ POR2X1_429/CTRL2 POR2X1_429/a_16_28# POR2X1_429/CTRL POR2X1_429/a_76_344# POR2X1_429/a_56_344#
+ POR2X1
XPOR2X1_418 VDD GND POR2X1_16/A POR2X1_52/A POR2X1_418/Y POR2X1_418/m4_208_n4# POR2X1_418/O
+ POR2X1_418/CTRL2 POR2X1_418/a_16_28# POR2X1_418/CTRL POR2X1_418/a_76_344# POR2X1_418/a_56_344#
+ POR2X1
XPOR2X1_215 VDD GND POR2X1_205/Y POR2X1_215/A POR2X1_215/Y POR2X1_215/m4_208_n4# POR2X1_215/O
+ POR2X1_215/CTRL2 POR2X1_215/a_16_28# POR2X1_215/CTRL POR2X1_215/a_76_344# POR2X1_215/a_56_344#
+ POR2X1
XPOR2X1_204 VDD GND PAND2X1_79/Y POR2X1_84/Y POR2X1_205/A POR2X1_204/m4_208_n4# POR2X1_204/O
+ POR2X1_204/CTRL2 POR2X1_204/a_16_28# POR2X1_204/CTRL POR2X1_204/a_76_344# POR2X1_204/a_56_344#
+ POR2X1
XPOR2X1_259 VDD GND POR2X1_259/B POR2X1_259/A POR2X1_555/B PAND2X1_89/m4_208_n4# POR2X1_259/O
+ POR2X1_259/CTRL2 POR2X1_259/a_16_28# POR2X1_259/CTRL POR2X1_259/a_76_344# POR2X1_259/a_56_344#
+ POR2X1
XPOR2X1_226 VDD GND POR2X1_20/B POR2X1_283/A POR2X1_226/Y POR2X1_226/m4_208_n4# POR2X1_226/O
+ POR2X1_226/CTRL2 POR2X1_226/a_16_28# POR2X1_226/CTRL POR2X1_226/a_76_344# POR2X1_226/a_56_344#
+ POR2X1
XPOR2X1_237 VDD GND POR2X1_83/B POR2X1_236/Y POR2X1_237/Y POR2X1_237/m4_208_n4# POR2X1_237/O
+ POR2X1_237/CTRL2 POR2X1_237/a_16_28# POR2X1_237/CTRL POR2X1_237/a_76_344# POR2X1_237/a_56_344#
+ POR2X1
XPOR2X1_248 VDD GND POR2X1_48/A POR2X1_248/A POR2X1_248/Y POR2X1_248/m4_208_n4# POR2X1_248/O
+ POR2X1_248/CTRL2 POR2X1_248/a_16_28# POR2X1_248/CTRL POR2X1_248/a_76_344# POR2X1_248/a_56_344#
+ POR2X1
XPOR2X1_760 VDD GND POR2X1_65/A POR2X1_760/A POR2X1_760/Y POR2X1_760/m4_208_n4# POR2X1_760/O
+ POR2X1_760/CTRL2 POR2X1_760/a_16_28# POR2X1_760/CTRL POR2X1_760/a_76_344# POR2X1_760/a_56_344#
+ POR2X1
XPOR2X1_771 VDD GND POR2X1_769/Y POR2X1_771/A POR2X1_774/B POR2X1_771/m4_208_n4# POR2X1_771/O
+ POR2X1_771/CTRL2 POR2X1_771/a_16_28# POR2X1_771/CTRL POR2X1_771/a_76_344# POR2X1_771/a_56_344#
+ POR2X1
XPOR2X1_782 VDD GND POR2X1_782/B POR2X1_782/A POR2X1_797/A POR2X1_782/m4_208_n4# POR2X1_782/O
+ POR2X1_782/CTRL2 POR2X1_782/a_16_28# POR2X1_782/CTRL POR2X1_782/a_76_344# POR2X1_782/a_56_344#
+ POR2X1
XPOR2X1_793 VDD GND POR2X1_789/Y POR2X1_793/A POR2X1_805/A POR2X1_793/m4_208_n4# POR2X1_793/O
+ POR2X1_793/CTRL2 POR2X1_793/a_16_28# POR2X1_793/CTRL POR2X1_793/a_76_344# POR2X1_793/a_56_344#
+ POR2X1
XPAND2X1_723 VDD GND PAND2X1_717/Y PAND2X1_723/A PAND2X1_723/Y PAND2X1_723/a_16_344#
+ PAND2X1_216/m4_208_n4# PAND2X1_723/O PAND2X1_723/a_56_28# PAND2X1_723/CTRL2 PAND2X1_723/CTRL
+ PAND2X1_723/a_76_28# PAND2X1
XPAND2X1_701 VDD GND POR2X1_383/A PAND2X1_57/B POR2X1_710/A PAND2X1_701/a_16_344#
+ PAND2X1_701/m4_208_n4# PAND2X1_701/O PAND2X1_701/a_56_28# PAND2X1_701/CTRL2 PAND2X1_701/CTRL
+ PAND2X1_701/a_76_28# PAND2X1
XPAND2X1_712 VDD GND PAND2X1_712/B PAND2X1_707/Y PAND2X1_725/A PAND2X1_712/a_16_344#
+ PAND2X1_712/m4_208_n4# PAND2X1_712/O PAND2X1_712/a_56_28# PAND2X1_712/CTRL2 PAND2X1_712/CTRL
+ PAND2X1_712/a_76_28# PAND2X1
XPAND2X1_734 VDD GND PAND2X1_734/B POR2X1_406/Y PAND2X1_737/B PAND2X1_734/a_16_344#
+ PAND2X1_734/m4_208_n4# PAND2X1_734/O PAND2X1_734/a_56_28# PAND2X1_734/CTRL2 PAND2X1_734/CTRL
+ PAND2X1_734/a_76_28# PAND2X1
XPAND2X1_745 VDD GND POR2X1_750/B PAND2X1_41/B POR2X1_781/B PAND2X1_745/a_16_344#
+ PAND2X1_745/m4_208_n4# PAND2X1_745/O PAND2X1_745/a_56_28# PAND2X1_745/CTRL2 PAND2X1_745/CTRL
+ PAND2X1_745/a_76_28# PAND2X1
XPAND2X1_756 VDD GND POR2X1_669/B POR2X1_411/B POR2X1_757/A PAND2X1_756/a_16_344#
+ PAND2X1_756/m4_208_n4# PAND2X1_756/O PAND2X1_756/a_56_28# PAND2X1_756/CTRL2 PAND2X1_756/CTRL
+ PAND2X1_756/a_76_28# PAND2X1
XPAND2X1_767 VDD GND POR2X1_78/Y POR2X1_66/B POR2X1_773/B PAND2X1_767/a_16_344# PAND2X1_491/m4_208_n4#
+ PAND2X1_767/O PAND2X1_767/a_56_28# PAND2X1_767/CTRL2 PAND2X1_767/CTRL PAND2X1_767/a_76_28#
+ PAND2X1
XPAND2X1_789 VDD GND POR2X1_751/Y POR2X1_748/Y PAND2X1_793/A PAND2X1_789/a_16_344#
+ PAND2X1_793/m4_208_n4# PAND2X1_789/O PAND2X1_789/a_56_28# PAND2X1_789/CTRL2 PAND2X1_789/CTRL
+ PAND2X1_789/a_76_28# PAND2X1
XPAND2X1_778 VDD GND POR2X1_496/Y POR2X1_372/A PAND2X1_778/Y PAND2X1_778/a_16_344#
+ PAND2X1_778/m4_208_n4# PAND2X1_778/O PAND2X1_778/a_56_28# PAND2X1_778/CTRL2 PAND2X1_778/CTRL
+ PAND2X1_778/a_76_28# PAND2X1
XPOR2X1_590 VDD GND PAND2X1_39/B POR2X1_590/A POR2X1_590/Y POR2X1_590/m4_208_n4# POR2X1_590/O
+ POR2X1_590/CTRL2 POR2X1_590/a_16_28# POR2X1_590/CTRL POR2X1_590/a_76_344# POR2X1_590/a_56_344#
+ POR2X1
XPAND2X1_531 VDD GND PAND2X1_73/Y PAND2X1_41/B POR2X1_549/B PAND2X1_531/a_16_344#
+ PAND2X1_531/m4_208_n4# PAND2X1_531/O PAND2X1_531/a_56_28# PAND2X1_531/CTRL2 PAND2X1_531/CTRL
+ PAND2X1_531/a_76_28# PAND2X1
XPAND2X1_520 VDD GND POR2X1_519/Y POR2X1_518/Y PAND2X1_642/B PAND2X1_520/a_16_344#
+ PAND2X1_520/m4_208_n4# PAND2X1_520/O PAND2X1_520/a_56_28# PAND2X1_520/CTRL2 PAND2X1_520/CTRL
+ PAND2X1_520/a_76_28# PAND2X1
XPAND2X1_553 VDD GND PAND2X1_553/B PAND2X1_553/A PAND2X1_563/A PAND2X1_553/a_16_344#
+ PAND2X1_553/m4_208_n4# PAND2X1_553/O PAND2X1_553/a_56_28# PAND2X1_553/CTRL2 PAND2X1_553/CTRL
+ PAND2X1_553/a_76_28# PAND2X1
XPAND2X1_542 VDD GND POR2X1_312/Y POR2X1_280/Y PAND2X1_552/A PAND2X1_542/a_16_344#
+ PAND2X1_542/m4_208_n4# PAND2X1_542/O PAND2X1_542/a_56_28# PAND2X1_542/CTRL2 PAND2X1_542/CTRL
+ PAND2X1_542/a_76_28# PAND2X1
XPAND2X1_564 VDD GND PAND2X1_564/B PAND2X1_551/Y PAND2X1_569/A PAND2X1_564/a_16_344#
+ PAND2X1_564/m4_208_n4# PAND2X1_564/O PAND2X1_564/a_56_28# PAND2X1_564/CTRL2 PAND2X1_564/CTRL
+ PAND2X1_564/a_76_28# PAND2X1
XPAND2X1_575 VDD GND PAND2X1_575/B PAND2X1_575/A PAND2X1_579/A PAND2X1_575/a_16_344#
+ PAND2X1_575/m4_208_n4# PAND2X1_575/O PAND2X1_575/a_56_28# PAND2X1_575/CTRL2 PAND2X1_575/CTRL
+ PAND2X1_575/a_76_28# PAND2X1
XPAND2X1_586 VDD GND POR2X1_130/A PAND2X1_72/A POR2X1_637/A PAND2X1_586/a_16_344#
+ PAND2X1_586/m4_208_n4# PAND2X1_586/O PAND2X1_586/a_56_28# PAND2X1_586/CTRL2 PAND2X1_586/CTRL
+ PAND2X1_586/a_76_28# PAND2X1
XPAND2X1_597 VDD GND POR2X1_596/Y POR2X1_294/B POR2X1_644/B PAND2X1_597/a_16_344#
+ PAND2X1_597/m4_208_n4# PAND2X1_597/O PAND2X1_597/a_56_28# PAND2X1_597/CTRL2 PAND2X1_597/CTRL
+ PAND2X1_597/a_76_28# PAND2X1
XPAND2X1_350 VDD GND PAND2X1_341/Y PAND2X1_350/A PAND2X1_358/A PAND2X1_350/a_16_344#
+ PAND2X1_350/m4_208_n4# PAND2X1_350/O PAND2X1_350/a_56_28# PAND2X1_350/CTRL2 PAND2X1_350/CTRL
+ PAND2X1_350/a_76_28# PAND2X1
XPAND2X1_361 VDD GND PAND2X1_473/B PAND2X1_267/Y PAND2X1_362/B PAND2X1_361/a_16_344#
+ PAND2X1_361/m4_208_n4# PAND2X1_361/O PAND2X1_361/a_56_28# PAND2X1_361/CTRL2 PAND2X1_361/CTRL
+ PAND2X1_361/a_76_28# PAND2X1
XPAND2X1_372 VDD GND POR2X1_778/B D_INPUT_1 POR2X1_458/B PAND2X1_372/a_16_344# PAND2X1_372/m4_208_n4#
+ PAND2X1_372/O PAND2X1_372/a_56_28# PAND2X1_372/CTRL2 PAND2X1_372/CTRL PAND2X1_372/a_76_28#
+ PAND2X1
XPAND2X1_383 VDD GND POR2X1_236/Y POR2X1_90/Y POR2X1_384/A PAND2X1_383/a_16_344# PAND2X1_383/m4_208_n4#
+ PAND2X1_383/O PAND2X1_383/a_56_28# PAND2X1_383/CTRL2 PAND2X1_383/CTRL PAND2X1_383/a_76_28#
+ PAND2X1
XPAND2X1_394 VDD GND POR2X1_532/A PAND2X1_48/B POR2X1_400/A PAND2X1_394/a_16_344#
+ PAND2X1_394/m4_208_n4# PAND2X1_394/O PAND2X1_394/a_56_28# PAND2X1_394/CTRL2 PAND2X1_394/CTRL
+ PAND2X1_394/a_76_28# PAND2X1
XPAND2X1_180 VDD GND POR2X1_177/Y POR2X1_176/Y PAND2X1_182/A PAND2X1_180/a_16_344#
+ PAND2X1_180/m4_208_n4# PAND2X1_180/O PAND2X1_180/a_56_28# PAND2X1_180/CTRL2 PAND2X1_180/CTRL
+ PAND2X1_180/a_76_28# PAND2X1
XPAND2X1_191 VDD GND PAND2X1_190/Y POR2X1_187/Y PAND2X1_191/Y PAND2X1_191/a_16_344#
+ PAND2X1_191/m4_208_n4# PAND2X1_191/O PAND2X1_191/a_56_28# PAND2X1_191/CTRL2 PAND2X1_191/CTRL
+ PAND2X1_191/a_76_28# PAND2X1
XPOR2X1_408 VDD GND INPUT_6 POR2X1_22/A POR2X1_408/Y POR2X1_408/m4_208_n4# POR2X1_408/O
+ POR2X1_408/CTRL2 POR2X1_408/a_16_28# POR2X1_408/CTRL POR2X1_408/a_76_344# POR2X1_408/a_56_344#
+ POR2X1
XPOR2X1_419 VDD GND POR2X1_39/B POR2X1_42/Y POR2X1_419/Y POR2X1_419/m4_208_n4# POR2X1_419/O
+ POR2X1_419/CTRL2 POR2X1_419/a_16_28# POR2X1_419/CTRL POR2X1_419/a_76_344# POR2X1_419/a_56_344#
+ POR2X1
XPOR2X1_205 VDD GND POR2X1_203/Y POR2X1_205/A POR2X1_205/Y POR2X1_205/m4_208_n4# POR2X1_205/O
+ POR2X1_205/CTRL2 POR2X1_205/a_16_28# POR2X1_205/CTRL POR2X1_205/a_76_344# POR2X1_205/a_56_344#
+ POR2X1
XPOR2X1_216 VDD GND POR2X1_101/Y POR2X1_116/Y POR2X1_216/Y POR2X1_216/m4_208_n4# POR2X1_216/O
+ POR2X1_216/CTRL2 POR2X1_216/a_16_28# POR2X1_216/CTRL POR2X1_216/a_76_344# POR2X1_216/a_56_344#
+ POR2X1
XPOR2X1_227 VDD GND POR2X1_227/B POR2X1_227/A POR2X1_509/B POR2X1_227/m4_208_n4# POR2X1_227/O
+ POR2X1_227/CTRL2 POR2X1_227/a_16_28# POR2X1_227/CTRL POR2X1_227/a_76_344# POR2X1_227/a_56_344#
+ POR2X1
XPOR2X1_238 VDD GND POR2X1_23/Y POR2X1_52/A POR2X1_238/Y POR2X1_238/m4_208_n4# POR2X1_238/O
+ POR2X1_238/CTRL2 POR2X1_238/a_16_28# POR2X1_238/CTRL POR2X1_238/a_76_344# POR2X1_238/a_56_344#
+ POR2X1
XPOR2X1_249 VDD GND PAND2X1_23/Y PAND2X1_39/B POR2X1_249/Y POR2X1_249/m4_208_n4# POR2X1_249/O
+ POR2X1_249/CTRL2 POR2X1_249/a_16_28# POR2X1_249/CTRL POR2X1_249/a_76_344# POR2X1_249/a_56_344#
+ POR2X1
XPOR2X1_761 VDD GND INPUT_0 POR2X1_761/A POR2X1_761/Y POR2X1_761/m4_208_n4# POR2X1_761/O
+ POR2X1_761/CTRL2 POR2X1_761/a_16_28# POR2X1_761/CTRL POR2X1_761/a_76_344# POR2X1_761/a_56_344#
+ POR2X1
XPOR2X1_750 VDD GND POR2X1_750/B POR2X1_750/A POR2X1_750/Y POR2X1_750/m4_208_n4# POR2X1_750/O
+ POR2X1_750/CTRL2 POR2X1_750/a_16_28# POR2X1_750/CTRL POR2X1_750/a_76_344# POR2X1_750/a_56_344#
+ POR2X1
XPOR2X1_772 VDD GND POR2X1_557/B POR2X1_768/Y POR2X1_773/A POR2X1_772/m4_208_n4# POR2X1_772/O
+ POR2X1_772/CTRL2 POR2X1_772/a_16_28# POR2X1_772/CTRL POR2X1_772/a_76_344# POR2X1_772/a_56_344#
+ POR2X1
XPOR2X1_783 VDD GND POR2X1_783/B POR2X1_783/A POR2X1_783/Y POR2X1_783/m4_208_n4# POR2X1_783/O
+ POR2X1_783/CTRL2 POR2X1_783/a_16_28# POR2X1_783/CTRL POR2X1_783/a_76_344# POR2X1_783/a_56_344#
+ POR2X1
XPOR2X1_794 VDD GND POR2X1_794/B POR2X1_788/Y POR2X1_804/B POR2X1_794/m4_208_n4# POR2X1_794/O
+ POR2X1_794/CTRL2 POR2X1_794/a_16_28# POR2X1_794/CTRL POR2X1_794/a_76_344# POR2X1_794/a_56_344#
+ POR2X1
XPAND2X1_702 VDD GND POR2X1_135/Y POR2X1_45/Y PAND2X1_715/B PAND2X1_702/a_16_344#
+ PAND2X1_702/m4_208_n4# PAND2X1_702/O PAND2X1_702/a_56_28# PAND2X1_702/CTRL2 PAND2X1_702/CTRL
+ PAND2X1_702/a_76_28# PAND2X1
XPAND2X1_713 VDD GND PAND2X1_713/B PAND2X1_713/A PAND2X1_725/B PAND2X1_713/a_16_344#
+ PAND2X1_713/m4_208_n4# PAND2X1_713/O PAND2X1_713/a_56_28# PAND2X1_713/CTRL2 PAND2X1_713/CTRL
+ PAND2X1_713/a_76_28# PAND2X1
XPAND2X1_735 VDD GND PAND2X1_658/B PAND2X1_573/B PAND2X1_735/Y PAND2X1_735/a_16_344#
+ PAND2X1_735/m4_208_n4# PAND2X1_735/O PAND2X1_735/a_56_28# PAND2X1_735/CTRL2 PAND2X1_735/CTRL
+ PAND2X1_735/a_76_28# PAND2X1
XPAND2X1_724 VDD GND PAND2X1_724/B PAND2X1_714/Y PAND2X1_732/A PAND2X1_724/a_16_344#
+ PAND2X1_724/m4_208_n4# PAND2X1_724/O PAND2X1_724/a_56_28# PAND2X1_724/CTRL2 PAND2X1_724/CTRL
+ PAND2X1_724/a_76_28# PAND2X1
XPAND2X1_746 VDD GND POR2X1_260/A PAND2X1_73/Y POR2X1_781/A PAND2X1_746/a_16_344#
+ PAND2X1_746/m4_208_n4# PAND2X1_746/O PAND2X1_746/a_56_28# PAND2X1_746/CTRL2 PAND2X1_746/CTRL
+ PAND2X1_746/a_76_28# PAND2X1
XPAND2X1_768 VDD GND POR2X1_134/Y POR2X1_103/Y PAND2X1_768/Y PAND2X1_768/a_16_344#
+ PAND2X1_768/m4_208_n4# PAND2X1_768/O PAND2X1_768/a_56_28# PAND2X1_768/CTRL2 PAND2X1_768/CTRL
+ PAND2X1_768/a_76_28# PAND2X1
XPAND2X1_757 VDD GND POR2X1_756/Y PAND2X1_57/B POR2X1_791/A PAND2X1_757/a_16_344#
+ PAND2X1_757/m4_208_n4# PAND2X1_757/O PAND2X1_757/a_56_28# PAND2X1_757/CTRL2 PAND2X1_757/CTRL
+ PAND2X1_757/a_76_28# PAND2X1
XPAND2X1_779 VDD GND POR2X1_697/Y POR2X1_511/Y PAND2X1_779/Y PAND2X1_779/a_16_344#
+ PAND2X1_779/m4_208_n4# PAND2X1_779/O PAND2X1_779/a_56_28# PAND2X1_779/CTRL2 PAND2X1_779/CTRL
+ PAND2X1_779/a_76_28# PAND2X1
XPOR2X1_580 VDD GND POR2X1_578/Y POR2X1_579/Y D_GATE_579 POR2X1_580/m4_208_n4# POR2X1_580/O
+ POR2X1_580/CTRL2 POR2X1_580/a_16_28# POR2X1_580/CTRL POR2X1_580/a_76_344# POR2X1_580/a_56_344#
+ POR2X1
XPOR2X1_591 VDD GND POR2X1_65/A POR2X1_591/A POR2X1_591/Y POR2X1_591/m4_208_n4# POR2X1_591/O
+ POR2X1_591/CTRL2 POR2X1_591/a_16_28# POR2X1_591/CTRL POR2X1_591/a_76_344# POR2X1_591/a_56_344#
+ POR2X1
XPAND2X1_521 VDD GND POR2X1_68/A PAND2X1_20/A POR2X1_523/B PAND2X1_521/a_16_344# PAND2X1_521/m4_208_n4#
+ PAND2X1_521/O PAND2X1_521/a_56_28# PAND2X1_521/CTRL2 PAND2X1_521/CTRL PAND2X1_521/a_76_28#
+ PAND2X1
XPAND2X1_510 VDD GND PAND2X1_510/B PAND2X1_508/Y PAND2X1_657/B PAND2X1_510/a_16_344#
+ PAND2X1_510/m4_208_n4# PAND2X1_510/O PAND2X1_510/a_56_28# PAND2X1_510/CTRL2 PAND2X1_510/CTRL
+ PAND2X1_510/a_76_28# PAND2X1
XPAND2X1_554 VDD GND PAND2X1_140/A POR2X1_106/Y PAND2X1_563/B PAND2X1_554/a_16_344#
+ PAND2X1_554/m4_208_n4# PAND2X1_554/O PAND2X1_554/a_56_28# PAND2X1_554/CTRL2 PAND2X1_554/CTRL
+ PAND2X1_554/a_76_28# PAND2X1
XPAND2X1_543 VDD GND POR2X1_369/Y POR2X1_315/Y PAND2X1_552/B PAND2X1_543/a_16_344#
+ PAND2X1_543/m4_208_n4# PAND2X1_543/O PAND2X1_543/a_56_28# PAND2X1_543/CTRL2 PAND2X1_543/CTRL
+ PAND2X1_543/a_76_28# PAND2X1
XPAND2X1_565 VDD GND PAND2X1_550/Y PAND2X1_565/A PAND2X1_569/B PAND2X1_565/a_16_344#
+ PAND2X1_565/m4_208_n4# PAND2X1_565/O PAND2X1_565/a_56_28# PAND2X1_565/CTRL2 PAND2X1_565/CTRL
+ PAND2X1_565/a_76_28# PAND2X1
XPAND2X1_532 VDD GND POR2X1_394/A POR2X1_102/Y POR2X1_533/A PAND2X1_532/a_16_344#
+ PAND2X1_791/m4_208_n4# PAND2X1_532/O PAND2X1_532/a_56_28# PAND2X1_532/CTRL2 PAND2X1_532/CTRL
+ PAND2X1_532/a_76_28# PAND2X1
XPAND2X1_576 VDD GND PAND2X1_576/B PAND2X1_571/Y PAND2X1_579/B PAND2X1_576/a_16_344#
+ PAND2X1_576/m4_208_n4# PAND2X1_576/O PAND2X1_576/a_56_28# PAND2X1_576/CTRL2 PAND2X1_576/CTRL
+ PAND2X1_576/a_76_28# PAND2X1
XPAND2X1_598 VDD GND POR2X1_293/Y POR2X1_46/Y POR2X1_599/A PAND2X1_598/a_16_344# PAND2X1_598/m4_208_n4#
+ PAND2X1_598/O PAND2X1_598/a_56_28# PAND2X1_598/CTRL2 PAND2X1_598/CTRL PAND2X1_598/a_76_28#
+ PAND2X1
XPAND2X1_587 VDD GND PAND2X1_47/B D_INPUT_7 PAND2X1_587/Y PAND2X1_587/a_16_344# PAND2X1_587/m4_208_n4#
+ PAND2X1_587/O PAND2X1_587/a_56_28# PAND2X1_587/CTRL2 PAND2X1_587/CTRL PAND2X1_587/a_76_28#
+ PAND2X1
XPAND2X1_340 VDD GND PAND2X1_340/B POR2X1_88/Y PAND2X1_350/A PAND2X1_340/a_16_344#
+ PAND2X1_340/m4_208_n4# PAND2X1_340/O PAND2X1_340/a_56_28# PAND2X1_340/CTRL2 PAND2X1_340/CTRL
+ PAND2X1_340/a_76_28# PAND2X1
XPAND2X1_351 VDD GND PAND2X1_339/Y PAND2X1_351/A PAND2X1_351/Y PAND2X1_351/a_16_344#
+ PAND2X1_351/m4_208_n4# PAND2X1_351/O PAND2X1_351/a_56_28# PAND2X1_351/CTRL2 PAND2X1_351/CTRL
+ PAND2X1_351/a_76_28# PAND2X1
XPAND2X1_362 VDD GND PAND2X1_362/B PAND2X1_362/A PAND2X1_366/A PAND2X1_362/a_16_344#
+ PAND2X1_806/m4_208_n4# PAND2X1_362/O PAND2X1_362/a_56_28# PAND2X1_362/CTRL2 PAND2X1_362/CTRL
+ PAND2X1_362/a_76_28# PAND2X1
XPAND2X1_373 VDD GND POR2X1_78/A POR2X1_66/A POR2X1_544/B PAND2X1_373/a_16_344# PAND2X1_373/m4_208_n4#
+ PAND2X1_373/O PAND2X1_373/a_56_28# PAND2X1_373/CTRL2 PAND2X1_373/CTRL PAND2X1_373/a_76_28#
+ PAND2X1
XPAND2X1_384 VDD GND POR2X1_383/Y PAND2X1_41/B POR2X1_391/A PAND2X1_384/a_16_344#
+ PAND2X1_384/m4_208_n4# PAND2X1_384/O PAND2X1_384/a_56_28# PAND2X1_384/CTRL2 PAND2X1_384/CTRL
+ PAND2X1_384/a_76_28# PAND2X1
XPAND2X1_395 VDD GND POR2X1_814/B PAND2X1_60/B POR2X1_401/B PAND2X1_395/a_16_344#
+ PAND2X1_395/m4_208_n4# PAND2X1_395/O PAND2X1_395/a_56_28# PAND2X1_395/CTRL2 PAND2X1_395/CTRL
+ PAND2X1_395/a_76_28# PAND2X1
XPAND2X1_181 VDD GND POR2X1_179/Y POR2X1_178/Y PAND2X1_182/B PAND2X1_181/a_16_344#
+ PAND2X1_181/m4_208_n4# PAND2X1_181/O PAND2X1_181/a_56_28# PAND2X1_181/CTRL2 PAND2X1_181/CTRL
+ PAND2X1_181/a_76_28# PAND2X1
XPAND2X1_170 VDD GND PAND2X1_169/Y PAND2X1_168/Y PAND2X1_211/A PAND2X1_170/a_16_344#
+ PAND2X1_170/m4_208_n4# PAND2X1_170/O PAND2X1_170/a_56_28# PAND2X1_170/CTRL2 PAND2X1_170/CTRL
+ PAND2X1_170/a_76_28# PAND2X1
XPAND2X1_192 VDD GND PAND2X1_191/Y POR2X1_189/Y PAND2X1_192/Y PAND2X1_192/a_16_344#
+ PAND2X1_192/m4_208_n4# PAND2X1_192/O PAND2X1_192/a_56_28# PAND2X1_192/CTRL2 PAND2X1_192/CTRL
+ PAND2X1_192/a_76_28# PAND2X1
XPOR2X1_409 VDD GND POR2X1_409/B POR2X1_408/Y POR2X1_409/Y POR2X1_409/m4_208_n4# POR2X1_409/O
+ POR2X1_409/CTRL2 POR2X1_409/a_16_28# POR2X1_409/CTRL POR2X1_409/a_76_344# POR2X1_409/a_56_344#
+ POR2X1
XPOR2X1_206 VDD GND POR2X1_201/Y POR2X1_206/A POR2X1_215/A POR2X1_206/m4_208_n4# POR2X1_206/O
+ POR2X1_206/CTRL2 POR2X1_206/a_16_28# POR2X1_206/CTRL POR2X1_206/a_76_344# POR2X1_206/a_56_344#
+ POR2X1
XPOR2X1_228 VDD GND PAND2X1_7/Y PAND2X1_52/Y POR2X1_228/Y POR2X1_228/m4_208_n4# POR2X1_228/O
+ POR2X1_228/CTRL2 POR2X1_228/a_16_28# POR2X1_228/CTRL POR2X1_228/a_76_344# POR2X1_228/a_56_344#
+ POR2X1
XPOR2X1_217 VDD GND POR2X1_572/B POR2X1_141/Y POR2X1_218/A POR2X1_217/m4_208_n4# POR2X1_217/O
+ POR2X1_217/CTRL2 POR2X1_217/a_16_28# POR2X1_217/CTRL POR2X1_217/a_76_344# POR2X1_217/a_56_344#
+ POR2X1
XPOR2X1_239 VDD GND POR2X1_52/A POR2X1_102/Y POR2X1_239/Y POR2X1_239/m4_208_n4# POR2X1_239/O
+ POR2X1_239/CTRL2 POR2X1_239/a_16_28# POR2X1_239/CTRL POR2X1_239/a_76_344# POR2X1_239/a_56_344#
+ POR2X1
XPOR2X1_751 VDD GND POR2X1_7/B POR2X1_751/A POR2X1_751/Y POR2X1_751/m4_208_n4# POR2X1_751/O
+ POR2X1_751/CTRL2 POR2X1_751/a_16_28# POR2X1_751/CTRL POR2X1_751/a_76_344# POR2X1_751/a_56_344#
+ POR2X1
XPOR2X1_762 VDD GND D_INPUT_6 POR2X1_12/A POR2X1_763/A POR2X1_762/m4_208_n4# POR2X1_762/O
+ POR2X1_762/CTRL2 POR2X1_762/a_16_28# POR2X1_762/CTRL POR2X1_762/a_76_344# POR2X1_762/a_56_344#
+ POR2X1
XPOR2X1_740 VDD GND POR2X1_738/Y POR2X1_740/A POR2X1_740/Y POR2X1_740/m4_208_n4# POR2X1_740/O
+ POR2X1_740/CTRL2 POR2X1_740/a_16_28# POR2X1_740/CTRL POR2X1_740/a_76_344# POR2X1_740/a_56_344#
+ POR2X1
XPOR2X1_795 VDD GND POR2X1_795/B POR2X1_786/Y POR2X1_804/A POR2X1_795/m4_208_n4# POR2X1_795/O
+ POR2X1_795/CTRL2 POR2X1_795/a_16_28# POR2X1_795/CTRL POR2X1_795/a_76_344# POR2X1_795/a_56_344#
+ POR2X1
XPOR2X1_784 VDD GND POR2X1_777/Y POR2X1_784/A POR2X1_796/A POR2X1_784/m4_208_n4# POR2X1_784/O
+ POR2X1_784/CTRL2 POR2X1_784/a_16_28# POR2X1_784/CTRL POR2X1_784/a_76_344# POR2X1_784/a_56_344#
+ POR2X1
XPOR2X1_773 VDD GND POR2X1_773/B POR2X1_773/A POR2X1_774/A POR2X1_773/m4_208_n4# POR2X1_773/O
+ POR2X1_773/CTRL2 POR2X1_773/a_16_28# POR2X1_773/CTRL POR2X1_773/a_76_344# POR2X1_773/a_56_344#
+ POR2X1
XPAND2X1_703 VDD GND POR2X1_312/Y POR2X1_167/Y PAND2X1_714/A PAND2X1_703/a_16_344#
+ PAND2X1_317/m4_208_n4# PAND2X1_703/O PAND2X1_703/a_56_28# PAND2X1_703/CTRL2 PAND2X1_703/CTRL
+ PAND2X1_703/a_76_28# PAND2X1
XPAND2X1_736 VDD GND PAND2X1_735/Y PAND2X1_736/A PAND2X1_736/Y PAND2X1_736/a_16_344#
+ PAND2X1_736/m4_208_n4# PAND2X1_736/O PAND2X1_736/a_56_28# PAND2X1_736/CTRL2 PAND2X1_736/CTRL
+ PAND2X1_736/a_76_28# PAND2X1
XPAND2X1_714 VDD GND PAND2X1_714/B PAND2X1_714/A PAND2X1_714/Y PAND2X1_714/a_16_344#
+ PAND2X1_714/m4_208_n4# PAND2X1_714/O PAND2X1_714/a_56_28# PAND2X1_714/CTRL2 PAND2X1_714/CTRL
+ PAND2X1_714/a_76_28# PAND2X1
XPAND2X1_747 VDD GND POR2X1_68/A PAND2X1_48/B POR2X1_782/B PAND2X1_747/a_16_344# PAND2X1_747/m4_208_n4#
+ PAND2X1_747/O PAND2X1_747/a_56_28# PAND2X1_747/CTRL2 PAND2X1_747/CTRL PAND2X1_747/a_76_28#
+ PAND2X1
XPAND2X1_725 VDD GND PAND2X1_725/B PAND2X1_725/A PAND2X1_725/Y PAND2X1_725/a_16_344#
+ PAND2X1_725/m4_208_n4# PAND2X1_725/O PAND2X1_725/a_56_28# PAND2X1_725/CTRL2 PAND2X1_725/CTRL
+ PAND2X1_725/a_76_28# PAND2X1
XPAND2X1_769 VDD GND POR2X1_764/Y POR2X1_763/Y PAND2X1_769/Y PAND2X1_769/a_16_344#
+ PAND2X1_769/m4_208_n4# PAND2X1_769/O PAND2X1_769/a_56_28# PAND2X1_769/CTRL2 PAND2X1_769/CTRL
+ PAND2X1_769/a_76_28# PAND2X1
XPAND2X1_758 VDD GND POR2X1_96/A POR2X1_40/Y POR2X1_759/A PAND2X1_758/a_16_344# PAND2X1_758/m4_208_n4#
+ PAND2X1_758/O PAND2X1_758/a_56_28# PAND2X1_758/CTRL2 PAND2X1_758/CTRL PAND2X1_758/a_76_28#
+ PAND2X1
XPOR2X1_570 VDD GND POR2X1_570/B POR2X1_563/Y POR2X1_570/Y POR2X1_570/m4_208_n4# POR2X1_570/O
+ POR2X1_570/CTRL2 POR2X1_570/a_16_28# POR2X1_570/CTRL POR2X1_570/a_76_344# POR2X1_570/a_56_344#
+ POR2X1
XPOR2X1_581 VDD GND D_INPUT_6 POR2X1_3/A POR2X1_582/A POR2X1_581/m4_208_n4# POR2X1_581/O
+ POR2X1_581/CTRL2 POR2X1_581/a_16_28# POR2X1_581/CTRL POR2X1_581/a_76_344# POR2X1_581/a_56_344#
+ POR2X1
XPOR2X1_592 VDD GND POR2X1_832/B POR2X1_592/A POR2X1_592/Y POR2X1_592/m4_208_n4# POR2X1_592/O
+ POR2X1_592/CTRL2 POR2X1_592/a_16_28# POR2X1_592/CTRL POR2X1_592/a_76_344# POR2X1_592/a_56_344#
+ POR2X1
XPAND2X1_522 VDD GND POR2X1_590/A PAND2X1_58/A POR2X1_523/A PAND2X1_522/a_16_344#
+ PAND2X1_522/m4_208_n4# PAND2X1_522/O PAND2X1_522/a_56_28# PAND2X1_522/CTRL2 PAND2X1_522/CTRL
+ PAND2X1_522/a_76_28# PAND2X1
XPAND2X1_500 VDD GND PAND2X1_499/Y POR2X1_497/Y PAND2X1_501/B PAND2X1_500/a_16_344#
+ PAND2X1_84/m4_208_n4# PAND2X1_500/O PAND2X1_500/a_56_28# PAND2X1_500/CTRL2 PAND2X1_500/CTRL
+ PAND2X1_500/a_76_28# PAND2X1
XPAND2X1_511 VDD GND PAND2X1_48/A PAND2X1_32/B POR2X1_513/B PAND2X1_511/a_16_344#
+ POR2X1_807/m4_208_n4# PAND2X1_511/O PAND2X1_511/a_56_28# PAND2X1_511/CTRL2 PAND2X1_511/CTRL
+ PAND2X1_511/a_76_28# PAND2X1
XPAND2X1_555 VDD GND POR2X1_481/Y PAND2X1_555/A PAND2X1_555/Y PAND2X1_555/a_16_344#
+ PAND2X1_555/m4_208_n4# PAND2X1_555/O PAND2X1_555/a_56_28# PAND2X1_555/CTRL2 PAND2X1_555/CTRL
+ PAND2X1_555/a_76_28# PAND2X1
XPAND2X1_533 VDD GND POR2X1_532/Y PAND2X1_96/B POR2X1_788/B PAND2X1_533/a_16_344#
+ PAND2X1_533/m4_208_n4# PAND2X1_533/O PAND2X1_533/a_56_28# PAND2X1_533/CTRL2 PAND2X1_533/CTRL
+ PAND2X1_533/a_76_28# PAND2X1
XPAND2X1_544 VDD GND POR2X1_438/Y POR2X1_373/Y PAND2X1_551/A PAND2X1_544/a_16_344#
+ PAND2X1_544/m4_208_n4# PAND2X1_544/O PAND2X1_544/a_56_28# PAND2X1_544/CTRL2 PAND2X1_544/CTRL
+ PAND2X1_544/a_76_28# PAND2X1
XPAND2X1_577 VDD GND PAND2X1_577/B PAND2X1_569/Y PAND2X1_577/Y PAND2X1_577/a_16_344#
+ PAND2X1_577/m4_208_n4# PAND2X1_577/O PAND2X1_577/a_56_28# PAND2X1_577/CTRL2 PAND2X1_577/CTRL
+ PAND2X1_577/a_76_28# PAND2X1
XPAND2X1_566 VDD GND PAND2X1_303/Y PAND2X1_211/A PAND2X1_566/Y PAND2X1_566/a_16_344#
+ PAND2X1_566/m4_208_n4# PAND2X1_566/O PAND2X1_566/a_56_28# PAND2X1_566/CTRL2 PAND2X1_566/CTRL
+ PAND2X1_566/a_76_28# PAND2X1
XPAND2X1_588 VDD GND PAND2X1_587/Y POR2X1_502/A POR2X1_638/B PAND2X1_588/a_16_344#
+ PAND2X1_588/m4_208_n4# PAND2X1_588/O PAND2X1_588/a_56_28# PAND2X1_588/CTRL2 PAND2X1_588/CTRL
+ PAND2X1_588/a_76_28# PAND2X1
XPAND2X1_599 VDD GND POR2X1_828/A PAND2X1_69/A POR2X1_644/A PAND2X1_599/a_16_344#
+ POR2X1_598/m4_208_n4# PAND2X1_599/O PAND2X1_599/a_56_28# PAND2X1_599/CTRL2 PAND2X1_599/CTRL
+ PAND2X1_599/a_76_28# PAND2X1
XPAND2X1_330 VDD GND POR2X1_72/B POR2X1_52/A POR2X1_331/A PAND2X1_330/a_16_344# PAND2X1_330/m4_208_n4#
+ PAND2X1_330/O PAND2X1_330/a_56_28# PAND2X1_330/CTRL2 PAND2X1_330/CTRL PAND2X1_330/a_76_28#
+ PAND2X1
XPAND2X1_341 VDD GND PAND2X1_341/B PAND2X1_341/A PAND2X1_341/Y PAND2X1_341/a_16_344#
+ PAND2X1_341/m4_208_n4# PAND2X1_341/O PAND2X1_341/a_56_28# PAND2X1_341/CTRL2 PAND2X1_341/CTRL
+ PAND2X1_341/a_76_28# PAND2X1
XPAND2X1_363 VDD GND PAND2X1_360/Y PAND2X1_359/Y PAND2X1_363/Y PAND2X1_363/a_16_344#
+ PAND2X1_363/m4_208_n4# PAND2X1_363/O PAND2X1_363/a_56_28# PAND2X1_363/CTRL2 PAND2X1_363/CTRL
+ PAND2X1_363/a_76_28# PAND2X1
XPAND2X1_352 VDD GND PAND2X1_352/B PAND2X1_352/A PAND2X1_352/Y PAND2X1_352/a_16_344#
+ PAND2X1_352/m4_208_n4# PAND2X1_352/O PAND2X1_352/a_56_28# PAND2X1_352/CTRL2 PAND2X1_352/CTRL
+ PAND2X1_352/a_76_28# PAND2X1
XPAND2X1_385 VDD GND POR2X1_814/B POR2X1_66/A POR2X1_537/B PAND2X1_385/a_16_344# PAND2X1_385/m4_208_n4#
+ PAND2X1_385/O PAND2X1_385/a_56_28# PAND2X1_385/CTRL2 PAND2X1_385/CTRL PAND2X1_385/a_76_28#
+ PAND2X1
XPAND2X1_374 VDD GND POR2X1_373/Y POR2X1_322/Y PAND2X1_717/A PAND2X1_374/a_16_344#
+ PAND2X1_374/m4_208_n4# PAND2X1_374/O PAND2X1_374/a_56_28# PAND2X1_374/CTRL2 PAND2X1_374/CTRL
+ PAND2X1_374/a_76_28# PAND2X1
XPAND2X1_396 VDD GND PAND2X1_69/A PAND2X1_23/Y POR2X1_401/A PAND2X1_396/a_16_344#
+ PAND2X1_396/m4_208_n4# PAND2X1_396/O PAND2X1_396/a_56_28# PAND2X1_396/CTRL2 PAND2X1_396/CTRL
+ PAND2X1_396/a_76_28# PAND2X1
XPAND2X1_160 VDD GND POR2X1_394/A POR2X1_23/Y PAND2X1_162/A PAND2X1_160/a_16_344#
+ PAND2X1_160/m4_208_n4# PAND2X1_160/O PAND2X1_160/a_56_28# PAND2X1_160/CTRL2 PAND2X1_160/CTRL
+ PAND2X1_160/a_76_28# PAND2X1
XPAND2X1_171 VDD GND PAND2X1_41/B PAND2X1_23/Y POR2X1_174/B PAND2X1_171/a_16_344#
+ POR2X1_567/m4_208_n4# PAND2X1_171/O PAND2X1_171/a_56_28# PAND2X1_171/CTRL2 PAND2X1_171/CTRL
+ PAND2X1_171/a_76_28# PAND2X1
XPAND2X1_193 VDD GND POR2X1_13/Y POR2X1_7/Y PAND2X1_193/Y PAND2X1_193/a_16_344# PAND2X1_193/m4_208_n4#
+ PAND2X1_193/O PAND2X1_193/a_56_28# PAND2X1_193/CTRL2 PAND2X1_193/CTRL PAND2X1_193/a_76_28#
+ PAND2X1
XPAND2X1_182 VDD GND PAND2X1_182/B PAND2X1_182/A PAND2X1_352/A PAND2X1_182/a_16_344#
+ PAND2X1_182/m4_208_n4# PAND2X1_182/O PAND2X1_182/a_56_28# PAND2X1_182/CTRL2 PAND2X1_182/CTRL
+ PAND2X1_182/a_76_28# PAND2X1
XPOR2X1_207 VDD GND POR2X1_207/B POR2X1_207/A POR2X1_214/B POR2X1_207/m4_208_n4# POR2X1_207/O
+ POR2X1_207/CTRL2 POR2X1_207/a_16_28# POR2X1_207/CTRL POR2X1_207/a_76_344# POR2X1_207/a_56_344#
+ POR2X1
XPOR2X1_229 VDD GND POR2X1_13/A POR2X1_23/Y POR2X1_229/Y POR2X1_229/m4_208_n4# POR2X1_229/O
+ POR2X1_229/CTRL2 POR2X1_229/a_16_28# POR2X1_229/CTRL POR2X1_229/a_76_344# POR2X1_229/a_56_344#
+ POR2X1
XPOR2X1_218 VDD GND POR2X1_216/Y POR2X1_218/A POR2X1_218/Y POR2X1_218/m4_208_n4# POR2X1_218/O
+ POR2X1_218/CTRL2 POR2X1_218/a_16_28# POR2X1_218/CTRL POR2X1_218/a_76_344# POR2X1_218/a_56_344#
+ POR2X1
XPOR2X1_763 VDD GND POR2X1_46/Y POR2X1_763/A POR2X1_763/Y POR2X1_763/m4_208_n4# POR2X1_763/O
+ POR2X1_763/CTRL2 POR2X1_763/a_16_28# POR2X1_763/CTRL POR2X1_763/a_76_344# POR2X1_763/a_56_344#
+ POR2X1
XPOR2X1_730 VDD GND POR2X1_730/B POR2X1_729/Y POR2X1_730/Y POR2X1_730/m4_208_n4# POR2X1_730/O
+ POR2X1_730/CTRL2 POR2X1_730/a_16_28# POR2X1_730/CTRL POR2X1_730/a_76_344# POR2X1_730/a_56_344#
+ POR2X1
XPOR2X1_752 VDD GND D_INPUT_5 POR2X1_51/A POR2X1_752/Y POR2X1_752/m4_208_n4# POR2X1_752/O
+ POR2X1_752/CTRL2 POR2X1_752/a_16_28# POR2X1_752/CTRL POR2X1_752/a_76_344# POR2X1_752/a_56_344#
+ POR2X1
XPOR2X1_741 VDD GND POR2X1_741/B POR2X1_741/A POR2X1_741/Y POR2X1_741/m4_208_n4# POR2X1_741/O
+ POR2X1_741/CTRL2 POR2X1_741/a_16_28# POR2X1_741/CTRL POR2X1_741/a_76_344# POR2X1_741/a_56_344#
+ POR2X1
XPOR2X1_785 VDD GND POR2X1_785/B POR2X1_785/A POR2X1_795/B POR2X1_785/m4_208_n4# POR2X1_785/O
+ POR2X1_785/CTRL2 POR2X1_785/a_16_28# POR2X1_785/CTRL POR2X1_785/a_76_344# POR2X1_785/a_56_344#
+ POR2X1
XPOR2X1_796 VDD GND POR2X1_783/Y POR2X1_796/A POR2X1_796/Y POR2X1_796/m4_208_n4# POR2X1_796/O
+ POR2X1_796/CTRL2 POR2X1_796/a_16_28# POR2X1_796/CTRL POR2X1_796/a_76_344# POR2X1_796/a_56_344#
+ POR2X1
XPOR2X1_774 VDD GND POR2X1_774/B POR2X1_774/A POR2X1_774/Y POR2X1_774/m4_208_n4# POR2X1_774/O
+ POR2X1_774/CTRL2 POR2X1_774/a_16_28# POR2X1_774/CTRL POR2X1_774/a_76_344# POR2X1_774/a_56_344#
+ POR2X1
XPAND2X1_704 VDD GND POR2X1_417/Y POR2X1_313/Y PAND2X1_714/B PAND2X1_704/a_16_344#
+ PAND2X1_704/m4_208_n4# PAND2X1_704/O PAND2X1_704/a_56_28# PAND2X1_704/CTRL2 PAND2X1_704/CTRL
+ PAND2X1_704/a_76_28# PAND2X1
XPAND2X1_737 VDD GND PAND2X1_737/B PAND2X1_733/Y PAND2X1_741/B PAND2X1_737/a_16_344#
+ PAND2X1_737/m4_208_n4# PAND2X1_737/O PAND2X1_737/a_56_28# PAND2X1_737/CTRL2 PAND2X1_737/CTRL
+ PAND2X1_737/a_76_28# PAND2X1
XPAND2X1_715 VDD GND PAND2X1_715/B PAND2X1_115/B PAND2X1_724/B PAND2X1_715/a_16_344#
+ PAND2X1_715/m4_208_n4# PAND2X1_715/O PAND2X1_715/a_56_28# PAND2X1_715/CTRL2 PAND2X1_715/CTRL
+ PAND2X1_715/a_76_28# PAND2X1
XPAND2X1_726 VDD GND PAND2X1_726/B POR2X1_152/Y PAND2X1_731/A PAND2X1_726/a_16_344#
+ PAND2X1_726/m4_208_n4# PAND2X1_726/O PAND2X1_726/a_56_28# PAND2X1_726/CTRL2 PAND2X1_726/CTRL
+ PAND2X1_726/a_76_28# PAND2X1
XPAND2X1_748 VDD GND POR2X1_709/A PAND2X1_6/A POR2X1_789/B PAND2X1_748/a_16_344# PAND2X1_748/m4_208_n4#
+ PAND2X1_748/O PAND2X1_748/a_56_28# PAND2X1_748/CTRL2 PAND2X1_748/CTRL PAND2X1_748/a_76_28#
+ PAND2X1
XPAND2X1_759 VDD GND POR2X1_758/Y POR2X1_383/A POR2X1_792/B PAND2X1_759/a_16_344#
+ PAND2X1_759/m4_208_n4# PAND2X1_759/O PAND2X1_759/a_56_28# PAND2X1_759/CTRL2 PAND2X1_759/CTRL
+ PAND2X1_759/a_76_28# PAND2X1
XPOR2X1_1 VDD GND INPUT_6 D_INPUT_7 POR2X1_3/B POR2X1_1/m4_208_n4# POR2X1_1/O POR2X1_1/CTRL2
+ POR2X1_1/a_16_28# POR2X1_1/CTRL POR2X1_1/a_76_344# POR2X1_1/a_56_344# POR2X1
XPOR2X1_571 VDD GND POR2X1_560/Y POR2X1_561/Y POR2X1_571/Y POR2X1_571/m4_208_n4# POR2X1_571/O
+ POR2X1_571/CTRL2 POR2X1_571/a_16_28# POR2X1_571/CTRL POR2X1_571/a_76_344# POR2X1_571/a_56_344#
+ POR2X1
XPOR2X1_560 VDD GND POR2X1_523/Y POR2X1_559/Y POR2X1_560/Y POR2X1_560/m4_208_n4# POR2X1_560/O
+ POR2X1_560/CTRL2 POR2X1_560/a_16_28# POR2X1_560/CTRL POR2X1_560/a_76_344# POR2X1_560/a_56_344#
+ POR2X1
XPOR2X1_582 VDD GND POR2X1_257/A POR2X1_582/A POR2X1_582/Y POR2X1_582/m4_208_n4# POR2X1_582/O
+ POR2X1_582/CTRL2 POR2X1_582/a_16_28# POR2X1_582/CTRL POR2X1_582/a_76_344# POR2X1_582/a_56_344#
+ POR2X1
XPOR2X1_593 VDD GND POR2X1_593/B POR2X1_592/Y POR2X1_652/A POR2X1_593/m4_208_n4# POR2X1_593/O
+ POR2X1_593/CTRL2 POR2X1_593/a_16_28# POR2X1_593/CTRL POR2X1_593/a_76_344# POR2X1_593/a_56_344#
+ POR2X1
XPAND2X1_501 VDD GND PAND2X1_501/B POR2X1_498/Y PAND2X1_573/B PAND2X1_501/a_16_344#
+ PAND2X1_501/m4_208_n4# PAND2X1_501/O PAND2X1_501/a_56_28# PAND2X1_501/CTRL2 PAND2X1_501/CTRL
+ PAND2X1_501/a_76_28# PAND2X1
XPAND2X1_512 VDD GND POR2X1_306/Y INPUT_0 PAND2X1_512/Y PAND2X1_512/a_16_344# PAND2X1_512/m4_208_n4#
+ PAND2X1_512/O PAND2X1_512/a_56_28# PAND2X1_512/CTRL2 PAND2X1_512/CTRL PAND2X1_512/a_76_28#
+ PAND2X1
XPAND2X1_523 VDD GND POR2X1_522/Y POR2X1_521/Y PAND2X1_844/B PAND2X1_523/a_16_344#
+ PAND2X1_523/m4_208_n4# PAND2X1_523/O PAND2X1_523/a_56_28# PAND2X1_523/CTRL2 PAND2X1_523/CTRL
+ PAND2X1_523/a_76_28# PAND2X1
XPAND2X1_534 VDD GND PAND2X1_60/B POR2X1_296/B POR2X1_535/A PAND2X1_534/a_16_344#
+ PAND2X1_534/m4_208_n4# PAND2X1_534/O PAND2X1_534/a_56_28# PAND2X1_534/CTRL2 PAND2X1_534/CTRL
+ PAND2X1_534/a_76_28# PAND2X1
XPAND2X1_545 VDD GND POR2X1_524/Y POR2X1_441/Y PAND2X1_545/Y PAND2X1_545/a_16_344#
+ PAND2X1_545/m4_208_n4# PAND2X1_545/O PAND2X1_545/a_56_28# PAND2X1_545/CTRL2 PAND2X1_545/CTRL
+ PAND2X1_545/a_76_28# PAND2X1
XPAND2X1_567 VDD GND PAND2X1_539/Y PAND2X1_535/Y PAND2X1_568/B PAND2X1_567/a_16_344#
+ PAND2X1_567/m4_208_n4# PAND2X1_567/O PAND2X1_567/a_56_28# PAND2X1_567/CTRL2 PAND2X1_567/CTRL
+ PAND2X1_567/a_76_28# PAND2X1
XPAND2X1_578 VDD GND PAND2X1_577/Y PAND2X1_578/A PAND2X1_578/Y PAND2X1_578/a_16_344#
+ PAND2X1_287/m4_208_n4# PAND2X1_578/O PAND2X1_578/a_56_28# PAND2X1_578/CTRL2 PAND2X1_578/CTRL
+ PAND2X1_578/a_76_28# PAND2X1
XPAND2X1_556 VDD GND PAND2X1_556/B PAND2X1_631/A PAND2X1_562/B PAND2X1_556/a_16_344#
+ POR2X1_183/m4_208_n4# PAND2X1_556/O PAND2X1_556/a_56_28# PAND2X1_556/CTRL2 PAND2X1_556/CTRL
+ PAND2X1_556/a_76_28# PAND2X1
XPAND2X1_589 VDD GND POR2X1_130/A PAND2X1_58/A POR2X1_592/A PAND2X1_589/a_16_344#
+ PAND2X1_589/m4_208_n4# PAND2X1_589/O PAND2X1_589/a_56_28# PAND2X1_589/CTRL2 PAND2X1_589/CTRL
+ PAND2X1_589/a_76_28# PAND2X1
XPOR2X1_390 VDD GND POR2X1_390/B POR2X1_389/Y POR2X1_392/B POR2X1_390/m4_208_n4# POR2X1_390/O
+ POR2X1_390/CTRL2 POR2X1_390/a_16_28# POR2X1_390/CTRL POR2X1_390/a_76_344# POR2X1_390/a_56_344#
+ POR2X1
XPAND2X1_320 VDD GND PAND2X1_90/Y PAND2X1_69/A POR2X1_324/B PAND2X1_320/a_16_344#
+ PAND2X1_320/m4_208_n4# PAND2X1_320/O PAND2X1_320/a_56_28# PAND2X1_320/CTRL2 PAND2X1_320/CTRL
+ PAND2X1_320/a_76_28# PAND2X1
XPAND2X1_364 VDD GND PAND2X1_364/B PAND2X1_357/Y PAND2X1_365/B PAND2X1_364/a_16_344#
+ PAND2X1_364/m4_208_n4# PAND2X1_364/O PAND2X1_364/a_56_28# PAND2X1_364/CTRL2 PAND2X1_364/CTRL
+ PAND2X1_364/a_76_28# PAND2X1
XPAND2X1_342 VDD GND POR2X1_248/Y POR2X1_246/Y PAND2X1_349/A PAND2X1_342/a_16_344#
+ PAND2X1_342/m4_208_n4# PAND2X1_342/O PAND2X1_342/a_56_28# PAND2X1_342/CTRL2 PAND2X1_342/CTRL
+ PAND2X1_342/a_76_28# PAND2X1
XPAND2X1_353 VDD GND PAND2X1_308/Y PAND2X1_303/Y PAND2X1_353/Y PAND2X1_353/a_16_344#
+ PAND2X1_353/m4_208_n4# PAND2X1_353/O PAND2X1_353/a_56_28# PAND2X1_353/CTRL2 PAND2X1_353/CTRL
+ PAND2X1_353/a_76_28# PAND2X1
XPAND2X1_331 VDD GND POR2X1_330/Y POR2X1_186/Y POR2X1_355/A PAND2X1_331/a_16_344#
+ PAND2X1_331/m4_208_n4# PAND2X1_331/O PAND2X1_331/a_56_28# PAND2X1_331/CTRL2 PAND2X1_331/CTRL
+ PAND2X1_331/a_76_28# PAND2X1
XPAND2X1_386 VDD GND PAND2X1_18/B D_INPUT_4 PAND2X1_386/Y PAND2X1_386/a_16_344# PAND2X1_386/m4_208_n4#
+ PAND2X1_386/O PAND2X1_386/a_56_28# PAND2X1_386/CTRL2 PAND2X1_386/CTRL PAND2X1_386/a_76_28#
+ PAND2X1
XPAND2X1_375 VDD GND POR2X1_416/B POR2X1_32/A POR2X1_376/A PAND2X1_375/a_16_344# PAND2X1_375/m4_208_n4#
+ PAND2X1_375/O PAND2X1_375/a_56_28# PAND2X1_375/CTRL2 PAND2X1_375/CTRL PAND2X1_375/a_76_28#
+ PAND2X1
XPAND2X1_397 VDD GND PAND2X1_82/Y POR2X1_66/B POR2X1_402/B PAND2X1_397/a_16_344# POR2X1_398/m4_208_n4#
+ PAND2X1_397/O PAND2X1_397/a_56_28# PAND2X1_397/CTRL2 PAND2X1_397/CTRL PAND2X1_397/a_76_28#
+ PAND2X1
XPAND2X1_150 VDD GND PAND2X1_63/B PAND2X1_90/A POR2X1_186/B PAND2X1_150/a_16_344#
+ PAND2X1_150/m4_208_n4# PAND2X1_150/O PAND2X1_150/a_56_28# PAND2X1_150/CTRL2 PAND2X1_150/CTRL
+ PAND2X1_150/a_76_28# PAND2X1
XPAND2X1_172 VDD GND POR2X1_590/A PAND2X1_72/A POR2X1_174/A PAND2X1_172/a_16_344#
+ PAND2X1_172/m4_208_n4# PAND2X1_172/O PAND2X1_172/a_56_28# PAND2X1_172/CTRL2 PAND2X1_172/CTRL
+ PAND2X1_172/a_76_28# PAND2X1
XPAND2X1_161 VDD GND POR2X1_669/B POR2X1_257/A PAND2X1_161/Y PAND2X1_161/a_16_344#
+ PAND2X1_161/m4_208_n4# PAND2X1_161/O PAND2X1_161/a_56_28# PAND2X1_161/CTRL2 PAND2X1_161/CTRL
+ PAND2X1_161/a_76_28# PAND2X1
XPAND2X1_183 VDD GND PAND2X1_41/B PAND2X1_6/Y POR2X1_540/A PAND2X1_183/a_16_344# PAND2X1_183/m4_208_n4#
+ PAND2X1_183/O PAND2X1_183/a_56_28# PAND2X1_183/CTRL2 PAND2X1_183/CTRL PAND2X1_183/a_76_28#
+ PAND2X1
XPAND2X1_194 VDD GND POR2X1_39/Y POR2X1_16/Y PAND2X1_200/B PAND2X1_194/a_16_344# PAND2X1_194/m4_208_n4#
+ PAND2X1_194/O PAND2X1_194/a_56_28# PAND2X1_194/CTRL2 PAND2X1_194/CTRL PAND2X1_194/a_76_28#
+ PAND2X1
XPOR2X1_208 VDD GND POR2X1_35/Y POR2X1_208/A POR2X1_208/Y POR2X1_208/m4_208_n4# POR2X1_208/O
+ POR2X1_208/CTRL2 POR2X1_208/a_16_28# POR2X1_208/CTRL POR2X1_208/a_76_344# POR2X1_208/a_56_344#
+ POR2X1
XPOR2X1_219 VDD GND POR2X1_219/B POR2X1_215/Y POR2X1_222/A POR2X1_219/m4_208_n4# POR2X1_219/O
+ POR2X1_219/CTRL2 POR2X1_219/a_16_28# POR2X1_219/CTRL POR2X1_219/a_76_344# POR2X1_219/a_56_344#
+ POR2X1
XPOR2X1_720 VDD GND POR2X1_720/B POR2X1_720/A POR2X1_720/Y POR2X1_720/m4_208_n4# POR2X1_720/O
+ POR2X1_720/CTRL2 POR2X1_720/a_16_28# POR2X1_720/CTRL POR2X1_720/a_76_344# POR2X1_720/a_56_344#
+ POR2X1
XPOR2X1_742 VDD GND POR2X1_740/Y POR2X1_741/Y D_GATE_741 POR2X1_742/m4_208_n4# POR2X1_742/O
+ POR2X1_742/CTRL2 POR2X1_742/a_16_28# POR2X1_742/CTRL POR2X1_742/a_76_344# POR2X1_742/a_56_344#
+ POR2X1
XPOR2X1_731 VDD GND POR2X1_726/Y POR2X1_731/A POR2X1_731/Y POR2X1_731/m4_208_n4# POR2X1_731/O
+ POR2X1_731/CTRL2 POR2X1_731/a_16_28# POR2X1_731/CTRL POR2X1_731/a_76_344# POR2X1_731/a_56_344#
+ POR2X1
XPOR2X1_753 VDD GND POR2X1_816/A POR2X1_752/Y POR2X1_753/Y POR2X1_753/m4_208_n4# POR2X1_753/O
+ POR2X1_753/CTRL2 POR2X1_753/a_16_28# POR2X1_753/CTRL POR2X1_753/a_76_344# POR2X1_753/a_56_344#
+ POR2X1
XPOR2X1_786 VDD GND POR2X1_84/Y POR2X1_786/A POR2X1_786/Y POR2X1_786/m4_208_n4# POR2X1_786/O
+ POR2X1_786/CTRL2 POR2X1_786/a_16_28# POR2X1_786/CTRL POR2X1_786/a_76_344# POR2X1_786/a_56_344#
+ POR2X1
XPOR2X1_775 VDD GND POR2X1_97/A POR2X1_775/A POR2X1_785/B POR2X1_785/m4_208_n4# POR2X1_775/O
+ POR2X1_775/CTRL2 POR2X1_775/a_16_28# POR2X1_775/CTRL POR2X1_775/a_76_344# POR2X1_775/a_56_344#
+ POR2X1
XPOR2X1_764 VDD GND POR2X1_40/Y POR2X1_394/A POR2X1_764/Y POR2X1_764/m4_208_n4# POR2X1_764/O
+ POR2X1_764/CTRL2 POR2X1_764/a_16_28# POR2X1_764/CTRL POR2X1_764/a_76_344# POR2X1_764/a_56_344#
+ POR2X1
XPOR2X1_797 VDD GND POR2X1_149/Y POR2X1_797/A POR2X1_803/A POR2X1_797/m4_208_n4# POR2X1_797/O
+ POR2X1_797/CTRL2 POR2X1_797/a_16_28# POR2X1_797/CTRL POR2X1_797/a_76_344# POR2X1_797/a_56_344#
+ POR2X1
XPAND2X1_716 VDD GND PAND2X1_716/B PAND2X1_341/A PAND2X1_723/A PAND2X1_716/a_16_344#
+ PAND2X1_716/m4_208_n4# PAND2X1_716/O PAND2X1_716/a_56_28# PAND2X1_716/CTRL2 PAND2X1_716/CTRL
+ PAND2X1_716/a_76_28# PAND2X1
XPAND2X1_727 VDD GND PAND2X1_444/Y PAND2X1_308/Y PAND2X1_731/B PAND2X1_727/a_16_344#
+ PAND2X1_727/m4_208_n4# PAND2X1_727/O PAND2X1_727/a_56_28# PAND2X1_727/CTRL2 PAND2X1_727/CTRL
+ PAND2X1_727/a_76_28# PAND2X1
XPAND2X1_738 VDD GND PAND2X1_738/B PAND2X1_738/A PAND2X1_738/Y PAND2X1_738/a_16_344#
+ PAND2X1_738/m4_208_n4# PAND2X1_738/O PAND2X1_738/a_56_28# PAND2X1_738/CTRL2 PAND2X1_738/CTRL
+ PAND2X1_738/a_76_28# PAND2X1
XPAND2X1_705 VDD GND POR2X1_526/Y POR2X1_485/Y PAND2X1_713/A PAND2X1_705/a_16_344#
+ PAND2X1_705/m4_208_n4# PAND2X1_705/O PAND2X1_705/a_56_28# PAND2X1_705/CTRL2 PAND2X1_705/CTRL
+ PAND2X1_705/a_76_28# PAND2X1
XPAND2X1_749 VDD GND PAND2X1_8/Y D_INPUT_0 POR2X1_750/A PAND2X1_749/a_16_344# PAND2X1_749/m4_208_n4#
+ PAND2X1_749/O PAND2X1_749/a_56_28# PAND2X1_749/CTRL2 PAND2X1_749/CTRL PAND2X1_749/a_76_28#
+ PAND2X1
XPOR2X1_2 VDD GND INPUT_4 INPUT_5 POR2X1_3/A POR2X1_2/m4_208_n4# POR2X1_2/O POR2X1_2/CTRL2
+ POR2X1_2/a_16_28# POR2X1_2/CTRL POR2X1_2/a_76_344# POR2X1_2/a_56_344# POR2X1
XPOR2X1_550 VDD GND POR2X1_550/B POR2X1_550/A POR2X1_550/Y POR2X1_550/m4_208_n4# POR2X1_550/O
+ POR2X1_550/CTRL2 POR2X1_550/a_16_28# POR2X1_550/CTRL POR2X1_550/a_76_344# POR2X1_550/a_56_344#
+ POR2X1
XPOR2X1_561 VDD GND POR2X1_561/B POR2X1_558/Y POR2X1_561/Y POR2X1_561/m4_208_n4# POR2X1_561/O
+ POR2X1_561/CTRL2 POR2X1_561/a_16_28# POR2X1_561/CTRL POR2X1_561/a_76_344# POR2X1_561/a_56_344#
+ POR2X1
XPOR2X1_594 VDD GND POR2X1_96/A POR2X1_594/A POR2X1_594/Y POR2X1_594/m4_208_n4# POR2X1_594/O
+ POR2X1_594/CTRL2 POR2X1_594/a_16_28# POR2X1_594/CTRL POR2X1_594/a_76_344# POR2X1_594/a_56_344#
+ POR2X1
XPOR2X1_572 VDD GND POR2X1_572/B POR2X1_267/Y POR2X1_572/Y POR2X1_572/m4_208_n4# POR2X1_572/O
+ POR2X1_572/CTRL2 POR2X1_572/a_16_28# POR2X1_572/CTRL POR2X1_572/a_76_344# POR2X1_572/a_56_344#
+ POR2X1
XPOR2X1_583 VDD GND POR2X1_32/A POR2X1_49/Y POR2X1_583/Y POR2X1_583/m4_208_n4# POR2X1_583/O
+ POR2X1_583/CTRL2 POR2X1_583/a_16_28# POR2X1_583/CTRL POR2X1_583/a_76_344# POR2X1_583/a_56_344#
+ POR2X1
XPAND2X1_502 VDD GND POR2X1_376/B POR2X1_77/Y POR2X1_503/A PAND2X1_502/a_16_344# PAND2X1_502/m4_208_n4#
+ PAND2X1_502/O PAND2X1_502/a_56_28# PAND2X1_502/CTRL2 PAND2X1_502/CTRL PAND2X1_502/a_76_28#
+ PAND2X1
XPAND2X1_513 VDD GND PAND2X1_512/Y POR2X1_511/Y POR2X1_516/B PAND2X1_513/a_16_344#
+ PAND2X1_513/m4_208_n4# PAND2X1_513/O PAND2X1_513/a_56_28# PAND2X1_513/CTRL2 PAND2X1_513/CTRL
+ PAND2X1_513/a_76_28# PAND2X1
XPAND2X1_524 VDD GND POR2X1_614/A PAND2X1_48/B POR2X1_545/A PAND2X1_524/a_16_344#
+ PAND2X1_524/m4_208_n4# PAND2X1_524/O PAND2X1_524/a_56_28# PAND2X1_524/CTRL2 PAND2X1_524/CTRL
+ PAND2X1_524/a_76_28# PAND2X1
XPAND2X1_546 VDD GND POR2X1_526/Y POR2X1_525/Y PAND2X1_546/Y PAND2X1_546/a_16_344#
+ PAND2X1_546/m4_208_n4# PAND2X1_546/O PAND2X1_546/a_56_28# PAND2X1_546/CTRL2 PAND2X1_546/CTRL
+ PAND2X1_546/a_76_28# PAND2X1
XPAND2X1_535 VDD GND POR2X1_534/Y POR2X1_533/Y PAND2X1_535/Y PAND2X1_535/a_16_344#
+ PAND2X1_855/m4_208_n4# PAND2X1_535/O PAND2X1_535/a_56_28# PAND2X1_535/CTRL2 PAND2X1_535/CTRL
+ PAND2X1_535/a_76_28# PAND2X1
XPAND2X1_557 VDD GND POR2X1_490/Y PAND2X1_557/A PAND2X1_561/A PAND2X1_557/a_16_344#
+ PAND2X1_473/m4_208_n4# PAND2X1_557/O PAND2X1_557/a_56_28# PAND2X1_557/CTRL2 PAND2X1_557/CTRL
+ PAND2X1_557/a_76_28# PAND2X1
XPAND2X1_579 VDD GND PAND2X1_579/B PAND2X1_579/A PAND2X1_580/B PAND2X1_579/a_16_344#
+ PAND2X1_579/m4_208_n4# PAND2X1_579/O PAND2X1_579/a_56_28# PAND2X1_579/CTRL2 PAND2X1_579/CTRL
+ PAND2X1_579/a_76_28# PAND2X1
XPAND2X1_568 VDD GND PAND2X1_568/B PAND2X1_566/Y PAND2X1_578/A PAND2X1_568/a_16_344#
+ PAND2X1_347/m4_208_n4# PAND2X1_568/O PAND2X1_568/a_56_28# PAND2X1_568/CTRL2 PAND2X1_568/CTRL
+ PAND2X1_568/a_76_28# PAND2X1
XPOR2X1_380 VDD GND POR2X1_394/A POR2X1_380/A POR2X1_380/Y POR2X1_380/m4_208_n4# POR2X1_380/O
+ POR2X1_380/CTRL2 POR2X1_380/a_16_28# POR2X1_380/CTRL POR2X1_380/a_76_344# POR2X1_380/a_56_344#
+ POR2X1
XPOR2X1_391 VDD GND POR2X1_391/B POR2X1_391/A POR2X1_391/Y POR2X1_391/m4_208_n4# POR2X1_391/O
+ POR2X1_391/CTRL2 POR2X1_391/a_16_28# POR2X1_391/CTRL POR2X1_391/a_76_344# POR2X1_391/a_56_344#
+ POR2X1
XPAND2X1_310 VDD GND PAND2X1_41/B POR2X1_68/B POR2X1_335/A PAND2X1_310/a_16_344# PAND2X1_310/m4_208_n4#
+ PAND2X1_310/O PAND2X1_310/a_56_28# PAND2X1_310/CTRL2 PAND2X1_310/CTRL PAND2X1_310/a_76_28#
+ PAND2X1
XPAND2X1_321 VDD GND PAND2X1_65/B POR2X1_294/B POR2X1_324/A PAND2X1_321/a_16_344#
+ PAND2X1_321/m4_208_n4# PAND2X1_321/O PAND2X1_321/a_56_28# PAND2X1_321/CTRL2 PAND2X1_321/CTRL
+ PAND2X1_321/a_76_28# PAND2X1
XPAND2X1_354 VDD GND PAND2X1_854/A PAND2X1_354/A PAND2X1_354/Y PAND2X1_354/a_16_344#
+ PAND2X1_354/m4_208_n4# PAND2X1_354/O PAND2X1_354/a_56_28# PAND2X1_354/CTRL2 PAND2X1_354/CTRL
+ PAND2X1_354/a_76_28# PAND2X1
XPAND2X1_343 VDD GND POR2X1_251/Y POR2X1_250/Y PAND2X1_349/B PAND2X1_343/a_16_344#
+ PAND2X1_343/m4_208_n4# PAND2X1_343/O PAND2X1_343/a_56_28# PAND2X1_343/CTRL2 PAND2X1_343/CTRL
+ PAND2X1_343/a_76_28# PAND2X1
XPAND2X1_332 VDD GND POR2X1_135/Y POR2X1_111/Y PAND2X1_332/Y PAND2X1_332/a_16_344#
+ PAND2X1_332/m4_208_n4# PAND2X1_332/O PAND2X1_332/a_56_28# PAND2X1_332/CTRL2 PAND2X1_332/CTRL
+ PAND2X1_332/a_76_28# PAND2X1
XPAND2X1_365 VDD GND PAND2X1_365/B PAND2X1_365/A PAND2X1_367/A PAND2X1_365/a_16_344#
+ PAND2X1_365/m4_208_n4# PAND2X1_365/O PAND2X1_365/a_56_28# PAND2X1_365/CTRL2 PAND2X1_365/CTRL
+ PAND2X1_365/a_76_28# PAND2X1
XPAND2X1_376 VDD GND POR2X1_375/Y POR2X1_502/A POR2X1_459/B PAND2X1_376/a_16_344#
+ PAND2X1_376/m4_208_n4# PAND2X1_376/O PAND2X1_376/a_56_28# PAND2X1_376/CTRL2 PAND2X1_376/CTRL
+ PAND2X1_376/a_76_28# PAND2X1
XPAND2X1_387 VDD GND PAND2X1_386/Y PAND2X1_93/B POR2X1_389/A PAND2X1_387/a_16_344#
+ PAND2X1_387/m4_208_n4# PAND2X1_387/O PAND2X1_387/a_56_28# PAND2X1_387/CTRL2 PAND2X1_387/CTRL
+ PAND2X1_387/a_76_28# PAND2X1
XPAND2X1_398 VDD GND POR2X1_293/Y POR2X1_16/A POR2X1_399/A PAND2X1_398/a_16_344# PAND2X1_398/m4_208_n4#
+ PAND2X1_398/O PAND2X1_398/a_56_28# PAND2X1_398/CTRL2 PAND2X1_398/CTRL PAND2X1_398/a_76_28#
+ PAND2X1
XPAND2X1_140 VDD GND POR2X1_131/Y PAND2X1_140/A PAND2X1_140/Y PAND2X1_140/a_16_344#
+ PAND2X1_140/m4_208_n4# PAND2X1_140/O PAND2X1_140/a_56_28# PAND2X1_140/CTRL2 PAND2X1_140/CTRL
+ PAND2X1_140/a_76_28# PAND2X1
XPAND2X1_151 VDD GND POR2X1_150/Y POR2X1_55/Y POR2X1_152/A PAND2X1_151/a_16_344# PAND2X1_151/m4_208_n4#
+ PAND2X1_151/O PAND2X1_151/a_56_28# PAND2X1_151/CTRL2 PAND2X1_151/CTRL PAND2X1_151/a_76_28#
+ PAND2X1
XPAND2X1_162 VDD GND PAND2X1_161/Y PAND2X1_162/A POR2X1_163/A PAND2X1_162/a_16_344#
+ PAND2X1_162/m4_208_n4# PAND2X1_162/O PAND2X1_162/a_56_28# PAND2X1_162/CTRL2 PAND2X1_162/CTRL
+ PAND2X1_162/a_76_28# PAND2X1
XPAND2X1_173 VDD GND POR2X1_186/B PAND2X1_72/A POR2X1_175/B PAND2X1_173/a_16_344#
+ PAND2X1_173/m4_208_n4# PAND2X1_173/O PAND2X1_173/a_56_28# PAND2X1_173/CTRL2 PAND2X1_173/CTRL
+ PAND2X1_173/a_76_28# PAND2X1
XPAND2X1_184 VDD GND PAND2X1_96/B PAND2X1_71/Y POR2X1_456/B PAND2X1_184/a_16_344#
+ PAND2X1_184/m4_208_n4# PAND2X1_184/O PAND2X1_184/a_56_28# PAND2X1_184/CTRL2 PAND2X1_184/CTRL
+ PAND2X1_184/a_76_28# PAND2X1
XPAND2X1_195 VDD GND POR2X1_43/Y POR2X1_41/Y PAND2X1_199/A PAND2X1_195/a_16_344# PAND2X1_195/m4_208_n4#
+ PAND2X1_195/O PAND2X1_195/a_56_28# PAND2X1_195/CTRL2 PAND2X1_195/CTRL PAND2X1_195/a_76_28#
+ PAND2X1
XPOR2X1_209 VDD GND POR2X1_149/Y POR2X1_209/A POR2X1_213/B POR2X1_209/m4_208_n4# POR2X1_209/O
+ POR2X1_209/CTRL2 POR2X1_209/a_16_28# POR2X1_209/CTRL POR2X1_209/a_76_344# POR2X1_209/a_56_344#
+ POR2X1
XPOR2X1_710 VDD GND POR2X1_710/B POR2X1_710/A POR2X1_710/Y POR2X1_710/m4_208_n4# POR2X1_710/O
+ POR2X1_710/CTRL2 POR2X1_710/a_16_28# POR2X1_710/CTRL POR2X1_710/a_76_344# POR2X1_710/a_56_344#
+ POR2X1
XPOR2X1_721 VDD GND POR2X1_673/Y POR2X1_720/Y POR2X1_734/A POR2X1_721/m4_208_n4# POR2X1_721/O
+ POR2X1_721/CTRL2 POR2X1_721/a_16_28# POR2X1_721/CTRL POR2X1_721/a_76_344# POR2X1_721/a_56_344#
+ POR2X1
XPOR2X1_743 VDD GND POR2X1_7/B POR2X1_153/Y POR2X1_743/Y POR2X1_743/m4_208_n4# POR2X1_743/O
+ POR2X1_743/CTRL2 POR2X1_743/a_16_28# POR2X1_743/CTRL POR2X1_743/a_76_344# POR2X1_743/a_56_344#
+ POR2X1
XPOR2X1_732 VDD GND POR2X1_732/B POR2X1_725/Y POR2X1_738/A POR2X1_732/m4_208_n4# POR2X1_732/O
+ POR2X1_732/CTRL2 POR2X1_732/a_16_28# POR2X1_732/CTRL POR2X1_732/a_76_344# POR2X1_732/a_56_344#
+ POR2X1
XPOR2X1_754 VDD GND POR2X1_39/B POR2X1_754/A POR2X1_754/Y POR2X1_754/m4_208_n4# POR2X1_754/O
+ POR2X1_754/CTRL2 POR2X1_754/a_16_28# POR2X1_754/CTRL POR2X1_754/a_76_344# POR2X1_754/a_56_344#
+ POR2X1
XPOR2X1_776 VDD GND POR2X1_776/B POR2X1_776/A POR2X1_785/A POR2X1_776/m4_208_n4# POR2X1_776/O
+ POR2X1_776/CTRL2 POR2X1_776/a_16_28# POR2X1_776/CTRL POR2X1_776/a_76_344# POR2X1_776/a_56_344#
+ POR2X1
XPOR2X1_765 VDD GND POR2X1_13/A POR2X1_16/A POR2X1_765/Y POR2X1_765/m4_208_n4# POR2X1_765/O
+ POR2X1_765/CTRL2 POR2X1_765/a_16_28# POR2X1_765/CTRL POR2X1_765/a_76_344# POR2X1_765/a_56_344#
+ POR2X1
XPOR2X1_787 VDD GND POR2X1_370/Y POR2X1_556/A POR2X1_794/B POR2X1_787/m4_208_n4# POR2X1_787/O
+ POR2X1_787/CTRL2 POR2X1_787/a_16_28# POR2X1_787/CTRL POR2X1_787/a_76_344# POR2X1_787/a_56_344#
+ POR2X1
XPOR2X1_798 VDD GND POR2X1_319/Y POR2X1_468/B POR2X1_802/B POR2X1_798/m4_208_n4# POR2X1_798/O
+ POR2X1_798/CTRL2 POR2X1_798/a_16_28# POR2X1_798/CTRL POR2X1_798/a_76_344# POR2X1_798/a_56_344#
+ POR2X1
XPAND2X1_717 VDD GND PAND2X1_493/Y PAND2X1_717/A PAND2X1_717/Y PAND2X1_717/a_16_344#
+ PAND2X1_717/m4_208_n4# PAND2X1_717/O PAND2X1_717/a_56_28# PAND2X1_717/CTRL2 PAND2X1_717/CTRL
+ PAND2X1_717/a_76_28# PAND2X1
XPAND2X1_728 VDD GND POR2X1_680/Y POR2X1_679/Y PAND2X1_730/A PAND2X1_728/a_16_344#
+ PAND2X1_728/m4_208_n4# PAND2X1_728/O PAND2X1_728/a_56_28# PAND2X1_728/CTRL2 PAND2X1_728/CTRL
+ PAND2X1_728/a_76_28# PAND2X1
XPAND2X1_706 VDD GND POR2X1_693/Y POR2X1_692/Y PAND2X1_713/B PAND2X1_706/a_16_344#
+ PAND2X1_706/m4_208_n4# PAND2X1_706/O PAND2X1_706/a_56_28# PAND2X1_706/CTRL2 PAND2X1_706/CTRL
+ PAND2X1_706/a_76_28# PAND2X1
XPAND2X1_739 VDD GND PAND2X1_739/B PAND2X1_192/Y PAND2X1_739/Y PAND2X1_739/a_16_344#
+ PAND2X1_739/m4_208_n4# PAND2X1_739/O PAND2X1_739/a_56_28# PAND2X1_739/CTRL2 PAND2X1_739/CTRL
+ PAND2X1_739/a_76_28# PAND2X1
XPOR2X1_3 VDD GND POR2X1_3/B POR2X1_3/A POR2X1_7/B POR2X1_3/m4_208_n4# POR2X1_3/O
+ POR2X1_3/CTRL2 POR2X1_3/a_16_28# POR2X1_3/CTRL POR2X1_3/a_76_344# POR2X1_3/a_56_344#
+ POR2X1
XPOR2X1_562 VDD GND POR2X1_562/B POR2X1_556/Y POR2X1_570/B POR2X1_562/m4_208_n4# POR2X1_562/O
+ POR2X1_562/CTRL2 POR2X1_562/a_16_28# POR2X1_562/CTRL POR2X1_562/a_76_344# POR2X1_562/a_56_344#
+ POR2X1
XPOR2X1_540 VDD GND POR2X1_181/B POR2X1_540/A POR2X1_540/Y POR2X1_540/m4_208_n4# POR2X1_540/O
+ POR2X1_540/CTRL2 POR2X1_540/a_16_28# POR2X1_540/CTRL POR2X1_540/a_76_344# POR2X1_540/a_56_344#
+ POR2X1
XPOR2X1_551 VDD GND POR2X1_544/Y POR2X1_551/A POR2X1_564/B POR2X1_551/m4_208_n4# POR2X1_551/O
+ POR2X1_551/CTRL2 POR2X1_551/a_16_28# POR2X1_551/CTRL POR2X1_551/a_76_344# POR2X1_551/a_56_344#
+ POR2X1
XPOR2X1_595 VDD GND POR2X1_83/B POR2X1_250/A POR2X1_595/Y POR2X1_595/m4_208_n4# POR2X1_595/O
+ POR2X1_595/CTRL2 POR2X1_595/a_16_28# POR2X1_595/CTRL POR2X1_595/a_76_344# POR2X1_595/a_56_344#
+ POR2X1
XPOR2X1_573 VDD GND POR2X1_404/Y POR2X1_573/A POR2X1_575/B POR2X1_573/m4_208_n4# POR2X1_573/O
+ POR2X1_573/CTRL2 POR2X1_573/a_16_28# POR2X1_573/CTRL POR2X1_573/a_76_344# POR2X1_573/a_56_344#
+ POR2X1
XPOR2X1_584 VDD GND POR2X1_7/A POR2X1_52/A POR2X1_584/Y POR2X1_584/m4_208_n4# POR2X1_584/O
+ POR2X1_584/CTRL2 POR2X1_584/a_16_28# POR2X1_584/CTRL POR2X1_584/a_76_344# POR2X1_584/a_56_344#
+ POR2X1
XPAND2X1_503 VDD GND POR2X1_502/Y PAND2X1_65/B POR2X1_509/A PAND2X1_503/a_16_344#
+ POR2X1_227/m4_208_n4# PAND2X1_503/O PAND2X1_503/a_56_28# PAND2X1_503/CTRL2 PAND2X1_503/CTRL
+ PAND2X1_503/a_76_28# PAND2X1
XPAND2X1_525 VDD GND PAND2X1_52/B POR2X1_294/B POR2X1_546/B PAND2X1_525/a_16_344#
+ POR2X1_546/m4_208_n4# PAND2X1_525/O PAND2X1_525/a_56_28# PAND2X1_525/CTRL2 PAND2X1_525/CTRL
+ PAND2X1_525/a_76_28# PAND2X1
XPAND2X1_536 VDD GND POR2X1_590/A POR2X1_260/B POR2X1_537/A PAND2X1_536/a_16_344#
+ PAND2X1_536/m4_208_n4# PAND2X1_536/O PAND2X1_536/a_56_28# PAND2X1_536/CTRL2 PAND2X1_536/CTRL
+ PAND2X1_536/a_76_28# PAND2X1
XPAND2X1_514 VDD GND POR2X1_136/Y D_INPUT_0 PAND2X1_514/Y PAND2X1_514/a_16_344# PAND2X1_514/m4_208_n4#
+ PAND2X1_514/O PAND2X1_514/a_56_28# PAND2X1_514/CTRL2 PAND2X1_514/CTRL PAND2X1_514/a_76_28#
+ PAND2X1
XPAND2X1_558 VDD GND POR2X1_494/Y PAND2X1_493/Y PAND2X1_558/Y PAND2X1_558/a_16_344#
+ PAND2X1_558/m4_208_n4# PAND2X1_558/O PAND2X1_558/a_56_28# PAND2X1_558/CTRL2 PAND2X1_558/CTRL
+ PAND2X1_558/a_76_28# PAND2X1
XPAND2X1_547 VDD GND POR2X1_528/Y POR2X1_527/Y PAND2X1_550/B PAND2X1_547/a_16_344#
+ PAND2X1_547/m4_208_n4# PAND2X1_547/O PAND2X1_547/a_56_28# PAND2X1_547/CTRL2 PAND2X1_547/CTRL
+ PAND2X1_547/a_76_28# PAND2X1
XPAND2X1_569 VDD GND PAND2X1_569/B PAND2X1_569/A PAND2X1_569/Y PAND2X1_569/a_16_344#
+ PAND2X1_770/m4_208_n4# PAND2X1_569/O PAND2X1_569/a_56_28# PAND2X1_569/CTRL2 PAND2X1_569/CTRL
+ PAND2X1_569/a_76_28# PAND2X1
XPOR2X1_370 VDD GND POR2X1_335/B POR2X1_543/A POR2X1_370/Y POR2X1_370/m4_208_n4# POR2X1_370/O
+ POR2X1_370/CTRL2 POR2X1_370/a_16_28# POR2X1_370/CTRL POR2X1_370/a_76_344# POR2X1_370/a_56_344#
+ POR2X1
XPOR2X1_381 VDD GND D_INPUT_3 POR2X1_13/A POR2X1_817/A POR2X1_381/m4_208_n4# POR2X1_381/O
+ POR2X1_381/CTRL2 POR2X1_381/a_16_28# POR2X1_381/CTRL POR2X1_381/a_76_344# POR2X1_381/a_56_344#
+ POR2X1
XPOR2X1_392 VDD GND POR2X1_392/B POR2X1_391/Y POR2X1_860/A POR2X1_392/m4_208_n4# POR2X1_392/O
+ POR2X1_392/CTRL2 POR2X1_392/a_16_28# POR2X1_392/CTRL POR2X1_392/a_76_344# POR2X1_392/a_56_344#
+ POR2X1
XPAND2X1_311 VDD GND POR2X1_590/A POR2X1_66/A POR2X1_538/A PAND2X1_311/a_16_344# PAND2X1_311/m4_208_n4#
+ PAND2X1_311/O PAND2X1_311/a_56_28# PAND2X1_311/CTRL2 PAND2X1_311/CTRL PAND2X1_311/a_76_28#
+ PAND2X1
XPAND2X1_300 VDD GND POR2X1_121/B PAND2X1_60/B POR2X1_301/A PAND2X1_300/a_16_344#
+ PAND2X1_300/m4_208_n4# PAND2X1_300/O PAND2X1_300/a_56_28# PAND2X1_300/CTRL2 PAND2X1_300/CTRL
+ PAND2X1_300/a_76_28# PAND2X1
XPAND2X1_355 VDD GND POR2X1_331/Y POR2X1_329/Y PAND2X1_356/B PAND2X1_355/a_16_344#
+ PAND2X1_355/m4_208_n4# PAND2X1_355/O PAND2X1_355/a_56_28# PAND2X1_355/CTRL2 PAND2X1_355/CTRL
+ PAND2X1_355/a_76_28# PAND2X1
XPAND2X1_333 VDD GND POR2X1_289/Y POR2X1_171/Y PAND2X1_333/Y PAND2X1_333/a_16_344#
+ PAND2X1_333/m4_208_n4# PAND2X1_333/O PAND2X1_333/a_56_28# PAND2X1_333/CTRL2 PAND2X1_333/CTRL
+ PAND2X1_333/a_76_28# PAND2X1
XPAND2X1_322 VDD GND POR2X1_502/A PAND2X1_57/B POR2X1_325/B PAND2X1_322/a_16_344#
+ PAND2X1_322/m4_208_n4# PAND2X1_322/O PAND2X1_322/a_56_28# PAND2X1_322/CTRL2 PAND2X1_322/CTRL
+ PAND2X1_322/a_76_28# PAND2X1
XPAND2X1_344 VDD GND POR2X1_256/Y PAND2X1_254/Y PAND2X1_348/A PAND2X1_344/a_16_344#
+ PAND2X1_344/m4_208_n4# PAND2X1_344/O PAND2X1_344/a_56_28# PAND2X1_344/CTRL2 PAND2X1_344/CTRL
+ PAND2X1_344/a_76_28# PAND2X1
XPAND2X1_366 VDD GND PAND2X1_363/Y PAND2X1_366/A PAND2X1_366/Y PAND2X1_366/a_16_344#
+ PAND2X1_366/m4_208_n4# PAND2X1_366/O PAND2X1_366/a_56_28# PAND2X1_366/CTRL2 PAND2X1_366/CTRL
+ PAND2X1_366/a_76_28# PAND2X1
XPAND2X1_377 VDD GND POR2X1_14/Y POR2X1_66/B PAND2X1_377/Y PAND2X1_377/a_16_344# PAND2X1_376/m4_208_n4#
+ PAND2X1_377/O PAND2X1_377/a_56_28# PAND2X1_377/CTRL2 PAND2X1_377/CTRL PAND2X1_377/a_76_28#
+ PAND2X1
XPAND2X1_388 VDD GND POR2X1_176/Y POR2X1_167/Y PAND2X1_388/Y PAND2X1_388/a_16_344#
+ PAND2X1_439/m4_208_n4# PAND2X1_388/O PAND2X1_388/a_56_28# PAND2X1_388/CTRL2 PAND2X1_388/CTRL
+ PAND2X1_388/a_76_28# PAND2X1
XPAND2X1_399 VDD GND POR2X1_398/Y PAND2X1_57/B POR2X1_403/B PAND2X1_399/a_16_344#
+ PAND2X1_399/m4_208_n4# PAND2X1_399/O PAND2X1_399/a_56_28# PAND2X1_399/CTRL2 PAND2X1_399/CTRL
+ PAND2X1_399/a_76_28# PAND2X1
XPAND2X1_130 VDD GND POR2X1_129/Y POR2X1_7/A POR2X1_131/A PAND2X1_130/a_16_344# PAND2X1_130/m4_208_n4#
+ PAND2X1_130/O PAND2X1_130/a_56_28# PAND2X1_130/CTRL2 PAND2X1_130/CTRL PAND2X1_130/a_76_28#
+ PAND2X1
XPAND2X1_141 VDD GND PAND2X1_140/Y PAND2X1_139/Y PAND2X1_217/B PAND2X1_141/a_16_344#
+ PAND2X1_141/m4_208_n4# PAND2X1_141/O PAND2X1_141/a_56_28# PAND2X1_141/CTRL2 PAND2X1_141/CTRL
+ PAND2X1_141/a_76_28# PAND2X1
XPAND2X1_152 VDD GND POR2X1_151/Y PAND2X1_48/B POR2X1_209/A PAND2X1_152/a_16_344#
+ PAND2X1_152/m4_208_n4# PAND2X1_152/O PAND2X1_152/a_56_28# PAND2X1_152/CTRL2 PAND2X1_152/CTRL
+ PAND2X1_152/a_76_28# PAND2X1
XPAND2X1_163 VDD GND POR2X1_162/Y PAND2X1_52/B POR2X1_210/A PAND2X1_163/a_16_344#
+ PAND2X1_163/m4_208_n4# PAND2X1_163/O PAND2X1_163/a_56_28# PAND2X1_163/CTRL2 PAND2X1_163/CTRL
+ PAND2X1_163/a_76_28# PAND2X1
XPAND2X1_185 VDD GND POR2X1_73/Y POR2X1_55/Y POR2X1_816/A PAND2X1_185/a_16_344# PAND2X1_185/m4_208_n4#
+ PAND2X1_185/O PAND2X1_185/a_56_28# PAND2X1_185/CTRL2 PAND2X1_185/CTRL PAND2X1_185/a_76_28#
+ PAND2X1
XPAND2X1_174 VDD GND POR2X1_172/Y POR2X1_171/Y PAND2X1_175/B PAND2X1_174/a_16_344#
+ PAND2X1_174/m4_208_n4# PAND2X1_174/O PAND2X1_174/a_56_28# PAND2X1_174/CTRL2 PAND2X1_174/CTRL
+ PAND2X1_174/a_76_28# PAND2X1
XPAND2X1_196 VDD GND POR2X1_48/Y POR2X1_45/Y PAND2X1_199/B PAND2X1_196/a_16_344# PAND2X1_196/m4_208_n4#
+ PAND2X1_196/O PAND2X1_196/a_56_28# PAND2X1_196/CTRL2 PAND2X1_196/CTRL PAND2X1_196/a_76_28#
+ PAND2X1
XPOR2X1_700 VDD GND POR2X1_60/A POR2X1_90/Y POR2X1_700/Y POR2X1_700/m4_208_n4# POR2X1_700/O
+ POR2X1_700/CTRL2 POR2X1_700/a_16_28# POR2X1_700/CTRL POR2X1_700/a_76_344# POR2X1_700/a_56_344#
+ POR2X1
XPOR2X1_711 VDD GND POR2X1_711/B POR2X1_710/Y POR2X1_711/Y POR2X1_711/m4_208_n4# POR2X1_711/O
+ POR2X1_711/CTRL2 POR2X1_711/a_16_28# POR2X1_711/CTRL POR2X1_711/a_76_344# POR2X1_711/a_56_344#
+ POR2X1
XPOR2X1_744 VDD GND POR2X1_57/A POR2X1_394/A POR2X1_744/Y POR2X1_744/m4_208_n4# POR2X1_744/O
+ POR2X1_744/CTRL2 POR2X1_744/a_16_28# POR2X1_744/CTRL POR2X1_744/a_76_344# POR2X1_744/a_56_344#
+ POR2X1
XPOR2X1_722 VDD GND POR2X1_722/B POR2X1_722/A POR2X1_722/Y POR2X1_722/m4_208_n4# POR2X1_722/O
+ POR2X1_722/CTRL2 POR2X1_722/a_16_28# POR2X1_722/CTRL POR2X1_722/a_76_344# POR2X1_722/a_56_344#
+ POR2X1
XPOR2X1_733 VDD GND POR2X1_722/Y POR2X1_733/A POR2X1_733/Y POR2X1_733/m4_208_n4# POR2X1_733/O
+ POR2X1_733/CTRL2 POR2X1_733/a_16_28# POR2X1_733/CTRL POR2X1_733/a_76_344# POR2X1_733/a_56_344#
+ POR2X1
XPOR2X1_755 VDD GND POR2X1_60/A POR2X1_665/A POR2X1_755/Y POR2X1_755/m4_208_n4# POR2X1_755/O
+ POR2X1_755/CTRL2 POR2X1_755/a_16_28# POR2X1_755/CTRL POR2X1_755/a_76_344# POR2X1_755/a_56_344#
+ POR2X1
XPOR2X1_766 VDD GND POR2X1_65/A POR2X1_90/Y POR2X1_766/Y POR2X1_766/m4_208_n4# POR2X1_766/O
+ POR2X1_766/CTRL2 POR2X1_766/a_16_28# POR2X1_766/CTRL POR2X1_766/a_76_344# POR2X1_766/a_56_344#
+ POR2X1
XPOR2X1_788 VDD GND POR2X1_788/B POR2X1_788/A POR2X1_788/Y POR2X1_788/m4_208_n4# POR2X1_788/O
+ POR2X1_788/CTRL2 POR2X1_788/a_16_28# POR2X1_788/CTRL POR2X1_788/a_76_344# POR2X1_788/a_56_344#
+ POR2X1
XPOR2X1_777 VDD GND POR2X1_777/B POR2X1_307/A POR2X1_777/Y POR2X1_777/m4_208_n4# POR2X1_777/O
+ POR2X1_777/CTRL2 POR2X1_777/a_16_28# POR2X1_777/CTRL POR2X1_777/a_76_344# POR2X1_777/a_56_344#
+ POR2X1
XPOR2X1_799 VDD GND POR2X1_567/A POR2X1_652/A POR2X1_802/A POR2X1_593/m4_208_n4# POR2X1_799/O
+ POR2X1_799/CTRL2 POR2X1_799/a_16_28# POR2X1_799/CTRL POR2X1_799/a_76_344# POR2X1_799/a_56_344#
+ POR2X1
XPAND2X1_729 VDD GND PAND2X1_691/Y PAND2X1_687/Y PAND2X1_730/B PAND2X1_729/a_16_344#
+ PAND2X1_729/m4_208_n4# PAND2X1_729/O PAND2X1_729/a_56_28# PAND2X1_729/CTRL2 PAND2X1_729/CTRL
+ PAND2X1_729/a_76_28# PAND2X1
XPAND2X1_707 VDD GND POR2X1_695/Y POR2X1_694/Y PAND2X1_707/Y PAND2X1_707/a_16_344#
+ PAND2X1_707/m4_208_n4# PAND2X1_707/O PAND2X1_707/a_56_28# PAND2X1_707/CTRL2 PAND2X1_707/CTRL
+ PAND2X1_707/a_76_28# PAND2X1
XPAND2X1_718 VDD GND PAND2X1_645/B POR2X1_591/Y PAND2X1_718/Y PAND2X1_718/a_16_344#
+ PAND2X1_718/m4_208_n4# PAND2X1_718/O PAND2X1_718/a_56_28# PAND2X1_718/CTRL2 PAND2X1_718/CTRL
+ PAND2X1_718/a_76_28# PAND2X1
XPOR2X1_4 VDD GND D_INPUT_0 INPUT_1 POR2X1_4/Y POR2X1_4/m4_208_n4# POR2X1_4/O POR2X1_4/CTRL2
+ POR2X1_4/a_16_28# POR2X1_4/CTRL POR2X1_4/a_76_344# POR2X1_4/a_56_344# POR2X1
XPOR2X1_541 VDD GND POR2X1_541/B POR2X1_274/B POR2X1_553/A POR2X1_541/m4_208_n4# POR2X1_541/O
+ POR2X1_541/CTRL2 POR2X1_541/a_16_28# POR2X1_541/CTRL POR2X1_541/a_76_344# POR2X1_541/a_56_344#
+ POR2X1
XPOR2X1_530 VDD GND POR2X1_39/B POR2X1_102/Y POR2X1_530/Y POR2X1_530/m4_208_n4# POR2X1_530/O
+ POR2X1_530/CTRL2 POR2X1_530/a_16_28# POR2X1_530/CTRL POR2X1_530/a_76_344# POR2X1_530/a_56_344#
+ POR2X1
XPOR2X1_552 VDD GND POR2X1_542/Y POR2X1_552/A POR2X1_552/Y POR2X1_552/m4_208_n4# POR2X1_552/O
+ POR2X1_552/CTRL2 POR2X1_552/a_16_28# POR2X1_552/CTRL POR2X1_552/a_76_344# POR2X1_552/a_56_344#
+ POR2X1
XPOR2X1_563 VDD GND POR2X1_553/Y POR2X1_554/Y POR2X1_563/Y POR2X1_563/m4_208_n4# POR2X1_563/O
+ POR2X1_563/CTRL2 POR2X1_563/a_16_28# POR2X1_563/CTRL POR2X1_563/a_76_344# POR2X1_563/a_56_344#
+ POR2X1
XPOR2X1_574 VDD GND POR2X1_510/Y POR2X1_574/A POR2X1_574/Y POR2X1_574/m4_208_n4# POR2X1_574/O
+ POR2X1_574/CTRL2 POR2X1_574/a_16_28# POR2X1_574/CTRL POR2X1_574/a_76_344# POR2X1_574/a_56_344#
+ POR2X1
XPOR2X1_596 VDD GND PAND2X1_57/B POR2X1_596/A POR2X1_596/Y POR2X1_596/m4_208_n4# POR2X1_596/O
+ POR2X1_596/CTRL2 POR2X1_596/a_16_28# POR2X1_596/CTRL POR2X1_596/a_76_344# POR2X1_596/a_56_344#
+ POR2X1
XPOR2X1_585 VDD GND POR2X1_43/B POR2X1_293/Y POR2X1_585/Y POR2X1_585/m4_208_n4# POR2X1_585/O
+ POR2X1_585/CTRL2 POR2X1_585/a_16_28# POR2X1_585/CTRL POR2X1_585/a_76_344# POR2X1_585/a_56_344#
+ POR2X1
XPAND2X1_504 VDD GND POR2X1_260/A POR2X1_294/B POR2X1_507/B PAND2X1_504/a_16_344#
+ PAND2X1_504/m4_208_n4# PAND2X1_504/O PAND2X1_504/a_56_28# PAND2X1_504/CTRL2 PAND2X1_504/CTRL
+ PAND2X1_504/a_76_28# PAND2X1
XPAND2X1_537 VDD GND POR2X1_536/Y POR2X1_385/Y PAND2X1_643/A PAND2X1_537/a_16_344#
+ PAND2X1_537/m4_208_n4# PAND2X1_537/O PAND2X1_537/a_56_28# PAND2X1_537/CTRL2 PAND2X1_537/CTRL
+ PAND2X1_537/a_76_28# PAND2X1
XPAND2X1_526 VDD GND POR2X1_750/B PAND2X1_32/B POR2X1_546/A PAND2X1_526/a_16_344#
+ PAND2X1_526/m4_208_n4# PAND2X1_526/O PAND2X1_526/a_56_28# PAND2X1_526/CTRL2 PAND2X1_526/CTRL
+ PAND2X1_526/a_76_28# PAND2X1
XPAND2X1_515 VDD GND PAND2X1_514/Y POR2X1_417/Y POR2X1_516/A PAND2X1_515/a_16_344#
+ PAND2X1_515/m4_208_n4# PAND2X1_515/O PAND2X1_515/a_56_28# PAND2X1_515/CTRL2 PAND2X1_515/CTRL
+ PAND2X1_515/a_76_28# PAND2X1
XPAND2X1_548 VDD GND POR2X1_530/Y POR2X1_529/Y PAND2X1_549/B PAND2X1_548/a_16_344#
+ PAND2X1_548/m4_208_n4# PAND2X1_548/O PAND2X1_548/a_56_28# PAND2X1_548/CTRL2 PAND2X1_548/CTRL
+ PAND2X1_548/a_76_28# PAND2X1
XPAND2X1_559 VDD GND PAND2X1_642/B POR2X1_517/Y PAND2X1_560/B PAND2X1_559/a_16_344#
+ PAND2X1_559/m4_208_n4# PAND2X1_559/O PAND2X1_559/a_56_28# PAND2X1_559/CTRL2 PAND2X1_559/CTRL
+ PAND2X1_559/a_76_28# PAND2X1
XPOR2X1_360 VDD GND POR2X1_244/Y POR2X1_360/A POR2X1_363/A POR2X1_360/m4_208_n4# POR2X1_360/O
+ POR2X1_360/CTRL2 POR2X1_360/a_16_28# POR2X1_360/CTRL POR2X1_360/a_76_344# POR2X1_360/a_56_344#
+ POR2X1
XPOR2X1_371 VDD GND POR2X1_5/Y POR2X1_32/A POR2X1_372/A POR2X1_371/m4_208_n4# POR2X1_371/O
+ POR2X1_371/CTRL2 POR2X1_371/a_16_28# POR2X1_371/CTRL POR2X1_371/a_76_344# POR2X1_371/a_56_344#
+ POR2X1
XPOR2X1_393 VDD GND POR2X1_38/Y POR2X1_40/Y POR2X1_393/Y POR2X1_393/m4_208_n4# POR2X1_393/O
+ POR2X1_393/CTRL2 POR2X1_393/a_16_28# POR2X1_393/CTRL POR2X1_393/a_76_344# POR2X1_393/a_56_344#
+ POR2X1
XPOR2X1_382 VDD GND POR2X1_38/B POR2X1_817/A POR2X1_382/Y POR2X1_382/m4_208_n4# POR2X1_382/O
+ POR2X1_382/CTRL2 POR2X1_382/a_16_28# POR2X1_382/CTRL POR2X1_382/a_76_344# POR2X1_382/a_56_344#
+ POR2X1
XPAND2X1_312 VDD GND PAND2X1_65/B PAND2X1_55/Y POR2X1_703/A PAND2X1_312/a_16_344#
+ PAND2X1_312/m4_208_n4# PAND2X1_312/O PAND2X1_312/a_56_28# PAND2X1_312/CTRL2 PAND2X1_312/CTRL
+ PAND2X1_312/a_76_28# PAND2X1
XPAND2X1_301 VDD GND POR2X1_300/Y POR2X1_75/Y PAND2X1_716/B PAND2X1_301/a_16_344#
+ PAND2X1_301/m4_208_n4# PAND2X1_301/O PAND2X1_301/a_56_28# PAND2X1_301/CTRL2 PAND2X1_301/CTRL
+ PAND2X1_301/a_76_28# PAND2X1
XPAND2X1_323 VDD GND PAND2X1_111/B PAND2X1_96/B POR2X1_325/A PAND2X1_323/a_16_344#
+ PAND2X1_323/m4_208_n4# PAND2X1_323/O PAND2X1_323/a_56_28# PAND2X1_323/CTRL2 PAND2X1_323/CTRL
+ PAND2X1_323/a_76_28# PAND2X1
XPAND2X1_345 VDD GND POR2X1_261/Y PAND2X1_555/A PAND2X1_345/Y PAND2X1_345/a_16_344#
+ PAND2X1_345/m4_208_n4# PAND2X1_345/O PAND2X1_345/a_56_28# PAND2X1_345/CTRL2 PAND2X1_345/CTRL
+ PAND2X1_345/a_76_28# PAND2X1
XPAND2X1_334 VDD GND POR2X1_291/Y POR2X1_290/Y PAND2X1_338/B PAND2X1_334/a_16_344#
+ PAND2X1_334/m4_208_n4# PAND2X1_334/O PAND2X1_334/a_56_28# PAND2X1_334/CTRL2 PAND2X1_334/CTRL
+ PAND2X1_334/a_76_28# PAND2X1
XPAND2X1_356 VDD GND PAND2X1_356/B PAND2X1_354/Y PAND2X1_365/A PAND2X1_356/a_16_344#
+ PAND2X1_356/m4_208_n4# PAND2X1_356/O PAND2X1_356/a_56_28# PAND2X1_356/CTRL2 PAND2X1_356/CTRL
+ PAND2X1_356/a_76_28# PAND2X1
XPAND2X1_367 VDD GND PAND2X1_366/Y PAND2X1_367/A GATE_366 PAND2X1_367/a_16_344# PAND2X1_367/m4_208_n4#
+ PAND2X1_367/O PAND2X1_367/a_56_28# PAND2X1_367/CTRL2 PAND2X1_367/CTRL PAND2X1_367/a_76_28#
+ PAND2X1
XPAND2X1_378 VDD GND PAND2X1_377/Y POR2X1_42/Y POR2X1_459/A PAND2X1_378/a_16_344#
+ PAND2X1_378/m4_208_n4# PAND2X1_378/O PAND2X1_378/a_56_28# PAND2X1_378/CTRL2 PAND2X1_378/CTRL
+ PAND2X1_378/a_76_28# PAND2X1
XPAND2X1_389 VDD GND POR2X1_387/Y POR2X1_385/Y PAND2X1_389/Y PAND2X1_389/a_16_344#
+ PAND2X1_389/m4_208_n4# PAND2X1_389/O PAND2X1_389/a_56_28# PAND2X1_389/CTRL2 PAND2X1_389/CTRL
+ PAND2X1_389/a_76_28# PAND2X1
XPOR2X1_190 VDD GND POR2X1_540/A POR2X1_456/B POR2X1_190/Y POR2X1_190/m4_208_n4# POR2X1_190/O
+ POR2X1_190/CTRL2 POR2X1_190/a_16_28# POR2X1_190/CTRL POR2X1_190/a_76_344# POR2X1_190/a_56_344#
+ POR2X1
XPAND2X1_120 VDD GND POR2X1_38/Y POR2X1_41/B POR2X1_666/A PAND2X1_120/a_16_344# PAND2X1_120/m4_208_n4#
+ PAND2X1_120/O PAND2X1_120/a_56_28# PAND2X1_120/CTRL2 PAND2X1_120/CTRL PAND2X1_120/a_76_28#
+ PAND2X1
XPAND2X1_131 VDD GND POR2X1_130/Y POR2X1_260/B POR2X1_140/A PAND2X1_131/a_16_344#
+ PAND2X1_131/m4_208_n4# PAND2X1_131/O PAND2X1_131/a_56_28# PAND2X1_131/CTRL2 PAND2X1_131/CTRL
+ PAND2X1_131/a_76_28# PAND2X1
XPAND2X1_153 VDD GND PAND2X1_90/A D_INPUT_1 POR2X1_407/A PAND2X1_153/a_16_344# PAND2X1_153/m4_208_n4#
+ PAND2X1_153/O PAND2X1_153/a_56_28# PAND2X1_153/CTRL2 PAND2X1_153/CTRL PAND2X1_153/a_76_28#
+ PAND2X1
XPAND2X1_142 VDD GND PAND2X1_65/B POR2X1_68/A POR2X1_830/A PAND2X1_142/a_16_344# PAND2X1_142/m4_208_n4#
+ PAND2X1_142/O PAND2X1_142/a_56_28# PAND2X1_142/CTRL2 PAND2X1_142/CTRL PAND2X1_142/a_76_28#
+ PAND2X1
XPAND2X1_164 VDD GND POR2X1_502/A PAND2X1_20/A POR2X1_776/B PAND2X1_164/a_16_344#
+ PAND2X1_164/m4_208_n4# PAND2X1_164/O PAND2X1_164/a_56_28# PAND2X1_164/CTRL2 PAND2X1_164/CTRL
+ PAND2X1_164/a_76_28# PAND2X1
XPAND2X1_197 VDD GND POR2X1_56/Y POR2X1_52/Y PAND2X1_197/Y PAND2X1_197/a_16_344# PAND2X1_197/m4_208_n4#
+ PAND2X1_197/O PAND2X1_197/a_56_28# PAND2X1_197/CTRL2 PAND2X1_197/CTRL PAND2X1_197/a_76_28#
+ PAND2X1
XPAND2X1_186 VDD GND POR2X1_816/A POR2X1_150/Y POR2X1_594/A PAND2X1_186/a_16_344#
+ PAND2X1_186/m4_208_n4# PAND2X1_186/O PAND2X1_186/a_56_28# PAND2X1_186/CTRL2 PAND2X1_186/CTRL
+ PAND2X1_186/a_76_28# PAND2X1
XPAND2X1_175 VDD GND PAND2X1_175/B POR2X1_173/Y PAND2X1_853/B PAND2X1_175/a_16_344#
+ PAND2X1_175/m4_208_n4# PAND2X1_175/O PAND2X1_175/a_56_28# PAND2X1_175/CTRL2 PAND2X1_175/CTRL
+ PAND2X1_175/a_76_28# PAND2X1
XPOR2X1_701 VDD GND POR2X1_57/A POR2X1_236/Y POR2X1_701/Y POR2X1_701/m4_208_n4# POR2X1_701/O
+ POR2X1_701/CTRL2 POR2X1_701/a_16_28# POR2X1_701/CTRL POR2X1_701/a_76_344# POR2X1_701/a_56_344#
+ POR2X1
XPOR2X1_723 VDD GND POR2X1_723/B POR2X1_717/Y POR2X1_733/A POR2X1_723/m4_208_n4# POR2X1_723/O
+ POR2X1_723/CTRL2 POR2X1_723/a_16_28# POR2X1_723/CTRL POR2X1_723/a_76_344# POR2X1_723/a_56_344#
+ POR2X1
XPOR2X1_745 VDD GND POR2X1_40/Y POR2X1_669/B POR2X1_745/Y POR2X1_745/m4_208_n4# POR2X1_745/O
+ POR2X1_745/CTRL2 POR2X1_745/a_16_28# POR2X1_745/CTRL POR2X1_745/a_76_344# POR2X1_745/a_56_344#
+ POR2X1
XPOR2X1_712 VDD GND POR2X1_707/Y POR2X1_712/A POR2X1_712/Y POR2X1_712/m4_208_n4# POR2X1_712/O
+ POR2X1_712/CTRL2 POR2X1_712/a_16_28# POR2X1_712/CTRL POR2X1_712/a_76_344# POR2X1_712/a_56_344#
+ POR2X1
XPOR2X1_734 VDD GND POR2X1_734/B POR2X1_734/A POR2X1_737/A POR2X1_734/m4_208_n4# POR2X1_734/O
+ POR2X1_734/CTRL2 POR2X1_734/a_16_28# POR2X1_734/CTRL POR2X1_734/a_76_344# POR2X1_734/a_56_344#
+ POR2X1
XPOR2X1_767 VDD GND POR2X1_7/B POR2X1_79/A POR2X1_767/Y POR2X1_767/m4_208_n4# POR2X1_767/O
+ POR2X1_767/CTRL2 POR2X1_767/a_16_28# POR2X1_767/CTRL POR2X1_767/a_76_344# POR2X1_767/a_56_344#
+ POR2X1
XPOR2X1_778 VDD GND POR2X1_778/B POR2X1_499/A POR2X1_784/A POR2X1_778/m4_208_n4# POR2X1_778/O
+ POR2X1_778/CTRL2 POR2X1_778/a_16_28# POR2X1_778/CTRL POR2X1_778/a_76_344# POR2X1_778/a_56_344#
+ POR2X1
XPOR2X1_756 VDD GND POR2X1_814/B POR2X1_750/B POR2X1_756/Y POR2X1_756/m4_208_n4# POR2X1_756/O
+ POR2X1_756/CTRL2 POR2X1_756/a_16_28# POR2X1_756/CTRL POR2X1_756/a_76_344# POR2X1_756/a_56_344#
+ POR2X1
XPOR2X1_789 VDD GND POR2X1_789/B POR2X1_789/A POR2X1_789/Y POR2X1_789/m4_208_n4# POR2X1_789/O
+ POR2X1_789/CTRL2 POR2X1_789/a_16_28# POR2X1_789/CTRL POR2X1_789/a_76_344# POR2X1_789/a_56_344#
+ POR2X1
XPAND2X1_708 VDD GND POR2X1_697/Y POR2X1_696/Y PAND2X1_712/B PAND2X1_708/a_16_344#
+ PAND2X1_708/m4_208_n4# PAND2X1_708/O PAND2X1_708/a_56_28# PAND2X1_708/CTRL2 PAND2X1_708/CTRL
+ PAND2X1_708/a_76_28# PAND2X1
XPAND2X1_719 VDD GND POR2X1_666/Y POR2X1_665/Y PAND2X1_719/Y PAND2X1_719/a_16_344#
+ PAND2X1_719/m4_208_n4# PAND2X1_719/O PAND2X1_719/a_56_28# PAND2X1_719/CTRL2 PAND2X1_719/CTRL
+ PAND2X1_719/a_76_28# PAND2X1
XPOR2X1_5 VDD GND INPUT_2 D_INPUT_3 POR2X1_5/Y POR2X1_5/m4_208_n4# POR2X1_5/O POR2X1_5/CTRL2
+ POR2X1_5/a_16_28# POR2X1_5/CTRL POR2X1_5/a_76_344# POR2X1_5/a_56_344# POR2X1
XPOR2X1_520 VDD GND POR2X1_520/B POR2X1_520/A POR2X1_559/A POR2X1_520/m4_208_n4# POR2X1_520/O
+ POR2X1_520/CTRL2 POR2X1_520/a_16_28# POR2X1_520/CTRL POR2X1_520/a_76_344# POR2X1_520/a_56_344#
+ POR2X1
XPOR2X1_553 VDD GND POR2X1_540/Y POR2X1_553/A POR2X1_553/Y POR2X1_553/m4_208_n4# POR2X1_553/O
+ POR2X1_553/CTRL2 POR2X1_553/a_16_28# POR2X1_553/CTRL POR2X1_553/a_76_344# POR2X1_553/a_56_344#
+ POR2X1
XPOR2X1_542 VDD GND POR2X1_542/B POR2X1_703/A POR2X1_542/Y POR2X1_542/m4_208_n4# POR2X1_542/O
+ POR2X1_542/CTRL2 POR2X1_542/a_16_28# POR2X1_542/CTRL POR2X1_542/a_76_344# POR2X1_542/a_56_344#
+ POR2X1
XPOR2X1_531 VDD GND POR2X1_40/Y POR2X1_73/Y POR2X1_531/Y POR2X1_531/m4_208_n4# POR2X1_531/O
+ POR2X1_531/CTRL2 POR2X1_531/a_16_28# POR2X1_531/CTRL POR2X1_531/a_76_344# POR2X1_531/a_56_344#
+ POR2X1
XPOR2X1_575 VDD GND POR2X1_575/B POR2X1_574/Y POR2X1_579/B POR2X1_575/m4_208_n4# POR2X1_575/O
+ POR2X1_575/CTRL2 POR2X1_575/a_16_28# POR2X1_575/CTRL POR2X1_575/a_76_344# POR2X1_575/a_56_344#
+ POR2X1
XPOR2X1_564 VDD GND POR2X1_564/B POR2X1_552/Y POR2X1_564/Y POR2X1_564/m4_208_n4# POR2X1_564/O
+ POR2X1_564/CTRL2 POR2X1_564/a_16_28# POR2X1_564/CTRL POR2X1_564/a_76_344# POR2X1_564/a_56_344#
+ POR2X1
XPOR2X1_586 VDD GND POR2X1_72/B POR2X1_129/Y POR2X1_586/Y POR2X1_586/m4_208_n4# POR2X1_586/O
+ POR2X1_586/CTRL2 POR2X1_586/a_16_28# POR2X1_586/CTRL POR2X1_586/a_76_344# POR2X1_586/a_56_344#
+ POR2X1
XPOR2X1_597 VDD GND POR2X1_41/B POR2X1_597/A POR2X1_597/Y POR2X1_597/m4_208_n4# POR2X1_597/O
+ POR2X1_597/CTRL2 POR2X1_597/a_16_28# POR2X1_597/CTRL POR2X1_597/a_76_344# POR2X1_597/a_56_344#
+ POR2X1
XPAND2X1_527 VDD GND PAND2X1_111/B PAND2X1_65/B POR2X1_547/B PAND2X1_527/a_16_344#
+ PAND2X1_527/m4_208_n4# PAND2X1_527/O PAND2X1_527/a_56_28# PAND2X1_527/CTRL2 PAND2X1_527/CTRL
+ PAND2X1_527/a_76_28# PAND2X1
XPAND2X1_516 VDD GND POR2X1_515/Y POR2X1_513/Y POR2X1_574/A PAND2X1_516/a_16_344#
+ PAND2X1_516/m4_208_n4# PAND2X1_516/O PAND2X1_516/a_56_28# PAND2X1_516/CTRL2 PAND2X1_516/CTRL
+ PAND2X1_516/a_76_28# PAND2X1
XPAND2X1_505 VDD GND PAND2X1_23/Y PAND2X1_20/A POR2X1_507/A PAND2X1_505/a_16_344#
+ PAND2X1_505/m4_208_n4# PAND2X1_505/O PAND2X1_505/a_56_28# PAND2X1_505/CTRL2 PAND2X1_505/CTRL
+ PAND2X1_505/a_76_28# PAND2X1
XPAND2X1_538 VDD GND POR2X1_311/Y POR2X1_13/Y PAND2X1_539/B PAND2X1_538/a_16_344#
+ PAND2X1_802/m4_208_n4# PAND2X1_538/O PAND2X1_538/a_56_28# PAND2X1_538/CTRL2 PAND2X1_538/CTRL
+ PAND2X1_538/a_76_28# PAND2X1
XPAND2X1_549 VDD GND PAND2X1_549/B POR2X1_531/Y PAND2X1_565/A PAND2X1_549/a_16_344#
+ PAND2X1_549/m4_208_n4# PAND2X1_549/O PAND2X1_549/a_56_28# PAND2X1_549/CTRL2 PAND2X1_549/CTRL
+ PAND2X1_549/a_76_28# PAND2X1
XPOR2X1_350 VDD GND POR2X1_350/B POR2X1_341/Y POR2X1_350/Y POR2X1_502/m4_208_n4# POR2X1_350/O
+ POR2X1_350/CTRL2 POR2X1_350/a_16_28# POR2X1_350/CTRL POR2X1_350/a_76_344# POR2X1_350/a_56_344#
+ POR2X1
XPOR2X1_361 VDD GND POR2X1_267/Y POR2X1_276/Y POR2X1_362/A POR2X1_361/m4_208_n4# POR2X1_361/O
+ POR2X1_361/CTRL2 POR2X1_361/a_16_28# POR2X1_361/CTRL POR2X1_361/a_76_344# POR2X1_361/a_56_344#
+ POR2X1
XPOR2X1_394 VDD GND POR2X1_48/A POR2X1_394/A POR2X1_394/Y POR2X1_394/m4_208_n4# POR2X1_394/O
+ POR2X1_394/CTRL2 POR2X1_394/a_16_28# POR2X1_394/CTRL POR2X1_394/a_76_344# POR2X1_394/a_56_344#
+ POR2X1
XPOR2X1_383 VDD GND PAND2X1_90/Y POR2X1_383/A POR2X1_383/Y POR2X1_383/m4_208_n4# POR2X1_383/O
+ POR2X1_383/CTRL2 POR2X1_383/a_16_28# POR2X1_383/CTRL POR2X1_383/a_76_344# POR2X1_383/a_56_344#
+ POR2X1
XPOR2X1_372 VDD GND INPUT_1 POR2X1_372/A POR2X1_372/Y POR2X1_372/m4_208_n4# POR2X1_372/O
+ POR2X1_372/CTRL2 POR2X1_372/a_16_28# POR2X1_372/CTRL POR2X1_372/a_76_344# POR2X1_372/a_56_344#
+ POR2X1
XPAND2X1_302 VDD GND POR2X1_299/Y POR2X1_298/Y PAND2X1_303/B PAND2X1_302/a_16_344#
+ PAND2X1_302/m4_208_n4# PAND2X1_302/O PAND2X1_302/a_56_28# PAND2X1_302/CTRL2 PAND2X1_302/CTRL
+ PAND2X1_302/a_76_28# PAND2X1
XPAND2X1_313 VDD GND PAND2X1_90/Y PAND2X1_72/A POR2X1_317/B PAND2X1_313/a_16_344#
+ PAND2X1_313/m4_208_n4# PAND2X1_313/O PAND2X1_313/a_56_28# PAND2X1_313/CTRL2 PAND2X1_313/CTRL
+ PAND2X1_313/a_76_28# PAND2X1
XPAND2X1_346 VDD GND POR2X1_295/Y POR2X1_292/Y PAND2X1_346/Y PAND2X1_346/a_16_344#
+ POR2X1_481/m4_208_n4# PAND2X1_346/O PAND2X1_346/a_56_28# PAND2X1_346/CTRL2 PAND2X1_346/CTRL
+ PAND2X1_346/a_76_28# PAND2X1
XPAND2X1_335 VDD GND POR2X1_310/Y POR2X1_309/Y PAND2X1_337/A PAND2X1_335/a_16_344#
+ PAND2X1_335/m4_208_n4# PAND2X1_335/O PAND2X1_335/a_56_28# PAND2X1_335/CTRL2 PAND2X1_335/CTRL
+ PAND2X1_335/a_76_28# PAND2X1
XPAND2X1_324 VDD GND POR2X1_321/Y POR2X1_320/Y PAND2X1_324/Y PAND2X1_324/a_16_344#
+ PAND2X1_324/m4_208_n4# PAND2X1_324/O PAND2X1_324/a_56_28# PAND2X1_324/CTRL2 PAND2X1_324/CTRL
+ PAND2X1_324/a_76_28# PAND2X1
XPAND2X1_368 VDD GND POR2X1_270/Y PAND2X1_6/Y POR2X1_457/B PAND2X1_368/a_16_344# PAND2X1_368/m4_208_n4#
+ PAND2X1_368/O PAND2X1_368/a_56_28# PAND2X1_368/CTRL2 PAND2X1_368/CTRL PAND2X1_368/a_76_28#
+ PAND2X1
XPAND2X1_357 VDD GND PAND2X1_353/Y PAND2X1_352/Y PAND2X1_357/Y PAND2X1_357/a_16_344#
+ PAND2X1_357/m4_208_n4# PAND2X1_357/O PAND2X1_357/a_56_28# PAND2X1_357/CTRL2 PAND2X1_357/CTRL
+ PAND2X1_357/a_76_28# PAND2X1
XPAND2X1_379 VDD GND POR2X1_83/B POR2X1_13/A POR2X1_380/A PAND2X1_379/a_16_344# PAND2X1_379/m4_208_n4#
+ PAND2X1_379/O PAND2X1_379/a_56_28# PAND2X1_379/CTRL2 PAND2X1_379/CTRL PAND2X1_379/a_76_28#
+ PAND2X1
XPOR2X1_180 VDD GND POR2X1_180/B POR2X1_180/A POR2X1_180/Y POR2X1_180/m4_208_n4# POR2X1_180/O
+ POR2X1_180/CTRL2 POR2X1_180/a_16_28# POR2X1_180/CTRL POR2X1_180/a_76_344# POR2X1_180/a_56_344#
+ POR2X1
XPOR2X1_191 VDD GND POR2X1_191/B POR2X1_190/Y POR2X1_191/Y POR2X1_191/m4_208_n4# POR2X1_191/O
+ POR2X1_191/CTRL2 POR2X1_191/a_16_28# POR2X1_191/CTRL POR2X1_191/a_76_344# POR2X1_191/a_56_344#
+ POR2X1
XPAND2X1_110 VDD GND PAND2X1_94/A D_INPUT_0 PAND2X1_111/B PAND2X1_110/a_16_344# PAND2X1_110/m4_208_n4#
+ PAND2X1_110/O PAND2X1_110/a_56_28# PAND2X1_110/CTRL2 PAND2X1_110/CTRL PAND2X1_110/a_76_28#
+ PAND2X1
XPAND2X1_121 VDD GND POR2X1_666/A POR2X1_119/Y POR2X1_122/A PAND2X1_121/a_16_344#
+ PAND2X1_121/m4_208_n4# PAND2X1_121/O PAND2X1_121/a_56_28# PAND2X1_121/CTRL2 PAND2X1_121/CTRL
+ PAND2X1_121/a_76_28# PAND2X1
XPAND2X1_143 VDD GND PAND2X1_8/Y D_INPUT_1 POR2X1_502/A PAND2X1_143/a_16_344# PAND2X1_143/m4_208_n4#
+ PAND2X1_143/O PAND2X1_143/a_56_28# PAND2X1_143/CTRL2 PAND2X1_143/CTRL PAND2X1_143/a_76_28#
+ PAND2X1
XPAND2X1_132 VDD GND PAND2X1_96/B PAND2X1_90/Y POR2X1_137/B PAND2X1_132/a_16_344#
+ PAND2X1_132/m4_208_n4# PAND2X1_132/O PAND2X1_132/a_56_28# PAND2X1_132/CTRL2 PAND2X1_132/CTRL
+ PAND2X1_132/a_76_28# PAND2X1
XPAND2X1_154 VDD GND POR2X1_38/Y POR2X1_7/A PAND2X1_156/A PAND2X1_154/a_16_344# PAND2X1_154/m4_208_n4#
+ PAND2X1_154/O PAND2X1_154/a_56_28# PAND2X1_154/CTRL2 PAND2X1_154/CTRL PAND2X1_154/a_76_28#
+ PAND2X1
XPAND2X1_165 VDD GND PAND2X1_73/Y PAND2X1_52/B POR2X1_168/A PAND2X1_165/a_16_344#
+ PAND2X1_165/m4_208_n4# PAND2X1_165/O PAND2X1_165/a_56_28# PAND2X1_165/CTRL2 PAND2X1_165/CTRL
+ PAND2X1_165/a_76_28# PAND2X1
XPAND2X1_176 VDD GND PAND2X1_90/Y POR2X1_66/A POR2X1_180/B PAND2X1_176/a_16_344# PAND2X1_176/m4_208_n4#
+ PAND2X1_176/O PAND2X1_176/a_56_28# PAND2X1_176/CTRL2 PAND2X1_176/CTRL PAND2X1_176/a_76_28#
+ PAND2X1
XPAND2X1_187 VDD GND POR2X1_186/Y PAND2X1_41/B POR2X1_191/B PAND2X1_187/a_16_344#
+ POR2X1_191/m4_208_n4# PAND2X1_187/O PAND2X1_187/a_56_28# PAND2X1_187/CTRL2 PAND2X1_187/CTRL
+ PAND2X1_187/a_76_28# PAND2X1
XPAND2X1_198 VDD GND PAND2X1_197/Y POR2X1_57/Y PAND2X1_198/Y PAND2X1_198/a_16_344#
+ PAND2X1_198/m4_208_n4# PAND2X1_198/O PAND2X1_198/a_56_28# PAND2X1_198/CTRL2 PAND2X1_198/CTRL
+ PAND2X1_198/a_76_28# PAND2X1
XPOR2X1_702 VDD GND POR2X1_702/B POR2X1_702/A POR2X1_715/A POR2X1_702/m4_208_n4# POR2X1_702/O
+ POR2X1_702/CTRL2 POR2X1_702/a_16_28# POR2X1_702/CTRL POR2X1_702/a_76_344# POR2X1_702/a_56_344#
+ POR2X1
XPOR2X1_735 VDD GND POR2X1_573/A POR2X1_632/Y POR2X1_736/A POR2X1_735/m4_208_n4# POR2X1_735/O
+ POR2X1_735/CTRL2 POR2X1_735/a_16_28# POR2X1_735/CTRL POR2X1_735/a_76_344# POR2X1_735/a_56_344#
+ POR2X1
XPOR2X1_724 VDD GND POR2X1_724/B POR2X1_724/A POR2X1_732/B POR2X1_724/m4_208_n4# POR2X1_724/O
+ POR2X1_724/CTRL2 POR2X1_724/a_16_28# POR2X1_724/CTRL POR2X1_724/a_76_344# POR2X1_724/a_56_344#
+ POR2X1
XPOR2X1_713 VDD GND POR2X1_713/B POR2X1_713/A POR2X1_713/Y POR2X1_713/m4_208_n4# POR2X1_713/O
+ POR2X1_713/CTRL2 POR2X1_713/a_16_28# POR2X1_713/CTRL POR2X1_713/a_76_344# POR2X1_713/a_56_344#
+ POR2X1
XPOR2X1_757 VDD GND POR2X1_57/A POR2X1_757/A POR2X1_757/Y POR2X1_755/m4_208_n4# POR2X1_757/O
+ POR2X1_757/CTRL2 POR2X1_757/a_16_28# POR2X1_757/CTRL POR2X1_757/a_76_344# POR2X1_757/a_56_344#
+ POR2X1
XPOR2X1_768 VDD GND POR2X1_113/B POR2X1_768/A POR2X1_768/Y POR2X1_768/m4_208_n4# POR2X1_768/O
+ POR2X1_768/CTRL2 POR2X1_768/a_16_28# POR2X1_768/CTRL POR2X1_768/a_76_344# POR2X1_768/a_56_344#
+ POR2X1
XPOR2X1_746 VDD GND POR2X1_73/Y POR2X1_416/B POR2X1_746/Y POR2X1_746/m4_208_n4# POR2X1_746/O
+ POR2X1_746/CTRL2 POR2X1_746/a_16_28# POR2X1_746/CTRL POR2X1_746/a_76_344# POR2X1_746/a_56_344#
+ POR2X1
XPOR2X1_779 VDD GND POR2X1_513/B POR2X1_779/A POR2X1_783/B POR2X1_779/m4_208_n4# POR2X1_779/O
+ POR2X1_779/CTRL2 POR2X1_779/a_16_28# POR2X1_779/CTRL POR2X1_779/a_76_344# POR2X1_779/a_56_344#
+ POR2X1
XPAND2X1_709 VDD GND POR2X1_748/A POR2X1_698/Y PAND2X1_711/A PAND2X1_709/a_16_344#
+ POR2X1_698/m4_208_n4# PAND2X1_709/O PAND2X1_709/a_56_28# PAND2X1_709/CTRL2 PAND2X1_709/CTRL
+ PAND2X1_709/a_76_28# PAND2X1
XPOR2X1_6 VDD GND POR2X1_4/Y POR2X1_5/Y POR2X1_7/A POR2X1_6/m4_208_n4# POR2X1_6/O
+ POR2X1_6/CTRL2 POR2X1_6/a_16_28# POR2X1_6/CTRL POR2X1_6/a_76_344# POR2X1_6/a_56_344#
+ POR2X1
XPOR2X1_510 VDD GND POR2X1_510/B POR2X1_510/A POR2X1_510/Y PAND2X1_52/m4_208_n4# POR2X1_510/O
+ POR2X1_510/CTRL2 POR2X1_510/a_16_28# POR2X1_510/CTRL POR2X1_510/a_76_344# POR2X1_510/a_56_344#
+ POR2X1
XPOR2X1_521 VDD GND POR2X1_20/B POR2X1_49/Y POR2X1_521/Y POR2X1_521/m4_208_n4# POR2X1_521/O
+ POR2X1_521/CTRL2 POR2X1_521/a_16_28# POR2X1_521/CTRL POR2X1_521/a_76_344# POR2X1_521/a_56_344#
+ POR2X1
XPOR2X1_543 VDD GND POR2X1_445/A POR2X1_543/A POR2X1_552/A POR2X1_543/m4_208_n4# POR2X1_543/O
+ POR2X1_543/CTRL2 POR2X1_543/a_16_28# POR2X1_543/CTRL POR2X1_543/a_76_344# POR2X1_543/a_56_344#
+ POR2X1
XPOR2X1_532 VDD GND POR2X1_590/A POR2X1_532/A POR2X1_532/Y POR2X1_532/m4_208_n4# POR2X1_532/O
+ POR2X1_532/CTRL2 POR2X1_532/a_16_28# POR2X1_532/CTRL POR2X1_532/a_76_344# POR2X1_532/a_56_344#
+ POR2X1
XPOR2X1_565 VDD GND POR2X1_565/B POR2X1_550/Y POR2X1_569/A POR2X1_565/m4_208_n4# POR2X1_565/O
+ POR2X1_565/CTRL2 POR2X1_565/a_16_28# POR2X1_565/CTRL POR2X1_565/a_76_344# POR2X1_565/a_56_344#
+ POR2X1
XPOR2X1_576 VDD GND POR2X1_571/Y POR2X1_572/Y POR2X1_576/Y POR2X1_576/m4_208_n4# POR2X1_576/O
+ POR2X1_576/CTRL2 POR2X1_576/a_16_28# POR2X1_576/CTRL POR2X1_576/a_76_344# POR2X1_576/a_56_344#
+ POR2X1
XPOR2X1_554 VDD GND POR2X1_554/B POR2X1_140/B POR2X1_554/Y POR2X1_554/m4_208_n4# POR2X1_554/O
+ POR2X1_554/CTRL2 POR2X1_554/a_16_28# POR2X1_554/CTRL POR2X1_554/a_76_344# POR2X1_554/a_56_344#
+ POR2X1
XPOR2X1_587 VDD GND INPUT_7 POR2X1_51/B POR2X1_587/Y POR2X1_587/m4_208_n4# POR2X1_587/O
+ POR2X1_587/CTRL2 POR2X1_587/a_16_28# POR2X1_587/CTRL POR2X1_587/a_76_344# POR2X1_587/a_56_344#
+ POR2X1
XPOR2X1_598 VDD GND PAND2X1_48/A POR2X1_294/A POR2X1_828/A POR2X1_598/m4_208_n4# POR2X1_598/O
+ POR2X1_598/CTRL2 POR2X1_598/a_16_28# POR2X1_598/CTRL POR2X1_598/a_76_344# POR2X1_598/a_56_344#
+ POR2X1
XPAND2X1_517 VDD GND POR2X1_264/Y PAND2X1_32/B POR2X1_559/B PAND2X1_517/a_16_344#
+ PAND2X1_517/m4_208_n4# PAND2X1_517/O PAND2X1_517/a_56_28# PAND2X1_517/CTRL2 PAND2X1_517/CTRL
+ PAND2X1_517/a_76_28# PAND2X1
XPAND2X1_506 VDD GND POR2X1_419/Y POR2X1_239/Y PAND2X1_506/Y PAND2X1_506/a_16_344#
+ PAND2X1_506/m4_208_n4# PAND2X1_506/O PAND2X1_506/a_56_28# PAND2X1_506/CTRL2 PAND2X1_506/CTRL
+ PAND2X1_506/a_76_28# PAND2X1
XPAND2X1_528 VDD GND PAND2X1_57/B PAND2X1_6/Y POR2X1_620/B PAND2X1_528/a_16_344# PAND2X1_528/m4_208_n4#
+ PAND2X1_528/O PAND2X1_528/a_56_28# PAND2X1_528/CTRL2 PAND2X1_528/CTRL PAND2X1_528/a_76_28#
+ PAND2X1
XPAND2X1_539 VDD GND PAND2X1_539/B PAND2X1_643/A PAND2X1_539/Y PAND2X1_539/a_16_344#
+ PAND2X1_539/m4_208_n4# PAND2X1_539/O PAND2X1_539/a_56_28# PAND2X1_539/CTRL2 PAND2X1_539/CTRL
+ PAND2X1_539/a_76_28# PAND2X1
XPOR2X1_340 VDD GND PAND2X1_88/Y POR2X1_509/B POR2X1_350/B POR2X1_340/m4_208_n4# POR2X1_340/O
+ POR2X1_340/CTRL2 POR2X1_340/a_16_28# POR2X1_340/CTRL POR2X1_340/a_76_344# POR2X1_340/a_56_344#
+ POR2X1
XPOR2X1_351 VDD GND POR2X1_351/B POR2X1_339/Y POR2X1_351/Y POR2X1_351/m4_208_n4# POR2X1_351/O
+ POR2X1_351/CTRL2 POR2X1_351/a_16_28# POR2X1_351/CTRL POR2X1_351/a_76_344# POR2X1_351/a_56_344#
+ POR2X1
XPOR2X1_362 VDD GND POR2X1_362/B POR2X1_362/A POR2X1_362/Y POR2X1_362/m4_208_n4# POR2X1_362/O
+ POR2X1_362/CTRL2 POR2X1_362/a_16_28# POR2X1_362/CTRL POR2X1_362/a_76_344# POR2X1_362/a_56_344#
+ POR2X1
XPOR2X1_395 VDD GND POR2X1_60/A POR2X1_411/B POR2X1_395/Y POR2X1_395/m4_208_n4# POR2X1_395/O
+ POR2X1_395/CTRL2 POR2X1_395/a_16_28# POR2X1_395/CTRL POR2X1_395/a_76_344# POR2X1_395/a_56_344#
+ POR2X1
XPOR2X1_384 VDD GND POR2X1_40/Y POR2X1_384/A POR2X1_384/Y POR2X1_384/m4_208_n4# POR2X1_384/O
+ POR2X1_384/CTRL2 POR2X1_384/a_16_28# POR2X1_384/CTRL POR2X1_384/a_76_344# POR2X1_384/a_56_344#
+ POR2X1
XPOR2X1_373 VDD GND POR2X1_83/B POR2X1_77/Y POR2X1_373/Y POR2X1_373/m4_208_n4# POR2X1_373/O
+ POR2X1_373/CTRL2 POR2X1_373/a_16_28# POR2X1_373/CTRL POR2X1_373/a_76_344# POR2X1_373/a_56_344#
+ POR2X1
XPAND2X1_303 VDD GND PAND2X1_303/B PAND2X1_716/B PAND2X1_303/Y PAND2X1_303/a_16_344#
+ PAND2X1_303/m4_208_n4# PAND2X1_303/O PAND2X1_303/a_56_28# PAND2X1_303/CTRL2 PAND2X1_303/CTRL
+ PAND2X1_303/a_76_28# PAND2X1
XPAND2X1_314 VDD GND PAND2X1_65/B POR2X1_78/B POR2X1_317/A PAND2X1_314/a_16_344# PAND2X1_314/m4_208_n4#
+ PAND2X1_314/O PAND2X1_314/a_56_28# PAND2X1_314/CTRL2 PAND2X1_314/CTRL PAND2X1_314/a_76_28#
+ PAND2X1
XPAND2X1_336 VDD GND POR2X1_312/Y POR2X1_311/Y PAND2X1_336/Y PAND2X1_336/a_16_344#
+ PAND2X1_336/m4_208_n4# PAND2X1_336/O PAND2X1_336/a_56_28# PAND2X1_336/CTRL2 PAND2X1_336/CTRL
+ PAND2X1_336/a_76_28# PAND2X1
XPAND2X1_325 VDD GND POR2X1_323/Y POR2X1_322/Y PAND2X1_326/B PAND2X1_325/a_16_344#
+ PAND2X1_565/m4_208_n4# PAND2X1_325/O PAND2X1_325/a_56_28# PAND2X1_325/CTRL2 PAND2X1_325/CTRL
+ PAND2X1_325/a_76_28# PAND2X1
XPAND2X1_358 VDD GND PAND2X1_351/Y PAND2X1_358/A PAND2X1_364/B PAND2X1_358/a_16_344#
+ PAND2X1_358/m4_208_n4# PAND2X1_358/O PAND2X1_358/a_56_28# PAND2X1_358/CTRL2 PAND2X1_358/CTRL
+ PAND2X1_358/a_76_28# PAND2X1
XPAND2X1_369 VDD GND POR2X1_121/B PAND2X1_58/A POR2X1_543/A PAND2X1_369/a_16_344#
+ PAND2X1_369/m4_208_n4# PAND2X1_369/O PAND2X1_369/a_56_28# PAND2X1_369/CTRL2 PAND2X1_369/CTRL
+ PAND2X1_369/a_76_28# PAND2X1
XPAND2X1_347 VDD GND PAND2X1_346/Y POR2X1_297/Y PAND2X1_347/Y PAND2X1_347/a_16_344#
+ PAND2X1_347/m4_208_n4# PAND2X1_347/O PAND2X1_347/a_56_28# PAND2X1_347/CTRL2 PAND2X1_347/CTRL
+ PAND2X1_347/a_76_28# PAND2X1
XPOR2X1_170 VDD GND POR2X1_170/B POR2X1_169/Y POR2X1_566/B POR2X1_170/m4_208_n4# POR2X1_170/O
+ POR2X1_170/CTRL2 POR2X1_170/a_16_28# POR2X1_170/CTRL POR2X1_170/a_76_344# POR2X1_170/a_56_344#
+ POR2X1
XPOR2X1_192 VDD GND POR2X1_192/B POR2X1_191/Y POR2X1_192/Y POR2X1_580/m4_208_n4# POR2X1_192/O
+ POR2X1_192/CTRL2 POR2X1_192/a_16_28# POR2X1_192/CTRL POR2X1_192/a_76_344# POR2X1_192/a_56_344#
+ POR2X1
XPOR2X1_181 VDD GND POR2X1_181/B POR2X1_181/A POR2X1_181/Y POR2X1_181/m4_208_n4# POR2X1_181/O
+ POR2X1_181/CTRL2 POR2X1_181/a_16_28# POR2X1_181/CTRL POR2X1_181/a_76_344# POR2X1_181/a_56_344#
+ POR2X1
XPAND2X1_111 VDD GND PAND2X1_111/B PAND2X1_32/B POR2X1_332/B PAND2X1_111/a_16_344#
+ PAND2X1_111/m4_208_n4# PAND2X1_111/O PAND2X1_111/a_56_28# PAND2X1_111/CTRL2 PAND2X1_111/CTRL
+ PAND2X1_111/a_76_28# PAND2X1
XPAND2X1_100 VDD GND POR2X1_88/Y POR2X1_86/Y PAND2X1_101/B PAND2X1_100/a_16_344# PAND2X1_100/m4_208_n4#
+ PAND2X1_100/O PAND2X1_100/a_56_28# PAND2X1_100/CTRL2 PAND2X1_100/CTRL PAND2X1_100/a_76_28#
+ PAND2X1
XPAND2X1_122 VDD GND POR2X1_121/Y PAND2X1_57/B POR2X1_124/B PAND2X1_122/a_16_344#
+ PAND2X1_122/m4_208_n4# PAND2X1_122/O PAND2X1_122/a_56_28# PAND2X1_122/CTRL2 PAND2X1_122/CTRL
+ PAND2X1_122/a_76_28# PAND2X1
XPAND2X1_144 VDD GND POR2X1_502/A PAND2X1_60/B POR2X1_147/A PAND2X1_144/a_16_344#
+ PAND2X1_144/m4_208_n4# PAND2X1_144/O PAND2X1_144/a_56_28# PAND2X1_144/CTRL2 PAND2X1_144/CTRL
+ PAND2X1_144/a_76_28# PAND2X1
XPAND2X1_133 VDD GND POR2X1_29/A PAND2X1_8/Y POR2X1_614/A PAND2X1_133/a_16_344# PAND2X1_133/m4_208_n4#
+ PAND2X1_133/O PAND2X1_133/a_56_28# PAND2X1_133/CTRL2 PAND2X1_133/CTRL PAND2X1_133/a_76_28#
+ PAND2X1
XPAND2X1_166 VDD GND PAND2X1_41/B POR2X1_78/B POR2X1_169/B PAND2X1_166/a_16_344# PAND2X1_166/m4_208_n4#
+ PAND2X1_166/O PAND2X1_166/a_56_28# PAND2X1_166/CTRL2 PAND2X1_166/CTRL PAND2X1_166/a_76_28#
+ PAND2X1
XPAND2X1_188 VDD GND POR2X1_816/A POR2X1_38/Y POR2X1_498/A PAND2X1_188/a_16_344# PAND2X1_188/m4_208_n4#
+ PAND2X1_188/O PAND2X1_188/a_56_28# PAND2X1_188/CTRL2 PAND2X1_188/CTRL PAND2X1_188/a_76_28#
+ PAND2X1
XPAND2X1_177 VDD GND PAND2X1_72/A POR2X1_68/A POR2X1_180/A PAND2X1_177/a_16_344# POR2X1_544/m4_208_n4#
+ PAND2X1_177/O PAND2X1_177/a_56_28# PAND2X1_177/CTRL2 PAND2X1_177/CTRL PAND2X1_177/a_76_28#
+ PAND2X1
XPAND2X1_155 VDD GND POR2X1_153/Y POR2X1_49/Y PAND2X1_156/B PAND2X1_155/a_16_344#
+ PAND2X1_155/m4_208_n4# PAND2X1_155/O PAND2X1_155/a_56_28# PAND2X1_155/CTRL2 PAND2X1_155/CTRL
+ PAND2X1_155/a_76_28# PAND2X1
XPAND2X1_199 VDD GND PAND2X1_199/B PAND2X1_199/A PAND2X1_207/A PAND2X1_199/a_16_344#
+ PAND2X1_199/m4_208_n4# PAND2X1_199/O PAND2X1_199/a_56_28# PAND2X1_199/CTRL2 PAND2X1_199/CTRL
+ PAND2X1_199/a_76_28# PAND2X1
XPOR2X1_714 VDD GND POR2X1_703/Y POR2X1_704/Y POR2X1_724/B POR2X1_714/m4_208_n4# POR2X1_714/O
+ POR2X1_714/CTRL2 POR2X1_714/a_16_28# POR2X1_714/CTRL POR2X1_714/a_76_344# POR2X1_714/a_56_344#
+ POR2X1
XPOR2X1_703 VDD GND POR2X1_169/A POR2X1_703/A POR2X1_703/Y POR2X1_703/m4_208_n4# POR2X1_703/O
+ POR2X1_703/CTRL2 POR2X1_703/a_16_28# POR2X1_703/CTRL POR2X1_703/a_76_344# POR2X1_703/a_56_344#
+ POR2X1
XPOR2X1_725 VDD GND POR2X1_712/Y POR2X1_713/Y POR2X1_725/Y POR2X1_725/m4_208_n4# POR2X1_725/O
+ POR2X1_725/CTRL2 POR2X1_725/a_16_28# POR2X1_725/CTRL POR2X1_725/a_76_344# POR2X1_725/a_56_344#
+ POR2X1
XPOR2X1_736 VDD GND POR2X1_675/Y POR2X1_736/A POR2X1_741/B POR2X1_741/m4_208_n4# POR2X1_736/O
+ POR2X1_736/CTRL2 POR2X1_736/a_16_28# POR2X1_736/CTRL POR2X1_736/a_76_344# POR2X1_736/a_56_344#
+ POR2X1
XPOR2X1_769 VDD GND POR2X1_769/B POR2X1_769/A POR2X1_769/Y POR2X1_769/m4_208_n4# POR2X1_769/O
+ POR2X1_769/CTRL2 POR2X1_769/a_16_28# POR2X1_769/CTRL POR2X1_769/a_76_344# POR2X1_769/a_56_344#
+ POR2X1
XPOR2X1_747 VDD GND POR2X1_48/A POR2X1_49/Y POR2X1_747/Y POR2X1_747/m4_208_n4# POR2X1_747/O
+ POR2X1_747/CTRL2 POR2X1_747/a_16_28# POR2X1_747/CTRL POR2X1_747/a_76_344# POR2X1_747/a_56_344#
+ POR2X1
XPOR2X1_758 VDD GND PAND2X1_41/B PAND2X1_96/B POR2X1_758/Y POR2X1_758/m4_208_n4# POR2X1_758/O
+ POR2X1_758/CTRL2 POR2X1_758/a_16_28# POR2X1_758/CTRL POR2X1_758/a_76_344# POR2X1_758/a_56_344#
+ POR2X1
XPOR2X1_7 VDD GND POR2X1_7/B POR2X1_7/A POR2X1_7/Y POR2X1_7/m4_208_n4# POR2X1_7/O
+ POR2X1_7/CTRL2 POR2X1_7/a_16_28# POR2X1_7/CTRL POR2X1_7/a_76_344# POR2X1_7/a_56_344#
+ POR2X1
XPOR2X1_500 VDD GND POR2X1_844/B POR2X1_500/A POR2X1_500/Y POR2X1_500/m4_208_n4# POR2X1_500/O
+ POR2X1_500/CTRL2 POR2X1_500/a_16_28# POR2X1_500/CTRL POR2X1_500/a_76_344# POR2X1_500/a_56_344#
+ POR2X1
XPOR2X1_511 VDD GND POR2X1_32/A POR2X1_46/Y POR2X1_511/Y POR2X1_511/m4_208_n4# POR2X1_511/O
+ POR2X1_511/CTRL2 POR2X1_511/a_16_28# POR2X1_511/CTRL POR2X1_511/a_76_344# POR2X1_511/a_56_344#
+ POR2X1
XPOR2X1_533 VDD GND POR2X1_96/A POR2X1_533/A POR2X1_533/Y POR2X1_533/m4_208_n4# POR2X1_533/O
+ POR2X1_533/CTRL2 POR2X1_533/a_16_28# POR2X1_533/CTRL POR2X1_533/a_76_344# POR2X1_533/a_56_344#
+ POR2X1
XPOR2X1_522 VDD GND POR2X1_43/B POR2X1_102/Y POR2X1_522/Y POR2X1_522/m4_208_n4# POR2X1_522/O
+ POR2X1_522/CTRL2 POR2X1_522/a_16_28# POR2X1_522/CTRL POR2X1_522/a_76_344# POR2X1_522/a_56_344#
+ POR2X1
XPOR2X1_544 VDD GND POR2X1_544/B POR2X1_544/A POR2X1_544/Y POR2X1_544/m4_208_n4# POR2X1_544/O
+ POR2X1_544/CTRL2 POR2X1_544/a_16_28# POR2X1_544/CTRL POR2X1_544/a_76_344# POR2X1_544/a_56_344#
+ POR2X1
XPOR2X1_566 VDD GND POR2X1_566/B POR2X1_566/A POR2X1_568/B POR2X1_566/m4_208_n4# POR2X1_566/O
+ POR2X1_566/CTRL2 POR2X1_566/a_16_28# POR2X1_566/CTRL POR2X1_566/a_76_344# POR2X1_566/a_56_344#
+ POR2X1
XPOR2X1_555 VDD GND POR2X1_555/B POR2X1_555/A POR2X1_562/B POR2X1_555/m4_208_n4# POR2X1_555/O
+ POR2X1_555/CTRL2 POR2X1_555/a_16_28# POR2X1_555/CTRL POR2X1_555/a_76_344# POR2X1_555/a_56_344#
+ POR2X1
XPOR2X1_577 VDD GND POR2X1_569/Y POR2X1_570/Y POR2X1_577/Y POR2X1_577/m4_208_n4# POR2X1_577/O
+ POR2X1_577/CTRL2 POR2X1_577/a_16_28# POR2X1_577/CTRL POR2X1_577/a_76_344# POR2X1_577/a_56_344#
+ POR2X1
XPOR2X1_599 VDD GND POR2X1_39/B POR2X1_599/A POR2X1_761/A POR2X1_599/m4_208_n4# POR2X1_599/O
+ POR2X1_599/CTRL2 POR2X1_599/a_16_28# POR2X1_599/CTRL POR2X1_599/a_76_344# POR2X1_599/a_56_344#
+ POR2X1
XPOR2X1_588 VDD GND POR2X1_376/B POR2X1_587/Y POR2X1_588/Y POR2X1_588/m4_208_n4# POR2X1_588/O
+ POR2X1_588/CTRL2 POR2X1_588/a_16_28# POR2X1_588/CTRL POR2X1_588/a_76_344# POR2X1_588/a_56_344#
+ POR2X1
XPAND2X1_518 VDD GND PAND2X1_73/Y PAND2X1_65/B POR2X1_520/B PAND2X1_518/a_16_344#
+ PAND2X1_518/m4_208_n4# PAND2X1_518/O PAND2X1_518/a_56_28# PAND2X1_518/CTRL2 PAND2X1_518/CTRL
+ PAND2X1_518/a_76_28# PAND2X1
XPAND2X1_507 VDD GND POR2X1_505/Y POR2X1_504/Y PAND2X1_508/B PAND2X1_507/a_16_344#
+ PAND2X1_507/m4_208_n4# PAND2X1_507/O PAND2X1_507/a_56_28# PAND2X1_507/CTRL2 PAND2X1_507/CTRL
+ PAND2X1_507/a_76_28# PAND2X1
XPAND2X1_529 VDD GND POR2X1_66/A INPUT_3 POR2X1_548/B PAND2X1_529/a_16_344# PAND2X1_529/m4_208_n4#
+ PAND2X1_529/O PAND2X1_529/a_56_28# PAND2X1_529/CTRL2 PAND2X1_529/CTRL PAND2X1_529/a_76_28#
+ PAND2X1
XPOR2X1_341 VDD GND POR2X1_228/Y POR2X1_341/A POR2X1_341/Y POR2X1_341/m4_208_n4# POR2X1_341/O
+ POR2X1_341/CTRL2 POR2X1_341/a_16_28# POR2X1_341/CTRL POR2X1_341/a_76_344# POR2X1_341/a_56_344#
+ POR2X1
XPOR2X1_352 VDD GND POR2X1_212/B POR2X1_337/Y POR2X1_357/B POR2X1_352/m4_208_n4# POR2X1_352/O
+ POR2X1_352/CTRL2 POR2X1_352/a_16_28# POR2X1_352/CTRL POR2X1_352/a_76_344# POR2X1_352/a_56_344#
+ POR2X1
XPOR2X1_330 VDD GND PAND2X1_52/B PAND2X1_72/A POR2X1_330/Y POR2X1_330/m4_208_n4# POR2X1_330/O
+ POR2X1_330/CTRL2 POR2X1_330/a_16_28# POR2X1_330/CTRL POR2X1_330/a_76_344# POR2X1_330/a_56_344#
+ POR2X1
XPOR2X1_363 VDD GND POR2X1_359/Y POR2X1_363/A POR2X1_366/A POR2X1_205/m4_208_n4# POR2X1_363/O
+ POR2X1_363/CTRL2 POR2X1_363/a_16_28# POR2X1_363/CTRL POR2X1_363/a_76_344# POR2X1_363/a_56_344#
+ POR2X1
XPOR2X1_385 VDD GND POR2X1_83/B POR2X1_411/B POR2X1_385/Y POR2X1_385/m4_208_n4# POR2X1_385/O
+ POR2X1_385/CTRL2 POR2X1_385/a_16_28# POR2X1_385/CTRL POR2X1_385/a_76_344# POR2X1_385/a_56_344#
+ POR2X1
XPOR2X1_374 VDD GND POR2X1_325/B POR2X1_544/B POR2X1_717/B POR2X1_374/m4_208_n4# POR2X1_374/O
+ POR2X1_374/CTRL2 POR2X1_374/a_16_28# POR2X1_374/CTRL POR2X1_374/a_76_344# POR2X1_374/a_56_344#
+ POR2X1
XPOR2X1_396 VDD GND POR2X1_23/Y POR2X1_39/B POR2X1_396/Y POR2X1_396/m4_208_n4# POR2X1_396/O
+ POR2X1_396/CTRL2 POR2X1_396/a_16_28# POR2X1_396/CTRL POR2X1_396/a_76_344# POR2X1_396/a_56_344#
+ POR2X1
XPAND2X1_315 VDD GND POR2X1_614/A PAND2X1_32/B POR2X1_445/A PAND2X1_315/a_16_344#
+ PAND2X1_315/m4_208_n4# PAND2X1_315/O PAND2X1_315/a_56_28# PAND2X1_315/CTRL2 PAND2X1_315/CTRL
+ PAND2X1_315/a_76_28# PAND2X1
XPAND2X1_337 VDD GND PAND2X1_336/Y PAND2X1_337/A PAND2X1_352/B PAND2X1_337/a_16_344#
+ PAND2X1_337/m4_208_n4# PAND2X1_337/O PAND2X1_337/a_56_28# PAND2X1_337/CTRL2 PAND2X1_337/CTRL
+ PAND2X1_337/a_76_28# PAND2X1
XPAND2X1_304 VDD GND POR2X1_383/A PAND2X1_56/A POR2X1_307/B PAND2X1_304/a_16_344#
+ PAND2X1_304/m4_208_n4# PAND2X1_304/O PAND2X1_304/a_56_28# PAND2X1_304/CTRL2 PAND2X1_304/CTRL
+ PAND2X1_304/a_76_28# PAND2X1
XPAND2X1_326 VDD GND PAND2X1_326/B PAND2X1_324/Y PAND2X1_854/A PAND2X1_326/a_16_344#
+ PAND2X1_326/m4_208_n4# PAND2X1_326/O PAND2X1_326/a_56_28# PAND2X1_326/CTRL2 PAND2X1_326/CTRL
+ PAND2X1_326/a_76_28# PAND2X1
XPAND2X1_359 VDD GND PAND2X1_359/B PAND2X1_348/Y PAND2X1_359/Y PAND2X1_359/a_16_344#
+ PAND2X1_359/m4_208_n4# PAND2X1_359/O PAND2X1_359/a_56_28# PAND2X1_359/CTRL2 PAND2X1_359/CTRL
+ PAND2X1_359/a_76_28# PAND2X1
XPAND2X1_348 VDD GND PAND2X1_345/Y PAND2X1_348/A PAND2X1_348/Y PAND2X1_348/a_16_344#
+ PAND2X1_348/m4_208_n4# PAND2X1_348/O PAND2X1_348/a_56_28# PAND2X1_348/CTRL2 PAND2X1_348/CTRL
+ PAND2X1_348/a_76_28# PAND2X1
XPAND2X1_860 VDD GND PAND2X1_474/A PAND2X1_860/A PAND2X1_861/B PAND2X1_860/a_16_344#
+ PAND2X1_860/m4_208_n4# PAND2X1_860/O PAND2X1_860/a_56_28# PAND2X1_860/CTRL2 PAND2X1_860/CTRL
+ PAND2X1_860/a_76_28# PAND2X1
XPOR2X1_160 VDD GND PAND2X1_23/Y POR2X1_532/A POR2X1_162/B POR2X1_356/m4_208_n4# POR2X1_160/O
+ POR2X1_160/CTRL2 POR2X1_160/a_16_28# POR2X1_160/CTRL POR2X1_160/a_76_344# POR2X1_160/a_56_344#
+ POR2X1
XPOR2X1_193 VDD GND PAND2X1_7/Y POR2X1_193/A POR2X1_193/Y POR2X1_193/m4_208_n4# POR2X1_193/O
+ POR2X1_193/CTRL2 POR2X1_193/a_16_28# POR2X1_193/CTRL POR2X1_193/a_76_344# POR2X1_193/a_56_344#
+ POR2X1
XPOR2X1_171 VDD GND POR2X1_23/Y POR2X1_40/Y POR2X1_171/Y POR2X1_171/m4_208_n4# POR2X1_171/O
+ POR2X1_171/CTRL2 POR2X1_171/a_16_28# POR2X1_171/CTRL POR2X1_171/a_76_344# POR2X1_171/a_56_344#
+ POR2X1
XPOR2X1_182 VDD GND POR2X1_180/Y POR2X1_181/Y POR2X1_212/B POR2X1_182/m4_208_n4# POR2X1_182/O
+ POR2X1_182/CTRL2 POR2X1_182/a_16_28# POR2X1_182/CTRL POR2X1_182/a_76_344# POR2X1_182/a_56_344#
+ POR2X1
XPAND2X1_101 VDD GND PAND2X1_101/B PAND2X1_99/Y PAND2X1_656/A PAND2X1_101/a_16_344#
+ POR2X1_86/m4_208_n4# PAND2X1_101/O PAND2X1_101/a_56_28# PAND2X1_101/CTRL2 PAND2X1_101/CTRL
+ PAND2X1_101/a_76_28# PAND2X1
XPAND2X1_112 VDD GND POR2X1_111/Y POR2X1_109/Y PAND2X1_115/B PAND2X1_112/a_16_344#
+ PAND2X1_112/m4_208_n4# PAND2X1_112/O PAND2X1_112/a_56_28# PAND2X1_112/CTRL2 PAND2X1_112/CTRL
+ PAND2X1_112/a_76_28# PAND2X1
XPAND2X1_134 VDD GND POR2X1_614/A PAND2X1_96/B POR2X1_768/A PAND2X1_134/a_16_344#
+ PAND2X1_107/m4_208_n4# PAND2X1_134/O PAND2X1_134/a_56_28# PAND2X1_134/CTRL2 PAND2X1_134/CTRL
+ PAND2X1_134/a_76_28# PAND2X1
XPAND2X1_145 VDD GND POR2X1_78/A PAND2X1_52/B POR2X1_148/B PAND2X1_145/a_16_344# PAND2X1_146/m4_208_n4#
+ PAND2X1_145/O PAND2X1_145/a_56_28# PAND2X1_145/CTRL2 PAND2X1_145/CTRL PAND2X1_145/a_76_28#
+ PAND2X1
XPAND2X1_123 VDD GND POR2X1_118/Y POR2X1_117/Y PAND2X1_123/Y PAND2X1_123/a_16_344#
+ POR2X1_117/m4_208_n4# PAND2X1_123/O PAND2X1_123/a_56_28# PAND2X1_123/CTRL2 PAND2X1_123/CTRL
+ PAND2X1_123/a_76_28# PAND2X1
XPAND2X1_167 VDD GND POR2X1_750/B PAND2X1_65/B POR2X1_169/A PAND2X1_167/a_16_344#
+ PAND2X1_167/m4_208_n4# PAND2X1_167/O PAND2X1_167/a_56_28# PAND2X1_167/CTRL2 PAND2X1_167/CTRL
+ PAND2X1_167/a_76_28# PAND2X1
XPAND2X1_178 VDD GND POR2X1_260/A PAND2X1_55/Y POR2X1_181/B PAND2X1_178/a_16_344#
+ PAND2X1_178/m4_208_n4# PAND2X1_178/O PAND2X1_178/a_56_28# PAND2X1_178/CTRL2 PAND2X1_178/CTRL
+ PAND2X1_178/a_76_28# PAND2X1
XPAND2X1_156 VDD GND PAND2X1_156/B PAND2X1_156/A POR2X1_158/B PAND2X1_156/a_16_344#
+ PAND2X1_156/m4_208_n4# PAND2X1_156/O PAND2X1_156/a_56_28# PAND2X1_156/CTRL2 PAND2X1_156/CTRL
+ PAND2X1_156/a_76_28# PAND2X1
XPAND2X1_189 VDD GND POR2X1_188/Y PAND2X1_96/B POR2X1_192/B PAND2X1_189/a_16_344#
+ PAND2X1_189/m4_208_n4# PAND2X1_189/O PAND2X1_189/a_56_28# PAND2X1_189/CTRL2 PAND2X1_189/CTRL
+ PAND2X1_189/a_76_28# PAND2X1
XPAND2X1_690 VDD GND POR2X1_634/A D_INPUT_0 POR2X1_691/A PAND2X1_690/a_16_344# PAND2X1_690/m4_208_n4#
+ PAND2X1_690/O PAND2X1_690/a_56_28# PAND2X1_690/CTRL2 PAND2X1_690/CTRL PAND2X1_690/a_76_28#
+ PAND2X1
XPOR2X1_715 VDD GND POR2X1_112/Y POR2X1_715/A POR2X1_724/A POR2X1_715/m4_208_n4# POR2X1_715/O
+ POR2X1_715/CTRL2 POR2X1_715/a_16_28# POR2X1_715/CTRL POR2X1_715/a_76_344# POR2X1_715/a_56_344#
+ POR2X1
XPOR2X1_704 VDD GND POR2X1_317/B POR2X1_446/B POR2X1_704/Y POR2X1_704/m4_208_n4# POR2X1_704/O
+ POR2X1_704/CTRL2 POR2X1_704/a_16_28# POR2X1_704/CTRL POR2X1_704/a_76_344# POR2X1_704/a_56_344#
+ POR2X1
XPOR2X1_726 VDD GND POR2X1_209/A POR2X1_711/Y POR2X1_726/Y POR2X1_726/m4_208_n4# POR2X1_726/O
+ POR2X1_726/CTRL2 POR2X1_726/a_16_28# POR2X1_726/CTRL POR2X1_726/a_76_344# POR2X1_726/a_56_344#
+ POR2X1
XPOR2X1_759 VDD GND POR2X1_236/Y POR2X1_759/A POR2X1_759/Y POR2X1_759/m4_208_n4# POR2X1_759/O
+ POR2X1_759/CTRL2 POR2X1_759/a_16_28# POR2X1_759/CTRL POR2X1_759/a_76_344# POR2X1_759/a_56_344#
+ POR2X1
XPOR2X1_748 VDD GND POR2X1_4/Y POR2X1_748/A POR2X1_748/Y POR2X1_748/m4_208_n4# POR2X1_748/O
+ POR2X1_748/CTRL2 POR2X1_748/a_16_28# POR2X1_748/CTRL POR2X1_748/a_76_344# POR2X1_748/a_56_344#
+ POR2X1
XPOR2X1_737 VDD GND POR2X1_733/Y POR2X1_737/A POR2X1_741/A POR2X1_737/m4_208_n4# POR2X1_737/O
+ POR2X1_737/CTRL2 POR2X1_737/a_16_28# POR2X1_737/CTRL POR2X1_737/a_76_344# POR2X1_737/a_56_344#
+ POR2X1
XPOR2X1_8 VDD GND D_INPUT_2 INPUT_3 POR2X1_8/Y POR2X1_8/m4_208_n4# POR2X1_8/O POR2X1_8/CTRL2
+ POR2X1_8/a_16_28# POR2X1_8/CTRL POR2X1_8/a_76_344# POR2X1_8/a_56_344# POR2X1
XPOR2X1_501 VDD GND POR2X1_501/B POR2X1_500/Y POR2X1_573/A POR2X1_501/m4_208_n4# POR2X1_501/O
+ POR2X1_501/CTRL2 POR2X1_501/a_16_28# POR2X1_501/CTRL POR2X1_501/a_76_344# POR2X1_501/a_56_344#
+ POR2X1
XPOR2X1_534 VDD GND POR2X1_42/Y POR2X1_60/A POR2X1_534/Y POR2X1_829/m4_208_n4# POR2X1_534/O
+ POR2X1_534/CTRL2 POR2X1_534/a_16_28# POR2X1_534/CTRL POR2X1_534/a_76_344# POR2X1_534/a_56_344#
+ POR2X1
XPOR2X1_523 VDD GND POR2X1_523/B POR2X1_523/A POR2X1_523/Y POR2X1_523/m4_208_n4# POR2X1_523/O
+ POR2X1_523/CTRL2 POR2X1_523/a_16_28# POR2X1_523/CTRL POR2X1_523/a_76_344# POR2X1_523/a_56_344#
+ POR2X1
XPOR2X1_512 VDD GND D_INPUT_0 POR2X1_308/B POR2X1_513/A POR2X1_512/m4_208_n4# POR2X1_512/O
+ POR2X1_512/CTRL2 POR2X1_512/a_16_28# POR2X1_512/CTRL POR2X1_512/a_76_344# POR2X1_512/a_56_344#
+ POR2X1
XPOR2X1_567 VDD GND POR2X1_567/B POR2X1_567/A POR2X1_568/A POR2X1_567/m4_208_n4# POR2X1_567/O
+ POR2X1_567/CTRL2 POR2X1_567/a_16_28# POR2X1_567/CTRL POR2X1_567/a_76_344# POR2X1_567/a_56_344#
+ POR2X1
XPOR2X1_556 VDD GND POR2X1_631/B POR2X1_556/A POR2X1_556/Y POR2X1_556/m4_208_n4# POR2X1_556/O
+ POR2X1_556/CTRL2 POR2X1_556/a_16_28# POR2X1_556/CTRL POR2X1_556/a_76_344# POR2X1_556/a_56_344#
+ POR2X1
XPOR2X1_578 VDD GND POR2X1_568/Y POR2X1_577/Y POR2X1_578/Y POR2X1_578/m4_208_n4# POR2X1_578/O
+ POR2X1_578/CTRL2 POR2X1_578/a_16_28# POR2X1_578/CTRL POR2X1_578/a_76_344# POR2X1_578/a_56_344#
+ POR2X1
XPOR2X1_545 VDD GND POR2X1_443/A POR2X1_545/A POR2X1_551/A POR2X1_545/m4_208_n4# POR2X1_545/O
+ POR2X1_545/CTRL2 POR2X1_545/a_16_28# POR2X1_545/CTRL POR2X1_545/a_76_344# POR2X1_545/a_56_344#
+ POR2X1
XPOR2X1_589 VDD GND POR2X1_43/B POR2X1_129/Y POR2X1_589/Y POR2X1_589/m4_208_n4# POR2X1_589/O
+ POR2X1_589/CTRL2 POR2X1_589/a_16_28# POR2X1_589/CTRL POR2X1_589/a_76_344# POR2X1_589/a_56_344#
+ POR2X1
XPAND2X1_519 VDD GND POR2X1_260/A PAND2X1_48/A POR2X1_520/A PAND2X1_519/a_16_344#
+ PAND2X1_492/m4_208_n4# PAND2X1_519/O PAND2X1_519/a_56_28# PAND2X1_519/CTRL2 PAND2X1_519/CTRL
+ PAND2X1_519/a_76_28# PAND2X1
XPAND2X1_508 VDD GND PAND2X1_508/B PAND2X1_506/Y PAND2X1_508/Y PAND2X1_508/a_16_344#
+ PAND2X1_508/m4_208_n4# PAND2X1_508/O PAND2X1_508/a_56_28# PAND2X1_508/CTRL2 PAND2X1_508/CTRL
+ PAND2X1_508/a_76_28# PAND2X1
XPOR2X1_342 VDD GND POR2X1_342/B POR2X1_342/A POR2X1_342/Y POR2X1_342/m4_208_n4# POR2X1_342/O
+ POR2X1_342/CTRL2 POR2X1_342/a_16_28# POR2X1_342/CTRL POR2X1_342/a_76_344# POR2X1_342/a_56_344#
+ POR2X1
XPOR2X1_331 VDD GND POR2X1_594/A POR2X1_331/A POR2X1_331/Y POR2X1_331/m4_208_n4# POR2X1_331/O
+ POR2X1_331/CTRL2 POR2X1_331/a_16_28# POR2X1_331/CTRL POR2X1_331/a_76_344# POR2X1_331/a_56_344#
+ POR2X1
XPOR2X1_353 VDD GND POR2X1_566/A POR2X1_353/A POR2X1_353/Y POR2X1_353/m4_208_n4# POR2X1_353/O
+ POR2X1_353/CTRL2 POR2X1_353/a_16_28# POR2X1_353/CTRL POR2X1_353/a_76_344# POR2X1_353/a_56_344#
+ POR2X1
XPOR2X1_320 VDD GND POR2X1_39/B POR2X1_90/Y POR2X1_320/Y POR2X1_320/m4_208_n4# POR2X1_320/O
+ POR2X1_320/CTRL2 POR2X1_320/a_16_28# POR2X1_320/CTRL POR2X1_320/a_76_344# POR2X1_320/a_56_344#
+ POR2X1
XPOR2X1_364 VDD GND POR2X1_357/Y POR2X1_364/A POR2X1_365/A POR2X1_364/m4_208_n4# POR2X1_364/O
+ POR2X1_364/CTRL2 POR2X1_364/a_16_28# POR2X1_364/CTRL POR2X1_364/a_76_344# POR2X1_364/a_56_344#
+ POR2X1
XPOR2X1_386 VDD GND INPUT_4 POR2X1_36/B POR2X1_386/Y POR2X1_386/m4_208_n4# POR2X1_386/O
+ POR2X1_386/CTRL2 POR2X1_386/a_16_28# POR2X1_386/CTRL POR2X1_386/a_76_344# POR2X1_386/a_56_344#
+ POR2X1
XPOR2X1_375 VDD GND PAND2X1_32/B POR2X1_260/A POR2X1_375/Y POR2X1_22/m4_208_n4# POR2X1_375/O
+ POR2X1_375/CTRL2 POR2X1_375/a_16_28# POR2X1_375/CTRL POR2X1_375/a_76_344# POR2X1_375/a_56_344#
+ POR2X1
XPOR2X1_397 VDD GND POR2X1_7/B POR2X1_83/A POR2X1_397/Y POR2X1_397/m4_208_n4# POR2X1_397/O
+ POR2X1_397/CTRL2 POR2X1_397/a_16_28# POR2X1_397/CTRL POR2X1_397/a_76_344# POR2X1_397/a_56_344#
+ POR2X1
XPAND2X1_327 VDD GND POR2X1_667/A POR2X1_63/Y POR2X1_760/A PAND2X1_327/a_16_344# PAND2X1_327/m4_208_n4#
+ PAND2X1_327/O PAND2X1_327/a_56_28# PAND2X1_327/CTRL2 PAND2X1_327/CTRL PAND2X1_327/a_76_28#
+ PAND2X1
XPAND2X1_316 VDD GND PAND2X1_81/B POR2X1_260/B POR2X1_318/A PAND2X1_316/a_16_344#
+ PAND2X1_316/m4_208_n4# PAND2X1_316/O PAND2X1_316/a_56_28# PAND2X1_316/CTRL2 PAND2X1_316/CTRL
+ PAND2X1_316/a_76_28# PAND2X1
XPAND2X1_305 VDD GND PAND2X1_90/Y POR2X1_66/B POR2X1_307/A PAND2X1_305/a_16_344# PAND2X1_305/m4_208_n4#
+ PAND2X1_305/O PAND2X1_305/a_56_28# PAND2X1_305/CTRL2 PAND2X1_305/CTRL PAND2X1_305/a_76_28#
+ PAND2X1
XPAND2X1_338 VDD GND PAND2X1_338/B PAND2X1_333/Y PAND2X1_351/A PAND2X1_338/a_16_344#
+ PAND2X1_338/m4_208_n4# PAND2X1_338/O PAND2X1_338/a_56_28# PAND2X1_338/CTRL2 PAND2X1_338/CTRL
+ PAND2X1_338/a_76_28# PAND2X1
XPAND2X1_349 VDD GND PAND2X1_349/B PAND2X1_349/A PAND2X1_359/B PAND2X1_349/a_16_344#
+ PAND2X1_349/m4_208_n4# PAND2X1_349/O PAND2X1_349/a_56_28# PAND2X1_349/CTRL2 PAND2X1_349/CTRL
+ PAND2X1_349/a_76_28# PAND2X1
XPAND2X1_850 VDD GND PAND2X1_843/Y PAND2X1_842/Y PAND2X1_850/Y PAND2X1_850/a_16_344#
+ PAND2X1_850/m4_208_n4# PAND2X1_850/O PAND2X1_850/a_56_28# PAND2X1_850/CTRL2 PAND2X1_850/CTRL
+ PAND2X1_850/a_76_28# PAND2X1
XPAND2X1_861 VDD GND PAND2X1_861/B PAND2X1_658/A PAND2X1_865/A PAND2X1_861/a_16_344#
+ PAND2X1_861/m4_208_n4# PAND2X1_861/O PAND2X1_861/a_56_28# PAND2X1_861/CTRL2 PAND2X1_861/CTRL
+ PAND2X1_861/a_76_28# PAND2X1
XPOR2X1_150 VDD GND POR2X1_37/Y POR2X1_62/Y POR2X1_150/Y POR2X1_150/m4_208_n4# POR2X1_150/O
+ POR2X1_150/CTRL2 POR2X1_150/a_16_28# POR2X1_150/CTRL POR2X1_150/a_76_344# POR2X1_150/a_56_344#
+ POR2X1
XPOR2X1_161 VDD GND POR2X1_614/A POR2X1_750/B POR2X1_161/Y POR2X1_161/m4_208_n4# POR2X1_161/O
+ POR2X1_161/CTRL2 POR2X1_161/a_16_28# POR2X1_161/CTRL POR2X1_161/a_76_344# POR2X1_161/a_56_344#
+ POR2X1
XPOR2X1_194 VDD GND POR2X1_194/B POR2X1_194/A POR2X1_200/A POR2X1_194/m4_208_n4# POR2X1_194/O
+ POR2X1_194/CTRL2 POR2X1_194/a_16_28# POR2X1_194/CTRL POR2X1_194/a_76_344# POR2X1_194/a_56_344#
+ POR2X1
XPOR2X1_172 VDD GND POR2X1_72/B POR2X1_102/Y POR2X1_172/Y POR2X1_172/m4_208_n4# POR2X1_172/O
+ POR2X1_172/CTRL2 POR2X1_172/a_16_28# POR2X1_172/CTRL POR2X1_172/a_76_344# POR2X1_172/a_56_344#
+ POR2X1
XPOR2X1_183 VDD GND POR2X1_7/A POR2X1_40/Y POR2X1_183/Y POR2X1_183/m4_208_n4# POR2X1_183/O
+ POR2X1_183/CTRL2 POR2X1_183/a_16_28# POR2X1_183/CTRL POR2X1_183/a_76_344# POR2X1_183/a_56_344#
+ POR2X1
XPAND2X1_102 VDD GND POR2X1_94/A PAND2X1_8/Y POR2X1_590/A PAND2X1_102/a_16_344# PAND2X1_102/m4_208_n4#
+ PAND2X1_102/O PAND2X1_102/a_56_28# PAND2X1_102/CTRL2 PAND2X1_102/CTRL PAND2X1_102/a_76_28#
+ PAND2X1
XPAND2X1_135 VDD GND POR2X1_614/A PAND2X1_60/B POR2X1_702/A PAND2X1_135/a_16_344#
+ PAND2X1_135/m4_208_n4# PAND2X1_135/O PAND2X1_135/a_56_28# PAND2X1_135/CTRL2 PAND2X1_135/CTRL
+ PAND2X1_135/a_76_28# PAND2X1
XPAND2X1_113 VDD GND POR2X1_107/Y POR2X1_103/Y PAND2X1_114/B PAND2X1_113/a_16_344#
+ PAND2X1_113/m4_208_n4# PAND2X1_113/O PAND2X1_113/a_56_28# PAND2X1_113/CTRL2 PAND2X1_113/CTRL
+ PAND2X1_113/a_76_28# PAND2X1
XPAND2X1_124 VDD GND PAND2X1_123/Y POR2X1_122/Y PAND2X1_124/Y PAND2X1_124/a_16_344#
+ PAND2X1_124/m4_208_n4# PAND2X1_124/O PAND2X1_124/a_56_28# PAND2X1_124/CTRL2 PAND2X1_124/CTRL
+ PAND2X1_124/a_76_28# PAND2X1
XPAND2X1_179 VDD GND POR2X1_814/B PAND2X1_69/A POR2X1_181/A PAND2X1_179/a_16_344#
+ PAND2X1_179/m4_208_n4# PAND2X1_179/O PAND2X1_179/a_56_28# PAND2X1_179/CTRL2 PAND2X1_179/CTRL
+ PAND2X1_179/a_76_28# PAND2X1
XPAND2X1_146 VDD GND POR2X1_532/A PAND2X1_69/A POR2X1_148/A PAND2X1_146/a_16_344#
+ PAND2X1_146/m4_208_n4# PAND2X1_146/O PAND2X1_146/a_56_28# PAND2X1_146/CTRL2 PAND2X1_146/CTRL
+ PAND2X1_146/a_76_28# PAND2X1
XPAND2X1_168 VDD GND POR2X1_165/Y POR2X1_164/Y PAND2X1_168/Y PAND2X1_168/a_16_344#
+ PAND2X1_168/m4_208_n4# PAND2X1_168/O PAND2X1_168/a_56_28# PAND2X1_168/CTRL2 PAND2X1_168/CTRL
+ PAND2X1_168/a_76_28# PAND2X1
XPAND2X1_157 VDD GND PAND2X1_18/B PAND2X1_3/B POR2X1_260/A PAND2X1_157/a_16_344# PAND2X1_157/m4_208_n4#
+ PAND2X1_157/O PAND2X1_157/a_56_28# PAND2X1_157/CTRL2 PAND2X1_157/CTRL PAND2X1_157/a_76_28#
+ PAND2X1
XPOR2X1_90 VDD GND POR2X1_37/Y POR2X1_54/Y POR2X1_90/Y POR2X1_90/m4_208_n4# POR2X1_90/O
+ POR2X1_90/CTRL2 POR2X1_90/a_16_28# POR2X1_90/CTRL POR2X1_90/a_76_344# POR2X1_90/a_56_344#
+ POR2X1
XPAND2X1_680 VDD GND POR2X1_186/Y PAND2X1_52/B POR2X1_728/A PAND2X1_680/a_16_344#
+ PAND2X1_680/m4_208_n4# PAND2X1_680/O PAND2X1_680/a_56_28# PAND2X1_680/CTRL2 PAND2X1_680/CTRL
+ PAND2X1_680/a_76_28# PAND2X1
XPAND2X1_691 VDD GND POR2X1_690/Y POR2X1_689/Y PAND2X1_691/Y PAND2X1_691/a_16_344#
+ PAND2X1_691/m4_208_n4# PAND2X1_691/O PAND2X1_691/a_56_28# PAND2X1_691/CTRL2 PAND2X1_691/CTRL
+ PAND2X1_691/a_76_28# PAND2X1
XPAND2X1_1 VDD GND INPUT_7 D_INPUT_6 PAND2X1_3/A PAND2X1_1/a_16_344# PAND2X1_1/m4_208_n4#
+ PAND2X1_1/O PAND2X1_1/a_56_28# PAND2X1_1/CTRL2 PAND2X1_1/CTRL PAND2X1_1/a_76_28#
+ PAND2X1
XPOR2X1_716 VDD GND POR2X1_228/Y POR2X1_303/B POR2X1_723/B POR2X1_301/m4_208_n4# POR2X1_716/O
+ POR2X1_716/CTRL2 POR2X1_716/a_16_28# POR2X1_716/CTRL POR2X1_716/a_76_344# POR2X1_716/a_56_344#
+ POR2X1
XPOR2X1_705 VDD GND POR2X1_705/B POR2X1_546/A POR2X1_713/B POR2X1_705/m4_208_n4# POR2X1_705/O
+ POR2X1_705/CTRL2 POR2X1_705/a_16_28# POR2X1_705/CTRL POR2X1_705/a_76_344# POR2X1_705/a_56_344#
+ POR2X1
XPOR2X1_727 VDD GND POR2X1_353/A POR2X1_444/Y POR2X1_731/A POR2X1_727/m4_208_n4# POR2X1_727/O
+ POR2X1_727/CTRL2 POR2X1_727/a_16_28# POR2X1_727/CTRL POR2X1_727/a_76_344# POR2X1_727/a_56_344#
+ POR2X1
XPOR2X1_749 VDD GND INPUT_0 POR2X1_8/Y POR2X1_749/Y POR2X1_749/m4_208_n4# POR2X1_749/O
+ POR2X1_749/CTRL2 POR2X1_749/a_16_28# POR2X1_749/CTRL POR2X1_749/a_76_344# POR2X1_749/a_56_344#
+ POR2X1
XPOR2X1_738 VDD GND POR2X1_731/Y POR2X1_738/A POR2X1_738/Y POR2X1_738/m4_208_n4# POR2X1_738/O
+ POR2X1_738/CTRL2 POR2X1_738/a_16_28# POR2X1_738/CTRL POR2X1_738/a_76_344# POR2X1_738/a_56_344#
+ POR2X1
XPOR2X1_9 VDD GND INPUT_0 INPUT_1 POR2X1_9/Y POR2X1_9/m4_208_n4# POR2X1_9/O POR2X1_9/CTRL2
+ POR2X1_9/a_16_28# POR2X1_9/CTRL POR2X1_9/a_76_344# POR2X1_9/a_56_344# POR2X1
XPOR2X1_502 VDD GND POR2X1_78/A POR2X1_502/A POR2X1_502/Y POR2X1_502/m4_208_n4# POR2X1_502/O
+ POR2X1_502/CTRL2 POR2X1_502/a_16_28# POR2X1_502/CTRL POR2X1_502/a_76_344# POR2X1_502/a_56_344#
+ POR2X1
XPOR2X1_524 VDD GND POR2X1_48/A POR2X1_257/A POR2X1_524/Y POR2X1_524/m4_208_n4# POR2X1_524/O
+ POR2X1_524/CTRL2 POR2X1_524/a_16_28# POR2X1_524/CTRL POR2X1_524/a_76_344# POR2X1_524/a_56_344#
+ POR2X1
XPOR2X1_535 VDD GND POR2X1_788/B POR2X1_535/A POR2X1_567/B POR2X1_535/m4_208_n4# POR2X1_535/O
+ POR2X1_535/CTRL2 POR2X1_535/a_16_28# POR2X1_535/CTRL POR2X1_535/a_76_344# POR2X1_535/a_56_344#
+ POR2X1
XPOR2X1_513 VDD GND POR2X1_513/B POR2X1_513/A POR2X1_513/Y POR2X1_513/m4_208_n4# POR2X1_513/O
+ POR2X1_513/CTRL2 POR2X1_513/a_16_28# POR2X1_513/CTRL POR2X1_513/a_76_344# POR2X1_513/a_56_344#
+ POR2X1
XPOR2X1_546 VDD GND POR2X1_546/B POR2X1_546/A POR2X1_550/B POR2X1_546/m4_208_n4# POR2X1_546/O
+ POR2X1_546/CTRL2 POR2X1_546/a_16_28# POR2X1_546/CTRL POR2X1_546/a_76_344# POR2X1_546/a_56_344#
+ POR2X1
XPOR2X1_557 VDD GND POR2X1_557/B POR2X1_557/A POR2X1_561/B POR2X1_558/m4_208_n4# POR2X1_557/O
+ POR2X1_557/CTRL2 POR2X1_557/a_16_28# POR2X1_557/CTRL POR2X1_557/a_76_344# POR2X1_557/a_56_344#
+ POR2X1
XPOR2X1_568 VDD GND POR2X1_568/B POR2X1_568/A POR2X1_568/Y POR2X1_568/m4_208_n4# POR2X1_568/O
+ POR2X1_568/CTRL2 POR2X1_568/a_16_28# POR2X1_568/CTRL POR2X1_568/a_76_344# POR2X1_568/a_56_344#
+ POR2X1
XPOR2X1_579 VDD GND POR2X1_579/B POR2X1_576/Y POR2X1_579/Y POR2X1_579/m4_208_n4# POR2X1_579/O
+ POR2X1_579/CTRL2 POR2X1_579/a_16_28# POR2X1_579/CTRL POR2X1_579/a_76_344# POR2X1_579/a_56_344#
+ POR2X1
XPAND2X1_509 VDD GND POR2X1_503/Y PAND2X1_340/B PAND2X1_510/B PAND2X1_509/a_16_344#
+ PAND2X1_509/m4_208_n4# PAND2X1_509/O PAND2X1_509/a_56_28# PAND2X1_509/CTRL2 PAND2X1_509/CTRL
+ PAND2X1_509/a_76_28# PAND2X1
XPOR2X1_310 VDD GND POR2X1_5/Y POR2X1_40/Y POR2X1_310/Y POR2X1_310/m4_208_n4# POR2X1_310/O
+ POR2X1_310/CTRL2 POR2X1_310/a_16_28# POR2X1_310/CTRL POR2X1_310/a_76_344# POR2X1_310/a_56_344#
+ POR2X1
XPOR2X1_332 VDD GND POR2X1_332/B POR2X1_702/A POR2X1_332/Y POR2X1_332/m4_208_n4# POR2X1_332/O
+ POR2X1_332/CTRL2 POR2X1_332/a_16_28# POR2X1_332/CTRL POR2X1_332/a_76_344# POR2X1_332/a_56_344#
+ POR2X1
XPOR2X1_343 VDD GND POR2X1_343/B POR2X1_343/A POR2X1_343/Y POR2X1_343/m4_208_n4# POR2X1_343/O
+ POR2X1_343/CTRL2 POR2X1_343/a_16_28# POR2X1_343/CTRL POR2X1_343/a_76_344# POR2X1_343/a_56_344#
+ POR2X1
XPOR2X1_321 VDD GND POR2X1_41/B POR2X1_65/A POR2X1_321/Y POR2X1_320/m4_208_n4# POR2X1_321/O
+ POR2X1_321/CTRL2 POR2X1_321/a_16_28# POR2X1_321/CTRL POR2X1_321/a_76_344# POR2X1_321/a_56_344#
+ POR2X1
XPOR2X1_376 VDD GND POR2X1_376/B POR2X1_376/A POR2X1_376/Y POR2X1_376/m4_208_n4# POR2X1_376/O
+ POR2X1_376/CTRL2 POR2X1_376/a_16_28# POR2X1_376/CTRL POR2X1_376/a_76_344# POR2X1_376/a_56_344#
+ POR2X1
XPOR2X1_365 VDD GND POR2X1_356/Y POR2X1_365/A POR2X1_365/Y POR2X1_365/m4_208_n4# POR2X1_365/O
+ POR2X1_365/CTRL2 POR2X1_365/a_16_28# POR2X1_365/CTRL POR2X1_365/a_76_344# POR2X1_365/a_56_344#
+ POR2X1
XPOR2X1_354 VDD GND POR2X1_319/Y POR2X1_854/B POR2X1_356/B POR2X1_354/m4_208_n4# POR2X1_354/O
+ POR2X1_354/CTRL2 POR2X1_354/a_16_28# POR2X1_354/CTRL POR2X1_354/a_76_344# POR2X1_354/a_56_344#
+ POR2X1
XPOR2X1_398 VDD GND POR2X1_78/B POR2X1_294/A POR2X1_398/Y POR2X1_398/m4_208_n4# POR2X1_398/O
+ POR2X1_398/CTRL2 POR2X1_398/a_16_28# POR2X1_398/CTRL POR2X1_398/a_76_344# POR2X1_398/a_56_344#
+ POR2X1
XPOR2X1_387 VDD GND POR2X1_93/A POR2X1_386/Y POR2X1_387/Y POR2X1_387/m4_208_n4# POR2X1_387/O
+ POR2X1_387/CTRL2 POR2X1_387/a_16_28# POR2X1_387/CTRL POR2X1_387/a_76_344# POR2X1_387/a_56_344#
+ POR2X1
XPAND2X1_306 VDD GND POR2X1_502/A PAND2X1_58/A POR2X1_308/B PAND2X1_306/a_16_344#
+ PAND2X1_306/m4_208_n4# PAND2X1_306/O PAND2X1_306/a_56_28# PAND2X1_306/CTRL2 PAND2X1_306/CTRL
+ PAND2X1_306/a_76_28# PAND2X1
XPAND2X1_317 VDD GND POR2X1_314/Y POR2X1_313/Y PAND2X1_317/Y PAND2X1_317/a_16_344#
+ PAND2X1_317/m4_208_n4# PAND2X1_317/O PAND2X1_317/a_56_28# PAND2X1_317/CTRL2 PAND2X1_317/CTRL
+ PAND2X1_317/a_76_28# PAND2X1
XPAND2X1_328 VDD GND PAND2X1_95/B D_INPUT_4 POR2X1_596/A PAND2X1_328/a_16_344# PAND2X1_328/m4_208_n4#
+ PAND2X1_328/O PAND2X1_328/a_56_28# PAND2X1_328/CTRL2 PAND2X1_328/CTRL PAND2X1_328/a_76_28#
+ PAND2X1
XPAND2X1_339 VDD GND PAND2X1_332/Y PAND2X1_61/Y PAND2X1_339/Y PAND2X1_339/a_16_344#
+ PAND2X1_339/m4_208_n4# PAND2X1_339/O PAND2X1_339/a_56_28# PAND2X1_339/CTRL2 PAND2X1_339/CTRL
+ PAND2X1_339/a_76_28# PAND2X1
XPAND2X1_840 VDD GND PAND2X1_840/B PAND2X1_840/A PAND2X1_840/Y PAND2X1_840/a_16_344#
+ PAND2X1_840/m4_208_n4# PAND2X1_840/O PAND2X1_840/a_56_28# PAND2X1_840/CTRL2 PAND2X1_840/CTRL
+ PAND2X1_840/a_76_28# PAND2X1
XPAND2X1_851 VDD GND PAND2X1_841/Y PAND2X1_840/Y PAND2X1_858/B PAND2X1_851/a_16_344#
+ PAND2X1_851/m4_208_n4# PAND2X1_851/O PAND2X1_851/a_56_28# PAND2X1_851/CTRL2 PAND2X1_851/CTRL
+ PAND2X1_851/a_76_28# PAND2X1
XPAND2X1_862 VDD GND PAND2X1_862/B PAND2X1_858/Y PAND2X1_862/Y PAND2X1_862/a_16_344#
+ PAND2X1_862/m4_208_n4# PAND2X1_862/O PAND2X1_862/a_56_28# PAND2X1_862/CTRL2 PAND2X1_862/CTRL
+ PAND2X1_862/a_76_28# PAND2X1
XPOR2X1_140 VDD GND POR2X1_140/B POR2X1_140/A POR2X1_141/A POR2X1_140/m4_208_n4# POR2X1_140/O
+ POR2X1_140/CTRL2 POR2X1_140/a_16_28# POR2X1_140/CTRL POR2X1_140/a_76_344# POR2X1_140/a_56_344#
+ POR2X1
XPOR2X1_151 VDD GND PAND2X1_55/Y POR2X1_186/B POR2X1_151/Y POR2X1_151/m4_208_n4# POR2X1_151/O
+ POR2X1_151/CTRL2 POR2X1_151/a_16_28# POR2X1_151/CTRL POR2X1_151/a_76_344# POR2X1_151/a_56_344#
+ POR2X1
XPOR2X1_195 VDD GND PAND2X1_41/Y POR2X1_195/A POR2X1_199/B POR2X1_195/m4_208_n4# POR2X1_195/O
+ POR2X1_195/CTRL2 POR2X1_195/a_16_28# POR2X1_195/CTRL POR2X1_195/a_76_344# POR2X1_195/a_56_344#
+ POR2X1
XPOR2X1_184 VDD GND POR2X1_71/Y POR2X1_96/A POR2X1_184/Y POR2X1_184/m4_208_n4# POR2X1_184/O
+ POR2X1_184/CTRL2 POR2X1_184/a_16_28# POR2X1_184/CTRL POR2X1_184/a_76_344# POR2X1_184/a_56_344#
+ POR2X1
XPOR2X1_173 VDD GND POR2X1_72/B POR2X1_150/Y POR2X1_173/Y POR2X1_173/m4_208_n4# POR2X1_173/O
+ POR2X1_173/CTRL2 POR2X1_173/a_16_28# POR2X1_173/CTRL POR2X1_173/a_76_344# POR2X1_173/a_56_344#
+ POR2X1
XPOR2X1_162 VDD GND POR2X1_162/B POR2X1_161/Y POR2X1_162/Y POR2X1_162/m4_208_n4# POR2X1_162/O
+ POR2X1_162/CTRL2 POR2X1_162/a_16_28# POR2X1_162/CTRL POR2X1_162/a_76_344# POR2X1_162/a_56_344#
+ POR2X1
XPAND2X1_103 VDD GND POR2X1_590/A PAND2X1_48/B POR2X1_113/B PAND2X1_103/a_16_344#
+ PAND2X1_103/m4_208_n4# PAND2X1_103/O PAND2X1_103/a_56_28# PAND2X1_103/CTRL2 PAND2X1_103/CTRL
+ PAND2X1_103/a_76_28# PAND2X1
XPAND2X1_136 VDD GND POR2X1_296/B POR2X1_66/B POR2X1_138/A PAND2X1_136/a_16_344# POR2X1_514/m4_208_n4#
+ PAND2X1_136/O PAND2X1_136/a_56_28# PAND2X1_136/CTRL2 PAND2X1_136/CTRL PAND2X1_136/a_76_28#
+ PAND2X1
XPAND2X1_125 VDD GND POR2X1_814/B PAND2X1_96/B POR2X1_128/B PAND2X1_125/a_16_344#
+ PAND2X1_125/m4_208_n4# PAND2X1_125/O PAND2X1_125/a_56_28# PAND2X1_125/CTRL2 PAND2X1_125/CTRL
+ PAND2X1_125/a_76_28# PAND2X1
XPAND2X1_114 VDD GND PAND2X1_114/B POR2X1_108/Y PAND2X1_114/Y PAND2X1_114/a_16_344#
+ PAND2X1_114/m4_208_n4# PAND2X1_114/O PAND2X1_114/a_56_28# PAND2X1_114/CTRL2 PAND2X1_114/CTRL
+ PAND2X1_114/a_76_28# PAND2X1
XPAND2X1_169 VDD GND POR2X1_167/Y POR2X1_166/Y PAND2X1_169/Y PAND2X1_169/a_16_344#
+ PAND2X1_169/m4_208_n4# PAND2X1_169/O PAND2X1_169/a_56_28# PAND2X1_169/CTRL2 PAND2X1_169/CTRL
+ PAND2X1_169/a_76_28# PAND2X1
XPAND2X1_147 VDD GND POR2X1_144/Y POR2X1_142/Y PAND2X1_149/A PAND2X1_147/a_16_344#
+ PAND2X1_147/m4_208_n4# PAND2X1_147/O PAND2X1_147/a_56_28# PAND2X1_147/CTRL2 PAND2X1_147/CTRL
+ PAND2X1_147/a_76_28# PAND2X1
XPAND2X1_158 VDD GND POR2X1_260/A POR2X1_156/Y POR2X1_210/B PAND2X1_158/a_16_344#
+ PAND2X1_158/m4_208_n4# PAND2X1_158/O PAND2X1_158/a_56_28# PAND2X1_158/CTRL2 PAND2X1_158/CTRL
+ PAND2X1_158/a_76_28# PAND2X1
XPOR2X1_80 VDD GND POR2X1_5/Y POR2X1_29/A POR2X1_81/A POR2X1_80/m4_208_n4# POR2X1_80/O
+ POR2X1_80/CTRL2 POR2X1_80/a_16_28# POR2X1_80/CTRL POR2X1_80/a_76_344# POR2X1_80/a_56_344#
+ POR2X1
XPOR2X1_91 VDD GND POR2X1_52/A POR2X1_90/Y POR2X1_91/Y POR2X1_91/m4_208_n4# POR2X1_91/O
+ POR2X1_91/CTRL2 POR2X1_91/a_16_28# POR2X1_91/CTRL POR2X1_91/a_76_344# POR2X1_91/a_56_344#
+ POR2X1
XPAND2X1_692 VDD GND PAND2X1_48/A PAND2X1_20/A POR2X1_706/B PAND2X1_692/a_16_344#
+ PAND2X1_692/m4_208_n4# PAND2X1_692/O PAND2X1_692/a_56_28# PAND2X1_692/CTRL2 PAND2X1_692/CTRL
+ PAND2X1_692/a_76_28# PAND2X1
XPAND2X1_681 VDD GND POR2X1_407/A PAND2X1_32/B POR2X1_685/B PAND2X1_681/a_16_344#
+ PAND2X1_681/m4_208_n4# PAND2X1_681/O PAND2X1_681/a_56_28# PAND2X1_681/CTRL2 PAND2X1_681/CTRL
+ PAND2X1_681/a_76_28# PAND2X1
XPAND2X1_670 VDD GND POR2X1_590/A PAND2X1_41/B POR2X1_673/B PAND2X1_670/a_16_344#
+ PAND2X1_54/m4_208_n4# PAND2X1_670/O PAND2X1_670/a_56_28# PAND2X1_670/CTRL2 PAND2X1_670/CTRL
+ PAND2X1_670/a_76_28# PAND2X1
XPAND2X1_2 VDD GND D_INPUT_5 D_INPUT_4 PAND2X1_3/B PAND2X1_2/a_16_344# PAND2X1_2/m4_208_n4#
+ PAND2X1_2/O PAND2X1_2/a_56_28# PAND2X1_2/CTRL2 PAND2X1_2/CTRL PAND2X1_2/a_76_28#
+ PAND2X1
C0 POR2X1_556/Y PAND2X1_60/B 0.02fF
C1 POR2X1_215/Y POR2X1_631/B 0.06fF
C2 POR2X1_567/A PAND2X1_90/Y 0.08fF
C3 PAND2X1_81/a_16_344# PAND2X1_60/B 0.02fF
C4 PAND2X1_777/CTRL POR2X1_293/Y 0.01fF
C5 POR2X1_188/A POR2X1_858/A 0.01fF
C6 PAND2X1_716/B VDD 0.74fF
C7 D_GATE_662 POR2X1_456/B 0.07fF
C8 PAND2X1_347/Y POR2X1_385/Y 0.05fF
C9 POR2X1_360/A POR2X1_334/A 0.09fF
C10 PAND2X1_686/O POR2X1_42/Y 0.02fF
C11 POR2X1_614/A PAND2X1_315/O 0.09fF
C12 PAND2X1_850/a_76_28# PAND2X1_842/Y 0.07fF
C13 POR2X1_96/A PAND2X1_156/A 0.05fF
C14 POR2X1_327/Y POR2X1_276/CTRL2 0.01fF
C15 POR2X1_16/A PAND2X1_401/O 0.01fF
C16 POR2X1_730/Y POR2X1_732/CTRL 0.01fF
C17 PAND2X1_54/O POR2X1_4/Y 0.09fF
C18 GATE_662 VDD 0.10fF
C19 POR2X1_8/Y D_INPUT_2 0.03fF
C20 PAND2X1_787/A PAND2X1_388/Y 0.08fF
C21 POR2X1_287/B PAND2X1_122/a_16_344# 0.01fF
C22 POR2X1_49/Y POR2X1_39/B 0.27fF
C23 POR2X1_540/Y VDD 1.05fF
C24 PAND2X1_90/Y POR2X1_542/O 0.04fF
C25 PAND2X1_138/m4_208_n4# POR2X1_39/B 0.15fF
C26 PAND2X1_687/CTRL2 POR2X1_829/A 0.00fF
C27 PAND2X1_644/O POR2X1_597/Y 0.04fF
C28 POR2X1_271/A POR2X1_256/m4_208_n4# 0.07fF
C29 POR2X1_16/A POR2X1_816/A 0.05fF
C30 POR2X1_502/A POR2X1_191/Y 0.13fF
C31 POR2X1_865/O POR2X1_101/Y 0.05fF
C32 D_INPUT_1 POR2X1_456/B 0.03fF
C33 PAND2X1_57/B POR2X1_4/Y 0.00fF
C34 PAND2X1_474/A POR2X1_77/Y 0.03fF
C35 PAND2X1_509/a_76_28# POR2X1_503/Y 0.07fF
C36 POR2X1_858/B POR2X1_840/B 0.04fF
C37 POR2X1_327/Y PAND2X1_152/a_76_28# 0.03fF
C38 PAND2X1_48/B POR2X1_726/CTRL2 0.01fF
C39 POR2X1_130/O PAND2X1_6/Y 0.01fF
C40 PAND2X1_90/Y POR2X1_779/CTRL2 0.03fF
C41 POR2X1_57/A POR2X1_744/CTRL2 0.01fF
C42 PAND2X1_90/m4_208_n4# POR2X1_546/A 0.08fF
C43 POR2X1_356/A POR2X1_447/B 0.03fF
C44 PAND2X1_737/CTRL2 POR2X1_7/B 0.01fF
C45 POR2X1_41/B PAND2X1_865/Y 0.07fF
C46 POR2X1_68/A POR2X1_593/O 0.02fF
C47 POR2X1_176/CTRL2 PAND2X1_566/Y 0.01fF
C48 POR2X1_456/B POR2X1_724/A 0.08fF
C49 POR2X1_537/Y POR2X1_740/Y 0.03fF
C50 PAND2X1_4/CTRL POR2X1_260/A 0.01fF
C51 PAND2X1_28/CTRL PAND2X1_63/B 0.01fF
C52 PAND2X1_469/B PAND2X1_357/O 0.27fF
C53 PAND2X1_95/B PAND2X1_328/O -0.00fF
C54 PAND2X1_197/Y POR2X1_7/Y 0.07fF
C55 PAND2X1_682/O POR2X1_809/A 0.00fF
C56 POR2X1_407/Y POR2X1_596/a_76_344# 0.00fF
C57 POR2X1_62/Y POR2X1_620/O 0.16fF
C58 POR2X1_313/a_16_28# POR2X1_313/Y 0.02fF
C59 PAND2X1_170/CTRL2 POR2X1_73/Y 0.01fF
C60 POR2X1_286/B POR2X1_649/O 0.00fF
C61 PAND2X1_274/O POR2X1_39/B 0.01fF
C62 POR2X1_711/B POR2X1_710/CTRL 0.01fF
C63 POR2X1_730/Y POR2X1_383/A 0.03fF
C64 POR2X1_16/A PAND2X1_854/A 0.04fF
C65 PAND2X1_620/O POR2X1_408/Y 0.05fF
C66 POR2X1_356/A POR2X1_510/O 0.01fF
C67 PAND2X1_553/B POR2X1_39/B 0.07fF
C68 INPUT_6 PAND2X1_2/CTRL2 0.01fF
C69 PAND2X1_687/m4_208_n4# POR2X1_761/m4_208_n4# 0.13fF
C70 POR2X1_416/B POR2X1_625/Y 0.00fF
C71 POR2X1_394/A PAND2X1_121/CTRL2 0.10fF
C72 POR2X1_52/A POR2X1_305/O 0.01fF
C73 POR2X1_27/CTRL POR2X1_669/B 0.01fF
C74 POR2X1_68/B PAND2X1_396/CTRL2 0.01fF
C75 VDD POR2X1_343/B 0.25fF
C76 POR2X1_681/CTRL POR2X1_32/A 0.01fF
C77 POR2X1_110/Y POR2X1_417/a_16_28# 0.03fF
C78 POR2X1_52/A PAND2X1_440/a_16_344# 0.02fF
C79 POR2X1_7/A PAND2X1_156/A 0.14fF
C80 PAND2X1_93/B POR2X1_276/B 0.01fF
C81 PAND2X1_341/B PAND2X1_338/B 0.03fF
C82 POR2X1_517/CTRL POR2X1_73/Y 0.04fF
C83 POR2X1_327/Y PAND2X1_534/a_76_28# 0.05fF
C84 POR2X1_158/Y PAND2X1_705/CTRL2 0.00fF
C85 POR2X1_624/CTRL POR2X1_94/A 0.13fF
C86 POR2X1_335/A POR2X1_343/Y 0.05fF
C87 POR2X1_135/CTRL2 POR2X1_7/A 0.03fF
C88 POR2X1_84/A POR2X1_243/B 0.03fF
C89 POR2X1_485/Y POR2X1_32/A 0.03fF
C90 POR2X1_257/A POR2X1_48/A 16.63fF
C91 POR2X1_673/CTRL2 POR2X1_624/B 0.10fF
C92 POR2X1_825/Y PAND2X1_673/Y 0.03fF
C93 POR2X1_520/B POR2X1_559/A 0.01fF
C94 POR2X1_669/B POR2X1_20/B 0.32fF
C95 POR2X1_83/a_16_28# POR2X1_153/Y 0.07fF
C96 PAND2X1_3/a_16_344# PAND2X1_3/B 0.05fF
C97 PAND2X1_682/O POR2X1_728/A 0.00fF
C98 POR2X1_666/O POR2X1_411/B 0.01fF
C99 POR2X1_54/Y PAND2X1_68/O 0.02fF
C100 POR2X1_446/B POR2X1_218/Y 0.00fF
C101 PAND2X1_611/CTRL POR2X1_389/Y 0.00fF
C102 POR2X1_327/Y POR2X1_186/B 0.03fF
C103 POR2X1_341/A POR2X1_296/B 0.07fF
C104 POR2X1_48/A POR2X1_612/B 0.01fF
C105 POR2X1_777/B PAND2X1_246/O 0.02fF
C106 PAND2X1_65/B POR2X1_260/CTRL2 0.00fF
C107 POR2X1_23/Y PAND2X1_477/O 0.13fF
C108 POR2X1_866/A POR2X1_811/CTRL 0.26fF
C109 POR2X1_359/B POR2X1_334/Y 0.02fF
C110 POR2X1_738/A POR2X1_738/a_16_28# 0.03fF
C111 POR2X1_307/A POR2X1_711/Y 0.06fF
C112 PAND2X1_403/B POR2X1_411/B 0.00fF
C113 POR2X1_116/A POR2X1_330/Y 0.05fF
C114 PAND2X1_483/O PAND2X1_631/A 0.15fF
C115 POR2X1_848/CTRL VDD 0.00fF
C116 POR2X1_416/B POR2X1_695/CTRL2 0.00fF
C117 POR2X1_410/Y PAND2X1_52/B 0.04fF
C118 POR2X1_465/a_16_28# POR2X1_186/Y 0.03fF
C119 INPUT_3 POR2X1_69/A 0.05fF
C120 PAND2X1_74/CTRL POR2X1_341/A 0.07fF
C121 PAND2X1_332/Y PAND2X1_858/Y 0.14fF
C122 POR2X1_411/B POR2X1_272/CTRL 0.03fF
C123 POR2X1_832/A PAND2X1_56/A 0.03fF
C124 POR2X1_67/Y PAND2X1_381/a_16_344# 0.01fF
C125 POR2X1_537/Y POR2X1_774/A 0.03fF
C126 POR2X1_458/Y PAND2X1_57/B 0.07fF
C127 POR2X1_343/B PAND2X1_32/B 0.80fF
C128 POR2X1_14/Y PAND2X1_407/O 0.01fF
C129 POR2X1_66/B POR2X1_66/Y 0.03fF
C130 POR2X1_416/B PAND2X1_551/a_16_344# 0.01fF
C131 POR2X1_286/O POR2X1_66/A 0.01fF
C132 POR2X1_210/Y POR2X1_568/A 0.03fF
C133 POR2X1_250/Y VDD 0.99fF
C134 POR2X1_409/B POR2X1_37/Y 0.09fF
C135 POR2X1_728/O POR2X1_814/A 0.37fF
C136 POR2X1_499/A POR2X1_573/CTRL2 0.08fF
C137 PAND2X1_175/B PAND2X1_862/CTRL2 0.01fF
C138 PAND2X1_388/O POR2X1_167/Y 0.02fF
C139 PAND2X1_454/B POR2X1_40/Y 0.03fF
C140 POR2X1_62/Y POR2X1_7/Y 0.00fF
C141 PAND2X1_637/CTRL PAND2X1_638/B 0.01fF
C142 PAND2X1_637/O POR2X1_585/Y -0.00fF
C143 PAND2X1_452/A POR2X1_158/Y 0.03fF
C144 POR2X1_617/Y POR2X1_616/Y 0.02fF
C145 PAND2X1_792/B PAND2X1_792/a_16_344# 0.02fF
C146 POR2X1_704/Y POR2X1_169/A 0.01fF
C147 POR2X1_566/B PAND2X1_52/B 0.03fF
C148 POR2X1_492/Y POR2X1_394/A 0.06fF
C149 POR2X1_192/B POR2X1_357/B 0.18fF
C150 POR2X1_49/Y PAND2X1_469/CTRL2 0.01fF
C151 POR2X1_180/A PAND2X1_52/B 0.03fF
C152 PAND2X1_57/B PAND2X1_45/O 0.01fF
C153 PAND2X1_10/CTRL POR2X1_296/B 0.01fF
C154 POR2X1_444/CTRL VDD 0.00fF
C155 POR2X1_490/Y PAND2X1_217/B 0.12fF
C156 POR2X1_20/B POR2X1_297/Y 0.14fF
C157 POR2X1_441/Y PAND2X1_738/Y 0.05fF
C158 POR2X1_23/Y POR2X1_40/Y 0.32fF
C159 POR2X1_278/Y POR2X1_262/Y 0.01fF
C160 POR2X1_158/Y PAND2X1_713/CTRL2 0.00fF
C161 PAND2X1_48/B POR2X1_462/CTRL 0.00fF
C162 PAND2X1_242/Y PAND2X1_175/B 0.00fF
C163 POR2X1_555/A POR2X1_454/A 0.10fF
C164 POR2X1_287/B POR2X1_458/CTRL 0.01fF
C165 POR2X1_65/A POR2X1_438/Y 0.03fF
C166 POR2X1_49/Y POR2X1_48/A 0.20fF
C167 POR2X1_604/Y POR2X1_603/Y 0.19fF
C168 POR2X1_866/B POR2X1_866/A 0.05fF
C169 POR2X1_832/A POR2X1_661/A 0.14fF
C170 POR2X1_445/A VDD 0.87fF
C171 POR2X1_812/CTRL POR2X1_452/Y 0.01fF
C172 POR2X1_848/A POR2X1_5/Y 1.12fF
C173 PAND2X1_405/O POR2X1_38/Y 0.17fF
C174 PAND2X1_844/Y POR2X1_20/B 0.01fF
C175 PAND2X1_73/Y PAND2X1_46/CTRL2 0.06fF
C176 POR2X1_537/Y PAND2X1_108/CTRL 0.01fF
C177 POR2X1_115/CTRL POR2X1_446/B 0.01fF
C178 POR2X1_38/CTRL VDD 0.00fF
C179 POR2X1_807/A D_INPUT_0 0.07fF
C180 POR2X1_490/Y VDD 0.49fF
C181 POR2X1_78/A POR2X1_264/O 0.12fF
C182 PAND2X1_282/a_16_344# PAND2X1_41/B 0.02fF
C183 POR2X1_833/CTRL POR2X1_541/B 0.08fF
C184 POR2X1_65/A POR2X1_487/O 0.07fF
C185 POR2X1_748/A POR2X1_420/Y 0.01fF
C186 PAND2X1_617/CTRL2 POR2X1_68/B 0.03fF
C187 PAND2X1_94/A PAND2X1_233/CTRL 0.00fF
C188 POR2X1_602/B POR2X1_811/B 0.03fF
C189 POR2X1_79/Y PAND2X1_205/CTRL2 0.01fF
C190 POR2X1_383/A PAND2X1_255/O 0.08fF
C191 PAND2X1_449/CTRL2 POR2X1_90/Y 0.01fF
C192 POR2X1_54/Y POR2X1_615/Y 0.01fF
C193 PAND2X1_865/Y POR2X1_77/Y 0.07fF
C194 POR2X1_502/A POR2X1_866/A 0.10fF
C195 POR2X1_669/B PAND2X1_381/CTRL2 0.16fF
C196 POR2X1_376/B PAND2X1_796/O 0.15fF
C197 POR2X1_150/Y POR2X1_183/Y 0.03fF
C198 PAND2X1_20/A POR2X1_489/CTRL 0.03fF
C199 POR2X1_377/CTRL2 POR2X1_54/Y 0.01fF
C200 POR2X1_23/Y PAND2X1_659/B 0.04fF
C201 POR2X1_801/O POR2X1_121/B 0.03fF
C202 POR2X1_296/CTRL PAND2X1_69/A 0.00fF
C203 POR2X1_60/A PAND2X1_140/O 0.03fF
C204 POR2X1_814/B POR2X1_243/A 0.02fF
C205 POR2X1_738/a_16_28# POR2X1_731/Y -0.00fF
C206 POR2X1_48/A POR2X1_481/CTRL 0.00fF
C207 POR2X1_65/A POR2X1_603/Y 0.01fF
C208 POR2X1_552/a_16_28# PAND2X1_72/A 0.03fF
C209 PAND2X1_407/O POR2X1_55/Y 0.25fF
C210 POR2X1_338/CTRL POR2X1_814/A 0.07fF
C211 POR2X1_508/B PAND2X1_52/B 0.00fF
C212 PAND2X1_624/CTRL POR2X1_29/A 0.01fF
C213 POR2X1_394/A POR2X1_321/CTRL 0.06fF
C214 POR2X1_817/O POR2X1_817/A 0.04fF
C215 PAND2X1_860/A POR2X1_153/Y 0.13fF
C216 POR2X1_68/CTRL2 PAND2X1_57/B 0.01fF
C217 POR2X1_661/m4_208_n4# POR2X1_78/A 0.09fF
C218 POR2X1_515/a_16_28# D_INPUT_0 0.01fF
C219 PAND2X1_841/Y PAND2X1_840/Y 0.02fF
C220 POR2X1_68/A POR2X1_446/B 0.05fF
C221 POR2X1_48/A PAND2X1_553/B 0.02fF
C222 PAND2X1_612/B PAND2X1_283/CTRL 0.00fF
C223 POR2X1_259/A POR2X1_186/Y 0.01fF
C224 POR2X1_460/CTRL2 POR2X1_260/B 0.03fF
C225 POR2X1_389/Y POR2X1_734/A 0.07fF
C226 POR2X1_231/CTRL POR2X1_66/A 0.00fF
C227 POR2X1_836/CTRL POR2X1_578/Y 0.03fF
C228 POR2X1_27/Y POR2X1_5/Y 0.01fF
C229 POR2X1_567/B POR2X1_466/O 0.01fF
C230 POR2X1_504/Y PAND2X1_620/Y 0.03fF
C231 POR2X1_409/B POR2X1_293/Y 0.03fF
C232 PAND2X1_61/CTRL POR2X1_58/Y 0.01fF
C233 POR2X1_278/Y POR2X1_498/Y 0.15fF
C234 POR2X1_210/O POR2X1_220/Y 0.00fF
C235 POR2X1_865/B POR2X1_475/O 0.01fF
C236 POR2X1_72/B PAND2X1_778/CTRL2 0.03fF
C237 POR2X1_566/A POR2X1_241/B 0.03fF
C238 D_INPUT_0 POR2X1_546/B 0.01fF
C239 PAND2X1_93/B PAND2X1_144/O 0.01fF
C240 POR2X1_334/Y PAND2X1_257/O 0.06fF
C241 PAND2X1_104/a_76_28# POR2X1_814/B 0.02fF
C242 POR2X1_719/A POR2X1_130/A -0.06fF
C243 POR2X1_646/Y POR2X1_784/A 0.03fF
C244 POR2X1_83/B PAND2X1_734/B 0.00fF
C245 PAND2X1_671/Y POR2X1_35/B 0.01fF
C246 POR2X1_429/O VDD 0.00fF
C247 POR2X1_490/O POR2X1_7/A 0.01fF
C248 POR2X1_640/O INPUT_0 0.04fF
C249 PAND2X1_56/Y POR2X1_218/Y 0.10fF
C250 POR2X1_308/m4_208_n4# POR2X1_794/B 0.08fF
C251 POR2X1_13/A PAND2X1_795/CTRL2 0.01fF
C252 PAND2X1_251/CTRL PAND2X1_69/A 0.01fF
C253 POR2X1_268/Y INPUT_0 0.11fF
C254 PAND2X1_81/CTRL2 POR2X1_66/A 0.03fF
C255 POR2X1_66/A POR2X1_391/Y 0.07fF
C256 POR2X1_97/A D_GATE_222 0.08fF
C257 POR2X1_78/B POR2X1_543/A 0.09fF
C258 PAND2X1_821/CTRL POR2X1_590/A 0.01fF
C259 POR2X1_689/A POR2X1_102/Y 0.00fF
C260 POR2X1_407/A D_INPUT_0 0.12fF
C261 PAND2X1_23/Y POR2X1_287/O 0.01fF
C262 PAND2X1_453/CTRL POR2X1_14/Y 0.01fF
C263 POR2X1_378/Y PAND2X1_459/CTRL 0.01fF
C264 D_INPUT_0 POR2X1_56/Y 0.07fF
C265 PAND2X1_205/Y VDD 0.34fF
C266 POR2X1_407/A POR2X1_811/A 0.03fF
C267 PAND2X1_23/Y PAND2X1_11/Y 0.01fF
C268 PAND2X1_39/B POR2X1_725/Y 0.07fF
C269 PAND2X1_248/O POR2X1_532/A 0.02fF
C270 POR2X1_482/Y POR2X1_252/CTRL 0.01fF
C271 POR2X1_629/B POR2X1_785/A 0.01fF
C272 POR2X1_299/O PAND2X1_776/Y 0.03fF
C273 POR2X1_763/A POR2X1_701/Y 0.04fF
C274 PAND2X1_61/Y INPUT_0 0.22fF
C275 POR2X1_667/A POR2X1_42/Y 0.03fF
C276 POR2X1_624/Y PAND2X1_133/CTRL2 0.01fF
C277 POR2X1_849/A D_INPUT_1 0.06fF
C278 POR2X1_647/CTRL PAND2X1_60/B 0.00fF
C279 PAND2X1_843/CTRL POR2X1_251/Y 0.01fF
C280 POR2X1_407/A POR2X1_287/CTRL2 0.01fF
C281 POR2X1_48/A PAND2X1_778/Y 0.03fF
C282 PAND2X1_784/CTRL2 POR2X1_72/B 0.03fF
C283 PAND2X1_403/B PAND2X1_398/CTRL2 0.10fF
C284 POR2X1_16/A INPUT_3 0.03fF
C285 POR2X1_702/B PAND2X1_57/B 0.01fF
C286 POR2X1_102/Y PAND2X1_398/O 0.02fF
C287 PAND2X1_467/Y POR2X1_694/Y 0.01fF
C288 POR2X1_68/A POR2X1_121/B 0.18fF
C289 PAND2X1_435/Y POR2X1_56/Y 0.00fF
C290 POR2X1_556/A POR2X1_216/Y 0.01fF
C291 PAND2X1_72/A POR2X1_181/A 0.10fF
C292 POR2X1_302/CTRL2 POR2X1_302/Y 0.00fF
C293 POR2X1_13/a_16_28# POR2X1_250/A 0.01fF
C294 POR2X1_29/A POR2X1_409/CTRL 0.01fF
C295 POR2X1_231/B POR2X1_186/Y 0.01fF
C296 POR2X1_2/O VDD 0.00fF
C297 PAND2X1_262/CTRL POR2X1_786/A 0.04fF
C298 POR2X1_54/Y PAND2X1_819/a_16_344# 0.02fF
C299 PAND2X1_390/Y POR2X1_55/Y 0.03fF
C300 PAND2X1_192/Y PAND2X1_191/CTRL2 0.01fF
C301 POR2X1_586/Y PAND2X1_69/A 0.00fF
C302 PAND2X1_787/CTRL POR2X1_7/B 0.01fF
C303 PAND2X1_47/B PAND2X1_587/O 0.02fF
C304 POR2X1_445/A POR2X1_543/CTRL2 0.03fF
C305 POR2X1_634/CTRL2 POR2X1_391/Y 0.01fF
C306 PAND2X1_96/B POR2X1_174/A 0.03fF
C307 POR2X1_850/B POR2X1_513/Y 0.03fF
C308 PAND2X1_90/Y PAND2X1_386/Y 0.03fF
C309 POR2X1_856/B POR2X1_510/Y 0.16fF
C310 POR2X1_13/A POR2X1_236/Y 0.23fF
C311 PAND2X1_20/A POR2X1_713/Y 0.04fF
C312 POR2X1_49/Y PAND2X1_197/Y 0.03fF
C313 POR2X1_33/O POR2X1_68/B 0.02fF
C314 PAND2X1_151/CTRL VDD 0.00fF
C315 POR2X1_409/B POR2X1_408/Y 0.16fF
C316 POR2X1_591/A POR2X1_591/a_16_28# 0.08fF
C317 POR2X1_93/A POR2X1_225/CTRL 0.03fF
C318 PAND2X1_696/CTRL POR2X1_648/Y 0.02fF
C319 POR2X1_475/A POR2X1_717/Y 0.03fF
C320 POR2X1_329/CTRL PAND2X1_362/B 0.01fF
C321 POR2X1_383/A POR2X1_218/Y 0.10fF
C322 POR2X1_114/Y VDD 0.02fF
C323 PAND2X1_90/A POR2X1_5/Y 0.06fF
C324 PAND2X1_421/O PAND2X1_65/B 0.01fF
C325 PAND2X1_474/Y POR2X1_81/Y 0.16fF
C326 POR2X1_60/A PAND2X1_509/O 0.00fF
C327 PAND2X1_152/CTRL VDD 0.00fF
C328 PAND2X1_387/CTRL2 POR2X1_712/Y 0.03fF
C329 PAND2X1_93/B POR2X1_456/B 0.06fF
C330 PAND2X1_258/CTRL2 POR2X1_260/A 0.03fF
C331 POR2X1_78/A PAND2X1_173/O 0.04fF
C332 PAND2X1_216/B PAND2X1_218/B 0.00fF
C333 POR2X1_814/B POR2X1_204/O 0.01fF
C334 POR2X1_750/B POR2X1_556/Y 0.05fF
C335 PAND2X1_243/B VDD 0.48fF
C336 POR2X1_60/A POR2X1_142/Y 0.09fF
C337 POR2X1_842/O POR2X1_675/Y 0.01fF
C338 POR2X1_834/Y POR2X1_66/A 0.03fF
C339 POR2X1_20/B PAND2X1_353/Y 0.03fF
C340 POR2X1_3/A POR2X1_748/A 0.79fF
C341 PAND2X1_48/B POR2X1_215/CTRL 0.01fF
C342 POR2X1_777/B POR2X1_68/B 0.07fF
C343 POR2X1_84/CTRL2 PAND2X1_57/B 0.03fF
C344 PAND2X1_642/O POR2X1_48/A 0.01fF
C345 PAND2X1_639/B VDD 0.01fF
C346 POR2X1_407/A PAND2X1_90/Y 0.08fF
C347 PAND2X1_850/Y POR2X1_150/Y 0.03fF
C348 POR2X1_847/A POR2X1_408/Y 0.02fF
C349 POR2X1_63/O POR2X1_236/Y 0.02fF
C350 PAND2X1_81/B POR2X1_786/O 0.01fF
C351 POR2X1_186/Y PAND2X1_88/Y 0.03fF
C352 PAND2X1_20/A POR2X1_725/Y 0.01fF
C353 PAND2X1_48/B POR2X1_76/Y 0.03fF
C354 POR2X1_278/Y PAND2X1_287/O 0.00fF
C355 POR2X1_248/CTRL POR2X1_5/Y 0.00fF
C356 POR2X1_390/B POR2X1_590/A 0.07fF
C357 POR2X1_423/Y POR2X1_91/Y 0.03fF
C358 PAND2X1_249/a_76_28# POR2X1_38/Y 0.03fF
C359 PAND2X1_197/CTRL PAND2X1_364/B 0.03fF
C360 POR2X1_474/CTRL2 POR2X1_101/Y 0.12fF
C361 POR2X1_255/CTRL PAND2X1_349/A 0.01fF
C362 POR2X1_567/B POR2X1_566/CTRL 0.03fF
C363 POR2X1_78/A POR2X1_456/B 0.06fF
C364 PAND2X1_477/B POR2X1_237/O 0.02fF
C365 PAND2X1_65/B POR2X1_68/B 2.47fF
C366 POR2X1_51/A POR2X1_22/A 0.34fF
C367 POR2X1_502/A PAND2X1_95/a_56_28# 0.00fF
C368 PAND2X1_817/CTRL POR2X1_750/Y 0.03fF
C369 POR2X1_748/A POR2X1_748/Y 0.01fF
C370 POR2X1_614/A POR2X1_370/Y 0.01fF
C371 POR2X1_468/a_16_28# POR2X1_468/B -0.00fF
C372 PAND2X1_738/CTRL2 PAND2X1_149/A 0.01fF
C373 POR2X1_734/A POR2X1_713/B 0.07fF
C374 PAND2X1_643/Y POR2X1_236/Y 0.07fF
C375 POR2X1_78/B POR2X1_243/CTRL 0.03fF
C376 POR2X1_57/A POR2X1_485/CTRL 0.01fF
C377 PAND2X1_635/Y POR2X1_386/Y 0.03fF
C378 POR2X1_376/Y POR2X1_376/A 0.01fF
C379 PAND2X1_472/A PAND2X1_673/Y 0.79fF
C380 PAND2X1_651/Y PAND2X1_573/CTRL2 0.06fF
C381 POR2X1_740/Y PAND2X1_152/O 0.00fF
C382 PAND2X1_63/Y VDD 1.57fF
C383 POR2X1_558/B POR2X1_294/A 0.03fF
C384 POR2X1_175/a_16_28# POR2X1_614/A 0.01fF
C385 POR2X1_388/CTRL POR2X1_566/A 0.01fF
C386 PAND2X1_48/B POR2X1_740/Y 0.11fF
C387 POR2X1_70/CTRL2 POR2X1_90/Y 0.12fF
C388 POR2X1_476/A POR2X1_113/B 0.03fF
C389 POR2X1_61/Y POR2X1_215/Y 0.01fF
C390 POR2X1_52/A POR2X1_289/CTRL 0.01fF
C391 POR2X1_462/B PAND2X1_57/B 0.03fF
C392 POR2X1_45/Y PAND2X1_215/B 0.07fF
C393 POR2X1_383/A POR2X1_710/A 0.01fF
C394 POR2X1_504/CTRL POR2X1_14/Y 0.00fF
C395 POR2X1_196/Y POR2X1_244/B 0.02fF
C396 POR2X1_814/B POR2X1_725/Y 0.07fF
C397 PAND2X1_676/CTRL VDD 0.00fF
C398 POR2X1_809/A POR2X1_801/B 0.01fF
C399 PAND2X1_852/CTRL POR2X1_42/Y 0.01fF
C400 PAND2X1_655/B VDD 0.03fF
C401 POR2X1_406/Y PAND2X1_560/CTRL2 0.04fF
C402 POR2X1_347/B PAND2X1_69/CTRL 0.05fF
C403 POR2X1_416/B POR2X1_411/B 1.05fF
C404 POR2X1_13/A PAND2X1_858/Y 0.01fF
C405 POR2X1_614/A PAND2X1_309/CTRL 0.01fF
C406 D_GATE_222 POR2X1_294/B 0.02fF
C407 POR2X1_446/B POR2X1_169/A 0.05fF
C408 POR2X1_658/m4_208_n4# POR2X1_554/m4_208_n4# 0.13fF
C409 PAND2X1_736/A PAND2X1_652/A 0.10fF
C410 POR2X1_46/Y POR2X1_90/Y 0.03fF
C411 PAND2X1_20/A POR2X1_559/A 0.03fF
C412 PAND2X1_460/CTRL2 PAND2X1_472/B 0.01fF
C413 POR2X1_102/Y PAND2X1_508/a_76_28# 0.00fF
C414 POR2X1_65/A PAND2X1_467/Y 0.03fF
C415 POR2X1_72/B PAND2X1_861/O 0.01fF
C416 PAND2X1_707/Y PAND2X1_725/A 0.06fF
C417 POR2X1_807/A POR2X1_590/a_76_344# 0.00fF
C418 POR2X1_587/CTRL POR2X1_587/Y 0.00fF
C419 POR2X1_355/B POR2X1_341/Y 0.03fF
C420 PAND2X1_57/B POR2X1_724/A 0.07fF
C421 PAND2X1_188/CTRL2 POR2X1_816/A 0.01fF
C422 POR2X1_680/Y POR2X1_816/A 0.03fF
C423 PAND2X1_534/CTRL VDD 0.00fF
C424 POR2X1_833/CTRL2 POR2X1_786/Y 0.02fF
C425 PAND2X1_535/a_16_344# POR2X1_236/Y 0.00fF
C426 POR2X1_364/A POR2X1_785/A 0.01fF
C427 POR2X1_111/O POR2X1_46/Y 0.02fF
C428 POR2X1_220/Y POR2X1_220/A 0.01fF
C429 PAND2X1_8/CTRL2 INPUT_2 0.05fF
C430 POR2X1_250/A PAND2X1_537/O 0.07fF
C431 PAND2X1_484/a_76_28# PAND2X1_73/Y 0.01fF
C432 PAND2X1_56/Y POR2X1_68/A 0.10fF
C433 POR2X1_22/A POR2X1_408/a_16_28# 0.05fF
C434 PAND2X1_675/A POR2X1_437/Y 0.01fF
C435 POR2X1_72/B PAND2X1_704/O 0.01fF
C436 PAND2X1_857/A VDD 0.18fF
C437 POR2X1_594/Y POR2X1_594/A 0.00fF
C438 PAND2X1_803/a_76_28# POR2X1_83/B 0.01fF
C439 POR2X1_573/CTRL POR2X1_456/B 0.01fF
C440 INPUT_1 POR2X1_627/CTRL2 0.10fF
C441 PAND2X1_696/O POR2X1_66/A 0.02fF
C442 POR2X1_334/Y POR2X1_330/Y 0.07fF
C443 POR2X1_685/A VDD 0.00fF
C444 POR2X1_446/A PAND2X1_72/A 0.06fF
C445 PAND2X1_65/B POR2X1_502/O 0.16fF
C446 PAND2X1_41/B POR2X1_544/B 0.03fF
C447 D_INPUT_3 POR2X1_7/B 0.03fF
C448 PAND2X1_374/O VDD 0.00fF
C449 POR2X1_241/Y POR2X1_566/B 0.26fF
C450 POR2X1_259/B PAND2X1_52/Y 0.69fF
C451 PAND2X1_651/Y PAND2X1_339/Y 0.03fF
C452 POR2X1_66/A POR2X1_383/Y 0.07fF
C453 PAND2X1_614/a_16_344# POR2X1_129/Y 0.01fF
C454 POR2X1_294/B POR2X1_702/CTRL2 0.01fF
C455 PAND2X1_726/B POR2X1_763/O 0.03fF
C456 POR2X1_25/Y POR2X1_748/A 0.03fF
C457 PAND2X1_65/B PAND2X1_103/m4_208_n4# 0.08fF
C458 POR2X1_220/Y POR2X1_569/A 0.07fF
C459 PAND2X1_63/Y PAND2X1_81/B 0.03fF
C460 PAND2X1_347/Y PAND2X1_343/CTRL 0.01fF
C461 INPUT_0 POR2X1_385/O 0.01fF
C462 POR2X1_234/A POR2X1_20/B 0.05fF
C463 POR2X1_368/a_16_28# POR2X1_283/A 0.09fF
C464 POR2X1_516/Y PAND2X1_851/a_76_28# 0.02fF
C465 PAND2X1_40/CTRL POR2X1_407/Y 0.01fF
C466 VDD POR2X1_260/A 4.16fF
C467 PAND2X1_645/B POR2X1_665/Y 0.03fF
C468 PAND2X1_592/Y POR2X1_283/A 0.03fF
C469 POR2X1_49/Y POR2X1_62/Y 0.10fF
C470 PAND2X1_567/O PAND2X1_568/B 0.00fF
C471 POR2X1_778/B PAND2X1_69/A 0.02fF
C472 POR2X1_532/A POR2X1_391/Y 0.10fF
C473 PAND2X1_216/a_76_28# PAND2X1_656/A 0.01fF
C474 POR2X1_404/Y POR2X1_569/A 0.07fF
C475 POR2X1_81/Y PAND2X1_510/B 0.08fF
C476 POR2X1_245/Y POR2X1_42/Y 0.02fF
C477 POR2X1_516/m4_208_n4# POR2X1_184/Y 0.12fF
C478 POR2X1_417/Y PAND2X1_352/CTRL 0.01fF
C479 PAND2X1_63/Y PAND2X1_32/B 0.08fF
C480 POR2X1_446/a_16_28# PAND2X1_72/A 0.00fF
C481 POR2X1_57/A PAND2X1_779/Y 0.01fF
C482 PAND2X1_536/O PAND2X1_60/B 0.03fF
C483 PAND2X1_854/A PAND2X1_324/Y 0.01fF
C484 PAND2X1_414/CTRL2 POR2X1_67/Y 0.01fF
C485 PAND2X1_292/CTRL POR2X1_66/A 0.01fF
C486 PAND2X1_568/B PAND2X1_566/Y 0.01fF
C487 PAND2X1_216/B PAND2X1_793/Y 0.03fF
C488 PAND2X1_579/B POR2X1_394/A 0.03fF
C489 POR2X1_697/Y PAND2X1_550/B 0.00fF
C490 POR2X1_3/A PAND2X1_635/O 0.17fF
C491 POR2X1_363/A VDD 0.22fF
C492 POR2X1_703/A PAND2X1_176/O 0.02fF
C493 PAND2X1_430/CTRL2 PAND2X1_3/B 0.01fF
C494 POR2X1_35/Y POR2X1_215/Y 0.01fF
C495 POR2X1_43/B PAND2X1_349/A 0.03fF
C496 PAND2X1_6/Y PAND2X1_60/B 11.36fF
C497 POR2X1_464/Y POR2X1_703/A 0.05fF
C498 POR2X1_43/B PAND2X1_63/B 0.03fF
C499 POR2X1_68/A POR2X1_383/A 0.27fF
C500 POR2X1_476/A POR2X1_768/A 0.01fF
C501 POR2X1_271/A POR2X1_13/A 0.02fF
C502 POR2X1_359/B POR2X1_349/Y -0.00fF
C503 POR2X1_131/CTRL2 PAND2X1_349/A 0.01fF
C504 POR2X1_334/B PAND2X1_94/A 0.26fF
C505 POR2X1_199/O PAND2X1_824/B 0.06fF
C506 POR2X1_113/Y PAND2X1_32/B 0.03fF
C507 PAND2X1_800/O PAND2X1_863/B 0.02fF
C508 POR2X1_614/A PAND2X1_63/B 0.11fF
C509 PAND2X1_85/Y POR2X1_4/Y 0.01fF
C510 PAND2X1_560/O PAND2X1_844/B -0.00fF
C511 POR2X1_504/CTRL POR2X1_55/Y 0.01fF
C512 POR2X1_186/Y POR2X1_568/B 0.12fF
C513 POR2X1_394/A POR2X1_763/Y 0.14fF
C514 POR2X1_741/Y POR2X1_260/A 2.77fF
C515 POR2X1_16/A PAND2X1_675/A 0.20fF
C516 POR2X1_43/Y POR2X1_669/B 0.07fF
C517 POR2X1_791/A PAND2X1_60/B 0.06fF
C518 POR2X1_42/Y PAND2X1_507/CTRL 0.01fF
C519 PAND2X1_539/Y PAND2X1_794/B 0.03fF
C520 POR2X1_685/A PAND2X1_32/B 0.00fF
C521 POR2X1_88/A PAND2X1_206/B 0.02fF
C522 POR2X1_416/B PAND2X1_742/O 0.04fF
C523 POR2X1_38/B PAND2X1_63/B 0.03fF
C524 POR2X1_776/B POR2X1_566/O 0.01fF
C525 PAND2X1_480/CTRL2 POR2X1_43/B 0.03fF
C526 PAND2X1_608/CTRL POR2X1_411/B 0.01fF
C527 POR2X1_164/O POR2X1_164/Y 0.01fF
C528 POR2X1_553/A POR2X1_112/Y 0.03fF
C529 POR2X1_302/Y POR2X1_188/Y 0.01fF
C530 POR2X1_532/A PAND2X1_528/CTRL2 0.01fF
C531 POR2X1_416/B POR2X1_24/CTRL2 0.15fF
C532 PAND2X1_94/A POR2X1_124/B 0.05fF
C533 POR2X1_51/A POR2X1_328/O 0.01fF
C534 POR2X1_110/Y POR2X1_693/CTRL 0.06fF
C535 PAND2X1_48/B POR2X1_774/A 0.03fF
C536 POR2X1_190/Y POR2X1_192/B 0.01fF
C537 POR2X1_96/A PAND2X1_858/a_56_28# 0.00fF
C538 PAND2X1_727/CTRL2 POR2X1_90/Y 0.00fF
C539 POR2X1_388/O POR2X1_703/A 0.03fF
C540 PAND2X1_610/CTRL VDD 0.00fF
C541 POR2X1_508/m4_208_n4# PAND2X1_824/m4_208_n4# 0.04fF
C542 POR2X1_161/Y POR2X1_162/Y 0.07fF
C543 POR2X1_73/Y PAND2X1_123/a_16_344# 0.02fF
C544 POR2X1_584/a_76_344# POR2X1_260/A 0.00fF
C545 PAND2X1_284/a_16_344# POR2X1_394/A 0.02fF
C546 POR2X1_260/A PAND2X1_32/B 0.51fF
C547 VDD PAND2X1_508/B 0.06fF
C548 PAND2X1_803/Y POR2X1_108/Y 0.06fF
C549 POR2X1_141/Y PAND2X1_72/A 0.12fF
C550 PAND2X1_631/A POR2X1_252/CTRL2 -0.00fF
C551 POR2X1_669/B POR2X1_321/CTRL 0.16fF
C552 POR2X1_834/Y POR2X1_532/A 0.03fF
C553 POR2X1_41/B PAND2X1_352/Y 0.01fF
C554 POR2X1_130/A PAND2X1_136/O 0.05fF
C555 PAND2X1_423/CTRL2 PAND2X1_72/A 0.01fF
C556 POR2X1_416/B POR2X1_376/B 0.07fF
C557 POR2X1_790/A POR2X1_720/CTRL 0.04fF
C558 PAND2X1_612/O POR2X1_472/B 0.02fF
C559 POR2X1_532/A PAND2X1_690/O 0.01fF
C560 POR2X1_680/O POR2X1_79/Y 0.01fF
C561 POR2X1_394/A POR2X1_73/Y 0.24fF
C562 POR2X1_5/Y POR2X1_80/O 0.01fF
C563 POR2X1_327/Y POR2X1_542/B 0.03fF
C564 POR2X1_675/A PAND2X1_72/A 0.01fF
C565 PAND2X1_294/CTRL2 POR2X1_150/Y 0.03fF
C566 POR2X1_258/Y PAND2X1_569/Y 0.07fF
C567 POR2X1_596/A POR2X1_596/a_16_28# 0.09fF
C568 POR2X1_326/O POR2X1_319/Y 0.01fF
C569 POR2X1_326/CTRL POR2X1_854/B -0.00fF
C570 POR2X1_567/A D_GATE_222 0.10fF
C571 PAND2X1_823/O POR2X1_854/B 0.02fF
C572 POR2X1_52/CTRL PAND2X1_215/B 0.03fF
C573 POR2X1_557/A POR2X1_569/A 0.07fF
C574 POR2X1_119/Y POR2X1_234/CTRL 0.04fF
C575 POR2X1_150/Y POR2X1_437/CTRL 0.01fF
C576 POR2X1_88/O POR2X1_88/A 0.14fF
C577 POR2X1_505/CTRL PAND2X1_632/B 0.01fF
C578 POR2X1_571/CTRL POR2X1_569/A 0.05fF
C579 POR2X1_614/A POR2X1_552/A 0.01fF
C580 POR2X1_20/B POR2X1_298/CTRL2 0.00fF
C581 POR2X1_52/A POR2X1_416/B 0.16fF
C582 PAND2X1_97/Y D_INPUT_0 0.08fF
C583 PAND2X1_409/CTRL2 PAND2X1_52/B 0.16fF
C584 POR2X1_494/Y POR2X1_77/Y 0.03fF
C585 POR2X1_673/Y POR2X1_260/A 0.01fF
C586 POR2X1_503/CTRL POR2X1_8/Y 0.00fF
C587 POR2X1_220/Y PAND2X1_72/A 0.10fF
C588 PAND2X1_244/B POR2X1_394/A 0.07fF
C589 POR2X1_43/B PAND2X1_860/a_76_28# 0.01fF
C590 POR2X1_116/A POR2X1_558/B 0.34fF
C591 POR2X1_287/A D_INPUT_0 0.00fF
C592 PAND2X1_5/O POR2X1_4/Y 0.02fF
C593 POR2X1_728/a_16_28# POR2X1_728/A 0.03fF
C594 POR2X1_43/CTRL2 POR2X1_43/B 0.01fF
C595 PAND2X1_60/a_76_28# PAND2X1_39/B 0.05fF
C596 PAND2X1_317/Y POR2X1_416/B 5.40fF
C597 POR2X1_404/Y PAND2X1_72/A 0.03fF
C598 PAND2X1_86/Y POR2X1_334/A 0.02fF
C599 PAND2X1_309/O POR2X1_717/B 0.02fF
C600 POR2X1_811/CTRL2 PAND2X1_39/B 0.01fF
C601 POR2X1_709/B PAND2X1_698/CTRL 0.00fF
C602 POR2X1_27/O POR2X1_27/Y 0.00fF
C603 POR2X1_343/A POR2X1_458/Y 0.05fF
C604 POR2X1_861/A POR2X1_383/A 0.24fF
C605 POR2X1_532/A POR2X1_383/Y 0.03fF
C606 POR2X1_716/O POR2X1_723/B 0.01fF
C607 INPUT_1 PAND2X1_156/A 0.01fF
C608 POR2X1_228/CTRL POR2X1_260/A 0.01fF
C609 PAND2X1_691/Y PAND2X1_687/O 0.08fF
C610 PAND2X1_645/Y POR2X1_600/Y 0.03fF
C611 POR2X1_858/B POR2X1_737/A 0.03fF
C612 PAND2X1_217/B POR2X1_329/A 0.05fF
C613 POR2X1_362/A POR2X1_294/A 0.03fF
C614 PAND2X1_10/O PAND2X1_9/Y 0.02fF
C615 D_INPUT_6 D_INPUT_4 0.95fF
C616 POR2X1_620/A POR2X1_624/Y 0.06fF
C617 POR2X1_342/Y POR2X1_532/A 0.01fF
C618 POR2X1_768/CTRL POR2X1_294/A 0.03fF
C619 POR2X1_38/Y PAND2X1_339/O 0.16fF
C620 PAND2X1_601/a_16_344# D_INPUT_0 0.01fF
C621 POR2X1_632/Y PAND2X1_60/B 0.03fF
C622 PAND2X1_23/Y POR2X1_303/B 0.03fF
C623 PAND2X1_681/O PAND2X1_32/B 0.02fF
C624 PAND2X1_39/B POR2X1_811/B 0.02fF
C625 PAND2X1_66/CTRL2 POR2X1_67/A 0.03fF
C626 POR2X1_159/CTRL INPUT_3 0.16fF
C627 PAND2X1_303/Y PAND2X1_353/Y 0.05fF
C628 POR2X1_329/A VDD 0.85fF
C629 POR2X1_150/Y PAND2X1_211/A 0.00fF
C630 POR2X1_865/B POR2X1_717/B 0.09fF
C631 PAND2X1_60/B POR2X1_500/CTRL 0.03fF
C632 PAND2X1_841/CTRL POR2X1_677/Y 0.00fF
C633 POR2X1_858/B POR2X1_858/A 0.07fF
C634 POR2X1_817/CTRL POR2X1_32/A 0.03fF
C635 PAND2X1_60/B PAND2X1_52/B 0.11fF
C636 PAND2X1_265/CTRL2 POR2X1_260/B 0.01fF
C637 POR2X1_54/Y PAND2X1_817/a_56_28# 0.00fF
C638 POR2X1_68/B POR2X1_8/a_76_344# 0.00fF
C639 POR2X1_83/B PAND2X1_66/O 0.00fF
C640 POR2X1_399/CTRL POR2X1_411/B 0.01fF
C641 POR2X1_20/B PAND2X1_499/Y 0.01fF
C642 PAND2X1_60/B PAND2X1_135/a_16_344# 0.02fF
C643 PAND2X1_97/Y PAND2X1_351/CTRL2 0.01fF
C644 PAND2X1_796/B POR2X1_5/Y 0.00fF
C645 PAND2X1_759/O PAND2X1_48/A 0.01fF
C646 POR2X1_60/A POR2X1_409/B 0.10fF
C647 POR2X1_29/A POR2X1_296/B 0.06fF
C648 POR2X1_275/Y VDD 0.03fF
C649 PAND2X1_206/B PAND2X1_341/CTRL 0.01fF
C650 POR2X1_16/a_16_28# POR2X1_73/Y 0.09fF
C651 POR2X1_76/B POR2X1_575/CTRL 0.01fF
C652 POR2X1_866/A POR2X1_862/B 0.03fF
C653 POR2X1_411/B PAND2X1_738/Y 0.05fF
C654 POR2X1_862/A POR2X1_286/Y 0.02fF
C655 PAND2X1_52/B POR2X1_353/A 0.03fF
C656 POR2X1_96/A POR2X1_150/Y 0.12fF
C657 POR2X1_41/B POR2X1_603/CTRL 0.06fF
C658 PAND2X1_432/a_56_28# POR2X1_866/A 0.00fF
C659 PAND2X1_72/A POR2X1_332/CTRL 0.01fF
C660 POR2X1_610/Y VDD 0.00fF
C661 POR2X1_366/Y PAND2X1_417/CTRL 0.05fF
C662 PAND2X1_224/a_16_344# PAND2X1_32/B 0.01fF
C663 POR2X1_864/A POR2X1_828/CTRL 0.00fF
C664 PAND2X1_58/A POR2X1_121/B 0.06fF
C665 POR2X1_150/Y PAND2X1_335/O 0.28fF
C666 POR2X1_60/A PAND2X1_794/CTRL 0.01fF
C667 PAND2X1_65/B POR2X1_848/A 0.15fF
C668 PAND2X1_23/Y POR2X1_705/B 0.09fF
C669 POR2X1_475/A POR2X1_734/B 0.12fF
C670 POR2X1_23/Y POR2X1_5/Y 0.13fF
C671 PAND2X1_613/O PAND2X1_8/Y 0.07fF
C672 PAND2X1_243/B PAND2X1_9/Y 0.03fF
C673 POR2X1_776/A POR2X1_578/Y 0.03fF
C674 POR2X1_353/Y POR2X1_444/A 0.01fF
C675 PAND2X1_31/CTRL2 VDD 0.00fF
C676 POR2X1_445/a_76_344# POR2X1_341/A 0.02fF
C677 PAND2X1_75/CTRL2 POR2X1_532/A 0.01fF
C678 PAND2X1_839/CTRL POR2X1_411/B 0.01fF
C679 POR2X1_814/A POR2X1_68/B 2.79fF
C680 PAND2X1_39/B POR2X1_783/B 0.02fF
C681 PAND2X1_8/CTRL INPUT_3 0.01fF
C682 PAND2X1_341/B POR2X1_85/Y 0.02fF
C683 POR2X1_445/A POR2X1_445/O 0.01fF
C684 POR2X1_54/Y POR2X1_294/B 0.03fF
C685 POR2X1_814/B POR2X1_499/m4_208_n4# 0.05fF
C686 POR2X1_753/a_16_28# POR2X1_752/Y 0.06fF
C687 POR2X1_273/Y POR2X1_411/B 0.10fF
C688 D_INPUT_3 PAND2X1_206/B 0.10fF
C689 PAND2X1_93/B PAND2X1_57/B 0.13fF
C690 PAND2X1_61/Y POR2X1_102/Y 0.03fF
C691 POR2X1_730/Y POR2X1_440/CTRL 0.01fF
C692 PAND2X1_23/Y PAND2X1_67/CTRL 0.01fF
C693 PAND2X1_459/CTRL POR2X1_750/B 0.00fF
C694 PAND2X1_216/CTRL2 PAND2X1_218/B 0.01fF
C695 POR2X1_78/A POR2X1_448/B 0.02fF
C696 POR2X1_490/Y PAND2X1_216/O 0.01fF
C697 POR2X1_692/m4_208_n4# POR2X1_692/Y 0.12fF
C698 POR2X1_655/A PAND2X1_385/CTRL 0.00fF
C699 POR2X1_29/A POR2X1_236/Y 0.08fF
C700 POR2X1_441/Y PAND2X1_724/O 0.01fF
C701 POR2X1_633/Y PAND2X1_73/Y 0.04fF
C702 POR2X1_260/B PAND2X1_55/Y 2.87fF
C703 POR2X1_78/A POR2X1_608/CTRL2 0.03fF
C704 POR2X1_41/Y POR2X1_43/Y 0.00fF
C705 POR2X1_102/Y POR2X1_760/CTRL 0.01fF
C706 POR2X1_454/A POR2X1_563/Y 0.03fF
C707 PAND2X1_63/Y PAND2X1_9/Y 1.36fF
C708 POR2X1_102/Y PAND2X1_778/O 0.05fF
C709 POR2X1_567/B POR2X1_579/Y 0.05fF
C710 POR2X1_243/A VDD 0.11fF
C711 POR2X1_490/O POR2X1_38/Y 0.01fF
C712 POR2X1_60/A POR2X1_272/Y 0.02fF
C713 PAND2X1_326/B PAND2X1_326/a_76_28# 0.04fF
C714 POR2X1_614/A POR2X1_676/O 0.17fF
C715 PAND2X1_85/CTRL2 POR2X1_260/A 0.01fF
C716 PAND2X1_212/CTRL PAND2X1_357/Y 0.01fF
C717 POR2X1_849/O POR2X1_750/B 0.01fF
C718 PAND2X1_477/O POR2X1_238/Y 0.04fF
C719 PAND2X1_218/B PAND2X1_218/O 0.00fF
C720 POR2X1_791/Y PAND2X1_41/B 0.00fF
C721 POR2X1_78/A PAND2X1_57/B 0.04fF
C722 POR2X1_473/O PAND2X1_32/B 0.31fF
C723 POR2X1_752/Y POR2X1_585/O 0.03fF
C724 POR2X1_820/O POR2X1_820/B -0.01fF
C725 POR2X1_60/A PAND2X1_788/O 0.01fF
C726 POR2X1_823/Y POR2X1_411/B 0.02fF
C727 PAND2X1_276/O PAND2X1_390/Y 0.02fF
C728 PAND2X1_831/a_76_28# PAND2X1_217/B 0.10fF
C729 POR2X1_12/A POR2X1_700/Y 0.03fF
C730 PAND2X1_96/B POR2X1_446/B 0.03fF
C731 PAND2X1_217/B PAND2X1_795/m4_208_n4# 0.06fF
C732 POR2X1_150/Y POR2X1_7/A 0.05fF
C733 POR2X1_645/O POR2X1_330/Y 0.34fF
C734 D_INPUT_0 POR2X1_42/Y 0.15fF
C735 POR2X1_136/Y POR2X1_411/B 0.06fF
C736 PAND2X1_23/Y POR2X1_610/m4_208_n4# 0.05fF
C737 POR2X1_427/Y POR2X1_763/A 0.17fF
C738 POR2X1_669/B POR2X1_763/Y 0.07fF
C739 POR2X1_133/CTRL2 POR2X1_40/Y 0.03fF
C740 POR2X1_814/B POR2X1_116/CTRL2 0.03fF
C741 POR2X1_150/Y PAND2X1_130/O 0.05fF
C742 PAND2X1_433/O D_INPUT_0 0.04fF
C743 POR2X1_862/A PAND2X1_69/A 0.07fF
C744 POR2X1_411/B PAND2X1_181/CTRL2 0.01fF
C745 D_INPUT_5 INPUT_6 0.04fF
C746 POR2X1_688/CTRL2 POR2X1_260/A 0.01fF
C747 POR2X1_220/Y PAND2X1_39/m4_208_n4# 0.08fF
C748 POR2X1_811/B POR2X1_513/B 0.31fF
C749 POR2X1_260/B POR2X1_407/Y 0.02fF
C750 POR2X1_614/A POR2X1_567/B 0.05fF
C751 POR2X1_212/A POR2X1_212/CTRL2 0.01fF
C752 POR2X1_260/a_16_28# POR2X1_260/A 0.04fF
C753 POR2X1_427/Y POR2X1_763/a_56_344# 0.00fF
C754 POR2X1_71/Y PAND2X1_657/a_76_28# 0.02fF
C755 POR2X1_287/O POR2X1_733/A 0.13fF
C756 PAND2X1_790/CTRL POR2X1_7/A 0.09fF
C757 PAND2X1_432/a_16_344# POR2X1_130/A 0.02fF
C758 POR2X1_265/a_56_344# POR2X1_73/Y 0.00fF
C759 POR2X1_116/A POR2X1_362/A 0.03fF
C760 POR2X1_383/A PAND2X1_271/CTRL 0.01fF
C761 PAND2X1_65/B POR2X1_480/A 0.07fF
C762 POR2X1_65/A PAND2X1_556/B 0.03fF
C763 PAND2X1_23/Y POR2X1_489/B 0.03fF
C764 POR2X1_43/B POR2X1_32/A 0.83fF
C765 POR2X1_368/CTRL2 POR2X1_5/Y 0.01fF
C766 PAND2X1_859/O VDD 0.00fF
C767 POR2X1_718/A VDD 0.14fF
C768 POR2X1_65/A PAND2X1_549/CTRL 0.01fF
C769 PAND2X1_31/CTRL INPUT_6 0.01fF
C770 POR2X1_174/B POR2X1_775/A 0.05fF
C771 POR2X1_355/B PAND2X1_41/B 0.06fF
C772 POR2X1_547/O POR2X1_78/A 0.01fF
C773 PAND2X1_208/O PAND2X1_35/Y 0.02fF
C774 POR2X1_568/A POR2X1_161/CTRL 0.03fF
C775 PAND2X1_667/CTRL2 VDD 0.00fF
C776 POR2X1_381/a_76_344# POR2X1_236/Y 0.09fF
C777 PAND2X1_56/Y PAND2X1_58/A 0.07fF
C778 PAND2X1_9/Y POR2X1_260/A 0.03fF
C779 POR2X1_834/Y POR2X1_648/CTRL2 0.07fF
C780 PAND2X1_733/O POR2X1_7/B 0.04fF
C781 POR2X1_65/A PAND2X1_254/Y 0.03fF
C782 POR2X1_49/Y POR2X1_597/A 0.01fF
C783 PAND2X1_23/Y POR2X1_202/CTRL2 0.00fF
C784 POR2X1_820/B VDD 0.01fF
C785 POR2X1_814/B POR2X1_247/CTRL2 0.00fF
C786 PAND2X1_90/A POR2X1_777/B 0.10fF
C787 POR2X1_814/B PAND2X1_176/CTRL 0.01fF
C788 PAND2X1_73/Y PAND2X1_69/A 0.16fF
C789 POR2X1_669/B POR2X1_73/Y 0.27fF
C790 PAND2X1_204/O PAND2X1_735/Y 0.05fF
C791 POR2X1_495/Y POR2X1_72/B 0.01fF
C792 POR2X1_52/A PAND2X1_192/Y 0.01fF
C793 PAND2X1_73/a_76_28# POR2X1_294/B 0.02fF
C794 POR2X1_821/O POR2X1_236/Y 0.00fF
C795 POR2X1_632/A POR2X1_220/Y 0.00fF
C796 POR2X1_514/a_56_344# PAND2X1_20/A 0.00fF
C797 POR2X1_41/B PAND2X1_192/O 0.05fF
C798 POR2X1_166/m4_208_n4# POR2X1_438/Y 0.12fF
C799 PAND2X1_6/Y PAND2X1_626/O 0.00fF
C800 POR2X1_43/B POR2X1_417/Y 0.05fF
C801 POR2X1_255/CTRL POR2X1_184/Y 0.00fF
C802 POR2X1_614/A POR2X1_806/O 0.01fF
C803 POR2X1_651/Y POR2X1_725/O 0.01fF
C804 POR2X1_43/B POR2X1_419/Y 0.00fF
C805 PAND2X1_63/Y POR2X1_267/A 0.05fF
C806 POR2X1_488/m4_208_n4# PAND2X1_738/Y 0.04fF
C807 POR2X1_65/A POR2X1_488/Y 0.00fF
C808 POR2X1_625/O POR2X1_7/B 0.01fF
C809 PAND2X1_96/B POR2X1_121/B 0.00fF
C810 PAND2X1_115/O PAND2X1_562/B 0.06fF
C811 POR2X1_122/O POR2X1_411/B 0.01fF
C812 POR2X1_422/Y POR2X1_93/A 0.00fF
C813 POR2X1_567/B POR2X1_440/Y 0.05fF
C814 POR2X1_651/Y PAND2X1_72/A 0.78fF
C815 PAND2X1_90/A PAND2X1_65/B 0.13fF
C816 POR2X1_840/B POR2X1_656/m4_208_n4# 0.04fF
C817 POR2X1_22/A POR2X1_12/CTRL2 0.01fF
C818 PAND2X1_453/CTRL POR2X1_511/Y 0.03fF
C819 PAND2X1_6/Y POR2X1_750/B 0.08fF
C820 POR2X1_244/B POR2X1_220/Y 0.03fF
C821 POR2X1_46/Y INPUT_0 0.03fF
C822 POR2X1_74/CTRL POR2X1_23/Y 0.04fF
C823 POR2X1_78/B POR2X1_193/A 0.10fF
C824 PAND2X1_96/B POR2X1_630/A 0.04fF
C825 POR2X1_294/a_16_28# POR2X1_507/A 0.09fF
C826 POR2X1_78/B POR2X1_579/Y 0.03fF
C827 POR2X1_52/A PAND2X1_512/Y 0.01fF
C828 POR2X1_66/B POR2X1_194/O 0.01fF
C829 POR2X1_818/Y POR2X1_260/A 0.03fF
C830 PAND2X1_23/a_16_344# PAND2X1_6/A 0.02fF
C831 POR2X1_197/a_16_28# POR2X1_244/B 0.02fF
C832 POR2X1_278/Y PAND2X1_205/B 0.02fF
C833 POR2X1_16/A PAND2X1_214/CTRL -0.01fF
C834 POR2X1_390/B POR2X1_66/A 0.04fF
C835 POR2X1_22/CTRL2 INPUT_5 0.00fF
C836 POR2X1_634/A POR2X1_711/a_56_344# 0.03fF
C837 POR2X1_590/A PAND2X1_63/B 0.03fF
C838 PAND2X1_488/CTRL2 POR2X1_68/B 0.03fF
C839 POR2X1_40/Y POR2X1_310/a_76_344# 0.00fF
C840 PAND2X1_697/CTRL PAND2X1_65/B 0.01fF
C841 POR2X1_96/A PAND2X1_364/B 0.02fF
C842 POR2X1_466/A PAND2X1_313/O 0.04fF
C843 POR2X1_48/A PAND2X1_563/A 0.04fF
C844 POR2X1_383/A PAND2X1_58/A 0.17fF
C845 POR2X1_467/Y PAND2X1_60/B 0.07fF
C846 POR2X1_57/A POR2X1_666/Y 0.16fF
C847 PAND2X1_641/Y POR2X1_263/Y 0.01fF
C848 PAND2X1_252/m4_208_n4# POR2X1_750/B 0.03fF
C849 PAND2X1_206/B PAND2X1_358/a_76_28# 0.02fF
C850 POR2X1_778/B POR2X1_778/CTRL2 0.03fF
C851 POR2X1_65/A PAND2X1_105/m4_208_n4# 0.07fF
C852 POR2X1_834/Y POR2X1_660/Y 0.00fF
C853 POR2X1_513/B POR2X1_783/B 0.01fF
C854 POR2X1_856/B POR2X1_317/B 0.02fF
C855 PAND2X1_249/a_76_28# POR2X1_591/Y 0.01fF
C856 POR2X1_201/CTRL POR2X1_201/Y 0.01fF
C857 PAND2X1_659/B PAND2X1_658/B 0.04fF
C858 POR2X1_299/Y POR2X1_394/A 0.03fF
C859 POR2X1_204/O VDD 0.00fF
C860 POR2X1_68/A INPUT_0 0.03fF
C861 POR2X1_78/B POR2X1_614/A 0.27fF
C862 POR2X1_616/Y PAND2X1_66/CTRL2 0.01fF
C863 POR2X1_722/A POR2X1_66/A 0.85fF
C864 PAND2X1_15/O POR2X1_260/A 0.09fF
C865 POR2X1_566/A D_GATE_741 0.10fF
C866 PAND2X1_56/Y PAND2X1_309/CTRL2 0.01fF
C867 POR2X1_510/B PAND2X1_41/B 0.03fF
C868 PAND2X1_90/Y POR2X1_736/CTRL 0.27fF
C869 PAND2X1_483/CTRL POR2X1_60/A 0.01fF
C870 POR2X1_65/A POR2X1_165/O 0.01fF
C871 POR2X1_43/B PAND2X1_35/Y 0.08fF
C872 POR2X1_48/A POR2X1_320/CTRL2 0.03fF
C873 POR2X1_20/B POR2X1_39/B 1.52fF
C874 PAND2X1_735/Y POR2X1_56/Y 0.46fF
C875 PAND2X1_55/Y POR2X1_205/Y 0.03fF
C876 POR2X1_72/B PAND2X1_723/A 0.07fF
C877 POR2X1_506/O POR2X1_506/B 0.00fF
C878 POR2X1_41/B PAND2X1_845/CTRL2 0.00fF
C879 PAND2X1_702/CTRL VDD 0.00fF
C880 POR2X1_333/A POR2X1_326/O 0.16fF
C881 POR2X1_57/A VDD 4.31fF
C882 POR2X1_725/a_76_344# POR2X1_712/Y 0.00fF
C883 PAND2X1_213/Y PAND2X1_543/O 0.02fF
C884 POR2X1_186/Y POR2X1_151/CTRL 0.04fF
C885 PAND2X1_55/Y POR2X1_363/O 0.06fF
C886 PAND2X1_232/CTRL PAND2X1_41/B 0.01fF
C887 POR2X1_68/B POR2X1_401/B 0.00fF
C888 POR2X1_133/CTRL POR2X1_93/A 0.01fF
C889 PAND2X1_94/A POR2X1_752/Y 0.03fF
C890 POR2X1_537/Y POR2X1_858/O 0.01fF
C891 POR2X1_368/Y POR2X1_293/Y 0.02fF
C892 POR2X1_808/A POR2X1_260/A 0.03fF
C893 POR2X1_814/B POR2X1_360/a_16_28# 0.02fF
C894 POR2X1_348/A POR2X1_348/a_16_28# 0.11fF
C895 POR2X1_584/CTRL POR2X1_42/Y 0.08fF
C896 POR2X1_100/O POR2X1_243/Y 0.03fF
C897 POR2X1_41/B POR2X1_248/O 0.05fF
C898 POR2X1_346/B POR2X1_194/A 0.02fF
C899 POR2X1_254/Y POR2X1_205/A 0.01fF
C900 POR2X1_119/Y POR2X1_609/Y 0.14fF
C901 PAND2X1_55/Y POR2X1_402/A 0.44fF
C902 PAND2X1_80/O PAND2X1_111/B 0.02fF
C903 POR2X1_719/CTRL2 POR2X1_502/A 0.02fF
C904 PAND2X1_350/O INPUT_0 0.06fF
C905 PAND2X1_550/B PAND2X1_712/B 0.01fF
C906 POR2X1_198/O POR2X1_68/A 0.02fF
C907 POR2X1_578/Y POR2X1_577/CTRL 0.00fF
C908 PAND2X1_58/A PAND2X1_71/Y 0.01fF
C909 PAND2X1_6/Y POR2X1_84/O 0.16fF
C910 POR2X1_41/B PAND2X1_270/CTRL2 0.04fF
C911 PAND2X1_631/O POR2X1_55/Y 0.01fF
C912 PAND2X1_220/O PAND2X1_566/Y 0.00fF
C913 PAND2X1_48/B POR2X1_638/Y 0.92fF
C914 POR2X1_377/CTRL2 D_INPUT_1 0.15fF
C915 POR2X1_740/Y PAND2X1_111/a_56_28# 0.00fF
C916 POR2X1_741/Y PAND2X1_111/a_16_344# 0.01fF
C917 PAND2X1_48/B POR2X1_196/Y 0.03fF
C918 POR2X1_43/B POR2X1_184/Y 0.05fF
C919 POR2X1_102/Y PAND2X1_141/CTRL2 0.01fF
C920 POR2X1_13/A POR2X1_597/O 0.03fF
C921 POR2X1_725/Y VDD -0.00fF
C922 POR2X1_254/Y POR2X1_366/A 0.12fF
C923 PAND2X1_110/O PAND2X1_32/B 0.07fF
C924 PAND2X1_390/Y POR2X1_129/Y 0.00fF
C925 POR2X1_584/Y VDD 0.04fF
C926 POR2X1_809/A POR2X1_605/B 0.24fF
C927 POR2X1_414/O POR2X1_4/Y 0.01fF
C928 POR2X1_140/B POR2X1_140/A 0.02fF
C929 POR2X1_315/CTRL2 POR2X1_90/Y 0.00fF
C930 PAND2X1_651/Y POR2X1_43/B 0.07fF
C931 POR2X1_52/A POR2X1_823/Y 0.01fF
C932 POR2X1_860/a_16_28# POR2X1_860/A 0.03fF
C933 POR2X1_54/Y POR2X1_8/CTRL 0.01fF
C934 POR2X1_566/A POR2X1_507/CTRL2 0.13fF
C935 POR2X1_16/A POR2X1_689/O 0.02fF
C936 POR2X1_7/B PAND2X1_347/a_76_28# 0.01fF
C937 PAND2X1_56/Y PAND2X1_96/B 0.05fF
C938 PAND2X1_96/B POR2X1_795/B 0.07fF
C939 POR2X1_543/A POR2X1_543/a_16_28# 0.03fF
C940 PAND2X1_834/CTRL POR2X1_37/Y 0.01fF
C941 POR2X1_501/CTRL POR2X1_573/A 0.01fF
C942 PAND2X1_117/CTRL2 POR2X1_383/A 0.00fF
C943 POR2X1_65/A PAND2X1_358/A 0.07fF
C944 PAND2X1_476/A POR2X1_14/Y 0.02fF
C945 PAND2X1_41/B POR2X1_195/CTRL2 0.03fF
C946 POR2X1_272/Y PAND2X1_301/CTRL 0.01fF
C947 POR2X1_741/a_16_28# POR2X1_741/B -0.00fF
C948 PAND2X1_111/a_16_344# PAND2X1_32/B 0.01fF
C949 PAND2X1_220/CTRL2 PAND2X1_388/Y 0.01fF
C950 PAND2X1_6/Y PAND2X1_275/m4_208_n4# 0.07fF
C951 PAND2X1_243/B PAND2X1_402/B 0.02fF
C952 POR2X1_614/A PAND2X1_495/CTRL2 0.04fF
C953 POR2X1_57/A PAND2X1_850/CTRL 0.01fF
C954 POR2X1_596/O VDD 0.00fF
C955 PAND2X1_95/B PAND2X1_60/B 0.02fF
C956 POR2X1_66/A PAND2X1_529/O 0.05fF
C957 PAND2X1_563/B POR2X1_394/A 0.04fF
C958 POR2X1_43/B PAND2X1_844/B 0.05fF
C959 POR2X1_814/B POR2X1_703/CTRL 0.05fF
C960 POR2X1_65/A PAND2X1_779/CTRL 0.00fF
C961 PAND2X1_798/B POR2X1_91/Y 0.03fF
C962 POR2X1_123/A PAND2X1_132/O 0.01fF
C963 POR2X1_111/Y VDD 0.35fF
C964 POR2X1_41/B POR2X1_310/Y 0.06fF
C965 POR2X1_7/B PAND2X1_112/CTRL 0.00fF
C966 PAND2X1_844/Y PAND2X1_244/B 0.01fF
C967 POR2X1_502/A INPUT_1 0.03fF
C968 POR2X1_96/A POR2X1_96/CTRL 0.01fF
C969 PAND2X1_723/Y PAND2X1_853/B 0.03fF
C970 PAND2X1_182/A POR2X1_176/Y 0.00fF
C971 PAND2X1_675/A PAND2X1_388/Y 0.01fF
C972 POR2X1_174/O POR2X1_192/Y 0.04fF
C973 POR2X1_68/A PAND2X1_393/CTRL2 0.02fF
C974 PAND2X1_6/Y PAND2X1_424/O 0.17fF
C975 POR2X1_266/A POR2X1_5/Y 0.05fF
C976 PAND2X1_652/CTRL PAND2X1_557/A 0.01fF
C977 POR2X1_394/A PAND2X1_738/a_76_28# 0.02fF
C978 POR2X1_559/A VDD 1.57fF
C979 PAND2X1_299/O POR2X1_188/Y 0.07fF
C980 PAND2X1_20/A PAND2X1_136/a_16_344# 0.02fF
C981 POR2X1_271/A POR2X1_256/CTRL 0.00fF
C982 POR2X1_468/CTRL2 POR2X1_444/Y 0.02fF
C983 PAND2X1_90/Y POR2X1_383/CTRL2 0.01fF
C984 PAND2X1_251/a_56_28# PAND2X1_52/B 0.00fF
C985 POR2X1_137/Y D_INPUT_1 0.03fF
C986 PAND2X1_785/Y POR2X1_394/A 1.22fF
C987 POR2X1_149/Y POR2X1_260/A 0.03fF
C988 POR2X1_710/O POR2X1_713/B 0.18fF
C989 POR2X1_66/B D_INPUT_4 1.07fF
C990 PAND2X1_603/O PAND2X1_72/A 0.04fF
C991 POR2X1_62/Y PAND2X1_8/Y 0.03fF
C992 INPUT_0 POR2X1_371/CTRL 0.02fF
C993 PAND2X1_659/B PAND2X1_657/B 0.00fF
C994 PAND2X1_140/A PAND2X1_113/CTRL 0.01fF
C995 POR2X1_804/A POR2X1_274/B 0.05fF
C996 POR2X1_750/B POR2X1_632/Y 0.05fF
C997 POR2X1_383/A PAND2X1_96/B 0.78fF
C998 POR2X1_220/B POR2X1_161/a_16_28# 0.02fF
C999 POR2X1_725/Y PAND2X1_32/B 0.07fF
C1000 POR2X1_295/O POR2X1_77/Y 0.07fF
C1001 POR2X1_255/O PAND2X1_840/Y 0.01fF
C1002 POR2X1_130/A POR2X1_557/O 0.01fF
C1003 POR2X1_13/A PAND2X1_851/CTRL 0.01fF
C1004 POR2X1_537/Y POR2X1_220/Y 0.03fF
C1005 POR2X1_13/A POR2X1_595/a_76_344# 0.02fF
C1006 POR2X1_753/Y POR2X1_90/CTRL2 0.09fF
C1007 POR2X1_754/Y POR2X1_90/O 0.08fF
C1008 PAND2X1_865/Y PAND2X1_580/B 0.66fF
C1009 POR2X1_16/A PAND2X1_578/A 0.01fF
C1010 POR2X1_276/Y POR2X1_501/B 0.03fF
C1011 POR2X1_416/B PAND2X1_733/CTRL 0.07fF
C1012 PAND2X1_232/CTRL2 POR2X1_68/B 0.03fF
C1013 PAND2X1_804/O PAND2X1_860/A 0.03fF
C1014 PAND2X1_139/CTRL2 POR2X1_13/A 0.01fF
C1015 INPUT_1 POR2X1_409/O 0.02fF
C1016 PAND2X1_640/B PAND2X1_403/O 0.12fF
C1017 POR2X1_313/Y POR2X1_90/Y 0.02fF
C1018 POR2X1_509/CTRL2 PAND2X1_41/B 0.10fF
C1019 VDD POR2X1_589/CTRL 0.00fF
C1020 POR2X1_833/A D_INPUT_1 0.04fF
C1021 INPUT_0 PAND2X1_517/O 0.14fF
C1022 POR2X1_750/B PAND2X1_52/B 0.31fF
C1023 POR2X1_517/CTRL2 POR2X1_13/A 0.01fF
C1024 PAND2X1_562/a_16_344# POR2X1_394/A 0.02fF
C1025 PAND2X1_824/B POR2X1_631/B 0.02fF
C1026 POR2X1_639/Y POR2X1_260/A 0.03fF
C1027 POR2X1_578/Y POR2X1_191/Y 0.05fF
C1028 POR2X1_572/B POR2X1_294/A 0.03fF
C1029 POR2X1_222/A POR2X1_569/A 0.07fF
C1030 POR2X1_141/O POR2X1_343/Y 0.00fF
C1031 POR2X1_559/A PAND2X1_32/B 0.03fF
C1032 POR2X1_294/B POR2X1_4/Y 0.22fF
C1033 PAND2X1_849/B POR2X1_7/A 0.06fF
C1034 PAND2X1_476/A POR2X1_55/Y 0.02fF
C1035 POR2X1_502/Y POR2X1_350/O 0.01fF
C1036 POR2X1_62/Y PAND2X1_341/a_76_28# 0.01fF
C1037 PAND2X1_643/A POR2X1_42/Y 0.03fF
C1038 POR2X1_685/A POR2X1_687/A 0.05fF
C1039 POR2X1_447/B PAND2X1_625/CTRL 0.08fF
C1040 POR2X1_789/A POR2X1_294/A 0.01fF
C1041 POR2X1_493/B POR2X1_383/A 0.00fF
C1042 POR2X1_7/A PAND2X1_154/a_76_28# 0.01fF
C1043 POR2X1_217/CTRL2 PAND2X1_72/A 0.04fF
C1044 POR2X1_614/A POR2X1_294/A 0.07fF
C1045 PAND2X1_483/O POR2X1_7/A 0.11fF
C1046 POR2X1_10/CTRL PAND2X1_63/B 0.01fF
C1047 POR2X1_684/Y POR2X1_683/Y 0.00fF
C1048 PAND2X1_96/B PAND2X1_71/Y 0.89fF
C1049 PAND2X1_96/B POR2X1_332/m4_208_n4# 0.08fF
C1050 PAND2X1_501/O PAND2X1_735/Y 0.09fF
C1051 PAND2X1_860/A POR2X1_72/B 0.05fF
C1052 POR2X1_81/A PAND2X1_658/A 0.03fF
C1053 POR2X1_848/A POR2X1_846/Y 0.07fF
C1054 POR2X1_659/A POR2X1_657/Y 0.04fF
C1055 POR2X1_804/A POR2X1_512/O 0.02fF
C1056 POR2X1_596/A PAND2X1_48/A 0.03fF
C1057 POR2X1_38/B POR2X1_294/A 0.00fF
C1058 POR2X1_560/O POR2X1_844/B 0.00fF
C1059 POR2X1_687/A POR2X1_260/A 0.01fF
C1060 PAND2X1_385/CTRL2 POR2X1_711/Y 0.02fF
C1061 POR2X1_703/A POR2X1_543/O 0.02fF
C1062 PAND2X1_172/O POR2X1_353/A 0.07fF
C1063 POR2X1_722/CTRL2 PAND2X1_60/B 0.01fF
C1064 POR2X1_41/Y POR2X1_73/Y 0.03fF
C1065 INPUT_0 POR2X1_138/A 0.09fF
C1066 POR2X1_316/Y POR2X1_56/Y 0.03fF
C1067 POR2X1_46/Y PAND2X1_327/a_76_28# 0.02fF
C1068 POR2X1_809/A POR2X1_855/B 0.04fF
C1069 POR2X1_446/B POR2X1_222/CTRL 0.01fF
C1070 POR2X1_648/Y PAND2X1_58/A 0.03fF
C1071 PAND2X1_98/a_16_344# POR2X1_93/Y 0.02fF
C1072 POR2X1_48/A POR2X1_20/B 2.60fF
C1073 POR2X1_612/O POR2X1_612/Y 0.02fF
C1074 POR2X1_351/Y POR2X1_568/B 0.01fF
C1075 POR2X1_81/A POR2X1_73/Y 0.03fF
C1076 PAND2X1_494/a_16_344# POR2X1_383/Y 0.01fF
C1077 POR2X1_324/a_76_344# POR2X1_568/Y 0.03fF
C1078 POR2X1_348/a_16_28# POR2X1_334/Y 0.07fF
C1079 POR2X1_673/Y POR2X1_559/A 1.62fF
C1080 PAND2X1_61/Y POR2X1_9/Y 0.03fF
C1081 POR2X1_343/Y POR2X1_833/a_76_344# 0.10fF
C1082 POR2X1_257/A PAND2X1_205/A 0.03fF
C1083 POR2X1_43/B PAND2X1_858/B 0.03fF
C1084 POR2X1_118/CTRL2 POR2X1_77/Y 0.00fF
C1085 POR2X1_63/Y POR2X1_263/Y 0.14fF
C1086 POR2X1_102/Y PAND2X1_449/CTRL2 0.00fF
C1087 PAND2X1_82/a_56_28# POR2X1_84/A 0.00fF
C1088 POR2X1_687/CTRL2 POR2X1_452/Y 0.01fF
C1089 POR2X1_394/A PAND2X1_348/A 0.01fF
C1090 POR2X1_327/Y POR2X1_244/Y 0.00fF
C1091 PAND2X1_717/A POR2X1_423/Y 0.03fF
C1092 PAND2X1_59/O D_INPUT_4 0.17fF
C1093 POR2X1_66/B POR2X1_66/CTRL 0.01fF
C1094 PAND2X1_233/O INPUT_0 0.03fF
C1095 POR2X1_184/O POR2X1_91/Y 0.01fF
C1096 PAND2X1_619/CTRL POR2X1_29/A 0.01fF
C1097 POR2X1_83/B PAND2X1_201/a_16_344# 0.00fF
C1098 POR2X1_248/O POR2X1_77/Y 0.01fF
C1099 POR2X1_311/Y POR2X1_150/Y 0.03fF
C1100 POR2X1_16/A POR2X1_397/CTRL2 0.01fF
C1101 POR2X1_416/B PAND2X1_324/a_16_344# 0.01fF
C1102 POR2X1_451/A INPUT_5 0.01fF
C1103 POR2X1_192/CTRL POR2X1_191/Y 0.09fF
C1104 POR2X1_192/O POR2X1_192/B 0.01fF
C1105 POR2X1_394/A POR2X1_300/Y 0.05fF
C1106 PAND2X1_39/B POR2X1_296/B 15.75fF
C1107 POR2X1_293/Y POR2X1_310/CTRL2 0.03fF
C1108 PAND2X1_645/Y PAND2X1_644/Y 1.08fF
C1109 POR2X1_81/A PAND2X1_244/B 0.01fF
C1110 POR2X1_24/Y POR2X1_29/A 0.01fF
C1111 POR2X1_866/A POR2X1_807/O 0.08fF
C1112 POR2X1_49/Y PAND2X1_447/O 0.02fF
C1113 POR2X1_814/A POR2X1_480/A 0.10fF
C1114 POR2X1_814/B POR2X1_621/a_16_28# 0.01fF
C1115 POR2X1_460/Y POR2X1_752/Y 0.02fF
C1116 PAND2X1_47/B POR2X1_635/A 0.01fF
C1117 POR2X1_77/CTRL2 POR2X1_14/Y 0.03fF
C1118 PAND2X1_43/CTRL POR2X1_330/Y 0.02fF
C1119 PAND2X1_366/a_16_344# PAND2X1_354/Y 0.01fF
C1120 PAND2X1_424/CTRL PAND2X1_72/A 0.01fF
C1121 POR2X1_83/A POR2X1_825/Y 0.00fF
C1122 POR2X1_99/CTRL PAND2X1_65/Y 0.00fF
C1123 PAND2X1_224/CTRL POR2X1_578/Y 0.11fF
C1124 POR2X1_169/A POR2X1_704/a_16_28# 0.02fF
C1125 POR2X1_65/A POR2X1_441/Y 0.06fF
C1126 PAND2X1_631/A POR2X1_394/A 0.10fF
C1127 POR2X1_612/Y POR2X1_413/O 0.05fF
C1128 POR2X1_135/a_56_344# POR2X1_394/A 0.03fF
C1129 POR2X1_567/B POR2X1_590/A 0.09fF
C1130 POR2X1_77/Y POR2X1_310/Y 0.02fF
C1131 POR2X1_260/B POR2X1_375/Y 0.00fF
C1132 POR2X1_811/a_16_28# POR2X1_811/A 0.03fF
C1133 POR2X1_422/a_16_28# POR2X1_422/Y 0.01fF
C1134 POR2X1_222/A PAND2X1_72/A 0.03fF
C1135 PAND2X1_35/A POR2X1_94/A 0.01fF
C1136 PAND2X1_809/A PAND2X1_809/O 0.02fF
C1137 PAND2X1_653/m4_208_n4# POR2X1_760/A 0.08fF
C1138 PAND2X1_303/Y POR2X1_39/B 0.03fF
C1139 POR2X1_298/Y POR2X1_32/A 0.01fF
C1140 PAND2X1_90/A POR2X1_814/A 0.04fF
C1141 POR2X1_257/A PAND2X1_76/Y 0.03fF
C1142 POR2X1_669/B POR2X1_753/Y 0.10fF
C1143 PAND2X1_678/O VDD 0.00fF
C1144 POR2X1_760/A PAND2X1_364/B 1.73fF
C1145 PAND2X1_628/CTRL POR2X1_532/A 0.01fF
C1146 POR2X1_455/a_56_344# POR2X1_341/A 0.00fF
C1147 POR2X1_37/CTRL D_INPUT_0 0.01fF
C1148 POR2X1_686/A POR2X1_260/B 0.01fF
C1149 PAND2X1_20/A POR2X1_296/B 0.14fF
C1150 POR2X1_37/Y PAND2X1_390/Y 0.03fF
C1151 POR2X1_417/Y POR2X1_298/Y 0.01fF
C1152 PAND2X1_255/CTRL2 PAND2X1_60/B 0.03fF
C1153 PAND2X1_444/CTRL POR2X1_236/Y 0.01fF
C1154 POR2X1_667/CTRL2 POR2X1_73/Y 0.02fF
C1155 POR2X1_730/Y POR2X1_863/A 0.03fF
C1156 PAND2X1_141/O POR2X1_39/B 0.05fF
C1157 POR2X1_416/B PAND2X1_716/B 0.03fF
C1158 PAND2X1_93/B PAND2X1_85/Y 0.01fF
C1159 POR2X1_63/Y PAND2X1_215/B 0.02fF
C1160 POR2X1_764/a_16_28# POR2X1_40/Y 0.01fF
C1161 POR2X1_220/CTRL POR2X1_220/Y 0.00fF
C1162 POR2X1_413/A POR2X1_20/B 0.09fF
C1163 POR2X1_590/A POR2X1_391/A 0.11fF
C1164 PAND2X1_817/CTRL2 POR2X1_750/B 0.02fF
C1165 PAND2X1_319/B PAND2X1_717/A 0.03fF
C1166 POR2X1_814/B POR2X1_296/B 0.13fF
C1167 POR2X1_862/A POR2X1_121/Y 0.08fF
C1168 POR2X1_188/A POR2X1_830/CTRL2 0.01fF
C1169 POR2X1_84/A PAND2X1_57/B 0.03fF
C1170 POR2X1_56/a_16_28# POR2X1_423/Y 0.02fF
C1171 PAND2X1_571/A INPUT_0 0.03fF
C1172 POR2X1_467/Y POR2X1_750/B 0.68fF
C1173 PAND2X1_847/O POR2X1_4/Y 0.01fF
C1174 POR2X1_274/O POR2X1_325/A 0.01fF
C1175 POR2X1_298/a_56_344# POR2X1_46/Y 0.03fF
C1176 POR2X1_792/O PAND2X1_90/Y 0.03fF
C1177 PAND2X1_666/O POR2X1_130/A 0.03fF
C1178 POR2X1_54/Y POR2X1_415/Y 0.05fF
C1179 PAND2X1_246/CTRL POR2X1_205/A 0.03fF
C1180 PAND2X1_9/Y POR2X1_204/O 0.16fF
C1181 POR2X1_63/Y PAND2X1_6/A 0.02fF
C1182 POR2X1_142/a_16_28# POR2X1_49/Y 0.05fF
C1183 POR2X1_106/a_16_28# POR2X1_106/Y 0.03fF
C1184 POR2X1_266/O POR2X1_294/B 0.02fF
C1185 POR2X1_296/B POR2X1_325/A 0.03fF
C1186 POR2X1_327/CTRL POR2X1_558/B 0.00fF
C1187 POR2X1_78/B POR2X1_590/A 0.19fF
C1188 POR2X1_846/a_76_344# POR2X1_129/Y 0.00fF
C1189 PAND2X1_236/a_16_344# POR2X1_29/A 0.03fF
C1190 POR2X1_150/Y POR2X1_38/Y 0.03fF
C1191 POR2X1_96/A POR2X1_626/O 0.18fF
C1192 POR2X1_66/B POR2X1_555/A 0.03fF
C1193 POR2X1_294/Y PAND2X1_58/a_76_28# 0.02fF
C1194 POR2X1_496/Y POR2X1_516/B 0.07fF
C1195 PAND2X1_462/CTRL2 POR2X1_416/B 0.01fF
C1196 POR2X1_654/B POR2X1_734/A 0.07fF
C1197 POR2X1_232/CTRL POR2X1_37/Y 0.03fF
C1198 POR2X1_808/A POR2X1_718/A 0.02fF
C1199 POR2X1_632/O POR2X1_222/Y 0.01fF
C1200 POR2X1_82/O POR2X1_14/Y 0.01fF
C1201 POR2X1_311/Y PAND2X1_553/A 0.00fF
C1202 PAND2X1_5/O INPUT_3 0.01fF
C1203 POR2X1_811/B VDD 0.35fF
C1204 POR2X1_186/Y PAND2X1_321/CTRL2 0.17fF
C1205 PAND2X1_58/A INPUT_0 0.07fF
C1206 D_INPUT_5 POR2X1_638/Y 0.02fF
C1207 POR2X1_181/CTRL POR2X1_181/A 0.01fF
C1208 PAND2X1_831/Y POR2X1_411/B 0.87fF
C1209 POR2X1_49/Y POR2X1_847/B 0.03fF
C1210 POR2X1_41/B POR2X1_225/CTRL 0.03fF
C1211 POR2X1_78/A PAND2X1_89/CTRL2 0.03fF
C1212 PAND2X1_263/O POR2X1_94/A 0.19fF
C1213 POR2X1_497/O PAND2X1_501/B 0.01fF
C1214 PAND2X1_94/A PAND2X1_699/CTRL2 0.00fF
C1215 POR2X1_186/Y POR2X1_213/B 0.05fF
C1216 POR2X1_296/B POR2X1_513/B 0.10fF
C1217 PAND2X1_853/CTRL POR2X1_23/Y 0.01fF
C1218 POR2X1_227/A POR2X1_566/B 0.03fF
C1219 PAND2X1_423/m4_208_n4# POR2X1_330/Y 0.06fF
C1220 POR2X1_852/CTRL2 POR2X1_852/B 0.05fF
C1221 POR2X1_493/A PAND2X1_519/O 0.01fF
C1222 PAND2X1_118/CTRL POR2X1_66/A 0.05fF
C1223 POR2X1_43/Y POR2X1_39/B 0.19fF
C1224 POR2X1_102/Y POR2X1_46/Y 0.15fF
C1225 POR2X1_556/A POR2X1_218/CTRL2 0.01fF
C1226 POR2X1_558/B POR2X1_218/A 0.19fF
C1227 POR2X1_20/B PAND2X1_840/O 0.07fF
C1228 PAND2X1_732/CTRL2 POR2X1_763/Y 0.05fF
C1229 POR2X1_297/CTRL PAND2X1_347/Y 0.01fF
C1230 PAND2X1_333/CTRL POR2X1_5/Y 0.03fF
C1231 PAND2X1_217/B PAND2X1_84/Y 0.05fF
C1232 POR2X1_265/m4_208_n4# POR2X1_406/m4_208_n4# 0.05fF
C1233 D_INPUT_0 POR2X1_565/CTRL 0.01fF
C1234 POR2X1_115/CTRL2 POR2X1_141/Y 0.00fF
C1235 POR2X1_311/Y PAND2X1_364/B 1.49fF
C1236 POR2X1_681/CTRL2 POR2X1_153/Y 0.03fF
C1237 PAND2X1_56/CTRL POR2X1_330/Y 0.28fF
C1238 POR2X1_83/B PAND2X1_364/O 0.04fF
C1239 POR2X1_389/A PAND2X1_609/CTRL 0.00fF
C1240 POR2X1_407/A POR2X1_644/B 0.10fF
C1241 POR2X1_555/B POR2X1_740/Y 0.05fF
C1242 POR2X1_632/O POR2X1_532/A 0.02fF
C1243 POR2X1_76/Y POR2X1_330/Y 0.03fF
C1244 POR2X1_444/a_76_344# POR2X1_568/Y 0.10fF
C1245 PAND2X1_56/CTRL2 POR2X1_593/B 0.01fF
C1246 POR2X1_293/a_16_28# POR2X1_5/Y 0.03fF
C1247 POR2X1_428/Y PAND2X1_710/CTRL2 0.01fF
C1248 POR2X1_655/A PAND2X1_60/B 0.03fF
C1249 POR2X1_315/Y POR2X1_257/A 0.10fF
C1250 PAND2X1_473/B PAND2X1_736/O 0.01fF
C1251 POR2X1_5/Y POR2X1_372/A 0.01fF
C1252 POR2X1_590/A PAND2X1_530/a_16_344# 0.01fF
C1253 POR2X1_56/B POR2X1_748/A 0.61fF
C1254 POR2X1_683/Y POR2X1_32/A 0.03fF
C1255 POR2X1_278/Y PAND2X1_61/Y 0.05fF
C1256 PAND2X1_20/A PAND2X1_79/CTRL2 0.03fF
C1257 POR2X1_41/B POR2X1_423/Y 0.12fF
C1258 POR2X1_242/O POR2X1_578/Y 0.01fF
C1259 POR2X1_558/O PAND2X1_20/A 0.01fF
C1260 POR2X1_96/A POR2X1_46/a_16_28# 0.07fF
C1261 PAND2X1_390/Y POR2X1_293/Y 0.03fF
C1262 PAND2X1_57/B PAND2X1_65/Y 0.03fF
C1263 PAND2X1_48/B POR2X1_141/Y 0.03fF
C1264 PAND2X1_738/Y PAND2X1_180/O 0.10fF
C1265 PAND2X1_53/O PAND2X1_48/A 0.07fF
C1266 PAND2X1_644/Y POR2X1_755/Y 0.03fF
C1267 PAND2X1_644/CTRL2 POR2X1_40/Y 0.01fF
C1268 PAND2X1_671/O POR2X1_54/Y 0.02fF
C1269 PAND2X1_859/a_76_28# INPUT_0 0.03fF
C1270 PAND2X1_95/B POR2X1_750/B 0.01fF
C1271 PAND2X1_13/CTRL2 POR2X1_294/B 0.01fF
C1272 PAND2X1_84/Y VDD 0.29fF
C1273 PAND2X1_667/O INPUT_0 0.16fF
C1274 PAND2X1_245/CTRL POR2X1_68/B 0.01fF
C1275 POR2X1_338/O POR2X1_567/B 0.08fF
C1276 PAND2X1_52/Y POR2X1_294/B 0.03fF
C1277 POR2X1_619/Y POR2X1_29/A 0.73fF
C1278 POR2X1_564/Y POR2X1_78/B 0.07fF
C1279 POR2X1_702/B POR2X1_294/B 0.00fF
C1280 POR2X1_672/A POR2X1_40/Y 0.05fF
C1281 POR2X1_810/O POR2X1_750/B 0.01fF
C1282 POR2X1_843/CTRL PAND2X1_60/B 0.01fF
C1283 POR2X1_66/A PAND2X1_63/B 4.96fF
C1284 POR2X1_62/Y POR2X1_20/B 0.03fF
C1285 POR2X1_41/B POR2X1_368/CTRL 0.04fF
C1286 PAND2X1_771/Y PAND2X1_569/B 0.29fF
C1287 POR2X1_137/Y POR2X1_78/A 0.02fF
C1288 PAND2X1_817/a_56_28# D_INPUT_1 0.00fF
C1289 PAND2X1_771/Y PAND2X1_578/a_16_344# 0.07fF
C1290 POR2X1_461/CTRL2 POR2X1_793/A 0.15fF
C1291 POR2X1_220/Y POR2X1_483/B 0.01fF
C1292 PAND2X1_216/B PAND2X1_267/Y 0.02fF
C1293 POR2X1_614/A POR2X1_94/A 0.05fF
C1294 POR2X1_403/CTRL2 POR2X1_35/Y 0.09fF
C1295 PAND2X1_808/Y POR2X1_488/O 0.01fF
C1296 PAND2X1_540/O POR2X1_183/Y 0.00fF
C1297 POR2X1_247/CTRL2 VDD 0.00fF
C1298 PAND2X1_658/O POR2X1_816/A 0.02fF
C1299 PAND2X1_96/B POR2X1_634/O 0.02fF
C1300 POR2X1_669/B PAND2X1_656/A 0.03fF
C1301 POR2X1_344/O PAND2X1_6/Y 0.07fF
C1302 POR2X1_120/CTRL POR2X1_294/B 0.01fF
C1303 POR2X1_748/A POR2X1_748/O 0.19fF
C1304 POR2X1_362/Y PAND2X1_106/CTRL2 0.01fF
C1305 PAND2X1_632/B POR2X1_482/CTRL 0.01fF
C1306 POR2X1_734/A POR2X1_705/CTRL 0.10fF
C1307 POR2X1_660/CTRL2 POR2X1_725/Y 0.04fF
C1308 VDD POR2X1_783/B 0.26fF
C1309 PAND2X1_812/O PAND2X1_805/A 0.02fF
C1310 POR2X1_423/Y POR2X1_256/Y 0.04fF
C1311 POR2X1_82/O POR2X1_55/Y 0.17fF
C1312 PAND2X1_472/A PAND2X1_721/CTRL2 0.02fF
C1313 POR2X1_119/Y POR2X1_63/Y 0.05fF
C1314 POR2X1_83/O D_INPUT_0 0.08fF
C1315 PAND2X1_669/O POR2X1_750/Y 0.01fF
C1316 PAND2X1_658/A PAND2X1_499/Y 0.75fF
C1317 POR2X1_48/A PAND2X1_715/B 0.01fF
C1318 POR2X1_71/Y PAND2X1_735/Y 0.07fF
C1319 POR2X1_94/A POR2X1_38/B 0.12fF
C1320 PAND2X1_469/B PAND2X1_787/a_76_28# 0.04fF
C1321 PAND2X1_831/Y POR2X1_271/Y 0.04fF
C1322 POR2X1_502/A POR2X1_794/m4_208_n4# 0.12fF
C1323 POR2X1_61/Y POR2X1_219/CTRL2 0.03fF
C1324 POR2X1_669/B PAND2X1_124/CTRL2 0.01fF
C1325 POR2X1_836/A POR2X1_854/B 0.05fF
C1326 POR2X1_61/Y PAND2X1_69/A 0.01fF
C1327 PAND2X1_585/a_16_344# PAND2X1_60/B 0.02fF
C1328 PAND2X1_23/Y POR2X1_192/Y 0.09fF
C1329 PAND2X1_48/B POR2X1_220/Y 0.06fF
C1330 POR2X1_416/B POR2X1_250/Y 10.29fF
C1331 POR2X1_197/CTRL2 PAND2X1_6/Y 0.00fF
C1332 PAND2X1_417/O POR2X1_169/A 0.09fF
C1333 POR2X1_40/Y POR2X1_387/Y 0.14fF
C1334 POR2X1_65/A PAND2X1_640/a_56_28# 0.00fF
C1335 POR2X1_43/B POR2X1_821/CTRL2 0.01fF
C1336 POR2X1_274/Y POR2X1_532/A 0.06fF
C1337 POR2X1_232/CTRL POR2X1_293/Y 0.01fF
C1338 POR2X1_329/A POR2X1_522/O 0.01fF
C1339 POR2X1_10/CTRL POR2X1_32/A 0.01fF
C1340 POR2X1_43/Y POR2X1_827/O 0.00fF
C1341 PAND2X1_478/CTRL PAND2X1_480/B 0.07fF
C1342 POR2X1_483/A POR2X1_804/A 0.01fF
C1343 POR2X1_558/B POR2X1_557/B 0.03fF
C1344 POR2X1_83/B POR2X1_59/CTRL2 0.00fF
C1345 PAND2X1_48/B POR2X1_404/Y 0.03fF
C1346 PAND2X1_651/Y PAND2X1_84/O 0.42fF
C1347 POR2X1_637/A PAND2X1_60/B 0.03fF
C1348 POR2X1_51/A POR2X1_43/B 0.00fF
C1349 PAND2X1_564/O PAND2X1_551/Y -0.00fF
C1350 PAND2X1_499/Y POR2X1_73/Y 0.05fF
C1351 POR2X1_84/CTRL2 POR2X1_294/B 0.01fF
C1352 PAND2X1_222/B POR2X1_250/A 0.03fF
C1353 PAND2X1_605/O POR2X1_604/Y 0.04fF
C1354 POR2X1_376/B POR2X1_376/A 0.00fF
C1355 POR2X1_334/B POR2X1_137/CTRL 0.05fF
C1356 POR2X1_537/Y POR2X1_841/B 0.03fF
C1357 PAND2X1_73/Y PAND2X1_413/CTRL2 0.01fF
C1358 PAND2X1_104/CTRL2 INPUT_1 0.00fF
C1359 PAND2X1_286/a_16_344# PAND2X1_568/B 0.01fF
C1360 VDD POR2X1_594/A 0.26fF
C1361 PAND2X1_600/O POR2X1_294/A 0.01fF
C1362 PAND2X1_418/O PAND2X1_52/B 0.06fF
C1363 PAND2X1_468/O PAND2X1_469/B 0.02fF
C1364 POR2X1_49/Y POR2X1_315/Y 1.15fF
C1365 POR2X1_46/Y POR2X1_531/Y 0.02fF
C1366 PAND2X1_96/B INPUT_0 0.37fF
C1367 D_INPUT_0 PAND2X1_48/A 0.10fF
C1368 POR2X1_29/A POR2X1_720/CTRL 0.03fF
C1369 PAND2X1_480/CTRL2 PAND2X1_478/B 0.01fF
C1370 POR2X1_861/CTRL2 POR2X1_572/B 0.01fF
C1371 POR2X1_52/A POR2X1_305/Y 0.04fF
C1372 PAND2X1_218/A PAND2X1_364/B 0.03fF
C1373 POR2X1_52/A POR2X1_823/O 0.02fF
C1374 POR2X1_685/CTRL2 POR2X1_729/Y 0.02fF
C1375 POR2X1_407/A PAND2X1_498/CTRL 0.01fF
C1376 PAND2X1_564/B POR2X1_394/A 0.08fF
C1377 PAND2X1_691/Y PAND2X1_729/a_16_344# 0.01fF
C1378 POR2X1_569/CTRL2 POR2X1_570/Y 0.02fF
C1379 POR2X1_68/A PAND2X1_273/CTRL2 0.03fF
C1380 PAND2X1_597/O POR2X1_796/A 0.01fF
C1381 POR2X1_137/CTRL2 PAND2X1_96/B 0.01fF
C1382 POR2X1_66/A POR2X1_552/A 0.01fF
C1383 PAND2X1_241/CTRL POR2X1_90/Y 0.01fF
C1384 VDD PAND2X1_149/A 0.24fF
C1385 POR2X1_558/A INPUT_0 0.04fF
C1386 POR2X1_590/A POR2X1_294/A 0.10fF
C1387 POR2X1_52/A PAND2X1_814/O 0.04fF
C1388 POR2X1_302/O POR2X1_383/A 0.05fF
C1389 POR2X1_853/A POR2X1_170/O 0.01fF
C1390 POR2X1_475/A POR2X1_362/A 0.01fF
C1391 POR2X1_423/Y PAND2X1_308/Y 0.00fF
C1392 POR2X1_41/B PAND2X1_319/B 0.03fF
C1393 POR2X1_38/Y PAND2X1_364/B 0.07fF
C1394 D_INPUT_1 POR2X1_294/B 0.10fF
C1395 POR2X1_341/A POR2X1_715/CTRL2 0.04fF
C1396 POR2X1_516/CTRL2 POR2X1_184/Y 0.09fF
C1397 POR2X1_96/B VDD 0.40fF
C1398 POR2X1_858/B POR2X1_362/B 0.01fF
C1399 PAND2X1_631/CTRL2 PAND2X1_6/A 0.07fF
C1400 POR2X1_244/B POR2X1_222/A 0.02fF
C1401 PAND2X1_631/A POR2X1_669/B 0.26fF
C1402 POR2X1_674/Y POR2X1_385/Y 0.05fF
C1403 POR2X1_198/CTRL2 PAND2X1_88/Y 0.01fF
C1404 PAND2X1_824/B POR2X1_61/Y 0.03fF
C1405 PAND2X1_207/O PAND2X1_207/A 0.02fF
C1406 PAND2X1_124/Y PAND2X1_198/O 0.01fF
C1407 PAND2X1_71/CTRL PAND2X1_111/B 0.01fF
C1408 POR2X1_35/Y POR2X1_219/CTRL2 0.01fF
C1409 POR2X1_252/CTRL2 POR2X1_7/A -0.03fF
C1410 INPUT_1 POR2X1_29/CTRL 0.01fF
C1411 POR2X1_805/Y PAND2X1_759/CTRL2 0.01fF
C1412 POR2X1_72/B PAND2X1_156/A 0.05fF
C1413 POR2X1_614/A POR2X1_804/B 0.01fF
C1414 PAND2X1_182/CTRL PAND2X1_357/Y 0.03fF
C1415 PAND2X1_69/A POR2X1_35/Y 0.03fF
C1416 PAND2X1_118/CTRL POR2X1_532/A 0.01fF
C1417 POR2X1_130/A POR2X1_664/CTRL2 0.08fF
C1418 POR2X1_757/A PAND2X1_645/B 0.01fF
C1419 POR2X1_493/B INPUT_0 0.04fF
C1420 PAND2X1_64/CTRL2 PAND2X1_52/B 0.33fF
C1421 POR2X1_489/CTRL2 POR2X1_113/B 0.01fF
C1422 POR2X1_72/B POR2X1_373/CTRL 0.01fF
C1423 POR2X1_790/A POR2X1_68/B 0.02fF
C1424 POR2X1_389/O POR2X1_537/B 0.12fF
C1425 POR2X1_752/CTRL2 INPUT_5 0.00fF
C1426 POR2X1_22/A INPUT_6 0.05fF
C1427 POR2X1_208/A POR2X1_198/B 0.01fF
C1428 POR2X1_590/A PAND2X1_102/CTRL 0.00fF
C1429 POR2X1_535/a_16_28# POR2X1_535/A 0.05fF
C1430 POR2X1_68/A POR2X1_544/a_56_344# 0.00fF
C1431 POR2X1_383/A PAND2X1_530/O 0.08fF
C1432 POR2X1_16/A PAND2X1_468/CTRL -0.02fF
C1433 POR2X1_8/Y POR2X1_13/A 0.03fF
C1434 POR2X1_366/CTRL PAND2X1_48/B 0.01fF
C1435 PAND2X1_6/Y POR2X1_318/A 0.12fF
C1436 PAND2X1_23/Y POR2X1_568/Y 0.05fF
C1437 POR2X1_853/A POR2X1_854/B 0.05fF
C1438 POR2X1_96/A PAND2X1_507/CTRL2 0.10fF
C1439 POR2X1_65/A PAND2X1_714/B 0.05fF
C1440 POR2X1_455/A POR2X1_510/Y 0.03fF
C1441 PAND2X1_90/Y PAND2X1_48/A 0.21fF
C1442 PAND2X1_48/B POR2X1_215/A 0.30fF
C1443 POR2X1_220/Y POR2X1_210/B 0.44fF
C1444 POR2X1_57/A PAND2X1_852/B 0.01fF
C1445 POR2X1_55/Y PAND2X1_514/CTRL 0.01fF
C1446 POR2X1_765/O POR2X1_765/Y 0.01fF
C1447 POR2X1_567/A PAND2X1_52/Y 0.05fF
C1448 POR2X1_43/Y POR2X1_48/A 0.03fF
C1449 POR2X1_327/Y POR2X1_302/Y 0.01fF
C1450 POR2X1_226/Y POR2X1_4/Y 0.03fF
C1451 POR2X1_865/B POR2X1_68/B 0.03fF
C1452 POR2X1_68/B PAND2X1_88/Y 0.01fF
C1453 POR2X1_513/Y POR2X1_228/Y 0.03fF
C1454 POR2X1_16/A POR2X1_689/A 0.00fF
C1455 D_INPUT_1 PAND2X1_111/B 0.04fF
C1456 POR2X1_209/A POR2X1_535/A 0.01fF
C1457 POR2X1_590/Y POR2X1_513/B 0.95fF
C1458 POR2X1_76/Y POR2X1_715/A 0.03fF
C1459 PAND2X1_55/Y POR2X1_407/a_76_344# 0.01fF
C1460 PAND2X1_798/B PAND2X1_574/O 0.03fF
C1461 PAND2X1_270/m4_208_n4# POR2X1_184/Y 0.12fF
C1462 PAND2X1_585/O PAND2X1_56/A 0.02fF
C1463 POR2X1_218/A POR2X1_362/A 0.02fF
C1464 POR2X1_527/Y POR2X1_90/Y 0.03fF
C1465 POR2X1_16/A PAND2X1_398/O 0.01fF
C1466 POR2X1_554/Y POR2X1_186/B 0.03fF
C1467 VDD POR2X1_726/O 0.00fF
C1468 PAND2X1_254/Y PAND2X1_508/Y 0.02fF
C1469 PAND2X1_389/Y PAND2X1_388/Y 0.46fF
C1470 POR2X1_664/CTRL POR2X1_712/Y 0.03fF
C1471 INPUT_6 POR2X1_1/CTRL2 0.04fF
C1472 PAND2X1_482/CTRL2 POR2X1_294/B 0.01fF
C1473 POR2X1_532/A PAND2X1_63/B 0.02fF
C1474 PAND2X1_65/B PAND2X1_179/O 0.03fF
C1475 POR2X1_16/A POR2X1_765/a_56_344# 0.00fF
C1476 POR2X1_423/Y POR2X1_77/Y 0.03fF
C1477 POR2X1_394/A PAND2X1_302/O 0.04fF
C1478 PAND2X1_824/B POR2X1_35/Y 0.51fF
C1479 POR2X1_327/Y POR2X1_861/CTRL 0.01fF
C1480 POR2X1_541/a_16_28# POR2X1_274/B 0.02fF
C1481 PAND2X1_849/B POR2X1_38/Y 0.02fF
C1482 POR2X1_840/B POR2X1_260/A 0.06fF
C1483 POR2X1_460/A POR2X1_752/O 0.06fF
C1484 POR2X1_750/B POR2X1_161/O 0.03fF
C1485 PAND2X1_6/Y POR2X1_574/Y 0.06fF
C1486 POR2X1_389/Y PAND2X1_52/B 0.03fF
C1487 PAND2X1_701/CTRL PAND2X1_69/A 0.01fF
C1488 POR2X1_13/A PAND2X1_346/CTRL 0.01fF
C1489 PAND2X1_234/CTRL2 POR2X1_66/A 0.01fF
C1490 POR2X1_489/CTRL2 POR2X1_768/A 0.06fF
C1491 PAND2X1_251/CTRL2 POR2X1_814/A 0.00fF
C1492 POR2X1_614/A POR2X1_334/Y 0.02fF
C1493 POR2X1_565/B POR2X1_4/Y 1.11fF
C1494 PAND2X1_630/B POR2X1_496/Y 0.06fF
C1495 POR2X1_327/Y POR2X1_501/B 0.03fF
C1496 POR2X1_537/Y POR2X1_114/B 0.05fF
C1497 POR2X1_567/A D_GATE_662 0.17fF
C1498 PAND2X1_467/Y PAND2X1_452/A 0.06fF
C1499 POR2X1_567/B POR2X1_440/B 0.05fF
C1500 POR2X1_468/B POR2X1_568/B 0.05fF
C1501 POR2X1_809/A POR2X1_605/A 0.43fF
C1502 POR2X1_16/A POR2X1_258/Y 0.03fF
C1503 PAND2X1_242/Y PAND2X1_390/Y 0.05fF
C1504 POR2X1_545/A POR2X1_551/A 0.35fF
C1505 POR2X1_7/A PAND2X1_507/CTRL2 0.03fF
C1506 INPUT_4 POR2X1_39/B 0.16fF
C1507 PAND2X1_858/CTRL PAND2X1_858/Y 0.00fF
C1508 POR2X1_865/CTRL PAND2X1_48/A 0.07fF
C1509 POR2X1_78/B POR2X1_147/O 0.03fF
C1510 POR2X1_334/Y POR2X1_360/CTRL2 0.01fF
C1511 POR2X1_43/B PAND2X1_338/O 0.01fF
C1512 PAND2X1_651/CTRL POR2X1_588/Y 0.01fF
C1513 PAND2X1_865/Y POR2X1_184/Y 0.02fF
C1514 PAND2X1_30/CTRL POR2X1_750/B 0.01fF
C1515 POR2X1_763/Y POR2X1_39/B 0.12fF
C1516 PAND2X1_798/Y POR2X1_42/Y 1.24fF
C1517 PAND2X1_23/Y POR2X1_486/B 0.10fF
C1518 PAND2X1_115/B POR2X1_39/B 0.52fF
C1519 POR2X1_270/Y POR2X1_659/a_16_28# 0.02fF
C1520 POR2X1_850/CTRL POR2X1_737/A 0.01fF
C1521 POR2X1_463/CTRL2 PAND2X1_58/A -0.00fF
C1522 PAND2X1_187/O POR2X1_191/B 0.00fF
C1523 POR2X1_213/B PAND2X1_146/CTRL 0.01fF
C1524 POR2X1_361/O PAND2X1_48/A 0.17fF
C1525 POR2X1_361/CTRL POR2X1_294/A 0.00fF
C1526 PAND2X1_94/A POR2X1_768/O 0.03fF
C1527 INPUT_1 PAND2X1_483/O 0.08fF
C1528 PAND2X1_658/A POR2X1_39/B 0.03fF
C1529 POR2X1_567/A POR2X1_724/A 0.15fF
C1530 PAND2X1_20/A PAND2X1_85/O 0.06fF
C1531 POR2X1_112/CTRL2 PAND2X1_60/B 0.01fF
C1532 POR2X1_327/Y POR2X1_539/CTRL 0.02fF
C1533 POR2X1_96/CTRL POR2X1_153/Y 0.01fF
C1534 PAND2X1_94/A PAND2X1_531/CTRL 0.01fF
C1535 GATE_222 PAND2X1_805/A 0.03fF
C1536 POR2X1_669/B POR2X1_669/Y 0.09fF
C1537 POR2X1_846/A POR2X1_752/Y 0.03fF
C1538 PAND2X1_440/CTRL PAND2X1_794/B 0.01fF
C1539 PAND2X1_132/a_16_344# PAND2X1_52/B 0.02fF
C1540 PAND2X1_39/B POR2X1_807/CTRL 0.01fF
C1541 POR2X1_99/A PAND2X1_86/CTRL2 0.00fF
C1542 POR2X1_150/Y PAND2X1_794/CTRL2 0.01fF
C1543 POR2X1_178/CTRL POR2X1_416/B 0.01fF
C1544 POR2X1_732/B PAND2X1_72/A 5.31fF
C1545 POR2X1_557/B POR2X1_768/CTRL 0.01fF
C1546 POR2X1_73/Y POR2X1_39/B 0.17fF
C1547 PAND2X1_649/A PAND2X1_656/A 0.03fF
C1548 POR2X1_97/CTRL POR2X1_97/B 0.01fF
C1549 POR2X1_77/Y PAND2X1_359/a_16_344# 0.01fF
C1550 POR2X1_7/O POR2X1_7/Y 0.02fF
C1551 POR2X1_814/B PAND2X1_85/O 0.01fF
C1552 POR2X1_54/Y POR2X1_754/Y 0.01fF
C1553 POR2X1_532/A POR2X1_342/A 0.01fF
C1554 PAND2X1_496/m4_208_n4# POR2X1_777/B 0.03fF
C1555 PAND2X1_43/a_16_344# POR2X1_296/B 0.02fF
C1556 POR2X1_632/Y POR2X1_318/A 0.17fF
C1557 PAND2X1_192/Y POR2X1_250/Y 0.09fF
C1558 POR2X1_862/A POR2X1_286/O 0.00fF
C1559 PAND2X1_563/A PAND2X1_554/CTRL2 0.01fF
C1560 PAND2X1_319/B POR2X1_77/Y 0.14fF
C1561 POR2X1_677/Y POR2X1_46/Y 0.05fF
C1562 POR2X1_274/A POR2X1_218/Y 0.07fF
C1563 PAND2X1_485/a_76_28# POR2X1_260/B 0.02fF
C1564 PAND2X1_449/O POR2X1_423/Y 0.02fF
C1565 PAND2X1_48/B POR2X1_651/Y 0.01fF
C1566 INPUT_2 POR2X1_8/CTRL2 0.01fF
C1567 POR2X1_68/A POR2X1_863/A 0.03fF
C1568 POR2X1_275/A PAND2X1_390/Y 0.00fF
C1569 POR2X1_500/CTRL POR2X1_318/A 0.02fF
C1570 POR2X1_862/Y POR2X1_590/A 0.06fF
C1571 POR2X1_60/A PAND2X1_407/O 0.02fF
C1572 POR2X1_188/Y POR2X1_741/A 0.01fF
C1573 POR2X1_411/B POR2X1_503/A 0.17fF
C1574 PAND2X1_166/m4_208_n4# POR2X1_854/B 0.04fF
C1575 POR2X1_260/B POR2X1_121/B 0.41fF
C1576 PAND2X1_11/O INPUT_5 0.07fF
C1577 PAND2X1_623/Y POR2X1_9/Y 0.07fF
C1578 POR2X1_65/A POR2X1_411/B 0.06fF
C1579 PAND2X1_52/B POR2X1_713/B 0.05fF
C1580 PAND2X1_237/CTRL POR2X1_241/B 0.01fF
C1581 PAND2X1_850/Y POR2X1_394/A 0.10fF
C1582 POR2X1_835/B VDD 0.20fF
C1583 PAND2X1_67/O POR2X1_330/Y 0.08fF
C1584 PAND2X1_793/Y POR2X1_67/Y 0.01fF
C1585 POR2X1_274/CTRL POR2X1_296/B 0.01fF
C1586 POR2X1_102/Y PAND2X1_571/A 0.03fF
C1587 PAND2X1_282/CTRL2 PAND2X1_73/Y 0.03fF
C1588 POR2X1_461/Y PAND2X1_90/Y 0.03fF
C1589 POR2X1_260/B POR2X1_267/a_16_28# 0.03fF
C1590 PAND2X1_93/B POR2X1_201/CTRL 0.01fF
C1591 PAND2X1_23/Y POR2X1_486/CTRL2 0.05fF
C1592 PAND2X1_48/B POR2X1_486/CTRL 0.01fF
C1593 POR2X1_416/B POR2X1_260/A 0.03fF
C1594 POR2X1_87/CTRL POR2X1_260/A 0.01fF
C1595 POR2X1_97/A POR2X1_78/A 0.13fF
C1596 POR2X1_326/A POR2X1_568/B 0.05fF
C1597 POR2X1_407/A POR2X1_458/Y 0.03fF
C1598 PAND2X1_341/B POR2X1_86/CTRL2 0.01fF
C1599 POR2X1_102/Y POR2X1_268/a_56_344# 0.00fF
C1600 PAND2X1_798/B PAND2X1_717/A 0.03fF
C1601 PAND2X1_217/a_16_344# INPUT_0 0.01fF
C1602 POR2X1_180/B POR2X1_863/A 0.03fF
C1603 POR2X1_257/A PAND2X1_480/B 0.10fF
C1604 POR2X1_66/A POR2X1_391/A 0.01fF
C1605 POR2X1_48/A PAND2X1_456/O 0.01fF
C1606 POR2X1_856/B POR2X1_856/O 0.08fF
C1607 POR2X1_55/CTRL2 POR2X1_94/A 0.01fF
C1608 PAND2X1_410/CTRL PAND2X1_404/A 0.00fF
C1609 POR2X1_84/A PAND2X1_85/Y 1.84fF
C1610 PAND2X1_9/Y POR2X1_247/CTRL2 0.02fF
C1611 POR2X1_48/A INPUT_7 0.02fF
C1612 POR2X1_188/A PAND2X1_282/a_16_344# 0.01fF
C1613 POR2X1_52/A PAND2X1_464/a_16_344# 0.03fF
C1614 POR2X1_163/Y PAND2X1_725/Y 0.05fF
C1615 POR2X1_102/Y POR2X1_251/CTRL 0.00fF
C1616 POR2X1_62/Y POR2X1_86/Y 0.00fF
C1617 POR2X1_23/Y PAND2X1_712/CTRL 0.01fF
C1618 POR2X1_94/A POR2X1_590/A 2.09fF
C1619 POR2X1_571/Y POR2X1_500/CTRL2 0.01fF
C1620 POR2X1_640/a_56_344# PAND2X1_73/Y 0.00fF
C1621 POR2X1_202/B POR2X1_202/O 0.00fF
C1622 PAND2X1_63/Y PAND2X1_246/CTRL2 0.00fF
C1623 PAND2X1_600/CTRL2 POR2X1_130/A 0.12fF
C1624 POR2X1_29/CTRL2 POR2X1_409/B 0.04fF
C1625 POR2X1_849/A POR2X1_849/a_16_28# 0.05fF
C1626 POR2X1_479/CTRL POR2X1_286/Y 0.16fF
C1627 POR2X1_60/A PAND2X1_390/Y 0.03fF
C1628 POR2X1_669/B POR2X1_763/A 0.07fF
C1629 PAND2X1_206/B PAND2X1_350/CTRL2 0.00fF
C1630 PAND2X1_58/A PAND2X1_23/O 0.01fF
C1631 POR2X1_78/B POR2X1_66/A 6.16fF
C1632 POR2X1_828/Y PAND2X1_73/Y 0.01fF
C1633 PAND2X1_20/A POR2X1_186/Y 22.06fF
C1634 POR2X1_54/Y POR2X1_42/Y 0.13fF
C1635 PAND2X1_485/CTRL POR2X1_546/A 0.02fF
C1636 PAND2X1_695/a_76_28# PAND2X1_59/B 0.02fF
C1637 POR2X1_504/Y POR2X1_14/Y 0.03fF
C1638 PAND2X1_216/CTRL2 PAND2X1_267/Y 0.01fF
C1639 POR2X1_650/A POR2X1_78/A 3.04fF
C1640 POR2X1_446/B PAND2X1_55/Y 0.03fF
C1641 POR2X1_257/A PAND2X1_162/CTRL 0.01fF
C1642 PAND2X1_836/CTRL2 POR2X1_411/B 0.01fF
C1643 POR2X1_12/A POR2X1_700/O 0.00fF
C1644 POR2X1_52/A POR2X1_815/Y 0.01fF
C1645 POR2X1_567/B PAND2X1_524/CTRL 0.00fF
C1646 POR2X1_121/A PAND2X1_39/B 0.01fF
C1647 POR2X1_274/O VDD 0.00fF
C1648 POR2X1_105/O POR2X1_814/B 0.07fF
C1649 PAND2X1_207/A POR2X1_39/B 0.03fF
C1650 POR2X1_102/Y PAND2X1_787/Y 0.05fF
C1651 D_INPUT_0 PAND2X1_734/B 0.03fF
C1652 PAND2X1_9/Y POR2X1_409/CTRL 0.01fF
C1653 POR2X1_415/A PAND2X1_6/A 0.08fF
C1654 PAND2X1_23/Y POR2X1_301/A 0.01fF
C1655 PAND2X1_437/CTRL POR2X1_186/B 0.01fF
C1656 POR2X1_722/B PAND2X1_93/B 0.01fF
C1657 POR2X1_296/B VDD 6.71fF
C1658 POR2X1_777/B POR2X1_734/A 0.10fF
C1659 POR2X1_567/B POR2X1_802/B 0.03fF
C1660 POR2X1_541/B POR2X1_541/O 0.01fF
C1661 POR2X1_43/B PAND2X1_444/CTRL2 0.03fF
C1662 POR2X1_48/A POR2X1_763/Y 0.10fF
C1663 PAND2X1_93/B POR2X1_294/B 0.63fF
C1664 POR2X1_186/Y POR2X1_776/CTRL2 0.01fF
C1665 POR2X1_366/Y PAND2X1_93/B 0.01fF
C1666 POR2X1_542/B POR2X1_663/B 0.05fF
C1667 PAND2X1_56/Y POR2X1_260/B 0.03fF
C1668 POR2X1_260/B POR2X1_795/B 0.11fF
C1669 POR2X1_356/A POR2X1_466/A 0.02fF
C1670 POR2X1_814/B POR2X1_186/Y 0.03fF
C1671 POR2X1_466/A PAND2X1_183/a_16_344# 0.06fF
C1672 PAND2X1_218/O PAND2X1_267/Y 0.02fF
C1673 PAND2X1_58/A PAND2X1_511/CTRL2 0.01fF
C1674 POR2X1_68/A POR2X1_274/A 0.03fF
C1675 PAND2X1_471/B POR2X1_669/B 1.07fF
C1676 POR2X1_45/Y PAND2X1_124/Y 0.03fF
C1677 POR2X1_130/A POR2X1_267/O 0.03fF
C1678 POR2X1_590/A PAND2X1_754/CTRL2 0.01fF
C1679 PAND2X1_209/A PAND2X1_213/O 0.03fF
C1680 POR2X1_54/Y POR2X1_15/CTRL2 0.30fF
C1681 POR2X1_16/A POR2X1_600/O 0.02fF
C1682 PAND2X1_65/B POR2X1_734/A 1.66fF
C1683 POR2X1_188/CTRL2 PAND2X1_39/B 0.03fF
C1684 POR2X1_65/A POR2X1_376/B 0.06fF
C1685 POR2X1_848/A POR2X1_790/A 0.20fF
C1686 POR2X1_590/A PAND2X1_110/CTRL2 0.01fF
C1687 POR2X1_407/A PAND2X1_251/O 0.01fF
C1688 PAND2X1_557/A PAND2X1_739/Y 0.08fF
C1689 POR2X1_32/A POR2X1_494/Y 0.07fF
C1690 POR2X1_49/Y PAND2X1_596/O 0.02fF
C1691 POR2X1_646/O POR2X1_121/B 0.01fF
C1692 POR2X1_568/A POR2X1_568/CTRL 0.01fF
C1693 POR2X1_847/a_16_28# POR2X1_283/A 0.03fF
C1694 POR2X1_3/A POR2X1_12/A 1.01fF
C1695 PAND2X1_90/A PAND2X1_245/CTRL 0.01fF
C1696 POR2X1_499/A POR2X1_101/Y 3.81fF
C1697 POR2X1_14/Y POR2X1_586/O 0.01fF
C1698 POR2X1_99/A INPUT_0 0.34fF
C1699 POR2X1_730/Y POR2X1_467/O 0.01fF
C1700 POR2X1_800/A POR2X1_801/B 0.03fF
C1701 POR2X1_863/A POR2X1_169/A 0.03fF
C1702 POR2X1_366/Y POR2X1_78/A 0.07fF
C1703 POR2X1_78/A POR2X1_294/B 13.82fF
C1704 POR2X1_17/CTRL VDD 0.00fF
C1705 PAND2X1_392/B POR2X1_236/Y 0.06fF
C1706 POR2X1_865/B POR2X1_458/CTRL2 0.03fF
C1707 POR2X1_679/A PAND2X1_175/B 0.19fF
C1708 PAND2X1_247/a_76_28# POR2X1_7/A 0.01fF
C1709 POR2X1_853/A PAND2X1_73/Y 0.01fF
C1710 POR2X1_499/O POR2X1_576/Y 0.01fF
C1711 PAND2X1_55/Y POR2X1_121/B 0.15fF
C1712 POR2X1_296/B POR2X1_741/Y 0.08fF
C1713 POR2X1_444/B POR2X1_319/Y 0.15fF
C1714 PAND2X1_401/CTRL2 POR2X1_14/Y 0.01fF
C1715 POR2X1_48/A POR2X1_73/Y 0.21fF
C1716 POR2X1_422/O POR2X1_93/A 0.08fF
C1717 POR2X1_49/Y PAND2X1_480/B 0.01fF
C1718 PAND2X1_81/B POR2X1_296/B 0.02fF
C1719 POR2X1_567/B POR2X1_532/A 0.05fF
C1720 PAND2X1_419/O PAND2X1_69/A -0.00fF
C1721 POR2X1_840/B POR2X1_656/CTRL2 0.18fF
C1722 POR2X1_45/Y POR2X1_83/B 0.03fF
C1723 POR2X1_333/A POR2X1_468/a_16_28# 0.04fF
C1724 POR2X1_121/A POR2X1_805/Y 0.05fF
C1725 PAND2X1_73/Y POR2X1_391/Y 0.07fF
C1726 POR2X1_49/Y POR2X1_754/A 0.03fF
C1727 PAND2X1_784/A POR2X1_42/Y 0.03fF
C1728 PAND2X1_219/A PAND2X1_219/a_16_344# 0.02fF
C1729 POR2X1_270/CTRL POR2X1_66/A 0.00fF
C1730 POR2X1_278/Y POR2X1_488/O 0.08fF
C1731 PAND2X1_93/B PAND2X1_111/B 0.03fF
C1732 POR2X1_52/A POR2X1_503/A 0.01fF
C1733 PAND2X1_554/a_76_28# POR2X1_7/B 0.01fF
C1734 POR2X1_471/A POR2X1_456/B 0.03fF
C1735 POR2X1_383/A POR2X1_260/B 0.37fF
C1736 POR2X1_45/CTRL2 PAND2X1_480/B 0.15fF
C1737 POR2X1_121/A PAND2X1_20/A 0.07fF
C1738 PAND2X1_222/A POR2X1_385/CTRL 0.00fF
C1739 PAND2X1_65/B PAND2X1_224/CTRL2 0.01fF
C1740 POR2X1_236/Y VDD 5.18fF
C1741 POR2X1_97/A POR2X1_775/a_76_344# 0.01fF
C1742 POR2X1_54/Y POR2X1_754/CTRL 0.05fF
C1743 POR2X1_278/Y PAND2X1_204/CTRL 0.06fF
C1744 POR2X1_464/CTRL VDD 0.00fF
C1745 PAND2X1_801/B PAND2X1_863/B 0.01fF
C1746 POR2X1_52/A POR2X1_65/A 0.22fF
C1747 POR2X1_547/B VDD 0.02fF
C1748 POR2X1_296/B PAND2X1_32/B 0.13fF
C1749 POR2X1_196/Y POR2X1_555/B 0.02fF
C1750 PAND2X1_47/CTRL PAND2X1_11/Y 0.02fF
C1751 POR2X1_504/Y POR2X1_55/Y 0.04fF
C1752 POR2X1_62/O POR2X1_750/B 0.01fF
C1753 POR2X1_52/A PAND2X1_558/CTRL 0.01fF
C1754 POR2X1_655/CTRL2 POR2X1_711/Y 0.05fF
C1755 POR2X1_407/Y POR2X1_121/B 0.03fF
C1756 POR2X1_57/A POR2X1_666/O 0.01fF
C1757 POR2X1_740/Y POR2X1_543/A 0.03fF
C1758 POR2X1_481/A POR2X1_295/Y 0.09fF
C1759 POR2X1_65/A POR2X1_152/A 0.03fF
C1760 POR2X1_98/B POR2X1_240/B 0.23fF
C1761 POR2X1_257/A PAND2X1_725/CTRL2 0.00fF
C1762 POR2X1_614/A POR2X1_254/CTRL2 0.03fF
C1763 POR2X1_65/A PAND2X1_105/CTRL2 0.10fF
C1764 PAND2X1_65/B POR2X1_828/O 0.01fF
C1765 PAND2X1_11/Y PAND2X1_26/O 0.04fF
C1766 POR2X1_188/A POR2X1_710/CTRL 0.01fF
C1767 PAND2X1_74/CTRL PAND2X1_32/B 0.01fF
C1768 INPUT_1 POR2X1_817/CTRL2 0.01fF
C1769 POR2X1_610/O POR2X1_260/A 0.09fF
C1770 PAND2X1_274/O PAND2X1_480/B 0.07fF
C1771 POR2X1_71/Y PAND2X1_501/B 0.03fF
C1772 POR2X1_121/A POR2X1_814/B 0.02fF
C1773 POR2X1_43/B POR2X1_39/O 0.02fF
C1774 PAND2X1_6/Y POR2X1_35/B 0.01fF
C1775 POR2X1_777/B POR2X1_786/Y 0.07fF
C1776 POR2X1_78/A PAND2X1_111/B 0.03fF
C1777 POR2X1_81/Y VDD 0.20fF
C1778 POR2X1_278/Y POR2X1_46/Y 0.10fF
C1779 PAND2X1_423/a_76_28# PAND2X1_55/Y 0.01fF
C1780 POR2X1_396/Y POR2X1_83/B 0.03fF
C1781 POR2X1_57/A PAND2X1_403/B 0.29fF
C1782 PAND2X1_662/CTRL2 PAND2X1_660/B 0.01fF
C1783 PAND2X1_436/CTRL POR2X1_129/Y 0.01fF
C1784 PAND2X1_820/CTRL2 POR2X1_669/B 0.05fF
C1785 POR2X1_166/CTRL POR2X1_40/Y 0.01fF
C1786 POR2X1_68/A POR2X1_797/CTRL 0.01fF
C1787 PAND2X1_480/B PAND2X1_553/B 0.05fF
C1788 POR2X1_62/Y POR2X1_624/Y 0.02fF
C1789 POR2X1_748/A POR2X1_93/A 0.03fF
C1790 POR2X1_793/O POR2X1_789/Y 0.00fF
C1791 POR2X1_672/A POR2X1_5/Y 0.01fF
C1792 POR2X1_78/B POR2X1_222/Y 0.07fF
C1793 POR2X1_376/B PAND2X1_565/O 0.16fF
C1794 POR2X1_416/B POR2X1_329/A 0.23fF
C1795 POR2X1_25/Y POR2X1_12/A 0.06fF
C1796 D_INPUT_3 POR2X1_40/Y 0.12fF
C1797 POR2X1_548/B POR2X1_502/A 0.01fF
C1798 PAND2X1_480/B PAND2X1_303/O 0.04fF
C1799 PAND2X1_65/B POR2X1_786/Y 0.07fF
C1800 PAND2X1_84/Y PAND2X1_717/O 0.02fF
C1801 PAND2X1_425/O INPUT_6 0.02fF
C1802 POR2X1_334/B PAND2X1_80/a_16_344# 0.03fF
C1803 VDD POR2X1_501/O 0.00fF
C1804 PAND2X1_803/A POR2X1_90/Y 0.04fF
C1805 POR2X1_332/B POR2X1_740/Y 0.05fF
C1806 PAND2X1_58/A POR2X1_796/A 0.03fF
C1807 POR2X1_684/CTRL POR2X1_7/B 0.01fF
C1808 PAND2X1_81/B POR2X1_547/B 0.06fF
C1809 POR2X1_258/a_16_28# POR2X1_312/Y 0.01fF
C1810 POR2X1_335/A POR2X1_302/Y 0.02fF
C1811 PAND2X1_241/Y POR2X1_423/Y 0.03fF
C1812 PAND2X1_580/CTRL VDD -0.00fF
C1813 PAND2X1_467/Y POR2X1_14/Y 4.02fF
C1814 POR2X1_78/B POR2X1_84/a_16_28# 0.00fF
C1815 PAND2X1_735/CTRL2 POR2X1_816/A 0.03fF
C1816 POR2X1_673/Y POR2X1_296/B 0.03fF
C1817 POR2X1_543/A PAND2X1_312/CTRL2 0.01fF
C1818 POR2X1_304/Y POR2X1_305/Y 0.00fF
C1819 POR2X1_346/B PAND2X1_39/O 0.00fF
C1820 POR2X1_267/Y VDD 0.11fF
C1821 POR2X1_327/CTRL POR2X1_572/B 0.01fF
C1822 POR2X1_311/Y PAND2X1_336/CTRL 0.02fF
C1823 PAND2X1_65/B POR2X1_788/B 1.37fF
C1824 POR2X1_8/Y POR2X1_29/A 0.03fF
C1825 POR2X1_437/O POR2X1_385/Y 0.02fF
C1826 PAND2X1_591/CTRL2 PAND2X1_48/A 0.04fF
C1827 POR2X1_355/B POR2X1_775/A 0.19fF
C1828 PAND2X1_722/CTRL POR2X1_394/A 0.01fF
C1829 POR2X1_232/Y VDD 0.12fF
C1830 POR2X1_178/CTRL PAND2X1_738/Y 0.13fF
C1831 PAND2X1_20/A POR2X1_664/CTRL 0.00fF
C1832 POR2X1_41/B PAND2X1_798/B 0.07fF
C1833 POR2X1_547/B PAND2X1_32/B 0.03fF
C1834 PAND2X1_839/O POR2X1_293/Y 0.15fF
C1835 POR2X1_790/B PAND2X1_753/CTRL 0.00fF
C1836 POR2X1_174/A POR2X1_704/Y 0.11fF
C1837 POR2X1_16/A PAND2X1_404/O 0.02fF
C1838 POR2X1_78/B POR2X1_532/A 0.21fF
C1839 POR2X1_339/O PAND2X1_20/A 0.01fF
C1840 D_GATE_222 POR2X1_776/B 0.06fF
C1841 VDD PAND2X1_858/Y 0.06fF
C1842 POR2X1_52/A PAND2X1_190/Y 0.01fF
C1843 POR2X1_505/Y PAND2X1_632/B 0.04fF
C1844 POR2X1_5/Y POR2X1_387/Y 0.11fF
C1845 POR2X1_13/Y POR2X1_42/Y 0.03fF
C1846 POR2X1_66/A POR2X1_294/A 1.24fF
C1847 POR2X1_514/a_16_28# INPUT_0 0.01fF
C1848 POR2X1_567/A PAND2X1_93/B 8.48fF
C1849 POR2X1_22/A POR2X1_22/a_16_28# 0.05fF
C1850 POR2X1_391/Y PAND2X1_132/CTRL2 0.02fF
C1851 PAND2X1_94/A PAND2X1_42/CTRL2 0.01fF
C1852 POR2X1_445/a_16_28# POR2X1_455/A 0.03fF
C1853 PAND2X1_56/Y PAND2X1_55/Y 0.07fF
C1854 PAND2X1_55/Y POR2X1_795/B 0.07fF
C1855 POR2X1_16/A POR2X1_492/CTRL2 0.19fF
C1856 PAND2X1_714/Y PAND2X1_731/B 0.04fF
C1857 PAND2X1_48/B POR2X1_114/B 0.03fF
C1858 POR2X1_243/Y PAND2X1_88/Y 0.06fF
C1859 POR2X1_34/A POR2X1_294/A 0.01fF
C1860 POR2X1_844/CTRL POR2X1_546/A 0.00fF
C1861 POR2X1_188/A POR2X1_675/Y 0.02fF
C1862 POR2X1_566/A POR2X1_341/Y 0.05fF
C1863 POR2X1_510/A POR2X1_294/B 0.02fF
C1864 POR2X1_856/CTRL2 POR2X1_260/A 0.02fF
C1865 POR2X1_582/CTRL2 INPUT_5 0.01fF
C1866 POR2X1_750/B POR2X1_156/Y 0.71fF
C1867 PAND2X1_38/O POR2X1_68/B 0.04fF
C1868 PAND2X1_7/O POR2X1_222/Y 0.01fF
C1869 PAND2X1_6/Y PAND2X1_275/CTRL2 0.09fF
C1870 POR2X1_572/B POR2X1_218/A 0.01fF
C1871 PAND2X1_631/O POR2X1_293/Y 0.07fF
C1872 PAND2X1_476/A POR2X1_37/Y 0.14fF
C1873 POR2X1_52/CTRL PAND2X1_124/Y 0.07fF
C1874 PAND2X1_651/Y POR2X1_494/Y 0.05fF
C1875 POR2X1_188/A POR2X1_851/CTRL2 0.01fF
C1876 POR2X1_800/A POR2X1_796/CTRL2 0.00fF
C1877 POR2X1_565/B D_INPUT_1 0.07fF
C1878 POR2X1_16/A PAND2X1_61/Y 0.00fF
C1879 POR2X1_394/A PAND2X1_545/O 0.10fF
C1880 PAND2X1_341/B POR2X1_32/A 0.01fF
C1881 POR2X1_567/B POR2X1_510/CTRL2 0.15fF
C1882 POR2X1_503/O POR2X1_65/A 0.18fF
C1883 POR2X1_591/Y PAND2X1_364/B 0.02fF
C1884 PAND2X1_556/B POR2X1_283/A 0.02fF
C1885 POR2X1_483/B POR2X1_222/A 0.01fF
C1886 POR2X1_852/B POR2X1_507/A 0.07fF
C1887 POR2X1_73/Y PAND2X1_197/Y 0.03fF
C1888 PAND2X1_48/B POR2X1_458/B 0.02fF
C1889 POR2X1_507/CTRL VDD 0.00fF
C1890 PAND2X1_859/A POR2X1_394/A 0.09fF
C1891 POR2X1_567/A POR2X1_78/A 0.07fF
C1892 PAND2X1_39/B POR2X1_717/B 0.02fF
C1893 POR2X1_558/O PAND2X1_32/B 0.01fF
C1894 PAND2X1_401/CTRL POR2X1_73/Y 0.00fF
C1895 PAND2X1_552/B PAND2X1_388/CTRL 0.01fF
C1896 POR2X1_575/B POR2X1_573/A 0.20fF
C1897 POR2X1_501/O PAND2X1_32/B 0.09fF
C1898 INPUT_1 POR2X1_58/O 0.02fF
C1899 POR2X1_327/Y PAND2X1_299/O 0.02fF
C1900 PAND2X1_470/O POR2X1_238/Y 0.01fF
C1901 PAND2X1_94/A POR2X1_87/Y 0.01fF
C1902 POR2X1_335/A POR2X1_501/B 0.09fF
C1903 POR2X1_502/A POR2X1_566/B 0.13fF
C1904 POR2X1_56/Y POR2X1_816/A 0.03fF
C1905 POR2X1_49/Y POR2X1_373/Y 0.03fF
C1906 PAND2X1_254/Y POR2X1_283/A 0.03fF
C1907 PAND2X1_652/CTRL2 POR2X1_83/B 0.01fF
C1908 POR2X1_407/A D_INPUT_1 0.03fF
C1909 POR2X1_502/A POR2X1_180/A 0.03fF
C1910 PAND2X1_839/B POR2X1_293/Y 0.02fF
C1911 POR2X1_16/A PAND2X1_404/A 0.12fF
C1912 POR2X1_68/A PAND2X1_424/CTRL2 0.05fF
C1913 VDD POR2X1_757/Y 0.09fF
C1914 POR2X1_267/Y PAND2X1_32/B 0.07fF
C1915 POR2X1_327/Y POR2X1_733/CTRL2 0.02fF
C1916 D_INPUT_3 PAND2X1_8/a_16_344# 0.02fF
C1917 POR2X1_447/B POR2X1_330/Y 0.07fF
C1918 POR2X1_383/A POR2X1_340/CTRL 0.00fF
C1919 POR2X1_140/B POR2X1_724/A 0.03fF
C1920 POR2X1_83/Y POR2X1_40/Y 0.02fF
C1921 POR2X1_383/A POR2X1_205/Y 0.02fF
C1922 PAND2X1_48/B POR2X1_222/A 0.01fF
C1923 POR2X1_72/B POR2X1_171/Y 0.00fF
C1924 POR2X1_804/A POR2X1_541/CTRL2 0.08fF
C1925 POR2X1_740/Y POR2X1_574/A 0.03fF
C1926 POR2X1_383/A PAND2X1_55/Y 2.48fF
C1927 POR2X1_559/O POR2X1_38/B 0.30fF
C1928 POR2X1_590/Y VDD 0.01fF
C1929 POR2X1_753/Y POR2X1_39/B 0.43fF
C1930 POR2X1_538/A POR2X1_740/Y 0.03fF
C1931 POR2X1_417/Y PAND2X1_352/Y 0.65fF
C1932 PAND2X1_787/A POR2X1_309/Y 0.02fF
C1933 PAND2X1_821/CTRL POR2X1_854/B 0.15fF
C1934 PAND2X1_5/a_76_28# D_INPUT_2 0.02fF
C1935 POR2X1_271/A VDD 0.21fF
C1936 POR2X1_186/Y PAND2X1_680/O 0.18fF
C1937 POR2X1_383/A POR2X1_205/O 0.10fF
C1938 POR2X1_110/Y PAND2X1_803/A 0.03fF
C1939 PAND2X1_4/CTRL2 POR2X1_38/B 0.01fF
C1940 PAND2X1_445/m4_208_n4# PAND2X1_457/m4_208_n4# 0.13fF
C1941 PAND2X1_865/Y PAND2X1_579/CTRL 0.01fF
C1942 PAND2X1_703/CTRL POR2X1_236/Y 0.01fF
C1943 POR2X1_466/A PAND2X1_72/A 0.10fF
C1944 POR2X1_631/A PAND2X1_69/A 0.00fF
C1945 POR2X1_546/A POR2X1_546/a_16_28# 0.05fF
C1946 PAND2X1_390/Y POR2X1_589/CTRL2 0.01fF
C1947 PAND2X1_48/B PAND2X1_103/O 0.02fF
C1948 PAND2X1_731/O PAND2X1_731/A 0.02fF
C1949 PAND2X1_56/Y POR2X1_337/A 0.10fF
C1950 POR2X1_507/CTRL2 D_GATE_741 0.02fF
C1951 POR2X1_313/a_16_28# POR2X1_90/Y 0.10fF
C1952 POR2X1_96/A POR2X1_394/A 1.06fF
C1953 POR2X1_387/Y POR2X1_310/O 0.06fF
C1954 POR2X1_814/B POR2X1_542/Y 0.01fF
C1955 PAND2X1_804/B PAND2X1_853/B 0.19fF
C1956 POR2X1_252/CTRL2 POR2X1_153/Y 0.14fF
C1957 PAND2X1_785/A POR2X1_91/Y 0.03fF
C1958 PAND2X1_764/CTRL PAND2X1_32/B 0.01fF
C1959 POR2X1_334/B PAND2X1_184/CTRL 0.01fF
C1960 PAND2X1_23/Y PAND2X1_481/CTRL2 0.01fF
C1961 POR2X1_62/Y PAND2X1_459/Y 0.02fF
C1962 POR2X1_383/A POR2X1_407/Y 0.03fF
C1963 POR2X1_73/Y PAND2X1_840/O 0.01fF
C1964 POR2X1_265/Y POR2X1_13/A 0.26fF
C1965 PAND2X1_266/CTRL POR2X1_262/Y 0.00fF
C1966 POR2X1_840/B POR2X1_725/Y 0.01fF
C1967 POR2X1_550/O POR2X1_550/Y 0.19fF
C1968 POR2X1_671/O POR2X1_4/Y 0.02fF
C1969 POR2X1_559/B POR2X1_68/B 0.00fF
C1970 POR2X1_569/O POR2X1_568/B 0.04fF
C1971 PAND2X1_846/O POR2X1_750/A 0.05fF
C1972 POR2X1_7/B PAND2X1_156/A 0.09fF
C1973 PAND2X1_476/A POR2X1_406/Y 0.18fF
C1974 POR2X1_662/Y POR2X1_186/B 0.02fF
C1975 PAND2X1_751/O POR2X1_294/A 0.04fF
C1976 PAND2X1_671/CTRL INPUT_2 0.00fF
C1977 POR2X1_532/A POR2X1_141/A 0.01fF
C1978 PAND2X1_563/A PAND2X1_566/Y 0.07fF
C1979 POR2X1_537/Y POR2X1_784/A 0.02fF
C1980 POR2X1_463/Y PAND2X1_69/A 0.06fF
C1981 PAND2X1_55/Y PAND2X1_71/Y 0.03fF
C1982 POR2X1_480/A POR2X1_568/B 0.10fF
C1983 PAND2X1_96/B PAND2X1_184/CTRL2 0.00fF
C1984 POR2X1_817/A POR2X1_4/Y 0.03fF
C1985 PAND2X1_96/B POR2X1_332/CTRL2 0.09fF
C1986 POR2X1_565/B POR2X1_620/B 0.00fF
C1987 POR2X1_857/m4_208_n4# PAND2X1_72/A 0.09fF
C1988 POR2X1_845/O POR2X1_7/A 0.01fF
C1989 POR2X1_616/Y POR2X1_617/CTRL 0.01fF
C1990 POR2X1_614/A POR2X1_724/B 0.00fF
C1991 PAND2X1_569/B PAND2X1_168/O 0.00fF
C1992 POR2X1_222/Y POR2X1_735/CTRL 0.10fF
C1993 POR2X1_686/CTRL POR2X1_260/A 0.01fF
C1994 POR2X1_316/Y PAND2X1_455/Y 0.10fF
C1995 PAND2X1_476/A POR2X1_293/Y 0.03fF
C1996 POR2X1_283/A PAND2X1_175/CTRL2 0.01fF
C1997 POR2X1_274/B POR2X1_569/A 0.04fF
C1998 POR2X1_798/O PAND2X1_52/B 0.01fF
C1999 POR2X1_346/A POR2X1_837/B 0.01fF
C2000 PAND2X1_182/B PAND2X1_182/a_16_344# 0.01fF
C2001 POR2X1_42/Y POR2X1_4/Y 0.20fF
C2002 PAND2X1_48/B PAND2X1_122/CTRL2 0.00fF
C2003 POR2X1_814/B POR2X1_717/B 0.06fF
C2004 D_GATE_222 POR2X1_192/B 0.10fF
C2005 PAND2X1_48/B PAND2X1_665/CTRL2 0.03fF
C2006 PAND2X1_824/B POR2X1_631/A 0.07fF
C2007 POR2X1_41/a_16_28# POR2X1_73/Y 0.07fF
C2008 POR2X1_10/CTRL2 POR2X1_7/A 0.03fF
C2009 INPUT_0 PAND2X1_136/a_76_28# 0.02fF
C2010 POR2X1_740/Y POR2X1_738/CTRL2 0.00fF
C2011 PAND2X1_785/Y POR2X1_39/B 0.03fF
C2012 POR2X1_43/B POR2X1_183/a_16_28# 0.02fF
C2013 PAND2X1_23/Y POR2X1_374/O 0.01fF
C2014 POR2X1_62/Y POR2X1_73/Y 0.06fF
C2015 PAND2X1_61/a_76_28# POR2X1_9/Y 0.02fF
C2016 PAND2X1_341/B PAND2X1_651/Y 0.05fF
C2017 POR2X1_9/Y PAND2X1_58/A 0.10fF
C2018 POR2X1_532/A POR2X1_735/CTRL 0.01fF
C2019 PAND2X1_862/B POR2X1_80/CTRL2 0.01fF
C2020 POR2X1_325/A POR2X1_717/B 0.04fF
C2021 PAND2X1_119/O POR2X1_294/A 0.22fF
C2022 POR2X1_738/A POR2X1_353/A 0.01fF
C2023 POR2X1_63/Y POR2X1_813/a_76_344# 0.01fF
C2024 PAND2X1_785/A POR2X1_109/Y 0.01fF
C2025 POR2X1_49/Y POR2X1_386/Y 0.07fF
C2026 POR2X1_394/A POR2X1_7/A 0.09fF
C2027 POR2X1_532/A POR2X1_294/A 0.83fF
C2028 POR2X1_112/a_16_28# POR2X1_775/A 0.05fF
C2029 PAND2X1_653/Y PAND2X1_737/CTRL 0.10fF
C2030 POR2X1_502/A POR2X1_325/B 0.01fF
C2031 PAND2X1_108/CTRL2 PAND2X1_55/Y 0.06fF
C2032 PAND2X1_465/B POR2X1_77/Y 0.03fF
C2033 POR2X1_338/O POR2X1_334/Y 0.06fF
C2034 PAND2X1_831/Y PAND2X1_716/B 0.01fF
C2035 PAND2X1_404/Y POR2X1_490/a_56_344# 0.00fF
C2036 POR2X1_313/Y PAND2X1_317/CTRL 0.01fF
C2037 POR2X1_776/B POR2X1_567/m4_208_n4# 0.10fF
C2038 POR2X1_493/A POR2X1_556/A 0.06fF
C2039 PAND2X1_96/B POR2X1_554/CTRL2 0.01fF
C2040 POR2X1_13/A POR2X1_167/Y 0.02fF
C2041 POR2X1_263/CTRL POR2X1_37/Y 0.01fF
C2042 PAND2X1_514/O PAND2X1_348/A 0.05fF
C2043 POR2X1_610/Y POR2X1_610/O 0.01fF
C2044 POR2X1_327/Y POR2X1_860/CTRL 0.01fF
C2045 PAND2X1_450/CTRL2 POR2X1_416/B 0.00fF
C2046 PAND2X1_798/B POR2X1_77/Y 0.02fF
C2047 PAND2X1_358/A PAND2X1_100/O 0.05fF
C2048 POR2X1_736/A PAND2X1_178/m4_208_n4# 0.07fF
C2049 PAND2X1_481/O POR2X1_260/A 0.01fF
C2050 POR2X1_863/A POR2X1_435/Y 0.20fF
C2051 POR2X1_62/Y PAND2X1_244/B 0.03fF
C2052 POR2X1_66/B POR2X1_814/Y 0.02fF
C2053 POR2X1_286/B POR2X1_66/A 0.01fF
C2054 POR2X1_276/B POR2X1_218/Y 0.03fF
C2055 POR2X1_394/A POR2X1_394/a_76_344# 0.01fF
C2056 PAND2X1_69/A POR2X1_736/A 0.05fF
C2057 POR2X1_814/A POR2X1_734/A 0.07fF
C2058 POR2X1_83/B POR2X1_271/B 0.03fF
C2059 POR2X1_149/B PAND2X1_72/A 0.05fF
C2060 PAND2X1_9/Y POR2X1_296/B 2.58fF
C2061 POR2X1_191/O POR2X1_319/Y 0.02fF
C2062 PAND2X1_287/Y PAND2X1_773/Y 0.03fF
C2063 POR2X1_496/Y PAND2X1_796/B 0.00fF
C2064 POR2X1_78/B PAND2X1_607/CTRL 0.01fF
C2065 POR2X1_68/A PAND2X1_96/O 0.17fF
C2066 PAND2X1_323/CTRL POR2X1_456/B 0.01fF
C2067 POR2X1_57/A POR2X1_416/B 0.41fF
C2068 POR2X1_846/Y POR2X1_734/A 0.05fF
C2069 PAND2X1_631/A PAND2X1_514/O 0.05fF
C2070 PAND2X1_535/CTRL POR2X1_533/Y 0.01fF
C2071 PAND2X1_438/O POR2X1_192/Y 0.02fF
C2072 PAND2X1_656/A POR2X1_39/B 0.03fF
C2073 PAND2X1_33/CTRL POR2X1_94/A 0.01fF
C2074 POR2X1_150/Y POR2X1_72/B 0.07fF
C2075 POR2X1_298/CTRL POR2X1_32/A 0.01fF
C2076 POR2X1_624/B POR2X1_5/Y 0.19fF
C2077 POR2X1_112/Y PAND2X1_135/CTRL 0.09fF
C2078 POR2X1_715/a_56_344# POR2X1_702/A 0.00fF
C2079 POR2X1_325/O POR2X1_736/A 0.03fF
C2080 POR2X1_16/A POR2X1_85/O 0.01fF
C2081 POR2X1_39/B PAND2X1_124/CTRL2 0.00fF
C2082 POR2X1_23/Y POR2X1_496/Y 0.09fF
C2083 POR2X1_773/A POR2X1_113/B 0.03fF
C2084 POR2X1_66/B POR2X1_659/A 0.01fF
C2085 PAND2X1_96/B POR2X1_863/A 0.03fF
C2086 POR2X1_48/A POR2X1_753/Y 0.07fF
C2087 POR2X1_847/B POR2X1_20/B 0.10fF
C2088 POR2X1_54/Y POR2X1_615/CTRL2 0.01fF
C2089 PAND2X1_600/CTRL PAND2X1_20/A -0.00fF
C2090 POR2X1_22/A PAND2X1_635/Y 0.06fF
C2091 POR2X1_754/O POR2X1_39/B 0.02fF
C2092 PAND2X1_76/Y POR2X1_20/B 0.03fF
C2093 POR2X1_54/Y PAND2X1_463/a_16_344# 0.02fF
C2094 POR2X1_423/Y POR2X1_253/a_16_28# 0.02fF
C2095 POR2X1_634/O POR2X1_260/B 0.01fF
C2096 POR2X1_417/Y POR2X1_298/CTRL 0.01fF
C2097 POR2X1_866/A POR2X1_866/a_56_344# 0.03fF
C2098 POR2X1_122/Y POR2X1_411/B 0.01fF
C2099 PAND2X1_348/A POR2X1_39/B 0.07fF
C2100 POR2X1_558/B POR2X1_474/CTRL 0.01fF
C2101 POR2X1_852/CTRL POR2X1_776/A 0.03fF
C2102 PAND2X1_9/Y POR2X1_236/Y 0.05fF
C2103 POR2X1_111/Y POR2X1_416/B 0.02fF
C2104 PAND2X1_834/O POR2X1_153/Y 0.12fF
C2105 POR2X1_65/A POR2X1_681/Y 0.03fF
C2106 POR2X1_23/Y PAND2X1_733/A 0.03fF
C2107 POR2X1_638/A POR2X1_66/A 0.05fF
C2108 POR2X1_96/A POR2X1_679/O 0.02fF
C2109 POR2X1_48/A PAND2X1_541/CTRL2 0.01fF
C2110 POR2X1_3/B D_INPUT_4 0.01fF
C2111 PAND2X1_823/a_16_344# PAND2X1_52/B 0.01fF
C2112 POR2X1_300/Y POR2X1_39/B 0.06fF
C2113 POR2X1_257/A PAND2X1_276/a_76_28# 0.02fF
C2114 PAND2X1_147/O POR2X1_142/Y 0.03fF
C2115 PAND2X1_475/O D_INPUT_0 0.06fF
C2116 POR2X1_62/Y PAND2X1_358/CTRL 0.01fF
C2117 PAND2X1_72/Y PAND2X1_72/A 0.01fF
C2118 PAND2X1_669/CTRL POR2X1_750/B 0.01fF
C2119 PAND2X1_638/B PAND2X1_58/A 0.05fF
C2120 POR2X1_805/CTRL PAND2X1_90/Y 0.05fF
C2121 POR2X1_24/Y VDD 0.18fF
C2122 POR2X1_124/O POR2X1_556/A 0.01fF
C2123 PAND2X1_285/a_16_344# PAND2X1_805/A 0.02fF
C2124 POR2X1_679/Y VDD 0.00fF
C2125 POR2X1_814/A POR2X1_786/Y 0.10fF
C2126 POR2X1_65/CTRL2 PAND2X1_6/A 0.02fF
C2127 POR2X1_661/A POR2X1_725/Y 0.01fF
C2128 POR2X1_119/Y POR2X1_184/a_16_28# 0.08fF
C2129 PAND2X1_267/B PAND2X1_215/B 0.04fF
C2130 POR2X1_77/CTRL POR2X1_13/A 0.01fF
C2131 POR2X1_66/B POR2X1_14/Y 0.00fF
C2132 PAND2X1_631/A POR2X1_39/B 0.03fF
C2133 POR2X1_769/O PAND2X1_52/B 0.01fF
C2134 POR2X1_648/Y POR2X1_407/Y 0.07fF
C2135 POR2X1_260/B INPUT_0 0.15fF
C2136 POR2X1_496/Y PAND2X1_513/CTRL 0.06fF
C2137 PAND2X1_90/A POR2X1_341/A 0.07fF
C2138 PAND2X1_57/B PAND2X1_248/CTRL2 0.03fF
C2139 PAND2X1_237/O VDD 0.00fF
C2140 POR2X1_665/CTRL PAND2X1_645/B 0.08fF
C2141 PAND2X1_454/O PAND2X1_454/B 0.00fF
C2142 POR2X1_18/a_76_344# D_INPUT_6 0.00fF
C2143 POR2X1_807/CTRL VDD 0.00fF
C2144 POR2X1_475/A POR2X1_590/A 0.06fF
C2145 PAND2X1_55/Y PAND2X1_67/CTRL2 0.01fF
C2146 POR2X1_636/a_16_28# POR2X1_750/B 0.03fF
C2147 POR2X1_841/a_16_28# POR2X1_733/A 0.08fF
C2148 POR2X1_78/A POR2X1_807/A 0.02fF
C2149 POR2X1_13/A PAND2X1_776/Y 0.09fF
C2150 POR2X1_848/O POR2X1_713/B 0.01fF
C2151 POR2X1_688/O PAND2X1_32/B 0.01fF
C2152 POR2X1_20/B PAND2X1_566/Y 0.03fF
C2153 POR2X1_814/A PAND2X1_163/CTRL 0.06fF
C2154 POR2X1_515/a_16_28# PAND2X1_93/B 0.03fF
C2155 POR2X1_634/A PAND2X1_41/B 0.63fF
C2156 POR2X1_141/Y POR2X1_330/Y 0.05fF
C2157 POR2X1_316/Y PAND2X1_840/Y 0.05fF
C2158 POR2X1_48/A PAND2X1_785/Y 0.03fF
C2159 PAND2X1_93/B PAND2X1_386/Y 0.04fF
C2160 PAND2X1_16/CTRL POR2X1_630/A 0.00fF
C2161 PAND2X1_23/Y POR2X1_76/A 0.02fF
C2162 POR2X1_633/A PAND2X1_278/a_16_344# 0.02fF
C2163 PAND2X1_277/O POR2X1_546/A 0.05fF
C2164 POR2X1_78/B POR2X1_660/Y 0.03fF
C2165 POR2X1_32/A POR2X1_497/Y 0.01fF
C2166 POR2X1_43/CTRL POR2X1_39/B 0.01fF
C2167 POR2X1_337/Y POR2X1_181/A 0.03fF
C2168 PAND2X1_72/A PAND2X1_179/CTRL2 0.02fF
C2169 PAND2X1_816/CTRL POR2X1_862/A 0.02fF
C2170 POR2X1_467/Y POR2X1_798/O 0.04fF
C2171 POR2X1_411/B PAND2X1_570/a_76_28# 0.01fF
C2172 POR2X1_201/O POR2X1_61/Y 0.00fF
C2173 POR2X1_84/A POR2X1_294/B 0.14fF
C2174 POR2X1_821/CTRL POR2X1_669/B 0.01fF
C2175 POR2X1_831/a_76_344# POR2X1_513/Y 0.01fF
C2176 PAND2X1_413/a_56_28# INPUT_0 0.00fF
C2177 POR2X1_267/A POR2X1_547/B 0.02fF
C2178 POR2X1_72/O POR2X1_72/B 0.19fF
C2179 POR2X1_596/A POR2X1_678/O 0.01fF
C2180 PAND2X1_425/Y INPUT_6 1.79fF
C2181 POR2X1_624/Y POR2X1_804/A 0.10fF
C2182 PAND2X1_265/CTRL2 INPUT_0 0.06fF
C2183 POR2X1_254/Y POR2X1_241/B 0.08fF
C2184 PAND2X1_849/O POR2X1_60/Y 0.02fF
C2185 POR2X1_96/A POR2X1_669/B 0.44fF
C2186 PAND2X1_471/CTRL2 POR2X1_14/Y 0.00fF
C2187 POR2X1_315/a_16_28# POR2X1_257/A 0.07fF
C2188 POR2X1_20/B POR2X1_245/O 0.09fF
C2189 POR2X1_220/Y POR2X1_555/B 0.03fF
C2190 POR2X1_314/a_56_344# POR2X1_48/A 0.00fF
C2191 POR2X1_633/A VDD 0.28fF
C2192 INPUT_2 POR2X1_126/CTRL 0.01fF
C2193 POR2X1_441/Y PAND2X1_551/O 0.02fF
C2194 POR2X1_556/A POR2X1_510/Y 0.06fF
C2195 POR2X1_728/CTRL2 POR2X1_330/Y 0.01fF
C2196 POR2X1_566/A PAND2X1_230/CTRL 0.29fF
C2197 POR2X1_76/CTRL POR2X1_573/A 0.01fF
C2198 POR2X1_407/A PAND2X1_93/B 0.07fF
C2199 PAND2X1_630/O POR2X1_48/A 0.04fF
C2200 POR2X1_251/A PAND2X1_553/A 0.03fF
C2201 POR2X1_511/Y PAND2X1_513/CTRL2 0.10fF
C2202 POR2X1_274/A PAND2X1_96/B 0.03fF
C2203 POR2X1_84/B POR2X1_84/Y 0.03fF
C2204 POR2X1_315/Y POR2X1_20/B 2.06fF
C2205 PAND2X1_607/CTRL POR2X1_294/A 0.03fF
C2206 POR2X1_565/B POR2X1_78/A -0.00fF
C2207 PAND2X1_241/CTRL POR2X1_102/Y 0.01fF
C2208 POR2X1_14/Y POR2X1_395/CTRL 0.01fF
C2209 POR2X1_855/B POR2X1_803/CTRL2 0.01fF
C2210 POR2X1_186/Y VDD 4.70fF
C2211 POR2X1_48/A PAND2X1_324/CTRL2 0.05fF
C2212 PAND2X1_771/Y PAND2X1_569/A 0.07fF
C2213 POR2X1_676/Y POR2X1_750/B 0.01fF
C2214 POR2X1_556/A POR2X1_276/Y 0.04fF
C2215 POR2X1_270/Y PAND2X1_69/A 0.03fF
C2216 POR2X1_220/Y POR2X1_330/Y 0.08fF
C2217 POR2X1_130/A PAND2X1_41/B 0.17fF
C2218 POR2X1_60/A PAND2X1_592/Y 0.03fF
C2219 PAND2X1_90/A PAND2X1_77/O 0.01fF
C2220 POR2X1_60/A PAND2X1_174/CTRL2 0.03fF
C2221 POR2X1_285/Y POR2X1_294/B 0.03fF
C2222 POR2X1_449/CTRL PAND2X1_90/Y 0.34fF
C2223 POR2X1_236/CTRL2 POR2X1_236/Y 0.01fF
C2224 POR2X1_41/B POR2X1_495/CTRL2 0.05fF
C2225 POR2X1_645/CTRL PAND2X1_90/Y 0.07fF
C2226 POR2X1_42/CTRL POR2X1_37/Y 0.01fF
C2227 POR2X1_760/A POR2X1_394/A 0.07fF
C2228 D_INPUT_0 POR2X1_576/Y 0.01fF
C2229 POR2X1_566/A PAND2X1_41/B 0.13fF
C2230 POR2X1_118/CTRL2 POR2X1_32/A 0.01fF
C2231 PAND2X1_463/CTRL POR2X1_7/B 0.01fF
C2232 POR2X1_96/A PAND2X1_231/CTRL 0.01fF
C2233 PAND2X1_96/B PAND2X1_594/CTRL2 0.01fF
C2234 POR2X1_72/B PAND2X1_364/B 0.07fF
C2235 POR2X1_66/B POR2X1_55/Y 0.03fF
C2236 POR2X1_777/B PAND2X1_372/O 0.02fF
C2237 POR2X1_49/Y POR2X1_627/Y 0.11fF
C2238 POR2X1_236/O VDD 0.00fF
C2239 POR2X1_407/A POR2X1_78/A 0.29fF
C2240 POR2X1_179/O POR2X1_102/Y 0.02fF
C2241 POR2X1_378/CTRL2 POR2X1_55/Y 0.00fF
C2242 PAND2X1_90/A POR2X1_500/A 0.03fF
C2243 POR2X1_504/Y POR2X1_628/CTRL2 0.01fF
C2244 PAND2X1_36/O PAND2X1_32/B 0.04fF
C2245 POR2X1_389/A POR2X1_66/A 0.04fF
C2246 POR2X1_423/Y POR2X1_256/a_16_28# 0.02fF
C2247 PAND2X1_472/A POR2X1_102/Y 0.03fF
C2248 POR2X1_96/A POR2X1_230/O 0.02fF
C2249 POR2X1_43/B PAND2X1_244/O 0.03fF
C2250 POR2X1_88/a_16_28# POR2X1_7/A 0.03fF
C2251 PAND2X1_20/A POR2X1_574/a_56_344# 0.00fF
C2252 POR2X1_60/A PAND2X1_370/CTRL 0.29fF
C2253 PAND2X1_845/O POR2X1_83/B 0.01fF
C2254 POR2X1_123/O PAND2X1_41/B 0.17fF
C2255 POR2X1_152/a_16_28# POR2X1_669/B 0.06fF
C2256 POR2X1_351/Y PAND2X1_20/A 0.07fF
C2257 POR2X1_29/A POR2X1_68/B 0.05fF
C2258 POR2X1_48/A PAND2X1_656/A 0.03fF
C2259 PAND2X1_848/CTRL2 POR2X1_38/B 0.03fF
C2260 PAND2X1_319/B PAND2X1_220/A 0.03fF
C2261 POR2X1_502/A POR2X1_794/CTRL2 0.11fF
C2262 POR2X1_201/O POR2X1_35/Y 0.01fF
C2263 POR2X1_188/A PAND2X1_816/a_56_28# 0.00fF
C2264 PAND2X1_51/O POR2X1_635/A 0.02fF
C2265 POR2X1_188/A PAND2X1_536/CTRL 0.01fF
C2266 POR2X1_590/A POR2X1_447/O 0.18fF
C2267 PAND2X1_520/O VDD 0.00fF
C2268 POR2X1_241/B POR2X1_341/Y 0.01fF
C2269 POR2X1_624/Y POR2X1_6/O 0.02fF
C2270 POR2X1_186/Y POR2X1_741/Y 0.19fF
C2271 POR2X1_864/CTRL2 PAND2X1_32/B 0.01fF
C2272 POR2X1_411/B PAND2X1_508/Y 0.03fF
C2273 PAND2X1_65/Y POR2X1_294/B 0.01fF
C2274 POR2X1_230/Y VDD 0.03fF
C2275 POR2X1_376/Y POR2X1_55/Y 0.02fF
C2276 PAND2X1_212/B PAND2X1_388/Y 0.05fF
C2277 POR2X1_52/A PAND2X1_209/CTRL 0.01fF
C2278 PAND2X1_712/CTRL2 PAND2X1_707/Y 0.01fF
C2279 POR2X1_96/A POR2X1_329/CTRL2 0.00fF
C2280 POR2X1_483/A POR2X1_795/CTRL 0.01fF
C2281 PAND2X1_20/A POR2X1_844/CTRL 0.01fF
C2282 POR2X1_3/A POR2X1_83/B 0.04fF
C2283 POR2X1_669/B POR2X1_7/A 0.24fF
C2284 PAND2X1_641/CTRL2 POR2X1_263/Y 0.01fF
C2285 PAND2X1_137/Y POR2X1_13/A 0.01fF
C2286 POR2X1_653/O POR2X1_661/B 0.01fF
C2287 POR2X1_653/a_56_344# POR2X1_652/Y 0.01fF
C2288 POR2X1_51/A POR2X1_22/O 0.01fF
C2289 PAND2X1_41/B POR2X1_844/B 0.03fF
C2290 POR2X1_135/Y POR2X1_42/Y 0.03fF
C2291 PAND2X1_94/A D_INPUT_0 0.10fF
C2292 PAND2X1_725/A PAND2X1_725/B 0.04fF
C2293 POR2X1_186/Y PAND2X1_32/B 0.03fF
C2294 PAND2X1_556/B POR2X1_55/Y 0.03fF
C2295 POR2X1_338/CTRL PAND2X1_20/A 0.01fF
C2296 PAND2X1_6/Y POR2X1_850/A 0.01fF
C2297 PAND2X1_55/Y INPUT_0 0.03fF
C2298 POR2X1_635/A PAND2X1_3/B 0.00fF
C2299 PAND2X1_94/A POR2X1_55/CTRL 0.01fF
C2300 POR2X1_76/Y POR2X1_193/A 0.03fF
C2301 POR2X1_549/A VDD 0.14fF
C2302 POR2X1_76/Y POR2X1_579/Y 0.02fF
C2303 POR2X1_48/A PAND2X1_348/A 0.07fF
C2304 PAND2X1_216/CTRL PAND2X1_364/B 0.03fF
C2305 PAND2X1_602/Y VDD 0.17fF
C2306 PAND2X1_90/A PAND2X1_38/O 0.01fF
C2307 POR2X1_459/CTRL POR2X1_459/A 0.00fF
C2308 POR2X1_121/A VDD 0.40fF
C2309 POR2X1_863/CTRL2 POR2X1_855/Y 0.01fF
C2310 POR2X1_508/CTRL POR2X1_192/Y 0.14fF
C2311 POR2X1_157/CTRL INPUT_5 0.01fF
C2312 PAND2X1_554/a_16_344# PAND2X1_348/Y 0.03fF
C2313 PAND2X1_211/CTRL PAND2X1_352/Y 0.01fF
C2314 PAND2X1_254/Y POR2X1_55/Y 0.05fF
C2315 PAND2X1_394/CTRL POR2X1_215/A 0.04fF
C2316 D_INPUT_3 POR2X1_611/CTRL 0.01fF
C2317 POR2X1_78/B PAND2X1_697/O 0.01fF
C2318 PAND2X1_651/Y POR2X1_497/Y 1.96fF
C2319 PAND2X1_48/B POR2X1_784/A 0.03fF
C2320 POR2X1_832/a_16_28# POR2X1_832/B -0.00fF
C2321 POR2X1_113/Y POR2X1_392/B 0.01fF
C2322 POR2X1_334/Y POR2X1_66/A 0.07fF
C2323 POR2X1_129/CTRL POR2X1_129/Y 0.08fF
C2324 POR2X1_23/Y POR2X1_75/Y 0.04fF
C2325 PAND2X1_242/CTRL2 POR2X1_7/B 0.00fF
C2326 PAND2X1_387/CTRL PAND2X1_60/B 0.01fF
C2327 POR2X1_672/O VDD 0.00fF
C2328 POR2X1_271/B PAND2X1_841/Y 0.03fF
C2329 POR2X1_119/Y PAND2X1_477/CTRL 0.01fF
C2330 POR2X1_423/Y PAND2X1_349/A 0.06fF
C2331 POR2X1_474/CTRL POR2X1_362/A 0.03fF
C2332 POR2X1_474/O POR2X1_276/Y 0.01fF
C2333 POR2X1_406/Y PAND2X1_734/CTRL 0.01fF
C2334 POR2X1_66/B PAND2X1_232/CTRL 0.01fF
C2335 POR2X1_579/Y POR2X1_740/Y 0.05fF
C2336 PAND2X1_845/CTRL2 PAND2X1_35/Y 0.01fF
C2337 POR2X1_57/A POR2X1_399/CTRL 0.05fF
C2338 POR2X1_390/B POR2X1_390/a_16_28# 0.07fF
C2339 D_INPUT_3 POR2X1_5/Y 0.82fF
C2340 POR2X1_120/a_16_28# POR2X1_712/Y 0.00fF
C2341 POR2X1_215/A POR2X1_330/Y 0.23fF
C2342 POR2X1_625/a_76_344# POR2X1_93/A 0.01fF
C2343 POR2X1_850/CTRL POR2X1_362/B 0.01fF
C2344 PAND2X1_52/a_56_28# PAND2X1_72/A 0.00fF
C2345 POR2X1_383/A POR2X1_860/A 0.04fF
C2346 POR2X1_366/Y POR2X1_317/O 0.03fF
C2347 POR2X1_656/CTRL2 POR2X1_737/A 0.01fF
C2348 POR2X1_782/m4_208_n4# POR2X1_260/A 0.09fF
C2349 POR2X1_119/Y POR2X1_118/Y 0.11fF
C2350 POR2X1_497/Y PAND2X1_844/B 0.58fF
C2351 PAND2X1_48/B POR2X1_732/B 0.03fF
C2352 POR2X1_614/A POR2X1_76/Y 0.02fF
C2353 POR2X1_278/Y PAND2X1_347/CTRL2 0.00fF
C2354 PAND2X1_440/O POR2X1_150/Y 0.03fF
C2355 POR2X1_835/B POR2X1_568/A 0.05fF
C2356 POR2X1_548/CTRL2 PAND2X1_63/B 0.01fF
C2357 POR2X1_590/A POR2X1_557/B 0.14fF
C2358 POR2X1_68/B POR2X1_546/A 0.03fF
C2359 POR2X1_619/Y VDD -0.00fF
C2360 POR2X1_73/Y PAND2X1_549/O 0.07fF
C2361 POR2X1_61/Y POR2X1_259/CTRL2 0.03fF
C2362 PAND2X1_679/CTRL2 POR2X1_687/A 0.03fF
C2363 PAND2X1_865/Y PAND2X1_489/O 0.00fF
C2364 POR2X1_52/A POR2X1_526/CTRL 0.03fF
C2365 POR2X1_57/A PAND2X1_738/Y 0.09fF
C2366 POR2X1_71/Y POR2X1_816/A 0.03fF
C2367 POR2X1_356/A POR2X1_535/a_16_28# 0.04fF
C2368 PAND2X1_631/A POR2X1_48/A 0.08fF
C2369 PAND2X1_402/B POR2X1_236/Y 0.01fF
C2370 POR2X1_633/m4_208_n4# PAND2X1_52/B 0.09fF
C2371 PAND2X1_471/O PAND2X1_241/Y 0.03fF
C2372 POR2X1_42/Y POR2X1_816/A 0.05fF
C2373 POR2X1_614/A POR2X1_740/Y 0.07fF
C2374 POR2X1_397/Y PAND2X1_720/O 0.01fF
C2375 PAND2X1_94/A PAND2X1_90/Y 0.10fF
C2376 POR2X1_25/Y POR2X1_83/B 2.73fF
C2377 POR2X1_566/A POR2X1_228/Y 0.01fF
C2378 POR2X1_502/A PAND2X1_60/B 0.15fF
C2379 POR2X1_356/A POR2X1_209/A 4.14fF
C2380 POR2X1_83/B POR2X1_701/CTRL 0.01fF
C2381 PAND2X1_434/CTRL2 VDD 0.00fF
C2382 POR2X1_542/B POR2X1_662/Y 0.00fF
C2383 PAND2X1_784/CTRL PAND2X1_778/Y 0.01fF
C2384 POR2X1_16/A PAND2X1_204/CTRL 0.25fF
C2385 POR2X1_186/Y PAND2X1_746/CTRL 0.01fF
C2386 PAND2X1_478/Y POR2X1_394/A 0.01fF
C2387 POR2X1_251/Y PAND2X1_843/Y 0.01fF
C2388 POR2X1_763/Y POR2X1_152/Y 0.05fF
C2389 PAND2X1_23/Y POR2X1_540/A 0.03fF
C2390 POR2X1_347/CTRL POR2X1_296/B 0.01fF
C2391 POR2X1_383/A POR2X1_327/CTRL2 0.01fF
C2392 PAND2X1_490/CTRL2 PAND2X1_6/Y 0.00fF
C2393 POR2X1_625/Y POR2X1_283/A 0.03fF
C2394 POR2X1_57/A PAND2X1_839/CTRL 0.01fF
C2395 POR2X1_504/Y POR2X1_129/Y 0.02fF
C2396 POR2X1_130/A POR2X1_561/CTRL 0.01fF
C2397 POR2X1_3/A PAND2X1_709/O 0.15fF
C2398 PAND2X1_562/B PAND2X1_853/B 0.19fF
C2399 POR2X1_141/O POR2X1_244/Y 0.02fF
C2400 PAND2X1_6/A PAND2X1_69/A 1.46fF
C2401 POR2X1_481/A PAND2X1_336/O 0.02fF
C2402 PAND2X1_476/A POR2X1_60/A 7.42fF
C2403 PAND2X1_858/O PAND2X1_390/Y 0.02fF
C2404 POR2X1_835/O POR2X1_835/B 0.01fF
C2405 POR2X1_463/Y PAND2X1_700/O 0.00fF
C2406 POR2X1_335/O POR2X1_260/A 0.18fF
C2407 POR2X1_514/Y POR2X1_137/Y 0.01fF
C2408 POR2X1_90/Y POR2X1_321/a_56_344# 0.00fF
C2409 POR2X1_36/B POR2X1_22/A 0.10fF
C2410 POR2X1_532/A POR2X1_804/B 0.01fF
C2411 PAND2X1_197/Y PAND2X1_656/A 0.01fF
C2412 PAND2X1_270/CTRL2 POR2X1_184/Y 0.10fF
C2413 POR2X1_376/B PAND2X1_508/Y 0.03fF
C2414 POR2X1_413/A PAND2X1_656/A 0.06fF
C2415 POR2X1_480/A PAND2X1_142/CTRL 0.03fF
C2416 POR2X1_93/A PAND2X1_6/A 0.81fF
C2417 POR2X1_41/B POR2X1_41/CTRL2 0.01fF
C2418 POR2X1_559/B PAND2X1_90/A 0.02fF
C2419 PAND2X1_531/CTRL POR2X1_549/B 0.02fF
C2420 POR2X1_218/A POR2X1_361/CTRL 0.01fF
C2421 POR2X1_572/B POR2X1_361/a_16_28# 0.02fF
C2422 POR2X1_539/A PAND2X1_23/Y 0.03fF
C2423 POR2X1_16/A POR2X1_46/Y 0.03fF
C2424 PAND2X1_182/B VDD 0.06fF
C2425 POR2X1_394/A PAND2X1_719/CTRL 0.03fF
C2426 POR2X1_614/A PAND2X1_312/CTRL2 0.03fF
C2427 POR2X1_68/A PAND2X1_306/a_16_344# 0.03fF
C2428 POR2X1_23/Y PAND2X1_332/Y 0.04fF
C2429 POR2X1_855/B POR2X1_800/A 3.39fF
C2430 POR2X1_440/Y POR2X1_740/Y 0.02fF
C2431 PAND2X1_219/B POR2X1_7/Y 0.01fF
C2432 POR2X1_740/Y POR2X1_702/a_16_28# 0.05fF
C2433 POR2X1_65/A POR2X1_518/CTRL2 0.03fF
C2434 PAND2X1_168/Y PAND2X1_326/B 0.34fF
C2435 POR2X1_123/A POR2X1_391/Y 0.07fF
C2436 POR2X1_13/A PAND2X1_853/B 0.03fF
C2437 PAND2X1_741/a_16_344# PAND2X1_853/B 0.02fF
C2438 PAND2X1_291/O PAND2X1_69/A 0.05fF
C2439 POR2X1_119/Y PAND2X1_403/Y 0.03fF
C2440 POR2X1_83/Y POR2X1_5/Y 0.00fF
C2441 PAND2X1_631/A PAND2X1_513/O 0.03fF
C2442 POR2X1_809/Y POR2X1_812/B 0.51fF
C2443 POR2X1_811/B PAND2X1_56/A 0.02fF
C2444 PAND2X1_548/O POR2X1_530/Y 0.00fF
C2445 POR2X1_833/CTRL POR2X1_260/A 0.01fF
C2446 POR2X1_366/A POR2X1_112/Y 0.34fF
C2447 POR2X1_228/Y POR2X1_573/A 0.03fF
C2448 POR2X1_30/CTRL2 POR2X1_260/A 0.02fF
C2449 POR2X1_57/A POR2X1_823/Y 0.00fF
C2450 POR2X1_57/A POR2X1_136/Y 0.00fF
C2451 POR2X1_614/A PAND2X1_253/CTRL 0.01fF
C2452 PAND2X1_358/A PAND2X1_341/CTRL2 0.01fF
C2453 POR2X1_68/A POR2X1_456/B 0.06fF
C2454 POR2X1_495/CTRL2 POR2X1_77/Y 0.01fF
C2455 PAND2X1_93/B PAND2X1_628/CTRL2 0.00fF
C2456 POR2X1_615/CTRL POR2X1_39/B 0.01fF
C2457 POR2X1_101/Y PAND2X1_69/A 0.12fF
C2458 POR2X1_8/Y PAND2X1_35/O 0.02fF
C2459 PAND2X1_358/A POR2X1_55/Y 0.10fF
C2460 POR2X1_220/Y POR2X1_337/Y 0.48fF
C2461 POR2X1_677/Y POR2X1_271/O 0.00fF
C2462 POR2X1_532/A POR2X1_710/Y 0.02fF
C2463 POR2X1_459/Y POR2X1_460/Y 0.08fF
C2464 POR2X1_719/O PAND2X1_60/B 0.01fF
C2465 PAND2X1_653/Y POR2X1_7/O 0.01fF
C2466 POR2X1_542/Y VDD 0.14fF
C2467 PAND2X1_96/O PAND2X1_58/A 0.17fF
C2468 POR2X1_579/Y PAND2X1_171/O 0.16fF
C2469 POR2X1_96/A PAND2X1_538/a_76_28# 0.01fF
C2470 POR2X1_49/Y PAND2X1_847/CTRL2 0.00fF
C2471 PAND2X1_185/O POR2X1_77/Y 0.04fF
C2472 POR2X1_567/B PAND2X1_437/O 0.02fF
C2473 POR2X1_8/Y PAND2X1_227/CTRL2 0.01fF
C2474 POR2X1_334/Y POR2X1_222/Y 0.07fF
C2475 POR2X1_265/Y POR2X1_406/O 0.13fF
C2476 PAND2X1_290/O PAND2X1_85/Y 0.11fF
C2477 POR2X1_43/Y PAND2X1_195/CTRL 0.02fF
C2478 POR2X1_257/A POR2X1_431/O 0.01fF
C2479 POR2X1_25/Y POR2X1_47/CTRL 0.01fF
C2480 PAND2X1_218/A POR2X1_394/A 0.01fF
C2481 POR2X1_10/CTRL2 POR2X1_38/Y 0.03fF
C2482 GATE_479 POR2X1_158/Y 0.03fF
C2483 PAND2X1_662/Y POR2X1_413/A 0.01fF
C2484 POR2X1_433/Y POR2X1_129/Y 0.00fF
C2485 POR2X1_767/Y VDD 0.00fF
C2486 POR2X1_654/B PAND2X1_52/B 0.03fF
C2487 POR2X1_358/a_56_344# POR2X1_192/B 0.00fF
C2488 POR2X1_358/CTRL POR2X1_191/Y 0.11fF
C2489 PAND2X1_349/A PAND2X1_840/a_16_344# 0.01fF
C2490 POR2X1_567/A POR2X1_661/B 0.03fF
C2491 POR2X1_666/A POR2X1_77/Y 0.01fF
C2492 POR2X1_177/Y POR2X1_77/Y 0.00fF
C2493 POR2X1_137/Y POR2X1_773/B 0.05fF
C2494 POR2X1_316/Y PAND2X1_445/Y 0.03fF
C2495 PAND2X1_219/CTRL POR2X1_7/Y 0.01fF
C2496 POR2X1_203/CTRL2 PAND2X1_72/Y 0.01fF
C2497 POR2X1_804/A POR2X1_186/B 0.04fF
C2498 PAND2X1_364/m4_208_n4# PAND2X1_355/m4_208_n4# 0.13fF
C2499 POR2X1_394/A PAND2X1_509/CTRL2 0.05fF
C2500 POR2X1_16/A PAND2X1_350/O 0.00fF
C2501 PAND2X1_809/A PAND2X1_539/O 0.09fF
C2502 PAND2X1_209/A PAND2X1_162/A 0.29fF
C2503 POR2X1_634/A POR2X1_635/B 0.00fF
C2504 POR2X1_38/Y POR2X1_394/A 2.72fF
C2505 POR2X1_186/CTRL2 POR2X1_725/Y 0.05fF
C2506 POR2X1_334/Y POR2X1_532/A 0.46fF
C2507 POR2X1_111/Y POR2X1_136/Y 0.02fF
C2508 PAND2X1_291/O PAND2X1_824/B 0.04fF
C2509 POR2X1_118/a_16_28# POR2X1_153/Y 0.09fF
C2510 POR2X1_54/Y POR2X1_461/Y 0.00fF
C2511 POR2X1_57/A POR2X1_122/O 0.01fF
C2512 PAND2X1_9/Y POR2X1_24/Y 0.01fF
C2513 POR2X1_13/A POR2X1_80/O 0.15fF
C2514 POR2X1_648/Y POR2X1_807/a_16_28# 0.02fF
C2515 POR2X1_16/A PAND2X1_727/CTRL2 0.01fF
C2516 POR2X1_62/Y POR2X1_15/O 0.01fF
C2517 VDD POR2X1_717/B 0.22fF
C2518 PAND2X1_271/CTRL2 POR2X1_76/A 0.01fF
C2519 POR2X1_36/B POR2X1_328/O 0.01fF
C2520 POR2X1_639/Y PAND2X1_328/a_76_28# 0.02fF
C2521 PAND2X1_724/CTRL2 PAND2X1_326/B 0.01fF
C2522 POR2X1_119/Y POR2X1_91/Y 0.23fF
C2523 POR2X1_62/Y PAND2X1_656/A 0.01fF
C2524 PAND2X1_728/O PAND2X1_853/B 0.04fF
C2525 PAND2X1_101/B PAND2X1_99/Y 0.04fF
C2526 PAND2X1_60/B POR2X1_188/Y 0.03fF
C2527 VDD PAND2X1_146/CTRL 0.00fF
C2528 PAND2X1_70/O POR2X1_451/A 0.03fF
C2529 POR2X1_369/Y PAND2X1_388/Y 0.02fF
C2530 INPUT_1 POR2X1_394/A 0.14fF
C2531 POR2X1_183/Y POR2X1_39/B 0.10fF
C2532 POR2X1_509/a_16_28# PAND2X1_52/B 0.01fF
C2533 PAND2X1_649/A POR2X1_689/Y 0.03fF
C2534 PAND2X1_339/Y POR2X1_522/CTRL 0.01fF
C2535 PAND2X1_271/O PAND2X1_93/B 0.04fF
C2536 POR2X1_680/a_76_344# POR2X1_594/A 0.00fF
C2537 PAND2X1_52/B PAND2X1_145/CTRL 0.01fF
C2538 POR2X1_38/Y PAND2X1_198/CTRL2 0.00fF
C2539 PAND2X1_51/CTRL2 PAND2X1_3/B 0.01fF
C2540 POR2X1_840/O POR2X1_513/A 0.00fF
C2541 POR2X1_394/A POR2X1_153/Y 0.21fF
C2542 PAND2X1_60/CTRL POR2X1_66/A 0.01fF
C2543 POR2X1_188/Y POR2X1_737/CTRL 0.01fF
C2544 POR2X1_741/Y POR2X1_717/B 0.03fF
C2545 PAND2X1_93/B POR2X1_632/CTRL 0.01fF
C2546 POR2X1_553/A POR2X1_540/Y 0.00fF
C2547 PAND2X1_407/O POR2X1_409/B 0.03fF
C2548 PAND2X1_466/B POR2X1_669/B 0.03fF
C2549 POR2X1_327/Y POR2X1_741/A 0.01fF
C2550 POR2X1_63/Y POR2X1_83/B 0.30fF
C2551 PAND2X1_9/Y PAND2X1_15/a_16_344# 0.02fF
C2552 POR2X1_9/Y POR2X1_415/CTRL 0.05fF
C2553 POR2X1_387/Y POR2X1_372/CTRL 0.05fF
C2554 POR2X1_37/Y POR2X1_289/Y 0.02fF
C2555 PAND2X1_469/CTRL POR2X1_32/A 0.02fF
C2556 POR2X1_528/Y POR2X1_305/CTRL2 0.03fF
C2557 POR2X1_711/Y POR2X1_513/O 0.03fF
C2558 POR2X1_48/A POR2X1_416/A 0.01fF
C2559 POR2X1_717/B PAND2X1_32/B 0.00fF
C2560 POR2X1_241/a_16_28# POR2X1_776/A 0.03fF
C2561 POR2X1_124/CTRL2 POR2X1_137/Y 0.00fF
C2562 PAND2X1_96/B PAND2X1_96/O 0.01fF
C2563 POR2X1_353/Y POR2X1_443/CTRL2 0.01fF
C2564 POR2X1_96/B POR2X1_416/B 0.05fF
C2565 POR2X1_87/B POR2X1_38/B 0.01fF
C2566 POR2X1_129/CTRL POR2X1_37/Y 0.01fF
C2567 POR2X1_456/B POR2X1_169/A 0.03fF
C2568 POR2X1_648/Y POR2X1_779/a_16_28# 0.03fF
C2569 PAND2X1_633/CTRL POR2X1_826/Y 0.15fF
C2570 POR2X1_119/Y POR2X1_109/Y 0.03fF
C2571 POR2X1_60/A PAND2X1_207/CTRL 0.01fF
C2572 POR2X1_19/a_76_344# POR2X1_5/Y 0.01fF
C2573 POR2X1_99/A POR2X1_99/Y 0.01fF
C2574 PAND2X1_47/B PAND2X1_31/O 0.08fF
C2575 POR2X1_814/A PAND2X1_372/O 0.04fF
C2576 POR2X1_647/B POR2X1_389/Y 0.03fF
C2577 PAND2X1_510/B POR2X1_80/O 0.00fF
C2578 PAND2X1_143/m4_208_n4# PAND2X1_133/m4_208_n4# 0.05fF
C2579 PAND2X1_472/CTRL POR2X1_77/Y 0.01fF
C2580 POR2X1_48/A PAND2X1_564/B 0.03fF
C2581 POR2X1_195/O PAND2X1_41/Y 0.00fF
C2582 POR2X1_814/A POR2X1_193/CTRL2 0.04fF
C2583 POR2X1_52/A PAND2X1_464/B 0.06fF
C2584 POR2X1_66/B POR2X1_476/A 11.01fF
C2585 POR2X1_83/B POR2X1_427/O 0.06fF
C2586 PAND2X1_340/B POR2X1_381/CTRL2 0.01fF
C2587 PAND2X1_255/CTRL PAND2X1_69/A 0.03fF
C2588 PAND2X1_480/B POR2X1_20/B 0.05fF
C2589 POR2X1_729/O POR2X1_814/A 0.08fF
C2590 POR2X1_48/A POR2X1_615/CTRL 0.07fF
C2591 POR2X1_20/B POR2X1_754/A 0.03fF
C2592 POR2X1_150/Y POR2X1_7/B 0.05fF
C2593 POR2X1_13/A PAND2X1_796/B 0.01fF
C2594 PAND2X1_417/O PAND2X1_55/Y 0.09fF
C2595 POR2X1_389/A PAND2X1_607/CTRL 0.00fF
C2596 POR2X1_120/a_16_28# PAND2X1_39/B -0.00fF
C2597 POR2X1_163/O POR2X1_23/Y 0.01fF
C2598 PAND2X1_473/CTRL2 POR2X1_329/A 0.01fF
C2599 PAND2X1_793/Y POR2X1_257/A 0.05fF
C2600 POR2X1_66/A POR2X1_404/a_16_28# 0.02fF
C2601 POR2X1_438/Y PAND2X1_544/CTRL 0.01fF
C2602 POR2X1_285/Y POR2X1_643/A 0.03fF
C2603 POR2X1_423/Y POR2X1_32/A 0.03fF
C2604 PAND2X1_96/B PAND2X1_89/a_76_28# 0.02fF
C2605 POR2X1_295/m4_208_n4# POR2X1_90/Y 0.17fF
C2606 PAND2X1_796/CTRL2 PAND2X1_783/Y 0.01fF
C2607 PAND2X1_57/B PAND2X1_26/A 0.02fF
C2608 POR2X1_20/B PAND2X1_398/CTRL 0.01fF
C2609 PAND2X1_657/O PAND2X1_217/B 0.03fF
C2610 PAND2X1_474/Y POR2X1_23/Y 0.03fF
C2611 INPUT_3 POR2X1_42/Y 0.05fF
C2612 POR2X1_241/B PAND2X1_41/B 0.03fF
C2613 PAND2X1_205/A PAND2X1_579/B 0.03fF
C2614 POR2X1_294/CTRL POR2X1_294/B 0.01fF
C2615 POR2X1_485/Y PAND2X1_565/A 0.01fF
C2616 PAND2X1_557/A POR2X1_40/Y 0.03fF
C2617 POR2X1_861/m4_208_n4# POR2X1_499/A 0.08fF
C2618 POR2X1_13/A POR2X1_23/Y 0.17fF
C2619 POR2X1_547/CTRL2 POR2X1_624/Y 0.01fF
C2620 POR2X1_491/CTRL2 PAND2X1_558/Y 0.00fF
C2621 POR2X1_496/Y POR2X1_372/A 0.00fF
C2622 POR2X1_102/Y PAND2X1_803/A 0.03fF
C2623 POR2X1_774/Y POR2X1_866/CTRL 0.01fF
C2624 PAND2X1_56/Y POR2X1_446/B 0.05fF
C2625 POR2X1_23/Y PAND2X1_214/B 0.04fF
C2626 POR2X1_471/a_76_344# POR2X1_66/A 0.01fF
C2627 PAND2X1_57/B POR2X1_218/Y 0.07fF
C2628 PAND2X1_223/B VDD 0.09fF
C2629 POR2X1_23/Y PAND2X1_775/O 0.13fF
C2630 POR2X1_677/CTRL2 PAND2X1_390/Y 0.01fF
C2631 PAND2X1_219/A PAND2X1_733/Y 0.01fF
C2632 POR2X1_800/A POR2X1_808/a_56_344# 0.01fF
C2633 POR2X1_72/B POR2X1_427/Y 0.01fF
C2634 PAND2X1_404/Y PAND2X1_339/Y 0.03fF
C2635 PAND2X1_865/O POR2X1_329/A 0.04fF
C2636 PAND2X1_23/Y PAND2X1_94/CTRL 0.00fF
C2637 POR2X1_175/a_76_344# POR2X1_78/A 0.00fF
C2638 POR2X1_466/A PAND2X1_152/O 0.35fF
C2639 D_INPUT_0 PAND2X1_351/O 0.24fF
C2640 PAND2X1_436/A POR2X1_677/a_16_28# 0.08fF
C2641 POR2X1_866/B POR2X1_750/B 0.01fF
C2642 POR2X1_78/B POR2X1_400/CTRL 0.01fF
C2643 PAND2X1_39/B POR2X1_68/B 0.20fF
C2644 POR2X1_275/O D_INPUT_0 0.01fF
C2645 PAND2X1_48/B POR2X1_466/A 0.09fF
C2646 D_INPUT_3 POR2X1_612/CTRL2 0.03fF
C2647 PAND2X1_95/B PAND2X1_3/A 0.12fF
C2648 POR2X1_52/A POR2X1_751/A 0.01fF
C2649 POR2X1_57/A PAND2X1_838/B 0.04fF
C2650 PAND2X1_271/a_16_344# POR2X1_804/A 0.03fF
C2651 POR2X1_502/A PAND2X1_279/CTRL2 0.02fF
C2652 POR2X1_68/A PAND2X1_94/CTRL2 0.06fF
C2653 POR2X1_814/B POR2X1_461/a_76_344# 0.00fF
C2654 POR2X1_272/O POR2X1_272/Y 0.02fF
C2655 POR2X1_368/CTRL POR2X1_417/Y 0.00fF
C2656 POR2X1_114/B POR2X1_734/B 0.02fF
C2657 POR2X1_411/B POR2X1_283/A 1.04fF
C2658 PAND2X1_90/A POR2X1_29/A 5.89fF
C2659 PAND2X1_725/Y VDD 0.11fF
C2660 POR2X1_411/B PAND2X1_121/CTRL 0.01fF
C2661 POR2X1_48/A POR2X1_183/Y 0.03fF
C2662 PAND2X1_600/CTRL PAND2X1_32/B 0.03fF
C2663 POR2X1_68/A POR2X1_849/A 0.00fF
C2664 POR2X1_222/O POR2X1_724/A 0.04fF
C2665 POR2X1_457/O POR2X1_220/Y 0.01fF
C2666 PAND2X1_34/a_16_344# POR2X1_42/Y 0.01fF
C2667 POR2X1_625/O POR2X1_5/Y 0.07fF
C2668 POR2X1_433/Y POR2X1_37/Y 0.01fF
C2669 POR2X1_811/A POR2X1_796/CTRL2 0.00fF
C2670 POR2X1_155/O POR2X1_750/B 0.01fF
C2671 POR2X1_590/A POR2X1_740/Y 0.11fF
C2672 POR2X1_496/Y PAND2X1_658/B 0.04fF
C2673 POR2X1_41/B POR2X1_748/A 0.07fF
C2674 PAND2X1_118/CTRL PAND2X1_73/Y 0.01fF
C2675 PAND2X1_118/CTRL2 POR2X1_78/A 0.01fF
C2676 POR2X1_502/A POR2X1_750/B 2.08fF
C2677 PAND2X1_420/CTRL2 POR2X1_294/B 0.04fF
C2678 POR2X1_668/CTRL2 VDD 0.00fF
C2679 POR2X1_864/A POR2X1_260/A 0.01fF
C2680 POR2X1_13/A POR2X1_312/Y 0.02fF
C2681 PAND2X1_643/CTRL2 POR2X1_102/Y 0.03fF
C2682 PAND2X1_433/O POR2X1_78/A 0.03fF
C2683 POR2X1_697/CTRL2 POR2X1_236/Y 0.00fF
C2684 POR2X1_49/Y PAND2X1_661/CTRL 0.01fF
C2685 POR2X1_663/B POR2X1_703/A 0.05fF
C2686 PAND2X1_57/B POR2X1_710/A 0.51fF
C2687 POR2X1_220/Y POR2X1_543/A 0.03fF
C2688 POR2X1_590/A POR2X1_732/O 0.10fF
C2689 POR2X1_750/B PAND2X1_176/O 0.04fF
C2690 PAND2X1_57/B PAND2X1_597/O 0.15fF
C2691 POR2X1_411/B POR2X1_385/a_16_28# 0.02fF
C2692 POR2X1_866/A POR2X1_777/Y 0.10fF
C2693 POR2X1_493/A PAND2X1_60/B 0.02fF
C2694 POR2X1_504/Y POR2X1_293/Y 0.03fF
C2695 PAND2X1_139/B PAND2X1_140/Y 0.04fF
C2696 POR2X1_254/CTRL2 POR2X1_222/Y 0.03fF
C2697 POR2X1_407/A POR2X1_307/O 0.02fF
C2698 POR2X1_260/B POR2X1_796/A 0.03fF
C2699 POR2X1_327/Y POR2X1_556/A 0.03fF
C2700 POR2X1_424/Y PAND2X1_308/Y 0.03fF
C2701 POR2X1_840/B POR2X1_296/B 0.03fF
C2702 POR2X1_263/Y PAND2X1_338/B 0.03fF
C2703 POR2X1_368/CTRL2 POR2X1_13/A 0.00fF
C2704 POR2X1_669/B POR2X1_38/Y 0.05fF
C2705 PAND2X1_23/O PAND2X1_55/Y 0.01fF
C2706 POR2X1_123/Y POR2X1_78/A 0.01fF
C2707 POR2X1_275/a_76_344# PAND2X1_390/Y 0.00fF
C2708 PAND2X1_137/a_76_28# PAND2X1_354/A 0.01fF
C2709 POR2X1_567/B POR2X1_854/B 0.05fF
C2710 POR2X1_37/Y PAND2X1_840/CTRL 0.01fF
C2711 PAND2X1_319/B POR2X1_32/A 0.03fF
C2712 POR2X1_263/Y POR2X1_235/CTRL 0.01fF
C2713 POR2X1_114/B POR2X1_330/Y 0.05fF
C2714 POR2X1_88/Y VDD 0.12fF
C2715 POR2X1_865/a_56_344# POR2X1_590/A 0.00fF
C2716 PAND2X1_573/a_76_28# PAND2X1_499/Y 0.03fF
C2717 POR2X1_23/Y PAND2X1_510/B 0.02fF
C2718 POR2X1_777/B PAND2X1_536/O 0.04fF
C2719 POR2X1_260/B POR2X1_332/CTRL2 0.01fF
C2720 POR2X1_423/Y POR2X1_184/Y 0.06fF
C2721 PAND2X1_20/A POR2X1_68/B 0.23fF
C2722 POR2X1_78/A POR2X1_216/CTRL 0.01fF
C2723 PAND2X1_16/O D_GATE_222 0.02fF
C2724 POR2X1_498/CTRL PAND2X1_735/Y 0.08fF
C2725 POR2X1_605/A POR2X1_605/a_16_28# 0.05fF
C2726 POR2X1_332/B POR2X1_220/Y 0.03fF
C2727 POR2X1_188/A POR2X1_513/Y 0.03fF
C2728 POR2X1_241/B POR2X1_228/Y 0.08fF
C2729 POR2X1_814/B PAND2X1_411/O 0.18fF
C2730 PAND2X1_651/Y POR2X1_423/Y 0.06fF
C2731 POR2X1_388/O POR2X1_750/B 0.02fF
C2732 POR2X1_555/B POR2X1_222/A 0.02fF
C2733 POR2X1_829/a_56_344# POR2X1_761/Y 0.00fF
C2734 PAND2X1_720/O POR2X1_667/Y 0.00fF
C2735 PAND2X1_73/Y PAND2X1_63/B 0.01fF
C2736 PAND2X1_58/A PAND2X1_306/a_16_344# 0.01fF
C2737 POR2X1_164/CTRL2 POR2X1_376/B 0.00fF
C2738 POR2X1_41/B POR2X1_79/Y 0.03fF
C2739 POR2X1_333/CTRL2 POR2X1_241/B 0.01fF
C2740 D_GATE_222 PAND2X1_164/CTRL 0.08fF
C2741 POR2X1_383/A POR2X1_121/B 0.14fF
C2742 PAND2X1_319/B POR2X1_417/Y 2.52fF
C2743 PAND2X1_90/A POR2X1_546/A 2.80fF
C2744 PAND2X1_652/A PAND2X1_804/A 0.01fF
C2745 POR2X1_302/CTRL POR2X1_114/B 0.01fF
C2746 POR2X1_539/a_16_28# PAND2X1_93/B 0.03fF
C2747 PAND2X1_6/Y PAND2X1_65/B 1.01fF
C2748 POR2X1_307/Y POR2X1_513/B 0.01fF
C2749 PAND2X1_231/CTRL POR2X1_38/Y 0.04fF
C2750 POR2X1_528/Y POR2X1_420/Y 0.00fF
C2751 POR2X1_865/B POR2X1_734/A 0.07fF
C2752 POR2X1_549/CTRL POR2X1_68/B 0.00fF
C2753 POR2X1_66/B POR2X1_366/A 0.03fF
C2754 POR2X1_814/B POR2X1_68/B 0.15fF
C2755 POR2X1_293/Y POR2X1_586/O 0.34fF
C2756 PAND2X1_798/B PAND2X1_580/B 0.01fF
C2757 POR2X1_322/Y PAND2X1_168/Y 0.33fF
C2758 POR2X1_461/A POR2X1_713/B 0.35fF
C2759 INPUT_1 POR2X1_669/B 0.32fF
C2760 PAND2X1_742/O POR2X1_283/A 0.05fF
C2761 POR2X1_241/B POR2X1_502/CTRL 0.01fF
C2762 PAND2X1_76/Y POR2X1_73/Y 2.53fF
C2763 POR2X1_750/B PAND2X1_158/CTRL2 0.01fF
C2764 PAND2X1_96/B POR2X1_573/O 0.16fF
C2765 POR2X1_417/O POR2X1_5/Y 0.02fF
C2766 PAND2X1_535/Y PAND2X1_805/A 0.05fF
C2767 POR2X1_378/A POR2X1_94/A 0.11fF
C2768 POR2X1_230/O POR2X1_38/Y -0.02fF
C2769 PAND2X1_23/Y PAND2X1_371/CTRL 0.06fF
C2770 PAND2X1_48/B PAND2X1_371/O 0.15fF
C2771 POR2X1_351/Y VDD -0.00fF
C2772 POR2X1_862/B PAND2X1_60/B 0.03fF
C2773 POR2X1_68/A PAND2X1_57/B 0.57fF
C2774 POR2X1_504/Y POR2X1_408/Y 0.03fF
C2775 POR2X1_208/A PAND2X1_41/B 0.04fF
C2776 POR2X1_593/B POR2X1_592/O 0.01fF
C2777 POR2X1_343/Y PAND2X1_256/a_56_28# 0.00fF
C2778 POR2X1_581/CTRL2 INPUT_5 0.01fF
C2779 POR2X1_850/O POR2X1_850/A 0.01fF
C2780 POR2X1_750/B POR2X1_799/CTRL 0.00fF
C2781 POR2X1_669/B POR2X1_153/Y 0.17fF
C2782 POR2X1_102/Y PAND2X1_722/CTRL2 0.01fF
C2783 PAND2X1_857/A POR2X1_65/A 0.01fF
C2784 PAND2X1_340/CTRL POR2X1_7/A 0.01fF
C2785 PAND2X1_213/Y POR2X1_236/Y 0.03fF
C2786 POR2X1_844/CTRL VDD -0.00fF
C2787 PAND2X1_294/CTRL2 POR2X1_39/B 0.03fF
C2788 POR2X1_349/Y POR2X1_532/A 0.11fF
C2789 POR2X1_573/a_16_28# POR2X1_573/A 0.10fF
C2790 POR2X1_575/B POR2X1_501/CTRL 0.02fF
C2791 POR2X1_590/A POR2X1_774/A 0.03fF
C2792 POR2X1_376/B POR2X1_283/A 0.04fF
C2793 POR2X1_433/Y POR2X1_293/Y 0.03fF
C2794 POR2X1_66/B PAND2X1_127/O 0.03fF
C2795 PAND2X1_675/A POR2X1_42/Y 0.03fF
C2796 POR2X1_96/A PAND2X1_734/O 0.01fF
C2797 POR2X1_25/Y POR2X1_59/a_16_28# -0.00fF
C2798 PAND2X1_836/CTRL POR2X1_293/Y 0.00fF
C2799 PAND2X1_469/B POR2X1_42/Y 0.03fF
C2800 VDD POR2X1_757/CTRL 0.00fF
C2801 PAND2X1_365/a_56_28# POR2X1_7/B 0.00fF
C2802 POR2X1_669/CTRL POR2X1_73/Y 0.10fF
C2803 POR2X1_590/A POR2X1_550/B 0.00fF
C2804 POR2X1_220/B POR2X1_551/A 0.03fF
C2805 PAND2X1_824/O VDD 0.00fF
C2806 POR2X1_78/B POR2X1_854/B 0.33fF
C2807 PAND2X1_48/B POR2X1_219/CTRL 0.01fF
C2808 PAND2X1_805/A PAND2X1_539/Y 0.01fF
C2809 PAND2X1_698/CTRL2 PAND2X1_65/B 0.00fF
C2810 PAND2X1_6/Y PAND2X1_599/O 0.17fF
C2811 PAND2X1_738/Y PAND2X1_149/A 0.01fF
C2812 POR2X1_650/A POR2X1_773/B 0.05fF
C2813 POR2X1_42/Y POR2X1_748/CTRL2 0.15fF
C2814 POR2X1_785/A POR2X1_570/B 0.03fF
C2815 PAND2X1_23/Y PAND2X1_69/A 2.82fF
C2816 POR2X1_41/B PAND2X1_186/a_76_28# 0.01fF
C2817 POR2X1_590/CTRL VDD 0.00fF
C2818 POR2X1_466/A POR2X1_181/CTRL 0.33fF
C2819 POR2X1_336/CTRL2 POR2X1_740/Y 0.01fF
C2820 POR2X1_417/Y PAND2X1_357/CTRL2 0.01fF
C2821 PAND2X1_90/A POR2X1_500/Y 0.03fF
C2822 PAND2X1_723/Y POR2X1_7/CTRL 0.01fF
C2823 POR2X1_16/A PAND2X1_787/Y 0.01fF
C2824 POR2X1_362/B POR2X1_260/A 0.03fF
C2825 POR2X1_277/CTRL POR2X1_278/A 0.00fF
C2826 PAND2X1_472/A PAND2X1_401/a_16_344# 0.01fF
C2827 POR2X1_400/CTRL POR2X1_294/A 0.01fF
C2828 PAND2X1_787/Y PAND2X1_175/a_76_28# 0.06fF
C2829 PAND2X1_279/CTRL2 POR2X1_188/Y 0.01fF
C2830 POR2X1_124/O PAND2X1_60/B 0.01fF
C2831 PAND2X1_701/O POR2X1_710/A 0.02fF
C2832 POR2X1_68/A POR2X1_828/A 0.08fF
C2833 PAND2X1_625/O PAND2X1_69/A 0.03fF
C2834 PAND2X1_789/O PAND2X1_793/A 0.01fF
C2835 PAND2X1_56/Y POR2X1_574/a_16_28# 0.13fF
C2836 PAND2X1_23/Y POR2X1_468/Y 0.01fF
C2837 PAND2X1_854/O PAND2X1_535/Y 0.00fF
C2838 PAND2X1_632/B INPUT_0 0.05fF
C2839 PAND2X1_593/Y INPUT_0 0.06fF
C2840 PAND2X1_58/CTRL2 POR2X1_507/A 0.03fF
C2841 POR2X1_52/A POR2X1_283/A 0.10fF
C2842 PAND2X1_724/B POR2X1_387/Y 0.04fF
C2843 INPUT_2 PAND2X1_472/A 0.02fF
C2844 POR2X1_502/A POR2X1_502/CTRL2 0.09fF
C2845 PAND2X1_804/B PAND2X1_175/CTRL 0.04fF
C2846 D_INPUT_3 D_INPUT_2 5.30fF
C2847 POR2X1_20/B POR2X1_386/Y 0.10fF
C2848 POR2X1_578/Y POR2X1_566/B 0.05fF
C2849 POR2X1_8/Y VDD 0.98fF
C2850 POR2X1_750/B POR2X1_188/Y 0.03fF
C2851 PAND2X1_381/Y POR2X1_39/B 0.03fF
C2852 PAND2X1_104/O POR2X1_4/Y 0.09fF
C2853 PAND2X1_48/B POR2X1_274/B 0.03fF
C2854 POR2X1_527/O POR2X1_96/A 0.00fF
C2855 PAND2X1_23/Y POR2X1_325/O 0.01fF
C2856 PAND2X1_641/a_16_344# POR2X1_13/A 0.03fF
C2857 POR2X1_332/B POR2X1_332/CTRL 0.03fF
C2858 POR2X1_84/Y POR2X1_786/Y 0.03fF
C2859 PAND2X1_55/Y POR2X1_796/A 0.07fF
C2860 PAND2X1_6/A PAND2X1_338/B 0.07fF
C2861 PAND2X1_108/CTRL POR2X1_590/A 0.01fF
C2862 PAND2X1_56/Y POR2X1_383/A 0.24fF
C2863 POR2X1_404/Y POR2X1_362/A 0.32fF
C2864 POR2X1_333/A POR2X1_568/B 0.02fF
C2865 POR2X1_96/CTRL POR2X1_7/B 0.01fF
C2866 POR2X1_296/B PAND2X1_56/A 0.03fF
C2867 PAND2X1_686/CTRL POR2X1_7/B 0.01fF
C2868 PAND2X1_71/CTRL2 POR2X1_244/Y 0.01fF
C2869 POR2X1_532/A POR2X1_140/CTRL 0.01fF
C2870 POR2X1_314/O POR2X1_16/A 0.01fF
C2871 POR2X1_57/A PAND2X1_724/O 0.03fF
C2872 POR2X1_270/CTRL2 POR2X1_724/A 0.02fF
C2873 PAND2X1_501/O POR2X1_498/Y -0.00fF
C2874 POR2X1_773/B POR2X1_294/B 0.22fF
C2875 POR2X1_333/a_16_28# POR2X1_578/Y 0.03fF
C2876 POR2X1_391/CTRL2 POR2X1_816/A 0.11fF
C2877 PAND2X1_862/Y VDD 0.14fF
C2878 POR2X1_708/CTRL2 POR2X1_294/A 0.01fF
C2879 PAND2X1_23/Y PAND2X1_823/O 0.04fF
C2880 PAND2X1_89/m4_208_n4# POR2X1_785/A 0.12fF
C2881 POR2X1_192/Y POR2X1_566/O 0.01fF
C2882 POR2X1_857/CTRL2 PAND2X1_72/A 0.10fF
C2883 POR2X1_732/a_16_28# PAND2X1_60/B 0.02fF
C2884 POR2X1_177/a_16_28# POR2X1_236/Y 0.02fF
C2885 PAND2X1_728/CTRL2 POR2X1_816/A 0.01fF
C2886 POR2X1_766/Y VDD 0.10fF
C2887 POR2X1_16/A POR2X1_315/CTRL2 0.01fF
C2888 POR2X1_399/Y POR2X1_411/B 0.01fF
C2889 POR2X1_385/Y VDD 2.14fF
C2890 POR2X1_60/A POR2X1_80/CTRL 0.01fF
C2891 POR2X1_333/A POR2X1_161/CTRL2 0.07fF
C2892 PAND2X1_23/Y PAND2X1_824/B 0.07fF
C2893 PAND2X1_6/Y POR2X1_259/O 0.18fF
C2894 POR2X1_748/A POR2X1_77/Y 0.03fF
C2895 PAND2X1_367/CTRL VDD -0.00fF
C2896 PAND2X1_853/B PAND2X1_335/a_16_344# 0.02fF
C2897 POR2X1_45/Y PAND2X1_579/A 0.00fF
C2898 PAND2X1_859/A POR2X1_39/B 0.05fF
C2899 PAND2X1_295/O POR2X1_837/B 0.01fF
C2900 PAND2X1_480/CTRL POR2X1_238/Y 0.01fF
C2901 POR2X1_275/a_56_344# POR2X1_394/A 0.03fF
C2902 POR2X1_407/Y POR2X1_796/A 0.03fF
C2903 PAND2X1_71/CTRL PAND2X1_48/A 0.01fF
C2904 D_INPUT_0 POR2X1_303/B 0.01fF
C2905 POR2X1_41/B PAND2X1_730/A 0.03fF
C2906 PAND2X1_178/O POR2X1_186/B 0.02fF
C2907 POR2X1_652/Y POR2X1_652/A 0.00fF
C2908 POR2X1_510/Y PAND2X1_60/B 0.03fF
C2909 POR2X1_9/Y POR2X1_260/B 0.07fF
C2910 PAND2X1_6/A PAND2X1_341/Y 0.01fF
C2911 POR2X1_796/A POR2X1_783/Y 0.01fF
C2912 POR2X1_62/Y PAND2X1_197/CTRL 0.01fF
C2913 POR2X1_180/B POR2X1_540/O 0.00fF
C2914 POR2X1_130/A PAND2X1_304/CTRL 0.01fF
C2915 PAND2X1_386/a_76_28# D_INPUT_4 0.01fF
C2916 PAND2X1_65/B POR2X1_632/Y 0.03fF
C2917 PAND2X1_96/B POR2X1_456/B 6.19fF
C2918 POR2X1_390/B POR2X1_335/B 0.00fF
C2919 POR2X1_777/B PAND2X1_52/B 0.05fF
C2920 POR2X1_456/B POR2X1_736/CTRL2 0.00fF
C2921 POR2X1_137/Y POR2X1_116/Y 0.00fF
C2922 POR2X1_502/A PAND2X1_665/CTRL 0.01fF
C2923 POR2X1_508/B POR2X1_578/Y 0.03fF
C2924 POR2X1_447/B POR2X1_579/Y 0.03fF
C2925 POR2X1_325/A POR2X1_374/a_16_28# 0.02fF
C2926 POR2X1_732/a_16_28# POR2X1_353/A 0.03fF
C2927 POR2X1_814/A POR2X1_647/CTRL 0.01fF
C2928 POR2X1_383/A PAND2X1_253/CTRL2 0.03fF
C2929 POR2X1_276/Y PAND2X1_60/B 0.37fF
C2930 POR2X1_661/A POR2X1_296/B 0.10fF
C2931 D_GATE_662 POR2X1_192/B 0.10fF
C2932 POR2X1_186/Y POR2X1_568/A 0.06fF
C2933 POR2X1_821/CTRL POR2X1_39/B 0.01fF
C2934 POR2X1_416/B POR2X1_236/Y 7.47fF
C2935 POR2X1_570/B POR2X1_186/B 0.03fF
C2936 PAND2X1_659/Y POR2X1_599/A 0.09fF
C2937 POR2X1_189/O PAND2X1_480/B 0.02fF
C2938 PAND2X1_65/B PAND2X1_52/B 7.67fF
C2939 POR2X1_145/O PAND2X1_797/Y 0.01fF
C2940 POR2X1_845/CTRL POR2X1_673/Y 0.01fF
C2941 POR2X1_809/A PAND2X1_69/A 0.05fF
C2942 PAND2X1_65/B POR2X1_212/B 0.07fF
C2943 POR2X1_96/A POR2X1_39/B 0.20fF
C2944 D_INPUT_1 PAND2X1_48/A 10.86fF
C2945 POR2X1_566/B POR2X1_192/CTRL 0.05fF
C2946 POR2X1_571/Y POR2X1_844/B 0.01fF
C2947 POR2X1_579/B POR2X1_573/A 0.01fF
C2948 POR2X1_503/O POR2X1_283/A 0.01fF
C2949 PAND2X1_860/A POR2X1_40/Y 0.03fF
C2950 POR2X1_257/A POR2X1_253/CTRL 0.01fF
C2951 POR2X1_110/Y POR2X1_90/Y 0.03fF
C2952 PAND2X1_723/CTRL POR2X1_7/Y 0.01fF
C2953 PAND2X1_90/A POR2X1_561/B 0.04fF
C2954 POR2X1_462/CTRL POR2X1_66/A 0.01fF
C2955 POR2X1_814/A POR2X1_210/CTRL 0.04fF
C2956 POR2X1_572/Y POR2X1_500/Y 0.02fF
C2957 POR2X1_48/A POR2X1_412/CTRL2 0.03fF
C2958 POR2X1_327/Y POR2X1_276/A 0.00fF
C2959 POR2X1_692/CTRL2 POR2X1_20/B 0.03fF
C2960 POR2X1_313/Y POR2X1_16/A 0.00fF
C2961 POR2X1_119/Y POR2X1_425/Y 0.02fF
C2962 POR2X1_567/A PAND2X1_504/m4_208_n4# 0.03fF
C2963 PAND2X1_628/CTRL POR2X1_61/Y 0.01fF
C2964 POR2X1_383/A PAND2X1_71/Y 0.03fF
C2965 PAND2X1_661/Y PAND2X1_120/O 0.01fF
C2966 PAND2X1_426/CTRL POR2X1_121/B 0.01fF
C2967 PAND2X1_649/A POR2X1_38/Y 0.01fF
C2968 PAND2X1_6/Y POR2X1_542/a_16_28# 0.02fF
C2969 PAND2X1_238/O PAND2X1_52/B 0.04fF
C2970 POR2X1_673/Y POR2X1_546/a_16_28# 0.01fF
C2971 POR2X1_51/O INPUT_6 0.01fF
C2972 POR2X1_43/B POR2X1_522/CTRL 0.00fF
C2973 PAND2X1_599/O PAND2X1_52/B 0.01fF
C2974 POR2X1_73/CTRL PAND2X1_341/B 0.01fF
C2975 POR2X1_274/A POR2X1_260/B 0.03fF
C2976 POR2X1_741/Y POR2X1_715/CTRL2 0.01fF
C2977 POR2X1_264/Y PAND2X1_72/A 0.02fF
C2978 POR2X1_416/B POR2X1_232/Y 0.01fF
C2979 POR2X1_741/B POR2X1_186/B 0.00fF
C2980 PAND2X1_69/A POR2X1_711/Y 0.07fF
C2981 POR2X1_846/A PAND2X1_90/Y 0.03fF
C2982 POR2X1_817/a_56_344# PAND2X1_340/B 0.00fF
C2983 PAND2X1_488/O POR2X1_814/A 0.03fF
C2984 PAND2X1_691/Y POR2X1_684/Y 0.05fF
C2985 POR2X1_510/Y POR2X1_554/O 0.18fF
C2986 POR2X1_23/Y POR2X1_437/O 0.01fF
C2987 POR2X1_182/O POR2X1_854/B 0.04fF
C2988 POR2X1_65/A POR2X1_329/A 0.07fF
C2989 PAND2X1_404/CTRL POR2X1_20/B 0.05fF
C2990 POR2X1_772/O POR2X1_113/B 0.01fF
C2991 POR2X1_66/B POR2X1_658/CTRL 0.01fF
C2992 PAND2X1_785/A POR2X1_77/Y 0.03fF
C2993 POR2X1_846/A POR2X1_793/O 0.16fF
C2994 POR2X1_14/Y POR2X1_411/B 0.09fF
C2995 POR2X1_76/CTRL2 POR2X1_296/B 0.03fF
C2996 PAND2X1_69/A POR2X1_728/A 0.00fF
C2997 POR2X1_634/A PAND2X1_47/O 0.20fF
C2998 PAND2X1_193/Y POR2X1_597/A 0.00fF
C2999 POR2X1_416/B PAND2X1_344/CTRL 0.01fF
C3000 POR2X1_434/CTRL POR2X1_434/A 0.01fF
C3001 POR2X1_557/A POR2X1_557/a_16_28# 0.03fF
C3002 POR2X1_431/CTRL POR2X1_5/Y 0.26fF
C3003 PAND2X1_76/O POR2X1_20/B 0.04fF
C3004 PAND2X1_603/CTRL2 POR2X1_260/B 0.01fF
C3005 POR2X1_257/A POR2X1_516/Y 0.01fF
C3006 POR2X1_7/A POR2X1_39/B 0.17fF
C3007 POR2X1_83/B POR2X1_415/A 0.02fF
C3008 PAND2X1_865/Y PAND2X1_216/B 0.07fF
C3009 PAND2X1_108/CTRL2 POR2X1_383/A 0.03fF
C3010 POR2X1_811/B POR2X1_435/B 0.00fF
C3011 POR2X1_54/Y POR2X1_104/O 0.01fF
C3012 PAND2X1_18/B PAND2X1_2/CTRL 0.00fF
C3013 POR2X1_83/B PAND2X1_222/A 0.03fF
C3014 POR2X1_848/CTRL2 POR2X1_859/A 0.01fF
C3015 POR2X1_623/Y POR2X1_5/Y 0.03fF
C3016 POR2X1_241/B POR2X1_454/A 0.03fF
C3017 POR2X1_433/Y PAND2X1_242/Y 0.05fF
C3018 POR2X1_814/A POR2X1_596/Y 0.02fF
C3019 PAND2X1_41/O POR2X1_330/Y 0.01fF
C3020 PAND2X1_798/Y PAND2X1_539/Y 0.12fF
C3021 PAND2X1_220/Y POR2X1_150/Y 0.03fF
C3022 PAND2X1_202/CTRL POR2X1_69/Y 0.01fF
C3023 PAND2X1_202/CTRL2 POR2X1_67/Y 0.01fF
C3024 PAND2X1_638/B POR2X1_260/B 0.02fF
C3025 POR2X1_343/Y POR2X1_569/A 0.10fF
C3026 POR2X1_20/B PAND2X1_541/a_16_344# 0.02fF
C3027 POR2X1_23/Y POR2X1_163/Y 0.01fF
C3028 POR2X1_23/Y POR2X1_29/A 2.40fF
C3029 PAND2X1_264/CTRL POR2X1_77/Y 0.01fF
C3030 POR2X1_48/A PAND2X1_381/Y 0.12fF
C3031 POR2X1_705/B PAND2X1_90/Y 0.03fF
C3032 POR2X1_96/Y PAND2X1_358/A 0.07fF
C3033 POR2X1_60/A POR2X1_289/Y 0.01fF
C3034 PAND2X1_628/CTRL POR2X1_35/Y 0.01fF
C3035 POR2X1_567/B PAND2X1_73/Y 0.05fF
C3036 PAND2X1_246/O VDD 0.00fF
C3037 POR2X1_260/A D_INPUT_4 0.10fF
C3038 POR2X1_81/A POR2X1_153/Y 0.30fF
C3039 PAND2X1_59/B PAND2X1_11/Y 1.04fF
C3040 PAND2X1_94/CTRL2 PAND2X1_58/A 0.00fF
C3041 POR2X1_35/B POR2X1_622/A 0.01fF
C3042 POR2X1_43/B PAND2X1_635/Y 0.03fF
C3043 POR2X1_679/CTRL VDD -0.00fF
C3044 POR2X1_441/Y POR2X1_524/Y 0.00fF
C3045 PAND2X1_251/a_76_28# POR2X1_296/B 0.02fF
C3046 POR2X1_351/O PAND2X1_72/A 0.01fF
C3047 POR2X1_397/Y POR2X1_20/B 0.01fF
C3048 PAND2X1_201/O INPUT_0 0.04fF
C3049 POR2X1_519/CTRL2 POR2X1_43/Y 0.00fF
C3050 POR2X1_257/A PAND2X1_738/O 0.07fF
C3051 POR2X1_78/A PAND2X1_595/O 0.07fF
C3052 POR2X1_654/B POR2X1_655/A 0.03fF
C3053 POR2X1_849/A PAND2X1_58/A 0.10fF
C3054 POR2X1_681/O POR2X1_829/A 0.00fF
C3055 PAND2X1_266/O PAND2X1_215/B 0.17fF
C3056 POR2X1_630/CTRL2 POR2X1_750/B 0.17fF
C3057 POR2X1_48/A PAND2X1_554/CTRL 0.00fF
C3058 POR2X1_590/Y PAND2X1_56/A 0.15fF
C3059 POR2X1_422/Y POR2X1_32/A 0.21fF
C3060 PAND2X1_39/B POR2X1_480/A 0.10fF
C3061 POR2X1_814/A POR2X1_730/CTRL 0.06fF
C3062 POR2X1_260/CTRL2 POR2X1_741/Y 0.01fF
C3063 POR2X1_623/B POR2X1_296/B 0.02fF
C3064 POR2X1_66/A POR2X1_200/CTRL2 0.01fF
C3065 POR2X1_604/O POR2X1_236/Y 0.03fF
C3066 POR2X1_814/B POR2X1_606/O 0.02fF
C3067 POR2X1_271/A POR2X1_416/B 0.03fF
C3068 PAND2X1_206/B PAND2X1_101/O 0.01fF
C3069 PAND2X1_658/A PAND2X1_414/CTRL2 0.01fF
C3070 POR2X1_632/O POR2X1_61/Y 0.05fF
C3071 POR2X1_415/A POR2X1_415/CTRL2 0.05fF
C3072 D_INPUT_0 POR2X1_780/CTRL 0.01fF
C3073 PAND2X1_472/B POR2X1_411/B 0.07fF
C3074 PAND2X1_39/B POR2X1_243/Y 0.07fF
C3075 PAND2X1_6/Y POR2X1_814/A 0.26fF
C3076 POR2X1_68/A PAND2X1_52/O 0.01fF
C3077 PAND2X1_818/CTRL2 PAND2X1_340/B 0.01fF
C3078 POR2X1_866/a_16_28# POR2X1_801/B 0.02fF
C3079 POR2X1_60/A POR2X1_603/Y 0.03fF
C3080 POR2X1_846/A POR2X1_789/O 0.18fF
C3081 PAND2X1_458/CTRL POR2X1_387/Y 0.06fF
C3082 POR2X1_37/Y PAND2X1_333/CTRL2 0.01fF
C3083 PAND2X1_326/B PAND2X1_169/CTRL2 0.01fF
C3084 POR2X1_832/Y VDD 0.08fF
C3085 POR2X1_411/B POR2X1_55/Y 0.13fF
C3086 POR2X1_16/A POR2X1_825/Y 0.03fF
C3087 POR2X1_656/CTRL2 POR2X1_362/B 0.00fF
C3088 PAND2X1_601/O PAND2X1_57/B 0.01fF
C3089 POR2X1_109/O VDD 0.00fF
C3090 PAND2X1_79/a_76_28# POR2X1_844/B 0.04fF
C3091 POR2X1_24/CTRL2 POR2X1_14/Y 0.03fF
C3092 POR2X1_83/B PAND2X1_168/Y 0.01fF
C3093 POR2X1_335/A POR2X1_556/A 0.01fF
C3094 POR2X1_366/Y POR2X1_471/A 0.07fF
C3095 PAND2X1_90/A PAND2X1_39/B 0.01fF
C3096 POR2X1_23/Y POR2X1_256/CTRL 0.13fF
C3097 POR2X1_467/Y POR2X1_448/a_16_28# 0.02fF
C3098 POR2X1_707/B POR2X1_750/B 0.02fF
C3099 POR2X1_768/A POR2X1_113/B 0.04fF
C3100 PAND2X1_240/O POR2X1_102/Y 0.03fF
C3101 PAND2X1_55/Y POR2X1_243/B 0.01fF
C3102 POR2X1_841/B POR2X1_284/CTRL 0.00fF
C3103 PAND2X1_450/CTRL POR2X1_257/A 0.01fF
C3104 POR2X1_96/A POR2X1_48/A 0.06fF
C3105 POR2X1_376/B POR2X1_14/Y 0.07fF
C3106 POR2X1_639/O POR2X1_750/B 0.00fF
C3107 POR2X1_251/A PAND2X1_540/O 0.02fF
C3108 POR2X1_841/B PAND2X1_369/CTRL2 0.05fF
C3109 POR2X1_462/B POR2X1_461/Y 0.01fF
C3110 PAND2X1_248/CTRL2 POR2X1_294/B 0.01fF
C3111 POR2X1_76/O POR2X1_741/Y 0.02fF
C3112 POR2X1_141/CTRL PAND2X1_20/A 0.01fF
C3113 POR2X1_805/Y POR2X1_480/A 0.00fF
C3114 POR2X1_376/B PAND2X1_453/A 0.05fF
C3115 POR2X1_78/B PAND2X1_73/Y 0.26fF
C3116 PAND2X1_9/a_76_28# POR2X1_94/A 0.05fF
C3117 POR2X1_734/B POR2X1_784/A 0.01fF
C3118 D_INPUT_0 POR2X1_217/a_16_28# 0.02fF
C3119 POR2X1_41/B POR2X1_263/Y 0.02fF
C3120 POR2X1_833/A PAND2X1_255/O 0.07fF
C3121 PAND2X1_58/A POR2X1_608/CTRL2 0.01fF
C3122 POR2X1_467/Y PAND2X1_65/B 0.03fF
C3123 PAND2X1_679/CTRL POR2X1_750/B 0.01fF
C3124 PAND2X1_718/Y POR2X1_666/A 0.00fF
C3125 PAND2X1_404/Y POR2X1_43/B 0.96fF
C3126 PAND2X1_717/A PAND2X1_112/O 0.02fF
C3127 POR2X1_605/B PAND2X1_90/Y 0.04fF
C3128 PAND2X1_849/B PAND2X1_206/B 0.07fF
C3129 POR2X1_119/CTRL2 POR2X1_37/Y 0.00fF
C3130 POR2X1_23/Y PAND2X1_445/CTRL 0.28fF
C3131 PAND2X1_287/O PAND2X1_771/Y 0.02fF
C3132 POR2X1_632/O POR2X1_35/Y 0.01fF
C3133 POR2X1_102/Y POR2X1_498/CTRL2 0.10fF
C3134 POR2X1_257/A PAND2X1_702/O 0.00fF
C3135 POR2X1_76/O PAND2X1_32/B 0.00fF
C3136 PAND2X1_279/O VDD -0.00fF
C3137 POR2X1_748/A PAND2X1_793/a_16_344# 0.02fF
C3138 PAND2X1_20/A POR2X1_243/Y 0.41fF
C3139 PAND2X1_319/B PAND2X1_211/CTRL 0.01fF
C3140 POR2X1_66/A POR2X1_740/Y 0.06fF
C3141 POR2X1_365/Y POR2X1_97/A 3.76fF
C3142 PAND2X1_58/A PAND2X1_57/B 1.12fF
C3143 POR2X1_324/B PAND2X1_320/O 0.00fF
C3144 POR2X1_193/Y PAND2X1_52/Y 0.03fF
C3145 POR2X1_697/Y POR2X1_427/O 0.01fF
C3146 PAND2X1_733/O PAND2X1_723/Y 0.03fF
C3147 POR2X1_343/Y PAND2X1_72/A 0.05fF
C3148 POR2X1_179/Y POR2X1_411/B 0.01fF
C3149 POR2X1_102/Y POR2X1_411/O 0.18fF
C3150 POR2X1_423/Y POR2X1_256/CTRL2 0.01fF
C3151 POR2X1_164/Y POR2X1_485/Y 0.06fF
C3152 POR2X1_52/A POR2X1_14/Y 3.60fF
C3153 POR2X1_814/B POR2X1_480/A 0.10fF
C3154 PAND2X1_832/O PAND2X1_499/Y 0.05fF
C3155 POR2X1_796/Y POR2X1_644/A 0.02fF
C3156 PAND2X1_558/Y PAND2X1_579/B 0.06fF
C3157 PAND2X1_771/Y PAND2X1_578/A 0.07fF
C3158 POR2X1_68/CTRL POR2X1_402/A 0.01fF
C3159 POR2X1_814/A PAND2X1_310/O 0.01fF
C3160 PAND2X1_831/Y POR2X1_271/CTRL2 0.01fF
C3161 POR2X1_52/A PAND2X1_453/A 0.07fF
C3162 PAND2X1_319/B PAND2X1_212/O 0.06fF
C3163 POR2X1_66/B POR2X1_415/a_16_28# 0.02fF
C3164 POR2X1_668/Y POR2X1_750/B 0.79fF
C3165 PAND2X1_798/B POR2X1_32/A 0.03fF
C3166 PAND2X1_90/A PAND2X1_20/A 0.10fF
C3167 POR2X1_66/B POR2X1_293/Y 0.19fF
C3168 POR2X1_168/A POR2X1_568/A 0.01fF
C3169 PAND2X1_137/Y PAND2X1_140/CTRL 0.04fF
C3170 POR2X1_220/a_16_28# POR2X1_210/Y 0.06fF
C3171 POR2X1_461/B PAND2X1_90/Y 0.05fF
C3172 PAND2X1_23/Y POR2X1_506/B 0.00fF
C3173 POR2X1_624/Y POR2X1_569/A 0.08fF
C3174 PAND2X1_476/O POR2X1_46/Y 0.01fF
C3175 PAND2X1_575/A PAND2X1_573/B 0.28fF
C3176 POR2X1_152/a_16_28# POR2X1_48/A 0.01fF
C3177 POR2X1_814/B POR2X1_243/Y 0.07fF
C3178 POR2X1_13/A POR2X1_250/A 0.67fF
C3179 PAND2X1_459/CTRL2 POR2X1_55/Y 0.00fF
C3180 PAND2X1_807/B PAND2X1_354/CTRL2 0.01fF
C3181 POR2X1_124/CTRL PAND2X1_41/B 0.01fF
C3182 PAND2X1_465/O POR2X1_7/B 0.15fF
C3183 POR2X1_781/O POR2X1_781/A 0.01fF
C3184 POR2X1_856/B POR2X1_535/A 0.01fF
C3185 POR2X1_48/A POR2X1_689/Y 0.00fF
C3186 PAND2X1_37/O PAND2X1_6/A 0.06fF
C3187 PAND2X1_94/A POR2X1_54/Y 0.91fF
C3188 POR2X1_404/CTRL POR2X1_404/Y 0.01fF
C3189 POR2X1_346/B PAND2X1_39/B 0.05fF
C3190 POR2X1_24/CTRL2 POR2X1_55/Y 0.00fF
C3191 POR2X1_717/a_56_344# POR2X1_558/B 0.01fF
C3192 POR2X1_119/Y PAND2X1_717/A 0.03fF
C3193 POR2X1_8/Y PAND2X1_9/Y 0.03fF
C3194 PAND2X1_279/O POR2X1_741/Y 0.01fF
C3195 PAND2X1_651/Y POR2X1_422/Y 0.03fF
C3196 PAND2X1_673/CTRL POR2X1_13/A 0.01fF
C3197 PAND2X1_82/CTRL2 POR2X1_66/A 0.03fF
C3198 PAND2X1_453/a_16_344# POR2X1_72/B 0.02fF
C3199 POR2X1_60/A POR2X1_433/Y 0.03fF
C3200 POR2X1_446/B POR2X1_704/a_16_28# 0.03fF
C3201 POR2X1_119/Y PAND2X1_266/O 0.08fF
C3202 POR2X1_141/Y POR2X1_572/B 0.03fF
C3203 PAND2X1_738/Y POR2X1_236/Y 0.05fF
C3204 POR2X1_196/Y POR2X1_590/A 0.03fF
C3205 POR2X1_137/Y POR2X1_218/Y 1.75fF
C3206 POR2X1_131/CTRL POR2X1_102/Y 0.01fF
C3207 PAND2X1_94/A POR2X1_202/A 0.04fF
C3208 POR2X1_458/Y POR2X1_343/CTRL2 0.01fF
C3209 PAND2X1_180/O PAND2X1_182/A 0.00fF
C3210 POR2X1_198/B PAND2X1_41/B 0.01fF
C3211 POR2X1_611/O POR2X1_293/Y 0.01fF
C3212 POR2X1_660/O POR2X1_840/B 0.00fF
C3213 POR2X1_68/A POR2X1_244/CTRL 0.16fF
C3214 POR2X1_48/A POR2X1_7/A 13.39fF
C3215 POR2X1_13/A POR2X1_372/A 0.93fF
C3216 PAND2X1_787/m4_208_n4# PAND2X1_715/m4_208_n4# 0.13fF
C3217 POR2X1_669/B POR2X1_591/Y 0.03fF
C3218 PAND2X1_90/A POR2X1_814/B 0.03fF
C3219 POR2X1_66/B POR2X1_460/a_16_28# 0.03fF
C3220 POR2X1_516/B VDD 0.04fF
C3221 PAND2X1_248/O POR2X1_101/Y 0.12fF
C3222 PAND2X1_48/B POR2X1_287/B 0.06fF
C3223 POR2X1_832/CTRL POR2X1_722/Y 0.01fF
C3224 POR2X1_480/A POR2X1_513/B 0.07fF
C3225 PAND2X1_48/Y POR2X1_205/Y 2.53fF
C3226 PAND2X1_230/O PAND2X1_32/B 0.01fF
C3227 POR2X1_376/B POR2X1_55/Y 0.16fF
C3228 PAND2X1_48/Y PAND2X1_55/Y 0.02fF
C3229 POR2X1_496/Y POR2X1_387/Y 0.09fF
C3230 POR2X1_855/B D_INPUT_0 0.03fF
C3231 PAND2X1_41/B D_GATE_741 0.01fF
C3232 PAND2X1_279/O PAND2X1_32/B 0.03fF
C3233 POR2X1_315/Y POR2X1_299/Y 0.01fF
C3234 POR2X1_866/O PAND2X1_32/B 0.01fF
C3235 PAND2X1_57/B POR2X1_435/Y 0.46fF
C3236 POR2X1_468/B VDD 0.19fF
C3237 POR2X1_855/B POR2X1_811/A 0.01fF
C3238 PAND2X1_95/B PAND2X1_65/B 0.06fF
C3239 PAND2X1_48/B POR2X1_483/A 0.03fF
C3240 POR2X1_37/Y POR2X1_235/a_16_28# 0.01fF
C3241 PAND2X1_48/B POR2X1_778/CTRL 0.05fF
C3242 POR2X1_832/CTRL2 POR2X1_832/B 0.03fF
C3243 POR2X1_113/Y POR2X1_390/CTRL 0.07fF
C3244 POR2X1_542/B POR2X1_794/B 0.01fF
C3245 PAND2X1_253/CTRL POR2X1_66/A 0.01fF
C3246 POR2X1_13/A PAND2X1_99/CTRL2 0.01fF
C3247 PAND2X1_556/B POR2X1_293/Y 0.02fF
C3248 POR2X1_814/A POR2X1_632/Y 0.07fF
C3249 PAND2X1_546/Y PAND2X1_712/B 0.23fF
C3250 PAND2X1_20/A PAND2X1_397/CTRL2 0.10fF
C3251 POR2X1_13/A POR2X1_290/Y 0.37fF
C3252 POR2X1_617/Y POR2X1_415/A 0.03fF
C3253 POR2X1_130/A POR2X1_664/Y 0.07fF
C3254 POR2X1_78/B PAND2X1_144/CTRL 0.01fF
C3255 POR2X1_60/a_16_28# POR2X1_60/A -0.00fF
C3256 PAND2X1_491/O PAND2X1_41/B 0.07fF
C3257 POR2X1_66/B POR2X1_21/O 0.10fF
C3258 PAND2X1_483/CTRL2 POR2X1_669/B 0.03fF
C3259 PAND2X1_563/B PAND2X1_566/Y 0.14fF
C3260 POR2X1_719/a_16_28# PAND2X1_73/Y 0.02fF
C3261 PAND2X1_691/Y POR2X1_32/A 0.03fF
C3262 POR2X1_193/A POR2X1_220/Y 0.03fF
C3263 POR2X1_220/Y POR2X1_579/Y 0.03fF
C3264 PAND2X1_207/O POR2X1_153/Y 0.04fF
C3265 POR2X1_410/CTRL POR2X1_790/B 0.03fF
C3266 POR2X1_135/CTRL POR2X1_257/A 0.01fF
C3267 PAND2X1_26/A PAND2X1_18/B 0.07fF
C3268 PAND2X1_254/Y POR2X1_293/Y 0.03fF
C3269 PAND2X1_63/Y PAND2X1_262/a_16_344# 0.04fF
C3270 POR2X1_159/CTRL2 PAND2X1_63/B 0.01fF
C3271 D_INPUT_0 PAND2X1_749/CTRL 0.01fF
C3272 POR2X1_57/A POR2X1_323/CTRL2 0.01fF
C3273 POR2X1_96/A PAND2X1_197/Y 0.02fF
C3274 POR2X1_57/A POR2X1_65/A 9.52fF
C3275 PAND2X1_632/B POR2X1_102/Y 0.03fF
C3276 POR2X1_862/A POR2X1_294/A 0.03fF
C3277 POR2X1_814/A PAND2X1_52/B 0.88fF
C3278 PAND2X1_632/a_16_344# POR2X1_496/Y 0.03fF
C3279 POR2X1_750/B POR2X1_510/Y 0.05fF
C3280 POR2X1_566/A POR2X1_775/A 0.03fF
C3281 POR2X1_13/A PAND2X1_658/B 0.72fF
C3282 POR2X1_52/A POR2X1_55/Y 0.08fF
C3283 POR2X1_356/A POR2X1_785/A 0.05fF
C3284 PAND2X1_797/Y POR2X1_257/A 0.03fF
C3285 POR2X1_515/a_16_28# POR2X1_514/Y -0.00fF
C3286 POR2X1_62/Y PAND2X1_28/a_16_344# 0.02fF
C3287 POR2X1_37/Y PAND2X1_358/A 0.07fF
C3288 PAND2X1_90/A POR2X1_327/O 0.01fF
C3289 PAND2X1_93/B PAND2X1_48/A 0.06fF
C3290 POR2X1_66/A POR2X1_774/A 0.06fF
C3291 PAND2X1_28/CTRL2 POR2X1_750/B 0.01fF
C3292 PAND2X1_48/CTRL POR2X1_786/Y 0.06fF
C3293 POR2X1_390/CTRL POR2X1_260/A 0.04fF
C3294 POR2X1_671/a_16_28# D_INPUT_2 0.02fF
C3295 PAND2X1_72/O VDD 0.00fF
C3296 POR2X1_16/A PAND2X1_78/CTRL2 0.01fF
C3297 POR2X1_572/B POR2X1_404/Y 0.03fF
C3298 PAND2X1_267/Y POR2X1_7/Y 0.01fF
C3299 POR2X1_365/Y POR2X1_366/Y 0.01fF
C3300 PAND2X1_392/B PAND2X1_383/CTRL 0.01fF
C3301 POR2X1_627/O POR2X1_93/A 0.02fF
C3302 POR2X1_652/a_16_28# PAND2X1_90/Y 0.09fF
C3303 POR2X1_65/A POR2X1_229/Y 0.03fF
C3304 POR2X1_526/Y PAND2X1_713/B 0.02fF
C3305 POR2X1_200/a_16_28# POR2X1_200/A 0.05fF
C3306 POR2X1_542/B POR2X1_663/a_76_344# 0.02fF
C3307 POR2X1_55/Y POR2X1_152/A 0.01fF
C3308 POR2X1_614/A POR2X1_220/Y 0.13fF
C3309 POR2X1_41/B PAND2X1_6/A 0.53fF
C3310 POR2X1_66/A POR2X1_550/B 0.03fF
C3311 POR2X1_68/B VDD 2.33fF
C3312 PAND2X1_513/O POR2X1_7/A 0.01fF
C3313 PAND2X1_783/O POR2X1_90/Y 0.01fF
C3314 POR2X1_804/A POR2X1_722/Y 0.03fF
C3315 POR2X1_20/B PAND2X1_861/B 0.72fF
C3316 POR2X1_96/A PAND2X1_359/O 0.05fF
C3317 POR2X1_532/A POR2X1_215/CTRL 0.01fF
C3318 PAND2X1_94/A PAND2X1_23/CTRL 0.01fF
C3319 INPUT_1 PAND2X1_73/a_16_344# 0.02fF
C3320 PAND2X1_96/B PAND2X1_57/B 0.15fF
C3321 POR2X1_823/Y POR2X1_236/Y 0.01fF
C3322 POR2X1_262/Y PAND2X1_339/m4_208_n4# 0.07fF
C3323 POR2X1_614/A POR2X1_404/Y 0.07fF
C3324 POR2X1_102/Y PAND2X1_532/a_76_28# 0.01fF
C3325 POR2X1_296/B POR2X1_737/A 0.05fF
C3326 PAND2X1_126/O POR2X1_5/Y 0.01fF
C3327 POR2X1_259/A POR2X1_259/a_16_28# 0.01fF
C3328 PAND2X1_48/B POR2X1_705/CTRL2 0.00fF
C3329 PAND2X1_139/B PAND2X1_130/CTRL2 0.00fF
C3330 PAND2X1_651/Y PAND2X1_465/B 0.02fF
C3331 POR2X1_502/A POR2X1_578/CTRL 0.00fF
C3332 PAND2X1_476/A POR2X1_409/B 0.06fF
C3333 POR2X1_650/A POR2X1_116/Y 0.03fF
C3334 POR2X1_78/A PAND2X1_48/A 0.13fF
C3335 PAND2X1_73/Y POR2X1_294/A 0.34fF
C3336 POR2X1_52/A PAND2X1_186/CTRL 0.01fF
C3337 POR2X1_65/A POR2X1_744/O 0.01fF
C3338 PAND2X1_786/O POR2X1_394/A 0.06fF
C3339 POR2X1_722/Y PAND2X1_306/CTRL2 0.01fF
C3340 POR2X1_706/B INPUT_1 0.02fF
C3341 PAND2X1_309/CTRL POR2X1_335/B 0.05fF
C3342 POR2X1_865/B PAND2X1_372/O 0.01fF
C3343 POR2X1_186/Y POR2X1_444/Y 0.04fF
C3344 POR2X1_706/A PAND2X1_94/A 0.01fF
C3345 PAND2X1_798/B POR2X1_184/Y 0.00fF
C3346 PAND2X1_553/B PAND2X1_702/O 0.03fF
C3347 POR2X1_481/Y PAND2X1_555/CTRL2 0.01fF
C3348 POR2X1_628/a_76_344# PAND2X1_6/A 0.00fF
C3349 PAND2X1_550/Y VDD 0.17fF
C3350 POR2X1_447/B POR2X1_590/A 0.09fF
C3351 POR2X1_236/Y POR2X1_172/CTRL2 0.03fF
C3352 PAND2X1_808/Y PAND2X1_773/CTRL 0.01fF
C3353 PAND2X1_69/A POR2X1_733/A 0.10fF
C3354 POR2X1_72/B POR2X1_394/A 0.56fF
C3355 POR2X1_383/A INPUT_0 0.08fF
C3356 PAND2X1_578/CTRL VDD 0.00fF
C3357 POR2X1_555/A POR2X1_260/A 0.01fF
C3358 POR2X1_334/B PAND2X1_69/A 0.03fF
C3359 POR2X1_346/CTRL2 PAND2X1_23/Y 0.00fF
C3360 POR2X1_332/B POR2X1_222/A 0.05fF
C3361 POR2X1_787/CTRL POR2X1_325/A 0.01fF
C3362 PAND2X1_83/CTRL POR2X1_35/Y 0.01fF
C3363 PAND2X1_562/a_16_344# PAND2X1_566/Y 0.04fF
C3364 PAND2X1_48/B POR2X1_209/A 0.01fF
C3365 POR2X1_477/A POR2X1_540/A 0.03fF
C3366 PAND2X1_94/A PAND2X1_14/O 0.00fF
C3367 PAND2X1_20/A POR2X1_572/Y 0.04fF
C3368 POR2X1_624/Y PAND2X1_72/A 0.19fF
C3369 POR2X1_40/Y PAND2X1_156/A 0.05fF
C3370 POR2X1_532/A POR2X1_740/Y 0.06fF
C3371 PAND2X1_215/O POR2X1_7/Y 0.02fF
C3372 POR2X1_370/Y PAND2X1_368/O 0.01fF
C3373 PAND2X1_21/CTRL POR2X1_260/A 0.01fF
C3374 PAND2X1_461/O D_INPUT_0 0.15fF
C3375 PAND2X1_275/CTRL POR2X1_573/A 0.01fF
C3376 POR2X1_43/B POR2X1_118/O 0.01fF
C3377 VDD POR2X1_172/O 0.00fF
C3378 PAND2X1_94/A PAND2X1_80/O 0.03fF
C3379 PAND2X1_659/Y PAND2X1_200/O 0.03fF
C3380 POR2X1_244/B POR2X1_259/CTRL 0.01fF
C3381 POR2X1_516/Y PAND2X1_865/A 0.05fF
C3382 PAND2X1_65/B POR2X1_216/Y 0.01fF
C3383 POR2X1_675/CTRL POR2X1_188/Y 0.01fF
C3384 POR2X1_765/O POR2X1_73/Y 0.06fF
C3385 POR2X1_104/O POR2X1_4/Y 0.01fF
C3386 PAND2X1_63/Y PAND2X1_316/O 0.01fF
C3387 POR2X1_564/Y POR2X1_714/a_16_28# 0.01fF
C3388 POR2X1_156/B POR2X1_407/A 0.00fF
C3389 PAND2X1_575/A POR2X1_91/Y 4.57fF
C3390 POR2X1_810/CTRL POR2X1_809/Y 0.01fF
C3391 PAND2X1_81/B POR2X1_68/B 0.01fF
C3392 POR2X1_539/A POR2X1_337/O 0.01fF
C3393 POR2X1_186/CTRL VDD -0.00fF
C3394 POR2X1_57/A PAND2X1_190/Y 0.05fF
C3395 POR2X1_124/B PAND2X1_69/A 0.01fF
C3396 PAND2X1_288/A PAND2X1_367/A 0.06fF
C3397 POR2X1_246/a_16_28# POR2X1_90/Y 0.03fF
C3398 PAND2X1_499/Y POR2X1_153/Y 0.03fF
C3399 PAND2X1_566/Y PAND2X1_347/a_16_344# 0.06fF
C3400 POR2X1_416/B POR2X1_626/CTRL 0.01fF
C3401 PAND2X1_495/CTRL POR2X1_786/Y 0.01fF
C3402 POR2X1_7/A PAND2X1_197/Y 0.03fF
C3403 POR2X1_57/A PAND2X1_836/CTRL2 0.03fF
C3404 POR2X1_85/Y POR2X1_263/Y 0.61fF
C3405 POR2X1_590/A POR2X1_510/O 0.17fF
C3406 PAND2X1_756/O POR2X1_394/A 0.01fF
C3407 POR2X1_192/Y POR2X1_192/O 0.01fF
C3408 PAND2X1_62/a_56_28# POR2X1_394/A 0.00fF
C3409 POR2X1_38/Y POR2X1_521/O 0.01fF
C3410 PAND2X1_553/B PAND2X1_114/CTRL 0.06fF
C3411 PAND2X1_390/CTRL POR2X1_283/A 0.00fF
C3412 POR2X1_16/A POR2X1_57/CTRL2 0.19fF
C3413 POR2X1_322/Y PAND2X1_565/CTRL2 0.00fF
C3414 PAND2X1_725/B PAND2X1_725/O 0.00fF
C3415 POR2X1_192/Y POR2X1_703/Y 0.21fF
C3416 POR2X1_68/B PAND2X1_32/B 4.66fF
C3417 PAND2X1_118/CTRL POR2X1_123/A 0.01fF
C3418 POR2X1_81/A PAND2X1_244/a_16_344# 0.04fF
C3419 POR2X1_7/B PAND2X1_336/CTRL 0.01fF
C3420 POR2X1_112/Y POR2X1_573/A 0.03fF
C3421 POR2X1_38/Y PAND2X1_734/O 0.17fF
C3422 POR2X1_596/A POR2X1_605/A 0.04fF
C3423 PAND2X1_660/Y POR2X1_413/A 0.01fF
C3424 PAND2X1_580/O PAND2X1_568/B 0.02fF
C3425 POR2X1_116/Y POR2X1_294/B 0.03fF
C3426 POR2X1_532/A POR2X1_711/CTRL2 0.16fF
C3427 POR2X1_828/CTRL2 POR2X1_260/A 0.01fF
C3428 POR2X1_539/CTRL POR2X1_662/Y 0.01fF
C3429 POR2X1_49/Y PAND2X1_797/Y 0.03fF
C3430 POR2X1_326/A VDD 0.47fF
C3431 POR2X1_7/B PAND2X1_507/CTRL2 0.03fF
C3432 POR2X1_730/Y POR2X1_294/B 0.07fF
C3433 POR2X1_832/A POR2X1_513/Y 0.01fF
C3434 PAND2X1_816/CTRL POR2X1_463/Y 0.02fF
C3435 POR2X1_119/Y PAND2X1_541/a_76_28# 0.01fF
C3436 POR2X1_625/Y POR2X1_129/Y 0.03fF
C3437 POR2X1_579/Y POR2X1_332/CTRL 0.00fF
C3438 INPUT_0 PAND2X1_71/Y 0.03fF
C3439 POR2X1_566/A POR2X1_339/Y 0.05fF
C3440 PAND2X1_631/A PAND2X1_76/Y 0.07fF
C3441 POR2X1_265/Y VDD 0.27fF
C3442 PAND2X1_560/B PAND2X1_364/B 0.07fF
C3443 POR2X1_767/CTRL VDD 0.00fF
C3444 POR2X1_416/B POR2X1_255/CTRL2 0.01fF
C3445 POR2X1_364/A POR2X1_566/B 0.03fF
C3446 PAND2X1_48/B PAND2X1_484/CTRL2 0.00fF
C3447 POR2X1_417/CTRL POR2X1_283/A 0.04fF
C3448 PAND2X1_476/A PAND2X1_721/a_76_28# 0.04fF
C3449 POR2X1_110/Y INPUT_0 0.04fF
C3450 PAND2X1_710/CTRL PAND2X1_711/A 0.01fF
C3451 POR2X1_356/A POR2X1_186/B 0.07fF
C3452 POR2X1_324/Y VDD 0.04fF
C3453 PAND2X1_658/CTRL2 POR2X1_77/Y 0.03fF
C3454 PAND2X1_727/a_16_344# POR2X1_152/A 0.02fF
C3455 PAND2X1_140/A PAND2X1_284/Y 0.01fF
C3456 POR2X1_333/CTRL PAND2X1_32/B 0.10fF
C3457 POR2X1_323/Y POR2X1_394/A 0.03fF
C3458 POR2X1_795/CTRL POR2X1_186/B 0.01fF
C3459 PAND2X1_264/CTRL2 POR2X1_73/Y 0.04fF
C3460 POR2X1_258/O POR2X1_258/Y 0.01fF
C3461 POR2X1_16/A POR2X1_518/Y 0.12fF
C3462 PAND2X1_684/CTRL POR2X1_149/B 0.01fF
C3463 POR2X1_557/A POR2X1_614/A 0.03fF
C3464 PAND2X1_422/CTRL PAND2X1_60/B 0.01fF
C3465 PAND2X1_23/Y POR2X1_54/CTRL2 0.00fF
C3466 POR2X1_81/CTRL POR2X1_494/Y 0.00fF
C3467 PAND2X1_832/O POR2X1_39/B 0.00fF
C3468 POR2X1_9/Y PAND2X1_66/CTRL 0.04fF
C3469 POR2X1_110/Y POR2X1_424/O 0.06fF
C3470 POR2X1_405/CTRL2 PAND2X1_52/B 0.01fF
C3471 POR2X1_814/B POR2X1_716/CTRL 0.01fF
C3472 POR2X1_705/O POR2X1_260/A 0.01fF
C3473 POR2X1_41/B POR2X1_119/Y 0.15fF
C3474 POR2X1_394/A PAND2X1_547/CTRL2 0.01fF
C3475 POR2X1_557/A POR2X1_38/B 0.07fF
C3476 POR2X1_300/O POR2X1_300/Y 0.05fF
C3477 POR2X1_54/Y POR2X1_462/CTRL2 0.03fF
C3478 POR2X1_135/CTRL PAND2X1_553/B 0.01fF
C3479 PAND2X1_59/CTRL POR2X1_260/A 0.01fF
C3480 PAND2X1_584/O PAND2X1_52/B 0.01fF
C3481 POR2X1_673/Y POR2X1_68/B 0.03fF
C3482 POR2X1_447/B POR2X1_857/B 0.03fF
C3483 POR2X1_326/A POR2X1_741/Y 0.03fF
C3484 POR2X1_42/Y POR2X1_397/CTRL2 0.01fF
C3485 PAND2X1_388/Y PAND2X1_114/O 0.08fF
C3486 POR2X1_732/B POR2X1_337/Y 0.15fF
C3487 POR2X1_513/B PAND2X1_304/O 0.05fF
C3488 POR2X1_41/B POR2X1_85/CTRL 0.00fF
C3489 POR2X1_690/O INPUT_0 0.05fF
C3490 POR2X1_193/A POR2X1_554/CTRL 0.00fF
C3491 PAND2X1_57/B POR2X1_342/B 0.03fF
C3492 PAND2X1_350/CTRL PAND2X1_341/Y 0.01fF
C3493 PAND2X1_853/O PAND2X1_659/Y 0.01fF
C3494 PAND2X1_641/O POR2X1_229/Y 0.00fF
C3495 PAND2X1_281/CTRL2 POR2X1_649/B 0.01fF
C3496 POR2X1_554/B POR2X1_76/A 0.03fF
C3497 POR2X1_181/B POR2X1_703/A 0.03fF
C3498 POR2X1_532/A POR2X1_774/A 0.03fF
C3499 PAND2X1_552/a_16_344# PAND2X1_569/Y 0.02fF
C3500 PAND2X1_90/O D_INPUT_1 0.11fF
C3501 POR2X1_327/Y PAND2X1_60/B 0.06fF
C3502 POR2X1_119/Y POR2X1_256/Y 0.03fF
C3503 POR2X1_853/A PAND2X1_165/m4_208_n4# 0.07fF
C3504 PAND2X1_94/A PAND2X1_748/O 0.15fF
C3505 PAND2X1_473/B POR2X1_589/Y 0.01fF
C3506 PAND2X1_607/O POR2X1_606/Y 0.02fF
C3507 PAND2X1_551/A PAND2X1_326/B 0.06fF
C3508 VDD POR2X1_167/Y 0.36fF
C3509 PAND2X1_832/CTRL2 POR2X1_677/Y 0.00fF
C3510 POR2X1_355/B POR2X1_181/Y 0.03fF
C3511 POR2X1_569/A POR2X1_186/B 0.07fF
C3512 POR2X1_85/Y PAND2X1_215/B 0.01fF
C3513 PAND2X1_373/O POR2X1_544/B 0.05fF
C3514 POR2X1_286/B POR2X1_862/A 0.03fF
C3515 PAND2X1_115/O POR2X1_416/B 0.02fF
C3516 POR2X1_416/B POR2X1_329/a_16_28# 0.00fF
C3517 POR2X1_62/Y POR2X1_7/A 0.10fF
C3518 POR2X1_730/Y PAND2X1_533/O 0.05fF
C3519 POR2X1_27/a_16_28# POR2X1_32/A 0.03fF
C3520 POR2X1_283/A PAND2X1_716/B 0.07fF
C3521 POR2X1_121/A PAND2X1_56/A 0.02fF
C3522 POR2X1_467/Y POR2X1_814/A 0.03fF
C3523 POR2X1_446/B POR2X1_446/a_56_344# 0.00fF
C3524 POR2X1_165/CTRL2 PAND2X1_326/B 0.01fF
C3525 PAND2X1_484/CTRL POR2X1_260/A 0.01fF
C3526 POR2X1_785/A PAND2X1_72/A 0.03fF
C3527 PAND2X1_640/CTRL2 POR2X1_77/Y 0.00fF
C3528 POR2X1_456/B POR2X1_180/CTRL2 0.01fF
C3529 POR2X1_644/CTRL2 POR2X1_260/B 0.01fF
C3530 POR2X1_507/a_16_28# POR2X1_507/A 0.11fF
C3531 PAND2X1_6/A POR2X1_77/Y 0.17fF
C3532 POR2X1_327/Y POR2X1_353/A 0.03fF
C3533 POR2X1_48/A PAND2X1_415/O 0.01fF
C3534 PAND2X1_731/CTRL2 POR2X1_77/Y 0.10fF
C3535 POR2X1_85/Y PAND2X1_6/A 0.02fF
C3536 POR2X1_101/A POR2X1_334/Y 0.05fF
C3537 PAND2X1_821/O PAND2X1_52/B 0.03fF
C3538 POR2X1_416/B PAND2X1_547/O 0.03fF
C3539 POR2X1_39/B PAND2X1_509/CTRL2 0.16fF
C3540 POR2X1_745/Y POR2X1_746/Y 0.01fF
C3541 PAND2X1_152/a_76_28# PAND2X1_72/A 0.02fF
C3542 PAND2X1_96/O PAND2X1_55/Y 0.02fF
C3543 PAND2X1_435/Y POR2X1_271/B 0.13fF
C3544 PAND2X1_254/Y PAND2X1_242/Y 0.27fF
C3545 POR2X1_38/Y POR2X1_39/B 0.21fF
C3546 PAND2X1_405/O POR2X1_5/Y 0.03fF
C3547 PAND2X1_273/O POR2X1_717/B 0.02fF
C3548 PAND2X1_630/B VDD 0.01fF
C3549 PAND2X1_863/B PAND2X1_193/Y 0.06fF
C3550 INPUT_3 POR2X1_614/Y 0.02fF
C3551 POR2X1_376/B POR2X1_441/CTRL 0.05fF
C3552 PAND2X1_94/A POR2X1_4/Y 0.10fF
C3553 POR2X1_435/B POR2X1_296/B 0.03fF
C3554 POR2X1_66/Y POR2X1_296/B 0.07fF
C3555 POR2X1_63/Y POR2X1_667/A 0.27fF
C3556 POR2X1_99/A POR2X1_99/CTRL 0.01fF
C3557 POR2X1_285/Y POR2X1_649/a_16_28# 0.03fF
C3558 PAND2X1_263/m4_208_n4# PAND2X1_202/m4_208_n4# 0.04fF
C3559 POR2X1_119/Y PAND2X1_308/Y 0.07fF
C3560 POR2X1_351/Y POR2X1_568/A 0.03fF
C3561 POR2X1_648/A VDD 0.00fF
C3562 PAND2X1_39/B POR2X1_400/CTRL2 0.01fF
C3563 POR2X1_840/B POR2X1_717/B 0.05fF
C3564 POR2X1_866/A POR2X1_646/Y 0.08fF
C3565 POR2X1_490/O POR2X1_40/Y 0.01fF
C3566 PAND2X1_269/a_76_28# POR2X1_236/Y 0.01fF
C3567 POR2X1_66/B POR2X1_473/CTRL 0.05fF
C3568 POR2X1_477/O POR2X1_186/Y 0.25fF
C3569 POR2X1_383/A POR2X1_862/O 0.02fF
C3570 POR2X1_493/CTRL PAND2X1_72/A 0.01fF
C3571 POR2X1_110/Y POR2X1_110/CTRL2 0.01fF
C3572 PAND2X1_127/a_76_28# POR2X1_567/A -0.02fF
C3573 POR2X1_147/a_16_28# POR2X1_532/A 0.02fF
C3574 POR2X1_49/Y PAND2X1_217/CTRL 0.02fF
C3575 POR2X1_609/Y D_INPUT_0 0.03fF
C3576 POR2X1_411/B PAND2X1_793/A 0.03fF
C3577 POR2X1_49/Y POR2X1_628/Y 0.03fF
C3578 POR2X1_263/CTRL2 POR2X1_236/Y 0.16fF
C3579 INPUT_1 POR2X1_39/B 0.47fF
C3580 POR2X1_137/Y POR2X1_138/A 0.00fF
C3581 POR2X1_485/Y PAND2X1_713/B 0.02fF
C3582 POR2X1_77/Y PAND2X1_112/O 0.03fF
C3583 POR2X1_102/Y PAND2X1_590/O 0.03fF
C3584 POR2X1_647/B POR2X1_654/B 0.03fF
C3585 POR2X1_441/Y PAND2X1_544/CTRL 0.01fF
C3586 POR2X1_416/B PAND2X1_155/O 0.02fF
C3587 PAND2X1_449/m4_208_n4# POR2X1_511/Y 0.15fF
C3588 PAND2X1_644/Y POR2X1_60/A 0.03fF
C3589 POR2X1_311/Y POR2X1_48/A 0.03fF
C3590 POR2X1_52/A POR2X1_815/CTRL2 0.01fF
C3591 POR2X1_842/O POR2X1_850/B 0.01fF
C3592 POR2X1_858/O POR2X1_590/A 0.01fF
C3593 POR2X1_454/A PAND2X1_229/CTRL2 0.03fF
C3594 PAND2X1_48/B POR2X1_630/B 0.01fF
C3595 POR2X1_503/m4_208_n4# POR2X1_236/Y 0.07fF
C3596 POR2X1_153/Y POR2X1_39/B 4.31fF
C3597 PAND2X1_207/O PAND2X1_214/A 0.02fF
C3598 POR2X1_384/A POR2X1_39/B 0.05fF
C3599 PAND2X1_404/Y PAND2X1_474/A 0.03fF
C3600 POR2X1_49/Y PAND2X1_267/Y 0.03fF
C3601 POR2X1_416/B PAND2X1_182/B 0.01fF
C3602 PAND2X1_414/O POR2X1_42/Y 0.02fF
C3603 PAND2X1_476/O PAND2X1_571/A 0.03fF
C3604 POR2X1_567/A POR2X1_542/CTRL 0.23fF
C3605 POR2X1_296/Y POR2X1_296/B 0.09fF
C3606 POR2X1_159/CTRL2 POR2X1_32/A 0.01fF
C3607 POR2X1_760/A PAND2X1_197/Y 0.03fF
C3608 PAND2X1_793/Y POR2X1_20/B 0.05fF
C3609 POR2X1_241/a_56_344# POR2X1_241/B 0.00fF
C3610 POR2X1_68/Y VDD 0.15fF
C3611 PAND2X1_826/CTRL VDD 0.00fF
C3612 POR2X1_453/CTRL2 POR2X1_590/A 0.33fF
C3613 PAND2X1_159/O POR2X1_29/A 0.02fF
C3614 PAND2X1_93/B POR2X1_193/Y 0.03fF
C3615 PAND2X1_244/CTRL POR2X1_102/Y 0.01fF
C3616 PAND2X1_404/Y PAND2X1_84/O 0.05fF
C3617 POR2X1_564/Y POR2X1_446/A 0.01fF
C3618 PAND2X1_72/A POR2X1_186/B 2.30fF
C3619 POR2X1_49/CTRL POR2X1_29/A 0.01fF
C3620 POR2X1_669/B POR2X1_72/B 0.12fF
C3621 PAND2X1_594/O POR2X1_186/Y 0.01fF
C3622 POR2X1_119/Y POR2X1_77/Y 0.08fF
C3623 POR2X1_67/Y POR2X1_38/B 0.07fF
C3624 POR2X1_66/B POR2X1_634/A 0.02fF
C3625 POR2X1_20/B PAND2X1_334/CTRL2 0.01fF
C3626 POR2X1_848/A VDD 0.17fF
C3627 PAND2X1_776/Y VDD 0.25fF
C3628 POR2X1_341/A POR2X1_715/a_76_344# 0.01fF
C3629 POR2X1_802/A PAND2X1_72/A 0.01fF
C3630 POR2X1_112/a_76_344# POR2X1_632/Y 0.00fF
C3631 POR2X1_814/A POR2X1_350/B 0.03fF
C3632 POR2X1_864/CTRL POR2X1_750/B 0.01fF
C3633 POR2X1_675/A POR2X1_590/A 0.01fF
C3634 POR2X1_188/A POR2X1_634/A 1.35fF
C3635 PAND2X1_770/O PAND2X1_771/Y 0.02fF
C3636 POR2X1_82/O POR2X1_409/B 0.01fF
C3637 POR2X1_57/A PAND2X1_837/CTRL 0.01fF
C3638 PAND2X1_124/Y PAND2X1_198/m4_208_n4# 0.09fF
C3639 PAND2X1_20/A POR2X1_402/CTRL2 0.10fF
C3640 POR2X1_32/A POR2X1_666/A 0.06fF
C3641 POR2X1_818/Y PAND2X1_751/CTRL2 0.01fF
C3642 POR2X1_443/A POR2X1_545/A 0.07fF
C3643 PAND2X1_214/CTRL2 PAND2X1_35/Y 0.01fF
C3644 POR2X1_445/A POR2X1_563/Y 0.01fF
C3645 POR2X1_692/CTRL2 POR2X1_763/Y 0.05fF
C3646 POR2X1_669/B PAND2X1_756/O 0.00fF
C3647 PAND2X1_655/B POR2X1_600/a_16_28# 0.03fF
C3648 PAND2X1_256/O POR2X1_205/A 0.12fF
C3649 POR2X1_250/Y POR2X1_283/A 0.25fF
C3650 POR2X1_333/A POR2X1_213/B 0.01fF
C3651 POR2X1_625/Y POR2X1_37/Y 0.01fF
C3652 PAND2X1_711/B VDD 0.01fF
C3653 POR2X1_257/A POR2X1_253/Y 0.02fF
C3654 POR2X1_676/CTRL2 POR2X1_828/A 0.01fF
C3655 PAND2X1_116/CTRL POR2X1_40/Y 0.01fF
C3656 POR2X1_278/Y PAND2X1_577/Y 0.03fF
C3657 POR2X1_862/B POR2X1_389/Y 0.03fF
C3658 PAND2X1_9/Y POR2X1_68/B 0.03fF
C3659 PAND2X1_761/O PAND2X1_32/B 0.03fF
C3660 PAND2X1_276/O POR2X1_271/Y 0.02fF
C3661 POR2X1_825/Y POR2X1_397/CTRL 0.00fF
C3662 PAND2X1_766/CTRL PAND2X1_90/Y 0.07fF
C3663 POR2X1_220/Y POR2X1_590/A 0.06fF
C3664 POR2X1_304/Y POR2X1_14/Y 0.00fF
C3665 POR2X1_484/O POR2X1_763/Y 0.05fF
C3666 POR2X1_753/Y POR2X1_754/A 0.00fF
C3667 POR2X1_304/Y PAND2X1_453/A 0.04fF
C3668 PAND2X1_68/CTRL POR2X1_42/Y 0.29fF
C3669 POR2X1_341/A POR2X1_541/a_76_344# 0.01fF
C3670 PAND2X1_48/B PAND2X1_282/CTRL 0.00fF
C3671 POR2X1_66/B POR2X1_130/A 0.69fF
C3672 POR2X1_220/B POR2X1_740/Y 0.03fF
C3673 POR2X1_295/O POR2X1_481/A 0.01fF
C3674 POR2X1_644/CTRL2 POR2X1_407/Y 0.01fF
C3675 POR2X1_634/O INPUT_0 0.02fF
C3676 POR2X1_614/A POR2X1_841/B 5.09fF
C3677 POR2X1_567/B POR2X1_35/Y 0.05fF
C3678 POR2X1_590/A POR2X1_404/Y 0.03fF
C3679 POR2X1_56/CTRL2 POR2X1_55/Y 0.00fF
C3680 POR2X1_330/Y PAND2X1_131/CTRL 0.06fF
C3681 POR2X1_606/O PAND2X1_32/B 0.02fF
C3682 POR2X1_440/Y POR2X1_477/CTRL2 0.01fF
C3683 POR2X1_41/B POR2X1_442/Y 0.02fF
C3684 POR2X1_458/CTRL2 PAND2X1_32/B 0.03fF
C3685 POR2X1_355/B POR2X1_466/Y 0.01fF
C3686 PAND2X1_254/Y POR2X1_60/A 0.01fF
C3687 PAND2X1_847/m4_208_n4# POR2X1_32/A 0.07fF
C3688 POR2X1_660/Y POR2X1_740/Y 0.03fF
C3689 POR2X1_188/A POR2X1_130/A 0.05fF
C3690 POR2X1_102/Y POR2X1_275/CTRL 0.00fF
C3691 PAND2X1_52/B POR2X1_180/Y 0.06fF
C3692 POR2X1_376/B POR2X1_511/Y 0.08fF
C3693 POR2X1_671/CTRL2 POR2X1_5/Y 0.03fF
C3694 POR2X1_423/a_16_28# POR2X1_372/Y 0.05fF
C3695 POR2X1_794/B POR2X1_722/Y 0.03fF
C3696 PAND2X1_217/CTRL2 PAND2X1_267/Y 0.01fF
C3697 PAND2X1_307/CTRL2 POR2X1_56/B 0.01fF
C3698 POR2X1_78/B POR2X1_61/Y 0.02fF
C3699 POR2X1_99/A PAND2X1_57/B 0.03fF
C3700 POR2X1_14/Y POR2X1_233/a_16_28# 0.02fF
C3701 POR2X1_854/CTRL POR2X1_854/B 0.01fF
C3702 POR2X1_490/Y PAND2X1_572/CTRL 0.01fF
C3703 PAND2X1_443/O POR2X1_91/Y 0.02fF
C3704 POR2X1_335/Y POR2X1_270/Y 0.04fF
C3705 POR2X1_734/A POR2X1_546/A 0.27fF
C3706 PAND2X1_23/Y POR2X1_836/A 0.03fF
C3707 POR2X1_775/A POR2X1_241/B 0.03fF
C3708 POR2X1_638/Y POR2X1_66/A 0.01fF
C3709 POR2X1_51/O PAND2X1_635/Y 0.01fF
C3710 PAND2X1_84/Y PAND2X1_558/CTRL 0.01fF
C3711 POR2X1_662/CTRL POR2X1_725/Y 0.08fF
C3712 POR2X1_141/CTRL VDD 0.00fF
C3713 POR2X1_48/A POR2X1_38/Y 0.15fF
C3714 PAND2X1_652/A PAND2X1_361/CTRL2 0.14fF
C3715 POR2X1_657/a_56_344# POR2X1_741/Y 0.00fF
C3716 POR2X1_657/a_16_28# POR2X1_740/Y 0.10fF
C3717 POR2X1_668/Y POR2X1_720/A 0.01fF
C3718 PAND2X1_769/CTRL2 VDD 0.00fF
C3719 PAND2X1_455/CTRL POR2X1_7/B 0.01fF
C3720 POR2X1_83/B PAND2X1_565/CTRL2 0.03fF
C3721 POR2X1_445/a_16_28# POR2X1_750/B 0.08fF
C3722 POR2X1_60/A POR2X1_599/A 0.06fF
C3723 POR2X1_480/A VDD 0.29fF
C3724 POR2X1_245/CTRL POR2X1_37/Y 0.01fF
C3725 POR2X1_558/a_16_28# POR2X1_78/A 0.07fF
C3726 INPUT_1 POR2X1_621/A 0.03fF
C3727 POR2X1_192/Y PAND2X1_90/Y 0.05fF
C3728 POR2X1_800/A POR2X1_783/CTRL 0.00fF
C3729 POR2X1_72/B PAND2X1_174/CTRL 0.01fF
C3730 POR2X1_417/Y PAND2X1_552/B 0.11fF
C3731 POR2X1_143/CTRL2 POR2X1_236/Y 0.32fF
C3732 POR2X1_179/CTRL2 POR2X1_40/Y 0.00fF
C3733 POR2X1_241/B POR2X1_112/Y 0.03fF
C3734 POR2X1_750/B POR2X1_803/A 0.03fF
C3735 PAND2X1_682/CTRL2 POR2X1_750/B 0.01fF
C3736 POR2X1_411/B POR2X1_129/Y 0.14fF
C3737 POR2X1_102/Y POR2X1_90/Y 0.03fF
C3738 INPUT_1 POR2X1_266/CTRL 0.09fF
C3739 PAND2X1_76/Y PAND2X1_775/CTRL 0.04fF
C3740 POR2X1_66/B PAND2X1_638/O 0.01fF
C3741 PAND2X1_3/A PAND2X1_1/CTRL2 0.01fF
C3742 POR2X1_79/A PAND2X1_580/B 0.00fF
C3743 PAND2X1_96/B POR2X1_479/O 0.01fF
C3744 POR2X1_243/Y VDD -0.00fF
C3745 POR2X1_104/O D_INPUT_1 0.02fF
C3746 PAND2X1_771/Y POR2X1_258/Y 0.05fF
C3747 POR2X1_83/B PAND2X1_341/A 0.03fF
C3748 POR2X1_389/A PAND2X1_73/Y 0.03fF
C3749 POR2X1_52/A POR2X1_511/Y 0.03fF
C3750 POR2X1_455/a_16_28# POR2X1_220/Y 0.02fF
C3751 POR2X1_278/Y PAND2X1_659/O 0.06fF
C3752 PAND2X1_717/A PAND2X1_326/B 0.03fF
C3753 POR2X1_267/A POR2X1_68/B 0.02fF
C3754 POR2X1_260/B POR2X1_456/B 0.10fF
C3755 PAND2X1_798/B PAND2X1_579/CTRL 0.01fF
C3756 PAND2X1_468/CTRL2 PAND2X1_580/B 0.00fF
C3757 POR2X1_278/Y POR2X1_498/CTRL2 0.03fF
C3758 PAND2X1_478/CTRL2 PAND2X1_803/A 0.00fF
C3759 PAND2X1_803/Y PAND2X1_212/B 0.44fF
C3760 PAND2X1_48/B POR2X1_663/CTRL 0.09fF
C3761 PAND2X1_23/Y POR2X1_663/CTRL2 0.01fF
C3762 POR2X1_525/a_16_28# POR2X1_52/A 0.07fF
C3763 POR2X1_83/B POR2X1_93/A 1.16fF
C3764 PAND2X1_190/Y PAND2X1_140/a_16_344# 0.06fF
C3765 POR2X1_390/B POR2X1_270/Y 0.03fF
C3766 POR2X1_553/Y VDD 0.09fF
C3767 POR2X1_217/CTRL2 POR2X1_572/B 0.01fF
C3768 PAND2X1_854/a_16_344# PAND2X1_805/A 0.02fF
C3769 PAND2X1_6/Y POR2X1_259/A 0.54fF
C3770 POR2X1_657/CTRL2 POR2X1_510/Y 0.09fF
C3771 POR2X1_634/A PAND2X1_59/O 0.15fF
C3772 PAND2X1_225/O POR2X1_38/B 0.11fF
C3773 POR2X1_124/B POR2X1_640/Y 0.05fF
C3774 PAND2X1_753/O VDD 0.00fF
C3775 PAND2X1_659/Y POR2X1_411/B 0.10fF
C3776 POR2X1_66/B POR2X1_573/A 0.00fF
C3777 POR2X1_96/A PAND2X1_549/O 0.00fF
C3778 POR2X1_13/A POR2X1_669/CTRL2 0.01fF
C3779 POR2X1_596/A POR2X1_678/A 0.02fF
C3780 PAND2X1_61/Y POR2X1_56/Y 0.03fF
C3781 INPUT_1 POR2X1_48/A 0.25fF
C3782 PAND2X1_254/Y PAND2X1_515/CTRL2 0.01fF
C3783 POR2X1_49/Y POR2X1_29/Y 0.09fF
C3784 PAND2X1_90/A VDD 2.17fF
C3785 PAND2X1_42/CTRL D_INPUT_1 0.03fF
C3786 POR2X1_593/B PAND2X1_69/A 0.03fF
C3787 POR2X1_613/Y POR2X1_20/B 0.11fF
C3788 POR2X1_41/B PAND2X1_486/CTRL2 0.01fF
C3789 POR2X1_626/Y POR2X1_93/A -0.01fF
C3790 POR2X1_312/Y PAND2X1_182/a_16_344# 0.02fF
C3791 POR2X1_780/O POR2X1_532/A 0.01fF
C3792 POR2X1_475/A POR2X1_778/B 0.03fF
C3793 PAND2X1_48/B PAND2X1_372/CTRL2 0.01fF
C3794 POR2X1_625/Y POR2X1_293/Y 0.07fF
C3795 POR2X1_244/B POR2X1_785/A 0.03fF
C3796 POR2X1_83/B PAND2X1_720/CTRL 0.01fF
C3797 POR2X1_102/Y POR2X1_757/a_16_28# 0.03fF
C3798 POR2X1_428/CTRL2 POR2X1_32/A 0.03fF
C3799 POR2X1_83/B PAND2X1_559/CTRL2 0.00fF
C3800 PAND2X1_218/CTRL INPUT_0 0.01fF
C3801 POR2X1_590/A POR2X1_215/A 0.01fF
C3802 PAND2X1_840/B VDD 0.00fF
C3803 PAND2X1_641/Y D_INPUT_0 3.06fF
C3804 D_INPUT_0 POR2X1_571/CTRL2 0.02fF
C3805 POR2X1_78/B POR2X1_35/Y 0.08fF
C3806 INPUT_1 POR2X1_225/CTRL2 0.01fF
C3807 POR2X1_121/B PAND2X1_305/m4_208_n4# 0.08fF
C3808 POR2X1_556/A POR2X1_362/a_16_28# 0.02fF
C3809 POR2X1_75/O PAND2X1_76/Y 0.07fF
C3810 POR2X1_300/CTRL POR2X1_13/A 0.01fF
C3811 POR2X1_48/A POR2X1_153/Y 0.12fF
C3812 POR2X1_823/O POR2X1_236/Y 0.03fF
C3813 POR2X1_557/A POR2X1_590/A 0.01fF
C3814 PAND2X1_422/CTRL POR2X1_750/B 0.00fF
C3815 POR2X1_159/a_16_28# POR2X1_38/Y 0.02fF
C3816 PAND2X1_281/O POR2X1_862/A 0.06fF
C3817 POR2X1_453/a_16_28# PAND2X1_60/B 0.02fF
C3818 PAND2X1_697/CTRL VDD 0.00fF
C3819 POR2X1_605/A PAND2X1_90/Y 0.02fF
C3820 POR2X1_57/A PAND2X1_139/a_16_344# 0.02fF
C3821 POR2X1_383/A PAND2X1_766/CTRL2 0.03fF
C3822 POR2X1_45/Y PAND2X1_735/Y 0.07fF
C3823 POR2X1_445/CTRL2 POR2X1_222/Y 0.01fF
C3824 POR2X1_659/A POR2X1_540/Y 0.05fF
C3825 PAND2X1_95/B INPUT_5 0.00fF
C3826 POR2X1_480/A PAND2X1_32/B 0.07fF
C3827 POR2X1_96/A PAND2X1_652/A 0.03fF
C3828 PAND2X1_23/Y PAND2X1_238/CTRL 0.01fF
C3829 PAND2X1_489/CTRL2 PAND2X1_557/A 0.01fF
C3830 POR2X1_330/Y POR2X1_274/B 0.10fF
C3831 POR2X1_3/A POR2X1_25/CTRL2 0.02fF
C3832 POR2X1_397/Y POR2X1_73/Y 0.07fF
C3833 PAND2X1_40/CTRL PAND2X1_57/B 0.01fF
C3834 PAND2X1_562/B POR2X1_387/Y 0.10fF
C3835 POR2X1_42/O VDD 0.00fF
C3836 PAND2X1_236/CTRL POR2X1_68/B 0.00fF
C3837 POR2X1_666/CTRL POR2X1_394/A 0.03fF
C3838 POR2X1_57/A POR2X1_122/Y 0.01fF
C3839 PAND2X1_810/A PAND2X1_810/CTRL 0.01fF
C3840 PAND2X1_308/CTRL POR2X1_14/Y 0.00fF
C3841 POR2X1_60/CTRL2 POR2X1_13/A 0.01fF
C3842 PAND2X1_473/CTRL VDD 0.00fF
C3843 POR2X1_78/B POR2X1_335/B 0.08fF
C3844 PAND2X1_308/CTRL PAND2X1_453/A 0.01fF
C3845 POR2X1_45/Y PAND2X1_493/Y 0.03fF
C3846 POR2X1_124/B POR2X1_121/Y 0.00fF
C3847 POR2X1_466/A POR2X1_337/Y 0.10fF
C3848 PAND2X1_820/CTRL2 POR2X1_847/B 0.03fF
C3849 PAND2X1_621/O POR2X1_750/B 0.06fF
C3850 POR2X1_447/B POR2X1_66/A 0.12fF
C3851 PAND2X1_90/A PAND2X1_81/B 0.04fF
C3852 GATE_479 PAND2X1_467/Y 0.03fF
C3853 POR2X1_68/A POR2X1_294/B 0.17fF
C3854 POR2X1_713/A POR2X1_383/A 0.05fF
C3855 PAND2X1_215/B POR2X1_52/Y 0.02fF
C3856 POR2X1_393/Y POR2X1_394/A 0.03fF
C3857 POR2X1_60/A PAND2X1_358/A 0.07fF
C3858 POR2X1_733/A POR2X1_723/B 0.10fF
C3859 PAND2X1_715/CTRL POR2X1_387/Y 0.05fF
C3860 POR2X1_335/CTRL2 POR2X1_337/A 0.01fF
C3861 POR2X1_788/Y PAND2X1_144/O 0.00fF
C3862 VDD PAND2X1_305/O 0.00fF
C3863 POR2X1_155/CTRL POR2X1_162/Y 0.03fF
C3864 POR2X1_700/CTRL2 POR2X1_700/Y 0.00fF
C3865 POR2X1_271/Y POR2X1_129/Y 0.21fF
C3866 POR2X1_60/A PAND2X1_337/a_56_28# 0.00fF
C3867 POR2X1_483/CTRL POR2X1_228/Y 0.04fF
C3868 PAND2X1_460/CTRL POR2X1_7/B 0.01fF
C3869 POR2X1_593/CTRL2 POR2X1_750/B 0.01fF
C3870 PAND2X1_90/A PAND2X1_32/B 7.83fF
C3871 POR2X1_13/A POR2X1_387/Y 0.16fF
C3872 PAND2X1_48/B POR2X1_541/CTRL2 0.03fF
C3873 PAND2X1_530/CTRL PAND2X1_69/A 0.01fF
C3874 POR2X1_16/A PAND2X1_803/A -0.00fF
C3875 POR2X1_110/Y POR2X1_102/Y 0.16fF
C3876 PAND2X1_116/m4_208_n4# POR2X1_283/A 0.15fF
C3877 POR2X1_327/Y POR2X1_750/B 0.31fF
C3878 POR2X1_614/A POR2X1_114/B 0.03fF
C3879 POR2X1_855/A POR2X1_260/A 0.01fF
C3880 POR2X1_38/Y PAND2X1_197/Y 0.10fF
C3881 POR2X1_325/a_16_28# POR2X1_325/A 0.03fF
C3882 PAND2X1_726/B PAND2X1_713/B 0.03fF
C3883 PAND2X1_17/O INPUT_6 0.03fF
C3884 PAND2X1_738/Y PAND2X1_336/CTRL2 0.14fF
C3885 PAND2X1_23/Y PAND2X1_505/O 0.00fF
C3886 POR2X1_346/B VDD 0.10fF
C3887 PAND2X1_498/a_76_28# POR2X1_840/B 0.03fF
C3888 POR2X1_97/A POR2X1_169/A 5.90fF
C3889 PAND2X1_494/O PAND2X1_32/B 0.03fF
C3890 POR2X1_516/A PAND2X1_254/Y 0.01fF
C3891 POR2X1_376/B POR2X1_129/Y 0.03fF
C3892 POR2X1_193/A POR2X1_222/A 0.03fF
C3893 POR2X1_528/Y POR2X1_56/B 0.67fF
C3894 POR2X1_579/Y POR2X1_222/A 0.03fF
C3895 POR2X1_740/A POR2X1_740/a_16_28# -0.00fF
C3896 D_INPUT_1 POR2X1_576/Y 0.03fF
C3897 POR2X1_549/CTRL POR2X1_266/A 0.01fF
C3898 POR2X1_330/Y POR2X1_512/O 0.02fF
C3899 POR2X1_832/A POR2X1_832/B 0.00fF
C3900 POR2X1_407/A PAND2X1_743/a_76_28# 0.02fF
C3901 POR2X1_60/CTRL PAND2X1_651/Y 0.01fF
C3902 POR2X1_566/A PAND2X1_313/CTRL 0.10fF
C3903 POR2X1_809/A POR2X1_828/Y 0.02fF
C3904 PAND2X1_450/O POR2X1_425/Y 0.02fF
C3905 POR2X1_71/Y PAND2X1_574/CTRL 0.01fF
C3906 POR2X1_78/CTRL PAND2X1_79/Y 0.00fF
C3907 PAND2X1_403/CTRL2 POR2X1_411/B 0.01fF
C3908 POR2X1_786/Y PAND2X1_150/CTRL 0.01fF
C3909 POR2X1_423/Y POR2X1_183/a_16_28# 0.02fF
C3910 POR2X1_335/A PAND2X1_60/B 0.03fF
C3911 PAND2X1_6/Y PAND2X1_88/Y 0.02fF
C3912 PAND2X1_751/O POR2X1_750/Y 0.00fF
C3913 PAND2X1_6/Y POR2X1_84/Y 0.03fF
C3914 POR2X1_5/Y PAND2X1_156/A 0.03fF
C3915 POR2X1_863/A POR2X1_446/B 0.03fF
C3916 POR2X1_61/Y POR2X1_294/A 0.02fF
C3917 POR2X1_68/A PAND2X1_111/B 0.03fF
C3918 POR2X1_345/O POR2X1_244/B 0.01fF
C3919 POR2X1_196/Y POR2X1_532/A 0.05fF
C3920 PAND2X1_319/B PAND2X1_182/O 0.09fF
C3921 PAND2X1_853/B VDD 0.66fF
C3922 POR2X1_754/A POR2X1_754/O 0.02fF
C3923 PAND2X1_480/B PAND2X1_348/A 0.10fF
C3924 PAND2X1_65/B PAND2X1_527/O 0.04fF
C3925 PAND2X1_537/O PAND2X1_364/B 0.06fF
C3926 PAND2X1_464/B POR2X1_329/A 0.03fF
C3927 POR2X1_315/Y PAND2X1_302/O 0.17fF
C3928 POR2X1_81/A POR2X1_72/B 0.03fF
C3929 POR2X1_40/Y POR2X1_524/O 0.01fF
C3930 POR2X1_566/A POR2X1_97/a_16_28# 0.07fF
C3931 POR2X1_244/B POR2X1_186/B 0.03fF
C3932 PAND2X1_803/Y PAND2X1_389/O 0.02fF
C3933 POR2X1_137/Y PAND2X1_96/B 0.04fF
C3934 PAND2X1_90/A POR2X1_673/Y 0.11fF
C3935 PAND2X1_55/Y POR2X1_456/B 0.08fF
C3936 POR2X1_740/Y POR2X1_308/B 0.10fF
C3937 PAND2X1_284/O POR2X1_280/Y 0.02fF
C3938 POR2X1_740/Y POR2X1_787/O 0.28fF
C3939 POR2X1_741/Y POR2X1_787/CTRL 0.00fF
C3940 POR2X1_614/A POR2X1_222/A 0.05fF
C3941 POR2X1_110/CTRL2 INPUT_0 0.09fF
C3942 POR2X1_96/Y POR2X1_376/B 0.00fF
C3943 POR2X1_66/A POR2X1_181/A 0.01fF
C3944 PAND2X1_305/O PAND2X1_32/B 0.05fF
C3945 POR2X1_740/A PAND2X1_23/Y 0.03fF
C3946 POR2X1_137/Y POR2X1_216/CTRL2 0.00fF
C3947 POR2X1_346/B POR2X1_741/Y 0.05fF
C3948 POR2X1_394/A POR2X1_7/B 0.81fF
C3949 POR2X1_52/A POR2X1_129/Y 0.03fF
C3950 POR2X1_814/B PAND2X1_179/O 0.02fF
C3951 POR2X1_545/A POR2X1_551/O 0.01fF
C3952 VDD POR2X1_572/Y 0.12fF
C3953 PAND2X1_850/Y PAND2X1_76/Y 0.12fF
C3954 PAND2X1_7/CTRL POR2X1_259/B 0.08fF
C3955 POR2X1_96/A PAND2X1_779/O 0.00fF
C3956 PAND2X1_535/Y PAND2X1_854/A 0.02fF
C3957 POR2X1_510/Y POR2X1_318/A 0.07fF
C3958 POR2X1_76/B D_INPUT_0 0.13fF
C3959 PAND2X1_79/Y POR2X1_569/A 0.01fF
C3960 POR2X1_628/m4_208_n4# POR2X1_260/A 0.08fF
C3961 POR2X1_562/CTRL POR2X1_186/B 0.00fF
C3962 PAND2X1_94/A D_INPUT_1 1.74fF
C3963 PAND2X1_105/CTRL PAND2X1_348/A 0.08fF
C3964 PAND2X1_572/CTRL2 PAND2X1_723/A 0.00fF
C3965 PAND2X1_472/O PAND2X1_472/A 0.06fF
C3966 POR2X1_72/B PAND2X1_327/O 0.05fF
C3967 POR2X1_237/Y PAND2X1_308/Y 0.02fF
C3968 PAND2X1_631/A PAND2X1_480/B 0.10fF
C3969 POR2X1_52/A PAND2X1_659/Y 0.03fF
C3970 PAND2X1_808/Y PAND2X1_360/Y 0.00fF
C3971 POR2X1_579/B POR2X1_501/CTRL 0.00fF
C3972 PAND2X1_773/B POR2X1_767/Y 0.09fF
C3973 VDD PAND2X1_304/O 0.00fF
C3974 POR2X1_669/B PAND2X1_147/CTRL 0.04fF
C3975 POR2X1_55/Y PAND2X1_716/B 0.03fF
C3976 POR2X1_68/B POR2X1_772/CTRL 0.06fF
C3977 POR2X1_833/A PAND2X1_96/B 0.00fF
C3978 POR2X1_366/CTRL2 POR2X1_383/A 0.03fF
C3979 POR2X1_537/Y PAND2X1_536/CTRL2 0.01fF
C3980 POR2X1_467/Y POR2X1_535/CTRL2 0.01fF
C3981 POR2X1_527/Y PAND2X1_549/B 0.00fF
C3982 POR2X1_249/Y PAND2X1_60/B 0.03fF
C3983 POR2X1_376/B PAND2X1_333/Y 0.21fF
C3984 POR2X1_383/A POR2X1_796/A 0.03fF
C3985 POR2X1_168/O POR2X1_578/Y 0.01fF
C3986 POR2X1_72/CTRL2 POR2X1_71/Y 0.01fF
C3987 POR2X1_41/B PAND2X1_326/B 0.03fF
C3988 PAND2X1_661/m4_208_n4# PAND2X1_659/Y 0.08fF
C3989 POR2X1_334/Y POR2X1_631/B 0.07fF
C3990 POR2X1_35/Y POR2X1_294/A 0.03fF
C3991 POR2X1_485/Y POR2X1_257/A 0.05fF
C3992 POR2X1_447/B POR2X1_222/Y 0.07fF
C3993 PAND2X1_539/Y PAND2X1_854/A 0.02fF
C3994 POR2X1_8/Y POR2X1_384/CTRL2 0.00fF
C3995 POR2X1_567/B PAND2X1_52/CTRL2 0.14fF
C3996 POR2X1_110/Y POR2X1_531/Y 0.01fF
C3997 POR2X1_590/a_16_28# POR2X1_796/A 0.02fF
C3998 POR2X1_264/Y PAND2X1_517/CTRL 0.01fF
C3999 POR2X1_567/A POR2X1_68/A 0.08fF
C4000 PAND2X1_6/Y POR2X1_508/A 0.17fF
C4001 PAND2X1_831/Y POR2X1_271/A 0.38fF
C4002 POR2X1_390/B POR2X1_101/Y 0.03fF
C4003 D_INPUT_5 POR2X1_20/B 0.02fF
C4004 PAND2X1_6/Y POR2X1_359/O 0.08fF
C4005 POR2X1_69/Y D_INPUT_0 0.15fF
C4006 POR2X1_119/Y POR2X1_52/Y 0.05fF
C4007 POR2X1_532/A PAND2X1_692/CTRL2 0.01fF
C4008 POR2X1_249/Y POR2X1_773/O 0.00fF
C4009 POR2X1_7/A POR2X1_6/O 0.01fF
C4010 POR2X1_62/Y POR2X1_38/Y 0.13fF
C4011 POR2X1_704/CTRL POR2X1_317/B 0.01fF
C4012 POR2X1_366/Y POR2X1_169/A 0.28fF
C4013 POR2X1_572/Y PAND2X1_32/B 0.01fF
C4014 POR2X1_303/O POR2X1_513/Y 0.10fF
C4015 PAND2X1_587/Y PAND2X1_52/B 0.01fF
C4016 POR2X1_188/CTRL2 POR2X1_737/A 0.01fF
C4017 POR2X1_486/CTRL POR2X1_590/A 0.01fF
C4018 PAND2X1_856/B PAND2X1_856/CTRL 0.00fF
C4019 POR2X1_416/B POR2X1_232/O 0.16fF
C4020 POR2X1_67/Y POR2X1_590/A 0.03fF
C4021 POR2X1_52/A PAND2X1_333/Y 0.03fF
C4022 PAND2X1_48/B POR2X1_343/Y 0.20fF
C4023 POR2X1_518/CTRL POR2X1_73/Y 0.08fF
C4024 POR2X1_415/A PAND2X1_66/CTRL2 0.00fF
C4025 POR2X1_16/A PAND2X1_722/CTRL2 0.01fF
C4026 POR2X1_382/Y POR2X1_4/Y 0.01fF
C4027 POR2X1_416/B POR2X1_743/Y 0.01fF
C4028 PAND2X1_650/A POR2X1_153/Y 0.03fF
C4029 PAND2X1_655/Y PAND2X1_691/CTRL2 0.01fF
C4030 POR2X1_369/Y PAND2X1_803/Y 0.02fF
C4031 POR2X1_234/A PAND2X1_520/CTRL2 0.01fF
C4032 POR2X1_274/A POR2X1_446/B 0.03fF
C4033 PAND2X1_193/Y PAND2X1_596/O 0.09fF
C4034 POR2X1_98/A PAND2X1_41/B 0.07fF
C4035 PAND2X1_117/O PAND2X1_72/A 0.02fF
C4036 POR2X1_468/B POR2X1_568/A 0.11fF
C4037 POR2X1_808/A POR2X1_648/A 0.02fF
C4038 POR2X1_364/m4_208_n4# POR2X1_365/m4_208_n4# 0.05fF
C4039 PAND2X1_658/A PAND2X1_861/B 0.02fF
C4040 POR2X1_411/B POR2X1_37/Y 0.21fF
C4041 PAND2X1_860/A PAND2X1_347/Y 0.09fF
C4042 POR2X1_51/O POR2X1_36/B 0.05fF
C4043 POR2X1_63/Y D_INPUT_0 0.08fF
C4044 POR2X1_20/B POR2X1_268/CTRL 0.01fF
C4045 PAND2X1_659/Y POR2X1_679/B 0.01fF
C4046 INPUT_1 POR2X1_62/Y 0.06fF
C4047 POR2X1_180/B POR2X1_567/A 0.03fF
C4048 PAND2X1_802/CTRL2 PAND2X1_539/Y 0.01fF
C4049 POR2X1_591/Y POR2X1_39/B 0.05fF
C4050 POR2X1_632/Y PAND2X1_88/Y 0.04fF
C4051 POR2X1_60/A POR2X1_441/Y 0.03fF
C4052 PAND2X1_612/B POR2X1_66/A 0.03fF
C4053 POR2X1_20/B POR2X1_516/Y 0.03fF
C4054 POR2X1_73/Y PAND2X1_861/B 0.01fF
C4055 POR2X1_48/A POR2X1_248/A 0.00fF
C4056 PAND2X1_30/O INPUT_4 0.03fF
C4057 POR2X1_67/Y POR2X1_668/O 0.01fF
C4058 POR2X1_537/O POR2X1_537/Y 0.00fF
C4059 PAND2X1_91/CTRL2 POR2X1_97/A 0.00fF
C4060 POR2X1_316/a_76_344# POR2X1_153/Y 0.03fF
C4061 POR2X1_62/Y POR2X1_153/Y 0.05fF
C4062 POR2X1_827/CTRL VDD -0.00fF
C4063 POR2X1_104/O INPUT_3 0.10fF
C4064 POR2X1_863/A POR2X1_795/B 0.01fF
C4065 POR2X1_150/Y POR2X1_40/Y 1.82fF
C4066 POR2X1_383/Y POR2X1_520/A 0.85fF
C4067 POR2X1_646/B PAND2X1_90/Y 0.05fF
C4068 PAND2X1_659/Y PAND2X1_557/CTRL 0.00fF
C4069 POR2X1_610/CTRL POR2X1_590/A 0.03fF
C4070 PAND2X1_73/O PAND2X1_9/Y 0.02fF
C4071 PAND2X1_85/CTRL2 POR2X1_243/Y 0.03fF
C4072 POR2X1_250/Y POR2X1_488/a_16_28# 0.03fF
C4073 POR2X1_648/Y PAND2X1_511/CTRL2 0.03fF
C4074 POR2X1_841/B POR2X1_590/A 0.18fF
C4075 PAND2X1_65/B POR2X1_227/A 0.02fF
C4076 POR2X1_722/A PAND2X1_696/CTRL2 0.03fF
C4077 PAND2X1_640/B POR2X1_669/B 0.07fF
C4078 POR2X1_48/A POR2X1_819/CTRL 0.01fF
C4079 POR2X1_647/B POR2X1_777/B 0.05fF
C4080 PAND2X1_629/CTRL POR2X1_628/Y 0.00fF
C4081 POR2X1_294/O POR2X1_355/A 0.01fF
C4082 POR2X1_834/Y POR2X1_711/Y 0.10fF
C4083 POR2X1_202/A POR2X1_202/CTRL2 0.05fF
C4084 PAND2X1_571/A PAND2X1_561/Y 0.02fF
C4085 POR2X1_56/CTRL POR2X1_496/Y 0.05fF
C4086 POR2X1_447/A POR2X1_186/Y 0.01fF
C4087 PAND2X1_23/Y PAND2X1_75/CTRL2 0.00fF
C4088 POR2X1_337/Y PAND2X1_179/CTRL2 0.02fF
C4089 POR2X1_8/Y POR2X1_416/B 0.07fF
C4090 POR2X1_14/Y PAND2X1_448/O 0.17fF
C4091 POR2X1_96/A PAND2X1_447/O 0.04fF
C4092 POR2X1_460/Y POR2X1_459/O 0.01fF
C4093 PAND2X1_689/CTRL2 POR2X1_812/A 0.04fF
C4094 POR2X1_66/B PAND2X1_609/m4_208_n4# 0.15fF
C4095 PAND2X1_207/O POR2X1_72/B 0.01fF
C4096 POR2X1_54/Y PAND2X1_62/a_16_344# 0.02fF
C4097 POR2X1_411/B PAND2X1_715/O 0.02fF
C4098 POR2X1_231/A POR2X1_454/A 0.01fF
C4099 POR2X1_629/O POR2X1_186/Y 0.02fF
C4100 POR2X1_555/CTRL POR2X1_186/B 0.08fF
C4101 PAND2X1_217/B POR2X1_23/Y 0.05fF
C4102 POR2X1_335/a_76_344# POR2X1_556/A 0.01fF
C4103 PAND2X1_796/B VDD 0.36fF
C4104 PAND2X1_45/CTRL POR2X1_740/Y 0.45fF
C4105 PAND2X1_33/CTRL2 POR2X1_7/B 0.03fF
C4106 PAND2X1_362/A PAND2X1_807/B 0.01fF
C4107 POR2X1_260/B POR2X1_448/B 0.02fF
C4108 POR2X1_853/A POR2X1_465/CTRL2 0.02fF
C4109 PAND2X1_454/B VDD 0.24fF
C4110 POR2X1_294/Y POR2X1_202/O 0.00fF
C4111 PAND2X1_267/a_76_28# POR2X1_72/B 0.01fF
C4112 POR2X1_760/A PAND2X1_652/A 0.05fF
C4113 POR2X1_84/B VDD 0.00fF
C4114 POR2X1_748/A POR2X1_32/A 0.06fF
C4115 POR2X1_567/A POR2X1_169/A 0.06fF
C4116 POR2X1_66/B POR2X1_241/B 0.03fF
C4117 POR2X1_89/a_16_28# POR2X1_376/B 0.04fF
C4118 PAND2X1_769/Y PAND2X1_769/O 0.00fF
C4119 POR2X1_333/A PAND2X1_20/A 0.45fF
C4120 POR2X1_411/B POR2X1_293/Y 2.04fF
C4121 PAND2X1_340/B INPUT_0 0.08fF
C4122 POR2X1_260/B PAND2X1_131/CTRL2 0.01fF
C4123 POR2X1_462/B POR2X1_462/CTRL2 0.01fF
C4124 PAND2X1_251/CTRL2 VDD 0.00fF
C4125 POR2X1_463/O POR2X1_532/A 0.08fF
C4126 POR2X1_376/B POR2X1_37/Y 0.16fF
C4127 POR2X1_60/A PAND2X1_200/O 0.03fF
C4128 POR2X1_416/B POR2X1_385/Y 0.05fF
C4129 PAND2X1_90/A PAND2X1_9/Y 0.36fF
C4130 PAND2X1_205/CTRL2 PAND2X1_735/Y 0.01fF
C4131 PAND2X1_65/B PAND2X1_65/a_16_344# 0.02fF
C4132 PAND2X1_798/a_16_344# PAND2X1_354/A 0.02fF
C4133 PAND2X1_794/O POR2X1_40/Y 0.05fF
C4134 PAND2X1_39/B POR2X1_828/O 0.35fF
C4135 POR2X1_78/A PAND2X1_42/CTRL 0.02fF
C4136 POR2X1_260/B PAND2X1_57/B 0.62fF
C4137 POR2X1_847/B PAND2X1_381/Y 0.01fF
C4138 POR2X1_311/Y PAND2X1_349/B 0.03fF
C4139 POR2X1_23/Y VDD 3.96fF
C4140 PAND2X1_474/CTRL2 POR2X1_43/B 0.03fF
C4141 POR2X1_270/Y POR2X1_370/Y 0.68fF
C4142 POR2X1_623/CTRL VDD 0.00fF
C4143 PAND2X1_603/CTRL PAND2X1_90/Y 0.03fF
C4144 PAND2X1_48/B POR2X1_624/Y 0.07fF
C4145 INPUT_2 PAND2X1_618/CTRL2 0.00fF
C4146 POR2X1_366/Y PAND2X1_271/CTRL 0.01fF
C4147 PAND2X1_20/A POR2X1_734/A 0.07fF
C4148 POR2X1_322/Y PAND2X1_717/A 0.67fF
C4149 POR2X1_654/m4_208_n4# POR2X1_774/A 0.15fF
C4150 POR2X1_748/A POR2X1_419/Y 0.05fF
C4151 POR2X1_41/B PAND2X1_852/A 0.01fF
C4152 POR2X1_77/Y PAND2X1_326/B 0.03fF
C4153 POR2X1_362/B POR2X1_296/B 5.35fF
C4154 POR2X1_96/A PAND2X1_205/A 0.03fF
C4155 POR2X1_683/Y POR2X1_604/CTRL2 0.00fF
C4156 POR2X1_416/B PAND2X1_346/CTRL 0.01fF
C4157 POR2X1_333/A POR2X1_814/B 0.10fF
C4158 POR2X1_614/A PAND2X1_761/CTRL2 0.03fF
C4159 POR2X1_307/B POR2X1_590/A 2.99fF
C4160 PAND2X1_781/CTRL2 POR2X1_745/Y 0.02fF
C4161 PAND2X1_404/Y POR2X1_494/Y 0.00fF
C4162 PAND2X1_601/O POR2X1_294/B -0.00fF
C4163 POR2X1_329/A POR2X1_283/A 0.10fF
C4164 POR2X1_324/Y POR2X1_568/A 0.01fF
C4165 POR2X1_696/CTRL2 POR2X1_376/B 0.01fF
C4166 POR2X1_792/a_16_28# POR2X1_791/Y 0.09fF
C4167 POR2X1_102/Y PAND2X1_756/CTRL2 0.01fF
C4168 POR2X1_788/A PAND2X1_90/Y 0.02fF
C4169 PAND2X1_6/Y POR2X1_341/A 0.07fF
C4170 POR2X1_220/Y POR2X1_66/A 0.06fF
C4171 INPUT_3 POR2X1_380/O 0.13fF
C4172 POR2X1_88/a_16_28# POR2X1_7/B 0.02fF
C4173 POR2X1_179/a_16_28# POR2X1_411/B 0.03fF
C4174 POR2X1_604/Y POR2X1_236/Y 0.01fF
C4175 POR2X1_260/B POR2X1_285/A 0.01fF
C4176 POR2X1_648/Y POR2X1_796/A 0.03fF
C4177 PAND2X1_39/B POR2X1_786/Y 0.07fF
C4178 POR2X1_796/Y PAND2X1_599/CTRL 0.01fF
C4179 POR2X1_356/A POR2X1_856/B 0.10fF
C4180 PAND2X1_94/CTRL2 PAND2X1_55/Y 0.01fF
C4181 POR2X1_52/A PAND2X1_448/CTRL 0.01fF
C4182 POR2X1_52/A POR2X1_37/Y 0.23fF
C4183 POR2X1_678/A PAND2X1_90/Y -0.02fF
C4184 PAND2X1_463/CTRL POR2X1_5/Y 0.04fF
C4185 POR2X1_66/A POR2X1_404/Y 0.51fF
C4186 POR2X1_668/CTRL POR2X1_750/B 0.11fF
C4187 PAND2X1_220/Y PAND2X1_540/O 0.09fF
C4188 POR2X1_708/CTRL POR2X1_121/B 0.15fF
C4189 POR2X1_568/B PAND2X1_52/B 0.08fF
C4190 POR2X1_814/B POR2X1_734/A 0.07fF
C4191 POR2X1_429/a_76_344# INPUT_7 0.03fF
C4192 POR2X1_322/O POR2X1_23/Y 0.02fF
C4193 POR2X1_102/Y INPUT_0 0.21fF
C4194 PAND2X1_413/a_56_28# PAND2X1_57/B 0.00fF
C4195 POR2X1_471/a_56_344# POR2X1_78/A 0.00fF
C4196 POR2X1_399/O PAND2X1_403/B 0.04fF
C4197 POR2X1_674/CTRL2 PAND2X1_652/A 0.16fF
C4198 PAND2X1_573/CTRL PAND2X1_573/B 0.01fF
C4199 PAND2X1_556/B PAND2X1_556/O 0.00fF
C4200 POR2X1_483/A POR2X1_330/Y 0.03fF
C4201 POR2X1_99/A PAND2X1_85/Y 0.02fF
C4202 POR2X1_188/A POR2X1_733/O 0.01fF
C4203 PAND2X1_206/A PAND2X1_341/A 1.03fF
C4204 POR2X1_72/B PAND2X1_499/Y 0.47fF
C4205 PAND2X1_489/O PAND2X1_798/B 0.06fF
C4206 POR2X1_83/B POR2X1_237/a_16_28# 0.03fF
C4207 POR2X1_411/B POR2X1_408/Y 0.05fF
C4208 POR2X1_669/B POR2X1_7/B 0.20fF
C4209 POR2X1_221/O POR2X1_186/Y 0.01fF
C4210 PAND2X1_217/B PAND2X1_558/O 0.02fF
C4211 POR2X1_863/B PAND2X1_73/Y 0.01fF
C4212 PAND2X1_653/Y PAND2X1_267/Y 1.17fF
C4213 PAND2X1_436/A INPUT_0 0.04fF
C4214 POR2X1_43/B POR2X1_420/O 0.01fF
C4215 PAND2X1_790/O POR2X1_93/A 0.17fF
C4216 PAND2X1_458/O PAND2X1_716/B 0.04fF
C4217 PAND2X1_93/O POR2X1_66/A 0.02fF
C4218 PAND2X1_294/CTRL POR2X1_387/Y 0.07fF
C4219 PAND2X1_39/B PAND2X1_27/CTRL2 0.01fF
C4220 POR2X1_596/A POR2X1_644/CTRL 0.01fF
C4221 POR2X1_859/A POR2X1_750/A 0.03fF
C4222 POR2X1_829/A PAND2X1_200/Y 0.00fF
C4223 POR2X1_312/Y VDD 0.25fF
C4224 POR2X1_65/A POR2X1_236/Y 0.33fF
C4225 PAND2X1_206/B POR2X1_394/A 0.10fF
C4226 D_INPUT_0 PAND2X1_744/O 0.06fF
C4227 PAND2X1_443/Y PAND2X1_724/B 0.04fF
C4228 PAND2X1_243/B POR2X1_14/Y 0.05fF
C4229 POR2X1_764/Y VDD 0.09fF
C4230 PAND2X1_57/O PAND2X1_41/B 0.02fF
C4231 PAND2X1_738/Y PAND2X1_540/CTRL 0.14fF
C4232 PAND2X1_782/CTRL2 POR2X1_747/Y 0.00fF
C4233 POR2X1_102/Y PAND2X1_717/CTRL2 0.01fF
C4234 POR2X1_505/CTRL2 POR2X1_20/B 0.03fF
C4235 PAND2X1_90/A POR2X1_267/A 0.20fF
C4236 PAND2X1_513/CTRL VDD 0.00fF
C4237 PAND2X1_58/A POR2X1_294/B 0.13fF
C4238 POR2X1_44/O VDD 0.00fF
C4239 PAND2X1_429/Y POR2X1_750/B 0.00fF
C4240 POR2X1_683/CTRL POR2X1_72/B 0.01fF
C4241 POR2X1_196/a_76_344# POR2X1_205/Y 0.01fF
C4242 POR2X1_250/O POR2X1_250/A 0.17fF
C4243 POR2X1_40/Y PAND2X1_364/B 0.07fF
C4244 POR2X1_72/O PAND2X1_659/B 0.00fF
C4245 D_INPUT_0 POR2X1_498/A 0.02fF
C4246 POR2X1_114/B POR2X1_590/A 0.04fF
C4247 POR2X1_120/O PAND2X1_90/Y 0.01fF
C4248 POR2X1_797/A POR2X1_797/a_16_28# 0.05fF
C4249 PAND2X1_212/B POR2X1_309/Y 0.01fF
C4250 POR2X1_855/B POR2X1_808/CTRL 0.01fF
C4251 POR2X1_118/Y POR2X1_278/A 0.08fF
C4252 PAND2X1_671/Y VDD 0.13fF
C4253 POR2X1_615/CTRL POR2X1_754/A 0.04fF
C4254 POR2X1_383/A POR2X1_274/A 0.03fF
C4255 POR2X1_110/a_16_28# POR2X1_372/Y 0.06fF
C4256 POR2X1_525/CTRL POR2X1_41/B 0.01fF
C4257 POR2X1_631/a_76_344# POR2X1_294/B 0.00fF
C4258 POR2X1_802/CTRL PAND2X1_93/B 0.10fF
C4259 POR2X1_502/A POR2X1_5/Y 0.03fF
C4260 POR2X1_257/A PAND2X1_726/B 0.07fF
C4261 POR2X1_667/Y POR2X1_73/Y 0.03fF
C4262 POR2X1_96/A PAND2X1_76/Y 0.03fF
C4263 POR2X1_13/A PAND2X1_596/CTRL 0.01fF
C4264 POR2X1_355/O POR2X1_356/A 0.01fF
C4265 PAND2X1_20/A POR2X1_786/Y 0.03fF
C4266 POR2X1_834/Y PAND2X1_601/CTRL 0.25fF
C4267 PAND2X1_12/CTRL POR2X1_260/A 0.00fF
C4268 POR2X1_838/B PAND2X1_96/B 0.00fF
C4269 PAND2X1_20/A POR2X1_775/O 0.01fF
C4270 POR2X1_54/Y PAND2X1_749/CTRL 0.05fF
C4271 POR2X1_590/A POR2X1_458/B 0.13fF
C4272 POR2X1_376/B POR2X1_293/Y 0.10fF
C4273 POR2X1_96/A POR2X1_297/A 0.01fF
C4274 POR2X1_775/A PAND2X1_229/CTRL2 0.01fF
C4275 POR2X1_482/Y PAND2X1_6/A 0.10fF
C4276 PAND2X1_571/A PAND2X1_717/Y 0.03fF
C4277 PAND2X1_625/CTRL2 POR2X1_852/B 0.02fF
C4278 PAND2X1_433/CTRL2 PAND2X1_65/B 0.03fF
C4279 POR2X1_441/Y POR2X1_373/CTRL2 0.01fF
C4280 POR2X1_856/B POR2X1_569/A 0.10fF
C4281 PAND2X1_404/A POR2X1_233/CTRL 0.00fF
C4282 POR2X1_263/Y PAND2X1_63/B 0.18fF
C4283 PAND2X1_651/Y POR2X1_748/A 0.03fF
C4284 POR2X1_717/a_56_344# POR2X1_590/A 0.00fF
C4285 POR2X1_2/a_56_344# INPUT_5 0.01fF
C4286 PAND2X1_483/CTRL2 POR2X1_48/A 0.01fF
C4287 PAND2X1_793/Y PAND2X1_579/B 0.00fF
C4288 POR2X1_297/Y POR2X1_7/B 0.06fF
C4289 POR2X1_423/CTRL2 POR2X1_7/A 0.03fF
C4290 POR2X1_383/A POR2X1_269/A 0.00fF
C4291 POR2X1_66/A POR2X1_773/CTRL 0.00fF
C4292 POR2X1_68/A POR2X1_807/A 1.11fF
C4293 POR2X1_83/B PAND2X1_338/B 0.03fF
C4294 POR2X1_673/Y POR2X1_623/CTRL 0.03fF
C4295 POR2X1_96/A PAND2X1_863/B 0.03fF
C4296 PAND2X1_58/A PAND2X1_111/B 0.01fF
C4297 POR2X1_57/A POR2X1_825/CTRL 0.01fF
C4298 POR2X1_557/A POR2X1_66/A 0.02fF
C4299 POR2X1_494/CTRL2 POR2X1_5/Y 0.02fF
C4300 POR2X1_814/B POR2X1_786/Y 0.03fF
C4301 POR2X1_652/CTRL2 PAND2X1_90/Y 0.14fF
C4302 PAND2X1_444/Y POR2X1_91/Y 0.02fF
C4303 PAND2X1_151/CTRL POR2X1_55/Y 0.01fF
C4304 POR2X1_722/B POR2X1_435/Y 0.10fF
C4305 POR2X1_532/A PAND2X1_766/O 0.01fF
C4306 PAND2X1_824/B POR2X1_630/O 0.04fF
C4307 PAND2X1_563/CTRL VDD 0.00fF
C4308 POR2X1_296/B POR2X1_553/A 0.00fF
C4309 POR2X1_96/A PAND2X1_191/O 0.04fF
C4310 POR2X1_471/CTRL POR2X1_732/B 0.07fF
C4311 PAND2X1_833/O PAND2X1_658/B -0.03fF
C4312 POR2X1_97/A PAND2X1_503/CTRL 0.01fF
C4313 POR2X1_333/A POR2X1_212/O 0.07fF
C4314 POR2X1_376/B PAND2X1_242/a_76_28# 0.02fF
C4315 PAND2X1_95/B PAND2X1_587/Y 0.20fF
C4316 PAND2X1_57/B POR2X1_205/Y 0.03fF
C4317 POR2X1_573/CTRL POR2X1_576/Y 0.01fF
C4318 PAND2X1_56/Y POR2X1_308/a_76_344# 0.03fF
C4319 PAND2X1_57/B PAND2X1_55/Y 0.29fF
C4320 PAND2X1_456/a_76_28# POR2X1_184/Y 0.02fF
C4321 POR2X1_10/m4_208_n4# POR2X1_48/A 0.07fF
C4322 POR2X1_650/A PAND2X1_96/B 0.09fF
C4323 POR2X1_52/A POR2X1_293/Y 0.33fF
C4324 POR2X1_409/O POR2X1_5/Y 0.02fF
C4325 PAND2X1_94/A POR2X1_78/A 0.14fF
C4326 POR2X1_590/A PAND2X1_103/O 0.00fF
C4327 POR2X1_65/A POR2X1_313/a_56_344# 0.00fF
C4328 POR2X1_316/Y POR2X1_271/B 0.03fF
C4329 PAND2X1_551/Y VDD 0.00fF
C4330 PAND2X1_65/B POR2X1_203/Y 0.00fF
C4331 POR2X1_49/Y PAND2X1_560/O 0.17fF
C4332 POR2X1_658/CTRL2 POR2X1_632/Y 0.01fF
C4333 PAND2X1_391/CTRL POR2X1_751/Y 0.01fF
C4334 PAND2X1_852/a_76_28# POR2X1_122/Y 0.02fF
C4335 POR2X1_753/Y POR2X1_753/CTRL2 0.10fF
C4336 POR2X1_121/B PAND2X1_300/a_16_344# 0.01fF
C4337 POR2X1_43/B POR2X1_278/m4_208_n4# 0.04fF
C4338 PAND2X1_57/B POR2X1_363/O 0.01fF
C4339 POR2X1_192/Y D_GATE_222 0.12fF
C4340 PAND2X1_341/B PAND2X1_404/Y 0.03fF
C4341 POR2X1_48/A PAND2X1_703/CTRL2 0.01fF
C4342 POR2X1_686/B PAND2X1_6/Y 0.03fF
C4343 POR2X1_199/O POR2X1_740/Y 0.02fF
C4344 PAND2X1_243/B POR2X1_55/Y 0.09fF
C4345 PAND2X1_793/Y PAND2X1_658/A 3.44fF
C4346 PAND2X1_61/Y PAND2X1_99/Y 0.02fF
C4347 POR2X1_118/Y POR2X1_117/Y 0.00fF
C4348 POR2X1_94/CTRL2 POR2X1_7/B 0.03fF
C4349 PAND2X1_398/CTRL2 POR2X1_293/Y 0.00fF
C4350 PAND2X1_48/B POR2X1_785/A 0.03fF
C4351 POR2X1_502/A POR2X1_775/CTRL2 0.01fF
C4352 POR2X1_515/a_16_28# POR2X1_68/A 0.02fF
C4353 POR2X1_14/Y POR2X1_260/A 0.06fF
C4354 PAND2X1_57/B POR2X1_402/A 0.04fF
C4355 PAND2X1_824/B POR2X1_240/B 0.02fF
C4356 POR2X1_840/B POR2X1_217/O 0.12fF
C4357 PAND2X1_23/Y PAND2X1_816/CTRL 0.10fF
C4358 POR2X1_96/A PAND2X1_566/Y 0.05fF
C4359 POR2X1_41/B PAND2X1_794/B 0.03fF
C4360 POR2X1_536/Y PAND2X1_593/Y 0.00fF
C4361 PAND2X1_90/Y POR2X1_704/CTRL2 0.03fF
C4362 POR2X1_154/O PAND2X1_6/Y 0.00fF
C4363 POR2X1_502/A POR2X1_705/CTRL 0.00fF
C4364 PAND2X1_55/Y POR2X1_285/A 0.03fF
C4365 POR2X1_376/B POR2X1_408/Y 0.09fF
C4366 PAND2X1_849/B POR2X1_40/Y 0.03fF
C4367 POR2X1_315/Y PAND2X1_211/A 0.03fF
C4368 POR2X1_197/a_56_344# POR2X1_196/Y 0.00fF
C4369 PAND2X1_821/CTRL PAND2X1_23/Y 0.02fF
C4370 POR2X1_188/A POR2X1_188/a_16_28# 0.08fF
C4371 POR2X1_167/CTRL PAND2X1_714/A 0.06fF
C4372 POR2X1_341/A POR2X1_632/Y 0.07fF
C4373 POR2X1_401/O POR2X1_68/B 0.01fF
C4374 PAND2X1_859/O POR2X1_283/A 0.01fF
C4375 POR2X1_78/B POR2X1_631/A 0.03fF
C4376 PAND2X1_593/O POR2X1_591/Y 0.02fF
C4377 POR2X1_471/O POR2X1_540/A 0.01fF
C4378 PAND2X1_48/Y POR2X1_383/A 0.03fF
C4379 POR2X1_83/B PAND2X1_337/CTRL2 0.03fF
C4380 PAND2X1_803/A PAND2X1_549/B 0.00fF
C4381 POR2X1_68/A POR2X1_546/B 0.03fF
C4382 POR2X1_408/O POR2X1_587/Y 0.01fF
C4383 PAND2X1_76/Y POR2X1_7/A 0.03fF
C4384 PAND2X1_57/B POR2X1_407/Y 0.07fF
C4385 POR2X1_51/B POR2X1_44/a_56_344# 0.01fF
C4386 POR2X1_376/B PAND2X1_374/CTRL 0.00fF
C4387 PAND2X1_488/CTRL POR2X1_260/A 0.01fF
C4388 POR2X1_750/B POR2X1_737/a_16_28# 0.00fF
C4389 POR2X1_220/Y POR2X1_532/A 0.10fF
C4390 POR2X1_16/A POR2X1_39/CTRL 0.02fF
C4391 PAND2X1_793/Y POR2X1_73/Y 0.03fF
C4392 PAND2X1_216/B POR2X1_423/Y 7.76fF
C4393 POR2X1_43/B PAND2X1_478/CTRL 0.01fF
C4394 PAND2X1_293/CTRL PAND2X1_60/B 0.01fF
C4395 VDD POR2X1_319/Y 0.80fF
C4396 POR2X1_16/A PAND2X1_240/O 0.03fF
C4397 PAND2X1_849/B PAND2X1_849/O 0.00fF
C4398 D_INPUT_3 POR2X1_13/A 0.04fF
C4399 POR2X1_57/A PAND2X1_182/A 0.00fF
C4400 POR2X1_130/A POR2X1_832/A 0.03fF
C4401 PAND2X1_69/A PAND2X1_369/CTRL 0.09fF
C4402 POR2X1_493/B POR2X1_650/A 0.03fF
C4403 POR2X1_254/Y POR2X1_228/Y 0.10fF
C4404 POR2X1_455/a_16_28# POR2X1_222/A 0.01fF
C4405 POR2X1_404/B PAND2X1_60/B 0.01fF
C4406 POR2X1_614/A POR2X1_732/B 0.03fF
C4407 POR2X1_38/Y POR2X1_597/A 0.02fF
C4408 POR2X1_532/A POR2X1_404/Y 0.03fF
C4409 PAND2X1_96/B POR2X1_294/B 0.19fF
C4410 POR2X1_366/Y PAND2X1_96/B 0.07fF
C4411 POR2X1_840/Y D_INPUT_0 0.01fF
C4412 POR2X1_578/Y POR2X1_578/CTRL 0.00fF
C4413 POR2X1_123/B POR2X1_123/CTRL 0.00fF
C4414 POR2X1_68/A POR2X1_407/A 0.12fF
C4415 PAND2X1_642/B PAND2X1_398/O 0.01fF
C4416 POR2X1_590/A POR2X1_362/O 0.01fF
C4417 POR2X1_177/CTRL POR2X1_72/B 0.01fF
C4418 POR2X1_41/B POR2X1_322/Y 0.09fF
C4419 POR2X1_267/A POR2X1_572/Y 0.02fF
C4420 POR2X1_23/CTRL POR2X1_4/Y 0.05fF
C4421 PAND2X1_631/A POR2X1_56/O 0.01fF
C4422 POR2X1_805/A POR2X1_710/O 0.10fF
C4423 PAND2X1_170/O PAND2X1_168/Y 0.01fF
C4424 POR2X1_122/a_16_28# POR2X1_102/Y 0.11fF
C4425 POR2X1_718/a_76_344# POR2X1_834/Y 0.04fF
C4426 POR2X1_596/A PAND2X1_604/O 0.02fF
C4427 POR2X1_800/A PAND2X1_69/A 0.03fF
C4428 POR2X1_578/Y POR2X1_785/m4_208_n4# 0.10fF
C4429 PAND2X1_633/Y VDD -0.00fF
C4430 POR2X1_640/a_16_28# POR2X1_559/A 0.14fF
C4431 POR2X1_360/A POR2X1_101/CTRL2 0.03fF
C4432 PAND2X1_593/Y PAND2X1_730/B 0.03fF
C4433 POR2X1_228/CTRL2 PAND2X1_7/Y 0.01fF
C4434 POR2X1_52/A POR2X1_408/Y 7.08fF
C4435 POR2X1_337/A PAND2X1_57/B 0.03fF
C4436 POR2X1_124/B POR2X1_391/Y 0.08fF
C4437 POR2X1_96/A POR2X1_315/Y 0.09fF
C4438 PAND2X1_242/Y POR2X1_411/B 0.05fF
C4439 PAND2X1_20/A PAND2X1_396/O 0.02fF
C4440 POR2X1_334/Y POR2X1_61/Y 0.07fF
C4441 POR2X1_78/B PAND2X1_232/a_76_28# 0.01fF
C4442 POR2X1_558/A POR2X1_294/B 0.05fF
C4443 POR2X1_16/A POR2X1_85/m4_208_n4# 0.22fF
C4444 PAND2X1_793/Y PAND2X1_244/B 0.03fF
C4445 PAND2X1_649/A POR2X1_393/Y 0.88fF
C4446 INPUT_6 POR2X1_587/O 0.01fF
C4447 POR2X1_96/A PAND2X1_472/CTRL2 0.01fF
C4448 PAND2X1_441/O POR2X1_854/B 0.04fF
C4449 POR2X1_43/Y POR2X1_827/Y 0.02fF
C4450 POR2X1_483/A POR2X1_715/A 0.01fF
C4451 POR2X1_358/CTRL POR2X1_566/B 0.17fF
C4452 D_INPUT_3 POR2X1_63/O 0.04fF
C4453 POR2X1_840/B PAND2X1_72/O 0.14fF
C4454 PAND2X1_866/a_76_28# PAND2X1_805/A 0.01fF
C4455 POR2X1_407/Y POR2X1_828/A 0.01fF
C4456 PAND2X1_472/O PAND2X1_673/Y 0.28fF
C4457 POR2X1_49/Y PAND2X1_338/CTRL2 -0.00fF
C4458 POR2X1_319/CTRL POR2X1_568/Y 0.31fF
C4459 POR2X1_740/Y POR2X1_854/B 0.03fF
C4460 POR2X1_382/Y POR2X1_816/A 0.00fF
C4461 POR2X1_306/CTRL POR2X1_90/Y 0.01fF
C4462 POR2X1_237/Y PAND2X1_241/Y 0.10fF
C4463 PAND2X1_23/Y PAND2X1_757/a_76_28# 0.02fF
C4464 PAND2X1_192/Y POR2X1_385/Y 0.05fF
C4465 POR2X1_856/B PAND2X1_72/A 0.10fF
C4466 POR2X1_66/B PAND2X1_136/O 0.03fF
C4467 POR2X1_435/Y PAND2X1_533/O 0.11fF
C4468 PAND2X1_824/B POR2X1_214/O 0.05fF
C4469 POR2X1_291/CTRL2 POR2X1_42/Y 0.01fF
C4470 POR2X1_198/CTRL POR2X1_215/A 0.02fF
C4471 PAND2X1_653/CTRL2 PAND2X1_557/A 0.01fF
C4472 POR2X1_390/B PAND2X1_23/Y 0.03fF
C4473 POR2X1_467/Y POR2X1_568/B 0.03fF
C4474 POR2X1_493/B POR2X1_294/B 0.06fF
C4475 POR2X1_5/Y POR2X1_171/Y 0.02fF
C4476 PAND2X1_384/CTRL POR2X1_546/A 0.00fF
C4477 POR2X1_614/A POR2X1_729/Y 0.02fF
C4478 POR2X1_703/A PAND2X1_178/O 0.03fF
C4479 POR2X1_266/A VDD 0.01fF
C4480 PAND2X1_6/A PAND2X1_63/B 0.05fF
C4481 POR2X1_693/Y PAND2X1_550/B 0.04fF
C4482 POR2X1_278/Y PAND2X1_360/Y 0.03fF
C4483 POR2X1_16/A POR2X1_591/CTRL2 0.01fF
C4484 POR2X1_834/Y PAND2X1_433/CTRL 0.27fF
C4485 POR2X1_55/Y POR2X1_260/A 0.03fF
C4486 PAND2X1_784/m4_208_n4# POR2X1_7/A 0.12fF
C4487 PAND2X1_737/B POR2X1_57/Y 0.01fF
C4488 PAND2X1_96/B PAND2X1_111/B 0.01fF
C4489 D_INPUT_1 POR2X1_361/a_76_344# 0.01fF
C4490 POR2X1_41/B POR2X1_144/CTRL2 0.13fF
C4491 PAND2X1_291/CTRL PAND2X1_88/Y 0.02fF
C4492 POR2X1_814/A POR2X1_227/A 0.00fF
C4493 D_GATE_222 POR2X1_785/B 0.09fF
C4494 POR2X1_67/Y POR2X1_816/CTRL 0.03fF
C4495 POR2X1_832/Y POR2X1_661/A 0.01fF
C4496 POR2X1_72/B POR2X1_39/B 0.72fF
C4497 POR2X1_416/B POR2X1_609/CTRL2 0.03fF
C4498 INPUT_6 POR2X1_582/A 0.00fF
C4499 PAND2X1_640/B POR2X1_234/A 0.03fF
C4500 PAND2X1_65/B PAND2X1_167/O 0.03fF
C4501 POR2X1_110/Y POR2X1_368/O 0.01fF
C4502 PAND2X1_109/O PAND2X1_41/B 0.11fF
C4503 PAND2X1_90/A POR2X1_558/Y 0.00fF
C4504 PAND2X1_299/m4_208_n4# D_INPUT_0 0.12fF
C4505 PAND2X1_48/B POR2X1_186/B 9.11fF
C4506 POR2X1_57/A POR2X1_283/A 0.06fF
C4507 POR2X1_48/Y POR2X1_153/Y 0.04fF
C4508 VDD POR2X1_691/A -0.00fF
C4509 POR2X1_741/Y POR2X1_507/A 0.10fF
C4510 POR2X1_57/A PAND2X1_121/CTRL 0.01fF
C4511 POR2X1_662/Y POR2X1_741/A 0.01fF
C4512 POR2X1_83/Y POR2X1_13/A 0.02fF
C4513 POR2X1_407/Y POR2X1_707/Y 0.01fF
C4514 POR2X1_481/Y POR2X1_394/A 0.03fF
C4515 POR2X1_505/O PAND2X1_6/A 0.03fF
C4516 POR2X1_651/Y POR2X1_66/A 0.01fF
C4517 POR2X1_635/B PAND2X1_762/m4_208_n4# 0.07fF
C4518 POR2X1_334/Y POR2X1_193/CTRL 0.06fF
C4519 POR2X1_532/A POR2X1_215/A 0.04fF
C4520 POR2X1_780/A POR2X1_796/A 0.01fF
C4521 PAND2X1_496/O PAND2X1_48/A 0.01fF
C4522 POR2X1_3/A POR2X1_158/B 0.05fF
C4523 POR2X1_539/A POR2X1_188/O 0.01fF
C4524 POR2X1_87/O PAND2X1_41/B 0.01fF
C4525 POR2X1_557/A POR2X1_532/A 0.04fF
C4526 PAND2X1_366/a_16_344# POR2X1_42/Y 0.02fF
C4527 POR2X1_68/B POR2X1_773/a_56_344# 0.00fF
C4528 PAND2X1_535/Y PAND2X1_856/B 0.25fF
C4529 POR2X1_407/Y POR2X1_771/A 0.03fF
C4530 PAND2X1_218/a_16_344# PAND2X1_853/B 0.01fF
C4531 POR2X1_216/O POR2X1_101/Y 0.02fF
C4532 PAND2X1_850/Y PAND2X1_480/B 0.10fF
C4533 POR2X1_72/Y POR2X1_119/Y 0.24fF
C4534 PAND2X1_55/Y POR2X1_512/CTRL2 0.00fF
C4535 PAND2X1_42/a_76_28# POR2X1_590/A 0.01fF
C4536 PAND2X1_6/Y PAND2X1_142/CTRL 0.01fF
C4537 PAND2X1_563/a_76_28# POR2X1_394/A 0.02fF
C4538 INPUT_0 POR2X1_761/A 0.06fF
C4539 POR2X1_189/Y PAND2X1_730/A 0.18fF
C4540 PAND2X1_473/B POR2X1_589/a_16_28# 0.07fF
C4541 POR2X1_411/B POR2X1_275/A 0.01fF
C4542 PAND2X1_96/B PAND2X1_533/O 0.03fF
C4543 POR2X1_78/B POR2X1_736/A 0.09fF
C4544 POR2X1_101/Y PAND2X1_63/B 0.03fF
C4545 PAND2X1_283/O POR2X1_294/A 0.26fF
C4546 PAND2X1_106/O POR2X1_276/Y 0.03fF
C4547 POR2X1_85/Y PAND2X1_206/CTRL 0.01fF
C4548 PAND2X1_382/CTRL POR2X1_260/A 0.02fF
C4549 POR2X1_43/B POR2X1_7/Y 0.26fF
C4550 POR2X1_351/B POR2X1_570/B 0.03fF
C4551 POR2X1_20/B POR2X1_628/Y 0.04fF
C4552 POR2X1_266/A PAND2X1_32/B 0.03fF
C4553 POR2X1_709/CTRL INPUT_1 0.01fF
C4554 POR2X1_118/a_16_28# PAND2X1_560/B 0.03fF
C4555 POR2X1_245/CTRL2 PAND2X1_156/A 0.07fF
C4556 POR2X1_369/Y POR2X1_309/Y 0.01fF
C4557 PAND2X1_294/O POR2X1_411/B 0.02fF
C4558 POR2X1_709/B POR2X1_532/A 0.03fF
C4559 POR2X1_78/B POR2X1_500/O 0.02fF
C4560 POR2X1_111/Y POR2X1_283/A 0.04fF
C4561 PAND2X1_771/O PAND2X1_769/Y 0.02fF
C4562 PAND2X1_510/O PAND2X1_510/B 0.00fF
C4563 POR2X1_480/A POR2X1_568/A 0.07fF
C4564 POR2X1_446/B POR2X1_276/B 0.00fF
C4565 POR2X1_244/Y POR2X1_569/A 0.07fF
C4566 PAND2X1_232/CTRL POR2X1_260/A 0.00fF
C4567 POR2X1_84/B PAND2X1_9/Y 0.01fF
C4568 POR2X1_294/B POR2X1_342/B 0.02fF
C4569 POR2X1_257/A PAND2X1_213/CTRL 0.01fF
C4570 PAND2X1_613/CTRL PAND2X1_9/Y 0.01fF
C4571 POR2X1_559/Y POR2X1_560/a_16_28# -0.00fF
C4572 POR2X1_86/CTRL2 PAND2X1_6/A -0.01fF
C4573 POR2X1_394/A PAND2X1_713/A 0.01fF
C4574 PAND2X1_643/Y PAND2X1_729/CTRL 0.13fF
C4575 POR2X1_631/A POR2X1_294/A 0.00fF
C4576 POR2X1_567/A PAND2X1_96/B 0.06fF
C4577 POR2X1_745/Y POR2X1_746/CTRL 0.00fF
C4578 POR2X1_669/B PAND2X1_206/B 0.10fF
C4579 POR2X1_282/a_16_28# POR2X1_102/Y 0.03fF
C4580 POR2X1_368/m4_208_n4# POR2X1_416/B 0.07fF
C4581 PAND2X1_38/O PAND2X1_52/B 0.04fF
C4582 POR2X1_691/A PAND2X1_32/B 0.13fF
C4583 POR2X1_567/A POR2X1_736/CTRL2 0.03fF
C4584 PAND2X1_96/B PAND2X1_323/O 0.09fF
C4585 POR2X1_722/Y PAND2X1_72/A 0.02fF
C4586 PAND2X1_6/Y POR2X1_592/Y 0.01fF
C4587 POR2X1_439/Y POR2X1_440/CTRL2 0.01fF
C4588 PAND2X1_547/CTRL2 POR2X1_39/B 0.00fF
C4589 POR2X1_83/B PAND2X1_717/A 0.01fF
C4590 POR2X1_14/Y POR2X1_329/A 0.09fF
C4591 POR2X1_624/B POR2X1_29/A 0.01fF
C4592 PAND2X1_171/O POR2X1_854/B 0.02fF
C4593 POR2X1_23/Y PAND2X1_9/Y 0.03fF
C4594 POR2X1_499/A D_INPUT_0 0.01fF
C4595 POR2X1_623/CTRL PAND2X1_9/Y 0.01fF
C4596 D_INPUT_3 PAND2X1_610/CTRL2 0.01fF
C4597 POR2X1_174/B POR2X1_835/B 0.01fF
C4598 POR2X1_54/Y POR2X1_77/a_16_28# 0.04fF
C4599 PAND2X1_310/CTRL2 POR2X1_260/A 0.00fF
C4600 POR2X1_326/A POR2X1_737/O 0.05fF
C4601 PAND2X1_568/B PAND2X1_367/O 0.02fF
C4602 PAND2X1_794/B POR2X1_77/Y 0.00fF
C4603 POR2X1_119/Y PAND2X1_349/A 0.03fF
C4604 POR2X1_461/A POR2X1_814/A 0.06fF
C4605 POR2X1_25/Y POR2X1_158/B 0.03fF
C4606 POR2X1_78/B PAND2X1_125/a_56_28# 0.00fF
C4607 PAND2X1_439/O POR2X1_72/B 0.01fF
C4608 PAND2X1_62/O POR2X1_9/Y 0.15fF
C4609 POR2X1_773/B PAND2X1_48/A 0.03fF
C4610 POR2X1_266/A POR2X1_673/Y 0.07fF
C4611 POR2X1_677/Y INPUT_0 0.04fF
C4612 POR2X1_52/A PAND2X1_242/Y 0.01fF
C4613 POR2X1_669/B POR2X1_604/CTRL 0.01fF
C4614 POR2X1_350/B POR2X1_568/B 0.03fF
C4615 PAND2X1_88/Y POR2X1_555/CTRL2 0.01fF
C4616 PAND2X1_480/CTRL2 POR2X1_119/Y 0.00fF
C4617 POR2X1_87/CTRL POR2X1_68/B 0.06fF
C4618 POR2X1_60/A POR2X1_411/B 0.16fF
C4619 POR2X1_9/Y INPUT_0 0.10fF
C4620 POR2X1_307/Y POR2X1_661/A 0.03fF
C4621 POR2X1_816/CTRL2 POR2X1_750/B 0.22fF
C4622 POR2X1_271/Y POR2X1_275/A 0.02fF
C4623 POR2X1_847/A POR2X1_847/a_16_28# 0.09fF
C4624 POR2X1_329/A POR2X1_237/CTRL 0.04fF
C4625 POR2X1_129/Y PAND2X1_716/B 0.03fF
C4626 POR2X1_411/B POR2X1_591/A 0.02fF
C4627 POR2X1_88/O POR2X1_669/B 0.04fF
C4628 PAND2X1_283/m4_208_n4# POR2X1_654/B 0.08fF
C4629 POR2X1_564/B POR2X1_564/CTRL 0.01fF
C4630 PAND2X1_48/B PAND2X1_628/O 0.03fF
C4631 POR2X1_34/a_16_28# POR2X1_34/B 0.02fF
C4632 PAND2X1_508/B PAND2X1_508/O 0.00fF
C4633 POR2X1_9/Y POR2X1_617/O 0.03fF
C4634 PAND2X1_611/CTRL VDD 0.00fF
C4635 POR2X1_68/A PAND2X1_628/CTRL2 0.01fF
C4636 POR2X1_416/B PAND2X1_181/O 0.05fF
C4637 POR2X1_397/Y POR2X1_669/Y 0.03fF
C4638 PAND2X1_659/Y PAND2X1_716/B 0.03fF
C4639 PAND2X1_213/Y POR2X1_167/Y 0.02fF
C4640 POR2X1_63/Y PAND2X1_231/O 0.02fF
C4641 PAND2X1_425/Y PAND2X1_581/Y 0.01fF
C4642 D_INPUT_3 POR2X1_49/a_56_344# 0.03fF
C4643 POR2X1_263/Y POR2X1_32/A 0.02fF
C4644 POR2X1_430/a_16_28# POR2X1_669/B 0.01fF
C4645 PAND2X1_436/CTRL PAND2X1_390/Y 0.01fF
C4646 POR2X1_651/Y POR2X1_532/A 0.03fF
C4647 POR2X1_329/A POR2X1_55/Y 0.03fF
C4648 D_INPUT_5 INPUT_7 0.63fF
C4649 POR2X1_846/Y POR2X1_790/CTRL 0.01fF
C4650 POR2X1_23/Y PAND2X1_208/CTRL2 0.01fF
C4651 POR2X1_379/a_16_28# PAND2X1_52/B 0.08fF
C4652 POR2X1_251/A POR2X1_48/A 1.34fF
C4653 POR2X1_728/CTRL2 POR2X1_452/Y 0.01fF
C4654 PAND2X1_70/CTRL POR2X1_635/A 0.01fF
C4655 POR2X1_48/A POR2X1_72/B 0.35fF
C4656 POR2X1_811/A POR2X1_783/CTRL 0.00fF
C4657 PAND2X1_287/Y PAND2X1_805/A 0.05fF
C4658 POR2X1_244/B POR2X1_776/A 0.01fF
C4659 POR2X1_837/B PAND2X1_505/CTRL 0.01fF
C4660 POR2X1_244/Y PAND2X1_72/A 0.03fF
C4661 POR2X1_67/Y POR2X1_619/a_76_344# 0.00fF
C4662 POR2X1_504/Y POR2X1_626/CTRL2 0.01fF
C4663 POR2X1_227/B POR2X1_776/B 0.03fF
C4664 POR2X1_20/B POR2X1_372/Y 0.03fF
C4665 POR2X1_243/B INPUT_0 0.02fF
C4666 PAND2X1_404/Y POR2X1_497/Y 0.09fF
C4667 POR2X1_56/a_16_28# POR2X1_83/B 0.00fF
C4668 POR2X1_24/CTRL POR2X1_29/A 0.01fF
C4669 PAND2X1_392/O PAND2X1_474/A 0.00fF
C4670 PAND2X1_317/a_76_28# POR2X1_167/Y 0.02fF
C4671 POR2X1_291/CTRL POR2X1_825/Y 0.00fF
C4672 POR2X1_625/CTRL POR2X1_37/Y 0.01fF
C4673 POR2X1_257/A PAND2X1_213/B 0.03fF
C4674 D_INPUT_5 INPUT_4 0.34fF
C4675 POR2X1_373/O POR2X1_77/Y 0.01fF
C4676 PAND2X1_73/Y PAND2X1_278/O 0.10fF
C4677 POR2X1_127/Y PAND2X1_577/Y 0.03fF
C4678 POR2X1_838/B POR2X1_355/A 0.03fF
C4679 POR2X1_78/B POR2X1_270/Y 0.10fF
C4680 PAND2X1_93/B POR2X1_215/CTRL2 0.00fF
C4681 POR2X1_813/O POR2X1_55/Y 0.03fF
C4682 POR2X1_180/a_16_28# POR2X1_181/Y 0.07fF
C4683 POR2X1_22/A POR2X1_20/B 0.03fF
C4684 PAND2X1_717/A PAND2X1_168/CTRL2 0.01fF
C4685 POR2X1_262/Y PAND2X1_716/CTRL 0.02fF
C4686 POR2X1_416/Y POR2X1_20/B 0.03fF
C4687 D_GATE_366 POR2X1_212/A 0.02fF
C4688 POR2X1_32/A PAND2X1_778/CTRL 0.01fF
C4689 POR2X1_856/B POR2X1_244/B 0.03fF
C4690 POR2X1_816/a_76_344# POR2X1_816/A 0.01fF
C4691 POR2X1_43/B POR2X1_257/A 0.10fF
C4692 PAND2X1_88/CTRL PAND2X1_41/B 0.01fF
C4693 POR2X1_67/O POR2X1_55/Y 0.03fF
C4694 POR2X1_376/B POR2X1_60/A 11.23fF
C4695 PAND2X1_862/B POR2X1_37/Y 0.04fF
C4696 POR2X1_263/Y PAND2X1_35/Y 0.04fF
C4697 POR2X1_220/Y POR2X1_220/B 0.01fF
C4698 PAND2X1_215/CTRL PAND2X1_723/Y 0.06fF
C4699 POR2X1_185/CTRL2 POR2X1_260/B 0.01fF
C4700 POR2X1_427/Y POR2X1_40/Y 0.01fF
C4701 PAND2X1_149/CTRL2 POR2X1_669/B 0.01fF
C4702 POR2X1_49/Y PAND2X1_208/O 0.01fF
C4703 POR2X1_182/a_16_28# POR2X1_180/Y -0.00fF
C4704 POR2X1_72/B PAND2X1_513/O 0.05fF
C4705 POR2X1_257/A PAND2X1_785/CTRL 0.05fF
C4706 POR2X1_20/B POR2X1_526/Y 0.05fF
C4707 POR2X1_441/Y POR2X1_142/Y 0.03fF
C4708 PAND2X1_23/Y PAND2X1_827/O 0.03fF
C4709 POR2X1_68/A POR2X1_632/CTRL 0.01fF
C4710 INPUT_3 POR2X1_382/Y 0.03fF
C4711 POR2X1_333/A VDD 9.23fF
C4712 PAND2X1_73/Y POR2X1_76/Y 1.06fF
C4713 PAND2X1_20/A PAND2X1_755/CTRL2 0.00fF
C4714 POR2X1_72/B PAND2X1_199/A 0.06fF
C4715 POR2X1_83/B PAND2X1_435/CTRL 0.02fF
C4716 POR2X1_855/CTRL POR2X1_803/A 0.01fF
C4717 POR2X1_49/CTRL2 POR2X1_236/Y 0.13fF
C4718 PAND2X1_217/B PAND2X1_475/m4_208_n4# 0.07fF
C4719 POR2X1_428/Y POR2X1_700/Y 0.01fF
C4720 POR2X1_817/Y POR2X1_817/CTRL 0.00fF
C4721 POR2X1_416/B PAND2X1_327/CTRL 0.30fF
C4722 POR2X1_29/A PAND2X1_375/CTRL2 0.07fF
C4723 POR2X1_56/CTRL2 POR2X1_293/Y 0.03fF
C4724 POR2X1_686/A POR2X1_448/B 0.02fF
C4725 PAND2X1_404/Y POR2X1_521/a_56_344# 0.00fF
C4726 POR2X1_590/A POR2X1_784/A 0.02fF
C4727 PAND2X1_623/Y POR2X1_754/Y 0.07fF
C4728 POR2X1_72/B PAND2X1_558/a_16_344# 0.05fF
C4729 POR2X1_41/B POR2X1_83/B 10.76fF
C4730 POR2X1_60/A PAND2X1_598/O 0.04fF
C4731 PAND2X1_404/CTRL2 POR2X1_293/Y 0.00fF
C4732 POR2X1_49/CTRL VDD 0.00fF
C4733 POR2X1_409/B POR2X1_599/A 0.01fF
C4734 PAND2X1_423/CTRL POR2X1_480/A 0.03fF
C4735 POR2X1_608/Y POR2X1_294/B 0.05fF
C4736 POR2X1_827/Y POR2X1_73/Y 0.02fF
C4737 POR2X1_383/A POR2X1_276/B 0.00fF
C4738 POR2X1_610/CTRL POR2X1_532/A 0.07fF
C4739 PAND2X1_6/Y POR2X1_678/Y 0.06fF
C4740 POR2X1_454/A POR2X1_341/Y 0.03fF
C4741 POR2X1_51/A POR2X1_748/A 0.03fF
C4742 POR2X1_41/B PAND2X1_215/a_16_344# 0.01fF
C4743 POR2X1_431/CTRL2 POR2X1_129/Y 0.01fF
C4744 POR2X1_52/A POR2X1_60/A 3.18fF
C4745 PAND2X1_206/A PAND2X1_338/B 0.03fF
C4746 POR2X1_734/A VDD 1.47fF
C4747 POR2X1_178/Y POR2X1_150/Y 0.19fF
C4748 PAND2X1_73/Y POR2X1_740/Y 0.05fF
C4749 PAND2X1_287/a_16_344# PAND2X1_577/Y 0.02fF
C4750 PAND2X1_673/CTRL2 POR2X1_236/Y 0.10fF
C4751 PAND2X1_58/A POR2X1_546/B 0.01fF
C4752 POR2X1_420/CTRL2 POR2X1_90/Y 0.01fF
C4753 POR2X1_416/B POR2X1_167/Y 0.03fF
C4754 POR2X1_16/A PAND2X1_201/O 0.00fF
C4755 POR2X1_590/A POR2X1_732/B 0.05fF
C4756 POR2X1_250/A VDD 0.08fF
C4757 POR2X1_66/B POR2X1_465/B 0.03fF
C4758 POR2X1_614/A POR2X1_466/A 0.03fF
C4759 POR2X1_13/A POR2X1_60/Y 0.01fF
C4760 PAND2X1_652/A PAND2X1_794/CTRL2 0.00fF
C4761 PAND2X1_512/a_56_28# INPUT_0 0.00fF
C4762 PAND2X1_651/Y POR2X1_263/Y 0.05fF
C4763 POR2X1_295/CTRL POR2X1_7/B 0.01fF
C4764 PAND2X1_205/A POR2X1_38/Y 0.03fF
C4765 PAND2X1_333/CTRL VDD 0.00fF
C4766 POR2X1_633/Y POR2X1_640/A 0.00fF
C4767 PAND2X1_480/B PAND2X1_579/O 0.02fF
C4768 POR2X1_122/Y POR2X1_236/Y 0.00fF
C4769 PAND2X1_6/A POR2X1_32/A 0.08fF
C4770 POR2X1_257/A PAND2X1_434/CTRL 0.01fF
C4771 POR2X1_54/Y POR2X1_773/CTRL2 0.03fF
C4772 POR2X1_649/B POR2X1_66/A 0.01fF
C4773 PAND2X1_631/CTRL POR2X1_669/B 0.04fF
C4774 PAND2X1_777/O POR2X1_90/Y 0.07fF
C4775 PAND2X1_69/CTRL2 POR2X1_296/B 0.00fF
C4776 POR2X1_403/A POR2X1_403/a_16_28# 0.05fF
C4777 POR2X1_528/Y POR2X1_613/CTRL2 0.05fF
C4778 POR2X1_422/CTRL POR2X1_7/A 0.00fF
C4779 POR2X1_13/A PAND2X1_778/CTRL2 0.00fF
C4780 POR2X1_692/a_56_344# POR2X1_526/Y 0.00fF
C4781 POR2X1_348/CTRL PAND2X1_93/B 0.10fF
C4782 PAND2X1_852/CTRL2 POR2X1_40/Y 0.00fF
C4783 PAND2X1_218/B PAND2X1_656/A 0.19fF
C4784 PAND2X1_599/CTRL POR2X1_330/Y 0.01fF
C4785 PAND2X1_811/CTRL VDD -0.00fF
C4786 POR2X1_304/a_16_28# POR2X1_236/Y 0.05fF
C4787 POR2X1_407/A PAND2X1_58/A 0.03fF
C4788 POR2X1_814/B PAND2X1_372/O 0.04fF
C4789 PAND2X1_816/a_76_28# POR2X1_634/A 0.03fF
C4790 POR2X1_596/A POR2X1_834/CTRL2 0.01fF
C4791 POR2X1_502/A PAND2X1_65/B 0.81fF
C4792 POR2X1_113/Y POR2X1_476/A 0.05fF
C4793 POR2X1_830/O POR2X1_741/Y 0.00fF
C4794 POR2X1_72/B PAND2X1_197/Y 0.03fF
C4795 POR2X1_355/A POR2X1_294/B 0.00fF
C4796 POR2X1_66/B D_GATE_741 0.02fF
C4797 POR2X1_389/CTRL POR2X1_389/Y 0.02fF
C4798 POR2X1_49/Y PAND2X1_624/A 0.01fF
C4799 POR2X1_567/B POR2X1_351/CTRL2 0.06fF
C4800 POR2X1_68/a_16_28# POR2X1_68/B 0.02fF
C4801 POR2X1_446/B POR2X1_456/B 0.03fF
C4802 PAND2X1_803/Y PAND2X1_352/A 0.02fF
C4803 POR2X1_294/Y PAND2X1_60/B 0.39fF
C4804 POR2X1_81/a_16_28# POR2X1_43/B 0.00fF
C4805 PAND2X1_807/a_76_28# PAND2X1_805/Y 0.07fF
C4806 POR2X1_5/Y PAND2X1_364/B 0.03fF
C4807 POR2X1_114/B PAND2X1_279/a_16_344# 0.01fF
C4808 PAND2X1_20/A POR2X1_556/Y 0.03fF
C4809 PAND2X1_224/CTRL2 VDD 0.00fF
C4810 POR2X1_465/B POR2X1_563/CTRL 0.01fF
C4811 POR2X1_590/A POR2X1_206/O 0.17fF
C4812 PAND2X1_65/B PAND2X1_176/O 0.03fF
C4813 POR2X1_516/Y POR2X1_73/Y 0.15fF
C4814 POR2X1_763/Y PAND2X1_738/O 0.08fF
C4815 POR2X1_333/A PAND2X1_32/B 0.05fF
C4816 POR2X1_119/Y POR2X1_411/A 0.07fF
C4817 PAND2X1_650/a_16_344# D_INPUT_0 0.01fF
C4818 PAND2X1_127/O POR2X1_445/A 0.01fF
C4819 POR2X1_278/Y INPUT_0 0.07fF
C4820 D_INPUT_3 POR2X1_29/A 0.14fF
C4821 PAND2X1_94/A POR2X1_84/A 0.09fF
C4822 POR2X1_264/CTRL2 PAND2X1_32/B 0.01fF
C4823 POR2X1_416/B PAND2X1_630/B 0.03fF
C4824 POR2X1_236/Y POR2X1_395/CTRL2 0.01fF
C4825 POR2X1_41/B PAND2X1_140/Y 0.03fF
C4826 PAND2X1_793/Y PAND2X1_804/A 0.03fF
C4827 POR2X1_49/Y POR2X1_43/B 3.37fF
C4828 POR2X1_66/B PAND2X1_491/O 0.04fF
C4829 PAND2X1_90/Y PAND2X1_132/O 0.04fF
C4830 POR2X1_108/O POR2X1_102/Y 0.07fF
C4831 POR2X1_440/Y POR2X1_466/A 0.05fF
C4832 POR2X1_57/A POR2X1_14/Y 0.05fF
C4833 PAND2X1_215/B PAND2X1_741/B 0.03fF
C4834 PAND2X1_653/CTRL POR2X1_329/A 0.02fF
C4835 POR2X1_114/O POR2X1_777/B 0.02fF
C4836 PAND2X1_85/Y PAND2X1_55/Y 0.07fF
C4837 PAND2X1_96/B POR2X1_643/A 0.01fF
C4838 POR2X1_96/A PAND2X1_480/B 0.05fF
C4839 POR2X1_49/Y PAND2X1_148/Y 0.03fF
C4840 POR2X1_290/Y VDD 0.13fF
C4841 PAND2X1_63/Y POR2X1_641/a_16_28# 0.07fF
C4842 POR2X1_57/A PAND2X1_453/A 0.04fF
C4843 POR2X1_829/A INPUT_0 0.03fF
C4844 POR2X1_16/A PAND2X1_590/O 0.00fF
C4845 POR2X1_330/Y POR2X1_541/CTRL2 0.03fF
C4846 POR2X1_404/a_16_28# POR2X1_35/Y 0.01fF
C4847 PAND2X1_382/O POR2X1_29/A 0.04fF
C4848 POR2X1_100/CTRL2 POR2X1_99/A 0.01fF
C4849 POR2X1_670/a_16_28# POR2X1_42/Y 0.03fF
C4850 POR2X1_147/A POR2X1_830/A 0.00fF
C4851 POR2X1_119/CTRL VDD 0.00fF
C4852 POR2X1_65/A PAND2X1_547/O 0.01fF
C4853 POR2X1_174/O POR2X1_567/B 0.04fF
C4854 POR2X1_734/A PAND2X1_32/B 0.33fF
C4855 PAND2X1_56/Y POR2X1_335/CTRL2 0.14fF
C4856 POR2X1_13/A PAND2X1_784/CTRL2 0.00fF
C4857 POR2X1_814/A POR2X1_343/a_76_344# 0.00fF
C4858 PAND2X1_862/B POR2X1_293/Y 0.03fF
C4859 POR2X1_135/Y POR2X1_45/Y 0.06fF
C4860 PAND2X1_93/B POR2X1_733/Y 0.03fF
C4861 PAND2X1_69/A POR2X1_585/CTRL 0.01fF
C4862 POR2X1_862/A POR2X1_774/A 0.03fF
C4863 POR2X1_188/A POR2X1_121/CTRL2 0.01fF
C4864 POR2X1_49/Y POR2X1_38/B 0.03fF
C4865 POR2X1_259/CTRL POR2X1_555/B 0.01fF
C4866 PAND2X1_205/a_16_344# PAND2X1_853/B 0.02fF
C4867 POR2X1_57/A POR2X1_279/Y 0.01fF
C4868 POR2X1_614/A PAND2X1_581/Y 0.01fF
C4869 POR2X1_238/Y VDD 0.13fF
C4870 PAND2X1_20/A PAND2X1_505/a_76_28# 0.01fF
C4871 POR2X1_667/A PAND2X1_559/CTRL2 0.01fF
C4872 PAND2X1_658/B VDD 1.20fF
C4873 POR2X1_70/a_16_28# POR2X1_96/A 0.05fF
C4874 POR2X1_55/Y PAND2X1_515/CTRL 0.01fF
C4875 POR2X1_14/Y POR2X1_584/Y 0.03fF
C4876 POR2X1_388/O PAND2X1_65/B 0.01fF
C4877 POR2X1_686/a_76_344# POR2X1_750/B 0.01fF
C4878 POR2X1_46/Y POR2X1_42/Y 0.05fF
C4879 PAND2X1_140/CTRL POR2X1_387/Y 0.00fF
C4880 PAND2X1_94/A POR2X1_285/Y 0.03fF
C4881 PAND2X1_222/O PAND2X1_643/A 0.01fF
C4882 POR2X1_549/B D_INPUT_1 0.03fF
C4883 POR2X1_723/CTRL POR2X1_723/B 0.01fF
C4884 PAND2X1_659/Y POR2X1_490/Y 0.03fF
C4885 PAND2X1_222/A PAND2X1_643/A 0.02fF
C4886 POR2X1_43/B POR2X1_586/CTRL2 0.03fF
C4887 POR2X1_786/Y VDD -0.00fF
C4888 POR2X1_23/Y PAND2X1_851/CTRL2 0.03fF
C4889 PAND2X1_671/O PAND2X1_58/A 0.02fF
C4890 PAND2X1_206/CTRL2 POR2X1_73/Y 0.01fF
C4891 POR2X1_775/O VDD 0.00fF
C4892 POR2X1_407/A POR2X1_435/Y 0.11fF
C4893 POR2X1_853/a_16_28# POR2X1_776/B 0.00fF
C4894 POR2X1_65/A POR2X1_597/O 0.01fF
C4895 POR2X1_669/B PAND2X1_560/B 0.02fF
C4896 POR2X1_497/Y POR2X1_521/a_16_28# 0.02fF
C4897 POR2X1_83/B PAND2X1_308/Y 0.03fF
C4898 POR2X1_43/B PAND2X1_553/B 0.07fF
C4899 VDD POR2X1_788/B 0.44fF
C4900 PAND2X1_65/Y POR2X1_360/O 0.01fF
C4901 POR2X1_185/CTRL2 PAND2X1_55/Y 0.03fF
C4902 PAND2X1_56/O POR2X1_804/A 0.04fF
C4903 POR2X1_43/B POR2X1_262/O 0.02fF
C4904 PAND2X1_735/Y POR2X1_498/A 0.02fF
C4905 PAND2X1_73/Y POR2X1_774/A 0.03fF
C4906 POR2X1_81/O POR2X1_153/Y 0.02fF
C4907 POR2X1_249/Y POR2X1_389/Y 0.03fF
C4908 PAND2X1_407/CTRL2 POR2X1_39/B 0.01fF
C4909 POR2X1_72/B POR2X1_530/O 0.01fF
C4910 PAND2X1_40/a_76_28# PAND2X1_587/Y 0.01fF
C4911 POR2X1_13/A POR2X1_417/O 0.18fF
C4912 POR2X1_316/Y PAND2X1_457/Y 0.01fF
C4913 PAND2X1_334/O POR2X1_42/Y 0.02fF
C4914 PAND2X1_732/A PAND2X1_169/Y 0.01fF
C4915 PAND2X1_624/CTRL POR2X1_283/A 0.02fF
C4916 POR2X1_793/CTRL POR2X1_713/B 0.01fF
C4917 PAND2X1_41/B POR2X1_502/CTRL 0.03fF
C4918 PAND2X1_91/CTRL POR2X1_169/A 0.02fF
C4919 POR2X1_199/O POR2X1_196/Y 0.02fF
C4920 PAND2X1_651/Y PAND2X1_215/B 0.05fF
C4921 PAND2X1_863/B POR2X1_38/Y 0.06fF
C4922 POR2X1_673/Y POR2X1_734/A 0.13fF
C4923 POR2X1_528/a_16_28# POR2X1_56/B 0.02fF
C4924 PAND2X1_320/O POR2X1_568/Y 0.04fF
C4925 PAND2X1_496/CTRL2 POR2X1_500/Y 0.00fF
C4926 POR2X1_417/CTRL POR2X1_293/Y 0.02fF
C4927 PAND2X1_665/CTRL2 POR2X1_66/A 0.01fF
C4928 POR2X1_119/Y POR2X1_32/A 0.34fF
C4929 POR2X1_416/B POR2X1_77/CTRL 0.12fF
C4930 PAND2X1_473/B PAND2X1_728/CTRL 0.02fF
C4931 POR2X1_597/A POR2X1_591/Y 0.00fF
C4932 POR2X1_260/Y POR2X1_203/Y 0.00fF
C4933 POR2X1_45/Y POR2X1_816/A 0.03fF
C4934 POR2X1_786/Y POR2X1_741/Y 0.07fF
C4935 PAND2X1_48/O POR2X1_366/A 0.13fF
C4936 POR2X1_614/A POR2X1_341/CTRL 0.01fF
C4937 PAND2X1_58/A PAND2X1_142/a_76_28# 0.01fF
C4938 PAND2X1_480/B POR2X1_7/A 0.05fF
C4939 PAND2X1_6/A POR2X1_184/Y 0.07fF
C4940 POR2X1_753/O POR2X1_752/Y 0.00fF
C4941 POR2X1_606/O PAND2X1_56/A 0.01fF
C4942 POR2X1_52/A POR2X1_583/a_56_344# 0.00fF
C4943 POR2X1_40/Y POR2X1_183/CTRL2 0.01fF
C4944 POR2X1_466/O POR2X1_209/A 0.03fF
C4945 POR2X1_341/A POR2X1_579/CTRL2 0.06fF
C4946 POR2X1_57/A POR2X1_55/Y 2.88fF
C4947 PAND2X1_738/Y PAND2X1_181/O 0.02fF
C4948 PAND2X1_682/CTRL PAND2X1_69/A 0.01fF
C4949 POR2X1_614/A POR2X1_559/Y 0.01fF
C4950 PAND2X1_640/B POR2X1_39/B 0.03fF
C4951 PAND2X1_48/B POR2X1_736/O 0.01fF
C4952 PAND2X1_69/A PAND2X1_146/O 0.04fF
C4953 PAND2X1_651/Y PAND2X1_6/A 0.10fF
C4954 POR2X1_566/A POR2X1_97/CTRL2 0.14fF
C4955 POR2X1_66/CTRL2 PAND2X1_69/A 0.01fF
C4956 PAND2X1_462/CTRL2 POR2X1_37/Y 0.03fF
C4957 POR2X1_140/B PAND2X1_96/B 0.64fF
C4958 POR2X1_480/A POR2X1_444/Y 0.07fF
C4959 PAND2X1_23/Y POR2X1_359/Y 0.01fF
C4960 POR2X1_740/Y PAND2X1_306/CTRL 0.00fF
C4961 PAND2X1_217/B PAND2X1_657/B 0.00fF
C4962 PAND2X1_76/Y POR2X1_153/Y 0.03fF
C4963 POR2X1_119/Y POR2X1_417/Y 0.05fF
C4964 POR2X1_41/B PAND2X1_196/CTRL 0.00fF
C4965 POR2X1_559/Y POR2X1_38/B 0.03fF
C4966 POR2X1_786/Y PAND2X1_32/B 0.07fF
C4967 PAND2X1_738/Y PAND2X1_343/CTRL 0.28fF
C4968 POR2X1_866/A PAND2X1_72/A 0.03fF
C4969 POR2X1_614/A POR2X1_644/A 0.03fF
C4970 POR2X1_775/O PAND2X1_32/B 0.01fF
C4971 PAND2X1_839/B PAND2X1_839/O 0.00fF
C4972 PAND2X1_808/CTRL POR2X1_283/A 0.01fF
C4973 POR2X1_567/A POR2X1_355/A 0.03fF
C4974 PAND2X1_476/A PAND2X1_231/CTRL2 0.00fF
C4975 POR2X1_156/O POR2X1_750/B 0.01fF
C4976 PAND2X1_48/B POR2X1_726/Y 0.01fF
C4977 INPUT_6 PAND2X1_587/O 0.15fF
C4978 POR2X1_596/A PAND2X1_69/A 0.43fF
C4979 INPUT_1 POR2X1_669/CTRL 0.00fF
C4980 POR2X1_532/A POR2X1_771/O 0.01fF
C4981 POR2X1_557/A POR2X1_786/A 0.04fF
C4982 PAND2X1_508/Y POR2X1_236/Y 0.03fF
C4983 PAND2X1_542/CTRL VDD 0.00fF
C4984 POR2X1_664/CTRL2 POR2X1_664/Y 0.01fF
C4985 PAND2X1_63/Y POR2X1_205/A 0.22fF
C4986 PAND2X1_847/CTRL POR2X1_32/A 0.11fF
C4987 PAND2X1_6/Y POR2X1_774/CTRL 0.01fF
C4988 POR2X1_390/B POR2X1_733/A 0.13fF
C4989 PAND2X1_60/CTRL2 PAND2X1_69/A 0.02fF
C4990 PAND2X1_476/A POR2X1_230/CTRL2 0.00fF
C4991 PAND2X1_241/CTRL2 PAND2X1_308/Y 0.01fF
C4992 POR2X1_83/B POR2X1_77/Y 2.27fF
C4993 POR2X1_170/CTRL POR2X1_566/B 0.01fF
C4994 PAND2X1_72/Y POR2X1_579/Y 0.00fF
C4995 POR2X1_65/A POR2X1_517/CTRL2 0.01fF
C4996 POR2X1_85/Y POR2X1_83/B 0.01fF
C4997 PAND2X1_358/A PAND2X1_351/Y 0.15fF
C4998 PAND2X1_657/B VDD 0.18fF
C4999 POR2X1_406/Y PAND2X1_716/B 0.06fF
C5000 POR2X1_111/Y POR2X1_55/Y 0.03fF
C5001 PAND2X1_651/Y POR2X1_588/Y 0.01fF
C5002 PAND2X1_56/Y POR2X1_456/B 0.06fF
C5003 PAND2X1_329/CTRL POR2X1_532/A 0.01fF
C5004 POR2X1_83/A POR2X1_16/A 0.03fF
C5005 POR2X1_192/Y POR2X1_564/CTRL 0.49fF
C5006 PAND2X1_216/B PAND2X1_798/B 0.03fF
C5007 POR2X1_101/O PAND2X1_69/A 0.03fF
C5008 POR2X1_383/A POR2X1_784/O 0.11fF
C5009 POR2X1_532/A POR2X1_222/A 0.04fF
C5010 POR2X1_416/B POR2X1_27/Y 0.00fF
C5011 POR2X1_9/Y PAND2X1_340/B 0.61fF
C5012 POR2X1_356/A POR2X1_351/B 0.05fF
C5013 PAND2X1_661/CTRL2 PAND2X1_659/Y 0.10fF
C5014 POR2X1_816/A POR2X1_171/O 0.01fF
C5015 POR2X1_172/Y POR2X1_530/Y 0.01fF
C5016 PAND2X1_850/Y PAND2X1_473/B 0.53fF
C5017 POR2X1_239/a_16_28# POR2X1_239/Y 0.02fF
C5018 PAND2X1_358/A PAND2X1_101/CTRL 0.02fF
C5019 POR2X1_537/Y POR2X1_722/Y 0.00fF
C5020 PAND2X1_553/B POR2X1_183/CTRL 0.04fF
C5021 POR2X1_575/B POR2X1_579/B 0.03fF
C5022 POR2X1_513/Y POR2X1_260/A 0.03fF
C5023 POR2X1_119/Y PAND2X1_35/Y 0.05fF
C5024 PAND2X1_691/Y PAND2X1_645/B 0.07fF
C5025 POR2X1_16/A POR2X1_90/Y 0.03fF
C5026 PAND2X1_723/a_76_28# PAND2X1_723/A 0.01fF
C5027 POR2X1_614/A PAND2X1_72/Y 0.63fF
C5028 POR2X1_316/CTRL POR2X1_43/B 0.01fF
C5029 POR2X1_293/Y PAND2X1_716/B 0.14fF
C5030 PAND2X1_403/CTRL POR2X1_37/Y 0.01fF
C5031 POR2X1_219/B POR2X1_260/A 0.07fF
C5032 POR2X1_440/Y POR2X1_478/B 0.14fF
C5033 PAND2X1_835/a_16_344# POR2X1_394/A 0.01fF
C5034 POR2X1_12/A POR2X1_18/CTRL 0.01fF
C5035 D_INPUT_5 POR2X1_18/O 0.01fF
C5036 POR2X1_365/Y POR2X1_192/B 1.41fF
C5037 POR2X1_178/O PAND2X1_348/A 0.03fF
C5038 PAND2X1_568/B PAND2X1_578/O 0.01fF
C5039 PAND2X1_23/Y POR2X1_359/CTRL 0.01fF
C5040 POR2X1_485/Y POR2X1_20/B 0.58fF
C5041 POR2X1_825/Y PAND2X1_721/B 0.05fF
C5042 POR2X1_85/CTRL PAND2X1_35/Y 0.01fF
C5043 POR2X1_755/Y POR2X1_757/Y 0.17fF
C5044 PAND2X1_797/Y POR2X1_763/Y 0.07fF
C5045 POR2X1_213/B PAND2X1_52/B 0.03fF
C5046 POR2X1_16/A POR2X1_167/CTRL2 0.01fF
C5047 PAND2X1_93/B PAND2X1_86/CTRL 0.09fF
C5048 PAND2X1_777/CTRL2 POR2X1_387/Y 0.06fF
C5049 POR2X1_383/A POR2X1_456/B 0.06fF
C5050 POR2X1_677/Y POR2X1_102/Y 0.03fF
C5051 POR2X1_332/Y POR2X1_556/Y 0.00fF
C5052 POR2X1_496/O POR2X1_20/B 0.01fF
C5053 POR2X1_366/A POR2X1_260/A 0.05fF
C5054 POR2X1_119/Y POR2X1_184/Y 0.03fF
C5055 POR2X1_362/B POR2X1_717/B 0.03fF
C5056 PAND2X1_446/Y POR2X1_424/Y 0.06fF
C5057 POR2X1_431/CTRL2 POR2X1_37/Y 0.01fF
C5058 POR2X1_516/a_16_28# PAND2X1_508/Y 0.09fF
C5059 POR2X1_407/Y PAND2X1_18/B 0.03fF
C5060 POR2X1_463/Y POR2X1_710/Y 0.01fF
C5061 POR2X1_614/A POR2X1_512/O 0.01fF
C5062 PAND2X1_658/A PAND2X1_860/CTRL 0.01fF
C5063 POR2X1_464/Y POR2X1_542/a_16_28# 0.03fF
C5064 POR2X1_7/B POR2X1_39/B 21.15fF
C5065 PAND2X1_462/CTRL2 POR2X1_293/Y 0.01fF
C5066 PAND2X1_137/Y POR2X1_416/B 0.03fF
C5067 POR2X1_65/CTRL2 D_INPUT_0 0.01fF
C5068 POR2X1_375/O POR2X1_260/A 0.02fF
C5069 PAND2X1_862/B PAND2X1_862/CTRL2 0.04fF
C5070 PAND2X1_436/A POR2X1_677/Y 0.03fF
C5071 PAND2X1_653/O POR2X1_594/Y -0.00fF
C5072 PAND2X1_659/Y PAND2X1_676/CTRL 0.00fF
C5073 POR2X1_13/A PAND2X1_351/A 0.06fF
C5074 POR2X1_518/a_76_344# POR2X1_519/Y 0.03fF
C5075 POR2X1_90/Y POR2X1_320/a_16_28# 0.03fF
C5076 POR2X1_38/Y PAND2X1_737/CTRL 0.01fF
C5077 PAND2X1_738/Y POR2X1_167/Y 0.03fF
C5078 POR2X1_270/Y POR2X1_116/A 0.00fF
C5079 INPUT_1 PAND2X1_701/CTRL2 0.01fF
C5080 PAND2X1_39/B POR2X1_647/CTRL 0.00fF
C5081 PAND2X1_797/Y POR2X1_73/Y 0.03fF
C5082 PAND2X1_259/O PAND2X1_771/Y 0.31fF
C5083 PAND2X1_242/CTRL POR2X1_77/Y 0.03fF
C5084 POR2X1_73/Y PAND2X1_860/CTRL 0.01fF
C5085 POR2X1_669/Y POR2X1_667/Y 0.06fF
C5086 POR2X1_813/CTRL2 POR2X1_263/Y 0.01fF
C5087 POR2X1_123/CTRL PAND2X1_72/A 0.04fF
C5088 POR2X1_661/A POR2X1_480/A 0.07fF
C5089 POR2X1_35/B POR2X1_621/CTRL2 0.01fF
C5090 POR2X1_129/Y POR2X1_260/A 0.03fF
C5091 POR2X1_44/a_76_344# PAND2X1_635/Y 0.00fF
C5092 POR2X1_447/B POR2X1_854/B 0.05fF
C5093 POR2X1_101/Y POR2X1_294/A 0.07fF
C5094 POR2X1_23/Y PAND2X1_407/CTRL 0.00fF
C5095 POR2X1_532/A PAND2X1_134/a_56_28# 0.00fF
C5096 PAND2X1_865/O PAND2X1_862/Y 0.01fF
C5097 POR2X1_383/CTRL POR2X1_520/A 0.01fF
C5098 PAND2X1_41/O POR2X1_66/A 0.02fF
C5099 POR2X1_861/CTRL PAND2X1_72/A 0.01fF
C5100 POR2X1_805/A PAND2X1_52/B 0.01fF
C5101 POR2X1_443/A POR2X1_220/B 0.01fF
C5102 PAND2X1_111/CTRL PAND2X1_72/A 0.00fF
C5103 POR2X1_65/A POR2X1_292/a_76_344# 0.01fF
C5104 PAND2X1_860/A PAND2X1_804/B 0.09fF
C5105 POR2X1_43/Y POR2X1_519/Y 0.66fF
C5106 POR2X1_319/A POR2X1_856/B 0.03fF
C5107 PAND2X1_796/B PAND2X1_796/O 0.00fF
C5108 POR2X1_567/A POR2X1_799/a_56_344# 0.00fF
C5109 PAND2X1_437/a_16_344# POR2X1_192/Y 0.04fF
C5110 POR2X1_506/CTRL POR2X1_508/B 0.00fF
C5111 POR2X1_38/CTRL POR2X1_37/Y 0.01fF
C5112 PAND2X1_206/B PAND2X1_340/CTRL 0.01fF
C5113 POR2X1_491/CTRL POR2X1_150/Y 0.01fF
C5114 POR2X1_814/B POR2X1_624/B 1.75fF
C5115 POR2X1_329/A POR2X1_511/Y 0.07fF
C5116 PAND2X1_72/A POR2X1_501/B 0.03fF
C5117 PAND2X1_403/CTRL POR2X1_293/Y 0.01fF
C5118 PAND2X1_159/O PAND2X1_9/Y 0.02fF
C5119 PAND2X1_640/B POR2X1_48/A 0.01fF
C5120 POR2X1_649/a_76_344# POR2X1_643/A 0.00fF
C5121 POR2X1_731/a_76_344# PAND2X1_52/B 0.01fF
C5122 POR2X1_480/O POR2X1_478/Y 0.00fF
C5123 PAND2X1_606/CTRL2 POR2X1_102/Y 0.00fF
C5124 POR2X1_49/CTRL PAND2X1_9/Y 0.01fF
C5125 POR2X1_378/CTRL PAND2X1_9/Y 0.01fF
C5126 POR2X1_475/CTRL2 POR2X1_734/A 0.02fF
C5127 POR2X1_663/B POR2X1_750/B 0.06fF
C5128 POR2X1_681/Y POR2X1_60/A 1.12fF
C5129 POR2X1_523/A POR2X1_523/B 0.02fF
C5130 POR2X1_774/CTRL PAND2X1_52/B 0.01fF
C5131 POR2X1_624/Y POR2X1_330/Y 0.07fF
C5132 PAND2X1_657/CTRL2 POR2X1_23/Y 0.00fF
C5133 POR2X1_502/A POR2X1_814/A 0.15fF
C5134 PAND2X1_23/Y POR2X1_837/A 0.21fF
C5135 PAND2X1_806/O PAND2X1_362/A 0.04fF
C5136 PAND2X1_3/A PAND2X1_36/a_16_344# 0.01fF
C5137 PAND2X1_47/B PAND2X1_59/B 0.03fF
C5138 PAND2X1_635/Y POR2X1_587/O 0.01fF
C5139 POR2X1_466/A POR2X1_590/A 0.05fF
C5140 POR2X1_568/A POR2X1_319/Y 0.03fF
C5141 POR2X1_477/O POR2X1_480/A 0.04fF
C5142 PAND2X1_357/a_76_28# PAND2X1_353/Y 0.02fF
C5143 POR2X1_502/A POR2X1_846/Y 0.04fF
C5144 POR2X1_48/A POR2X1_393/Y 0.01fF
C5145 POR2X1_450/CTRL POR2X1_121/B 0.08fF
C5146 POR2X1_66/B PAND2X1_666/O 0.01fF
C5147 POR2X1_411/B PAND2X1_719/O 0.03fF
C5148 PAND2X1_817/CTRL PAND2X1_381/Y 0.01fF
C5149 PAND2X1_817/CTRL2 POR2X1_29/A 0.01fF
C5150 POR2X1_650/A POR2X1_260/B 0.02fF
C5151 POR2X1_416/B PAND2X1_853/B 0.10fF
C5152 POR2X1_497/CTRL POR2X1_32/A 0.01fF
C5153 PAND2X1_437/CTRL PAND2X1_60/B 0.01fF
C5154 POR2X1_78/A POR2X1_474/CTRL2 0.01fF
C5155 PAND2X1_416/O VDD 0.00fF
C5156 PAND2X1_802/O PAND2X1_798/Y 0.08fF
C5157 POR2X1_41/B PAND2X1_838/O 0.04fF
C5158 POR2X1_661/A PAND2X1_305/O 0.06fF
C5159 PAND2X1_61/CTRL2 PAND2X1_61/Y 0.01fF
C5160 POR2X1_96/A PAND2X1_203/O 0.03fF
C5161 POR2X1_805/a_16_28# POR2X1_805/B 0.02fF
C5162 POR2X1_605/B POR2X1_78/A 0.05fF
C5163 POR2X1_411/B PAND2X1_269/CTRL2 0.01fF
C5164 POR2X1_830/O POR2X1_830/Y 0.01fF
C5165 PAND2X1_57/B POR2X1_446/B 0.03fF
C5166 POR2X1_502/A POR2X1_444/B 0.00fF
C5167 PAND2X1_73/Y POR2X1_780/O 0.01fF
C5168 POR2X1_490/Y POR2X1_406/Y 0.03fF
C5169 POR2X1_119/Y PAND2X1_858/B 0.10fF
C5170 POR2X1_322/a_56_344# POR2X1_441/Y 0.00fF
C5171 POR2X1_654/CTRL POR2X1_121/B 0.01fF
C5172 POR2X1_559/a_16_28# POR2X1_814/A 0.02fF
C5173 PAND2X1_773/Y PAND2X1_580/B 0.30fF
C5174 POR2X1_852/B POR2X1_202/B 0.10fF
C5175 POR2X1_415/A POR2X1_617/CTRL 0.08fF
C5176 POR2X1_65/A PAND2X1_223/B 0.16fF
C5177 POR2X1_857/A POR2X1_795/B 0.04fF
C5178 POR2X1_496/Y POR2X1_627/CTRL2 0.05fF
C5179 POR2X1_20/B PAND2X1_339/Y 0.02fF
C5180 POR2X1_335/CTRL POR2X1_66/A 0.00fF
C5181 POR2X1_302/B PAND2X1_279/O 0.02fF
C5182 POR2X1_290/O POR2X1_83/B 0.03fF
C5183 POR2X1_665/CTRL2 POR2X1_665/A 0.01fF
C5184 PAND2X1_304/O PAND2X1_56/A 0.04fF
C5185 POR2X1_104/CTRL2 POR2X1_5/Y 0.00fF
C5186 PAND2X1_863/O POR2X1_102/Y 0.05fF
C5187 PAND2X1_201/CTRL PAND2X1_341/A 0.01fF
C5188 POR2X1_516/CTRL2 POR2X1_257/A 0.01fF
C5189 POR2X1_556/A POR2X1_804/A 0.03fF
C5190 POR2X1_158/O POR2X1_416/B 0.22fF
C5191 POR2X1_856/a_16_28# PAND2X1_73/Y 0.02fF
C5192 POR2X1_678/CTRL2 PAND2X1_69/A 0.01fF
C5193 PAND2X1_576/B POR2X1_46/Y 0.03fF
C5194 PAND2X1_20/A POR2X1_849/O 0.01fF
C5195 POR2X1_78/A POR2X1_549/B 0.04fF
C5196 POR2X1_436/B VDD 0.11fF
C5197 POR2X1_260/B POR2X1_294/B 2.17fF
C5198 POR2X1_68/A POR2X1_676/CTRL 0.03fF
C5199 POR2X1_407/A POR2X1_676/CTRL2 0.03fF
C5200 PAND2X1_830/Y POR2X1_48/A 0.02fF
C5201 POR2X1_81/a_16_28# PAND2X1_474/A 0.02fF
C5202 PAND2X1_485/a_76_28# PAND2X1_57/B 0.03fF
C5203 POR2X1_609/Y POR2X1_607/Y 0.01fF
C5204 PAND2X1_6/Y PAND2X1_39/B 1.19fF
C5205 PAND2X1_249/a_76_28# PAND2X1_733/A 0.01fF
C5206 POR2X1_48/A POR2X1_7/B 0.19fF
C5207 POR2X1_862/B POR2X1_777/B 0.05fF
C5208 PAND2X1_474/Y POR2X1_497/CTRL2 0.00fF
C5209 POR2X1_48/A POR2X1_277/O 0.01fF
C5210 PAND2X1_23/Y POR2X1_567/B 0.08fF
C5211 PAND2X1_48/B POR2X1_856/B 0.06fF
C5212 PAND2X1_650/CTRL2 PAND2X1_9/Y 0.01fF
C5213 PAND2X1_73/Y POR2X1_445/CTRL2 0.01fF
C5214 POR2X1_20/B PAND2X1_344/O 0.05fF
C5215 PAND2X1_602/Y PAND2X1_645/Y 0.26fF
C5216 PAND2X1_240/CTRL2 POR2X1_5/Y 0.01fF
C5217 POR2X1_411/B POR2X1_142/Y 0.03fF
C5218 POR2X1_555/A POR2X1_186/Y 0.23fF
C5219 PAND2X1_195/CTRL2 VDD 0.00fF
C5220 POR2X1_278/Y POR2X1_102/Y 0.12fF
C5221 POR2X1_264/Y POR2X1_558/B 0.12fF
C5222 PAND2X1_57/B POR2X1_121/B 0.03fF
C5223 POR2X1_657/Y POR2X1_228/Y 0.12fF
C5224 POR2X1_114/B POR2X1_458/O 0.01fF
C5225 GATE_479 POR2X1_376/B 0.03fF
C5226 POR2X1_66/A POR2X1_732/B 0.12fF
C5227 POR2X1_865/B POR2X1_647/B 0.02fF
C5228 POR2X1_411/B PAND2X1_175/B 0.03fF
C5229 PAND2X1_862/B POR2X1_60/A 0.03fF
C5230 PAND2X1_124/Y POR2X1_52/Y 0.33fF
C5231 POR2X1_536/Y INPUT_0 0.00fF
C5232 D_INPUT_3 PAND2X1_415/a_16_344# 0.02fF
C5233 POR2X1_264/O INPUT_0 0.06fF
C5234 POR2X1_555/B POR2X1_785/A 0.03fF
C5235 POR2X1_413/A PAND2X1_647/B 0.01fF
C5236 POR2X1_116/A POR2X1_101/Y 0.10fF
C5237 PAND2X1_90/A POR2X1_623/B 0.02fF
C5238 POR2X1_96/A PAND2X1_76/O 0.01fF
C5239 POR2X1_329/A POR2X1_129/Y 0.03fF
C5240 POR2X1_270/a_76_344# POR2X1_445/A 0.00fF
C5241 PAND2X1_463/O PAND2X1_460/Y 0.06fF
C5242 POR2X1_838/B PAND2X1_55/Y 0.00fF
C5243 PAND2X1_793/Y PAND2X1_78/O 0.03fF
C5244 POR2X1_78/B PAND2X1_597/CTRL 0.01fF
C5245 POR2X1_427/CTRL2 PAND2X1_565/A 0.00fF
C5246 POR2X1_458/O POR2X1_458/B 0.00fF
C5247 POR2X1_146/CTRL POR2X1_257/A 0.00fF
C5248 PAND2X1_58/A POR2X1_42/Y 0.07fF
C5249 PAND2X1_478/Y PAND2X1_480/B 0.04fF
C5250 POR2X1_52/A POR2X1_750/A 0.03fF
C5251 D_INPUT_0 PAND2X1_69/A 0.53fF
C5252 POR2X1_61/Y POR2X1_215/CTRL 0.03fF
C5253 POR2X1_65/A POR2X1_88/Y 0.01fF
C5254 POR2X1_49/Y PAND2X1_350/A 0.01fF
C5255 POR2X1_20/B PAND2X1_726/B 0.08fF
C5256 PAND2X1_319/B POR2X1_298/a_16_28# 0.02fF
C5257 PAND2X1_454/a_16_344# POR2X1_60/A 0.01fF
C5258 PAND2X1_360/CTRL POR2X1_42/Y 0.01fF
C5259 PAND2X1_512/O POR2X1_7/B 0.15fF
C5260 POR2X1_811/A PAND2X1_69/A 0.03fF
C5261 D_INPUT_0 PAND2X1_341/A 0.05fF
C5262 POR2X1_750/B POR2X1_554/Y 0.05fF
C5263 POR2X1_96/A PAND2X1_541/a_16_344# 0.01fF
C5264 POR2X1_66/B PAND2X1_385/O 0.01fF
C5265 POR2X1_52/A POR2X1_306/Y 0.04fF
C5266 PAND2X1_659/Y POR2X1_329/A 0.03fF
C5267 POR2X1_669/B POR2X1_747/Y 0.01fF
C5268 PAND2X1_206/A PAND2X1_100/CTRL2 0.01fF
C5269 POR2X1_360/A PAND2X1_41/B 0.03fF
C5270 PAND2X1_478/B PAND2X1_478/CTRL 0.01fF
C5271 PAND2X1_65/O POR2X1_205/A 0.07fF
C5272 POR2X1_685/A POR2X1_676/a_16_28# 0.02fF
C5273 POR2X1_814/A POR2X1_188/Y 0.03fF
C5274 POR2X1_60/a_56_344# D_INPUT_0 0.01fF
C5275 PAND2X1_472/A PAND2X1_721/B 0.03fF
C5276 PAND2X1_814/CTRL POR2X1_669/B 0.32fF
C5277 POR2X1_52/A GATE_479 0.03fF
C5278 PAND2X1_20/A POR2X1_78/CTRL2 0.01fF
C5279 POR2X1_48/Y POR2X1_72/B 0.01fF
C5280 PAND2X1_791/O POR2X1_757/Y 0.00fF
C5281 POR2X1_814/B PAND2X1_183/O 0.32fF
C5282 PAND2X1_6/Y PAND2X1_20/A 0.10fF
C5283 POR2X1_590/A POR2X1_550/CTRL2 0.01fF
C5284 POR2X1_663/m4_208_n4# PAND2X1_90/Y 0.06fF
C5285 POR2X1_300/CTRL PAND2X1_217/B 0.04fF
C5286 POR2X1_252/CTRL2 POR2X1_5/Y 0.08fF
C5287 POR2X1_862/Y POR2X1_101/Y 0.00fF
C5288 INPUT_0 PAND2X1_730/B 0.03fF
C5289 POR2X1_508/CTRL2 POR2X1_852/B 0.06fF
C5290 POR2X1_275/Y POR2X1_129/Y 0.01fF
C5291 POR2X1_718/a_16_28# POR2X1_435/Y 0.01fF
C5292 POR2X1_96/A PAND2X1_473/B 0.03fF
C5293 PAND2X1_193/CTRL2 POR2X1_7/B 0.01fF
C5294 POR2X1_763/CTRL POR2X1_46/Y 0.01fF
C5295 PAND2X1_652/A POR2X1_72/B 0.05fF
C5296 INPUT_2 POR2X1_102/Y 0.01fF
C5297 POR2X1_65/A PAND2X1_453/O 0.01fF
C5298 POR2X1_355/CTRL PAND2X1_23/Y 0.01fF
C5299 PAND2X1_435/a_16_344# POR2X1_236/Y 0.02fF
C5300 PAND2X1_41/B POR2X1_350/CTRL2 0.04fF
C5301 PAND2X1_116/O PAND2X1_114/Y 0.00fF
C5302 POR2X1_186/Y PAND2X1_145/O 0.04fF
C5303 PAND2X1_362/A PAND2X1_362/a_76_28# 0.01fF
C5304 POR2X1_355/A PAND2X1_504/CTRL 0.01fF
C5305 POR2X1_237/Y POR2X1_417/Y 0.06fF
C5306 PAND2X1_824/B POR2X1_240/CTRL 0.01fF
C5307 POR2X1_306/CTRL POR2X1_102/Y 0.01fF
C5308 PAND2X1_836/O PAND2X1_403/B 0.00fF
C5309 POR2X1_61/Y POR2X1_740/Y 0.10fF
C5310 POR2X1_296/Y POR2X1_68/B 0.15fF
C5311 POR2X1_32/A PAND2X1_350/CTRL 0.00fF
C5312 POR2X1_94/A PAND2X1_6/A 0.21fF
C5313 POR2X1_483/A POR2X1_193/A 0.03fF
C5314 PAND2X1_860/A PAND2X1_332/Y 0.03fF
C5315 POR2X1_669/CTRL2 VDD 0.00fF
C5316 POR2X1_443/CTRL2 POR2X1_191/Y 0.11fF
C5317 INPUT_1 POR2X1_422/CTRL 0.01fF
C5318 POR2X1_832/B PAND2X1_589/CTRL 0.01fF
C5319 POR2X1_463/Y POR2X1_805/O 0.00fF
C5320 POR2X1_828/Y POR2X1_800/A 0.00fF
C5321 PAND2X1_137/Y PAND2X1_738/Y 0.05fF
C5322 PAND2X1_787/Y POR2X1_42/Y 0.01fF
C5323 POR2X1_43/B POR2X1_278/CTRL 0.28fF
C5324 PAND2X1_651/Y PAND2X1_456/CTRL2 0.30fF
C5325 POR2X1_192/Y POR2X1_223/O 0.01fF
C5326 POR2X1_221/CTRL POR2X1_221/Y 0.01fF
C5327 POR2X1_447/B POR2X1_66/a_16_28# 0.05fF
C5328 POR2X1_538/O POR2X1_814/B 0.01fF
C5329 PAND2X1_241/Y POR2X1_83/B 0.04fF
C5330 POR2X1_22/A INPUT_7 0.03fF
C5331 POR2X1_61/CTRL2 POR2X1_66/A 0.01fF
C5332 POR2X1_20/B PAND2X1_338/CTRL2 0.01fF
C5333 POR2X1_657/O POR2X1_228/Y 0.01fF
C5334 PAND2X1_137/CTRL2 POR2X1_96/A 0.03fF
C5335 POR2X1_78/B PAND2X1_23/Y 0.09fF
C5336 POR2X1_13/Y PAND2X1_193/O -0.00fF
C5337 PAND2X1_6/Y POR2X1_814/B 0.21fF
C5338 POR2X1_20/B PAND2X1_352/CTRL 0.01fF
C5339 POR2X1_809/A POR2X1_676/O 0.01fF
C5340 PAND2X1_206/B POR2X1_39/B 0.09fF
C5341 PAND2X1_41/B POR2X1_758/CTRL2 0.03fF
C5342 POR2X1_300/CTRL VDD 0.00fF
C5343 POR2X1_833/A POR2X1_499/a_56_344# 0.00fF
C5344 PAND2X1_470/CTRL2 PAND2X1_803/A 0.00fF
C5345 POR2X1_96/B POR2X1_14/Y 0.06fF
C5346 POR2X1_68/B POR2X1_392/B 0.09fF
C5347 POR2X1_852/A POR2X1_578/Y 0.01fF
C5348 POR2X1_68/A PAND2X1_525/a_76_28# 0.01fF
C5349 PAND2X1_48/B POR2X1_722/Y 0.01fF
C5350 POR2X1_763/A PAND2X1_711/A 0.07fF
C5351 PAND2X1_705/CTRL VDD 0.00fF
C5352 POR2X1_278/Y PAND2X1_808/Y 0.03fF
C5353 POR2X1_614/A POR2X1_483/A 0.05fF
C5354 PAND2X1_217/B PAND2X1_572/a_16_344# 0.10fF
C5355 PAND2X1_865/Y POR2X1_257/A 0.03fF
C5356 PAND2X1_90/Y PAND2X1_69/A 0.35fF
C5357 POR2X1_254/Y POR2X1_775/A 0.03fF
C5358 PAND2X1_6/Y POR2X1_325/A 4.34fF
C5359 D_GATE_662 POR2X1_192/Y 0.10fF
C5360 POR2X1_672/A VDD 0.00fF
C5361 POR2X1_491/Y POR2X1_150/Y 0.01fF
C5362 PAND2X1_794/B PAND2X1_580/B 0.00fF
C5363 POR2X1_680/Y PAND2X1_191/Y 0.03fF
C5364 PAND2X1_63/Y POR2X1_786/CTRL 0.02fF
C5365 POR2X1_646/O POR2X1_294/B 0.01fF
C5366 POR2X1_814/B POR2X1_791/A 0.01fF
C5367 PAND2X1_65/B PAND2X1_26/CTRL2 0.01fF
C5368 POR2X1_215/CTRL POR2X1_35/Y 0.01fF
C5369 PAND2X1_56/Y PAND2X1_57/B 0.56fF
C5370 POR2X1_537/Y POR2X1_866/A 0.03fF
C5371 POR2X1_333/Y POR2X1_97/A 0.03fF
C5372 POR2X1_319/A POR2X1_191/Y 0.24fF
C5373 POR2X1_614/A PAND2X1_8/Y 0.06fF
C5374 POR2X1_652/Y POR2X1_740/Y 0.00fF
C5375 POR2X1_22/A INPUT_4 0.06fF
C5376 POR2X1_722/B PAND2X1_55/Y 0.03fF
C5377 POR2X1_402/CTRL PAND2X1_60/B 0.01fF
C5378 POR2X1_567/A POR2X1_260/B 0.05fF
C5379 POR2X1_57/A POR2X1_511/Y 0.10fF
C5380 PAND2X1_55/Y POR2X1_294/B 0.35fF
C5381 POR2X1_102/Y POR2X1_530/a_16_28# 0.09fF
C5382 PAND2X1_377/Y POR2X1_42/Y 0.04fF
C5383 POR2X1_366/Y PAND2X1_55/Y 0.07fF
C5384 POR2X1_41/B PAND2X1_357/Y 0.03fF
C5385 POR2X1_750/m4_208_n4# POR2X1_720/A 0.01fF
C5386 POR2X1_218/Y PAND2X1_48/A 0.10fF
C5387 POR2X1_614/A POR2X1_812/O 0.01fF
C5388 POR2X1_38/B PAND2X1_8/Y 0.08fF
C5389 POR2X1_193/A POR2X1_795/m4_208_n4# 0.09fF
C5390 POR2X1_122/CTRL2 POR2X1_102/Y 0.01fF
C5391 POR2X1_407/A POR2X1_708/B 0.00fF
C5392 POR2X1_800/A PAND2X1_599/CTRL2 0.00fF
C5393 PAND2X1_65/B POR2X1_510/Y 0.03fF
C5394 POR2X1_578/Y POR2X1_775/CTRL2 0.10fF
C5395 POR2X1_496/Y PAND2X1_156/A 0.10fF
C5396 POR2X1_777/B POR2X1_276/Y 0.03fF
C5397 POR2X1_28/O POR2X1_4/Y 0.06fF
C5398 POR2X1_403/m4_208_n4# PAND2X1_60/B 0.08fF
C5399 D_INPUT_0 POR2X1_512/CTRL 0.01fF
C5400 POR2X1_788/Y POR2X1_294/B 0.03fF
C5401 PAND2X1_308/Y PAND2X1_444/Y 0.09fF
C5402 PAND2X1_95/B PAND2X1_95/a_76_28# 0.01fF
C5403 POR2X1_49/Y PAND2X1_714/Y 0.07fF
C5404 INPUT_1 POR2X1_24/O 0.02fF
C5405 POR2X1_35/Y POR2X1_740/Y 0.05fF
C5406 POR2X1_387/Y VDD 5.88fF
C5407 POR2X1_283/A POR2X1_236/Y 0.13fF
C5408 POR2X1_345/O POR2X1_330/Y 0.09fF
C5409 POR2X1_764/O POR2X1_40/Y 0.03fF
C5410 PAND2X1_863/B POR2X1_591/Y 0.03fF
C5411 POR2X1_20/CTRL2 POR2X1_38/B 0.00fF
C5412 POR2X1_102/CTRL2 POR2X1_37/Y 0.00fF
C5413 POR2X1_73/Y POR2X1_372/Y 0.07fF
C5414 PAND2X1_56/Y POR2X1_715/m4_208_n4# 0.06fF
C5415 POR2X1_38/Y PAND2X1_598/a_56_28# 0.00fF
C5416 POR2X1_337/O POR2X1_335/Y 0.04fF
C5417 POR2X1_409/CTRL POR2X1_55/Y 0.01fF
C5418 PAND2X1_649/A PAND2X1_400/CTRL2 0.01fF
C5419 POR2X1_599/A PAND2X1_717/a_16_344# 0.01fF
C5420 PAND2X1_65/B POR2X1_276/Y 0.03fF
C5421 PAND2X1_572/CTRL2 PAND2X1_364/B 0.05fF
C5422 POR2X1_239/CTRL POR2X1_55/Y 0.03fF
C5423 POR2X1_394/A POR2X1_40/Y 0.51fF
C5424 POR2X1_85/Y PAND2X1_206/A 0.02fF
C5425 POR2X1_504/CTRL POR2X1_504/Y 0.01fF
C5426 POR2X1_330/Y POR2X1_186/B 0.03fF
C5427 POR2X1_41/B POR2X1_278/A 0.00fF
C5428 PAND2X1_39/B PAND2X1_52/B 0.18fF
C5429 D_INPUT_7 PAND2X1_11/CTRL 0.01fF
C5430 POR2X1_8/Y POR2X1_65/A 0.06fF
C5431 POR2X1_407/Y POR2X1_294/B 0.00fF
C5432 POR2X1_60/A PAND2X1_716/B 7.27fF
C5433 POR2X1_90/Y PAND2X1_324/Y 1.28fF
C5434 POR2X1_763/Y POR2X1_526/Y 0.07fF
C5435 POR2X1_383/A PAND2X1_57/B 0.20fF
C5436 POR2X1_316/a_56_344# PAND2X1_390/Y 0.00fF
C5437 POR2X1_66/B POR2X1_113/B 0.03fF
C5438 POR2X1_55/Y POR2X1_9/CTRL2 0.16fF
C5439 PAND2X1_858/O POR2X1_271/Y 0.00fF
C5440 POR2X1_627/Y POR2X1_7/A 0.04fF
C5441 POR2X1_602/B POR2X1_722/CTRL2 0.01fF
C5442 POR2X1_335/B POR2X1_740/Y 0.03fF
C5443 POR2X1_96/B PAND2X1_472/B 0.01fF
C5444 POR2X1_519/Y POR2X1_73/Y 0.07fF
C5445 POR2X1_32/A PAND2X1_326/B 0.02fF
C5446 PAND2X1_702/a_16_344# POR2X1_42/Y 0.00fF
C5447 POR2X1_176/CTRL POR2X1_312/Y 0.01fF
C5448 POR2X1_347/A POR2X1_402/a_16_28# 0.02fF
C5449 POR2X1_574/CTRL2 POR2X1_724/A 0.01fF
C5450 POR2X1_693/CTRL PAND2X1_550/B 0.01fF
C5451 POR2X1_416/B POR2X1_23/Y 0.77fF
C5452 PAND2X1_55/Y PAND2X1_111/B 0.03fF
C5453 POR2X1_327/Y POR2X1_850/A 0.12fF
C5454 POR2X1_68/B PAND2X1_19/CTRL2 0.01fF
C5455 PAND2X1_784/CTRL POR2X1_7/A 0.09fF
C5456 INPUT_0 POR2X1_456/B 0.03fF
C5457 POR2X1_16/A INPUT_0 0.06fF
C5458 PAND2X1_506/CTRL POR2X1_239/Y 0.01fF
C5459 D_GATE_222 POR2X1_775/a_16_28# 0.05fF
C5460 POR2X1_78/B POR2X1_719/B 0.10fF
C5461 POR2X1_376/B PAND2X1_156/B 0.01fF
C5462 POR2X1_131/Y POR2X1_13/A 0.13fF
C5463 POR2X1_840/CTRL POR2X1_513/Y 0.02fF
C5464 POR2X1_660/Y POR2X1_513/A 0.01fF
C5465 PAND2X1_639/B POR2X1_408/Y 0.35fF
C5466 POR2X1_72/B PAND2X1_506/Y 0.03fF
C5467 PAND2X1_41/B POR2X1_571/Y 0.03fF
C5468 POR2X1_724/CTRL2 POR2X1_703/Y 0.01fF
C5469 POR2X1_65/A POR2X1_176/O 0.01fF
C5470 PAND2X1_275/O PAND2X1_60/B 0.08fF
C5471 POR2X1_336/CTRL PAND2X1_69/A 0.01fF
C5472 POR2X1_68/A PAND2X1_747/O 0.01fF
C5473 POR2X1_383/A POR2X1_341/CTRL2 0.03fF
C5474 POR2X1_334/B PAND2X1_63/B 0.03fF
C5475 POR2X1_123/Y PAND2X1_96/B 0.01fF
C5476 INPUT_1 POR2X1_754/A 0.29fF
C5477 PAND2X1_90/A POR2X1_561/CTRL2 0.03fF
C5478 POR2X1_390/B POR2X1_337/O 0.00fF
C5479 PAND2X1_48/B POR2X1_151/CTRL2 0.03fF
C5480 POR2X1_48/a_16_28# POR2X1_153/Y 0.09fF
C5481 PAND2X1_384/CTRL VDD 0.00fF
C5482 PAND2X1_96/B POR2X1_736/CTRL 0.01fF
C5483 PAND2X1_638/CTRL2 POR2X1_588/Y 0.01fF
C5484 D_GATE_662 POR2X1_568/Y 0.10fF
C5485 POR2X1_635/B PAND2X1_762/CTRL2 0.10fF
C5486 POR2X1_293/Y POR2X1_260/A 0.07fF
C5487 POR2X1_65/A POR2X1_177/m4_208_n4# 0.07fF
C5488 PAND2X1_480/B POR2X1_153/Y 0.05fF
C5489 POR2X1_740/Y PAND2X1_368/O 0.05fF
C5490 POR2X1_52/A PAND2X1_620/O 0.05fF
C5491 POR2X1_36/B POR2X1_582/CTRL 0.01fF
C5492 D_INPUT_3 PAND2X1_509/CTRL 0.02fF
C5493 INPUT_1 PAND2X1_341/O 0.01fF
C5494 PAND2X1_812/A PAND2X1_366/Y 0.01fF
C5495 POR2X1_356/A POR2X1_782/O 0.03fF
C5496 POR2X1_725/Y POR2X1_513/Y 0.07fF
C5497 POR2X1_90/Y PAND2X1_549/B 0.03fF
C5498 POR2X1_662/Y POR2X1_353/A 0.01fF
C5499 PAND2X1_48/B POR2X1_244/Y 0.03fF
C5500 PAND2X1_20/A POR2X1_725/CTRL 0.01fF
C5501 POR2X1_750/B POR2X1_39/B 0.10fF
C5502 POR2X1_416/B PAND2X1_221/O 0.05fF
C5503 PAND2X1_841/CTRL2 POR2X1_153/Y 0.00fF
C5504 PAND2X1_20/A POR2X1_500/CTRL 0.01fF
C5505 PAND2X1_94/A PAND2X1_283/a_16_344# 0.04fF
C5506 POR2X1_36/B POR2X1_582/A 0.03fF
C5507 POR2X1_16/A POR2X1_234/CTRL2 0.01fF
C5508 PAND2X1_20/A PAND2X1_52/B 0.14fF
C5509 PAND2X1_69/A PAND2X1_133/CTRL 0.01fF
C5510 POR2X1_378/Y POR2X1_62/Y 0.02fF
C5511 POR2X1_730/B POR2X1_730/Y 0.09fF
C5512 POR2X1_394/A PAND2X1_188/a_16_344# 0.04fF
C5513 POR2X1_461/Y POR2X1_848/a_16_28# 0.03fF
C5514 POR2X1_62/Y POR2X1_7/B 0.03fF
C5515 POR2X1_440/Y POR2X1_209/A 0.69fF
C5516 POR2X1_566/A POR2X1_540/Y 0.08fF
C5517 POR2X1_416/B POR2X1_312/Y 0.79fF
C5518 POR2X1_328/CTRL INPUT_5 0.01fF
C5519 POR2X1_328/O INPUT_4 0.02fF
C5520 POR2X1_333/A POR2X1_568/A 0.07fF
C5521 PAND2X1_106/CTRL2 POR2X1_383/A 0.03fF
C5522 POR2X1_301/A POR2X1_458/Y 0.01fF
C5523 POR2X1_111/a_16_28# POR2X1_283/A 0.08fF
C5524 PAND2X1_23/Y POR2X1_294/A 0.16fF
C5525 POR2X1_677/a_76_344# POR2X1_77/Y 0.01fF
C5526 POR2X1_65/A PAND2X1_326/CTRL2 0.03fF
C5527 POR2X1_416/B PAND2X1_740/O 0.01fF
C5528 PAND2X1_850/Y PAND2X1_592/CTRL 0.01fF
C5529 POR2X1_567/A PAND2X1_280/a_16_344# -0.02fF
C5530 POR2X1_616/Y PAND2X1_623/Y 0.03fF
C5531 POR2X1_549/CTRL PAND2X1_52/B 0.29fF
C5532 POR2X1_814/B PAND2X1_52/B 2.55fF
C5533 POR2X1_78/B POR2X1_711/Y 0.07fF
C5534 POR2X1_567/A PAND2X1_55/Y 0.08fF
C5535 POR2X1_68/A PAND2X1_48/A 0.03fF
C5536 POR2X1_383/A POR2X1_707/Y 1.57fF
C5537 PAND2X1_625/O POR2X1_294/A 0.17fF
C5538 PAND2X1_734/O PAND2X1_560/B 0.01fF
C5539 POR2X1_21/O POR2X1_260/A 0.01fF
C5540 PAND2X1_610/CTRL POR2X1_293/Y 0.01fF
C5541 PAND2X1_20/A PAND2X1_125/a_16_344# 0.01fF
C5542 POR2X1_302/A POR2X1_188/Y 0.50fF
C5543 POR2X1_83/A POR2X1_397/CTRL 0.01fF
C5544 POR2X1_343/Y POR2X1_723/CTRL2 0.00fF
C5545 POR2X1_829/A POR2X1_761/A 0.03fF
C5546 POR2X1_57/A POR2X1_129/Y 0.03fF
C5547 POR2X1_622/CTRL POR2X1_29/A 0.01fF
C5548 PAND2X1_227/O PAND2X1_340/B 0.01fF
C5549 POR2X1_73/Y PAND2X1_325/CTRL2 0.01fF
C5550 POR2X1_444/Y POR2X1_319/Y 0.06fF
C5551 POR2X1_48/A PAND2X1_206/B 0.07fF
C5552 POR2X1_341/Y POR2X1_339/Y 0.87fF
C5553 POR2X1_329/A POR2X1_37/Y 0.07fF
C5554 PAND2X1_652/CTRL PAND2X1_652/A 0.04fF
C5555 PAND2X1_849/B PAND2X1_100/CTRL 0.01fF
C5556 POR2X1_329/A PAND2X1_561/CTRL 0.01fF
C5557 POR2X1_540/A POR2X1_552/O 0.02fF
C5558 POR2X1_249/Y POR2X1_734/CTRL2 0.01fF
C5559 PAND2X1_413/CTRL POR2X1_814/A 0.01fF
C5560 POR2X1_190/CTRL2 POR2X1_188/Y 0.01fF
C5561 POR2X1_61/A PAND2X1_69/A 0.04fF
C5562 POR2X1_383/A PAND2X1_701/O 0.06fF
C5563 POR2X1_416/B POR2X1_481/a_16_28# 0.00fF
C5564 POR2X1_54/Y POR2X1_415/A 0.10fF
C5565 PAND2X1_476/A PAND2X1_734/CTRL 0.00fF
C5566 POR2X1_333/Y POR2X1_351/CTRL 0.30fF
C5567 POR2X1_57/A PAND2X1_659/Y 0.06fF
C5568 POR2X1_814/B PAND2X1_125/a_16_344# 0.02fF
C5569 POR2X1_102/Y POR2X1_498/m4_208_n4# 0.12fF
C5570 POR2X1_66/B POR2X1_98/A 0.41fF
C5571 POR2X1_130/A POR2X1_343/B 0.32fF
C5572 POR2X1_246/CTRL POR2X1_39/B 0.01fF
C5573 POR2X1_540/Y POR2X1_573/A 0.02fF
C5574 PAND2X1_109/O POR2X1_775/A 0.03fF
C5575 POR2X1_709/B POR2X1_710/B 0.03fF
C5576 POR2X1_316/Y PAND2X1_457/CTRL 0.01fF
C5577 POR2X1_334/Y POR2X1_101/Y 0.04fF
C5578 POR2X1_110/Y PAND2X1_549/B 0.06fF
C5579 POR2X1_99/B POR2X1_228/Y 0.02fF
C5580 POR2X1_411/B POR2X1_409/B 0.07fF
C5581 PAND2X1_440/O PAND2X1_652/A 0.05fF
C5582 POR2X1_432/CTRL2 POR2X1_271/B 0.01fF
C5583 PAND2X1_357/Y POR2X1_77/Y 0.03fF
C5584 POR2X1_802/a_16_28# POR2X1_802/A 0.03fF
C5585 POR2X1_503/a_16_28# POR2X1_411/B 0.02fF
C5586 POR2X1_741/B POR2X1_741/A 0.01fF
C5587 POR2X1_13/A PAND2X1_860/A 0.03fF
C5588 D_GATE_662 POR2X1_356/Y 0.04fF
C5589 POR2X1_814/A POR2X1_862/B 0.05fF
C5590 POR2X1_467/CTRL2 PAND2X1_52/B 0.01fF
C5591 PAND2X1_301/CTRL PAND2X1_716/B 0.01fF
C5592 POR2X1_23/Y POR2X1_265/CTRL 0.01fF
C5593 POR2X1_715/A POR2X1_186/B 0.03fF
C5594 POR2X1_48/A PAND2X1_606/O 0.06fF
C5595 POR2X1_750/O POR2X1_39/B 0.01fF
C5596 POR2X1_505/CTRL2 PAND2X1_631/A 0.01fF
C5597 PAND2X1_213/Y PAND2X1_169/a_16_344# 0.01fF
C5598 PAND2X1_737/B PAND2X1_737/O 0.06fF
C5599 POR2X1_435/O PAND2X1_72/A 0.01fF
C5600 POR2X1_16/A POR2X1_767/a_16_28# 0.03fF
C5601 POR2X1_278/A POR2X1_77/Y 0.18fF
C5602 POR2X1_12/A POR2X1_32/A 0.07fF
C5603 POR2X1_825/Y POR2X1_42/Y 0.13fF
C5604 PAND2X1_663/a_76_28# PAND2X1_659/Y 0.01fF
C5605 PAND2X1_295/a_76_28# POR2X1_294/Y 0.04fF
C5606 POR2X1_738/A POR2X1_568/B 0.05fF
C5607 PAND2X1_140/A POR2X1_77/Y 0.01fF
C5608 PAND2X1_458/CTRL2 POR2X1_372/Y 0.01fF
C5609 POR2X1_337/Y POR2X1_186/B 0.07fF
C5610 POR2X1_257/A PAND2X1_478/B 0.01fF
C5611 POR2X1_356/m4_208_n4# POR2X1_356/B 0.14fF
C5612 POR2X1_11/CTRL INPUT_7 0.01fF
C5613 POR2X1_406/Y POR2X1_329/A 0.43fF
C5614 PAND2X1_439/CTRL PAND2X1_738/Y 0.13fF
C5615 POR2X1_760/A PAND2X1_473/B 0.05fF
C5616 PAND2X1_290/O PAND2X1_94/A 0.17fF
C5617 PAND2X1_856/O PAND2X1_863/A 0.01fF
C5618 PAND2X1_798/Y PAND2X1_356/a_76_28# 0.03fF
C5619 POR2X1_106/CTRL POR2X1_48/A 0.01fF
C5620 PAND2X1_419/CTRL2 POR2X1_296/B 0.00fF
C5621 PAND2X1_267/CTRL POR2X1_102/Y 0.01fF
C5622 POR2X1_662/a_16_28# POR2X1_661/Y 0.02fF
C5623 POR2X1_490/Y POR2X1_60/A 0.03fF
C5624 POR2X1_624/B VDD 0.77fF
C5625 PAND2X1_467/Y POR2X1_158/Y 0.03fF
C5626 PAND2X1_499/O POR2X1_20/B 0.00fF
C5627 POR2X1_420/CTRL2 POR2X1_102/Y 0.01fF
C5628 POR2X1_260/B POR2X1_643/A 0.00fF
C5629 POR2X1_329/A POR2X1_293/Y 0.14fF
C5630 PAND2X1_613/CTRL2 PAND2X1_41/B 0.01fF
C5631 POR2X1_96/O POR2X1_77/Y 0.17fF
C5632 PAND2X1_94/A POR2X1_124/CTRL2 0.16fF
C5633 POR2X1_88/A VDD -0.00fF
C5634 POR2X1_411/B POR2X1_272/Y 0.15fF
C5635 PAND2X1_560/B POR2X1_39/B 0.12fF
C5636 POR2X1_431/Y VDD 0.04fF
C5637 POR2X1_115/O POR2X1_554/B 0.01fF
C5638 POR2X1_860/CTRL PAND2X1_72/A 0.01fF
C5639 POR2X1_257/A PAND2X1_210/O 0.15fF
C5640 POR2X1_11/CTRL INPUT_4 0.01fF
C5641 PAND2X1_205/A POR2X1_72/B 0.03fF
C5642 POR2X1_83/B PAND2X1_220/A 0.00fF
C5643 POR2X1_119/Y POR2X1_150/a_16_28# 0.09fF
C5644 PAND2X1_827/CTRL POR2X1_355/A 0.01fF
C5645 POR2X1_24/CTRL2 POR2X1_409/B 0.03fF
C5646 POR2X1_567/A POR2X1_741/O 0.01fF
C5647 POR2X1_192/B POR2X1_169/A 2.51fF
C5648 POR2X1_78/B PAND2X1_601/CTRL 0.04fF
C5649 POR2X1_485/Y POR2X1_763/Y 0.08fF
C5650 PAND2X1_689/a_56_28# POR2X1_121/B 0.00fF
C5651 PAND2X1_486/CTRL POR2X1_484/Y 0.01fF
C5652 POR2X1_48/A PAND2X1_220/Y 0.03fF
C5653 PAND2X1_357/a_76_28# POR2X1_39/B 0.02fF
C5654 D_INPUT_7 D_INPUT_6 0.10fF
C5655 POR2X1_69/Y D_INPUT_1 0.03fF
C5656 POR2X1_294/A POR2X1_711/Y 0.03fF
C5657 POR2X1_35/B POR2X1_34/B 0.00fF
C5658 POR2X1_517/a_16_28# PAND2X1_404/Y 0.02fF
C5659 POR2X1_669/B POR2X1_40/Y 3.71fF
C5660 PAND2X1_586/CTRL PAND2X1_72/A 0.01fF
C5661 POR2X1_150/Y PAND2X1_724/B 0.03fF
C5662 PAND2X1_23/Y POR2X1_116/A 0.03fF
C5663 POR2X1_66/B POR2X1_267/O 0.01fF
C5664 PAND2X1_624/A POR2X1_20/B 0.06fF
C5665 PAND2X1_859/O POR2X1_37/Y 0.13fF
C5666 POR2X1_188/A POR2X1_858/a_76_344# 0.00fF
C5667 POR2X1_566/A POR2X1_445/A 0.12fF
C5668 POR2X1_536/Y POR2X1_102/Y 0.04fF
C5669 PAND2X1_464/B PAND2X1_785/CTRL2 0.03fF
C5670 PAND2X1_420/CTRL POR2X1_630/A 0.02fF
C5671 POR2X1_814/B POR2X1_288/CTRL 0.03fF
C5672 POR2X1_496/CTRL POR2X1_55/Y 0.01fF
C5673 PAND2X1_48/B POR2X1_472/B 0.07fF
C5674 PAND2X1_41/B PAND2X1_531/O 0.02fF
C5675 PAND2X1_793/Y POR2X1_437/CTRL 0.01fF
C5676 PAND2X1_793/CTRL2 POR2X1_29/A 0.01fF
C5677 POR2X1_43/B POR2X1_20/B 1.64fF
C5678 POR2X1_287/B POR2X1_590/A 0.10fF
C5679 POR2X1_801/A POR2X1_801/B 0.30fF
C5680 PAND2X1_645/O POR2X1_48/A 0.15fF
C5681 POR2X1_312/O POR2X1_20/B 0.17fF
C5682 PAND2X1_48/A POR2X1_138/A 0.03fF
C5683 POR2X1_428/Y POR2X1_700/O 0.02fF
C5684 POR2X1_814/A POR2X1_510/Y 0.07fF
C5685 POR2X1_49/Y PAND2X1_478/B 0.09fF
C5686 PAND2X1_52/B PAND2X1_680/O 0.06fF
C5687 POR2X1_274/A PAND2X1_131/m4_208_n4# 0.07fF
C5688 PAND2X1_630/O POR2X1_628/Y 0.01fF
C5689 POR2X1_568/B POR2X1_568/O 0.06fF
C5690 POR2X1_485/Y POR2X1_73/Y 0.98fF
C5691 POR2X1_138/CTRL2 POR2X1_260/B 0.01fF
C5692 POR2X1_458/O POR2X1_784/A 0.03fF
C5693 PAND2X1_48/B POR2X1_866/A 0.03fF
C5694 POR2X1_210/CTRL VDD 0.00fF
C5695 PAND2X1_605/a_76_28# INPUT_0 0.02fF
C5696 PAND2X1_221/O PAND2X1_192/Y 0.03fF
C5697 PAND2X1_221/a_16_344# PAND2X1_220/Y 0.04fF
C5698 POR2X1_383/A PAND2X1_52/O 0.01fF
C5699 PAND2X1_838/CTRL POR2X1_73/Y 0.04fF
C5700 POR2X1_624/Y POR2X1_501/a_76_344# 0.01fF
C5701 POR2X1_20/B POR2X1_38/B 0.03fF
C5702 POR2X1_820/Y POR2X1_32/A 0.03fF
C5703 POR2X1_590/A PAND2X1_8/Y 0.23fF
C5704 POR2X1_14/Y POR2X1_236/Y 3.20fF
C5705 POR2X1_123/B POR2X1_556/A 0.02fF
C5706 PAND2X1_39/B PAND2X1_743/O 0.05fF
C5707 POR2X1_814/A POR2X1_276/Y 0.03fF
C5708 PAND2X1_96/B POR2X1_649/a_16_28# 0.01fF
C5709 D_INPUT_0 POR2X1_522/a_76_344# 0.02fF
C5710 POR2X1_102/Y PAND2X1_730/B 0.02fF
C5711 POR2X1_140/B POR2X1_260/B 0.02fF
C5712 POR2X1_78/A POR2X1_192/Y 0.03fF
C5713 PAND2X1_73/Y POR2X1_220/Y 0.06fF
C5714 PAND2X1_721/B PAND2X1_673/Y 0.01fF
C5715 POR2X1_812/CTRL2 POR2X1_121/B 0.03fF
C5716 POR2X1_814/A POR2X1_768/CTRL2 0.08fF
C5717 POR2X1_407/A POR2X1_260/B 0.10fF
C5718 POR2X1_428/Y PAND2X1_711/CTRL 0.09fF
C5719 PAND2X1_48/B POR2X1_269/CTRL2 0.01fF
C5720 PAND2X1_735/Y PAND2X1_573/B 0.25fF
C5721 POR2X1_642/O POR2X1_66/A 0.01fF
C5722 PAND2X1_717/A PAND2X1_579/A 0.00fF
C5723 PAND2X1_6/Y PAND2X1_258/CTRL2 0.00fF
C5724 PAND2X1_221/O PAND2X1_738/Y 0.04fF
C5725 POR2X1_254/Y POR2X1_66/B 0.07fF
C5726 PAND2X1_73/Y POR2X1_404/Y 0.40fF
C5727 POR2X1_21/CTRL D_INPUT_5 0.01fF
C5728 POR2X1_850/O PAND2X1_39/B 0.05fF
C5729 POR2X1_36/B POR2X1_582/Y 0.01fF
C5730 POR2X1_66/A POR2X1_341/CTRL 0.06fF
C5731 PAND2X1_217/CTRL PAND2X1_656/A 0.01fF
C5732 POR2X1_3/A POR2X1_428/Y 0.04fF
C5733 POR2X1_41/B POR2X1_667/A 0.00fF
C5734 POR2X1_296/B POR2X1_55/Y 0.00fF
C5735 PAND2X1_339/O PAND2X1_332/Y -0.00fF
C5736 POR2X1_405/O VDD 0.00fF
C5737 PAND2X1_631/CTRL POR2X1_48/A 0.01fF
C5738 PAND2X1_116/O POR2X1_106/Y 0.02fF
C5739 POR2X1_452/Y POR2X1_729/Y 1.23fF
C5740 POR2X1_459/CTRL POR2X1_750/B 0.01fF
C5741 POR2X1_435/a_16_28# POR2X1_796/A 0.03fF
C5742 POR2X1_366/Y POR2X1_174/A 0.07fF
C5743 POR2X1_567/B POR2X1_340/m4_208_n4# 0.06fF
C5744 POR2X1_28/O D_INPUT_1 0.01fF
C5745 PAND2X1_58/A POR2X1_791/CTRL 0.01fF
C5746 PAND2X1_575/A POR2X1_32/A 0.05fF
C5747 D_INPUT_0 POR2X1_723/B 0.03fF
C5748 POR2X1_52/A POR2X1_847/A 0.01fF
C5749 POR2X1_62/O POR2X1_29/A 0.04fF
C5750 PAND2X1_787/CTRL VDD -0.00fF
C5751 PAND2X1_462/B POR2X1_102/Y 0.21fF
C5752 POR2X1_226/CTRL POR2X1_42/Y 0.03fF
C5753 PAND2X1_403/B POR2X1_290/Y 0.23fF
C5754 POR2X1_356/A POR2X1_436/CTRL2 0.04fF
C5755 PAND2X1_84/CTRL POR2X1_5/Y 0.01fF
C5756 POR2X1_610/a_16_28# PAND2X1_69/A 0.03fF
C5757 PAND2X1_159/a_16_344# POR2X1_7/B 0.02fF
C5758 PAND2X1_20/A PAND2X1_95/B 0.06fF
C5759 PAND2X1_848/B POR2X1_669/B 0.18fF
C5760 POR2X1_65/A POR2X1_516/B 0.03fF
C5761 POR2X1_66/A POR2X1_194/CTRL2 0.01fF
C5762 PAND2X1_90/A PAND2X1_73/CTRL2 0.03fF
C5763 POR2X1_23/Y PAND2X1_575/O 0.01fF
C5764 POR2X1_96/A PAND2X1_78/a_76_28# 0.01fF
C5765 POR2X1_696/Y VDD 0.00fF
C5766 POR2X1_62/Y PAND2X1_206/B 0.10fF
C5767 PAND2X1_700/O PAND2X1_90/Y 0.06fF
C5768 PAND2X1_23/Y POR2X1_638/A 0.01fF
C5769 PAND2X1_96/B POR2X1_479/B 1.16fF
C5770 PAND2X1_685/O POR2X1_60/A 0.03fF
C5771 PAND2X1_740/O PAND2X1_738/Y 0.04fF
C5772 PAND2X1_58/A POR2X1_565/CTRL 0.01fF
C5773 POR2X1_301/O POR2X1_590/A 0.01fF
C5774 POR2X1_590/A POR2X1_705/CTRL2 0.01fF
C5775 POR2X1_594/Y PAND2X1_557/A 0.16fF
C5776 PAND2X1_55/Y POR2X1_643/A 0.01fF
C5777 PAND2X1_787/Y PAND2X1_139/Y 0.02fF
C5778 PAND2X1_23/Y POR2X1_242/CTRL 0.01fF
C5779 POR2X1_76/O POR2X1_553/A 0.08fF
C5780 POR2X1_493/CTRL POR2X1_558/B 0.00fF
C5781 POR2X1_493/O POR2X1_493/A 0.01fF
C5782 PAND2X1_793/Y PAND2X1_579/O 0.02fF
C5783 PAND2X1_96/B PAND2X1_595/O 0.02fF
C5784 POR2X1_25/a_16_28# INPUT_7 0.03fF
C5785 PAND2X1_267/Y PAND2X1_656/A 0.02fF
C5786 POR2X1_57/A POR2X1_37/Y 0.17fF
C5787 POR2X1_17/O INPUT_5 0.02fF
C5788 POR2X1_346/B POR2X1_66/Y 0.00fF
C5789 POR2X1_174/B POR2X1_351/Y 0.03fF
C5790 POR2X1_83/B PAND2X1_337/A 0.00fF
C5791 POR2X1_662/Y POR2X1_750/B 0.03fF
C5792 PAND2X1_23/Y POR2X1_94/A 0.00fF
C5793 PAND2X1_54/O INPUT_0 0.15fF
C5794 POR2X1_178/CTRL POR2X1_60/A 0.01fF
C5795 POR2X1_7/B POR2X1_595/Y 0.00fF
C5796 PAND2X1_96/B POR2X1_792/O 0.01fF
C5797 POR2X1_664/Y PAND2X1_41/B 0.03fF
C5798 PAND2X1_16/CTRL POR2X1_294/B 0.00fF
C5799 PAND2X1_341/B POR2X1_65/CTRL 0.01fF
C5800 POR2X1_383/A POR2X1_647/a_16_28# 0.03fF
C5801 POR2X1_605/A POR2X1_78/A 0.00fF
C5802 PAND2X1_288/A PAND2X1_805/A 3.60fF
C5803 PAND2X1_90/A POR2X1_392/B 0.35fF
C5804 POR2X1_596/Y VDD 0.13fF
C5805 D_INPUT_0 PAND2X1_338/B 0.03fF
C5806 POR2X1_16/A PAND2X1_340/B 0.00fF
C5807 POR2X1_41/B PAND2X1_712/B 0.02fF
C5808 POR2X1_573/CTRL2 POR2X1_404/Y 0.04fF
C5809 POR2X1_186/Y POR2X1_563/Y 0.03fF
C5810 POR2X1_57/A POR2X1_279/CTRL 0.01fF
C5811 PAND2X1_472/B POR2X1_236/Y 0.10fF
C5812 PAND2X1_65/B POR2X1_578/Y 0.03fF
C5813 POR2X1_48/A PAND2X1_713/A 0.01fF
C5814 POR2X1_807/A PAND2X1_55/Y 0.05fF
C5815 POR2X1_775/A PAND2X1_41/B 0.03fF
C5816 PAND2X1_225/CTRL D_INPUT_1 0.01fF
C5817 POR2X1_274/CTRL2 POR2X1_569/A 0.03fF
C5818 PAND2X1_57/B INPUT_0 7.02fF
C5819 POR2X1_646/Y PAND2X1_60/B 0.17fF
C5820 POR2X1_322/Y POR2X1_32/A 0.02fF
C5821 POR2X1_114/Y POR2X1_130/A 0.02fF
C5822 POR2X1_537/CTRL POR2X1_260/B 0.01fF
C5823 POR2X1_502/A PAND2X1_587/Y 0.01fF
C5824 PAND2X1_90/Y PAND2X1_145/CTRL2 0.01fF
C5825 POR2X1_346/B POR2X1_629/O 0.00fF
C5826 POR2X1_356/A POR2X1_781/CTRL 0.04fF
C5827 POR2X1_13/CTRL2 POR2X1_7/B 0.01fF
C5828 POR2X1_164/O POR2X1_72/B 0.01fF
C5829 PAND2X1_786/CTRL2 POR2X1_91/Y 0.02fF
C5830 POR2X1_443/m4_208_n4# POR2X1_545/m4_208_n4# 0.13fF
C5831 POR2X1_163/A VDD 0.00fF
C5832 POR2X1_55/Y POR2X1_236/Y 0.15fF
C5833 POR2X1_62/Y POR2X1_65/Y 0.00fF
C5834 PAND2X1_673/O POR2X1_670/Y 0.02fF
C5835 PAND2X1_20/A POR2X1_350/B 0.02fF
C5836 POR2X1_68/A POR2X1_193/Y 0.03fF
C5837 POR2X1_78/B POR2X1_733/A 0.03fF
C5838 POR2X1_405/O PAND2X1_32/B 0.01fF
C5839 POR2X1_66/B PAND2X1_697/m4_208_n4# 0.20fF
C5840 POR2X1_502/A POR2X1_853/O 0.02fF
C5841 D_INPUT_0 POR2X1_576/CTRL 0.01fF
C5842 POR2X1_96/A PAND2X1_793/Y 0.06fF
C5843 PAND2X1_126/O POR2X1_29/A 0.00fF
C5844 PAND2X1_377/CTRL2 POR2X1_42/Y 0.01fF
C5845 POR2X1_78/B POR2X1_334/B 0.12fF
C5846 POR2X1_13/A POR2X1_684/CTRL 0.01fF
C5847 POR2X1_504/Y PAND2X1_631/O 0.02fF
C5848 POR2X1_669/B PAND2X1_559/O 0.15fF
C5849 POR2X1_640/A POR2X1_391/Y 0.00fF
C5850 POR2X1_83/B PAND2X1_349/A 0.03fF
C5851 POR2X1_748/A INPUT_6 0.06fF
C5852 POR2X1_83/B PAND2X1_63/B 0.03fF
C5853 PAND2X1_865/CTRL2 POR2X1_102/Y 0.01fF
C5854 PAND2X1_857/A POR2X1_60/A 0.03fF
C5855 POR2X1_712/A PAND2X1_65/B 0.04fF
C5856 POR2X1_196/Y POR2X1_61/Y 0.02fF
C5857 PAND2X1_652/A PAND2X1_192/a_76_28# 0.01fF
C5858 POR2X1_750/B POR2X1_194/a_16_28# 0.10fF
C5859 POR2X1_62/Y POR2X1_88/O 0.01fF
C5860 POR2X1_415/A POR2X1_4/Y 0.06fF
C5861 POR2X1_48/A PAND2X1_560/B 0.03fF
C5862 POR2X1_557/A PAND2X1_73/Y 0.07fF
C5863 PAND2X1_91/CTRL2 POR2X1_192/B 0.07fF
C5864 POR2X1_316/Y PAND2X1_464/CTRL 0.01fF
C5865 PAND2X1_536/O VDD 0.00fF
C5866 POR2X1_111/CTRL2 POR2X1_5/Y 0.01fF
C5867 POR2X1_407/Y PAND2X1_597/a_16_344# 0.01fF
C5868 POR2X1_834/Y PAND2X1_591/m4_208_n4# 0.04fF
C5869 POR2X1_119/Y PAND2X1_444/CTRL2 0.00fF
C5870 POR2X1_408/O INPUT_5 0.18fF
C5871 POR2X1_783/CTRL2 POR2X1_796/A 0.01fF
C5872 POR2X1_107/O POR2X1_90/Y 0.04fF
C5873 PAND2X1_258/O POR2X1_186/B 0.04fF
C5874 PAND2X1_855/O POR2X1_236/Y 0.04fF
C5875 PAND2X1_460/CTRL POR2X1_5/Y 0.01fF
C5876 PAND2X1_6/Y VDD 2.87fF
C5877 POR2X1_41/B PAND2X1_852/CTRL 0.01fF
C5878 POR2X1_16/A POR2X1_102/Y 1.59fF
C5879 PAND2X1_118/O POR2X1_502/A 0.02fF
C5880 POR2X1_140/B PAND2X1_516/CTRL 0.00fF
C5881 POR2X1_510/A POR2X1_192/Y 0.05fF
C5882 POR2X1_266/A POR2X1_266/a_16_28# 0.03fF
C5883 POR2X1_283/m4_208_n4# PAND2X1_356/m4_208_n4# 0.13fF
C5884 POR2X1_99/B POR2X1_454/A 0.01fF
C5885 PAND2X1_818/m4_208_n4# POR2X1_42/Y 0.06fF
C5886 PAND2X1_484/CTRL2 POR2X1_590/A 0.01fF
C5887 PAND2X1_48/B PAND2X1_280/a_76_28# 0.01fF
C5888 PAND2X1_471/O PAND2X1_464/Y 0.01fF
C5889 PAND2X1_63/Y POR2X1_130/A 0.10fF
C5890 POR2X1_416/B PAND2X1_634/CTRL 0.01fF
C5891 POR2X1_383/A POR2X1_343/A 0.06fF
C5892 POR2X1_832/Y POR2X1_512/a_76_344# 0.01fF
C5893 POR2X1_41/B PAND2X1_546/CTRL2 0.01fF
C5894 POR2X1_466/A POR2X1_552/CTRL 0.01fF
C5895 POR2X1_706/B POR2X1_713/B 0.01fF
C5896 POR2X1_634/A POR2X1_260/A 2.02fF
C5897 POR2X1_333/A POR2X1_444/Y 0.05fF
C5898 PAND2X1_96/B POR2X1_194/B 0.06fF
C5899 PAND2X1_499/CTRL POR2X1_283/A 0.01fF
C5900 POR2X1_532/A PAND2X1_131/CTRL 0.01fF
C5901 POR2X1_178/Y PAND2X1_540/O 0.02fF
C5902 PAND2X1_674/CTRL POR2X1_732/B 0.11fF
C5903 PAND2X1_543/O POR2X1_142/Y 0.09fF
C5904 POR2X1_845/O POR2X1_5/Y 0.00fF
C5905 D_INPUT_3 VDD 3.25fF
C5906 POR2X1_128/O PAND2X1_96/B 0.01fF
C5907 POR2X1_52/A POR2X1_93/O 0.02fF
C5908 POR2X1_475/A POR2X1_101/Y 0.04fF
C5909 POR2X1_407/A PAND2X1_55/Y 0.19fF
C5910 POR2X1_186/Y POR2X1_675/Y 0.03fF
C5911 POR2X1_113/Y POR2X1_130/A 0.10fF
C5912 PAND2X1_575/A POR2X1_184/Y 0.00fF
C5913 POR2X1_66/A PAND2X1_179/CTRL2 0.03fF
C5914 PAND2X1_472/A POR2X1_42/Y 0.03fF
C5915 PAND2X1_735/Y POR2X1_91/Y 0.07fF
C5916 POR2X1_850/A POR2X1_249/Y 0.02fF
C5917 POR2X1_795/CTRL2 PAND2X1_32/B 0.03fF
C5918 PAND2X1_349/A PAND2X1_140/Y 0.01fF
C5919 PAND2X1_65/B POR2X1_598/CTRL 0.01fF
C5920 POR2X1_729/CTRL2 POR2X1_614/A 0.03fF
C5921 POR2X1_323/O POR2X1_164/Y 0.07fF
C5922 POR2X1_829/A POR2X1_761/Y 0.00fF
C5923 POR2X1_197/Y POR2X1_244/B 0.06fF
C5924 PAND2X1_65/B POR2X1_407/O 0.01fF
C5925 PAND2X1_252/CTRL2 PAND2X1_55/Y 0.01fF
C5926 PAND2X1_661/Y PAND2X1_688/O 0.01fF
C5927 PAND2X1_58/A PAND2X1_48/A 0.11fF
C5928 POR2X1_856/B PAND2X1_167/a_16_344# 0.06fF
C5929 PAND2X1_382/O VDD 0.00fF
C5930 POR2X1_42/Y POR2X1_396/a_16_28# 0.02fF
C5931 PAND2X1_48/B POR2X1_501/B 0.12fF
C5932 INPUT_0 PAND2X1_549/B 0.14fF
C5933 POR2X1_614/A POR2X1_264/Y 0.03fF
C5934 POR2X1_447/CTRL2 POR2X1_294/B 0.01fF
C5935 PAND2X1_803/A PAND2X1_727/CTRL 0.00fF
C5936 PAND2X1_6/Y POR2X1_741/Y 0.07fF
C5937 POR2X1_57/A POR2X1_293/Y 3.94fF
C5938 POR2X1_32/Y POR2X1_42/Y 0.01fF
C5939 PAND2X1_862/B PAND2X1_175/B 0.03fF
C5940 POR2X1_186/Y POR2X1_544/B 0.07fF
C5941 PAND2X1_371/a_16_344# POR2X1_68/B 0.01fF
C5942 POR2X1_327/Y POR2X1_777/B 0.03fF
C5943 POR2X1_102/Y PAND2X1_336/Y 0.00fF
C5944 POR2X1_220/Y PAND2X1_163/O 0.00fF
C5945 POR2X1_222/Y POR2X1_194/CTRL2 0.03fF
C5946 POR2X1_55/Y PAND2X1_344/CTRL 0.01fF
C5947 POR2X1_114/B POR2X1_778/B 0.02fF
C5948 D_GATE_222 PAND2X1_69/A 0.06fF
C5949 POR2X1_41/B POR2X1_245/Y 0.07fF
C5950 PAND2X1_63/Y POR2X1_204/CTRL 0.01fF
C5951 POR2X1_502/A PAND2X1_373/CTRL2 0.01fF
C5952 VDD POR2X1_7/CTRL 0.00fF
C5953 PAND2X1_470/CTRL POR2X1_43/B 0.01fF
C5954 POR2X1_543/A POR2X1_186/B 0.03fF
C5955 VDD POR2X1_569/Y 0.10fF
C5956 POR2X1_196/Y POR2X1_35/Y 0.02fF
C5957 POR2X1_62/Y POR2X1_750/B 11.37fF
C5958 PAND2X1_339/Y POR2X1_73/Y 0.07fF
C5959 POR2X1_138/m4_208_n4# PAND2X1_32/B 0.08fF
C5960 POR2X1_390/B POR2X1_723/CTRL 0.00fF
C5961 POR2X1_157/O POR2X1_36/B 0.01fF
C5962 PAND2X1_857/O POR2X1_83/B 0.05fF
C5963 POR2X1_507/B POR2X1_355/A 0.01fF
C5964 PAND2X1_105/a_16_344# POR2X1_90/Y 0.01fF
C5965 POR2X1_635/B PAND2X1_47/O 0.00fF
C5966 POR2X1_188/A POR2X1_711/B 0.02fF
C5967 POR2X1_229/Y POR2X1_293/Y 0.05fF
C5968 POR2X1_394/A POR2X1_5/Y 0.12fF
C5969 PAND2X1_6/Y PAND2X1_32/B 0.31fF
C5970 POR2X1_407/A POR2X1_407/Y 0.03fF
C5971 POR2X1_130/A POR2X1_260/A 0.08fF
C5972 POR2X1_141/O POR2X1_574/Y 0.00fF
C5973 POR2X1_149/B POR2X1_532/A 0.01fF
C5974 POR2X1_327/Y PAND2X1_65/B 0.10fF
C5975 PAND2X1_4/CTRL2 PAND2X1_6/A 0.01fF
C5976 POR2X1_816/A POR2X1_498/A 0.01fF
C5977 POR2X1_559/Y POR2X1_532/A 0.01fF
C5978 POR2X1_840/B POR2X1_786/Y 0.03fF
C5979 PAND2X1_209/CTRL2 POR2X1_394/A 0.01fF
C5980 PAND2X1_115/O POR2X1_283/A 0.05fF
C5981 POR2X1_329/a_16_28# POR2X1_283/A 0.01fF
C5982 POR2X1_502/A PAND2X1_376/O 0.03fF
C5983 POR2X1_566/A POR2X1_260/A 0.05fF
C5984 POR2X1_865/B POR2X1_114/O 0.01fF
C5985 POR2X1_778/B POR2X1_458/B 0.01fF
C5986 POR2X1_49/Y PAND2X1_341/B 0.03fF
C5987 POR2X1_316/CTRL2 INPUT_0 0.09fF
C5988 POR2X1_782/A PAND2X1_747/O 0.01fF
C5989 POR2X1_139/a_16_28# PAND2X1_32/B 0.01fF
C5990 PAND2X1_777/a_76_28# POR2X1_39/B 0.01fF
C5991 POR2X1_532/A POR2X1_219/CTRL 0.01fF
C5992 PAND2X1_216/B POR2X1_79/Y 0.03fF
C5993 PAND2X1_23/Y POR2X1_710/Y 0.02fF
C5994 POR2X1_416/B PAND2X1_34/CTRL2 0.04fF
C5995 PAND2X1_649/A POR2X1_40/Y 0.00fF
C5996 POR2X1_68/A PAND2X1_670/O 0.15fF
C5997 POR2X1_13/A PAND2X1_301/a_16_344# 0.01fF
C5998 POR2X1_532/A POR2X1_644/A 0.03fF
C5999 POR2X1_93/CTRL D_INPUT_3 0.03fF
C6000 POR2X1_537/Y POR2X1_733/CTRL2 0.01fF
C6001 PAND2X1_635/O INPUT_6 0.01fF
C6002 POR2X1_242/m4_208_n4# POR2X1_192/B 0.04fF
C6003 POR2X1_447/B POR2X1_61/Y 0.06fF
C6004 PAND2X1_48/B POR2X1_703/A 0.03fF
C6005 PAND2X1_308/B POR2X1_153/Y 0.03fF
C6006 PAND2X1_57/B POR2X1_398/CTRL2 0.01fF
C6007 PAND2X1_731/B PAND2X1_326/B 0.02fF
C6008 PAND2X1_836/O POR2X1_823/Y -0.00fF
C6009 PAND2X1_726/B POR2X1_763/Y 2.24fF
C6010 POR2X1_804/A PAND2X1_60/B 0.03fF
C6011 POR2X1_548/O POR2X1_620/B 0.02fF
C6012 POR2X1_751/a_76_344# POR2X1_816/A 0.00fF
C6013 POR2X1_332/B POR2X1_186/B 0.10fF
C6014 PAND2X1_182/A PAND2X1_182/B 0.02fF
C6015 POR2X1_637/O PAND2X1_72/A 0.01fF
C6016 GATE_741 PAND2X1_354/Y 0.03fF
C6017 POR2X1_228/Y POR2X1_112/Y 0.35fF
C6018 PAND2X1_560/O POR2X1_73/Y 0.01fF
C6019 POR2X1_111/Y POR2X1_293/Y 0.02fF
C6020 POR2X1_667/A POR2X1_77/Y 0.04fF
C6021 POR2X1_73/CTRL PAND2X1_6/A 0.03fF
C6022 PAND2X1_565/O PAND2X1_550/Y 0.00fF
C6023 POR2X1_537/CTRL PAND2X1_55/Y 0.03fF
C6024 PAND2X1_808/Y POR2X1_16/A 0.03fF
C6025 POR2X1_367/O POR2X1_191/Y 0.08fF
C6026 POR2X1_101/Y POR2X1_218/A 0.11fF
C6027 POR2X1_13/A PAND2X1_156/A 0.03fF
C6028 PAND2X1_93/B POR2X1_76/B 0.03fF
C6029 PAND2X1_659/Y PAND2X1_84/Y 0.00fF
C6030 POR2X1_435/Y PAND2X1_48/A 0.07fF
C6031 POR2X1_366/Y POR2X1_704/Y 0.01fF
C6032 POR2X1_183/Y PAND2X1_114/CTRL 0.00fF
C6033 PAND2X1_838/B POR2X1_827/CTRL 0.01fF
C6034 PAND2X1_643/A PAND2X1_539/B 0.13fF
C6035 POR2X1_197/CTRL POR2X1_99/B 0.00fF
C6036 PAND2X1_863/B POR2X1_595/CTRL 0.01fF
C6037 POR2X1_204/CTRL POR2X1_260/A 0.00fF
C6038 POR2X1_83/Y VDD 0.52fF
C6039 POR2X1_271/A POR2X1_55/Y 0.17fF
C6040 POR2X1_208/A PAND2X1_291/CTRL2 0.00fF
C6041 POR2X1_43/B PAND2X1_715/B 0.03fF
C6042 PAND2X1_117/CTRL2 PAND2X1_48/A -0.00fF
C6043 PAND2X1_560/B PAND2X1_197/Y 0.03fF
C6044 POR2X1_778/B PAND2X1_103/O 0.02fF
C6045 PAND2X1_824/B D_GATE_222 0.07fF
C6046 POR2X1_720/A POR2X1_39/B 0.03fF
C6047 POR2X1_5/Y PAND2X1_198/CTRL2 0.01fF
C6048 POR2X1_119/Y PAND2X1_659/a_16_344# 0.04fF
C6049 PAND2X1_23/Y POR2X1_334/Y 0.07fF
C6050 POR2X1_383/A POR2X1_137/Y 0.03fF
C6051 POR2X1_40/Y PAND2X1_327/O 0.01fF
C6052 POR2X1_52/A POR2X1_150/CTRL 0.01fF
C6053 POR2X1_339/CTRL2 POR2X1_556/Y 0.00fF
C6054 POR2X1_359/a_16_28# POR2X1_349/Y 0.03fF
C6055 POR2X1_416/B POR2X1_250/A 6.37fF
C6056 PAND2X1_317/Y PAND2X1_703/O 0.01fF
C6057 POR2X1_720/B POR2X1_720/CTRL2 0.10fF
C6058 POR2X1_566/A POR2X1_181/CTRL2 0.16fF
C6059 POR2X1_707/O POR2X1_407/Y 0.01fF
C6060 POR2X1_81/A PAND2X1_659/B 0.03fF
C6061 POR2X1_16/A POR2X1_821/Y 0.02fF
C6062 POR2X1_7/B PAND2X1_506/Y 0.01fF
C6063 POR2X1_567/B PAND2X1_438/O 0.27fF
C6064 POR2X1_834/Y POR2X1_596/A 0.04fF
C6065 PAND2X1_73/Y POR2X1_651/Y 0.03fF
C6066 POR2X1_334/B POR2X1_294/A 0.50fF
C6067 POR2X1_508/A POR2X1_508/CTRL2 0.01fF
C6068 PAND2X1_150/O POR2X1_260/A 0.03fF
C6069 PAND2X1_352/CTRL2 POR2X1_55/Y 0.01fF
C6070 POR2X1_741/Y POR2X1_195/O 0.06fF
C6071 PAND2X1_673/CTRL POR2X1_416/B 0.01fF
C6072 PAND2X1_162/A PAND2X1_162/a_76_28# 0.07fF
C6073 POR2X1_275/A POR2X1_275/Y 0.09fF
C6074 POR2X1_188/CTRL2 POR2X1_675/Y 0.01fF
C6075 POR2X1_363/A POR2X1_363/a_16_28# 0.02fF
C6076 VDD POR2X1_632/Y 0.40fF
C6077 PAND2X1_6/Y POR2X1_228/CTRL 0.01fF
C6078 POR2X1_502/A POR2X1_568/B 0.03fF
C6079 POR2X1_406/Y PAND2X1_339/CTRL 0.04fF
C6080 PAND2X1_271/CTRL2 POR2X1_116/A 0.00fF
C6081 POR2X1_65/A POR2X1_167/Y 0.77fF
C6082 PAND2X1_650/O PAND2X1_641/Y 0.02fF
C6083 POR2X1_655/O POR2X1_646/Y 0.02fF
C6084 POR2X1_551/O POR2X1_854/B 0.34fF
C6085 POR2X1_725/Y POR2X1_151/O 0.03fF
C6086 POR2X1_71/CTRL POR2X1_91/Y 0.02fF
C6087 PAND2X1_665/O POR2X1_664/Y -0.00fF
C6088 POR2X1_124/B POR2X1_294/A 0.12fF
C6089 POR2X1_119/Y PAND2X1_716/O 0.08fF
C6090 POR2X1_760/A PAND2X1_218/B 0.03fF
C6091 POR2X1_383/A POR2X1_833/A 0.07fF
C6092 POR2X1_11/a_16_28# D_INPUT_5 0.05fF
C6093 POR2X1_411/B POR2X1_679/A 0.08fF
C6094 PAND2X1_96/B PAND2X1_48/A 0.25fF
C6095 POR2X1_239/Y POR2X1_153/Y 0.05fF
C6096 POR2X1_709/m4_208_n4# POR2X1_713/B 0.06fF
C6097 VDD PAND2X1_52/B 7.78fF
C6098 PAND2X1_23/Y POR2X1_343/CTRL 0.03fF
C6099 PAND2X1_20/A PAND2X1_19/Y 0.01fF
C6100 VDD POR2X1_212/B 0.08fF
C6101 VDD POR2X1_759/O 0.00fF
C6102 POR2X1_188/A POR2X1_643/CTRL2 0.01fF
C6103 PAND2X1_163/CTRL POR2X1_210/A 0.01fF
C6104 POR2X1_9/Y POR2X1_69/A 0.03fF
C6105 POR2X1_416/B POR2X1_290/Y 4.83fF
C6106 POR2X1_343/Y POR2X1_579/Y 0.05fF
C6107 POR2X1_630/B POR2X1_590/A 0.02fF
C6108 POR2X1_274/A POR2X1_276/B 0.00fF
C6109 POR2X1_16/A PAND2X1_317/CTRL 0.01fF
C6110 POR2X1_157/CTRL POR2X1_416/B 0.01fF
C6111 POR2X1_96/A PAND2X1_862/O 0.01fF
C6112 PAND2X1_372/CTRL POR2X1_717/B 0.01fF
C6113 POR2X1_654/B POR2X1_643/O 0.03fF
C6114 POR2X1_661/O POR2X1_661/A 0.04fF
C6115 POR2X1_343/Y POR2X1_572/B 0.05fF
C6116 PAND2X1_175/B PAND2X1_716/B 0.03fF
C6117 POR2X1_60/A POR2X1_329/A 0.17fF
C6118 PAND2X1_838/a_76_28# POR2X1_827/Y 0.07fF
C6119 PAND2X1_270/a_76_28# PAND2X1_508/Y 0.01fF
C6120 POR2X1_864/CTRL POR2X1_814/A 0.28fF
C6121 POR2X1_416/B POR2X1_238/Y 0.03fF
C6122 POR2X1_156/CTRL POR2X1_162/Y 0.01fF
C6123 POR2X1_624/Y POR2X1_499/CTRL 0.01fF
C6124 POR2X1_20/B POR2X1_298/Y 0.01fF
C6125 POR2X1_632/Y PAND2X1_32/B 0.03fF
C6126 PAND2X1_481/O POR2X1_507/A 0.02fF
C6127 POR2X1_493/B PAND2X1_48/A 0.00fF
C6128 POR2X1_614/A POR2X1_343/Y 0.05fF
C6129 POR2X1_394/A POR2X1_599/CTRL 0.11fF
C6130 PAND2X1_94/CTRL POR2X1_202/A 0.03fF
C6131 POR2X1_508/B PAND2X1_823/CTRL2 0.00fF
C6132 POR2X1_833/A PAND2X1_71/Y 0.03fF
C6133 POR2X1_344/Y POR2X1_363/A 0.07fF
C6134 PAND2X1_641/CTRL PAND2X1_341/B 0.02fF
C6135 POR2X1_359/B POR2X1_244/Y 0.01fF
C6136 POR2X1_112/a_76_344# POR2X1_510/Y 0.00fF
C6137 POR2X1_456/B POR2X1_564/O 0.02fF
C6138 POR2X1_43/Y POR2X1_43/B 0.16fF
C6139 POR2X1_600/Y POR2X1_601/CTRL 0.03fF
C6140 PAND2X1_469/B POR2X1_173/a_56_344# 0.00fF
C6141 PAND2X1_212/CTRL PAND2X1_352/A 0.01fF
C6142 POR2X1_389/A POR2X1_711/Y 0.15fF
C6143 POR2X1_622/A POR2X1_29/A 0.00fF
C6144 PAND2X1_52/B PAND2X1_32/B 0.27fF
C6145 POR2X1_62/Y PAND2X1_560/B 1.42fF
C6146 POR2X1_60/A POR2X1_813/O 0.01fF
C6147 PAND2X1_459/CTRL PAND2X1_9/Y 0.01fF
C6148 POR2X1_14/Y POR2X1_24/Y 0.95fF
C6149 POR2X1_245/Y POR2X1_77/Y 0.05fF
C6150 POR2X1_48/A PAND2X1_400/CTRL2 0.02fF
C6151 POR2X1_610/Y POR2X1_634/A 0.01fF
C6152 POR2X1_567/A POR2X1_339/m4_208_n4# 0.03fF
C6153 POR2X1_527/CTRL2 POR2X1_39/B 0.00fF
C6154 POR2X1_24/CTRL PAND2X1_9/Y 0.01fF
C6155 PAND2X1_124/Y POR2X1_32/A 0.03fF
C6156 PAND2X1_217/B PAND2X1_203/CTRL 0.01fF
C6157 PAND2X1_488/m4_208_n4# POR2X1_486/m4_208_n4# 0.05fF
C6158 POR2X1_634/A PAND2X1_59/a_76_28# 0.06fF
C6159 PAND2X1_20/A POR2X1_655/A 0.59fF
C6160 PAND2X1_33/CTRL2 POR2X1_5/Y 0.06fF
C6161 POR2X1_818/O POR2X1_734/A 0.30fF
C6162 PAND2X1_93/B POR2X1_788/A 0.03fF
C6163 POR2X1_77/O POR2X1_40/Y 0.09fF
C6164 INPUT_1 PAND2X1_462/CTRL 0.11fF
C6165 POR2X1_846/B POR2X1_846/A 0.37fF
C6166 PAND2X1_282/CTRL POR2X1_590/A 0.01fF
C6167 POR2X1_863/A PAND2X1_173/O 0.01fF
C6168 PAND2X1_603/CTRL POR2X1_78/A 0.01fF
C6169 POR2X1_422/CTRL POR2X1_72/B 0.01fF
C6170 PAND2X1_207/O POR2X1_40/Y 0.01fF
C6171 POR2X1_338/a_16_28# PAND2X1_72/A 0.03fF
C6172 POR2X1_673/Y PAND2X1_529/a_76_28# 0.01fF
C6173 POR2X1_411/B PAND2X1_756/a_16_344# 0.02fF
C6174 POR2X1_814/B POR2X1_655/A 0.84fF
C6175 PAND2X1_245/O POR2X1_296/B 0.00fF
C6176 POR2X1_150/Y PAND2X1_804/B 0.07fF
C6177 POR2X1_83/B POR2X1_32/A 5.25fF
C6178 POR2X1_859/a_76_344# INPUT_0 0.02fF
C6179 PAND2X1_58/A POR2X1_614/Y 0.17fF
C6180 PAND2X1_61/a_16_344# POR2X1_60/A 0.01fF
C6181 PAND2X1_98/a_16_344# INPUT_0 0.04fF
C6182 POR2X1_175/A POR2X1_856/B 0.03fF
C6183 POR2X1_78/A POR2X1_788/A 0.03fF
C6184 POR2X1_78/B POR2X1_222/CTRL2 0.05fF
C6185 PAND2X1_48/B PAND2X1_85/m4_208_n4# 0.15fF
C6186 PAND2X1_746/CTRL PAND2X1_52/B 0.02fF
C6187 POR2X1_568/B POR2X1_188/Y 0.03fF
C6188 INPUT_3 POR2X1_618/CTRL2 0.08fF
C6189 POR2X1_150/Y PAND2X1_390/CTRL2 0.01fF
C6190 POR2X1_863/A POR2X1_456/B 0.06fF
C6191 POR2X1_669/B PAND2X1_706/O 0.04fF
C6192 POR2X1_287/B POR2X1_66/A 1.97fF
C6193 POR2X1_51/A POR2X1_12/A 0.03fF
C6194 PAND2X1_472/B POR2X1_24/Y 0.02fF
C6195 PAND2X1_850/Y POR2X1_589/O 0.03fF
C6196 POR2X1_83/B POR2X1_417/Y 0.08fF
C6197 POR2X1_353/Y POR2X1_220/B 0.04fF
C6198 PAND2X1_611/CTRL2 POR2X1_68/B 0.00fF
C6199 POR2X1_111/CTRL PAND2X1_717/A 0.01fF
C6200 POR2X1_66/B PAND2X1_88/CTRL 0.01fF
C6201 PAND2X1_618/O PAND2X1_6/A 0.05fF
C6202 POR2X1_806/a_56_344# POR2X1_330/Y 0.03fF
C6203 POR2X1_66/B POR2X1_476/CTRL2 0.01fF
C6204 PAND2X1_82/Y POR2X1_98/A 0.02fF
C6205 PAND2X1_85/Y PAND2X1_15/CTRL2 0.04fF
C6206 POR2X1_539/A POR2X1_458/Y 0.07fF
C6207 POR2X1_54/Y POR2X1_642/CTRL 0.01fF
C6208 POR2X1_413/A PAND2X1_634/a_76_28# 0.04fF
C6209 POR2X1_669/B POR2X1_5/Y 0.14fF
C6210 POR2X1_24/Y POR2X1_55/Y 0.01fF
C6211 PAND2X1_20/A POR2X1_637/A 0.00fF
C6212 PAND2X1_625/CTRL2 PAND2X1_39/B 0.01fF
C6213 POR2X1_676/Y POR2X1_678/Y 0.00fF
C6214 PAND2X1_35/Y PAND2X1_124/Y 0.03fF
C6215 POR2X1_366/Y POR2X1_446/B 0.09fF
C6216 POR2X1_66/A PAND2X1_8/Y 0.01fF
C6217 POR2X1_441/Y POR2X1_438/CTRL 0.01fF
C6218 POR2X1_499/A D_INPUT_1 0.03fF
C6219 PAND2X1_462/B PAND2X1_606/CTRL2 0.01fF
C6220 POR2X1_484/CTRL VDD 0.00fF
C6221 POR2X1_66/B PAND2X1_41/B 2.70fF
C6222 POR2X1_491/a_16_28# POR2X1_102/Y 0.01fF
C6223 PAND2X1_6/Y PAND2X1_9/Y 0.03fF
C6224 POR2X1_16/A POR2X1_9/Y 0.07fF
C6225 PAND2X1_558/Y POR2X1_72/B 0.01fF
C6226 POR2X1_523/Y POR2X1_54/Y 0.05fF
C6227 POR2X1_657/Y POR2X1_112/Y 0.07fF
C6228 POR2X1_516/A POR2X1_329/A 0.16fF
C6229 POR2X1_411/B POR2X1_234/a_16_28# 0.02fF
C6230 POR2X1_57/A POR2X1_412/O 0.03fF
C6231 POR2X1_188/A PAND2X1_41/B 0.03fF
C6232 POR2X1_14/Y POR2X1_236/O 0.00fF
C6233 POR2X1_413/A PAND2X1_646/O 0.02fF
C6234 POR2X1_52/A POR2X1_626/CTRL2 0.01fF
C6235 PAND2X1_557/A PAND2X1_363/Y 0.02fF
C6236 POR2X1_478/Y VDD 0.10fF
C6237 POR2X1_120/O POR2X1_78/A 0.03fF
C6238 POR2X1_41/B D_INPUT_0 0.03fF
C6239 POR2X1_415/A POR2X1_816/A 0.13fF
C6240 PAND2X1_117/O POR2X1_558/B 0.00fF
C6241 POR2X1_775/A POR2X1_454/A 0.03fF
C6242 POR2X1_639/A POR2X1_639/O 0.02fF
C6243 PAND2X1_795/B POR2X1_32/A 0.03fF
C6244 POR2X1_614/A POR2X1_624/Y 0.07fF
C6245 POR2X1_590/A PAND2X1_372/CTRL2 0.00fF
C6246 POR2X1_54/Y PAND2X1_69/A 13.78fF
C6247 POR2X1_257/A POR2X1_248/O 0.05fF
C6248 POR2X1_285/a_16_28# POR2X1_590/A 0.03fF
C6249 POR2X1_567/B POR2X1_477/A 0.05fF
C6250 PAND2X1_239/a_56_28# POR2X1_578/Y 0.00fF
C6251 POR2X1_365/O POR2X1_356/Y 0.00fF
C6252 POR2X1_270/Y POR2X1_740/Y 0.04fF
C6253 POR2X1_626/CTRL POR2X1_55/Y 0.01fF
C6254 POR2X1_508/CTRL POR2X1_567/B 0.10fF
C6255 D_INPUT_3 PAND2X1_9/Y 0.05fF
C6256 POR2X1_624/Y POR2X1_38/B 0.07fF
C6257 POR2X1_811/A PAND2X1_599/CTRL2 0.00fF
C6258 POR2X1_467/Y VDD 0.36fF
C6259 PAND2X1_218/A PAND2X1_218/B 0.08fF
C6260 POR2X1_202/A PAND2X1_69/A 0.07fF
C6261 POR2X1_707/B PAND2X1_587/Y 0.01fF
C6262 POR2X1_669/B POR2X1_747/a_16_28# 0.03fF
C6263 POR2X1_83/B PAND2X1_35/Y 0.04fF
C6264 POR2X1_60/A POR2X1_256/O 0.17fF
C6265 PAND2X1_169/O POR2X1_167/Y 0.00fF
C6266 POR2X1_311/Y PAND2X1_793/Y 0.03fF
C6267 POR2X1_556/A POR2X1_569/A 0.07fF
C6268 POR2X1_857/a_76_344# POR2X1_192/Y 0.04fF
C6269 POR2X1_47/CTRL POR2X1_32/A 0.01fF
C6270 POR2X1_49/Y POR2X1_497/Y 0.00fF
C6271 PAND2X1_557/A POR2X1_250/O 0.01fF
C6272 POR2X1_78/B POR2X1_593/B 0.03fF
C6273 POR2X1_60/Y VDD 0.32fF
C6274 POR2X1_649/B POR2X1_862/A 0.41fF
C6275 POR2X1_327/Y POR2X1_814/A 0.06fF
C6276 POR2X1_97/A POR2X1_795/B 0.03fF
C6277 PAND2X1_476/O INPUT_0 0.05fF
C6278 POR2X1_102/Y PAND2X1_188/CTRL2 0.01fF
C6279 POR2X1_121/B POR2X1_294/B 0.03fF
C6280 PAND2X1_480/B POR2X1_72/B 0.08fF
C6281 PAND2X1_475/O POR2X1_46/Y 0.02fF
C6282 POR2X1_859/A PAND2X1_225/a_76_28# 0.01fF
C6283 POR2X1_330/Y POR2X1_722/Y 0.03fF
C6284 POR2X1_264/Y POR2X1_590/A 0.00fF
C6285 POR2X1_683/CTRL POR2X1_40/Y 0.01fF
C6286 PAND2X1_640/O D_INPUT_0 0.01fF
C6287 POR2X1_52/A PAND2X1_465/CTRL 0.00fF
C6288 PAND2X1_862/B PAND2X1_659/A 0.00fF
C6289 PAND2X1_220/A PAND2X1_357/Y 0.01fF
C6290 POR2X1_355/B POR2X1_186/Y 0.10fF
C6291 POR2X1_602/O PAND2X1_60/B 0.01fF
C6292 POR2X1_511/Y POR2X1_236/Y 0.03fF
C6293 POR2X1_63/CTRL POR2X1_83/B 0.01fF
C6294 PAND2X1_543/CTRL POR2X1_236/Y 0.01fF
C6295 POR2X1_526/CTRL2 POR2X1_669/B 0.05fF
C6296 POR2X1_630/A POR2X1_294/B 3.53fF
C6297 PAND2X1_425/Y PAND2X1_157/CTRL 0.01fF
C6298 POR2X1_679/B POR2X1_679/A 0.04fF
C6299 POR2X1_828/Y PAND2X1_760/O 0.17fF
C6300 PAND2X1_65/B PAND2X1_760/CTRL2 0.01fF
C6301 POR2X1_65/A PAND2X1_137/Y 0.03fF
C6302 PAND2X1_23/Y PAND2X1_96/CTRL2 0.00fF
C6303 POR2X1_220/Y POR2X1_61/Y 0.07fF
C6304 POR2X1_709/A POR2X1_789/B 0.01fF
C6305 PAND2X1_85/Y INPUT_0 0.03fF
C6306 POR2X1_288/CTRL PAND2X1_32/B 0.00fF
C6307 POR2X1_632/a_56_344# POR2X1_510/Y 0.00fF
C6308 PAND2X1_229/CTRL POR2X1_231/B 0.00fF
C6309 POR2X1_66/B POR2X1_130/Y 0.01fF
C6310 PAND2X1_659/B PAND2X1_499/Y 0.05fF
C6311 PAND2X1_93/B POR2X1_215/Y 0.01fF
C6312 PAND2X1_23/Y PAND2X1_250/CTRL2 0.05fF
C6313 PAND2X1_48/B PAND2X1_250/CTRL 0.00fF
C6314 POR2X1_175/CTRL POR2X1_566/A 0.31fF
C6315 PAND2X1_651/Y POR2X1_83/B 0.03fF
C6316 PAND2X1_223/a_16_344# POR2X1_7/B 0.02fF
C6317 POR2X1_657/O POR2X1_112/Y 0.01fF
C6318 PAND2X1_454/CTRL2 PAND2X1_803/A 0.00fF
C6319 POR2X1_241/Y VDD 0.00fF
C6320 PAND2X1_639/B PAND2X1_639/O 0.06fF
C6321 POR2X1_383/A POR2X1_286/CTRL 0.01fF
C6322 PAND2X1_76/Y POR2X1_7/B 0.00fF
C6323 POR2X1_83/B PAND2X1_243/CTRL 0.01fF
C6324 POR2X1_66/Y POR2X1_507/A 0.00fF
C6325 POR2X1_68/B POR2X1_390/CTRL 0.01fF
C6326 POR2X1_669/B POR2X1_665/A 0.06fF
C6327 POR2X1_763/A PAND2X1_709/CTRL 0.03fF
C6328 PAND2X1_23/Y POR2X1_475/A 0.07fF
C6329 POR2X1_96/B POR2X1_37/Y 0.06fF
C6330 PAND2X1_46/CTRL2 D_INPUT_1 0.01fF
C6331 PAND2X1_6/Y POR2X1_808/A 0.08fF
C6332 POR2X1_383/A POR2X1_97/A 0.03fF
C6333 PAND2X1_865/O POR2X1_23/Y 0.01fF
C6334 POR2X1_57/A POR2X1_60/A 0.19fF
C6335 PAND2X1_687/O POR2X1_597/Y 0.03fF
C6336 POR2X1_60/A POR2X1_534/CTRL2 0.01fF
C6337 PAND2X1_495/a_16_344# PAND2X1_20/A 0.02fF
C6338 PAND2X1_84/Y POR2X1_293/Y 0.02fF
C6339 POR2X1_102/Y PAND2X1_388/Y 0.03fF
C6340 POR2X1_52/A PAND2X1_520/CTRL 0.01fF
C6341 POR2X1_860/CTRL2 POR2X1_218/Y 0.10fF
C6342 POR2X1_296/B POR2X1_366/A 0.03fF
C6343 PAND2X1_668/O PAND2X1_673/Y 0.12fF
C6344 PAND2X1_73/Y POR2X1_222/A 0.03fF
C6345 POR2X1_653/CTRL2 POR2X1_740/Y 0.00fF
C6346 POR2X1_73/a_56_344# POR2X1_37/Y 0.01fF
C6347 POR2X1_263/Y PAND2X1_737/B 0.01fF
C6348 POR2X1_329/A PAND2X1_339/CTRL2 0.01fF
C6349 PAND2X1_345/CTRL PAND2X1_555/A 0.01fF
C6350 POR2X1_57/A POR2X1_591/A 0.02fF
C6351 PAND2X1_833/O POR2X1_495/Y 0.15fF
C6352 POR2X1_260/B POR2X1_596/a_16_28# 0.02fF
C6353 POR2X1_347/A PAND2X1_94/CTRL 0.01fF
C6354 POR2X1_291/O D_INPUT_0 0.07fF
C6355 PAND2X1_57/B PAND2X1_322/a_16_344# 0.02fF
C6356 POR2X1_106/Y PAND2X1_357/Y 0.03fF
C6357 POR2X1_590/A PAND2X1_528/CTRL 0.02fF
C6358 PAND2X1_95/B VDD 0.76fF
C6359 POR2X1_834/Y D_INPUT_0 0.00fF
C6360 PAND2X1_865/Y POR2X1_20/B 0.07fF
C6361 PAND2X1_23/Y POR2X1_349/Y 0.00fF
C6362 POR2X1_102/Y PAND2X1_549/B 0.06fF
C6363 PAND2X1_96/B POR2X1_288/A 0.02fF
C6364 POR2X1_83/B POR2X1_9/a_16_28# 0.01fF
C6365 PAND2X1_90/Y POR2X1_391/Y 0.44fF
C6366 PAND2X1_863/B POR2X1_7/B 0.03fF
C6367 POR2X1_66/B POR2X1_228/Y 0.10fF
C6368 POR2X1_83/B POR2X1_503/Y 0.05fF
C6369 POR2X1_454/A POR2X1_339/Y 0.01fF
C6370 POR2X1_687/A POR2X1_687/a_16_28# 0.04fF
C6371 PAND2X1_673/Y POR2X1_42/Y 0.03fF
C6372 POR2X1_65/O POR2X1_39/B 0.27fF
C6373 D_INPUT_0 PAND2X1_690/O 0.15fF
C6374 PAND2X1_658/B PAND2X1_512/Y 0.00fF
C6375 POR2X1_43/B PAND2X1_735/CTRL 0.02fF
C6376 POR2X1_212/A POR2X1_191/Y 0.05fF
C6377 POR2X1_184/Y PAND2X1_140/Y 0.02fF
C6378 POR2X1_68/A POR2X1_284/B 0.03fF
C6379 PAND2X1_140/A POR2X1_251/O 0.02fF
C6380 POR2X1_287/B POR2X1_532/A 0.03fF
C6381 PAND2X1_93/CTRL2 PAND2X1_57/B 0.11fF
C6382 POR2X1_567/A POR2X1_446/B 0.03fF
C6383 PAND2X1_436/A PAND2X1_549/B 0.12fF
C6384 PAND2X1_357/Y PAND2X1_580/B 0.03fF
C6385 POR2X1_174/B POR2X1_502/O 0.00fF
C6386 PAND2X1_795/B POR2X1_184/Y 0.57fF
C6387 POR2X1_13/A POR2X1_494/CTRL2 0.00fF
C6388 POR2X1_579/Y POR2X1_785/A 0.03fF
C6389 POR2X1_625/m4_208_n4# POR2X1_90/Y 0.07fF
C6390 PAND2X1_750/a_76_28# POR2X1_749/Y 0.05fF
C6391 PAND2X1_59/B PAND2X1_3/B 0.05fF
C6392 POR2X1_220/Y POR2X1_35/Y 0.03fF
C6393 POR2X1_231/CTRL2 POR2X1_795/B 0.05fF
C6394 POR2X1_538/CTRL2 POR2X1_193/A 0.03fF
C6395 POR2X1_814/B PAND2X1_757/O 0.03fF
C6396 PAND2X1_137/Y PAND2X1_190/Y 0.10fF
C6397 POR2X1_483/A POR2X1_532/A 0.03fF
C6398 PAND2X1_688/CTRL2 POR2X1_38/Y 0.01fF
C6399 PAND2X1_129/O POR2X1_68/B 0.03fF
C6400 PAND2X1_90/Y POR2X1_712/CTRL2 0.06fF
C6401 PAND2X1_766/CTRL2 POR2X1_707/Y 0.00fF
C6402 PAND2X1_743/O VDD 0.00fF
C6403 POR2X1_68/A POR2X1_855/Y 0.01fF
C6404 POR2X1_241/Y PAND2X1_32/B 0.07fF
C6405 POR2X1_60/A PAND2X1_301/O 0.17fF
C6406 INPUT_1 PAND2X1_77/m4_208_n4# 0.12fF
C6407 POR2X1_46/Y PAND2X1_546/O 0.03fF
C6408 PAND2X1_140/A POR2X1_106/Y 0.01fF
C6409 POR2X1_35/Y POR2X1_404/Y 0.04fF
C6410 POR2X1_383/A POR2X1_650/A 0.03fF
C6411 POR2X1_777/B POR2X1_249/Y 0.05fF
C6412 POR2X1_856/B POR2X1_337/Y 0.10fF
C6413 POR2X1_532/A PAND2X1_8/Y 0.03fF
C6414 POR2X1_43/B PAND2X1_115/B 0.53fF
C6415 PAND2X1_700/a_16_344# POR2X1_532/A 0.01fF
C6416 POR2X1_366/Y PAND2X1_56/Y 0.05fF
C6417 PAND2X1_56/Y POR2X1_294/B 0.03fF
C6418 POR2X1_795/B POR2X1_294/B 0.14fF
C6419 PAND2X1_742/B POR2X1_331/a_16_28# 0.01fF
C6420 PAND2X1_566/Y POR2X1_7/B 1.51fF
C6421 POR2X1_627/CTRL POR2X1_7/A 0.01fF
C6422 POR2X1_131/Y PAND2X1_140/CTRL 0.01fF
C6423 PAND2X1_584/O POR2X1_774/B 0.04fF
C6424 PAND2X1_96/B PAND2X1_516/O 0.03fF
C6425 POR2X1_778/B POR2X1_784/A 0.01fF
C6426 POR2X1_236/Y POR2X1_511/a_56_344# 0.00fF
C6427 VDD POR2X1_350/B 0.29fF
C6428 POR2X1_137/Y INPUT_0 0.25fF
C6429 POR2X1_61/Y POR2X1_215/A 0.45fF
C6430 PAND2X1_206/CTRL2 POR2X1_7/A 0.01fF
C6431 POR2X1_357/a_16_28# POR2X1_97/A 0.03fF
C6432 POR2X1_634/A POR2X1_559/A 0.12fF
C6433 PAND2X1_811/O PAND2X1_568/B 0.02fF
C6434 POR2X1_316/CTRL2 PAND2X1_436/A 0.03fF
C6435 POR2X1_556/A PAND2X1_72/A 0.26fF
C6436 PAND2X1_108/O PAND2X1_60/B 0.04fF
C6437 POR2X1_614/A POR2X1_785/A 0.06fF
C6438 POR2X1_43/B PAND2X1_658/A 0.03fF
C6439 POR2X1_13/A POR2X1_9/CTRL 0.01fF
C6440 POR2X1_41/B POR2X1_111/CTRL 0.08fF
C6441 POR2X1_150/Y PAND2X1_332/Y 0.03fF
C6442 PAND2X1_365/B POR2X1_42/Y 0.05fF
C6443 PAND2X1_755/CTRL PAND2X1_60/B 0.01fF
C6444 POR2X1_376/B PAND2X1_155/CTRL 0.01fF
C6445 PAND2X1_9/Y PAND2X1_52/B 0.05fF
C6446 POR2X1_660/Y POR2X1_512/O 0.02fF
C6447 PAND2X1_65/B POR2X1_249/Y 0.00fF
C6448 POR2X1_327/Y POR2X1_405/CTRL2 0.01fF
C6449 POR2X1_20/O POR2X1_68/B 0.01fF
C6450 PAND2X1_462/B INPUT_2 0.17fF
C6451 POR2X1_105/Y POR2X1_260/A 0.03fF
C6452 POR2X1_717/Y POR2X1_501/B 0.03fF
C6453 POR2X1_124/a_16_28# POR2X1_124/B -0.00fF
C6454 POR2X1_802/B POR2X1_209/A 0.03fF
C6455 PAND2X1_651/Y PAND2X1_242/CTRL 0.00fF
C6456 PAND2X1_95/B PAND2X1_32/B 0.19fF
C6457 POR2X1_65/A POR2X1_766/a_16_28# 0.01fF
C6458 PAND2X1_682/O POR2X1_68/A 0.05fF
C6459 POR2X1_130/A POR2X1_725/Y 0.10fF
C6460 PAND2X1_20/A PAND2X1_527/O 0.05fF
C6461 POR2X1_392/a_16_28# PAND2X1_32/B 0.01fF
C6462 PAND2X1_716/CTRL2 POR2X1_52/Y 0.00fF
C6463 POR2X1_583/CTRL2 POR2X1_42/Y 0.03fF
C6464 POR2X1_834/Y PAND2X1_90/Y 0.15fF
C6465 VDD PAND2X1_112/CTRL 0.00fF
C6466 POR2X1_72/B POR2X1_373/Y 0.41fF
C6467 POR2X1_719/CTRL2 PAND2X1_48/B 0.03fF
C6468 POR2X1_13/A PAND2X1_196/CTRL2 0.00fF
C6469 POR2X1_236/Y PAND2X1_124/O 0.02fF
C6470 POR2X1_518/Y PAND2X1_642/B 0.00fF
C6471 PAND2X1_484/O PAND2X1_41/B 0.01fF
C6472 PAND2X1_291/CTRL2 POR2X1_198/B 0.03fF
C6473 POR2X1_71/CTRL2 POR2X1_5/Y 0.00fF
C6474 POR2X1_677/CTRL POR2X1_129/Y 0.01fF
C6475 POR2X1_49/Y POR2X1_177/O 0.01fF
C6476 D_GATE_662 POR2X1_540/A 0.07fF
C6477 PAND2X1_57/B POR2X1_796/A 0.03fF
C6478 POR2X1_697/Y POR2X1_511/CTRL 0.01fF
C6479 POR2X1_43/B POR2X1_73/Y 0.17fF
C6480 POR2X1_197/Y PAND2X1_48/B 0.03fF
C6481 POR2X1_174/CTRL VDD 0.00fF
C6482 PAND2X1_678/CTRL PAND2X1_860/A 0.01fF
C6483 POR2X1_493/CTRL POR2X1_572/B 0.00fF
C6484 POR2X1_78/A POR2X1_374/O 0.20fF
C6485 POR2X1_311/a_16_28# POR2X1_481/A 0.02fF
C6486 POR2X1_861/a_16_28# POR2X1_501/B 0.00fF
C6487 POR2X1_88/Y PAND2X1_100/O 0.00fF
C6488 POR2X1_278/Y POR2X1_16/A 0.20fF
C6489 D_INPUT_0 POR2X1_77/Y 0.06fF
C6490 POR2X1_833/A INPUT_0 0.07fF
C6491 POR2X1_383/A POR2X1_294/B 0.45fF
C6492 PAND2X1_723/Y POR2X1_394/A 0.01fF
C6493 POR2X1_366/Y POR2X1_383/A 0.01fF
C6494 PAND2X1_743/O PAND2X1_32/B 0.08fF
C6495 PAND2X1_56/Y PAND2X1_111/B 0.01fF
C6496 POR2X1_216/Y VDD 0.10fF
C6497 POR2X1_32/A PAND2X1_841/Y 0.12fF
C6498 POR2X1_85/Y D_INPUT_0 0.25fF
C6499 POR2X1_337/CTRL2 POR2X1_260/A 0.00fF
C6500 POR2X1_129/Y POR2X1_236/Y 0.40fF
C6501 POR2X1_36/B POR2X1_581/O 0.01fF
C6502 POR2X1_3/A POR2X1_581/a_56_344# 0.01fF
C6503 POR2X1_114/CTRL2 POR2X1_113/Y 0.02fF
C6504 POR2X1_680/CTRL2 POR2X1_40/Y 0.03fF
C6505 PAND2X1_666/CTRL2 PAND2X1_72/A 0.01fF
C6506 PAND2X1_472/CTRL2 POR2X1_7/B 0.03fF
C6507 POR2X1_760/A PAND2X1_405/a_16_344# 0.02fF
C6508 POR2X1_66/B PAND2X1_665/O 0.16fF
C6509 POR2X1_330/Y POR2X1_330/CTRL 0.08fF
C6510 POR2X1_16/A POR2X1_829/A 0.03fF
C6511 POR2X1_228/Y POR2X1_556/m4_208_n4# 0.08fF
C6512 PAND2X1_109/a_56_28# POR2X1_97/A 0.00fF
C6513 POR2X1_78/A PAND2X1_179/a_76_28# 0.01fF
C6514 POR2X1_728/a_16_28# POR2X1_730/Y 0.02fF
C6515 POR2X1_522/Y PAND2X1_844/B 0.03fF
C6516 PAND2X1_94/A PAND2X1_92/a_76_28# 0.01fF
C6517 POR2X1_590/a_16_28# POR2X1_294/B 0.03fF
C6518 POR2X1_343/Y POR2X1_590/A 0.05fF
C6519 PAND2X1_564/O POR2X1_394/A 0.01fF
C6520 PAND2X1_357/Y PAND2X1_349/A 0.08fF
C6521 PAND2X1_342/CTRL2 POR2X1_248/Y 0.01fF
C6522 POR2X1_687/A POR2X1_730/CTRL 0.01fF
C6523 PAND2X1_48/B INPUT_1 0.03fF
C6524 PAND2X1_549/B POR2X1_531/Y 0.00fF
C6525 POR2X1_722/CTRL2 VDD 0.00fF
C6526 POR2X1_43/B PAND2X1_244/B 0.03fF
C6527 POR2X1_244/B POR2X1_228/CTRL2 0.01fF
C6528 PAND2X1_41/B POR2X1_199/B 0.01fF
C6529 POR2X1_494/CTRL2 PAND2X1_510/B 0.01fF
C6530 POR2X1_272/Y PAND2X1_716/B 0.52fF
C6531 PAND2X1_723/CTRL POR2X1_7/A 0.01fF
C6532 PAND2X1_569/B PAND2X1_551/A 0.00fF
C6533 PAND2X1_659/Y POR2X1_236/Y 0.07fF
C6534 PAND2X1_69/A POR2X1_148/B 0.02fF
C6535 PAND2X1_793/Y POR2X1_153/Y 0.03fF
C6536 PAND2X1_508/Y POR2X1_516/B 1.29fF
C6537 POR2X1_814/CTRL2 POR2X1_260/B 0.01fF
C6538 POR2X1_215/A POR2X1_35/Y 0.00fF
C6539 POR2X1_339/a_76_344# POR2X1_785/A 0.01fF
C6540 PAND2X1_841/B POR2X1_153/Y 0.04fF
C6541 POR2X1_840/CTRL2 POR2X1_725/Y 0.05fF
C6542 POR2X1_40/Y POR2X1_39/B 1.90fF
C6543 POR2X1_68/A PAND2X1_94/A 0.33fF
C6544 POR2X1_762/CTRL INPUT_4 0.01fF
C6545 PAND2X1_787/A POR2X1_91/Y 0.03fF
C6546 POR2X1_123/B PAND2X1_60/B 0.22fF
C6547 POR2X1_156/B POR2X1_855/B 0.12fF
C6548 PAND2X1_6/Y POR2X1_687/A 0.02fF
C6549 POR2X1_510/Y PAND2X1_88/Y 0.03fF
C6550 PAND2X1_661/B PAND2X1_196/CTRL2 0.01fF
C6551 POR2X1_193/A POR2X1_186/B 0.57fF
C6552 PAND2X1_702/O POR2X1_7/A 0.01fF
C6553 PAND2X1_182/B POR2X1_55/Y 3.09fF
C6554 PAND2X1_54/a_16_344# POR2X1_4/Y 0.02fF
C6555 POR2X1_579/Y POR2X1_186/B 0.03fF
C6556 POR2X1_114/CTRL2 POR2X1_260/A 0.00fF
C6557 PAND2X1_113/O POR2X1_107/Y -0.00fF
C6558 PAND2X1_687/B POR2X1_236/Y 0.03fF
C6559 POR2X1_7/B POR2X1_523/B 0.00fF
C6560 POR2X1_13/A POR2X1_171/Y 0.02fF
C6561 PAND2X1_687/CTRL POR2X1_829/A 0.00fF
C6562 POR2X1_791/CTRL2 PAND2X1_48/A 0.32fF
C6563 POR2X1_68/A POR2X1_782/CTRL 0.01fF
C6564 PAND2X1_854/Y VDD 0.00fF
C6565 POR2X1_687/Y POR2X1_729/Y 0.12fF
C6566 PAND2X1_90/Y POR2X1_383/Y 0.05fF
C6567 PAND2X1_455/O POR2X1_77/Y 0.03fF
C6568 PAND2X1_738/B POR2X1_77/Y 0.03fF
C6569 POR2X1_829/A POR2X1_599/a_16_28# 0.05fF
C6570 POR2X1_327/Y POR2X1_302/A 0.01fF
C6571 POR2X1_383/A PAND2X1_111/B 0.03fF
C6572 POR2X1_16/A INPUT_2 0.00fF
C6573 PAND2X1_805/Y PAND2X1_221/Y 0.03fF
C6574 POR2X1_425/Y POR2X1_158/B 0.01fF
C6575 POR2X1_275/a_16_28# POR2X1_129/Y 0.03fF
C6576 PAND2X1_140/A PAND2X1_349/A 0.00fF
C6577 POR2X1_865/B POR2X1_276/Y 0.03fF
C6578 PAND2X1_90/Y POR2X1_779/CTRL 0.03fF
C6579 POR2X1_57/A POR2X1_744/CTRL 0.01fF
C6580 POR2X1_697/Y PAND2X1_708/a_16_344# 0.03fF
C6581 POR2X1_536/CTRL2 PAND2X1_222/B 0.01fF
C6582 POR2X1_465/B POR2X1_540/Y 0.00fF
C6583 PAND2X1_737/CTRL POR2X1_7/B 0.01fF
C6584 POR2X1_52/A PAND2X1_639/Y 0.12fF
C6585 PAND2X1_427/a_76_28# PAND2X1_72/A 0.01fF
C6586 PAND2X1_140/A PAND2X1_114/B 0.03fF
C6587 POR2X1_276/A POR2X1_569/A 0.03fF
C6588 POR2X1_614/A POR2X1_186/B 0.20fF
C6589 PAND2X1_439/CTRL2 POR2X1_438/Y 0.03fF
C6590 PAND2X1_4/O POR2X1_260/A 0.01fF
C6591 POR2X1_307/CTRL2 POR2X1_661/A 0.05fF
C6592 POR2X1_294/B POR2X1_788/CTRL 0.06fF
C6593 POR2X1_527/Y PAND2X1_550/B 0.01fF
C6594 POR2X1_129/Y PAND2X1_858/Y 0.01fF
C6595 PAND2X1_170/CTRL POR2X1_73/Y 0.01fF
C6596 POR2X1_472/Y PAND2X1_52/B 0.01fF
C6597 POR2X1_567/A POR2X1_795/B 0.10fF
C6598 PAND2X1_341/B PAND2X1_341/a_76_28# 0.01fF
C6599 POR2X1_178/Y PAND2X1_181/a_16_344# 0.03fF
C6600 PAND2X1_236/CTRL PAND2X1_52/B 0.28fF
C6601 POR2X1_8/Y POR2X1_283/A 0.10fF
C6602 POR2X1_72/B POR2X1_386/Y 0.00fF
C6603 INPUT_3 POR2X1_415/A 0.01fF
C6604 VDD PAND2X1_351/A 0.00fF
C6605 PAND2X1_824/B POR2X1_201/Y 0.02fF
C6606 PAND2X1_69/A POR2X1_4/Y 0.35fF
C6607 POR2X1_54/a_16_28# D_INPUT_1 0.00fF
C6608 POR2X1_27/O POR2X1_669/B 0.01fF
C6609 PAND2X1_635/Y POR2X1_748/A 0.04fF
C6610 PAND2X1_71/Y PAND2X1_111/B 3.87fF
C6611 INPUT_1 POR2X1_376/CTRL 0.01fF
C6612 POR2X1_68/B PAND2X1_396/CTRL 0.01fF
C6613 POR2X1_447/B POR2X1_631/A 0.04fF
C6614 POR2X1_394/A PAND2X1_346/Y 7.39fF
C6615 PAND2X1_800/O PAND2X1_691/Y 0.03fF
C6616 POR2X1_93/A POR2X1_4/Y 0.03fF
C6617 POR2X1_702/a_16_28# POR2X1_186/B 0.01fF
C6618 PAND2X1_631/A PAND2X1_344/O 0.10fF
C6619 POR2X1_624/O POR2X1_94/A 0.01fF
C6620 POR2X1_283/A POR2X1_385/Y 0.05fF
C6621 POR2X1_135/CTRL POR2X1_7/A 0.01fF
C6622 PAND2X1_351/a_76_28# PAND2X1_351/A 0.02fF
C6623 POR2X1_416/B POR2X1_672/A 0.02fF
C6624 POR2X1_567/A POR2X1_383/A 0.30fF
C6625 PAND2X1_566/O PAND2X1_303/Y 0.00fF
C6626 POR2X1_171/Y PAND2X1_510/B 0.02fF
C6627 PAND2X1_93/B POR2X1_76/A 0.03fF
C6628 POR2X1_14/O INPUT_3 0.01fF
C6629 POR2X1_499/A POR2X1_78/A 0.03fF
C6630 POR2X1_306/Y POR2X1_329/A 0.02fF
C6631 POR2X1_160/CTRL2 POR2X1_356/B 0.07fF
C6632 PAND2X1_20/A POR2X1_227/A 0.00fF
C6633 POR2X1_760/A PAND2X1_361/a_16_344# 0.01fF
C6634 POR2X1_860/CTRL2 POR2X1_861/A 0.01fF
C6635 POR2X1_514/CTRL2 POR2X1_138/A 0.00fF
C6636 POR2X1_119/Y PAND2X1_737/B 0.05fF
C6637 POR2X1_394/A PAND2X1_123/Y 0.03fF
C6638 PAND2X1_50/O D_INPUT_7 0.04fF
C6639 POR2X1_449/A POR2X1_652/A 0.01fF
C6640 PAND2X1_19/Y VDD 0.12fF
C6641 PAND2X1_611/O POR2X1_389/Y 0.02fF
C6642 POR2X1_327/Y POR2X1_151/Y 0.10fF
C6643 POR2X1_309/a_16_28# POR2X1_411/B 0.02fF
C6644 POR2X1_777/B PAND2X1_246/a_16_344# 0.02fF
C6645 PAND2X1_65/B POR2X1_260/CTRL 0.01fF
C6646 POR2X1_23/Y PAND2X1_477/a_16_344# 0.03fF
C6647 POR2X1_866/A POR2X1_811/O 0.02fF
C6648 PAND2X1_478/B POR2X1_20/B 0.03fF
C6649 POR2X1_624/Y POR2X1_590/A 1.67fF
C6650 POR2X1_838/B PAND2X1_67/CTRL2 0.00fF
C6651 POR2X1_9/Y PAND2X1_57/B 0.10fF
C6652 PAND2X1_686/O POR2X1_684/Y 0.00fF
C6653 POR2X1_639/Y PAND2X1_52/B 0.03fF
C6654 POR2X1_416/B POR2X1_387/Y 0.15fF
C6655 POR2X1_416/B POR2X1_695/CTRL 0.01fF
C6656 POR2X1_158/Y POR2X1_695/CTRL2 0.00fF
C6657 PAND2X1_74/O POR2X1_341/A 0.05fF
C6658 POR2X1_579/CTRL2 PAND2X1_32/B 0.01fF
C6659 POR2X1_411/B POR2X1_272/O 0.02fF
C6660 POR2X1_411/B PAND2X1_390/Y 0.03fF
C6661 PAND2X1_26/A PAND2X1_11/Y 0.78fF
C6662 POR2X1_319/A POR2X1_454/B 0.06fF
C6663 POR2X1_431/CTRL VDD 0.00fF
C6664 POR2X1_150/Y PAND2X1_562/B 0.07fF
C6665 POR2X1_416/B PAND2X1_551/a_56_28# 0.00fF
C6666 PAND2X1_717/A PAND2X1_735/Y 0.07fF
C6667 PAND2X1_175/B PAND2X1_862/CTRL 0.01fF
C6668 POR2X1_499/A POR2X1_573/CTRL 0.01fF
C6669 PAND2X1_771/Y PAND2X1_577/Y 3.75fF
C6670 POR2X1_257/A POR2X1_423/Y 0.07fF
C6671 POR2X1_35/B POR2X1_621/A 0.00fF
C6672 POR2X1_623/Y VDD 0.00fF
C6673 PAND2X1_637/O PAND2X1_638/B 0.02fF
C6674 POR2X1_491/Y POR2X1_394/A 0.05fF
C6675 POR2X1_769/Y PAND2X1_52/B 0.01fF
C6676 POR2X1_49/Y PAND2X1_469/CTRL 0.01fF
C6677 POR2X1_647/B POR2X1_814/B 0.03fF
C6678 POR2X1_809/a_16_28# POR2X1_121/B 0.09fF
C6679 POR2X1_35/B POR2X1_34/CTRL2 0.01fF
C6680 POR2X1_180/A PAND2X1_72/A 0.05fF
C6681 POR2X1_687/A PAND2X1_52/B 0.02fF
C6682 POR2X1_837/B POR2X1_402/A 0.01fF
C6683 PAND2X1_812/A PAND2X1_865/Y 0.02fF
C6684 POR2X1_648/Y POR2X1_294/B 0.06fF
C6685 PAND2X1_717/A PAND2X1_493/Y 0.06fF
C6686 POR2X1_566/A POR2X1_318/CTRL2 0.32fF
C6687 POR2X1_169/a_16_28# POR2X1_169/A 0.03fF
C6688 POR2X1_352/O PAND2X1_52/B 0.10fF
C6689 PAND2X1_623/a_16_344# POR2X1_669/B 0.10fF
C6690 POR2X1_416/B POR2X1_419/a_16_28# 0.01fF
C6691 POR2X1_13/A POR2X1_150/Y 0.03fF
C6692 PAND2X1_235/CTRL2 POR2X1_296/B 0.00fF
C6693 POR2X1_357/B POR2X1_182/O 0.05fF
C6694 POR2X1_352/O POR2X1_212/B 0.01fF
C6695 POR2X1_48/A POR2X1_40/Y 10.76fF
C6696 PAND2X1_48/B POR2X1_462/O 0.01fF
C6697 POR2X1_16/A POR2X1_824/m4_208_n4# 0.09fF
C6698 POR2X1_685/a_16_28# POR2X1_452/Y 0.03fF
C6699 POR2X1_458/Y PAND2X1_69/A 0.13fF
C6700 POR2X1_287/B POR2X1_458/O 0.00fF
C6701 POR2X1_65/A POR2X1_23/Y 0.13fF
C6702 POR2X1_32/A PAND2X1_444/Y 0.13fF
C6703 POR2X1_96/A POR2X1_628/Y 0.16fF
C6704 POR2X1_812/O POR2X1_452/Y 0.00fF
C6705 POR2X1_137/B PAND2X1_132/O 0.07fF
C6706 POR2X1_655/A VDD 0.12fF
C6707 POR2X1_20/B POR2X1_494/Y 0.02fF
C6708 PAND2X1_73/Y PAND2X1_46/CTRL 0.03fF
C6709 PAND2X1_841/CTRL POR2X1_271/B 0.01fF
C6710 POR2X1_54/Y POR2X1_121/Y 0.03fF
C6711 POR2X1_45/CTRL POR2X1_23/Y 0.01fF
C6712 POR2X1_801/O POR2X1_801/B 0.00fF
C6713 POR2X1_515/a_16_28# POR2X1_446/B -0.00fF
C6714 POR2X1_416/Y POR2X1_412/CTRL2 0.01fF
C6715 POR2X1_83/B PAND2X1_249/O 0.04fF
C6716 POR2X1_833/O POR2X1_541/B 0.06fF
C6717 POR2X1_416/B PAND2X1_737/CTRL2 0.03fF
C6718 POR2X1_630/B POR2X1_532/A 0.01fF
C6719 POR2X1_83/B PAND2X1_731/B 0.03fF
C6720 PAND2X1_617/CTRL POR2X1_68/B 0.03fF
C6721 PAND2X1_476/O POR2X1_102/Y 0.03fF
C6722 PAND2X1_94/A PAND2X1_233/O 0.08fF
C6723 POR2X1_445/A POR2X1_465/B 0.03fF
C6724 POR2X1_79/Y PAND2X1_205/CTRL 0.01fF
C6725 POR2X1_96/A POR2X1_271/CTRL 0.02fF
C6726 PAND2X1_449/CTRL POR2X1_90/Y 0.01fF
C6727 POR2X1_37/Y POR2X1_236/Y 1.78fF
C6728 POR2X1_669/B PAND2X1_381/CTRL 0.12fF
C6729 POR2X1_682/CTRL2 POR2X1_60/A 0.01fF
C6730 PAND2X1_721/B PAND2X1_721/CTRL2 0.01fF
C6731 POR2X1_852/B POR2X1_629/B 0.06fF
C6732 POR2X1_377/CTRL POR2X1_54/Y 0.01fF
C6733 POR2X1_296/O PAND2X1_69/A 0.01fF
C6734 POR2X1_19/CTRL2 POR2X1_38/B 0.00fF
C6735 POR2X1_271/Y PAND2X1_390/Y 0.00fF
C6736 POR2X1_48/A POR2X1_481/O 0.11fF
C6737 POR2X1_329/A PAND2X1_175/B 0.03fF
C6738 PAND2X1_407/a_16_344# POR2X1_55/Y 0.04fF
C6739 PAND2X1_624/O POR2X1_29/A 0.03fF
C6740 PAND2X1_58/A POR2X1_585/O 0.02fF
C6741 PAND2X1_232/O POR2X1_98/A 0.08fF
C6742 PAND2X1_463/O POR2X1_94/A 0.01fF
C6743 PAND2X1_772/O PAND2X1_768/Y 0.00fF
C6744 POR2X1_68/CTRL PAND2X1_57/B 0.01fF
C6745 POR2X1_356/A POR2X1_446/m4_208_n4# 0.06fF
C6746 POR2X1_78/B POR2X1_240/B 0.07fF
C6747 POR2X1_814/B POR2X1_461/A 0.03fF
C6748 PAND2X1_717/A PAND2X1_569/B 0.52fF
C6749 POR2X1_814/A POR2X1_249/Y 0.03fF
C6750 PAND2X1_612/B PAND2X1_283/O 0.00fF
C6751 POR2X1_460/CTRL POR2X1_260/B 0.01fF
C6752 PAND2X1_443/Y VDD 0.05fF
C6753 POR2X1_81/Y POR2X1_37/Y 0.02fF
C6754 PAND2X1_843/CTRL PAND2X1_220/Y 0.15fF
C6755 POR2X1_269/A PAND2X1_57/B 0.00fF
C6756 POR2X1_284/B PAND2X1_58/A 0.03fF
C6757 POR2X1_65/A POR2X1_312/Y 0.03fF
C6758 PAND2X1_243/B POR2X1_409/B 0.03fF
C6759 POR2X1_836/O POR2X1_578/Y 0.02fF
C6760 PAND2X1_695/O POR2X1_634/A 0.28fF
C6761 POR2X1_376/B PAND2X1_390/Y 0.05fF
C6762 POR2X1_60/A PAND2X1_84/Y 0.01fF
C6763 POR2X1_130/A POR2X1_811/B 0.02fF
C6764 POR2X1_582/CTRL POR2X1_257/A 0.01fF
C6765 POR2X1_92/CTRL INPUT_3 0.05fF
C6766 PAND2X1_833/a_16_344# POR2X1_60/A 0.00fF
C6767 PAND2X1_793/Y PAND2X1_794/CTRL2 0.01fF
C6768 POR2X1_323/CTRL POR2X1_65/A 0.01fF
C6769 POR2X1_72/B PAND2X1_473/B 0.03fF
C6770 PAND2X1_319/B POR2X1_257/A 0.03fF
C6771 PAND2X1_23/Y POR2X1_637/CTRL 0.10fF
C6772 POR2X1_23/Y PAND2X1_190/Y 0.05fF
C6773 POR2X1_655/A PAND2X1_32/B 0.03fF
C6774 PAND2X1_557/A VDD 0.19fF
C6775 POR2X1_264/Y POR2X1_66/A 0.03fF
C6776 POR2X1_346/CTRL2 POR2X1_202/A 0.03fF
C6777 POR2X1_266/O PAND2X1_69/A 0.13fF
C6778 PAND2X1_489/O PAND2X1_794/B 0.04fF
C6779 PAND2X1_287/Y PAND2X1_578/A 0.17fF
C6780 POR2X1_257/A POR2X1_582/A 0.00fF
C6781 PAND2X1_848/B POR2X1_48/A 0.02fF
C6782 POR2X1_341/A POR2X1_510/Y 0.07fF
C6783 POR2X1_346/B POR2X1_66/CTRL 0.00fF
C6784 POR2X1_302/Y POR2X1_330/Y 0.05fF
C6785 POR2X1_590/A POR2X1_785/A 0.03fF
C6786 POR2X1_697/Y POR2X1_32/A 0.06fF
C6787 PAND2X1_480/B POR2X1_272/CTRL2 0.26fF
C6788 PAND2X1_652/Y POR2X1_83/B 0.01fF
C6789 PAND2X1_251/O PAND2X1_69/A 0.03fF
C6790 POR2X1_590/A PAND2X1_536/CTRL2 0.01fF
C6791 POR2X1_628/Y POR2X1_7/A 0.66fF
C6792 POR2X1_637/A VDD 0.00fF
C6793 POR2X1_502/A POR2X1_602/B 1.92fF
C6794 POR2X1_66/B POR2X1_360/A 0.03fF
C6795 POR2X1_68/A POR2X1_801/B 0.03fF
C6796 PAND2X1_453/O POR2X1_14/Y 0.15fF
C6797 POR2X1_378/Y PAND2X1_459/O 0.03fF
C6798 POR2X1_232/Y POR2X1_37/Y 0.03fF
C6799 PAND2X1_479/CTRL VDD 0.00fF
C6800 POR2X1_13/A PAND2X1_244/a_76_28# 0.01fF
C6801 POR2X1_482/Y POR2X1_252/O 0.01fF
C6802 POR2X1_68/CTRL2 PAND2X1_69/A 0.03fF
C6803 POR2X1_494/CTRL2 POR2X1_29/A 0.01fF
C6804 POR2X1_43/B POR2X1_753/Y 0.04fF
C6805 POR2X1_52/A PAND2X1_455/CTRL2 0.03fF
C6806 POR2X1_645/a_16_28# POR2X1_718/A 0.03fF
C6807 POR2X1_650/A INPUT_0 0.03fF
C6808 POR2X1_647/O PAND2X1_60/B 0.01fF
C6809 PAND2X1_52/B POR2X1_568/A 0.05fF
C6810 PAND2X1_843/O POR2X1_251/Y 0.09fF
C6811 POR2X1_260/B POR2X1_537/B 3.15fF
C6812 POR2X1_83/A PAND2X1_721/B 0.03fF
C6813 POR2X1_407/A POR2X1_287/CTRL 0.00fF
C6814 PAND2X1_94/A POR2X1_709/A 0.01fF
C6815 POR2X1_260/B POR2X1_391/CTRL2 0.02fF
C6816 POR2X1_212/B POR2X1_568/A 0.04fF
C6817 POR2X1_423/Y PAND2X1_553/B 1.39fF
C6818 PAND2X1_784/CTRL POR2X1_72/B 0.01fF
C6819 POR2X1_346/CTRL2 POR2X1_346/A 0.01fF
C6820 PAND2X1_48/Y PAND2X1_57/B 0.02fF
C6821 POR2X1_407/A POR2X1_121/B 0.06fF
C6822 PAND2X1_267/Y POR2X1_7/A 0.01fF
C6823 PAND2X1_222/A PAND2X1_537/CTRL2 0.00fF
C6824 PAND2X1_90/A POR2X1_720/Y 0.01fF
C6825 POR2X1_302/CTRL POR2X1_302/Y 0.00fF
C6826 POR2X1_29/A POR2X1_409/O 0.01fF
C6827 POR2X1_505/Y POR2X1_42/Y 0.30fF
C6828 POR2X1_297/Y PAND2X1_347/Y 0.01fF
C6829 POR2X1_750/B PAND2X1_178/O 0.05fF
C6830 POR2X1_66/B PAND2X1_697/CTRL2 0.12fF
C6831 PAND2X1_787/O POR2X1_7/B 0.15fF
C6832 PAND2X1_573/B POR2X1_816/A 0.00fF
C6833 PAND2X1_192/Y PAND2X1_191/CTRL 0.01fF
C6834 POR2X1_330/Y PAND2X1_369/a_76_28# 0.05fF
C6835 POR2X1_585/Y PAND2X1_69/A 0.01fF
C6836 POR2X1_539/A PAND2X1_93/B 0.03fF
C6837 POR2X1_634/CTRL POR2X1_391/Y 0.07fF
C6838 GATE_741 PAND2X1_730/B 0.06fF
C6839 POR2X1_519/a_16_28# PAND2X1_838/B 0.02fF
C6840 POR2X1_78/A POR2X1_540/A 0.03fF
C6841 PAND2X1_479/A VDD -0.00fF
C6842 PAND2X1_592/CTRL2 VDD -0.00fF
C6843 POR2X1_460/A PAND2X1_11/Y 0.01fF
C6844 POR2X1_93/A POR2X1_225/O 0.09fF
C6845 POR2X1_646/Y POR2X1_784/a_16_28# 0.03fF
C6846 POR2X1_417/Y PAND2X1_357/Y 0.01fF
C6847 POR2X1_278/A POR2X1_32/A 0.15fF
C6848 POR2X1_776/A POR2X1_566/CTRL 0.01fF
C6849 PAND2X1_658/A PAND2X1_474/A 0.12fF
C6850 POR2X1_106/O POR2X1_387/Y 0.05fF
C6851 POR2X1_54/CTRL2 POR2X1_54/Y 0.13fF
C6852 POR2X1_293/Y POR2X1_236/Y 0.10fF
C6853 POR2X1_834/Y PAND2X1_591/CTRL2 0.16fF
C6854 PAND2X1_387/CTRL POR2X1_712/Y 0.02fF
C6855 PAND2X1_129/O PAND2X1_90/A 0.04fF
C6856 PAND2X1_641/O POR2X1_23/Y 0.05fF
C6857 POR2X1_65/A PAND2X1_551/Y 0.07fF
C6858 PAND2X1_341/B POR2X1_20/B 0.03fF
C6859 PAND2X1_220/Y PAND2X1_566/Y 0.23fF
C6860 POR2X1_528/Y POR2X1_32/A 0.03fF
C6861 PAND2X1_6/Y PAND2X1_423/CTRL 0.01fF
C6862 POR2X1_43/B PAND2X1_276/CTRL2 0.00fF
C6863 POR2X1_648/Y POR2X1_779/CTRL2 0.01fF
C6864 POR2X1_390/B D_INPUT_0 0.03fF
C6865 POR2X1_13/A PAND2X1_364/B 0.02fF
C6866 POR2X1_566/A PAND2X1_176/CTRL 0.01fF
C6867 PAND2X1_480/B POR2X1_7/B 0.05fF
C6868 POR2X1_539/A POR2X1_78/A 0.03fF
C6869 POR2X1_88/Y PAND2X1_341/CTRL2 0.00fF
C6870 PAND2X1_429/Y INPUT_5 0.04fF
C6871 PAND2X1_115/a_76_28# PAND2X1_787/Y 0.03fF
C6872 INPUT_0 POR2X1_294/B 1.78fF
C6873 POR2X1_96/A POR2X1_372/Y 0.03fF
C6874 POR2X1_278/Y POR2X1_680/Y 0.03fF
C6875 POR2X1_495/Y VDD 0.01fF
C6876 POR2X1_20/B PAND2X1_352/Y 0.05fF
C6877 POR2X1_865/B POR2X1_474/m4_208_n4# 0.15fF
C6878 PAND2X1_48/B POR2X1_215/O 0.01fF
C6879 POR2X1_88/Y POR2X1_55/Y 0.05fF
C6880 PAND2X1_474/A POR2X1_73/Y 0.03fF
C6881 POR2X1_754/A POR2X1_7/B 0.00fF
C6882 POR2X1_275/O POR2X1_46/Y 0.26fF
C6883 PAND2X1_23/Y POR2X1_76/Y 1.73fF
C6884 POR2X1_72/B POR2X1_239/Y 0.03fF
C6885 POR2X1_81/Y POR2X1_293/Y 0.00fF
C6886 POR2X1_260/B PAND2X1_48/A 0.94fF
C6887 POR2X1_383/A POR2X1_643/A 0.05fF
C6888 POR2X1_57/A GATE_479 0.03fF
C6889 POR2X1_68/A POR2X1_215/CTRL2 0.01fF
C6890 PAND2X1_734/O POR2X1_5/Y 0.03fF
C6891 POR2X1_496/Y PAND2X1_507/CTRL2 0.04fF
C6892 PAND2X1_267/CTRL2 POR2X1_7/Y 0.01fF
C6893 PAND2X1_219/B POR2X1_591/Y 0.03fF
C6894 PAND2X1_197/O PAND2X1_364/B 0.05fF
C6895 POR2X1_474/CTRL POR2X1_101/Y 0.18fF
C6896 POR2X1_255/O PAND2X1_349/A 0.01fF
C6897 POR2X1_567/B POR2X1_566/O 0.16fF
C6898 PAND2X1_94/A PAND2X1_58/A 0.11fF
C6899 POR2X1_271/A POR2X1_271/a_16_28# 0.05fF
C6900 POR2X1_528/Y POR2X1_419/Y 0.09fF
C6901 POR2X1_186/Y POR2X1_736/a_56_344# 0.00fF
C6902 PAND2X1_289/CTRL2 POR2X1_568/B 0.03fF
C6903 POR2X1_857/B POR2X1_785/A 0.42fF
C6904 POR2X1_43/B PAND2X1_785/Y 0.10fF
C6905 PAND2X1_349/A PAND2X1_141/a_16_344# 0.01fF
C6906 POR2X1_502/A PAND2X1_95/a_76_28# 0.01fF
C6907 PAND2X1_817/O POR2X1_750/Y 0.08fF
C6908 POR2X1_537/O POR2X1_590/A 0.00fF
C6909 POR2X1_72/B POR2X1_511/a_16_28# 0.02fF
C6910 POR2X1_502/A POR2X1_712/Y 0.07fF
C6911 POR2X1_78/B POR2X1_243/O 0.03fF
C6912 PAND2X1_65/B PAND2X1_314/a_16_344# 0.01fF
C6913 POR2X1_57/A POR2X1_485/O 0.02fF
C6914 PAND2X1_651/Y PAND2X1_573/CTRL 0.01fF
C6915 PAND2X1_217/B PAND2X1_723/A 0.00fF
C6916 POR2X1_8/Y POR2X1_14/Y 0.13fF
C6917 PAND2X1_23/Y POR2X1_740/Y 0.27fF
C6918 POR2X1_16/A POR2X1_69/A 0.69fF
C6919 POR2X1_70/CTRL POR2X1_90/Y 0.00fF
C6920 POR2X1_355/B POR2X1_351/Y 0.01fF
C6921 POR2X1_66/B POR2X1_61/O 0.17fF
C6922 POR2X1_383/A POR2X1_807/A 0.03fF
C6923 POR2X1_61/Y POR2X1_222/A 0.02fF
C6924 POR2X1_814/B POR2X1_218/CTRL2 0.11fF
C6925 POR2X1_590/A POR2X1_186/B 2.36fF
C6926 PAND2X1_700/CTRL2 PAND2X1_60/B 0.01fF
C6927 POR2X1_669/B PAND2X1_123/Y 0.00fF
C6928 PAND2X1_631/O POR2X1_625/Y 0.12fF
C6929 POR2X1_186/Y PAND2X1_172/CTRL2 0.01fF
C6930 PAND2X1_244/B PAND2X1_474/A 0.03fF
C6931 POR2X1_516/Y POR2X1_153/Y 0.03fF
C6932 POR2X1_347/B PAND2X1_69/O 0.01fF
C6933 POR2X1_296/B PAND2X1_527/CTRL 0.00fF
C6934 POR2X1_65/A PAND2X1_633/Y 0.06fF
C6935 POR2X1_57/A PAND2X1_719/O 0.01fF
C6936 PAND2X1_625/CTRL2 POR2X1_741/Y 0.14fF
C6937 PAND2X1_625/O POR2X1_740/Y 0.13fF
C6938 POR2X1_232/Y POR2X1_293/Y 0.06fF
C6939 PAND2X1_90/A PAND2X1_316/O 0.05fF
C6940 POR2X1_32/A POR2X1_117/Y 0.00fF
C6941 POR2X1_49/Y PAND2X1_477/A 0.02fF
C6942 POR2X1_853/A D_GATE_222 0.12fF
C6943 PAND2X1_512/Y POR2X1_387/Y 0.07fF
C6944 INPUT_0 PAND2X1_111/B 0.03fF
C6945 PAND2X1_188/CTRL POR2X1_816/A 0.01fF
C6946 PAND2X1_866/A PAND2X1_866/O 0.00fF
C6947 POR2X1_481/Y PAND2X1_566/Y 0.03fF
C6948 PAND2X1_56/Y POR2X1_140/B 0.05fF
C6949 POR2X1_833/CTRL POR2X1_786/Y 0.06fF
C6950 POR2X1_29/A POR2X1_171/Y 0.02fF
C6951 PAND2X1_8/CTRL INPUT_2 0.05fF
C6952 POR2X1_346/B POR2X1_555/A 0.03fF
C6953 POR2X1_278/A PAND2X1_35/Y 0.00fF
C6954 POR2X1_802/CTRL POR2X1_435/Y 0.07fF
C6955 PAND2X1_213/A PAND2X1_161/Y 0.00fF
C6956 PAND2X1_6/Y PAND2X1_273/O 0.15fF
C6957 PAND2X1_370/CTRL2 PAND2X1_566/Y 0.00fF
C6958 PAND2X1_726/B POR2X1_763/A 0.22fF
C6959 POR2X1_41/a_16_28# POR2X1_40/Y 0.08fF
C6960 POR2X1_573/O POR2X1_456/B 0.01fF
C6961 INPUT_1 POR2X1_627/CTRL 0.00fF
C6962 PAND2X1_82/Y POR2X1_402/B 0.01fF
C6963 PAND2X1_717/Y INPUT_0 0.03fF
C6964 POR2X1_775/A POR2X1_112/Y 0.56fF
C6965 PAND2X1_633/CTRL POR2X1_153/Y 0.05fF
C6966 POR2X1_242/CTRL2 POR2X1_192/B 0.17fF
C6967 POR2X1_297/Y PAND2X1_346/Y 0.00fF
C6968 POR2X1_523/Y D_INPUT_1 0.03fF
C6969 POR2X1_356/A PAND2X1_60/B 0.05fF
C6970 PAND2X1_807/a_56_28# POR2X1_7/B 0.00fF
C6971 PAND2X1_563/a_76_28# PAND2X1_566/Y 0.03fF
C6972 POR2X1_264/Y POR2X1_532/A 0.03fF
C6973 POR2X1_62/Y POR2X1_40/Y 0.06fF
C6974 POR2X1_383/A PAND2X1_386/Y 0.01fF
C6975 POR2X1_687/B POR2X1_729/Y 0.01fF
C6976 POR2X1_131/Y VDD 0.02fF
C6977 POR2X1_7/A POR2X1_372/Y 0.04fF
C6978 POR2X1_532/A POR2X1_710/CTRL2 0.01fF
C6979 PAND2X1_90/Y POR2X1_209/CTRL2 0.01fF
C6980 POR2X1_66/B POR2X1_99/B 0.03fF
C6981 POR2X1_83/CTRL PAND2X1_734/B 0.01fF
C6982 POR2X1_57/A POR2X1_396/CTRL2 0.03fF
C6983 PAND2X1_55/Y POR2X1_537/B 0.07fF
C6984 POR2X1_41/B PAND2X1_569/B 0.07fF
C6985 PAND2X1_6/Y POR2X1_840/B 0.03fF
C6986 POR2X1_462/B PAND2X1_69/A 0.04fF
C6987 POR2X1_614/A POR2X1_542/B 0.03fF
C6988 D_INPUT_1 PAND2X1_69/A 0.13fF
C6989 PAND2X1_23/Y POR2X1_348/O 0.05fF
C6990 PAND2X1_686/CTRL POR2X1_13/A 0.01fF
C6991 PAND2X1_206/CTRL2 POR2X1_153/Y 0.12fF
C6992 PAND2X1_96/B POR2X1_576/Y 0.00fF
C6993 POR2X1_614/A PAND2X1_79/Y 0.07fF
C6994 POR2X1_596/A POR2X1_770/CTRL2 0.01fF
C6995 POR2X1_93/A POR2X1_816/A 0.03fF
C6996 PAND2X1_90/Y POR2X1_652/A 0.07fF
C6997 POR2X1_68/A POR2X1_348/CTRL 0.29fF
C6998 POR2X1_43/B PAND2X1_656/A 0.08fF
C6999 POR2X1_816/A POR2X1_91/Y 0.03fF
C7000 PAND2X1_414/CTRL POR2X1_67/Y 0.01fF
C7001 POR2X1_8/Y PAND2X1_472/B 0.07fF
C7002 PAND2X1_69/A POR2X1_724/A 0.15fF
C7003 POR2X1_619/O POR2X1_283/A 0.07fF
C7004 PAND2X1_598/CTRL2 POR2X1_394/A 0.05fF
C7005 POR2X1_804/A POR2X1_318/A 0.10fF
C7006 PAND2X1_430/CTRL PAND2X1_3/B 0.01fF
C7007 POR2X1_83/A POR2X1_235/Y 0.03fF
C7008 POR2X1_35/Y POR2X1_222/A 0.01fF
C7009 PAND2X1_632/B POR2X1_42/Y 0.03fF
C7010 PAND2X1_803/Y POR2X1_90/Y 0.01fF
C7011 POR2X1_356/A POR2X1_353/A 0.05fF
C7012 POR2X1_407/A POR2X1_383/A 0.11fF
C7013 POR2X1_253/Y POR2X1_7/A 0.00fF
C7014 POR2X1_16/A PAND2X1_462/B 0.02fF
C7015 POR2X1_43/B PAND2X1_124/CTRL2 0.01fF
C7016 POR2X1_333/Y POR2X1_776/B 0.03fF
C7017 POR2X1_528/Y PAND2X1_651/Y 0.00fF
C7018 POR2X1_8/Y POR2X1_55/Y 0.12fF
C7019 POR2X1_51/O INPUT_7 0.17fF
C7020 POR2X1_57/A POR2X1_142/Y 0.03fF
C7021 POR2X1_57/a_16_28# PAND2X1_737/B 0.01fF
C7022 PAND2X1_474/Y POR2X1_150/O 0.00fF
C7023 POR2X1_271/A POR2X1_293/Y 0.02fF
C7024 PAND2X1_714/A PAND2X1_169/CTRL2 0.01fF
C7025 D_GATE_741 POR2X1_260/A 0.09fF
C7026 POR2X1_16/A POR2X1_437/Y 0.03fF
C7027 POR2X1_366/O PAND2X1_6/Y 0.18fF
C7028 POR2X1_685/A POR2X1_685/B 0.02fF
C7029 POR2X1_43/B POR2X1_754/O 0.03fF
C7030 POR2X1_123/A PAND2X1_518/a_16_344# 0.01fF
C7031 PAND2X1_608/O POR2X1_411/B 0.01fF
C7032 POR2X1_557/A POR2X1_78/O 0.01fF
C7033 POR2X1_93/m4_208_n4# PAND2X1_509/m4_208_n4# 0.13fF
C7034 POR2X1_532/A PAND2X1_528/CTRL 0.01fF
C7035 POR2X1_416/B POR2X1_24/CTRL 0.25fF
C7036 POR2X1_110/Y POR2X1_693/O 0.37fF
C7037 PAND2X1_865/Y PAND2X1_579/B 0.00fF
C7038 POR2X1_72/B PAND2X1_861/B 0.05fF
C7039 POR2X1_43/B PAND2X1_348/A 0.07fF
C7040 POR2X1_96/A PAND2X1_858/a_76_28# 0.01fF
C7041 PAND2X1_94/A PAND2X1_96/B 9.82fF
C7042 PAND2X1_727/CTRL POR2X1_90/Y 0.01fF
C7043 POR2X1_334/B POR2X1_557/B 0.07fF
C7044 POR2X1_510/B PAND2X1_824/O 0.01fF
C7045 POR2X1_493/a_16_28# PAND2X1_60/B 0.02fF
C7046 PAND2X1_714/Y POR2X1_73/Y 0.10fF
C7047 POR2X1_5/Y POR2X1_39/B 0.13fF
C7048 POR2X1_554/B POR2X1_116/A 0.03fF
C7049 POR2X1_3/CTRL2 POR2X1_260/A 0.05fF
C7050 POR2X1_569/A PAND2X1_60/B 0.21fF
C7051 PAND2X1_23/Y PAND2X1_171/O 0.03fF
C7052 POR2X1_760/A PAND2X1_217/CTRL 0.03fF
C7053 PAND2X1_55/Y PAND2X1_48/A 0.28fF
C7054 POR2X1_246/Y POR2X1_248/Y 0.04fF
C7055 PAND2X1_9/Y POR2X1_623/Y 0.01fF
C7056 PAND2X1_631/A POR2X1_252/CTRL 0.01fF
C7057 POR2X1_39/Y POR2X1_73/Y 0.02fF
C7058 POR2X1_334/Y POR2X1_562/B 0.03fF
C7059 POR2X1_438/CTRL2 POR2X1_373/Y 0.00fF
C7060 POR2X1_804/A POR2X1_574/Y 0.03fF
C7061 PAND2X1_549/CTRL2 POR2X1_39/B 0.00fF
C7062 POR2X1_556/A POR2X1_658/a_76_344# 0.00fF
C7063 POR2X1_416/B POR2X1_290/a_16_28# 0.01fF
C7064 POR2X1_124/B POR2X1_557/B 0.03fF
C7065 POR2X1_41/B POR2X1_316/Y 0.07fF
C7066 PAND2X1_545/Y PAND2X1_854/A 0.00fF
C7067 POR2X1_158/Y PAND2X1_712/O 0.00fF
C7068 PAND2X1_294/CTRL POR2X1_150/Y 0.04fF
C7069 POR2X1_730/Y POR2X1_855/B 0.00fF
C7070 POR2X1_327/Y POR2X1_865/B 0.04fF
C7071 POR2X1_150/Y PAND2X1_211/O 0.17fF
C7072 POR2X1_505/O POR2X1_245/Y 0.01fF
C7073 POR2X1_760/A PAND2X1_267/Y 0.08fF
C7074 PAND2X1_464/B PAND2X1_776/Y 0.02fF
C7075 POR2X1_57/A PAND2X1_156/B 0.15fF
C7076 PAND2X1_631/A POR2X1_43/B 0.23fF
C7077 POR2X1_119/Y POR2X1_234/O 0.13fF
C7078 PAND2X1_69/A POR2X1_620/B 0.67fF
C7079 POR2X1_407/Y PAND2X1_48/A 0.08fF
C7080 POR2X1_728/CTRL PAND2X1_52/B 0.00fF
C7081 POR2X1_294/B POR2X1_510/CTRL 0.01fF
C7082 PAND2X1_217/B PAND2X1_860/A 0.05fF
C7083 POR2X1_150/Y POR2X1_437/O 0.02fF
C7084 POR2X1_240/A POR2X1_66/A 0.02fF
C7085 POR2X1_257/A POR2X1_582/Y 0.01fF
C7086 POR2X1_571/O POR2X1_569/A 0.04fF
C7087 POR2X1_20/B POR2X1_298/CTRL 0.01fF
C7088 POR2X1_802/B POR2X1_532/a_16_28# 0.05fF
C7089 PAND2X1_341/A PAND2X1_101/B 0.01fF
C7090 POR2X1_52/A POR2X1_158/Y 0.00fF
C7091 PAND2X1_859/B POR2X1_77/Y 0.03fF
C7092 POR2X1_760/A POR2X1_674/a_16_28# 0.00fF
C7093 PAND2X1_434/CTRL2 POR2X1_129/Y 0.01fF
C7094 POR2X1_643/a_16_28# POR2X1_643/A 0.01fF
C7095 PAND2X1_409/CTRL PAND2X1_52/B 0.11fF
C7096 POR2X1_740/Y POR2X1_711/Y 0.00fF
C7097 PAND2X1_242/Y POR2X1_236/Y 3.42fF
C7098 POR2X1_43/CTRL POR2X1_43/B 0.01fF
C7099 PAND2X1_174/O POR2X1_77/Y 0.09fF
C7100 POR2X1_499/CTRL2 POR2X1_341/A 0.02fF
C7101 POR2X1_43/B POR2X1_589/a_16_28# 0.02fF
C7102 POR2X1_738/A POR2X1_726/CTRL 0.01fF
C7103 PAND2X1_860/A VDD 0.69fF
C7104 POR2X1_454/a_16_28# POR2X1_454/A 0.03fF
C7105 POR2X1_811/CTRL PAND2X1_39/B 0.02fF
C7106 POR2X1_709/B PAND2X1_698/O 0.00fF
C7107 POR2X1_287/A POR2X1_121/B 0.03fF
C7108 POR2X1_326/A POR2X1_675/Y 0.03fF
C7109 PAND2X1_644/Y POR2X1_600/Y 0.03fF
C7110 POR2X1_228/O POR2X1_260/A 0.01fF
C7111 POR2X1_703/A POR2X1_703/O 0.14fF
C7112 POR2X1_158/a_16_28# POR2X1_425/Y 0.01fF
C7113 POR2X1_607/A POR2X1_411/A 0.00fF
C7114 POR2X1_460/Y PAND2X1_58/A 0.04fF
C7115 POR2X1_624/Y POR2X1_66/A 0.07fF
C7116 PAND2X1_10/a_16_344# PAND2X1_9/Y 0.01fF
C7117 POR2X1_703/A POR2X1_337/Y 0.09fF
C7118 POR2X1_16/A POR2X1_599/a_16_28# -0.01fF
C7119 PAND2X1_632/B POR2X1_252/Y 0.02fF
C7120 POR2X1_532/A POR2X1_532/a_16_28# 0.04fF
C7121 POR2X1_648/Y POR2X1_807/A 0.03fF
C7122 POR2X1_343/Y POR2X1_532/A 0.11fF
C7123 POR2X1_768/O POR2X1_294/A 0.03fF
C7124 POR2X1_326/A POR2X1_544/B 0.00fF
C7125 POR2X1_7/B POR2X1_386/Y 0.01fF
C7126 PAND2X1_404/Y POR2X1_263/Y 0.03fF
C7127 POR2X1_461/a_16_28# POR2X1_814/A 0.03fF
C7128 POR2X1_576/a_56_344# POR2X1_572/Y 0.01fF
C7129 POR2X1_513/Y POR2X1_717/B 0.03fF
C7130 POR2X1_54/Y PAND2X1_37/O 0.02fF
C7131 D_INPUT_3 POR2X1_416/B 0.03fF
C7132 POR2X1_333/Y POR2X1_192/B 0.03fF
C7133 PAND2X1_341/Y POR2X1_4/Y 0.03fF
C7134 POR2X1_129/Y PAND2X1_851/CTRL 0.01fF
C7135 POR2X1_188/A POR2X1_841/CTRL2 0.01fF
C7136 PAND2X1_66/CTRL POR2X1_67/A 0.03fF
C7137 POR2X1_159/O INPUT_3 0.24fF
C7138 POR2X1_68/A POR2X1_303/B 0.05fF
C7139 PAND2X1_841/O POR2X1_677/Y -0.00fF
C7140 POR2X1_817/O POR2X1_32/A 0.02fF
C7141 POR2X1_736/A POR2X1_737/CTRL2 0.23fF
C7142 PAND2X1_265/CTRL POR2X1_260/B 0.01fF
C7143 POR2X1_54/Y PAND2X1_817/a_76_28# 0.03fF
C7144 PAND2X1_60/B PAND2X1_72/A 12.91fF
C7145 PAND2X1_771/B VDD 0.17fF
C7146 PAND2X1_569/B POR2X1_77/Y 0.08fF
C7147 POR2X1_113/CTRL POR2X1_768/A 0.02fF
C7148 POR2X1_298/Y POR2X1_299/Y 0.01fF
C7149 POR2X1_544/a_16_28# PAND2X1_52/B 0.02fF
C7150 PAND2X1_6/Y POR2X1_661/A 0.07fF
C7151 POR2X1_191/a_16_28# POR2X1_444/Y 0.03fF
C7152 POR2X1_39/a_16_28# POR2X1_38/Y 0.05fF
C7153 PAND2X1_65/B POR2X1_663/B 0.03fF
C7154 PAND2X1_789/CTRL POR2X1_39/B 0.01fF
C7155 POR2X1_568/B POR2X1_317/B 0.03fF
C7156 POR2X1_337/Y PAND2X1_167/CTRL2 0.01fF
C7157 POR2X1_20/B POR2X1_497/Y 0.02fF
C7158 POR2X1_544/B POR2X1_374/a_16_28# 0.03fF
C7159 POR2X1_261/A POR2X1_411/B 0.00fF
C7160 PAND2X1_97/Y PAND2X1_351/CTRL 0.01fF
C7161 POR2X1_23/Y POR2X1_49/CTRL2 0.01fF
C7162 PAND2X1_779/CTRL2 POR2X1_39/B 0.00fF
C7163 PAND2X1_206/B PAND2X1_341/O 0.00fF
C7164 POR2X1_609/Y PAND2X1_404/O 0.00fF
C7165 PAND2X1_39/B POR2X1_403/Y 0.01fF
C7166 POR2X1_96/A POR2X1_485/Y 0.23fF
C7167 PAND2X1_85/Y POR2X1_243/B 0.01fF
C7168 POR2X1_774/A POR2X1_711/Y 0.03fF
C7169 POR2X1_667/A POR2X1_32/A 0.04fF
C7170 POR2X1_34/B POR2X1_34/Y 0.02fF
C7171 D_INPUT_5 POR2X1_25/O 0.03fF
C7172 PAND2X1_72/A POR2X1_353/A 0.03fF
C7173 POR2X1_56/B PAND2X1_466/A 0.02fF
C7174 PAND2X1_798/Y PAND2X1_366/a_56_28# 0.00fF
C7175 PAND2X1_487/a_16_344# POR2X1_287/B 0.01fF
C7176 PAND2X1_432/a_76_28# POR2X1_866/A 0.03fF
C7177 POR2X1_41/B POR2X1_603/O 0.35fF
C7178 PAND2X1_72/A POR2X1_332/O 0.17fF
C7179 POR2X1_304/a_16_28# PAND2X1_454/B 0.02fF
C7180 POR2X1_647/B VDD 0.46fF
C7181 PAND2X1_58/A PAND2X1_11/Y 0.01fF
C7182 POR2X1_407/A POR2X1_648/Y 0.06fF
C7183 POR2X1_67/CTRL POR2X1_236/Y 0.09fF
C7184 POR2X1_366/Y PAND2X1_417/O 0.11fF
C7185 PAND2X1_58/A POR2X1_606/Y 0.84fF
C7186 POR2X1_864/A POR2X1_828/O 0.00fF
C7187 POR2X1_502/A PAND2X1_39/B 0.10fF
C7188 PAND2X1_205/O PAND2X1_473/B 0.04fF
C7189 PAND2X1_39/B POR2X1_783/A 0.02fF
C7190 POR2X1_23/Y POR2X1_278/O 0.01fF
C7191 POR2X1_255/O POR2X1_32/A 0.02fF
C7192 PAND2X1_48/B POR2X1_556/A 2.77fF
C7193 POR2X1_274/Y D_INPUT_0 0.31fF
C7194 POR2X1_48/A POR2X1_5/Y 0.15fF
C7195 POR2X1_210/A PAND2X1_52/B 0.09fF
C7196 POR2X1_41/B POR2X1_54/Y 0.05fF
C7197 POR2X1_260/B PAND2X1_378/CTRL2 0.03fF
C7198 POR2X1_776/A POR2X1_579/Y 0.03fF
C7199 POR2X1_644/CTRL2 PAND2X1_57/B 0.00fF
C7200 PAND2X1_839/O POR2X1_411/B 0.03fF
C7201 PAND2X1_331/a_56_28# POR2X1_330/Y 0.00fF
C7202 POR2X1_49/Y POR2X1_422/Y 4.14fF
C7203 POR2X1_241/B POR2X1_254/O 0.02fF
C7204 PAND2X1_341/B POR2X1_86/Y 0.01fF
C7205 POR2X1_275/a_16_28# POR2X1_275/A 0.01fF
C7206 PAND2X1_8/O INPUT_3 0.13fF
C7207 PAND2X1_608/a_76_28# POR2X1_73/Y 0.02fF
C7208 POR2X1_729/CTRL2 POR2X1_452/Y 0.01fF
C7209 PAND2X1_787/A PAND2X1_717/A 0.07fF
C7210 POR2X1_157/O POR2X1_257/A 0.01fF
C7211 POR2X1_434/A POR2X1_480/A 0.21fF
C7212 POR2X1_257/A PAND2X1_707/Y 0.01fF
C7213 INPUT_1 PAND2X1_54/a_76_28# 0.01fF
C7214 POR2X1_227/A PAND2X1_32/B 0.03fF
C7215 POR2X1_730/Y POR2X1_440/O 0.01fF
C7216 POR2X1_32/A PAND2X1_712/B 0.01fF
C7217 POR2X1_566/A PAND2X1_258/CTRL 0.13fF
C7218 PAND2X1_23/Y PAND2X1_67/O 0.03fF
C7219 POR2X1_523/Y INPUT_3 0.84fF
C7220 PAND2X1_404/Y PAND2X1_215/B 0.03fF
C7221 POR2X1_270/Y POR2X1_220/Y 0.03fF
C7222 PAND2X1_459/O POR2X1_750/B 0.06fF
C7223 PAND2X1_216/CTRL PAND2X1_218/B 0.01fF
C7224 POR2X1_257/A PAND2X1_798/B 0.03fF
C7225 POR2X1_609/Y PAND2X1_404/A 1.17fF
C7226 POR2X1_316/Y POR2X1_77/Y 0.03fF
C7227 POR2X1_29/CTRL POR2X1_29/A 0.01fF
C7228 POR2X1_66/B POR2X1_504/Y 0.14fF
C7229 PAND2X1_211/CTRL PAND2X1_357/Y 0.01fF
C7230 PAND2X1_96/B PAND2X1_43/CTRL2 0.02fF
C7231 INPUT_1 POR2X1_624/CTRL 0.01fF
C7232 POR2X1_831/O POR2X1_804/A 0.31fF
C7233 POR2X1_78/A POR2X1_608/CTRL 0.03fF
C7234 PAND2X1_73/Y POR2X1_608/O 0.10fF
C7235 INPUT_3 PAND2X1_69/A 0.07fF
C7236 POR2X1_102/Y POR2X1_760/O 0.01fF
C7237 POR2X1_130/A POR2X1_296/B 0.10fF
C7238 PAND2X1_318/a_16_344# PAND2X1_776/Y 0.03fF
C7239 PAND2X1_661/Y POR2X1_681/O 0.04fF
C7240 POR2X1_60/A POR2X1_236/Y 3.22fF
C7241 POR2X1_856/B POR2X1_579/Y 0.03fF
C7242 PAND2X1_270/CTRL2 POR2X1_20/B 0.01fF
C7243 POR2X1_83/B POR2X1_250/CTRL 0.01fF
C7244 POR2X1_49/Y POR2X1_743/CTRL2 0.01fF
C7245 POR2X1_614/A POR2X1_676/a_56_344# 0.00fF
C7246 PAND2X1_85/CTRL POR2X1_260/A 0.00fF
C7247 POR2X1_647/B PAND2X1_32/B 0.03fF
C7248 PAND2X1_404/Y PAND2X1_6/A 0.15fF
C7249 PAND2X1_139/a_76_28# POR2X1_40/Y 0.01fF
C7250 PAND2X1_212/O PAND2X1_357/Y 0.02fF
C7251 POR2X1_66/A POR2X1_785/A 0.06fF
C7252 POR2X1_65/A POR2X1_250/A 0.01fF
C7253 INPUT_3 POR2X1_93/A 0.02fF
C7254 PAND2X1_58/A PAND2X1_56/CTRL2 0.01fF
C7255 PAND2X1_218/A PAND2X1_267/Y 0.01fF
C7256 POR2X1_147/A PAND2X1_93/B 0.01fF
C7257 POR2X1_240/CTRL2 PAND2X1_88/Y 0.01fF
C7258 POR2X1_538/CTRL2 POR2X1_66/A 0.00fF
C7259 POR2X1_624/Y POR2X1_532/A 0.18fF
C7260 POR2X1_558/a_16_28# POR2X1_260/B 0.03fF
C7261 PAND2X1_678/O PAND2X1_175/B 0.02fF
C7262 PAND2X1_839/B POR2X1_411/B 0.03fF
C7263 PAND2X1_276/a_16_344# PAND2X1_390/Y 0.01fF
C7264 POR2X1_411/B PAND2X1_348/Y 0.07fF
C7265 PAND2X1_96/B PAND2X1_406/CTRL2 0.01fF
C7266 POR2X1_502/A PAND2X1_20/A 0.08fF
C7267 POR2X1_461/A VDD 0.00fF
C7268 POR2X1_667/A PAND2X1_35/Y 0.01fF
C7269 POR2X1_814/B POR2X1_116/CTRL 0.01fF
C7270 POR2X1_159/a_16_28# POR2X1_5/Y 0.00fF
C7271 POR2X1_78/B PAND2X1_16/CTRL2 0.01fF
C7272 POR2X1_862/A POR2X1_649/CTRL 0.00fF
C7273 POR2X1_56/B POR2X1_423/O 0.02fF
C7274 POR2X1_297/Y PAND2X1_354/A 0.06fF
C7275 POR2X1_150/Y PAND2X1_130/a_16_344# 0.02fF
C7276 POR2X1_411/B PAND2X1_181/CTRL 0.01fF
C7277 PAND2X1_433/a_16_344# D_INPUT_0 0.02fF
C7278 PAND2X1_93/B POR2X1_219/CTRL2 0.00fF
C7279 POR2X1_12/A INPUT_6 0.06fF
C7280 POR2X1_719/O PAND2X1_39/B 0.05fF
C7281 POR2X1_688/CTRL POR2X1_260/A 0.01fF
C7282 PAND2X1_93/B PAND2X1_69/A 0.41fF
C7283 POR2X1_81/Y POR2X1_60/A 0.00fF
C7284 POR2X1_440/B POR2X1_186/B 0.01fF
C7285 POR2X1_614/A POR2X1_856/B 0.04fF
C7286 POR2X1_212/A POR2X1_212/CTRL 0.01fF
C7287 POR2X1_820/CTRL2 POR2X1_42/Y 0.18fF
C7288 POR2X1_269/m4_208_n4# POR2X1_740/Y 0.06fF
C7289 POR2X1_383/A PAND2X1_271/O 0.01fF
C7290 POR2X1_754/A POR2X1_750/B 0.03fF
C7291 PAND2X1_793/Y POR2X1_72/B 0.06fF
C7292 PAND2X1_792/CTRL POR2X1_759/Y 0.00fF
C7293 POR2X1_66/B POR2X1_664/Y 0.01fF
C7294 POR2X1_548/CTRL2 PAND2X1_8/Y 0.00fF
C7295 POR2X1_448/Y POR2X1_435/Y 0.07fF
C7296 PAND2X1_619/CTRL2 POR2X1_260/A 0.03fF
C7297 PAND2X1_31/O INPUT_6 0.15fF
C7298 POR2X1_356/A POR2X1_750/B 0.02fF
C7299 POR2X1_502/A POR2X1_814/B 5.85fF
C7300 POR2X1_754/Y POR2X1_90/Y 0.01fF
C7301 POR2X1_568/A POR2X1_161/O 0.10fF
C7302 POR2X1_381/a_16_28# POR2X1_236/Y 0.13fF
C7303 POR2X1_695/Y POR2X1_425/Y 0.13fF
C7304 POR2X1_590/A POR2X1_208/Y 0.01fF
C7305 INPUT_1 POR2X1_628/Y 0.03fF
C7306 POR2X1_834/Y POR2X1_648/CTRL 0.17fF
C7307 POR2X1_66/B POR2X1_775/A 0.03fF
C7308 PAND2X1_23/Y POR2X1_202/CTRL 0.00fF
C7309 POR2X1_274/O POR2X1_573/A 0.02fF
C7310 POR2X1_848/A POR2X1_283/A 0.07fF
C7311 POR2X1_814/B POR2X1_247/CTRL 0.00fF
C7312 POR2X1_78/A POR2X1_649/CTRL2 0.08fF
C7313 PAND2X1_73/Y POR2X1_644/A 0.03fF
C7314 POR2X1_78/A PAND2X1_69/A 0.58fF
C7315 POR2X1_814/B PAND2X1_176/O 0.01fF
C7316 PAND2X1_652/A POR2X1_40/Y 0.06fF
C7317 POR2X1_814/B POR2X1_464/Y 0.08fF
C7318 POR2X1_29/A PAND2X1_670/CTRL2 0.01fF
C7319 POR2X1_590/A PAND2X1_79/Y 0.09fF
C7320 POR2X1_296/B POR2X1_573/A 3.55fF
C7321 POR2X1_502/A POR2X1_325/A 0.02fF
C7322 POR2X1_760/CTRL2 POR2X1_7/B 0.01fF
C7323 POR2X1_376/B PAND2X1_174/CTRL2 0.08fF
C7324 POR2X1_676/Y VDD -0.00fF
C7325 POR2X1_68/A POR2X1_202/CTRL2 0.01fF
C7326 PAND2X1_164/CTRL2 POR2X1_776/B 0.01fF
C7327 POR2X1_255/O POR2X1_184/Y 0.03fF
C7328 POR2X1_260/B POR2X1_789/B 0.03fF
C7329 D_INPUT_0 PAND2X1_349/A 0.03fF
C7330 POR2X1_54/Y POR2X1_753/O 0.04fF
C7331 POR2X1_66/B POR2X1_112/Y 0.03fF
C7332 POR2X1_856/B POR2X1_440/Y 0.03fF
C7333 D_INPUT_0 PAND2X1_63/B 0.08fF
C7334 POR2X1_68/A PAND2X1_279/a_76_28# -0.04fF
C7335 POR2X1_688/a_16_28# POR2X1_294/A 0.00fF
C7336 POR2X1_814/A PAND2X1_122/a_16_344# 0.01fF
C7337 POR2X1_22/A POR2X1_12/CTRL 0.01fF
C7338 POR2X1_197/Y POR2X1_555/B 0.30fF
C7339 POR2X1_5/Y PAND2X1_197/Y 0.14fF
C7340 PAND2X1_453/O POR2X1_511/Y 0.08fF
C7341 POR2X1_114/B POR2X1_405/a_56_344# 0.00fF
C7342 POR2X1_178/Y POR2X1_48/A 0.00fF
C7343 POR2X1_245/Y POR2X1_32/A 0.20fF
C7344 POR2X1_684/CTRL VDD 0.00fF
C7345 PAND2X1_401/CTRL POR2X1_5/Y 0.01fF
C7346 POR2X1_83/B POR2X1_172/Y 0.05fF
C7347 POR2X1_448/CTRL PAND2X1_60/B 0.01fF
C7348 POR2X1_502/A POR2X1_513/B 0.03fF
C7349 POR2X1_16/A PAND2X1_214/O 0.01fF
C7350 POR2X1_271/CTRL POR2X1_153/Y 0.01fF
C7351 POR2X1_22/CTRL INPUT_5 0.01fF
C7352 POR2X1_355/B POR2X1_468/B 0.03fF
C7353 PAND2X1_824/B PAND2X1_93/B 0.16fF
C7354 PAND2X1_73/Y POR2X1_274/B 0.00fF
C7355 POR2X1_634/A POR2X1_711/a_76_344# 0.03fF
C7356 PAND2X1_675/a_16_344# POR2X1_250/Y 0.04fF
C7357 PAND2X1_488/CTRL POR2X1_68/B 0.01fF
C7358 POR2X1_567/B POR2X1_703/Y 0.05fF
C7359 POR2X1_325/O POR2X1_78/A 0.18fF
C7360 PAND2X1_812/CTRL2 VDD 0.00fF
C7361 POR2X1_287/B POR2X1_778/B 0.01fF
C7362 POR2X1_433/CTRL PAND2X1_549/B 0.11fF
C7363 PAND2X1_661/B POR2X1_117/CTRL2 0.03fF
C7364 POR2X1_614/Y PAND2X1_28/O 0.00fF
C7365 POR2X1_230/Y POR2X1_293/Y 0.03fF
C7366 POR2X1_388/O POR2X1_814/B 0.01fF
C7367 POR2X1_379/CTRL PAND2X1_20/A 0.00fF
C7368 POR2X1_634/A PAND2X1_764/CTRL 0.07fF
C7369 POR2X1_614/A POR2X1_786/CTRL2 0.03fF
C7370 POR2X1_516/B POR2X1_55/Y 0.02fF
C7371 PAND2X1_39/B POR2X1_188/Y 0.31fF
C7372 POR2X1_210/Y PAND2X1_41/B 0.03fF
C7373 POR2X1_220/A POR2X1_750/B 0.05fF
C7374 POR2X1_857/B POR2X1_853/CTRL 0.01fF
C7375 POR2X1_102/Y PAND2X1_717/Y 0.04fF
C7376 POR2X1_537/O POR2X1_66/A 0.05fF
C7377 POR2X1_43/B PAND2X1_715/CTRL2 0.00fF
C7378 POR2X1_197/Y POR2X1_330/Y 0.03fF
C7379 PAND2X1_568/a_56_28# POR2X1_7/B 0.00fF
C7380 POR2X1_647/CTRL POR2X1_737/A 0.01fF
C7381 POR2X1_52/A PAND2X1_592/Y 10.57fF
C7382 PAND2X1_207/O PAND2X1_123/Y 0.05fF
C7383 POR2X1_778/B POR2X1_778/CTRL 0.01fF
C7384 POR2X1_65/A PAND2X1_650/CTRL2 0.02fF
C7385 POR2X1_154/O POR2X1_803/A 0.01fF
C7386 POR2X1_332/B PAND2X1_111/CTRL 0.01fF
C7387 PAND2X1_95/B PAND2X1_409/CTRL 0.02fF
C7388 POR2X1_201/O POR2X1_201/Y 0.01fF
C7389 POR2X1_210/Y POR2X1_781/A 0.07fF
C7390 POR2X1_23/Y PAND2X1_508/Y 0.07fF
C7391 POR2X1_41/B POR2X1_13/Y 0.00fF
C7392 POR2X1_853/CTRL2 POR2X1_795/B 0.01fF
C7393 POR2X1_66/A POR2X1_186/B 0.13fF
C7394 POR2X1_130/A POR2X1_267/Y 0.03fF
C7395 INPUT_0 POR2X1_56/Y 0.07fF
C7396 POR2X1_119/Y PAND2X1_404/Y 0.02fF
C7397 POR2X1_616/Y PAND2X1_66/CTRL 0.01fF
C7398 POR2X1_389/m4_208_n4# POR2X1_130/A 0.03fF
C7399 PAND2X1_844/a_16_344# D_INPUT_0 0.04fF
C7400 PAND2X1_842/O PAND2X1_389/Y 0.01fF
C7401 POR2X1_131/O PAND2X1_140/Y 0.01fF
C7402 POR2X1_750/B POR2X1_569/A 0.10fF
C7403 POR2X1_804/A PAND2X1_131/O 0.15fF
C7404 PAND2X1_48/B PAND2X1_751/m4_208_n4# 0.08fF
C7405 POR2X1_203/Y VDD 0.18fF
C7406 PAND2X1_819/CTRL POR2X1_750/B 0.03fF
C7407 POR2X1_78/B POR2X1_596/A 0.19fF
C7408 POR2X1_40/O POR2X1_40/Y 0.01fF
C7409 POR2X1_614/A POR2X1_722/Y 0.03fF
C7410 POR2X1_740/Y POR2X1_733/A 0.07fF
C7411 PAND2X1_6/CTRL2 POR2X1_35/B 0.01fF
C7412 POR2X1_807/a_16_28# PAND2X1_48/A 0.01fF
C7413 POR2X1_166/CTRL PAND2X1_738/Y 0.01fF
C7414 POR2X1_724/CTRL2 POR2X1_724/A 0.01fF
C7415 POR2X1_725/a_16_28# POR2X1_712/Y -0.00fF
C7416 PAND2X1_663/CTRL2 PAND2X1_660/B 0.01fF
C7417 POR2X1_83/A POR2X1_42/Y 0.59fF
C7418 POR2X1_271/A POR2X1_60/A 0.06fF
C7419 POR2X1_186/Y POR2X1_151/O 0.03fF
C7420 PAND2X1_232/O PAND2X1_41/B 0.03fF
C7421 PAND2X1_854/A PAND2X1_539/B 0.25fF
C7422 PAND2X1_472/B POR2X1_68/B 0.02fF
C7423 PAND2X1_803/O POR2X1_60/A 0.18fF
C7424 POR2X1_108/Y POR2X1_106/Y 0.02fF
C7425 POR2X1_477/O PAND2X1_52/B 0.02fF
C7426 POR2X1_543/A POR2X1_703/A 0.58fF
C7427 POR2X1_16/A POR2X1_127/Y 0.13fF
C7428 POR2X1_344/A POR2X1_205/A 0.19fF
C7429 PAND2X1_604/CTRL2 PAND2X1_69/A 0.01fF
C7430 POR2X1_235/Y POR2X1_230/a_16_28# 0.00fF
C7431 POR2X1_730/Y POR2X1_439/Y 0.00fF
C7432 PAND2X1_79/CTRL2 POR2X1_844/B 0.02fF
C7433 POR2X1_208/Y POR2X1_214/B 0.09fF
C7434 PAND2X1_733/A POR2X1_394/A -0.05fF
C7435 POR2X1_96/A PAND2X1_344/O 0.05fF
C7436 POR2X1_494/Y POR2X1_73/Y 0.03fF
C7437 PAND2X1_202/CTRL2 POR2X1_7/A 0.01fF
C7438 POR2X1_41/B PAND2X1_270/CTRL 0.07fF
C7439 POR2X1_90/Y POR2X1_42/Y 0.18fF
C7440 POR2X1_41/B PAND2X1_787/A 0.03fF
C7441 POR2X1_467/Y POR2X1_210/A 0.04fF
C7442 POR2X1_377/CTRL D_INPUT_1 0.01fF
C7443 POR2X1_86/CTRL2 D_INPUT_0 0.01fF
C7444 POR2X1_27/CTRL2 POR2X1_9/Y 0.01fF
C7445 PAND2X1_496/a_16_344# D_INPUT_1 0.01fF
C7446 POR2X1_155/Y POR2X1_162/Y 0.01fF
C7447 POR2X1_738/A VDD -0.00fF
C7448 POR2X1_532/A POR2X1_785/A 0.03fF
C7449 PAND2X1_752/Y POR2X1_459/A 0.23fF
C7450 POR2X1_68/B POR2X1_55/Y 0.00fF
C7451 PAND2X1_318/CTRL PAND2X1_787/A 0.01fF
C7452 POR2X1_707/a_16_28# PAND2X1_41/B 0.02fF
C7453 PAND2X1_523/a_76_28# POR2X1_522/Y 0.02fF
C7454 PAND2X1_252/O POR2X1_222/Y 0.01fF
C7455 POR2X1_832/a_16_28# POR2X1_832/A 0.03fF
C7456 POR2X1_7/B POR2X1_239/Y 0.76fF
C7457 POR2X1_555/A POR2X1_507/A 0.03fF
C7458 PAND2X1_810/CTRL VDD 0.00fF
C7459 POR2X1_54/Y POR2X1_8/O 0.01fF
C7460 POR2X1_566/A POR2X1_507/CTRL 0.15fF
C7461 POR2X1_501/O POR2X1_573/A 0.02fF
C7462 PAND2X1_41/B POR2X1_195/CTRL 0.01fF
C7463 POR2X1_272/Y PAND2X1_301/O 0.02fF
C7464 PAND2X1_390/Y PAND2X1_716/B 0.03fF
C7465 PAND2X1_664/CTRL PAND2X1_645/B 0.04fF
C7466 PAND2X1_220/CTRL PAND2X1_388/Y 0.01fF
C7467 PAND2X1_69/A PAND2X1_145/a_76_28# 0.01fF
C7468 POR2X1_66/A PAND2X1_529/a_16_344# 0.01fF
C7469 POR2X1_860/A PAND2X1_48/A 0.03fF
C7470 PAND2X1_216/O PAND2X1_723/A 0.00fF
C7471 POR2X1_730/Y POR2X1_192/Y 0.01fF
C7472 POR2X1_40/Y PAND2X1_506/Y 0.01fF
C7473 PAND2X1_57/B POR2X1_456/B 0.06fF
C7474 POR2X1_65/A POR2X1_103/m4_208_n4# 0.07fF
C7475 POR2X1_101/Y POR2X1_404/Y 4.06fF
C7476 POR2X1_407/A POR2X1_780/A 0.05fF
C7477 POR2X1_722/B POR2X1_796/A 0.04fF
C7478 PAND2X1_6/Y POR2X1_686/CTRL 0.08fF
C7479 PAND2X1_713/O PAND2X1_713/B 0.01fF
C7480 POR2X1_365/Y POR2X1_568/Y 0.05fF
C7481 PAND2X1_244/B POR2X1_494/Y 0.03fF
C7482 POR2X1_130/A POR2X1_590/Y 0.00fF
C7483 POR2X1_29/Y POR2X1_38/Y 0.13fF
C7484 PAND2X1_13/a_76_28# POR2X1_186/B 0.02fF
C7485 PAND2X1_181/O POR2X1_55/Y 0.01fF
C7486 POR2X1_796/A POR2X1_294/B 11.92fF
C7487 POR2X1_68/A PAND2X1_393/CTRL 0.03fF
C7488 POR2X1_62/Y POR2X1_5/Y 0.19fF
C7489 POR2X1_305/Y POR2X1_387/Y 0.01fF
C7490 POR2X1_7/B POR2X1_534/Y 0.03fF
C7491 PAND2X1_803/a_76_28# PAND2X1_803/A 0.05fF
C7492 POR2X1_617/a_16_28# POR2X1_408/Y 0.01fF
C7493 POR2X1_187/Y PAND2X1_192/Y 0.17fF
C7494 PAND2X1_551/A PAND2X1_854/A 0.19fF
C7495 POR2X1_327/Y POR2X1_686/B 0.12fF
C7496 POR2X1_468/CTRL POR2X1_444/Y 0.01fF
C7497 POR2X1_380/O POR2X1_380/Y 0.01fF
C7498 PAND2X1_251/a_76_28# PAND2X1_52/B 0.01fF
C7499 PAND2X1_90/Y POR2X1_383/CTRL 0.01fF
C7500 POR2X1_271/A PAND2X1_515/CTRL2 0.19fF
C7501 POR2X1_68/A POR2X1_855/B 0.11fF
C7502 PAND2X1_156/A VDD 3.08fF
C7503 POR2X1_283/A POR2X1_248/CTRL 0.01fF
C7504 POR2X1_579/Y POR2X1_244/Y 0.06fF
C7505 PAND2X1_603/a_16_344# PAND2X1_72/A 0.02fF
C7506 POR2X1_113/Y PAND2X1_153/O 0.17fF
C7507 POR2X1_355/B POR2X1_326/A 0.03fF
C7508 POR2X1_365/Y POR2X1_357/CTRL2 0.00fF
C7509 PAND2X1_140/A PAND2X1_113/O 0.02fF
C7510 POR2X1_327/CTRL2 PAND2X1_48/A 0.00fF
C7511 INPUT_1 POR2X1_416/Y 0.06fF
C7512 POR2X1_619/Y POR2X1_408/Y 0.03fF
C7513 PAND2X1_830/Y POR2X1_131/A 0.00fF
C7514 POR2X1_16/Y POR2X1_42/Y 0.01fF
C7515 POR2X1_709/O PAND2X1_69/A 0.18fF
C7516 POR2X1_13/A PAND2X1_851/O 0.01fF
C7517 POR2X1_516/a_16_28# POR2X1_516/A 0.05fF
C7518 POR2X1_142/Y PAND2X1_149/A 0.01fF
C7519 D_GATE_479 POR2X1_356/Y 0.09fF
C7520 POR2X1_132/CTRL POR2X1_7/B 0.01fF
C7521 POR2X1_753/Y POR2X1_90/CTRL 0.03fF
C7522 PAND2X1_284/Y POR2X1_258/Y 0.01fF
C7523 POR2X1_313/CTRL2 POR2X1_313/Y 0.01fF
C7524 PAND2X1_360/Y POR2X1_42/Y 0.90fF
C7525 INPUT_1 POR2X1_29/Y 0.11fF
C7526 POR2X1_416/B PAND2X1_733/O 0.09fF
C7527 POR2X1_802/B POR2X1_802/A 0.01fF
C7528 POR2X1_362/A POR2X1_501/B 0.15fF
C7529 PAND2X1_232/CTRL POR2X1_68/B -0.01fF
C7530 POR2X1_62/Y POR2X1_522/a_16_28# 0.01fF
C7531 POR2X1_222/Y POR2X1_186/B 0.03fF
C7532 POR2X1_96/Y POR2X1_88/Y 0.03fF
C7533 PAND2X1_139/CTRL POR2X1_13/A 0.01fF
C7534 POR2X1_865/B POR2X1_249/Y 0.05fF
C7535 POR2X1_614/A POR2X1_244/Y 2.23fF
C7536 POR2X1_509/CTRL PAND2X1_41/B 0.00fF
C7537 D_INPUT_2 POR2X1_5/CTRL2 0.01fF
C7538 POR2X1_550/A POR2X1_550/Y 0.02fF
C7539 POR2X1_750/B PAND2X1_72/A 0.29fF
C7540 POR2X1_517/CTRL POR2X1_13/A 0.01fF
C7541 PAND2X1_41/B POR2X1_181/Y 0.03fF
C7542 PAND2X1_21/O D_INPUT_4 0.15fF
C7543 PAND2X1_23/Y POR2X1_447/B 0.12fF
C7544 PAND2X1_736/A PAND2X1_330/CTRL2 0.05fF
C7545 POR2X1_54/CTRL2 D_INPUT_1 0.01fF
C7546 VDD POR2X1_731/Y 0.10fF
C7547 PAND2X1_714/CTRL2 PAND2X1_326/B 0.01fF
C7548 VDD POR2X1_568/O 0.00fF
C7549 PAND2X1_390/m4_208_n4# PAND2X1_853/B 0.15fF
C7550 POR2X1_239/O POR2X1_153/Y 0.06fF
C7551 PAND2X1_639/Y PAND2X1_639/B 0.02fF
C7552 PAND2X1_6/Y POR2X1_737/A 0.03fF
C7553 POR2X1_346/O POR2X1_507/A 0.03fF
C7554 POR2X1_360/CTRL2 POR2X1_244/Y 0.00fF
C7555 POR2X1_538/A POR2X1_703/A 0.07fF
C7556 POR2X1_108/Y PAND2X1_114/B 0.00fF
C7557 POR2X1_447/B PAND2X1_625/O 0.09fF
C7558 POR2X1_532/A POR2X1_186/B 0.10fF
C7559 POR2X1_388/CTRL2 POR2X1_337/Y 0.00fF
C7560 PAND2X1_213/Y PAND2X1_704/O 0.01fF
C7561 PAND2X1_798/B PAND2X1_865/A 0.02fF
C7562 POR2X1_10/O PAND2X1_63/B 0.01fF
C7563 PAND2X1_81/CTRL2 POR2X1_4/Y 0.01fF
C7564 POR2X1_598/CTRL2 POR2X1_260/A 0.01fF
C7565 POR2X1_23/Y PAND2X1_464/B 0.05fF
C7566 PAND2X1_403/B PAND2X1_403/O 0.01fF
C7567 POR2X1_441/CTRL2 POR2X1_669/B 0.03fF
C7568 POR2X1_846/A PAND2X1_58/A 0.05fF
C7569 PAND2X1_850/Y POR2X1_43/B 0.22fF
C7570 POR2X1_596/A POR2X1_294/A 0.03fF
C7571 PAND2X1_341/B POR2X1_73/Y 0.01fF
C7572 PAND2X1_440/O PAND2X1_793/Y 0.02fF
C7573 PAND2X1_715/B POR2X1_310/Y 0.00fF
C7574 POR2X1_283/A PAND2X1_853/B 0.08fF
C7575 POR2X1_520/CTRL2 POR2X1_559/A 0.01fF
C7576 POR2X1_520/O POR2X1_520/B 0.01fF
C7577 POR2X1_441/Y POR2X1_438/Y 0.01fF
C7578 POR2X1_416/B POR2X1_628/CTRL 0.01fF
C7579 POR2X1_722/CTRL PAND2X1_60/B 0.01fF
C7580 POR2X1_537/Y PAND2X1_60/B 0.04fF
C7581 POR2X1_446/B POR2X1_222/O 0.01fF
C7582 POR2X1_628/a_16_28# POR2X1_39/B 0.01fF
C7583 POR2X1_324/a_16_28# POR2X1_568/Y 0.11fF
C7584 POR2X1_303/O POR2X1_228/Y 0.01fF
C7585 POR2X1_343/Y POR2X1_833/a_16_28# 0.11fF
C7586 POR2X1_102/Y PAND2X1_449/CTRL 0.01fF
C7587 PAND2X1_82/a_76_28# POR2X1_84/A 0.01fF
C7588 POR2X1_431/CTRL2 PAND2X1_390/Y 0.01fF
C7589 PAND2X1_341/B PAND2X1_244/B 0.03fF
C7590 PAND2X1_20/A PAND2X1_612/O 0.02fF
C7591 POR2X1_4/Y PAND2X1_528/CTRL2 0.02fF
C7592 POR2X1_186/O POR2X1_186/B 0.06fF
C7593 POR2X1_687/CTRL POR2X1_452/Y 0.01fF
C7594 POR2X1_68/B PAND2X1_517/a_76_28# 0.01fF
C7595 POR2X1_245/CTRL2 POR2X1_39/B 0.02fF
C7596 POR2X1_556/A POR2X1_269/a_16_28# 0.02fF
C7597 PAND2X1_611/CTRL2 POR2X1_734/A 0.05fF
C7598 POR2X1_614/A PAND2X1_681/CTRL2 0.03fF
C7599 PAND2X1_435/CTRL2 POR2X1_677/Y 0.00fF
C7600 POR2X1_66/B POR2X1_66/O 0.01fF
C7601 PAND2X1_233/a_16_344# INPUT_0 0.02fF
C7602 PAND2X1_619/O POR2X1_29/A 0.01fF
C7603 POR2X1_822/Y POR2X1_77/Y 0.03fF
C7604 POR2X1_532/O PAND2X1_60/B 0.01fF
C7605 PAND2X1_72/CTRL2 PAND2X1_72/A 0.00fF
C7606 POR2X1_776/A POR2X1_590/A 0.03fF
C7607 POR2X1_16/A POR2X1_397/CTRL 0.00fF
C7608 POR2X1_652/CTRL PAND2X1_72/A 0.01fF
C7609 POR2X1_366/Y POR2X1_863/A 0.07fF
C7610 POR2X1_863/A POR2X1_294/B 0.07fF
C7611 POR2X1_416/B PAND2X1_324/a_56_28# 0.00fF
C7612 PAND2X1_639/Y POR2X1_260/A 0.08fF
C7613 PAND2X1_787/A POR2X1_77/Y 0.03fF
C7614 POR2X1_470/m4_208_n4# POR2X1_477/m4_208_n4# 0.15fF
C7615 POR2X1_477/B POR2X1_477/CTRL2 0.00fF
C7616 POR2X1_135/Y PAND2X1_717/A 0.06fF
C7617 PAND2X1_177/O PAND2X1_52/B 0.04fF
C7618 POR2X1_714/CTRL2 PAND2X1_72/A 0.01fF
C7619 POR2X1_166/CTRL2 POR2X1_167/Y 0.00fF
C7620 POR2X1_20/B POR2X1_423/Y 0.06fF
C7621 POR2X1_77/CTRL POR2X1_14/Y 0.01fF
C7622 PAND2X1_43/O POR2X1_330/Y 0.03fF
C7623 POR2X1_60/A POR2X1_679/Y 0.10fF
C7624 PAND2X1_424/O PAND2X1_72/A 0.03fF
C7625 POR2X1_257/A POR2X1_495/CTRL2 0.05fF
C7626 PAND2X1_630/B POR2X1_55/Y 0.03fF
C7627 POR2X1_99/O PAND2X1_65/Y 0.11fF
C7628 PAND2X1_803/CTRL2 PAND2X1_797/Y 0.03fF
C7629 POR2X1_73/Y POR2X1_166/Y 0.01fF
C7630 PAND2X1_72/A POR2X1_704/CTRL 0.00fF
C7631 INPUT_3 POR2X1_293/O 0.01fF
C7632 PAND2X1_245/CTRL2 POR2X1_66/A 0.01fF
C7633 POR2X1_856/B POR2X1_590/A 0.06fF
C7634 POR2X1_862/B PAND2X1_39/B 0.03fF
C7635 POR2X1_848/A POR2X1_14/Y 0.07fF
C7636 D_INPUT_0 POR2X1_32/A 0.13fF
C7637 PAND2X1_20/A POR2X1_493/A 0.03fF
C7638 PAND2X1_58/A PAND2X1_591/CTRL 0.01fF
C7639 POR2X1_228/Y PAND2X1_135/O 0.02fF
C7640 POR2X1_801/a_16_28# POR2X1_452/Y 0.03fF
C7641 POR2X1_669/B POR2X1_496/Y 0.07fF
C7642 PAND2X1_299/CTRL2 POR2X1_260/B 0.01fF
C7643 POR2X1_647/B POR2X1_472/Y 0.01fF
C7644 PAND2X1_628/O POR2X1_532/A 0.04fF
C7645 POR2X1_455/a_76_344# POR2X1_341/A 0.02fF
C7646 POR2X1_39/B PAND2X1_123/Y 0.23fF
C7647 POR2X1_37/O D_INPUT_0 0.15fF
C7648 PAND2X1_47/B PAND2X1_25/O 0.02fF
C7649 POR2X1_608/Y POR2X1_606/Y 0.05fF
C7650 POR2X1_476/A POR2X1_476/CTRL 0.00fF
C7651 POR2X1_768/A POR2X1_260/A 0.00fF
C7652 POR2X1_78/B POR2X1_240/CTRL 0.03fF
C7653 PAND2X1_120/O POR2X1_77/Y 0.17fF
C7654 POR2X1_711/Y PAND2X1_692/CTRL2 0.01fF
C7655 POR2X1_67/Y PAND2X1_6/A 0.03fF
C7656 POR2X1_174/B POR2X1_333/A 1.13fF
C7657 POR2X1_54/Y PAND2X1_460/Y 0.01fF
C7658 POR2X1_688/Y VDD 0.01fF
C7659 PAND2X1_443/CTRL VDD 0.00fF
C7660 POR2X1_294/Y POR2X1_852/B 0.02fF
C7661 PAND2X1_717/A POR2X1_816/A 0.03fF
C7662 POR2X1_669/B PAND2X1_733/A 0.03fF
C7663 PAND2X1_496/O POR2X1_499/A 0.02fF
C7664 PAND2X1_444/O POR2X1_236/Y 0.02fF
C7665 POR2X1_394/A PAND2X1_332/Y 0.75fF
C7666 POR2X1_667/CTRL POR2X1_73/Y -0.01fF
C7667 POR2X1_254/Y POR2X1_445/A 0.04fF
C7668 POR2X1_567/B PAND2X1_90/Y 0.05fF
C7669 POR2X1_848/Y POR2X1_859/A 0.03fF
C7670 POR2X1_554/B POR2X1_218/A 0.03fF
C7671 POR2X1_640/Y POR2X1_78/A 0.09fF
C7672 POR2X1_737/A PAND2X1_52/B 0.03fF
C7673 POR2X1_416/B PAND2X1_708/m4_208_n4# 0.07fF
C7674 PAND2X1_817/CTRL POR2X1_750/B 0.00fF
C7675 POR2X1_105/Y POR2X1_296/B 0.20fF
C7676 POR2X1_257/A PAND2X1_552/B 0.03fF
C7677 POR2X1_188/A POR2X1_830/CTRL 0.01fF
C7678 POR2X1_78/B D_INPUT_0 5.69fF
C7679 POR2X1_66/B POR2X1_188/A 0.03fF
C7680 POR2X1_48/A PAND2X1_564/O 0.08fF
C7681 PAND2X1_104/CTRL2 POR2X1_814/B 0.00fF
C7682 PAND2X1_246/O POR2X1_205/A 0.06fF
C7683 POR2X1_803/a_16_28# POR2X1_803/A 0.08fF
C7684 POR2X1_37/Y POR2X1_88/Y 0.02fF
C7685 POR2X1_366/Y POR2X1_274/A 0.03fF
C7686 POR2X1_98/A POR2X1_260/A 0.06fF
C7687 POR2X1_102/Y POR2X1_238/O 0.07fF
C7688 D_INPUT_0 PAND2X1_35/Y 0.03fF
C7689 POR2X1_202/B VDD 0.05fF
C7690 PAND2X1_73/Y PAND2X1_8/Y 0.04fF
C7691 POR2X1_78/A POR2X1_724/CTRL2 0.01fF
C7692 PAND2X1_319/B POR2X1_20/B 0.11fF
C7693 POR2X1_262/Y POR2X1_91/Y 0.02fF
C7694 POR2X1_232/O POR2X1_37/Y 0.03fF
C7695 POR2X1_20/B POR2X1_751/O 0.02fF
C7696 POR2X1_23/Y PAND2X1_705/CTRL2 0.00fF
C7697 POR2X1_64/CTRL2 POR2X1_39/B 0.00fF
C7698 POR2X1_814/B POR2X1_862/B 0.03fF
C7699 POR2X1_590/A POR2X1_722/Y 0.03fF
C7700 POR2X1_49/Y PAND2X1_828/CTRL2 0.03fF
C7701 POR2X1_688/Y PAND2X1_32/B 0.06fF
C7702 POR2X1_78/A POR2X1_121/Y 0.03fF
C7703 POR2X1_41/B POR2X1_225/O 0.04fF
C7704 POR2X1_45/Y PAND2X1_571/A 0.03fF
C7705 D_INPUT_2 POR2X1_48/A 0.07fF
C7706 PAND2X1_263/a_16_344# POR2X1_94/A 0.04fF
C7707 POR2X1_260/B PAND2X1_385/m4_208_n4# 0.15fF
C7708 PAND2X1_719/Y INPUT_0 0.23fF
C7709 PAND2X1_94/A PAND2X1_699/CTRL 0.01fF
C7710 POR2X1_270/CTRL2 POR2X1_446/B 0.01fF
C7711 PAND2X1_575/B INPUT_0 0.06fF
C7712 POR2X1_49/Y POR2X1_177/Y 0.04fF
C7713 PAND2X1_6/Y POR2X1_629/O 0.01fF
C7714 POR2X1_428/Y POR2X1_425/Y 0.03fF
C7715 POR2X1_306/Y POR2X1_236/Y 0.01fF
C7716 POR2X1_852/CTRL POR2X1_852/B 0.06fF
C7717 POR2X1_443/CTRL POR2X1_568/Y 0.31fF
C7718 POR2X1_41/B PAND2X1_219/A 0.03fF
C7719 POR2X1_66/B POR2X1_859/A 0.07fF
C7720 PAND2X1_476/CTRL PAND2X1_473/Y 0.01fF
C7721 POR2X1_556/A POR2X1_218/CTRL 0.01fF
C7722 PAND2X1_732/CTRL POR2X1_763/Y 0.08fF
C7723 POR2X1_77/Y POR2X1_80/a_16_28# 0.00fF
C7724 POR2X1_366/Y POR2X1_269/A 0.04fF
C7725 POR2X1_297/O PAND2X1_347/Y 0.02fF
C7726 POR2X1_260/B POR2X1_140/CTRL2 0.01fF
C7727 POR2X1_43/B PAND2X1_61/CTRL 0.01fF
C7728 PAND2X1_333/O POR2X1_5/Y 0.10fF
C7729 POR2X1_23/CTRL2 POR2X1_42/Y 0.01fF
C7730 POR2X1_298/Y PAND2X1_302/O 0.02fF
C7731 POR2X1_334/B PAND2X1_15/CTRL 0.05fF
C7732 PAND2X1_637/CTRL PAND2X1_69/A 0.01fF
C7733 GATE_479 POR2X1_236/Y 0.01fF
C7734 POR2X1_78/A PAND2X1_145/CTRL2 0.02fF
C7735 D_INPUT_0 POR2X1_184/Y 0.03fF
C7736 POR2X1_407/A POR2X1_858/CTRL 0.00fF
C7737 POR2X1_681/CTRL POR2X1_153/Y 0.06fF
C7738 POR2X1_244/B POR2X1_750/B 0.05fF
C7739 PAND2X1_56/O POR2X1_330/Y 0.04fF
C7740 POR2X1_602/A POR2X1_294/B 0.01fF
C7741 POR2X1_322/CTRL POR2X1_83/B 0.01fF
C7742 POR2X1_389/A PAND2X1_609/O 0.09fF
C7743 POR2X1_444/a_16_28# POR2X1_568/Y 0.12fF
C7744 PAND2X1_56/CTRL POR2X1_593/B 0.01fF
C7745 PAND2X1_116/CTRL VDD 0.00fF
C7746 POR2X1_566/A POR2X1_186/Y 0.07fF
C7747 PAND2X1_651/Y D_INPUT_0 0.10fF
C7748 POR2X1_185/CTRL PAND2X1_73/Y 0.08fF
C7749 POR2X1_78/B PAND2X1_90/Y 0.21fF
C7750 POR2X1_485/O POR2X1_236/Y 0.01fF
C7751 POR2X1_866/B VDD 0.01fF
C7752 POR2X1_476/A POR2X1_68/B 0.03fF
C7753 PAND2X1_182/A POR2X1_312/Y 0.05fF
C7754 POR2X1_504/Y POR2X1_625/Y 0.00fF
C7755 POR2X1_590/A POR2X1_565/O 0.02fF
C7756 PAND2X1_20/A PAND2X1_79/CTRL 0.02fF
C7757 PAND2X1_39/B POR2X1_276/Y 0.02fF
C7758 PAND2X1_57/B POR2X1_398/Y 0.05fF
C7759 POR2X1_66/A PAND2X1_79/Y 0.02fF
C7760 PAND2X1_40/CTRL PAND2X1_11/Y 0.01fF
C7761 POR2X1_569/O POR2X1_355/B 0.10fF
C7762 PAND2X1_659/B PAND2X1_76/Y 0.01fF
C7763 PAND2X1_659/A PAND2X1_659/a_76_28# 0.01fF
C7764 POR2X1_413/A POR2X1_607/O 0.01fF
C7765 POR2X1_65/A PAND2X1_564/a_56_28# 0.00fF
C7766 POR2X1_67/A POR2X1_90/Y 0.07fF
C7767 POR2X1_102/Y POR2X1_56/Y 0.03fF
C7768 PAND2X1_23/Y POR2X1_141/Y 0.03fF
C7769 POR2X1_23/Y POR2X1_283/A 0.20fF
C7770 PAND2X1_9/CTRL2 PAND2X1_69/A 0.01fF
C7771 POR2X1_270/Y POR2X1_222/A 0.00fF
C7772 POR2X1_285/Y POR2X1_649/CTRL2 0.01fF
C7773 POR2X1_20/B PAND2X1_357/CTRL2 0.00fF
C7774 POR2X1_355/B POR2X1_480/A 0.07fF
C7775 PAND2X1_245/O POR2X1_68/B 0.17fF
C7776 POR2X1_49/Y PAND2X1_552/B 0.73fF
C7777 PAND2X1_94/A POR2X1_260/B 0.14fF
C7778 POR2X1_338/O POR2X1_856/B 0.02fF
C7779 PAND2X1_824/a_16_344# POR2X1_856/B 0.06fF
C7780 POR2X1_502/A VDD 4.82fF
C7781 POR2X1_40/Y PAND2X1_566/Y 0.06fF
C7782 POR2X1_284/CTRL2 POR2X1_325/A 0.01fF
C7783 PAND2X1_436/A POR2X1_56/Y 0.07fF
C7784 D_INPUT_3 POR2X1_14/a_76_344# 0.01fF
C7785 PAND2X1_48/Y POR2X1_294/B 0.01fF
C7786 POR2X1_783/A VDD -0.00fF
C7787 PAND2X1_17/O INPUT_7 0.01fF
C7788 POR2X1_5/Y POR2X1_395/O 0.16fF
C7789 POR2X1_254/Y PAND2X1_48/O 0.03fF
C7790 PAND2X1_84/CTRL2 POR2X1_293/Y 0.09fF
C7791 POR2X1_498/Y POR2X1_91/Y 0.03fF
C7792 PAND2X1_124/Y PAND2X1_737/B 0.03fF
C7793 POR2X1_43/B PAND2X1_211/A 0.12fF
C7794 PAND2X1_6/Y POR2X1_302/B 0.03fF
C7795 PAND2X1_769/O POR2X1_763/Y 0.00fF
C7796 POR2X1_164/O POR2X1_40/Y 0.02fF
C7797 PAND2X1_269/CTRL2 POR2X1_236/Y 0.01fF
C7798 POR2X1_83/B INPUT_6 0.03fF
C7799 PAND2X1_817/a_76_28# D_INPUT_1 0.01fF
C7800 PAND2X1_485/CTRL2 POR2X1_260/A 0.01fF
C7801 POR2X1_461/CTRL POR2X1_793/A 0.00fF
C7802 POR2X1_304/O POR2X1_329/A -0.01fF
C7803 POR2X1_528/a_16_28# POR2X1_419/Y 0.03fF
C7804 POR2X1_403/CTRL POR2X1_35/Y 0.00fF
C7805 POR2X1_67/A PAND2X1_154/CTRL 0.05fF
C7806 PAND2X1_803/Y POR2X1_102/Y 0.03fF
C7807 POR2X1_247/CTRL VDD 0.00fF
C7808 PAND2X1_658/a_16_344# POR2X1_816/A 0.01fF
C7809 PAND2X1_96/B POR2X1_202/CTRL2 0.03fF
C7810 POR2X1_147/m4_208_n4# POR2X1_788/m4_208_n4# 0.05fF
C7811 PAND2X1_90/Y PAND2X1_176/a_76_28# 0.01fF
C7812 POR2X1_121/B POR2X1_537/B 0.26fF
C7813 PAND2X1_824/B POR2X1_84/A 0.03fF
C7814 POR2X1_362/Y PAND2X1_106/CTRL -0.02fF
C7815 POR2X1_464/Y VDD 0.00fF
C7816 PAND2X1_632/B POR2X1_482/O 0.01fF
C7817 PAND2X1_651/Y PAND2X1_455/O 0.00fF
C7818 PAND2X1_812/a_16_344# PAND2X1_805/A 0.02fF
C7819 POR2X1_734/A POR2X1_705/O 0.10fF
C7820 POR2X1_660/CTRL POR2X1_725/Y 0.08fF
C7821 VDD PAND2X1_709/CTRL2 0.00fF
C7822 POR2X1_717/CTRL2 POR2X1_777/B 0.04fF
C7823 VDD POR2X1_532/Y 0.01fF
C7824 POR2X1_693/Y POR2X1_692/Y 0.02fF
C7825 PAND2X1_472/A PAND2X1_721/CTRL 0.00fF
C7826 POR2X1_30/O INPUT_7 0.18fF
C7827 POR2X1_23/Y PAND2X1_713/CTRL2 0.01fF
C7828 PAND2X1_20/A POR2X1_510/Y 0.02fF
C7829 INPUT_0 POR2X1_42/Y 0.13fF
C7830 POR2X1_99/A POR2X1_98/B 0.02fF
C7831 PAND2X1_859/A POR2X1_38/B 0.03fF
C7832 POR2X1_277/CTRL POR2X1_46/Y 0.01fF
C7833 POR2X1_61/Y POR2X1_219/CTRL 0.03fF
C7834 PAND2X1_97/O POR2X1_394/A 0.09fF
C7835 PAND2X1_118/CTRL2 INPUT_0 0.03fF
C7836 POR2X1_83/B PAND2X1_154/O 0.15fF
C7837 PAND2X1_793/Y POR2X1_7/B 0.06fF
C7838 POR2X1_669/B PAND2X1_124/CTRL 0.01fF
C7839 POR2X1_8/Y POR2X1_37/Y 0.45fF
C7840 PAND2X1_65/B PAND2X1_518/CTRL2 0.01fF
C7841 PAND2X1_595/a_76_28# POR2X1_249/Y 0.05fF
C7842 PAND2X1_23/Y POR2X1_220/Y 0.10fF
C7843 PAND2X1_795/CTRL2 PAND2X1_175/B 0.01fF
C7844 POR2X1_846/Y POR2X1_39/B 0.22fF
C7845 PAND2X1_137/Y POR2X1_55/Y 0.03fF
C7846 POR2X1_866/B PAND2X1_32/B 0.04fF
C7847 POR2X1_121/A POR2X1_130/A 0.06fF
C7848 POR2X1_43/B POR2X1_821/CTRL 0.01fF
C7849 POR2X1_232/O POR2X1_293/Y 0.01fF
C7850 PAND2X1_227/CTRL POR2X1_236/Y 0.29fF
C7851 POR2X1_302/CTRL2 PAND2X1_32/B 0.01fF
C7852 POR2X1_102/Y PAND2X1_508/CTRL2 0.04fF
C7853 POR2X1_10/O POR2X1_32/A 0.01fF
C7854 POR2X1_194/A POR2X1_194/a_16_28# 0.01fF
C7855 POR2X1_860/O POR2X1_296/B 0.01fF
C7856 PAND2X1_478/O PAND2X1_480/B 0.08fF
C7857 POR2X1_502/A POR2X1_741/Y 0.03fF
C7858 POR2X1_52/A PAND2X1_213/A 0.01fF
C7859 POR2X1_48/A PAND2X1_123/Y 0.03fF
C7860 POR2X1_510/A POR2X1_510/a_16_28# 0.02fF
C7861 POR2X1_52/A PAND2X1_776/O 0.03fF
C7862 POR2X1_68/A POR2X1_192/Y 0.05fF
C7863 POR2X1_83/B POR2X1_59/CTRL 0.01fF
C7864 PAND2X1_546/Y POR2X1_46/Y 0.01fF
C7865 PAND2X1_769/O POR2X1_73/Y 0.02fF
C7866 POR2X1_659/m4_208_n4# POR2X1_736/A 0.05fF
C7867 POR2X1_96/A POR2X1_43/B 2.37fF
C7868 POR2X1_267/O POR2X1_260/A 0.01fF
C7869 POR2X1_65/A POR2X1_387/Y 0.09fF
C7870 POR2X1_315/Y POR2X1_40/Y 0.08fF
C7871 PAND2X1_90/A POR2X1_55/Y 0.03fF
C7872 PAND2X1_372/CTRL2 POR2X1_778/B 0.03fF
C7873 POR2X1_795/B POR2X1_776/B 0.03fF
C7874 PAND2X1_661/Y POR2X1_39/CTRL 0.00fF
C7875 PAND2X1_50/O D_INPUT_6 0.00fF
C7876 POR2X1_673/CTRL POR2X1_260/A 0.01fF
C7877 POR2X1_579/Y PAND2X1_111/CTRL 0.00fF
C7878 POR2X1_477/A POR2X1_740/Y 0.03fF
C7879 POR2X1_102/a_16_28# POR2X1_54/Y 0.10fF
C7880 POR2X1_260/B PAND2X1_136/CTRL2 0.01fF
C7881 POR2X1_43/B PAND2X1_335/O 0.05fF
C7882 PAND2X1_356/B PAND2X1_356/O 0.00fF
C7883 POR2X1_509/a_76_344# POR2X1_509/A 0.01fF
C7884 D_INPUT_0 POR2X1_294/A 0.22fF
C7885 POR2X1_236/Y POR2X1_142/Y 0.03fF
C7886 POR2X1_502/A PAND2X1_32/B 0.21fF
C7887 PAND2X1_740/O POR2X1_283/A 0.08fF
C7888 POR2X1_861/CTRL POR2X1_572/B 0.01fF
C7889 POR2X1_555/B POR2X1_228/CTRL2 0.01fF
C7890 POR2X1_242/a_16_28# POR2X1_566/B 0.04fF
C7891 POR2X1_259/CTRL2 PAND2X1_52/Y 0.01fF
C7892 POR2X1_811/A POR2X1_294/A 0.09fF
C7893 POR2X1_307/Y POR2X1_513/Y 0.40fF
C7894 POR2X1_57/A PAND2X1_520/CTRL 0.02fF
C7895 PAND2X1_371/CTRL2 PAND2X1_69/A 0.01fF
C7896 POR2X1_807/A POR2X1_796/A 0.03fF
C7897 POR2X1_407/A PAND2X1_498/O 0.04fF
C7898 POR2X1_685/CTRL POR2X1_729/Y 0.02fF
C7899 POR2X1_96/A POR2X1_38/B 0.03fF
C7900 POR2X1_814/B POR2X1_276/Y 0.03fF
C7901 PAND2X1_597/a_16_344# POR2X1_796/A 0.02fF
C7902 POR2X1_143/CTRL2 D_INPUT_3 0.12fF
C7903 POR2X1_423/Y PAND2X1_715/B 0.04fF
C7904 POR2X1_227/A POR2X1_568/A 0.03fF
C7905 POR2X1_477/A POR2X1_732/O 0.02fF
C7906 POR2X1_368/CTRL2 POR2X1_283/A 0.03fF
C7907 PAND2X1_55/Y POR2X1_435/CTRL2 0.01fF
C7908 POR2X1_137/CTRL PAND2X1_96/B 0.05fF
C7909 POR2X1_719/O VDD 0.00fF
C7910 PAND2X1_241/O POR2X1_90/Y 0.02fF
C7911 POR2X1_549/a_16_28# POR2X1_383/A 0.02fF
C7912 POR2X1_121/B PAND2X1_48/A 1.24fF
C7913 PAND2X1_55/Y POR2X1_576/Y 0.01fF
C7914 POR2X1_517/Y POR2X1_73/Y 0.05fF
C7915 PAND2X1_831/CTRL2 POR2X1_153/Y 0.00fF
C7916 POR2X1_90/Y PAND2X1_302/CTRL2 0.00fF
C7917 POR2X1_341/A POR2X1_715/CTRL 0.03fF
C7918 POR2X1_88/Y POR2X1_408/Y 0.14fF
C7919 POR2X1_516/CTRL POR2X1_184/Y 0.00fF
C7920 POR2X1_590/A POR2X1_191/Y 0.05fF
C7921 POR2X1_614/A PAND2X1_111/CTRL 0.01fF
C7922 POR2X1_572/B POR2X1_501/B 0.03fF
C7923 POR2X1_68/A PAND2X1_29/O 0.19fF
C7924 PAND2X1_572/CTRL2 PAND2X1_197/Y 0.00fF
C7925 POR2X1_83/A PAND2X1_243/CTRL2 0.00fF
C7926 POR2X1_35/Y POR2X1_219/CTRL 0.01fF
C7927 POR2X1_343/Y PAND2X1_251/CTRL 0.01fF
C7928 PAND2X1_137/a_76_28# POR2X1_132/Y 0.02fF
C7929 POR2X1_537/a_16_28# POR2X1_389/Y 0.01fF
C7930 POR2X1_394/A PAND2X1_562/B 0.08fF
C7931 INPUT_1 POR2X1_29/O 0.02fF
C7932 POR2X1_252/CTRL POR2X1_7/A 0.02fF
C7933 PAND2X1_152/O PAND2X1_60/B 0.06fF
C7934 POR2X1_85/a_16_28# POR2X1_23/Y 0.03fF
C7935 PAND2X1_182/O PAND2X1_357/Y 0.02fF
C7936 POR2X1_57/A POR2X1_312/CTRL2 0.03fF
C7937 POR2X1_5/Y POR2X1_6/O 0.02fF
C7938 PAND2X1_278/CTRL2 POR2X1_294/A 0.06fF
C7939 POR2X1_676/Y POR2X1_687/A 0.01fF
C7940 PAND2X1_216/B PAND2X1_140/Y 0.03fF
C7941 PAND2X1_48/B PAND2X1_60/B 0.24fF
C7942 POR2X1_130/A POR2X1_664/CTRL 0.03fF
C7943 PAND2X1_57/B POR2X1_707/Y 0.01fF
C7944 POR2X1_134/Y PAND2X1_566/Y 0.03fF
C7945 POR2X1_163/O POR2X1_394/A 0.01fF
C7946 POR2X1_38/Y PAND2X1_339/Y 0.15fF
C7947 POR2X1_729/CTRL2 POR2X1_687/Y 0.00fF
C7948 POR2X1_296/B PAND2X1_136/O 0.06fF
C7949 POR2X1_45/Y PAND2X1_702/a_16_344# 0.02fF
C7950 POR2X1_489/CTRL POR2X1_113/B 0.04fF
C7951 POR2X1_614/A PAND2X1_150/CTRL2 0.04fF
C7952 POR2X1_254/Y POR2X1_260/A 0.03fF
C7953 PAND2X1_865/Y PAND2X1_78/O 0.00fF
C7954 POR2X1_57/A PAND2X1_547/CTRL 0.01fF
C7955 PAND2X1_199/A PAND2X1_123/Y 0.00fF
C7956 PAND2X1_318/m4_208_n4# POR2X1_91/Y 0.12fF
C7957 PAND2X1_57/B POR2X1_771/A 0.01fF
C7958 POR2X1_590/A PAND2X1_102/O 0.00fF
C7959 PAND2X1_474/Y POR2X1_394/A 0.03fF
C7960 PAND2X1_190/Y POR2X1_387/Y 0.10fF
C7961 POR2X1_16/A PAND2X1_468/O 0.11fF
C7962 POR2X1_567/A POR2X1_456/CTRL 0.18fF
C7963 POR2X1_43/B POR2X1_7/A 0.21fF
C7964 PAND2X1_115/B POR2X1_310/Y 0.01fF
C7965 PAND2X1_90/Y POR2X1_294/A 0.24fF
C7966 POR2X1_464/Y POR2X1_543/CTRL2 0.00fF
C7967 PAND2X1_23/Y POR2X1_215/A 0.03fF
C7968 PAND2X1_797/Y POR2X1_72/B 0.03fF
C7969 POR2X1_7/B POR2X1_376/CTRL 0.09fF
C7970 PAND2X1_641/Y POR2X1_46/Y 0.00fF
C7971 PAND2X1_57/B PAND2X1_701/O 0.02fF
C7972 POR2X1_13/A POR2X1_394/A 0.24fF
C7973 PAND2X1_94/A PAND2X1_55/Y 1.71fF
C7974 PAND2X1_270/CTRL2 POR2X1_73/Y 0.01fF
C7975 PAND2X1_119/a_16_344# PAND2X1_96/B 0.02fF
C7976 POR2X1_51/B POR2X1_22/A 0.10fF
C7977 POR2X1_614/A POR2X1_7/A 0.03fF
C7978 POR2X1_162/O POR2X1_161/Y 0.03fF
C7979 PAND2X1_84/Y POR2X1_150/CTRL 0.04fF
C7980 PAND2X1_48/B POR2X1_353/A 0.03fF
C7981 POR2X1_719/O PAND2X1_32/B 0.01fF
C7982 POR2X1_114/B POR2X1_101/Y 0.07fF
C7983 POR2X1_407/A POR2X1_796/A 0.06fF
C7984 POR2X1_661/A POR2X1_655/A 0.08fF
C7985 PAND2X1_175/B PAND2X1_858/Y 0.00fF
C7986 PAND2X1_23/Y POR2X1_332/CTRL 0.01fF
C7987 POR2X1_809/A POR2X1_220/Y 0.10fF
C7988 PAND2X1_41/B PAND2X1_166/O 0.06fF
C7989 POR2X1_12/A PAND2X1_635/Y 0.01fF
C7990 VDD POR2X1_171/Y 0.31fF
C7991 POR2X1_38/B POR2X1_7/A 0.06fF
C7992 PAND2X1_585/a_16_344# PAND2X1_56/A 0.01fF
C7993 VDD POR2X1_188/Y 1.01fF
C7994 POR2X1_416/B PAND2X1_557/A 0.03fF
C7995 PAND2X1_550/B POR2X1_90/Y 0.03fF
C7996 POR2X1_68/A POR2X1_546/CTRL2 0.00fF
C7997 POR2X1_252/Y INPUT_0 0.03fF
C7998 POR2X1_664/O POR2X1_712/Y 0.04fF
C7999 POR2X1_522/Y POR2X1_521/Y 0.02fF
C8000 POR2X1_614/A POR2X1_703/A 0.07fF
C8001 POR2X1_55/Y PAND2X1_853/B 0.16fF
C8002 POR2X1_458/B POR2X1_101/Y 0.01fF
C8003 PAND2X1_674/CTRL POR2X1_186/B 0.01fF
C8004 PAND2X1_534/O PAND2X1_60/B 0.01fF
C8005 POR2X1_327/Y POR2X1_861/O 0.01fF
C8006 POR2X1_569/A POR2X1_318/A 0.07fF
C8007 PAND2X1_714/A POR2X1_77/Y 0.07fF
C8008 POR2X1_833/a_16_28# POR2X1_186/B 0.02fF
C8009 PAND2X1_658/B PAND2X1_508/Y 0.34fF
C8010 PAND2X1_127/CTRL POR2X1_532/A 0.01fF
C8011 POR2X1_569/CTRL PAND2X1_52/B 0.03fF
C8012 POR2X1_559/a_16_28# POR2X1_673/Y 0.04fF
C8013 POR2X1_462/B POR2X1_753/O 0.00fF
C8014 PAND2X1_234/CTRL POR2X1_66/A 0.01fF
C8015 POR2X1_489/CTRL POR2X1_768/A 0.05fF
C8016 PAND2X1_850/Y POR2X1_275/CTRL2 0.03fF
C8017 PAND2X1_440/CTRL2 PAND2X1_580/B 0.00fF
C8018 POR2X1_190/a_76_344# POR2X1_456/B 0.02fF
C8019 PAND2X1_661/B POR2X1_394/A 0.03fF
C8020 PAND2X1_643/Y POR2X1_394/A 0.07fF
C8021 POR2X1_192/Y POR2X1_169/A 0.05fF
C8022 POR2X1_795/B POR2X1_192/B 0.21fF
C8023 POR2X1_423/Y POR2X1_589/Y 0.01fF
C8024 POR2X1_96/B POR2X1_96/CTRL2 0.13fF
C8025 POR2X1_741/Y POR2X1_188/Y 0.03fF
C8026 PAND2X1_501/a_16_344# PAND2X1_501/B 0.02fF
C8027 POR2X1_8/Y POR2X1_408/Y 0.03fF
C8028 PAND2X1_224/CTRL POR2X1_590/A 0.01fF
C8029 POR2X1_38/B POR2X1_384/Y 0.01fF
C8030 POR2X1_220/Y POR2X1_711/Y 0.07fF
C8031 INPUT_5 POR2X1_39/B 0.01fF
C8032 PAND2X1_858/O PAND2X1_858/Y 0.00fF
C8033 POR2X1_140/B POR2X1_554/CTRL2 0.01fF
C8034 POR2X1_460/Y POR2X1_260/B 0.04fF
C8035 PAND2X1_30/O POR2X1_750/B 0.02fF
C8036 PAND2X1_348/A PAND2X1_348/CTRL2 0.03fF
C8037 POR2X1_48/A POR2X1_846/Y 0.38fF
C8038 POR2X1_188/Y PAND2X1_32/B 0.03fF
C8039 POR2X1_391/Y PAND2X1_134/O 0.06fF
C8040 PAND2X1_724/B POR2X1_39/B 0.01fF
C8041 POR2X1_220/Y POR2X1_728/A 2.79fF
C8042 POR2X1_862/m4_208_n4# POR2X1_130/A 0.05fF
C8043 POR2X1_574/Y POR2X1_569/A 0.19fF
C8044 POR2X1_850/O POR2X1_737/A 0.01fF
C8045 PAND2X1_39/B PAND2X1_609/CTRL2 0.00fF
C8046 POR2X1_463/CTRL PAND2X1_58/A 0.01fF
C8047 POR2X1_678/O POR2X1_260/B 0.00fF
C8048 POR2X1_394/A PAND2X1_510/B 0.04fF
C8049 PAND2X1_619/O PAND2X1_618/Y -0.00fF
C8050 POR2X1_361/O POR2X1_294/A 0.08fF
C8051 POR2X1_833/A POR2X1_456/B 0.00fF
C8052 POR2X1_394/A POR2X1_321/Y 0.03fF
C8053 POR2X1_101/O POR2X1_334/Y 0.01fF
C8054 POR2X1_54/Y POR2X1_126/O 0.01fF
C8055 POR2X1_278/Y PAND2X1_349/CTRL 0.01fF
C8056 POR2X1_353/A POR2X1_151/a_16_28# 0.03fF
C8057 PAND2X1_93/B PAND2X1_268/CTRL2 0.01fF
C8058 POR2X1_383/A PAND2X1_48/A 3.48fF
C8059 POR2X1_116/A D_INPUT_0 0.03fF
C8060 POR2X1_189/CTRL POR2X1_816/A 0.01fF
C8061 POR2X1_502/Y POR2X1_854/B 0.16fF
C8062 PAND2X1_6/Y POR2X1_716/CTRL2 0.15fF
C8063 POR2X1_616/Y PAND2X1_154/CTRL 0.01fF
C8064 POR2X1_9/Y POR2X1_226/Y 0.50fF
C8065 POR2X1_129/CTRL POR2X1_411/B 0.00fF
C8066 POR2X1_260/B PAND2X1_406/CTRL2 0.01fF
C8067 POR2X1_110/Y PAND2X1_550/B 0.09fF
C8068 POR2X1_62/Y PAND2X1_100/CTRL 0.01fF
C8069 PAND2X1_132/a_56_28# PAND2X1_52/B 0.00fF
C8070 PAND2X1_269/O POR2X1_268/Y 0.00fF
C8071 PAND2X1_39/B POR2X1_807/O 0.15fF
C8072 PAND2X1_604/a_16_344# PAND2X1_72/A 0.01fF
C8073 POR2X1_77/Y POR2X1_816/A 0.03fF
C8074 POR2X1_329/A PAND2X1_390/Y 0.03fF
C8075 POR2X1_99/A PAND2X1_86/CTRL 0.01fF
C8076 POR2X1_343/Y POR2X1_778/B 0.04fF
C8077 POR2X1_557/B POR2X1_768/O 0.18fF
C8078 POR2X1_814/A PAND2X1_7/Y -0.00fF
C8079 POR2X1_68/A POR2X1_716/a_76_344# 0.03fF
C8080 POR2X1_20/B POR2X1_422/Y 0.05fF
C8081 POR2X1_808/B POR2X1_808/O 0.00fF
C8082 POR2X1_77/Y PAND2X1_359/a_56_28# 0.00fF
C8083 POR2X1_316/Y PAND2X1_349/A 0.03fF
C8084 POR2X1_75/m4_208_n4# POR2X1_416/B 0.07fF
C8085 POR2X1_14/Y PAND2X1_796/B 0.02fF
C8086 POR2X1_556/A POR2X1_330/Y 0.05fF
C8087 INPUT_2 POR2X1_8/CTRL 0.01fF
C8088 PAND2X1_217/B POR2X1_150/Y 0.05fF
C8089 PAND2X1_453/A PAND2X1_796/B 0.02fF
C8090 PAND2X1_609/CTRL2 POR2X1_805/Y 0.03fF
C8091 POR2X1_275/Y PAND2X1_390/Y 0.01fF
C8092 POR2X1_119/Y POR2X1_122/CTRL -0.02fF
C8093 POR2X1_614/CTRL2 POR2X1_614/Y 0.04fF
C8094 PAND2X1_71/Y PAND2X1_48/A 0.04fF
C8095 POR2X1_68/A POR2X1_76/B 0.03fF
C8096 POR2X1_856/B POR2X1_66/A 4.82fF
C8097 POR2X1_66/B PAND2X1_416/CTRL 0.00fF
C8098 POR2X1_866/A POR2X1_590/A 0.04fF
C8099 POR2X1_257/A POR2X1_748/A 0.07fF
C8100 POR2X1_60/A PAND2X1_407/a_16_344# 0.02fF
C8101 PAND2X1_72/A POR2X1_318/A 0.07fF
C8102 POR2X1_260/B PAND2X1_11/Y 0.03fF
C8103 POR2X1_49/Y POR2X1_442/CTRL 0.06fF
C8104 POR2X1_260/B POR2X1_606/Y 0.03fF
C8105 POR2X1_49/Y POR2X1_424/Y 0.07fF
C8106 POR2X1_34/CTRL2 POR2X1_34/Y 0.00fF
C8107 PAND2X1_237/O POR2X1_241/B 0.04fF
C8108 POR2X1_66/A PAND2X1_595/a_56_28# 0.00fF
C8109 PAND2X1_173/a_76_28# PAND2X1_72/A 0.02fF
C8110 POR2X1_357/a_16_28# POR2X1_192/B 0.05fF
C8111 POR2X1_9/Y POR2X1_415/Y 0.02fF
C8112 POR2X1_23/Y POR2X1_14/Y 0.08fF
C8113 POR2X1_677/Y POR2X1_56/Y 0.03fF
C8114 PAND2X1_58/A POR2X1_606/a_16_28# 0.02fF
C8115 POR2X1_807/O POR2X1_805/Y 0.04fF
C8116 PAND2X1_476/A PAND2X1_716/B 0.06fF
C8117 PAND2X1_282/CTRL PAND2X1_73/Y 0.06fF
C8118 POR2X1_326/A POR2X1_532/CTRL2 0.00fF
C8119 PAND2X1_93/B POR2X1_201/O 0.16fF
C8120 POR2X1_150/Y VDD 1.07fF
C8121 PAND2X1_23/Y POR2X1_486/CTRL 0.05fF
C8122 PAND2X1_48/B POR2X1_486/O 0.19fF
C8123 POR2X1_87/O POR2X1_260/A 0.01fF
C8124 POR2X1_738/A POR2X1_568/A 0.03fF
C8125 POR2X1_3/A POR2X1_698/Y 0.20fF
C8126 POR2X1_396/Y POR2X1_825/Y 0.17fF
C8127 POR2X1_416/B PAND2X1_196/m4_208_n4# 0.06fF
C8128 PAND2X1_666/a_16_344# PAND2X1_20/A 0.01fF
C8129 POR2X1_37/Y POR2X1_609/CTRL2 0.00fF
C8130 PAND2X1_341/B POR2X1_86/CTRL 0.01fF
C8131 PAND2X1_429/O PAND2X1_11/Y 0.01fF
C8132 POR2X1_102/Y POR2X1_268/a_76_344# 0.00fF
C8133 POR2X1_647/CTRL POR2X1_362/B 0.06fF
C8134 POR2X1_434/CTRL2 POR2X1_480/A 0.03fF
C8135 POR2X1_859/a_76_344# PAND2X1_57/B 0.01fF
C8136 POR2X1_848/A POR2X1_625/CTRL2 0.01fF
C8137 D_INPUT_0 POR2X1_94/A 6.41fF
C8138 POR2X1_49/Y PAND2X1_68/CTRL2 0.03fF
C8139 PAND2X1_633/CTRL PAND2X1_640/B 0.02fF
C8140 PAND2X1_286/B POR2X1_283/Y 0.01fF
C8141 POR2X1_63/Y POR2X1_46/Y 0.01fF
C8142 POR2X1_674/a_16_28# POR2X1_72/B 0.00fF
C8143 POR2X1_554/B POR2X1_740/Y 0.01fF
C8144 PAND2X1_23/Y PAND2X1_45/a_76_28# 0.01fF
C8145 POR2X1_574/Y PAND2X1_72/A 0.03fF
C8146 POR2X1_55/CTRL POR2X1_94/A 0.01fF
C8147 POR2X1_102/Y PAND2X1_719/Y 0.01fF
C8148 POR2X1_692/CTRL POR2X1_692/Y 0.00fF
C8149 PAND2X1_9/Y POR2X1_247/CTRL 0.00fF
C8150 POR2X1_13/A POR2X1_604/a_16_28# 0.00fF
C8151 PAND2X1_10/O PAND2X1_41/B 0.03fF
C8152 POR2X1_48/A PAND2X1_712/CTRL 0.01fF
C8153 POR2X1_695/Y PAND2X1_712/CTRL2 0.04fF
C8154 PAND2X1_41/CTRL2 POR2X1_294/B 0.01fF
C8155 PAND2X1_75/CTRL2 POR2X1_724/A 0.10fF
C8156 POR2X1_366/Y POR2X1_276/B 0.00fF
C8157 POR2X1_698/a_16_28# POR2X1_394/A 0.06fF
C8158 PAND2X1_63/Y PAND2X1_246/CTRL 0.01fF
C8159 PAND2X1_340/B POR2X1_817/A 0.84fF
C8160 PAND2X1_600/CTRL POR2X1_130/A 0.02fF
C8161 POR2X1_241/B POR2X1_186/Y 0.03fF
C8162 PAND2X1_231/O POR2X1_32/A 0.01fF
C8163 PAND2X1_93/B POR2X1_653/a_56_344# 0.00fF
C8164 PAND2X1_796/B POR2X1_55/Y 0.03fF
C8165 POR2X1_409/B POR2X1_236/Y 0.10fF
C8166 POR2X1_812/A POR2X1_750/B 0.03fF
C8167 PAND2X1_557/A POR2X1_487/Y 0.01fF
C8168 PAND2X1_6/Y POR2X1_864/A 0.14fF
C8169 PAND2X1_576/B INPUT_0 0.03fF
C8170 POR2X1_23/Y PAND2X1_735/O 0.03fF
C8171 POR2X1_137/B POR2X1_391/Y 1.08fF
C8172 PAND2X1_39/B POR2X1_803/A 0.02fF
C8173 POR2X1_423/CTRL2 POR2X1_5/Y 0.01fF
C8174 PAND2X1_485/O POR2X1_546/A 0.13fF
C8175 PAND2X1_640/CTRL2 POR2X1_826/Y 0.01fF
C8176 POR2X1_52/A POR2X1_289/Y 0.01fF
C8177 PAND2X1_216/CTRL PAND2X1_267/Y 0.01fF
C8178 POR2X1_663/CTRL2 POR2X1_78/A 0.00fF
C8179 PAND2X1_771/O POR2X1_73/Y 0.06fF
C8180 PAND2X1_340/B POR2X1_42/Y 0.05fF
C8181 POR2X1_257/A PAND2X1_162/O 0.15fF
C8182 POR2X1_590/A POR2X1_207/A 0.02fF
C8183 PAND2X1_836/CTRL POR2X1_411/B 0.01fF
C8184 PAND2X1_585/O PAND2X1_41/B 0.04fF
C8185 PAND2X1_472/B POR2X1_23/Y 0.07fF
C8186 POR2X1_864/CTRL2 POR2X1_774/Y 0.01fF
C8187 POR2X1_621/A PAND2X1_49/CTRL2 0.00fF
C8188 POR2X1_136/O POR2X1_411/B 0.08fF
C8189 POR2X1_49/Y POR2X1_748/A 0.10fF
C8190 PAND2X1_23/Y POR2X1_610/CTRL -0.00fF
C8191 PAND2X1_413/CTRL VDD -0.00fF
C8192 D_INPUT_7 POR2X1_1/a_16_28# 0.05fF
C8193 POR2X1_49/Y PAND2X1_476/CTRL 0.01fF
C8194 POR2X1_567/B PAND2X1_524/O 0.04fF
C8195 POR2X1_297/O PAND2X1_354/A 0.02fF
C8196 POR2X1_832/Y POR2X1_832/B 0.01fF
C8197 D_INPUT_7 POR2X1_260/A 0.06fF
C8198 POR2X1_66/A POR2X1_722/Y 0.01fF
C8199 PAND2X1_267/O PAND2X1_215/B 0.06fF
C8200 PAND2X1_9/Y POR2X1_409/O 0.01fF
C8201 POR2X1_117/a_16_28# POR2X1_667/A 0.02fF
C8202 PAND2X1_557/A PAND2X1_192/Y 0.03fF
C8203 PAND2X1_23/Y POR2X1_841/B 0.03fF
C8204 PAND2X1_84/CTRL2 POR2X1_60/A 0.01fF
C8205 PAND2X1_437/O POR2X1_186/B 0.09fF
C8206 PAND2X1_738/B PAND2X1_731/B 0.16fF
C8207 POR2X1_856/B POR2X1_802/B 0.03fF
C8208 POR2X1_302/Y POR2X1_590/A 0.02fF
C8209 POR2X1_23/Y POR2X1_55/Y 2.72fF
C8210 POR2X1_13/A POR2X1_669/B 0.26fF
C8211 POR2X1_32/A PAND2X1_735/Y 0.10fF
C8212 POR2X1_25/Y POR2X1_698/Y 0.01fF
C8213 POR2X1_23/Y PAND2X1_726/CTRL2 0.10fF
C8214 POR2X1_274/A POR2X1_140/B 0.03fF
C8215 POR2X1_776/A POR2X1_532/A 0.03fF
C8216 POR2X1_471/A POR2X1_540/A 0.03fF
C8217 PAND2X1_58/A PAND2X1_511/CTRL 0.01fF
C8218 POR2X1_68/A POR2X1_301/A 0.02fF
C8219 POR2X1_257/A PAND2X1_785/A 0.01fF
C8220 PAND2X1_808/Y PAND2X1_771/Y 0.64fF
C8221 POR2X1_590/A POR2X1_723/a_16_28# 0.00fF
C8222 POR2X1_590/A PAND2X1_754/CTRL 0.01fF
C8223 POR2X1_362/B POR2X1_405/O 0.02fF
C8224 POR2X1_707/B VDD 0.47fF
C8225 POR2X1_376/B PAND2X1_513/CTRL2 0.15fF
C8226 POR2X1_30/a_16_28# D_INPUT_5 0.03fF
C8227 POR2X1_54/Y POR2X1_15/CTRL 0.01fF
C8228 POR2X1_60/A POR2X1_88/Y 0.03fF
C8229 POR2X1_567/B D_GATE_222 0.10fF
C8230 POR2X1_465/B POR2X1_296/B 0.31fF
C8231 POR2X1_285/Y POR2X1_121/Y 0.03fF
C8232 POR2X1_123/A POR2X1_633/a_16_28# 0.01fF
C8233 POR2X1_188/CTRL PAND2X1_39/B 0.01fF
C8234 POR2X1_695/O POR2X1_425/Y 0.02fF
C8235 PAND2X1_35/A POR2X1_38/Y 0.03fF
C8236 PAND2X1_347/Y PAND2X1_349/B 0.01fF
C8237 POR2X1_568/A POR2X1_731/Y 0.01fF
C8238 PAND2X1_557/A PAND2X1_738/Y 0.44fF
C8239 PAND2X1_40/O PAND2X1_59/B 0.02fF
C8240 POR2X1_32/A PAND2X1_493/Y 0.04fF
C8241 PAND2X1_735/a_76_28# PAND2X1_573/B 0.05fF
C8242 POR2X1_541/B POR2X1_203/a_16_28# 0.01fF
C8243 POR2X1_568/A POR2X1_568/O 0.01fF
C8244 POR2X1_319/A POR2X1_714/CTRL2 0.00fF
C8245 POR2X1_36/B POR2X1_12/A 0.40fF
C8246 PAND2X1_90/A PAND2X1_245/O 0.01fF
C8247 D_INPUT_5 PAND2X1_60/B 0.02fF
C8248 POR2X1_865/O POR2X1_260/B 0.01fF
C8249 PAND2X1_76/Y POR2X1_5/Y 0.03fF
C8250 PAND2X1_20/A POR2X1_578/Y 10.02fF
C8251 PAND2X1_480/B POR2X1_40/Y 0.05fF
C8252 PAND2X1_601/CTRL2 PAND2X1_60/B 0.01fF
C8253 POR2X1_493/A PAND2X1_32/B 0.03fF
C8254 POR2X1_862/B VDD 0.03fF
C8255 POR2X1_264/Y PAND2X1_73/Y 0.05fF
C8256 POR2X1_502/A POR2X1_808/A 0.02fF
C8257 PAND2X1_259/a_16_344# PAND2X1_569/Y 0.02fF
C8258 POR2X1_865/B POR2X1_458/CTRL 0.03fF
C8259 POR2X1_54/Y PAND2X1_63/B 0.03fF
C8260 POR2X1_102/Y POR2X1_42/Y 0.77fF
C8261 PAND2X1_453/O POR2X1_60/A 0.05fF
C8262 POR2X1_853/A POR2X1_78/A 0.03fF
C8263 POR2X1_52/A PAND2X1_512/CTRL 0.01fF
C8264 POR2X1_63/O POR2X1_669/B 0.01fF
C8265 PAND2X1_455/a_16_344# PAND2X1_445/Y 0.02fF
C8266 POR2X1_72/B POR2X1_531/CTRL 0.01fF
C8267 POR2X1_648/Y PAND2X1_48/A 5.13fF
C8268 D_INPUT_3 POR2X1_612/Y 0.35fF
C8269 PAND2X1_39/B POR2X1_598/CTRL 0.04fF
C8270 POR2X1_856/B POR2X1_532/A 0.06fF
C8271 PAND2X1_217/B PAND2X1_364/B 0.36fF
C8272 POR2X1_78/A POR2X1_391/Y 0.14fF
C8273 PAND2X1_801/a_76_28# POR2X1_236/Y 0.00fF
C8274 POR2X1_41/B PAND2X1_842/CTRL 0.02fF
C8275 POR2X1_651/Y POR2X1_711/Y 0.03fF
C8276 POR2X1_264/O POR2X1_294/B 0.03fF
C8277 PAND2X1_793/Y PAND2X1_220/Y 0.03fF
C8278 POR2X1_270/O POR2X1_66/A 0.01fF
C8279 POR2X1_52/A POR2X1_504/Y 0.04fF
C8280 PAND2X1_48/B POR2X1_750/B 0.11fF
C8281 POR2X1_264/Y POR2X1_264/CTRL 0.01fF
C8282 PAND2X1_89/CTRL POR2X1_61/Y 0.02fF
C8283 PAND2X1_222/A POR2X1_385/O 0.00fF
C8284 PAND2X1_341/O POR2X1_40/Y 0.01fF
C8285 PAND2X1_90/A PAND2X1_412/CTRL2 0.01fF
C8286 POR2X1_464/O VDD 0.00fF
C8287 POR2X1_701/Y VDD 0.01fF
C8288 POR2X1_197/CTRL2 POR2X1_244/B 0.01fF
C8289 POR2X1_278/Y PAND2X1_204/O 0.12fF
C8290 PAND2X1_643/Y POR2X1_669/B 0.03fF
C8291 PAND2X1_85/Y PAND2X1_57/B 0.04fF
C8292 POR2X1_60/A POR2X1_289/O 0.02fF
C8293 POR2X1_312/Y POR2X1_55/Y 0.03fF
C8294 PAND2X1_362/B PAND2X1_730/B 0.08fF
C8295 PAND2X1_73/Y POR2X1_541/CTRL2 0.01fF
C8296 POR2X1_590/A POR2X1_501/B 0.05fF
C8297 POR2X1_283/Y PAND2X1_794/B 0.03fF
C8298 GATE_741 PAND2X1_362/B 0.00fF
C8299 PAND2X1_738/Y PAND2X1_544/O 0.04fF
C8300 INPUT_1 PAND2X1_35/A 0.02fF
C8301 POR2X1_392/B POR2X1_392/a_16_28# 0.01fF
C8302 POR2X1_407/Y PAND2X1_11/Y 2.28fF
C8303 POR2X1_43/B PAND2X1_639/CTRL 0.01fF
C8304 POR2X1_668/Y VDD 0.03fF
C8305 POR2X1_655/CTRL POR2X1_711/Y 0.06fF
C8306 POR2X1_327/Y PAND2X1_39/B 0.20fF
C8307 POR2X1_707/B PAND2X1_32/B 0.02fF
C8308 PAND2X1_478/Y POR2X1_43/B 0.01fF
C8309 PAND2X1_74/O PAND2X1_32/B 0.02fF
C8310 INPUT_1 POR2X1_817/CTRL 0.01fF
C8311 POR2X1_834/Y PAND2X1_93/B 0.05fF
C8312 POR2X1_399/O POR2X1_293/Y 0.18fF
C8313 VDD PAND2X1_364/B 3.20fF
C8314 POR2X1_124/O VDD 0.00fF
C8315 INPUT_7 POR2X1_587/O 0.16fF
C8316 POR2X1_416/B PAND2X1_405/O 0.18fF
C8317 PAND2X1_262/CTRL2 PAND2X1_69/A 0.00fF
C8318 POR2X1_614/A POR2X1_549/CTRL2 0.03fF
C8319 POR2X1_466/CTRL VDD -0.00fF
C8320 POR2X1_29/A PAND2X1_133/CTRL2 0.03fF
C8321 POR2X1_748/A PAND2X1_778/Y 0.03fF
C8322 POR2X1_376/B POR2X1_433/Y 0.03fF
C8323 POR2X1_657/Y POR2X1_540/Y 0.05fF
C8324 POR2X1_516/B POR2X1_293/Y 0.03fF
C8325 PAND2X1_63/Y PAND2X1_41/B 0.09fF
C8326 POR2X1_178/O PAND2X1_220/Y 0.04fF
C8327 POR2X1_423/Y POR2X1_73/Y 8.76fF
C8328 POR2X1_39/CTRL2 POR2X1_38/Y 0.00fF
C8329 POR2X1_862/B PAND2X1_32/B 0.03fF
C8330 POR2X1_32/A PAND2X1_569/B 0.02fF
C8331 POR2X1_32/A POR2X1_158/B 0.03fF
C8332 POR2X1_96/A PAND2X1_758/CTRL2 0.03fF
C8333 POR2X1_496/Y PAND2X1_748/CTRL 0.03fF
C8334 POR2X1_523/Y POR2X1_849/a_16_28# 0.02fF
C8335 VDD PAND2X1_101/O 0.00fF
C8336 PAND2X1_6/Y POR2X1_362/B 0.03fF
C8337 POR2X1_78/B D_GATE_222 0.13fF
C8338 PAND2X1_460/O POR2X1_94/A 0.03fF
C8339 PAND2X1_96/B POR2X1_439/Y 0.22fF
C8340 POR2X1_539/CTRL POR2X1_590/A 0.01fF
C8341 POR2X1_651/O PAND2X1_386/Y 0.02fF
C8342 PAND2X1_65/B POR2X1_804/A 0.05fF
C8343 PAND2X1_84/Y PAND2X1_717/a_16_344# 0.01fF
C8344 PAND2X1_42/O POR2X1_38/B 0.27fF
C8345 POR2X1_65/A POR2X1_166/CTRL 0.01fF
C8346 POR2X1_153/a_56_344# POR2X1_48/A 0.00fF
C8347 POR2X1_334/B PAND2X1_80/a_56_28# 0.00fF
C8348 POR2X1_185/CTRL2 PAND2X1_57/B 0.01fF
C8349 POR2X1_684/O POR2X1_7/B 0.01fF
C8350 POR2X1_323/O POR2X1_73/Y 0.01fF
C8351 POR2X1_614/A POR2X1_155/CTRL2 0.00fF
C8352 VDD POR2X1_357/Y 0.02fF
C8353 POR2X1_66/B PAND2X1_82/Y 0.24fF
C8354 POR2X1_731/CTRL2 VDD 0.00fF
C8355 POR2X1_481/A PAND2X1_357/Y 0.03fF
C8356 POR2X1_834/Y POR2X1_78/A 0.05fF
C8357 PAND2X1_20/A PAND2X1_297/CTRL 0.00fF
C8358 POR2X1_849/a_16_28# PAND2X1_69/A 0.02fF
C8359 POR2X1_708/CTRL POR2X1_407/A 0.01fF
C8360 POR2X1_748/A POR2X1_245/a_16_28# 0.02fF
C8361 POR2X1_65/A D_INPUT_3 0.03fF
C8362 POR2X1_543/A PAND2X1_312/CTRL 0.01fF
C8363 PAND2X1_65/B POR2X1_705/a_16_28# 0.00fF
C8364 POR2X1_83/A PAND2X1_734/B 0.05fF
C8365 POR2X1_567/A POR2X1_629/CTRL2 0.01fF
C8366 POR2X1_311/Y PAND2X1_336/O 0.04fF
C8367 PAND2X1_65/B POR2X1_535/A 0.01fF
C8368 POR2X1_126/O POR2X1_4/Y 0.04fF
C8369 PAND2X1_722/O POR2X1_394/A 0.03fF
C8370 POR2X1_614/A PAND2X1_257/CTRL2 0.03fF
C8371 PAND2X1_20/A POR2X1_664/O 0.00fF
C8372 POR2X1_383/A POR2X1_288/A 0.03fF
C8373 INPUT_7 POR2X1_582/A 0.00fF
C8374 POR2X1_389/A PAND2X1_90/Y 0.07fF
C8375 PAND2X1_104/CTRL2 POR2X1_673/Y 0.08fF
C8376 PAND2X1_865/Y POR2X1_437/CTRL 0.01fF
C8377 POR2X1_794/a_16_28# POR2X1_788/Y 0.02fF
C8378 POR2X1_41/B PAND2X1_469/B 0.10fF
C8379 POR2X1_29/A POR2X1_394/A 0.03fF
C8380 POR2X1_163/Y POR2X1_394/A 0.01fF
C8381 PAND2X1_476/A POR2X1_490/Y 0.03fF
C8382 POR2X1_283/A POR2X1_250/A 0.40fF
C8383 PAND2X1_651/Y PAND2X1_735/Y 0.10fF
C8384 POR2X1_101/CTRL POR2X1_814/B 0.01fF
C8385 PAND2X1_824/B PAND2X1_420/CTRL2 0.05fF
C8386 PAND2X1_445/Y POR2X1_90/Y 0.01fF
C8387 POR2X1_55/m4_208_n4# POR2X1_673/Y 0.08fF
C8388 PAND2X1_88/CTRL POR2X1_260/A 0.01fF
C8389 PAND2X1_808/Y POR2X1_42/Y 0.03fF
C8390 POR2X1_260/B PAND2X1_526/CTRL2 0.03fF
C8391 POR2X1_76/Y POR2X1_702/A 0.99fF
C8392 PAND2X1_96/B POR2X1_192/Y 0.05fF
C8393 POR2X1_391/Y PAND2X1_132/CTRL 0.03fF
C8394 POR2X1_188/A POR2X1_858/B 0.00fF
C8395 POR2X1_294/B PAND2X1_144/O 0.07fF
C8396 POR2X1_263/Y POR2X1_7/Y 0.06fF
C8397 POR2X1_864/A PAND2X1_52/B 0.03fF
C8398 POR2X1_781/A PAND2X1_747/a_76_28# 0.04fF
C8399 POR2X1_46/Y POR2X1_498/A 0.39fF
C8400 POR2X1_16/A POR2X1_492/CTRL -0.02fF
C8401 POR2X1_502/A POR2X1_639/Y 0.15fF
C8402 PAND2X1_23/Y POR2X1_114/B 0.07fF
C8403 POR2X1_844/O POR2X1_546/A 0.10fF
C8404 POR2X1_856/CTRL POR2X1_260/A 0.02fF
C8405 PAND2X1_467/Y POR2X1_376/B 0.07fF
C8406 POR2X1_43/a_16_28# PAND2X1_838/B 0.04fF
C8407 PAND2X1_696/O PAND2X1_93/B 0.03fF
C8408 PAND2X1_41/B POR2X1_260/A 0.38fF
C8409 PAND2X1_811/O PAND2X1_811/Y 0.00fF
C8410 POR2X1_750/B POR2X1_210/B 0.01fF
C8411 POR2X1_510/Y VDD 0.56fF
C8412 PAND2X1_793/Y PAND2X1_575/CTRL 0.01fF
C8413 POR2X1_800/A POR2X1_796/CTRL 0.00fF
C8414 POR2X1_740/Y POR2X1_731/CTRL 0.00fF
C8415 PAND2X1_689/CTRL POR2X1_691/A 0.01fF
C8416 POR2X1_505/Y PAND2X1_507/O 0.16fF
C8417 PAND2X1_6/Y POR2X1_691/CTRL 0.01fF
C8418 POR2X1_740/Y POR2X1_702/A 0.49fF
C8419 PAND2X1_90/a_16_344# POR2X1_590/A 0.01fF
C8420 POR2X1_96/CTRL2 POR2X1_236/Y 0.30fF
C8421 PAND2X1_663/CTRL2 VDD 0.00fF
C8422 PAND2X1_624/A POR2X1_38/Y 0.06fF
C8423 POR2X1_373/Y POR2X1_40/Y 0.03fF
C8424 PAND2X1_813/CTRL POR2X1_5/Y 0.15fF
C8425 PAND2X1_96/B POR2X1_574/CTRL2 0.01fF
C8426 POR2X1_821/Y POR2X1_42/Y 0.40fF
C8427 PAND2X1_23/Y POR2X1_458/B 0.12fF
C8428 POR2X1_60/A POR2X1_385/Y 0.43fF
C8429 PAND2X1_350/A POR2X1_7/A 0.08fF
C8430 POR2X1_93/Y POR2X1_77/Y 0.01fF
C8431 POR2X1_780/CTRL2 POR2X1_294/A 0.03fF
C8432 PAND2X1_849/B VDD 0.31fF
C8433 POR2X1_536/CTRL2 POR2X1_13/A 0.11fF
C8434 POR2X1_276/Y VDD 0.10fF
C8435 POR2X1_415/CTRL2 POR2X1_750/Y 0.03fF
C8436 POR2X1_327/Y POR2X1_814/B 0.08fF
C8437 POR2X1_78/B POR2X1_592/A 0.00fF
C8438 PAND2X1_795/a_76_28# POR2X1_394/A 0.06fF
C8439 POR2X1_43/B POR2X1_38/Y 0.27fF
C8440 POR2X1_389/CTRL2 POR2X1_725/Y 0.01fF
C8441 POR2X1_327/Y POR2X1_733/CTRL 0.06fF
C8442 POR2X1_537/Y POR2X1_389/Y 0.03fF
C8443 POR2X1_785/A POR2X1_854/B 0.05fF
C8444 POR2X1_496/Y POR2X1_39/B 0.12fF
C8445 PAND2X1_23/Y POR2X1_222/A 0.03fF
C8446 POR2X1_78/A POR2X1_383/Y 0.04fF
C8447 POR2X1_101/Y POR2X1_784/A 0.07fF
C8448 PAND2X1_594/CTRL POR2X1_711/Y 0.02fF
C8449 POR2X1_407/O POR2X1_513/B 0.02fF
C8450 POR2X1_432/CTRL2 POR2X1_77/Y 0.03fF
C8451 POR2X1_804/A POR2X1_541/CTRL 0.02fF
C8452 PAND2X1_275/CTRL2 POR2X1_569/A 0.02fF
C8453 POR2X1_327/Y POR2X1_325/A 0.06fF
C8454 POR2X1_741/Y POR2X1_510/Y 0.10fF
C8455 PAND2X1_491/a_16_344# PAND2X1_32/B 0.02fF
C8456 PAND2X1_810/O POR2X1_7/B 0.03fF
C8457 POR2X1_283/A PAND2X1_658/B 0.03fF
C8458 POR2X1_68/A POR2X1_215/Y 0.01fF
C8459 PAND2X1_472/A POR2X1_396/Y 0.02fF
C8460 POR2X1_343/Y PAND2X1_73/Y 0.05fF
C8461 POR2X1_38/Y POR2X1_38/B 0.04fF
C8462 POR2X1_322/Y PAND2X1_565/A 0.00fF
C8463 POR2X1_344/A POR2X1_344/Y 0.04fF
C8464 PAND2X1_363/a_16_344# POR2X1_42/Y 0.01fF
C8465 PAND2X1_703/O POR2X1_236/Y 0.02fF
C8466 POR2X1_316/Y POR2X1_417/Y 0.02fF
C8467 PAND2X1_855/CTRL2 PAND2X1_854/A 0.01fF
C8468 PAND2X1_390/Y POR2X1_589/CTRL 0.01fF
C8469 POR2X1_366/Y POR2X1_456/B 0.07fF
C8470 POR2X1_507/CTRL D_GATE_741 0.02fF
C8471 POR2X1_45/Y PAND2X1_196/O 0.07fF
C8472 POR2X1_860/CTRL POR2X1_572/B 0.01fF
C8473 POR2X1_71/a_16_28# PAND2X1_84/Y 0.03fF
C8474 PAND2X1_709/a_76_28# POR2X1_158/B 0.00fF
C8475 PAND2X1_373/a_76_28# POR2X1_732/B 0.10fF
C8476 POR2X1_510/Y PAND2X1_32/B 0.03fF
C8477 POR2X1_252/CTRL POR2X1_153/Y 0.24fF
C8478 INPUT_0 PAND2X1_48/A 8.44fF
C8479 POR2X1_265/Y POR2X1_406/Y 0.16fF
C8480 PAND2X1_733/A POR2X1_39/B 0.03fF
C8481 POR2X1_334/B PAND2X1_184/O 0.02fF
C8482 POR2X1_580/CTRL2 POR2X1_191/Y 0.12fF
C8483 PAND2X1_57/B PAND2X1_18/B 0.03fF
C8484 POR2X1_210/Y POR2X1_162/Y 0.03fF
C8485 PAND2X1_23/Y PAND2X1_481/CTRL 0.01fF
C8486 POR2X1_327/Y POR2X1_327/O 0.01fF
C8487 INPUT_1 POR2X1_43/B 1.04fF
C8488 PAND2X1_266/O POR2X1_262/Y -0.00fF
C8489 VDD POR2X1_749/Y 0.00fF
C8490 POR2X1_837/A POR2X1_202/A 0.01fF
C8491 POR2X1_569/a_56_344# POR2X1_568/B 0.03fF
C8492 POR2X1_390/B D_INPUT_1 0.05fF
C8493 PAND2X1_639/Y PAND2X1_636/CTRL 0.03fF
C8494 POR2X1_315/Y POR2X1_299/O 0.23fF
C8495 POR2X1_614/A INPUT_1 0.07fF
C8496 POR2X1_276/Y PAND2X1_32/B 0.05fF
C8497 PAND2X1_469/B PAND2X1_308/Y 0.84fF
C8498 POR2X1_773/B PAND2X1_69/A 0.10fF
C8499 POR2X1_567/B POR2X1_440/CTRL2 0.30fF
C8500 POR2X1_48/Y PAND2X1_123/Y 0.06fF
C8501 PAND2X1_671/O INPUT_2 0.07fF
C8502 POR2X1_846/A POR2X1_260/B 0.03fF
C8503 POR2X1_326/A POR2X1_832/B 0.06fF
C8504 PAND2X1_31/CTRL2 D_INPUT_7 0.01fF
C8505 PAND2X1_354/Y POR2X1_42/Y 4.15fF
C8506 POR2X1_542/B POR2X1_787/O 0.01fF
C8507 POR2X1_110/O POR2X1_372/Y 0.06fF
C8508 POR2X1_43/B POR2X1_153/Y 4.04fF
C8509 POR2X1_717/CTRL POR2X1_390/B 0.00fF
C8510 PAND2X1_865/Y POR2X1_96/A 0.09fF
C8511 PAND2X1_96/B PAND2X1_184/CTRL 0.01fF
C8512 INPUT_1 POR2X1_38/B 0.37fF
C8513 POR2X1_167/m4_208_n4# POR2X1_90/Y 0.07fF
C8514 PAND2X1_215/B POR2X1_7/Y 0.07fF
C8515 POR2X1_119/Y PAND2X1_549/a_76_28# 0.02fF
C8516 POR2X1_844/B POR2X1_546/a_16_28# 0.01fF
C8517 POR2X1_81/A POR2X1_13/A 4.20fF
C8518 POR2X1_616/Y POR2X1_617/O 0.01fF
C8519 PAND2X1_858/CTRL2 POR2X1_43/B 0.00fF
C8520 INPUT_0 PAND2X1_102/CTRL2 0.00fF
C8521 POR2X1_834/Y POR2X1_513/CTRL2 0.18fF
C8522 PAND2X1_460/O POR2X1_409/Y 0.00fF
C8523 PAND2X1_531/CTRL2 PAND2X1_32/B 0.01fF
C8524 POR2X1_571/a_16_28# POR2X1_844/B 0.01fF
C8525 POR2X1_686/O POR2X1_260/A 0.02fF
C8526 POR2X1_108/CTRL2 PAND2X1_348/A 0.03fF
C8527 PAND2X1_408/CTRL2 PAND2X1_18/B 0.00fF
C8528 POR2X1_739/O POR2X1_444/Y 0.03fF
C8529 POR2X1_532/A POR2X1_244/Y 0.06fF
C8530 PAND2X1_359/Y PAND2X1_357/Y 0.11fF
C8531 POR2X1_283/A PAND2X1_175/CTRL 0.03fF
C8532 PAND2X1_794/B PAND2X1_365/A 0.00fF
C8533 POR2X1_119/Y PAND2X1_478/CTRL 0.01fF
C8534 POR2X1_9/Y POR2X1_754/Y 0.07fF
C8535 POR2X1_228/Y POR2X1_260/A 0.01fF
C8536 POR2X1_38/B POR2X1_153/Y 0.03fF
C8537 PAND2X1_23/Y PAND2X1_122/CTRL2 0.05fF
C8538 PAND2X1_48/B PAND2X1_122/CTRL 0.01fF
C8539 POR2X1_362/B PAND2X1_52/B 10.12fF
C8540 POR2X1_105/Y POR2X1_717/B 0.00fF
C8541 INPUT_0 PAND2X1_840/Y 0.00fF
C8542 POR2X1_38/B POR2X1_384/A 0.04fF
C8543 PAND2X1_48/B PAND2X1_665/CTRL 0.01fF
C8544 POR2X1_187/Y PAND2X1_190/Y 0.01fF
C8545 PAND2X1_763/CTRL2 PAND2X1_52/B 0.03fF
C8546 POR2X1_10/CTRL POR2X1_7/A 0.01fF
C8547 POR2X1_740/Y POR2X1_738/CTRL 0.00fF
C8548 POR2X1_731/a_16_28# POR2X1_731/A 0.03fF
C8549 POR2X1_741/CTRL2 POR2X1_741/Y 0.00fF
C8550 POR2X1_83/B PAND2X1_635/Y 0.02fF
C8551 POR2X1_130/CTRL2 POR2X1_141/A 0.01fF
C8552 POR2X1_68/B PAND2X1_527/CTRL 0.01fF
C8553 PAND2X1_221/Y POR2X1_283/Y 0.12fF
C8554 D_INPUT_6 POR2X1_3/B 0.01fF
C8555 POR2X1_348/CTRL2 POR2X1_334/Y 0.03fF
C8556 PAND2X1_830/CTRL2 PAND2X1_348/A 0.03fF
C8557 POR2X1_407/Y PAND2X1_328/CTRL2 0.01fF
C8558 POR2X1_614/A PAND2X1_680/CTRL 0.01fF
C8559 PAND2X1_862/B POR2X1_80/CTRL 0.01fF
C8560 POR2X1_702/O POR2X1_715/A 0.01fF
C8561 PAND2X1_659/Y PAND2X1_473/CTRL 0.00fF
C8562 PAND2X1_661/Y POR2X1_16/Y 0.06fF
C8563 POR2X1_145/Y POR2X1_146/Y 0.47fF
C8564 PAND2X1_653/Y PAND2X1_737/O 0.01fF
C8565 POR2X1_271/O POR2X1_271/B 0.00fF
C8566 POR2X1_532/A POR2X1_191/Y 0.05fF
C8567 POR2X1_338/O POR2X1_351/B 0.01fF
C8568 PAND2X1_220/CTRL2 POR2X1_77/Y 0.01fF
C8569 POR2X1_313/Y PAND2X1_317/O 0.03fF
C8570 POR2X1_558/B POR2X1_556/A 0.10fF
C8571 PAND2X1_434/O POR2X1_431/Y 0.00fF
C8572 POR2X1_394/A POR2X1_744/CTRL2 0.01fF
C8573 POR2X1_502/A POR2X1_568/A 0.10fF
C8574 POR2X1_263/O POR2X1_37/Y 0.01fF
C8575 POR2X1_316/Y PAND2X1_651/Y 0.15fF
C8576 POR2X1_499/A POR2X1_218/Y 0.07fF
C8577 PAND2X1_58/A POR2X1_646/B 0.00fF
C8578 PAND2X1_675/A POR2X1_77/Y 0.03fF
C8579 POR2X1_445/A POR2X1_454/A 0.09fF
C8580 PAND2X1_450/CTRL2 POR2X1_158/Y 0.00fF
C8581 PAND2X1_469/B POR2X1_77/Y 0.05fF
C8582 PAND2X1_810/B PAND2X1_223/B 0.03fF
C8583 PAND2X1_242/Y POR2X1_516/B 0.05fF
C8584 POR2X1_703/Y POR2X1_724/B 0.01fF
C8585 PAND2X1_127/m4_208_n4# POR2X1_456/B 0.15fF
C8586 POR2X1_66/B PAND2X1_75/O 0.03fF
C8587 POR2X1_13/A POR2X1_234/A 0.05fF
C8588 POR2X1_472/B POR2X1_66/A 0.00fF
C8589 POR2X1_691/CTRL PAND2X1_52/B 0.01fF
C8590 PAND2X1_63/B POR2X1_4/Y 0.06fF
C8591 D_INPUT_1 PAND2X1_529/O 0.02fF
C8592 POR2X1_617/Y POR2X1_750/Y 0.12fF
C8593 POR2X1_394/A POR2X1_394/a_16_28# 0.01fF
C8594 POR2X1_707/B PAND2X1_426/a_76_28# 0.05fF
C8595 POR2X1_813/CTRL POR2X1_669/B 0.01fF
C8596 POR2X1_333/a_56_344# POR2X1_192/B 0.00fF
C8597 POR2X1_333/O POR2X1_191/Y 0.26fF
C8598 POR2X1_24/Y POR2X1_409/B 0.02fF
C8599 POR2X1_196/CTRL2 POR2X1_334/Y 0.05fF
C8600 POR2X1_444/A POR2X1_444/B 0.08fF
C8601 POR2X1_567/B POR2X1_446/O 0.10fF
C8602 POR2X1_169/A POR2X1_704/CTRL2 0.07fF
C8603 POR2X1_48/A PAND2X1_750/a_76_28# 0.01fF
C8604 POR2X1_460/Y POR2X1_375/Y 0.00fF
C8605 POR2X1_772/a_16_28# POR2X1_768/Y 0.03fF
C8606 POR2X1_129/Y PAND2X1_853/B 0.01fF
C8607 POR2X1_49/Y POR2X1_441/a_16_28# 0.02fF
C8608 POR2X1_630/B POR2X1_61/Y 0.01fF
C8609 POR2X1_78/B PAND2X1_607/O 0.01fF
C8610 POR2X1_76/A POR2X1_218/Y 0.07fF
C8611 POR2X1_864/A POR2X1_467/Y 0.03fF
C8612 POR2X1_54/Y POR2X1_32/A 3.35fF
C8613 POR2X1_567/A POR2X1_456/B 0.06fF
C8614 POR2X1_81/A PAND2X1_510/B 0.01fF
C8615 PAND2X1_73/Y POR2X1_624/Y 0.86fF
C8616 POR2X1_866/A POR2X1_66/A 0.01fF
C8617 PAND2X1_323/O POR2X1_456/B 0.03fF
C8618 POR2X1_458/Y POR2X1_370/Y 0.15fF
C8619 POR2X1_485/Y POR2X1_72/B 0.03fF
C8620 POR2X1_848/A POR2X1_37/Y 0.03fF
C8621 POR2X1_195/A POR2X1_66/A 0.02fF
C8622 PAND2X1_535/O POR2X1_533/Y 0.15fF
C8623 PAND2X1_33/O POR2X1_94/A 0.03fF
C8624 POR2X1_9/Y POR2X1_817/A 0.38fF
C8625 PAND2X1_659/Y PAND2X1_853/B 0.03fF
C8626 PAND2X1_630/B POR2X1_293/Y 0.05fF
C8627 POR2X1_298/O POR2X1_32/A 0.04fF
C8628 POR2X1_112/Y PAND2X1_135/O 0.01fF
C8629 POR2X1_13/A POR2X1_667/CTRL2 0.01fF
C8630 POR2X1_553/A POR2X1_632/Y 0.07fF
C8631 POR2X1_681/Y POR2X1_603/Y 0.03fF
C8632 POR2X1_556/A POR2X1_543/A 0.03fF
C8633 PAND2X1_404/Y POR2X1_83/B 0.02fF
C8634 PAND2X1_612/O POR2X1_472/Y 0.05fF
C8635 POR2X1_39/B PAND2X1_124/CTRL 0.01fF
C8636 POR2X1_48/A POR2X1_496/Y 0.10fF
C8637 POR2X1_9/Y POR2X1_42/Y 0.32fF
C8638 D_INPUT_5 POR2X1_750/B 8.21fF
C8639 POR2X1_290/Y POR2X1_399/Y 0.01fF
C8640 POR2X1_610/Y PAND2X1_41/B 0.01fF
C8641 PAND2X1_96/B POR2X1_76/B 0.04fF
C8642 POR2X1_434/A POR2X1_436/B 0.01fF
C8643 POR2X1_102/Y PAND2X1_576/B 0.03fF
C8644 POR2X1_20/B POR2X1_666/A 0.01fF
C8645 POR2X1_814/B POR2X1_240/CTRL2 0.02fF
C8646 POR2X1_605/B POR2X1_260/B 0.01fF
C8647 POR2X1_119/Y POR2X1_7/Y 0.05fF
C8648 POR2X1_329/A PAND2X1_592/Y 0.03fF
C8649 POR2X1_417/Y POR2X1_298/O 0.01fF
C8650 POR2X1_866/A POR2X1_866/a_76_344# 0.03fF
C8651 POR2X1_558/B POR2X1_474/O 0.07fF
C8652 POR2X1_482/a_16_28# POR2X1_669/B 0.09fF
C8653 POR2X1_29/CTRL PAND2X1_9/Y 0.01fF
C8654 POR2X1_624/Y POR2X1_573/CTRL2 0.01fF
C8655 POR2X1_669/B POR2X1_29/A 0.08fF
C8656 POR2X1_827/a_16_28# POR2X1_42/Y 0.08fF
C8657 POR2X1_13/A POR2X1_603/CTRL2 0.01fF
C8658 POR2X1_852/O POR2X1_776/A 0.02fF
C8659 POR2X1_411/B PAND2X1_556/B 0.02fF
C8660 POR2X1_332/B POR2X1_556/A 0.03fF
C8661 POR2X1_461/Y INPUT_0 0.03fF
C8662 POR2X1_102/Y POR2X1_67/A 0.19fF
C8663 POR2X1_78/B POR2X1_648/CTRL 0.10fF
C8664 PAND2X1_147/a_16_344# POR2X1_142/Y 0.02fF
C8665 POR2X1_630/B POR2X1_35/Y 0.01fF
C8666 POR2X1_15/CTRL2 POR2X1_9/Y 0.01fF
C8667 POR2X1_62/Y PAND2X1_358/O 0.02fF
C8668 POR2X1_848/A POR2X1_615/O 0.02fF
C8669 PAND2X1_39/B PAND2X1_760/CTRL2 0.01fF
C8670 PAND2X1_224/CTRL POR2X1_532/A 0.01fF
C8671 POR2X1_106/a_56_344# POR2X1_60/A 0.00fF
C8672 PAND2X1_58/A POR2X1_788/A 0.03fF
C8673 PAND2X1_669/O POR2X1_750/B 0.03fF
C8674 POR2X1_32/A PAND2X1_784/A 0.85fF
C8675 POR2X1_49/Y POR2X1_263/Y 0.13fF
C8676 PAND2X1_115/CTRL POR2X1_150/Y 0.03fF
C8677 POR2X1_805/O PAND2X1_90/Y 0.00fF
C8678 POR2X1_416/B PAND2X1_156/A 0.05fF
C8679 PAND2X1_299/CTRL D_INPUT_0 0.08fF
C8680 POR2X1_323/Y POR2X1_485/Y 0.01fF
C8681 POR2X1_814/A POR2X1_804/A 0.05fF
C8682 POR2X1_655/Y POR2X1_590/A 0.03fF
C8683 POR2X1_119/CTRL2 POR2X1_411/B 0.01fF
C8684 POR2X1_65/CTRL PAND2X1_6/A 0.03fF
C8685 POR2X1_461/B POR2X1_260/B 0.01fF
C8686 POR2X1_582/Y INPUT_4 0.01fF
C8687 POR2X1_23/Y POR2X1_511/Y 0.07fF
C8688 POR2X1_115/CTRL POR2X1_76/A 0.00fF
C8689 POR2X1_77/O POR2X1_13/A 0.01fF
C8690 POR2X1_628/Y POR2X1_7/B 0.03fF
C8691 POR2X1_294/Y PAND2X1_58/CTRL2 0.00fF
C8692 POR2X1_66/A POR2X1_207/A 0.01fF
C8693 POR2X1_150/Y PAND2X1_717/O 0.02fF
C8694 POR2X1_590/A PAND2X1_525/CTRL2 0.01fF
C8695 PAND2X1_299/CTRL2 POR2X1_121/B 0.01fF
C8696 POR2X1_49/CTRL POR2X1_14/Y 0.01fF
C8697 POR2X1_496/Y PAND2X1_513/O 0.06fF
C8698 POR2X1_13/A PAND2X1_436/O 0.01fF
C8699 PAND2X1_318/a_76_28# POR2X1_20/B 0.01fF
C8700 PAND2X1_623/Y POR2X1_415/A 0.03fF
C8701 PAND2X1_57/B PAND2X1_248/CTRL 0.01fF
C8702 PAND2X1_42/O POR2X1_590/A 0.03fF
C8703 POR2X1_665/O PAND2X1_645/B 0.05fF
C8704 POR2X1_78/B POR2X1_644/B 0.03fF
C8705 PAND2X1_55/Y PAND2X1_67/CTRL 0.01fF
C8706 POR2X1_590/A POR2X1_733/CTRL2 0.03fF
C8707 POR2X1_278/Y PAND2X1_771/Y 0.06fF
C8708 POR2X1_335/A PAND2X1_39/B 0.02fF
C8709 POR2X1_98/CTRL VDD 0.00fF
C8710 POR2X1_644/Y POR2X1_513/B 0.01fF
C8711 POR2X1_423/Y PAND2X1_541/CTRL2 0.01fF
C8712 POR2X1_670/Y POR2X1_672/Y 0.00fF
C8713 PAND2X1_16/O POR2X1_630/A 0.03fF
C8714 PAND2X1_622/a_76_28# PAND2X1_381/Y 0.03fF
C8715 PAND2X1_464/B POR2X1_387/Y 0.04fF
C8716 POR2X1_78/B POR2X1_661/Y 0.03fF
C8717 POR2X1_32/A PAND2X1_501/B 0.03fF
C8718 POR2X1_848/A POR2X1_293/Y 0.18fF
C8719 POR2X1_257/A PAND2X1_6/A 0.07fF
C8720 POR2X1_711/Y POR2X1_513/A 0.02fF
C8721 POR2X1_43/O POR2X1_39/B 0.17fF
C8722 PAND2X1_816/O POR2X1_862/A 0.02fF
C8723 POR2X1_590/A POR2X1_206/A 0.03fF
C8724 POR2X1_814/B POR2X1_673/O 0.01fF
C8725 PAND2X1_404/O PAND2X1_403/Y 0.00fF
C8726 POR2X1_201/O PAND2X1_65/Y 0.03fF
C8727 POR2X1_841/B POR2X1_733/A 0.07fF
C8728 POR2X1_821/O POR2X1_669/B 0.01fF
C8729 POR2X1_65/A POR2X1_60/Y 0.05fF
C8730 POR2X1_831/a_16_28# POR2X1_513/Y 0.02fF
C8731 PAND2X1_413/a_76_28# INPUT_0 0.03fF
C8732 POR2X1_613/a_16_28# POR2X1_55/Y 0.10fF
C8733 POR2X1_660/Y POR2X1_722/Y 0.02fF
C8734 PAND2X1_55/Y PAND2X1_591/CTRL 0.01fF
C8735 PAND2X1_6/Y PAND2X1_422/a_56_28# 0.00fF
C8736 POR2X1_293/CTRL2 POR2X1_5/Y 0.03fF
C8737 POR2X1_102/Y PAND2X1_139/Y 0.07fF
C8738 PAND2X1_265/CTRL INPUT_0 0.07fF
C8739 PAND2X1_52/B D_INPUT_4 0.05fF
C8740 PAND2X1_849/CTRL PAND2X1_61/Y 0.01fF
C8741 PAND2X1_221/Y PAND2X1_365/A 0.01fF
C8742 PAND2X1_471/CTRL POR2X1_14/Y 0.01fF
C8743 PAND2X1_473/B POR2X1_40/Y 0.03fF
C8744 POR2X1_60/A POR2X1_516/B 0.02fF
C8745 POR2X1_441/Y PAND2X1_551/a_16_344# 0.01fF
C8746 POR2X1_126/O D_INPUT_1 0.02fF
C8747 POR2X1_640/O POR2X1_633/Y 0.00fF
C8748 POR2X1_376/B PAND2X1_333/CTRL2 0.08fF
C8749 POR2X1_538/A POR2X1_556/A 0.03fF
C8750 POR2X1_39/B PAND2X1_332/Y 0.03fF
C8751 POR2X1_76/O POR2X1_573/A 0.01fF
C8752 POR2X1_566/A PAND2X1_230/O 0.02fF
C8753 POR2X1_416/Y PAND2X1_640/B 0.01fF
C8754 PAND2X1_840/B POR2X1_37/Y 0.01fF
C8755 PAND2X1_104/O INPUT_0 0.02fF
C8756 PAND2X1_465/O VDD 0.00fF
C8757 POR2X1_630/m4_208_n4# POR2X1_222/Y 0.08fF
C8758 POR2X1_96/A PAND2X1_478/B 0.03fF
C8759 POR2X1_376/B POR2X1_376/Y 0.01fF
C8760 POR2X1_511/Y PAND2X1_513/CTRL 0.00fF
C8761 POR2X1_290/Y POR2X1_14/Y 0.02fF
C8762 PAND2X1_607/O POR2X1_294/A 0.03fF
C8763 PAND2X1_241/O POR2X1_102/Y 0.03fF
C8764 POR2X1_866/A POR2X1_532/A 0.05fF
C8765 POR2X1_855/B POR2X1_803/CTRL 0.01fF
C8766 POR2X1_48/A PAND2X1_324/CTRL 0.01fF
C8767 POR2X1_728/B POR2X1_750/B 0.01fF
C8768 POR2X1_192/Y POR2X1_355/A 0.04fF
C8769 POR2X1_556/A POR2X1_362/A 1.08fF
C8770 PAND2X1_795/a_16_344# INPUT_0 0.01fF
C8771 POR2X1_423/Y PAND2X1_785/Y 0.03fF
C8772 POR2X1_655/A PAND2X1_305/CTRL2 -0.00fF
C8773 POR2X1_427/Y VDD 0.18fF
C8774 PAND2X1_487/a_76_28# PAND2X1_96/B 0.02fF
C8775 PAND2X1_472/A POR2X1_609/Y 0.03fF
C8776 POR2X1_670/Y POR2X1_83/B 0.09fF
C8777 POR2X1_236/CTRL POR2X1_236/Y 0.01fF
C8778 PAND2X1_466/A PAND2X1_308/Y 0.02fF
C8779 POR2X1_41/B POR2X1_495/CTRL 0.06fF
C8780 POR2X1_645/O PAND2X1_90/Y 0.09fF
C8781 POR2X1_593/B POR2X1_220/Y 0.06fF
C8782 POR2X1_42/O POR2X1_37/Y 0.03fF
C8783 POR2X1_376/B PAND2X1_556/B 0.02fF
C8784 PAND2X1_32/CTRL2 POR2X1_294/A 0.00fF
C8785 POR2X1_257/A POR2X1_280/Y 0.06fF
C8786 POR2X1_439/a_16_28# POR2X1_544/A 0.03fF
C8787 POR2X1_691/B POR2X1_866/A 0.03fF
C8788 PAND2X1_159/O POR2X1_55/Y 0.17fF
C8789 PAND2X1_404/A PAND2X1_403/Y 0.01fF
C8790 PAND2X1_39/B POR2X1_249/Y 0.03fF
C8791 PAND2X1_139/B PAND2X1_787/Y 0.16fF
C8792 POR2X1_748/A PAND2X1_790/Y 4.16fF
C8793 POR2X1_257/A PAND2X1_112/O 0.18fF
C8794 PAND2X1_474/Y PAND2X1_499/Y 0.00fF
C8795 POR2X1_297/A PAND2X1_347/Y 0.01fF
C8796 PAND2X1_4/CTRL2 D_INPUT_0 0.00fF
C8797 POR2X1_465/B POR2X1_186/Y 0.08fF
C8798 POR2X1_848/A POR2X1_408/Y 0.10fF
C8799 PAND2X1_55/Y POR2X1_202/CTRL2 0.01fF
C8800 POR2X1_49/CTRL POR2X1_55/Y 0.00fF
C8801 POR2X1_378/CTRL POR2X1_55/Y 0.01fF
C8802 POR2X1_49/Y PAND2X1_215/B 0.07fF
C8803 POR2X1_614/A POR2X1_454/B 0.03fF
C8804 PAND2X1_648/a_76_28# PAND2X1_645/Y 0.02fF
C8805 PAND2X1_669/m4_208_n4# D_INPUT_1 0.08fF
C8806 PAND2X1_520/CTRL POR2X1_236/Y 0.01fF
C8807 POR2X1_102/Y PAND2X1_642/B 1.43fF
C8808 PAND2X1_464/Y POR2X1_83/B 0.06fF
C8809 PAND2X1_48/B POR2X1_389/Y 0.02fF
C8810 POR2X1_411/B PAND2X1_789/O 0.01fF
C8811 POR2X1_48/A POR2X1_280/m4_208_n4# 0.08fF
C8812 POR2X1_13/A PAND2X1_499/Y 0.03fF
C8813 POR2X1_83/B PAND2X1_565/A 0.03fF
C8814 PAND2X1_9/O PAND2X1_6/A 0.16fF
C8815 POR2X1_407/A POR2X1_783/CTRL2 0.09fF
C8816 POR2X1_754/A POR2X1_5/Y 0.03fF
C8817 PAND2X1_456/O PAND2X1_465/B 0.01fF
C8818 POR2X1_46/Y POR2X1_692/Y 0.01fF
C8819 POR2X1_364/A PAND2X1_20/A 0.00fF
C8820 POR2X1_94/CTRL POR2X1_94/A 0.01fF
C8821 PAND2X1_848/CTRL POR2X1_38/B 0.01fF
C8822 POR2X1_188/A PAND2X1_816/a_76_28# 0.01fF
C8823 POR2X1_400/A POR2X1_214/CTRL 0.00fF
C8824 POR2X1_792/CTRL2 PAND2X1_60/B 0.01fF
C8825 POR2X1_66/A POR2X1_7/A 0.03fF
C8826 PAND2X1_787/A POR2X1_32/A 0.21fF
C8827 POR2X1_809/A PAND2X1_761/CTRL2 0.01fF
C8828 POR2X1_454/A POR2X1_260/A 0.02fF
C8829 POR2X1_186/Y D_GATE_741 0.08fF
C8830 POR2X1_477/A POR2X1_675/A 0.12fF
C8831 POR2X1_653/B POR2X1_740/Y 0.00fF
C8832 POR2X1_864/CTRL PAND2X1_32/B 0.01fF
C8833 PAND2X1_283/CTRL POR2X1_654/B 0.02fF
C8834 POR2X1_78/B PAND2X1_322/O 0.04fF
C8835 PAND2X1_286/B PAND2X1_568/B 0.19fF
C8836 POR2X1_130/CTRL POR2X1_260/B 0.01fF
C8837 POR2X1_73/CTRL D_INPUT_0 0.01fF
C8838 POR2X1_740/Y POR2X1_830/A 0.06fF
C8839 POR2X1_634/A POR2X1_68/B 0.06fF
C8840 POR2X1_52/A PAND2X1_209/O 0.01fF
C8841 POR2X1_49/Y PAND2X1_6/A 0.23fF
C8842 PAND2X1_64/CTRL POR2X1_260/A 0.01fF
C8843 POR2X1_36/B POR2X1_83/B 0.14fF
C8844 POR2X1_483/A POR2X1_795/O 0.01fF
C8845 PAND2X1_20/A POR2X1_844/O 0.01fF
C8846 POR2X1_251/a_16_28# PAND2X1_190/Y 0.04fF
C8847 POR2X1_52/A PAND2X1_556/B 1.95fF
C8848 PAND2X1_751/CTRL POR2X1_546/A 0.13fF
C8849 POR2X1_121/B POR2X1_307/A 0.01fF
C8850 POR2X1_578/Y VDD 0.49fF
C8851 POR2X1_480/A POR2X1_832/B 0.01fF
C8852 POR2X1_55/Y POR2X1_372/A 0.03fF
C8853 PAND2X1_641/CTRL POR2X1_263/Y 0.01fF
C8854 POR2X1_66/A POR2X1_703/A 0.56fF
C8855 POR2X1_52/A POR2X1_859/A 0.03fF
C8856 PAND2X1_852/CTRL2 VDD -0.00fF
C8857 PAND2X1_512/CTRL2 POR2X1_239/Y 0.01fF
C8858 POR2X1_774/Y PAND2X1_583/CTRL 0.01fF
C8859 POR2X1_489/CTRL2 POR2X1_68/B 0.03fF
C8860 POR2X1_639/Y POR2X1_639/O 0.01fF
C8861 PAND2X1_297/CTRL2 POR2X1_296/B 0.00fF
C8862 POR2X1_54/Y POR2X1_294/A 0.05fF
C8863 PAND2X1_6/Y POR2X1_555/A 0.03fF
C8864 PAND2X1_742/B PAND2X1_740/Y 0.14fF
C8865 PAND2X1_556/B POR2X1_152/A 0.03fF
C8866 POR2X1_335/A POR2X1_325/A 0.03fF
C8867 POR2X1_417/Y PAND2X1_787/A 0.19fF
C8868 POR2X1_119/Y POR2X1_257/A 0.20fF
C8869 PAND2X1_94/A POR2X1_55/O 0.16fF
C8870 POR2X1_722/A PAND2X1_93/B 0.59fF
C8871 POR2X1_96/A POR2X1_494/Y 1.38fF
C8872 POR2X1_278/Y POR2X1_42/Y 0.03fF
C8873 PAND2X1_57/B POR2X1_294/B 0.47fF
C8874 PAND2X1_56/Y POR2X1_284/B 0.03fF
C8875 POR2X1_366/Y PAND2X1_57/B 0.03fF
C8876 PAND2X1_61/Y PAND2X1_341/A 0.09fF
C8877 POR2X1_330/Y PAND2X1_60/B 0.06fF
C8878 PAND2X1_90/A PAND2X1_92/CTRL2 0.03fF
C8879 PAND2X1_216/O PAND2X1_364/B 0.05fF
C8880 POR2X1_40/Y POR2X1_239/Y 0.01fF
C8881 POR2X1_102/Y PAND2X1_550/B 0.03fF
C8882 POR2X1_23/Y POR2X1_129/Y 0.03fF
C8883 POR2X1_455/a_16_28# POR2X1_455/A 0.02fF
C8884 POR2X1_43/B POR2X1_421/O 0.01fF
C8885 POR2X1_390/B POR2X1_78/A 0.00fF
C8886 PAND2X1_347/Y PAND2X1_566/Y 0.00fF
C8887 POR2X1_863/CTRL POR2X1_855/Y 0.01fF
C8888 PAND2X1_65/B POR2X1_570/B 0.02fF
C8889 POR2X1_508/O POR2X1_192/Y 0.04fF
C8890 INPUT_1 POR2X1_590/A 8.01fF
C8891 PAND2X1_554/a_56_28# PAND2X1_348/Y 0.00fF
C8892 PAND2X1_394/O POR2X1_215/A 0.16fF
C8893 POR2X1_262/O PAND2X1_215/B 0.18fF
C8894 POR2X1_829/A POR2X1_42/Y 0.04fF
C8895 PAND2X1_823/CTRL POR2X1_836/A 0.01fF
C8896 POR2X1_69/a_16_28# POR2X1_7/A 0.02fF
C8897 POR2X1_16/A PAND2X1_721/B 0.03fF
C8898 PAND2X1_231/CTRL2 POR2X1_229/Y 0.00fF
C8899 PAND2X1_23/Y POR2X1_784/A 0.14fF
C8900 POR2X1_826/CTRL2 PAND2X1_338/B 0.08fF
C8901 PAND2X1_673/CTRL2 D_INPUT_3 0.14fF
C8902 POR2X1_383/A PAND2X1_299/CTRL2 0.08fF
C8903 POR2X1_351/B POR2X1_66/A 0.01fF
C8904 POR2X1_517/a_16_28# POR2X1_73/Y 0.04fF
C8905 POR2X1_474/O POR2X1_362/A 0.02fF
C8906 POR2X1_66/B PAND2X1_232/O 0.02fF
C8907 POR2X1_567/B POR2X1_564/CTRL 0.01fF
C8908 POR2X1_807/A PAND2X1_306/a_16_344# 0.03fF
C8909 PAND2X1_20/A POR2X1_398/m4_208_n4# 0.19fF
C8910 POR2X1_52/A POR2X1_599/A 0.08fF
C8911 PAND2X1_659/Y POR2X1_23/Y 0.03fF
C8912 PAND2X1_840/B POR2X1_293/Y 0.05fF
C8913 POR2X1_614/A PAND2X1_56/O 0.06fF
C8914 POR2X1_22/A POR2X1_7/B 0.10fF
C8915 POR2X1_596/A POR2X1_770/A 0.54fF
C8916 PAND2X1_569/B PAND2X1_731/B 0.03fF
C8917 POR2X1_850/O POR2X1_362/B 0.18fF
C8918 POR2X1_78/A POR2X1_209/CTRL2 0.03fF
C8919 POR2X1_23/Y PAND2X1_708/a_76_28# 0.02fF
C8920 PAND2X1_52/a_76_28# PAND2X1_72/A 0.01fF
C8921 POR2X1_625/a_16_28# POR2X1_93/A 0.02fF
C8922 POR2X1_49/Y POR2X1_419/CTRL2 0.05fF
C8923 PAND2X1_23/Y POR2X1_732/B 0.05fF
C8924 PAND2X1_73/Y POR2X1_186/B 0.03fF
C8925 PAND2X1_41/B PAND2X1_670/a_76_28# 0.01fF
C8926 POR2X1_130/A POR2X1_68/B 0.06fF
C8927 PAND2X1_244/CTRL2 POR2X1_153/Y 0.05fF
C8928 PAND2X1_480/B POR2X1_310/O 0.02fF
C8929 POR2X1_445/CTRL2 POR2X1_702/A 0.00fF
C8930 POR2X1_294/B POR2X1_193/O 0.04fF
C8931 POR2X1_278/Y PAND2X1_347/CTRL 0.01fF
C8932 PAND2X1_658/B POR2X1_55/Y 0.01fF
C8933 PAND2X1_250/O POR2X1_249/Y -0.00fF
C8934 PAND2X1_137/CTRL2 POR2X1_134/Y 0.01fF
C8935 POR2X1_327/Y POR2X1_149/A 0.00fF
C8936 POR2X1_96/Y POR2X1_23/Y 0.03fF
C8937 POR2X1_548/CTRL PAND2X1_63/B 0.01fF
C8938 POR2X1_840/CTRL2 POR2X1_307/Y 0.01fF
C8939 POR2X1_176/CTRL2 POR2X1_83/B 0.03fF
C8940 POR2X1_32/A POR2X1_701/CTRL2 0.03fF
C8941 POR2X1_669/A POR2X1_669/a_16_28# 0.03fF
C8942 POR2X1_146/Y POR2X1_669/B 0.01fF
C8943 POR2X1_61/Y POR2X1_259/CTRL 0.02fF
C8944 PAND2X1_679/CTRL POR2X1_687/A 0.01fF
C8945 POR2X1_8/Y POR2X1_750/A 0.03fF
C8946 PAND2X1_69/A POR2X1_208/CTRL2 0.04fF
C8947 POR2X1_114/B POR2X1_733/A 0.06fF
C8948 POR2X1_814/B POR2X1_249/Y 0.03fF
C8949 POR2X1_72/Y POR2X1_816/A 0.01fF
C8950 POR2X1_220/B POR2X1_191/Y 0.05fF
C8951 PAND2X1_821/CTRL POR2X1_510/A 0.00fF
C8952 POR2X1_578/Y PAND2X1_32/B 0.03fF
C8953 POR2X1_750/A POR2X1_749/CTRL2 0.03fF
C8954 POR2X1_239/O POR2X1_7/B 0.17fF
C8955 PAND2X1_499/Y PAND2X1_510/B 0.03fF
C8956 POR2X1_383/A POR2X1_284/B 0.02fF
C8957 PAND2X1_465/B POR2X1_73/Y 0.03fF
C8958 PAND2X1_580/B PAND2X1_854/A 0.02fF
C8959 POR2X1_499/A POR2X1_138/A 0.03fF
C8960 PAND2X1_23/Y POR2X1_249/O 0.01fF
C8961 POR2X1_41/B PAND2X1_389/Y 0.03fF
C8962 POR2X1_817/Y PAND2X1_6/A 0.94fF
C8963 POR2X1_32/A POR2X1_4/Y 9.50fF
C8964 PAND2X1_228/CTRL2 PAND2X1_341/A 0.01fF
C8965 POR2X1_537/a_76_344# POR2X1_188/A 0.00fF
C8966 POR2X1_43/B PAND2X1_449/Y 0.01fF
C8967 POR2X1_57/A PAND2X1_592/Y 0.87fF
C8968 POR2X1_265/Y POR2X1_60/A 0.03fF
C8969 POR2X1_750/Y PAND2X1_526/m4_208_n4# 0.02fF
C8970 POR2X1_83/B POR2X1_701/O 0.18fF
C8971 PAND2X1_41/B POR2X1_559/A 0.10fF
C8972 POR2X1_750/B POR2X1_553/CTRL 0.33fF
C8973 POR2X1_468/O POR2X1_478/B 0.00fF
C8974 POR2X1_16/A PAND2X1_204/O -0.01fF
C8975 POR2X1_761/Y POR2X1_42/Y 0.03fF
C8976 PAND2X1_652/A PAND2X1_186/CTRL2 0.31fF
C8977 POR2X1_16/A POR2X1_238/O 0.02fF
C8978 POR2X1_514/Y POR2X1_139/A 0.00fF
C8979 PAND2X1_715/CTRL2 POR2X1_310/Y 0.01fF
C8980 PAND2X1_48/B POR2X1_318/A 0.07fF
C8981 POR2X1_57/A PAND2X1_839/O 0.01fF
C8982 PAND2X1_798/B POR2X1_73/Y 1.08fF
C8983 POR2X1_853/CTRL POR2X1_854/B 0.15fF
C8984 PAND2X1_799/a_16_344# PAND2X1_364/B 0.02fF
C8985 POR2X1_774/B VDD 0.06fF
C8986 POR2X1_130/A POR2X1_561/O 0.01fF
C8987 POR2X1_311/Y PAND2X1_865/Y 0.07fF
C8988 POR2X1_51/A POR2X1_158/B 0.50fF
C8989 POR2X1_68/A POR2X1_540/A 0.03fF
C8990 POR2X1_376/B PAND2X1_358/A 0.02fF
C8991 PAND2X1_858/a_16_344# PAND2X1_390/Y 0.01fF
C8992 POR2X1_590/O POR2X1_513/B 0.02fF
C8993 POR2X1_43/B POR2X1_591/Y 0.03fF
C8994 PAND2X1_48/B POR2X1_713/B 0.04fF
C8995 PAND2X1_126/CTRL PAND2X1_90/A 0.01fF
C8996 POR2X1_68/B POR2X1_844/B 0.03fF
C8997 POR2X1_722/Y POR2X1_308/B 0.01fF
C8998 PAND2X1_270/CTRL POR2X1_184/Y 0.00fF
C8999 POR2X1_725/Y POR2X1_777/CTRL 0.08fF
C9000 PAND2X1_318/O POR2X1_315/Y 0.02fF
C9001 POR2X1_57/Y PAND2X1_656/A 0.01fF
C9002 POR2X1_618/a_76_344# POR2X1_7/A 0.01fF
C9003 POR2X1_49/Y POR2X1_119/Y 0.59fF
C9004 POR2X1_218/A POR2X1_361/O 0.00fF
C9005 VDD POR2X1_317/B 0.01fF
C9006 PAND2X1_644/Y POR2X1_759/CTRL 0.00fF
C9007 POR2X1_224/CTRL2 POR2X1_394/A 0.05fF
C9008 POR2X1_43/B PAND2X1_470/A 0.01fF
C9009 PAND2X1_170/CTRL2 VDD -0.00fF
C9010 PAND2X1_631/A POR2X1_423/Y 0.03fF
C9011 POR2X1_502/A POR2X1_444/Y 0.01fF
C9012 POR2X1_327/Y VDD 2.39fF
C9013 POR2X1_614/A PAND2X1_312/CTRL 0.01fF
C9014 POR2X1_713/A PAND2X1_48/A 0.00fF
C9015 POR2X1_360/A POR2X1_260/A 0.10fF
C9016 POR2X1_383/A PAND2X1_519/CTRL 0.01fF
C9017 POR2X1_717/CTRL2 POR2X1_865/B 0.01fF
C9018 PAND2X1_18/O PAND2X1_18/B 0.01fF
C9019 PAND2X1_20/A POR2X1_554/a_76_344# 0.00fF
C9020 PAND2X1_211/A PAND2X1_352/Y 0.37fF
C9021 POR2X1_539/A POR2X1_68/A 0.03fF
C9022 POR2X1_619/A POR2X1_382/Y 0.03fF
C9023 PAND2X1_772/O POR2X1_77/Y 0.05fF
C9024 PAND2X1_511/CTRL2 PAND2X1_48/A 0.11fF
C9025 POR2X1_833/O POR2X1_260/A 0.01fF
C9026 PAND2X1_550/B POR2X1_531/Y 0.00fF
C9027 D_INPUT_1 PAND2X1_63/B 0.03fF
C9028 POR2X1_174/B PAND2X1_52/B 0.12fF
C9029 PAND2X1_566/Y PAND2X1_346/Y 0.33fF
C9030 POR2X1_293/Y PAND2X1_853/B 0.03fF
C9031 POR2X1_78/B POR2X1_4/Y 0.03fF
C9032 POR2X1_57/A PAND2X1_839/B 0.03fF
C9033 POR2X1_532/A POR2X1_7/A 0.06fF
C9034 PAND2X1_697/CTRL2 POR2X1_260/A 0.00fF
C9035 PAND2X1_48/B POR2X1_574/Y 0.03fF
C9036 POR2X1_565/B POR2X1_6/a_76_344# 0.02fF
C9037 PAND2X1_800/a_76_28# POR2X1_96/A 0.01fF
C9038 POR2X1_495/CTRL POR2X1_77/Y 0.01fF
C9039 PAND2X1_93/B PAND2X1_628/CTRL 0.01fF
C9040 POR2X1_68/A PAND2X1_6/O 0.01fF
C9041 POR2X1_8/Y PAND2X1_35/a_16_344# 0.02fF
C9042 POR2X1_855/B POR2X1_783/Y 0.01fF
C9043 PAND2X1_562/B POR2X1_39/B 0.11fF
C9044 POR2X1_96/A PAND2X1_341/B 0.49fF
C9045 POR2X1_180/B POR2X1_540/A 0.00fF
C9046 POR2X1_383/A POR2X1_307/A 0.03fF
C9047 POR2X1_774/B PAND2X1_32/B 0.01fF
C9048 POR2X1_730/Y PAND2X1_69/A 0.03fF
C9049 PAND2X1_35/O POR2X1_394/A 0.02fF
C9050 PAND2X1_90/A PAND2X1_527/CTRL 0.03fF
C9051 POR2X1_327/Y POR2X1_741/Y 0.03fF
C9052 POR2X1_283/A POR2X1_387/Y 0.15fF
C9053 POR2X1_49/Y PAND2X1_847/CTRL 0.01fF
C9054 POR2X1_554/Y POR2X1_735/O 0.03fF
C9055 POR2X1_8/Y PAND2X1_227/CTRL 0.00fF
C9056 PAND2X1_185/a_16_344# POR2X1_77/Y 0.02fF
C9057 PAND2X1_149/CTRL2 PAND2X1_797/Y 0.01fF
C9058 POR2X1_334/Y D_GATE_222 0.07fF
C9059 POR2X1_265/Y POR2X1_406/a_56_344# 0.00fF
C9060 POR2X1_43/Y PAND2X1_195/O 0.05fF
C9061 POR2X1_57/A PAND2X1_343/CTRL2 0.03fF
C9062 POR2X1_25/Y POR2X1_47/O 0.01fF
C9063 PAND2X1_227/CTRL2 POR2X1_394/A 0.05fF
C9064 POR2X1_10/CTRL POR2X1_38/Y 0.04fF
C9065 POR2X1_322/Y POR2X1_164/Y 0.00fF
C9066 D_INPUT_6 PAND2X1_1/a_76_28# 0.02fF
C9067 POR2X1_358/O POR2X1_191/Y 0.28fF
C9068 POR2X1_43/B PAND2X1_566/a_76_28# 0.02fF
C9069 POR2X1_38/Y POR2X1_39/Y 0.01fF
C9070 POR2X1_136/a_16_28# PAND2X1_348/A 0.07fF
C9071 PAND2X1_715/CTRL POR2X1_39/B 0.11fF
C9072 PAND2X1_219/O POR2X1_7/Y 0.02fF
C9073 POR2X1_16/A PAND2X1_803/Y 0.01fF
C9074 POR2X1_203/CTRL PAND2X1_72/Y 0.01fF
C9075 POR2X1_860/CTRL2 POR2X1_383/A 0.10fF
C9076 POR2X1_327/Y PAND2X1_32/B 2.33fF
C9077 PAND2X1_476/A POR2X1_406/a_76_344# 0.00fF
C9078 POR2X1_502/A PAND2X1_109/CTRL -0.00fF
C9079 POR2X1_394/A PAND2X1_509/CTRL 0.05fF
C9080 PAND2X1_94/A POR2X1_383/A 1.54fF
C9081 POR2X1_35/Y POR2X1_502/Y 0.05fF
C9082 POR2X1_13/A POR2X1_39/B 0.28fF
C9083 POR2X1_9/Y POR2X1_67/A 0.18fF
C9084 POR2X1_96/A POR2X1_533/Y 0.04fF
C9085 POR2X1_596/A POR2X1_774/A 0.03fF
C9086 PAND2X1_173/CTRL2 POR2X1_186/B 0.03fF
C9087 POR2X1_569/A POR2X1_576/O 0.01fF
C9088 POR2X1_502/A PAND2X1_56/A 0.01fF
C9089 PAND2X1_63/Y POR2X1_571/Y 0.05fF
C9090 PAND2X1_503/a_16_344# POR2X1_854/B 0.06fF
C9091 POR2X1_54/Y POR2X1_286/B 0.01fF
C9092 POR2X1_544/A PAND2X1_52/B 0.01fF
C9093 PAND2X1_653/CTRL2 PAND2X1_652/A 0.03fF
C9094 POR2X1_527/a_76_344# PAND2X1_550/B 0.00fF
C9095 POR2X1_840/B POR2X1_188/Y 0.04fF
C9096 POR2X1_16/A PAND2X1_727/CTRL 0.01fF
C9097 PAND2X1_95/B D_INPUT_4 0.28fF
C9098 POR2X1_124/B PAND2X1_122/CTRL2 0.00fF
C9099 POR2X1_38/B POR2X1_560/CTRL2 0.01fF
C9100 PAND2X1_641/Y POR2X1_83/CTRL 0.02fF
C9101 POR2X1_529/O POR2X1_39/B 0.30fF
C9102 POR2X1_542/B POR2X1_374/CTRL2 0.03fF
C9103 PAND2X1_639/Y POR2X1_584/a_16_28# 0.02fF
C9104 POR2X1_196/O POR2X1_814/A 0.07fF
C9105 PAND2X1_271/CTRL POR2X1_76/A 0.04fF
C9106 POR2X1_416/B PAND2X1_709/CTRL2 0.01fF
C9107 PAND2X1_862/Y PAND2X1_175/B 0.01fF
C9108 POR2X1_566/B POR2X1_566/CTRL 0.02fF
C9109 POR2X1_567/A POR2X1_540/O 0.02fF
C9110 PAND2X1_257/O POR2X1_750/B 0.15fF
C9111 PAND2X1_803/Y PAND2X1_336/Y 0.02fF
C9112 POR2X1_532/A POR2X1_342/a_16_28# 0.01fF
C9113 PAND2X1_63/B POR2X1_620/B 0.03fF
C9114 POR2X1_796/A PAND2X1_48/A 0.07fF
C9115 PAND2X1_341/B POR2X1_7/A 0.03fF
C9116 PAND2X1_94/A PAND2X1_71/Y 2.25fF
C9117 POR2X1_540/A POR2X1_181/O 0.02fF
C9118 PAND2X1_32/CTRL2 POR2X1_94/A 0.03fF
C9119 POR2X1_539/O POR2X1_326/A 0.01fF
C9120 PAND2X1_165/O POR2X1_854/B 0.04fF
C9121 PAND2X1_52/B PAND2X1_145/O 0.09fF
C9122 PAND2X1_476/A POR2X1_229/Y 0.00fF
C9123 PAND2X1_661/B POR2X1_39/B 0.03fF
C9124 PAND2X1_510/O PAND2X1_508/Y 0.01fF
C9125 POR2X1_34/B PAND2X1_39/B 0.02fF
C9126 POR2X1_824/CTRL2 POR2X1_16/A 0.10fF
C9127 POR2X1_309/a_76_344# POR2X1_150/Y 0.01fF
C9128 PAND2X1_60/O POR2X1_66/A 0.01fF
C9129 POR2X1_773/A POR2X1_773/a_16_28# 0.03fF
C9130 POR2X1_188/Y POR2X1_737/O 0.02fF
C9131 PAND2X1_93/B POR2X1_632/O 0.18fF
C9132 POR2X1_502/A POR2X1_661/A 0.07fF
C9133 POR2X1_250/Y PAND2X1_740/CTRL 0.15fF
C9134 POR2X1_78/B POR2X1_458/Y 0.07fF
C9135 PAND2X1_52/B POR2X1_705/O 0.07fF
C9136 POR2X1_554/B POR2X1_141/Y 1.92fF
C9137 POR2X1_394/A PAND2X1_345/Y 0.03fF
C9138 POR2X1_99/B POR2X1_260/A 0.03fF
C9139 POR2X1_9/Y POR2X1_415/O 0.03fF
C9140 PAND2X1_469/O POR2X1_32/A 0.05fF
C9141 POR2X1_748/A POR2X1_20/B 6.92fF
C9142 POR2X1_257/A POR2X1_279/a_16_28# 0.06fF
C9143 PAND2X1_431/O POR2X1_466/A 0.36fF
C9144 POR2X1_23/Y POR2X1_37/Y 0.81fF
C9145 PAND2X1_406/CTRL2 POR2X1_121/B 0.00fF
C9146 PAND2X1_108/O POR2X1_814/A 0.19fF
C9147 PAND2X1_163/CTRL2 PAND2X1_52/B 0.01fF
C9148 PAND2X1_649/A POR2X1_394/a_16_28# 0.02fF
C9149 POR2X1_544/Y POR2X1_551/A 0.01fF
C9150 POR2X1_376/B POR2X1_441/Y 1.31fF
C9151 POR2X1_161/CTRL POR2X1_162/Y 0.01fF
C9152 PAND2X1_479/B POR2X1_329/A 0.02fF
C9153 POR2X1_54/Y POR2X1_94/A 1.19fF
C9154 POR2X1_282/Y VDD 0.13fF
C9155 POR2X1_19/a_16_28# POR2X1_5/Y 0.01fF
C9156 PAND2X1_63/O POR2X1_296/B 0.05fF
C9157 POR2X1_333/A PAND2X1_91/a_76_28# 0.03fF
C9158 POR2X1_4/Y POR2X1_294/A 0.03fF
C9159 PAND2X1_510/B POR2X1_80/a_56_344# 0.00fF
C9160 POR2X1_209/A POR2X1_535/a_56_344# 0.00fF
C9161 POR2X1_257/A PAND2X1_725/B 0.02fF
C9162 POR2X1_801/B POR2X1_121/B 0.06fF
C9163 PAND2X1_20/A POR2X1_34/B 0.02fF
C9164 POR2X1_20/B POR2X1_79/A 0.37fF
C9165 POR2X1_728/B POR2X1_467/a_16_28# 0.03fF
C9166 PAND2X1_340/B POR2X1_381/CTRL 0.01fF
C9167 PAND2X1_219/A POR2X1_32/A 0.03fF
C9168 PAND2X1_255/O PAND2X1_69/A 0.06fF
C9169 POR2X1_471/A POR2X1_724/CTRL2 0.01fF
C9170 PAND2X1_93/B POR2X1_274/Y 0.05fF
C9171 PAND2X1_557/A POR2X1_487/CTRL 0.08fF
C9172 POR2X1_476/A POR2X1_734/A 0.07fF
C9173 POR2X1_292/Y POR2X1_7/B 0.03fF
C9174 POR2X1_804/a_76_344# POR2X1_330/Y 0.03fF
C9175 POR2X1_556/A POR2X1_193/A 12.58fF
C9176 POR2X1_48/A PAND2X1_562/B 0.07fF
C9177 POR2X1_556/A POR2X1_579/Y 0.03fF
C9178 POR2X1_60/A POR2X1_432/a_76_344# 0.01fF
C9179 POR2X1_389/A PAND2X1_607/O 0.01fF
C9180 PAND2X1_805/O PAND2X1_287/Y 0.02fF
C9181 POR2X1_163/O POR2X1_48/A 0.00fF
C9182 POR2X1_555/B POR2X1_750/B 0.05fF
C9183 POR2X1_556/A POR2X1_572/B 0.04fF
C9184 PAND2X1_865/O PAND2X1_860/A 0.04fF
C9185 POR2X1_130/A POR2X1_606/O 0.32fF
C9186 POR2X1_708/a_16_28# PAND2X1_39/B 0.03fF
C9187 PAND2X1_796/B POR2X1_293/Y 0.02fF
C9188 POR2X1_644/Y VDD 0.04fF
C9189 POR2X1_287/A POR2X1_249/CTRL 0.01fF
C9190 PAND2X1_319/a_16_344# POR2X1_48/A 0.02fF
C9191 PAND2X1_831/O POR2X1_102/Y 0.03fF
C9192 POR2X1_49/Y POR2X1_442/Y 0.02fF
C9193 POR2X1_66/A POR2X1_206/A 0.02fF
C9194 POR2X1_294/O POR2X1_294/B 0.17fF
C9195 POR2X1_648/Y POR2X1_307/A 0.00fF
C9196 POR2X1_68/A POR2X1_831/CTRL2 0.01fF
C9197 PAND2X1_48/B PAND2X1_487/CTRL2 0.00fF
C9198 POR2X1_474/CTRL2 POR2X1_860/A 0.01fF
C9199 POR2X1_614/A POR2X1_556/A 0.22fF
C9200 POR2X1_262/Y POR2X1_52/Y 0.03fF
C9201 PAND2X1_478/Y PAND2X1_478/B 0.01fF
C9202 POR2X1_547/CTRL POR2X1_624/Y 0.00fF
C9203 POR2X1_491/CTRL PAND2X1_558/Y 0.00fF
C9204 POR2X1_13/A POR2X1_48/A 0.43fF
C9205 POR2X1_750/B POR2X1_330/Y 0.05fF
C9206 PAND2X1_71/a_76_28# PAND2X1_39/B 0.01fF
C9207 POR2X1_39/CTRL2 POR2X1_72/B 0.03fF
C9208 PAND2X1_656/CTRL VDD 0.00fF
C9209 POR2X1_499/A PAND2X1_96/B 0.00fF
C9210 POR2X1_774/Y POR2X1_866/O 0.02fF
C9211 PAND2X1_37/CTRL2 PAND2X1_8/Y 0.02fF
C9212 POR2X1_65/A PAND2X1_557/A 0.03fF
C9213 POR2X1_23/Y POR2X1_293/Y 0.30fF
C9214 POR2X1_471/a_16_28# POR2X1_66/A 0.02fF
C9215 POR2X1_341/A POR2X1_341/a_76_344# 0.03fF
C9216 POR2X1_649/B POR2X1_649/a_56_344# 0.01fF
C9217 PAND2X1_466/A PAND2X1_241/Y 0.01fF
C9218 POR2X1_677/CTRL PAND2X1_390/Y 0.01fF
C9219 POR2X1_20/B PAND2X1_785/A 0.05fF
C9220 PAND2X1_219/A PAND2X1_741/B 0.01fF
C9221 PAND2X1_793/Y POR2X1_487/CTRL2 0.01fF
C9222 POR2X1_20/B POR2X1_291/Y 0.01fF
C9223 POR2X1_270/Y POR2X1_659/CTRL2 0.01fF
C9224 POR2X1_231/A POR2X1_186/Y 0.01fF
C9225 PAND2X1_865/a_16_344# POR2X1_329/A 0.01fF
C9226 POR2X1_56/CTRL2 PAND2X1_254/Y 0.01fF
C9227 PAND2X1_23/Y PAND2X1_94/O 0.00fF
C9228 POR2X1_629/B VDD 0.13fF
C9229 POR2X1_175/a_16_28# POR2X1_78/A 0.01fF
C9230 POR2X1_416/Y PAND2X1_606/O 0.02fF
C9231 D_INPUT_0 PAND2X1_351/a_16_344# 0.06fF
C9232 POR2X1_849/A POR2X1_546/B 0.11fF
C9233 POR2X1_78/B POR2X1_400/O 0.02fF
C9234 PAND2X1_445/Y POR2X1_102/Y 0.01fF
C9235 PAND2X1_23/Y POR2X1_466/A 0.03fF
C9236 POR2X1_567/B D_GATE_662 0.10fF
C9237 D_INPUT_3 POR2X1_612/CTRL 0.01fF
C9238 POR2X1_188/A POR2X1_285/CTRL 0.01fF
C9239 POR2X1_68/A POR2X1_849/B 0.01fF
C9240 PAND2X1_95/B PAND2X1_51/a_16_344# 0.02fF
C9241 POR2X1_502/A PAND2X1_279/CTRL 0.01fF
C9242 PAND2X1_96/B POR2X1_76/A 0.03fF
C9243 POR2X1_68/A PAND2X1_94/CTRL 0.07fF
C9244 PAND2X1_390/Y POR2X1_236/Y 0.12fF
C9245 PAND2X1_787/A PAND2X1_211/CTRL 0.00fF
C9246 PAND2X1_219/A PAND2X1_35/Y 0.01fF
C9247 PAND2X1_475/O INPUT_0 0.05fF
C9248 POR2X1_360/A POR2X1_243/A 0.01fF
C9249 PAND2X1_659/CTRL POR2X1_72/B 0.01fF
C9250 PAND2X1_137/Y POR2X1_60/A 0.07fF
C9251 POR2X1_605/A POR2X1_260/B 0.03fF
C9252 PAND2X1_695/O PAND2X1_41/B 0.01fF
C9253 POR2X1_121/A PAND2X1_666/O 0.00fF
C9254 POR2X1_609/CTRL POR2X1_609/A 0.01fF
C9255 POR2X1_78/B POR2X1_456/CTRL2 0.19fF
C9256 POR2X1_388/CTRL2 POR2X1_66/A 0.00fF
C9257 POR2X1_776/A POR2X1_854/B 0.05fF
C9258 INPUT_3 PAND2X1_63/B 0.03fF
C9259 POR2X1_296/B POR2X1_575/B 0.17fF
C9260 POR2X1_616/Y POR2X1_9/Y 0.22fF
C9261 POR2X1_78/B PAND2X1_52/Y 0.05fF
C9262 POR2X1_811/A POR2X1_796/CTRL 0.00fF
C9263 POR2X1_397/Y POR2X1_5/Y 0.02fF
C9264 POR2X1_48/A PAND2X1_553/CTRL2 0.01fF
C9265 PAND2X1_661/B POR2X1_48/A 0.00fF
C9266 PAND2X1_118/CTRL POR2X1_78/A 0.01fF
C9267 PAND2X1_793/Y POR2X1_40/Y 0.03fF
C9268 PAND2X1_420/CTRL POR2X1_294/B 0.02fF
C9269 POR2X1_48/A PAND2X1_643/Y 0.00fF
C9270 POR2X1_222/CTRL2 POR2X1_222/A 0.01fF
C9271 POR2X1_432/Y VDD 0.00fF
C9272 PAND2X1_90/Y POR2X1_770/A 0.02fF
C9273 POR2X1_697/CTRL POR2X1_236/Y 0.01fF
C9274 PAND2X1_733/A POR2X1_597/A 0.00fF
C9275 POR2X1_52/A POR2X1_491/O 0.16fF
C9276 POR2X1_49/Y PAND2X1_661/O 0.02fF
C9277 POR2X1_32/A POR2X1_816/A 0.06fF
C9278 PAND2X1_90/Y POR2X1_793/a_76_344# 0.09fF
C9279 POR2X1_719/CTRL2 POR2X1_66/A 0.01fF
C9280 POR2X1_130/A POR2X1_480/A 0.10fF
C9281 PAND2X1_7/CTRL2 POR2X1_750/B 0.14fF
C9282 POR2X1_558/B PAND2X1_60/B 0.03fF
C9283 POR2X1_66/B POR2X1_790/B 0.03fF
C9284 POR2X1_96/A PAND2X1_192/O 0.03fF
C9285 D_INPUT_2 POR2X1_293/CTRL2 0.01fF
C9286 POR2X1_677/Y PAND2X1_840/Y 0.03fF
C9287 POR2X1_669/B POR2X1_321/a_16_28# 0.09fF
C9288 PAND2X1_73/Y PAND2X1_79/Y 0.07fF
C9289 POR2X1_128/A POR2X1_222/Y 0.07fF
C9290 POR2X1_22/A POR2X1_750/B 0.01fF
C9291 POR2X1_356/A PAND2X1_65/B 0.15fF
C9292 POR2X1_856/B POR2X1_854/B 0.01fF
C9293 POR2X1_43/B POR2X1_72/B 1.37fF
C9294 POR2X1_263/Y POR2X1_235/O 0.01fF
C9295 PAND2X1_658/A PAND2X1_185/O 0.01fF
C9296 PAND2X1_429/Y VDD 0.12fF
C9297 POR2X1_7/B PAND2X1_366/Y 0.03fF
C9298 POR2X1_48/A POR2X1_321/Y 0.05fF
C9299 POR2X1_368/CTRL2 POR2X1_293/Y 0.01fF
C9300 PAND2X1_7/O PAND2X1_52/Y 0.02fF
C9301 POR2X1_423/Y POR2X1_183/Y 0.04fF
C9302 POR2X1_78/A POR2X1_216/O 0.02fF
C9303 PAND2X1_85/Y POR2X1_294/B 0.00fF
C9304 PAND2X1_90/Y POR2X1_740/Y 0.05fF
C9305 POR2X1_840/B PAND2X1_74/O 0.10fF
C9306 PAND2X1_621/O POR2X1_818/Y 0.01fF
C9307 POR2X1_15/CTRL2 POR2X1_69/A 0.01fF
C9308 PAND2X1_211/a_16_344# PAND2X1_853/B 0.02fF
C9309 POR2X1_498/O PAND2X1_735/Y 0.06fF
C9310 PAND2X1_675/A POR2X1_106/Y 0.03fF
C9311 POR2X1_391/A POR2X1_816/A 0.03fF
C9312 POR2X1_16/A PAND2X1_571/CTRL2 0.21fF
C9313 PAND2X1_390/Y PAND2X1_858/Y 0.17fF
C9314 POR2X1_14/Y POR2X1_387/Y 0.02fF
C9315 POR2X1_7/B POR2X1_295/Y 1.19fF
C9316 POR2X1_829/a_76_344# POR2X1_761/Y 0.00fF
C9317 POR2X1_433/CTRL2 PAND2X1_349/A 0.01fF
C9318 INPUT_1 POR2X1_66/A 0.07fF
C9319 POR2X1_78/A PAND2X1_63/B 0.03fF
C9320 PAND2X1_94/A PAND2X1_15/CTRL2 0.00fF
C9321 PAND2X1_90/A POR2X1_130/A 0.08fF
C9322 PAND2X1_658/B POR2X1_511/Y 1.68fF
C9323 PAND2X1_58/A PAND2X1_306/a_56_28# 0.00fF
C9324 POR2X1_164/CTRL POR2X1_376/B 0.01fF
C9325 PAND2X1_730/B POR2X1_42/Y 0.39fF
C9326 PAND2X1_23/Y PAND2X1_131/CTRL 0.01fF
C9327 PAND2X1_48/B PAND2X1_131/O 0.04fF
C9328 POR2X1_128/A POR2X1_532/A 0.01fF
C9329 POR2X1_333/CTRL POR2X1_241/B 0.01fF
C9330 GATE_741 POR2X1_42/Y 0.03fF
C9331 POR2X1_580/a_16_28# POR2X1_579/Y 0.03fF
C9332 D_GATE_222 PAND2X1_164/O 0.09fF
C9333 POR2X1_710/A PAND2X1_69/A 0.01fF
C9334 PAND2X1_661/Y POR2X1_102/Y 0.03fF
C9335 PAND2X1_185/O POR2X1_73/Y 0.15fF
C9336 POR2X1_8/Y POR2X1_409/B 0.07fF
C9337 PAND2X1_798/B PAND2X1_804/A 0.02fF
C9338 POR2X1_13/A PAND2X1_197/Y 0.16fF
C9339 PAND2X1_675/A PAND2X1_580/B 0.03fF
C9340 PAND2X1_257/CTRL2 POR2X1_222/Y 0.03fF
C9341 PAND2X1_469/B PAND2X1_580/B 0.02fF
C9342 POR2X1_750/a_16_28# POR2X1_750/A 0.04fF
C9343 POR2X1_65/A PAND2X1_553/O 0.08fF
C9344 POR2X1_710/A POR2X1_710/a_16_28# 0.12fF
C9345 POR2X1_164/Y POR2X1_83/B 0.01fF
C9346 POR2X1_399/a_16_28# POR2X1_399/A 0.03fF
C9347 POR2X1_254/O POR2X1_228/Y 0.03fF
C9348 POR2X1_241/B POR2X1_502/O 0.03fF
C9349 PAND2X1_6/A PAND2X1_8/Y 0.72fF
C9350 POR2X1_174/B POR2X1_174/CTRL 0.05fF
C9351 POR2X1_859/A POR2X1_790/B 0.13fF
C9352 POR2X1_502/A PAND2X1_411/CTRL2 0.03fF
C9353 POR2X1_41/B POR2X1_846/B 0.02fF
C9354 POR2X1_750/B PAND2X1_158/CTRL 0.01fF
C9355 POR2X1_78/B D_INPUT_1 0.07fF
C9356 POR2X1_140/B PAND2X1_57/B 0.03fF
C9357 PAND2X1_61/Y PAND2X1_338/B 0.00fF
C9358 PAND2X1_23/Y PAND2X1_371/O 0.10fF
C9359 POR2X1_137/Y POR2X1_650/A 0.03fF
C9360 POR2X1_364/A VDD 0.45fF
C9361 POR2X1_407/A PAND2X1_57/B 0.07fF
C9362 INPUT_0 POR2X1_576/Y 0.03fF
C9363 POR2X1_777/B POR2X1_569/A 0.10fF
C9364 PAND2X1_845/O PAND2X1_673/Y 0.00fF
C9365 POR2X1_813/CTRL POR2X1_39/B 0.25fF
C9366 POR2X1_343/Y PAND2X1_256/a_76_28# 0.02fF
C9367 POR2X1_581/CTRL INPUT_5 0.01fF
C9368 POR2X1_750/B POR2X1_799/O 0.01fF
C9369 PAND2X1_434/CTRL POR2X1_72/B 0.00fF
C9370 POR2X1_416/B POR2X1_150/Y 0.03fF
C9371 POR2X1_78/B POR2X1_724/A 1.13fF
C9372 PAND2X1_671/CTRL2 POR2X1_35/B 0.01fF
C9373 D_INPUT_0 POR2X1_550/B 0.02fF
C9374 PAND2X1_391/O POR2X1_384/Y 0.07fF
C9375 POR2X1_590/A POR2X1_741/A 0.00fF
C9376 POR2X1_14/Y POR2X1_419/a_16_28# 0.08fF
C9377 POR2X1_62/Y PAND2X1_10/CTRL 0.01fF
C9378 POR2X1_220/Y POR2X1_702/A 0.03fF
C9379 PAND2X1_340/O POR2X1_7/A 0.01fF
C9380 POR2X1_550/A PAND2X1_525/O 0.02fF
C9381 POR2X1_802/a_16_28# POR2X1_750/B 0.02fF
C9382 POR2X1_844/O VDD 0.00fF
C9383 PAND2X1_294/CTRL POR2X1_39/B 0.01fF
C9384 POR2X1_575/B POR2X1_501/O 0.04fF
C9385 POR2X1_327/Y POR2X1_830/Y 0.03fF
C9386 PAND2X1_453/A POR2X1_419/a_16_28# 0.01fF
C9387 POR2X1_174/A POR2X1_564/B 0.03fF
C9388 POR2X1_35/Y POR2X1_785/A 0.06fF
C9389 PAND2X1_643/CTRL POR2X1_13/Y 0.01fF
C9390 POR2X1_262/CTRL2 POR2X1_73/Y 0.01fF
C9391 PAND2X1_610/CTRL2 POR2X1_48/A 0.03fF
C9392 POR2X1_287/B POR2X1_101/Y 0.03fF
C9393 POR2X1_60/A PAND2X1_853/B 0.03fF
C9394 PAND2X1_65/B POR2X1_569/A 0.07fF
C9395 PAND2X1_836/O POR2X1_293/Y 0.15fF
C9396 POR2X1_548/B POR2X1_614/A 0.03fF
C9397 POR2X1_67/CTRL2 POR2X1_39/B 0.16fF
C9398 PAND2X1_90/A POR2X1_844/B 0.03fF
C9399 PAND2X1_592/Y POR2X1_594/A 0.06fF
C9400 PAND2X1_469/Y VDD -0.00fF
C9401 POR2X1_504/Y POR2X1_260/A 0.03fF
C9402 POR2X1_455/A POR2X1_222/Y 0.03fF
C9403 PAND2X1_653/Y PAND2X1_215/B 0.07fF
C9404 POR2X1_669/O POR2X1_73/Y 0.02fF
C9405 PAND2X1_55/Y PAND2X1_29/O 0.01fF
C9406 PAND2X1_481/CTRL2 POR2X1_355/A 0.01fF
C9407 POR2X1_496/Y PAND2X1_506/Y 1.51fF
C9408 POR2X1_332/B PAND2X1_60/B 1.09fF
C9409 PAND2X1_48/B POR2X1_219/O 0.01fF
C9410 PAND2X1_698/CTRL PAND2X1_65/B 0.01fF
C9411 POR2X1_46/Y POR2X1_91/Y 0.03fF
C9412 POR2X1_68/A POR2X1_523/Y 0.94fF
C9413 POR2X1_189/Y POR2X1_816/A 0.04fF
C9414 PAND2X1_96/B PAND2X1_132/O 0.01fF
C9415 PAND2X1_621/Y POR2X1_619/Y 0.01fF
C9416 PAND2X1_217/B POR2X1_394/A 0.19fF
C9417 POR2X1_42/Y POR2X1_748/CTRL 0.13fF
C9418 POR2X1_666/Y POR2X1_394/A 0.12fF
C9419 POR2X1_336/CTRL POR2X1_740/Y 0.01fF
C9420 POR2X1_417/Y PAND2X1_357/CTRL 0.01fF
C9421 PAND2X1_865/Y PAND2X1_794/CTRL2 0.00fF
C9422 PAND2X1_90/A PAND2X1_150/O 0.01fF
C9423 PAND2X1_723/Y POR2X1_7/O 0.15fF
C9424 POR2X1_78/A POR2X1_552/A 0.05fF
C9425 POR2X1_68/A POR2X1_219/CTRL2 0.01fF
C9426 POR2X1_400/O POR2X1_294/A 0.16fF
C9427 PAND2X1_279/CTRL POR2X1_188/Y 0.01fF
C9428 POR2X1_249/Y VDD 0.19fF
C9429 POR2X1_370/CTRL2 POR2X1_543/A 0.01fF
C9430 POR2X1_68/A PAND2X1_69/A 0.27fF
C9431 POR2X1_407/A POR2X1_828/A 0.43fF
C9432 POR2X1_137/Y POR2X1_294/B 0.05fF
C9433 POR2X1_54/a_16_28# PAND2X1_58/A 0.02fF
C9434 PAND2X1_94/A INPUT_0 3.32fF
C9435 PAND2X1_23/Y POR2X1_478/B 0.03fF
C9436 PAND2X1_651/Y POR2X1_816/A 0.05fF
C9437 POR2X1_55/Y POR2X1_387/Y 0.21fF
C9438 PAND2X1_539/Y INPUT_0 0.09fF
C9439 POR2X1_66/B POR2X1_540/Y 0.02fF
C9440 POR2X1_672/CTRL2 POR2X1_38/B 0.01fF
C9441 POR2X1_278/Y POR2X1_187/O 0.05fF
C9442 POR2X1_114/CTRL2 POR2X1_68/B 0.01fF
C9443 POR2X1_313/CTRL2 POR2X1_90/Y 0.03fF
C9444 PAND2X1_174/O POR2X1_172/Y 0.00fF
C9445 POR2X1_781/a_16_28# POR2X1_568/Y 0.07fF
C9446 POR2X1_466/A POR2X1_711/Y 0.10fF
C9447 PAND2X1_804/B PAND2X1_175/O 0.04fF
C9448 PAND2X1_386/Y POR2X1_707/Y 0.15fF
C9449 POR2X1_750/B POR2X1_337/Y 0.09fF
C9450 PAND2X1_106/O PAND2X1_48/B 0.15fF
C9451 PAND2X1_90/Y POR2X1_774/A 0.14fF
C9452 POR2X1_90/Y POR2X1_700/Y 0.73fF
C9453 POR2X1_707/O PAND2X1_57/B 0.18fF
C9454 PAND2X1_658/A POR2X1_530/Y 0.02fF
C9455 POR2X1_29/A POR2X1_39/B 0.20fF
C9456 PAND2X1_104/a_16_344# POR2X1_4/Y 0.00fF
C9457 POR2X1_94/A POR2X1_4/Y 0.16fF
C9458 PAND2X1_23/Y POR2X1_274/B 0.05fF
C9459 POR2X1_315/Y PAND2X1_724/B 0.07fF
C9460 POR2X1_460/A PAND2X1_69/A 0.03fF
C9461 POR2X1_394/A VDD 9.94fF
C9462 POR2X1_332/B POR2X1_332/O 0.03fF
C9463 POR2X1_574/CTRL POR2X1_574/A 0.01fF
C9464 POR2X1_528/CTRL POR2X1_528/Y 0.01fF
C9465 PAND2X1_96/B POR2X1_540/A 0.00fF
C9466 PAND2X1_675/A PAND2X1_349/A 0.03fF
C9467 PAND2X1_469/B PAND2X1_349/A 0.03fF
C9468 POR2X1_333/Y POR2X1_192/Y 0.05fF
C9469 POR2X1_118/O POR2X1_278/A 0.04fF
C9470 PAND2X1_850/Y POR2X1_423/Y 0.09fF
C9471 POR2X1_687/A POR2X1_803/A 0.35fF
C9472 POR2X1_48/a_16_28# PAND2X1_123/Y 0.02fF
C9473 POR2X1_119/Y POR2X1_122/A 0.02fF
C9474 POR2X1_532/A POR2X1_140/O 0.02fF
C9475 POR2X1_545/A POR2X1_180/A 0.07fF
C9476 POR2X1_270/CTRL POR2X1_724/A 0.05fF
C9477 PAND2X1_759/m4_208_n4# PAND2X1_48/A 0.04fF
C9478 PAND2X1_675/A PAND2X1_114/B 0.15fF
C9479 POR2X1_62/Y PAND2X1_474/Y 0.02fF
C9480 POR2X1_391/CTRL POR2X1_816/A 0.00fF
C9481 POR2X1_49/Y PAND2X1_326/B 0.06fF
C9482 POR2X1_16/A POR2X1_42/Y 0.43fF
C9483 POR2X1_786/Y POR2X1_366/A 0.07fF
C9484 POR2X1_491/Y PAND2X1_558/Y 0.02fF
C9485 PAND2X1_199/A PAND2X1_199/O 0.00fF
C9486 POR2X1_833/A POR2X1_294/B 0.27fF
C9487 POR2X1_529/Y PAND2X1_548/O 0.00fF
C9488 POR2X1_167/CTRL POR2X1_90/Y 0.08fF
C9489 POR2X1_197/Y POR2X1_532/A 0.02fF
C9490 POR2X1_3/A POR2X1_3/a_16_28# 0.02fF
C9491 POR2X1_23/Y PAND2X1_242/Y 0.10fF
C9492 POR2X1_62/Y POR2X1_13/A 0.02fF
C9493 POR2X1_131/Y PAND2X1_190/Y 0.33fF
C9494 POR2X1_356/A POR2X1_174/a_16_28# 0.12fF
C9495 POR2X1_502/A POR2X1_737/A 0.03fF
C9496 PAND2X1_6/Y PAND2X1_528/O 0.03fF
C9497 PAND2X1_4/m4_208_n4# D_INPUT_1 0.01fF
C9498 POR2X1_494/Y POR2X1_153/Y 0.03fF
C9499 POR2X1_60/A POR2X1_80/O 0.01fF
C9500 POR2X1_773/B POR2X1_391/Y 0.10fF
C9501 POR2X1_383/A POR2X1_865/O 0.02fF
C9502 PAND2X1_803/Y PAND2X1_388/Y 0.02fF
C9503 POR2X1_180/B PAND2X1_69/A 0.01fF
C9504 POR2X1_802/O POR2X1_532/A 0.01fF
C9505 POR2X1_46/Y POR2X1_109/Y 0.05fF
C9506 PAND2X1_738/CTRL2 POR2X1_39/B 0.04fF
C9507 POR2X1_249/Y PAND2X1_32/B 0.10fF
C9508 D_INPUT_3 POR2X1_283/A 0.03fF
C9509 POR2X1_59/CTRL2 POR2X1_90/Y 0.01fF
C9510 POR2X1_68/A PAND2X1_824/B 0.07fF
C9511 POR2X1_840/B POR2X1_276/Y 0.05fF
C9512 POR2X1_652/Y POR2X1_802/A 0.01fF
C9513 PAND2X1_845/a_76_28# POR2X1_813/Y 0.07fF
C9514 POR2X1_826/CTRL2 POR2X1_77/Y 0.00fF
C9515 POR2X1_41/CTRL2 POR2X1_73/Y 0.03fF
C9516 POR2X1_24/a_76_344# POR2X1_77/Y 0.01fF
C9517 PAND2X1_658/B POR2X1_129/Y 0.03fF
C9518 POR2X1_62/Y PAND2X1_197/O 0.02fF
C9519 POR2X1_130/A PAND2X1_304/O 0.04fF
C9520 POR2X1_57/A POR2X1_527/CTRL 0.01fF
C9521 POR2X1_299/CTRL2 PAND2X1_308/Y 0.01fF
C9522 POR2X1_35/Y POR2X1_186/B 0.03fF
C9523 INPUT_1 POR2X1_532/A 0.08fF
C9524 PAND2X1_6/Y POR2X1_544/B 0.03fF
C9525 POR2X1_777/B PAND2X1_72/A 0.05fF
C9526 POR2X1_456/B POR2X1_736/CTRL 0.01fF
C9527 D_INPUT_6 POR2X1_260/A 0.03fF
C9528 PAND2X1_727/CTRL2 POR2X1_91/Y 0.01fF
C9529 PAND2X1_801/CTRL PAND2X1_863/B 0.01fF
C9530 POR2X1_305/Y PAND2X1_156/A 0.08fF
C9531 POR2X1_809/A POR2X1_149/B 0.02fF
C9532 POR2X1_49/Y POR2X1_387/a_16_28# 0.03fF
C9533 PAND2X1_661/Y PAND2X1_194/a_56_28# 0.00fF
C9534 POR2X1_814/A POR2X1_647/O 0.60fF
C9535 PAND2X1_449/a_16_344# POR2X1_424/Y 0.02fF
C9536 PAND2X1_631/A PAND2X1_465/B 0.01fF
C9537 PAND2X1_744/CTRL2 POR2X1_294/A 0.02fF
C9538 POR2X1_63/O POR2X1_62/Y 0.03fF
C9539 POR2X1_260/B POR2X1_646/B 0.10fF
C9540 POR2X1_821/O POR2X1_39/B 0.16fF
C9541 POR2X1_546/A POR2X1_39/B 0.01fF
C9542 POR2X1_833/A PAND2X1_111/B 0.03fF
C9543 PAND2X1_65/B PAND2X1_72/A 6.41fF
C9544 POR2X1_162/Y POR2X1_260/A 0.00fF
C9545 POR2X1_447/B POR2X1_66/CTRL2 0.04fF
C9546 POR2X1_845/O POR2X1_673/Y 0.01fF
C9547 POR2X1_294/A POR2X1_816/A 0.06fF
C9548 PAND2X1_632/A PAND2X1_508/CTRL 0.01fF
C9549 POR2X1_809/A POR2X1_644/A 0.28fF
C9550 D_INPUT_1 POR2X1_294/A 23.85fF
C9551 POR2X1_410/CTRL PAND2X1_52/B 0.01fF
C9552 POR2X1_366/O POR2X1_276/Y 0.09fF
C9553 POR2X1_257/A POR2X1_253/O 0.01fF
C9554 POR2X1_68/B POR2X1_773/A 0.03fF
C9555 PAND2X1_723/O POR2X1_7/Y 0.02fF
C9556 POR2X1_863/A POR2X1_436/a_16_28# 0.03fF
C9557 PAND2X1_127/CTRL2 POR2X1_456/B 0.11fF
C9558 POR2X1_462/O POR2X1_66/A 0.01fF
C9559 POR2X1_416/B PAND2X1_364/B 0.07fF
C9560 POR2X1_814/A POR2X1_210/O 0.33fF
C9561 POR2X1_304/CTRL POR2X1_43/B 0.01fF
C9562 POR2X1_12/A POR2X1_257/A 0.03fF
C9563 PAND2X1_621/a_16_344# POR2X1_750/Y 0.02fF
C9564 PAND2X1_341/B POR2X1_38/Y 0.91fF
C9565 POR2X1_48/A POR2X1_412/CTRL 0.00fF
C9566 PAND2X1_65/B POR2X1_535/O 0.02fF
C9567 PAND2X1_831/O POR2X1_677/Y 0.00fF
C9568 POR2X1_76/Y POR2X1_715/O 0.02fF
C9569 PAND2X1_634/CTRL POR2X1_37/Y 0.03fF
C9570 PAND2X1_628/O POR2X1_61/Y 0.01fF
C9571 PAND2X1_426/O POR2X1_121/B 0.02fF
C9572 POR2X1_263/Y POR2X1_20/B 0.03fF
C9573 POR2X1_814/B PAND2X1_607/CTRL2 0.01fF
C9574 POR2X1_146/a_16_28# POR2X1_394/A 0.03fF
C9575 POR2X1_311/CTRL2 PAND2X1_336/Y 0.01fF
C9576 VDD POR2X1_91/CTRL -0.00fF
C9577 PAND2X1_69/A POR2X1_169/A 0.03fF
C9578 POR2X1_667/a_16_28# POR2X1_667/A 0.03fF
C9579 POR2X1_59/O POR2X1_394/A 0.01fF
C9580 POR2X1_848/CTRL2 POR2X1_734/A 0.03fF
C9581 POR2X1_864/A PAND2X1_829/CTRL2 0.00fF
C9582 PAND2X1_508/Y PAND2X1_861/O 0.04fF
C9583 POR2X1_741/Y POR2X1_715/CTRL 0.01fF
C9584 POR2X1_740/Y POR2X1_715/O 0.06fF
C9585 POR2X1_556/A POR2X1_590/A 0.01fF
C9586 POR2X1_817/a_76_344# PAND2X1_340/B 0.00fF
C9587 INPUT_3 POR2X1_32/A 0.10fF
C9588 PAND2X1_846/CTRL2 POR2X1_38/B 0.03fF
C9589 POR2X1_14/Y POR2X1_88/A 0.05fF
C9590 POR2X1_568/Y POR2X1_738/O 0.38fF
C9591 POR2X1_51/O POR2X1_51/B 0.01fF
C9592 POR2X1_621/A POR2X1_29/A 0.00fF
C9593 POR2X1_66/B POR2X1_658/O 0.01fF
C9594 POR2X1_76/CTRL POR2X1_296/B 0.01fF
C9595 POR2X1_428/Y POR2X1_32/A 0.01fF
C9596 POR2X1_685/CTRL2 POR2X1_814/A 0.02fF
C9597 PAND2X1_661/Y POR2X1_761/A 0.36fF
C9598 POR2X1_434/O POR2X1_434/A 0.03fF
C9599 POR2X1_715/CTRL PAND2X1_32/B 0.16fF
C9600 POR2X1_431/O POR2X1_5/Y 0.02fF
C9601 POR2X1_271/Y POR2X1_411/B 0.01fF
C9602 PAND2X1_76/a_16_344# POR2X1_20/B 0.01fF
C9603 POR2X1_467/a_16_28# POR2X1_330/Y 0.04fF
C9604 PAND2X1_603/CTRL POR2X1_260/B 0.01fF
C9605 POR2X1_651/Y POR2X1_725/m4_208_n4# 0.08fF
C9606 POR2X1_90/Y PAND2X1_326/a_76_28# 0.02fF
C9607 POR2X1_343/Y POR2X1_575/CTRL 0.11fF
C9608 PAND2X1_613/O POR2X1_29/A 0.06fF
C9609 POR2X1_60/A PAND2X1_454/B 0.05fF
C9610 PAND2X1_341/B POR2X1_153/Y 0.05fF
C9611 PAND2X1_832/CTRL2 POR2X1_271/B 0.01fF
C9612 POR2X1_848/CTRL POR2X1_859/A 0.05fF
C9613 POR2X1_744/CTRL2 POR2X1_39/B 0.00fF
C9614 POR2X1_554/B POR2X1_217/CTRL2 0.03fF
C9615 PAND2X1_809/B PAND2X1_539/Y 0.72fF
C9616 POR2X1_66/B POR2X1_445/A 0.09fF
C9617 PAND2X1_737/B PAND2X1_198/CTRL 0.01fF
C9618 PAND2X1_202/CTRL POR2X1_67/Y 0.01fF
C9619 PAND2X1_202/O POR2X1_69/Y 0.01fF
C9620 PAND2X1_404/Y POR2X1_667/A 0.08fF
C9621 POR2X1_560/Y POR2X1_561/Y 0.00fF
C9622 POR2X1_66/B POR2X1_643/Y 0.00fF
C9623 POR2X1_48/A POR2X1_29/A 0.06fF
C9624 POR2X1_48/A POR2X1_163/Y 0.01fF
C9625 PAND2X1_862/a_16_344# POR2X1_91/Y 0.01fF
C9626 POR2X1_737/A POR2X1_188/Y 0.01fF
C9627 POR2X1_376/B PAND2X1_449/m4_208_n4# 0.15fF
C9628 POR2X1_814/B POR2X1_663/B 0.03fF
C9629 POR2X1_849/B PAND2X1_58/A 0.01fF
C9630 PAND2X1_628/O POR2X1_35/Y 0.02fF
C9631 POR2X1_376/B POR2X1_411/B 0.08fF
C9632 POR2X1_856/B PAND2X1_73/Y 0.03fF
C9633 POR2X1_567/B POR2X1_78/A 0.05fF
C9634 PAND2X1_96/CTRL2 POR2X1_202/A 0.02fF
C9635 PAND2X1_94/CTRL PAND2X1_58/A 0.01fF
C9636 POR2X1_678/A POR2X1_260/B 0.09fF
C9637 POR2X1_188/A POR2X1_643/Y 0.01fF
C9638 POR2X1_356/A POR2X1_814/A 0.10fF
C9639 POR2X1_23/Y POR2X1_60/A 7.47fF
C9640 POR2X1_679/O VDD 0.00fF
C9641 POR2X1_323/a_16_28# POR2X1_485/Y 0.02fF
C9642 POR2X1_90/Y POR2X1_91/a_16_28# 0.03fF
C9643 POR2X1_34/O POR2X1_94/A 0.07fF
C9644 POR2X1_582/Y POR2X1_763/A 0.01fF
C9645 PAND2X1_201/a_16_344# INPUT_0 0.04fF
C9646 POR2X1_519/CTRL POR2X1_43/Y 0.00fF
C9647 POR2X1_83/B PAND2X1_392/O 0.01fF
C9648 POR2X1_150/Y PAND2X1_738/Y 0.05fF
C9649 POR2X1_846/Y POR2X1_754/A 0.30fF
C9650 POR2X1_630/CTRL POR2X1_750/B 0.14fF
C9651 POR2X1_260/B PAND2X1_13/CTRL 0.01fF
C9652 POR2X1_669/B POR2X1_819/O 0.09fF
C9653 POR2X1_48/A PAND2X1_554/O 0.10fF
C9654 POR2X1_541/B PAND2X1_48/O 0.01fF
C9655 PAND2X1_848/O POR2X1_669/B 0.19fF
C9656 POR2X1_260/O POR2X1_740/Y 0.02fF
C9657 POR2X1_260/CTRL POR2X1_741/Y 0.00fF
C9658 POR2X1_66/A POR2X1_200/CTRL 0.01fF
C9659 PAND2X1_658/A PAND2X1_414/CTRL 0.01fF
C9660 GATE_479 PAND2X1_776/Y 0.37fF
C9661 POR2X1_48/A POR2X1_820/A 0.01fF
C9662 POR2X1_48/A PAND2X1_738/CTRL2 0.03fF
C9663 POR2X1_415/A POR2X1_415/CTRL 0.06fF
C9664 POR2X1_127/Y PAND2X1_771/Y 0.03fF
C9665 D_INPUT_0 POR2X1_780/O 0.16fF
C9666 POR2X1_38/O POR2X1_5/Y 0.01fF
C9667 POR2X1_544/B PAND2X1_52/B 0.08fF
C9668 POR2X1_52/A POR2X1_411/B 0.08fF
C9669 POR2X1_485/a_56_344# PAND2X1_550/B 0.00fF
C9670 POR2X1_324/A POR2X1_220/B 0.01fF
C9671 PAND2X1_458/O POR2X1_387/Y 0.07fF
C9672 POR2X1_37/Y PAND2X1_333/CTRL 0.06fF
C9673 POR2X1_609/Y PAND2X1_240/O 0.00fF
C9674 GATE_579 VDD 0.00fF
C9675 PAND2X1_475/O POR2X1_102/Y 0.05fF
C9676 POR2X1_20/B POR2X1_628/O 0.01fF
C9677 POR2X1_411/B PAND2X1_398/CTRL2 0.01fF
C9678 PAND2X1_326/B PAND2X1_169/CTRL 0.01fF
C9679 POR2X1_78/B PAND2X1_93/B 0.58fF
C9680 PAND2X1_244/CTRL2 POR2X1_72/B 0.02fF
C9681 PAND2X1_41/B POR2X1_296/B 0.07fF
C9682 POR2X1_638/Y PAND2X1_53/O 0.15fF
C9683 PAND2X1_216/B POR2X1_173/Y 0.02fF
C9684 POR2X1_24/CTRL POR2X1_14/Y 0.01fF
C9685 POR2X1_814/A POR2X1_220/A 0.02fF
C9686 POR2X1_274/A PAND2X1_516/O 0.04fF
C9687 POR2X1_843/O POR2X1_287/B 0.01fF
C9688 PAND2X1_35/A POR2X1_7/B 0.01fF
C9689 POR2X1_853/A POR2X1_471/A 0.01fF
C9690 POR2X1_48/A POR2X1_256/CTRL 0.01fF
C9691 POR2X1_20/B PAND2X1_6/A 0.45fF
C9692 POR2X1_23/Y PAND2X1_515/CTRL2 0.22fF
C9693 POR2X1_116/A D_INPUT_1 0.03fF
C9694 POR2X1_706/B PAND2X1_20/A 0.01fF
C9695 POR2X1_41/B POR2X1_692/CTRL 0.01fF
C9696 POR2X1_197/CTRL2 POR2X1_555/B 0.01fF
C9697 PAND2X1_236/CTRL2 POR2X1_590/A 0.00fF
C9698 POR2X1_34/B VDD 0.00fF
C9699 POR2X1_620/A VDD 0.00fF
C9700 POR2X1_336/CTRL2 POR2X1_556/A 0.00fF
C9701 POR2X1_664/m4_208_n4# PAND2X1_387/m4_208_n4# 0.13fF
C9702 PAND2X1_65/B POR2X1_448/CTRL 0.01fF
C9703 PAND2X1_450/O POR2X1_257/A 0.01fF
C9704 POR2X1_569/a_16_28# POR2X1_174/A 0.03fF
C9705 POR2X1_814/A POR2X1_569/A 0.10fF
C9706 POR2X1_841/B PAND2X1_369/CTRL 0.02fF
C9707 PAND2X1_65/B PAND2X1_245/a_76_28# 0.02fF
C9708 PAND2X1_248/CTRL POR2X1_294/B 0.01fF
C9709 POR2X1_669/B VDD 5.17fF
C9710 POR2X1_141/O PAND2X1_20/A 0.01fF
C9711 POR2X1_78/B POR2X1_78/A 26.02fF
C9712 POR2X1_400/A POR2X1_590/A 0.03fF
C9713 POR2X1_341/A POR2X1_804/A 0.51fF
C9714 POR2X1_102/Y PAND2X1_719/CTRL2 0.01fF
C9715 POR2X1_750/B POR2X1_543/A 0.03fF
C9716 POR2X1_748/A INPUT_7 0.06fF
C9717 PAND2X1_307/a_76_28# POR2X1_40/Y 0.00fF
C9718 POR2X1_97/CTRL POR2X1_814/A 0.03fF
C9719 POR2X1_709/A PAND2X1_69/A 0.02fF
C9720 PAND2X1_613/a_76_28# PAND2X1_55/Y 0.04fF
C9721 PAND2X1_580/CTRL PAND2X1_578/Y 0.01fF
C9722 PAND2X1_58/A POR2X1_608/CTRL 0.01fF
C9723 POR2X1_290/Y POR2X1_37/Y 0.17fF
C9724 POR2X1_41/B PAND2X1_623/CTRL2 0.02fF
C9725 PAND2X1_679/O POR2X1_750/B 0.01fF
C9726 PAND2X1_714/A PAND2X1_731/B 0.16fF
C9727 POR2X1_490/Y POR2X1_599/A 0.05fF
C9728 POR2X1_192/Y POR2X1_174/A 0.06fF
C9729 PAND2X1_717/A PAND2X1_112/a_16_344# 0.02fF
C9730 POR2X1_119/CTRL POR2X1_37/Y 0.01fF
C9731 POR2X1_302/CTRL2 POR2X1_302/B 0.01fF
C9732 POR2X1_96/A POR2X1_487/a_16_28# 0.03fF
C9733 PAND2X1_250/m4_208_n4# POR2X1_389/Y 0.01fF
C9734 PAND2X1_287/a_16_344# PAND2X1_771/Y 0.04fF
C9735 POR2X1_48/A PAND2X1_506/O 0.05fF
C9736 PAND2X1_206/CTRL2 POR2X1_40/Y 0.03fF
C9737 POR2X1_102/Y POR2X1_498/CTRL 0.00fF
C9738 POR2X1_437/a_76_344# PAND2X1_190/Y 0.04fF
C9739 PAND2X1_39/B POR2X1_249/a_16_28# 0.07fF
C9740 PAND2X1_620/Y POR2X1_627/CTRL2 0.00fF
C9741 POR2X1_150/Y PAND2X1_181/CTRL2 0.01fF
C9742 POR2X1_366/Y POR2X1_97/A 0.50fF
C9743 POR2X1_37/Y PAND2X1_658/B 0.05fF
C9744 POR2X1_842/a_56_344# POR2X1_741/Y 0.00fF
C9745 POR2X1_464/a_56_344# POR2X1_750/B 0.00fF
C9746 PAND2X1_41/B POR2X1_547/B 0.07fF
C9747 PAND2X1_278/CTRL INPUT_0 0.47fF
C9748 PAND2X1_20/A POR2X1_554/Y 0.01fF
C9749 POR2X1_679/B POR2X1_411/B 0.09fF
C9750 POR2X1_332/B POR2X1_750/B 0.05fF
C9751 POR2X1_46/Y PAND2X1_706/CTRL2 0.11fF
C9752 POR2X1_49/Y POR2X1_820/Y 0.68fF
C9753 POR2X1_748/A INPUT_4 0.08fF
C9754 PAND2X1_863/B PAND2X1_733/A 0.03fF
C9755 POR2X1_68/O POR2X1_402/A 0.01fF
C9756 POR2X1_502/A POR2X1_302/B 0.02fF
C9757 POR2X1_475/CTRL2 POR2X1_249/Y 0.01fF
C9758 POR2X1_781/B VDD 0.03fF
C9759 POR2X1_436/CTRL2 POR2X1_802/B 0.01fF
C9760 POR2X1_96/A POR2X1_423/Y 0.03fF
C9761 PAND2X1_6/Y PAND2X1_689/CTRL 0.01fF
C9762 POR2X1_186/Y POR2X1_742/a_16_28# 0.03fF
C9763 POR2X1_541/B POR2X1_260/A 0.04fF
C9764 PAND2X1_137/Y PAND2X1_140/O 0.02fF
C9765 PAND2X1_220/O POR2X1_83/B 0.01fF
C9766 POR2X1_96/A POR2X1_297/a_56_344# 0.00fF
C9767 POR2X1_503/O POR2X1_411/B 0.02fF
C9768 PAND2X1_59/B INPUT_6 0.01fF
C9769 PAND2X1_459/CTRL POR2X1_55/Y 0.01fF
C9770 POR2X1_788/A POR2X1_788/Y 0.01fF
C9771 PAND2X1_362/A PAND2X1_354/CTRL 0.01fF
C9772 POR2X1_147/A PAND2X1_58/A 0.01fF
C9773 POR2X1_523/Y PAND2X1_58/A 0.03fF
C9774 PAND2X1_65/B POR2X1_244/B 0.06fF
C9775 POR2X1_65/A POR2X1_314/CTRL2 0.01fF
C9776 POR2X1_783/a_16_28# POR2X1_783/B -0.00fF
C9777 POR2X1_404/O POR2X1_404/Y 0.05fF
C9778 POR2X1_356/A POR2X1_852/B 0.03fF
C9779 POR2X1_24/CTRL POR2X1_55/Y 0.01fF
C9780 PAND2X1_82/CTRL POR2X1_66/A 0.01fF
C9781 PAND2X1_798/B PAND2X1_78/O 0.06fF
C9782 PAND2X1_48/B POR2X1_654/B 0.03fF
C9783 POR2X1_297/Y VDD 0.00fF
C9784 POR2X1_769/A PAND2X1_32/B 0.01fF
C9785 PAND2X1_793/Y POR2X1_5/Y 0.05fF
C9786 POR2X1_207/B POR2X1_590/A 0.02fF
C9787 POR2X1_52/A POR2X1_376/B 0.16fF
C9788 PAND2X1_9/Y POR2X1_394/A 0.03fF
C9789 POR2X1_458/Y POR2X1_343/CTRL 0.01fF
C9790 PAND2X1_660/CTRL POR2X1_413/A 0.01fF
C9791 PAND2X1_805/Y PAND2X1_854/A 0.52fF
C9792 PAND2X1_58/A PAND2X1_69/A 7.68fF
C9793 POR2X1_718/a_16_28# PAND2X1_57/B 0.03fF
C9794 POR2X1_417/Y PAND2X1_469/B 0.03fF
C9795 POR2X1_516/A POR2X1_23/Y 0.05fF
C9796 POR2X1_404/B VDD 0.19fF
C9797 POR2X1_805/Y POR2X1_758/CTRL 0.01fF
C9798 POR2X1_650/A POR2X1_294/B 0.03fF
C9799 PAND2X1_23/Y POR2X1_287/B 0.15fF
C9800 POR2X1_683/Y POR2X1_72/B 0.01fF
C9801 POR2X1_413/A PAND2X1_660/B 2.20fF
C9802 POR2X1_66/B PAND2X1_63/Y 0.06fF
C9803 POR2X1_673/CTRL2 POR2X1_38/B 0.01fF
C9804 POR2X1_132/O POR2X1_20/B 0.02fF
C9805 POR2X1_376/B POR2X1_152/A 0.03fF
C9806 PAND2X1_474/a_76_28# POR2X1_153/Y 0.05fF
C9807 PAND2X1_751/CTRL VDD 0.00fF
C9808 PAND2X1_479/CTRL2 POR2X1_599/A 0.16fF
C9809 PAND2X1_535/Y POR2X1_102/Y 0.05fF
C9810 POR2X1_116/A POR2X1_362/CTRL2 0.00fF
C9811 POR2X1_296/B POR2X1_228/Y 0.03fF
C9812 POR2X1_333/A POR2X1_577/O 0.03fF
C9813 POR2X1_293/Y POR2X1_372/A 0.03fF
C9814 POR2X1_678/A POR2X1_407/Y 0.00fF
C9815 POR2X1_41/O PAND2X1_852/A 0.01fF
C9816 PAND2X1_55/Y POR2X1_402/a_16_28# 0.02fF
C9817 POR2X1_407/A POR2X1_343/A 0.09fF
C9818 PAND2X1_23/Y POR2X1_483/A 0.03fF
C9819 PAND2X1_76/Y PAND2X1_514/Y 0.03fF
C9820 POR2X1_94/A D_INPUT_1 0.33fF
C9821 D_INPUT_3 POR2X1_14/Y 0.34fF
C9822 PAND2X1_48/B POR2X1_778/O 0.31fF
C9823 PAND2X1_284/a_76_28# POR2X1_279/Y 0.01fF
C9824 PAND2X1_844/Y VDD -0.00fF
C9825 POR2X1_119/Y POR2X1_20/B 0.14fF
C9826 POR2X1_113/Y POR2X1_390/O 0.01fF
C9827 POR2X1_13/A PAND2X1_99/CTRL 0.01fF
C9828 POR2X1_813/Y POR2X1_669/B 0.04fF
C9829 PAND2X1_854/CTRL VDD -0.00fF
C9830 PAND2X1_6/A PAND2X1_381/CTRL2 0.01fF
C9831 PAND2X1_702/O POR2X1_40/Y 0.00fF
C9832 PAND2X1_180/CTRL2 PAND2X1_566/Y 0.00fF
C9833 POR2X1_859/A POR2X1_415/m4_208_n4# 0.05fF
C9834 POR2X1_13/A POR2X1_597/A 0.01fF
C9835 POR2X1_400/A POR2X1_214/B 0.00fF
C9836 POR2X1_590/A POR2X1_566/B 0.03fF
C9837 POR2X1_61/Y POR2X1_208/Y 0.04fF
C9838 PAND2X1_65/B POR2X1_793/A 3.79fF
C9839 POR2X1_66/B POR2X1_113/Y 0.03fF
C9840 PAND2X1_421/a_76_28# PAND2X1_90/Y 0.01fF
C9841 POR2X1_102/Y POR2X1_246/Y 0.01fF
C9842 POR2X1_186/Y POR2X1_341/Y 0.03fF
C9843 POR2X1_330/Y POR2X1_318/A 0.09fF
C9844 POR2X1_221/Y VDD 0.07fF
C9845 PAND2X1_635/O INPUT_7 0.08fF
C9846 POR2X1_402/A POR2X1_402/a_16_28# 0.03fF
C9847 PAND2X1_643/Y POR2X1_595/Y 0.03fF
C9848 POR2X1_48/A POR2X1_394/a_16_28# -0.00fF
C9849 POR2X1_13/A POR2X1_48/Y 0.18fF
C9850 PAND2X1_319/B PAND2X1_211/A 0.07fF
C9851 POR2X1_290/Y POR2X1_293/Y 0.10fF
C9852 POR2X1_572/B POR2X1_572/O 0.02fF
C9853 POR2X1_817/Y POR2X1_820/Y 0.18fF
C9854 PAND2X1_433/O PAND2X1_57/B 0.02fF
C9855 POR2X1_147/A POR2X1_435/Y 0.06fF
C9856 POR2X1_814/A PAND2X1_72/A 0.20fF
C9857 POR2X1_79/Y PAND2X1_730/CTRL2 0.01fF
C9858 POR2X1_38/Y PAND2X1_340/O 0.04fF
C9859 POR2X1_791/A POR2X1_791/Y 0.01fF
C9860 PAND2X1_682/CTRL POR2X1_220/Y 0.10fF
C9861 POR2X1_423/Y POR2X1_7/A 0.15fF
C9862 POR2X1_722/B POR2X1_294/B 0.06fF
C9863 PAND2X1_93/B POR2X1_294/A 0.10fF
C9864 POR2X1_791/A POR2X1_637/B 0.03fF
C9865 PAND2X1_370/O VDD 0.00fF
C9866 POR2X1_23/Y POR2X1_373/CTRL2 0.01fF
C9867 POR2X1_390/O POR2X1_260/A 0.08fF
C9868 PAND2X1_28/CTRL POR2X1_750/B 0.00fF
C9869 PAND2X1_73/Y POR2X1_244/Y 0.03fF
C9870 POR2X1_853/A POR2X1_570/a_16_28# 0.03fF
C9871 POR2X1_198/CTRL2 POR2X1_198/B 0.01fF
C9872 POR2X1_16/A PAND2X1_78/CTRL 0.01fF
C9873 PAND2X1_434/CTRL2 PAND2X1_390/Y 0.01fF
C9874 PAND2X1_124/Y POR2X1_7/Y 0.03fF
C9875 POR2X1_49/Y POR2X1_583/a_16_28# 0.11fF
C9876 POR2X1_78/A PAND2X1_142/CTRL2 0.01fF
C9877 POR2X1_43/B POR2X1_7/B 0.33fF
C9878 POR2X1_66/B POR2X1_260/A 1.30fF
C9879 POR2X1_435/Y PAND2X1_69/A 0.07fF
C9880 POR2X1_41/B POR2X1_255/Y 0.10fF
C9881 POR2X1_113/O PAND2X1_65/B 0.01fF
C9882 POR2X1_511/Y POR2X1_387/Y 0.07fF
C9883 PAND2X1_73/Y PAND2X1_527/CTRL2 0.02fF
C9884 PAND2X1_592/Y PAND2X1_850/O 0.15fF
C9885 POR2X1_43/B POR2X1_277/O 0.08fF
C9886 POR2X1_647/Y POR2X1_101/Y 0.01fF
C9887 PAND2X1_635/O INPUT_4 0.02fF
C9888 POR2X1_532/A POR2X1_215/O 0.02fF
C9889 PAND2X1_94/A PAND2X1_23/O 0.06fF
C9890 INPUT_1 PAND2X1_23/CTRL2 0.00fF
C9891 POR2X1_853/A POR2X1_853/a_16_28# 0.02fF
C9892 POR2X1_96/A PAND2X1_359/a_16_344# 0.02fF
C9893 POR2X1_306/a_16_28# POR2X1_236/Y 0.03fF
C9894 PAND2X1_661/O PAND2X1_653/Y 0.04fF
C9895 POR2X1_347/A PAND2X1_96/CTRL2 0.01fF
C9896 POR2X1_188/A POR2X1_260/A 3.06fF
C9897 POR2X1_143/a_16_28# POR2X1_43/B 0.00fF
C9898 POR2X1_62/Y POR2X1_29/A 0.20fF
C9899 POR2X1_383/A POR2X1_549/B 0.03fF
C9900 POR2X1_596/A POR2X1_220/Y 0.03fF
C9901 POR2X1_659/A POR2X1_632/Y 0.01fF
C9902 POR2X1_480/A POR2X1_799/CTRL2 0.03fF
C9903 POR2X1_72/B POR2X1_39/Y 0.01fF
C9904 PAND2X1_48/B POR2X1_705/CTRL 0.01fF
C9905 PAND2X1_785/CTRL POR2X1_7/B 0.01fF
C9906 POR2X1_502/A POR2X1_578/O 0.11fF
C9907 POR2X1_78/A POR2X1_294/A 0.17fF
C9908 POR2X1_52/A PAND2X1_186/O 0.15fF
C9909 POR2X1_327/Y POR2X1_453/O 0.08fF
C9910 POR2X1_330/Y POR2X1_574/Y 0.05fF
C9911 POR2X1_38/B POR2X1_7/B 0.06fF
C9912 POR2X1_514/Y POR2X1_139/CTRL2 0.00fF
C9913 POR2X1_730/Y POR2X1_828/Y 0.02fF
C9914 PAND2X1_69/A PAND2X1_377/Y 0.01fF
C9915 D_INPUT_3 PAND2X1_472/B 0.10fF
C9916 PAND2X1_825/CTRL VDD 0.00fF
C9917 POR2X1_722/Y PAND2X1_306/CTRL 0.01fF
C9918 POR2X1_713/A PAND2X1_94/A 0.01fF
C9919 PAND2X1_469/B POR2X1_184/Y 0.03fF
C9920 POR2X1_481/Y PAND2X1_555/CTRL 0.01fF
C9921 POR2X1_68/A POR2X1_723/B 0.05fF
C9922 POR2X1_566/A POR2X1_319/Y 0.07fF
C9923 POR2X1_346/B PAND2X1_16/a_76_28# 0.04fF
C9924 POR2X1_236/Y POR2X1_172/CTRL 0.06fF
C9925 PAND2X1_808/Y PAND2X1_773/O 0.02fF
C9926 POR2X1_188/O POR2X1_220/Y 0.02fF
C9927 PAND2X1_661/B POR2X1_48/Y 0.03fF
C9928 POR2X1_49/Y PAND2X1_844/CTRL 0.00fF
C9929 POR2X1_83/B POR2X1_7/Y 0.03fF
C9930 POR2X1_346/CTRL PAND2X1_23/Y 0.00fF
C9931 POR2X1_251/Y PAND2X1_140/A 0.01fF
C9932 POR2X1_49/Y POR2X1_144/CTRL2 0.01fF
C9933 POR2X1_326/A POR2X1_436/CTRL 0.01fF
C9934 PAND2X1_477/B POR2X1_43/B 0.04fF
C9935 POR2X1_8/Y POR2X1_58/CTRL2 0.10fF
C9936 POR2X1_193/A PAND2X1_60/B 8.46fF
C9937 D_INPUT_3 POR2X1_55/Y 0.05fF
C9938 POR2X1_579/Y PAND2X1_60/B 0.07fF
C9939 POR2X1_244/B POR2X1_259/O 0.01fF
C9940 POR2X1_346/CTRL2 POR2X1_68/A 0.01fF
C9941 PAND2X1_852/O POR2X1_821/Y 0.05fF
C9942 POR2X1_294/B PAND2X1_111/B 0.08fF
C9943 POR2X1_675/O POR2X1_188/Y 0.02fF
C9944 POR2X1_255/Y POR2X1_256/Y 0.04fF
C9945 PAND2X1_661/Y POR2X1_829/A 0.34fF
C9946 POR2X1_618/a_16_28# POR2X1_382/Y 0.01fF
C9947 PAND2X1_390/Y PAND2X1_851/CTRL 0.01fF
C9948 POR2X1_537/Y POR2X1_777/B 0.05fF
C9949 POR2X1_810/O POR2X1_809/Y 0.02fF
C9950 POR2X1_572/B PAND2X1_60/B 0.04fF
C9951 POR2X1_315/CTRL2 POR2X1_91/Y 0.01fF
C9952 PAND2X1_56/Y POR2X1_702/CTRL 0.13fF
C9953 POR2X1_360/A POR2X1_360/a_16_28# 0.04fF
C9954 POR2X1_41/B POR2X1_385/O 0.02fF
C9955 POR2X1_302/B POR2X1_188/Y 0.00fF
C9956 POR2X1_859/A POR2X1_260/A 0.07fF
C9957 POR2X1_416/B POR2X1_626/O 0.01fF
C9958 PAND2X1_216/B PAND2X1_735/Y 0.07fF
C9959 D_INPUT_0 POR2X1_522/CTRL 0.07fF
C9960 POR2X1_665/A POR2X1_665/Y 0.15fF
C9961 PAND2X1_96/B PAND2X1_69/A 0.38fF
C9962 POR2X1_537/Y POR2X1_660/A 0.12fF
C9963 POR2X1_57/A PAND2X1_836/CTRL 0.01fF
C9964 PAND2X1_76/Y POR2X1_75/Y 0.10fF
C9965 PAND2X1_865/Y POR2X1_72/B 0.03fF
C9966 PAND2X1_205/A PAND2X1_332/Y 0.10fF
C9967 PAND2X1_388/Y POR2X1_309/Y 0.03fF
C9968 POR2X1_322/Y PAND2X1_565/CTRL 0.00fF
C9969 POR2X1_322/CTRL PAND2X1_569/B 0.03fF
C9970 POR2X1_192/Y POR2X1_704/Y 0.28fF
C9971 PAND2X1_797/Y POR2X1_40/Y 0.03fF
C9972 POR2X1_573/O PAND2X1_48/A 0.05fF
C9973 POR2X1_7/B PAND2X1_336/O 0.17fF
C9974 POR2X1_300/a_56_344# PAND2X1_349/A 0.00fF
C9975 PAND2X1_41/B PAND2X1_759/CTRL2 0.03fF
C9976 POR2X1_449/A POR2X1_220/Y 0.07fF
C9977 INPUT_1 POR2X1_786/A 0.03fF
C9978 POR2X1_503/O POR2X1_52/A 0.01fF
C9979 POR2X1_614/A PAND2X1_60/B 0.22fF
C9980 PAND2X1_631/m4_208_n4# POR2X1_90/Y 0.07fF
C9981 POR2X1_463/O POR2X1_459/Y 0.04fF
C9982 PAND2X1_284/O POR2X1_258/Y 0.03fF
C9983 PAND2X1_20/A POR2X1_39/B 0.03fF
C9984 POR2X1_532/A POR2X1_711/CTRL 0.02fF
C9985 POR2X1_828/CTRL POR2X1_260/A 0.01fF
C9986 POR2X1_166/O POR2X1_73/Y 0.01fF
C9987 PAND2X1_689/CTRL PAND2X1_52/B 0.01fF
C9988 POR2X1_552/CTRL2 VDD 0.00fF
C9989 POR2X1_791/B POR2X1_791/A 0.00fF
C9990 POR2X1_417/CTRL2 POR2X1_387/Y 0.06fF
C9991 POR2X1_41/CTRL POR2X1_42/Y 0.01fF
C9992 PAND2X1_816/O POR2X1_463/Y 0.02fF
C9993 POR2X1_579/Y POR2X1_332/O 0.00fF
C9994 POR2X1_325/CTRL2 POR2X1_542/B 0.03fF
C9995 PAND2X1_534/CTRL2 POR2X1_788/B 0.03fF
C9996 POR2X1_390/B POR2X1_301/CTRL2 0.00fF
C9997 POR2X1_222/A POR2X1_702/A 0.03fF
C9998 POR2X1_368/a_16_28# POR2X1_271/A 0.03fF
C9999 POR2X1_116/Y POR2X1_391/Y 0.01fF
C10000 POR2X1_359/CTRL2 PAND2X1_57/B 0.03fF
C10001 POR2X1_417/O POR2X1_283/A 0.03fF
C10002 POR2X1_567/A POR2X1_653/O 0.03fF
C10003 PAND2X1_658/CTRL POR2X1_77/Y 0.02fF
C10004 PAND2X1_574/CTRL2 POR2X1_73/Y 0.00fF
C10005 POR2X1_203/O PAND2X1_111/B 0.01fF
C10006 POR2X1_795/O POR2X1_186/B 0.01fF
C10007 PAND2X1_353/Y VDD 0.01fF
C10008 PAND2X1_264/CTRL POR2X1_73/Y 0.07fF
C10009 POR2X1_16/A PAND2X1_642/B 0.03fF
C10010 POR2X1_13/A PAND2X1_506/Y 0.06fF
C10011 PAND2X1_422/O PAND2X1_60/B 0.17fF
C10012 PAND2X1_649/A VDD 0.00fF
C10013 POR2X1_9/Y PAND2X1_66/O 0.09fF
C10014 POR2X1_57/A PAND2X1_467/Y 0.03fF
C10015 POR2X1_642/a_16_28# POR2X1_559/A -0.00fF
C10016 POR2X1_405/CTRL PAND2X1_52/B 0.00fF
C10017 POR2X1_81/A VDD 1.25fF
C10018 INPUT_1 POR2X1_248/O 0.02fF
C10019 POR2X1_567/A POR2X1_231/CTRL2 0.13fF
C10020 POR2X1_118/CTRL2 POR2X1_153/Y 0.04fF
C10021 POR2X1_416/B POR2X1_427/Y 0.00fF
C10022 POR2X1_307/A PAND2X1_305/m4_208_n4# 0.02fF
C10023 POR2X1_796/A POR2X1_307/A 0.13fF
C10024 POR2X1_440/Y PAND2X1_60/B 0.03fF
C10025 POR2X1_54/Y POR2X1_462/CTRL 0.01fF
C10026 PAND2X1_59/O POR2X1_260/A 0.02fF
C10027 POR2X1_508/B POR2X1_857/B 0.03fF
C10028 POR2X1_493/CTRL2 POR2X1_773/B 0.00fF
C10029 POR2X1_339/O POR2X1_341/Y 0.00fF
C10030 PAND2X1_833/O POR2X1_39/B 0.01fF
C10031 PAND2X1_824/B PAND2X1_96/B 0.08fF
C10032 POR2X1_614/A POR2X1_370/CTRL2 0.03fF
C10033 POR2X1_42/Y POR2X1_397/CTRL 0.01fF
C10034 POR2X1_566/A PAND2X1_179/O 0.08fF
C10035 POR2X1_567/A POR2X1_294/B 0.05fF
C10036 POR2X1_366/Y POR2X1_567/A 0.07fF
C10037 PAND2X1_852/B POR2X1_394/A 3.68fF
C10038 POR2X1_383/A PAND2X1_298/CTRL2 0.12fF
C10039 POR2X1_248/O POR2X1_153/Y 0.04fF
C10040 POR2X1_327/Y POR2X1_840/B 0.09fF
C10041 POR2X1_513/B PAND2X1_304/a_16_344# 0.01fF
C10042 POR2X1_662/CTRL2 POR2X1_353/A 0.01fF
C10043 POR2X1_41/B POR2X1_85/O 0.00fF
C10044 POR2X1_193/A POR2X1_554/O 0.01fF
C10045 PAND2X1_350/O PAND2X1_341/Y 0.01fF
C10046 PAND2X1_76/Y PAND2X1_332/Y 0.09fF
C10047 POR2X1_840/Y PAND2X1_55/Y 0.01fF
C10048 PAND2X1_543/m4_208_n4# POR2X1_77/Y 0.12fF
C10049 POR2X1_416/B POR2X1_411/CTRL2 0.01fF
C10050 POR2X1_440/Y POR2X1_353/A 0.01fF
C10051 POR2X1_499/A POR2X1_260/B 0.03fF
C10052 PAND2X1_94/A PAND2X1_184/CTRL2 0.01fF
C10053 PAND2X1_470/CTRL POR2X1_119/Y 0.01fF
C10054 POR2X1_3/A POR2X1_762/O 0.22fF
C10055 PAND2X1_175/B PAND2X1_853/B 0.06fF
C10056 POR2X1_116/A PAND2X1_93/B 0.03fF
C10057 POR2X1_355/B PAND2X1_52/B 31.86fF
C10058 PAND2X1_832/CTRL POR2X1_677/Y 0.00fF
C10059 POR2X1_304/CTRL2 POR2X1_90/Y 0.01fF
C10060 POR2X1_472/B POR2X1_862/A 0.09fF
C10061 POR2X1_673/Y POR2X1_721/O 0.14fF
C10062 POR2X1_845/A POR2X1_7/A 0.02fF
C10063 POR2X1_556/A POR2X1_66/A 0.03fF
C10064 POR2X1_730/Y PAND2X1_533/a_16_344# 0.01fF
C10065 POR2X1_234/A VDD 0.39fF
C10066 POR2X1_119/Y PAND2X1_121/CTRL2 0.00fF
C10067 PAND2X1_779/Y POR2X1_39/B 0.01fF
C10068 POR2X1_76/A POR2X1_260/B 0.15fF
C10069 PAND2X1_484/O POR2X1_260/A 0.01fF
C10070 POR2X1_252/Y PAND2X1_549/B 0.03fF
C10071 PAND2X1_640/CTRL POR2X1_77/Y 0.00fF
C10072 POR2X1_456/B POR2X1_180/CTRL 0.00fF
C10073 POR2X1_644/CTRL POR2X1_260/B 0.01fF
C10074 PAND2X1_20/A POR2X1_296/CTRL2 0.01fF
C10075 POR2X1_774/O POR2X1_691/A 0.01fF
C10076 POR2X1_174/B POR2X1_227/A 0.03fF
C10077 PAND2X1_448/a_76_28# POR2X1_20/B 0.02fF
C10078 PAND2X1_731/CTRL POR2X1_77/Y 0.00fF
C10079 POR2X1_620/A PAND2X1_9/Y 0.01fF
C10080 POR2X1_855/Y POR2X1_863/A 0.04fF
C10081 POR2X1_281/Y VDD 0.14fF
C10082 POR2X1_86/Y PAND2X1_6/A 0.03fF
C10083 D_INPUT_5 PAND2X1_3/A 1.52fF
C10084 POR2X1_116/A POR2X1_78/A 0.03fF
C10085 POR2X1_456/B PAND2X1_48/A 0.03fF
C10086 PAND2X1_821/a_16_344# PAND2X1_52/B 0.01fF
C10087 POR2X1_39/B PAND2X1_509/CTRL 0.18fF
C10088 POR2X1_814/B POR2X1_646/a_16_28# 0.01fF
C10089 POR2X1_669/B PAND2X1_9/Y 0.03fF
C10090 PAND2X1_404/CTRL2 POR2X1_411/B 0.01fF
C10091 POR2X1_87/CTRL2 POR2X1_38/B 0.01fF
C10092 POR2X1_376/B POR2X1_441/O 0.02fF
C10093 POR2X1_209/A POR2X1_711/Y 0.03fF
C10094 POR2X1_286/B POR2X1_78/A 0.03fF
C10095 PAND2X1_826/CTRL2 POR2X1_296/B 0.02fF
C10096 PAND2X1_404/Y D_INPUT_0 0.07fF
C10097 POR2X1_837/B PAND2X1_57/B 0.04fF
C10098 PAND2X1_1/CTRL2 D_INPUT_4 0.01fF
C10099 PAND2X1_31/CTRL PAND2X1_3/A 0.00fF
C10100 POR2X1_99/A POR2X1_99/O 0.02fF
C10101 POR2X1_257/A POR2X1_83/B 1.92fF
C10102 POR2X1_597/a_16_28# POR2X1_761/A 0.02fF
C10103 POR2X1_199/B POR2X1_260/A 0.06fF
C10104 POR2X1_66/B POR2X1_610/Y 0.20fF
C10105 POR2X1_139/A POR2X1_138/A 0.02fF
C10106 PAND2X1_287/Y PAND2X1_577/Y 0.02fF
C10107 POR2X1_313/O POR2X1_167/Y 0.01fF
C10108 POR2X1_866/A PAND2X1_73/Y 0.05fF
C10109 POR2X1_831/O POR2X1_330/Y 0.02fF
C10110 INPUT_3 POR2X1_94/A 0.12fF
C10111 PAND2X1_20/A POR2X1_34/CTRL2 0.01fF
C10112 POR2X1_66/B POR2X1_473/O 0.02fF
C10113 POR2X1_493/O PAND2X1_72/A 0.01fF
C10114 POR2X1_110/Y POR2X1_110/CTRL 0.01fF
C10115 POR2X1_306/Y PAND2X1_796/B 0.70fF
C10116 POR2X1_49/Y PAND2X1_217/O 0.01fF
C10117 POR2X1_306/Y PAND2X1_454/B 0.06fF
C10118 PAND2X1_717/A POR2X1_46/Y 0.03fF
C10119 PAND2X1_254/Y POR2X1_329/A 0.03fF
C10120 PAND2X1_717/A PAND2X1_151/a_76_28# 0.02fF
C10121 POR2X1_263/CTRL POR2X1_236/Y 0.15fF
C10122 PAND2X1_436/a_76_28# PAND2X1_435/Y 0.03fF
C10123 PAND2X1_659/Y PAND2X1_737/CTRL2 0.03fF
C10124 POR2X1_606/a_16_28# POR2X1_121/B 0.03fF
C10125 POR2X1_814/B POR2X1_621/A 0.07fF
C10126 POR2X1_590/A POR2X1_458/m4_208_n4# 0.08fF
C10127 POR2X1_61/A POR2X1_447/B 0.02fF
C10128 POR2X1_705/B INPUT_0 0.05fF
C10129 PAND2X1_267/Y POR2X1_40/Y 0.03fF
C10130 POR2X1_416/B PAND2X1_507/CTRL2 0.01fF
C10131 POR2X1_49/Y PAND2X1_443/O 0.01fF
C10132 PAND2X1_39/B POR2X1_403/m4_208_n4# 0.01fF
C10133 PAND2X1_694/CTRL PAND2X1_425/Y 0.01fF
C10134 POR2X1_292/CTRL POR2X1_90/Y 0.10fF
C10135 POR2X1_864/A POR2X1_783/A 0.08fF
C10136 POR2X1_663/B VDD 0.51fF
C10137 POR2X1_736/A POR2X1_186/B 0.07fF
C10138 PAND2X1_652/O POR2X1_385/Y 0.04fF
C10139 POR2X1_329/A POR2X1_599/A 0.05fF
C10140 POR2X1_602/m4_208_n4# POR2X1_330/Y 0.06fF
C10141 POR2X1_319/A PAND2X1_65/B 0.06fF
C10142 PAND2X1_58/A POR2X1_720/O 0.01fF
C10143 POR2X1_567/A POR2X1_542/O 0.01fF
C10144 PAND2X1_5/CTRL2 POR2X1_612/A 0.00fF
C10145 POR2X1_43/B PAND2X1_206/B 0.07fF
C10146 POR2X1_814/A POR2X1_793/A 0.05fF
C10147 POR2X1_141/Y D_INPUT_0 0.04fF
C10148 POR2X1_634/a_16_28# POR2X1_66/A 0.00fF
C10149 POR2X1_119/Y POR2X1_518/a_76_344# 0.02fF
C10150 GATE_479 POR2X1_23/Y 0.03fF
C10151 PAND2X1_826/O VDD 0.00fF
C10152 POR2X1_614/Y POR2X1_69/A 0.02fF
C10153 POR2X1_453/CTRL POR2X1_590/A 0.31fF
C10154 POR2X1_98/CTRL2 PAND2X1_41/B 0.01fF
C10155 POR2X1_834/O POR2X1_330/Y 0.08fF
C10156 PAND2X1_404/Y PAND2X1_84/a_16_344# 0.01fF
C10157 PAND2X1_72/A POR2X1_151/Y 0.04fF
C10158 POR2X1_78/B POR2X1_84/A 0.01fF
C10159 POR2X1_23/Y POR2X1_485/O 0.02fF
C10160 POR2X1_846/Y POR2X1_793/A 0.01fF
C10161 POR2X1_78/A POR2X1_94/A 0.05fF
C10162 POR2X1_106/a_16_28# POR2X1_251/A 0.01fF
C10163 D_INPUT_3 POR2X1_612/A 0.01fF
C10164 PAND2X1_48/B PAND2X1_416/CTRL2 0.00fF
C10165 POR2X1_850/A POR2X1_656/CTRL 0.01fF
C10166 POR2X1_20/B PAND2X1_334/CTRL 0.01fF
C10167 PAND2X1_48/B PAND2X1_268/CTRL 0.01fF
C10168 POR2X1_268/CTRL POR2X1_5/Y 0.01fF
C10169 POR2X1_856/B POR2X1_552/Y 0.02fF
C10170 POR2X1_49/Y POR2X1_83/B 0.20fF
C10171 POR2X1_112/a_16_28# POR2X1_632/Y 0.01fF
C10172 PAND2X1_703/O POR2X1_167/Y 0.02fF
C10173 PAND2X1_459/m4_208_n4# PAND2X1_58/A 0.15fF
C10174 PAND2X1_865/Y PAND2X1_440/O 0.00fF
C10175 POR2X1_864/O POR2X1_750/B 0.01fF
C10176 POR2X1_518/O POR2X1_77/Y 0.01fF
C10177 POR2X1_294/Y VDD 0.16fF
C10178 PAND2X1_770/a_16_344# PAND2X1_771/Y 0.04fF
C10179 POR2X1_105/O PAND2X1_41/B 0.01fF
C10180 POR2X1_634/A POR2X1_734/A 0.10fF
C10181 PAND2X1_638/B POR2X1_585/O 0.00fF
C10182 POR2X1_776/A POR2X1_35/Y 0.12fF
C10183 POR2X1_57/A PAND2X1_837/O 0.01fF
C10184 POR2X1_48/A PAND2X1_818/O 0.01fF
C10185 POR2X1_119/Y POR2X1_43/Y 0.05fF
C10186 PAND2X1_20/A POR2X1_402/CTRL 0.00fF
C10187 POR2X1_818/Y PAND2X1_751/CTRL 0.01fF
C10188 POR2X1_689/O POR2X1_32/A 0.01fF
C10189 PAND2X1_214/CTRL PAND2X1_35/Y 0.01fF
C10190 POR2X1_260/B PAND2X1_132/O 0.01fF
C10191 POR2X1_692/O POR2X1_46/Y 0.01fF
C10192 PAND2X1_57/CTRL2 POR2X1_590/A 0.00fF
C10193 POR2X1_114/B POR2X1_475/a_76_344# 0.00fF
C10194 PAND2X1_860/A PAND2X1_508/Y 0.03fF
C10195 POR2X1_556/A POR2X1_532/A 0.03fF
C10196 POR2X1_262/Y PAND2X1_844/B 0.06fF
C10197 POR2X1_186/Y PAND2X1_41/B 0.19fF
C10198 PAND2X1_798/B POR2X1_437/CTRL 0.04fF
C10199 PAND2X1_406/m4_208_n4# POR2X1_784/A 0.08fF
C10200 POR2X1_52/A POR2X1_484/CTRL2 0.00fF
C10201 POR2X1_13/A POR2X1_423/CTRL2 0.00fF
C10202 POR2X1_676/CTRL POR2X1_828/A 0.01fF
C10203 POR2X1_676/CTRL2 PAND2X1_69/A 0.01fF
C10204 PAND2X1_577/B PAND2X1_577/O -0.00fF
C10205 D_INPUT_0 POR2X1_404/Y 0.03fF
C10206 POR2X1_538/CTRL2 POR2X1_270/Y 0.08fF
C10207 PAND2X1_57/B POR2X1_792/O 0.07fF
C10208 POR2X1_548/B POR2X1_66/A 0.01fF
C10209 POR2X1_66/A PAND2X1_385/CTRL 0.01fF
C10210 POR2X1_400/CTRL POR2X1_206/A 0.10fF
C10211 POR2X1_825/Y POR2X1_397/O 0.00fF
C10212 PAND2X1_766/O PAND2X1_90/Y 0.20fF
C10213 POR2X1_477/A POR2X1_466/A 0.33fF
C10214 POR2X1_660/CTRL POR2X1_307/Y 0.03fF
C10215 D_GATE_865 POR2X1_750/B 0.01fF
C10216 POR2X1_754/Y POR2X1_615/Y 0.03fF
C10217 POR2X1_305/a_56_344# POR2X1_416/B 0.00fF
C10218 POR2X1_360/A POR2X1_296/B 0.01fF
C10219 PAND2X1_68/O POR2X1_42/Y 0.07fF
C10220 PAND2X1_48/B PAND2X1_282/O 0.01fF
C10221 POR2X1_333/A POR2X1_566/A 0.10fF
C10222 POR2X1_48/A PAND2X1_35/O 0.05fF
C10223 POR2X1_123/CTRL2 POR2X1_78/A 0.01fF
C10224 POR2X1_294/Y POR2X1_741/Y 0.05fF
C10225 PAND2X1_35/B VDD 0.02fF
C10226 POR2X1_644/CTRL POR2X1_407/Y 0.01fF
C10227 POR2X1_856/B POR2X1_35/Y 0.03fF
C10228 POR2X1_56/CTRL POR2X1_55/Y 0.01fF
C10229 POR2X1_330/Y PAND2X1_131/O 0.03fF
C10230 PAND2X1_570/O PAND2X1_771/Y 0.02fF
C10231 POR2X1_440/Y POR2X1_477/CTRL 0.01fF
C10232 POR2X1_458/CTRL PAND2X1_32/B 0.01fF
C10233 POR2X1_355/B POR2X1_467/Y 0.01fF
C10234 POR2X1_846/Y POR2X1_753/CTRL2 0.01fF
C10235 POR2X1_661/Y POR2X1_740/Y 0.33fF
C10236 POR2X1_102/Y POR2X1_275/O 0.01fF
C10237 PAND2X1_449/CTRL2 PAND2X1_308/Y 0.01fF
C10238 POR2X1_130/A POR2X1_734/A 0.10fF
C10239 POR2X1_283/CTRL2 PAND2X1_365/B 0.01fF
C10240 PAND2X1_97/CTRL2 POR2X1_91/Y 0.01fF
C10241 PAND2X1_217/CTRL2 PAND2X1_124/Y 0.03fF
C10242 POR2X1_854/O POR2X1_854/B 0.02fF
C10243 POR2X1_706/B VDD 0.01fF
C10244 POR2X1_490/Y PAND2X1_572/O 0.01fF
C10245 POR2X1_40/Y POR2X1_531/CTRL 0.01fF
C10246 POR2X1_447/A POR2X1_510/Y 0.01fF
C10247 POR2X1_389/A PAND2X1_93/B 0.02fF
C10248 POR2X1_263/Y POR2X1_73/Y 0.00fF
C10249 PAND2X1_267/CTRL2 POR2X1_7/A 0.01fF
C10250 POR2X1_537/Y POR2X1_814/A 0.05fF
C10251 POR2X1_141/O VDD 0.00fF
C10252 POR2X1_624/Y POR2X1_101/Y 0.05fF
C10253 PAND2X1_72/A PAND2X1_135/CTRL2 0.00fF
C10254 POR2X1_643/A POR2X1_294/B 0.25fF
C10255 PAND2X1_652/A PAND2X1_361/CTRL 0.11fF
C10256 POR2X1_657/a_76_344# POR2X1_741/Y 0.00fF
C10257 PAND2X1_769/CTRL VDD -0.00fF
C10258 POR2X1_750/B POR2X1_579/Y 0.05fF
C10259 POR2X1_60/A PAND2X1_658/B 0.92fF
C10260 PAND2X1_862/B POR2X1_376/B 0.03fF
C10261 PAND2X1_65/B POR2X1_483/B 0.02fF
C10262 PAND2X1_499/Y VDD 1.56fF
C10263 POR2X1_23/Y POR2X1_142/Y 0.04fF
C10264 POR2X1_72/B POR2X1_494/Y 0.08fF
C10265 POR2X1_83/B PAND2X1_565/CTRL 0.00fF
C10266 POR2X1_260/B POR2X1_537/A 0.01fF
C10267 POR2X1_13/A PAND2X1_76/Y 0.06fF
C10268 PAND2X1_94/A POR2X1_243/B 0.01fF
C10269 PAND2X1_480/B PAND2X1_276/CTRL 0.27fF
C10270 PAND2X1_48/B POR2X1_777/B 0.10fF
C10271 PAND2X1_416/CTRL POR2X1_260/A 0.06fF
C10272 POR2X1_220/Y PAND2X1_90/Y 0.07fF
C10273 POR2X1_23/Y PAND2X1_175/B 0.03fF
C10274 POR2X1_800/A POR2X1_783/O 0.00fF
C10275 POR2X1_431/Y POR2X1_129/Y 0.01fF
C10276 PAND2X1_630/O POR2X1_748/A 0.10fF
C10277 POR2X1_179/CTRL POR2X1_40/Y 0.01fF
C10278 POR2X1_78/Y POR2X1_557/B 0.18fF
C10279 POR2X1_806/CTRL2 PAND2X1_69/A 0.01fF
C10280 PAND2X1_284/Y PAND2X1_577/Y 8.31fF
C10281 POR2X1_840/B POR2X1_858/a_16_28# 0.08fF
C10282 PAND2X1_116/O PAND2X1_553/B 0.06fF
C10283 POR2X1_639/Y POR2X1_769/A 0.03fF
C10284 POR2X1_96/A PAND2X1_687/Y 0.06fF
C10285 PAND2X1_673/m4_208_n4# POR2X1_236/Y 0.09fF
C10286 POR2X1_420/Y POR2X1_90/Y 0.01fF
C10287 PAND2X1_76/Y PAND2X1_775/O 0.05fF
C10288 POR2X1_807/A POR2X1_294/B 0.02fF
C10289 POR2X1_43/B POR2X1_750/B 4.15fF
C10290 POR2X1_346/CTRL2 PAND2X1_58/A 0.00fF
C10291 POR2X1_66/A PAND2X1_393/O 0.01fF
C10292 INPUT_2 POR2X1_104/O 0.01fF
C10293 POR2X1_278/a_16_28# PAND2X1_734/B 0.05fF
C10294 POR2X1_104/a_56_344# D_INPUT_1 0.00fF
C10295 POR2X1_287/B POR2X1_733/A 0.05fF
C10296 POR2X1_614/A POR2X1_254/A 0.01fF
C10297 INPUT_1 POR2X1_28/CTRL2 0.00fF
C10298 POR2X1_253/CTRL2 PAND2X1_508/Y 0.00fF
C10299 POR2X1_389/A POR2X1_78/A 0.03fF
C10300 PAND2X1_48/B PAND2X1_65/B 0.32fF
C10301 PAND2X1_420/O PAND2X1_96/B 0.01fF
C10302 PAND2X1_88/CTRL2 POR2X1_38/B 0.01fF
C10303 PAND2X1_798/B PAND2X1_579/O 0.03fF
C10304 PAND2X1_468/CTRL PAND2X1_580/B 0.00fF
C10305 POR2X1_278/Y POR2X1_498/CTRL 0.08fF
C10306 PAND2X1_413/O POR2X1_713/B 0.29fF
C10307 PAND2X1_454/a_16_344# POR2X1_376/B 0.02fF
C10308 POR2X1_590/A PAND2X1_60/B 2.68fF
C10309 PAND2X1_244/B POR2X1_263/Y 0.03fF
C10310 PAND2X1_23/Y POR2X1_663/CTRL 0.01fF
C10311 POR2X1_614/A POR2X1_750/B 0.41fF
C10312 POR2X1_411/B PAND2X1_716/B 0.03fF
C10313 POR2X1_54/Y POR2X1_774/A 0.01fF
C10314 POR2X1_848/Y POR2X1_559/A 0.06fF
C10315 POR2X1_859/A POR2X1_790/CTRL2 0.02fF
C10316 PAND2X1_480/B PAND2X1_804/B 0.05fF
C10317 POR2X1_273/CTRL POR2X1_129/Y 0.12fF
C10318 PAND2X1_863/B POR2X1_13/A 0.02fF
C10319 PAND2X1_643/O POR2X1_595/Y 0.02fF
C10320 POR2X1_554/Y VDD 0.22fF
C10321 POR2X1_99/A PAND2X1_69/A 0.03fF
C10322 POR2X1_657/CTRL POR2X1_510/Y 0.00fF
C10323 POR2X1_68/A POR2X1_828/Y 0.05fF
C10324 POR2X1_141/a_16_28# POR2X1_139/Y -0.00fF
C10325 POR2X1_422/Y POR2X1_7/A 0.03fF
C10326 POR2X1_13/A POR2X1_669/CTRL 0.01fF
C10327 PAND2X1_562/B PAND2X1_566/Y 0.18fF
C10328 POR2X1_239/O POR2X1_40/Y 0.00fF
C10329 POR2X1_640/Y PAND2X1_96/B 0.03fF
C10330 PAND2X1_493/a_76_28# POR2X1_411/B 0.02fF
C10331 PAND2X1_254/Y PAND2X1_515/CTRL 0.01fF
C10332 PAND2X1_801/B PAND2X1_794/B 0.00fF
C10333 POR2X1_38/B POR2X1_750/B 0.07fF
C10334 POR2X1_557/A D_INPUT_0 0.03fF
C10335 POR2X1_114/B POR2X1_830/A 0.08fF
C10336 POR2X1_49/Y POR2X1_522/Y 0.12fF
C10337 POR2X1_41/B POR2X1_46/Y 0.13fF
C10338 POR2X1_37/Y PAND2X1_100/a_16_344# 0.01fF
C10339 POR2X1_124/B POR2X1_287/B 0.01fF
C10340 POR2X1_780/CTRL POR2X1_780/A 0.01fF
C10341 POR2X1_832/a_56_344# PAND2X1_55/Y 0.00fF
C10342 POR2X1_83/B PAND2X1_720/O 0.15fF
C10343 POR2X1_717/CTRL2 POR2X1_814/B 0.01fF
C10344 POR2X1_428/CTRL POR2X1_32/A 0.01fF
C10345 POR2X1_83/B PAND2X1_559/CTRL 0.01fF
C10346 POR2X1_465/B POR2X1_553/Y 0.01fF
C10347 POR2X1_81/O PAND2X1_510/B 0.01fF
C10348 POR2X1_334/Y PAND2X1_93/B 0.07fF
C10349 POR2X1_45/Y INPUT_0 0.03fF
C10350 POR2X1_270/Y POR2X1_186/B 0.03fF
C10351 D_INPUT_0 POR2X1_571/CTRL 0.01fF
C10352 PAND2X1_857/A PAND2X1_200/O 0.02fF
C10353 INPUT_1 POR2X1_225/CTRL 0.01fF
C10354 PAND2X1_731/A PAND2X1_731/B 0.04fF
C10355 POR2X1_300/O POR2X1_13/A 0.02fF
C10356 POR2X1_41/B PAND2X1_623/Y 0.03fF
C10357 POR2X1_66/B POR2X1_725/Y 0.07fF
C10358 PAND2X1_581/O PAND2X1_3/B 0.01fF
C10359 POR2X1_823/a_56_344# POR2X1_236/Y 0.00fF
C10360 INPUT_1 POR2X1_586/Y 0.01fF
C10361 PAND2X1_557/A POR2X1_283/A 0.51fF
C10362 D_INPUT_0 PAND2X1_514/a_76_28# 0.01fF
C10363 PAND2X1_449/CTRL2 POR2X1_77/Y 0.01fF
C10364 PAND2X1_422/O POR2X1_750/B 0.09fF
C10365 POR2X1_717/CTRL POR2X1_475/A 0.07fF
C10366 POR2X1_192/Y POR2X1_795/B 0.05fF
C10367 POR2X1_335/a_16_28# POR2X1_740/Y 0.06fF
C10368 POR2X1_383/A PAND2X1_766/CTRL 0.01fF
C10369 POR2X1_84/A POR2X1_294/A 0.03fF
C10370 POR2X1_590/A POR2X1_353/A 0.03fF
C10371 POR2X1_445/CTRL POR2X1_222/Y 0.00fF
C10372 POR2X1_96/A PAND2X1_798/B 0.29fF
C10373 PAND2X1_263/m4_208_n4# D_INPUT_1 0.01fF
C10374 GATE_741 PAND2X1_362/CTRL2 0.01fF
C10375 POR2X1_628/CTRL POR2X1_55/Y 0.01fF
C10376 POR2X1_565/B POR2X1_294/B 0.00fF
C10377 POR2X1_188/A POR2X1_725/Y 0.10fF
C10378 POR2X1_13/A PAND2X1_566/Y 0.05fF
C10379 POR2X1_66/A POR2X1_721/m4_208_n4# 0.09fF
C10380 POR2X1_41/B PAND2X1_840/A 0.04fF
C10381 POR2X1_87/B PAND2X1_32/CTRL2 0.00fF
C10382 PAND2X1_694/CTRL POR2X1_614/A 0.01fF
C10383 PAND2X1_236/O POR2X1_68/B 0.02fF
C10384 PAND2X1_94/A PAND2X1_616/O 0.02fF
C10385 PAND2X1_65/B POR2X1_577/a_76_344# 0.01fF
C10386 PAND2X1_810/A PAND2X1_810/O 0.03fF
C10387 POR2X1_666/O POR2X1_394/A 0.01fF
C10388 PAND2X1_472/a_16_344# POR2X1_83/B 0.02fF
C10389 POR2X1_400/A POR2X1_532/A 0.01fF
C10390 POR2X1_96/A POR2X1_759/Y 0.01fF
C10391 PAND2X1_473/O VDD 0.00fF
C10392 POR2X1_691/O POR2X1_783/B 0.03fF
C10393 POR2X1_814/B POR2X1_181/B 0.03fF
C10394 POR2X1_683/Y POR2X1_7/B 0.00fF
C10395 POR2X1_594/Y PAND2X1_652/A 0.02fF
C10396 POR2X1_57/A PAND2X1_556/B 0.03fF
C10397 POR2X1_334/Y POR2X1_78/A 0.09fF
C10398 POR2X1_546/A POR2X1_705/a_16_28# 0.05fF
C10399 PAND2X1_322/CTRL2 PAND2X1_32/B 0.01fF
C10400 PAND2X1_65/B PAND2X1_534/O 0.04fF
C10401 PAND2X1_72/CTRL2 POR2X1_579/Y 0.00fF
C10402 POR2X1_57/A PAND2X1_549/CTRL 0.01fF
C10403 POR2X1_722/B POR2X1_407/A 0.03fF
C10404 POR2X1_72/B POR2X1_172/a_76_344# 0.00fF
C10405 POR2X1_57/A POR2X1_822/a_16_28# 0.03fF
C10406 POR2X1_54/CTRL2 PAND2X1_58/A 0.01fF
C10407 PAND2X1_731/CTRL2 POR2X1_763/Y 0.03fF
C10408 PAND2X1_863/B PAND2X1_643/Y 0.11fF
C10409 PAND2X1_96/B POR2X1_121/Y 0.07fF
C10410 PAND2X1_23/Y POR2X1_469/a_16_28# 0.01fF
C10411 POR2X1_407/A POR2X1_294/B 0.10fF
C10412 POR2X1_364/A POR2X1_785/a_16_28# 0.01fF
C10413 POR2X1_48/A POR2X1_524/CTRL2 0.03fF
C10414 PAND2X1_228/CTRL2 POR2X1_52/Y 0.00fF
C10415 PAND2X1_736/A PAND2X1_357/Y 0.01fF
C10416 PAND2X1_715/O POR2X1_387/Y 0.09fF
C10417 POR2X1_22/A POR2X1_587/Y 0.03fF
C10418 PAND2X1_824/B POR2X1_99/A 0.02fF
C10419 PAND2X1_403/O POR2X1_399/Y -0.00fF
C10420 PAND2X1_421/CTRL2 POR2X1_596/A 0.01fF
C10421 POR2X1_358/CTRL PAND2X1_32/B 0.10fF
C10422 PAND2X1_658/A PAND2X1_6/A 0.00fF
C10423 POR2X1_777/Y VDD 0.09fF
C10424 PAND2X1_215/B POR2X1_73/Y 0.04fF
C10425 POR2X1_60/A PAND2X1_337/a_76_28# 0.05fF
C10426 POR2X1_700/CTRL POR2X1_700/Y 0.00fF
C10427 POR2X1_700/O POR2X1_90/Y 0.00fF
C10428 POR2X1_285/Y POR2X1_294/A 0.03fF
C10429 POR2X1_355/B POR2X1_350/B 0.03fF
C10430 POR2X1_483/O POR2X1_228/Y 0.02fF
C10431 POR2X1_593/CTRL POR2X1_750/B 0.00fF
C10432 PAND2X1_48/B POR2X1_541/CTRL 0.03fF
C10433 POR2X1_548/B POR2X1_532/A 0.06fF
C10434 PAND2X1_530/O PAND2X1_69/A 0.03fF
C10435 POR2X1_423/Y POR2X1_153/Y 0.11fF
C10436 PAND2X1_592/CTRL2 POR2X1_283/A 0.03fF
C10437 POR2X1_383/A POR2X1_192/Y 0.05fF
C10438 POR2X1_176/Y POR2X1_236/Y 0.00fF
C10439 POR2X1_614/A PAND2X1_72/CTRL2 0.03fF
C10440 POR2X1_271/Y PAND2X1_716/B 0.03fF
C10441 POR2X1_350/Y POR2X1_351/Y 0.01fF
C10442 PAND2X1_839/a_76_28# PAND2X1_835/Y 0.04fF
C10443 POR2X1_335/A POR2X1_840/B 0.05fF
C10444 POR2X1_38/Y POR2X1_57/Y 0.01fF
C10445 POR2X1_315/Y POR2X1_13/A 0.68fF
C10446 D_INPUT_1 POR2X1_218/A 0.07fF
C10447 POR2X1_293/Y POR2X1_387/Y 0.16fF
C10448 PAND2X1_6/Y POR2X1_513/Y 0.06fF
C10449 PAND2X1_738/Y PAND2X1_336/CTRL 0.14fF
C10450 PAND2X1_793/Y PAND2X1_489/CTRL2 0.01fF
C10451 PAND2X1_465/B POR2X1_7/A 0.01fF
C10452 PAND2X1_6/A POR2X1_73/Y 0.10fF
C10453 PAND2X1_691/Y POR2X1_96/A 0.03fF
C10454 POR2X1_504/Y PAND2X1_507/a_76_28# 0.04fF
C10455 POR2X1_177/CTRL2 POR2X1_236/Y 0.01fF
C10456 PAND2X1_63/Y PAND2X1_81/O 0.08fF
C10457 POR2X1_351/Y POR2X1_341/Y 0.22fF
C10458 POR2X1_680/Y PAND2X1_728/CTRL2 0.00fF
C10459 PAND2X1_631/A POR2X1_748/A 0.01fF
C10460 POR2X1_276/O POR2X1_366/A 0.01fF
C10461 POR2X1_327/Y POR2X1_217/CTRL 0.01fF
C10462 POR2X1_293/Y PAND2X1_121/O 0.06fF
C10463 POR2X1_853/A POR2X1_577/a_16_28# 0.05fF
C10464 POR2X1_78/O PAND2X1_79/Y 0.00fF
C10465 PAND2X1_389/Y POR2X1_184/Y 0.03fF
C10466 PAND2X1_55/Y POR2X1_537/A 0.02fF
C10467 PAND2X1_4/CTRL2 D_INPUT_1 0.02fF
C10468 PAND2X1_403/CTRL POR2X1_411/B 0.01fF
C10469 POR2X1_786/Y PAND2X1_150/O 0.09fF
C10470 POR2X1_495/Y POR2X1_283/A 0.02fF
C10471 POR2X1_709/B PAND2X1_90/Y 0.29fF
C10472 PAND2X1_6/Y POR2X1_205/A 0.07fF
C10473 POR2X1_346/CTRL2 PAND2X1_96/B 0.03fF
C10474 POR2X1_860/A POR2X1_362/CTRL 0.00fF
C10475 POR2X1_574/Y PAND2X1_516/CTRL2 0.01fF
C10476 POR2X1_46/Y PAND2X1_308/Y 0.03fF
C10477 PAND2X1_65/B PAND2X1_527/a_16_344# 0.01fF
C10478 PAND2X1_353/a_16_344# POR2X1_152/A 0.02fF
C10479 POR2X1_519/O POR2X1_42/Y 0.01fF
C10480 POR2X1_859/A POR2X1_559/A 0.01fF
C10481 PAND2X1_447/CTRL2 POR2X1_329/A 0.02fF
C10482 PAND2X1_264/O POR2X1_42/Y 0.09fF
C10483 POR2X1_68/B PAND2X1_153/O 0.02fF
C10484 POR2X1_669/B POR2X1_747/O 0.01fF
C10485 POR2X1_5/CTRL2 VDD -0.00fF
C10486 POR2X1_123/Y POR2X1_137/Y 0.02fF
C10487 POR2X1_774/Y POR2X1_691/A 0.01fF
C10488 PAND2X1_6/Y POR2X1_366/A 0.03fF
C10489 POR2X1_790/A PAND2X1_382/a_16_344# 0.02fF
C10490 PAND2X1_148/CTRL PAND2X1_209/A 0.01fF
C10491 PAND2X1_284/a_16_344# POR2X1_280/Y 0.02fF
C10492 POR2X1_110/CTRL INPUT_0 0.05fF
C10493 PAND2X1_80/a_16_344# PAND2X1_71/Y 0.01fF
C10494 POR2X1_190/Y POR2X1_191/B 0.08fF
C10495 PAND2X1_244/B PAND2X1_6/A 0.07fF
C10496 PAND2X1_6/O PAND2X1_55/Y 0.01fF
C10497 PAND2X1_65/B PAND2X1_517/CTRL 0.01fF
C10498 PAND2X1_305/a_16_344# PAND2X1_32/B 0.01fF
C10499 POR2X1_57/A POR2X1_165/O 0.02fF
C10500 POR2X1_137/Y POR2X1_216/CTRL 0.00fF
C10501 PAND2X1_57/B PAND2X1_48/A 0.12fF
C10502 POR2X1_327/Y PAND2X1_421/CTRL 0.01fF
C10503 PAND2X1_217/B POR2X1_39/B 0.05fF
C10504 POR2X1_276/A POR2X1_532/A 0.02fF
C10505 PAND2X1_297/CTRL2 POR2X1_68/B 0.01fF
C10506 POR2X1_532/A POR2X1_566/B 0.25fF
C10507 POR2X1_158/Y PAND2X1_725/Y 0.18fF
C10508 POR2X1_562/O POR2X1_186/B 0.01fF
C10509 PAND2X1_651/O POR2X1_43/B 0.05fF
C10510 POR2X1_840/B POR2X1_249/Y 0.05fF
C10511 POR2X1_52/A PAND2X1_716/B 0.03fF
C10512 POR2X1_416/B PAND2X1_540/O 0.04fF
C10513 PAND2X1_572/CTRL PAND2X1_723/A 0.01fF
C10514 POR2X1_72/B PAND2X1_327/a_16_344# 0.01fF
C10515 POR2X1_289/CTRL POR2X1_394/A 0.08fF
C10516 PAND2X1_311/CTRL2 POR2X1_260/A 0.00fF
C10517 POR2X1_43/B PAND2X1_560/B 0.03fF
C10518 PAND2X1_476/A POR2X1_230/Y 0.00fF
C10519 POR2X1_771/a_16_28# POR2X1_769/Y 0.02fF
C10520 POR2X1_356/A POR2X1_508/A 0.02fF
C10521 POR2X1_579/B POR2X1_501/O 0.00fF
C10522 POR2X1_814/A POR2X1_220/CTRL 0.01fF
C10523 POR2X1_68/B POR2X1_772/O 0.02fF
C10524 POR2X1_65/Y PAND2X1_201/CTRL2 0.09fF
C10525 PAND2X1_79/CTRL2 POR2X1_571/Y 0.01fF
C10526 PAND2X1_865/Y POR2X1_7/B 0.07fF
C10527 PAND2X1_550/B PAND2X1_549/B 1.17fF
C10528 VDD POR2X1_39/B 6.21fF
C10529 POR2X1_96/A POR2X1_184/O 0.08fF
C10530 POR2X1_333/O POR2X1_566/B 0.03fF
C10531 POR2X1_447/B D_GATE_222 0.07fF
C10532 POR2X1_780/B POR2X1_260/A 0.60fF
C10533 POR2X1_567/A PAND2X1_504/CTRL 0.21fF
C10534 POR2X1_567/B PAND2X1_52/CTRL 0.09fF
C10535 PAND2X1_661/Y POR2X1_16/A 0.07fF
C10536 POR2X1_614/A POR2X1_156/CTRL2 0.00fF
C10537 PAND2X1_213/Y POR2X1_394/A 0.05fF
C10538 POR2X1_356/A POR2X1_568/B 0.10fF
C10539 POR2X1_67/Y D_INPUT_0 0.03fF
C10540 POR2X1_12/A POR2X1_20/B 0.01fF
C10541 POR2X1_57/A PAND2X1_779/CTRL 0.01fF
C10542 POR2X1_46/Y POR2X1_77/Y 0.05fF
C10543 POR2X1_103/CTRL2 PAND2X1_349/A 0.01fF
C10544 PAND2X1_610/O D_INPUT_2 0.04fF
C10545 POR2X1_68/B POR2X1_113/B 0.06fF
C10546 POR2X1_574/A POR2X1_574/Y 0.23fF
C10547 POR2X1_119/Y POR2X1_73/Y 0.20fF
C10548 POR2X1_188/CTRL POR2X1_737/A 0.01fF
C10549 POR2X1_490/Y POR2X1_411/B 0.03fF
C10550 POR2X1_486/O POR2X1_590/A 0.00fF
C10551 POR2X1_14/Y PAND2X1_87/O 0.01fF
C10552 PAND2X1_23/Y POR2X1_343/Y 0.02fF
C10553 POR2X1_651/Y PAND2X1_90/Y 0.07fF
C10554 POR2X1_101/Y POR2X1_186/B 0.05fF
C10555 POR2X1_415/A PAND2X1_66/CTRL 0.01fF
C10556 POR2X1_788/CTRL2 PAND2X1_60/B 0.00fF
C10557 POR2X1_407/A POR2X1_779/CTRL2 0.00fF
C10558 POR2X1_231/B PAND2X1_72/A 0.01fF
C10559 PAND2X1_655/Y PAND2X1_691/CTRL 0.01fF
C10560 POR2X1_431/Y POR2X1_37/Y 0.01fF
C10561 POR2X1_847/O POR2X1_67/A 0.01fF
C10562 POR2X1_93/CTRL POR2X1_39/B 0.28fF
C10563 POR2X1_250/Y PAND2X1_742/O 0.11fF
C10564 POR2X1_20/B POR2X1_268/O 0.01fF
C10565 POR2X1_39/B PAND2X1_32/B 0.03fF
C10566 POR2X1_730/Y POR2X1_652/A 0.03fF
C10567 PAND2X1_742/B POR2X1_331/O 0.01fF
C10568 POR2X1_190/O POR2X1_568/B 0.16fF
C10569 PAND2X1_659/Y POR2X1_7/CTRL 0.00fF
C10570 POR2X1_220/A POR2X1_568/B 0.05fF
C10571 POR2X1_542/B POR2X1_736/A 0.05fF
C10572 PAND2X1_118/O PAND2X1_72/A 0.02fF
C10573 POR2X1_362/Y POR2X1_116/A 0.00fF
C10574 PAND2X1_484/O POR2X1_559/A 0.13fF
C10575 PAND2X1_802/CTRL PAND2X1_539/Y 0.01fF
C10576 PAND2X1_39/B POR2X1_646/Y 0.03fF
C10577 POR2X1_863/O POR2X1_863/A 0.08fF
C10578 POR2X1_736/A POR2X1_736/O 0.03fF
C10579 PAND2X1_30/a_16_344# INPUT_4 0.01fF
C10580 POR2X1_311/Y PAND2X1_222/CTRL2 0.00fF
C10581 PAND2X1_91/CTRL POR2X1_97/A 0.00fF
C10582 POR2X1_485/Y POR2X1_40/Y 0.03fF
C10583 POR2X1_327/Y POR2X1_737/A 0.11fF
C10584 POR2X1_168/a_16_28# POR2X1_566/B 0.02fF
C10585 POR2X1_834/CTRL2 POR2X1_260/B 0.01fF
C10586 PAND2X1_613/CTRL2 POR2X1_296/B 0.01fF
C10587 POR2X1_827/O VDD 0.00fF
C10588 POR2X1_569/A POR2X1_568/B 0.18fF
C10589 POR2X1_220/A POR2X1_161/CTRL2 0.03fF
C10590 POR2X1_23/Y POR2X1_409/B 0.57fF
C10591 PAND2X1_79/Y POR2X1_500/O 0.00fF
C10592 POR2X1_646/A PAND2X1_90/Y 0.05fF
C10593 PAND2X1_63/CTRL2 POR2X1_66/A 0.03fF
C10594 PAND2X1_659/Y PAND2X1_557/O 0.01fF
C10595 POR2X1_865/B PAND2X1_72/A 0.04fF
C10596 POR2X1_68/B POR2X1_768/A 0.03fF
C10597 POR2X1_499/A POR2X1_860/A 0.03fF
C10598 POR2X1_257/A PAND2X1_444/Y 0.06fF
C10599 PAND2X1_497/CTRL2 POR2X1_590/A 0.04fF
C10600 POR2X1_654/B POR2X1_649/O 0.03fF
C10601 PAND2X1_85/CTRL POR2X1_243/Y -0.01fF
C10602 POR2X1_846/Y POR2X1_615/a_76_344# 0.00fF
C10603 POR2X1_648/Y PAND2X1_511/CTRL 0.02fF
C10604 POR2X1_65/A PAND2X1_838/CTRL2 0.03fF
C10605 POR2X1_568/B POR2X1_570/Y 0.10fF
C10606 POR2X1_411/B PAND2X1_205/Y 0.06fF
C10607 POR2X1_623/CTRL2 POR2X1_296/B 0.01fF
C10608 POR2X1_301/A POR2X1_121/B 0.01fF
C10609 POR2X1_722/A PAND2X1_696/CTRL 0.04fF
C10610 POR2X1_150/Y PAND2X1_558/CTRL 0.01fF
C10611 POR2X1_23/Y PAND2X1_794/CTRL 0.01fF
C10612 POR2X1_48/A POR2X1_819/O 0.01fF
C10613 PAND2X1_206/B PAND2X1_350/A 0.00fF
C10614 POR2X1_717/a_16_28# POR2X1_717/B 0.03fF
C10615 POR2X1_458/Y POR2X1_740/Y 0.10fF
C10616 POR2X1_202/A POR2X1_202/CTRL 0.05fF
C10617 PAND2X1_373/CTRL2 PAND2X1_72/A 0.00fF
C10618 POR2X1_373/Y POR2X1_373/a_16_28# 0.02fF
C10619 POR2X1_228/Y POR2X1_556/CTRL 0.03fF
C10620 POR2X1_479/B POR2X1_479/O 0.01fF
C10621 PAND2X1_48/B POR2X1_814/A 1.13fF
C10622 POR2X1_56/O POR2X1_496/Y 0.07fF
C10623 POR2X1_431/CTRL POR2X1_55/Y 0.01fF
C10624 PAND2X1_242/Y POR2X1_387/Y 0.07fF
C10625 D_INPUT_5 PAND2X1_65/B 0.03fF
C10626 POR2X1_646/Y POR2X1_805/Y 0.03fF
C10627 POR2X1_478/a_16_28# PAND2X1_41/B 0.03fF
C10628 POR2X1_13/A PAND2X1_98/CTRL2 0.01fF
C10629 POR2X1_416/B POR2X1_394/A 0.34fF
C10630 PAND2X1_862/B PAND2X1_203/CTRL2 0.01fF
C10631 POR2X1_461/Y PAND2X1_57/B 0.03fF
C10632 POR2X1_621/A VDD 0.00fF
C10633 PAND2X1_477/CTRL PAND2X1_803/A 0.00fF
C10634 PAND2X1_58/A PAND2X1_37/O 0.01fF
C10635 POR2X1_72/CTRL POR2X1_23/Y 0.01fF
C10636 PAND2X1_45/O POR2X1_740/Y 0.04fF
C10637 PAND2X1_45/CTRL2 POR2X1_741/Y 0.10fF
C10638 PAND2X1_33/CTRL POR2X1_7/B 0.01fF
C10639 PAND2X1_860/A POR2X1_283/A 1.50fF
C10640 POR2X1_98/A POR2X1_68/B 0.09fF
C10641 PAND2X1_88/CTRL2 POR2X1_590/A 0.00fF
C10642 POR2X1_9/Y POR2X1_382/Y 0.05fF
C10643 POR2X1_333/A POR2X1_241/B 0.02fF
C10644 POR2X1_853/A POR2X1_465/CTRL 0.01fF
C10645 PAND2X1_243/B POR2X1_411/B 0.03fF
C10646 PAND2X1_613/O VDD 0.00fF
C10647 POR2X1_23/Y POR2X1_29/CTRL2 0.00fF
C10648 POR2X1_590/A POR2X1_750/B 0.11fF
C10649 POR2X1_462/B POR2X1_462/CTRL 0.01fF
C10650 POR2X1_807/CTRL2 POR2X1_480/A 0.03fF
C10651 POR2X1_23/Y POR2X1_272/Y 0.03fF
C10652 PAND2X1_9/CTRL2 POR2X1_94/A 0.00fF
C10653 PAND2X1_825/O PAND2X1_94/Y 0.00fF
C10654 PAND2X1_205/CTRL PAND2X1_735/Y 0.10fF
C10655 PAND2X1_404/Y PAND2X1_735/Y 0.01fF
C10656 POR2X1_349/Y PAND2X1_93/B 0.00fF
C10657 POR2X1_150/Y PAND2X1_190/Y 0.26fF
C10658 POR2X1_566/A POR2X1_454/m4_208_n4# 0.06fF
C10659 PAND2X1_594/CTRL PAND2X1_90/Y 0.09fF
C10660 PAND2X1_73/Y PAND2X1_42/O 0.07fF
C10661 POR2X1_847/B POR2X1_29/A 0.01fF
C10662 POR2X1_257/A POR2X1_697/Y 0.01fF
C10663 PAND2X1_722/CTRL POR2X1_666/A 0.01fF
C10664 POR2X1_48/A VDD 5.65fF
C10665 PAND2X1_474/CTRL POR2X1_43/B 0.01fF
C10666 POR2X1_623/O VDD 0.00fF
C10667 PAND2X1_603/O PAND2X1_90/Y 0.08fF
C10668 POR2X1_20/B PAND2X1_794/B 0.03fF
C10669 INPUT_2 PAND2X1_618/CTRL 0.00fF
C10670 PAND2X1_23/Y POR2X1_624/Y 0.90fF
C10671 POR2X1_366/Y PAND2X1_271/O 0.03fF
C10672 POR2X1_260/B POR2X1_410/a_16_28# 0.03fF
C10673 POR2X1_440/B PAND2X1_60/B 0.01fF
C10674 POR2X1_78/A POR2X1_475/A 0.01fF
C10675 POR2X1_517/O POR2X1_83/B 0.18fF
C10676 POR2X1_52/A POR2X1_490/Y 0.02fF
C10677 POR2X1_66/B POR2X1_254/O 0.01fF
C10678 POR2X1_126/CTRL2 D_INPUT_2 0.01fF
C10679 POR2X1_422/CTRL2 POR2X1_293/Y 0.01fF
C10680 POR2X1_683/Y POR2X1_604/CTRL 0.00fF
C10681 POR2X1_49/Y PAND2X1_444/Y 0.02fF
C10682 PAND2X1_781/CTRL POR2X1_745/Y 0.00fF
C10683 POR2X1_416/B PAND2X1_198/CTRL2 0.04fF
C10684 POR2X1_696/CTRL POR2X1_376/B 0.01fF
C10685 POR2X1_102/Y PAND2X1_756/CTRL 0.01fF
C10686 POR2X1_283/Y PAND2X1_805/A 0.03fF
C10687 POR2X1_43/B PAND2X1_436/CTRL2 0.00fF
C10688 POR2X1_603/Y POR2X1_236/Y 0.07fF
C10689 POR2X1_97/A POR2X1_853/CTRL2 0.01fF
C10690 POR2X1_115/O POR2X1_218/Y 0.03fF
C10691 POR2X1_57/A POR2X1_441/Y 0.03fF
C10692 POR2X1_10/a_76_344# POR2X1_9/Y 0.02fF
C10693 PAND2X1_39/B POR2X1_804/A 0.03fF
C10694 PAND2X1_531/O POR2X1_547/B 0.00fF
C10695 POR2X1_748/A POR2X1_763/A 0.02fF
C10696 POR2X1_796/Y PAND2X1_599/O 0.04fF
C10697 PAND2X1_655/B POR2X1_411/B 0.00fF
C10698 PAND2X1_360/CTRL2 PAND2X1_347/Y 0.01fF
C10699 PAND2X1_94/CTRL PAND2X1_55/Y 0.01fF
C10700 POR2X1_52/A PAND2X1_448/O 0.03fF
C10701 POR2X1_668/O POR2X1_750/B 0.00fF
C10702 PAND2X1_220/Y PAND2X1_540/a_16_344# 0.04fF
C10703 POR2X1_496/Y POR2X1_627/Y 0.05fF
C10704 PAND2X1_766/m4_208_n4# PAND2X1_41/B 0.09fF
C10705 POR2X1_568/B PAND2X1_72/A 0.11fF
C10706 PAND2X1_255/CTRL POR2X1_186/B 0.01fF
C10707 POR2X1_49/Y PAND2X1_783/Y 0.01fF
C10708 PAND2X1_413/a_76_28# PAND2X1_57/B 0.01fF
C10709 POR2X1_174/B POR2X1_502/A 0.10fF
C10710 POR2X1_220/CTRL2 POR2X1_210/Y 0.01fF
C10711 POR2X1_674/CTRL PAND2X1_652/A 0.14fF
C10712 PAND2X1_573/O PAND2X1_573/B 0.02fF
C10713 PAND2X1_556/B PAND2X1_556/a_16_344# 0.05fF
C10714 POR2X1_440/B POR2X1_353/A 0.37fF
C10715 POR2X1_637/B POR2X1_637/A 0.00fF
C10716 POR2X1_814/A POR2X1_210/B 0.04fF
C10717 PAND2X1_95/B PAND2X1_752/CTRL2 0.01fF
C10718 POR2X1_368/Y PAND2X1_776/Y 0.13fF
C10719 PAND2X1_78/O POR2X1_79/A 0.01fF
C10720 POR2X1_260/B PAND2X1_69/A 0.45fF
C10721 POR2X1_689/A POR2X1_32/A 0.01fF
C10722 POR2X1_32/A PAND2X1_375/O -0.00fF
C10723 PAND2X1_512/O VDD 0.00fF
C10724 POR2X1_648/a_16_28# POR2X1_532/A 0.03fF
C10725 PAND2X1_140/A POR2X1_257/A 0.03fF
C10726 POR2X1_23/Y POR2X1_229/CTRL2 0.01fF
C10727 PAND2X1_139/O PAND2X1_140/Y 0.01fF
C10728 PAND2X1_458/a_16_344# PAND2X1_716/B 0.02fF
C10729 PAND2X1_294/O POR2X1_387/Y 0.09fF
C10730 POR2X1_114/B D_INPUT_0 0.03fF
C10731 PAND2X1_863/CTRL2 VDD 0.00fF
C10732 PAND2X1_39/B PAND2X1_27/CTRL 0.07fF
C10733 POR2X1_596/A POR2X1_644/O 0.01fF
C10734 PAND2X1_7/Y VDD 0.01fF
C10735 PAND2X1_275/CTRL POR2X1_296/B 0.01fF
C10736 POR2X1_83/B PAND2X1_790/Y 0.03fF
C10737 POR2X1_609/Y POR2X1_234/CTRL2 0.00fF
C10738 POR2X1_341/A POR2X1_569/A 0.07fF
C10739 PAND2X1_738/Y PAND2X1_540/O 0.04fF
C10740 PAND2X1_782/CTRL POR2X1_747/Y 0.00fF
C10741 POR2X1_259/A POR2X1_244/B 0.01fF
C10742 PAND2X1_93/B POR2X1_140/CTRL 0.09fF
C10743 POR2X1_556/A POR2X1_787/O 0.03fF
C10744 POR2X1_693/Y POR2X1_32/A 0.05fF
C10745 PAND2X1_542/O PAND2X1_552/B 0.16fF
C10746 PAND2X1_513/O VDD 0.00fF
C10747 PAND2X1_793/Y PAND2X1_354/A 0.03fF
C10748 PAND2X1_467/B PAND2X1_707/Y 0.01fF
C10749 POR2X1_683/O POR2X1_72/B 0.01fF
C10750 PAND2X1_73/Y POR2X1_455/A 0.01fF
C10751 POR2X1_753/Y PAND2X1_6/A 0.07fF
C10752 POR2X1_45/Y POR2X1_102/Y 0.08fF
C10753 PAND2X1_199/A VDD 0.11fF
C10754 PAND2X1_73/Y PAND2X1_519/O 0.12fF
C10755 POR2X1_162/B POR2X1_356/Y 0.35fF
C10756 PAND2X1_854/a_16_344# POR2X1_102/Y 0.01fF
C10757 POR2X1_78/A POR2X1_218/A 0.00fF
C10758 POR2X1_311/Y PAND2X1_798/B 0.07fF
C10759 POR2X1_45/m4_208_n4# POR2X1_272/m4_208_n4# 0.13fF
C10760 POR2X1_855/B POR2X1_808/O 0.01fF
C10761 POR2X1_54/Y POR2X1_750/Y 0.05fF
C10762 POR2X1_834/CTRL2 POR2X1_407/Y 0.01fF
C10763 POR2X1_102/Y POR2X1_234/CTRL 0.01fF
C10764 POR2X1_708/O PAND2X1_90/Y 0.07fF
C10765 PAND2X1_58/A POR2X1_391/Y 0.02fF
C10766 POR2X1_52/A PAND2X1_205/Y 0.03fF
C10767 POR2X1_296/B POR2X1_112/Y 0.03fF
C10768 POR2X1_525/O POR2X1_41/B 0.02fF
C10769 POR2X1_777/B POR2X1_717/Y 0.03fF
C10770 PAND2X1_844/CTRL POR2X1_20/B 0.01fF
C10771 POR2X1_65/A PAND2X1_364/B 0.03fF
C10772 D_INPUT_3 POR2X1_37/Y 0.30fF
C10773 POR2X1_631/a_16_28# POR2X1_294/B 0.01fF
C10774 PAND2X1_217/B PAND2X1_197/Y 0.00fF
C10775 POR2X1_13/A PAND2X1_596/O 0.17fF
C10776 PAND2X1_34/O POR2X1_38/Y 0.05fF
C10777 POR2X1_66/A PAND2X1_60/B 11.81fF
C10778 PAND2X1_804/B PAND2X1_473/B 0.07fF
C10779 PAND2X1_129/O POR2X1_502/A 0.04fF
C10780 POR2X1_41/B PAND2X1_787/Y 0.14fF
C10781 POR2X1_130/A PAND2X1_755/CTRL2 0.12fF
C10782 PAND2X1_653/Y POR2X1_83/B 0.20fF
C10783 PAND2X1_20/A POR2X1_804/A 0.03fF
C10784 POR2X1_5/Y POR2X1_372/Y 0.01fF
C10785 POR2X1_834/Y PAND2X1_601/O 0.02fF
C10786 POR2X1_260/B PAND2X1_765/a_76_28# 0.02fF
C10787 PAND2X1_12/O POR2X1_260/A 0.08fF
C10788 INPUT_0 POR2X1_572/CTRL 0.07fF
C10789 PAND2X1_213/Y POR2X1_669/B 0.07fF
C10790 POR2X1_740/a_16_28# POR2X1_738/Y -0.00fF
C10791 PAND2X1_625/CTRL POR2X1_852/B 0.03fF
C10792 PAND2X1_404/A POR2X1_233/O 0.00fF
C10793 PAND2X1_13/CTRL POR2X1_795/B 0.03fF
C10794 POR2X1_502/A POR2X1_544/A 0.01fF
C10795 GATE_479 POR2X1_238/Y 0.00fF
C10796 POR2X1_13/A PAND2X1_480/B 0.05fF
C10797 PAND2X1_483/CTRL POR2X1_23/Y 0.03fF
C10798 PAND2X1_105/CTRL PAND2X1_562/B 0.06fF
C10799 PAND2X1_752/Y POR2X1_750/B 0.02fF
C10800 POR2X1_351/Y PAND2X1_41/B 0.03fF
C10801 PAND2X1_401/CTRL2 POR2X1_236/Y 0.01fF
C10802 POR2X1_423/CTRL POR2X1_7/A 0.03fF
C10803 PAND2X1_583/O POR2X1_750/B 0.02fF
C10804 POR2X1_407/A POR2X1_807/A 0.03fF
C10805 POR2X1_673/Y POR2X1_623/O 0.09fF
C10806 PAND2X1_137/Y PAND2X1_768/O 0.02fF
C10807 POR2X1_57/A POR2X1_825/O 0.02fF
C10808 POR2X1_60/A POR2X1_387/Y 2.48fF
C10809 POR2X1_416/Y POR2X1_5/Y 0.03fF
C10810 POR2X1_494/CTRL POR2X1_5/Y 0.02fF
C10811 POR2X1_662/Y VDD 0.23fF
C10812 PAND2X1_319/a_56_28# PAND2X1_317/Y 0.00fF
C10813 POR2X1_814/B POR2X1_804/A 0.05fF
C10814 POR2X1_413/A VDD 0.04fF
C10815 PAND2X1_197/Y VDD 0.08fF
C10816 POR2X1_102/CTRL2 POR2X1_411/B 0.01fF
C10817 PAND2X1_151/O POR2X1_55/Y 0.01fF
C10818 POR2X1_848/CTRL2 PAND2X1_52/B 0.10fF
C10819 PAND2X1_635/O POR2X1_763/A 0.03fF
C10820 PAND2X1_486/CTRL2 POR2X1_763/Y 0.03fF
C10821 D_INPUT_3 POR2X1_37/a_16_28# 0.03fF
C10822 POR2X1_66/A POR2X1_546/O 0.02fF
C10823 POR2X1_471/O POR2X1_732/B 0.15fF
C10824 POR2X1_97/A PAND2X1_503/O 0.05fF
C10825 PAND2X1_205/Y PAND2X1_186/O 0.05fF
C10826 PAND2X1_84/Y POR2X1_599/A 0.03fF
C10827 PAND2X1_275/O VDD 0.00fF
C10828 POR2X1_433/Y POR2X1_236/Y 0.11fF
C10829 POR2X1_29/Y POR2X1_5/Y 5.33fF
C10830 PAND2X1_261/a_16_344# POR2X1_260/Y 0.01fF
C10831 PAND2X1_23/Y POR2X1_738/Y 0.01fF
C10832 POR2X1_573/O POR2X1_576/Y 0.01fF
C10833 PAND2X1_56/Y POR2X1_308/a_16_28# 0.08fF
C10834 POR2X1_515/CTRL PAND2X1_6/Y 0.00fF
C10835 INPUT_1 PAND2X1_73/Y 0.00fF
C10836 INPUT_1 POR2X1_422/Y 0.01fF
C10837 POR2X1_78/B POR2X1_538/a_76_344# 0.00fF
C10838 POR2X1_658/CTRL POR2X1_632/Y 0.01fF
C10839 POR2X1_447/B POR2X1_202/A 0.12fF
C10840 POR2X1_804/A POR2X1_325/A 0.03fF
C10841 POR2X1_536/O POR2X1_102/Y 0.04fF
C10842 PAND2X1_6/CTRL2 PAND2X1_20/A 0.01fF
C10843 PAND2X1_23/Y POR2X1_276/CTRL2 0.03fF
C10844 PAND2X1_219/A PAND2X1_737/B 0.08fF
C10845 PAND2X1_318/a_76_28# POR2X1_96/A 0.01fF
C10846 POR2X1_834/Y PAND2X1_58/A 0.05fF
C10847 POR2X1_48/A PAND2X1_703/CTRL 0.01fF
C10848 POR2X1_199/CTRL POR2X1_741/Y 0.01fF
C10849 POR2X1_547/a_16_28# POR2X1_547/B 0.08fF
C10850 PAND2X1_824/O PAND2X1_41/B 0.01fF
C10851 POR2X1_500/A POR2X1_569/A 0.05fF
C10852 POR2X1_730/Y PAND2X1_829/a_16_344# 0.02fF
C10853 POR2X1_632/A PAND2X1_88/Y 0.00fF
C10854 PAND2X1_803/A POR2X1_91/Y 1.88fF
C10855 PAND2X1_48/B POR2X1_260/Y 0.06fF
C10856 POR2X1_532/A POR2X1_794/CTRL2 0.01fF
C10857 PAND2X1_23/Y POR2X1_785/A 0.03fF
C10858 POR2X1_502/A POR2X1_775/CTRL 0.03fF
C10859 POR2X1_186/Y POR2X1_727/CTRL 0.30fF
C10860 POR2X1_49/Y POR2X1_528/Y 0.15fF
C10861 POR2X1_302/a_16_28# PAND2X1_6/Y 0.02fF
C10862 PAND2X1_9/Y POR2X1_39/B 0.03fF
C10863 PAND2X1_23/Y PAND2X1_816/O 0.05fF
C10864 POR2X1_637/B PAND2X1_757/O 0.00fF
C10865 POR2X1_718/O POR2X1_832/A 0.11fF
C10866 POR2X1_43/B PAND2X1_466/CTRL2 0.03fF
C10867 POR2X1_502/A POR2X1_705/O 0.01fF
C10868 POR2X1_46/Y POR2X1_52/Y 0.03fF
C10869 PAND2X1_553/B PAND2X1_357/Y 0.15fF
C10870 PAND2X1_58/A POR2X1_753/O 0.02fF
C10871 POR2X1_662/Y POR2X1_741/Y 0.03fF
C10872 POR2X1_693/CTRL2 POR2X1_73/Y 0.01fF
C10873 POR2X1_334/B POR2X1_264/Y 0.05fF
C10874 POR2X1_691/CTRL2 POR2X1_800/A 0.00fF
C10875 POR2X1_25/a_76_344# D_INPUT_6 0.00fF
C10876 POR2X1_83/B PAND2X1_337/CTRL 0.01fF
C10877 POR2X1_78/A POR2X1_557/B 0.14fF
C10878 POR2X1_529/a_56_344# POR2X1_55/Y 0.03fF
C10879 POR2X1_244/B PAND2X1_88/Y 0.00fF
C10880 PAND2X1_55/Y PAND2X1_178/m4_208_n4# 0.15fF
C10881 POR2X1_376/B PAND2X1_374/O 0.15fF
C10882 POR2X1_65/A PAND2X1_849/B 0.03fF
C10883 PAND2X1_23/Y PAND2X1_504/O 0.03fF
C10884 POR2X1_548/O POR2X1_383/A 0.01fF
C10885 PAND2X1_347/Y PAND2X1_843/Y 0.00fF
C10886 POR2X1_256/a_16_28# POR2X1_255/Y 0.03fF
C10887 POR2X1_76/Y POR2X1_724/A 0.01fF
C10888 PAND2X1_6/Y POR2X1_832/B 0.11fF
C10889 POR2X1_43/B PAND2X1_478/O 0.01fF
C10890 POR2X1_566/A POR2X1_854/CTRL2 0.01fF
C10891 PAND2X1_293/O PAND2X1_60/B 0.02fF
C10892 POR2X1_376/B POR2X1_376/CTRL2 0.03fF
C10893 POR2X1_147/A POR2X1_788/Y 0.21fF
C10894 PAND2X1_69/A PAND2X1_369/O 0.01fF
C10895 POR2X1_307/B POR2X1_590/a_76_344# 0.01fF
C10896 PAND2X1_281/O POR2X1_285/Y 0.02fF
C10897 PAND2X1_408/m4_208_n4# PAND2X1_52/B 0.06fF
C10898 POR2X1_669/B POR2X1_701/a_56_344# 0.00fF
C10899 POR2X1_341/A PAND2X1_72/A 0.13fF
C10900 PAND2X1_55/Y PAND2X1_69/A 0.33fF
C10901 PAND2X1_467/Y POR2X1_236/Y 0.03fF
C10902 POR2X1_181/B VDD 0.01fF
C10903 POR2X1_504/a_56_344# POR2X1_750/B 0.01fF
C10904 POR2X1_43/B PAND2X1_734/CTRL2 0.30fF
C10905 POR2X1_327/Y POR2X1_302/B 0.97fF
C10906 PAND2X1_248/O POR2X1_342/B 0.00fF
C10907 POR2X1_655/A POR2X1_725/CTRL2 0.04fF
C10908 POR2X1_316/Y PAND2X1_436/a_76_28# 0.01fF
C10909 PAND2X1_76/m4_208_n4# PAND2X1_301/m4_208_n4# 0.05fF
C10910 POR2X1_578/Y POR2X1_578/O 0.01fF
C10911 POR2X1_818/Y POR2X1_39/B 0.03fF
C10912 PAND2X1_41/B PAND2X1_184/m4_208_n4# 0.09fF
C10913 POR2X1_41/B POR2X1_248/Y 0.03fF
C10914 POR2X1_177/O POR2X1_72/B 0.02fF
C10915 D_INPUT_3 POR2X1_293/Y 0.04fF
C10916 POR2X1_262/CTRL2 POR2X1_7/A 0.01fF
C10917 POR2X1_193/A POR2X1_318/A 0.07fF
C10918 POR2X1_23/O POR2X1_4/Y 0.09fF
C10919 PAND2X1_553/O POR2X1_55/Y 0.02fF
C10920 POR2X1_792/B PAND2X1_60/B 0.10fF
C10921 POR2X1_800/A POR2X1_644/A 0.03fF
C10922 POR2X1_477/A POR2X1_209/A 0.13fF
C10923 POR2X1_802/B PAND2X1_60/B 0.07fF
C10924 POR2X1_36/B POR2X1_425/a_16_28# 0.03fF
C10925 POR2X1_743/CTRL2 POR2X1_153/Y 0.01fF
C10926 PAND2X1_650/A VDD -0.00fF
C10927 POR2X1_788/A POR2X1_788/CTRL 0.01fF
C10928 POR2X1_740/Y POR2X1_724/A 2.58fF
C10929 D_INPUT_0 POR2X1_513/A 0.02fF
C10930 POR2X1_228/CTRL PAND2X1_7/Y 0.01fF
C10931 POR2X1_402/A PAND2X1_69/A 0.01fF
C10932 PAND2X1_215/B PAND2X1_656/A 0.07fF
C10933 POR2X1_334/CTRL INPUT_0 0.03fF
C10934 PAND2X1_96/B POR2X1_391/Y 0.42fF
C10935 POR2X1_237/Y POR2X1_73/Y 0.03fF
C10936 POR2X1_304/CTRL2 POR2X1_102/Y 0.01fF
C10937 POR2X1_334/Y PAND2X1_65/Y 0.03fF
C10938 POR2X1_383/A PAND2X1_71/O 0.01fF
C10939 POR2X1_773/A POR2X1_734/A 0.13fF
C10940 PAND2X1_562/O PAND2X1_555/Y 0.03fF
C10941 POR2X1_834/Y POR2X1_435/Y 0.05fF
C10942 PAND2X1_352/A POR2X1_77/Y 0.03fF
C10943 POR2X1_52/CTRL POR2X1_102/Y 0.01fF
C10944 POR2X1_222/Y PAND2X1_60/B 0.03fF
C10945 PAND2X1_649/A PAND2X1_403/B 0.04fF
C10946 POR2X1_116/Y POR2X1_392/CTRL2 0.03fF
C10947 POR2X1_96/A PAND2X1_472/CTRL 0.01fF
C10948 PAND2X1_812/CTRL PAND2X1_811/Y 0.01fF
C10949 POR2X1_858/A POR2X1_858/a_16_28# 0.07fF
C10950 POR2X1_358/O POR2X1_566/B 0.03fF
C10951 POR2X1_41/B PAND2X1_114/O 0.01fF
C10952 POR2X1_407/Y PAND2X1_69/A 0.03fF
C10953 POR2X1_325/O PAND2X1_55/Y 0.02fF
C10954 POR2X1_857/B POR2X1_502/CTRL2 0.04fF
C10955 PAND2X1_48/B POR2X1_472/a_16_28# 0.02fF
C10956 POR2X1_99/B POR2X1_186/Y 0.01fF
C10957 POR2X1_319/O POR2X1_568/Y 0.04fF
C10958 POR2X1_306/O POR2X1_90/Y 0.01fF
C10959 POR2X1_96/Y POR2X1_60/Y 0.00fF
C10960 POR2X1_416/B POR2X1_669/B 0.53fF
C10961 POR2X1_52/A POR2X1_260/A 0.04fF
C10962 PAND2X1_738/Y POR2X1_394/A 0.10fF
C10963 POR2X1_133/CTRL POR2X1_384/A 0.01fF
C10964 POR2X1_419/CTRL POR2X1_42/Y 0.01fF
C10965 POR2X1_514/Y POR2X1_141/A 0.00fF
C10966 PAND2X1_865/Y PAND2X1_220/Y 0.10fF
C10967 POR2X1_291/CTRL POR2X1_42/Y 0.01fF
C10968 PAND2X1_653/CTRL PAND2X1_557/A 0.01fF
C10969 POR2X1_51/B POR2X1_587/O 0.01fF
C10970 POR2X1_255/Y PAND2X1_349/A 0.01fF
C10971 PAND2X1_384/O POR2X1_546/A 0.01fF
C10972 PAND2X1_138/O POR2X1_135/Y 0.00fF
C10973 POR2X1_62/Y VDD 1.14fF
C10974 POR2X1_8/Y POR2X1_618/O 0.17fF
C10975 POR2X1_16/A POR2X1_591/CTRL 0.00fF
C10976 POR2X1_93/a_16_28# POR2X1_93/A 0.05fF
C10977 D_INPUT_1 POR2X1_361/a_16_28# 0.02fF
C10978 POR2X1_41/B POR2X1_144/CTRL 0.04fF
C10979 POR2X1_829/A PAND2X1_200/B 0.00fF
C10980 POR2X1_532/A PAND2X1_60/B 0.36fF
C10981 POR2X1_67/Y POR2X1_816/O 0.10fF
C10982 POR2X1_390/B POR2X1_68/A 0.03fF
C10983 PAND2X1_824/B PAND2X1_55/Y 0.07fF
C10984 POR2X1_274/B POR2X1_702/A 0.00fF
C10985 PAND2X1_816/a_76_28# POR2X1_260/A 0.01fF
C10986 D_INPUT_2 POR2X1_4/CTRL2 0.01fF
C10987 POR2X1_732/B POR2X1_703/Y 0.01fF
C10988 POR2X1_337/A PAND2X1_69/A 0.40fF
C10989 POR2X1_411/B POR2X1_329/A 0.06fF
C10990 PAND2X1_152/O POR2X1_151/Y -0.00fF
C10991 PAND2X1_502/CTRL2 POR2X1_42/Y 0.11fF
C10992 PAND2X1_499/CTRL2 POR2X1_39/B 0.03fF
C10993 D_GATE_222 POR2X1_332/CTRL 0.01fF
C10994 POR2X1_119/Y PAND2X1_785/Y 0.07fF
C10995 PAND2X1_23/Y POR2X1_186/B 0.94fF
C10996 PAND2X1_48/B POR2X1_151/Y 0.20fF
C10997 PAND2X1_71/O PAND2X1_71/Y 0.02fF
C10998 D_GATE_741 POR2X1_507/A 0.03fF
C10999 PAND2X1_216/B POR2X1_816/A 0.03fF
C11000 POR2X1_456/B POR2X1_576/Y 0.04fF
C11001 PAND2X1_226/CTRL2 POR2X1_192/B 0.07fF
C11002 POR2X1_60/Y PAND2X1_333/Y 0.00fF
C11003 POR2X1_62/Y PAND2X1_101/CTRL2 0.01fF
C11004 POR2X1_577/O POR2X1_569/Y 0.00fF
C11005 PAND2X1_633/O POR2X1_77/Y 0.17fF
C11006 POR2X1_285/B POR2X1_285/CTRL2 0.00fF
C11007 POR2X1_36/B POR2X1_158/B 0.01fF
C11008 POR2X1_83/Y POR2X1_293/Y 0.06fF
C11009 POR2X1_78/B PAND2X1_290/O 0.09fF
C11010 POR2X1_216/O POR2X1_116/Y 0.10fF
C11011 POR2X1_509/B PAND2X1_52/B 0.10fF
C11012 PAND2X1_55/Y POR2X1_512/CTRL 0.01fF
C11013 PAND2X1_787/Y POR2X1_77/Y 0.01fF
C11014 POR2X1_68/A POR2X1_652/A 0.05fF
C11015 POR2X1_83/Y PAND2X1_197/a_16_344# 0.04fF
C11016 POR2X1_855/B POR2X1_796/A -0.00fF
C11017 POR2X1_244/B POR2X1_568/B 0.03fF
C11018 PAND2X1_96/B PAND2X1_533/a_16_344# 0.02fF
C11019 POR2X1_739/a_16_28# POR2X1_730/Y 0.03fF
C11020 POR2X1_7/B PAND2X1_539/a_56_28# 0.00fF
C11021 POR2X1_85/Y PAND2X1_206/O 0.02fF
C11022 PAND2X1_575/O POR2X1_394/A 0.18fF
C11023 PAND2X1_469/B POR2X1_183/a_16_28# 0.02fF
C11024 PAND2X1_779/Y PAND2X1_779/O 0.02fF
C11025 POR2X1_62/Y PAND2X1_32/B 0.03fF
C11026 PAND2X1_819/CTRL2 POR2X1_260/A 0.01fF
C11027 PAND2X1_593/Y PAND2X1_537/CTRL 0.01fF
C11028 PAND2X1_631/A PAND2X1_6/A 0.03fF
C11029 POR2X1_686/B PAND2X1_72/A 0.01fF
C11030 PAND2X1_232/O POR2X1_260/A 0.01fF
C11031 POR2X1_137/Y PAND2X1_48/A 0.06fF
C11032 POR2X1_257/A PAND2X1_213/O 0.17fF
C11033 PAND2X1_613/O PAND2X1_9/Y 0.02fF
C11034 PAND2X1_109/CTRL2 D_GATE_222 0.04fF
C11035 POR2X1_72/CTRL2 PAND2X1_651/Y 0.05fF
C11036 POR2X1_86/CTRL PAND2X1_6/A 0.02fF
C11037 PAND2X1_134/CTRL PAND2X1_32/B 0.01fF
C11038 POR2X1_745/Y POR2X1_746/O 0.01fF
C11039 PAND2X1_467/Y PAND2X1_451/CTRL2 0.01fF
C11040 POR2X1_154/O PAND2X1_72/A 0.01fF
C11041 POR2X1_54/Y PAND2X1_612/B 0.01fF
C11042 POR2X1_567/A POR2X1_736/CTRL 0.03fF
C11043 POR2X1_283/A PAND2X1_156/A 0.03fF
C11044 PAND2X1_464/Y POR2X1_316/Y 0.05fF
C11045 PAND2X1_865/Y PAND2X1_575/CTRL 0.00fF
C11046 POR2X1_76/A POR2X1_446/B 0.03fF
C11047 POR2X1_439/Y POR2X1_440/CTRL 0.01fF
C11048 POR2X1_1/O PAND2X1_18/B 0.04fF
C11049 PAND2X1_349/A PAND2X1_141/CTRL2 0.01fF
C11050 POR2X1_186/O POR2X1_353/A 0.01fF
C11051 POR2X1_73/Y PAND2X1_326/B 4.70fF
C11052 POR2X1_48/A PAND2X1_9/Y 0.03fF
C11053 POR2X1_623/O PAND2X1_9/Y 0.01fF
C11054 POR2X1_119/Y PAND2X1_656/A 0.12fF
C11055 PAND2X1_761/CTRL2 D_INPUT_0 0.02fF
C11056 PAND2X1_310/CTRL POR2X1_260/A 0.01fF
C11057 POR2X1_826/Y D_INPUT_0 0.03fF
C11058 POR2X1_249/Y POR2X1_737/A 0.03fF
C11059 POR2X1_23/Y POR2X1_679/A 0.03fF
C11060 PAND2X1_26/CTRL2 D_INPUT_4 0.00fF
C11061 PAND2X1_404/O POR2X1_411/A 0.01fF
C11062 POR2X1_13/A POR2X1_386/Y 0.14fF
C11063 POR2X1_773/B POR2X1_294/A 0.10fF
C11064 POR2X1_62/Y POR2X1_673/Y 3.08fF
C11065 POR2X1_737/A POR2X1_737/a_16_28# 0.03fF
C11066 POR2X1_814/A POR2X1_489/O 0.02fF
C11067 POR2X1_83/B POR2X1_20/B 0.33fF
C11068 POR2X1_669/B POR2X1_604/O 0.01fF
C11069 POR2X1_122/O POR2X1_394/A 0.03fF
C11070 POR2X1_634/A POR2X1_859/CTRL2 0.04fF
C11071 PAND2X1_88/Y POR2X1_555/CTRL 0.01fF
C11072 POR2X1_376/B POR2X1_329/A 0.16fF
C11073 POR2X1_87/O POR2X1_68/B 0.06fF
C11074 POR2X1_644/O D_INPUT_0 0.02fF
C11075 POR2X1_139/CTRL2 POR2X1_138/A 0.00fF
C11076 POR2X1_48/A POR2X1_818/Y 1.20fF
C11077 POR2X1_816/CTRL POR2X1_750/B 0.00fF
C11078 POR2X1_271/Y POR2X1_275/Y 0.09fF
C11079 POR2X1_20/B POR2X1_626/Y -0.00fF
C11080 POR2X1_248/Y POR2X1_77/Y 0.01fF
C11081 POR2X1_126/a_16_28# POR2X1_37/Y 0.09fF
C11082 POR2X1_13/A PAND2X1_458/a_76_28# 0.02fF
C11083 POR2X1_564/B POR2X1_564/O 0.07fF
C11084 POR2X1_539/a_16_28# POR2X1_567/A 0.02fF
C11085 PAND2X1_48/A PAND2X1_18/B 0.11fF
C11086 POR2X1_20/B POR2X1_752/Y 0.03fF
C11087 PAND2X1_39/B POR2X1_794/B 0.12fF
C11088 POR2X1_34/a_16_28# POR2X1_34/A 0.07fF
C11089 POR2X1_119/Y POR2X1_300/Y 0.01fF
C11090 POR2X1_728/B POR2X1_814/A 0.04fF
C11091 PAND2X1_415/CTRL2 POR2X1_414/Y 0.00fF
C11092 POR2X1_45/Y POR2X1_677/Y 0.03fF
C11093 POR2X1_68/A PAND2X1_628/CTRL 0.01fF
C11094 PAND2X1_319/CTRL2 POR2X1_20/B 0.00fF
C11095 PAND2X1_404/A POR2X1_411/A 0.02fF
C11096 POR2X1_629/O POR2X1_629/B 0.01fF
C11097 PAND2X1_643/A PAND2X1_538/O 0.02fF
C11098 POR2X1_814/a_16_28# POR2X1_790/B 0.00fF
C11099 POR2X1_52/A POR2X1_329/A 0.08fF
C11100 POR2X1_751/Y POR2X1_39/B 0.00fF
C11101 POR2X1_814/A POR2X1_717/Y 0.03fF
C11102 POR2X1_119/Y PAND2X1_631/A 0.07fF
C11103 POR2X1_257/A PAND2X1_712/B 0.12fF
C11104 PAND2X1_199/B PAND2X1_199/a_76_28# 0.07fF
C11105 PAND2X1_88/CTRL2 POR2X1_66/A 0.30fF
C11106 POR2X1_609/Y POR2X1_102/Y 0.04fF
C11107 POR2X1_12/A INPUT_7 0.11fF
C11108 POR2X1_846/Y POR2X1_790/O 0.01fF
C11109 POR2X1_78/B POR2X1_471/A 0.07fF
C11110 POR2X1_254/A POR2X1_66/A 0.01fF
C11111 POR2X1_610/a_56_344# PAND2X1_41/B 0.00fF
C11112 PAND2X1_108/O PAND2X1_39/B 0.03fF
C11113 POR2X1_427/CTRL2 POR2X1_72/B 0.01fF
C11114 POR2X1_811/A POR2X1_783/O 0.00fF
C11115 POR2X1_542/CTRL POR2X1_552/A 0.11fF
C11116 POR2X1_49/CTRL POR2X1_409/B 0.02fF
C11117 POR2X1_66/A POR2X1_750/B 0.11fF
C11118 POR2X1_60/Y POR2X1_37/Y 0.03fF
C11119 POR2X1_66/B POR2X1_296/B 0.07fF
C11120 POR2X1_504/Y POR2X1_626/CTRL 0.01fF
C11121 POR2X1_102/Y POR2X1_420/Y 0.01fF
C11122 POR2X1_88/CTRL2 INPUT_0 0.04fF
C11123 PAND2X1_142/CTRL PAND2X1_72/A 0.01fF
C11124 PAND2X1_20/A POR2X1_33/a_16_28# 0.02fF
C11125 POR2X1_417/Y PAND2X1_212/B 0.03fF
C11126 POR2X1_188/A POR2X1_296/B 0.03fF
C11127 POR2X1_24/O POR2X1_29/A 0.01fF
C11128 POR2X1_291/O POR2X1_825/Y 0.00fF
C11129 PAND2X1_644/Y POR2X1_236/Y 0.04fF
C11130 POR2X1_486/O POR2X1_532/A 0.02fF
C11131 POR2X1_625/O POR2X1_37/Y 0.16fF
C11132 POR2X1_590/A POR2X1_389/Y 0.19fF
C11133 POR2X1_257/A PAND2X1_254/CTRL2 0.01fF
C11134 D_INPUT_5 INPUT_5 0.10fF
C11135 POR2X1_12/A INPUT_4 1.48fF
C11136 PAND2X1_844/a_76_28# PAND2X1_351/A 0.01fF
C11137 POR2X1_32/A PAND2X1_733/a_76_28# 0.02fF
C11138 PAND2X1_93/B POR2X1_215/CTRL 0.01fF
C11139 PAND2X1_571/A PAND2X1_571/Y 0.46fF
C11140 POR2X1_28/O INPUT_0 0.00fF
C11141 POR2X1_260/B POR2X1_121/Y 0.01fF
C11142 PAND2X1_20/A PAND2X1_20/CTRL2 0.01fF
C11143 PAND2X1_717/A PAND2X1_168/CTRL 0.01fF
C11144 POR2X1_262/Y PAND2X1_716/O 0.04fF
C11145 POR2X1_444/A VDD 0.04fF
C11146 POR2X1_334/B POR2X1_624/Y 0.03fF
C11147 POR2X1_27/a_16_28# POR2X1_38/Y 0.09fF
C11148 POR2X1_39/CTRL2 POR2X1_40/Y 0.01fF
C11149 POR2X1_32/A PAND2X1_778/O 0.02fF
C11150 POR2X1_816/a_16_28# POR2X1_816/A 0.01fF
C11151 PAND2X1_208/O POR2X1_40/Y 0.01fF
C11152 PAND2X1_602/Y POR2X1_600/Y 0.02fF
C11153 POR2X1_646/Y VDD 0.35fF
C11154 POR2X1_41/B PAND2X1_444/a_76_28# 0.02fF
C11155 POR2X1_330/O PAND2X1_52/B 0.01fF
C11156 PAND2X1_60/O POR2X1_35/Y 0.01fF
C11157 POR2X1_669/B PAND2X1_738/Y 0.10fF
C11158 POR2X1_814/A PAND2X1_503/CTRL2 0.05fF
C11159 PAND2X1_215/O PAND2X1_723/Y 0.14fF
C11160 POR2X1_57/A POR2X1_411/B 0.23fF
C11161 PAND2X1_93/B POR2X1_740/Y 0.11fF
C11162 PAND2X1_65/B POR2X1_330/Y 0.12fF
C11163 POR2X1_72/B PAND2X1_513/a_16_344# 0.01fF
C11164 POR2X1_67/a_16_28# PAND2X1_658/A 0.02fF
C11165 POR2X1_97/A POR2X1_776/B 0.00fF
C11166 POR2X1_68/A POR2X1_632/O 0.01fF
C11167 PAND2X1_810/A PAND2X1_366/Y 0.00fF
C11168 PAND2X1_460/Y PAND2X1_58/A 0.03fF
C11169 POR2X1_333/A POR2X1_781/O 0.34fF
C11170 POR2X1_43/B PAND2X1_477/O 0.01fF
C11171 PAND2X1_20/A PAND2X1_755/CTRL 0.00fF
C11172 POR2X1_855/O POR2X1_803/A 0.01fF
C11173 POR2X1_794/B POR2X1_325/A 0.03fF
C11174 POR2X1_383/A POR2X1_499/A 0.03fF
C11175 POR2X1_817/Y POR2X1_817/O 0.00fF
C11176 POR2X1_416/B PAND2X1_327/O 0.04fF
C11177 POR2X1_29/A PAND2X1_375/CTRL 0.03fF
C11178 PAND2X1_793/CTRL2 PAND2X1_793/A 0.01fF
C11179 PAND2X1_595/O POR2X1_294/B 0.16fF
C11180 POR2X1_56/CTRL POR2X1_293/Y 0.03fF
C11181 POR2X1_307/CTRL POR2X1_513/B 0.01fF
C11182 POR2X1_491/O PAND2X1_84/Y 0.01fF
C11183 POR2X1_260/B PAND2X1_536/a_76_28# 0.01fF
C11184 POR2X1_139/A POR2X1_260/B 0.01fF
C11185 POR2X1_836/B POR2X1_776/B 0.01fF
C11186 PAND2X1_863/a_16_344# PAND2X1_805/A 0.02fF
C11187 PAND2X1_784/O POR2X1_32/A 0.02fF
C11188 POR2X1_864/A POR2X1_598/CTRL 0.00fF
C11189 PAND2X1_349/B VDD 0.00fF
C11190 PAND2X1_852/A POR2X1_73/Y 0.03fF
C11191 PAND2X1_423/O POR2X1_480/A 0.06fF
C11192 POR2X1_257/A POR2X1_245/Y 0.12fF
C11193 POR2X1_96/A POR2X1_748/A 0.03fF
C11194 POR2X1_41/B PAND2X1_215/a_56_28# 0.00fF
C11195 POR2X1_431/CTRL POR2X1_129/Y 0.02fF
C11196 POR2X1_359/B POR2X1_814/A 0.02fF
C11197 POR2X1_116/O PAND2X1_65/B 0.01fF
C11198 POR2X1_78/A POR2X1_740/Y 0.03fF
C11199 PAND2X1_721/B POR2X1_42/Y 0.06fF
C11200 PAND2X1_318/CTRL2 POR2X1_417/Y 0.01fF
C11201 POR2X1_71/Y POR2X1_497/O 0.02fF
C11202 POR2X1_420/CTRL POR2X1_90/Y 0.01fF
C11203 POR2X1_595/Y VDD 0.01fF
C11204 PAND2X1_798/B PAND2X1_794/CTRL2 0.02fF
C11205 PAND2X1_650/A PAND2X1_9/Y 0.00fF
C11206 POR2X1_295/O POR2X1_7/B 0.16fF
C11207 PAND2X1_333/O VDD 0.00fF
C11208 PAND2X1_853/CTRL2 POR2X1_83/B 0.01fF
C11209 POR2X1_383/A POR2X1_76/A 0.04fF
C11210 D_GATE_811 POR2X1_121/B 0.03fF
C11211 POR2X1_97/A POR2X1_577/CTRL2 0.01fF
C11212 POR2X1_286/B POR2X1_773/B 0.04fF
C11213 POR2X1_255/Y POR2X1_32/A 0.03fF
C11214 POR2X1_54/Y POR2X1_773/CTRL 0.01fF
C11215 POR2X1_60/Y POR2X1_293/Y 0.03fF
C11216 POR2X1_416/B POR2X1_234/A 0.03fF
C11217 POR2X1_463/Y POR2X1_472/B 0.01fF
C11218 PAND2X1_650/CTRL2 POR2X1_409/B 0.01fF
C11219 POR2X1_528/Y POR2X1_613/CTRL 0.08fF
C11220 PAND2X1_556/B POR2X1_236/Y 0.03fF
C11221 PAND2X1_341/B PAND2X1_206/B 0.22fF
C11222 POR2X1_422/O POR2X1_7/A 0.01fF
C11223 POR2X1_327/Y POR2X1_864/A 0.00fF
C11224 POR2X1_348/O PAND2X1_93/B 0.01fF
C11225 POR2X1_315/Y PAND2X1_444/CTRL 0.04fF
C11226 PAND2X1_599/O POR2X1_330/Y 0.02fF
C11227 POR2X1_596/A POR2X1_834/CTRL 0.01fF
C11228 POR2X1_254/A POR2X1_222/Y 0.11fF
C11229 POR2X1_814/B PAND2X1_372/a_16_344# 0.02fF
C11230 POR2X1_387/O POR2X1_386/Y 0.03fF
C11231 POR2X1_257/A PAND2X1_579/A 0.00fF
C11232 PAND2X1_741/a_16_344# PAND2X1_473/B 0.02fF
C11233 POR2X1_52/A PAND2X1_859/O 0.03fF
C11234 POR2X1_811/CTRL2 POR2X1_780/B 0.04fF
C11235 POR2X1_525/CTRL POR2X1_763/Y 0.07fF
C11236 POR2X1_13/A POR2X1_397/Y 0.03fF
C11237 POR2X1_502/A POR2X1_663/O 0.02fF
C11238 PAND2X1_36/O D_INPUT_6 0.02fF
C11239 POR2X1_222/Y POR2X1_750/B 0.22fF
C11240 POR2X1_416/B POR2X1_281/Y 0.01fF
C11241 PAND2X1_272/m4_208_n4# POR2X1_112/Y 0.09fF
C11242 POR2X1_66/B POR2X1_267/Y 0.01fF
C11243 PAND2X1_470/CTRL POR2X1_83/B 0.00fF
C11244 POR2X1_43/B POR2X1_40/Y 0.33fF
C11245 PAND2X1_852/CTRL2 POR2X1_65/A 0.02fF
C11246 PAND2X1_778/CTRL2 POR2X1_293/Y 0.01fF
C11247 INPUT_0 PAND2X1_558/a_76_28# 0.02fF
C11248 POR2X1_284/B PAND2X1_57/B 0.01fF
C11249 PAND2X1_254/Y POR2X1_236/Y 0.03fF
C11250 POR2X1_775/A POR2X1_186/Y 0.03fF
C11251 POR2X1_226/Y POR2X1_42/Y 0.02fF
C11252 PAND2X1_787/Y PAND2X1_592/a_76_28# 0.06fF
C11253 POR2X1_465/B POR2X1_563/O 0.18fF
C11254 POR2X1_677/CTRL2 PAND2X1_658/B 0.08fF
C11255 PAND2X1_127/a_16_344# POR2X1_445/A 0.02fF
C11256 PAND2X1_607/CTRL2 PAND2X1_56/A 0.01fF
C11257 PAND2X1_650/a_56_28# D_INPUT_0 0.00fF
C11258 POR2X1_389/CTRL2 POR2X1_480/A 0.10fF
C11259 POR2X1_236/Y POR2X1_395/CTRL 0.01fF
C11260 PAND2X1_357/Y POR2X1_331/Y 0.09fF
C11261 POR2X1_66/A POR2X1_200/A 0.05fF
C11262 PAND2X1_433/O POR2X1_807/A 0.02fF
C11263 PAND2X1_13/O POR2X1_222/Y 0.01fF
C11264 POR2X1_62/Y PAND2X1_9/Y 0.07fF
C11265 POR2X1_615/CTRL PAND2X1_6/A 0.03fF
C11266 POR2X1_68/A POR2X1_274/Y 0.03fF
C11267 POR2X1_413/Y VDD 0.12fF
C11268 PAND2X1_90/Y POR2X1_732/B 0.06fF
C11269 PAND2X1_644/Y POR2X1_757/Y 0.03fF
C11270 POR2X1_590/A POR2X1_713/B 0.01fF
C11271 PAND2X1_88/CTRL POR2X1_68/B 0.04fF
C11272 POR2X1_730/Y POR2X1_567/B 0.05fF
C11273 POR2X1_495/Y POR2X1_511/Y 0.03fF
C11274 POR2X1_43/B PAND2X1_849/O 0.01fF
C11275 POR2X1_96/A POR2X1_79/Y 0.04fF
C11276 POR2X1_330/Y POR2X1_541/CTRL 0.02fF
C11277 POR2X1_38/B POR2X1_40/Y 0.03fF
C11278 PAND2X1_339/Y POR2X1_5/Y 0.06fF
C11279 POR2X1_100/CTRL POR2X1_99/A 0.01fF
C11280 PAND2X1_651/Y PAND2X1_61/Y 0.03fF
C11281 POR2X1_532/A POR2X1_750/B 0.14fF
C11282 POR2X1_48/Y VDD 0.01fF
C11283 POR2X1_686/A PAND2X1_69/A 0.02fF
C11284 POR2X1_13/A PAND2X1_784/CTRL 0.01fF
C11285 POR2X1_467/Y PAND2X1_534/CTRL2 0.01fF
C11286 POR2X1_811/B POR2X1_780/B 0.11fF
C11287 PAND2X1_341/B POR2X1_65/Y 0.01fF
C11288 POR2X1_68/B PAND2X1_41/B 1.64fF
C11289 POR2X1_196/Y PAND2X1_52/Y 0.31fF
C11290 POR2X1_649/B POR2X1_476/a_76_344# 0.01fF
C11291 PAND2X1_48/B PAND2X1_321/m4_208_n4# 0.07fF
C11292 POR2X1_466/A POR2X1_703/Y 0.05fF
C11293 POR2X1_259/O POR2X1_555/B 0.02fF
C11294 PAND2X1_652/A VDD 0.82fF
C11295 POR2X1_220/B POR2X1_353/A 5.09fF
C11296 PAND2X1_675/A POR2X1_481/A 0.03fF
C11297 PAND2X1_93/B POR2X1_774/A 0.07fF
C11298 POR2X1_667/A PAND2X1_559/CTRL 0.02fF
C11299 PAND2X1_23/CTRL2 PAND2X1_60/B 0.01fF
C11300 PAND2X1_61/Y PAND2X1_844/B 0.02fF
C11301 POR2X1_68/A POR2X1_370/Y 0.01fF
C11302 PAND2X1_55/Y POR2X1_121/Y 0.03fF
C11303 PAND2X1_784/CTRL2 POR2X1_293/Y 0.01fF
C11304 POR2X1_55/Y PAND2X1_515/O 0.17fF
C11305 POR2X1_748/A POR2X1_7/A 3.27fF
C11306 POR2X1_278/Y POR2X1_45/Y 0.07fF
C11307 POR2X1_686/a_16_28# POR2X1_750/B 0.02fF
C11308 POR2X1_43/B PAND2X1_659/B 0.03fF
C11309 POR2X1_660/Y POR2X1_353/A 0.00fF
C11310 POR2X1_483/A POR2X1_702/A 0.00fF
C11311 POR2X1_490/Y PAND2X1_716/B 0.73fF
C11312 PAND2X1_140/O POR2X1_387/Y 0.14fF
C11313 POR2X1_509/B POR2X1_350/B 0.06fF
C11314 POR2X1_57/A POR2X1_376/B 0.16fF
C11315 POR2X1_344/CTRL POR2X1_383/A 0.07fF
C11316 PAND2X1_6/Y POR2X1_130/A 0.03fF
C11317 POR2X1_723/O POR2X1_723/B 0.01fF
C11318 POR2X1_357/CTRL POR2X1_220/B 0.12fF
C11319 POR2X1_538/O POR2X1_566/A 0.01fF
C11320 POR2X1_186/Y POR2X1_162/Y 0.00fF
C11321 POR2X1_43/B POR2X1_586/CTRL 0.01fF
C11322 POR2X1_804/A VDD 4.35fF
C11323 POR2X1_197/Y POR2X1_61/Y 0.02fF
C11324 PAND2X1_206/CTRL POR2X1_73/Y 0.01fF
C11325 POR2X1_459/O POR2X1_459/B 0.00fF
C11326 PAND2X1_21/a_16_344# PAND2X1_32/B 0.02fF
C11327 PAND2X1_6/Y POR2X1_566/A 0.09fF
C11328 POR2X1_163/Y PAND2X1_725/CTRL2 0.11fF
C11329 PAND2X1_309/CTRL POR2X1_68/A 0.01fF
C11330 POR2X1_223/a_16_28# POR2X1_222/Y 0.02fF
C11331 POR2X1_406/A POR2X1_46/Y 0.04fF
C11332 POR2X1_247/a_16_28# POR2X1_294/B 0.05fF
C11333 POR2X1_555/A POR2X1_510/Y 0.03fF
C11334 POR2X1_304/O PAND2X1_454/B 0.00fF
C11335 PAND2X1_55/Y POR2X1_556/O 0.01fF
C11336 PAND2X1_116/CTRL POR2X1_283/A 0.00fF
C11337 VDD POR2X1_535/A 0.00fF
C11338 POR2X1_119/Y POR2X1_271/a_76_344# 0.02fF
C11339 INPUT_1 POR2X1_495/CTRL2 0.00fF
C11340 POR2X1_66/A PAND2X1_143/CTRL2 0.03fF
C11341 POR2X1_294/B POR2X1_565/CTRL 0.01fF
C11342 POR2X1_152/Y VDD 0.22fF
C11343 POR2X1_78/A POR2X1_774/A 0.03fF
C11344 PAND2X1_3/a_16_344# POR2X1_750/B 0.02fF
C11345 POR2X1_62/CTRL2 PAND2X1_6/A 0.00fF
C11346 PAND2X1_407/CTRL POR2X1_39/B 0.08fF
C11347 POR2X1_327/a_16_28# POR2X1_264/Y 0.03fF
C11348 PAND2X1_48/B POR2X1_790/A 0.03fF
C11349 PAND2X1_8/Y PAND2X1_670/CTRL 0.07fF
C11350 POR2X1_97/A POR2X1_192/B 0.19fF
C11351 PAND2X1_659/O POR2X1_91/Y 0.07fF
C11352 POR2X1_319/A POR2X1_568/B 0.03fF
C11353 PAND2X1_624/O POR2X1_283/A 0.08fF
C11354 POR2X1_480/A POR2X1_590/CTRL2 0.05fF
C11355 POR2X1_96/A PAND2X1_785/A 0.01fF
C11356 PAND2X1_23/Y POR2X1_515/Y 0.01fF
C11357 PAND2X1_41/B POR2X1_502/O 0.08fF
C11358 POR2X1_56/B POR2X1_90/Y 0.02fF
C11359 PAND2X1_91/O POR2X1_169/A 0.06fF
C11360 PAND2X1_140/A POR2X1_107/a_56_344# 0.00fF
C11361 POR2X1_865/CTRL POR2X1_784/A 0.04fF
C11362 POR2X1_85/Y POR2X1_490/a_16_28# 0.01fF
C11363 POR2X1_186/O POR2X1_750/B 0.02fF
C11364 POR2X1_14/Y PAND2X1_156/A 0.05fF
C11365 PAND2X1_23/Y POR2X1_208/Y 0.15fF
C11366 PAND2X1_182/A PAND2X1_182/a_76_28# 0.02fF
C11367 POR2X1_417/O POR2X1_293/Y 0.16fF
C11368 PAND2X1_665/CTRL POR2X1_66/A 0.01fF
C11369 PAND2X1_453/A PAND2X1_156/A 0.05fF
C11370 POR2X1_351/Y POR2X1_350/CTRL2 0.01fF
C11371 PAND2X1_220/Y PAND2X1_343/O 0.08fF
C11372 POR2X1_57/A POR2X1_52/A 0.22fF
C11373 PAND2X1_661/Y PAND2X1_596/a_76_28# 0.05fF
C11374 POR2X1_416/B POR2X1_77/O 0.01fF
C11375 PAND2X1_473/B PAND2X1_728/O 0.04fF
C11376 PAND2X1_710/O POR2X1_701/Y 0.15fF
C11377 PAND2X1_23/Y POR2X1_542/B 0.02fF
C11378 POR2X1_346/CTRL2 PAND2X1_55/Y 0.01fF
C11379 POR2X1_804/A POR2X1_741/Y 2.01fF
C11380 PAND2X1_48/B POR2X1_865/B 0.07fF
C11381 POR2X1_614/A POR2X1_341/O 0.00fF
C11382 PAND2X1_48/B PAND2X1_88/Y 0.07fF
C11383 PAND2X1_94/A PAND2X1_54/O 0.05fF
C11384 PAND2X1_46/CTRL2 PAND2X1_71/Y 0.01fF
C11385 PAND2X1_575/A POR2X1_73/Y 0.03fF
C11386 POR2X1_57/A PAND2X1_398/CTRL2 0.03fF
C11387 POR2X1_78/CTRL2 POR2X1_844/B 0.01fF
C11388 POR2X1_57/A PAND2X1_317/Y 0.00fF
C11389 PAND2X1_175/O VDD 0.00fF
C11390 POR2X1_40/Y POR2X1_183/CTRL 0.01fF
C11391 POR2X1_57/A POR2X1_152/A 0.03fF
C11392 POR2X1_46/Y PAND2X1_349/A 0.05fF
C11393 POR2X1_84/O POR2X1_532/A 0.01fF
C11394 POR2X1_814/A PAND2X1_257/O 0.14fF
C11395 POR2X1_786/A PAND2X1_60/B 0.04fF
C11396 POR2X1_341/A POR2X1_579/CTRL 0.06fF
C11397 POR2X1_83/Y POR2X1_60/A 0.02fF
C11398 POR2X1_65/A PAND2X1_170/CTRL2 0.02fF
C11399 POR2X1_186/Y POR2X1_339/Y 0.10fF
C11400 POR2X1_355/B POR2X1_738/A 0.03fF
C11401 PAND2X1_803/Y POR2X1_42/Y 0.03fF
C11402 POR2X1_780/B POR2X1_783/B 0.25fF
C11403 POR2X1_334/B POR2X1_493/CTRL 0.28fF
C11404 PAND2X1_848/B POR2X1_38/B 1.40fF
C11405 PAND2X1_94/A PAND2X1_57/B 0.10fF
C11406 POR2X1_547/B POR2X1_6/CTRL 0.00fF
C11407 PAND2X1_313/O VDD 0.00fF
C11408 POR2X1_740/Y PAND2X1_306/O 0.01fF
C11409 POR2X1_327/Y POR2X1_362/B 0.02fF
C11410 POR2X1_41/B PAND2X1_196/O 0.03fF
C11411 POR2X1_804/A PAND2X1_32/B 0.16fF
C11412 PAND2X1_674/CTRL PAND2X1_60/B 0.01fF
C11413 POR2X1_48/A POR2X1_747/O 0.01fF
C11414 POR2X1_41/B POR2X1_83/CTRL 0.00fF
C11415 PAND2X1_442/a_76_28# POR2X1_444/Y 0.04fF
C11416 PAND2X1_6/Y POR2X1_573/A 0.03fF
C11417 POR2X1_43/a_16_28# POR2X1_37/Y 0.05fF
C11418 POR2X1_502/A POR2X1_675/Y 0.03fF
C11419 PAND2X1_358/A POR2X1_236/Y 0.10fF
C11420 POR2X1_324/Y PAND2X1_41/B 0.01fF
C11421 POR2X1_650/A PAND2X1_48/A 0.03fF
C11422 POR2X1_677/Y POR2X1_271/B 2.54fF
C11423 PAND2X1_70/CTRL2 PAND2X1_3/B 0.00fF
C11424 POR2X1_197/Y POR2X1_35/Y 0.02fF
C11425 POR2X1_43/Y PAND2X1_124/Y 0.45fF
C11426 PAND2X1_631/A PAND2X1_456/CTRL2 0.01fF
C11427 POR2X1_7/B POR2X1_310/Y 0.04fF
C11428 PAND2X1_127/a_76_28# POR2X1_78/B 0.02fF
C11429 PAND2X1_126/CTRL2 PAND2X1_6/A 0.02fF
C11430 INPUT_1 POR2X1_669/O 0.01fF
C11431 POR2X1_596/A POR2X1_644/A 0.00fF
C11432 PAND2X1_840/A PAND2X1_349/A 0.00fF
C11433 POR2X1_119/Y POR2X1_763/A 0.07fF
C11434 POR2X1_68/A PAND2X1_63/B 0.03fF
C11435 PAND2X1_65/B POR2X1_337/Y 0.71fF
C11436 POR2X1_664/CTRL POR2X1_664/Y 0.01fF
C11437 POR2X1_207/A POR2X1_195/a_76_344# 0.01fF
C11438 POR2X1_502/A POR2X1_544/B 1.43fF
C11439 PAND2X1_55/Y POR2X1_576/CTRL 0.01fF
C11440 PAND2X1_6/Y POR2X1_774/O 0.16fF
C11441 POR2X1_169/B PAND2X1_65/B 0.01fF
C11442 PAND2X1_476/A POR2X1_230/CTRL 0.00fF
C11443 PAND2X1_241/CTRL PAND2X1_308/Y 0.01fF
C11444 POR2X1_271/A PAND2X1_254/Y 0.03fF
C11445 POR2X1_93/A POR2X1_619/A 0.04fF
C11446 PAND2X1_785/O POR2X1_91/Y 0.02fF
C11447 POR2X1_322/Y POR2X1_73/Y 0.12fF
C11448 POR2X1_575/CTRL2 POR2X1_573/A 0.01fF
C11449 POR2X1_170/O POR2X1_566/B 0.02fF
C11450 POR2X1_65/A POR2X1_517/CTRL 0.01fF
C11451 POR2X1_13/A POR2X1_131/A 0.01fF
C11452 POR2X1_691/a_76_344# POR2X1_855/B 0.02fF
C11453 PAND2X1_552/a_76_28# PAND2X1_552/B 0.02fF
C11454 VDD PAND2X1_506/Y 0.09fF
C11455 PAND2X1_329/O POR2X1_532/A 0.05fF
C11456 POR2X1_674/Y POR2X1_331/CTRL 0.01fF
C11457 POR2X1_383/A POR2X1_540/A 0.05fF
C11458 PAND2X1_778/Y POR2X1_245/Y 0.03fF
C11459 POR2X1_192/Y POR2X1_564/O 0.04fF
C11460 POR2X1_750/Y POR2X1_816/A 0.08fF
C11461 POR2X1_387/Y POR2X1_142/Y 0.07fF
C11462 POR2X1_416/B PAND2X1_35/B 0.05fF
C11463 POR2X1_569/A POR2X1_500/Y 0.12fF
C11464 POR2X1_96/A PAND2X1_730/A 0.04fF
C11465 POR2X1_816/A POR2X1_171/a_56_344# 0.00fF
C11466 D_INPUT_1 POR2X1_750/Y 0.13fF
C11467 POR2X1_43/Y POR2X1_83/B 0.03fF
C11468 POR2X1_634/A PAND2X1_52/B 0.17fF
C11469 PAND2X1_553/B POR2X1_183/O 0.03fF
C11470 POR2X1_119/Y POR2X1_234/Y 0.03fF
C11471 POR2X1_68/B POR2X1_561/CTRL 0.01fF
C11472 POR2X1_55/Y PAND2X1_156/A 0.05fF
C11473 POR2X1_54/Y POR2X1_67/Y 0.03fF
C11474 PAND2X1_724/CTRL PAND2X1_714/Y -0.01fF
C11475 POR2X1_294/B PAND2X1_48/A 0.35fF
C11476 PAND2X1_351/m4_208_n4# POR2X1_293/Y 0.12fF
C11477 POR2X1_602/B PAND2X1_72/A 0.01fF
C11478 PAND2X1_403/O POR2X1_37/Y 0.25fF
C11479 POR2X1_12/A POR2X1_18/O 0.01fF
C11480 PAND2X1_6/Y POR2X1_344/Y 0.03fF
C11481 POR2X1_567/A POR2X1_776/B 0.00fF
C11482 POR2X1_493/B POR2X1_493/CTRL2 0.13fF
C11483 POR2X1_539/A POR2X1_383/A 0.07fF
C11484 POR2X1_366/Y POR2X1_192/B 0.36fF
C11485 POR2X1_404/Y POR2X1_4/Y 0.03fF
C11486 PAND2X1_824/B POR2X1_447/CTRL2 0.04fF
C11487 PAND2X1_48/B POR2X1_359/O 0.01fF
C11488 POR2X1_566/B POR2X1_854/B 0.39fF
C11489 POR2X1_180/A POR2X1_854/B 0.05fF
C11490 POR2X1_95/a_16_28# POR2X1_51/A 0.05fF
C11491 PAND2X1_566/Y PAND2X1_345/Y 0.03fF
C11492 POR2X1_184/Y PAND2X1_141/CTRL2 0.00fF
C11493 POR2X1_85/O PAND2X1_35/Y 0.01fF
C11494 PAND2X1_6/Y POR2X1_349/CTRL2 0.00fF
C11495 POR2X1_16/A POR2X1_167/CTRL 0.01fF
C11496 POR2X1_762/CTRL2 D_INPUT_6 0.05fF
C11497 PAND2X1_777/CTRL POR2X1_387/Y 0.04fF
C11498 POR2X1_164/Y PAND2X1_569/B 0.01fF
C11499 PAND2X1_96/B POR2X1_652/A 0.03fF
C11500 POR2X1_68/A POR2X1_552/A 0.01fF
C11501 PAND2X1_466/B POR2X1_424/Y 0.14fF
C11502 PAND2X1_206/A POR2X1_20/B 0.03fF
C11503 PAND2X1_63/B POR2X1_376/O 0.01fF
C11504 POR2X1_431/CTRL POR2X1_37/Y 0.01fF
C11505 PAND2X1_833/a_76_28# POR2X1_77/Y 0.02fF
C11506 POR2X1_439/Y POR2X1_863/A 0.09fF
C11507 POR2X1_681/a_16_28# POR2X1_681/Y 0.02fF
C11508 POR2X1_407/Y PAND2X1_3/B 0.03fF
C11509 PAND2X1_48/B POR2X1_568/B 0.05fF
C11510 POR2X1_130/A PAND2X1_52/B 0.05fF
C11511 PAND2X1_658/A PAND2X1_860/O 0.01fF
C11512 PAND2X1_785/O POR2X1_109/Y 0.01fF
C11513 POR2X1_271/CTRL2 POR2X1_411/B 0.01fF
C11514 POR2X1_452/A POR2X1_750/B 0.01fF
C11515 POR2X1_65/CTRL D_INPUT_0 0.01fF
C11516 PAND2X1_862/B PAND2X1_862/CTRL 0.01fF
C11517 POR2X1_566/A PAND2X1_52/B 0.07fF
C11518 PAND2X1_632/A POR2X1_153/Y 0.05fF
C11519 POR2X1_71/Y PAND2X1_501/O 0.01fF
C11520 PAND2X1_659/Y PAND2X1_676/O 0.16fF
C11521 POR2X1_203/O PAND2X1_48/A 0.01fF
C11522 POR2X1_270/CTRL2 POR2X1_567/A -0.00fF
C11523 PAND2X1_111/B PAND2X1_48/A 0.01fF
C11524 POR2X1_38/Y PAND2X1_737/O 0.15fF
C11525 INPUT_1 PAND2X1_701/CTRL 0.01fF
C11526 PAND2X1_39/B POR2X1_647/O 0.01fF
C11527 PAND2X1_793/Y PAND2X1_332/Y 0.03fF
C11528 POR2X1_293/Y PAND2X1_351/A 0.03fF
C11529 POR2X1_456/B POR2X1_733/Y 0.33fF
C11530 PAND2X1_242/O POR2X1_77/Y 0.04fF
C11531 PAND2X1_472/CTRL POR2X1_153/Y 0.01fF
C11532 POR2X1_73/Y PAND2X1_860/O 0.17fF
C11533 POR2X1_16/A PAND2X1_200/B 0.02fF
C11534 PAND2X1_338/B PAND2X1_338/CTRL 0.04fF
C11535 POR2X1_260/A POR2X1_673/B 0.05fF
C11536 POR2X1_74/O POR2X1_271/A 0.01fF
C11537 POR2X1_334/Y POR2X1_97/O 0.04fF
C11538 POR2X1_814/A POR2X1_330/Y 0.15fF
C11539 POR2X1_518/Y POR2X1_77/Y 0.01fF
C11540 POR2X1_508/B POR2X1_854/B 0.05fF
C11541 PAND2X1_472/A POR2X1_77/Y 0.03fF
C11542 POR2X1_23/Y PAND2X1_407/O 0.05fF
C11543 POR2X1_383/O POR2X1_520/A 0.01fF
C11544 PAND2X1_483/O PAND2X1_508/Y 0.00fF
C11545 PAND2X1_73/Y POR2X1_556/A 0.08fF
C11546 POR2X1_257/A D_INPUT_0 0.03fF
C11547 POR2X1_329/A PAND2X1_733/CTRL 0.02fF
C11548 POR2X1_861/O PAND2X1_72/A 0.02fF
C11549 POR2X1_725/O POR2X1_712/Y 0.02fF
C11550 POR2X1_632/Y POR2X1_573/A 0.03fF
C11551 PAND2X1_838/B POR2X1_669/B 0.56fF
C11552 POR2X1_712/Y PAND2X1_72/A 0.03fF
C11553 POR2X1_844/B PAND2X1_52/B 0.03fF
C11554 PAND2X1_213/Y POR2X1_39/B 0.03fF
C11555 POR2X1_557/A POR2X1_4/Y 0.03fF
C11556 POR2X1_675/Y POR2X1_188/Y 0.39fF
C11557 PAND2X1_717/A PAND2X1_803/A 0.03fF
C11558 POR2X1_506/O POR2X1_508/B 0.01fF
C11559 PAND2X1_437/a_56_28# POR2X1_192/Y 0.00fF
C11560 POR2X1_540/Y POR2X1_260/A 0.00fF
C11561 PAND2X1_282/CTRL2 POR2X1_260/B 0.01fF
C11562 PAND2X1_206/B PAND2X1_340/O 0.00fF
C11563 POR2X1_452/a_16_28# POR2X1_121/B 0.09fF
C11564 PAND2X1_403/O POR2X1_293/Y 0.17fF
C11565 PAND2X1_63/B PAND2X1_529/CTRL 0.01fF
C11566 POR2X1_602/CTRL2 POR2X1_296/B 0.03fF
C11567 POR2X1_32/CTRL2 POR2X1_29/Y 0.03fF
C11568 PAND2X1_60/B POR2X1_716/O 0.01fF
C11569 POR2X1_649/a_16_28# POR2X1_643/A 0.00fF
C11570 PAND2X1_212/B PAND2X1_212/O 0.00fF
C11571 POR2X1_458/Y POR2X1_220/Y 0.07fF
C11572 POR2X1_270/Y POR2X1_269/CTRL2 0.00fF
C11573 PAND2X1_269/O INPUT_0 0.15fF
C11574 POR2X1_304/Y POR2X1_329/A 0.01fF
C11575 PAND2X1_606/CTRL POR2X1_102/Y 0.01fF
C11576 PAND2X1_221/Y PAND2X1_730/CTRL2 0.00fF
C11577 POR2X1_475/CTRL POR2X1_734/A 0.02fF
C11578 PAND2X1_96/B PAND2X1_125/CTRL2 0.01fF
C11579 PAND2X1_862/B POR2X1_329/A 0.03fF
C11580 PAND2X1_657/CTRL POR2X1_23/Y 0.02fF
C11581 PAND2X1_666/CTRL2 PAND2X1_73/Y 0.03fF
C11582 POR2X1_774/O PAND2X1_52/B 0.01fF
C11583 PAND2X1_352/A PAND2X1_220/A 0.07fF
C11584 POR2X1_703/A POR2X1_736/A 0.05fF
C11585 PAND2X1_447/O VDD 0.00fF
C11586 POR2X1_265/Y PAND2X1_476/A 0.03fF
C11587 POR2X1_416/B PAND2X1_514/O 0.02fF
C11588 PAND2X1_492/CTRL POR2X1_556/A 0.01fF
C11589 PAND2X1_20/A POR2X1_33/A 0.02fF
C11590 POR2X1_497/CTRL2 POR2X1_37/Y 0.03fF
C11591 POR2X1_68/A POR2X1_837/A 0.01fF
C11592 PAND2X1_96/B PAND2X1_628/CTRL 0.10fF
C11593 POR2X1_864/A PAND2X1_760/CTRL2 0.00fF
C11594 POR2X1_499/A INPUT_0 0.03fF
C11595 POR2X1_411/B PAND2X1_84/Y 0.03fF
C11596 POR2X1_559/A PAND2X1_517/m4_208_n4# 0.08fF
C11597 POR2X1_48/A PAND2X1_403/B 0.08fF
C11598 PAND2X1_678/CTRL PAND2X1_480/B 0.27fF
C11599 POR2X1_567/B POR2X1_439/CTRL 0.15fF
C11600 PAND2X1_9/O D_INPUT_0 0.02fF
C11601 POR2X1_66/B POR2X1_98/CTRL2 0.02fF
C11602 PAND2X1_217/B PAND2X1_205/A 0.05fF
C11603 POR2X1_119/Y PAND2X1_850/Y 0.23fF
C11604 POR2X1_23/Y PAND2X1_390/Y 0.03fF
C11605 POR2X1_450/O POR2X1_121/B 0.06fF
C11606 POR2X1_558/B POR2X1_777/B 0.01fF
C11607 POR2X1_51/A POR2X1_744/Y 0.01fF
C11608 PAND2X1_817/CTRL POR2X1_29/A 0.01fF
C11609 PAND2X1_817/O PAND2X1_381/Y 0.15fF
C11610 POR2X1_257/A POR2X1_697/a_16_28# 0.03fF
C11611 POR2X1_41/B POR2X1_484/Y 0.01fF
C11612 PAND2X1_437/O PAND2X1_60/B 0.15fF
C11613 POR2X1_220/B POR2X1_750/B 0.03fF
C11614 POR2X1_78/A POR2X1_474/CTRL 0.01fF
C11615 PAND2X1_222/O INPUT_0 0.05fF
C11616 PAND2X1_802/a_16_344# PAND2X1_798/Y 0.03fF
C11617 POR2X1_49/Y D_INPUT_0 0.95fF
C11618 D_INPUT_5 PAND2X1_587/Y 0.00fF
C11619 PAND2X1_222/A INPUT_0 1.23fF
C11620 POR2X1_96/A PAND2X1_203/a_16_344# 0.03fF
C11621 PAND2X1_65/B POR2X1_558/B 0.03fF
C11622 POR2X1_326/a_76_344# POR2X1_568/A 0.00fF
C11623 POR2X1_23/Y POR2X1_697/CTRL 0.08fF
C11624 PAND2X1_860/A PAND2X1_861/CTRL 0.01fF
C11625 POR2X1_422/Y POR2X1_72/B 0.01fF
C11626 POR2X1_278/Y PAND2X1_205/CTRL2 0.03fF
C11627 POR2X1_466/A PAND2X1_90/Y 0.05fF
C11628 PAND2X1_48/B POR2X1_341/A 0.07fF
C11629 PAND2X1_23/Y POR2X1_776/A 0.90fF
C11630 POR2X1_415/A POR2X1_617/O 0.05fF
C11631 POR2X1_496/Y POR2X1_627/CTRL 0.07fF
C11632 PAND2X1_288/m4_208_n4# POR2X1_7/B 0.09fF
C11633 POR2X1_20/B PAND2X1_357/Y 0.01fF
C11634 POR2X1_60/A PAND2X1_541/O 0.17fF
C11635 POR2X1_624/Y POR2X1_565/CTRL2 0.05fF
C11636 POR2X1_665/CTRL POR2X1_665/A 0.01fF
C11637 PAND2X1_304/a_16_344# PAND2X1_56/A 0.01fF
C11638 POR2X1_83/B INPUT_7 0.03fF
C11639 POR2X1_556/A POR2X1_631/B 0.03fF
C11640 POR2X1_517/O POR2X1_667/A 0.03fF
C11641 POR2X1_516/CTRL POR2X1_257/A 0.01fF
C11642 POR2X1_83/B POR2X1_237/CTRL2 0.03fF
C11643 PAND2X1_201/O PAND2X1_341/A 0.02fF
C11644 PAND2X1_73/O PAND2X1_41/B 0.01fF
C11645 POR2X1_678/CTRL PAND2X1_69/A 0.01fF
C11646 POR2X1_83/B POR2X1_48/CTRL2 0.01fF
C11647 POR2X1_852/B POR2X1_330/Y 0.07fF
C11648 POR2X1_694/CTRL2 POR2X1_257/A 0.00fF
C11649 POR2X1_48/A POR2X1_232/CTRL2 0.03fF
C11650 POR2X1_68/A POR2X1_676/O 0.02fF
C11651 POR2X1_407/A POR2X1_676/CTRL 0.04fF
C11652 PAND2X1_474/A POR2X1_40/Y 0.00fF
C11653 POR2X1_416/B POR2X1_39/B 17.13fF
C11654 POR2X1_41/B PAND2X1_264/a_76_28# 0.01fF
C11655 PAND2X1_808/Y PAND2X1_287/Y 0.03fF
C11656 POR2X1_196/O VDD -0.00fF
C11657 POR2X1_13/A POR2X1_667/Y 0.16fF
C11658 PAND2X1_139/B POR2X1_102/Y 0.02fF
C11659 D_INPUT_0 PAND2X1_553/B 0.03fF
C11660 POR2X1_569/O PAND2X1_41/B 0.01fF
C11661 PAND2X1_23/Y POR2X1_856/B 0.05fF
C11662 POR2X1_32/A POR2X1_46/Y 0.60fF
C11663 PAND2X1_430/CTRL2 POR2X1_750/B 0.01fF
C11664 PAND2X1_650/CTRL PAND2X1_9/Y 0.01fF
C11665 PAND2X1_73/Y POR2X1_445/CTRL 0.01fF
C11666 POR2X1_446/B PAND2X1_69/A 0.00fF
C11667 POR2X1_260/B POR2X1_391/Y 0.04fF
C11668 POR2X1_54/Y POR2X1_649/B 0.01fF
C11669 PAND2X1_612/B POR2X1_462/B 0.00fF
C11670 POR2X1_20/B PAND2X1_344/a_16_344# 0.02fF
C11671 PAND2X1_57/B PAND2X1_11/Y 0.05fF
C11672 PAND2X1_602/Y PAND2X1_644/Y 7.72fF
C11673 PAND2X1_240/CTRL POR2X1_5/Y 0.00fF
C11674 PAND2X1_282/CTRL2 PAND2X1_55/Y 0.02fF
C11675 PAND2X1_195/CTRL VDD -0.00fF
C11676 PAND2X1_140/A POR2X1_20/B 0.03fF
C11677 D_INPUT_0 PAND2X1_188/O 0.02fF
C11678 POR2X1_150/Y POR2X1_283/A 18.41fF
C11679 POR2X1_691/CTRL2 POR2X1_811/A 0.00fF
C11680 POR2X1_794/B VDD 0.50fF
C11681 POR2X1_311/Y POR2X1_79/Y 0.03fF
C11682 PAND2X1_65/B POR2X1_543/A 0.00fF
C11683 POR2X1_68/A POR2X1_567/B 0.09fF
C11684 POR2X1_528/Y POR2X1_20/B 0.07fF
C11685 POR2X1_480/A PAND2X1_41/B 0.07fF
C11686 PAND2X1_309/CTRL PAND2X1_58/A 0.01fF
C11687 POR2X1_356/A PAND2X1_20/A 0.05fF
C11688 POR2X1_96/A PAND2X1_76/a_16_344# 0.02fF
C11689 PAND2X1_787/Y POR2X1_106/Y 0.52fF
C11690 POR2X1_196/Y PAND2X1_93/B 0.06fF
C11691 POR2X1_270/a_16_28# POR2X1_445/A -0.01fF
C11692 PAND2X1_463/O PAND2X1_459/Y 0.02fF
C11693 POR2X1_557/A POR2X1_78/Y 1.50fF
C11694 POR2X1_417/Y POR2X1_46/Y 0.03fF
C11695 POR2X1_71/Y PAND2X1_575/B 0.01fF
C11696 POR2X1_78/B PAND2X1_597/O 0.01fF
C11697 PAND2X1_39/B POR2X1_569/A 0.07fF
C11698 POR2X1_427/CTRL PAND2X1_565/A 0.00fF
C11699 PAND2X1_659/B PAND2X1_474/A 0.04fF
C11700 POR2X1_146/O POR2X1_257/A 0.01fF
C11701 POR2X1_847/B VDD 0.25fF
C11702 PAND2X1_6/A PAND2X1_381/Y 0.04fF
C11703 POR2X1_196/O POR2X1_741/Y 0.02fF
C11704 PAND2X1_412/O POR2X1_546/A 0.10fF
C11705 PAND2X1_833/a_16_344# POR2X1_376/B 0.03fF
C11706 PAND2X1_658/A POR2X1_83/B 0.03fF
C11707 POR2X1_329/A PAND2X1_716/B 0.03fF
C11708 D_INPUT_0 POR2X1_550/CTRL2 0.01fF
C11709 PAND2X1_76/Y VDD 0.42fF
C11710 PAND2X1_95/B POR2X1_634/A 0.05fF
C11711 POR2X1_61/Y POR2X1_215/O 0.05fF
C11712 D_INPUT_0 POR2X1_644/A 0.13fF
C11713 INPUT_2 POR2X1_609/Y 0.01fF
C11714 POR2X1_220/Y PAND2X1_52/Y 0.03fF
C11715 POR2X1_811/A POR2X1_644/A 0.40fF
C11716 PAND2X1_787/Y PAND2X1_580/B 0.03fF
C11717 POR2X1_423/Y POR2X1_7/B 0.03fF
C11718 PAND2X1_852/A PAND2X1_656/A 0.03fF
C11719 POR2X1_48/A PAND2X1_213/Y 0.03fF
C11720 PAND2X1_6/Y POR2X1_241/B 0.03fF
C11721 POR2X1_260/Y POR2X1_330/Y 0.03fF
C11722 POR2X1_457/B POR2X1_370/Y 0.02fF
C11723 PAND2X1_478/B PAND2X1_478/O 0.11fF
C11724 POR2X1_68/A POR2X1_806/O 0.27fF
C11725 POR2X1_66/A POR2X1_318/A 0.07fF
C11726 POR2X1_63/a_16_28# POR2X1_32/A 0.03fF
C11727 POR2X1_67/Y POR2X1_4/Y 0.03fF
C11728 POR2X1_41/B PAND2X1_803/A 0.03fF
C11729 POR2X1_356/A POR2X1_814/B 0.10fF
C11730 PAND2X1_96/B PAND2X1_39/CTRL2 0.01fF
C11731 PAND2X1_814/O POR2X1_669/B 0.04fF
C11732 POR2X1_741/Y POR2X1_794/B 0.03fF
C11733 PAND2X1_90/A PAND2X1_41/B 0.16fF
C11734 PAND2X1_20/A POR2X1_78/CTRL 0.01fF
C11735 PAND2X1_108/O VDD 0.00fF
C11736 POR2X1_590/A POR2X1_550/CTRL 0.01fF
C11737 POR2X1_300/O PAND2X1_217/B 0.10fF
C11738 POR2X1_866/A POR2X1_101/Y 0.02fF
C11739 POR2X1_252/CTRL POR2X1_5/Y 0.00fF
C11740 POR2X1_567/B PAND2X1_315/CTRL2 0.16fF
C11741 POR2X1_750/B POR2X1_756/a_16_28# 0.03fF
C11742 PAND2X1_23/Y PAND2X1_395/CTRL2 0.00fF
C11743 POR2X1_102/Y PAND2X1_575/CTRL2 0.01fF
C11744 POR2X1_763/O POR2X1_46/Y 0.01fF
C11745 PAND2X1_798/B POR2X1_72/B 0.03fF
C11746 PAND2X1_208/CTRL POR2X1_599/A 0.01fF
C11747 POR2X1_83/B POR2X1_73/Y 0.20fF
C11748 POR2X1_355/O PAND2X1_23/Y 0.01fF
C11749 POR2X1_263/Y POR2X1_7/A 0.07fF
C11750 POR2X1_121/A POR2X1_188/A 0.03fF
C11751 POR2X1_683/Y POR2X1_40/Y 0.01fF
C11752 PAND2X1_95/B PAND2X1_588/CTRL2 0.01fF
C11753 PAND2X1_41/B POR2X1_350/CTRL 0.03fF
C11754 POR2X1_632/B PAND2X1_88/Y 0.00fF
C11755 POR2X1_834/Y POR2X1_260/B 0.01fF
C11756 PAND2X1_863/B VDD 0.00fF
C11757 PAND2X1_824/B POR2X1_240/O 0.01fF
C11758 POR2X1_306/O POR2X1_102/Y 0.01fF
C11759 PAND2X1_836/a_16_344# PAND2X1_403/B 0.02fF
C11760 POR2X1_257/A PAND2X1_162/A 0.00fF
C11761 POR2X1_630/A PAND2X1_69/A 0.01fF
C11762 POR2X1_32/A PAND2X1_350/O 0.08fF
C11763 POR2X1_669/CTRL VDD 0.00fF
C11764 POR2X1_52/A PAND2X1_84/Y 0.05fF
C11765 INPUT_1 POR2X1_422/O 0.01fF
C11766 POR2X1_832/B PAND2X1_589/O 0.03fF
C11767 PAND2X1_859/A PAND2X1_6/A 0.03fF
C11768 POR2X1_794/B PAND2X1_32/B 0.02fF
C11769 POR2X1_270/Y POR2X1_703/A 0.07fF
C11770 PAND2X1_65/B POR2X1_205/CTRL2 0.00fF
C11771 PAND2X1_808/Y PAND2X1_768/Y 0.00fF
C11772 POR2X1_189/m4_208_n4# PAND2X1_480/B 0.04fF
C11773 POR2X1_41/B PAND2X1_673/Y 0.00fF
C11774 PAND2X1_661/CTRL POR2X1_13/A 0.01fF
C11775 POR2X1_355/B POR2X1_502/A 0.03fF
C11776 POR2X1_221/O POR2X1_221/Y 0.01fF
C11777 PAND2X1_191/O VDD -0.00fF
C11778 POR2X1_290/CTRL PAND2X1_642/B 0.01fF
C11779 POR2X1_273/O POR2X1_153/Y 0.23fF
C11780 POR2X1_56/B INPUT_0 0.10fF
C11781 PAND2X1_793/Y POR2X1_13/A 0.03fF
C11782 POR2X1_335/A POR2X1_362/B 0.01fF
C11783 POR2X1_416/B POR2X1_827/O 0.03fF
C11784 POR2X1_61/CTRL POR2X1_66/A 0.01fF
C11785 PAND2X1_287/CTRL VDD -0.00fF
C11786 POR2X1_300/CTRL POR2X1_272/Y 0.01fF
C11787 PAND2X1_35/Y POR2X1_46/Y 0.03fF
C11788 PAND2X1_48/B PAND2X1_48/CTRL 0.00fF
C11789 POR2X1_43/B POR2X1_5/Y 0.25fF
C11790 PAND2X1_6/Y POR2X1_774/Y 0.01fF
C11791 POR2X1_49/Y POR2X1_528/a_16_28# 0.07fF
C11792 POR2X1_614/A PAND2X1_262/O 0.07fF
C11793 POR2X1_178/O PAND2X1_562/B 0.05fF
C11794 VDD PAND2X1_178/O 0.00fF
C11795 POR2X1_149/B PAND2X1_90/Y 0.59fF
C11796 POR2X1_809/A POR2X1_676/a_56_344# 0.00fF
C11797 PAND2X1_567/O VDD 0.00fF
C11798 POR2X1_141/Y POR2X1_724/A 0.06fF
C11799 PAND2X1_58/A PAND2X1_63/B 0.03fF
C11800 POR2X1_753/Y POR2X1_754/CTRL2 0.09fF
C11801 POR2X1_96/A PAND2X1_215/B 0.02fF
C11802 POR2X1_614/A POR2X1_5/Y 0.09fF
C11803 PAND2X1_96/B POR2X1_274/Y 0.03fF
C11804 POR2X1_566/A POR2X1_562/CTRL2 0.16fF
C11805 POR2X1_635/B POR2X1_451/A 0.01fF
C11806 POR2X1_78/B POR2X1_68/A 0.18fF
C11807 PAND2X1_20/A POR2X1_569/A 0.88fF
C11808 POR2X1_83/B PAND2X1_244/B 0.01fF
C11809 POR2X1_119/Y POR2X1_299/a_16_28# 0.09fF
C11810 POR2X1_280/Y PAND2X1_542/O 0.09fF
C11811 POR2X1_283/Y PAND2X1_854/A 0.02fF
C11812 PAND2X1_262/O POR2X1_38/B 0.04fF
C11813 PAND2X1_736/A PAND2X1_735/Y 0.00fF
C11814 PAND2X1_804/A PAND2X1_794/B 0.01fF
C11815 POR2X1_855/B POR2X1_783/CTRL2 0.01fF
C11816 POR2X1_638/B VDD 0.10fF
C11817 POR2X1_652/O POR2X1_480/A 0.03fF
C11818 PAND2X1_481/O POR2X1_294/Y -0.00fF
C11819 PAND2X1_566/Y VDD 2.23fF
C11820 POR2X1_256/CTRL2 POR2X1_255/Y 0.01fF
C11821 POR2X1_97/CTRL PAND2X1_20/A 0.01fF
C11822 POR2X1_38/B POR2X1_5/Y 2.34fF
C11823 PAND2X1_63/Y POR2X1_786/O 0.01fF
C11824 POR2X1_376/B POR2X1_9/CTRL2 0.01fF
C11825 PAND2X1_65/B PAND2X1_26/CTRL 0.01fF
C11826 POR2X1_58/Y POR2X1_55/Y 0.05fF
C11827 POR2X1_215/O POR2X1_35/Y 0.01fF
C11828 POR2X1_50/O INPUT_6 0.01fF
C11829 POR2X1_40/Y POR2X1_384/O 0.02fF
C11830 POR2X1_343/Y POR2X1_554/B 0.03fF
C11831 POR2X1_495/Y POR2X1_293/Y 0.06fF
C11832 POR2X1_661/B POR2X1_740/Y 0.00fF
C11833 POR2X1_22/A INPUT_5 0.02fF
C11834 POR2X1_402/O PAND2X1_60/B 0.01fF
C11835 POR2X1_184/Y POR2X1_46/Y 0.05fF
C11836 POR2X1_570/B VDD 0.23fF
C11837 POR2X1_96/A PAND2X1_6/A 0.04fF
C11838 PAND2X1_239/CTRL2 POR2X1_191/Y 0.11fF
C11839 PAND2X1_239/O POR2X1_192/B 0.14fF
C11840 POR2X1_383/A POR2X1_286/Y 0.01fF
C11841 POR2X1_49/Y POR2X1_146/O 0.06fF
C11842 PAND2X1_525/O POR2X1_550/Y 0.18fF
C11843 PAND2X1_564/B PAND2X1_569/a_16_344# 0.05fF
C11844 INPUT_1 POR2X1_748/A 0.03fF
C11845 POR2X1_120/CTRL2 PAND2X1_60/B 0.01fF
C11846 POR2X1_814/B POR2X1_569/A 0.10fF
C11847 POR2X1_218/Y POR2X1_294/A 1.75fF
C11848 PAND2X1_714/Y POR2X1_40/Y 0.08fF
C11849 PAND2X1_651/Y POR2X1_46/Y 0.00fF
C11850 POR2X1_123/B VDD 0.00fF
C11851 PAND2X1_613/m4_208_n4# POR2X1_4/Y 0.05fF
C11852 POR2X1_578/Y POR2X1_775/CTRL 0.00fF
C11853 POR2X1_800/A PAND2X1_599/CTRL 0.00fF
C11854 POR2X1_777/B POR2X1_362/A 0.03fF
C11855 POR2X1_81/CTRL2 PAND2X1_573/B 0.01fF
C11856 PAND2X1_787/Y PAND2X1_349/A 0.05fF
C11857 D_INPUT_0 POR2X1_512/O 0.01fF
C11858 PAND2X1_824/B POR2X1_630/A 0.09fF
C11859 POR2X1_346/B PAND2X1_41/B 0.01fF
C11860 POR2X1_52/A POR2X1_239/CTRL 0.01fF
C11861 POR2X1_52/A POR2X1_594/A 0.73fF
C11862 POR2X1_327/Y POR2X1_830/CTRL2 0.02fF
C11863 POR2X1_39/Y POR2X1_40/Y 0.01fF
C11864 POR2X1_48/A PAND2X1_346/CTRL2 0.01fF
C11865 POR2X1_260/B POR2X1_383/Y 3.30fF
C11866 POR2X1_220/Y POR2X1_724/A 0.07fF
C11867 POR2X1_391/A POR2X1_391/B 0.06fF
C11868 POR2X1_78/B PAND2X1_315/CTRL2 0.05fF
C11869 POR2X1_360/A POR2X1_68/B 0.07fF
C11870 POR2X1_20/CTRL POR2X1_38/B 0.00fF
C11871 PAND2X1_865/Y POR2X1_487/CTRL2 0.00fF
C11872 POR2X1_325/A POR2X1_569/A 0.14fF
C11873 POR2X1_102/CTRL POR2X1_37/Y 0.01fF
C11874 POR2X1_362/B POR2X1_249/Y 0.03fF
C11875 POR2X1_38/Y PAND2X1_598/a_76_28# 0.01fF
C11876 PAND2X1_212/CTRL2 POR2X1_77/Y 0.01fF
C11877 POR2X1_409/O POR2X1_55/Y 0.18fF
C11878 PAND2X1_649/A PAND2X1_400/CTRL 0.01fF
C11879 PAND2X1_36/a_76_28# PAND2X1_18/B 0.02fF
C11880 PAND2X1_655/Y POR2X1_689/Y 0.07fF
C11881 POR2X1_106/Y PAND2X1_114/O 0.02fF
C11882 PAND2X1_572/CTRL PAND2X1_364/B 0.07fF
C11883 POR2X1_113/Y POR2X1_114/Y 0.02fF
C11884 POR2X1_654/CTRL2 POR2X1_774/A 0.12fF
C11885 PAND2X1_94/A PAND2X1_85/Y 0.74fF
C11886 POR2X1_86/Y PAND2X1_206/A 0.03fF
C11887 POR2X1_311/Y PAND2X1_730/A 1.20fF
C11888 PAND2X1_39/B PAND2X1_72/A 0.06fF
C11889 POR2X1_315/Y VDD 0.10fF
C11890 POR2X1_567/B POR2X1_169/A 0.05fF
C11891 D_INPUT_7 PAND2X1_11/O 0.15fF
C11892 POR2X1_751/O POR2X1_7/B 0.01fF
C11893 PAND2X1_137/Y PAND2X1_348/Y 0.02fF
C11894 PAND2X1_823/CTRL2 VDD 0.00fF
C11895 POR2X1_865/B POR2X1_717/Y 0.03fF
C11896 PAND2X1_56/Y PAND2X1_69/A 0.11fF
C11897 PAND2X1_803/A PAND2X1_308/Y 0.03fF
C11898 PAND2X1_486/a_16_344# POR2X1_526/Y 0.01fF
C11899 POR2X1_334/B PAND2X1_79/Y 0.03fF
C11900 POR2X1_55/Y POR2X1_9/CTRL 0.30fF
C11901 POR2X1_65/A POR2X1_394/A 10.79fF
C11902 PAND2X1_672/CTRL POR2X1_35/B 0.01fF
C11903 POR2X1_602/B POR2X1_722/CTRL 0.01fF
C11904 POR2X1_532/A POR2X1_713/CTRL2 0.02fF
C11905 INPUT_0 PAND2X1_537/CTRL 0.01fF
C11906 POR2X1_96/A POR2X1_419/CTRL2 0.03fF
C11907 POR2X1_856/B POR2X1_711/Y 0.10fF
C11908 POR2X1_394/A PAND2X1_558/CTRL 0.07fF
C11909 PAND2X1_215/B POR2X1_7/A 2.58fF
C11910 POR2X1_514/CTRL2 POR2X1_137/Y 0.01fF
C11911 POR2X1_693/O PAND2X1_550/B 0.01fF
C11912 POR2X1_303/CTRL POR2X1_330/Y 0.31fF
C11913 PAND2X1_793/Y PAND2X1_510/B 0.00fF
C11914 POR2X1_158/Y POR2X1_23/Y 0.00fF
C11915 POR2X1_416/B POR2X1_48/A 4.69fF
C11916 PAND2X1_111/B PAND2X1_111/CTRL2 0.01fF
C11917 PAND2X1_490/CTRL2 POR2X1_38/B 0.00fF
C11918 POR2X1_68/B PAND2X1_19/CTRL 0.01fF
C11919 POR2X1_222/Y POR2X1_318/A 0.07fF
C11920 PAND2X1_401/O POR2X1_395/Y 0.00fF
C11921 PAND2X1_506/O POR2X1_239/Y 0.02fF
C11922 PAND2X1_242/O PAND2X1_241/Y 0.00fF
C11923 PAND2X1_48/O POR2X1_260/A 0.04fF
C11924 POR2X1_108/Y PAND2X1_553/B 0.11fF
C11925 PAND2X1_615/CTRL2 D_INPUT_1 0.03fF
C11926 POR2X1_541/CTRL2 POR2X1_702/A 0.00fF
C11927 VDD POR2X1_741/B 0.01fF
C11928 POR2X1_807/A PAND2X1_48/A 0.10fF
C11929 POR2X1_570/B PAND2X1_32/B 0.09fF
C11930 POR2X1_724/CTRL POR2X1_703/Y 0.01fF
C11931 POR2X1_119/Y PAND2X1_211/A 0.02fF
C11932 PAND2X1_865/Y POR2X1_40/Y 0.07fF
C11933 POR2X1_336/O PAND2X1_69/A 0.01fF
C11934 POR2X1_114/Y POR2X1_260/A 0.01fF
C11935 POR2X1_523/Y POR2X1_844/a_16_28# 0.04fF
C11936 POR2X1_250/Y POR2X1_329/A 0.17fF
C11937 POR2X1_93/A POR2X1_90/Y 0.06fF
C11938 PAND2X1_90/A POR2X1_561/CTRL 0.01fF
C11939 PAND2X1_48/B POR2X1_151/CTRL 0.03fF
C11940 POR2X1_90/Y POR2X1_91/Y 0.11fF
C11941 POR2X1_377/CTRL2 PAND2X1_94/A 0.00fF
C11942 POR2X1_861/CTRL POR2X1_101/Y 0.25fF
C11943 PAND2X1_384/O VDD 0.00fF
C11944 POR2X1_205/A POR2X1_203/Y 0.01fF
C11945 PAND2X1_6/A POR2X1_7/A 1.50fF
C11946 PAND2X1_638/CTRL POR2X1_588/Y 0.01fF
C11947 POR2X1_635/B PAND2X1_762/CTRL 0.00fF
C11948 POR2X1_541/a_16_28# PAND2X1_32/B 0.02fF
C11949 VDD POR2X1_523/B 0.05fF
C11950 PAND2X1_823/a_16_344# POR2X1_857/B 0.01fF
C11951 POR2X1_274/A POR2X1_76/B 0.29fF
C11952 POR2X1_740/Y PAND2X1_368/a_16_344# 0.02fF
C11953 PAND2X1_61/Y PAND2X1_338/O 0.02fF
C11954 POR2X1_185/CTRL2 PAND2X1_94/A 0.02fF
C11955 POR2X1_834/Y PAND2X1_55/Y 0.12fF
C11956 POR2X1_170/B POR2X1_169/a_76_344# 0.01fF
C11957 PAND2X1_723/O PAND2X1_656/A 0.05fF
C11958 POR2X1_532/A POR2X1_318/A 0.02fF
C11959 POR2X1_36/B POR2X1_582/O 0.01fF
C11960 PAND2X1_593/CTRL2 POR2X1_385/Y 0.01fF
C11961 D_INPUT_3 PAND2X1_509/O 0.05fF
C11962 POR2X1_383/A POR2X1_649/CTRL2 0.01fF
C11963 PAND2X1_630/a_76_28# POR2X1_7/A 0.02fF
C11964 POR2X1_722/A POR2X1_708/B 0.03fF
C11965 POR2X1_383/A PAND2X1_69/A 0.17fF
C11966 POR2X1_241/B PAND2X1_52/B 0.03fF
C11967 PAND2X1_23/Y POR2X1_244/Y 0.09fF
C11968 PAND2X1_56/Y PAND2X1_368/a_76_28# 0.03fF
C11969 POR2X1_532/A POR2X1_713/B 0.37fF
C11970 PAND2X1_20/A POR2X1_725/O 0.01fF
C11971 POR2X1_49/Y PAND2X1_198/CTRL 0.03fF
C11972 POR2X1_416/B PAND2X1_221/a_16_344# 0.01fF
C11973 POR2X1_88/CTRL2 POR2X1_9/Y 0.01fF
C11974 PAND2X1_57/B PAND2X1_328/CTRL2 0.00fF
C11975 PAND2X1_737/CTRL VDD 0.00fF
C11976 POR2X1_16/A POR2X1_234/CTRL 0.01fF
C11977 POR2X1_128/A POR2X1_736/A 0.12fF
C11978 PAND2X1_20/A PAND2X1_72/A 1.91fF
C11979 POR2X1_741/Y POR2X1_741/B 0.02fF
C11980 POR2X1_862/CTRL POR2X1_389/Y 0.03fF
C11981 POR2X1_101/Y PAND2X1_150/CTRL2 0.11fF
C11982 POR2X1_477/A POR2X1_186/B 0.03fF
C11983 PAND2X1_477/A PAND2X1_477/B 0.00fF
C11984 POR2X1_557/A D_INPUT_1 0.07fF
C11985 PAND2X1_48/a_76_28# PAND2X1_48/A 0.01fF
C11986 PAND2X1_94/A POR2X1_78/a_56_344# 0.00fF
C11987 POR2X1_394/A PAND2X1_188/a_56_28# 0.00fF
C11988 POR2X1_119/Y POR2X1_96/A 23.62fF
C11989 POR2X1_355/B POR2X1_188/Y 0.03fF
C11990 POR2X1_68/A PAND2X1_142/CTRL2 0.03fF
C11991 PAND2X1_94/A PAND2X1_49/m4_208_n4# 0.01fF
C11992 POR2X1_328/O INPUT_5 0.18fF
C11993 PAND2X1_63/Y POR2X1_260/A 0.10fF
C11994 PAND2X1_552/B PAND2X1_703/CTRL2 0.00fF
C11995 PAND2X1_106/CTRL POR2X1_383/A 0.01fF
C11996 POR2X1_710/B PAND2X1_60/B 0.01fF
C11997 POR2X1_833/A POR2X1_576/Y 0.00fF
C11998 POR2X1_388/a_16_28# POR2X1_180/B 0.03fF
C11999 POR2X1_834/Y POR2X1_407/Y 0.01fF
C12000 POR2X1_118/CTRL2 PAND2X1_560/B 0.03fF
C12001 POR2X1_13/Y PAND2X1_538/O 0.03fF
C12002 POR2X1_38/B POR2X1_6/CTRL2 0.02fF
C12003 PAND2X1_118/a_16_344# POR2X1_559/A 0.04fF
C12004 PAND2X1_803/A POR2X1_77/Y 0.02fF
C12005 POR2X1_841/B POR2X1_458/Y 0.07fF
C12006 POR2X1_698/Y POR2X1_32/A 0.01fF
C12007 POR2X1_588/Y POR2X1_7/A 0.03fF
C12008 POR2X1_416/B PAND2X1_193/CTRL2 0.05fF
C12009 PAND2X1_94/A POR2X1_137/Y 0.05fF
C12010 PAND2X1_349/A POR2X1_103/Y 0.02fF
C12011 POR2X1_677/a_16_28# POR2X1_77/Y 0.02fF
C12012 POR2X1_65/A PAND2X1_326/CTRL 0.01fF
C12013 POR2X1_562/B POR2X1_186/B 0.03fF
C12014 PAND2X1_495/O POR2X1_260/A 0.10fF
C12015 PAND2X1_75/CTRL2 POR2X1_260/B 0.01fF
C12016 PAND2X1_850/Y PAND2X1_592/O 0.03fF
C12017 POR2X1_55/Y POR2X1_171/Y 0.02fF
C12018 POR2X1_278/Y POR2X1_680/O 0.03fF
C12019 POR2X1_774/Y PAND2X1_52/B 0.01fF
C12020 PAND2X1_23/Y POR2X1_191/Y 0.08fF
C12021 POR2X1_105/Y PAND2X1_52/B 0.02fF
C12022 POR2X1_814/B PAND2X1_72/A 0.11fF
C12023 PAND2X1_569/B POR2X1_765/Y 0.04fF
C12024 PAND2X1_288/A PAND2X1_367/a_16_344# 0.05fF
C12025 POR2X1_113/Y POR2X1_260/A 0.27fF
C12026 POR2X1_407/A PAND2X1_48/A 0.10fF
C12027 POR2X1_68/A POR2X1_294/A 0.06fF
C12028 PAND2X1_738/Y POR2X1_39/B 0.01fF
C12029 PAND2X1_628/a_16_344# POR2X1_555/B 0.05fF
C12030 POR2X1_467/a_16_28# POR2X1_452/Y 0.01fF
C12031 POR2X1_83/A POR2X1_397/O 0.01fF
C12032 POR2X1_343/Y POR2X1_723/CTRL -0.00fF
C12033 POR2X1_49/Y POR2X1_90/O 0.02fF
C12034 PAND2X1_6/Y POR2X1_593/a_16_28# 0.01fF
C12035 PAND2X1_673/Y POR2X1_77/Y 0.03fF
C12036 POR2X1_265/Y PAND2X1_734/CTRL 0.01fF
C12037 POR2X1_622/O POR2X1_29/A 0.01fF
C12038 POR2X1_73/Y PAND2X1_325/CTRL 0.01fF
C12039 POR2X1_353/A POR2X1_854/B 0.03fF
C12040 PAND2X1_675/CTRL2 PAND2X1_736/A 0.01fF
C12041 POR2X1_722/Y POR2X1_711/Y 0.22fF
C12042 PAND2X1_849/B PAND2X1_100/O 0.03fF
C12043 POR2X1_329/A PAND2X1_561/O 0.02fF
C12044 POR2X1_249/Y POR2X1_734/CTRL 0.01fF
C12045 PAND2X1_413/O POR2X1_814/A 0.02fF
C12046 PAND2X1_94/A POR2X1_833/A 1.54fF
C12047 INPUT_1 POR2X1_463/Y 0.03fF
C12048 POR2X1_110/Y POR2X1_91/Y 0.03fF
C12049 POR2X1_57/A POR2X1_518/CTRL2 0.03fF
C12050 POR2X1_513/B PAND2X1_72/A 0.03fF
C12051 POR2X1_416/B PAND2X1_197/Y 0.02fF
C12052 PAND2X1_854/A PAND2X1_365/A 0.02fF
C12053 POR2X1_413/A POR2X1_416/B 0.02fF
C12054 POR2X1_240/B POR2X1_240/A 0.12fF
C12055 POR2X1_273/Y POR2X1_39/B 0.04fF
C12056 POR2X1_316/Y PAND2X1_457/O 0.04fF
C12057 POR2X1_457/Y POR2X1_750/B 0.04fF
C12058 POR2X1_327/O PAND2X1_72/A 0.02fF
C12059 POR2X1_116/A POR2X1_218/Y 0.02fF
C12060 PAND2X1_196/CTRL2 PAND2X1_199/B 0.00fF
C12061 POR2X1_132/a_76_344# PAND2X1_140/A 0.00fF
C12062 POR2X1_119/Y POR2X1_7/A 0.08fF
C12063 POR2X1_773/B POR2X1_557/B 0.05fF
C12064 PAND2X1_440/O PAND2X1_798/B 0.06fF
C12065 POR2X1_56/Y PAND2X1_840/Y 0.00fF
C12066 POR2X1_564/B POR2X1_456/B 0.94fF
C12067 POR2X1_121/a_16_28# POR2X1_537/Y 0.01fF
C12068 POR2X1_119/Y PAND2X1_344/a_76_28# 0.01fF
C12069 POR2X1_274/A POR2X1_301/A 0.56fF
C12070 POR2X1_66/Y POR2X1_294/Y 0.00fF
C12071 POR2X1_539/CTRL2 POR2X1_567/A 0.01fF
C12072 POR2X1_707/O PAND2X1_48/A 0.02fF
C12073 POR2X1_343/Y POR2X1_702/A 0.05fF
C12074 PAND2X1_479/CTRL2 POR2X1_329/A 0.01fF
C12075 POR2X1_329/A PAND2X1_205/Y 0.11fF
C12076 POR2X1_814/A POR2X1_543/A 0.59fF
C12077 POR2X1_467/CTRL PAND2X1_52/B 0.01fF
C12078 POR2X1_496/Y POR2X1_628/Y 0.02fF
C12079 PAND2X1_301/O PAND2X1_716/B 0.06fF
C12080 POR2X1_23/Y POR2X1_265/O 0.01fF
C12081 POR2X1_20/B POR2X1_667/A 0.01fF
C12082 PAND2X1_860/A POR2X1_293/Y 0.03fF
C12083 POR2X1_607/A POR2X1_20/B 0.06fF
C12084 POR2X1_644/O POR2X1_644/B 0.00fF
C12085 POR2X1_129/Y PAND2X1_156/A 0.03fF
C12086 PAND2X1_213/Y PAND2X1_169/a_56_28# 0.00fF
C12087 PAND2X1_425/Y PAND2X1_582/CTRL2 0.01fF
C12088 POR2X1_495/Y PAND2X1_242/Y 0.16fF
C12089 POR2X1_228/Y POR2X1_716/CTRL 0.01fF
C12090 POR2X1_846/A PAND2X1_57/B 0.03fF
C12091 PAND2X1_63/B POR2X1_342/B 0.05fF
C12092 POR2X1_9/Y POR2X1_618/CTRL2 0.14fF
C12093 PAND2X1_612/B POR2X1_78/A 0.03fF
C12094 PAND2X1_458/CTRL POR2X1_372/Y 0.01fF
C12095 POR2X1_11/O INPUT_7 0.01fF
C12096 PAND2X1_439/O PAND2X1_738/Y 0.08fF
C12097 POR2X1_520/a_16_28# POR2X1_383/Y 0.01fF
C12098 POR2X1_379/CTRL2 PAND2X1_52/B 0.15fF
C12099 POR2X1_106/O POR2X1_48/A 0.03fF
C12100 POR2X1_16/A PAND2X1_440/CTRL 0.06fF
C12101 POR2X1_685/A PAND2X1_681/O 0.02fF
C12102 POR2X1_420/CTRL POR2X1_102/Y 0.01fF
C12103 POR2X1_754/Y POR2X1_67/A 0.01fF
C12104 POR2X1_411/B POR2X1_236/Y 7.15fF
C12105 PAND2X1_613/CTRL PAND2X1_41/B 0.01fF
C12106 POR2X1_681/Y POR2X1_682/CTRL2 0.01fF
C12107 POR2X1_705/B PAND2X1_57/B 0.19fF
C12108 POR2X1_12/A POR2X1_763/A 0.48fF
C12109 PAND2X1_93/B POR2X1_141/Y 0.03fF
C12110 POR2X1_11/O INPUT_4 0.02fF
C12111 POR2X1_604/Y POR2X1_669/B 0.10fF
C12112 POR2X1_52/CTRL2 POR2X1_7/Y 0.01fF
C12113 POR2X1_760/A PAND2X1_215/B 0.07fF
C12114 POR2X1_636/B POR2X1_750/B 0.81fF
C12115 POR2X1_261/Y VDD 0.01fF
C12116 POR2X1_554/B POR2X1_276/CTRL2 0.03fF
C12117 PAND2X1_827/O POR2X1_355/A 0.02fF
C12118 PAND2X1_96/B POR2X1_837/A 0.01fF
C12119 POR2X1_278/Y POR2X1_63/Y 0.05fF
C12120 PAND2X1_571/A PAND2X1_576/CTRL2 0.01fF
C12121 PAND2X1_434/a_16_344# PAND2X1_390/Y 0.01fF
C12122 POR2X1_417/Y PAND2X1_352/A 0.91fF
C12123 POR2X1_24/CTRL POR2X1_409/B 0.04fF
C12124 POR2X1_847/B POR2X1_818/Y 0.02fF
C12125 POR2X1_257/A PAND2X1_735/Y 0.09fF
C12126 POR2X1_78/B PAND2X1_601/O 0.31fF
C12127 PAND2X1_689/a_76_28# POR2X1_121/B 0.03fF
C12128 PAND2X1_486/O POR2X1_484/Y 0.02fF
C12129 POR2X1_67/Y POR2X1_816/A 7.48fF
C12130 POR2X1_446/B POR2X1_724/CTRL2 0.01fF
C12131 POR2X1_754/Y POR2X1_615/CTRL2 0.02fF
C12132 POR2X1_35/B POR2X1_34/A 0.00fF
C12133 POR2X1_67/Y D_INPUT_1 0.18fF
C12134 POR2X1_150/Y POR2X1_55/Y 0.17fF
C12135 POR2X1_809/A PAND2X1_681/CTRL2 0.01fF
C12136 POR2X1_130/A POR2X1_655/A 0.05fF
C12137 PAND2X1_622/a_16_344# POR2X1_48/A 0.02fF
C12138 POR2X1_753/Y POR2X1_752/Y 0.01fF
C12139 POR2X1_259/A POR2X1_555/B 0.01fF
C12140 POR2X1_332/Y PAND2X1_72/A 0.01fF
C12141 PAND2X1_268/CTRL POR2X1_193/A 0.08fF
C12142 PAND2X1_423/CTRL2 POR2X1_78/A 0.01fF
C12143 POR2X1_654/B POR2X1_590/A 0.10fF
C12144 POR2X1_671/CTRL2 POR2X1_37/Y 0.01fF
C12145 PAND2X1_420/O POR2X1_630/A 0.05fF
C12146 POR2X1_65/A POR2X1_669/B 0.15fF
C12147 PAND2X1_793/Y POR2X1_67/CTRL2 0.01fF
C12148 POR2X1_57/A POR2X1_250/Y 0.02fF
C12149 POR2X1_68/A POR2X1_116/A 0.05fF
C12150 POR2X1_55/CTRL2 POR2X1_5/Y 0.03fF
C12151 PAND2X1_633/O POR2X1_32/A 0.04fF
C12152 PAND2X1_220/Y POR2X1_487/a_16_28# 0.04fF
C12153 PAND2X1_58/A POR2X1_391/A 0.03fF
C12154 PAND2X1_793/Y POR2X1_437/O 0.01fF
C12155 POR2X1_20/B PAND2X1_546/CTRL2 0.03fF
C12156 POR2X1_442/Y PAND2X1_211/A 0.02fF
C12157 POR2X1_20/B PAND2X1_182/CTRL2 0.00fF
C12158 PAND2X1_93/B POR2X1_220/Y 0.10fF
C12159 PAND2X1_73/Y POR2X1_455/CTRL2 0.01fF
C12160 POR2X1_48/A PAND2X1_738/Y 0.06fF
C12161 D_INPUT_0 PAND2X1_8/Y 0.14fF
C12162 POR2X1_411/B POR2X1_232/Y 0.00fF
C12163 POR2X1_538/A POR2X1_814/A 0.01fF
C12164 PAND2X1_810/a_76_28# PAND2X1_221/Y 0.02fF
C12165 PAND2X1_11/Y PAND2X1_18/O 0.00fF
C12166 PAND2X1_93/B POR2X1_404/Y 0.06fF
C12167 POR2X1_138/CTRL POR2X1_260/B 0.01fF
C12168 POR2X1_368/a_16_28# POR2X1_23/Y 0.06fF
C12169 POR2X1_342/B POR2X1_342/A 0.04fF
C12170 POR2X1_210/O VDD 0.00fF
C12171 POR2X1_23/Y PAND2X1_592/Y 0.03fF
C12172 PAND2X1_838/O POR2X1_73/Y 0.05fF
C12173 POR2X1_624/Y POR2X1_501/a_16_28# 0.02fF
C12174 POR2X1_335/B POR2X1_556/A 0.03fF
C12175 PAND2X1_338/a_76_28# PAND2X1_333/Y 0.02fF
C12176 PAND2X1_272/O PAND2X1_57/B 0.08fF
C12177 POR2X1_247/Y INPUT_0 0.00fF
C12178 POR2X1_78/B PAND2X1_58/A 0.08fF
C12179 PAND2X1_776/Y PAND2X1_776/O 0.01fF
C12180 PAND2X1_615/CTRL2 INPUT_3 0.04fF
C12181 PAND2X1_611/CTRL2 POR2X1_249/Y 0.01fF
C12182 POR2X1_624/Y POR2X1_702/A 0.08fF
C12183 PAND2X1_78/CTRL2 PAND2X1_580/B 0.00fF
C12184 PAND2X1_429/CTRL2 INPUT_5 0.03fF
C12185 POR2X1_78/A POR2X1_220/Y 0.06fF
C12186 PAND2X1_721/B PAND2X1_734/B 0.01fF
C12187 PAND2X1_793/Y POR2X1_29/A 0.04fF
C12188 POR2X1_177/Y POR2X1_72/B 0.02fF
C12189 POR2X1_686/A POR2X1_828/Y 0.14fF
C12190 POR2X1_13/A POR2X1_516/Y 0.03fF
C12191 POR2X1_812/CTRL POR2X1_121/B 0.04fF
C12192 PAND2X1_206/A POR2X1_73/Y 0.05fF
C12193 POR2X1_814/A POR2X1_768/CTRL 0.01fF
C12194 POR2X1_489/B PAND2X1_57/B 0.01fF
C12195 POR2X1_14/Y POR2X1_668/Y 0.03fF
C12196 POR2X1_20/B POR2X1_245/Y 0.10fF
C12197 PAND2X1_48/B POR2X1_269/CTRL 0.01fF
C12198 POR2X1_861/CTRL2 POR2X1_218/Y 0.09fF
C12199 PAND2X1_613/CTRL2 POR2X1_68/B 0.01fF
C12200 POR2X1_123/A POR2X1_556/A 0.04fF
C12201 POR2X1_179/Y POR2X1_150/Y 0.02fF
C12202 PAND2X1_474/A POR2X1_5/Y 0.23fF
C12203 PAND2X1_459/O VDD 0.00fF
C12204 POR2X1_472/CTRL2 POR2X1_472/B 0.03fF
C12205 POR2X1_78/A POR2X1_404/Y 0.00fF
C12206 POR2X1_66/A POR2X1_341/O 0.01fF
C12207 PAND2X1_217/O PAND2X1_656/A 0.02fF
C12208 PAND2X1_558/Y VDD 0.04fF
C12209 POR2X1_67/A POR2X1_42/Y 0.10fF
C12210 POR2X1_56/B POR2X1_102/Y 0.17fF
C12211 POR2X1_78/A PAND2X1_322/a_76_28# 0.00fF
C12212 POR2X1_306/a_16_28# PAND2X1_454/B 0.01fF
C12213 POR2X1_376/B POR2X1_236/Y 0.38fF
C12214 PAND2X1_217/B PAND2X1_480/B 0.10fF
C12215 POR2X1_853/A POR2X1_174/A 0.03fF
C12216 POR2X1_302/B PAND2X1_322/CTRL2 0.01fF
C12217 PAND2X1_787/O VDD 0.00fF
C12218 POR2X1_356/A POR2X1_209/a_16_28# 0.02fF
C12219 POR2X1_659/A POR2X1_510/Y 0.03fF
C12220 POR2X1_567/B PAND2X1_96/B 0.05fF
C12221 POR2X1_400/A POR2X1_61/Y 0.03fF
C12222 POR2X1_226/O POR2X1_42/Y 0.08fF
C12223 PAND2X1_84/O POR2X1_5/Y 0.17fF
C12224 POR2X1_257/A PAND2X1_569/B 0.07fF
C12225 POR2X1_257/A POR2X1_158/B 0.04fF
C12226 POR2X1_495/Y POR2X1_60/A 0.06fF
C12227 POR2X1_253/Y POR2X1_496/Y 0.14fF
C12228 POR2X1_66/A POR2X1_194/CTRL 0.01fF
C12229 PAND2X1_90/A PAND2X1_73/CTRL 0.01fF
C12230 PAND2X1_244/B PAND2X1_206/A 0.03fF
C12231 POR2X1_130/A PAND2X1_589/O -0.00fF
C12232 POR2X1_263/Y POR2X1_38/Y 0.05fF
C12233 POR2X1_78/B POR2X1_457/B 0.01fF
C12234 POR2X1_814/A POR2X1_342/O 0.02fF
C12235 POR2X1_278/Y PAND2X1_768/Y 0.02fF
C12236 PAND2X1_48/B POR2X1_602/B 0.02fF
C12237 POR2X1_590/A POR2X1_705/CTRL 0.01fF
C12238 PAND2X1_224/m4_208_n4# POR2X1_192/B 0.02fF
C12239 POR2X1_76/a_16_28# POR2X1_274/B 0.02fF
C12240 POR2X1_493/O POR2X1_558/B 0.00fF
C12241 PAND2X1_23/Y POR2X1_242/O 0.16fF
C12242 PAND2X1_124/Y PAND2X1_656/A 0.62fF
C12243 PAND2X1_859/a_16_344# POR2X1_13/A 0.02fF
C12244 PAND2X1_467/Y PAND2X1_452/CTRL 0.01fF
C12245 POR2X1_610/Y POR2X1_260/A 0.03fF
C12246 D_INPUT_3 POR2X1_409/B 0.10fF
C12247 POR2X1_121/m4_208_n4# POR2X1_655/A 0.01fF
C12248 PAND2X1_350/A POR2X1_5/Y 0.00fF
C12249 POR2X1_743/CTRL2 POR2X1_7/B 0.03fF
C12250 POR2X1_238/a_16_28# POR2X1_236/Y 0.03fF
C12251 POR2X1_136/Y POR2X1_48/A 0.03fF
C12252 POR2X1_475/m4_208_n4# POR2X1_101/Y 0.02fF
C12253 POR2X1_41/B PAND2X1_833/CTRL2 0.05fF
C12254 POR2X1_49/Y PAND2X1_859/B 0.01fF
C12255 PAND2X1_6/Y POR2X1_457/CTRL2 0.01fF
C12256 POR2X1_271/A POR2X1_411/B 0.23fF
C12257 POR2X1_72/B PAND2X1_552/B 0.42fF
C12258 POR2X1_777/B POR2X1_572/B 0.03fF
C12259 POR2X1_78/B POR2X1_435/Y 0.07fF
C12260 PAND2X1_78/O PAND2X1_794/B 0.04fF
C12261 PAND2X1_16/O POR2X1_294/B 0.09fF
C12262 PAND2X1_341/B POR2X1_65/O 0.01fF
C12263 PAND2X1_860/A PAND2X1_862/CTRL2 0.01fF
C12264 PAND2X1_390/Y PAND2X1_658/B 0.05fF
C12265 POR2X1_555/B PAND2X1_88/Y 0.02fF
C12266 POR2X1_573/CTRL POR2X1_404/Y 0.00fF
C12267 POR2X1_366/CTRL PAND2X1_93/B 0.01fF
C12268 POR2X1_68/B PAND2X1_531/O 0.02fF
C12269 PAND2X1_480/B VDD 3.50fF
C12270 PAND2X1_558/CTRL2 PAND2X1_493/Y 0.01fF
C12271 POR2X1_57/A POR2X1_279/O 0.01fF
C12272 PAND2X1_65/B POR2X1_193/A 0.03fF
C12273 PAND2X1_25/O INPUT_6 0.17fF
C12274 PAND2X1_65/B POR2X1_579/Y 0.03fF
C12275 POR2X1_614/A PAND2X1_582/CTRL2 0.00fF
C12276 PAND2X1_93/B POR2X1_215/A 0.13fF
C12277 POR2X1_68/A POR2X1_94/A 0.14fF
C12278 POR2X1_862/B PAND2X1_536/CTRL 0.00fF
C12279 PAND2X1_48/B POR2X1_213/B 0.03fF
C12280 POR2X1_52/A POR2X1_236/Y 5.54fF
C12281 PAND2X1_225/O D_INPUT_1 0.16fF
C12282 POR2X1_274/CTRL POR2X1_569/A 0.03fF
C12283 PAND2X1_394/CTRL PAND2X1_88/Y 0.01fF
C12284 PAND2X1_785/Y PAND2X1_795/B 0.01fF
C12285 POR2X1_254/A POR2X1_341/a_16_28# 0.02fF
C12286 PAND2X1_73/Y PAND2X1_60/B 0.21fF
C12287 PAND2X1_65/B POR2X1_572/B 0.03fF
C12288 POR2X1_614/A POR2X1_777/B 0.10fF
C12289 POR2X1_509/B POR2X1_340/a_16_28# 0.02fF
C12290 PAND2X1_63/Y PAND2X1_265/m4_208_n4# 0.03fF
C12291 PAND2X1_242/CTRL2 POR2X1_511/Y 0.03fF
C12292 POR2X1_96/A POR2X1_693/CTRL2 0.00fF
C12293 POR2X1_29/CTRL POR2X1_55/Y 0.01fF
C12294 POR2X1_356/A VDD 8.80fF
C12295 POR2X1_13/CTRL POR2X1_7/B 0.01fF
C12296 POR2X1_855/A POR2X1_803/A 0.44fF
C12297 PAND2X1_317/Y POR2X1_236/Y 0.11fF
C12298 POR2X1_814/B POR2X1_793/A 0.06fF
C12299 POR2X1_152/A POR2X1_236/Y 0.03fF
C12300 POR2X1_213/O POR2X1_213/B 0.00fF
C12301 PAND2X1_805/A PAND2X1_567/a_76_28# 0.01fF
C12302 PAND2X1_553/A POR2X1_55/Y 0.00fF
C12303 POR2X1_83/B PAND2X1_656/A 0.03fF
C12304 POR2X1_330/Y PAND2X1_88/Y 0.03fF
C12305 POR2X1_537/Y PAND2X1_39/B 0.03fF
C12306 POR2X1_631/A POR2X1_200/CTRL 0.11fF
C12307 PAND2X1_659/B POR2X1_494/Y 2.45fF
C12308 POR2X1_13/A POR2X1_684/O 0.18fF
C12309 PAND2X1_377/CTRL POR2X1_42/Y 0.05fF
C12310 PAND2X1_787/Y POR2X1_184/Y 0.05fF
C12311 POR2X1_634/A PAND2X1_757/O 0.28fF
C12312 PAND2X1_23/Y POR2X1_302/Y 0.02fF
C12313 POR2X1_497/Y POR2X1_521/CTRL2 0.00fF
C12314 PAND2X1_48/B POR2X1_546/A 0.00fF
C12315 POR2X1_16/A POR2X1_609/Y 0.05fF
C12316 POR2X1_614/A PAND2X1_65/B 2.89fF
C12317 POR2X1_317/Y PAND2X1_65/B 0.01fF
C12318 POR2X1_52/A POR2X1_81/Y 0.00fF
C12319 PAND2X1_6/Y POR2X1_464/CTRL2 0.01fF
C12320 POR2X1_302/CTRL2 POR2X1_513/Y 0.01fF
C12321 PAND2X1_283/CTRL VDD -0.00fF
C12322 POR2X1_809/A POR2X1_866/A 0.05fF
C12323 POR2X1_400/A POR2X1_35/Y 0.01fF
C12324 POR2X1_57/A PAND2X1_205/Y 0.03fF
C12325 POR2X1_60/A PAND2X1_723/A 0.00fF
C12326 PAND2X1_550/a_56_28# PAND2X1_546/Y 0.00fF
C12327 POR2X1_722/Y POR2X1_733/A 0.01fF
C12328 POR2X1_70/O POR2X1_697/Y 0.02fF
C12329 POR2X1_41/B PAND2X1_35/CTRL2 0.00fF
C12330 PAND2X1_319/B PAND2X1_220/Y 0.07fF
C12331 POR2X1_557/A POR2X1_78/A 0.06fF
C12332 PAND2X1_91/CTRL POR2X1_192/B 0.04fF
C12333 POR2X1_72/B POR2X1_530/Y 0.01fF
C12334 PAND2X1_465/B POR2X1_7/B 0.02fF
C12335 POR2X1_316/Y PAND2X1_464/O 0.04fF
C12336 POR2X1_360/A PAND2X1_90/A 0.03fF
C12337 POR2X1_263/Y POR2X1_153/Y 0.05fF
C12338 POR2X1_523/Y INPUT_0 0.05fF
C12339 PAND2X1_627/CTRL2 PAND2X1_69/A 0.00fF
C12340 POR2X1_401/A POR2X1_401/B 0.02fF
C12341 PAND2X1_42/CTRL PAND2X1_111/B 0.01fF
C12342 POR2X1_509/a_16_28# POR2X1_857/B 0.06fF
C12343 POR2X1_783/CTRL POR2X1_796/A 0.01fF
C12344 PAND2X1_258/a_16_344# POR2X1_186/B 0.00fF
C12345 PAND2X1_41/B POR2X1_319/Y 0.03fF
C12346 POR2X1_528/CTRL2 POR2X1_56/B 0.01fF
C12347 POR2X1_131/Y POR2X1_60/A 0.94fF
C12348 PAND2X1_90/Y POR2X1_209/A 0.03fF
C12349 POR2X1_78/B PAND2X1_96/B 0.43fF
C12350 POR2X1_140/B PAND2X1_516/O 0.00fF
C12351 POR2X1_254/Y POR2X1_786/Y 0.91fF
C12352 POR2X1_37/Y PAND2X1_156/A 0.03fF
C12353 POR2X1_316/Y POR2X1_257/A 0.06fF
C12354 PAND2X1_69/A INPUT_0 0.13fF
C12355 PAND2X1_52/Y POR2X1_222/A 0.02fF
C12356 POR2X1_832/Y POR2X1_512/a_16_28# 0.08fF
C12357 POR2X1_41/B PAND2X1_546/CTRL 0.01fF
C12358 POR2X1_416/B PAND2X1_634/O 0.04fF
C12359 POR2X1_260/Y POR2X1_205/CTRL2 0.00fF
C12360 POR2X1_466/A POR2X1_552/O 0.03fF
C12361 PAND2X1_341/A INPUT_0 0.02fF
C12362 POR2X1_278/Y POR2X1_498/A 0.08fF
C12363 PAND2X1_838/B POR2X1_39/B 0.01fF
C12364 POR2X1_49/Y PAND2X1_569/B 0.14fF
C12365 POR2X1_378/A POR2X1_378/a_16_28# 0.05fF
C12366 POR2X1_532/A PAND2X1_131/O 0.04fF
C12367 POR2X1_313/Y POR2X1_417/Y 0.12fF
C12368 POR2X1_51/A POR2X1_36/CTRL2 0.01fF
C12369 POR2X1_32/A PAND2X1_708/O 0.01fF
C12370 PAND2X1_476/A POR2X1_23/Y 0.05fF
C12371 POR2X1_220/A VDD 0.44fF
C12372 PAND2X1_492/CTRL PAND2X1_60/B 0.01fF
C12373 PAND2X1_461/CTRL2 POR2X1_612/Y 0.05fF
C12374 PAND2X1_48/B POR2X1_712/Y 0.03fF
C12375 POR2X1_278/Y PAND2X1_284/Y 0.10fF
C12376 INPUT_0 POR2X1_91/Y 0.07fF
C12377 POR2X1_62/Y POR2X1_623/B 0.01fF
C12378 POR2X1_237/Y PAND2X1_445/CTRL2 0.01fF
C12379 POR2X1_623/A POR2X1_5/Y 0.00fF
C12380 POR2X1_66/B POR2X1_752/m4_208_n4# 0.15fF
C12381 POR2X1_356/A PAND2X1_32/B 0.05fF
C12382 PAND2X1_303/B VDD 0.03fF
C12383 PAND2X1_94/A POR2X1_650/A 0.05fF
C12384 PAND2X1_11/Y PAND2X1_18/B 5.62fF
C12385 POR2X1_43/B PAND2X1_228/a_16_344# 0.04fF
C12386 POR2X1_439/Y POR2X1_456/B 0.02fF
C12387 POR2X1_52/A POR2X1_584/a_16_28# 0.01fF
C12388 POR2X1_119/Y PAND2X1_446/CTRL 0.02fF
C12389 POR2X1_795/CTRL PAND2X1_32/B 0.01fF
C12390 POR2X1_614/A PAND2X1_599/O 0.04fF
C12391 PAND2X1_252/CTRL PAND2X1_55/Y 0.01fF
C12392 PAND2X1_58/A POR2X1_294/A 0.10fF
C12393 PAND2X1_215/B POR2X1_38/Y 0.03fF
C12394 POR2X1_57/A PAND2X1_243/B 0.03fF
C12395 POR2X1_447/CTRL POR2X1_294/B 0.01fF
C12396 POR2X1_697/Y POR2X1_73/Y 0.00fF
C12397 POR2X1_866/A POR2X1_711/Y 0.07fF
C12398 PAND2X1_428/CTRL PAND2X1_48/A 0.30fF
C12399 POR2X1_235/Y PAND2X1_734/B 0.00fF
C12400 PAND2X1_551/A POR2X1_90/Y 0.09fF
C12401 POR2X1_383/A POR2X1_121/Y 2.07fF
C12402 D_INPUT_2 POR2X1_38/B 0.00fF
C12403 POR2X1_222/Y POR2X1_194/CTRL 0.02fF
C12404 POR2X1_503/O POR2X1_236/Y 0.02fF
C12405 PAND2X1_631/A POR2X1_83/B 0.03fF
C12406 POR2X1_396/Y POR2X1_669/a_76_344# 0.01fF
C12407 PAND2X1_63/Y POR2X1_204/O 0.01fF
C12408 POR2X1_502/A PAND2X1_373/CTRL 0.01fF
C12409 PAND2X1_470/O POR2X1_43/B 0.01fF
C12410 PAND2X1_229/O POR2X1_186/B 0.01fF
C12411 POR2X1_365/Y POR2X1_212/CTRL2 0.04fF
C12412 POR2X1_23/Y PAND2X1_327/CTRL2 0.01fF
C12413 POR2X1_390/B POR2X1_723/O 0.00fF
C12414 POR2X1_266/A PAND2X1_41/B 0.06fF
C12415 POR2X1_93/A POR2X1_618/a_16_28# 0.02fF
C12416 PAND2X1_550/CTRL2 POR2X1_394/A 0.01fF
C12417 PAND2X1_341/B POR2X1_40/Y 0.03fF
C12418 PAND2X1_144/CTRL PAND2X1_60/B 0.01fF
C12419 PAND2X1_96/B PAND2X1_767/CTRL 0.00fF
C12420 POR2X1_72/B PAND2X1_330/CTRL2 0.01fF
C12421 POR2X1_38/Y PAND2X1_6/A 0.09fF
C12422 POR2X1_122/Y POR2X1_394/A 0.07fF
C12423 PAND2X1_109/CTRL2 POR2X1_78/A 0.08fF
C12424 PAND2X1_792/m4_208_n4# POR2X1_533/m4_208_n4# 0.13fF
C12425 POR2X1_299/CTRL POR2X1_90/Y 0.01fF
C12426 PAND2X1_209/CTRL POR2X1_394/A 0.01fF
C12427 POR2X1_96/CTRL PAND2X1_472/B 0.04fF
C12428 PAND2X1_691/Y POR2X1_7/B 0.06fF
C12429 POR2X1_83/A PAND2X1_338/B 0.03fF
C12430 PAND2X1_478/Y POR2X1_119/Y 0.01fF
C12431 POR2X1_537/Y POR2X1_814/B 0.03fF
C12432 POR2X1_40/Y PAND2X1_352/Y 0.03fF
C12433 POR2X1_82/m4_208_n4# POR2X1_16/A 0.15fF
C12434 PAND2X1_784/a_16_344# POR2X1_245/Y 0.02fF
C12435 PAND2X1_216/B PAND2X1_205/B 0.01fF
C12436 POR2X1_416/B PAND2X1_34/CTRL 0.06fF
C12437 POR2X1_532/A POR2X1_219/O 0.02fF
C12438 POR2X1_569/A POR2X1_501/CTRL2 0.04fF
C12439 POR2X1_438/Y POR2X1_167/Y 0.52fF
C12440 POR2X1_25/CTRL PAND2X1_18/B 0.02fF
C12441 PAND2X1_174/a_16_344# PAND2X1_549/B 0.02fF
C12442 POR2X1_368/Y POR2X1_387/Y 0.03fF
C12443 POR2X1_239/CTRL2 POR2X1_239/Y 0.01fF
C12444 POR2X1_440/Y POR2X1_468/a_16_28# 0.11fF
C12445 POR2X1_741/Y POR2X1_569/A 0.07fF
C12446 PAND2X1_94/A POR2X1_294/B 0.26fF
C12447 POR2X1_93/O D_INPUT_3 0.03fF
C12448 POR2X1_537/Y POR2X1_733/CTRL 0.01fF
C12449 POR2X1_373/Y VDD 0.01fF
C12450 PAND2X1_358/A POR2X1_88/Y 0.01fF
C12451 POR2X1_65/A POR2X1_41/Y 0.01fF
C12452 POR2X1_514/CTRL POR2X1_101/Y 0.30fF
C12453 PAND2X1_483/O POR2X1_55/Y 0.04fF
C12454 PAND2X1_211/A PAND2X1_326/B 0.01fF
C12455 PAND2X1_84/Y PAND2X1_716/B 0.03fF
C12456 POR2X1_415/A POR2X1_9/Y 1.09fF
C12457 POR2X1_855/B POR2X1_828/A 0.03fF
C12458 POR2X1_569/A PAND2X1_32/B 0.79fF
C12459 PAND2X1_838/B POR2X1_827/O 0.01fF
C12460 PAND2X1_177/CTRL POR2X1_854/B 0.31fF
C12461 PAND2X1_863/B POR2X1_595/O 0.01fF
C12462 POR2X1_204/O POR2X1_260/A 0.01fF
C12463 POR2X1_337/A POR2X1_335/Y 0.02fF
C12464 POR2X1_57/A PAND2X1_857/A 7.24fF
C12465 POR2X1_119/Y POR2X1_609/A 0.17fF
C12466 INPUT_1 PAND2X1_6/A 3.69fF
C12467 POR2X1_208/A PAND2X1_291/CTRL 0.01fF
C12468 POR2X1_222/A POR2X1_724/A 0.20fF
C12469 POR2X1_293/Y PAND2X1_156/A 0.10fF
C12470 POR2X1_206/O POR2X1_201/Y 0.02fF
C12471 INPUT_3 POR2X1_67/Y 0.04fF
C12472 POR2X1_99/B POR2X1_243/Y 0.04fF
C12473 POR2X1_43/Y POR2X1_667/A 0.02fF
C12474 POR2X1_322/Y PAND2X1_374/CTRL2 0.00fF
C12475 POR2X1_322/O POR2X1_373/Y 0.01fF
C12476 PAND2X1_801/O POR2X1_236/Y 0.05fF
C12477 POR2X1_570/Y PAND2X1_32/B 0.46fF
C12478 POR2X1_339/CTRL POR2X1_556/Y 0.01fF
C12479 POR2X1_49/a_16_28# POR2X1_29/A 0.02fF
C12480 PAND2X1_640/CTRL2 POR2X1_153/Y 0.02fF
C12481 POR2X1_825/Y POR2X1_32/A 0.03fF
C12482 POR2X1_416/B POR2X1_595/Y 0.02fF
C12483 POR2X1_167/a_16_28# POR2X1_73/Y 0.06fF
C12484 PAND2X1_6/A POR2X1_153/Y 0.19fF
C12485 PAND2X1_90/A POR2X1_571/Y 0.07fF
C12486 POR2X1_720/B POR2X1_720/CTRL 0.00fF
C12487 POR2X1_68/A POR2X1_334/Y 0.10fF
C12488 D_INPUT_3 POR2X1_96/CTRL2 0.12fF
C12489 POR2X1_43/B PAND2X1_123/Y 0.23fF
C12490 PAND2X1_686/O POR2X1_73/Y 0.01fF
C12491 POR2X1_307/Y POR2X1_512/a_16_28# 0.02fF
C12492 POR2X1_661/A POR2X1_646/Y 0.07fF
C12493 POR2X1_78/A POR2X1_651/Y 0.03fF
C12494 POR2X1_616/Y POR2X1_42/Y 0.03fF
C12495 PAND2X1_94/A PAND2X1_111/B 2.91fF
C12496 POR2X1_96/Y POR2X1_58/Y 0.03fF
C12497 POR2X1_13/Y POR2X1_7/Y 0.01fF
C12498 POR2X1_40/Y POR2X1_166/Y 0.18fF
C12499 POR2X1_188/CTRL POR2X1_675/Y 0.01fF
C12500 POR2X1_702/A POR2X1_186/B 0.10fF
C12501 POR2X1_83/B PAND2X1_193/Y 0.02fF
C12502 POR2X1_293/Y PAND2X1_860/CTRL2 0.03fF
C12503 PAND2X1_6/Y POR2X1_342/CTRL2 0.00fF
C12504 PAND2X1_6/Y POR2X1_228/O 0.17fF
C12505 POR2X1_416/B POR2X1_13/CTRL2 0.01fF
C12506 POR2X1_406/Y PAND2X1_339/O 0.04fF
C12507 PAND2X1_175/B PAND2X1_861/O 0.02fF
C12508 POR2X1_318/CTRL2 POR2X1_445/A 0.01fF
C12509 PAND2X1_271/CTRL POR2X1_116/A 0.00fF
C12510 POR2X1_61/A POR2X1_61/B 0.01fF
C12511 POR2X1_390/B POR2X1_337/A 0.05fF
C12512 PAND2X1_704/O POR2X1_142/Y 0.01fF
C12513 POR2X1_71/O POR2X1_91/Y 0.16fF
C12514 POR2X1_411/B POR2X1_24/Y 0.03fF
C12515 POR2X1_73/Y POR2X1_117/Y 0.97fF
C12516 POR2X1_465/B POR2X1_632/Y 0.03fF
C12517 PAND2X1_96/B POR2X1_294/A 5.75fF
C12518 POR2X1_513/Y POR2X1_188/Y 0.03fF
C12519 POR2X1_509/O VDD 0.00fF
C12520 VDD PAND2X1_72/A 2.15fF
C12521 PAND2X1_683/CTRL POR2X1_596/A 0.01fF
C12522 POR2X1_65/A POR2X1_234/A 0.02fF
C12523 POR2X1_346/B POR2X1_61/O 0.00fF
C12524 POR2X1_119/Y POR2X1_38/Y 0.33fF
C12525 POR2X1_188/A POR2X1_643/CTRL 0.01fF
C12526 POR2X1_16/A PAND2X1_317/O 0.05fF
C12527 POR2X1_591/CTRL2 POR2X1_77/Y 0.00fF
C12528 POR2X1_332/B PAND2X1_135/CTRL2 0.01fF
C12529 POR2X1_550/A POR2X1_266/A 0.01fF
C12530 POR2X1_504/Y PAND2X1_630/B 0.02fF
C12531 POR2X1_322/Y PAND2X1_325/a_76_28# 0.02fF
C12532 POR2X1_78/A POR2X1_646/A 0.01fF
C12533 POR2X1_305/Y POR2X1_39/B 0.04fF
C12534 PAND2X1_490/a_76_28# POR2X1_4/Y 0.01fF
C12535 POR2X1_559/A POR2X1_260/A 0.19fF
C12536 POR2X1_329/A PAND2X1_361/O 0.05fF
C12537 VDD POR2X1_535/O 0.00fF
C12538 POR2X1_20/B D_INPUT_0 0.13fF
C12539 POR2X1_864/O POR2X1_814/A 0.04fF
C12540 POR2X1_274/A POR2X1_76/A 0.05fF
C12541 POR2X1_327/Y POR2X1_675/Y 0.03fF
C12542 PAND2X1_838/B POR2X1_48/A 0.03fF
C12543 VDD POR2X1_386/Y 0.29fF
C12544 POR2X1_832/CTRL POR2X1_661/A 0.08fF
C12545 POR2X1_8/Y PAND2X1_358/A 0.19fF
C12546 POR2X1_83/B POR2X1_669/Y 0.13fF
C12547 POR2X1_296/Y POR2X1_296/CTRL2 0.03fF
C12548 POR2X1_624/Y POR2X1_499/O 0.01fF
C12549 POR2X1_741/Y PAND2X1_72/A 0.03fF
C12550 POR2X1_568/B POR2X1_148/A 0.03fF
C12551 PAND2X1_435/Y POR2X1_20/B 0.07fF
C12552 POR2X1_447/B PAND2X1_823/CTRL 0.01fF
C12553 PAND2X1_94/O POR2X1_202/A 0.06fF
C12554 POR2X1_112/a_16_28# POR2X1_510/Y 0.00fF
C12555 PAND2X1_785/O POR2X1_77/Y 0.03fF
C12556 PAND2X1_831/Y POR2X1_39/B 0.01fF
C12557 POR2X1_119/Y INPUT_1 0.07fF
C12558 POR2X1_796/Y POR2X1_678/Y 0.05fF
C12559 POR2X1_60/A POR2X1_253/CTRL2 0.00fF
C12560 PAND2X1_212/O PAND2X1_352/A 0.02fF
C12561 POR2X1_101/Y PAND2X1_136/CTRL 0.30fF
C12562 PAND2X1_72/A PAND2X1_32/B 3.58fF
C12563 POR2X1_567/CTRL2 POR2X1_854/B 0.09fF
C12564 POR2X1_812/A PAND2X1_39/B 0.02fF
C12565 POR2X1_327/Y PAND2X1_683/O 0.06fF
C12566 POR2X1_119/Y POR2X1_153/Y 0.12fF
C12567 PAND2X1_459/O PAND2X1_9/Y 0.01fF
C12568 POR2X1_341/A POR2X1_330/Y 0.07fF
C12569 POR2X1_48/A PAND2X1_400/CTRL 0.01fF
C12570 PAND2X1_294/a_16_344# POR2X1_60/A 0.06fF
C12571 POR2X1_24/O PAND2X1_9/Y 0.01fF
C12572 PAND2X1_444/O PAND2X1_443/Y 0.00fF
C12573 PAND2X1_217/B PAND2X1_203/O 0.03fF
C12574 PAND2X1_488/a_16_344# POR2X1_556/A 0.02fF
C12575 POR2X1_458/Y POR2X1_784/A 0.11fF
C12576 POR2X1_88/CTRL2 POR2X1_69/A 0.01fF
C12577 PAND2X1_33/CTRL POR2X1_5/Y 0.01fF
C12578 POR2X1_6/a_16_28# POR2X1_4/Y 0.01fF
C12579 POR2X1_602/B PAND2X1_601/CTRL2 0.01fF
C12580 POR2X1_741/CTRL POR2X1_186/B 0.01fF
C12581 POR2X1_863/A POR2X1_540/A 0.03fF
C12582 POR2X1_571/Y POR2X1_572/Y 0.20fF
C12583 POR2X1_49/Y POR2X1_54/Y 0.26fF
C12584 POR2X1_126/CTRL POR2X1_94/A 0.08fF
C12585 POR2X1_520/CTRL2 PAND2X1_52/B 0.10fF
C12586 POR2X1_661/A POR2X1_804/A 0.10fF
C12587 POR2X1_814/A POR2X1_193/A 0.12fF
C12588 POR2X1_814/A POR2X1_579/Y 0.07fF
C12589 PAND2X1_282/O POR2X1_590/A 0.04fF
C12590 POR2X1_188/A POR2X1_832/Y 0.03fF
C12591 D_INPUT_7 PAND2X1_587/CTRL2 0.01fF
C12592 PAND2X1_603/O POR2X1_78/A 0.01fF
C12593 POR2X1_814/A POR2X1_572/B 0.03fF
C12594 POR2X1_422/O POR2X1_72/B 0.01fF
C12595 POR2X1_448/CTRL2 POR2X1_296/B 0.05fF
C12596 POR2X1_502/A POR2X1_444/CTRL2 0.01fF
C12597 POR2X1_387/Y POR2X1_310/CTRL2 0.06fF
C12598 POR2X1_661/A PAND2X1_306/CTRL2 0.05fF
C12599 POR2X1_857/A POR2X1_192/Y 0.24fF
C12600 POR2X1_736/A POR2X1_741/A 0.03fF
C12601 POR2X1_267/B POR2X1_260/B 0.01fF
C12602 POR2X1_559/CTRL2 POR2X1_814/A 0.01fF
C12603 POR2X1_567/B POR2X1_355/A 0.03fF
C12604 PAND2X1_687/O POR2X1_761/A 0.05fF
C12605 POR2X1_355/CTRL2 POR2X1_567/B 0.01fF
C12606 POR2X1_859/a_16_28# INPUT_0 0.04fF
C12607 POR2X1_533/O POR2X1_533/Y 0.01fF
C12608 POR2X1_814/A POR2X1_789/A 0.03fF
C12609 POR2X1_568/B POR2X1_337/Y 0.10fF
C12610 POR2X1_78/B POR2X1_222/CTRL 0.08fF
C12611 POR2X1_647/B POR2X1_130/A 0.05fF
C12612 POR2X1_654/B POR2X1_66/A 0.03fF
C12613 POR2X1_614/A POR2X1_814/A 1.16fF
C12614 PAND2X1_717/A POR2X1_90/Y 0.03fF
C12615 PAND2X1_206/A PAND2X1_206/a_76_28# 0.05fF
C12616 POR2X1_556/A POR2X1_795/O 0.06fF
C12617 POR2X1_43/B POR2X1_846/Y 0.00fF
C12618 PAND2X1_57/B POR2X1_648/a_56_344# 0.00fF
C12619 PAND2X1_73/Y POR2X1_750/B 0.08fF
C12620 POR2X1_76/B POR2X1_456/B 0.01fF
C12621 POR2X1_846/Y POR2X1_789/A 0.03fF
C12622 POR2X1_777/B POR2X1_590/A 0.06fF
C12623 POR2X1_814/A POR2X1_38/B 0.01fF
C12624 POR2X1_66/A POR2X1_5/Y 0.07fF
C12625 POR2X1_57/A POR2X1_329/A 0.10fF
C12626 POR2X1_111/O PAND2X1_717/A 0.16fF
C12627 PAND2X1_58/A POR2X1_94/A 0.58fF
C12628 PAND2X1_48/B PAND2X1_39/B 0.10fF
C12629 POR2X1_660/A POR2X1_590/A 0.03fF
C12630 POR2X1_814/A POR2X1_360/CTRL2 0.04fF
C12631 PAND2X1_258/CTRL2 POR2X1_244/B 0.01fF
C12632 PAND2X1_618/a_16_344# PAND2X1_6/A 0.02fF
C12633 PAND2X1_859/B PAND2X1_98/a_76_28# 0.01fF
C12634 POR2X1_66/B POR2X1_476/CTRL 0.00fF
C12635 POR2X1_333/A PAND2X1_41/B 7.76fF
C12636 POR2X1_54/Y POR2X1_642/O 0.01fF
C12637 POR2X1_46/a_16_28# POR2X1_14/Y 0.00fF
C12638 POR2X1_669/B PAND2X1_550/CTRL2 0.03fF
C12639 PAND2X1_65/B POR2X1_590/A 0.08fF
C12640 PAND2X1_625/CTRL PAND2X1_39/B 0.01fF
C12641 POR2X1_748/A POR2X1_72/B 0.03fF
C12642 POR2X1_122/Y POR2X1_669/B 0.29fF
C12643 POR2X1_441/Y POR2X1_438/O 0.01fF
C12644 PAND2X1_462/B PAND2X1_606/CTRL 0.01fF
C12645 POR2X1_484/O VDD 0.00fF
C12646 POR2X1_307/B POR2X1_78/A 0.03fF
C12647 POR2X1_814/B POR2X1_439/CTRL2 0.00fF
C12648 POR2X1_78/B POR2X1_608/Y 0.01fF
C12649 PAND2X1_790/a_16_344# POR2X1_42/Y 0.05fF
C12650 POR2X1_65/A POR2X1_295/CTRL 0.03fF
C12651 POR2X1_333/A POR2X1_781/A 0.03fF
C12652 POR2X1_78/B POR2X1_400/B 0.01fF
C12653 PAND2X1_752/O VDD 0.00fF
C12654 POR2X1_57/A POR2X1_412/a_56_344# 0.01fF
C12655 POR2X1_717/O POR2X1_499/A 0.03fF
C12656 PAND2X1_65/B POR2X1_267/a_76_344# 0.01fF
C12657 POR2X1_52/A POR2X1_626/CTRL 0.00fF
C12658 PAND2X1_41/B POR2X1_734/A 0.15fF
C12659 POR2X1_355/CTRL POR2X1_355/A 0.01fF
C12660 POR2X1_286/B PAND2X1_96/B 0.05fF
C12661 PAND2X1_418/O POR2X1_854/B 0.06fF
C12662 POR2X1_437/CTRL PAND2X1_794/B 0.01fF
C12663 POR2X1_555/A PAND2X1_626/m4_208_n4# 0.15fF
C12664 POR2X1_856/B POR2X1_477/A 0.03fF
C12665 POR2X1_16/A POR2X1_827/m4_208_n4# 0.09fF
C12666 PAND2X1_239/a_76_28# POR2X1_578/Y 0.04fF
C12667 POR2X1_515/a_56_344# PAND2X1_20/A 0.00fF
C12668 POR2X1_626/O POR2X1_55/Y 0.01fF
C12669 POR2X1_508/O POR2X1_567/B 0.01fF
C12670 POR2X1_271/B PAND2X1_549/B 0.05fF
C12671 PAND2X1_262/a_56_28# PAND2X1_41/B 0.00fF
C12672 PAND2X1_471/B POR2X1_83/B 0.11fF
C12673 POR2X1_811/A PAND2X1_599/CTRL 0.00fF
C12674 PAND2X1_58/A PAND2X1_754/CTRL2 0.01fF
C12675 PAND2X1_492/CTRL2 PAND2X1_41/B 0.00fF
C12676 POR2X1_257/A PAND2X1_787/A 0.10fF
C12677 PAND2X1_48/CTRL POR2X1_330/Y 0.02fF
C12678 POR2X1_305/Y POR2X1_48/A 0.07fF
C12679 POR2X1_118/CTRL POR2X1_118/Y 0.01fF
C12680 POR2X1_47/O POR2X1_32/A 0.01fF
C12681 PAND2X1_58/A PAND2X1_110/CTRL2 0.01fF
C12682 POR2X1_40/Y POR2X1_743/m4_208_n4# 0.09fF
C12683 PAND2X1_48/B POR2X1_805/Y 0.03fF
C12684 POR2X1_218/Y POR2X1_218/A 0.09fF
C12685 PAND2X1_90/A PAND2X1_531/O 0.01fF
C12686 PAND2X1_476/a_16_344# INPUT_0 0.01fF
C12687 POR2X1_102/Y PAND2X1_188/CTRL 0.00fF
C12688 POR2X1_718/CTRL2 POR2X1_435/Y 0.01fF
C12689 PAND2X1_795/O PAND2X1_785/Y 0.03fF
C12690 PAND2X1_48/B PAND2X1_20/A 0.10fF
C12691 PAND2X1_206/A PAND2X1_656/A 0.15fF
C12692 POR2X1_752/Y PAND2X1_377/O 0.02fF
C12693 POR2X1_683/O POR2X1_40/Y 0.01fF
C12694 POR2X1_60/Y PAND2X1_351/Y 0.02fF
C12695 POR2X1_143/O POR2X1_40/Y 0.01fF
C12696 PAND2X1_392/O POR2X1_816/A 0.02fF
C12697 POR2X1_60/A POR2X1_406/a_16_28# 0.01fF
C12698 POR2X1_865/B POR2X1_558/B 0.68fF
C12699 POR2X1_16/A POR2X1_63/Y 0.03fF
C12700 POR2X1_788/A PAND2X1_144/O 0.02fF
C12701 POR2X1_644/B POR2X1_644/A 0.00fF
C12702 POR2X1_110/Y PAND2X1_717/A 0.01fF
C12703 PAND2X1_552/A VDD 0.00fF
C12704 PAND2X1_543/O POR2X1_236/Y 0.02fF
C12705 POR2X1_526/CTRL POR2X1_669/B 0.07fF
C12706 PAND2X1_425/Y PAND2X1_157/O 0.02fF
C12707 PAND2X1_473/B VDD 0.28fF
C12708 PAND2X1_65/B PAND2X1_760/CTRL 0.01fF
C12709 POR2X1_43/B POR2X1_421/Y 0.01fF
C12710 POR2X1_55/a_76_344# PAND2X1_6/A 0.00fF
C12711 POR2X1_397/Y VDD 0.05fF
C12712 PAND2X1_793/Y PAND2X1_363/Y 0.02fF
C12713 PAND2X1_16/CTRL2 POR2X1_785/A 0.11fF
C12714 POR2X1_852/B POR2X1_579/Y 0.07fF
C12715 POR2X1_411/B PAND2X1_182/B 0.01fF
C12716 PAND2X1_752/O PAND2X1_32/B 0.04fF
C12717 POR2X1_564/Y PAND2X1_65/B 0.02fF
C12718 PAND2X1_93/B POR2X1_222/A 0.01fF
C12719 PAND2X1_667/CTRL POR2X1_546/A 0.00fF
C12720 PAND2X1_23/Y PAND2X1_250/CTRL 0.06fF
C12721 PAND2X1_48/B PAND2X1_250/O 0.06fF
C12722 PAND2X1_6/Y POR2X1_850/B 0.10fF
C12723 PAND2X1_309/O POR2X1_543/A 0.03fF
C12724 POR2X1_175/O POR2X1_566/A 0.04fF
C12725 POR2X1_16/A POR2X1_88/CTRL2 0.00fF
C12726 PAND2X1_128/CTRL POR2X1_127/Y 0.02fF
C12727 PAND2X1_140/A POR2X1_127/CTRL2 0.01fF
C12728 POR2X1_68/A PAND2X1_96/CTRL2 0.06fF
C12729 PAND2X1_223/a_56_28# POR2X1_7/B 0.00fF
C12730 PAND2X1_48/B POR2X1_814/B 0.28fF
C12731 POR2X1_686/CTRL2 PAND2X1_73/Y 0.01fF
C12732 PAND2X1_826/CTRL2 POR2X1_507/A 0.03fF
C12733 PAND2X1_454/CTRL PAND2X1_803/A 0.00fF
C12734 POR2X1_244/B VDD 0.04fF
C12735 PAND2X1_558/Y PAND2X1_717/O 0.00fF
C12736 POR2X1_857/B PAND2X1_65/B 0.03fF
C12737 PAND2X1_308/B VDD 0.04fF
C12738 POR2X1_448/Y POR2X1_294/B 0.03fF
C12739 POR2X1_341/A POR2X1_715/A 0.04fF
C12740 POR2X1_383/A POR2X1_286/O 0.02fF
C12741 POR2X1_667/A POR2X1_73/Y 0.27fF
C12742 POR2X1_68/B POR2X1_390/O 0.00fF
C12743 POR2X1_83/B PAND2X1_243/O 0.01fF
C12744 POR2X1_494/Y POR2X1_5/Y 0.01fF
C12745 POR2X1_114/B POR2X1_830/a_16_28# 0.03fF
C12746 POR2X1_763/Y PAND2X1_712/B 0.03fF
C12747 POR2X1_16/A PAND2X1_287/Y 0.06fF
C12748 PAND2X1_695/CTRL PAND2X1_48/B 0.01fF
C12749 POR2X1_763/A PAND2X1_709/O 0.05fF
C12750 POR2X1_627/Y VDD 0.10fF
C12751 POR2X1_102/Y POR2X1_93/A 0.06fF
C12752 PAND2X1_659/Y POR2X1_150/Y 0.03fF
C12753 PAND2X1_798/B PAND2X1_220/Y 0.10fF
C12754 POR2X1_356/A POR2X1_856/m4_208_n4# 0.06fF
C12755 POR2X1_389/A PAND2X1_58/A 0.03fF
C12756 PAND2X1_46/CTRL D_INPUT_1 0.00fF
C12757 POR2X1_102/Y POR2X1_91/Y 0.03fF
C12758 POR2X1_66/B POR2X1_68/B 0.28fF
C12759 POR2X1_233/a_16_28# POR2X1_236/Y 0.03fF
C12760 PAND2X1_254/Y POR2X1_516/B 0.16fF
C12761 PAND2X1_48/B POR2X1_325/A 0.03fF
C12762 POR2X1_264/Y PAND2X1_90/Y 0.02fF
C12763 POR2X1_60/A POR2X1_534/CTRL 0.01fF
C12764 POR2X1_778/B POR2X1_389/Y 0.02fF
C12765 POR2X1_811/CTRL2 POR2X1_260/A 0.01fF
C12766 PAND2X1_778/Y PAND2X1_784/A 0.00fF
C12767 POR2X1_52/A PAND2X1_520/O 0.04fF
C12768 PAND2X1_3/a_16_344# PAND2X1_3/A 0.02fF
C12769 POR2X1_653/CTRL POR2X1_740/Y 0.00fF
C12770 POR2X1_315/CTRL PAND2X1_803/A 0.00fF
C12771 PAND2X1_862/B POR2X1_81/Y 0.01fF
C12772 POR2X1_329/A PAND2X1_339/CTRL 0.01fF
C12773 POR2X1_445/A POR2X1_703/CTRL 0.05fF
C12774 POR2X1_13/A POR2X1_372/Y 0.98fF
C12775 PAND2X1_73/m4_208_n4# PAND2X1_69/A 0.07fF
C12776 POR2X1_562/CTRL VDD 0.00fF
C12777 PAND2X1_345/O PAND2X1_555/A 0.06fF
C12778 POR2X1_347/A PAND2X1_94/O 0.00fF
C12779 PAND2X1_116/O POR2X1_183/Y 0.00fF
C12780 POR2X1_83/B PAND2X1_374/CTRL2 0.03fF
C12781 PAND2X1_119/O POR2X1_654/B 0.01fF
C12782 PAND2X1_412/O PAND2X1_32/B 0.15fF
C12783 POR2X1_661/B POR2X1_220/Y 0.03fF
C12784 POR2X1_383/A POR2X1_836/A 0.01fF
C12785 POR2X1_41/B PAND2X1_191/Y 0.03fF
C12786 POR2X1_267/A POR2X1_569/A 0.07fF
C12787 PAND2X1_654/CTRL2 POR2X1_46/Y 0.01fF
C12788 POR2X1_502/A POR2X1_832/B 0.03fF
C12789 POR2X1_612/Y POR2X1_5/CTRL2 -0.00fF
C12790 POR2X1_252/CTRL2 POR2X1_55/Y 0.03fF
C12791 POR2X1_567/B POR2X1_180/CTRL2 0.06fF
C12792 PAND2X1_48/B POR2X1_513/B 0.03fF
C12793 POR2X1_244/B POR2X1_741/Y 0.04fF
C12794 POR2X1_68/A POR2X1_349/Y 0.02fF
C12795 POR2X1_286/CTRL2 POR2X1_774/A 0.01fF
C12796 POR2X1_96/A PAND2X1_575/A 0.03fF
C12797 POR2X1_793/A VDD 0.04fF
C12798 POR2X1_356/A POR2X1_149/Y 0.08fF
C12799 POR2X1_734/A PAND2X1_518/a_76_28# 0.01fF
C12800 PAND2X1_93/CTRL PAND2X1_57/B 0.00fF
C12801 PAND2X1_480/B PAND2X1_717/O 0.06fF
C12802 POR2X1_22/A POR2X1_13/A 0.10fF
C12803 POR2X1_532/A POR2X1_5/Y 0.03fF
C12804 PAND2X1_97/a_76_28# POR2X1_153/Y 0.05fF
C12805 POR2X1_251/Y PAND2X1_675/A 2.28fF
C12806 POR2X1_331/A POR2X1_331/a_16_28# 0.02fF
C12807 POR2X1_13/A POR2X1_494/CTRL 0.01fF
C12808 POR2X1_435/Y POR2X1_804/B 0.08fF
C12809 POR2X1_41/B POR2X1_83/A 0.00fF
C12810 POR2X1_96/A PAND2X1_794/B 0.08fF
C12811 POR2X1_811/B POR2X1_260/A 0.02fF
C12812 POR2X1_612/B POR2X1_4/Y 0.02fF
C12813 POR2X1_231/CTRL POR2X1_795/B 0.08fF
C12814 POR2X1_793/A POR2X1_793/a_16_28# 0.03fF
C12815 PAND2X1_90/Y POR2X1_712/CTRL 0.07fF
C12816 PAND2X1_766/CTRL POR2X1_707/Y 0.01fF
C12817 POR2X1_483/A POR2X1_702/CTRL2 0.01fF
C12818 PAND2X1_688/CTRL POR2X1_38/Y 0.01fF
C12819 POR2X1_43/B INPUT_5 0.00fF
C12820 POR2X1_296/B POR2X1_673/B 0.05fF
C12821 PAND2X1_335/CTRL2 POR2X1_309/Y 0.01fF
C12822 POR2X1_479/B PAND2X1_48/A 0.03fF
C12823 POR2X1_52/A POR2X1_617/a_16_28# 0.00fF
C12824 POR2X1_441/Y PAND2X1_326/CTRL2 0.01fF
C12825 POR2X1_763/Y PAND2X1_546/CTRL2 0.05fF
C12826 PAND2X1_862/B PAND2X1_858/Y 0.15fF
C12827 POR2X1_669/B PAND2X1_508/Y 0.03fF
C12828 POR2X1_43/B PAND2X1_724/B 0.04fF
C12829 POR2X1_770/a_16_28# POR2X1_770/A 0.03fF
C12830 POR2X1_41/B POR2X1_90/Y 0.22fF
C12831 D_GATE_662 POR2X1_732/B 0.10fF
C12832 PAND2X1_61/Y POR2X1_521/Y 0.01fF
C12833 POR2X1_859/A POR2X1_68/B 0.06fF
C12834 POR2X1_37/Y POR2X1_171/Y 0.04fF
C12835 PAND2X1_665/CTRL2 PAND2X1_93/B 0.02fF
C12836 POR2X1_627/O POR2X1_7/A 0.02fF
C12837 PAND2X1_493/CTRL2 POR2X1_60/A 0.01fF
C12838 POR2X1_131/Y PAND2X1_140/O 0.08fF
C12839 POR2X1_312/Y POR2X1_176/Y 0.01fF
C12840 POR2X1_853/A POR2X1_795/B 0.06fF
C12841 PAND2X1_631/A POR2X1_482/CTRL2 0.01fF
C12842 POR2X1_608/Y POR2X1_294/A 0.02fF
C12843 POR2X1_57/A POR2X1_821/a_56_344# 0.00fF
C12844 PAND2X1_206/CTRL POR2X1_7/A 0.01fF
C12845 POR2X1_669/B POR2X1_320/CTRL 0.10fF
C12846 POR2X1_400/B POR2X1_294/A 0.01fF
C12847 POR2X1_66/A PAND2X1_41/Y 0.01fF
C12848 POR2X1_13/A POR2X1_9/O 0.01fF
C12849 POR2X1_41/B POR2X1_111/O 0.05fF
C12850 POR2X1_65/A POR2X1_527/O 0.01fF
C12851 POR2X1_616/Y POR2X1_67/A 0.50fF
C12852 PAND2X1_755/O PAND2X1_60/B 0.03fF
C12853 POR2X1_376/B PAND2X1_155/O 0.17fF
C12854 POR2X1_685/CTRL2 POR2X1_687/A 0.01fF
C12855 PAND2X1_273/CTRL2 PAND2X1_69/A 0.01fF
C12856 POR2X1_820/Y POR2X1_7/A 0.03fF
C12857 POR2X1_112/CTRL2 POR2X1_241/B 0.08fF
C12858 PAND2X1_653/Y PAND2X1_218/CTRL2 0.04fF
C12859 POR2X1_327/Y POR2X1_405/CTRL 0.02fF
C12860 POR2X1_52/A POR2X1_619/Y 0.03fF
C12861 POR2X1_116/CTRL2 POR2X1_260/A 0.14fF
C12862 PAND2X1_480/CTRL2 PAND2X1_803/A 0.00fF
C12863 PAND2X1_651/Y PAND2X1_242/O 0.00fF
C12864 PAND2X1_682/O POR2X1_407/A 0.06fF
C12865 PAND2X1_20/A PAND2X1_527/a_16_344# 0.01fF
C12866 POR2X1_124/a_16_28# PAND2X1_96/B 0.02fF
C12867 PAND2X1_219/A POR2X1_7/Y 0.03fF
C12868 PAND2X1_64/O D_INPUT_4 0.16fF
C12869 PAND2X1_852/CTRL POR2X1_73/Y 0.04fF
C12870 PAND2X1_117/a_76_28# PAND2X1_32/B 0.01fF
C12871 POR2X1_20/B POR2X1_90/O 0.01fF
C12872 POR2X1_16/A PAND2X1_645/CTRL 0.01fF
C12873 PAND2X1_291/CTRL POR2X1_198/B 0.01fF
C12874 POR2X1_492/a_16_28# POR2X1_394/A 0.12fF
C12875 POR2X1_65/A PAND2X1_120/CTRL 0.01fF
C12876 POR2X1_677/O POR2X1_129/Y 0.00fF
C12877 VDD POR2X1_534/Y 0.03fF
C12878 POR2X1_732/B POR2X1_724/A 0.01fF
C12879 POR2X1_65/CTRL2 POR2X1_9/Y 0.02fF
C12880 POR2X1_697/Y POR2X1_511/O 0.01fF
C12881 POR2X1_99/A POR2X1_294/A 0.13fF
C12882 PAND2X1_798/B PAND2X1_575/CTRL 0.01fF
C12883 POR2X1_68/A POR2X1_140/CTRL 0.00fF
C12884 POR2X1_493/O POR2X1_572/B 0.07fF
C12885 PAND2X1_344/O PAND2X1_514/Y 0.01fF
C12886 PAND2X1_86/Y POR2X1_243/Y 0.02fF
C12887 PAND2X1_636/CTRL POR2X1_260/A 0.08fF
C12888 POR2X1_83/CTRL PAND2X1_35/Y 0.01fF
C12889 PAND2X1_490/CTRL2 POR2X1_532/A 0.01fF
C12890 PAND2X1_480/O POR2X1_236/Y 0.02fF
C12891 POR2X1_334/CTRL PAND2X1_57/B 0.03fF
C12892 POR2X1_407/Y POR2X1_770/CTRL2 0.01fF
C12893 POR2X1_343/Y D_INPUT_0 0.05fF
C12894 PAND2X1_237/CTRL2 PAND2X1_72/A 0.10fF
C12895 PAND2X1_579/A PAND2X1_579/B 0.00fF
C12896 PAND2X1_341/Y INPUT_0 0.01fF
C12897 PAND2X1_55/Y PAND2X1_63/B 0.03fF
C12898 PAND2X1_776/a_76_28# POR2X1_91/Y 0.02fF
C12899 PAND2X1_661/Y POR2X1_42/Y 0.03fF
C12900 POR2X1_86/Y D_INPUT_0 0.01fF
C12901 PAND2X1_213/Y PAND2X1_566/Y 0.00fF
C12902 POR2X1_35/Y PAND2X1_60/B 0.03fF
C12903 POR2X1_114/CTRL POR2X1_113/Y 0.06fF
C12904 POR2X1_49/Y POR2X1_4/Y 0.03fF
C12905 POR2X1_51/A POR2X1_744/a_16_28# 0.02fF
C12906 POR2X1_41/B PAND2X1_732/A 0.07fF
C12907 PAND2X1_666/CTRL PAND2X1_72/A 0.01fF
C12908 PAND2X1_472/CTRL POR2X1_7/B 0.01fF
C12909 PAND2X1_109/a_76_28# POR2X1_97/A 0.01fF
C12910 POR2X1_786/Y POR2X1_228/Y 0.10fF
C12911 POR2X1_783/B POR2X1_260/A 0.02fF
C12912 PAND2X1_564/a_16_344# POR2X1_394/A 0.02fF
C12913 POR2X1_355/B POR2X1_317/B 0.03fF
C12914 PAND2X1_342/CTRL POR2X1_248/Y 0.03fF
C12915 PAND2X1_23/Y INPUT_1 0.06fF
C12916 POR2X1_730/Y POR2X1_740/Y 0.03fF
C12917 POR2X1_409/O POR2X1_408/Y 0.05fF
C12918 POR2X1_494/CTRL PAND2X1_510/B 0.01fF
C12919 POR2X1_722/CTRL VDD 0.00fF
C12920 POR2X1_244/B POR2X1_228/CTRL 0.01fF
C12921 PAND2X1_723/O POR2X1_7/A 0.03fF
C12922 PAND2X1_569/A POR2X1_765/Y 0.01fF
C12923 POR2X1_143/CTRL2 POR2X1_62/Y 0.01fF
C12924 POR2X1_537/Y VDD 0.09fF
C12925 POR2X1_814/CTRL POR2X1_260/B 0.00fF
C12926 PAND2X1_483/CTRL2 PAND2X1_6/A 0.03fF
C12927 POR2X1_111/CTRL2 POR2X1_283/A 0.03fF
C12928 POR2X1_339/a_16_28# POR2X1_785/A 0.03fF
C12929 POR2X1_840/CTRL POR2X1_725/Y 0.07fF
C12930 POR2X1_655/Y POR2X1_711/Y 0.03fF
C12931 POR2X1_327/Y POR2X1_276/CTRL 0.01fF
C12932 PAND2X1_824/B PAND2X1_93/CTRL2 0.01fF
C12933 POR2X1_730/Y POR2X1_732/O 0.01fF
C12934 POR2X1_114/CTRL POR2X1_260/A 0.01fF
C12935 POR2X1_383/A POR2X1_712/CTRL2 0.03fF
C12936 POR2X1_394/A PAND2X1_705/CTRL2 0.01fF
C12937 POR2X1_65/A POR2X1_39/B 4.26fF
C12938 POR2X1_41/B POR2X1_110/Y 0.09fF
C12939 PAND2X1_843/CTRL POR2X1_416/B 0.10fF
C12940 PAND2X1_687/O POR2X1_829/A 0.00fF
C12941 PAND2X1_644/a_16_344# POR2X1_597/Y 0.02fF
C12942 POR2X1_791/CTRL PAND2X1_48/A 0.01fF
C12943 PAND2X1_863/A VDD 0.10fF
C12944 PAND2X1_659/Y PAND2X1_364/B 0.07fF
C12945 POR2X1_776/B POR2X1_192/B 0.03fF
C12946 POR2X1_123/A PAND2X1_60/B 0.00fF
C12947 PAND2X1_357/Y PAND2X1_348/A 0.07fF
C12948 PAND2X1_721/CTRL2 POR2X1_77/Y -0.00fF
C12949 POR2X1_865/B POR2X1_362/A 0.15fF
C12950 PAND2X1_48/B POR2X1_726/CTRL 0.01fF
C12951 POR2X1_710/B POR2X1_713/B 0.00fF
C12952 PAND2X1_854/A POR2X1_765/Y 0.02fF
C12953 PAND2X1_308/Y POR2X1_90/Y 2.33fF
C12954 PAND2X1_90/Y POR2X1_779/O 0.05fF
C12955 POR2X1_57/A POR2X1_744/O 0.03fF
C12956 PAND2X1_820/m4_208_n4# POR2X1_617/m4_208_n4# 0.05fF
C12957 POR2X1_16/A PAND2X1_284/Y 0.01fF
C12958 PAND2X1_737/O POR2X1_7/B 0.04fF
C12959 POR2X1_416/B PAND2X1_76/Y 12.19fF
C12960 PAND2X1_94/A PAND2X1_491/m4_208_n4# 0.07fF
C12961 POR2X1_176/CTRL PAND2X1_566/Y 0.03fF
C12962 POR2X1_537/Y POR2X1_741/Y 1.20fF
C12963 PAND2X1_28/O PAND2X1_63/B 0.02fF
C12964 PAND2X1_439/CTRL POR2X1_438/Y 0.01fF
C12965 POR2X1_486/B PAND2X1_57/B 0.13fF
C12966 POR2X1_276/Y POR2X1_366/A 0.57fF
C12967 PAND2X1_462/CTRL VDD 0.00fF
C12968 POR2X1_307/CTRL POR2X1_661/A 0.08fF
C12969 PAND2X1_96/B POR2X1_543/a_16_28# 0.02fF
C12970 POR2X1_285/B VDD 0.04fF
C12971 POR2X1_334/Y PAND2X1_96/B 0.07fF
C12972 PAND2X1_170/O POR2X1_73/Y 0.02fF
C12973 POR2X1_553/CTRL2 POR2X1_573/A 0.00fF
C12974 POR2X1_804/A POR2X1_737/A 0.03fF
C12975 VDD PAND2X1_861/B 0.10fF
C12976 POR2X1_155/CTRL2 POR2X1_728/A 0.00fF
C12977 POR2X1_711/B POR2X1_710/O 0.01fF
C12978 POR2X1_861/A POR2X1_218/A 0.01fF
C12979 PAND2X1_236/O PAND2X1_52/B 0.02fF
C12980 POR2X1_661/A POR2X1_794/B 0.07fF
C12981 POR2X1_537/Y PAND2X1_32/B 0.03fF
C12982 INPUT_6 PAND2X1_2/CTRL 0.01fF
C12983 POR2X1_283/A POR2X1_394/A 0.13fF
C12984 POR2X1_394/A PAND2X1_121/CTRL 0.03fF
C12985 POR2X1_814/A POR2X1_590/A 0.20fF
C12986 POR2X1_814/B PAND2X1_233/CTRL2 0.05fF
C12987 POR2X1_159/O POR2X1_9/Y 0.02fF
C12988 POR2X1_257/A PAND2X1_469/O 0.06fF
C12989 POR2X1_466/A POR2X1_453/Y 0.16fF
C12990 PAND2X1_351/Y PAND2X1_351/A 0.02fF
C12991 POR2X1_675/Y POR2X1_737/a_16_28# 0.02fF
C12992 POR2X1_537/B PAND2X1_48/A 0.01fF
C12993 POR2X1_329/A PAND2X1_215/CTRL2 0.03fF
C12994 POR2X1_270/Y POR2X1_556/A 0.12fF
C12995 POR2X1_681/O POR2X1_32/A 0.02fF
C12996 PAND2X1_453/m4_208_n4# POR2X1_77/Y 0.08fF
C12997 POR2X1_119/Y PAND2X1_470/A 0.15fF
C12998 POR2X1_83/A POR2X1_77/Y 0.02fF
C12999 POR2X1_356/A POR2X1_568/A 0.07fF
C13000 POR2X1_158/Y PAND2X1_705/CTRL 0.00fF
C13001 POR2X1_193/A PAND2X1_135/CTRL2 0.00fF
C13002 POR2X1_579/Y PAND2X1_135/CTRL2 0.00fF
C13003 PAND2X1_713/CTRL2 POR2X1_394/A 0.01fF
C13004 POR2X1_416/B PAND2X1_566/Y 0.12fF
C13005 POR2X1_55/a_16_28# POR2X1_623/Y 0.02fF
C13006 POR2X1_257/A POR2X1_695/Y 0.08fF
C13007 POR2X1_673/CTRL POR2X1_624/B 0.04fF
C13008 POR2X1_90/Y POR2X1_77/Y 9.16fF
C13009 POR2X1_160/CTRL POR2X1_356/B 0.01fF
C13010 POR2X1_624/Y D_INPUT_0 0.11fF
C13011 PAND2X1_865/Y PAND2X1_489/CTRL2 0.00fF
C13012 POR2X1_760/A PAND2X1_361/a_56_28# 0.00fF
C13013 POR2X1_96/A PAND2X1_221/Y 0.01fF
C13014 POR2X1_449/A POR2X1_802/A 0.03fF
C13015 POR2X1_110/Y PAND2X1_308/Y 0.03fF
C13016 POR2X1_622/O VDD 0.00fF
C13017 POR2X1_383/A POR2X1_383/Y 0.06fF
C13018 POR2X1_614/A PAND2X1_135/CTRL2 0.03fF
C13019 POR2X1_838/B PAND2X1_67/CTRL 0.00fF
C13020 POR2X1_431/CTRL2 POR2X1_236/Y 0.03fF
C13021 PAND2X1_60/CTRL PAND2X1_58/A 0.01fF
C13022 POR2X1_329/A PAND2X1_84/Y 0.03fF
C13023 POR2X1_431/Y PAND2X1_390/Y 0.01fF
C13024 POR2X1_417/Y PAND2X1_211/CTRL2 0.01fF
C13025 PAND2X1_20/A D_INPUT_5 0.01fF
C13026 POR2X1_158/Y POR2X1_695/CTRL 0.00fF
C13027 POR2X1_65/A POR2X1_65/a_16_28# 0.02fF
C13028 PAND2X1_74/a_16_344# POR2X1_341/A 0.03fF
C13029 POR2X1_579/CTRL PAND2X1_32/B 0.01fF
C13030 POR2X1_486/CTRL2 PAND2X1_57/B 0.01fF
C13031 POR2X1_863/A PAND2X1_69/A 0.03fF
C13032 POR2X1_416/B PAND2X1_551/a_76_28# 0.01fF
C13033 POR2X1_315/Y POR2X1_416/B 0.03fF
C13034 POR2X1_119/Y POR2X1_150/CTRL2 0.13fF
C13035 POR2X1_220/A POR2X1_568/A 0.03fF
C13036 POR2X1_837/A PAND2X1_55/Y 0.15fF
C13037 POR2X1_536/Y PAND2X1_222/A 0.06fF
C13038 POR2X1_499/A POR2X1_573/O 0.00fF
C13039 POR2X1_417/Y PAND2X1_212/CTRL2 0.01fF
C13040 POR2X1_602/a_16_28# POR2X1_602/A 0.05fF
C13041 POR2X1_857/B POR2X1_814/A 0.07fF
C13042 POR2X1_317/A PAND2X1_52/B 0.04fF
C13043 POR2X1_66/B POR2X1_848/A 0.07fF
C13044 POR2X1_49/Y PAND2X1_469/O 0.13fF
C13045 POR2X1_146/Y PAND2X1_797/Y 0.04fF
C13046 POR2X1_35/B POR2X1_34/CTRL 0.01fF
C13047 POR2X1_150/Y PAND2X1_151/CTRL2 0.03fF
C13048 PAND2X1_10/O POR2X1_296/B 0.03fF
C13049 POR2X1_842/CTRL POR2X1_794/B 0.03fF
C13050 POR2X1_260/B POR2X1_391/A 0.02fF
C13051 POR2X1_566/A POR2X1_318/CTRL 0.30fF
C13052 PAND2X1_56/Y PAND2X1_75/CTRL2 0.03fF
C13053 POR2X1_135/Y POR2X1_257/A 0.11fF
C13054 POR2X1_9/Y PAND2X1_69/A 0.07fF
C13055 POR2X1_13/A POR2X1_292/Y 0.23fF
C13056 POR2X1_411/B POR2X1_88/Y 0.03fF
C13057 POR2X1_20/B PAND2X1_735/Y 0.33fF
C13058 POR2X1_427/CTRL2 POR2X1_40/Y 0.01fF
C13059 POR2X1_158/Y PAND2X1_713/CTRL 0.00fF
C13060 POR2X1_630/B D_GATE_222 0.09fF
C13061 POR2X1_9/Y PAND2X1_341/A 0.03fF
C13062 PAND2X1_860/A PAND2X1_175/B 0.03fF
C13063 POR2X1_677/Y POR2X1_91/Y 0.03fF
C13064 POR2X1_332/B POR2X1_341/A 0.02fF
C13065 POR2X1_777/B POR2X1_66/A 0.08fF
C13066 POR2X1_54/Y PAND2X1_8/Y 0.36fF
C13067 PAND2X1_620/Y POR2X1_48/A 0.03fF
C13068 POR2X1_9/Y POR2X1_93/A 0.09fF
C13069 PAND2X1_783/B PAND2X1_783/O 0.00fF
C13070 POR2X1_150/Y POR2X1_293/Y 0.04fF
C13071 PAND2X1_222/A PAND2X1_730/B 0.03fF
C13072 POR2X1_220/CTRL VDD 0.00fF
C13073 POR2X1_65/A POR2X1_48/A 0.26fF
C13074 POR2X1_66/A POR2X1_194/A 0.10fF
C13075 POR2X1_705/B POR2X1_294/B 0.02fF
C13076 POR2X1_479/B POR2X1_288/A 0.07fF
C13077 PAND2X1_58/A POR2X1_753/m4_208_n4# 0.05fF
C13078 PAND2X1_431/m4_208_n4# POR2X1_453/m4_208_n4# 0.13fF
C13079 POR2X1_78/B POR2X1_260/B 6.00fF
C13080 POR2X1_329/A POR2X1_594/A 0.53fF
C13081 POR2X1_319/A VDD 0.13fF
C13082 POR2X1_110/Y POR2X1_77/Y 0.03fF
C13083 PAND2X1_73/Y PAND2X1_46/O 0.11fF
C13084 PAND2X1_841/O POR2X1_271/B 0.02fF
C13085 PAND2X1_96/CTRL2 PAND2X1_58/A 0.00fF
C13086 POR2X1_115/O POR2X1_446/B 0.01fF
C13087 POR2X1_38/O VDD 0.00fF
C13088 PAND2X1_65/B POR2X1_66/A 3.62fF
C13089 POR2X1_416/Y POR2X1_412/CTRL 0.01fF
C13090 PAND2X1_218/B VDD 0.08fF
C13091 PAND2X1_282/a_76_28# PAND2X1_41/B 0.02fF
C13092 POR2X1_833/a_56_344# POR2X1_541/B 0.00fF
C13093 POR2X1_566/A POR2X1_854/a_16_28# 0.02fF
C13094 PAND2X1_431/CTRL VDD -0.00fF
C13095 POR2X1_416/B PAND2X1_737/CTRL 0.02fF
C13096 PAND2X1_39/B POR2X1_717/Y 0.06fF
C13097 POR2X1_257/A PAND2X1_274/m4_208_n4# 0.09fF
C13098 PAND2X1_617/O POR2X1_68/B 0.03fF
C13099 PAND2X1_859/A POR2X1_83/B 0.03fF
C13100 POR2X1_79/Y PAND2X1_205/O 0.02fF
C13101 PAND2X1_449/O POR2X1_90/Y 0.02fF
C13102 POR2X1_848/A POR2X1_859/A 0.87fF
C13103 PAND2X1_803/A POR2X1_32/A 0.03fF
C13104 POR2X1_682/CTRL POR2X1_60/A 0.01fF
C13105 POR2X1_35/B PAND2X1_616/CTRL2 0.01fF
C13106 PAND2X1_721/B PAND2X1_721/CTRL 0.01fF
C13107 PAND2X1_20/A POR2X1_489/O 0.02fF
C13108 POR2X1_19/CTRL POR2X1_38/B 0.00fF
C13109 PAND2X1_169/Y PAND2X1_168/Y 0.14fF
C13110 POR2X1_338/O POR2X1_814/A 0.10fF
C13111 POR2X1_179/a_16_28# POR2X1_150/Y 0.02fF
C13112 POR2X1_423/Y POR2X1_40/Y 0.07fF
C13113 POR2X1_667/Y VDD -0.00fF
C13114 PAND2X1_677/CTRL2 POR2X1_718/A 0.01fF
C13115 POR2X1_68/O PAND2X1_57/B 0.01fF
C13116 POR2X1_257/A POR2X1_816/A 0.05fF
C13117 POR2X1_257/A PAND2X1_569/A 0.09fF
C13118 POR2X1_413/A POR2X1_612/Y 0.10fF
C13119 POR2X1_567/B POR2X1_340/CTRL 0.02fF
C13120 POR2X1_61/B POR2X1_202/A 0.03fF
C13121 POR2X1_417/Y PAND2X1_803/A 0.02fF
C13122 POR2X1_61/Y POR2X1_750/B 0.10fF
C13123 POR2X1_460/O POR2X1_260/B 0.01fF
C13124 POR2X1_66/B POR2X1_480/A 0.03fF
C13125 PAND2X1_843/O PAND2X1_220/Y 0.03fF
C13126 POR2X1_231/O POR2X1_66/A 0.01fF
C13127 POR2X1_49/Y PAND2X1_714/A 0.07fF
C13128 POR2X1_812/A VDD 0.10fF
C13129 PAND2X1_61/O POR2X1_58/Y 0.03fF
C13130 POR2X1_640/m4_208_n4# PAND2X1_41/B 0.12fF
C13131 PAND2X1_10/CTRL2 PAND2X1_55/Y 0.03fF
C13132 POR2X1_582/O POR2X1_257/A 0.02fF
C13133 POR2X1_72/B PAND2X1_778/CTRL 0.01fF
C13134 POR2X1_188/A POR2X1_480/A 0.03fF
C13135 POR2X1_96/A POR2X1_83/B 0.15fF
C13136 POR2X1_218/Y POR2X1_740/Y 0.10fF
C13137 PAND2X1_23/Y POR2X1_637/O 0.01fF
C13138 D_GATE_662 POR2X1_466/A 0.10fF
C13139 POR2X1_274/A PAND2X1_69/A 0.01fF
C13140 POR2X1_142/a_16_28# PAND2X1_738/Y 0.02fF
C13141 POR2X1_346/CTRL POR2X1_202/A 0.04fF
C13142 POR2X1_502/A POR2X1_634/A 0.14fF
C13143 POR2X1_346/B POR2X1_66/O 0.00fF
C13144 POR2X1_801/CTRL2 VDD 0.00fF
C13145 POR2X1_556/A POR2X1_101/Y 0.01fF
C13146 PAND2X1_96/B POR2X1_805/O 0.00fF
C13147 PAND2X1_480/B POR2X1_272/CTRL -0.00fF
C13148 POR2X1_58/Y POR2X1_60/A 0.08fF
C13149 POR2X1_96/A POR2X1_626/Y 0.00fF
C13150 POR2X1_403/CTRL2 POR2X1_403/B 0.03fF
C13151 POR2X1_13/A PAND2X1_795/CTRL 0.01fF
C13152 POR2X1_66/B POR2X1_553/Y 0.01fF
C13153 PAND2X1_81/CTRL POR2X1_66/A 0.03fF
C13154 POR2X1_43/B POR2X1_496/Y 0.07fF
C13155 POR2X1_499/A POR2X1_456/B 0.57fF
C13156 POR2X1_489/B POR2X1_294/B 0.03fF
C13157 POR2X1_135/Y POR2X1_45/CTRL2 0.01fF
C13158 POR2X1_78/A POR2X1_732/B 1.96fF
C13159 POR2X1_407/A POR2X1_801/B 0.01fF
C13160 PAND2X1_821/O POR2X1_590/A 0.15fF
C13161 PAND2X1_479/O VDD 0.00fF
C13162 PAND2X1_23/Y POR2X1_287/a_56_344# 0.00fF
C13163 POR2X1_497/Y POR2X1_5/Y 0.03fF
C13164 POR2X1_554/B POR2X1_244/Y 0.10fF
C13165 PAND2X1_219/B VDD 0.03fF
C13166 POR2X1_748/A POR2X1_7/B 0.05fF
C13167 POR2X1_68/CTRL PAND2X1_69/A 0.01fF
C13168 POR2X1_494/CTRL POR2X1_29/A 0.01fF
C13169 PAND2X1_793/Y PAND2X1_217/B 0.05fF
C13170 POR2X1_66/B PAND2X1_90/A 0.03fF
C13171 POR2X1_52/A PAND2X1_725/Y 0.03fF
C13172 PAND2X1_859/A POR2X1_224/a_16_28# 0.02fF
C13173 POR2X1_14/Y POR2X1_584/CTRL2 0.00fF
C13174 POR2X1_652/Y POR2X1_750/B 0.03fF
C13175 POR2X1_624/Y PAND2X1_133/CTRL 0.00fF
C13176 D_INPUT_0 POR2X1_73/Y 0.26fF
C13177 POR2X1_188/A PAND2X1_753/O 0.00fF
C13178 POR2X1_502/A PAND2X1_588/CTRL2 0.01fF
C13179 POR2X1_376/B POR2X1_88/Y 0.05fF
C13180 POR2X1_407/A POR2X1_287/O 0.01fF
C13181 PAND2X1_215/B POR2X1_72/B 0.07fF
C13182 POR2X1_8/Y POR2X1_411/B 0.07fF
C13183 POR2X1_260/B POR2X1_391/CTRL 0.01fF
C13184 POR2X1_29/Y POR2X1_29/A 0.46fF
C13185 PAND2X1_403/B PAND2X1_398/CTRL 0.01fF
C13186 POR2X1_346/CTRL POR2X1_346/A 0.01fF
C13187 POR2X1_466/A POR2X1_724/A 0.09fF
C13188 POR2X1_311/Y PAND2X1_794/B 0.03fF
C13189 PAND2X1_124/Y POR2X1_7/A 0.03fF
C13190 POR2X1_857/B POR2X1_852/B 0.04fF
C13191 POR2X1_500/A POR2X1_500/a_16_28# 0.03fF
C13192 POR2X1_60/a_16_28# POR2X1_23/Y 0.03fF
C13193 PAND2X1_63/Y POR2X1_296/B 0.03fF
C13194 PAND2X1_282/O POR2X1_532/A 0.13fF
C13195 PAND2X1_738/B POR2X1_763/Y 0.07fF
C13196 PAND2X1_58/O VDD 0.00fF
C13197 POR2X1_260/B POR2X1_141/A 0.48fF
C13198 PAND2X1_262/O POR2X1_786/A 0.11fF
C13199 PAND2X1_862/B PAND2X1_659/CTRL2 0.01fF
C13200 POR2X1_750/B PAND2X1_178/a_16_344# 0.02fF
C13201 POR2X1_66/B PAND2X1_697/CTRL 0.00fF
C13202 PAND2X1_192/Y PAND2X1_191/O 0.03fF
C13203 PAND2X1_638/B PAND2X1_69/A 0.09fF
C13204 PAND2X1_435/Y POR2X1_73/Y 0.95fF
C13205 POR2X1_514/Y POR2X1_141/Y 0.01fF
C13206 PAND2X1_612/B POR2X1_773/B 0.00fF
C13207 POR2X1_445/A POR2X1_543/CTRL 0.03fF
C13208 POR2X1_43/B PAND2X1_733/A 0.03fF
C13209 POR2X1_634/O POR2X1_391/Y 0.04fF
C13210 POR2X1_483/B VDD 0.19fF
C13211 POR2X1_682/Y VDD 0.01fF
C13212 POR2X1_814/B POR2X1_717/Y 0.99fF
C13213 PAND2X1_9/O D_INPUT_1 0.04fF
C13214 PAND2X1_453/O POR2X1_376/B 0.04fF
C13215 POR2X1_750/B POR2X1_35/Y 0.05fF
C13216 POR2X1_52/A PAND2X1_84/CTRL2 0.03fF
C13217 PAND2X1_592/CTRL VDD 0.00fF
C13218 POR2X1_222/Y POR2X1_194/A 0.03fF
C13219 POR2X1_812/A PAND2X1_32/B 0.03fF
C13220 PAND2X1_696/O POR2X1_648/Y 0.01fF
C13221 POR2X1_502/A POR2X1_130/A 0.03fF
C13222 POR2X1_376/B POR2X1_743/Y 0.01fF
C13223 POR2X1_52/A POR2X1_697/O 0.06fF
C13224 POR2X1_666/Y POR2X1_665/Y 0.07fF
C13225 PAND2X1_6/A POR2X1_72/B 0.07fF
C13226 POR2X1_776/A POR2X1_566/O 0.01fF
C13227 POR2X1_135/Y PAND2X1_553/B 0.01fF
C13228 POR2X1_329/O PAND2X1_362/B 0.01fF
C13229 PAND2X1_243/B POR2X1_236/Y 0.02fF
C13230 PAND2X1_793/Y VDD 0.07fF
C13231 POR2X1_13/A POR2X1_295/Y 0.11fF
C13232 PAND2X1_724/CTRL2 PAND2X1_169/Y 0.00fF
C13233 PAND2X1_11/a_16_344# D_INPUT_4 0.02fF
C13234 POR2X1_41/B INPUT_0 0.44fF
C13235 POR2X1_96/A PAND2X1_795/B 0.19fF
C13236 PAND2X1_244/B D_INPUT_0 0.03fF
C13237 POR2X1_566/A POR2X1_502/A 0.19fF
C13238 PAND2X1_35/Y PAND2X1_673/Y 0.00fF
C13239 POR2X1_302/B POR2X1_804/A 0.03fF
C13240 POR2X1_406/Y PAND2X1_364/B 0.07fF
C13241 PAND2X1_96/B PAND2X1_96/CTRL2 0.03fF
C13242 POR2X1_60/A POR2X1_9/CTRL 0.02fF
C13243 PAND2X1_841/B VDD 0.02fF
C13244 POR2X1_49/Y POR2X1_816/A 0.03fF
C13245 PAND2X1_152/O VDD 0.00fF
C13246 PAND2X1_65/B POR2X1_222/Y 0.03fF
C13247 PAND2X1_849/B POR2X1_37/Y 3.02fF
C13248 PAND2X1_258/CTRL POR2X1_260/A 0.01fF
C13249 POR2X1_78/B PAND2X1_55/Y 0.23fF
C13250 POR2X1_79/A POR2X1_7/B 0.01fF
C13251 PAND2X1_6/Y PAND2X1_423/O 0.17fF
C13252 PAND2X1_48/B VDD 2.38fF
C13253 POR2X1_43/B PAND2X1_276/CTRL 0.00fF
C13254 POR2X1_648/Y POR2X1_779/CTRL 0.01fF
C13255 POR2X1_254/Y POR2X1_795/CTRL2 0.08fF
C13256 POR2X1_83/B POR2X1_7/A 2.24fF
C13257 POR2X1_566/A PAND2X1_176/O 0.03fF
C13258 PAND2X1_319/B POR2X1_40/Y 0.07fF
C13259 POR2X1_66/B PAND2X1_397/CTRL2 0.02fF
C13260 PAND2X1_736/A PAND2X1_740/Y 0.10fF
C13261 POR2X1_311/Y POR2X1_107/Y 0.00fF
C13262 PAND2X1_232/CTRL2 POR2X1_590/A 0.00fF
C13263 PAND2X1_837/CTRL POR2X1_39/B 0.01fF
C13264 POR2X1_78/B POR2X1_788/Y 0.02fF
C13265 POR2X1_84/CTRL PAND2X1_57/B 0.01fF
C13266 PAND2X1_138/a_16_344# POR2X1_136/Y 0.02fF
C13267 PAND2X1_436/O PAND2X1_508/Y 0.04fF
C13268 PAND2X1_707/Y PAND2X1_707/O 0.01fF
C13269 POR2X1_127/Y PAND2X1_284/Y 0.03fF
C13270 POR2X1_94/A POR2X1_380/Y 0.05fF
C13271 POR2X1_626/Y POR2X1_7/A 0.00fF
C13272 POR2X1_325/CTRL2 POR2X1_750/B 0.03fF
C13273 POR2X1_248/O POR2X1_5/Y 0.06fF
C13274 POR2X1_260/B POR2X1_294/A 0.18fF
C13275 POR2X1_296/B POR2X1_260/A 0.22fF
C13276 POR2X1_316/Y POR2X1_20/B 0.10fF
C13277 PAND2X1_20/A PAND2X1_503/CTRL2 0.00fF
C13278 POR2X1_42/a_56_344# POR2X1_5/Y 0.00fF
C13279 POR2X1_68/A POR2X1_215/CTRL 0.01fF
C13280 INPUT_0 POR2X1_391/Y 0.10fF
C13281 POR2X1_474/O POR2X1_101/Y 0.15fF
C13282 POR2X1_860/A POR2X1_216/O 0.03fF
C13283 POR2X1_13/A PAND2X1_339/Y 0.97fF
C13284 PAND2X1_65/B POR2X1_532/A 1.48fF
C13285 PAND2X1_496/CTRL2 POR2X1_575/B 0.12fF
C13286 POR2X1_186/Y POR2X1_736/a_76_344# 0.00fF
C13287 PAND2X1_738/Y PAND2X1_566/Y 0.10fF
C13288 POR2X1_728/B POR2X1_467/CTRL2 0.03fF
C13289 PAND2X1_63/Y POR2X1_547/B 0.09fF
C13290 POR2X1_213/B POR2X1_148/A 0.21fF
C13291 PAND2X1_738/CTRL PAND2X1_149/A 0.01fF
C13292 POR2X1_403/B PAND2X1_69/A 0.03fF
C13293 POR2X1_78/B POR2X1_407/Y 0.02fF
C13294 POR2X1_822/Y POR2X1_822/O 0.00fF
C13295 PAND2X1_632/B POR2X1_482/Y 0.01fF
C13296 VDD PAND2X1_711/A 0.00fF
C13297 PAND2X1_811/Y PAND2X1_805/A 0.06fF
C13298 POR2X1_514/Y POR2X1_404/Y 0.01fF
C13299 POR2X1_66/B POR2X1_346/B 0.06fF
C13300 POR2X1_502/A POR2X1_844/B 0.05fF
C13301 PAND2X1_821/O POR2X1_857/B 0.05fF
C13302 INPUT_0 PAND2X1_548/O 0.05fF
C13303 PAND2X1_651/Y PAND2X1_573/O 0.47fF
C13304 POR2X1_137/CTRL2 POR2X1_391/Y 0.03fF
C13305 POR2X1_685/A PAND2X1_679/CTRL2 0.01fF
C13306 PAND2X1_48/B POR2X1_741/Y 0.11fF
C13307 POR2X1_388/O POR2X1_566/A 0.01fF
C13308 PAND2X1_243/CTRL2 PAND2X1_734/B 0.01fF
C13309 POR2X1_52/A POR2X1_289/O 0.01fF
C13310 POR2X1_814/B POR2X1_218/CTRL 0.01fF
C13311 PAND2X1_776/O POR2X1_238/Y 0.04fF
C13312 POR2X1_378/A POR2X1_5/Y 0.01fF
C13313 POR2X1_504/O POR2X1_14/Y 0.12fF
C13314 POR2X1_278/Y PAND2X1_341/A 0.10fF
C13315 POR2X1_186/Y PAND2X1_172/CTRL 0.01fF
C13316 POR2X1_14/Y POR2X1_394/A 0.19fF
C13317 POR2X1_37/Y POR2X1_150/O 0.00fF
C13318 POR2X1_68/A PAND2X1_441/O 0.06fF
C13319 PAND2X1_852/O POR2X1_42/Y 0.02fF
C13320 POR2X1_406/Y PAND2X1_560/CTRL 0.03fF
C13321 PAND2X1_736/A PAND2X1_675/A 0.15fF
C13322 POR2X1_614/A PAND2X1_309/O 0.01fF
C13323 PAND2X1_739/B PAND2X1_739/a_76_28# 0.02fF
C13324 POR2X1_68/A POR2X1_740/Y 0.07fF
C13325 PAND2X1_625/a_16_344# POR2X1_740/Y 0.04fF
C13326 PAND2X1_625/CTRL POR2X1_741/Y 0.08fF
C13327 PAND2X1_90/A PAND2X1_316/a_16_344# 0.01fF
C13328 PAND2X1_460/CTRL PAND2X1_472/B 0.01fF
C13329 PAND2X1_402/B POR2X1_397/Y 0.07fF
C13330 PAND2X1_857/A POR2X1_236/Y 0.07fF
C13331 POR2X1_278/Y POR2X1_91/Y 0.17fF
C13332 PAND2X1_35/Y POR2X1_229/a_16_28# 0.02fF
C13333 POR2X1_587/O POR2X1_587/Y 0.00fF
C13334 PAND2X1_188/O POR2X1_816/A 0.02fF
C13335 POR2X1_97/B POR2X1_78/A 0.62fF
C13336 PAND2X1_534/O VDD 0.00fF
C13337 POR2X1_833/O POR2X1_786/Y 0.34fF
C13338 PAND2X1_48/B PAND2X1_32/B 1.14fF
C13339 PAND2X1_785/A POR2X1_7/B 0.01fF
C13340 PAND2X1_535/a_76_28# POR2X1_236/Y 0.00fF
C13341 POR2X1_78/B POR2X1_337/A 0.03fF
C13342 POR2X1_327/Y POR2X1_269/Y 0.00fF
C13343 PAND2X1_8/O INPUT_2 0.13fF
C13344 POR2X1_537/Y POR2X1_830/Y 0.28fF
C13345 POR2X1_279/Y POR2X1_394/A 0.96fF
C13346 POR2X1_82/CTRL2 POR2X1_16/A 0.10fF
C13347 POR2X1_693/Y PAND2X1_565/A 1.77fF
C13348 POR2X1_8/Y POR2X1_376/B 0.03fF
C13349 INPUT_1 POR2X1_627/O 0.01fF
C13350 PAND2X1_434/O POR2X1_39/B 0.01fF
C13351 PAND2X1_48/B POR2X1_711/O 0.01fF
C13352 POR2X1_794/B POR2X1_737/A 0.03fF
C13353 POR2X1_60/A POR2X1_171/Y 0.05fF
C13354 POR2X1_362/Y POR2X1_362/O 0.00fF
C13355 PAND2X1_744/CTRL2 POR2X1_644/A 0.02fF
C13356 PAND2X1_845/a_76_28# POR2X1_55/Y 0.04fF
C13357 POR2X1_865/B POR2X1_572/B 0.04fF
C13358 POR2X1_471/A POR2X1_181/A 0.03fF
C13359 PAND2X1_219/O POR2X1_591/Y 0.05fF
C13360 POR2X1_66/B POR2X1_572/Y 0.02fF
C13361 PAND2X1_807/a_76_28# POR2X1_7/B 0.01fF
C13362 POR2X1_294/B POR2X1_702/CTRL 0.01fF
C13363 POR2X1_575/B POR2X1_575/CTRL2 0.08fF
C13364 POR2X1_359/B POR2X1_814/B 0.01fF
C13365 INPUT_0 POR2X1_385/a_56_344# 0.00fF
C13366 POR2X1_119/Y PAND2X1_786/O 0.19fF
C13367 PAND2X1_347/Y PAND2X1_343/O 0.04fF
C13368 POR2X1_288/A PAND2X1_48/A 0.03fF
C13369 POR2X1_408/O POR2X1_408/Y 0.00fF
C13370 PAND2X1_90/Y POR2X1_209/CTRL 0.01fF
C13371 POR2X1_38/B POR2X1_790/A 0.02fF
C13372 POR2X1_83/O PAND2X1_734/B 0.01fF
C13373 POR2X1_57/A POR2X1_396/CTRL 0.01fF
C13374 PAND2X1_90/Y POR2X1_186/B 0.09fF
C13375 VDD POR2X1_210/B 0.00fF
C13376 PAND2X1_40/O POR2X1_407/Y 0.01fF
C13377 POR2X1_119/Y POR2X1_72/B 0.12fF
C13378 POR2X1_65/A POR2X1_62/Y 0.03fF
C13379 PAND2X1_6/Y POR2X1_341/Y 0.03fF
C13380 POR2X1_68/A PAND2X1_312/CTRL2 0.01fF
C13381 D_INPUT_1 POR2X1_550/CTRL2 0.01fF
C13382 PAND2X1_737/B POR2X1_46/Y 0.51fF
C13383 PAND2X1_206/CTRL POR2X1_153/Y 0.08fF
C13384 PAND2X1_359/O PAND2X1_359/B 0.00fF
C13385 POR2X1_417/Y PAND2X1_352/O 0.03fF
C13386 PAND2X1_865/Y PAND2X1_354/A 0.07fF
C13387 POR2X1_377/O POR2X1_378/A 0.02fF
C13388 PAND2X1_716/CTRL2 PAND2X1_656/A 0.01fF
C13389 POR2X1_16/A PAND2X1_776/CTRL2 0.01fF
C13390 PAND2X1_812/A PAND2X1_805/A 0.03fF
C13391 POR2X1_68/A POR2X1_348/O 0.04fF
C13392 PAND2X1_414/O POR2X1_67/Y 0.02fF
C13393 PAND2X1_292/O POR2X1_66/A 0.02fF
C13394 PAND2X1_48/B POR2X1_543/CTRL2 0.01fF
C13395 POR2X1_317/m4_208_n4# POR2X1_854/B 0.04fF
C13396 PAND2X1_568/B PAND2X1_578/A 0.01fF
C13397 PAND2X1_241/Y POR2X1_90/Y 0.01fF
C13398 PAND2X1_598/CTRL POR2X1_394/A 0.06fF
C13399 POR2X1_703/A PAND2X1_176/a_16_344# 0.03fF
C13400 PAND2X1_316/m4_208_n4# POR2X1_318/A 0.09fF
C13401 POR2X1_52/A POR2X1_8/Y 0.08fF
C13402 PAND2X1_714/Y PAND2X1_724/B 0.01fF
C13403 PAND2X1_329/CTRL2 PAND2X1_69/A 0.01fF
C13404 PAND2X1_430/O PAND2X1_3/B 0.10fF
C13405 POR2X1_46/Y POR2X1_117/m4_208_n4# 0.07fF
C13406 PAND2X1_539/Y POR2X1_42/Y 0.03fF
C13407 PAND2X1_472/B POR2X1_394/A 0.10fF
C13408 POR2X1_131/CTRL PAND2X1_349/A 0.01fF
C13409 POR2X1_390/B PAND2X1_56/Y 0.03fF
C13410 POR2X1_43/B PAND2X1_124/CTRL 0.01fF
C13411 PAND2X1_117/CTRL2 POR2X1_557/B 0.00fF
C13412 PAND2X1_137/Y POR2X1_103/a_16_28# 0.03fF
C13413 POR2X1_504/O POR2X1_55/Y 0.01fF
C13414 PAND2X1_714/A PAND2X1_169/CTRL 0.04fF
C13415 POR2X1_394/A POR2X1_55/Y 0.15fF
C13416 POR2X1_840/B POR2X1_569/A 0.10fF
C13417 POR2X1_613/Y VDD 0.12fF
C13418 PAND2X1_8/Y POR2X1_4/Y 0.30fF
C13419 POR2X1_42/Y PAND2X1_507/O 0.13fF
C13420 POR2X1_57/A POR2X1_96/B 0.07fF
C13421 POR2X1_383/A POR2X1_493/CTRL2 0.01fF
C13422 POR2X1_416/B PAND2X1_742/a_16_344# 0.02fF
C13423 PAND2X1_480/CTRL POR2X1_43/B 0.01fF
C13424 POR2X1_274/B POR2X1_724/A 0.02fF
C13425 POR2X1_93/a_16_28# POR2X1_503/Y 0.02fF
C13426 VDD PAND2X1_517/CTRL 0.00fF
C13427 POR2X1_416/B POR2X1_24/O 0.02fF
C13428 VDD POR2X1_181/CTRL 0.00fF
C13429 POR2X1_52/A POR2X1_385/Y 0.15fF
C13430 PAND2X1_610/O VDD 0.00fF
C13431 POR2X1_20/CTRL2 POR2X1_4/Y 0.06fF
C13432 POR2X1_3/CTRL POR2X1_260/A 0.05fF
C13433 POR2X1_540/A POR2X1_456/B 0.74fF
C13434 POR2X1_508/A POR2X1_579/Y 0.03fF
C13435 POR2X1_122/Y POR2X1_39/B 0.26fF
C13436 PAND2X1_23/Y PAND2X1_171/a_16_344# 0.01fF
C13437 POR2X1_760/A PAND2X1_217/O 0.05fF
C13438 POR2X1_584/a_16_28# POR2X1_260/A 0.01fF
C13439 PAND2X1_55/Y POR2X1_294/A 0.15fF
C13440 PAND2X1_551/CTRL2 PAND2X1_569/B 0.00fF
C13441 POR2X1_244/Y POR2X1_702/A 0.03fF
C13442 INPUT_0 POR2X1_383/Y 0.53fF
C13443 PAND2X1_631/A POR2X1_252/O 0.16fF
C13444 POR2X1_327/Y POR2X1_513/Y 0.06fF
C13445 PAND2X1_423/CTRL PAND2X1_72/A 0.01fF
C13446 POR2X1_556/A POR2X1_658/a_16_28# 0.00fF
C13447 PAND2X1_612/a_16_344# POR2X1_472/B 0.02fF
C13448 POR2X1_68/A POR2X1_550/B 0.01fF
C13449 POR2X1_463/Y PAND2X1_60/B 0.03fF
C13450 POR2X1_254/Y POR2X1_632/Y 0.07fF
C13451 POR2X1_390/B POR2X1_383/A 0.03fF
C13452 POR2X1_409/Y POR2X1_380/Y 0.25fF
C13453 POR2X1_793/CTRL2 PAND2X1_52/B 0.01fF
C13454 POR2X1_311/Y PAND2X1_221/Y 0.06fF
C13455 POR2X1_5/Y POR2X1_80/a_76_344# 0.01fF
C13456 PAND2X1_684/m4_208_n4# PAND2X1_421/m4_208_n4# 0.13fF
C13457 PAND2X1_96/B POR2X1_557/B 0.04fF
C13458 INPUT_0 POR2X1_77/Y 0.32fF
C13459 POR2X1_379/Y PAND2X1_752/Y 0.24fF
C13460 POR2X1_547/a_16_28# POR2X1_266/A 0.02fF
C13461 PAND2X1_294/O POR2X1_150/Y 0.05fF
C13462 POR2X1_539/A POR2X1_456/B 0.03fF
C13463 POR2X1_305/Y PAND2X1_506/Y 0.02fF
C13464 POR2X1_54/Y POR2X1_20/B 0.03fF
C13465 POR2X1_814/A POR2X1_66/A 0.19fF
C13466 POR2X1_305/a_16_28# POR2X1_39/B 0.03fF
C13467 POR2X1_326/O POR2X1_854/B 0.18fF
C13468 POR2X1_760/A PAND2X1_124/Y 0.04fF
C13469 POR2X1_52/O PAND2X1_215/B 0.03fF
C13470 PAND2X1_187/O POR2X1_444/Y 0.02fF
C13471 POR2X1_416/B PAND2X1_480/B 0.03fF
C13472 POR2X1_579/Y POR2X1_568/B 24.79fF
C13473 PAND2X1_213/Y POR2X1_373/Y 0.03fF
C13474 POR2X1_407/Y POR2X1_294/A 0.03fF
C13475 POR2X1_119/Y PAND2X1_835/Y 0.01fF
C13476 POR2X1_424/O POR2X1_77/Y 0.00fF
C13477 POR2X1_3/A PAND2X1_18/B 0.17fF
C13478 POR2X1_564/Y POR2X1_180/Y 0.02fF
C13479 POR2X1_327/Y POR2X1_366/A 1.27fF
C13480 POR2X1_257/A POR2X1_428/Y 0.03fF
C13481 PAND2X1_634/CTRL2 POR2X1_48/A 0.03fF
C13482 POR2X1_505/O PAND2X1_632/B 0.01fF
C13483 POR2X1_20/B POR2X1_298/O 0.17fF
C13484 POR2X1_545/A POR2X1_568/B 0.03fF
C13485 POR2X1_163/A POR2X1_158/Y 0.00fF
C13486 POR2X1_110/Y PAND2X1_241/Y 0.03fF
C13487 PAND2X1_713/O PAND2X1_713/A -0.00fF
C13488 PAND2X1_175/CTRL2 PAND2X1_853/B 0.01fF
C13489 POR2X1_244/B POR2X1_568/A 0.05fF
C13490 PAND2X1_717/A POR2X1_102/Y 0.07fF
C13491 POR2X1_503/O POR2X1_8/Y 0.23fF
C13492 POR2X1_681/CTRL2 POR2X1_60/A 0.01fF
C13493 POR2X1_43/O POR2X1_43/B 0.02fF
C13494 POR2X1_614/A POR2X1_568/B 0.05fF
C13495 D_INPUT_3 POR2X1_5/a_16_28# 0.03fF
C13496 POR2X1_499/CTRL POR2X1_341/A 0.06fF
C13497 POR2X1_760/A POR2X1_83/B 0.15fF
C13498 PAND2X1_631/A POR2X1_245/Y 0.03fF
C13499 POR2X1_837/O POR2X1_837/A 0.02fF
C13500 POR2X1_811/O PAND2X1_39/B 0.12fF
C13501 POR2X1_287/B POR2X1_458/Y 0.04fF
C13502 PAND2X1_844/CTRL POR2X1_153/Y 0.28fF
C13503 POR2X1_14/Y PAND2X1_33/CTRL2 0.00fF
C13504 POR2X1_257/A POR2X1_432/CTRL2 0.03fF
C13505 POR2X1_52/A POR2X1_91/CTRL2 0.01fF
C13506 POR2X1_43/B PAND2X1_332/Y 0.03fF
C13507 POR2X1_60/A POR2X1_150/Y 0.25fF
C13508 PAND2X1_687/A POR2X1_761/A 0.06fF
C13509 POR2X1_68/A POR2X1_87/B 0.01fF
C13510 POR2X1_48/A PAND2X1_645/Y 0.01fF
C13511 POR2X1_411/B POR2X1_609/CTRL2 0.02fF
C13512 PAND2X1_156/A PAND2X1_156/B 0.03fF
C13513 PAND2X1_601/a_76_28# D_INPUT_0 0.02fF
C13514 POR2X1_840/B PAND2X1_72/A 0.33fF
C13515 POR2X1_673/Y PAND2X1_517/CTRL 0.28fF
C13516 POR2X1_341/Y PAND2X1_52/B 0.03fF
C13517 POR2X1_329/A POR2X1_236/Y 0.17fF
C13518 POR2X1_440/Y POR2X1_568/B 0.05fF
C13519 POR2X1_129/Y PAND2X1_851/O 0.02fF
C13520 POR2X1_859/CTRL2 PAND2X1_41/B 0.03fF
C13521 POR2X1_188/A POR2X1_841/CTRL 0.01fF
C13522 PAND2X1_66/O POR2X1_67/A 0.07fF
C13523 PAND2X1_39/B POR2X1_330/Y 0.17fF
C13524 POR2X1_673/Y PAND2X1_529/CTRL2 0.03fF
C13525 POR2X1_95/O POR2X1_394/A 0.08fF
C13526 POR2X1_519/CTRL2 POR2X1_416/B 0.01fF
C13527 PAND2X1_60/B POR2X1_500/O 0.04fF
C13528 POR2X1_49/Y INPUT_3 0.29fF
C13529 POR2X1_736/A POR2X1_737/CTRL 0.03fF
C13530 PAND2X1_404/Y PAND2X1_404/O 0.01fF
C13531 PAND2X1_265/O POR2X1_260/B 0.02fF
C13532 POR2X1_567/B POR2X1_174/A 0.05fF
C13533 POR2X1_327/Y POR2X1_532/CTRL2 0.17fF
C13534 POR2X1_635/A POR2X1_750/B 2.15fF
C13535 POR2X1_153/Y PAND2X1_860/O 0.11fF
C13536 POR2X1_130/CTRL2 POR2X1_343/Y 0.00fF
C13537 POR2X1_445/A POR2X1_186/Y 0.03fF
C13538 POR2X1_78/A POR2X1_466/A 0.72fF
C13539 POR2X1_399/O POR2X1_411/B 0.01fF
C13540 POR2X1_805/Y POR2X1_792/CTRL2 0.01fF
C13541 PAND2X1_435/CTRL2 POR2X1_271/B 0.01fF
C13542 POR2X1_663/O POR2X1_663/B 0.04fF
C13543 PAND2X1_97/Y PAND2X1_351/O 0.02fF
C13544 POR2X1_329/a_16_28# POR2X1_250/Y 0.05fF
C13545 PAND2X1_404/Y PAND2X1_61/Y 0.03fF
C13546 PAND2X1_472/B PAND2X1_33/CTRL2 0.02fF
C13547 POR2X1_777/B POR2X1_458/O 0.06fF
C13548 POR2X1_814/A POR2X1_222/Y 0.07fF
C13549 POR2X1_14/Y POR2X1_669/B 0.43fF
C13550 POR2X1_76/B POR2X1_575/O 0.13fF
C13551 PAND2X1_508/Y POR2X1_39/B 0.04fF
C13552 POR2X1_658/CTRL2 POR2X1_193/A 0.04fF
C13553 POR2X1_34/A POR2X1_34/Y 0.00fF
C13554 PAND2X1_52/B POR2X1_731/A 0.13fF
C13555 D_INPUT_5 POR2X1_25/a_56_344# 0.01fF
C13556 POR2X1_12/A POR2X1_25/O 0.00fF
C13557 PAND2X1_798/Y PAND2X1_366/a_76_28# 0.03fF
C13558 D_INPUT_5 VDD 1.19fF
C13559 PAND2X1_91/a_16_344# PAND2X1_90/Y 0.02fF
C13560 POR2X1_311/Y POR2X1_83/B 0.03fF
C13561 POR2X1_67/O POR2X1_236/Y 0.01fF
C13562 PAND2X1_679/O POR2X1_678/Y 0.00fF
C13563 POR2X1_43/B POR2X1_262/m4_208_n4# 0.04fF
C13564 PAND2X1_205/a_16_344# PAND2X1_473/B 0.02fF
C13565 POR2X1_60/A PAND2X1_794/O 0.03fF
C13566 PAND2X1_404/Y PAND2X1_404/A 0.02fF
C13567 PAND2X1_23/Y POR2X1_556/A 0.17fF
C13568 POR2X1_827/Y VDD 0.00fF
C13569 POR2X1_193/A POR2X1_341/A 0.07fF
C13570 POR2X1_210/A PAND2X1_72/A 0.00fF
C13571 PAND2X1_48/B PAND2X1_9/Y 3.62fF
C13572 POR2X1_341/A POR2X1_579/Y 0.09fF
C13573 POR2X1_796/Y VDD 0.29fF
C13574 POR2X1_814/A POR2X1_532/A 0.29fF
C13575 POR2X1_707/B POR2X1_634/A 0.03fF
C13576 PAND2X1_613/a_16_344# PAND2X1_8/Y 0.05fF
C13577 POR2X1_260/B PAND2X1_378/CTRL 0.03fF
C13578 POR2X1_644/CTRL PAND2X1_57/B 0.01fF
C13579 PAND2X1_31/CTRL VDD -0.00fF
C13580 POR2X1_96/A POR2X1_79/O 0.00fF
C13581 POR2X1_660/Y POR2X1_660/A 0.02fF
C13582 PAND2X1_20/A POR2X1_330/Y 0.05fF
C13583 PAND2X1_75/CTRL POR2X1_532/A 0.01fF
C13584 PAND2X1_331/a_76_28# POR2X1_330/Y 0.01fF
C13585 POR2X1_291/a_16_28# POR2X1_234/A 0.04fF
C13586 POR2X1_51/A POR2X1_260/B 0.02fF
C13587 POR2X1_241/B POR2X1_254/a_56_344# 0.00fF
C13588 POR2X1_718/A POR2X1_296/B 0.07fF
C13589 POR2X1_285/CTRL2 POR2X1_590/A 0.01fF
C13590 POR2X1_302/B POR2X1_794/B 0.02fF
C13591 PAND2X1_248/CTRL2 POR2X1_404/Y 0.03fF
C13592 POR2X1_78/a_16_28# POR2X1_844/B 0.02fF
C13593 PAND2X1_669/O VDD 0.00fF
C13594 POR2X1_718/m4_208_n4# D_INPUT_0 0.12fF
C13595 PAND2X1_216/O PAND2X1_218/B 0.05fF
C13596 POR2X1_470/CTRL VDD 0.00fF
C13597 POR2X1_257/A PAND2X1_469/B 0.12fF
C13598 POR2X1_413/Y POR2X1_612/Y 0.03fF
C13599 POR2X1_23/Y PAND2X1_254/Y 0.06fF
C13600 POR2X1_29/O POR2X1_29/A 0.01fF
C13601 POR2X1_655/A PAND2X1_385/O 0.15fF
C13602 POR2X1_411/CTRL2 POR2X1_37/Y 0.03fF
C13603 POR2X1_614/A POR2X1_341/A 0.02fF
C13604 POR2X1_78/B POR2X1_174/A 0.07fF
C13605 POR2X1_97/A POR2X1_192/Y 0.05fF
C13606 POR2X1_9/Y PAND2X1_341/Y 0.10fF
C13607 POR2X1_814/B POR2X1_330/Y 0.05fF
C13608 PAND2X1_96/B PAND2X1_43/CTRL 0.05fF
C13609 PAND2X1_75/m4_208_n4# POR2X1_724/A 0.12fF
C13610 POR2X1_624/Y POR2X1_140/A 0.03fF
C13611 PAND2X1_48/B POR2X1_818/Y 0.03fF
C13612 INPUT_1 POR2X1_624/O 0.01fF
C13613 POR2X1_632/B VDD 0.01fF
C13614 POR2X1_78/A POR2X1_608/O 0.03fF
C13615 PAND2X1_73/Y POR2X1_608/a_56_344# 0.00fF
C13616 POR2X1_65/A PAND2X1_349/B 0.07fF
C13617 POR2X1_866/A POR2X1_800/A 0.05fF
C13618 POR2X1_102/Y PAND2X1_778/a_16_344# 0.01fF
C13619 POR2X1_516/Y VDD 0.20fF
C13620 POR2X1_60/A POR2X1_701/Y 0.07fF
C13621 PAND2X1_270/CTRL POR2X1_20/B 0.01fF
C13622 PAND2X1_787/A POR2X1_20/B 0.90fF
C13623 POR2X1_41/B POR2X1_309/CTRL2 0.01fF
C13624 D_INPUT_5 PAND2X1_32/B 0.05fF
C13625 PAND2X1_109/O PAND2X1_52/B 0.02fF
C13626 POR2X1_502/A POR2X1_241/B 0.03fF
C13627 PAND2X1_85/O POR2X1_260/A 0.09fF
C13628 POR2X1_423/Y POR2X1_5/Y 0.04fF
C13629 PAND2X1_58/A PAND2X1_56/CTRL 0.01fF
C13630 POR2X1_861/O POR2X1_558/B 0.00fF
C13631 POR2X1_330/Y POR2X1_325/A 0.05fF
C13632 POR2X1_23/Y POR2X1_599/A 0.05fF
C13633 POR2X1_629/CTRL2 PAND2X1_69/A 0.00fF
C13634 POR2X1_43/B PAND2X1_97/O 0.02fF
C13635 POR2X1_149/B PAND2X1_93/B 0.02fF
C13636 POR2X1_63/Y POR2X1_235/CTRL2 0.01fF
C13637 POR2X1_454/A POR2X1_556/Y 0.03fF
C13638 POR2X1_774/Y POR2X1_866/B 0.01fF
C13639 POR2X1_38/CTRL2 POR2X1_38/B 0.01fF
C13640 POR2X1_645/a_76_344# POR2X1_330/Y 0.03fF
C13641 POR2X1_41/B POR2X1_102/Y 0.13fF
C13642 PAND2X1_96/B PAND2X1_406/CTRL 0.01fF
C13643 POR2X1_502/A POR2X1_719/A 0.02fF
C13644 PAND2X1_72/A PAND2X1_56/A 0.05fF
C13645 POR2X1_460/Y PAND2X1_376/CTRL2 0.01fF
C13646 POR2X1_133/CTRL POR2X1_40/Y 0.01fF
C13647 POR2X1_814/B POR2X1_116/O 0.08fF
C13648 POR2X1_669/B POR2X1_55/Y 0.32fF
C13649 POR2X1_165/Y PAND2X1_717/A 0.13fF
C13650 POR2X1_271/A POR2X1_329/A 0.00fF
C13651 POR2X1_78/B PAND2X1_16/CTRL 0.01fF
C13652 POR2X1_32/O POR2X1_32/A 0.02fF
C13653 PAND2X1_798/B POR2X1_487/CTRL2 0.05fF
C13654 PAND2X1_785/m4_208_n4# POR2X1_91/Y 0.12fF
C13655 POR2X1_411/B PAND2X1_181/O 0.04fF
C13656 PAND2X1_48/B PAND2X1_15/O 0.05fF
C13657 PAND2X1_93/B POR2X1_219/CTRL 0.01fF
C13658 POR2X1_722/A POR2X1_648/Y 0.07fF
C13659 POR2X1_60/A PAND2X1_364/B 0.07fF
C13660 POR2X1_702/B POR2X1_483/A 0.02fF
C13661 POR2X1_688/O POR2X1_260/A 0.02fF
C13662 POR2X1_130/A POR2X1_862/B 0.05fF
C13663 POR2X1_38/Y PAND2X1_124/Y 0.03fF
C13664 PAND2X1_581/O INPUT_6 0.01fF
C13665 POR2X1_212/A POR2X1_212/O 0.04fF
C13666 POR2X1_389/A POR2X1_260/B 0.05fF
C13667 POR2X1_427/Y POR2X1_763/a_16_28# 0.00fF
C13668 PAND2X1_206/A POR2X1_7/A 0.04fF
C13669 POR2X1_76/CTRL2 POR2X1_569/A 0.05fF
C13670 PAND2X1_58/A POR2X1_740/Y 0.03fF
C13671 POR2X1_330/Y POR2X1_513/B 0.05fF
C13672 POR2X1_94/CTRL2 POR2X1_14/Y 0.00fF
C13673 PAND2X1_790/O POR2X1_7/A 0.11fF
C13674 PAND2X1_794/CTRL2 PAND2X1_794/B 0.01fF
C13675 POR2X1_97/A POR2X1_502/m4_208_n4# 0.10fF
C13676 POR2X1_368/CTRL POR2X1_5/Y 0.01fF
C13677 POR2X1_548/CTRL PAND2X1_8/Y 0.01fF
C13678 POR2X1_65/A PAND2X1_549/O 0.01fF
C13679 POR2X1_590/A POR2X1_790/A 0.01fF
C13680 POR2X1_149/B POR2X1_78/A 0.78fF
C13681 POR2X1_51/B POR2X1_12/A 0.03fF
C13682 PAND2X1_619/CTRL POR2X1_260/A 0.03fF
C13683 POR2X1_333/A POR2X1_775/A 0.20fF
C13684 D_INPUT_0 PAND2X1_79/Y 0.01fF
C13685 PAND2X1_667/CTRL VDD -0.00fF
C13686 POR2X1_717/B POR2X1_343/B 0.00fF
C13687 POR2X1_130/CTRL2 POR2X1_624/Y 0.00fF
C13688 POR2X1_722/Y POR2X1_830/A 0.03fF
C13689 PAND2X1_55/Y POR2X1_94/A 0.03fF
C13690 POR2X1_834/Y POR2X1_648/O 0.16fF
C13691 POR2X1_673/CTRL2 PAND2X1_6/A 0.05fF
C13692 POR2X1_673/A PAND2X1_8/Y 0.02fF
C13693 POR2X1_65/A POR2X1_597/A 0.03fF
C13694 PAND2X1_23/Y POR2X1_202/O 0.00fF
C13695 POR2X1_596/A POR2X1_770/B 0.01fF
C13696 POR2X1_814/B POR2X1_247/O 0.11fF
C13697 POR2X1_78/A POR2X1_649/CTRL 0.00fF
C13698 POR2X1_31/m4_208_n4# POR2X1_12/A 0.12fF
C13699 PAND2X1_798/B POR2X1_40/Y 0.07fF
C13700 POR2X1_482/CTRL2 POR2X1_7/A 0.00fF
C13701 POR2X1_514/a_76_344# PAND2X1_20/A 0.00fF
C13702 PAND2X1_653/Y PAND2X1_219/A 0.03fF
C13703 POR2X1_626/O POR2X1_408/Y 0.02fF
C13704 POR2X1_865/B POR2X1_590/A 5.09fF
C13705 POR2X1_590/A PAND2X1_88/Y 0.01fF
C13706 POR2X1_41/B PAND2X1_192/a_16_344# 0.01fF
C13707 POR2X1_467/CTRL2 POR2X1_330/Y 0.02fF
C13708 D_INPUT_0 PAND2X1_656/A 0.05fF
C13709 POR2X1_728/B VDD 0.05fF
C13710 POR2X1_68/A POR2X1_202/CTRL 0.01fF
C13711 PAND2X1_164/CTRL POR2X1_776/B 0.01fF
C13712 PAND2X1_20/A PAND2X1_519/a_76_28# 0.02fF
C13713 PAND2X1_579/B PAND2X1_735/Y 0.07fF
C13714 POR2X1_852/B POR2X1_222/Y 0.07fF
C13715 POR2X1_83/B POR2X1_38/Y 0.31fF
C13716 POR2X1_49/Y PAND2X1_469/B 0.01fF
C13717 POR2X1_79/Y PAND2X1_739/Y 0.02fF
C13718 POR2X1_502/A PAND2X1_438/CTRL2 0.01fF
C13719 POR2X1_814/A PAND2X1_122/a_56_28# 0.00fF
C13720 PAND2X1_656/O PAND2X1_656/A 0.01fF
C13721 PAND2X1_211/A PAND2X1_357/Y 0.00fF
C13722 POR2X1_22/A POR2X1_12/O 0.01fF
C13723 POR2X1_262/Y POR2X1_7/Y 0.01fF
C13724 POR2X1_5/Y POR2X1_57/Y 0.01fF
C13725 PAND2X1_6/Y PAND2X1_41/B 0.12fF
C13726 POR2X1_114/B POR2X1_405/a_76_344# 0.00fF
C13727 PAND2X1_832/CTRL2 PAND2X1_651/Y 0.47fF
C13728 POR2X1_97/A POR2X1_568/Y 0.05fF
C13729 POR2X1_74/O POR2X1_23/Y 0.15fF
C13730 PAND2X1_288/A GATE_741 0.03fF
C13731 POR2X1_448/O PAND2X1_60/B 0.17fF
C13732 PAND2X1_216/B PAND2X1_571/A 0.02fF
C13733 POR2X1_296/B POR2X1_725/Y 0.10fF
C13734 PAND2X1_23/Y POR2X1_400/A 0.03fF
C13735 POR2X1_20/B POR2X1_4/Y 0.31fF
C13736 PAND2X1_488/CTRL2 POR2X1_532/A 0.33fF
C13737 POR2X1_22/O INPUT_5 0.17fF
C13738 D_INPUT_7 PAND2X1_52/B 0.48fF
C13739 PAND2X1_579/B PAND2X1_493/Y 0.70fF
C13740 POR2X1_98/CTRL2 POR2X1_260/A 0.02fF
C13741 POR2X1_634/A POR2X1_711/a_16_28# 0.11fF
C13742 POR2X1_333/A POR2X1_162/Y 0.14fF
C13743 POR2X1_856/B POR2X1_703/Y 0.03fF
C13744 PAND2X1_124/Y POR2X1_153/Y 0.07fF
C13745 POR2X1_14/Y POR2X1_750/m4_208_n4# 0.08fF
C13746 POR2X1_92/CTRL2 POR2X1_49/Y 0.01fF
C13747 POR2X1_433/O PAND2X1_549/B 0.01fF
C13748 PAND2X1_661/B POR2X1_117/CTRL 0.01fF
C13749 POR2X1_242/a_16_28# PAND2X1_32/B 0.01fF
C13750 PAND2X1_697/O PAND2X1_65/B 0.03fF
C13751 POR2X1_192/Y POR2X1_294/B 0.05fF
C13752 POR2X1_366/Y POR2X1_192/Y 0.10fF
C13753 PAND2X1_56/Y POR2X1_370/Y 0.03fF
C13754 POR2X1_106/Y POR2X1_90/Y 0.03fF
C13755 POR2X1_857/B POR2X1_853/O 0.00fF
C13756 POR2X1_43/B PAND2X1_474/Y 0.04fF
C13757 POR2X1_270/Y POR2X1_370/CTRL2 0.03fF
C13758 POR2X1_43/B PAND2X1_715/CTRL 0.01fF
C13759 PAND2X1_61/Y POR2X1_521/a_16_28# 0.02fF
C13760 POR2X1_96/A POR2X1_697/Y 0.03fF
C13761 POR2X1_647/O POR2X1_737/A 0.02fF
C13762 D_INPUT_0 PAND2X1_348/A 0.13fF
C13763 PAND2X1_309/CTRL2 POR2X1_740/Y 0.34fF
C13764 POR2X1_94/CTRL2 PAND2X1_472/B 0.04fF
C13765 POR2X1_778/B POR2X1_778/O 0.01fF
C13766 POR2X1_270/a_16_28# POR2X1_186/Y 0.01fF
C13767 POR2X1_65/A PAND2X1_650/CTRL 0.00fF
C13768 POR2X1_43/B POR2X1_13/A 3.12fF
C13769 POR2X1_48/A PAND2X1_508/Y 0.03fF
C13770 POR2X1_273/Y PAND2X1_480/B 0.20fF
C13771 PAND2X1_723/CTRL VDD 0.00fF
C13772 INPUT_1 POR2X1_83/B 0.14fF
C13773 POR2X1_616/Y PAND2X1_66/O 0.04fF
C13774 PAND2X1_190/O POR2X1_184/Y 0.00fF
C13775 POR2X1_131/CTRL2 POR2X1_13/A 0.00fF
C13776 PAND2X1_685/a_76_28# INPUT_0 0.02fF
C13777 D_INPUT_1 PAND2X1_8/Y 0.15fF
C13778 PAND2X1_56/Y PAND2X1_309/CTRL 0.01fF
C13779 D_INPUT_0 POR2X1_300/Y 0.03fF
C13780 PAND2X1_842/O PAND2X1_388/Y 0.05fF
C13781 POR2X1_96/A PAND2X1_357/Y 0.06fF
C13782 PAND2X1_831/Y PAND2X1_76/Y 0.03fF
C13783 PAND2X1_90/Y POR2X1_736/O 0.02fF
C13784 PAND2X1_483/O POR2X1_60/A 0.02fF
C13785 POR2X1_68/A PAND2X1_293/m4_208_n4# 0.07fF
C13786 POR2X1_48/A POR2X1_320/CTRL 0.01fF
C13787 POR2X1_102/Y PAND2X1_308/Y 0.05fF
C13788 PAND2X1_691/Y POR2X1_40/Y 0.03fF
C13789 PAND2X1_675/A PAND2X1_553/B 0.07fF
C13790 POR2X1_57/A POR2X1_236/Y 0.22fF
C13791 PAND2X1_469/B PAND2X1_553/B 0.10fF
C13792 POR2X1_41/B PAND2X1_845/CTRL 0.00fF
C13793 POR2X1_119/Y PAND2X1_640/B 0.07fF
C13794 PAND2X1_51/CTRL2 POR2X1_750/B 0.01fF
C13795 PAND2X1_801/B PAND2X1_854/A 0.25fF
C13796 PAND2X1_6/A POR2X1_7/B 4.93fF
C13797 POR2X1_376/B PAND2X1_550/Y 0.00fF
C13798 PAND2X1_735/Y POR2X1_73/Y 0.07fF
C13799 POR2X1_83/B POR2X1_153/Y 5.71fF
C13800 POR2X1_13/A POR2X1_38/B 0.03fF
C13801 POR2X1_20/CTRL2 D_INPUT_1 0.03fF
C13802 POR2X1_832/A POR2X1_480/A 0.09fF
C13803 POR2X1_83/B POR2X1_384/A 0.06fF
C13804 POR2X1_463/Y POR2X1_750/B 0.01fF
C13805 POR2X1_66/B POR2X1_507/A 0.01fF
C13806 POR2X1_724/CTRL POR2X1_724/A 0.01fF
C13807 PAND2X1_296/CTRL2 PAND2X1_359/Y 0.01fF
C13808 PAND2X1_58/A POR2X1_774/A 0.03fF
C13809 POR2X1_133/O POR2X1_93/A 0.01fF
C13810 POR2X1_283/A PAND2X1_499/Y 0.04fF
C13811 INPUT_1 POR2X1_752/Y 0.03fF
C13812 POR2X1_186/Y POR2X1_260/A 0.03fF
C13813 POR2X1_584/O POR2X1_42/Y 0.03fF
C13814 POR2X1_41/B POR2X1_821/Y 0.03fF
C13815 VDD PAND2X1_843/Y 0.00fF
C13816 PAND2X1_631/A D_INPUT_0 0.17fF
C13817 PAND2X1_604/CTRL PAND2X1_69/A 0.01fF
C13818 POR2X1_719/CTRL POR2X1_502/A -0.01fF
C13819 POR2X1_433/Y PAND2X1_658/B 0.05fF
C13820 PAND2X1_340/B POR2X1_77/Y 0.03fF
C13821 PAND2X1_58/A POR2X1_550/B 0.02fF
C13822 POR2X1_548/a_16_28# POR2X1_548/A 0.07fF
C13823 PAND2X1_350/a_16_344# INPUT_0 0.00fF
C13824 PAND2X1_79/CTRL POR2X1_844/B 0.01fF
C13825 POR2X1_136/Y PAND2X1_480/B 0.05fF
C13826 POR2X1_578/Y POR2X1_577/O 0.00fF
C13827 PAND2X1_6/Y POR2X1_130/Y 0.67fF
C13828 POR2X1_96/A PAND2X1_344/a_16_344# 0.01fF
C13829 POR2X1_566/A POR2X1_510/Y 0.05fF
C13830 PAND2X1_717/A POR2X1_677/Y 0.09fF
C13831 PAND2X1_202/CTRL POR2X1_7/A 0.01fF
C13832 POR2X1_218/CTRL VDD 0.00fF
C13833 POR2X1_86/CTRL D_INPUT_0 0.01fF
C13834 PAND2X1_48/B POR2X1_639/Y 0.12fF
C13835 POR2X1_335/A POR2X1_513/Y 0.05fF
C13836 POR2X1_562/CTRL2 POR2X1_341/Y 0.01fF
C13837 POR2X1_16/A PAND2X1_403/Y 0.01fF
C13838 POR2X1_740/Y PAND2X1_111/a_76_28# 0.06fF
C13839 POR2X1_102/Y PAND2X1_141/CTRL 0.01fF
C13840 PAND2X1_140/A POR2X1_96/A 0.00fF
C13841 PAND2X1_707/Y PAND2X1_705/a_76_28# 0.07fF
C13842 PAND2X1_96/B POR2X1_740/Y 0.16fF
C13843 POR2X1_345/A POR2X1_334/Y 0.04fF
C13844 VDD PAND2X1_114/CTRL -0.00fF
C13845 POR2X1_728/CTRL2 POR2X1_730/Y 0.01fF
C13846 POR2X1_528/Y POR2X1_96/A 0.10fF
C13847 POR2X1_382/Y POR2X1_42/Y 0.38fF
C13848 POR2X1_78/A PAND2X1_179/CTRL2 0.03fF
C13849 POR2X1_40/Y POR2X1_599/a_76_344# 0.01fF
C13850 POR2X1_659/CTRL2 POR2X1_724/A 0.03fF
C13851 POR2X1_72/B POR2X1_371/CTRL2 0.03fF
C13852 POR2X1_315/CTRL POR2X1_90/Y 0.01fF
C13853 PAND2X1_661/B POR2X1_43/B 0.05fF
C13854 POR2X1_193/a_76_344# POR2X1_631/B 0.00fF
C13855 PAND2X1_687/A POR2X1_829/A 0.00fF
C13856 POR2X1_130/A POR2X1_276/Y 0.06fF
C13857 POR2X1_68/A POR2X1_196/Y 0.03fF
C13858 PAND2X1_834/O POR2X1_37/Y 0.04fF
C13859 POR2X1_56/B PAND2X1_549/B 0.07fF
C13860 PAND2X1_117/CTRL POR2X1_383/A 0.01fF
C13861 PAND2X1_41/B POR2X1_195/O 0.01fF
C13862 PAND2X1_491/CTRL2 PAND2X1_96/B 0.01fF
C13863 POR2X1_179/CTRL2 POR2X1_142/Y 0.01fF
C13864 POR2X1_588/Y POR2X1_7/B 0.01fF
C13865 PAND2X1_482/CTRL2 POR2X1_483/A 0.01fF
C13866 POR2X1_219/O POR2X1_631/B 0.02fF
C13867 POR2X1_614/A PAND2X1_495/CTRL 0.03fF
C13868 POR2X1_57/A PAND2X1_850/O 0.01fF
C13869 POR2X1_319/A POR2X1_568/A 0.03fF
C13870 POR2X1_590/A POR2X1_568/B 0.08fF
C13871 PAND2X1_23/Y PAND2X1_393/O 0.06fF
C13872 POR2X1_730/Y POR2X1_220/Y 0.89fF
C13873 POR2X1_860/A POR2X1_294/A 0.03fF
C13874 POR2X1_394/A POR2X1_524/Y 0.03fF
C13875 PAND2X1_23/Y POR2X1_276/A 0.03fF
C13876 POR2X1_814/B POR2X1_703/O 0.01fF
C13877 POR2X1_65/A PAND2X1_779/O 0.01fF
C13878 PAND2X1_220/Y PAND2X1_730/A 0.00fF
C13879 PAND2X1_6/Y POR2X1_686/O 0.01fF
C13880 PAND2X1_23/Y POR2X1_566/B 0.03fF
C13881 POR2X1_96/A POR2X1_96/O 0.02fF
C13882 POR2X1_7/B PAND2X1_112/O 0.15fF
C13883 POR2X1_814/B POR2X1_337/Y 0.08fF
C13884 PAND2X1_23/Y POR2X1_180/A 0.03fF
C13885 POR2X1_38/Y POR2X1_522/Y 0.02fF
C13886 PAND2X1_6/A PAND2X1_60/B 0.03fF
C13887 POR2X1_845/A POR2X1_5/Y 0.06fF
C13888 PAND2X1_652/O PAND2X1_557/A 0.02fF
C13889 PAND2X1_860/A POR2X1_679/A 0.01fF
C13890 PAND2X1_6/Y POR2X1_228/Y 0.04fF
C13891 POR2X1_359/B VDD 0.26fF
C13892 POR2X1_72/B PAND2X1_326/B 0.03fF
C13893 POR2X1_271/A POR2X1_256/O 0.01fF
C13894 PAND2X1_90/Y POR2X1_383/O 0.02fF
C13895 POR2X1_814/A PAND2X1_417/CTRL2 0.03fF
C13896 POR2X1_271/A PAND2X1_515/CTRL 0.05fF
C13897 POR2X1_407/A POR2X1_855/B 0.03fF
C13898 POR2X1_102/Y POR2X1_77/Y 1.59fF
C13899 POR2X1_43/B PAND2X1_510/B 0.03fF
C13900 POR2X1_327/Y POR2X1_302/a_16_28# 0.03fF
C13901 POR2X1_164/Y POR2X1_693/Y 0.26fF
C13902 POR2X1_341/Y POR2X1_350/B 0.01fF
C13903 PAND2X1_8/Y POR2X1_620/B 0.07fF
C13904 PAND2X1_739/Y PAND2X1_730/A 0.02fF
C13905 POR2X1_548/A POR2X1_68/B 0.10fF
C13906 POR2X1_465/B POR2X1_553/CTRL2 0.00fF
C13907 INPUT_0 POR2X1_371/O 0.02fF
C13908 POR2X1_510/Y POR2X1_573/A 0.09fF
C13909 POR2X1_316/Y PAND2X1_456/O 0.01fF
C13910 PAND2X1_140/A PAND2X1_113/a_16_344# 0.01fF
C13911 PAND2X1_436/A POR2X1_77/Y 0.07fF
C13912 POR2X1_593/CTRL2 POR2X1_832/B 0.01fF
C13913 POR2X1_559/B POR2X1_38/B 0.04fF
C13914 POR2X1_750/B POR2X1_736/A 0.05fF
C13915 PAND2X1_200/B POR2X1_42/Y 0.01fF
C13916 POR2X1_334/Y POR2X1_205/Y 0.07fF
C13917 PAND2X1_569/B POR2X1_73/Y 0.98fF
C13918 POR2X1_334/Y PAND2X1_55/Y 0.07fF
C13919 POR2X1_132/O POR2X1_7/B 0.01fF
C13920 PAND2X1_176/CTRL2 POR2X1_337/Y 0.01fF
C13921 POR2X1_814/A POR2X1_452/Y 0.22fF
C13922 POR2X1_567/A POR2X1_192/Y 0.08fF
C13923 POR2X1_753/Y POR2X1_90/O 0.02fF
C13924 POR2X1_147/a_16_28# PAND2X1_58/A 0.01fF
C13925 PAND2X1_797/Y VDD 0.26fF
C13926 PAND2X1_69/A POR2X1_456/B 0.03fF
C13927 PAND2X1_232/O POR2X1_68/B 0.04fF
C13928 D_GATE_222 POR2X1_186/B 0.08fF
C13929 PAND2X1_82/Y PAND2X1_397/CTRL2 0.03fF
C13930 POR2X1_119/Y POR2X1_7/B 0.03fF
C13931 POR2X1_16/A PAND2X1_341/A 0.00fF
C13932 POR2X1_81/A PAND2X1_735/O 0.01fF
C13933 PAND2X1_853/O PAND2X1_853/B 0.02fF
C13934 POR2X1_528/Y POR2X1_7/A 0.00fF
C13935 D_INPUT_2 POR2X1_5/CTRL 0.01fF
C13936 POR2X1_101/Y PAND2X1_60/B 0.10fF
C13937 PAND2X1_41/B PAND2X1_52/B 23.81fF
C13938 POR2X1_383/A PAND2X1_63/B 0.11fF
C13939 POR2X1_514/CTRL2 PAND2X1_48/A 0.03fF
C13940 PAND2X1_562/a_76_28# POR2X1_394/A 0.02fF
C13941 POR2X1_416/B POR2X1_760/CTRL2 0.01fF
C13942 PAND2X1_41/B POR2X1_212/B 0.03fF
C13943 PAND2X1_824/B POR2X1_206/CTRL2 0.05fF
C13944 POR2X1_16/A POR2X1_91/Y 0.01fF
C13945 PAND2X1_23/Y POR2X1_508/B 0.03fF
C13946 POR2X1_55/Y PAND2X1_353/Y 0.15fF
C13947 PAND2X1_724/B PAND2X1_352/Y 0.06fF
C13948 PAND2X1_714/CTRL PAND2X1_326/B 0.01fF
C13949 POR2X1_41/B POR2X1_761/A 0.03fF
C13950 POR2X1_564/Y POR2X1_568/B 1.97fF
C13951 POR2X1_239/a_56_344# POR2X1_153/Y 0.00fF
C13952 PAND2X1_96/B POR2X1_774/A 0.03fF
C13953 PAND2X1_271/CTRL2 POR2X1_556/A 0.01fF
C13954 PAND2X1_6/Y PAND2X1_482/a_16_344# 0.01fF
C13955 POR2X1_447/B POR2X1_68/A 0.10fF
C13956 PAND2X1_48/A POR2X1_576/Y 0.03fF
C13957 POR2X1_702/CTRL2 POR2X1_186/B 0.01fF
C13958 PAND2X1_213/Y PAND2X1_704/a_16_344# 0.02fF
C13959 POR2X1_217/CTRL PAND2X1_72/A 0.04fF
C13960 POR2X1_857/B POR2X1_568/B 0.05fF
C13961 PAND2X1_563/A PAND2X1_854/A 0.02fF
C13962 POR2X1_814/A POR2X1_220/B 0.64fF
C13963 POR2X1_379/Y POR2X1_532/A 0.04fF
C13964 POR2X1_119/Y PAND2X1_477/B 0.00fF
C13965 POR2X1_486/B POR2X1_294/B 0.09fF
C13966 POR2X1_537/Y POR2X1_840/B 0.05fF
C13967 POR2X1_334/O POR2X1_101/Y 0.02fF
C13968 POR2X1_441/CTRL POR2X1_669/B 0.04fF
C13969 POR2X1_108/Y PAND2X1_348/A 0.01fF
C13970 POR2X1_257/A POR2X1_695/O 0.07fF
C13971 POR2X1_307/A PAND2X1_48/A 0.03fF
C13972 POR2X1_466/a_16_28# POR2X1_436/B 0.08fF
C13973 POR2X1_119/Y PAND2X1_711/O 0.06fF
C13974 POR2X1_16/A POR2X1_134/a_16_28# 0.03fF
C13975 PAND2X1_385/CTRL POR2X1_711/Y -0.03fF
C13976 POR2X1_57/A PAND2X1_352/CTRL2 0.03fF
C13977 POR2X1_520/CTRL POR2X1_559/A 0.04fF
C13978 POR2X1_23/Y POR2X1_441/Y 0.03fF
C13979 POR2X1_722/O PAND2X1_60/B 0.01fF
C13980 PAND2X1_63/B PAND2X1_71/Y 0.00fF
C13981 PAND2X1_808/Y POR2X1_77/Y 0.03fF
C13982 POR2X1_394/A PAND2X1_124/O 0.04fF
C13983 PAND2X1_23/Y POR2X1_325/B 0.02fF
C13984 POR2X1_316/Y POR2X1_73/Y 0.06fF
C13985 PAND2X1_696/CTRL2 PAND2X1_60/B 0.01fF
C13986 PAND2X1_94/A PAND2X1_48/A 0.05fF
C13987 POR2X1_102/Y PAND2X1_449/O 0.03fF
C13988 POR2X1_118/CTRL POR2X1_77/Y 0.01fF
C13989 POR2X1_567/B POR2X1_446/B 0.05fF
C13990 POR2X1_431/CTRL PAND2X1_390/Y 0.01fF
C13991 PAND2X1_317/Y POR2X1_167/Y 0.01fF
C13992 POR2X1_796/A POR2X1_722/a_16_28# 0.02fF
C13993 POR2X1_4/Y PAND2X1_528/CTRL 0.05fF
C13994 POR2X1_687/O POR2X1_452/Y 0.01fF
C13995 POR2X1_394/A POR2X1_129/Y 0.05fF
C13996 POR2X1_614/A PAND2X1_681/CTRL 0.01fF
C13997 PAND2X1_435/CTRL POR2X1_677/Y 0.00fF
C13998 PAND2X1_438/CTRL VDD 0.00fF
C13999 POR2X1_821/Y POR2X1_77/Y 0.12fF
C14000 POR2X1_83/B PAND2X1_201/a_76_28# 0.00fF
C14001 POR2X1_16/A POR2X1_397/O 0.01fF
C14002 POR2X1_416/B PAND2X1_324/a_76_28# 0.01fF
C14003 POR2X1_632/Y POR2X1_228/Y 0.07fF
C14004 POR2X1_853/A POR2X1_863/A 0.03fF
C14005 PAND2X1_35/A POR2X1_29/A 0.02fF
C14006 POR2X1_866/A POR2X1_807/a_76_344# 0.01fF
C14007 POR2X1_477/B POR2X1_477/CTRL 0.00fF
C14008 POR2X1_857/A POR2X1_857/a_16_28# 0.03fF
C14009 POR2X1_849/B POR2X1_849/A 0.04fF
C14010 POR2X1_283/A POR2X1_39/B 1.48fF
C14011 POR2X1_49/Y PAND2X1_466/A 0.05fF
C14012 PAND2X1_659/Y POR2X1_394/A 0.10fF
C14013 POR2X1_41/B POR2X1_9/Y 0.01fF
C14014 POR2X1_146/a_16_28# PAND2X1_797/Y 0.02fF
C14015 PAND2X1_177/a_16_344# PAND2X1_52/B 0.01fF
C14016 POR2X1_49/Y POR2X1_262/Y 0.03fF
C14017 PAND2X1_116/CTRL2 POR2X1_150/Y 0.01fF
C14018 POR2X1_169/a_16_28# POR2X1_192/B 0.02fF
C14019 POR2X1_77/O POR2X1_14/Y 0.01fF
C14020 PAND2X1_366/a_56_28# PAND2X1_354/Y 0.00fF
C14021 POR2X1_116/A POR2X1_860/A 0.15fF
C14022 POR2X1_846/O PAND2X1_6/A 0.08fF
C14023 POR2X1_257/A POR2X1_495/CTRL 0.03fF
C14024 POR2X1_278/Y PAND2X1_717/A 0.07fF
C14025 PAND2X1_224/O POR2X1_578/Y 0.01fF
C14026 PAND2X1_23/Y PAND2X1_94/Y 0.02fF
C14027 PAND2X1_803/CTRL PAND2X1_797/Y 0.01fF
C14028 POR2X1_411/B PAND2X1_340/CTRL2 0.09fF
C14029 POR2X1_113/Y POR2X1_717/B 0.05fF
C14030 POR2X1_800/a_16_28# POR2X1_452/Y 0.03fF
C14031 POR2X1_550/A PAND2X1_52/B 0.00fF
C14032 PAND2X1_95/B D_INPUT_7 0.04fF
C14033 PAND2X1_245/CTRL POR2X1_66/A 0.05fF
C14034 PAND2X1_446/Y PAND2X1_803/A 0.02fF
C14035 PAND2X1_48/A PAND2X1_136/CTRL2 0.03fF
C14036 POR2X1_486/CTRL2 POR2X1_294/B 0.03fF
C14037 POR2X1_848/Y POR2X1_734/A 0.03fF
C14038 POR2X1_49/Y PAND2X1_477/CTRL2 0.01fF
C14039 POR2X1_153/Y PAND2X1_841/Y 0.01fF
C14040 POR2X1_796/Y POR2X1_808/A 0.00fF
C14041 POR2X1_329/a_16_28# POR2X1_329/A 0.03fF
C14042 POR2X1_83/Y PAND2X1_476/A 0.02fF
C14043 PAND2X1_217/B PAND2X1_267/Y 0.14fF
C14044 PAND2X1_299/CTRL POR2X1_260/B 0.01fF
C14045 POR2X1_654/B POR2X1_862/A 0.03fF
C14046 PAND2X1_214/CTRL2 POR2X1_40/Y 0.03fF
C14047 POR2X1_646/B POR2X1_294/B 0.05fF
C14048 POR2X1_180/B POR2X1_181/A 0.02fF
C14049 POR2X1_270/Y POR2X1_750/B 0.05fF
C14050 POR2X1_257/A POR2X1_257/a_16_28# 0.03fF
C14051 INPUT_3 PAND2X1_8/Y 0.09fF
C14052 POR2X1_717/B POR2X1_260/A 0.03fF
C14053 PAND2X1_200/Y POR2X1_32/A 0.01fF
C14054 POR2X1_476/A POR2X1_476/O 0.06fF
C14055 POR2X1_394/A PAND2X1_333/Y 0.07fF
C14056 POR2X1_78/B POR2X1_446/B 0.06fF
C14057 POR2X1_212/A VDD 0.36fF
C14058 POR2X1_141/Y POR2X1_218/Y 0.05fF
C14059 POR2X1_78/B POR2X1_240/O 0.09fF
C14060 POR2X1_632/m4_208_n4# POR2X1_750/B 0.07fF
C14061 POR2X1_814/B POR2X1_558/B 0.06fF
C14062 PAND2X1_206/B PAND2X1_6/A 0.16fF
C14063 POR2X1_54/Y PAND2X1_459/Y 0.18fF
C14064 PAND2X1_39/B POR2X1_646/CTRL2 0.00fF
C14065 PAND2X1_255/CTRL PAND2X1_60/B 0.01fF
C14066 POR2X1_483/A PAND2X1_93/B 0.03fF
C14067 POR2X1_667/O POR2X1_73/Y 0.02fF
C14068 POR2X1_334/B POR2X1_556/A 0.05fF
C14069 POR2X1_856/B PAND2X1_90/Y 0.06fF
C14070 POR2X1_83/B PAND2X1_214/A 0.03fF
C14071 PAND2X1_267/Y VDD 0.38fF
C14072 POR2X1_654/B PAND2X1_73/Y 0.27fF
C14073 POR2X1_220/O POR2X1_220/Y 0.00fF
C14074 POR2X1_343/Y POR2X1_4/Y 0.14fF
C14075 POR2X1_65/A POR2X1_423/CTRL2 0.01fF
C14076 PAND2X1_404/Y POR2X1_46/Y 0.03fF
C14077 POR2X1_734/B VDD 0.11fF
C14078 POR2X1_855/a_16_28# POR2X1_855/A 0.09fF
C14079 POR2X1_659/A POR2X1_554/Y 0.36fF
C14080 PAND2X1_817/O POR2X1_750/B 0.07fF
C14081 POR2X1_287/B POR2X1_78/A 0.03fF
C14082 POR2X1_271/B POR2X1_56/Y 0.03fF
C14083 PAND2X1_408/O PAND2X1_32/B 0.03fF
C14084 POR2X1_117/CTRL2 POR2X1_60/A 0.03fF
C14085 POR2X1_640/CTRL2 PAND2X1_41/B 0.11fF
C14086 POR2X1_188/A POR2X1_830/O 0.01fF
C14087 POR2X1_66/B POR2X1_734/A 0.07fF
C14088 POR2X1_669/B POR2X1_511/Y 0.07fF
C14089 POR2X1_541/B POR2X1_786/Y 0.09fF
C14090 POR2X1_20/B POR2X1_816/A 0.05fF
C14091 POR2X1_124/B POR2X1_556/A 0.00fF
C14092 POR2X1_49/Y PAND2X1_623/m4_208_n4# 0.12fF
C14093 POR2X1_298/a_16_28# POR2X1_46/Y 0.02fF
C14094 POR2X1_52/A POR2X1_848/A 0.07fF
C14095 POR2X1_20/B D_INPUT_1 0.73fF
C14096 POR2X1_52/A PAND2X1_776/Y 0.01fF
C14097 POR2X1_65/Y PAND2X1_6/A 0.02fF
C14098 POR2X1_142/a_16_28# POR2X1_65/A 0.03fF
C14099 POR2X1_42/O POR2X1_411/B 0.02fF
C14100 POR2X1_43/B PAND2X1_211/O 0.04fF
C14101 PAND2X1_865/Y PAND2X1_332/Y 0.03fF
C14102 D_INPUT_0 POR2X1_722/Y 0.03fF
C14103 POR2X1_56/CTRL2 POR2X1_516/B 0.00fF
C14104 POR2X1_555/B VDD 0.53fF
C14105 POR2X1_327/O POR2X1_558/B 0.00fF
C14106 POR2X1_78/B POR2X1_121/B 0.03fF
C14107 POR2X1_49/Y PAND2X1_849/CTRL2 0.00fF
C14108 POR2X1_376/B POR2X1_27/Y 0.01fF
C14109 POR2X1_769/B PAND2X1_52/B 0.03fF
C14110 POR2X1_499/A POR2X1_137/Y 0.03fF
C14111 POR2X1_78/A PAND2X1_8/Y 0.04fF
C14112 POR2X1_150/Y POR2X1_142/Y 0.03fF
C14113 PAND2X1_462/CTRL POR2X1_416/B 0.01fF
C14114 POR2X1_78/A POR2X1_724/CTRL 0.04fF
C14115 POR2X1_65/A POR2X1_176/m4_208_n4# 0.07fF
C14116 POR2X1_218/Y POR2X1_404/Y 0.07fF
C14117 PAND2X1_57/B POR2X1_247/Y 0.03fF
C14118 PAND2X1_6/Y POR2X1_454/A 0.02fF
C14119 POR2X1_78/B POR2X1_630/A 0.03fF
C14120 POR2X1_48/A PAND2X1_705/CTRL2 0.01fF
C14121 PAND2X1_20/A PAND2X1_516/CTRL2 0.01fF
C14122 POR2X1_64/CTRL POR2X1_39/B 0.01fF
C14123 POR2X1_150/Y PAND2X1_175/B 0.02fF
C14124 PAND2X1_5/a_16_344# INPUT_3 0.03fF
C14125 POR2X1_646/CTRL2 POR2X1_805/Y 0.03fF
C14126 POR2X1_186/Y PAND2X1_321/CTRL 0.12fF
C14127 POR2X1_181/O POR2X1_181/A 0.01fF
C14128 POR2X1_567/B POR2X1_795/B 0.05fF
C14129 POR2X1_49/Y PAND2X1_828/CTRL 0.04fF
C14130 POR2X1_416/B POR2X1_43/m4_208_n4# 0.07fF
C14131 POR2X1_653/CTRL2 POR2X1_750/B 0.12fF
C14132 POR2X1_78/A PAND2X1_89/CTRL 0.01fF
C14133 PAND2X1_263/a_56_28# POR2X1_94/A 0.00fF
C14134 PAND2X1_718/Y INPUT_0 0.16fF
C14135 PAND2X1_94/A PAND2X1_699/O 0.15fF
C14136 POR2X1_20/B PAND2X1_854/A 0.02fF
C14137 POR2X1_270/CTRL POR2X1_446/B 0.01fF
C14138 POR2X1_482/Y INPUT_0 0.16fF
C14139 PAND2X1_853/O POR2X1_23/Y 0.03fF
C14140 POR2X1_330/Y VDD 5.77fF
C14141 POR2X1_829/A PAND2X1_200/CTRL2 0.00fF
C14142 PAND2X1_624/A POR2X1_29/A 0.12fF
C14143 POR2X1_60/A POR2X1_252/CTRL2 0.01fF
C14144 POR2X1_852/O POR2X1_852/B 0.08fF
C14145 PAND2X1_118/O POR2X1_66/A 0.01fF
C14146 POR2X1_175/A VDD -0.00fF
C14147 POR2X1_556/A POR2X1_218/O 0.01fF
C14148 PAND2X1_740/Y POR2X1_331/Y 0.00fF
C14149 POR2X1_523/Y POR2X1_849/A 0.02fF
C14150 PAND2X1_732/O POR2X1_763/Y 0.09fF
C14151 PAND2X1_808/B VDD 0.11fF
C14152 POR2X1_614/A POR2X1_678/Y 0.00fF
C14153 POR2X1_260/B POR2X1_140/CTRL 0.01fF
C14154 POR2X1_66/A POR2X1_790/A 0.03fF
C14155 POR2X1_23/CTRL POR2X1_42/Y 0.01fF
C14156 D_INPUT_0 POR2X1_565/O 0.01fF
C14157 POR2X1_115/CTRL POR2X1_141/Y 0.01fF
C14158 PAND2X1_637/O PAND2X1_69/A 0.17fF
C14159 POR2X1_596/A POR2X1_866/A 0.05fF
C14160 POR2X1_262/CTRL2 POR2X1_40/Y 0.03fF
C14161 POR2X1_329/A POR2X1_594/CTRL2 0.01fF
C14162 POR2X1_788/A POR2X1_294/B 0.08fF
C14163 POR2X1_519/CTRL2 PAND2X1_838/B 0.01fF
C14164 POR2X1_814/B POR2X1_723/CTRL2 0.02fF
C14165 POR2X1_105/CTRL2 POR2X1_717/Y 0.01fF
C14166 POR2X1_734/B PAND2X1_32/B 0.01fF
C14167 POR2X1_555/B POR2X1_741/Y 0.03fF
C14168 PAND2X1_83/O POR2X1_66/A -0.00fF
C14169 POR2X1_859/A POR2X1_734/A 0.66fF
C14170 PAND2X1_56/O POR2X1_593/B 0.02fF
C14171 POR2X1_708/CTRL2 PAND2X1_65/B 0.01fF
C14172 PAND2X1_834/O PAND2X1_242/Y 0.05fF
C14173 POR2X1_428/Y PAND2X1_710/CTRL 0.01fF
C14174 POR2X1_849/A PAND2X1_69/A 0.00fF
C14175 POR2X1_833/A POR2X1_499/A 0.02fF
C14176 POR2X1_267/B INPUT_0 0.04fF
C14177 POR2X1_185/O PAND2X1_73/Y 0.04fF
C14178 POR2X1_13/A PAND2X1_474/A 5.10fF
C14179 POR2X1_669/B POR2X1_745/a_16_28# 0.04fF
C14180 POR2X1_614/A POR2X1_29/A 0.05fF
C14181 PAND2X1_20/A PAND2X1_79/O 0.06fF
C14182 POR2X1_65/A PAND2X1_863/B 0.03fF
C14183 POR2X1_119/Y PAND2X1_608/CTRL2 0.03fF
C14184 PAND2X1_96/CTRL2 PAND2X1_55/Y 0.01fF
C14185 POR2X1_66/A PAND2X1_88/Y 0.09fF
C14186 PAND2X1_20/A POR2X1_401/A 0.01fF
C14187 POR2X1_695/CTRL2 POR2X1_23/Y 0.01fF
C14188 POR2X1_33/CTRL D_INPUT_1 0.02fF
C14189 POR2X1_66/A POR2X1_84/Y 0.08fF
C14190 PAND2X1_431/O PAND2X1_60/B 0.06fF
C14191 POR2X1_32/A POR2X1_90/Y 0.19fF
C14192 POR2X1_311/Y PAND2X1_357/Y 38.07fF
C14193 PAND2X1_58/A POR2X1_459/B 0.02fF
C14194 POR2X1_102/Y POR2X1_52/Y 0.04fF
C14195 INPUT_2 PAND2X1_37/O 0.00fF
C14196 POR2X1_38/B POR2X1_29/A 0.15fF
C14197 POR2X1_72/B PAND2X1_575/A 0.03fF
C14198 POR2X1_355/A POR2X1_740/Y 0.03fF
C14199 POR2X1_411/B PAND2X1_853/B 0.06fF
C14200 PAND2X1_13/CTRL POR2X1_294/B 0.01fF
C14201 PAND2X1_95/B PAND2X1_41/B 0.73fF
C14202 POR2X1_383/A POR2X1_567/B 0.03fF
C14203 PAND2X1_430/CTRL2 INPUT_5 0.03fF
C14204 POR2X1_236/Y POR2X1_531/CTRL2 0.00fF
C14205 POR2X1_635/B PAND2X1_52/B 0.03fF
C14206 PAND2X1_9/CTRL PAND2X1_69/A 0.01fF
C14207 POR2X1_48/A POR2X1_283/A 4.10fF
C14208 POR2X1_855/B POR2X1_808/B 0.01fF
C14209 POR2X1_687/A POR2X1_796/Y 0.16fF
C14210 POR2X1_566/A POR2X1_471/CTRL2 0.15fF
C14211 POR2X1_285/Y POR2X1_649/CTRL 0.01fF
C14212 POR2X1_20/B PAND2X1_357/CTRL 0.01fF
C14213 POR2X1_829/Y POR2X1_7/B 0.03fF
C14214 POR2X1_68/A POR2X1_141/Y 0.05fF
C14215 PAND2X1_465/B POR2X1_5/Y 0.03fF
C14216 POR2X1_78/A POR2X1_209/A 0.06fF
C14217 POR2X1_409/B PAND2X1_196/CTRL2 0.01fF
C14218 POR2X1_9/Y POR2X1_77/Y 0.47fF
C14219 POR2X1_284/CTRL POR2X1_325/A 0.01fF
C14220 POR2X1_83/B POR2X1_591/Y 0.03fF
C14221 PAND2X1_6/A POR2X1_750/B 0.06fF
C14222 PAND2X1_84/CTRL POR2X1_293/Y 0.03fF
C14223 POR2X1_226/O POR2X1_382/Y 0.12fF
C14224 POR2X1_843/O PAND2X1_60/B 0.18fF
C14225 POR2X1_419/Y POR2X1_90/Y 0.00fF
C14226 POR2X1_417/Y POR2X1_90/Y 0.07fF
C14227 POR2X1_283/A POR2X1_225/CTRL2 0.01fF
C14228 POR2X1_777/B POR2X1_778/B 0.03fF
C14229 POR2X1_41/B POR2X1_368/O 0.02fF
C14230 PAND2X1_241/Y POR2X1_102/Y 0.01fF
C14231 POR2X1_330/Y PAND2X1_32/B 0.08fF
C14232 POR2X1_343/Y POR2X1_458/Y 0.03fF
C14233 POR2X1_461/O POR2X1_793/A 0.01fF
C14234 POR2X1_41/B POR2X1_278/Y 0.12fF
C14235 PAND2X1_485/CTRL POR2X1_260/A 0.01fF
C14236 POR2X1_403/O POR2X1_35/Y 0.01fF
C14237 POR2X1_65/A PAND2X1_566/Y 0.07fF
C14238 POR2X1_47/CTRL2 VDD -0.00fF
C14239 POR2X1_175/A PAND2X1_32/B 0.03fF
C14240 PAND2X1_96/B POR2X1_202/CTRL 0.01fF
C14241 POR2X1_51/A POR2X1_64/O 0.01fF
C14242 POR2X1_120/O POR2X1_294/B 0.01fF
C14243 POR2X1_311/Y PAND2X1_140/A 0.03fF
C14244 POR2X1_660/O POR2X1_725/Y 0.05fF
C14245 PAND2X1_39/B POR2X1_342/O 0.07fF
C14246 POR2X1_52/A PAND2X1_137/Y 0.07fF
C14247 PAND2X1_472/A PAND2X1_721/O 0.10fF
C14248 PAND2X1_20/A POR2X1_574/A 0.01fF
C14249 POR2X1_41/B POR2X1_829/A 0.12fF
C14250 POR2X1_48/A PAND2X1_713/CTRL2 0.01fF
C14251 POR2X1_260/B POR2X1_557/B 0.03fF
C14252 POR2X1_78/B POR2X1_795/B 0.10fF
C14253 POR2X1_785/CTRL2 POR2X1_785/A 0.00fF
C14254 PAND2X1_406/CTRL2 PAND2X1_48/A 0.03fF
C14255 POR2X1_61/Y POR2X1_219/O 0.03fF
C14256 PAND2X1_65/B POR2X1_778/B 0.07fF
C14257 POR2X1_89/a_16_28# POR2X1_394/A 0.06fF
C14258 POR2X1_757/A VDD 0.00fF
C14259 PAND2X1_118/CTRL INPUT_0 0.01fF
C14260 POR2X1_51/B POR2X1_83/B 0.02fF
C14261 POR2X1_669/B PAND2X1_124/O 0.02fF
C14262 POR2X1_22/A VDD 0.59fF
C14263 POR2X1_448/B PAND2X1_69/A 0.01fF
C14264 POR2X1_519/Y VDD 0.16fF
C14265 PAND2X1_65/B PAND2X1_518/CTRL 0.01fF
C14266 D_INPUT_0 POR2X1_244/Y 0.03fF
C14267 PAND2X1_585/a_76_28# PAND2X1_60/B 0.01fF
C14268 PAND2X1_695/CTRL2 POR2X1_407/Y 0.01fF
C14269 POR2X1_322/Y POR2X1_72/B 0.40fF
C14270 PAND2X1_221/a_16_344# POR2X1_283/A 0.01fF
C14271 POR2X1_197/CTRL PAND2X1_6/Y 0.01fF
C14272 POR2X1_37/Y POR2X1_394/A 0.78fF
C14273 POR2X1_263/Y PAND2X1_560/B 0.03fF
C14274 POR2X1_65/A PAND2X1_640/a_76_28# 0.01fF
C14275 POR2X1_43/B POR2X1_821/O 0.02fF
C14276 PAND2X1_58/A POR2X1_750/Y 0.02fF
C14277 POR2X1_302/CTRL PAND2X1_32/B 0.01fF
C14278 POR2X1_194/A POR2X1_194/m4_208_n4# 0.01fF
C14279 POR2X1_253/Y VDD 0.18fF
C14280 POR2X1_119/Y POR2X1_265/CTRL2 0.13fF
C14281 POR2X1_789/A POR2X1_546/A 0.07fF
C14282 POR2X1_13/A POR2X1_683/Y 0.12fF
C14283 POR2X1_588/Y POR2X1_750/B 0.03fF
C14284 POR2X1_68/A POR2X1_220/Y 0.21fF
C14285 POR2X1_83/A PAND2X1_35/Y 0.00fF
C14286 POR2X1_29/Y VDD 0.18fF
C14287 POR2X1_189/Y PAND2X1_191/Y 0.00fF
C14288 PAND2X1_769/a_16_344# POR2X1_73/Y 0.02fF
C14289 POR2X1_634/A POR2X1_774/B 0.04fF
C14290 POR2X1_84/CTRL POR2X1_294/B 0.01fF
C14291 POR2X1_334/B POR2X1_137/O 0.05fF
C14292 POR2X1_186/Y POR2X1_725/Y 0.20fF
C14293 POR2X1_526/O PAND2X1_556/B 0.08fF
C14294 POR2X1_383/A PAND2X1_386/CTRL 0.10fF
C14295 POR2X1_669/B POR2X1_129/Y 0.05fF
C14296 PAND2X1_104/CTRL INPUT_1 0.01fF
C14297 POR2X1_538/A POR2X1_814/B 0.04fF
C14298 POR2X1_608/Y POR2X1_774/A 0.00fF
C14299 PAND2X1_57/B PAND2X1_69/A 0.22fF
C14300 PAND2X1_6/Y POR2X1_832/a_16_28# 0.03fF
C14301 POR2X1_43/B PAND2X1_335/a_16_344# 0.01fF
C14302 PAND2X1_474/A PAND2X1_510/B 0.03fF
C14303 VDD POR2X1_148/A 0.00fF
C14304 POR2X1_45/Y POR2X1_42/Y 1.68fF
C14305 POR2X1_38/B POR2X1_546/A 0.07fF
C14306 POR2X1_273/CTRL2 POR2X1_39/B 0.03fF
C14307 PAND2X1_480/CTRL PAND2X1_478/B 0.01fF
C14308 POR2X1_861/O POR2X1_572/B 0.01fF
C14309 POR2X1_526/Y VDD 0.44fF
C14310 POR2X1_696/CTRL2 POR2X1_394/A 0.01fF
C14311 PAND2X1_65/B POR2X1_854/B 0.14fF
C14312 POR2X1_555/B POR2X1_228/CTRL 0.01fF
C14313 POR2X1_259/CTRL PAND2X1_52/Y 0.01fF
C14314 POR2X1_57/A PAND2X1_520/O 0.04fF
C14315 PAND2X1_65/B POR2X1_710/B 0.10fF
C14316 POR2X1_685/O POR2X1_729/Y 0.01fF
C14317 POR2X1_569/CTRL POR2X1_570/Y 0.03fF
C14318 PAND2X1_512/Y POR2X1_239/Y 0.01fF
C14319 POR2X1_140/B POR2X1_574/CTRL2 0.00fF
C14320 POR2X1_348/a_16_28# POR2X1_814/B 0.02fF
C14321 POR2X1_68/A PAND2X1_273/CTRL 0.01fF
C14322 POR2X1_814/B POR2X1_362/A 0.03fF
C14323 POR2X1_110/Y POR2X1_32/A 0.02fF
C14324 POR2X1_96/B POR2X1_236/Y 0.20fF
C14325 PAND2X1_659/Y POR2X1_669/B 0.03fF
C14326 POR2X1_78/B POR2X1_383/A 0.17fF
C14327 POR2X1_111/CTRL2 POR2X1_293/Y -0.02fF
C14328 PAND2X1_55/Y POR2X1_435/CTRL 0.00fF
C14329 PAND2X1_47/B PAND2X1_18/B 0.01fF
C14330 PAND2X1_90/Y POR2X1_151/CTRL2 0.31fF
C14331 PAND2X1_241/a_16_344# POR2X1_90/Y 0.01fF
C14332 PAND2X1_579/A PAND2X1_579/O -0.00fF
C14333 POR2X1_606/Y PAND2X1_48/A 0.11fF
C14334 POR2X1_121/B POR2X1_294/A 0.10fF
C14335 INPUT_0 PAND2X1_349/A 0.40fF
C14336 PAND2X1_48/B POR2X1_840/B 0.05fF
C14337 PAND2X1_850/Y D_INPUT_0 0.07fF
C14338 PAND2X1_41/B POR2X1_216/Y 0.01fF
C14339 PAND2X1_831/CTRL POR2X1_153/Y 0.01fF
C14340 PAND2X1_770/O POR2X1_765/Y 0.01fF
C14341 INPUT_0 PAND2X1_63/B 0.03fF
C14342 POR2X1_435/B PAND2X1_72/A 0.01fF
C14343 POR2X1_96/Y POR2X1_669/B 0.03fF
C14344 POR2X1_96/A POR2X1_245/Y 0.01fF
C14345 PAND2X1_687/B POR2X1_669/B 0.02fF
C14346 POR2X1_447/B PAND2X1_58/A 0.09fF
C14347 POR2X1_230/Y POR2X1_229/Y 0.14fF
C14348 PAND2X1_631/CTRL PAND2X1_6/A 0.03fF
C14349 POR2X1_68/A PAND2X1_29/a_16_344# 0.02fF
C14350 POR2X1_455/A POR2X1_702/A 0.00fF
C14351 POR2X1_586/Y POR2X1_585/CTRL2 0.01fF
C14352 PAND2X1_762/CTRL2 PAND2X1_52/B 0.03fF
C14353 POR2X1_198/CTRL PAND2X1_88/Y 0.01fF
C14354 PAND2X1_572/CTRL PAND2X1_197/Y 0.00fF
C14355 PAND2X1_71/O PAND2X1_111/B 0.02fF
C14356 PAND2X1_477/B POR2X1_237/Y 0.18fF
C14357 POR2X1_35/Y POR2X1_219/O 0.01fF
C14358 POR2X1_83/A PAND2X1_243/CTRL 0.01fF
C14359 POR2X1_343/Y PAND2X1_251/O 0.34fF
C14360 POR2X1_46/Y PAND2X1_123/CTRL2 0.03fF
C14361 POR2X1_366/Y POR2X1_704/CTRL2 0.02fF
C14362 POR2X1_252/O POR2X1_7/A 0.11fF
C14363 POR2X1_805/Y PAND2X1_759/CTRL 0.01fF
C14364 POR2X1_222/Y PAND2X1_88/Y 0.03fF
C14365 POR2X1_110/Y POR2X1_417/Y 0.55fF
C14366 POR2X1_322/Y POR2X1_323/Y 0.00fF
C14367 POR2X1_683/Y PAND2X1_643/Y 0.03fF
C14368 POR2X1_728/B POR2X1_687/A 0.01fF
C14369 POR2X1_396/Y POR2X1_42/Y 0.15fF
C14370 PAND2X1_254/CTRL2 POR2X1_7/A 0.05fF
C14371 PAND2X1_118/O POR2X1_532/A 0.15fF
C14372 PAND2X1_23/Y PAND2X1_60/B 0.56fF
C14373 POR2X1_130/A POR2X1_664/O 0.02fF
C14374 PAND2X1_90/A POR2X1_548/A 0.00fF
C14375 POR2X1_356/A PAND2X1_173/m4_208_n4# 0.03fF
C14376 PAND2X1_651/Y POR2X1_90/Y 0.03fF
C14377 POR2X1_828/A PAND2X1_69/A 3.95fF
C14378 PAND2X1_64/CTRL PAND2X1_52/B 0.01fF
C14379 POR2X1_614/A PAND2X1_150/CTRL 0.06fF
C14380 POR2X1_72/B POR2X1_373/O 0.01fF
C14381 POR2X1_57/CTRL2 PAND2X1_737/B 0.01fF
C14382 POR2X1_57/A PAND2X1_547/O 0.03fF
C14383 PAND2X1_737/O POR2X1_40/Y 0.02fF
C14384 POR2X1_752/CTRL INPUT_5 0.01fF
C14385 POR2X1_416/B POR2X1_699/a_16_28# 0.03fF
C14386 PAND2X1_824/B PAND2X1_57/B 0.03fF
C14387 VDD POR2X1_715/A 0.14fF
C14388 POR2X1_327/Y POR2X1_130/A 0.03fF
C14389 POR2X1_366/O PAND2X1_48/B 0.01fF
C14390 POR2X1_567/A POR2X1_456/O 0.01fF
C14391 POR2X1_96/A PAND2X1_507/CTRL 0.05fF
C14392 PAND2X1_724/B POR2X1_310/Y 0.64fF
C14393 POR2X1_14/Y POR2X1_39/B 28.69fF
C14394 POR2X1_78/B PAND2X1_71/Y 0.04fF
C14395 POR2X1_153/CTRL2 POR2X1_7/B 0.03fF
C14396 POR2X1_121/A POR2X1_725/Y 0.09fF
C14397 POR2X1_532/A PAND2X1_88/Y 0.03fF
C14398 POR2X1_546/B POR2X1_546/CTRL2 0.02fF
C14399 POR2X1_36/B POR2X1_36/CTRL2 0.02fF
C14400 POR2X1_532/A POR2X1_84/Y 0.04fF
C14401 PAND2X1_270/CTRL POR2X1_73/Y 0.01fF
C14402 PAND2X1_453/A POR2X1_39/B 0.03fF
C14403 POR2X1_327/Y POR2X1_566/A 0.03fF
C14404 POR2X1_399/CTRL2 POR2X1_119/Y 0.01fF
C14405 POR2X1_46/Y PAND2X1_514/a_76_28# 0.03fF
C14406 POR2X1_55/Y PAND2X1_514/O 0.17fF
C14407 PAND2X1_119/a_56_28# PAND2X1_96/B 0.00fF
C14408 POR2X1_662/Y POR2X1_675/Y 0.03fF
C14409 PAND2X1_545/Y PAND2X1_324/Y 0.00fF
C14410 VDD POR2X1_703/O 0.00fF
C14411 PAND2X1_786/m4_208_n4# POR2X1_150/m4_208_n4# 0.13fF
C14412 POR2X1_37/Y POR2X1_90/CTRL2 0.00fF
C14413 PAND2X1_23/Y POR2X1_353/A 0.03fF
C14414 POR2X1_68/A POR2X1_215/A 0.61fF
C14415 POR2X1_332/B POR2X1_332/Y 0.02fF
C14416 POR2X1_108/Y POR2X1_183/Y 0.00fF
C14417 PAND2X1_481/CTRL2 POR2X1_294/B 0.00fF
C14418 POR2X1_394/A POR2X1_293/Y 0.27fF
C14419 POR2X1_52/A PAND2X1_853/B 0.03fF
C14420 POR2X1_643/CTRL POR2X1_643/Y 0.05fF
C14421 PAND2X1_23/Y POR2X1_332/O 0.02fF
C14422 VDD POR2X1_337/Y 0.00fF
C14423 PAND2X1_215/B PAND2X1_560/B 0.03fF
C14424 PAND2X1_23/Y POR2X1_787/a_16_28# 0.03fF
C14425 POR2X1_169/B VDD 0.10fF
C14426 POR2X1_662/Y POR2X1_544/B 0.04fF
C14427 POR2X1_447/a_16_28# POR2X1_510/Y 0.02fF
C14428 POR2X1_68/A POR2X1_546/CTRL 0.01fF
C14429 POR2X1_224/Y POR2X1_394/A 0.04fF
C14430 PAND2X1_482/CTRL POR2X1_294/B 0.01fF
C14431 PAND2X1_56/Y PAND2X1_142/CTRL2 0.01fF
C14432 PAND2X1_551/CTRL2 PAND2X1_854/A 0.00fF
C14433 POR2X1_394/A PAND2X1_302/a_16_344# 0.01fF
C14434 POR2X1_596/A POR2X1_596/CTRL2 0.01fF
C14435 POR2X1_245/Y POR2X1_7/A 0.10fF
C14436 POR2X1_297/a_16_28# POR2X1_77/Y 0.02fF
C14437 POR2X1_614/A POR2X1_520/B 0.08fF
C14438 POR2X1_119/Y PAND2X1_839/CTRL2 0.01fF
C14439 POR2X1_750/B POR2X1_161/a_56_344# 0.01fF
C14440 PAND2X1_701/O PAND2X1_69/A 0.15fF
C14441 POR2X1_13/A PAND2X1_346/O 0.02fF
C14442 PAND2X1_234/O POR2X1_66/A 0.02fF
C14443 POR2X1_537/CTRL2 PAND2X1_60/B 0.01fF
C14444 POR2X1_715/A PAND2X1_32/B 0.01fF
C14445 PAND2X1_251/CTRL POR2X1_814/A 0.01fF
C14446 PAND2X1_797/Y PAND2X1_714/O 0.01fF
C14447 PAND2X1_93/B POR2X1_630/B 0.01fF
C14448 INPUT_3 POR2X1_20/B 0.20fF
C14449 POR2X1_360/A PAND2X1_290/CTRL2 0.05fF
C14450 POR2X1_16/A POR2X1_235/CTRL 0.10fF
C14451 POR2X1_57/A PAND2X1_182/B 0.03fF
C14452 POR2X1_463/Y POR2X1_713/B 0.03fF
C14453 POR2X1_556/Y POR2X1_339/Y 0.22fF
C14454 PAND2X1_658/A POR2X1_4/Y 0.03fF
C14455 POR2X1_78/CTRL2 POR2X1_571/Y 0.01fF
C14456 POR2X1_719/B PAND2X1_60/B 0.01fF
C14457 POR2X1_278/Y POR2X1_77/Y 0.03fF
C14458 POR2X1_278/A POR2X1_153/Y 0.09fF
C14459 POR2X1_116/A POR2X1_446/B 0.01fF
C14460 POR2X1_110/Y PAND2X1_651/Y 0.08fF
C14461 PAND2X1_69/A POR2X1_512/CTRL2 0.00fF
C14462 POR2X1_7/A PAND2X1_507/CTRL 0.01fF
C14463 PAND2X1_6/Y POR2X1_99/B 0.03fF
C14464 POR2X1_865/O PAND2X1_48/A 0.01fF
C14465 POR2X1_334/Y POR2X1_360/CTRL 0.01fF
C14466 PAND2X1_94/A POR2X1_789/B 0.01fF
C14467 POR2X1_416/B PAND2X1_793/Y 0.03fF
C14468 POR2X1_343/Y PAND2X1_71/CTRL 0.28fF
C14469 PAND2X1_651/O POR2X1_588/Y 0.02fF
C14470 POR2X1_447/B PAND2X1_96/B 0.12fF
C14471 POR2X1_55/Y POR2X1_39/B 0.94fF
C14472 PAND2X1_242/Y POR2X1_432/Y 0.05fF
C14473 POR2X1_809/A PAND2X1_60/B 0.02fF
C14474 PAND2X1_726/CTRL2 POR2X1_39/B 0.01fF
C14475 POR2X1_860/m4_208_n4# POR2X1_383/A 0.12fF
C14476 PAND2X1_48/B PAND2X1_56/A 0.01fF
C14477 PAND2X1_39/B PAND2X1_609/CTRL 0.01fF
C14478 POR2X1_463/O PAND2X1_58/A 0.16fF
C14479 POR2X1_722/A POR2X1_796/A 0.03fF
C14480 POR2X1_16/A PAND2X1_341/Y 0.00fF
C14481 PAND2X1_844/Y PAND2X1_333/Y 0.12fF
C14482 POR2X1_23/Y POR2X1_411/B 0.10fF
C14483 POR2X1_16/A POR2X1_599/CTRL2 0.14fF
C14484 POR2X1_119/Y POR2X1_824/Y 0.02fF
C14485 POR2X1_383/A POR2X1_294/A 0.06fF
C14486 POR2X1_175/B POR2X1_186/B 0.01fF
C14487 POR2X1_112/CTRL PAND2X1_60/B 0.01fF
C14488 POR2X1_327/Y POR2X1_539/O 0.15fF
C14489 POR2X1_189/O POR2X1_816/A 0.01fF
C14490 POR2X1_96/O POR2X1_153/Y 0.01fF
C14491 POR2X1_20/B POR2X1_432/CTRL2 0.01fF
C14492 POR2X1_494/Y PAND2X1_332/Y 0.03fF
C14493 POR2X1_260/B PAND2X1_406/CTRL 0.01fF
C14494 POR2X1_404/Y POR2X1_138/A 0.03fF
C14495 PAND2X1_440/O PAND2X1_794/B 0.02fF
C14496 POR2X1_532/A POR2X1_568/B 0.08fF
C14497 POR2X1_62/Y PAND2X1_100/O 0.02fF
C14498 POR2X1_178/O POR2X1_416/B 0.05fF
C14499 POR2X1_150/Y PAND2X1_794/CTRL 0.03fF
C14500 POR2X1_210/A POR2X1_210/B 0.04fF
C14501 POR2X1_557/B POR2X1_768/a_56_344# 0.00fF
C14502 POR2X1_97/O POR2X1_97/B 0.02fF
C14503 PAND2X1_353/O PAND2X1_353/Y 0.00fF
C14504 POR2X1_858/B POR2X1_851/m4_208_n4# 0.01fF
C14505 INPUT_2 PAND2X1_462/a_16_344# 0.03fF
C14506 POR2X1_77/Y PAND2X1_359/a_76_28# 0.01fF
C14507 POR2X1_54/Y POR2X1_753/Y 0.33fF
C14508 POR2X1_635/CTRL2 POR2X1_750/B 0.01fF
C14509 POR2X1_736/A POR2X1_318/A 0.03fF
C14510 PAND2X1_798/Y PAND2X1_366/A 0.08fF
C14511 POR2X1_866/A D_INPUT_0 0.03fF
C14512 POR2X1_153/Y POR2X1_117/Y 0.13fF
C14513 PAND2X1_60/B POR2X1_711/Y 0.10fF
C14514 D_INPUT_0 PAND2X1_28/a_16_344# 0.02fF
C14515 POR2X1_97/A POR2X1_212/a_76_344# 0.01fF
C14516 POR2X1_192/B POR2X1_545/a_16_28# 0.10fF
C14517 INPUT_2 POR2X1_8/O 0.01fF
C14518 PAND2X1_337/CTRL2 PAND2X1_336/Y 0.01fF
C14519 PAND2X1_609/CTRL POR2X1_805/Y 0.03fF
C14520 PAND2X1_71/Y POR2X1_294/A 0.03fF
C14521 POR2X1_614/CTRL POR2X1_614/Y 0.03fF
C14522 POR2X1_66/B PAND2X1_416/O 0.02fF
C14523 POR2X1_500/O POR2X1_318/A 0.01fF
C14524 POR2X1_862/Y POR2X1_121/B 0.00fF
C14525 POR2X1_49/Y POR2X1_442/O 0.03fF
C14526 POR2X1_34/CTRL POR2X1_34/Y 0.01fF
C14527 POR2X1_669/B POR2X1_37/Y 0.13fF
C14528 POR2X1_81/A POR2X1_129/Y 0.09fF
C14529 POR2X1_66/A PAND2X1_595/a_76_28# 0.01fF
C14530 POR2X1_48/A POR2X1_14/Y 0.10fF
C14531 POR2X1_274/O POR2X1_296/B 0.01fF
C14532 POR2X1_408/Y POR2X1_90/CTRL2 0.01fF
C14533 POR2X1_376/B PAND2X1_796/B 0.00fF
C14534 POR2X1_485/Y VDD 0.28fF
C14535 POR2X1_326/A POR2X1_532/CTRL 0.01fF
C14536 PAND2X1_282/O PAND2X1_73/Y 0.11fF
C14537 POR2X1_48/A PAND2X1_453/A 0.03fF
C14538 POR2X1_45/O POR2X1_411/B 0.02fF
C14539 POR2X1_376/B PAND2X1_454/B 0.02fF
C14540 PAND2X1_659/Y PAND2X1_649/A 0.03fF
C14541 PAND2X1_23/Y POR2X1_486/O 0.04fF
C14542 PAND2X1_124/Y POR2X1_72/B 0.03fF
C14543 POR2X1_590/A POR2X1_29/A 0.03fF
C14544 POR2X1_149/CTRL VDD -0.00fF
C14545 POR2X1_24/CTRL2 POR2X1_23/Y 0.01fF
C14546 POR2X1_98/O PAND2X1_20/A 0.02fF
C14547 PAND2X1_666/a_56_28# PAND2X1_20/A 0.00fF
C14548 POR2X1_630/a_16_28# POR2X1_630/A -0.00fF
C14549 PAND2X1_633/O PAND2X1_404/Y 0.00fF
C14550 POR2X1_696/CTRL2 POR2X1_669/B 0.03fF
C14551 PAND2X1_429/a_16_344# PAND2X1_11/Y 0.02fF
C14552 PAND2X1_341/B POR2X1_86/O 0.01fF
C14553 POR2X1_537/Y POR2X1_858/A 0.16fF
C14554 POR2X1_102/Y POR2X1_268/a_16_28# 0.01fF
C14555 POR2X1_68/A POR2X1_67/Y 0.03fF
C14556 POR2X1_647/O POR2X1_362/B 0.07fF
C14557 POR2X1_434/CTRL POR2X1_480/A 0.04fF
C14558 POR2X1_866/A PAND2X1_90/Y 0.10fF
C14559 POR2X1_848/A POR2X1_625/CTRL 0.05fF
C14560 POR2X1_859/a_16_28# PAND2X1_57/B 0.02fF
C14561 POR2X1_814/B POR2X1_499/CTRL 0.13fF
C14562 PAND2X1_591/O POR2X1_593/B 0.00fF
C14563 POR2X1_49/Y PAND2X1_68/CTRL 0.01fF
C14564 PAND2X1_631/A POR2X1_316/Y 0.03fF
C14565 POR2X1_814/A POR2X1_778/B 1.26fF
C14566 POR2X1_23/Y POR2X1_376/B 0.19fF
C14567 PAND2X1_416/O POR2X1_859/A 0.06fF
C14568 POR2X1_99/B POR2X1_632/Y 0.03fF
C14569 POR2X1_55/O POR2X1_94/A 0.02fF
C14570 POR2X1_102/Y PAND2X1_718/Y 0.50fF
C14571 PAND2X1_410/O PAND2X1_404/A 0.01fF
C14572 PAND2X1_48/B POR2X1_477/O 0.07fF
C14573 POR2X1_482/Y POR2X1_102/Y 0.03fF
C14574 PAND2X1_9/Y POR2X1_247/O 0.01fF
C14575 PAND2X1_285/CTRL2 VDD 0.00fF
C14576 POR2X1_52/A PAND2X1_796/B 0.02fF
C14577 PAND2X1_73/Y POR2X1_777/B 0.11fF
C14578 POR2X1_102/Y POR2X1_251/O 0.01fF
C14579 POR2X1_9/Y PAND2X1_350/a_16_344# 0.06fF
C14580 POR2X1_23/Y PAND2X1_712/O 0.03fF
C14581 PAND2X1_43/CTRL PAND2X1_55/Y 0.09fF
C14582 POR2X1_3/A POR2X1_18/CTRL2 0.02fF
C14583 PAND2X1_41/CTRL POR2X1_294/B 0.01fF
C14584 POR2X1_571/Y POR2X1_500/CTRL 0.01fF
C14585 POR2X1_218/Y POR2X1_217/CTRL2 0.09fF
C14586 POR2X1_189/Y POR2X1_679/a_16_28# 0.02fF
C14587 POR2X1_83/B POR2X1_72/B 0.20fF
C14588 POR2X1_86/Y PAND2X1_101/B 0.01fF
C14589 PAND2X1_63/Y PAND2X1_246/O 0.03fF
C14590 PAND2X1_675/A POR2X1_20/B 0.03fF
C14591 POR2X1_260/B POR2X1_76/Y 0.03fF
C14592 POR2X1_29/CTRL POR2X1_409/B 0.07fF
C14593 POR2X1_558/B VDD 0.15fF
C14594 PAND2X1_438/O POR2X1_180/A 0.07fF
C14595 PAND2X1_39/B POR2X1_572/B 0.11fF
C14596 PAND2X1_469/B POR2X1_20/B 0.05fF
C14597 POR2X1_471/A POR2X1_732/B 0.03fF
C14598 POR2X1_687/Y POR2X1_814/A 0.12fF
C14599 POR2X1_341/A POR2X1_222/Y 0.07fF
C14600 POR2X1_479/O POR2X1_286/Y 0.05fF
C14601 POR2X1_748/A POR2X1_40/Y 0.03fF
C14602 PAND2X1_206/B PAND2X1_350/CTRL 0.01fF
C14603 PAND2X1_65/B PAND2X1_73/Y 4.56fF
C14604 POR2X1_423/CTRL POR2X1_5/Y 0.01fF
C14605 PAND2X1_640/CTRL POR2X1_826/Y 0.01fF
C14606 POR2X1_20/a_16_28# POR2X1_20/A 0.05fF
C14607 POR2X1_693/Y POR2X1_257/A 0.73fF
C14608 POR2X1_366/Y POR2X1_76/A 0.03fF
C14609 POR2X1_808/A POR2X1_330/Y 0.10fF
C14610 PAND2X1_216/O PAND2X1_267/Y 0.02fF
C14611 POR2X1_663/CTRL POR2X1_78/A 0.01fF
C14612 POR2X1_102/Y POR2X1_106/Y 0.03fF
C14613 POR2X1_230/a_16_28# POR2X1_32/A 0.05fF
C14614 POR2X1_658/CTRL2 POR2X1_532/A 0.01fF
C14615 POR2X1_814/A POR2X1_854/B 0.10fF
C14616 PAND2X1_836/O POR2X1_411/B 0.04fF
C14617 PAND2X1_472/B POR2X1_48/A 0.07fF
C14618 POR2X1_864/CTRL POR2X1_774/Y 0.01fF
C14619 PAND2X1_585/a_16_344# PAND2X1_41/B 0.01fF
C14620 PAND2X1_217/B PAND2X1_795/CTRL 0.28fF
C14621 POR2X1_621/A PAND2X1_49/CTRL 0.00fF
C14622 POR2X1_847/O POR2X1_93/A 0.05fF
C14623 PAND2X1_413/O VDD 0.00fF
C14624 POR2X1_29/Y PAND2X1_9/Y 0.04fF
C14625 POR2X1_52/A POR2X1_23/Y 9.98fF
C14626 POR2X1_296/B POR2X1_547/B 0.95fF
C14627 POR2X1_265/a_16_28# PAND2X1_35/Y 0.02fF
C14628 POR2X1_96/A D_INPUT_0 0.08fF
C14629 POR2X1_614/A PAND2X1_39/B 0.17fF
C14630 POR2X1_260/B POR2X1_740/Y 0.01fF
C14631 POR2X1_32/A INPUT_0 10.22fF
C14632 POR2X1_83/B PAND2X1_520/CTRL2 0.03fF
C14633 PAND2X1_84/CTRL POR2X1_60/A 0.01fF
C14634 POR2X1_590/A POR2X1_546/A 0.03fF
C14635 POR2X1_43/B PAND2X1_444/CTRL 0.01fF
C14636 POR2X1_624/Y D_INPUT_1 0.10fF
C14637 POR2X1_48/A POR2X1_55/Y 2.50fF
C14638 POR2X1_389/a_76_344# POR2X1_260/B 0.01fF
C14639 POR2X1_186/Y POR2X1_776/CTRL 0.01fF
C14640 POR2X1_341/A POR2X1_532/A 0.07fF
C14641 POR2X1_623/O POR2X1_55/Y 0.03fF
C14642 PAND2X1_39/B POR2X1_38/B 0.05fF
C14643 POR2X1_48/A PAND2X1_726/CTRL2 0.03fF
C14644 POR2X1_23/Y PAND2X1_726/CTRL 0.00fF
C14645 POR2X1_16/A PAND2X1_717/A 0.03fF
C14646 POR2X1_848/A POR2X1_790/B 0.07fF
C14647 POR2X1_67/Y POR2X1_391/B 0.00fF
C14648 PAND2X1_58/A PAND2X1_511/O 0.02fF
C14649 POR2X1_68/A POR2X1_841/B 0.01fF
C14650 POR2X1_45/Y PAND2X1_576/B 0.03fF
C14651 PAND2X1_491/CTRL2 POR2X1_260/B 0.01fF
C14652 POR2X1_860/A POR2X1_475/A 0.01fF
C14653 POR2X1_590/A PAND2X1_754/O 0.03fF
C14654 POR2X1_502/A POR2X1_850/B 0.03fF
C14655 POR2X1_383/A POR2X1_116/A 0.03fF
C14656 POR2X1_457/O VDD 0.00fF
C14657 POR2X1_376/B PAND2X1_513/CTRL 0.08fF
C14658 PAND2X1_612/B PAND2X1_96/B 0.03fF
C14659 POR2X1_669/B POR2X1_293/Y 0.21fF
C14660 POR2X1_54/Y POR2X1_15/O 0.04fF
C14661 POR2X1_624/Y POR2X1_724/A 0.07fF
C14662 POR2X1_65/A POR2X1_107/CTRL2 0.03fF
C14663 POR2X1_856/B D_GATE_222 0.10fF
C14664 PAND2X1_48/B PAND2X1_594/O 0.01fF
C14665 POR2X1_241/B POR2X1_578/Y 0.03fF
C14666 PAND2X1_655/a_76_28# PAND2X1_655/B 0.02fF
C14667 POR2X1_32/A PAND2X1_717/CTRL2 0.03fF
C14668 POR2X1_319/A PAND2X1_314/CTRL2 0.00fF
C14669 POR2X1_590/A PAND2X1_110/CTRL 0.01fF
C14670 PAND2X1_66/CTRL2 POR2X1_38/Y 0.03fF
C14671 POR2X1_63/Y POR2X1_235/Y 0.01fF
C14672 POR2X1_383/A POR2X1_286/B 0.34fF
C14673 POR2X1_263/Y PAND2X1_734/CTRL2 0.01fF
C14674 PAND2X1_795/B POR2X1_72/B 0.03fF
C14675 PAND2X1_20/A POR2X1_193/A 0.03fF
C14676 PAND2X1_20/A POR2X1_579/Y 0.06fF
C14677 PAND2X1_793/Y POR2X1_487/Y 0.04fF
C14678 PAND2X1_601/CTRL PAND2X1_60/B 0.01fF
C14679 POR2X1_79/Y POR2X1_40/Y 0.03fF
C14680 POR2X1_558/B PAND2X1_32/B 0.03fF
C14681 POR2X1_257/A POR2X1_258/Y 0.03fF
C14682 POR2X1_41/B PAND2X1_169/Y 0.03fF
C14683 POR2X1_68/A PAND2X1_603/O 0.07fF
C14684 POR2X1_166/CTRL POR2X1_438/Y 0.09fF
C14685 POR2X1_264/Y POR2X1_78/A 0.04fF
C14686 POR2X1_865/B POR2X1_458/O 0.01fF
C14687 POR2X1_96/B POR2X1_24/Y 0.03fF
C14688 PAND2X1_862/Y POR2X1_329/A 0.09fF
C14689 PAND2X1_453/a_16_344# POR2X1_60/A 0.01fF
C14690 POR2X1_25/Y POR2X1_18/CTRL2 0.01fF
C14691 POR2X1_488/CTRL PAND2X1_738/Y 0.32fF
C14692 PAND2X1_557/A PAND2X1_592/Y 0.03fF
C14693 PAND2X1_401/CTRL POR2X1_14/Y 0.01fF
C14694 PAND2X1_39/B PAND2X1_393/a_76_28# 0.01fF
C14695 POR2X1_422/a_76_344# POR2X1_93/A 0.00fF
C14696 POR2X1_78/A POR2X1_562/m4_208_n4# 0.09fF
C14697 PAND2X1_721/O PAND2X1_673/Y 0.00fF
C14698 POR2X1_840/B POR2X1_656/CTRL 0.28fF
C14699 POR2X1_383/A POR2X1_862/Y 0.01fF
C14700 POR2X1_329/A POR2X1_385/Y 0.03fF
C14701 PAND2X1_266/CTRL2 POR2X1_7/Y 0.01fF
C14702 PAND2X1_366/Y VDD 0.30fF
C14703 POR2X1_287/B PAND2X1_371/CTRL2 0.01fF
C14704 PAND2X1_741/B INPUT_0 0.03fF
C14705 POR2X1_275/A POR2X1_394/A 0.04fF
C14706 PAND2X1_23/Y POR2X1_750/B 0.08fF
C14707 POR2X1_45/CTRL PAND2X1_480/B 0.14fF
C14708 POR2X1_78/B INPUT_0 0.03fF
C14709 PAND2X1_90/A PAND2X1_412/CTRL 0.02fF
C14710 POR2X1_723/CTRL2 VDD -0.00fF
C14711 POR2X1_54/Y POR2X1_754/O 0.02fF
C14712 PAND2X1_317/Y POR2X1_312/Y 0.07fF
C14713 POR2X1_814/B POR2X1_193/A 0.33fF
C14714 POR2X1_614/A PAND2X1_20/A 0.21fF
C14715 PAND2X1_73/Y POR2X1_541/CTRL 0.01fF
C14716 PAND2X1_346/a_76_28# POR2X1_295/Y 0.03fF
C14717 PAND2X1_52/Y POR2X1_785/A 0.03fF
C14718 POR2X1_390/B POR2X1_274/A 0.03fF
C14719 POR2X1_687/Y POR2X1_687/O 0.00fF
C14720 POR2X1_295/Y VDD 0.17fF
C14721 POR2X1_332/B VDD 0.00fF
C14722 POR2X1_814/B POR2X1_572/B 0.05fF
C14723 D_INPUT_0 POR2X1_7/A 0.16fF
C14724 POR2X1_52/A PAND2X1_558/O 0.17fF
C14725 POR2X1_559/B POR2X1_66/A 0.07fF
C14726 POR2X1_655/O POR2X1_711/Y 0.06fF
C14727 POR2X1_66/B POR2X1_556/Y 0.03fF
C14728 PAND2X1_20/A POR2X1_38/B 0.03fF
C14729 POR2X1_19/CTRL2 POR2X1_4/Y 0.06fF
C14730 POR2X1_741/Y POR2X1_543/A 0.03fF
C14731 POR2X1_257/A PAND2X1_725/CTRL 0.01fF
C14732 POR2X1_614/A POR2X1_254/CTRL 0.01fF
C14733 POR2X1_389/A POR2X1_121/B 0.23fF
C14734 POR2X1_220/Y POR2X1_435/Y 0.07fF
C14735 POR2X1_669/B POR2X1_408/Y 0.12fF
C14736 PAND2X1_280/a_76_28# PAND2X1_90/Y 0.06fF
C14737 POR2X1_65/A PAND2X1_105/CTRL 0.00fF
C14738 POR2X1_709/B POR2X1_709/A 0.31fF
C14739 POR2X1_860/A POR2X1_218/A 0.16fF
C14740 POR2X1_188/A POR2X1_710/O 0.01fF
C14741 INPUT_1 POR2X1_817/O 0.01fF
C14742 PAND2X1_793/Y PAND2X1_738/Y 0.26fF
C14743 PAND2X1_845/a_76_28# POR2X1_60/A 0.00fF
C14744 PAND2X1_57/B POR2X1_121/Y 0.01fF
C14745 PAND2X1_274/a_16_344# PAND2X1_480/B 0.06fF
C14746 POR2X1_814/B POR2X1_789/A 0.03fF
C14747 PAND2X1_731/B POR2X1_90/Y 0.01fF
C14748 POR2X1_614/A POR2X1_549/CTRL 0.04fF
C14749 POR2X1_614/A POR2X1_814/B 0.10fF
C14750 POR2X1_389/CTRL POR2X1_130/A 0.32fF
C14751 POR2X1_466/O VDD 0.00fF
C14752 POR2X1_379/a_16_28# POR2X1_66/A 0.04fF
C14753 PAND2X1_662/CTRL PAND2X1_660/B 0.01fF
C14754 POR2X1_343/A PAND2X1_69/A 0.01fF
C14755 PAND2X1_436/O POR2X1_129/Y 0.02fF
C14756 PAND2X1_820/CTRL POR2X1_669/B 0.01fF
C14757 POR2X1_102/Y PAND2X1_349/A 0.04fF
C14758 POR2X1_624/Y POR2X1_620/B 0.02fF
C14759 PAND2X1_39/B POR2X1_398/a_16_28# 0.09fF
C14760 POR2X1_121/a_16_28# POR2X1_590/A 0.02fF
C14761 PAND2X1_480/O PAND2X1_776/Y 0.06fF
C14762 POR2X1_260/B POR2X1_774/A 0.03fF
C14763 POR2X1_166/O POR2X1_40/Y 0.01fF
C14764 POR2X1_68/A POR2X1_797/O 0.01fF
C14765 POR2X1_13/A POR2X1_494/Y 0.04fF
C14766 PAND2X1_808/Y PAND2X1_580/B 0.02fF
C14767 POR2X1_96/A PAND2X1_758/CTRL 0.01fF
C14768 PAND2X1_46/CTRL2 PAND2X1_111/B 0.01fF
C14769 POR2X1_72/B PAND2X1_168/CTRL2 0.01fF
C14770 PAND2X1_65/B POR2X1_631/B 0.01fF
C14771 PAND2X1_714/A POR2X1_73/Y 0.00fF
C14772 POR2X1_814/B POR2X1_38/B 0.10fF
C14773 PAND2X1_30/CTRL2 POR2X1_451/A 0.01fF
C14774 POR2X1_102/Y PAND2X1_114/B 0.03fF
C14775 POR2X1_401/A VDD -0.00fF
C14776 PAND2X1_96/B POR2X1_675/A 0.04fF
C14777 PAND2X1_339/Y VDD 0.00fF
C14778 PAND2X1_564/B PAND2X1_569/B 0.08fF
C14779 POR2X1_303/CTRL2 POR2X1_274/A 0.02fF
C14780 POR2X1_332/B POR2X1_741/Y 0.03fF
C14781 POR2X1_614/A POR2X1_325/A 0.03fF
C14782 PAND2X1_473/CTRL2 PAND2X1_473/B 0.03fF
C14783 POR2X1_814/B POR2X1_360/CTRL2 0.01fF
C14784 PAND2X1_580/O VDD 0.00fF
C14785 PAND2X1_735/CTRL POR2X1_816/A 0.01fF
C14786 PAND2X1_20/A PAND2X1_297/O 0.04fF
C14787 POR2X1_383/A POR2X1_94/A 0.01fF
C14788 POR2X1_817/A POR2X1_382/O 0.03fF
C14789 POR2X1_543/A PAND2X1_312/O 0.02fF
C14790 PAND2X1_579/B POR2X1_816/A 0.03fF
C14791 POR2X1_327/O POR2X1_572/B 0.01fF
C14792 PAND2X1_591/CTRL PAND2X1_48/A 0.03fF
C14793 PAND2X1_408/Y VDD 0.10fF
C14794 PAND2X1_651/Y INPUT_0 0.13fF
C14795 POR2X1_407/Y POR2X1_770/A 0.00fF
C14796 PAND2X1_107/CTRL2 POR2X1_640/Y 0.01fF
C14797 POR2X1_178/O PAND2X1_738/Y 0.12fF
C14798 POR2X1_278/Y POR2X1_52/Y 0.05fF
C14799 POR2X1_136/CTRL PAND2X1_480/B 0.28fF
C14800 POR2X1_687/A POR2X1_330/Y 0.17fF
C14801 POR2X1_852/B POR2X1_854/B 0.10fF
C14802 PAND2X1_865/Y POR2X1_437/O 0.00fF
C14803 POR2X1_790/B PAND2X1_753/O 0.01fF
C14804 PAND2X1_55/Y POR2X1_740/Y 0.08fF
C14805 POR2X1_332/B PAND2X1_32/B 0.12fF
C14806 PAND2X1_498/a_16_344# POR2X1_733/A 0.02fF
C14807 POR2X1_254/Y POR2X1_203/Y 0.03fF
C14808 PAND2X1_794/B POR2X1_7/B 0.03fF
C14809 PAND2X1_824/B PAND2X1_420/CTRL 0.05fF
C14810 POR2X1_538/a_16_28# PAND2X1_57/B 0.01fF
C14811 PAND2X1_562/B PAND2X1_348/CTRL2 0.03fF
C14812 POR2X1_65/A PAND2X1_264/CTRL2 0.03fF
C14813 POR2X1_382/O POR2X1_42/Y 0.34fF
C14814 POR2X1_78/B PAND2X1_393/CTRL2 0.01fF
C14815 POR2X1_646/CTRL2 PAND2X1_32/B 0.03fF
C14816 PAND2X1_96/B POR2X1_220/Y 0.10fF
C14817 PAND2X1_94/A PAND2X1_42/CTRL 0.01fF
C14818 POR2X1_667/A POR2X1_153/Y 0.07fF
C14819 POR2X1_60/A POR2X1_394/A 1.61fF
C14820 POR2X1_130/A POR2X1_361/CTRL2 0.12fF
C14821 PAND2X1_632/A POR2X1_5/Y 0.03fF
C14822 PAND2X1_216/B PAND2X1_561/A 0.00fF
C14823 POR2X1_864/A PAND2X1_72/A 0.03fF
C14824 POR2X1_114/Y POR2X1_68/B 0.15fF
C14825 POR2X1_16/A POR2X1_492/O 0.01fF
C14826 PAND2X1_732/A PAND2X1_731/B 0.01fF
C14827 POR2X1_763/A POR2X1_158/B 0.07fF
C14828 POR2X1_432/a_16_28# POR2X1_129/Y 0.09fF
C14829 PAND2X1_551/A PAND2X1_324/Y 0.01fF
C14830 PAND2X1_556/B POR2X1_387/Y 0.03fF
C14831 POR2X1_66/A POR2X1_703/m4_208_n4# 0.08fF
C14832 PAND2X1_569/B PAND2X1_544/CTRL2 0.01fF
C14833 PAND2X1_564/CTRL2 POR2X1_765/Y 0.01fF
C14834 POR2X1_591/A POR2X1_394/A 0.02fF
C14835 POR2X1_582/CTRL INPUT_5 0.01fF
C14836 POR2X1_582/O INPUT_4 0.01fF
C14837 INPUT_1 POR2X1_585/CTRL 0.01fF
C14838 PAND2X1_865/Y PAND2X1_811/A 0.44fF
C14839 PAND2X1_96/B POR2X1_404/Y 0.40fF
C14840 PAND2X1_6/Y PAND2X1_275/CTRL 0.00fF
C14841 PAND2X1_793/Y PAND2X1_575/O 0.02fF
C14842 POR2X1_52/O PAND2X1_124/Y 0.01fF
C14843 POR2X1_62/Y POR2X1_14/Y 0.03fF
C14844 POR2X1_43/B PAND2X1_523/m4_208_n4# 0.04fF
C14845 POR2X1_538/A VDD 0.05fF
C14846 POR2X1_188/A POR2X1_851/CTRL 0.01fF
C14847 POR2X1_800/A POR2X1_796/O 0.00fF
C14848 POR2X1_68/A POR2X1_114/B 0.05fF
C14849 POR2X1_567/B POR2X1_510/CTRL 0.13fF
C14850 PAND2X1_658/A POR2X1_816/A 0.04fF
C14851 PAND2X1_689/O POR2X1_691/A 0.01fF
C14852 POR2X1_786/A POR2X1_84/Y 0.01fF
C14853 POR2X1_154/CTRL2 POR2X1_855/B 0.01fF
C14854 PAND2X1_6/Y POR2X1_691/O 0.16fF
C14855 POR2X1_582/A INPUT_5 0.01fF
C14856 PAND2X1_13/CTRL2 POR2X1_186/B 0.01fF
C14857 PAND2X1_813/O POR2X1_5/Y 0.01fF
C14858 PAND2X1_319/B PAND2X1_724/B 0.02fF
C14859 PAND2X1_613/CTRL2 PAND2X1_52/B 0.12fF
C14860 POR2X1_507/O VDD 0.00fF
C14861 POR2X1_809/A POR2X1_750/B 0.02fF
C14862 POR2X1_465/B POR2X1_510/Y 0.03fF
C14863 POR2X1_130/A POR2X1_249/Y 0.05fF
C14864 PAND2X1_55/Y PAND2X1_312/CTRL2 0.01fF
C14865 POR2X1_220/B POR2X1_568/B 0.20fF
C14866 PAND2X1_401/O POR2X1_73/Y 0.08fF
C14867 PAND2X1_552/B PAND2X1_388/O 0.17fF
C14868 PAND2X1_52/Y POR2X1_186/B 0.03fF
C14869 POR2X1_362/A VDD 0.00fF
C14870 POR2X1_415/CTRL POR2X1_750/Y 0.01fF
C14871 POR2X1_212/A POR2X1_568/A 0.01fF
C14872 POR2X1_702/B POR2X1_186/B 0.00fF
C14873 POR2X1_40/Y PAND2X1_730/A 0.00fF
C14874 POR2X1_383/A PAND2X1_110/CTRL2 0.09fF
C14875 PAND2X1_652/CTRL POR2X1_83/B 0.01fF
C14876 PAND2X1_726/B VDD 0.02fF
C14877 POR2X1_733/A PAND2X1_60/B 0.05fF
C14878 POR2X1_164/a_16_28# POR2X1_693/Y 0.02fF
C14879 POR2X1_68/A PAND2X1_424/CTRL 0.08fF
C14880 PAND2X1_47/CTRL2 PAND2X1_32/B 0.01fF
C14881 POR2X1_334/B PAND2X1_60/B 0.05fF
C14882 POR2X1_164/Y POR2X1_46/Y 0.03fF
C14883 POR2X1_8/Y POR2X1_381/m4_208_n4# 0.12fF
C14884 POR2X1_124/CTRL POR2X1_276/Y 0.16fF
C14885 POR2X1_73/Y POR2X1_816/A 0.04fF
C14886 POR2X1_327/Y POR2X1_733/O 0.37fF
C14887 POR2X1_22/CTRL2 POR2X1_260/A 0.04fF
C14888 PAND2X1_569/A POR2X1_73/Y 0.03fF
C14889 PAND2X1_408/Y PAND2X1_32/B 0.01fF
C14890 PAND2X1_499/Y POR2X1_129/Y 0.03fF
C14891 POR2X1_112/CTRL POR2X1_750/B 0.27fF
C14892 POR2X1_383/A POR2X1_340/O 0.01fF
C14893 POR2X1_78/B POR2X1_398/CTRL2 0.01fF
C14894 POR2X1_383/A POR2X1_861/CTRL2 0.01fF
C14895 POR2X1_458/CTRL2 POR2X1_343/B 0.01fF
C14896 POR2X1_494/Y PAND2X1_510/B 0.02fF
C14897 PAND2X1_63/Y POR2X1_68/B 0.03fF
C14898 POR2X1_41/B POR2X1_16/A 3.17fF
C14899 POR2X1_804/A POR2X1_541/O 0.05fF
C14900 POR2X1_844/O POR2X1_844/B 0.00fF
C14901 POR2X1_305/Y POR2X1_239/Y 0.01fF
C14902 POR2X1_741/Y POR2X1_574/A 0.03fF
C14903 POR2X1_220/B POR2X1_161/CTRL2 0.03fF
C14904 POR2X1_337/A POR2X1_740/Y 0.10fF
C14905 POR2X1_538/A POR2X1_741/Y 0.03fF
C14906 PAND2X1_821/O POR2X1_854/B 0.02fF
C14907 PAND2X1_199/A PAND2X1_199/B 0.18fF
C14908 PAND2X1_382/CTRL2 POR2X1_816/A 0.10fF
C14909 PAND2X1_632/B POR2X1_252/a_16_28# 0.02fF
C14910 POR2X1_68/A POR2X1_222/A 0.01fF
C14911 POR2X1_186/Y PAND2X1_680/a_16_344# 0.04fF
C14912 PAND2X1_4/CTRL POR2X1_38/B 0.01fF
C14913 PAND2X1_489/CTRL2 PAND2X1_798/B 0.02fF
C14914 PAND2X1_363/a_56_28# POR2X1_42/Y 0.00fF
C14915 PAND2X1_404/Y POR2X1_825/Y 0.02fF
C14916 POR2X1_416/B POR2X1_516/Y 0.03fF
C14917 POR2X1_71/CTRL2 POR2X1_293/Y 0.13fF
C14918 POR2X1_730/Y POR2X1_732/B 0.00fF
C14919 POR2X1_113/Y POR2X1_68/B 0.23fF
C14920 POR2X1_208/Y POR2X1_201/Y 0.07fF
C14921 PAND2X1_23/Y PAND2X1_300/m4_208_n4# 0.07fF
C14922 PAND2X1_840/A PAND2X1_840/a_76_28# 0.05fF
C14923 POR2X1_252/O POR2X1_153/Y 0.02fF
C14924 INPUT_0 POR2X1_294/A 0.20fF
C14925 PAND2X1_764/O PAND2X1_32/B 0.03fF
C14926 PAND2X1_854/A POR2X1_73/Y 0.03fF
C14927 PAND2X1_244/B POR2X1_816/A 0.03fF
C14928 POR2X1_580/CTRL POR2X1_191/Y 0.11fF
C14929 PAND2X1_662/O PAND2X1_660/Y -0.00fF
C14930 PAND2X1_41/B POR2X1_182/a_16_28# 0.02fF
C14931 POR2X1_68/A POR2X1_551/O 0.08fF
C14932 PAND2X1_57/B PAND2X1_3/B 0.16fF
C14933 POR2X1_220/A POR2X1_161/Y 0.01fF
C14934 POR2X1_750/B POR2X1_711/Y 0.07fF
C14935 POR2X1_234/A POR2X1_37/Y 0.05fF
C14936 PAND2X1_469/B PAND2X1_715/B 0.25fF
C14937 D_INPUT_7 PAND2X1_581/CTRL2 0.03fF
C14938 PAND2X1_778/a_76_28# PAND2X1_506/Y 0.05fF
C14939 PAND2X1_390/CTRL PAND2X1_853/B 0.12fF
C14940 PAND2X1_793/A POR2X1_39/B 0.01fF
C14941 PAND2X1_385/CTRL2 PAND2X1_48/A 0.01fF
C14942 PAND2X1_55/Y POR2X1_774/A 0.07fF
C14943 POR2X1_625/CTRL2 POR2X1_39/B 0.03fF
C14944 PAND2X1_639/Y PAND2X1_636/O 0.00fF
C14945 POR2X1_62/Y PAND2X1_341/CTRL2 0.01fF
C14946 PAND2X1_469/B PAND2X1_303/Y 0.34fF
C14947 POR2X1_804/A POR2X1_675/Y 0.03fF
C14948 POR2X1_567/B POR2X1_440/CTRL 0.27fF
C14949 PAND2X1_242/Y POR2X1_669/B 0.10fF
C14950 POR2X1_750/B POR2X1_728/A 0.01fF
C14951 POR2X1_554/B POR2X1_556/A 0.03fF
C14952 POR2X1_96/A PAND2X1_643/A 0.03fF
C14953 PAND2X1_56/Y POR2X1_334/Y 0.10fF
C14954 POR2X1_62/Y POR2X1_55/Y 0.23fF
C14955 POR2X1_101/Y POR2X1_318/A 0.10fF
C14956 POR2X1_541/B PAND2X1_256/a_16_344# 0.02fF
C14957 POR2X1_833/A PAND2X1_69/A 0.01fF
C14958 POR2X1_717/O POR2X1_390/B 0.00fF
C14959 POR2X1_119/Y PAND2X1_466/CTRL2 0.03fF
C14960 POR2X1_68/B POR2X1_260/A 0.23fF
C14961 POR2X1_511/Y POR2X1_39/B 0.43fF
C14962 PAND2X1_535/Y PAND2X1_539/Y 0.01fF
C14963 PAND2X1_96/B PAND2X1_184/O 0.19fF
C14964 PAND2X1_96/B POR2X1_332/CTRL 0.00fF
C14965 POR2X1_814/A POR2X1_862/A 0.45fF
C14966 INPUT_0 PAND2X1_102/CTRL 0.01fF
C14967 PAND2X1_858/CTRL POR2X1_43/B 0.01fF
C14968 POR2X1_222/Y POR2X1_735/O 0.01fF
C14969 POR2X1_834/Y POR2X1_513/CTRL 0.30fF
C14970 PAND2X1_569/B PAND2X1_374/CTRL2 0.00fF
C14971 PAND2X1_6/Y POR2X1_339/Y 0.03fF
C14972 PAND2X1_649/A POR2X1_293/Y 0.00fF
C14973 POR2X1_651/Y PAND2X1_58/A 0.03fF
C14974 POR2X1_108/CTRL PAND2X1_348/A 0.04fF
C14975 PAND2X1_408/CTRL PAND2X1_18/B 0.01fF
C14976 POR2X1_283/A PAND2X1_175/O 0.04fF
C14977 POR2X1_614/A POR2X1_332/Y 0.02fF
C14978 POR2X1_553/A POR2X1_569/A 0.07fF
C14979 POR2X1_119/Y PAND2X1_478/O 0.17fF
C14980 POR2X1_594/CTRL2 POR2X1_594/A 0.01fF
C14981 POR2X1_23/Y POR2X1_441/O 0.02fF
C14982 INPUT_1 POR2X1_245/Y 0.03fF
C14983 POR2X1_407/Y POR2X1_774/A 0.03fF
C14984 PAND2X1_23/Y PAND2X1_122/CTRL 0.06fF
C14985 D_GATE_222 POR2X1_191/Y 0.10fF
C14986 INPUT_0 PAND2X1_858/B 0.08fF
C14987 POR2X1_150/Y POR2X1_679/A 0.00fF
C14988 POR2X1_10/O POR2X1_7/A 0.01fF
C14989 POR2X1_740/Y POR2X1_738/O 0.00fF
C14990 POR2X1_724/A POR2X1_186/B 0.07fF
C14991 POR2X1_43/B PAND2X1_500/CTRL2 0.01fF
C14992 POR2X1_16/A PAND2X1_100/CTRL2 0.00fF
C14993 PAND2X1_830/CTRL PAND2X1_348/A 0.02fF
C14994 POR2X1_407/Y PAND2X1_328/CTRL 0.01fF
C14995 POR2X1_614/A PAND2X1_680/O 0.17fF
C14996 POR2X1_532/A POR2X1_735/O 0.02fF
C14997 PAND2X1_862/B POR2X1_80/O 0.00fF
C14998 POR2X1_738/A POR2X1_731/A 0.00fF
C14999 PAND2X1_659/Y PAND2X1_473/O 0.01fF
C15000 POR2X1_780/A POR2X1_294/A 0.18fF
C15001 PAND2X1_73/Y POR2X1_814/A 0.18fF
C15002 POR2X1_383/A POR2X1_334/Y 0.19fF
C15003 POR2X1_57/A POR2X1_385/Y 0.05fF
C15004 PAND2X1_804/B POR2X1_173/CTRL2 0.05fF
C15005 PAND2X1_108/CTRL PAND2X1_55/Y 0.05fF
C15006 PAND2X1_393/CTRL2 POR2X1_294/A 0.00fF
C15007 PAND2X1_138/CTRL2 POR2X1_7/A 0.00fF
C15008 POR2X1_775/A POR2X1_632/Y 0.03fF
C15009 PAND2X1_404/Y POR2X1_490/a_16_28# 0.00fF
C15010 PAND2X1_220/CTRL POR2X1_77/Y 0.00fF
C15011 POR2X1_16/A PAND2X1_308/Y 0.00fF
C15012 POR2X1_67/Y PAND2X1_58/A 0.06fF
C15013 POR2X1_394/A POR2X1_744/CTRL 0.01fF
C15014 PAND2X1_835/CTRL2 POR2X1_77/Y 0.00fF
C15015 PAND2X1_96/B POR2X1_554/CTRL 0.01fF
C15016 POR2X1_383/A PAND2X1_281/O 0.02fF
C15017 POR2X1_263/a_56_344# POR2X1_37/Y 0.00fF
C15018 PAND2X1_600/O PAND2X1_39/B 0.06fF
C15019 PAND2X1_93/B POR2X1_624/Y 0.07fF
C15020 POR2X1_327/Y POR2X1_860/O 0.01fF
C15021 PAND2X1_450/CTRL POR2X1_416/B 0.01fF
C15022 PAND2X1_797/Y PAND2X1_213/Y 0.02fF
C15023 POR2X1_102/Y POR2X1_411/A 0.12fF
C15024 POR2X1_632/Y POR2X1_112/Y 0.03fF
C15025 POR2X1_471/A POR2X1_466/A 1.16fF
C15026 POR2X1_539/A POR2X1_567/A 0.08fF
C15027 POR2X1_775/A PAND2X1_52/B 0.03fF
C15028 POR2X1_669/B PAND2X1_750/CTRL2 0.43fF
C15029 POR2X1_691/O PAND2X1_52/B 0.01fF
C15030 PAND2X1_476/A PAND2X1_723/A 0.01fF
C15031 PAND2X1_482/CTRL2 POR2X1_186/B 0.01fF
C15032 POR2X1_234/A POR2X1_293/Y 0.00fF
C15033 POR2X1_856/B POR2X1_446/O 0.04fF
C15034 POR2X1_66/A PAND2X1_27/a_16_344# 0.09fF
C15035 PAND2X1_287/Y PAND2X1_771/Y 0.05fF
C15036 PAND2X1_39/B POR2X1_590/A 1.14fF
C15037 PAND2X1_860/A PAND2X1_592/Y 0.03fF
C15038 POR2X1_78/A POR2X1_624/Y 0.06fF
C15039 PAND2X1_340/B POR2X1_32/A 0.03fF
C15040 POR2X1_294/A POR2X1_398/CTRL2 0.00fF
C15041 PAND2X1_221/Y POR2X1_7/B 11.34fF
C15042 PAND2X1_849/CTRL2 POR2X1_20/B 0.01fF
C15043 POR2X1_13/A POR2X1_667/CTRL 0.01fF
C15044 POR2X1_502/A PAND2X1_53/CTRL2 0.02fF
C15045 POR2X1_39/B PAND2X1_124/O 0.15fF
C15046 PAND2X1_52/B POR2X1_162/Y 0.05fF
C15047 POR2X1_841/B PAND2X1_58/A 0.03fF
C15048 POR2X1_568/Y POR2X1_568/m4_208_n4# 0.07fF
C15049 POR2X1_846/A POR2X1_789/Y 0.01fF
C15050 POR2X1_66/A POR2X1_29/A 0.05fF
C15051 POR2X1_54/Y POR2X1_615/CTRL 0.01fF
C15052 POR2X1_687/B POR2X1_814/A 0.05fF
C15053 PAND2X1_640/B POR2X1_83/B 0.03fF
C15054 POR2X1_54/Y PAND2X1_395/CTRL2 0.09fF
C15055 POR2X1_16/A POR2X1_77/Y 0.40fF
C15056 PAND2X1_600/O PAND2X1_20/A 0.15fF
C15057 POR2X1_23/Y PAND2X1_76/CTRL2 0.03fF
C15058 POR2X1_16/A POR2X1_85/Y 0.03fF
C15059 PAND2X1_425/Y VDD 0.07fF
C15060 POR2X1_133/CTRL2 POR2X1_411/B 0.01fF
C15061 POR2X1_624/Y POR2X1_573/CTRL 0.01fF
C15062 POR2X1_29/O PAND2X1_9/Y 0.01fF
C15063 POR2X1_129/Y POR2X1_39/B 0.26fF
C15064 POR2X1_13/A POR2X1_603/CTRL 0.01fF
C15065 POR2X1_102/Y POR2X1_32/A 0.19fF
C15066 POR2X1_805/Y POR2X1_590/A 0.00fF
C15067 POR2X1_509/A POR2X1_814/A 0.02fF
C15068 POR2X1_48/A PAND2X1_541/CTRL 0.01fF
C15069 POR2X1_78/B POR2X1_648/O 0.01fF
C15070 POR2X1_60/A POR2X1_669/B 0.14fF
C15071 POR2X1_263/Y POR2X1_40/Y 0.07fF
C15072 POR2X1_602/B POR2X1_66/A 0.06fF
C15073 PAND2X1_20/A POR2X1_590/A 0.13fF
C15074 POR2X1_421/Y POR2X1_422/Y 0.01fF
C15075 POR2X1_15/CTRL POR2X1_9/Y 0.01fF
C15076 PAND2X1_475/a_16_344# D_INPUT_0 0.02fF
C15077 POR2X1_304/Y PAND2X1_454/B 0.13fF
C15078 PAND2X1_39/B PAND2X1_760/CTRL 0.01fF
C15079 PAND2X1_600/O POR2X1_814/B 0.06fF
C15080 PAND2X1_659/Y POR2X1_39/B 0.03fF
C15081 POR2X1_263/a_16_28# PAND2X1_35/Y 0.02fF
C15082 PAND2X1_669/a_16_344# POR2X1_750/B 0.01fF
C15083 POR2X1_634/A POR2X1_769/A 0.04fF
C15084 POR2X1_290/Y POR2X1_411/B 0.03fF
C15085 POR2X1_864/a_16_28# POR2X1_801/B 0.05fF
C15086 POR2X1_117/CTRL2 POR2X1_409/B 0.01fF
C15087 POR2X1_814/A POR2X1_631/B 0.07fF
C15088 PAND2X1_35/A VDD 0.15fF
C15089 D_INPUT_0 PAND2X1_525/CTRL2 0.01fF
C15090 PAND2X1_299/O D_INPUT_0 0.01fF
C15091 POR2X1_46/a_16_28# POR2X1_409/B 0.02fF
C15092 PAND2X1_285/a_76_28# PAND2X1_805/A 0.01fF
C15093 POR2X1_49/Y PAND2X1_623/CTRL2 0.10fF
C15094 POR2X1_677/Y PAND2X1_349/A 0.02fF
C15095 POR2X1_814/A POR2X1_784/CTRL2 0.06fF
C15096 POR2X1_496/Y POR2X1_423/Y 1.01fF
C15097 POR2X1_119/CTRL POR2X1_411/B 0.01fF
C15098 POR2X1_65/O PAND2X1_6/A 0.02fF
C15099 POR2X1_77/Y PAND2X1_336/Y 0.03fF
C15100 PAND2X1_68/CTRL2 POR2X1_5/Y 0.05fF
C15101 POR2X1_417/Y POR2X1_102/Y 0.02fF
C15102 POR2X1_102/Y POR2X1_419/Y 0.23fF
C15103 POR2X1_96/Y POR2X1_39/B 0.03fF
C15104 POR2X1_48/A POR2X1_511/Y 0.03fF
C15105 POR2X1_582/Y INPUT_5 0.01fF
C15106 POR2X1_428/Y INPUT_4 0.03fF
C15107 PAND2X1_240/a_16_344# D_INPUT_0 0.02fF
C15108 POR2X1_9/Y PAND2X1_63/B 0.07fF
C15109 POR2X1_48/A POR2X1_524/Y 0.01fF
C15110 POR2X1_156/CTRL2 POR2X1_728/A 0.00fF
C15111 POR2X1_590/A PAND2X1_525/CTRL 0.01fF
C15112 POR2X1_37/Y PAND2X1_499/Y 0.08fF
C15113 PAND2X1_299/CTRL POR2X1_121/B 0.01fF
C15114 POR2X1_411/B PAND2X1_658/B 0.05fF
C15115 POR2X1_19/CTRL2 D_INPUT_1 0.03fF
C15116 POR2X1_814/B POR2X1_590/A 0.26fF
C15117 POR2X1_496/Y PAND2X1_513/a_16_344# 0.03fF
C15118 POR2X1_407/A POR2X1_499/A 0.03fF
C15119 POR2X1_670/CTRL2 POR2X1_102/Y 0.00fF
C15120 POR2X1_499/CTRL VDD 0.00fF
C15121 PAND2X1_832/O PAND2X1_435/Y 0.01fF
C15122 POR2X1_68/A PAND2X1_761/CTRL2 0.10fF
C15123 PAND2X1_57/B PAND2X1_248/O 0.01fF
C15124 PAND2X1_42/a_16_344# POR2X1_590/A 0.01fF
C15125 PAND2X1_658/A INPUT_3 0.59fF
C15126 POR2X1_699/CTRL2 POR2X1_7/B 0.03fF
C15127 PAND2X1_862/B POR2X1_23/Y 0.06fF
C15128 POR2X1_415/A POR2X1_415/Y 0.02fF
C15129 PAND2X1_6/Y POR2X1_541/B 0.09fF
C15130 PAND2X1_55/Y PAND2X1_67/O 0.02fF
C15131 POR2X1_590/A POR2X1_733/CTRL 0.01fF
C15132 POR2X1_814/A PAND2X1_163/O 0.37fF
C15133 POR2X1_556/A POR2X1_702/A 0.03fF
C15134 POR2X1_66/A POR2X1_546/A 0.09fF
C15135 POR2X1_841/O POR2X1_513/Y 0.07fF
C15136 POR2X1_846/A POR2X1_789/B 0.02fF
C15137 POR2X1_411/B PAND2X1_577/O 0.02fF
C15138 POR2X1_169/B POR2X1_568/A 0.01fF
C15139 POR2X1_590/A POR2X1_325/A 0.03fF
C15140 POR2X1_428/Y POR2X1_426/CTRL 0.09fF
C15141 POR2X1_307/B PAND2X1_58/A 0.10fF
C15142 POR2X1_78/Y PAND2X1_79/Y 0.10fF
C15143 PAND2X1_72/A PAND2X1_179/CTRL 0.00fF
C15144 POR2X1_257/A POR2X1_255/Y 0.61fF
C15145 PAND2X1_816/a_16_344# POR2X1_862/A 0.04fF
C15146 PAND2X1_93/B POR2X1_785/A 0.03fF
C15147 POR2X1_102/Y PAND2X1_741/B 0.02fF
C15148 POR2X1_498/a_56_344# D_INPUT_0 0.00fF
C15149 POR2X1_140/B POR2X1_76/A 0.03fF
C15150 POR2X1_748/A POR2X1_5/Y 0.03fF
C15151 POR2X1_315/Y PAND2X1_464/B 0.01fF
C15152 POR2X1_49/Y PAND2X1_61/Y 2.01fF
C15153 POR2X1_687/B POR2X1_687/O 0.00fF
C15154 POR2X1_554/B POR2X1_276/A 0.03fF
C15155 POR2X1_661/Y POR2X1_722/Y 0.17fF
C15156 PAND2X1_6/Y PAND2X1_422/a_76_28# 0.01fF
C15157 POR2X1_658/a_16_28# POR2X1_318/A 0.08fF
C15158 PAND2X1_265/O INPUT_0 0.17fF
C15159 PAND2X1_72/A D_INPUT_4 0.03fF
C15160 INPUT_2 POR2X1_126/O 0.01fF
C15161 POR2X1_835/Y POR2X1_506/B 0.68fF
C15162 POR2X1_65/A POR2X1_760/CTRL2 0.00fF
C15163 POR2X1_376/B PAND2X1_333/CTRL 0.05fF
C15164 POR2X1_41/B POR2X1_142/CTRL2 0.13fF
C15165 POR2X1_728/CTRL POR2X1_330/Y 0.04fF
C15166 POR2X1_66/A POR2X1_204/CTRL2 0.02fF
C15167 POR2X1_29/A POR2X1_494/Y 0.01fF
C15168 POR2X1_81/A PAND2X1_242/Y 0.12fF
C15169 POR2X1_174/B POR2X1_356/A 0.23fF
C15170 POR2X1_83/B POR2X1_7/B 0.98fF
C15171 POR2X1_247/Y POR2X1_294/B 0.01fF
C15172 POR2X1_94/A INPUT_0 1.06fF
C15173 POR2X1_78/A POR2X1_785/A 0.10fF
C15174 PAND2X1_240/CTRL VDD 0.00fF
C15175 POR2X1_66/A POR2X1_712/Y 0.03fF
C15176 POR2X1_511/Y PAND2X1_513/O 0.03fF
C15177 PAND2X1_20/A POR2X1_857/B 0.03fF
C15178 POR2X1_863/A PAND2X1_167/a_76_28# 0.01fF
C15179 POR2X1_174/A POR2X1_740/Y 0.02fF
C15180 POR2X1_14/Y POR2X1_395/O 0.01fF
C15181 PAND2X1_82/m4_208_n4# PAND2X1_83/m4_208_n4# 0.05fF
C15182 POR2X1_855/B POR2X1_803/O 0.01fF
C15183 POR2X1_48/A PAND2X1_324/O 0.08fF
C15184 POR2X1_220/Y POR2X1_355/A 0.03fF
C15185 POR2X1_60/A PAND2X1_174/CTRL 0.02fF
C15186 POR2X1_655/A PAND2X1_305/CTRL 0.01fF
C15187 POR2X1_449/O PAND2X1_90/Y 0.04fF
C15188 POR2X1_236/O POR2X1_236/Y 0.02fF
C15189 POR2X1_41/B POR2X1_495/O 0.06fF
C15190 PAND2X1_340/B POR2X1_503/Y 0.02fF
C15191 PAND2X1_32/CTRL POR2X1_294/A 0.01fF
C15192 PAND2X1_284/Y PAND2X1_771/Y 0.20fF
C15193 POR2X1_148/a_16_28# POR2X1_148/A 0.06fF
C15194 POR2X1_99/A POR2X1_404/Y 0.03fF
C15195 POR2X1_118/CTRL POR2X1_32/A 0.01fF
C15196 PAND2X1_463/O POR2X1_7/B 0.15fF
C15197 PAND2X1_215/B POR2X1_40/Y 1.72fF
C15198 PAND2X1_630/B PAND2X1_508/B 0.28fF
C15199 POR2X1_96/A PAND2X1_231/O 0.01fF
C15200 POR2X1_849/O POR2X1_859/A 0.02fF
C15201 POR2X1_753/Y POR2X1_816/A 0.14fF
C15202 PAND2X1_96/B PAND2X1_594/CTRL 0.01fF
C15203 POR2X1_102/Y POR2X1_184/Y 0.07fF
C15204 D_INPUT_0 POR2X1_38/Y 0.17fF
C15205 D_GATE_865 VDD 0.05fF
C15206 POR2X1_462/B POR2X1_753/Y 0.10fF
C15207 POR2X1_96/A PAND2X1_805/A 0.03fF
C15208 PAND2X1_474/Y POR2X1_497/Y 0.03fF
C15209 POR2X1_114/B PAND2X1_58/A 0.04fF
C15210 D_INPUT_0 POR2X1_140/O 0.07fF
C15211 POR2X1_832/Y POR2X1_725/Y 0.12fF
C15212 PAND2X1_55/Y POR2X1_202/CTRL 0.01fF
C15213 POR2X1_364/A POR2X1_241/B 0.03fF
C15214 POR2X1_697/Y POR2X1_72/B 1.19fF
C15215 PAND2X1_467/B POR2X1_694/CTRL2 0.01fF
C15216 PAND2X1_349/B POR2X1_55/Y 0.09fF
C15217 POR2X1_504/Y POR2X1_628/CTRL 0.01fF
C15218 PAND2X1_520/O POR2X1_236/Y 0.02fF
C15219 PAND2X1_477/B POR2X1_83/B 0.47fF
C15220 PAND2X1_859/A PAND2X1_859/B 0.44fF
C15221 PAND2X1_651/Y POR2X1_102/Y 0.08fF
C15222 PAND2X1_23/Y POR2X1_389/Y 0.07fF
C15223 POR2X1_13/A POR2X1_497/Y 0.03fF
C15224 POR2X1_532/A POR2X1_29/A 0.04fF
C15225 POR2X1_376/Y PAND2X1_375/CTRL2 0.03fF
C15226 PAND2X1_20/A POR2X1_574/a_76_344# 0.00fF
C15227 POR2X1_407/A POR2X1_783/CTRL 0.00fF
C15228 POR2X1_60/A PAND2X1_370/O 0.04fF
C15229 PAND2X1_466/m4_208_n4# PAND2X1_446/m4_208_n4# 0.05fF
C15230 POR2X1_260/B POR2X1_750/Y 0.05fF
C15231 PAND2X1_20/A PAND2X1_752/Y 0.28fF
C15232 POR2X1_66/B PAND2X1_6/Y 0.21fF
C15233 POR2X1_763/A POR2X1_700/CTRL2 0.05fF
C15234 PAND2X1_798/B PAND2X1_354/A 0.02fF
C15235 POR2X1_278/Y PAND2X1_580/B 0.03fF
C15236 PAND2X1_848/O POR2X1_38/B 0.01fF
C15237 POR2X1_365/Y POR2X1_353/Y 0.00fF
C15238 POR2X1_502/A POR2X1_794/CTRL 0.00fF
C15239 POR2X1_251/A PAND2X1_357/Y 0.09fF
C15240 POR2X1_188/A PAND2X1_536/O 0.02fF
C15241 POR2X1_43/B PAND2X1_217/B 0.05fF
C15242 POR2X1_400/A POR2X1_214/O 0.00fF
C15243 POR2X1_792/CTRL PAND2X1_60/B 0.01fF
C15244 PAND2X1_626/CTRL PAND2X1_96/B 0.00fF
C15245 PAND2X1_6/A POR2X1_40/Y 0.19fF
C15246 PAND2X1_805/CTRL POR2X1_7/B 0.09fF
C15247 POR2X1_760/A PAND2X1_643/A 0.03fF
C15248 PAND2X1_422/CTRL2 POR2X1_296/B 0.05fF
C15249 PAND2X1_830/Y PAND2X1_140/Y 0.03fF
C15250 POR2X1_333/A POR2X1_210/Y 0.43fF
C15251 POR2X1_188/A PAND2X1_6/Y 0.03fF
C15252 POR2X1_864/O PAND2X1_32/B 0.01fF
C15253 POR2X1_35/B PAND2X1_6/A 0.21fF
C15254 PAND2X1_283/O POR2X1_654/B 0.01fF
C15255 POR2X1_78/B PAND2X1_322/a_16_344# 0.02fF
C15256 PAND2X1_473/Y POR2X1_46/Y 0.03fF
C15257 POR2X1_446/B POR2X1_724/B 0.01fF
C15258 POR2X1_252/CTRL VDD 0.00fF
C15259 PAND2X1_479/A PAND2X1_479/B 0.02fF
C15260 POR2X1_566/A PAND2X1_524/CTRL2 0.12fF
C15261 POR2X1_848/A POR2X1_260/A 0.07fF
C15262 POR2X1_335/A POR2X1_105/Y 0.03fF
C15263 POR2X1_20/B POR2X1_397/CTRL2 0.01fF
C15264 POR2X1_835/Y POR2X1_836/Y 0.55fF
C15265 POR2X1_96/A PAND2X1_735/Y 0.02fF
C15266 PAND2X1_213/B VDD 0.04fF
C15267 POR2X1_376/B PAND2X1_658/B 0.44fF
C15268 PAND2X1_220/Y PAND2X1_794/B 0.03fF
C15269 PAND2X1_712/CTRL PAND2X1_707/Y 0.01fF
C15270 POR2X1_96/A POR2X1_329/CTRL 0.01fF
C15271 POR2X1_193/A VDD 0.48fF
C15272 PAND2X1_751/O POR2X1_546/A 0.01fF
C15273 POR2X1_579/Y VDD 1.36fF
C15274 POR2X1_110/Y PAND2X1_446/Y 0.03fF
C15275 POR2X1_48/O POR2X1_48/Y 0.01fF
C15276 POR2X1_461/B POR2X1_789/Y 0.02fF
C15277 POR2X1_192/Y POR2X1_776/B 0.03fF
C15278 POR2X1_602/B POR2X1_532/A 0.03fF
C15279 POR2X1_730/Y POR2X1_466/A 0.05fF
C15280 PAND2X1_65/B POR2X1_35/Y 3.80fF
C15281 POR2X1_490/Y PAND2X1_853/B 0.03fF
C15282 INPUT_1 D_INPUT_0 0.29fF
C15283 POR2X1_572/B VDD 0.16fF
C15284 POR2X1_489/CTRL POR2X1_68/B 0.01fF
C15285 POR2X1_517/Y POR2X1_13/A 0.01fF
C15286 POR2X1_336/CTRL2 POR2X1_814/B 0.03fF
C15287 PAND2X1_711/CTRL2 POR2X1_763/A 0.05fF
C15288 POR2X1_338/O PAND2X1_20/A 0.18fF
C15289 POR2X1_467/Y POR2X1_162/Y 0.05fF
C15290 PAND2X1_93/B POR2X1_186/B 0.03fF
C15291 POR2X1_52/A POR2X1_290/Y 0.04fF
C15292 POR2X1_66/A POR2X1_520/B 0.01fF
C15293 POR2X1_108/CTRL2 PAND2X1_562/B 0.03fF
C15294 POR2X1_41/B POR2X1_680/Y 1.71fF
C15295 POR2X1_545/A VDD -0.00fF
C15296 PAND2X1_90/A PAND2X1_92/CTRL 0.01fF
C15297 POR2X1_43/B VDD 4.65fF
C15298 POR2X1_48/A POR2X1_129/Y 0.02fF
C15299 POR2X1_383/A POR2X1_254/CTRL2 0.03fF
C15300 PAND2X1_602/Y PAND2X1_788/a_16_344# 0.02fF
C15301 POR2X1_789/A VDD 0.14fF
C15302 POR2X1_459/O POR2X1_459/A 0.01fF
C15303 POR2X1_863/O POR2X1_855/Y 0.01fF
C15304 D_INPUT_0 POR2X1_153/Y 0.13fF
C15305 PAND2X1_148/Y VDD 0.02fF
C15306 POR2X1_157/O INPUT_5 0.10fF
C15307 D_GATE_865 PAND2X1_32/B 0.01fF
C15308 PAND2X1_554/a_76_28# PAND2X1_348/Y 0.03fF
C15309 PAND2X1_211/O PAND2X1_352/Y 0.09fF
C15310 POR2X1_532/A POR2X1_213/B 1.02fF
C15311 POR2X1_614/A VDD 3.42fF
C15312 D_INPUT_3 POR2X1_611/O 0.02fF
C15313 POR2X1_317/Y VDD 0.05fF
C15314 PAND2X1_57/B POR2X1_391/Y 0.20fF
C15315 POR2X1_383/A PAND2X1_299/CTRL 0.04fF
C15316 POR2X1_23/Y PAND2X1_716/B 0.06fF
C15317 POR2X1_129/O POR2X1_129/Y 0.04fF
C15318 PAND2X1_242/CTRL POR2X1_7/B 0.01fF
C15319 POR2X1_52/A POR2X1_238/Y 0.06fF
C15320 PAND2X1_387/O PAND2X1_60/B 0.02fF
C15321 POR2X1_271/B PAND2X1_840/Y 0.03fF
C15322 PAND2X1_41/B POR2X1_218/CTRL2 0.00fF
C15323 POR2X1_225/CTRL2 POR2X1_129/Y 0.01fF
C15324 POR2X1_119/Y PAND2X1_477/O 0.17fF
C15325 POR2X1_406/Y PAND2X1_734/O 0.02fF
C15326 PAND2X1_182/A PAND2X1_566/Y 0.17fF
C15327 POR2X1_416/Y POR2X1_232/CTRL2 0.01fF
C15328 POR2X1_567/B POR2X1_564/O 0.59fF
C15329 POR2X1_579/Y POR2X1_741/Y 0.03fF
C15330 POR2X1_38/B VDD 1.80fF
C15331 POR2X1_578/Y D_GATE_741 0.01fF
C15332 PAND2X1_830/CTRL2 PAND2X1_562/B 0.05fF
C15333 PAND2X1_41/B POR2X1_738/A 0.09fF
C15334 PAND2X1_659/Y POR2X1_48/A 0.03fF
C15335 PAND2X1_845/CTRL PAND2X1_35/Y 0.01fF
C15336 POR2X1_57/A POR2X1_399/O 0.06fF
C15337 PAND2X1_435/Y POR2X1_153/Y 0.01fF
C15338 POR2X1_188/A PAND2X1_698/CTRL2 0.01fF
C15339 POR2X1_71/CTRL2 POR2X1_60/A 0.01fF
C15340 POR2X1_78/A POR2X1_209/CTRL 0.01fF
C15341 POR2X1_656/CTRL POR2X1_737/A 0.01fF
C15342 POR2X1_794/B POR2X1_675/Y 0.03fF
C15343 POR2X1_78/A POR2X1_186/B 0.74fF
C15344 PAND2X1_469/B PAND2X1_115/B 0.05fF
C15345 POR2X1_445/CTRL POR2X1_702/A 0.00fF
C15346 POR2X1_278/Y PAND2X1_347/O 0.15fF
C15347 POR2X1_147/A POR2X1_294/B 0.03fF
C15348 PAND2X1_563/B PAND2X1_854/A 0.25fF
C15349 POR2X1_123/A PAND2X1_65/B 4.95fF
C15350 POR2X1_439/O POR2X1_456/B 0.01fF
C15351 PAND2X1_477/B PAND2X1_241/CTRL2 0.00fF
C15352 PAND2X1_76/Y POR2X1_283/A 0.07fF
C15353 POR2X1_523/Y POR2X1_294/B 0.02fF
C15354 PAND2X1_250/a_16_344# POR2X1_249/Y 0.05fF
C15355 POR2X1_563/CTRL2 POR2X1_569/A 0.02fF
C15356 POR2X1_840/CTRL POR2X1_307/Y 0.01fF
C15357 PAND2X1_679/O POR2X1_687/A 0.01fF
C15358 POR2X1_61/Y POR2X1_259/O 0.08fF
C15359 PAND2X1_69/A POR2X1_208/CTRL 0.03fF
C15360 POR2X1_40/Y PAND2X1_124/m4_208_n4# 0.01fF
C15361 POR2X1_416/B POR2X1_628/Y 0.04fF
C15362 POR2X1_52/A POR2X1_526/O 0.02fF
C15363 POR2X1_68/A POR2X1_732/B 0.03fF
C15364 POR2X1_79/Y PAND2X1_739/B 0.10fF
C15365 POR2X1_219/CTRL2 POR2X1_294/B 0.03fF
C15366 POR2X1_193/A PAND2X1_32/B 0.07fF
C15367 POR2X1_287/B POR2X1_773/B 0.05fF
C15368 POR2X1_579/Y PAND2X1_32/B 1.79fF
C15369 PAND2X1_90/A PAND2X1_63/Y 0.10fF
C15370 POR2X1_750/A POR2X1_749/CTRL 0.02fF
C15371 POR2X1_649/CTRL2 POR2X1_294/B 0.16fF
C15372 POR2X1_366/Y PAND2X1_69/A 0.42fF
C15373 PAND2X1_69/A POR2X1_294/B 0.30fF
C15374 POR2X1_40/a_56_344# INPUT_7 0.00fF
C15375 POR2X1_78/B POR2X1_796/A 0.03fF
C15376 POR2X1_614/A POR2X1_741/Y 0.06fF
C15377 POR2X1_390/B POR2X1_335/CTRL2 0.00fF
C15378 POR2X1_41/B PAND2X1_388/Y 13.65fF
C15379 POR2X1_278/Y PAND2X1_349/A 0.02fF
C15380 POR2X1_440/Y VDD 0.33fF
C15381 INPUT_1 PAND2X1_90/Y 0.05fF
C15382 PAND2X1_228/CTRL PAND2X1_341/A 0.01fF
C15383 POR2X1_730/Y POR2X1_448/A 0.01fF
C15384 POR2X1_563/Y POR2X1_570/B 0.01fF
C15385 PAND2X1_831/Y PAND2X1_841/B 0.03fF
C15386 POR2X1_330/Y POR2X1_210/A 0.04fF
C15387 POR2X1_614/A PAND2X1_81/B 0.03fF
C15388 POR2X1_68/B PAND2X1_110/O 0.04fF
C15389 POR2X1_750/B POR2X1_553/O 0.02fF
C15390 PAND2X1_434/CTRL VDD 0.00fF
C15391 PAND2X1_784/O PAND2X1_778/Y 0.03fF
C15392 PAND2X1_95/B D_INPUT_6 0.05fF
C15393 PAND2X1_856/O PAND2X1_805/A 0.06fF
C15394 POR2X1_186/Y PAND2X1_746/O 0.04fF
C15395 GATE_479 POR2X1_394/A 0.03fF
C15396 PAND2X1_652/A PAND2X1_186/CTRL 0.02fF
C15397 POR2X1_763/Y PAND2X1_731/A 0.13fF
C15398 PAND2X1_715/CTRL POR2X1_310/Y 0.01fF
C15399 POR2X1_43/B PAND2X1_32/B 0.03fF
C15400 POR2X1_41/B PAND2X1_549/B 0.07fF
C15401 POR2X1_347/O POR2X1_296/B 0.16fF
C15402 PAND2X1_726/CTRL2 POR2X1_152/Y 0.01fF
C15403 POR2X1_334/a_16_28# POR2X1_814/B 0.02fF
C15404 POR2X1_383/A POR2X1_327/CTRL 0.01fF
C15405 POR2X1_311/Y PAND2X1_643/A 0.93fF
C15406 PAND2X1_490/CTRL PAND2X1_6/Y 0.01fF
C15407 PAND2X1_90/A POR2X1_113/Y 0.02fF
C15408 PAND2X1_23/Y POR2X1_318/A 0.08fF
C15409 POR2X1_16/A PAND2X1_571/Y 0.05fF
C15410 POR2X1_853/O POR2X1_854/B 0.31fF
C15411 POR2X1_72/B POR2X1_117/Y 0.00fF
C15412 POR2X1_37/Y POR2X1_39/B 2.20fF
C15413 POR2X1_114/B PAND2X1_96/B 0.03fF
C15414 POR2X1_307/Y POR2X1_725/Y 0.06fF
C15415 POR2X1_532/A POR2X1_805/A 0.07fF
C15416 POR2X1_477/A PAND2X1_60/B 0.03fF
C15417 POR2X1_32/A POR2X1_761/A 0.03fF
C15418 POR2X1_614/A PAND2X1_32/B 0.28fF
C15419 POR2X1_119/Y POR2X1_40/Y 0.18fF
C15420 PAND2X1_23/Y POR2X1_713/B 0.01fF
C15421 POR2X1_243/Y POR2X1_260/A 0.07fF
C15422 POR2X1_78/B PAND2X1_399/CTRL2 0.01fF
C15423 POR2X1_834/Y PAND2X1_57/B 1.46fF
C15424 POR2X1_81/A POR2X1_60/A 0.01fF
C15425 POR2X1_785/B POR2X1_776/B 0.16fF
C15426 POR2X1_100/CTRL2 PAND2X1_69/A 0.02fF
C15427 PAND2X1_649/A POR2X1_591/A 0.01fF
C15428 POR2X1_865/B POR2X1_778/B 0.03fF
C15429 PAND2X1_472/A POR2X1_395/Y 0.06fF
C15430 POR2X1_480/A PAND2X1_142/O 0.06fF
C15431 PAND2X1_79/Y D_INPUT_1 0.46fF
C15432 POR2X1_38/B PAND2X1_32/B 0.10fF
C15433 POR2X1_41/B POR2X1_41/CTRL 0.01fF
C15434 PAND2X1_96/B POR2X1_649/B 0.27fF
C15435 POR2X1_222/Y POR2X1_128/B 0.03fF
C15436 POR2X1_563/a_16_28# POR2X1_186/B 0.03fF
C15437 POR2X1_224/CTRL POR2X1_394/A 0.05fF
C15438 PAND2X1_170/CTRL VDD 0.00fF
C15439 POR2X1_394/A PAND2X1_719/O 0.01fF
C15440 POR2X1_614/A PAND2X1_312/O 0.01fF
C15441 POR2X1_94/A PAND2X1_379/CTRL2 0.01fF
C15442 POR2X1_68/A PAND2X1_306/a_76_28# 0.01fF
C15443 POR2X1_180/B POR2X1_732/B 0.03fF
C15444 POR2X1_383/A POR2X1_218/A 0.03fF
C15445 PAND2X1_546/Y PAND2X1_550/B 0.00fF
C15446 POR2X1_139/A POR2X1_137/Y 0.00fF
C15447 POR2X1_362/Y POR2X1_343/Y 0.10fF
C15448 POR2X1_65/A POR2X1_518/CTRL 0.01fF
C15449 PAND2X1_90/A POR2X1_260/A 0.07fF
C15450 VDD POR2X1_183/CTRL 0.00fF
C15451 PAND2X1_865/Y PAND2X1_363/Y 0.02fF
C15452 POR2X1_66/B POR2X1_632/Y 1.02fF
C15453 PAND2X1_824/B POR2X1_208/CTRL 0.09fF
C15454 PAND2X1_308/Y PAND2X1_303/CTRL2 0.01fF
C15455 POR2X1_702/O POR2X1_702/A 0.01fF
C15456 PAND2X1_82/O POR2X1_38/B -0.00fF
C15457 POR2X1_96/A PAND2X1_355/CTRL2 0.00fF
C15458 PAND2X1_511/CTRL PAND2X1_48/A 0.05fF
C15459 POR2X1_477/A POR2X1_353/A 0.03fF
C15460 PAND2X1_824/B POR2X1_294/B 0.14fF
C15461 PAND2X1_96/B POR2X1_222/A 0.03fF
C15462 POR2X1_61/A POR2X1_206/A 0.02fF
C15463 POR2X1_296/B POR2X1_717/B 0.03fF
C15464 POR2X1_294/B PAND2X1_528/m4_208_n4# 0.04fF
C15465 POR2X1_174/B PAND2X1_72/A 0.07fF
C15466 POR2X1_730/Y POR2X1_149/B 0.03fF
C15467 POR2X1_639/Y PAND2X1_764/O 0.02fF
C15468 POR2X1_30/CTRL POR2X1_260/A 0.00fF
C15469 PAND2X1_697/CTRL POR2X1_260/A 0.00fF
C15470 POR2X1_192/Y POR2X1_192/B 0.05fF
C15471 POR2X1_119/Y PAND2X1_659/B 0.62fF
C15472 PAND2X1_23/Y POR2X1_574/Y 0.03fF
C15473 POR2X1_614/A POR2X1_543/CTRL2 0.03fF
C15474 PAND2X1_41/B POR2X1_731/Y 0.04fF
C15475 POR2X1_614/A PAND2X1_253/O 0.01fF
C15476 PAND2X1_358/A PAND2X1_341/CTRL 0.01fF
C15477 POR2X1_495/O POR2X1_77/Y 0.01fF
C15478 PAND2X1_93/B PAND2X1_628/O 0.17fF
C15479 POR2X1_785/O POR2X1_192/B 0.16fF
C15480 POR2X1_66/B PAND2X1_52/B 1.90fF
C15481 POR2X1_3/A POR2X1_1/O 0.20fF
C15482 POR2X1_614/A POR2X1_673/Y 0.03fF
C15483 POR2X1_615/O POR2X1_39/B 0.02fF
C15484 POR2X1_562/CTRL2 POR2X1_339/Y 0.01fF
C15485 POR2X1_46/Y POR2X1_7/Y 0.03fF
C15486 POR2X1_712/CTRL2 POR2X1_707/Y 0.00fF
C15487 PAND2X1_35/a_16_344# POR2X1_394/A 0.04fF
C15488 POR2X1_188/A PAND2X1_52/B 0.10fF
C15489 POR2X1_673/Y POR2X1_38/B 0.10fF
C15490 POR2X1_651/Y POR2X1_608/Y 0.08fF
C15491 POR2X1_343/Y PAND2X1_65/Y 0.02fF
C15492 POR2X1_265/Y POR2X1_406/a_76_344# 0.01fF
C15493 POR2X1_48/Y PAND2X1_199/B 0.06fF
C15494 POR2X1_57/A PAND2X1_343/CTRL 0.01fF
C15495 PAND2X1_227/CTRL POR2X1_394/A 0.08fF
C15496 POR2X1_10/O POR2X1_38/Y 0.02fF
C15497 PAND2X1_659/Y POR2X1_413/A 0.03fF
C15498 PAND2X1_808/CTRL POR2X1_385/Y 0.50fF
C15499 POR2X1_447/B PAND2X1_55/Y 0.12fF
C15500 POR2X1_862/a_16_28# POR2X1_862/B 0.07fF
C15501 POR2X1_55/Y PAND2X1_506/Y 0.01fF
C15502 POR2X1_358/a_16_28# POR2X1_192/B 0.02fF
C15503 POR2X1_677/Y POR2X1_32/A 0.03fF
C15504 POR2X1_532/A POR2X1_520/B 0.05fF
C15505 PAND2X1_715/O POR2X1_39/B 0.01fF
C15506 POR2X1_96/A POR2X1_316/Y 0.02fF
C15507 POR2X1_96/A PAND2X1_798/Y 1.85fF
C15508 POR2X1_68/B POR2X1_559/A 0.14fF
C15509 POR2X1_502/A PAND2X1_109/O 0.17fF
C15510 POR2X1_394/A PAND2X1_509/O 0.09fF
C15511 PAND2X1_683/CTRL2 PAND2X1_69/A 0.01fF
C15512 POR2X1_9/Y POR2X1_32/A 1.68fF
C15513 PAND2X1_632/A PAND2X1_632/O 0.00fF
C15514 POR2X1_23/Y POR2X1_250/Y 0.10fF
C15515 POR2X1_342/Y PAND2X1_57/B 0.04fF
C15516 D_INPUT_3 PAND2X1_358/A 0.10fF
C15517 PAND2X1_612/B PAND2X1_612/a_56_28# 0.00fF
C15518 POR2X1_186/CTRL POR2X1_725/Y 0.02fF
C15519 PAND2X1_173/CTRL POR2X1_186/B 0.01fF
C15520 POR2X1_8/Y POR2X1_96/B 0.03fF
C15521 PAND2X1_308/Y PAND2X1_549/B 0.03fF
C15522 PAND2X1_99/B PAND2X1_97/Y 0.27fF
C15523 POR2X1_661/A POR2X1_330/Y 0.10fF
C15524 POR2X1_385/Y POR2X1_594/A 0.03fF
C15525 POR2X1_293/Y POR2X1_39/B 1.23fF
C15526 POR2X1_394/A PAND2X1_175/B 0.05fF
C15527 POR2X1_54/Y POR2X1_472/B -0.00fF
C15528 POR2X1_732/B POR2X1_181/O 0.04fF
C15529 POR2X1_765/Y PAND2X1_569/a_56_28# 0.00fF
C15530 PAND2X1_480/a_76_28# POR2X1_91/Y 0.02fF
C15531 POR2X1_567/A PAND2X1_69/A 4.45fF
C15532 PAND2X1_9/Y PAND2X1_35/A 0.02fF
C15533 POR2X1_544/A PAND2X1_72/A 0.03fF
C15534 POR2X1_732/B POR2X1_169/A 0.02fF
C15535 POR2X1_859/A PAND2X1_52/B 0.07fF
C15536 PAND2X1_653/CTRL PAND2X1_652/A 0.08fF
C15537 POR2X1_856/B POR2X1_453/Y 0.03fF
C15538 POR2X1_346/B POR2X1_260/A 0.03fF
C15539 POR2X1_416/B POR2X1_372/Y 0.03fF
C15540 POR2X1_124/B PAND2X1_122/CTRL 0.00fF
C15541 PAND2X1_641/Y POR2X1_83/O 0.04fF
C15542 POR2X1_38/B POR2X1_560/CTRL 0.00fF
C15543 POR2X1_383/A POR2X1_557/B 0.03fF
C15544 PAND2X1_96/B PAND2X1_122/CTRL2 0.03fF
C15545 POR2X1_542/B POR2X1_374/CTRL 0.01fF
C15546 POR2X1_78/B POR2X1_863/A 0.07fF
C15547 PAND2X1_838/B POR2X1_827/Y 0.04fF
C15548 POR2X1_416/B PAND2X1_709/CTRL 0.03fF
C15549 PAND2X1_271/O POR2X1_76/A 0.07fF
C15550 POR2X1_326/A POR2X1_725/Y 0.07fF
C15551 POR2X1_566/B POR2X1_566/O 0.20fF
C15552 POR2X1_858/B POR2X1_851/CTRL 0.01fF
C15553 POR2X1_83/B PAND2X1_206/B 0.07fF
C15554 POR2X1_675/Y POR2X1_741/B 0.01fF
C15555 POR2X1_713/CTRL2 POR2X1_711/Y 0.01fF
C15556 PAND2X1_724/CTRL PAND2X1_326/B 0.01fF
C15557 PAND2X1_728/a_16_344# PAND2X1_853/B 0.01fF
C15558 POR2X1_735/a_16_28# POR2X1_318/A 0.09fF
C15559 POR2X1_416/B POR2X1_519/Y 0.01fF
C15560 PAND2X1_221/O POR2X1_250/Y 0.07fF
C15561 POR2X1_796/A POR2X1_294/A 0.07fF
C15562 POR2X1_416/Y POR2X1_416/B 0.01fF
C15563 PAND2X1_39/B POR2X1_66/A 0.36fF
C15564 PAND2X1_32/CTRL POR2X1_94/A 0.02fF
C15565 PAND2X1_339/Y POR2X1_522/O 0.18fF
C15566 POR2X1_680/a_16_28# POR2X1_594/A 0.03fF
C15567 POR2X1_678/Y POR2X1_808/CTRL2 0.03fF
C15568 POR2X1_38/Y PAND2X1_198/CTRL 0.01fF
C15569 PAND2X1_221/Y PAND2X1_739/Y 0.33fF
C15570 POR2X1_648/A POR2X1_718/A 0.01fF
C15571 POR2X1_416/B POR2X1_29/Y 0.51fF
C15572 PAND2X1_51/CTRL PAND2X1_3/B 0.01fF
C15573 POR2X1_52/CTRL2 POR2X1_7/A 0.01fF
C15574 POR2X1_34/A PAND2X1_39/B 0.04fF
C15575 POR2X1_768/CTRL2 POR2X1_113/B 0.01fF
C15576 POR2X1_309/a_16_28# POR2X1_150/Y 0.02fF
C15577 POR2X1_490/Y POR2X1_23/Y 0.17fF
C15578 POR2X1_814/A POR2X1_61/Y 0.07fF
C15579 POR2X1_54/Y PAND2X1_381/Y 0.05fF
C15580 POR2X1_316/Y POR2X1_7/A 0.07fF
C15581 PAND2X1_166/CTRL POR2X1_854/B 0.33fF
C15582 PAND2X1_399/CTRL2 POR2X1_294/A 0.00fF
C15583 POR2X1_250/Y PAND2X1_740/O 0.03fF
C15584 PAND2X1_508/O PAND2X1_506/Y 0.00fF
C15585 POR2X1_65/Y POR2X1_83/B 0.03fF
C15586 POR2X1_408/Y POR2X1_39/B 0.01fF
C15587 POR2X1_568/B POR2X1_854/B 0.01fF
C15588 PAND2X1_388/Y POR2X1_77/Y 0.06fF
C15589 PAND2X1_22/CTRL2 PAND2X1_11/Y 0.01fF
C15590 POR2X1_567/A PAND2X1_824/B 0.10fF
C15591 PAND2X1_469/a_16_344# POR2X1_32/A 0.01fF
C15592 POR2X1_711/Y POR2X1_713/B 0.01fF
C15593 POR2X1_244/Y POR2X1_4/Y 0.03fF
C15594 POR2X1_804/A PAND2X1_135/CTRL 0.12fF
C15595 POR2X1_528/Y POR2X1_305/CTRL 0.04fF
C15596 PAND2X1_696/m4_208_n4# POR2X1_648/Y 0.08fF
C15597 POR2X1_48/A POR2X1_37/Y 0.55fF
C15598 PAND2X1_549/B POR2X1_77/Y 0.03fF
C15599 POR2X1_260/B POR2X1_267/CTRL2 0.01fF
C15600 PAND2X1_406/CTRL POR2X1_121/B 0.01fF
C15601 PAND2X1_18/B PAND2X1_3/B 0.13fF
C15602 POR2X1_353/Y POR2X1_443/CTRL 0.01fF
C15603 POR2X1_129/O POR2X1_37/Y 0.01fF
C15604 POR2X1_841/B POR2X1_806/CTRL2 0.01fF
C15605 POR2X1_537/Y POR2X1_851/a_16_28# 0.01fF
C15606 POR2X1_161/O POR2X1_162/Y 0.01fF
C15607 POR2X1_677/Y POR2X1_184/Y 0.02fF
C15608 PAND2X1_633/O POR2X1_826/Y 0.01fF
C15609 POR2X1_35/B PAND2X1_24/O 0.01fF
C15610 POR2X1_60/A PAND2X1_207/O 0.03fF
C15611 PAND2X1_63/a_16_344# POR2X1_296/B 0.01fF
C15612 POR2X1_96/Y POR2X1_62/Y 0.03fF
C15613 POR2X1_805/Y POR2X1_66/A 0.01fF
C15614 PAND2X1_510/B POR2X1_80/a_76_344# 0.00fF
C15615 PAND2X1_472/O POR2X1_77/Y 0.15fF
C15616 PAND2X1_651/Y POR2X1_677/Y 0.05fF
C15617 PAND2X1_20/A POR2X1_66/A 0.92fF
C15618 PAND2X1_313/CTRL2 PAND2X1_72/A 0.00fF
C15619 POR2X1_814/A POR2X1_193/CTRL 0.05fF
C15620 PAND2X1_2/CTRL2 D_INPUT_4 0.01fF
C15621 PAND2X1_20/A POR2X1_34/A 0.03fF
C15622 PAND2X1_384/a_76_28# POR2X1_383/Y 0.04fF
C15623 PAND2X1_340/B POR2X1_381/O 0.01fF
C15624 POR2X1_814/A POR2X1_35/Y 0.07fF
C15625 POR2X1_760/A PAND2X1_218/CTRL2 0.02fF
C15626 POR2X1_566/A POR2X1_663/B 0.03fF
C15627 POR2X1_471/A POR2X1_724/CTRL 0.00fF
C15628 PAND2X1_557/A POR2X1_487/O 0.02fF
C15629 POR2X1_48/A POR2X1_615/O 0.01fF
C15630 POR2X1_856/B PAND2X1_52/Y 0.15fF
C15631 POR2X1_456/B PAND2X1_125/CTRL2 0.01fF
C15632 POR2X1_804/a_16_28# POR2X1_330/Y 0.09fF
C15633 POR2X1_814/B POR2X1_66/A 9.59fF
C15634 POR2X1_257/A POR2X1_46/Y 0.17fF
C15635 POR2X1_68/A PAND2X1_441/a_76_28# 0.02fF
C15636 POR2X1_60/A POR2X1_432/a_16_28# 0.01fF
C15637 PAND2X1_473/CTRL POR2X1_329/A 0.01fF
C15638 POR2X1_263/Y POR2X1_5/Y 0.02fF
C15639 POR2X1_438/Y PAND2X1_544/O 0.07fF
C15640 PAND2X1_404/Y PAND2X1_573/O 0.04fF
C15641 POR2X1_335/B POR2X1_814/A 0.04fF
C15642 POR2X1_220/B POR2X1_213/B 0.03fF
C15643 GATE_479 POR2X1_669/B 0.07fF
C15644 PAND2X1_796/CTRL PAND2X1_783/Y 0.01fF
C15645 POR2X1_667/A POR2X1_72/B 2.00fF
C15646 POR2X1_260/B POR2X1_220/Y 0.06fF
C15647 POR2X1_693/Y POR2X1_20/B 0.03fF
C15648 POR2X1_20/B PAND2X1_398/O 0.03fF
C15649 PAND2X1_790/O POR2X1_7/B 0.02fF
C15650 POR2X1_32/A PAND2X1_736/CTRL2 0.03fF
C15651 PAND2X1_473/Y PAND2X1_571/A 0.00fF
C15652 PAND2X1_73/Y POR2X1_285/CTRL2 0.04fF
C15653 POR2X1_83/B PAND2X1_220/Y -0.00fF
C15654 POR2X1_43/B PAND2X1_9/Y 0.02fF
C15655 POR2X1_848/A POR2X1_790/CTRL2 0.04fF
C15656 POR2X1_68/A POR2X1_831/CTRL 0.01fF
C15657 PAND2X1_48/B PAND2X1_487/CTRL 0.01fF
C15658 PAND2X1_23/Y PAND2X1_487/CTRL2 0.05fF
C15659 POR2X1_474/CTRL POR2X1_860/A 0.01fF
C15660 PAND2X1_464/m4_208_n4# PAND2X1_241/m4_208_n4# 0.13fF
C15661 POR2X1_446/B POR2X1_740/Y 0.03fF
C15662 POR2X1_260/B POR2X1_404/Y 0.03fF
C15663 POR2X1_20/B POR2X1_299/CTRL2 0.02fF
C15664 POR2X1_123/A POR2X1_814/A 0.03fF
C15665 POR2X1_78/B POR2X1_269/A 0.00fF
C15666 POR2X1_262/Y POR2X1_73/Y 9.61fF
C15667 POR2X1_750/B POR2X1_752/Y 0.03fF
C15668 PAND2X1_37/CTRL PAND2X1_8/Y 0.02fF
C15669 POR2X1_66/A PAND2X1_176/CTRL2 0.00fF
C15670 PAND2X1_243/B POR2X1_23/Y 0.00fF
C15671 POR2X1_78/B POR2X1_602/A 0.03fF
C15672 POR2X1_590/A VDD 3.62fF
C15673 POR2X1_554/B PAND2X1_60/B 0.03fF
C15674 POR2X1_66/A POR2X1_513/B 0.03fF
C15675 POR2X1_341/A POR2X1_341/a_16_28# 0.01fF
C15676 POR2X1_48/A POR2X1_293/Y 0.30fF
C15677 PAND2X1_217/B POR2X1_272/a_16_28# 0.01fF
C15678 POR2X1_649/B POR2X1_649/a_76_344# 0.01fF
C15679 POR2X1_23/Y PAND2X1_775/a_16_344# 0.03fF
C15680 POR2X1_278/Y POR2X1_32/A 0.05fF
C15681 PAND2X1_9/Y POR2X1_38/B 0.03fF
C15682 POR2X1_677/O PAND2X1_390/Y 0.00fF
C15683 PAND2X1_362/B POR2X1_594/CTRL 0.01fF
C15684 PAND2X1_793/Y POR2X1_487/CTRL 0.03fF
C15685 POR2X1_800/A POR2X1_808/a_16_28# 0.03fF
C15686 POR2X1_356/A POR2X1_434/A 0.01fF
C15687 POR2X1_174/B POR2X1_244/B 0.01fF
C15688 POR2X1_56/CTRL PAND2X1_254/Y 0.01fF
C15689 PAND2X1_39/B POR2X1_532/A 0.12fF
C15690 PAND2X1_63/Y POR2X1_84/B 0.01fF
C15691 POR2X1_829/A POR2X1_32/A 0.03fF
C15692 POR2X1_411/B POR2X1_387/Y 0.09fF
C15693 POR2X1_413/A POR2X1_37/Y 0.00fF
C15694 POR2X1_225/CTRL2 POR2X1_293/Y 0.01fF
C15695 POR2X1_856/B D_GATE_662 0.10fF
C15696 D_INPUT_3 POR2X1_612/O 0.01fF
C15697 POR2X1_648/Y POR2X1_407/a_16_28# 0.03fF
C15698 POR2X1_68/A POR2X1_855/CTRL2 0.03fF
C15699 PAND2X1_271/a_76_28# POR2X1_804/A 0.02fF
C15700 POR2X1_818/Y POR2X1_789/A 0.03fF
C15701 PAND2X1_623/O POR2X1_615/Y 0.01fF
C15702 POR2X1_72/B POR2X1_372/O 0.02fF
C15703 POR2X1_50/O INPUT_7 0.03fF
C15704 POR2X1_366/CTRL2 POR2X1_116/A 0.00fF
C15705 POR2X1_68/A PAND2X1_94/O 0.12fF
C15706 POR2X1_805/Y POR2X1_792/B 0.01fF
C15707 PAND2X1_676/a_76_28# POR2X1_257/A 0.02fF
C15708 POR2X1_9/Y POR2X1_294/A 0.01fF
C15709 POR2X1_368/O POR2X1_417/Y 0.02fF
C15710 POR2X1_68/A POR2X1_466/A 0.05fF
C15711 POR2X1_96/A PAND2X1_784/A 0.03fF
C15712 POR2X1_329/A PAND2X1_853/B 0.03fF
C15713 POR2X1_609/O POR2X1_609/A 0.01fF
C15714 POR2X1_78/B POR2X1_456/CTRL 0.00fF
C15715 POR2X1_411/B PAND2X1_121/O 0.03fF
C15716 PAND2X1_90/A POR2X1_243/A 0.02fF
C15717 POR2X1_542/B PAND2X1_93/B 0.03fF
C15718 POR2X1_54/Y POR2X1_7/A 0.15fF
C15719 POR2X1_128/CTRL2 POR2X1_750/B 0.14fF
C15720 PAND2X1_474/A VDD 0.10fF
C15721 PAND2X1_600/O PAND2X1_32/B 0.10fF
C15722 POR2X1_811/A POR2X1_796/O 0.00fF
C15723 POR2X1_13/A POR2X1_423/Y 0.10fF
C15724 INPUT_1 PAND2X1_33/O 0.01fF
C15725 POR2X1_590/A POR2X1_741/Y 0.06fF
C15726 POR2X1_75/a_16_28# POR2X1_23/Y 0.09fF
C15727 PAND2X1_242/Y POR2X1_39/B 0.05fF
C15728 POR2X1_48/A PAND2X1_553/CTRL 0.01fF
C15729 PAND2X1_118/O PAND2X1_73/Y 0.04fF
C15730 POR2X1_502/A PAND2X1_41/B 3.50fF
C15731 PAND2X1_420/O POR2X1_294/B 0.05fF
C15732 POR2X1_65/A POR2X1_682/Y 0.00fF
C15733 POR2X1_222/CTRL POR2X1_222/A 0.08fF
C15734 POR2X1_668/O VDD 0.00fF
C15735 PAND2X1_217/B POR2X1_275/CTRL2 0.32fF
C15736 PAND2X1_643/CTRL POR2X1_102/Y 0.01fF
C15737 POR2X1_49/Y POR2X1_46/Y 0.10fF
C15738 POR2X1_829/A POR2X1_829/a_16_28# 0.03fF
C15739 POR2X1_697/O POR2X1_236/Y 0.19fF
C15740 PAND2X1_20/A POR2X1_222/Y 0.02fF
C15741 POR2X1_646/B PAND2X1_48/A 0.00fF
C15742 POR2X1_709/a_56_344# POR2X1_709/A 0.00fF
C15743 POR2X1_83/B PAND2X1_370/CTRL2 0.03fF
C15744 PAND2X1_640/B POR2X1_278/A 0.09fF
C15745 POR2X1_65/A PAND2X1_793/Y 0.03fF
C15746 PAND2X1_496/CTRL POR2X1_777/B 0.29fF
C15747 PAND2X1_99/B PAND2X1_99/Y 0.11fF
C15748 PAND2X1_629/O POR2X1_627/Y 0.00fF
C15749 POR2X1_782/A POR2X1_782/a_16_28# 0.04fF
C15750 POR2X1_78/B POR2X1_403/B 0.60fF
C15751 PAND2X1_573/B POR2X1_56/Y 0.03fF
C15752 POR2X1_590/A PAND2X1_32/B 9.30fF
C15753 POR2X1_48/A POR2X1_408/Y 0.06fF
C15754 POR2X1_614/A POR2X1_267/A 0.02fF
C15755 POR2X1_88/Y POR2X1_236/Y 0.05fF
C15756 PAND2X1_857/A POR2X1_23/Y 0.05fF
C15757 POR2X1_498/Y POR2X1_73/Y 0.05fF
C15758 PAND2X1_564/B PAND2X1_569/A 0.01fF
C15759 POR2X1_542/B POR2X1_78/A 1.66fF
C15760 POR2X1_254/CTRL POR2X1_222/Y 0.01fF
C15761 POR2X1_448/CTRL2 POR2X1_788/B 0.03fF
C15762 PAND2X1_859/A POR2X1_382/CTRL2 0.01fF
C15763 POR2X1_283/Y PAND2X1_365/B 0.10fF
C15764 POR2X1_89/Y POR2X1_91/Y 0.06fF
C15765 POR2X1_78/A PAND2X1_79/Y 0.01fF
C15766 POR2X1_368/CTRL POR2X1_13/A 0.01fF
C15767 POR2X1_805/Y POR2X1_532/A 0.03fF
C15768 PAND2X1_215/B POR2X1_5/Y 0.02fF
C15769 POR2X1_37/Y PAND2X1_840/O 0.04fF
C15770 POR2X1_267/A POR2X1_38/B 0.02fF
C15771 POR2X1_263/Y POR2X1_235/a_56_344# 0.00fF
C15772 PAND2X1_96/B POR2X1_675/CTRL2 0.01fF
C15773 POR2X1_669/B POR2X1_142/Y 0.03fF
C15774 POR2X1_564/Y VDD 0.52fF
C15775 PAND2X1_48/B POR2X1_362/B 0.07fF
C15776 PAND2X1_90/A PAND2X1_667/CTRL2 0.12fF
C15777 PAND2X1_76/Y POR2X1_55/Y 0.03fF
C15778 PAND2X1_20/A POR2X1_532/A 0.10fF
C15779 POR2X1_649/CTRL2 POR2X1_643/A 0.05fF
C15780 POR2X1_614/A POR2X1_808/A 0.07fF
C15781 POR2X1_260/B POR2X1_332/CTRL 0.01fF
C15782 POR2X1_180/B POR2X1_466/A 0.05fF
C15783 POR2X1_641/CTRL2 POR2X1_318/A 0.03fF
C15784 POR2X1_278/Y PAND2X1_35/Y 0.03fF
C15785 POR2X1_857/B VDD 0.37fF
C15786 POR2X1_840/B PAND2X1_74/a_16_344# 0.03fF
C15787 POR2X1_15/CTRL POR2X1_69/A 0.01fF
C15788 POR2X1_483/CTRL2 POR2X1_193/A 0.02fF
C15789 POR2X1_814/B PAND2X1_411/a_56_28# 0.00fF
C15790 POR2X1_16/A PAND2X1_571/CTRL 0.27fF
C15791 POR2X1_37/Y PAND2X1_559/m4_208_n4# 0.04fF
C15792 PAND2X1_798/Y POR2X1_760/A 0.03fF
C15793 POR2X1_214/B VDD 0.00fF
C15794 POR2X1_433/CTRL PAND2X1_349/A 0.01fF
C15795 POR2X1_406/Y PAND2X1_197/Y 0.03fF
C15796 PAND2X1_6/A POR2X1_5/Y 0.21fF
C15797 PAND2X1_58/A PAND2X1_306/a_76_28# 0.01fF
C15798 POR2X1_294/B POR2X1_510/a_16_28# 0.02fF
C15799 PAND2X1_23/Y PAND2X1_131/O 0.11fF
C15800 PAND2X1_553/B POR2X1_46/Y 0.05fF
C15801 POR2X1_807/A PAND2X1_69/A 0.03fF
C15802 POR2X1_302/O POR2X1_114/B 0.01fF
C15803 POR2X1_41/B POR2X1_615/Y 0.00fF
C15804 POR2X1_455/CTRL2 POR2X1_702/A 0.00fF
C15805 PAND2X1_55/Y POR2X1_220/Y 0.06fF
C15806 POR2X1_294/B POR2X1_121/Y 0.03fF
C15807 POR2X1_814/B POR2X1_532/A 0.17fF
C15808 PAND2X1_231/O POR2X1_38/Y 0.01fF
C15809 PAND2X1_685/CTRL2 POR2X1_829/A 0.00fF
C15810 PAND2X1_253/a_16_344# POR2X1_186/B 0.00fF
C15811 PAND2X1_55/Y POR2X1_207/a_16_28# 0.02fF
C15812 POR2X1_437/Y PAND2X1_580/B 0.00fF
C15813 POR2X1_96/A POR2X1_13/Y 2.29fF
C15814 POR2X1_549/O POR2X1_68/B 0.01fF
C15815 PAND2X1_787/A PAND2X1_211/A 0.02fF
C15816 POR2X1_409/B POR2X1_394/A 0.10fF
C15817 POR2X1_673/Y POR2X1_590/A 0.03fF
C15818 POR2X1_38/B POR2X1_236/CTRL2 0.03fF
C15819 POR2X1_61/CTRL2 PAND2X1_58/A 0.01fF
C15820 POR2X1_46/Y PAND2X1_188/O 0.28fF
C15821 PAND2X1_865/O POR2X1_516/Y 0.04fF
C15822 PAND2X1_96/B POR2X1_741/a_16_28# 0.01fF
C15823 POR2X1_72/B POR2X1_245/Y 0.03fF
C15824 PAND2X1_662/CTRL VDD -0.00fF
C15825 PAND2X1_56/Y POR2X1_76/Y 0.32fF
C15826 PAND2X1_742/a_16_344# POR2X1_283/A 0.01fF
C15827 POR2X1_66/A POR2X1_703/CTRL2 0.10fF
C15828 POR2X1_502/A PAND2X1_411/CTRL 0.02fF
C15829 POR2X1_287/a_16_28# POR2X1_249/Y 0.01fF
C15830 POR2X1_750/B PAND2X1_158/O 0.02fF
C15831 POR2X1_275/A POR2X1_39/B 0.01fF
C15832 PAND2X1_617/O PAND2X1_52/B 0.18fF
C15833 PAND2X1_752/Y VDD 0.30fF
C15834 POR2X1_614/A POR2X1_483/CTRL2 0.05fF
C15835 POR2X1_481/A POR2X1_90/Y 0.03fF
C15836 PAND2X1_793/Y PAND2X1_190/Y 0.05fF
C15837 POR2X1_159/a_16_28# POR2X1_408/Y 0.03fF
C15838 POR2X1_78/B POR2X1_341/m4_208_n4# 0.03fF
C15839 POR2X1_532/A POR2X1_325/A 0.03fF
C15840 POR2X1_376/B POR2X1_387/Y 0.10fF
C15841 POR2X1_393/Y POR2X1_394/CTRL2 0.01fF
C15842 POR2X1_416/B POR2X1_485/Y 0.06fF
C15843 PAND2X1_90/A PAND2X1_110/O 0.01fF
C15844 POR2X1_16/A PAND2X1_718/Y 0.05fF
C15845 POR2X1_62/Y POR2X1_37/Y 0.06fF
C15846 POR2X1_581/O INPUT_5 0.01fF
C15847 PAND2X1_4/CTRL2 INPUT_0 0.00fF
C15848 POR2X1_416/B POR2X1_292/Y 0.06fF
C15849 PAND2X1_357/Y POR2X1_7/B 0.03fF
C15850 POR2X1_335/Y PAND2X1_57/B 0.01fF
C15851 POR2X1_523/Y POR2X1_546/B 0.26fF
C15852 POR2X1_83/B PAND2X1_560/B 0.01fF
C15853 POR2X1_55/Y PAND2X1_349/a_76_28# 0.01fF
C15854 POR2X1_564/Y PAND2X1_32/B 2.98fF
C15855 PAND2X1_56/Y POR2X1_740/Y 0.05fF
C15856 PAND2X1_294/O POR2X1_39/B 0.01fF
C15857 POR2X1_121/B POR2X1_774/A 3.01fF
C15858 POR2X1_38/Y PAND2X1_735/Y 0.07fF
C15859 POR2X1_327/Y POR2X1_850/B 0.03fF
C15860 POR2X1_278/Y PAND2X1_844/B 0.02fF
C15861 INPUT_0 POR2X1_172/Y 0.17fF
C15862 PAND2X1_96/B POR2X1_405/Y 0.01fF
C15863 PAND2X1_319/B POR2X1_13/A 0.04fF
C15864 POR2X1_72/B PAND2X1_579/A 0.12fF
C15865 POR2X1_480/A POR2X1_725/Y 0.07fF
C15866 PAND2X1_96/B POR2X1_784/A 0.03fF
C15867 POR2X1_67/CTRL POR2X1_39/B 0.06fF
C15868 POR2X1_57/A PAND2X1_137/Y 0.15fF
C15869 POR2X1_339/O POR2X1_186/Y 0.06fF
C15870 POR2X1_383/A POR2X1_770/A 0.01fF
C15871 POR2X1_532/A POR2X1_513/B 0.03fF
C15872 PAND2X1_365/a_76_28# POR2X1_7/B 0.01fF
C15873 POR2X1_96/A PAND2X1_787/A 0.03fF
C15874 PAND2X1_481/CTRL POR2X1_355/A 0.01fF
C15875 POR2X1_254/Y POR2X1_510/Y 0.07fF
C15876 POR2X1_554/Y POR2X1_573/A 0.02fF
C15877 POR2X1_68/A POR2X1_149/B 0.10fF
C15878 PAND2X1_698/O PAND2X1_65/B 0.23fF
C15879 PAND2X1_65/B POR2X1_463/Y 0.03fF
C15880 PAND2X1_149/O PAND2X1_149/A -0.00fF
C15881 POR2X1_42/Y POR2X1_748/O 0.11fF
C15882 INPUT_1 POR2X1_621/B 0.01fF
C15883 PAND2X1_721/B POR2X1_397/O 0.02fF
C15884 POR2X1_38/Y PAND2X1_493/Y 0.09fF
C15885 PAND2X1_671/Y POR2X1_260/A 0.00fF
C15886 POR2X1_466/A POR2X1_181/O 0.04fF
C15887 POR2X1_537/Y POR2X1_830/CTRL2 0.01fF
C15888 PAND2X1_480/B POR2X1_283/A 0.10fF
C15889 PAND2X1_96/B POR2X1_732/B 0.05fF
C15890 POR2X1_336/O POR2X1_740/Y 0.51fF
C15891 POR2X1_417/Y PAND2X1_357/O 0.03fF
C15892 PAND2X1_94/A POR2X1_461/B 0.02fF
C15893 POR2X1_779/A POR2X1_712/A 0.22fF
C15894 PAND2X1_90/Y POR2X1_758/Y 0.07fF
C15895 POR2X1_466/A POR2X1_169/A 0.05fF
C15896 PAND2X1_114/Y PAND2X1_388/Y 0.03fF
C15897 POR2X1_330/Y POR2X1_737/A 0.05fF
C15898 PAND2X1_231/O POR2X1_153/Y 0.19fF
C15899 POR2X1_68/A POR2X1_219/CTRL 0.01fF
C15900 PAND2X1_472/A PAND2X1_401/a_56_28# 0.00fF
C15901 POR2X1_277/O POR2X1_278/A 0.00fF
C15902 POR2X1_754/A POR2X1_283/A 0.10fF
C15903 PAND2X1_140/A POR2X1_7/B 0.06fF
C15904 PAND2X1_57/B PAND2X1_757/a_76_28# 0.02fF
C15905 POR2X1_68/A POR2X1_644/A 0.04fF
C15906 POR2X1_407/A PAND2X1_69/A 0.32fF
C15907 PAND2X1_714/Y VDD 0.04fF
C15908 POR2X1_567/A PAND2X1_420/O 0.25fF
C15909 PAND2X1_738/A POR2X1_763/Y 0.14fF
C15910 POR2X1_617/Y POR2X1_750/B 0.03fF
C15911 POR2X1_16/A PAND2X1_580/B 0.03fF
C15912 POR2X1_528/Y POR2X1_7/B 0.13fF
C15913 PAND2X1_56/Y POR2X1_336/a_56_344# 0.03fF
C15914 POR2X1_390/B PAND2X1_57/B 0.03fF
C15915 POR2X1_114/CTRL POR2X1_68/B 0.01fF
C15916 POR2X1_826/Y POR2X1_825/Y 0.00fF
C15917 PAND2X1_58/CTRL POR2X1_507/A 0.03fF
C15918 PAND2X1_61/O POR2X1_39/B 0.11fF
C15919 POR2X1_502/A POR2X1_502/CTRL 0.03fF
C15920 PAND2X1_73/Y POR2X1_568/B 0.08fF
C15921 POR2X1_39/Y VDD 0.03fF
C15922 POR2X1_41/B PAND2X1_264/O 0.05fF
C15923 POR2X1_272/Y POR2X1_394/A 0.03fF
C15924 PAND2X1_583/O PAND2X1_32/B 0.00fF
C15925 POR2X1_383/A POR2X1_740/Y 0.23fF
C15926 PAND2X1_50/CTRL2 PAND2X1_18/B 0.05fF
C15927 POR2X1_137/Y POR2X1_391/Y 0.02fF
C15928 POR2X1_56/Y POR2X1_91/Y 0.07fF
C15929 PAND2X1_641/Y PAND2X1_734/B 0.03fF
C15930 PAND2X1_88/Y POR2X1_631/B 0.03fF
C15931 PAND2X1_650/A POR2X1_293/Y 0.03fF
C15932 PAND2X1_865/Y PAND2X1_217/B 0.05fF
C15933 PAND2X1_859/A POR2X1_4/Y 0.03fF
C15934 POR2X1_190/Y POR2X1_353/A 0.46fF
C15935 POR2X1_205/Y POR2X1_215/A 0.01fF
C15936 POR2X1_563/Y POR2X1_569/A 0.19fF
C15937 PAND2X1_665/m4_208_n4# PAND2X1_666/m4_208_n4# 0.13fF
C15938 PAND2X1_55/Y POR2X1_215/A 0.00fF
C15939 POR2X1_40/Y PAND2X1_326/B 0.05fF
C15940 PAND2X1_6/Y POR2X1_832/A 0.05fF
C15941 POR2X1_60/A POR2X1_39/B 2.87fF
C15942 POR2X1_96/O POR2X1_7/B 0.01fF
C15943 POR2X1_557/B INPUT_0 0.07fF
C15944 VDD POR2X1_314/Y 0.13fF
C15945 POR2X1_119/Y POR2X1_5/Y 0.15fF
C15946 PAND2X1_686/O POR2X1_7/B 0.01fF
C15947 PAND2X1_672/CTRL VDD -0.00fF
C15948 PAND2X1_60/B POR2X1_702/A 0.06fF
C15949 PAND2X1_71/CTRL POR2X1_244/Y 0.00fF
C15950 POR2X1_270/O POR2X1_724/A 0.05fF
C15951 PAND2X1_575/B POR2X1_184/a_16_28# 0.02fF
C15952 POR2X1_804/A POR2X1_366/A 0.10fF
C15953 POR2X1_391/O POR2X1_816/A 0.01fF
C15954 POR2X1_264/Y POR2X1_773/B 0.06fF
C15955 POR2X1_403/B POR2X1_294/A 0.60fF
C15956 PAND2X1_659/Y POR2X1_393/CTRL2 0.01fF
C15957 POR2X1_708/CTRL POR2X1_294/A 0.00fF
C15958 POR2X1_356/A POR2X1_544/B 0.03fF
C15959 PAND2X1_199/A PAND2X1_199/a_16_344# 0.02fF
C15960 POR2X1_48/A PAND2X1_242/Y 0.05fF
C15961 PAND2X1_728/CTRL POR2X1_816/A 0.01fF
C15962 PAND2X1_832/O POR2X1_316/Y 0.05fF
C15963 POR2X1_614/A POR2X1_687/A 1.39fF
C15964 POR2X1_814/A POR2X1_859/O 0.07fF
C15965 PAND2X1_90/A POR2X1_559/A 0.07fF
C15966 POR2X1_701/a_76_344# POR2X1_236/Y 0.01fF
C15967 POR2X1_16/A POR2X1_315/CTRL 0.01fF
C15968 PAND2X1_645/B POR2X1_757/a_16_28# 0.01fF
C15969 POR2X1_333/A POR2X1_161/CTRL 0.02fF
C15970 PAND2X1_367/O VDD 0.00fF
C15971 PAND2X1_865/Y VDD 0.36fF
C15972 PAND2X1_480/O POR2X1_238/Y 0.04fF
C15973 PAND2X1_675/A PAND2X1_348/A 0.07fF
C15974 POR2X1_316/a_76_344# POR2X1_293/Y 0.01fF
C15975 POR2X1_329/A PAND2X1_796/B 0.02fF
C15976 POR2X1_62/Y POR2X1_293/Y 0.10fF
C15977 POR2X1_51/O VDD 0.00fF
C15978 PAND2X1_469/B PAND2X1_348/A 0.10fF
C15979 PAND2X1_71/O PAND2X1_48/A 0.02fF
C15980 POR2X1_59/CTRL POR2X1_90/Y 0.00fF
C15981 PAND2X1_454/B POR2X1_329/A 0.03fF
C15982 POR2X1_24/a_16_28# POR2X1_77/Y 0.03fF
C15983 PAND2X1_119/a_16_344# PAND2X1_94/A 0.02fF
C15984 PAND2X1_65/B POR2X1_736/A 0.05fF
C15985 PAND2X1_206/A PAND2X1_206/B 0.39fF
C15986 POR2X1_702/A POR2X1_332/O 0.14fF
C15987 PAND2X1_862/B POR2X1_184/CTRL2 0.02fF
C15988 PAND2X1_727/CTRL POR2X1_91/Y 0.01fF
C15989 POR2X1_502/A PAND2X1_665/O 0.12fF
C15990 POR2X1_822/CTRL2 POR2X1_77/Y 0.00fF
C15991 PAND2X1_799/CTRL2 PAND2X1_539/Y 0.01fF
C15992 POR2X1_43/B PAND2X1_851/CTRL2 0.00fF
C15993 POR2X1_260/B POR2X1_67/Y 0.00fF
C15994 POR2X1_107/O POR2X1_77/Y 0.12fF
C15995 POR2X1_383/A PAND2X1_253/CTRL 0.03fF
C15996 PAND2X1_661/Y PAND2X1_194/a_76_28# 0.01fF
C15997 PAND2X1_744/CTRL POR2X1_294/A -0.00fF
C15998 POR2X1_112/CTRL2 POR2X1_775/A 0.01fF
C15999 D_INPUT_1 PAND2X1_527/CTRL2 0.01fF
C16000 D_GATE_662 POR2X1_191/Y 0.07fF
C16001 PAND2X1_365/B PAND2X1_365/A 0.02fF
C16002 POR2X1_23/Y POR2X1_329/A 0.13fF
C16003 POR2X1_57/A PAND2X1_853/B 0.06fF
C16004 POR2X1_162/Y POR2X1_156/Y 0.01fF
C16005 PAND2X1_337/A PAND2X1_336/Y 0.00fF
C16006 POR2X1_416/B POR2X1_295/Y 0.21fF
C16007 POR2X1_566/B POR2X1_192/O 0.25fF
C16008 PAND2X1_631/A PAND2X1_469/B 0.44fF
C16009 POR2X1_673/Y POR2X1_623/A 0.03fF
C16010 POR2X1_112/CTRL2 POR2X1_112/Y 0.00fF
C16011 POR2X1_635/a_16_28# POR2X1_635/A 0.03fF
C16012 POR2X1_116/A POR2X1_274/A 0.03fF
C16013 PAND2X1_48/B D_INPUT_4 0.03fF
C16014 POR2X1_714/a_16_28# POR2X1_704/Y 0.09fF
C16015 POR2X1_471/A POR2X1_454/O 0.08fF
C16016 POR2X1_176/a_16_28# POR2X1_90/Y 0.07fF
C16017 POR2X1_707/B D_INPUT_7 0.00fF
C16018 POR2X1_383/A POR2X1_774/A 0.06fF
C16019 POR2X1_317/a_16_28# POR2X1_169/A 0.03fF
C16020 POR2X1_48/A POR2X1_412/O 0.01fF
C16021 POR2X1_317/A POR2X1_317/B 0.00fF
C16022 POR2X1_692/CTRL POR2X1_20/B 0.01fF
C16023 POR2X1_62/Y POR2X1_408/Y 0.03fF
C16024 VDD POR2X1_90/CTRL 0.00fF
C16025 PAND2X1_634/O POR2X1_37/Y 0.08fF
C16026 POR2X1_507/A POR2X1_260/A 0.02fF
C16027 POR2X1_514/Y POR2X1_343/Y 0.05fF
C16028 VDD POR2X1_354/CTRL 0.00fF
C16029 POR2X1_556/A D_INPUT_0 0.03fF
C16030 POR2X1_814/B PAND2X1_607/CTRL 0.01fF
C16031 VDD POR2X1_91/O 0.00fF
C16032 POR2X1_7/A POR2X1_4/Y 0.03fF
C16033 POR2X1_579/Y POR2X1_568/A 0.02fF
C16034 POR2X1_294/A PAND2X1_103/CTRL2 0.02fF
C16035 POR2X1_848/CTRL POR2X1_734/A 0.06fF
C16036 POR2X1_864/A PAND2X1_829/CTRL 0.00fF
C16037 PAND2X1_432/O POR2X1_648/Y 0.06fF
C16038 POR2X1_43/B POR2X1_522/O 0.21fF
C16039 POR2X1_73/O PAND2X1_341/B 0.01fF
C16040 PAND2X1_212/B POR2X1_20/B 0.03fF
C16041 POR2X1_475/CTRL2 POR2X1_590/A 0.09fF
C16042 POR2X1_81/A PAND2X1_175/B 0.03fF
C16043 PAND2X1_9/Y POR2X1_590/A 0.16fF
C16044 PAND2X1_798/B PAND2X1_332/Y 0.03fF
C16045 POR2X1_152/m4_208_n4# POR2X1_39/B 0.15fF
C16046 PAND2X1_846/CTRL POR2X1_38/B 0.01fF
C16047 PAND2X1_488/a_16_344# POR2X1_814/A 0.01fF
C16048 PAND2X1_73/Y POR2X1_341/A 0.09fF
C16049 POR2X1_545/A POR2X1_568/A 0.03fF
C16050 POR2X1_415/A POR2X1_67/A 0.04fF
C16051 POR2X1_446/A POR2X1_174/A 0.01fF
C16052 POR2X1_243/A POR2X1_243/a_16_28# 0.03fF
C16053 PAND2X1_404/O POR2X1_20/B 0.17fF
C16054 PAND2X1_826/CTRL2 POR2X1_202/B 0.01fF
C16055 POR2X1_76/O POR2X1_296/B 0.01fF
C16056 POR2X1_691/A POR2X1_260/A 0.01fF
C16057 POR2X1_685/CTRL POR2X1_814/A 0.06fF
C16058 PAND2X1_360/Y PAND2X1_359/Y 1.01fF
C16059 POR2X1_302/Y POR2X1_458/Y 0.02fF
C16060 POR2X1_416/B PAND2X1_344/O 0.02fF
C16061 POR2X1_317/Y POR2X1_568/A 0.01fF
C16062 PAND2X1_603/O POR2X1_260/B 0.03fF
C16063 POR2X1_444/Y POR2X1_738/CTRL2 0.03fF
C16064 POR2X1_130/A POR2X1_646/a_16_28# 0.09fF
C16065 POR2X1_20/B POR2X1_268/Y 0.04fF
C16066 PAND2X1_108/CTRL POR2X1_383/A 0.03fF
C16067 POR2X1_85/Y POR2X1_235/CTRL2 0.00fF
C16068 PAND2X1_832/CTRL POR2X1_271/B 0.01fF
C16069 POR2X1_440/B VDD 0.11fF
C16070 POR2X1_707/CTRL2 D_INPUT_4 0.02fF
C16071 PAND2X1_18/B PAND2X1_2/O 0.01fF
C16072 POR2X1_848/O POR2X1_859/A 0.32fF
C16073 D_INPUT_0 PAND2X1_591/O 0.05fF
C16074 POR2X1_66/Y POR2X1_330/Y 0.03fF
C16075 PAND2X1_61/Y POR2X1_20/B 0.02fF
C16076 POR2X1_744/CTRL POR2X1_39/B 0.01fF
C16077 POR2X1_818/Y POR2X1_590/A 0.03fF
C16078 PAND2X1_798/Y PAND2X1_802/B 0.14fF
C16079 PAND2X1_202/O POR2X1_67/Y 0.09fF
C16080 POR2X1_4/Y POR2X1_384/Y 0.08fF
C16081 POR2X1_66/B POR2X1_655/A 0.04fF
C16082 POR2X1_12/A POR2X1_40/Y 0.12fF
C16083 PAND2X1_264/O POR2X1_77/Y 0.03fF
C16084 POR2X1_669/B POR2X1_409/B 0.03fF
C16085 POR2X1_856/B POR2X1_78/A 0.06fF
C16086 POR2X1_316/Y POR2X1_153/Y 0.03fF
C16087 POR2X1_341/A POR2X1_573/CTRL2 0.06fF
C16088 PAND2X1_94/O PAND2X1_58/A 0.17fF
C16089 POR2X1_188/A POR2X1_655/A 0.03fF
C16090 POR2X1_32/A PAND2X1_777/O 0.02fF
C16091 PAND2X1_640/B POR2X1_667/A 0.03fF
C16092 POR2X1_48/A POR2X1_60/A 0.41fF
C16093 POR2X1_416/B PAND2X1_726/B 0.07fF
C16094 PAND2X1_852/A POR2X1_40/Y 0.51fF
C16095 PAND2X1_809/m4_208_n4# POR2X1_7/B 0.09fF
C16096 POR2X1_78/B PAND2X1_41/CTRL2 0.01fF
C16097 PAND2X1_404/A POR2X1_20/B 0.05fF
C16098 POR2X1_428/Y POR2X1_763/A 0.08fF
C16099 POR2X1_440/Y POR2X1_568/A 0.10fF
C16100 POR2X1_48/A POR2X1_591/A 0.01fF
C16101 POR2X1_65/A POR2X1_827/Y 0.00fF
C16102 POR2X1_630/O POR2X1_750/B 0.02fF
C16103 PAND2X1_864/B POR2X1_282/Y 0.03fF
C16104 PAND2X1_848/a_16_344# POR2X1_669/B 0.04fF
C16105 POR2X1_830/Y POR2X1_590/A 0.01fF
C16106 POR2X1_814/A POR2X1_730/O 0.37fF
C16107 POR2X1_66/A POR2X1_200/O 0.01fF
C16108 POR2X1_493/A PAND2X1_41/B 0.04fF
C16109 POR2X1_590/A POR2X1_267/A 6.90fF
C16110 POR2X1_49/Y PAND2X1_571/A 1.26fF
C16111 PAND2X1_283/O POR2X1_814/A 0.01fF
C16112 POR2X1_63/Y PAND2X1_734/B 0.25fF
C16113 PAND2X1_318/CTRL2 POR2X1_20/B 0.00fF
C16114 PAND2X1_658/A PAND2X1_414/O 0.02fF
C16115 D_INPUT_0 POR2X1_72/B 8.08fF
C16116 POR2X1_78/B POR2X1_644/CTRL2 0.01fF
C16117 POR2X1_150/Y PAND2X1_592/Y 0.03fF
C16118 POR2X1_415/A POR2X1_415/O 0.06fF
C16119 POR2X1_836/B POR2X1_836/A 0.02fF
C16120 POR2X1_474/a_56_344# POR2X1_590/A 0.00fF
C16121 POR2X1_544/B PAND2X1_72/A 1.92fF
C16122 POR2X1_38/a_56_344# POR2X1_5/Y 0.00fF
C16123 POR2X1_202/A POR2X1_206/A 0.02fF
C16124 PAND2X1_818/CTRL PAND2X1_340/B 0.01fF
C16125 POR2X1_413/A POR2X1_412/O 0.01fF
C16126 POR2X1_485/a_76_344# PAND2X1_550/B 0.00fF
C16127 POR2X1_814/B POR2X1_220/B 0.07fF
C16128 PAND2X1_55/Y POR2X1_296/a_16_28# 0.03fF
C16129 PAND2X1_622/CTRL2 POR2X1_29/A 0.01fF
C16130 POR2X1_37/Y PAND2X1_333/O 0.12fF
C16131 POR2X1_777/B POR2X1_288/O 0.03fF
C16132 PAND2X1_457/Y PAND2X1_445/Y 0.03fF
C16133 POR2X1_366/Y PAND2X1_268/CTRL2 0.01fF
C16134 POR2X1_851/A VDD 0.00fF
C16135 POR2X1_319/A POR2X1_724/a_56_344# 0.00fF
C16136 POR2X1_656/CTRL POR2X1_362/B 0.01fF
C16137 POR2X1_24/O POR2X1_14/Y 0.01fF
C16138 POR2X1_296/a_16_28# POR2X1_402/A 0.02fF
C16139 POR2X1_66/A VDD 6.19fF
C16140 POR2X1_23/Y POR2X1_256/O 0.29fF
C16141 PAND2X1_93/B POR2X1_722/Y 0.01fF
C16142 POR2X1_20/B POR2X1_255/Y 0.02fF
C16143 PAND2X1_838/B POR2X1_519/Y 0.03fF
C16144 POR2X1_302/B POR2X1_330/Y 0.05fF
C16145 PAND2X1_97/Y POR2X1_91/Y 0.02fF
C16146 POR2X1_23/Y PAND2X1_515/CTRL 0.21fF
C16147 POR2X1_514/Y POR2X1_624/Y 0.03fF
C16148 POR2X1_60/A PAND2X1_513/O 0.05fF
C16149 PAND2X1_236/CTRL POR2X1_590/A 0.00fF
C16150 POR2X1_336/CTRL POR2X1_556/A 0.00fF
C16151 PAND2X1_65/B POR2X1_448/O 0.02fF
C16152 POR2X1_841/B POR2X1_284/O 0.10fF
C16153 POR2X1_12/A POR2X1_587/Y 1.20fF
C16154 POR2X1_60/A PAND2X1_199/A 0.06fF
C16155 POR2X1_841/B PAND2X1_369/O 0.08fF
C16156 POR2X1_462/B POR2X1_472/B 0.00fF
C16157 PAND2X1_248/O POR2X1_294/B 0.02fF
C16158 POR2X1_811/B POR2X1_480/A 0.01fF
C16159 POR2X1_717/O POR2X1_116/A 0.04fF
C16160 PAND2X1_58/A POR2X1_608/O 0.01fF
C16161 POR2X1_41/B PAND2X1_623/CTRL 0.03fF
C16162 POR2X1_13/A POR2X1_422/Y 0.03fF
C16163 POR2X1_259/A POR2X1_61/Y 0.03fF
C16164 D_INPUT_3 POR2X1_411/B 0.03fF
C16165 POR2X1_114/B POR2X1_260/B 0.29fF
C16166 PAND2X1_733/A POR2X1_666/A 0.00fF
C16167 POR2X1_413/A PAND2X1_656/B 0.01fF
C16168 PAND2X1_332/Y POR2X1_184/O 0.06fF
C16169 POR2X1_41/B POR2X1_484/a_16_28# 0.07fF
C16170 POR2X1_119/O POR2X1_37/Y 0.16fF
C16171 POR2X1_629/A POR2X1_629/a_16_28# 0.03fF
C16172 POR2X1_23/Y PAND2X1_445/O 0.04fF
C16173 POR2X1_78/A POR2X1_722/Y 0.16fF
C16174 PAND2X1_478/B VDD 0.02fF
C16175 POR2X1_54/Y POR2X1_38/Y 0.14fF
C16176 POR2X1_302/CTRL POR2X1_302/B 0.01fF
C16177 POR2X1_262/Y PAND2X1_656/A 0.03fF
C16178 PAND2X1_427/O VDD -0.00fF
C16179 POR2X1_257/A POR2X1_280/O 0.07fF
C16180 PAND2X1_206/CTRL POR2X1_40/Y 0.01fF
C16181 POR2X1_102/Y POR2X1_498/O 0.01fF
C16182 POR2X1_437/a_16_28# PAND2X1_190/Y 0.09fF
C16183 POR2X1_257/A PAND2X1_702/a_16_344# 0.02fF
C16184 PAND2X1_404/A PAND2X1_404/a_56_28# 0.00fF
C16185 PAND2X1_620/Y POR2X1_627/CTRL 0.00fF
C16186 POR2X1_150/Y PAND2X1_181/CTRL 0.01fF
C16187 POR2X1_609/CTRL VDD 0.00fF
C16188 PAND2X1_319/B PAND2X1_211/O -0.02fF
C16189 POR2X1_66/A POR2X1_741/Y 1.22fF
C16190 POR2X1_116/m4_208_n4# POR2X1_390/m4_208_n4# 0.13fF
C16191 POR2X1_14/Y POR2X1_754/A 0.03fF
C16192 POR2X1_853/A POR2X1_97/A 0.06fF
C16193 POR2X1_16/A POR2X1_411/A 0.11fF
C16194 POR2X1_842/a_76_344# POR2X1_741/Y 0.00fF
C16195 POR2X1_257/A POR2X1_248/Y 0.04fF
C16196 POR2X1_376/B POR2X1_696/Y 0.07fF
C16197 PAND2X1_81/B POR2X1_66/A 0.08fF
C16198 POR2X1_65/A PAND2X1_206/CTRL2 0.00fF
C16199 POR2X1_79/A PAND2X1_354/A 0.04fF
C16200 PAND2X1_471/a_76_28# POR2X1_83/B 0.02fF
C16201 POR2X1_801/A POR2X1_801/a_16_28# 0.10fF
C16202 D_INPUT_2 POR2X1_414/CTRL2 0.01fF
C16203 POR2X1_487/CTRL2 PAND2X1_794/B 0.01fF
C16204 POR2X1_643/A POR2X1_121/Y 0.03fF
C16205 POR2X1_423/Y POR2X1_256/CTRL 0.01fF
C16206 PAND2X1_278/O INPUT_0 0.04fF
C16207 POR2X1_623/A PAND2X1_9/Y 0.01fF
C16208 POR2X1_291/CTRL2 POR2X1_20/B 0.05fF
C16209 PAND2X1_420/CTRL2 POR2X1_785/A 0.02fF
C16210 PAND2X1_832/a_16_344# PAND2X1_499/Y 0.01fF
C16211 POR2X1_48/A PAND2X1_702/CTRL2 0.01fF
C16212 POR2X1_152/CTRL2 POR2X1_669/B 0.04fF
C16213 PAND2X1_831/Y POR2X1_271/CTRL 0.01fF
C16214 POR2X1_475/CTRL POR2X1_249/Y 0.01fF
C16215 POR2X1_783/A POR2X1_783/a_16_28# 0.09fF
C16216 POR2X1_66/A PAND2X1_125/a_76_28# 0.01fF
C16217 POR2X1_311/Y POR2X1_13/Y 0.10fF
C16218 PAND2X1_609/O PAND2X1_60/B 0.04fF
C16219 POR2X1_60/A PAND2X1_197/Y 0.03fF
C16220 POR2X1_66/A PAND2X1_32/B 0.23fF
C16221 POR2X1_57/A POR2X1_23/Y 0.15fF
C16222 PAND2X1_6/Y PAND2X1_689/O 0.15fF
C16223 PAND2X1_96/B POR2X1_466/A 0.05fF
C16224 PAND2X1_381/Y POR2X1_816/A 0.03fF
C16225 POR2X1_220/a_16_28# POR2X1_220/A 0.05fF
C16226 PAND2X1_557/A POR2X1_488/Y 0.02fF
C16227 POR2X1_366/a_16_28# POR2X1_556/A 0.01fF
C16228 PAND2X1_381/Y D_INPUT_1 0.04fF
C16229 POR2X1_260/B POR2X1_222/A 0.03fF
C16230 PAND2X1_210/O VDD 0.00fF
C16231 PAND2X1_459/O POR2X1_55/Y 0.15fF
C16232 POR2X1_124/O PAND2X1_41/B 0.16fF
C16233 POR2X1_66/B PAND2X1_625/CTRL2 0.03fF
C16234 PAND2X1_362/A PAND2X1_354/O 0.02fF
C16235 PAND2X1_807/B PAND2X1_354/CTRL 0.01fF
C16236 POR2X1_856/B PAND2X1_173/CTRL 0.25fF
C16237 POR2X1_567/B PAND2X1_173/O 0.23fF
C16238 INPUT_1 POR2X1_54/Y 0.20fF
C16239 POR2X1_860/A POR2X1_404/Y 0.00fF
C16240 POR2X1_24/O POR2X1_55/Y 0.18fF
C16241 POR2X1_336/a_16_28# POR2X1_66/A 0.02fF
C16242 POR2X1_516/B POR2X1_236/Y 0.03fF
C16243 POR2X1_23/Y POR2X1_229/Y 0.01fF
C16244 PAND2X1_673/O POR2X1_13/A 0.02fF
C16245 POR2X1_754/Y POR2X1_93/A 0.22fF
C16246 PAND2X1_82/O POR2X1_66/A 0.01fF
C16247 PAND2X1_23/Y POR2X1_654/B 0.07fF
C16248 POR2X1_68/B POR2X1_296/B 0.08fF
C16249 POR2X1_800/A POR2X1_750/B 0.03fF
C16250 POR2X1_52/A POR2X1_696/Y 0.01fF
C16251 POR2X1_517/a_16_28# POR2X1_13/A 0.02fF
C16252 POR2X1_8/Y POR2X1_24/Y 0.01fF
C16253 POR2X1_131/O POR2X1_102/Y 0.01fF
C16254 PAND2X1_787/Y PAND2X1_553/B 0.10fF
C16255 PAND2X1_58/A POR2X1_550/CTRL2 0.01fF
C16256 POR2X1_499/A PAND2X1_48/A 0.03fF
C16257 PAND2X1_794/B POR2X1_40/Y 0.03fF
C16258 POR2X1_516/A POR2X1_48/A 0.06fF
C16259 POR2X1_417/Y PAND2X1_457/CTRL2 0.01fF
C16260 PAND2X1_57/B POR2X1_370/Y 0.03fF
C16261 POR2X1_68/A POR2X1_244/O 0.01fF
C16262 PAND2X1_220/A PAND2X1_388/Y 0.00fF
C16263 POR2X1_66/B PAND2X1_7/a_76_28# 0.02fF
C16264 PAND2X1_48/B POR2X1_555/A 0.16fF
C16265 POR2X1_634/CTRL2 PAND2X1_32/B 0.00fF
C16266 POR2X1_805/Y POR2X1_758/O 0.02fF
C16267 PAND2X1_524/CTRL VDD 0.00fF
C16268 POR2X1_149/A POR2X1_532/A 0.04fF
C16269 PAND2X1_23/Y POR2X1_850/A 0.02fF
C16270 POR2X1_832/O POR2X1_722/Y 0.01fF
C16271 POR2X1_278/a_16_28# PAND2X1_35/Y 0.01fF
C16272 POR2X1_814/B POR2X1_756/a_16_28# 0.03fF
C16273 POR2X1_362/B POR2X1_717/Y 0.68fF
C16274 PAND2X1_215/B PAND2X1_723/Y 0.14fF
C16275 PAND2X1_479/CTRL POR2X1_599/A 0.14fF
C16276 POR2X1_257/A PAND2X1_708/O 0.07fF
C16277 POR2X1_855/B POR2X1_801/B 0.02fF
C16278 PAND2X1_41/CTRL2 POR2X1_294/A 0.00fF
C16279 POR2X1_102/Y POR2X1_172/Y 0.02fF
C16280 POR2X1_792/B VDD 0.04fF
C16281 POR2X1_334/Y POR2X1_99/Y 0.27fF
C16282 POR2X1_750/B POR2X1_702/A 0.05fF
C16283 PAND2X1_825/CTRL2 POR2X1_296/B 0.00fF
C16284 POR2X1_612/Y POR2X1_4/CTRL2 0.03fF
C16285 PAND2X1_632/A POR2X1_496/Y 0.06fF
C16286 POR2X1_802/B VDD 0.03fF
C16287 PAND2X1_220/Y PAND2X1_357/Y 0.03fF
C16288 PAND2X1_93/B POR2X1_799/a_16_28# 0.03fF
C16289 INPUT_2 POR2X1_94/A 0.03fF
C16290 PAND2X1_651/Y PAND2X1_500/O 0.47fF
C16291 POR2X1_832/CTRL POR2X1_832/B 0.01fF
C16292 PAND2X1_253/O POR2X1_66/A 0.02fF
C16293 POR2X1_494/Y VDD 0.18fF
C16294 POR2X1_650/A POR2X1_391/Y 0.19fF
C16295 PAND2X1_575/B POR2X1_91/Y 0.03fF
C16296 PAND2X1_93/B POR2X1_244/Y 0.11fF
C16297 POR2X1_111/Y POR2X1_23/Y 0.02fF
C16298 POR2X1_673/Y POR2X1_66/A 13.33fF
C16299 POR2X1_814/A POR2X1_736/A 0.05fF
C16300 PAND2X1_6/A PAND2X1_381/CTRL 0.01fF
C16301 PAND2X1_180/CTRL PAND2X1_566/Y 0.01fF
C16302 POR2X1_13/A PAND2X1_465/B 0.02fF
C16303 PAND2X1_20/A PAND2X1_397/CTRL 0.01fF
C16304 POR2X1_355/B POR2X1_356/A 0.05fF
C16305 POR2X1_68/A POR2X1_483/A 0.05fF
C16306 POR2X1_616/Y POR2X1_415/A 0.08fF
C16307 POR2X1_120/CTRL2 POR2X1_712/Y 0.03fF
C16308 POR2X1_78/B PAND2X1_144/O 0.15fF
C16309 PAND2X1_844/Y PAND2X1_351/Y 0.02fF
C16310 PAND2X1_480/B POR2X1_55/Y 0.05fF
C16311 POR2X1_222/Y VDD 0.75fF
C16312 POR2X1_57/A POR2X1_312/Y 0.04fF
C16313 PAND2X1_659/B PAND2X1_575/A 0.03fF
C16314 PAND2X1_483/CTRL POR2X1_669/B 0.04fF
C16315 POR2X1_456/a_76_344# POR2X1_702/A 0.01fF
C16316 POR2X1_322/Y POR2X1_40/Y 0.01fF
C16317 POR2X1_52/A POR2X1_163/A 0.08fF
C16318 POR2X1_16/A POR2X1_32/A 1.80fF
C16319 PAND2X1_592/Y PAND2X1_364/B 0.09fF
C16320 POR2X1_135/O POR2X1_257/A 0.01fF
C16321 POR2X1_410/O POR2X1_790/B 0.09fF
C16322 POR2X1_482/Y PAND2X1_549/B 0.03fF
C16323 POR2X1_631/A POR2X1_852/B -0.02fF
C16324 POR2X1_68/A PAND2X1_8/Y 0.10fF
C16325 POR2X1_159/CTRL PAND2X1_63/B 0.01fF
C16326 D_INPUT_0 PAND2X1_749/O 0.15fF
C16327 POR2X1_61/Y PAND2X1_88/Y 0.03fF
C16328 POR2X1_57/A POR2X1_323/CTRL 0.01fF
C16329 PAND2X1_848/B POR2X1_820/Y 0.00fF
C16330 POR2X1_460/A PAND2X1_21/CTRL2 0.00fF
C16331 PAND2X1_739/Y PAND2X1_357/Y 0.08fF
C16332 POR2X1_13/A PAND2X1_798/B 0.01fF
C16333 POR2X1_79/Y PAND2X1_730/CTRL 0.01fF
C16334 POR2X1_149/B POR2X1_435/Y 0.03fF
C16335 POR2X1_38/Y PAND2X1_340/a_16_344# 0.02fF
C16336 PAND2X1_491/CTRL2 INPUT_0 0.06fF
C16337 POR2X1_62/Y PAND2X1_28/a_76_28# 0.02fF
C16338 D_INPUT_3 POR2X1_376/B 0.19fF
C16339 PAND2X1_140/A PAND2X1_220/Y 0.03fF
C16340 PAND2X1_568/O PAND2X1_566/Y 0.02fF
C16341 PAND2X1_48/O POR2X1_786/Y 0.30fF
C16342 PAND2X1_659/Y PAND2X1_205/A 0.14fF
C16343 PAND2X1_388/Y POR2X1_106/Y 0.03fF
C16344 POR2X1_68/B POR2X1_547/B 0.51fF
C16345 PAND2X1_57/B POR2X1_770/CTRL2 0.00fF
C16346 PAND2X1_392/B PAND2X1_383/O 0.03fF
C16347 POR2X1_777/B POR2X1_101/Y 0.13fF
C16348 POR2X1_96/A POR2X1_816/A 3.74fF
C16349 POR2X1_627/a_76_344# POR2X1_93/A 0.01fF
C16350 POR2X1_502/A PAND2X1_144/a_76_28# 0.02fF
C16351 PAND2X1_48/B PAND2X1_145/O 0.04fF
C16352 PAND2X1_770/O POR2X1_73/Y 0.02fF
C16353 POR2X1_532/A VDD 5.81fF
C16354 POR2X1_16/A POR2X1_417/Y 0.00fF
C16355 POR2X1_502/A POR2X1_544/CTRL2 0.01fF
C16356 PAND2X1_41/B POR2X1_276/Y 2.70fF
C16357 D_INPUT_5 D_INPUT_4 3.84fF
C16358 PAND2X1_90/Y POR2X1_407/CTRL2 0.03fF
C16359 PAND2X1_499/Y PAND2X1_175/B 0.03fF
C16360 INPUT_1 PAND2X1_23/CTRL 0.01fF
C16361 PAND2X1_94/A PAND2X1_23/a_16_344# 0.01fF
C16362 POR2X1_114/B PAND2X1_55/Y 0.04fF
C16363 POR2X1_294/B POR2X1_391/Y 0.10fF
C16364 INPUT_1 PAND2X1_73/a_76_28# 0.02fF
C16365 POR2X1_308/CTRL2 POR2X1_725/Y 0.02fF
C16366 POR2X1_283/A PAND2X1_473/B 2.98fF
C16367 POR2X1_49/Y POR2X1_313/Y 0.03fF
C16368 POR2X1_135/Y POR2X1_7/A 0.24fF
C16369 POR2X1_734/A POR2X1_260/A 0.12fF
C16370 POR2X1_691/B VDD 0.14fF
C16371 PAND2X1_65/B POR2X1_101/Y 0.12fF
C16372 PAND2X1_48/B POR2X1_705/O 0.17fF
C16373 POR2X1_708/m4_208_n4# PAND2X1_32/B 0.15fF
C16374 PAND2X1_139/B PAND2X1_130/CTRL 0.00fF
C16375 POR2X1_832/B POR2X1_804/A 0.05fF
C16376 POR2X1_840/B POR2X1_579/Y 0.03fF
C16377 PAND2X1_57/B POR2X1_359/Y 0.04fF
C16378 POR2X1_206/A POR2X1_201/Y 0.01fF
C16379 POR2X1_722/Y POR2X1_513/CTRL2 0.01fF
C16380 POR2X1_327/Y POR2X1_453/a_56_344# 0.03fF
C16381 POR2X1_514/Y POR2X1_139/CTRL 0.01fF
C16382 POR2X1_68/A POR2X1_61/B 0.01fF
C16383 PAND2X1_444/O POR2X1_39/B 0.04fF
C16384 PAND2X1_69/A POR2X1_42/Y 0.07fF
C16385 POR2X1_62/Y POR2X1_60/A 0.07fF
C16386 POR2X1_722/Y PAND2X1_306/O 0.02fF
C16387 POR2X1_416/B PAND2X1_35/A 0.03fF
C16388 PAND2X1_309/O POR2X1_335/B 0.02fF
C16389 POR2X1_706/A INPUT_1 0.04fF
C16390 POR2X1_52/A D_INPUT_3 0.03fF
C16391 POR2X1_301/O POR2X1_68/A 0.06fF
C16392 POR2X1_71/Y POR2X1_91/Y 0.01fF
C16393 POR2X1_236/Y POR2X1_172/O 0.07fF
C16394 POR2X1_628/a_16_28# PAND2X1_6/A 0.00fF
C16395 POR2X1_840/B POR2X1_572/B 0.05fF
C16396 POR2X1_49/Y PAND2X1_844/O 0.15fF
C16397 POR2X1_222/Y PAND2X1_32/B 0.03fF
C16398 POR2X1_96/A PAND2X1_854/A 0.02fF
C16399 POR2X1_49/Y POR2X1_144/CTRL 0.01fF
C16400 POR2X1_787/O POR2X1_325/A 0.01fF
C16401 POR2X1_326/A POR2X1_436/O 0.18fF
C16402 PAND2X1_56/Y POR2X1_196/Y 0.08fF
C16403 POR2X1_93/A POR2X1_42/Y 0.07fF
C16404 PAND2X1_83/O POR2X1_35/Y 0.02fF
C16405 PAND2X1_562/a_76_28# PAND2X1_566/Y 0.03fF
C16406 POR2X1_78/B POR2X1_456/B 0.15fF
C16407 POR2X1_647/CTRL2 PAND2X1_52/B 0.01fF
C16408 POR2X1_693/Y POR2X1_73/Y 0.01fF
C16409 POR2X1_83/B PAND2X1_352/B 0.01fF
C16410 POR2X1_532/A POR2X1_741/Y 0.06fF
C16411 POR2X1_245/Y POR2X1_7/B 0.05fF
C16412 PAND2X1_21/O POR2X1_260/A 0.02fF
C16413 PAND2X1_275/O POR2X1_573/A 0.04fF
C16414 PAND2X1_691/Y POR2X1_13/A 0.03fF
C16415 POR2X1_447/B POR2X1_630/A 0.06fF
C16416 POR2X1_346/CTRL POR2X1_68/A 0.01fF
C16417 POR2X1_690/Y POR2X1_689/Y 0.09fF
C16418 PAND2X1_676/O POR2X1_599/A 0.00fF
C16419 POR2X1_35/Y PAND2X1_88/Y 6.79fF
C16420 PAND2X1_76/Y POR2X1_129/Y 0.03fF
C16421 PAND2X1_216/B INPUT_0 0.02fF
C16422 PAND2X1_390/Y PAND2X1_851/O 0.02fF
C16423 POR2X1_614/A POR2X1_840/B 0.03fF
C16424 PAND2X1_602/Y POR2X1_757/CTRL 0.02fF
C16425 PAND2X1_55/Y POR2X1_222/A 0.03fF
C16426 POR2X1_355/B POR2X1_570/Y 0.07fF
C16427 POR2X1_294/B PAND2X1_528/CTRL2 0.14fF
C16428 POR2X1_16/A PAND2X1_35/Y 0.08fF
C16429 POR2X1_529/Y PAND2X1_658/A 0.00fF
C16430 PAND2X1_495/O POR2X1_786/Y 0.03fF
C16431 POR2X1_371/CTRL2 POR2X1_5/Y 0.01fF
C16432 POR2X1_57/A PAND2X1_836/O 0.01fF
C16433 POR2X1_709/a_16_28# POR2X1_502/A 0.02fF
C16434 PAND2X1_62/a_76_28# POR2X1_394/A 0.04fF
C16435 PAND2X1_190/Y PAND2X1_843/Y 0.05fF
C16436 POR2X1_532/A PAND2X1_32/B 0.30fF
C16437 PAND2X1_390/O POR2X1_283/A 0.09fF
C16438 PAND2X1_553/B PAND2X1_114/O 0.10fF
C16439 PAND2X1_388/Y PAND2X1_337/A 0.01fF
C16440 POR2X1_16/A POR2X1_57/CTRL -0.02fF
C16441 PAND2X1_25/CTRL2 PAND2X1_52/B 0.03fF
C16442 PAND2X1_118/O POR2X1_123/A 0.02fF
C16443 POR2X1_81/A PAND2X1_244/a_56_28# 0.00fF
C16444 POR2X1_855/B POR2X1_796/CTRL2 0.01fF
C16445 POR2X1_599/A PAND2X1_723/A 0.10fF
C16446 POR2X1_210/CTRL2 PAND2X1_52/B 0.01fF
C16447 POR2X1_532/A POR2X1_711/O 0.25fF
C16448 POR2X1_828/O POR2X1_260/A 0.02fF
C16449 POR2X1_834/Y POR2X1_294/B 0.10fF
C16450 PAND2X1_433/m4_208_n4# POR2X1_832/A 0.07fF
C16451 POR2X1_539/O POR2X1_662/Y 0.18fF
C16452 PAND2X1_689/O PAND2X1_52/B 0.01fF
C16453 POR2X1_7/A POR2X1_816/A 0.03fF
C16454 POR2X1_552/CTRL VDD -0.00fF
C16455 POR2X1_7/B PAND2X1_507/CTRL 0.02fF
C16456 POR2X1_417/CTRL POR2X1_387/Y 0.07fF
C16457 POR2X1_65/A PAND2X1_797/Y 0.03fF
C16458 PAND2X1_341/A PAND2X1_99/Y 0.13fF
C16459 D_INPUT_1 POR2X1_7/A 0.07fF
C16460 POR2X1_38/B POR2X1_384/CTRL2 0.01fF
C16461 POR2X1_16/A POR2X1_189/Y 0.05fF
C16462 POR2X1_750/A POR2X1_39/B 0.03fF
C16463 PAND2X1_534/CTRL POR2X1_788/B 0.01fF
C16464 POR2X1_325/CTRL POR2X1_542/B 0.01fF
C16465 POR2X1_383/A POR2X1_638/Y 0.03fF
C16466 POR2X1_48/Y PAND2X1_196/a_76_28# 0.02fF
C16467 POR2X1_390/B POR2X1_301/CTRL 0.00fF
C16468 PAND2X1_341/B VDD 0.42fF
C16469 PAND2X1_500/CTRL2 POR2X1_497/Y 0.01fF
C16470 PAND2X1_793/Y PAND2X1_508/Y 0.06fF
C16471 D_INPUT_6 PAND2X1_1/CTRL2 0.01fF
C16472 POR2X1_416/B POR2X1_255/CTRL 0.01fF
C16473 PAND2X1_48/B PAND2X1_484/CTRL 0.01fF
C16474 POR2X1_359/CTRL PAND2X1_57/B 0.01fF
C16475 POR2X1_590/A POR2X1_568/A 0.03fF
C16476 PAND2X1_710/O PAND2X1_711/A 0.02fF
C16477 PAND2X1_658/O POR2X1_77/Y 0.04fF
C16478 PAND2X1_574/CTRL POR2X1_73/Y 0.01fF
C16479 POR2X1_333/O PAND2X1_32/B 0.01fF
C16480 PAND2X1_83/a_56_28# PAND2X1_82/Y 0.00fF
C16481 PAND2X1_352/Y VDD 0.00fF
C16482 POR2X1_510/Y POR2X1_228/Y 0.10fF
C16483 POR2X1_786/Y POR2X1_260/A 0.04fF
C16484 PAND2X1_684/O POR2X1_149/B 0.02fF
C16485 PAND2X1_388/Y PAND2X1_349/A 0.03fF
C16486 PAND2X1_23/Y POR2X1_54/CTRL 0.00fF
C16487 POR2X1_9/Y PAND2X1_66/a_16_344# 0.04fF
C16488 POR2X1_537/B POR2X1_537/A 0.02fF
C16489 POR2X1_52/A POR2X1_83/Y 0.04fF
C16490 POR2X1_814/B POR2X1_716/O 0.01fF
C16491 POR2X1_394/A PAND2X1_547/CTRL 0.01fF
C16492 POR2X1_101/O PAND2X1_60/B 0.08fF
C16493 POR2X1_567/A POR2X1_231/CTRL 0.13fF
C16494 PAND2X1_349/A PAND2X1_549/B 0.03fF
C16495 POR2X1_270/CTRL POR2X1_456/B 0.02fF
C16496 POR2X1_293/Y PAND2X1_506/Y 0.07fF
C16497 POR2X1_158/Y POR2X1_427/Y 0.00fF
C16498 POR2X1_673/Y POR2X1_532/A 0.03fF
C16499 PAND2X1_476/A PAND2X1_364/B 0.07fF
C16500 POR2X1_54/Y POR2X1_462/O 0.01fF
C16501 POR2X1_135/O PAND2X1_553/B 0.01fF
C16502 POR2X1_722/B POR2X1_722/a_16_28# 0.02fF
C16503 POR2X1_493/CTRL POR2X1_773/B 0.03fF
C16504 PAND2X1_23/Y PAND2X1_396/CTRL2 -0.00fF
C16505 PAND2X1_6/A PAND2X1_502/O 0.07fF
C16506 VDD POR2X1_533/Y 0.08fF
C16507 POR2X1_42/Y POR2X1_397/O 0.01fF
C16508 POR2X1_540/Y PAND2X1_178/CTRL 0.01fF
C16509 POR2X1_116/A POR2X1_276/B 0.02fF
C16510 POR2X1_14/Y POR2X1_386/Y 0.03fF
C16511 POR2X1_384/Y POR2X1_816/A 0.00fF
C16512 POR2X1_707/B POR2X1_635/B 0.05fF
C16513 POR2X1_513/B PAND2X1_304/a_56_28# 0.00fF
C16514 POR2X1_270/Y POR2X1_814/A 0.40fF
C16515 PAND2X1_639/Y POR2X1_584/CTRL2 0.06fF
C16516 PAND2X1_57/B POR2X1_342/A 0.01fF
C16517 POR2X1_736/a_16_28# POR2X1_675/Y 0.03fF
C16518 PAND2X1_281/CTRL POR2X1_649/B 0.01fF
C16519 POR2X1_278/A PAND2X1_560/B 0.03fF
C16520 POR2X1_38/Y PAND2X1_120/O 0.01fF
C16521 POR2X1_472/a_16_28# POR2X1_463/Y 0.05fF
C16522 POR2X1_294/B POR2X1_383/Y 0.06fF
C16523 POR2X1_416/B POR2X1_411/CTRL 0.01fF
C16524 PAND2X1_269/CTRL2 POR2X1_39/B 0.01fF
C16525 POR2X1_236/Y POR2X1_167/Y 0.24fF
C16526 PAND2X1_850/Y PAND2X1_469/B 0.07fF
C16527 PAND2X1_55/Y POR2X1_513/A 0.04fF
C16528 PAND2X1_94/A PAND2X1_184/CTRL 0.00fF
C16529 PAND2X1_470/O POR2X1_119/Y 0.17fF
C16530 POR2X1_446/B POR2X1_446/A -0.01fF
C16531 POR2X1_342/Y POR2X1_294/B 0.03fF
C16532 PAND2X1_73/Y POR2X1_828/a_16_28# 0.02fF
C16533 POR2X1_355/B PAND2X1_72/A 0.10fF
C16534 POR2X1_38/Y POR2X1_4/Y 0.14fF
C16535 PAND2X1_716/B POR2X1_387/Y 0.07fF
C16536 POR2X1_35/Y POR2X1_568/B 0.03fF
C16537 POR2X1_396/CTRL2 POR2X1_39/B 0.00fF
C16538 POR2X1_126/a_16_28# POR2X1_411/B 0.01fF
C16539 PAND2X1_272/CTRL2 POR2X1_556/A 0.01fF
C16540 POR2X1_97/O POR2X1_186/B 0.02fF
C16541 POR2X1_554/B POR2X1_657/CTRL2 0.03fF
C16542 POR2X1_416/B POR2X1_43/B 0.16fF
C16543 POR2X1_447/B POR2X1_383/A 0.00fF
C16544 PAND2X1_9/Y POR2X1_66/A 0.05fF
C16545 PAND2X1_532/O POR2X1_394/A 0.00fF
C16546 PAND2X1_323/a_16_344# PAND2X1_111/B 0.01fF
C16547 POR2X1_165/CTRL PAND2X1_326/B 0.01fF
C16548 PAND2X1_189/CTRL POR2X1_353/A 0.05fF
C16549 POR2X1_456/B POR2X1_180/O 0.10fF
C16550 POR2X1_644/O POR2X1_260/B 0.01fF
C16551 PAND2X1_20/A POR2X1_296/CTRL 0.01fF
C16552 PAND2X1_731/O POR2X1_77/Y 0.01fF
C16553 POR2X1_863/B POR2X1_863/A 0.13fF
C16554 POR2X1_456/B POR2X1_294/A 0.03fF
C16555 POR2X1_416/B PAND2X1_547/a_16_344# 0.00fF
C16556 POR2X1_39/B PAND2X1_509/O 0.04fF
C16557 POR2X1_866/A PAND2X1_93/B 0.10fF
C16558 POR2X1_166/a_16_28# PAND2X1_326/B 0.01fF
C16559 POR2X1_461/B POR2X1_846/A 0.02fF
C16560 POR2X1_416/B POR2X1_38/B 0.05fF
C16561 PAND2X1_69/A POR2X1_343/m4_208_n4# 0.08fF
C16562 POR2X1_87/CTRL POR2X1_38/B 0.01fF
C16563 POR2X1_537/Y POR2X1_851/CTRL2 0.01fF
C16564 INPUT_1 POR2X1_4/Y 16.84fF
C16565 PAND2X1_826/CTRL POR2X1_296/B 0.02fF
C16566 POR2X1_68/Y POR2X1_296/B 0.01fF
C16567 PAND2X1_464/CTRL2 POR2X1_417/Y 0.01fF
C16568 POR2X1_71/a_16_28# POR2X1_394/A 0.07fF
C16569 POR2X1_864/A POR2X1_330/Y 0.05fF
C16570 POR2X1_383/A POR2X1_510/O 0.01fF
C16571 PAND2X1_31/O PAND2X1_3/A 0.04fF
C16572 POR2X1_210/Y PAND2X1_52/B 0.04fF
C16573 POR2X1_791/B PAND2X1_72/A 0.01fF
C16574 PAND2X1_288/A GATE_222 0.01fF
C16575 POR2X1_667/CTRL VDD 0.00fF
C16576 PAND2X1_39/B POR2X1_400/CTRL 0.01fF
C16577 PAND2X1_93/B POR2X1_269/CTRL2 0.01fF
C16578 POR2X1_66/B POR2X1_647/B 0.52fF
C16579 POR2X1_594/CTRL2 POR2X1_385/Y 0.01fF
C16580 POR2X1_866/A POR2X1_78/A 0.03fF
C16581 POR2X1_313/a_56_344# POR2X1_167/Y 0.00fF
C16582 POR2X1_707/B PAND2X1_762/CTRL2 0.01fF
C16583 POR2X1_265/CTRL2 POR2X1_667/A 0.00fF
C16584 PAND2X1_20/A POR2X1_34/CTRL 0.01fF
C16585 POR2X1_569/A POR2X1_500/CTRL2 0.02fF
C16586 POR2X1_669/B POR2X1_626/CTRL2 0.03fF
C16587 PAND2X1_73/Y POR2X1_678/Y 0.03fF
C16588 POR2X1_550/Y PAND2X1_52/B 0.11fF
C16589 PAND2X1_611/O POR2X1_130/A 0.05fF
C16590 POR2X1_510/B PAND2X1_72/A 0.07fF
C16591 POR2X1_141/Y POR2X1_446/B 0.10fF
C16592 PAND2X1_620/Y POR2X1_628/Y 0.03fF
C16593 POR2X1_614/A POR2X1_661/A 0.07fF
C16594 POR2X1_263/O POR2X1_236/Y 0.04fF
C16595 POR2X1_129/CTRL2 POR2X1_83/B 0.00fF
C16596 PAND2X1_659/Y PAND2X1_737/CTRL 0.01fF
C16597 PAND2X1_605/a_76_28# POR2X1_32/A 0.02fF
C16598 POR2X1_102/Y PAND2X1_590/a_16_344# 0.01fF
C16599 POR2X1_441/Y PAND2X1_544/O 0.02fF
C16600 PAND2X1_467/B POR2X1_695/Y 0.02fF
C16601 POR2X1_52/A POR2X1_815/CTRL 0.01fF
C16602 PAND2X1_124/Y POR2X1_40/Y 0.03fF
C16603 POR2X1_78/B PAND2X1_81/a_76_28# 0.00fF
C16604 POR2X1_454/A PAND2X1_229/CTRL 0.02fF
C16605 POR2X1_120/CTRL2 PAND2X1_39/B 0.00fF
C16606 POR2X1_837/B PAND2X1_69/A 0.00fF
C16607 PAND2X1_859/A POR2X1_93/Y 0.02fF
C16608 PAND2X1_502/CTRL2 POR2X1_77/Y 0.01fF
C16609 POR2X1_452/Y VDD 0.00fF
C16610 POR2X1_68/A POR2X1_630/B 0.01fF
C16611 POR2X1_808/A POR2X1_66/A 0.02fF
C16612 POR2X1_20/B POR2X1_46/Y 0.08fF
C16613 PAND2X1_116/CTRL2 POR2X1_48/A 0.01fF
C16614 POR2X1_748/A POR2X1_496/Y 0.10fF
C16615 POR2X1_159/CTRL POR2X1_32/A 0.01fF
C16616 POR2X1_655/CTRL2 POR2X1_307/A 0.00fF
C16617 GATE_479 POR2X1_48/A 0.03fF
C16618 POR2X1_67/a_16_28# POR2X1_5/Y 0.07fF
C16619 PAND2X1_55/Y POR2X1_659/m4_208_n4# 0.08fF
C16620 PAND2X1_860/A PAND2X1_175/CTRL2 0.01fF
C16621 POR2X1_453/O POR2X1_590/A 0.04fF
C16622 POR2X1_98/CTRL PAND2X1_41/B 0.01fF
C16623 POR2X1_834/a_56_344# POR2X1_330/Y 0.03fF
C16624 PAND2X1_833/a_76_28# POR2X1_257/A 0.02fF
C16625 PAND2X1_244/O POR2X1_102/Y 0.01fF
C16626 POR2X1_734/B POR2X1_362/B 0.12fF
C16627 POR2X1_479/B POR2X1_286/Y 0.00fF
C16628 PAND2X1_266/CTRL2 POR2X1_73/Y 0.03fF
C16629 PAND2X1_404/Y PAND2X1_84/a_56_28# 0.00fF
C16630 POR2X1_446/B POR2X1_220/Y 0.03fF
C16631 PAND2X1_776/Y POR2X1_236/Y 0.02fF
C16632 POR2X1_846/Y PAND2X1_6/A 0.03fF
C16633 POR2X1_838/B POR2X1_837/Y 0.04fF
C16634 POR2X1_83/B POR2X1_40/Y 7.72fF
C16635 POR2X1_76/A PAND2X1_516/O 0.07fF
C16636 PAND2X1_454/O POR2X1_424/Y 0.07fF
C16637 POR2X1_23/Y PAND2X1_84/Y 0.10fF
C16638 POR2X1_67/Y POR2X1_619/A 0.03fF
C16639 POR2X1_850/A POR2X1_656/O 0.01fF
C16640 POR2X1_66/B POR2X1_461/A 0.01fF
C16641 POR2X1_863/A POR2X1_724/B 0.01fF
C16642 POR2X1_20/B PAND2X1_334/O 0.04fF
C16643 PAND2X1_48/B PAND2X1_268/O 0.02fF
C16644 POR2X1_268/O POR2X1_5/Y 0.08fF
C16645 POR2X1_260/B POR2X1_405/Y 0.01fF
C16646 POR2X1_175/CTRL2 PAND2X1_73/Y 0.01fF
C16647 POR2X1_688/CTRL2 POR2X1_532/A 0.03fF
C16648 POR2X1_260/B POR2X1_784/A 0.03fF
C16649 POR2X1_220/B VDD 0.99fF
C16650 PAND2X1_811/O PAND2X1_811/A 0.00fF
C16651 POR2X1_105/a_56_344# PAND2X1_41/B 0.00fF
C16652 PAND2X1_169/Y PAND2X1_731/B 0.06fF
C16653 POR2X1_480/A POR2X1_296/B 0.10fF
C16654 PAND2X1_80/CTRL2 POR2X1_296/B 0.00fF
C16655 PAND2X1_20/A POR2X1_402/O 0.01fF
C16656 POR2X1_818/Y PAND2X1_751/O 0.02fF
C16657 POR2X1_814/B PAND2X1_616/CTRL2 0.02fF
C16658 POR2X1_566/A POR2X1_444/A 0.04fF
C16659 POR2X1_120/CTRL2 POR2X1_805/Y 0.03fF
C16660 POR2X1_60/A PAND2X1_333/O 0.05fF
C16661 POR2X1_306/Y PAND2X1_512/O 0.00fF
C16662 POR2X1_541/B POR2X1_203/Y 0.03fF
C16663 PAND2X1_214/O PAND2X1_35/Y 0.02fF
C16664 POR2X1_660/Y VDD 0.34fF
C16665 POR2X1_692/CTRL POR2X1_763/Y 0.08fF
C16666 PAND2X1_57/CTRL POR2X1_590/A 0.01fF
C16667 PAND2X1_655/B POR2X1_600/m4_208_n4# 0.09fF
C16668 POR2X1_814/A POR2X1_101/Y 0.22fF
C16669 POR2X1_397/Y POR2X1_14/Y 0.03fF
C16670 PAND2X1_675/A POR2X1_437/CTRL 0.01fF
C16671 POR2X1_653/B POR2X1_750/B 0.03fF
C16672 PAND2X1_798/B POR2X1_437/O 0.01fF
C16673 PAND2X1_9/Y POR2X1_532/A 0.06fF
C16674 POR2X1_52/A POR2X1_484/CTRL 0.01fF
C16675 D_INPUT_0 POR2X1_7/B 0.03fF
C16676 POR2X1_102/Y POR2X1_481/A 0.02fF
C16677 PAND2X1_116/O POR2X1_40/Y 0.03fF
C16678 POR2X1_13/A POR2X1_423/CTRL 0.01fF
C16679 POR2X1_676/O POR2X1_828/A 0.08fF
C16680 POR2X1_676/CTRL PAND2X1_69/A 0.01fF
C16681 PAND2X1_58/A PAND2X1_8/Y 0.07fF
C16682 PAND2X1_561/Y PAND2X1_571/Y 0.02fF
C16683 POR2X1_362/B POR2X1_330/Y 0.28fF
C16684 PAND2X1_402/CTRL POR2X1_5/Y 0.02fF
C16685 POR2X1_48/A PAND2X1_649/CTRL2 0.00fF
C16686 POR2X1_400/O POR2X1_206/A 0.01fF
C16687 PAND2X1_766/a_16_344# PAND2X1_90/Y 0.02fF
C16688 PAND2X1_308/B POR2X1_14/Y 0.03fF
C16689 POR2X1_636/O POR2X1_636/A 0.08fF
C16690 POR2X1_660/O POR2X1_307/Y 0.00fF
C16691 POR2X1_423/CTRL2 POR2X1_293/Y 0.01fF
C16692 POR2X1_40/Y PAND2X1_140/Y 0.03fF
C16693 POR2X1_181/a_16_28# PAND2X1_72/A 0.00fF
C16694 PAND2X1_308/B PAND2X1_453/A 0.04fF
C16695 POR2X1_451/CTRL2 POR2X1_635/Y 0.02fF
C16696 POR2X1_48/A PAND2X1_35/a_16_344# 0.01fF
C16697 PAND2X1_57/B PAND2X1_701/m4_208_n4# 0.07fF
C16698 PAND2X1_287/Y PAND2X1_773/O 0.08fF
C16699 POR2X1_123/CTRL POR2X1_78/A 0.01fF
C16700 POR2X1_294/Y D_GATE_741 0.04fF
C16701 POR2X1_644/O POR2X1_407/Y 0.01fF
C16702 INPUT_3 POR2X1_7/A 0.23fF
C16703 PAND2X1_90/A POR2X1_296/B 0.08fF
C16704 PAND2X1_473/Y PAND2X1_561/A 0.35fF
C16705 POR2X1_56/O POR2X1_55/Y 0.17fF
C16706 POR2X1_81/O POR2X1_293/Y 0.02fF
C16707 POR2X1_440/Y POR2X1_477/O 0.02fF
C16708 POR2X1_614/A POR2X1_266/a_16_28# 0.09fF
C16709 POR2X1_458/O PAND2X1_32/B 0.01fF
C16710 POR2X1_78/B POR2X1_398/Y 0.01fF
C16711 POR2X1_72/B PAND2X1_735/Y 0.19fF
C16712 PAND2X1_52/B POR2X1_181/Y 0.06fF
C16713 PAND2X1_449/CTRL PAND2X1_308/Y 0.01fF
C16714 PAND2X1_676/CTRL2 PAND2X1_205/A 0.00fF
C16715 POR2X1_283/CTRL PAND2X1_365/B 0.01fF
C16716 POR2X1_671/CTRL POR2X1_5/Y 0.01fF
C16717 PAND2X1_307/CTRL POR2X1_56/B 0.01fF
C16718 PAND2X1_73/Y POR2X1_805/A 0.68fF
C16719 POR2X1_48/Y POR2X1_60/A 0.01fF
C16720 POR2X1_329/A PAND2X1_657/B 0.04fF
C16721 POR2X1_454/A POR2X1_510/Y 0.03fF
C16722 PAND2X1_73/Y POR2X1_712/Y 0.03fF
C16723 POR2X1_186/Y POR2X1_468/B 0.05fF
C16724 POR2X1_98/CTRL2 POR2X1_68/B 0.04fF
C16725 POR2X1_639/Y POR2X1_66/A 0.12fF
C16726 POR2X1_820/Y POR2X1_5/Y 0.01fF
C16727 PAND2X1_80/CTRL2 POR2X1_547/B 0.01fF
C16728 PAND2X1_84/Y PAND2X1_558/O 0.02fF
C16729 POR2X1_60/A PAND2X1_652/A 0.06fF
C16730 POR2X1_662/O POR2X1_725/Y 0.05fF
C16731 POR2X1_78/B POR2X1_608/CTRL2 0.03fF
C16732 PAND2X1_72/A PAND2X1_135/CTRL 0.01fF
C16733 POR2X1_832/B POR2X1_794/B 0.03fF
C16734 POR2X1_13/A PAND2X1_828/CTRL2 0.00fF
C16735 PAND2X1_58/A POR2X1_61/B 0.01fF
C16736 POR2X1_657/a_16_28# POR2X1_741/Y 0.01fF
C16737 PAND2X1_769/O VDD 0.00fF
C16738 PAND2X1_455/O POR2X1_7/B 0.17fF
C16739 POR2X1_497/Y VDD 0.02fF
C16740 POR2X1_72/B PAND2X1_493/Y 0.06fF
C16741 POR2X1_625/CTRL2 POR2X1_754/A 0.00fF
C16742 PAND2X1_480/B PAND2X1_276/O 0.02fF
C16743 PAND2X1_23/Y POR2X1_777/B 0.10fF
C16744 POR2X1_245/O POR2X1_37/Y 0.16fF
C16745 POR2X1_65/A POR2X1_372/Y 0.08fF
C16746 PAND2X1_416/O POR2X1_260/A 0.03fF
C16747 POR2X1_840/B POR2X1_590/A 0.09fF
C16748 PAND2X1_802/CTRL2 POR2X1_760/A 0.01fF
C16749 POR2X1_72/B PAND2X1_174/O 0.01fF
C16750 POR2X1_78/A POR2X1_501/B 0.03fF
C16751 D_INPUT_0 PAND2X1_60/B 0.10fF
C16752 POR2X1_683/CTRL2 POR2X1_236/Y 0.10fF
C16753 POR2X1_78/B PAND2X1_57/B 16.96fF
C16754 POR2X1_143/CTRL POR2X1_236/Y 0.01fF
C16755 PAND2X1_682/CTRL POR2X1_750/B 0.01fF
C16756 POR2X1_67/A POR2X1_93/A 1.98fF
C16757 POR2X1_806/CTRL PAND2X1_69/A 0.01fF
C16758 PAND2X1_76/Y POR2X1_293/Y 0.07fF
C16759 INPUT_1 POR2X1_266/O 0.01fF
C16760 PAND2X1_3/A PAND2X1_1/CTRL 0.01fF
C16761 POR2X1_102/Y PAND2X1_645/B 0.03fF
C16762 POR2X1_346/CTRL PAND2X1_58/A 0.01fF
C16763 POR2X1_334/B PAND2X1_262/O 0.19fF
C16764 POR2X1_422/Y POR2X1_583/O 0.01fF
C16765 PAND2X1_219/A POR2X1_38/Y 1.88fF
C16766 POR2X1_3/A PAND2X1_11/Y 0.12fF
C16767 PAND2X1_568/B PAND2X1_577/Y 0.03fF
C16768 INPUT_1 POR2X1_28/CTRL 0.01fF
C16769 POR2X1_253/CTRL PAND2X1_508/Y 0.00fF
C16770 PAND2X1_93/B POR2X1_703/A 0.07fF
C16771 PAND2X1_23/Y PAND2X1_65/B 0.27fF
C16772 POR2X1_633/A POR2X1_68/B 0.09fF
C16773 PAND2X1_216/CTRL2 INPUT_0 0.01fF
C16774 POR2X1_65/A POR2X1_519/Y 0.12fF
C16775 PAND2X1_468/O PAND2X1_580/B 0.00fF
C16776 POR2X1_355/B POR2X1_244/B 0.03fF
C16777 POR2X1_809/Y POR2X1_812/A 0.01fF
C16778 POR2X1_278/Y POR2X1_498/O 0.05fF
C16779 PAND2X1_478/CTRL PAND2X1_803/A 0.00fF
C16780 PAND2X1_48/B POR2X1_663/O 0.01fF
C16781 POR2X1_786/A VDD 0.19fF
C16782 POR2X1_859/A POR2X1_790/CTRL 0.06fF
C16783 PAND2X1_190/Y PAND2X1_140/a_76_28# 0.06fF
C16784 PAND2X1_250/O POR2X1_778/B 0.03fF
C16785 POR2X1_217/CTRL POR2X1_572/B 0.01fF
C16786 PAND2X1_90/A POR2X1_547/B 0.04fF
C16787 POR2X1_657/O POR2X1_510/Y 0.12fF
C16788 POR2X1_124/B POR2X1_654/B 0.23fF
C16789 POR2X1_356/A POR2X1_570/CTRL2 0.51fF
C16790 POR2X1_13/A POR2X1_669/O 0.01fF
C16791 POR2X1_814/B POR2X1_778/B 0.03fF
C16792 POR2X1_566/A POR2X1_724/m4_208_n4# 0.06fF
C16793 POR2X1_742/CTRL POR2X1_741/Y 0.01fF
C16794 PAND2X1_254/Y PAND2X1_515/O 0.02fF
C16795 PAND2X1_840/B POR2X1_236/Y 0.10fF
C16796 POR2X1_808/A POR2X1_532/A 0.01fF
C16797 POR2X1_596/A POR2X1_750/B 0.03fF
C16798 PAND2X1_42/O D_INPUT_1 0.05fF
C16799 POR2X1_41/B PAND2X1_486/CTRL 0.01fF
C16800 PAND2X1_674/CTRL VDD 0.00fF
C16801 POR2X1_40/Y PAND2X1_168/CTRL2 0.01fF
C16802 PAND2X1_61/Y POR2X1_73/Y 0.03fF
C16803 PAND2X1_20/A POR2X1_854/B 0.05fF
C16804 POR2X1_60/A POR2X1_437/CTRL2 0.02fF
C16805 POR2X1_502/A POR2X1_664/Y 0.04fF
C16806 POR2X1_417/Y PAND2X1_388/Y 0.06fF
C16807 POR2X1_780/O POR2X1_780/A 0.03fF
C16808 PAND2X1_48/B PAND2X1_372/CTRL -0.06fF
C16809 POR2X1_287/B PAND2X1_96/B 0.03fF
C16810 POR2X1_83/B PAND2X1_559/O 0.17fF
C16811 POR2X1_428/O POR2X1_32/A 0.01fF
C16812 POR2X1_13/A PAND2X1_552/B 0.02fF
C16813 PAND2X1_218/O INPUT_0 0.02fF
C16814 POR2X1_465/B POR2X1_554/Y 0.02fF
C16815 PAND2X1_661/B PAND2X1_828/CTRL2 0.01fF
C16816 POR2X1_197/a_56_344# POR2X1_741/Y 0.00fF
C16817 POR2X1_346/B POR2X1_296/B 0.00fF
C16818 D_INPUT_0 POR2X1_571/O 0.01fF
C16819 POR2X1_389/m4_208_n4# POR2X1_480/A 0.08fF
C16820 PAND2X1_857/A PAND2X1_200/a_16_344# 0.02fF
C16821 INPUT_1 POR2X1_225/O 0.02fF
C16822 POR2X1_48/A PAND2X1_156/B 0.01fF
C16823 INPUT_1 POR2X1_585/Y 0.04fF
C16824 POR2X1_502/A POR2X1_775/A 0.04fF
C16825 PAND2X1_449/CTRL POR2X1_77/Y 0.00fF
C16826 POR2X1_717/O POR2X1_475/A 0.07fF
C16827 PAND2X1_55/Y POR2X1_784/A 0.02fF
C16828 POR2X1_650/A POR2X1_493/CTRL2 0.04fF
C16829 POR2X1_220/Y POR2X1_795/B 0.07fF
C16830 POR2X1_289/Y POR2X1_171/Y 0.04fF
C16831 POR2X1_383/A PAND2X1_766/O 0.01fF
C16832 POR2X1_96/A PAND2X1_675/A 0.29fF
C16833 POR2X1_445/O POR2X1_222/Y 0.01fF
C16834 PAND2X1_216/B POR2X1_102/Y 0.03fF
C16835 POR2X1_197/a_16_28# PAND2X1_56/Y 0.13fF
C16836 PAND2X1_73/Y POR2X1_520/B 0.02fF
C16837 PAND2X1_564/CTRL2 POR2X1_73/Y 0.05fF
C16838 POR2X1_130/A POR2X1_804/A 0.05fF
C16839 PAND2X1_23/Y PAND2X1_238/O 0.15fF
C16840 GATE_741 PAND2X1_362/CTRL 0.01fF
C16841 PAND2X1_489/CTRL PAND2X1_557/A 0.01fF
C16842 POR2X1_3/A POR2X1_25/CTRL 0.06fF
C16843 POR2X1_248/O VDD 0.00fF
C16844 PAND2X1_40/O PAND2X1_57/B 0.16fF
C16845 POR2X1_847/B POR2X1_408/Y 0.03fF
C16846 POR2X1_87/B PAND2X1_32/CTRL 0.02fF
C16847 POR2X1_189/Y POR2X1_680/Y 0.02fF
C16848 POR2X1_72/B PAND2X1_569/B 0.09fF
C16849 POR2X1_814/A POR2X1_579/O 0.02fF
C16850 PAND2X1_23/Y POR2X1_638/a_16_28# 0.01fF
C16851 POR2X1_814/B POR2X1_854/B 0.10fF
C16852 POR2X1_41/B POR2X1_56/Y 0.02fF
C16853 POR2X1_566/A POR2X1_804/A 0.34fF
C16854 PAND2X1_90/Y PAND2X1_60/B 0.16fF
C16855 POR2X1_814/B POR2X1_710/B 0.01fF
C16856 PAND2X1_81/B POR2X1_786/A 0.03fF
C16857 POR2X1_547/a_16_28# POR2X1_502/A 0.08fF
C16858 PAND2X1_308/O POR2X1_14/Y 0.15fF
C16859 POR2X1_708/a_16_28# POR2X1_779/A 0.07fF
C16860 POR2X1_60/CTRL POR2X1_13/A 0.01fF
C16861 PAND2X1_61/Y PAND2X1_244/B 0.03fF
C16862 INPUT_0 POR2X1_597/CTRL2 0.02fF
C16863 PAND2X1_837/CTRL2 POR2X1_42/Y 0.01fF
C16864 PAND2X1_308/O PAND2X1_453/A 0.03fF
C16865 POR2X1_97/m4_208_n4# PAND2X1_258/m4_208_n4# 0.13fF
C16866 POR2X1_16/A PAND2X1_731/B 0.01fF
C16867 POR2X1_667/A PAND2X1_560/B 0.03fF
C16868 PAND2X1_322/CTRL PAND2X1_32/B 0.01fF
C16869 PAND2X1_820/CTRL POR2X1_847/B 0.01fF
C16870 PAND2X1_731/CTRL POR2X1_763/Y 0.08fF
C16871 PAND2X1_621/a_16_344# POR2X1_750/B 0.01fF
C16872 POR2X1_455/m4_208_n4# PAND2X1_60/B 0.09fF
C16873 POR2X1_48/A POR2X1_524/CTRL 0.01fF
C16874 PAND2X1_490/CTRL2 POR2X1_334/B 0.05fF
C16875 POR2X1_449/A POR2X1_750/B 0.03fF
C16876 PAND2X1_228/CTRL POR2X1_52/Y 0.01fF
C16877 POR2X1_378/A VDD -0.00fF
C16878 POR2X1_834/Y POR2X1_807/A 0.05fF
C16879 PAND2X1_41/B POR2X1_352/a_76_344# 0.01fF
C16880 PAND2X1_775/CTRL2 POR2X1_91/Y 0.01fF
C16881 POR2X1_358/O PAND2X1_32/B 0.01fF
C16882 POR2X1_335/CTRL POR2X1_337/A 0.04fF
C16883 PAND2X1_390/Y POR2X1_394/A 0.03fF
C16884 POR2X1_57/A POR2X1_290/Y 0.00fF
C16885 POR2X1_155/O POR2X1_162/Y 0.05fF
C16886 POR2X1_700/O POR2X1_700/Y 0.02fF
C16887 POR2X1_532/A POR2X1_149/Y 0.03fF
C16888 POR2X1_101/A POR2X1_814/B 0.02fF
C16889 PAND2X1_658/A PAND2X1_548/CTRL2 0.01fF
C16890 PAND2X1_717/Y PAND2X1_571/Y 0.03fF
C16891 PAND2X1_460/O POR2X1_7/B 0.17fF
C16892 PAND2X1_41/B POR2X1_317/B 0.03fF
C16893 PAND2X1_48/B POR2X1_541/O 0.09fF
C16894 POR2X1_734/A POR2X1_559/A 0.53fF
C16895 POR2X1_570/CTRL2 POR2X1_569/A 0.05fF
C16896 PAND2X1_592/CTRL POR2X1_283/A 0.03fF
C16897 POR2X1_383/A POR2X1_220/Y 0.14fF
C16898 PAND2X1_90/Y POR2X1_353/A 0.05fF
C16899 PAND2X1_65/Y POR2X1_244/Y 0.10fF
C16900 PAND2X1_255/CTRL POR2X1_814/A 0.26fF
C16901 POR2X1_493/CTRL2 POR2X1_294/B 0.10fF
C16902 POR2X1_185/a_16_28# POR2X1_805/A 0.03fF
C16903 POR2X1_62/Y POR2X1_750/A 0.02fF
C16904 VDD POR2X1_310/Y 0.01fF
C16905 PAND2X1_793/Y POR2X1_283/A 0.03fF
C16906 PAND2X1_96/B PAND2X1_316/CTRL2 0.00fF
C16907 POR2X1_326/A POR2X1_186/Y 0.05fF
C16908 POR2X1_41/B POR2X1_235/Y 0.29fF
C16909 VDD POR2X1_308/B 0.00fF
C16910 PAND2X1_96/B POR2X1_61/B 0.01fF
C16911 POR2X1_296/B PAND2X1_304/O 0.24fF
C16912 POR2X1_409/B POR2X1_39/B 0.10fF
C16913 POR2X1_16/A POR2X1_821/CTRL2 0.01fF
C16914 POR2X1_382/O POR2X1_382/Y 0.01fF
C16915 POR2X1_55/Y POR2X1_239/Y 0.99fF
C16916 POR2X1_500/m4_208_n4# POR2X1_318/A 0.08fF
C16917 POR2X1_383/A POR2X1_404/Y 0.03fF
C16918 PAND2X1_338/B POR2X1_42/Y 0.00fF
C16919 POR2X1_480/A POR2X1_590/Y 0.03fF
C16920 POR2X1_333/CTRL2 POR2X1_578/Y 0.03fF
C16921 PAND2X1_738/Y PAND2X1_336/O 0.10fF
C16922 POR2X1_65/A PAND2X1_325/CTRL2 0.03fF
C16923 POR2X1_622/O POR2X1_622/B 0.04fF
C16924 POR2X1_255/Y POR2X1_73/Y 0.02fF
C16925 PAND2X1_73/Y POR2X1_561/B 0.32fF
C16926 POR2X1_115/a_16_28# POR2X1_366/A 0.03fF
C16927 POR2X1_343/Y POR2X1_218/Y 0.10fF
C16928 POR2X1_549/O POR2X1_266/A 0.01fF
C16929 POR2X1_38/Y POR2X1_816/A 0.04fF
C16930 POR2X1_398/Y POR2X1_294/A 0.05fF
C16931 POR2X1_60/O PAND2X1_651/Y 0.02fF
C16932 POR2X1_566/A PAND2X1_313/O 0.17fF
C16933 POR2X1_809/A PAND2X1_65/B 0.02fF
C16934 PAND2X1_522/CTRL INPUT_0 0.33fF
C16935 POR2X1_8/Y POR2X1_88/Y 0.12fF
C16936 POR2X1_71/Y PAND2X1_574/O 0.06fF
C16937 POR2X1_804/A POR2X1_573/A 0.05fF
C16938 PAND2X1_403/O POR2X1_411/B 0.02fF
C16939 PAND2X1_388/Y POR2X1_184/Y 1.84fF
C16940 POR2X1_136/Y POR2X1_43/B 0.03fF
C16941 POR2X1_346/CTRL PAND2X1_96/B 0.01fF
C16942 POR2X1_41/B PAND2X1_374/a_76_28# 0.02fF
C16943 POR2X1_860/A POR2X1_362/O 0.02fF
C16944 PAND2X1_57/B PAND2X1_142/CTRL2 0.01fF
C16945 PAND2X1_469/B POR2X1_7/A 0.21fF
C16946 POR2X1_590/A PAND2X1_56/A -0.00fF
C16947 POR2X1_144/a_16_28# POR2X1_376/B 0.01fF
C16948 POR2X1_3/A POR2X1_700/Y 0.16fF
C16949 D_GATE_222 POR2X1_566/B 0.10fF
C16950 PAND2X1_721/B POR2X1_77/Y 0.00fF
C16951 POR2X1_87/CTRL POR2X1_590/A 0.05fF
C16952 D_INPUT_0 POR2X1_716/a_16_28# 0.00fF
C16953 PAND2X1_480/B POR2X1_129/Y 0.05fF
C16954 PAND2X1_864/B PAND2X1_864/a_16_344# 0.02fF
C16955 POR2X1_608/CTRL2 POR2X1_294/A 0.08fF
C16956 PAND2X1_447/CTRL POR2X1_329/A 0.03fF
C16957 PAND2X1_48/B POR2X1_675/Y 0.03fF
C16958 POR2X1_5/CTRL VDD 0.00fF
C16959 POR2X1_276/A POR2X1_140/A 0.03fF
C16960 POR2X1_447/B PAND2X1_627/CTRL2 0.04fF
C16961 PAND2X1_651/Y PAND2X1_549/B 0.03fF
C16962 PAND2X1_148/O PAND2X1_209/A 0.03fF
C16963 POR2X1_754/A POR2X1_129/Y 0.01fF
C16964 PAND2X1_201/CTRL PAND2X1_206/B 0.00fF
C16965 POR2X1_741/Y POR2X1_787/O 0.01fF
C16966 PAND2X1_6/Y PAND2X1_373/O 0.01fF
C16967 INPUT_1 PAND2X1_401/O 0.04fF
C16968 POR2X1_137/Y POR2X1_216/O 0.00fF
C16969 POR2X1_722/B POR2X1_722/A 0.02fF
C16970 PAND2X1_48/B POR2X1_544/B 0.07fF
C16971 POR2X1_325/A POR2X1_374/CTRL2 0.01fF
C16972 POR2X1_732/CTRL2 POR2X1_353/A 0.01fF
C16973 PAND2X1_57/B POR2X1_294/A 4.18fF
C16974 PAND2X1_775/CTRL2 POR2X1_109/Y 0.03fF
C16975 POR2X1_707/a_16_28# PAND2X1_95/B 0.01fF
C16976 PAND2X1_659/Y PAND2X1_480/B 0.03fF
C16977 PAND2X1_658/A PAND2X1_861/a_56_28# 0.00fF
C16978 POR2X1_722/A POR2X1_294/B 0.09fF
C16979 POR2X1_383/A PAND2X1_824/CTRL2 0.01fF
C16980 PAND2X1_71/Y POR2X1_404/Y 0.03fF
C16981 PAND2X1_797/Y PAND2X1_209/CTRL 0.01fF
C16982 PAND2X1_7/O POR2X1_259/B 0.03fF
C16983 INPUT_1 POR2X1_816/A 0.03fF
C16984 POR2X1_532/A POR2X1_769/Y 0.03fF
C16985 INPUT_1 D_INPUT_1 2.29fF
C16986 PAND2X1_651/a_16_344# POR2X1_43/B 0.01fF
C16987 PAND2X1_105/O PAND2X1_348/A 0.08fF
C16988 PAND2X1_780/O POR2X1_744/Y 0.00fF
C16989 POR2X1_162/Y PAND2X1_158/CTRL2 0.01fF
C16990 POR2X1_416/B PAND2X1_540/a_16_344# 0.02fF
C16991 PAND2X1_572/O PAND2X1_723/A 0.00fF
C16992 POR2X1_226/Y POR2X1_77/Y 0.03fF
C16993 POR2X1_72/B PAND2X1_327/a_56_28# 0.00fF
C16994 PAND2X1_311/CTRL POR2X1_260/A 0.01fF
C16995 PAND2X1_808/Y PAND2X1_359/Y 0.00fF
C16996 PAND2X1_372/a_76_28# PAND2X1_48/A 0.02fF
C16997 POR2X1_816/A POR2X1_153/Y 0.03fF
C16998 POR2X1_569/A POR2X1_366/A 0.07fF
C16999 POR2X1_272/Y POR2X1_39/B 0.03fF
C17000 POR2X1_669/B PAND2X1_147/O 0.03fF
C17001 POR2X1_119/Y PAND2X1_724/B 0.03fF
C17002 POR2X1_7/B PAND2X1_643/A 0.09fF
C17003 POR2X1_384/A POR2X1_816/A 0.01fF
C17004 POR2X1_714/CTRL2 POR2X1_703/Y 0.01fF
C17005 POR2X1_661/A POR2X1_590/A 0.07fF
C17006 POR2X1_65/Y PAND2X1_201/CTRL 0.00fF
C17007 PAND2X1_79/CTRL POR2X1_571/Y 0.01fF
C17008 POR2X1_651/Y POR2X1_121/B 0.07fF
C17009 POR2X1_366/CTRL POR2X1_383/A 0.01fF
C17010 POR2X1_537/Y PAND2X1_536/CTRL 0.01fF
C17011 POR2X1_467/Y POR2X1_535/CTRL 0.01fF
C17012 POR2X1_176/CTRL2 POR2X1_90/Y 0.01fF
C17013 POR2X1_614/A POR2X1_737/A 0.03fF
C17014 POR2X1_332/Y POR2X1_341/a_16_28# 0.03fF
C17015 POR2X1_712/a_16_28# POR2X1_260/A 0.02fF
C17016 POR2X1_110/Y PAND2X1_464/Y 0.03fF
C17017 POR2X1_653/a_16_28# POR2X1_711/Y 0.06fF
C17018 PAND2X1_765/CTRL2 POR2X1_260/A 0.03fF
C17019 POR2X1_7/B PAND2X1_346/a_16_344# 0.02fF
C17020 PAND2X1_69/A PAND2X1_48/A 0.07fF
C17021 POR2X1_394/A POR2X1_757/CTRL2 0.13fF
C17022 POR2X1_8/Y POR2X1_384/CTRL 0.01fF
C17023 POR2X1_567/B PAND2X1_52/O 0.15fF
C17024 POR2X1_110/Y PAND2X1_565/A 0.02fF
C17025 POR2X1_833/A PAND2X1_63/B 0.07fF
C17026 POR2X1_262/Y PAND2X1_560/a_56_28# 0.00fF
C17027 PAND2X1_810/A PAND2X1_221/Y 0.05fF
C17028 POR2X1_264/Y PAND2X1_517/O 0.03fF
C17029 POR2X1_327/Y POR2X1_228/Y 0.03fF
C17030 PAND2X1_206/B D_INPUT_0 0.23fF
C17031 PAND2X1_357/Y PAND2X1_352/B 0.02fF
C17032 POR2X1_103/CTRL PAND2X1_349/A 0.01fF
C17033 POR2X1_532/A PAND2X1_692/CTRL 0.01fF
C17034 POR2X1_704/O POR2X1_317/B 0.17fF
C17035 POR2X1_616/Y POR2X1_93/A 0.01fF
C17036 POR2X1_136/Y POR2X1_183/CTRL 0.00fF
C17037 PAND2X1_856/B PAND2X1_856/O 0.05fF
C17038 POR2X1_152/CTRL2 POR2X1_39/B 0.12fF
C17039 POR2X1_43/Y POR2X1_46/Y 0.00fF
C17040 POR2X1_518/O POR2X1_73/Y 0.04fF
C17041 POR2X1_415/A PAND2X1_66/O 0.17fF
C17042 POR2X1_646/B POR2X1_606/Y 0.03fF
C17043 POR2X1_407/A POR2X1_779/CTRL 0.01fF
C17044 POR2X1_730/Y POR2X1_186/B 0.00fF
C17045 PAND2X1_129/CTRL2 POR2X1_68/B 0.01fF
C17046 PAND2X1_352/A POR2X1_20/B 0.01fF
C17047 POR2X1_99/B POR2X1_510/Y 0.03fF
C17048 POR2X1_234/A PAND2X1_520/CTRL 0.01fF
C17049 POR2X1_8/Y POR2X1_749/CTRL2 0.00fF
C17050 POR2X1_93/O POR2X1_39/B 0.02fF
C17051 POR2X1_557/A PAND2X1_71/Y 0.03fF
C17052 POR2X1_65/Y D_INPUT_0 0.01fF
C17053 POR2X1_790/B PAND2X1_52/B 0.03fF
C17054 PAND2X1_184/O PAND2X1_71/Y 0.04fF
C17055 PAND2X1_659/Y POR2X1_7/O 0.01fF
C17056 POR2X1_624/Y POR2X1_218/Y 0.18fF
C17057 POR2X1_20/B PAND2X1_58/A 0.05fF
C17058 PAND2X1_802/O PAND2X1_539/Y 0.02fF
C17059 PAND2X1_73/Y PAND2X1_39/B 0.09fF
C17060 POR2X1_459/Y POR2X1_750/B 0.01fF
C17061 POR2X1_863/A POR2X1_740/Y 0.03fF
C17062 POR2X1_1/CTRL2 D_INPUT_4 0.05fF
C17063 POR2X1_457/Y VDD 0.10fF
C17064 PAND2X1_803/Y POR2X1_77/Y 0.02fF
C17065 POR2X1_311/Y PAND2X1_222/CTRL 0.01fF
C17066 PAND2X1_91/O POR2X1_97/A 0.05fF
C17067 POR2X1_527/a_16_28# POR2X1_110/Y -0.00fF
C17068 POR2X1_316/a_16_28# POR2X1_153/Y 0.00fF
C17069 PAND2X1_613/CTRL POR2X1_296/B 0.01fF
C17070 POR2X1_834/CTRL POR2X1_260/B 0.01fF
C17071 POR2X1_678/A POR2X1_678/O 0.01fF
C17072 POR2X1_323/CTRL2 POR2X1_485/Y 0.01fF
C17073 POR2X1_68/B POR2X1_717/B 0.03fF
C17074 PAND2X1_429/Y D_INPUT_7 0.03fF
C17075 POR2X1_48/A POR2X1_409/B 1.35fF
C17076 PAND2X1_63/CTRL POR2X1_66/A 0.22fF
C17077 POR2X1_65/A POR2X1_485/Y 0.00fF
C17078 POR2X1_610/O POR2X1_590/A 0.02fF
C17079 POR2X1_532/A POR2X1_568/A 0.06fF
C17080 PAND2X1_497/CTRL POR2X1_590/A 0.04fF
C17081 PAND2X1_85/O POR2X1_243/Y 0.07fF
C17082 POR2X1_85/Y POR2X1_235/Y 0.17fF
C17083 POR2X1_648/Y PAND2X1_511/O 0.05fF
C17084 POR2X1_65/A PAND2X1_838/CTRL 0.01fF
C17085 POR2X1_590/Y PAND2X1_304/O 0.05fF
C17086 PAND2X1_864/B POR2X1_282/O 0.02fF
C17087 PAND2X1_20/A POR2X1_862/A 0.07fF
C17088 POR2X1_623/CTRL POR2X1_296/B 0.01fF
C17089 POR2X1_532/A PAND2X1_146/CTRL2 0.02fF
C17090 PAND2X1_206/A POR2X1_40/Y 0.00fF
C17091 POR2X1_234/A POR2X1_234/a_16_28# 0.03fF
C17092 POR2X1_567/A POR2X1_652/A 0.00fF
C17093 PAND2X1_72/A POR2X1_366/A 0.03fF
C17094 POR2X1_808/A POR2X1_808/CTRL2 0.05fF
C17095 POR2X1_296/CTRL VDD 0.00fF
C17096 POR2X1_60/A PAND2X1_205/A 0.03fF
C17097 PAND2X1_629/O POR2X1_628/Y 0.00fF
C17098 PAND2X1_86/CTRL2 POR2X1_404/Y 0.14fF
C17099 PAND2X1_373/CTRL PAND2X1_72/A 0.01fF
C17100 POR2X1_202/A POR2X1_202/O 0.07fF
C17101 POR2X1_257/A PAND2X1_803/A 0.07fF
C17102 POR2X1_257/A POR2X1_677/a_16_28# 0.03fF
C17103 PAND2X1_23/Y POR2X1_814/A 0.24fF
C17104 POR2X1_174/CTRL2 PAND2X1_72/A 0.09fF
C17105 POR2X1_709/A POR2X1_410/CTRL2 0.01fF
C17106 PAND2X1_23/Y PAND2X1_75/CTRL 0.01fF
C17107 POR2X1_337/Y PAND2X1_179/CTRL 0.05fF
C17108 POR2X1_431/O POR2X1_55/Y 0.01fF
C17109 PAND2X1_796/B POR2X1_236/Y 0.02fF
C17110 PAND2X1_221/Y PAND2X1_739/B 0.12fF
C17111 PAND2X1_73/Y POR2X1_805/Y 0.03fF
C17112 PAND2X1_454/B POR2X1_236/Y 0.88fF
C17113 PAND2X1_689/CTRL POR2X1_812/A 0.11fF
C17114 POR2X1_20/B POR2X1_233/CTRL2 0.02fF
C17115 POR2X1_672/Y POR2X1_5/Y 0.01fF
C17116 PAND2X1_448/a_76_28# POR2X1_421/Y 0.02fF
C17117 POR2X1_13/A PAND2X1_98/CTRL 0.01fF
C17118 POR2X1_555/O POR2X1_186/B 0.01fF
C17119 PAND2X1_20/A PAND2X1_73/Y 1.27fF
C17120 POR2X1_335/a_16_28# POR2X1_556/A 0.03fF
C17121 PAND2X1_862/B PAND2X1_203/CTRL 0.00fF
C17122 PAND2X1_246/m4_208_n4# POR2X1_404/Y 0.08fF
C17123 D_INPUT_0 POR2X1_750/B 0.03fF
C17124 POR2X1_849/A POR2X1_94/A 0.09fF
C17125 PAND2X1_45/CTRL POR2X1_741/Y 0.00fF
C17126 PAND2X1_33/O POR2X1_7/B 0.01fF
C17127 POR2X1_853/A POR2X1_465/O 0.00fF
C17128 POR2X1_467/Y POR2X1_448/CTRL2 0.01fF
C17129 PAND2X1_124/Y POR2X1_5/Y 0.03fF
C17130 POR2X1_35/a_16_28# POR2X1_34/Y -0.00fF
C17131 POR2X1_67/Y POR2X1_90/Y 0.03fF
C17132 POR2X1_540/Y POR2X1_632/Y 0.23fF
C17133 PAND2X1_96/B POR2X1_630/B 0.02fF
C17134 POR2X1_260/B PAND2X1_131/CTRL 0.01fF
C17135 POR2X1_416/Y PAND2X1_634/CTRL2 0.01fF
C17136 POR2X1_383/A POR2X1_655/CTRL 0.09fF
C17137 POR2X1_462/B POR2X1_462/O 0.01fF
C17138 POR2X1_23/Y POR2X1_236/Y 0.21fF
C17139 POR2X1_261/Y PAND2X1_555/A 0.00fF
C17140 POR2X1_466/Y POR2X1_467/Y 0.02fF
C17141 PAND2X1_251/CTRL VDD 0.00fF
C17142 PAND2X1_545/CTRL2 POR2X1_40/Y 0.01fF
C17143 POR2X1_174/B POR2X1_175/A 0.04fF
C17144 POR2X1_807/CTRL POR2X1_480/A 0.03fF
C17145 PAND2X1_9/CTRL POR2X1_94/A 0.07fF
C17146 POR2X1_48/A POR2X1_272/Y 0.11fF
C17147 POR2X1_355/B POR2X1_319/A 0.03fF
C17148 PAND2X1_205/O PAND2X1_735/Y 0.05fF
C17149 POR2X1_549/CTRL2 POR2X1_78/A 0.03fF
C17150 PAND2X1_307/CTRL2 POR2X1_40/Y 0.04fF
C17151 PAND2X1_798/a_76_28# PAND2X1_354/A 0.01fF
C17152 POR2X1_814/B PAND2X1_73/Y 0.28fF
C17153 POR2X1_636/B VDD 0.00fF
C17154 PAND2X1_865/Y POR2X1_416/B 0.07fF
C17155 PAND2X1_557/A PAND2X1_742/O 0.08fF
C17156 POR2X1_804/CTRL VDD 0.00fF
C17157 POR2X1_78/A PAND2X1_42/O 0.02fF
C17158 POR2X1_555/A POR2X1_555/B 0.00fF
C17159 PAND2X1_722/O POR2X1_666/A 0.17fF
C17160 PAND2X1_474/O POR2X1_43/B 0.05fF
C17161 POR2X1_329/A POR2X1_387/Y 0.07fF
C17162 POR2X1_72/B PAND2X1_784/A 0.01fF
C17163 POR2X1_27/CTRL2 PAND2X1_63/B 0.01fF
C17164 POR2X1_812/A POR2X1_800/m4_208_n4# 0.15fF
C17165 INPUT_2 PAND2X1_618/O 0.03fF
C17166 POR2X1_499/A POR2X1_576/Y 0.55fF
C17167 PAND2X1_23/Y POR2X1_444/B 0.02fF
C17168 PAND2X1_838/B POR2X1_43/B 0.00fF
C17169 PAND2X1_39/B POR2X1_249/CTRL2 0.01fF
C17170 POR2X1_422/CTRL POR2X1_293/Y 0.05fF
C17171 POR2X1_83/B POR2X1_5/Y 0.08fF
C17172 POR2X1_683/Y POR2X1_604/O 0.00fF
C17173 POR2X1_416/B PAND2X1_346/O 0.02fF
C17174 POR2X1_614/A PAND2X1_761/CTRL 0.01fF
C17175 PAND2X1_73/Y POR2X1_325/A 0.01fF
C17176 POR2X1_68/A POR2X1_624/Y 0.10fF
C17177 POR2X1_60/A PAND2X1_76/Y 0.06fF
C17178 POR2X1_814/A POR2X1_520/A 0.03fF
C17179 POR2X1_696/O POR2X1_376/B 0.01fF
C17180 POR2X1_586/Y VDD 0.19fF
C17181 POR2X1_754/A POR2X1_37/Y 0.00fF
C17182 PAND2X1_39/B POR2X1_784/CTRL2 0.11fF
C17183 POR2X1_78/B PAND2X1_420/CTRL 0.13fF
C17184 POR2X1_276/CTRL2 POR2X1_218/Y 0.09fF
C17185 INPUT_3 POR2X1_38/Y 0.09fF
C17186 PAND2X1_94/O PAND2X1_55/Y 0.02fF
C17187 PAND2X1_106/CTRL2 POR2X1_116/A 0.00fF
C17188 PAND2X1_106/O POR2X1_554/B 0.01fF
C17189 PAND2X1_210/CTRL2 PAND2X1_725/Y 0.00fF
C17190 POR2X1_66/B POR2X1_403/Y 0.00fF
C17191 POR2X1_149/B POR2X1_260/B 0.04fF
C17192 PAND2X1_463/O POR2X1_5/Y 0.08fF
C17193 PAND2X1_90/Y POR2X1_750/B 0.09fF
C17194 PAND2X1_220/Y PAND2X1_540/a_56_28# 0.00fF
C17195 POR2X1_708/O POR2X1_121/B 0.02fF
C17196 POR2X1_96/A POR2X1_498/Y 0.02fF
C17197 PAND2X1_255/O POR2X1_186/B 0.02fF
C17198 POR2X1_760/A PAND2X1_537/CTRL2 0.03fF
C17199 POR2X1_49/Y PAND2X1_803/A 0.05fF
C17200 PAND2X1_616/CTRL2 VDD -0.00fF
C17201 POR2X1_471/a_16_28# POR2X1_78/A 0.01fF
C17202 PAND2X1_594/CTRL2 POR2X1_740/Y 0.00fF
C17203 POR2X1_450/B VDD 0.22fF
C17204 POR2X1_262/Y POR2X1_7/A 0.06fF
C17205 POR2X1_674/O PAND2X1_652/A 0.14fF
C17206 POR2X1_388/CTRL2 PAND2X1_93/B 0.09fF
C17207 PAND2X1_489/a_76_28# POR2X1_488/Y 0.04fF
C17208 POR2X1_96/A PAND2X1_772/O 0.05fF
C17209 POR2X1_480/A POR2X1_186/Y 0.10fF
C17210 POR2X1_188/A POR2X1_733/a_56_344# 0.00fF
C17211 POR2X1_72/B PAND2X1_501/B 0.16fF
C17212 POR2X1_378/A PAND2X1_9/Y 0.00fF
C17213 POR2X1_52/A POR2X1_497/CTRL2 0.00fF
C17214 POR2X1_312/Y POR2X1_236/Y 0.00fF
C17215 PAND2X1_95/B PAND2X1_752/CTRL 0.01fF
C17216 POR2X1_624/B POR2X1_260/A 0.03fF
C17217 POR2X1_260/B POR2X1_644/A 0.31fF
C17218 POR2X1_66/B POR2X1_502/A 0.23fF
C17219 POR2X1_13/A POR2X1_748/A 0.01fF
C17220 POR2X1_423/Y VDD 0.46fF
C17221 POR2X1_786/A POR2X1_267/A 0.04fF
C17222 POR2X1_23/Y POR2X1_229/CTRL 0.01fF
C17223 PAND2X1_863/CTRL VDD 0.00fF
C17224 POR2X1_188/A POR2X1_502/A 0.06fF
C17225 PAND2X1_48/B POR2X1_14/Y 0.03fF
C17226 POR2X1_609/Y POR2X1_234/CTRL 0.00fF
C17227 POR2X1_442/Y PAND2X1_724/B 0.00fF
C17228 POR2X1_809/A POR2X1_814/A 0.05fF
C17229 PAND2X1_93/B POR2X1_140/O 0.01fF
C17230 POR2X1_446/B POR2X1_222/A 0.03fF
C17231 POR2X1_102/Y PAND2X1_717/CTRL 0.01fF
C17232 POR2X1_505/CTRL POR2X1_20/B 0.01fF
C17233 POR2X1_496/Y PAND2X1_6/A 0.09fF
C17234 POR2X1_719/CTRL2 PAND2X1_93/B 0.02fF
C17235 POR2X1_687/A POR2X1_452/Y 1.66fF
C17236 POR2X1_78/B PAND2X1_85/Y 0.20fF
C17237 POR2X1_196/a_16_28# POR2X1_205/Y 0.03fF
C17238 POR2X1_41/B PAND2X1_361/a_76_28# 0.02fF
C17239 POR2X1_311/Y PAND2X1_675/A 0.03fF
C17240 INPUT_1 INPUT_3 0.20fF
C17241 PAND2X1_854/a_56_28# POR2X1_102/Y 0.00fF
C17242 PAND2X1_73/Y PAND2X1_519/a_16_344# 0.06fF
C17243 POR2X1_197/Y PAND2X1_93/B 0.02fF
C17244 POR2X1_114/B POR2X1_121/B 0.03fF
C17245 POR2X1_509/A PAND2X1_20/A 0.01fF
C17246 POR2X1_855/B POR2X1_808/a_56_344# 0.00fF
C17247 POR2X1_834/CTRL POR2X1_407/Y 0.01fF
C17248 POR2X1_567/B POR2X1_190/a_76_344# 0.03fF
C17249 POR2X1_697/Y POR2X1_40/Y 2.63fF
C17250 POR2X1_356/A POR2X1_509/B 0.13fF
C17251 POR2X1_615/O POR2X1_754/A 0.01fF
C17252 POR2X1_260/B POR2X1_274/B 0.01fF
C17253 POR2X1_614/Y PAND2X1_69/A 0.01fF
C17254 POR2X1_383/A POR2X1_841/B 0.07fF
C17255 POR2X1_102/Y POR2X1_234/O 0.01fF
C17256 POR2X1_60/A PAND2X1_566/Y 0.05fF
C17257 POR2X1_52/A POR2X1_238/CTRL2 0.01fF
C17258 PAND2X1_844/O POR2X1_20/B 0.04fF
C17259 PAND2X1_674/CTRL2 POR2X1_186/Y 0.03fF
C17260 POR2X1_802/O PAND2X1_93/B 0.01fF
C17261 POR2X1_47/m4_208_n4# POR2X1_748/A 0.12fF
C17262 PAND2X1_23/Y POR2X1_852/B 0.10fF
C17263 PAND2X1_272/CTRL2 PAND2X1_60/B 0.03fF
C17264 POR2X1_225/a_16_28# POR2X1_90/Y 0.03fF
C17265 PAND2X1_34/a_16_344# POR2X1_38/Y 0.01fF
C17266 PAND2X1_23/Y PAND2X1_55/CTRL2 0.00fF
C17267 POR2X1_130/A PAND2X1_755/CTRL 0.05fF
C17268 PAND2X1_48/B POR2X1_791/Y 0.03fF
C17269 POR2X1_660/A POR2X1_733/A 0.07fF
C17270 POR2X1_223/CTRL VDD -0.00fF
C17271 PAND2X1_818/a_76_28# POR2X1_5/Y 0.01fF
C17272 POR2X1_54/Y PAND2X1_749/O 0.13fF
C17273 PAND2X1_357/Y POR2X1_40/Y 0.06fF
C17274 POR2X1_54/Y PAND2X1_522/O 0.23fF
C17275 PAND2X1_48/B POR2X1_637/B 0.03fF
C17276 POR2X1_775/A PAND2X1_229/CTRL 0.01fF
C17277 POR2X1_322/a_16_28# POR2X1_40/Y 0.01fF
C17278 PAND2X1_593/CTRL2 PAND2X1_364/B 0.06fF
C17279 PAND2X1_625/O POR2X1_852/B 0.08fF
C17280 POR2X1_495/Y POR2X1_376/B 0.15fF
C17281 POR2X1_235/CTRL2 POR2X1_32/A 0.01fF
C17282 PAND2X1_219/A POR2X1_591/Y 3.03fF
C17283 PAND2X1_433/CTRL PAND2X1_65/B 0.01fF
C17284 POR2X1_441/Y POR2X1_373/CTRL 0.01fF
C17285 POR2X1_614/A POR2X1_302/B 0.03fF
C17286 POR2X1_502/A POR2X1_859/A 0.07fF
C17287 POR2X1_605/B POR2X1_605/A 0.12fF
C17288 POR2X1_334/B PAND2X1_65/B 0.07fF
C17289 POR2X1_2/a_16_28# INPUT_5 0.03fF
C17290 POR2X1_679/Y PAND2X1_853/B 0.06fF
C17291 PAND2X1_798/B PAND2X1_363/Y 0.02fF
C17292 POR2X1_16/A PAND2X1_489/O 0.37fF
C17293 PAND2X1_483/CTRL POR2X1_48/A 0.01fF
C17294 POR2X1_322/m4_208_n4# POR2X1_49/Y 0.15fF
C17295 POR2X1_130/A PAND2X1_372/a_16_344# 0.02fF
C17296 POR2X1_655/Y POR2X1_784/CTRL 0.12fF
C17297 PAND2X1_650/A POR2X1_409/B 0.02fF
C17298 POR2X1_812/B POR2X1_636/a_16_28# 0.00fF
C17299 POR2X1_423/O POR2X1_7/A 0.07fF
C17300 POR2X1_814/A POR2X1_711/Y 0.10fF
C17301 PAND2X1_480/B POR2X1_293/Y 0.05fF
C17302 POR2X1_367/a_16_28# POR2X1_365/Y -0.00fF
C17303 POR2X1_49/Y POR2X1_583/CTRL2 0.02fF
C17304 POR2X1_294/O POR2X1_294/A 0.10fF
C17305 POR2X1_490/Y PAND2X1_557/O 0.00fF
C17306 POR2X1_494/O POR2X1_5/Y 0.06fF
C17307 PAND2X1_319/a_76_28# PAND2X1_317/Y 0.01fF
C17308 POR2X1_623/A POR2X1_623/B 0.01fF
C17309 POR2X1_57/Y VDD 0.00fF
C17310 POR2X1_652/CTRL PAND2X1_90/Y 0.13fF
C17311 POR2X1_330/Y PAND2X1_163/CTRL2 0.03fF
C17312 POR2X1_102/CTRL POR2X1_411/B 0.01fF
C17313 PAND2X1_23/Y POR2X1_401/B 0.33fF
C17314 POR2X1_271/A POR2X1_23/Y 2.10fF
C17315 POR2X1_848/CTRL PAND2X1_52/B 0.00fF
C17316 POR2X1_754/A POR2X1_293/Y 0.03fF
C17317 POR2X1_46/Y POR2X1_763/Y 0.20fF
C17318 PAND2X1_809/A PAND2X1_863/B 0.01fF
C17319 POR2X1_124/B PAND2X1_65/B 0.03fF
C17320 POR2X1_355/B PAND2X1_48/B 0.03fF
C17321 POR2X1_66/A POR2X1_546/a_56_344# 0.00fF
C17322 PAND2X1_205/Y PAND2X1_186/a_16_344# 0.01fF
C17323 POR2X1_486/B POR2X1_705/B 0.09fF
C17324 VDD POR2X1_587/O -0.00fF
C17325 POR2X1_315/Y POR2X1_60/A 0.10fF
C17326 D_INPUT_5 PAND2X1_2/a_56_28# 0.00fF
C17327 PAND2X1_115/Y PAND2X1_114/Y 0.06fF
C17328 POR2X1_814/A POR2X1_728/A 0.02fF
C17329 POR2X1_861/A POR2X1_624/Y 0.17fF
C17330 PAND2X1_793/Y POR2X1_55/Y 0.04fF
C17331 POR2X1_41/B POR2X1_42/Y 0.18fF
C17332 POR2X1_777/B PAND2X1_150/m4_208_n4# 0.15fF
C17333 POR2X1_515/O PAND2X1_6/Y 0.03fF
C17334 PAND2X1_95/a_16_344# PAND2X1_57/B 0.04fF
C17335 POR2X1_409/a_76_344# POR2X1_5/Y 0.01fF
C17336 INPUT_1 POR2X1_78/A 0.04fF
C17337 PAND2X1_297/O POR2X1_296/Y 0.00fF
C17338 POR2X1_528/Y POR2X1_40/Y 0.49fF
C17339 POR2X1_658/O POR2X1_632/Y 0.01fF
C17340 PAND2X1_391/O POR2X1_751/Y 0.02fF
C17341 PAND2X1_472/CTRL2 POR2X1_60/A 0.03fF
C17342 POR2X1_536/a_56_344# POR2X1_102/Y 0.01fF
C17343 POR2X1_778/B VDD 0.09fF
C17344 POR2X1_753/Y POR2X1_753/CTRL 0.02fF
C17345 POR2X1_48/A PAND2X1_703/O 0.03fF
C17346 POR2X1_199/O POR2X1_741/Y 0.59fF
C17347 POR2X1_296/B POR2X1_507/A 0.09fF
C17348 PAND2X1_73/Y POR2X1_598/a_16_28# 0.03fF
C17349 POR2X1_94/CTRL POR2X1_7/B 0.01fF
C17350 PAND2X1_398/CTRL POR2X1_293/Y 0.01fF
C17351 PAND2X1_23/Y POR2X1_260/Y 0.03fF
C17352 POR2X1_153/a_16_28# POR2X1_37/Y 0.07fF
C17353 POR2X1_186/Y POR2X1_727/O 0.02fF
C17354 POR2X1_41/B POR2X1_309/Y 0.01fF
C17355 POR2X1_549/A PAND2X1_90/A 0.01fF
C17356 POR2X1_433/CTRL2 POR2X1_153/Y 0.05fF
C17357 PAND2X1_90/Y POR2X1_704/CTRL 0.01fF
C17358 PAND2X1_319/B VDD 0.01fF
C17359 PAND2X1_821/O PAND2X1_23/Y 0.03fF
C17360 POR2X1_167/O PAND2X1_714/A 0.36fF
C17361 POR2X1_68/A POR2X1_785/A 0.03fF
C17362 POR2X1_693/CTRL POR2X1_73/Y 0.01fF
C17363 POR2X1_83/B PAND2X1_337/O 0.01fF
C17364 POR2X1_346/B POR2X1_186/Y 0.01fF
C17365 POR2X1_78/A POR2X1_768/Y 0.01fF
C17366 POR2X1_383/A POR2X1_307/B 0.01fF
C17367 POR2X1_529/a_76_344# POR2X1_55/Y 0.03fF
C17368 POR2X1_46/Y POR2X1_73/Y 0.23fF
C17369 POR2X1_447/B POR2X1_629/a_16_28# 0.05fF
C17370 POR2X1_687/Y VDD 0.11fF
C17371 POR2X1_460/A INPUT_4 0.05fF
C17372 POR2X1_51/B POR2X1_44/a_16_28# 0.05fF
C17373 PAND2X1_488/O POR2X1_260/A 0.04fF
C17374 POR2X1_618/CTRL2 POR2X1_382/Y 0.01fF
C17375 POR2X1_16/A POR2X1_39/O 0.15fF
C17376 VDD POR2X1_854/B 6.52fF
C17377 PAND2X1_849/B PAND2X1_849/a_16_344# 0.03fF
C17378 POR2X1_710/B VDD 0.24fF
C17379 POR2X1_307/B POR2X1_590/a_16_28# 0.03fF
C17380 POR2X1_362/B POR2X1_362/A 0.02fF
C17381 PAND2X1_90/Y POR2X1_721/CTRL2 0.05fF
C17382 POR2X1_246/CTRL2 POR2X1_90/Y 0.01fF
C17383 POR2X1_220/CTRL2 PAND2X1_52/B 0.01fF
C17384 POR2X1_712/A PAND2X1_697/CTRL2 0.01fF
C17385 POR2X1_264/Y PAND2X1_96/B 0.03fF
C17386 POR2X1_123/B POR2X1_123/O 0.11fF
C17387 PAND2X1_117/m4_208_n4# POR2X1_123/m4_208_n4# 0.13fF
C17388 POR2X1_754/A POR2X1_408/Y 0.03fF
C17389 POR2X1_590/A POR2X1_362/a_56_344# 0.00fF
C17390 PAND2X1_824/B POR2X1_193/Y 0.07fF
C17391 POR2X1_785/CTRL2 POR2X1_566/B 0.09fF
C17392 POR2X1_643/Y PAND2X1_52/B 0.05fF
C17393 PAND2X1_170/a_56_28# PAND2X1_168/Y 0.00fF
C17394 PAND2X1_57/B POR2X1_710/Y 0.01fF
C17395 POR2X1_56/Y POR2X1_52/Y 0.01fF
C17396 POR2X1_718/a_16_28# POR2X1_834/Y 0.08fF
C17397 POR2X1_360/A POR2X1_101/CTRL 0.03fF
C17398 PAND2X1_433/CTRL2 POR2X1_832/A 0.09fF
C17399 POR2X1_228/O PAND2X1_7/Y 0.01fF
C17400 POR2X1_228/CTRL2 PAND2X1_52/Y 0.01fF
C17401 POR2X1_624/Y POR2X1_138/A 0.04fF
C17402 POR2X1_825/Y POR2X1_20/B 0.04fF
C17403 POR2X1_278/Y PAND2X1_737/B 0.25fF
C17404 PAND2X1_228/CTRL2 PAND2X1_656/A 0.01fF
C17405 PAND2X1_703/a_16_344# POR2X1_312/Y 0.02fF
C17406 POR2X1_778/B PAND2X1_32/B 0.01fF
C17407 PAND2X1_860/A POR2X1_411/B 0.03fF
C17408 POR2X1_52/A PAND2X1_723/A 0.03fF
C17409 POR2X1_66/A PAND2X1_56/A 0.04fF
C17410 POR2X1_858/A POR2X1_590/A 0.01fF
C17411 POR2X1_558/A POR2X1_264/Y 0.01fF
C17412 POR2X1_297/a_16_28# PAND2X1_359/Y 0.03fF
C17413 PAND2X1_562/a_16_344# PAND2X1_555/Y 0.02fF
C17414 POR2X1_278/Y PAND2X1_216/B 0.07fF
C17415 PAND2X1_865/Y POR2X1_487/Y 0.00fF
C17416 POR2X1_188/A POR2X1_188/Y 0.00fF
C17417 PAND2X1_63/B POR2X1_294/B 0.03fF
C17418 PAND2X1_473/B POR2X1_129/Y 0.17fF
C17419 D_GATE_222 PAND2X1_60/B 2.17fF
C17420 POR2X1_116/Y POR2X1_392/CTRL 0.01fF
C17421 POR2X1_775/A POR2X1_510/Y 0.03fF
C17422 PAND2X1_793/Y PAND2X1_510/CTRL2 0.01fF
C17423 POR2X1_502/A POR2X1_6/CTRL 0.33fF
C17424 POR2X1_840/B PAND2X1_72/a_16_344# 0.03fF
C17425 POR2X1_706/B PAND2X1_692/O 0.00fF
C17426 POR2X1_407/Y POR2X1_644/A 0.03fF
C17427 POR2X1_49/Y PAND2X1_338/CTRL 0.01fF
C17428 POR2X1_795/B POR2X1_222/A 1.05fF
C17429 POR2X1_840/B POR2X1_532/A 3.53fF
C17430 POR2X1_140/A PAND2X1_60/B 0.01fF
C17431 PAND2X1_357/CTRL2 VDD 0.00fF
C17432 PAND2X1_605/CTRL2 POR2X1_42/Y 0.01fF
C17433 POR2X1_114/B POR2X1_383/A 0.06fF
C17434 PAND2X1_85/Y POR2X1_294/A 0.00fF
C17435 PAND2X1_29/a_76_28# POR2X1_68/B 0.02fF
C17436 POR2X1_158/Y POR2X1_669/B 0.10fF
C17437 POR2X1_81/A PAND2X1_390/Y 0.03fF
C17438 POR2X1_266/A POR2X1_547/B 0.02fF
C17439 POR2X1_419/O POR2X1_42/Y 0.10fF
C17440 PAND2X1_659/Y PAND2X1_473/B 0.06fF
C17441 POR2X1_458/Y POR2X1_556/A 0.07fF
C17442 PAND2X1_243/CTRL2 PAND2X1_338/B 0.03fF
C17443 POR2X1_291/O POR2X1_42/Y 0.01fF
C17444 POR2X1_198/O POR2X1_215/A 0.02fF
C17445 POR2X1_486/CTRL2 POR2X1_705/B 0.00fF
C17446 PAND2X1_489/CTRL2 PAND2X1_794/B 0.01fF
C17447 POR2X1_510/Y POR2X1_112/Y 0.10fF
C17448 POR2X1_192/Y POR2X1_564/B 0.05fF
C17449 POR2X1_493/B POR2X1_264/Y 0.01fF
C17450 POR2X1_220/B POR2X1_568/A 46.86fF
C17451 POR2X1_834/Y PAND2X1_433/O 0.04fF
C17452 POR2X1_16/A POR2X1_591/O 0.01fF
C17453 POR2X1_251/Y PAND2X1_360/Y 0.03fF
C17454 POR2X1_278/Y PAND2X1_359/Y 0.01fF
C17455 PAND2X1_236/CTRL2 POR2X1_4/Y 0.06fF
C17456 POR2X1_438/CTRL2 PAND2X1_569/B 0.01fF
C17457 PAND2X1_291/O PAND2X1_88/Y 0.02fF
C17458 POR2X1_416/B PAND2X1_478/B 0.01fF
C17459 POR2X1_854/B PAND2X1_32/B 0.05fF
C17460 POR2X1_57/A POR2X1_387/Y 0.07fF
C17461 POR2X1_390/B POR2X1_407/A 2.25fF
C17462 POR2X1_383/A POR2X1_649/B 0.16fF
C17463 D_INPUT_2 POR2X1_4/CTRL 0.01fF
C17464 POR2X1_62/Y PAND2X1_351/Y 0.03fF
C17465 PAND2X1_94/Y POR2X1_202/A 0.06fF
C17466 POR2X1_416/B POR2X1_609/CTRL 0.03fF
C17467 POR2X1_514/Y POR2X1_244/Y 0.03fF
C17468 PAND2X1_115/O PAND2X1_853/B 0.04fF
C17469 D_GATE_222 POR2X1_332/O 0.02fF
C17470 PAND2X1_6/Y POR2X1_260/A 3.33fF
C17471 PAND2X1_865/Y PAND2X1_738/Y 0.10fF
C17472 POR2X1_57/A PAND2X1_121/O 0.01fF
C17473 POR2X1_356/A POR2X1_180/a_16_28# 0.10fF
C17474 POR2X1_865/B POR2X1_101/Y 2.37fF
C17475 PAND2X1_63/B PAND2X1_111/B 0.81fF
C17476 POR2X1_661/A POR2X1_66/A 1.49fF
C17477 POR2X1_334/Y POR2X1_193/O 0.05fF
C17478 PAND2X1_226/CTRL POR2X1_192/B 0.10fF
C17479 PAND2X1_469/B POR2X1_153/Y 0.03fF
C17480 POR2X1_62/Y PAND2X1_101/CTRL 0.01fF
C17481 POR2X1_540/CTRL POR2X1_703/A 0.12fF
C17482 POR2X1_68/A POR2X1_186/B 0.09fF
C17483 POR2X1_383/A POR2X1_222/A 0.07fF
C17484 PAND2X1_6/Y POR2X1_363/A 0.25fF
C17485 POR2X1_8/Y POR2X1_68/B 0.03fF
C17486 POR2X1_216/a_56_344# POR2X1_116/Y 0.00fF
C17487 POR2X1_509/B PAND2X1_72/A 0.03fF
C17488 POR2X1_734/a_16_28# PAND2X1_32/B 0.03fF
C17489 PAND2X1_55/Y POR2X1_512/O 0.18fF
C17490 POR2X1_548/B POR2X1_4/Y 0.26fF
C17491 PAND2X1_6/Y PAND2X1_142/O 0.17fF
C17492 PAND2X1_466/A PAND2X1_466/B 0.16fF
C17493 POR2X1_614/A PAND2X1_313/m4_208_n4# 0.09fF
C17494 PAND2X1_175/B PAND2X1_175/O 0.00fF
C17495 POR2X1_253/Y PAND2X1_508/Y 0.00fF
C17496 POR2X1_68/A POR2X1_802/A 0.01fF
C17497 POR2X1_119/Y PAND2X1_514/Y 0.03fF
C17498 POR2X1_227/B POR2X1_776/A 0.03fF
C17499 POR2X1_283/A PAND2X1_130/a_76_28# 0.02fF
C17500 POR2X1_316/Y POR2X1_7/B 0.03fF
C17501 POR2X1_111/Y POR2X1_387/Y 0.04fF
C17502 POR2X1_461/Y POR2X1_859/a_16_28# 0.03fF
C17503 PAND2X1_382/O POR2X1_260/A 0.03fF
C17504 PAND2X1_724/B PAND2X1_326/B 0.00fF
C17505 POR2X1_537/Y POR2X1_513/Y 0.03fF
C17506 PAND2X1_129/CTRL2 PAND2X1_90/A 0.03fF
C17507 PAND2X1_661/Y PAND2X1_121/a_76_28# 0.02fF
C17508 POR2X1_709/O INPUT_1 0.01fF
C17509 POR2X1_245/CTRL PAND2X1_156/A 0.06fF
C17510 POR2X1_817/A POR2X1_77/Y 0.05fF
C17511 POR2X1_27/CTRL2 POR2X1_32/A 0.01fF
C17512 POR2X1_318/m4_208_n4# POR2X1_471/A 0.09fF
C17513 POR2X1_123/A POR2X1_520/B 0.01fF
C17514 PAND2X1_246/CTRL2 POR2X1_66/A -0.02fF
C17515 PAND2X1_437/CTRL2 POR2X1_186/Y 0.03fF
C17516 PAND2X1_454/CTRL2 POR2X1_77/Y 0.19fF
C17517 PAND2X1_69/A POR2X1_342/a_76_344# 0.01fF
C17518 POR2X1_137/Y POR2X1_294/A 0.03fF
C17519 POR2X1_294/B POR2X1_342/A 0.01fF
C17520 PAND2X1_193/Y PAND2X1_733/a_76_28# 0.07fF
C17521 POR2X1_57/A PAND2X1_737/CTRL2 0.01fF
C17522 POR2X1_86/O PAND2X1_6/A 0.05fF
C17523 PAND2X1_322/m4_208_n4# POR2X1_374/m4_208_n4# 0.13fF
C17524 PAND2X1_643/Y PAND2X1_729/O 0.01fF
C17525 PAND2X1_467/Y PAND2X1_451/CTRL 0.01fF
C17526 POR2X1_42/Y POR2X1_77/Y 0.60fF
C17527 POR2X1_180/B POR2X1_186/B 0.00fF
C17528 POR2X1_52/A POR2X1_387/a_76_344# 0.01fF
C17529 PAND2X1_865/Y PAND2X1_575/O 0.00fF
C17530 POR2X1_439/Y POR2X1_440/O 0.07fF
C17531 PAND2X1_547/CTRL POR2X1_39/B 0.01fF
C17532 D_INPUT_3 PAND2X1_610/CTRL 0.01fF
C17533 POR2X1_411/B POR2X1_268/CTRL2 0.01fF
C17534 POR2X1_309/Y POR2X1_77/Y 0.43fF
C17535 POR2X1_832/B PAND2X1_72/A 0.04fF
C17536 PAND2X1_310/O POR2X1_260/A 0.16fF
C17537 PAND2X1_578/Y GATE_579 0.01fF
C17538 POR2X1_23/Y POR2X1_24/Y 0.11fF
C17539 POR2X1_597/CTRL2 POR2X1_761/A 0.01fF
C17540 PAND2X1_23/Y PAND2X1_135/CTRL2 0.01fF
C17541 PAND2X1_26/CTRL D_INPUT_4 0.01fF
C17542 POR2X1_334/Y POR2X1_259/B 0.02fF
C17543 POR2X1_66/B PAND2X1_612/O 0.17fF
C17544 POR2X1_845/A POR2X1_673/Y 0.00fF
C17545 POR2X1_343/Y PAND2X1_96/B 0.05fF
C17546 POR2X1_833/A POR2X1_294/A 4.20fF
C17547 PAND2X1_848/CTRL INPUT_3 0.49fF
C17548 POR2X1_532/A PAND2X1_56/A 0.03fF
C17549 POR2X1_52/A PAND2X1_860/A 0.03fF
C17550 POR2X1_634/A POR2X1_859/CTRL 0.08fF
C17551 POR2X1_293/Y POR2X1_386/Y 0.01fF
C17552 POR2X1_440/O POR2X1_192/Y 0.04fF
C17553 PAND2X1_480/CTRL POR2X1_119/Y 0.01fF
C17554 POR2X1_139/CTRL POR2X1_138/A 0.01fF
C17555 POR2X1_816/O POR2X1_750/B 0.06fF
C17556 POR2X1_48/A POR2X1_626/CTRL2 0.01fF
C17557 PAND2X1_58/A POR2X1_624/Y 0.00fF
C17558 POR2X1_590/A POR2X1_447/A 0.54fF
C17559 POR2X1_329/A POR2X1_237/O 0.03fF
C17560 POR2X1_311/CTRL2 POR2X1_77/Y 0.02fF
C17561 POR2X1_61/a_16_28# POR2X1_447/B 0.06fF
C17562 POR2X1_67/Y INPUT_0 0.07fF
C17563 POR2X1_97/A POR2X1_567/B 0.05fF
C17564 POR2X1_130/a_16_28# POR2X1_260/B 0.03fF
C17565 POR2X1_369/a_16_28# POR2X1_119/Y 0.03fF
C17566 POR2X1_119/Y POR2X1_75/Y 0.06fF
C17567 PAND2X1_474/O PAND2X1_474/A 0.04fF
C17568 PAND2X1_415/CTRL POR2X1_414/Y 0.01fF
C17569 POR2X1_632/Y POR2X1_260/A 0.03fF
C17570 POR2X1_68/A PAND2X1_628/O 0.02fF
C17571 POR2X1_294/A POR2X1_195/m4_208_n4# 0.09fF
C17572 POR2X1_685/A PAND2X1_52/B 0.02fF
C17573 PAND2X1_213/Y POR2X1_166/Y 0.05fF
C17574 PAND2X1_39/B POR2X1_61/Y 0.02fF
C17575 POR2X1_66/B POR2X1_493/A 0.03fF
C17576 POR2X1_169/A POR2X1_186/B 0.03fF
C17577 POR2X1_150/Y PAND2X1_556/B 0.07fF
C17578 PAND2X1_436/O PAND2X1_390/Y 0.01fF
C17579 POR2X1_416/B PAND2X1_343/O 0.03fF
C17580 PAND2X1_624/a_16_344# POR2X1_20/B 0.02fF
C17581 POR2X1_495/a_16_28# POR2X1_283/A 0.02fF
C17582 POR2X1_814/A POR2X1_733/A 0.03fF
C17583 PAND2X1_464/B POR2X1_372/Y 0.01fF
C17584 POR2X1_334/B POR2X1_814/A 0.07fF
C17585 POR2X1_567/A POR2X1_552/A 0.13fF
C17586 POR2X1_666/CTRL2 POR2X1_102/Y 0.01fF
C17587 PAND2X1_52/B POR2X1_260/A 0.18fF
C17588 POR2X1_23/Y PAND2X1_208/CTRL 0.01fF
C17589 POR2X1_408/Y POR2X1_386/Y 0.13fF
C17590 POR2X1_383/CTRL2 POR2X1_383/Y 0.01fF
C17591 POR2X1_78/A POR2X1_454/B 0.03fF
C17592 POR2X1_711/Y POR2X1_151/Y 0.04fF
C17593 POR2X1_728/CTRL POR2X1_452/Y 0.01fF
C17594 PAND2X1_70/O POR2X1_635/A 0.02fF
C17595 POR2X1_66/B PAND2X1_413/CTRL 0.01fF
C17596 POR2X1_427/CTRL POR2X1_72/B 0.01fF
C17597 POR2X1_542/O POR2X1_552/A 0.00fF
C17598 POR2X1_593/m4_208_n4# PAND2X1_72/A 0.22fF
C17599 POR2X1_582/Y VDD 0.30fF
C17600 POR2X1_483/A POR2X1_260/B 0.03fF
C17601 POR2X1_837/B PAND2X1_505/O 0.01fF
C17602 POR2X1_748/A POR2X1_29/A 0.73fF
C17603 POR2X1_124/B POR2X1_814/A 2.01fF
C17604 POR2X1_504/Y POR2X1_626/O 0.01fF
C17605 POR2X1_620/A PAND2X1_41/B 0.01fF
C17606 POR2X1_88/CTRL INPUT_0 0.07fF
C17607 POR2X1_862/A VDD 1.24fF
C17608 PAND2X1_655/B POR2X1_600/CTRL2 0.01fF
C17609 POR2X1_252/Y POR2X1_77/Y 0.05fF
C17610 POR2X1_502/A POR2X1_602/CTRL2 0.01fF
C17611 POR2X1_54/Y POR2X1_7/B 0.13fF
C17612 POR2X1_378/a_16_28# D_INPUT_0 0.03fF
C17613 D_INPUT_0 PAND2X1_332/O 0.05fF
C17614 PAND2X1_402/CTRL2 POR2X1_14/Y 0.01fF
C17615 POR2X1_150/Y POR2X1_599/A 0.03fF
C17616 POR2X1_12/A INPUT_5 0.07fF
C17617 POR2X1_667/A POR2X1_40/Y 0.77fF
C17618 POR2X1_257/A PAND2X1_254/CTRL 0.01fF
C17619 POR2X1_60/A PAND2X1_558/Y 0.03fF
C17620 POR2X1_79/a_16_28# POR2X1_79/A 0.00fF
C17621 PAND2X1_93/B POR2X1_215/O 0.18fF
C17622 POR2X1_48/A PAND2X1_62/a_76_28# 0.02fF
C17623 PAND2X1_571/A PAND2X1_579/B 0.01fF
C17624 PAND2X1_571/CTRL2 PAND2X1_571/Y 0.00fF
C17625 POR2X1_614/A POR2X1_864/A 0.21fF
C17626 PAND2X1_20/A PAND2X1_20/CTRL 0.01fF
C17627 POR2X1_832/Y POR2X1_307/Y 0.05fF
C17628 PAND2X1_717/A PAND2X1_168/O 0.02fF
C17629 POR2X1_9/Y POR2X1_750/Y 0.01fF
C17630 PAND2X1_472/A POR2X1_20/B 0.10fF
C17631 POR2X1_440/CTRL2 POR2X1_353/A 0.00fF
C17632 POR2X1_119/Y PAND2X1_332/Y 0.07fF
C17633 PAND2X1_20/A POR2X1_61/Y 0.03fF
C17634 POR2X1_556/A D_INPUT_1 0.03fF
C17635 POR2X1_866/a_16_28# POR2X1_750/B 0.03fF
C17636 POR2X1_446/B POR2X1_732/B 0.01fF
C17637 PAND2X1_39/B POR2X1_35/Y 0.09fF
C17638 POR2X1_13/A POR2X1_263/Y 0.02fF
C17639 POR2X1_348/A POR2X1_244/CTRL 0.01fF
C17640 PAND2X1_88/O PAND2X1_41/B 0.03fF
C17641 POR2X1_347/A PAND2X1_94/Y 0.03fF
C17642 POR2X1_32/A PAND2X1_362/B 0.10fF
C17643 PAND2X1_621/Y POR2X1_48/A 0.01fF
C17644 POR2X1_262/Y POR2X1_38/Y 0.07fF
C17645 POR2X1_83/B PAND2X1_723/Y 0.03fF
C17646 PAND2X1_73/Y VDD 4.78fF
C17647 POR2X1_188/A POR2X1_862/B 0.01fF
C17648 POR2X1_422/Y VDD 0.13fF
C17649 POR2X1_556/A POR2X1_724/A 0.03fF
C17650 PAND2X1_564/B PAND2X1_564/CTRL2 0.03fF
C17651 PAND2X1_438/CTRL POR2X1_544/B 0.01fF
C17652 POR2X1_72/B PAND2X1_714/A 0.07fF
C17653 POR2X1_185/CTRL POR2X1_260/B 0.01fF
C17654 POR2X1_366/Y POR2X1_567/B 0.10fF
C17655 POR2X1_567/B POR2X1_294/B 0.05fF
C17656 PAND2X1_48/B POR2X1_476/A 0.03fF
C17657 PAND2X1_149/CTRL POR2X1_669/B 0.02fF
C17658 POR2X1_182/a_16_28# POR2X1_181/Y 0.03fF
C17659 PAND2X1_96/B POR2X1_624/Y 0.11fF
C17660 POR2X1_257/A PAND2X1_785/O 0.14fF
C17661 POR2X1_20/B POR2X1_380/Y 0.02fF
C17662 POR2X1_48/Y POR2X1_409/B 0.03fF
C17663 PAND2X1_20/A PAND2X1_755/O 0.00fF
C17664 POR2X1_83/B PAND2X1_435/O 0.05fF
C17665 POR2X1_186/Y POR2X1_798/a_76_344# 0.04fF
C17666 PAND2X1_390/Y PAND2X1_499/Y 0.03fF
C17667 POR2X1_49/CTRL POR2X1_236/Y 0.12fF
C17668 POR2X1_846/Y POR2X1_754/CTRL2 0.01fF
C17669 POR2X1_60/A PAND2X1_480/B 0.03fF
C17670 POR2X1_121/B POR2X1_405/Y 0.03fF
C17671 POR2X1_56/O POR2X1_293/Y 0.08fF
C17672 POR2X1_781/B POR2X1_781/A 0.00fF
C17673 PAND2X1_58/A INPUT_4 0.02fF
C17674 POR2X1_150/Y PAND2X1_175/CTRL2 0.10fF
C17675 POR2X1_121/B POR2X1_784/A 0.03fF
C17676 PAND2X1_623/Y POR2X1_753/Y 0.07fF
C17677 POR2X1_814/B PAND2X1_54/CTRL2 0.03fF
C17678 POR2X1_72/B PAND2X1_558/a_56_28# 0.00fF
C17679 POR2X1_296/B PAND2X1_144/CTRL2 0.05fF
C17680 POR2X1_836/A POR2X1_776/B 0.03fF
C17681 PAND2X1_404/CTRL POR2X1_293/Y 0.01fF
C17682 POR2X1_558/CTRL2 POR2X1_78/A 0.03fF
C17683 POR2X1_815/Y POR2X1_38/B -0.00fF
C17684 POR2X1_610/O POR2X1_532/A 0.07fF
C17685 POR2X1_41/B PAND2X1_215/a_76_28# 0.01fF
C17686 POR2X1_431/O POR2X1_129/Y 0.02fF
C17687 PAND2X1_73/Y POR2X1_741/Y 0.03fF
C17688 POR2X1_202/A PAND2X1_60/B 0.34fF
C17689 PAND2X1_784/A POR2X1_7/B 0.03fF
C17690 POR2X1_341/A POR2X1_101/Y 0.10fF
C17691 POR2X1_244/B POR2X1_509/B 0.01fF
C17692 POR2X1_420/O POR2X1_90/Y 0.01fF
C17693 POR2X1_863/a_16_28# PAND2X1_73/Y 0.02fF
C17694 PAND2X1_652/A PAND2X1_794/CTRL 0.01fF
C17695 PAND2X1_512/a_76_28# INPUT_0 0.01fF
C17696 PAND2X1_81/B PAND2X1_73/Y 0.03fF
C17697 PAND2X1_340/CTRL2 POR2X1_88/Y 0.00fF
C17698 POR2X1_439/Y POR2X1_192/Y 0.13fF
C17699 PAND2X1_853/CTRL POR2X1_83/B 0.01fF
C17700 PAND2X1_20/A POR2X1_231/a_16_28# 0.01fF
C17701 POR2X1_73/a_16_28# POR2X1_20/B 0.00fF
C17702 POR2X1_133/CTRL2 POR2X1_236/Y 0.01fF
C17703 PAND2X1_695/CTRL2 PAND2X1_57/B 0.00fF
C17704 PAND2X1_48/B POR2X1_269/Y 0.07fF
C17705 POR2X1_859/CTRL2 POR2X1_559/A 0.02fF
C17706 POR2X1_54/Y POR2X1_773/O 0.01fF
C17707 PAND2X1_631/O POR2X1_669/B 0.04fF
C17708 PAND2X1_687/Y VDD 0.15fF
C17709 PAND2X1_69/CTRL POR2X1_296/B 0.01fF
C17710 PAND2X1_626/O D_GATE_222 0.06fF
C17711 PAND2X1_20/A POR2X1_35/Y 0.07fF
C17712 PAND2X1_793/Y PAND2X1_793/A 0.44fF
C17713 PAND2X1_650/CTRL POR2X1_409/B 0.01fF
C17714 POR2X1_377/CTRL2 POR2X1_94/A 0.01fF
C17715 POR2X1_660/Y POR2X1_840/B 0.24fF
C17716 POR2X1_748/A PAND2X1_506/O 0.05fF
C17717 POR2X1_528/Y POR2X1_613/O 0.05fF
C17718 PAND2X1_73/Y PAND2X1_32/B 0.47fF
C17719 POR2X1_692/a_76_344# POR2X1_526/Y -0.00fF
C17720 POR2X1_13/A PAND2X1_778/CTRL 0.01fF
C17721 D_INPUT_0 POR2X1_318/A 0.10fF
C17722 PAND2X1_852/CTRL POR2X1_40/Y 0.01fF
C17723 PAND2X1_736/a_16_344# PAND2X1_735/Y 0.02fF
C17724 POR2X1_315/Y PAND2X1_444/O 0.12fF
C17725 POR2X1_254/A D_GATE_222 0.03fF
C17726 POR2X1_569/a_16_28# POR2X1_192/Y 0.04fF
C17727 PAND2X1_811/O VDD 0.00fF
C17728 POR2X1_121/B POR2X1_249/O 0.07fF
C17729 POR2X1_596/A POR2X1_834/O 0.01fF
C17730 POR2X1_241/B POR2X1_570/B 0.02fF
C17731 POR2X1_133/CTRL VDD 0.00fF
C17732 POR2X1_804/a_16_28# POR2X1_532/A 0.03fF
C17733 POR2X1_296/B POR2X1_788/B 0.05fF
C17734 PAND2X1_610/O POR2X1_612/A 0.03fF
C17735 POR2X1_811/CTRL POR2X1_780/B 0.03fF
C17736 PAND2X1_115/Y POR2X1_106/Y 0.06fF
C17737 POR2X1_389/O POR2X1_389/Y 0.00fF
C17738 POR2X1_525/O POR2X1_763/Y 0.05fF
C17739 POR2X1_41/B PAND2X1_733/Y 0.09fF
C17740 POR2X1_567/B POR2X1_351/CTRL 0.01fF
C17741 POR2X1_346/A PAND2X1_60/B 0.03fF
C17742 PAND2X1_470/O POR2X1_83/B 0.04fF
C17743 PAND2X1_217/B PAND2X1_798/B 0.05fF
C17744 POR2X1_349/Y PAND2X1_57/B 0.01fF
C17745 POR2X1_78/B POR2X1_231/CTRL2 0.03fF
C17746 PAND2X1_354/A PAND2X1_794/B 0.03fF
C17747 POR2X1_636/A VDD 0.08fF
C17748 PAND2X1_787/Y PAND2X1_115/B 0.15fF
C17749 POR2X1_290/Y POR2X1_236/Y 0.04fF
C17750 POR2X1_677/CTRL PAND2X1_658/B 0.09fF
C17751 PAND2X1_607/CTRL PAND2X1_56/A 0.01fF
C17752 POR2X1_40/Y POR2X1_321/O 0.02fF
C17753 POR2X1_264/CTRL PAND2X1_32/B 0.01fF
C17754 POR2X1_556/A POR2X1_362/CTRL2 0.01fF
C17755 POR2X1_859/A POR2X1_668/Y 0.05fF
C17756 POR2X1_72/B POR2X1_816/A 1.57fF
C17757 INPUT_1 PAND2X1_637/CTRL 0.01fF
C17758 PAND2X1_433/a_16_344# POR2X1_807/A 0.01fF
C17759 POR2X1_65/A POR2X1_43/B 0.06fF
C17760 POR2X1_452/Y POR2X1_210/A 0.08fF
C17761 POR2X1_686/A POR2X1_149/B 0.01fF
C17762 POR2X1_687/B VDD 0.10fF
C17763 POR2X1_327/a_16_28# PAND2X1_65/B 0.02fF
C17764 PAND2X1_48/CTRL2 POR2X1_294/B 0.01fF
C17765 PAND2X1_653/O POR2X1_329/A 0.01fF
C17766 POR2X1_366/Y POR2X1_78/B 0.03fF
C17767 POR2X1_78/B POR2X1_294/B 1.44fF
C17768 PAND2X1_465/B VDD 0.22fF
C17769 POR2X1_730/Y POR2X1_856/B 0.03fF
C17770 POR2X1_330/Y POR2X1_541/O 0.02fF
C17771 POR2X1_32/A PAND2X1_717/Y 0.01fF
C17772 POR2X1_356/A POR2X1_566/A 0.10fF
C17773 POR2X1_238/Y POR2X1_236/Y 0.78fF
C17774 PAND2X1_55/Y PAND2X1_8/Y 0.09fF
C17775 POR2X1_13/A PAND2X1_215/B 0.02fF
C17776 PAND2X1_658/B POR2X1_236/Y 0.05fF
C17777 POR2X1_341/A PAND2X1_323/CTRL2 0.06fF
C17778 PAND2X1_56/Y POR2X1_335/CTRL 0.15fF
C17779 POR2X1_123/A PAND2X1_20/A 0.03fF
C17780 POR2X1_814/A POR2X1_343/a_16_28# 0.00fF
C17781 PAND2X1_803/Y PAND2X1_360/O 0.01fF
C17782 POR2X1_467/Y PAND2X1_534/CTRL 0.01fF
C17783 POR2X1_66/B POR2X1_510/Y 0.06fF
C17784 POR2X1_649/B POR2X1_476/a_16_28# 0.09fF
C17785 POR2X1_188/A POR2X1_121/CTRL 0.01fF
C17786 PAND2X1_69/A POR2X1_585/O 0.12fF
C17787 PAND2X1_124/Y PAND2X1_123/Y 0.03fF
C17788 POR2X1_220/B POR2X1_444/Y 0.03fF
C17789 PAND2X1_798/B VDD 0.22fF
C17790 POR2X1_509/A VDD 0.03fF
C17791 POR2X1_667/A PAND2X1_559/O 0.03fF
C17792 PAND2X1_771/Y PAND2X1_569/a_76_28# 0.02fF
C17793 PAND2X1_23/CTRL PAND2X1_60/B 0.01fF
C17794 PAND2X1_784/CTRL POR2X1_293/Y 0.01fF
C17795 D_INPUT_0 POR2X1_574/Y 0.12fF
C17796 POR2X1_661/Y POR2X1_353/A 0.02fF
C17797 VDD POR2X1_759/Y 0.00fF
C17798 POR2X1_96/A POR2X1_693/Y 0.02fF
C17799 PAND2X1_425/Y D_INPUT_4 0.03fF
C17800 PAND2X1_23/Y POR2X1_231/B 0.00fF
C17801 POR2X1_603/a_16_28# POR2X1_761/A 0.02fF
C17802 VDD POR2X1_631/B 0.18fF
C17803 POR2X1_13/Y POR2X1_7/B 1.67fF
C17804 POR2X1_853/A POR2X1_776/B 0.22fF
C17805 PAND2X1_808/B POR2X1_283/A 0.01fF
C17806 POR2X1_284/B PAND2X1_69/A 0.07fF
C17807 POR2X1_23/Y PAND2X1_851/CTRL 0.03fF
C17808 POR2X1_195/A POR2X1_195/a_16_28# 0.03fF
C17809 PAND2X1_206/O POR2X1_73/Y 0.02fF
C17810 PAND2X1_803/Y POR2X1_106/Y 0.26fF
C17811 POR2X1_599/A PAND2X1_364/B 0.10fF
C17812 POR2X1_356/A POR2X1_340/a_76_344# 0.10fF
C17813 PAND2X1_55/Y POR2X1_659/CTRL2 0.10fF
C17814 PAND2X1_293/CTRL2 POR2X1_68/B 0.06fF
C17815 POR2X1_467/Y POR2X1_260/A 0.03fF
C17816 POR2X1_66/B POR2X1_768/CTRL2 0.01fF
C17817 PAND2X1_287/Y POR2X1_767/m4_208_n4# 0.08fF
C17818 PAND2X1_691/Y POR2X1_666/Y 1.51fF
C17819 PAND2X1_76/Y PAND2X1_175/B 0.03fF
C17820 PAND2X1_90/Y POR2X1_713/B 1.56fF
C17821 POR2X1_567/A POR2X1_567/B 0.67fF
C17822 POR2X1_330/Y POR2X1_675/Y 0.04fF
C17823 INPUT_1 POR2X1_495/CTRL 0.00fF
C17824 POR2X1_185/CTRL PAND2X1_55/Y 0.03fF
C17825 POR2X1_78/B PAND2X1_111/B 0.03fF
C17826 POR2X1_41/B PAND2X1_243/CTRL2 0.00fF
C17827 PAND2X1_55/Y POR2X1_61/B 0.01fF
C17828 POR2X1_81/a_56_344# POR2X1_153/Y 0.03fF
C17829 PAND2X1_407/O POR2X1_39/B 0.11fF
C17830 POR2X1_83/B PAND2X1_123/Y 0.03fF
C17831 PAND2X1_132/CTRL2 PAND2X1_32/B 0.00fF
C17832 PAND2X1_80/O PAND2X1_60/B 0.01fF
C17833 POR2X1_793/O POR2X1_713/B 0.02fF
C17834 POR2X1_480/A POR2X1_590/CTRL 0.08fF
C17835 POR2X1_60/A POR2X1_373/Y 0.03fF
C17836 PAND2X1_48/B POR2X1_513/Y 0.03fF
C17837 POR2X1_651/O POR2X1_638/Y 0.00fF
C17838 PAND2X1_91/a_16_344# POR2X1_169/A 0.02fF
C17839 POR2X1_548/B D_INPUT_1 0.01fF
C17840 PAND2X1_140/A POR2X1_107/a_76_344# 0.00fF
C17841 PAND2X1_734/B PAND2X1_338/B 0.03fF
C17842 POR2X1_115/CTRL2 POR2X1_366/A 0.01fF
C17843 PAND2X1_48/B POR2X1_219/B 0.07fF
C17844 POR2X1_476/Y POR2X1_249/Y 0.02fF
C17845 POR2X1_186/Y POR2X1_507/A 0.07fF
C17846 POR2X1_16/A PAND2X1_721/O 0.01fF
C17847 PAND2X1_96/B POR2X1_785/A 0.69fF
C17848 PAND2X1_496/CTRL POR2X1_500/Y 0.01fF
C17849 POR2X1_351/Y POR2X1_350/CTRL 0.01fF
C17850 POR2X1_766/CTRL VDD -0.00fF
C17851 POR2X1_853/A POR2X1_577/CTRL2 0.01fF
C17852 PAND2X1_182/B POR2X1_312/Y 1.53fF
C17853 PAND2X1_476/A POR2X1_669/B 0.12fF
C17854 POR2X1_759/A POR2X1_759/a_16_28# 0.05fF
C17855 POR2X1_346/CTRL PAND2X1_55/Y 0.01fF
C17856 POR2X1_202/a_16_28# POR2X1_507/A 0.09fF
C17857 PAND2X1_787/A POR2X1_7/B 0.05fF
C17858 POR2X1_525/Y POR2X1_526/Y 0.01fF
C17859 POR2X1_750/A POR2X1_523/B 0.28fF
C17860 POR2X1_627/Y POR2X1_408/Y 0.02fF
C17861 POR2X1_45/Y POR2X1_498/A 0.01fF
C17862 POR2X1_514/Y POR2X1_501/B 0.05fF
C17863 PAND2X1_23/Y POR2X1_865/B 0.07fF
C17864 PAND2X1_23/Y PAND2X1_88/Y 0.03fF
C17865 POR2X1_46/Y PAND2X1_656/A 0.03fF
C17866 PAND2X1_94/A PAND2X1_54/a_16_344# 0.02fF
C17867 PAND2X1_691/Y VDD 0.34fF
C17868 PAND2X1_46/CTRL PAND2X1_71/Y 0.01fF
C17869 POR2X1_13/A POR2X1_588/Y 6.52fF
C17870 POR2X1_606/a_56_344# PAND2X1_56/A 0.00fF
C17871 POR2X1_566/A POR2X1_569/A 0.10fF
C17872 POR2X1_3/A POR2X1_700/O 0.03fF
C17873 POR2X1_78/CTRL POR2X1_844/B 0.01fF
C17874 PAND2X1_391/a_76_28# POR2X1_4/Y 0.01fF
C17875 POR2X1_831/a_16_28# POR2X1_717/B 0.01fF
C17876 POR2X1_383/A POR2X1_405/Y 0.10fF
C17877 POR2X1_40/Y POR2X1_183/O 0.01fF
C17878 POR2X1_466/a_76_344# POR2X1_209/A 0.01fF
C17879 POR2X1_341/A POR2X1_579/O 0.05fF
C17880 POR2X1_65/A PAND2X1_170/CTRL 0.01fF
C17881 PAND2X1_682/O PAND2X1_69/A 0.03fF
C17882 POR2X1_68/A POR2X1_542/B 0.03fF
C17883 POR2X1_376/B PAND2X1_708/CTRL2 0.01fF
C17884 POR2X1_425/CTRL2 POR2X1_158/B 0.01fF
C17885 POR2X1_383/A POR2X1_784/A 0.03fF
C17886 POR2X1_283/A POR2X1_372/Y 0.68fF
C17887 POR2X1_566/A POR2X1_97/CTRL 0.14fF
C17888 PAND2X1_462/CTRL POR2X1_37/Y -0.00fF
C17889 POR2X1_334/B POR2X1_493/O 0.02fF
C17890 POR2X1_769/A POR2X1_769/B 0.00fF
C17891 PAND2X1_48/B POR2X1_366/A 0.05fF
C17892 POR2X1_332/Y POR2X1_61/Y 0.00fF
C17893 PAND2X1_251/CTRL2 POR2X1_717/B 0.01fF
C17894 POR2X1_376/B PAND2X1_156/A 0.05fF
C17895 POR2X1_76/Y POR2X1_456/B 1.10fF
C17896 PAND2X1_738/Y PAND2X1_343/O 0.02fF
C17897 POR2X1_41/B POR2X1_83/O 0.00fF
C17898 POR2X1_48/A POR2X1_747/a_56_344# 0.00fF
C17899 POR2X1_193/A POR2X1_553/A 0.03fF
C17900 PAND2X1_23/Y PAND2X1_373/CTRL2 0.01fF
C17901 PAND2X1_274/CTRL2 POR2X1_153/Y 0.00fF
C17902 PAND2X1_566/Y POR2X1_142/Y 0.07fF
C17903 PAND2X1_808/O POR2X1_283/A 0.02fF
C17904 PAND2X1_476/A PAND2X1_231/CTRL 0.00fF
C17905 PAND2X1_173/CTRL2 PAND2X1_32/B 0.01fF
C17906 POR2X1_364/A POR2X1_578/a_56_344# 0.00fF
C17907 D_GATE_662 POR2X1_180/A 0.07fF
C17908 POR2X1_124/m4_208_n4# POR2X1_493/m4_208_n4# 0.13fF
C17909 POR2X1_46/Y PAND2X1_348/A 0.10fF
C17910 POR2X1_628/CTRL POR2X1_260/A 0.01fF
C17911 PAND2X1_467/CTRL2 PAND2X1_725/A 0.00fF
C17912 POR2X1_664/O POR2X1_664/Y 0.05fF
C17913 PAND2X1_349/A POR2X1_56/Y 0.03fF
C17914 PAND2X1_65/B POR2X1_357/B 0.01fF
C17915 PAND2X1_847/O POR2X1_32/A 0.01fF
C17916 POR2X1_334/Y PAND2X1_89/CTRL2 0.03fF
C17917 POR2X1_740/Y POR2X1_456/B 0.05fF
C17918 PAND2X1_6/Y POR2X1_725/Y 0.07fF
C17919 PAND2X1_95/B POR2X1_260/A 0.05fF
C17920 PAND2X1_241/O PAND2X1_308/Y 0.03fF
C17921 PAND2X1_476/A POR2X1_230/O 0.00fF
C17922 POR2X1_569/A POR2X1_844/B 0.23fF
C17923 PAND2X1_308/Y PAND2X1_302/CTRL2 0.01fF
C17924 POR2X1_119/Y PAND2X1_474/Y 0.05fF
C17925 POR2X1_435/Y POR2X1_802/A 0.09fF
C17926 PAND2X1_390/Y POR2X1_39/B 0.08fF
C17927 POR2X1_46/Y POR2X1_300/Y 0.05fF
C17928 POR2X1_78/B POR2X1_567/A 0.13fF
C17929 POR2X1_481/A PAND2X1_336/Y 0.01fF
C17930 POR2X1_463/Y POR2X1_805/A 0.00fF
C17931 POR2X1_326/A POR2X1_468/B 0.58fF
C17932 PAND2X1_213/A POR2X1_394/A 0.01fF
C17933 POR2X1_52/A PAND2X1_156/A 0.05fF
C17934 POR2X1_569/A POR2X1_573/A 0.05fF
C17935 POR2X1_119/Y POR2X1_13/A 0.25fF
C17936 PAND2X1_661/CTRL PAND2X1_659/Y 0.00fF
C17937 PAND2X1_94/A PAND2X1_69/A 3.32fF
C17938 POR2X1_634/A PAND2X1_72/A 0.05fF
C17939 POR2X1_172/Y PAND2X1_549/B 0.01fF
C17940 PAND2X1_803/Y PAND2X1_349/A 0.03fF
C17941 PAND2X1_481/O POR2X1_222/Y 0.04fF
C17942 PAND2X1_358/A PAND2X1_101/O 0.07fF
C17943 POR2X1_324/Y POR2X1_468/B 0.00fF
C17944 POR2X1_68/B POR2X1_561/O 0.00fF
C17945 POR2X1_54/Y PAND2X1_206/B 0.05fF
C17946 PAND2X1_724/O PAND2X1_714/Y 0.06fF
C17947 VDD POR2X1_365/CTRL -0.00fF
C17948 POR2X1_316/O POR2X1_43/B 0.18fF
C17949 POR2X1_16/A PAND2X1_645/B 0.05fF
C17950 PAND2X1_803/Y PAND2X1_114/B 0.03fF
C17951 POR2X1_294/B POR2X1_294/A 2.41fF
C17952 PAND2X1_631/A POR2X1_46/Y 0.10fF
C17953 PAND2X1_835/a_76_28# POR2X1_394/A 0.02fF
C17954 POR2X1_7/B POR2X1_4/Y 0.03fF
C17955 POR2X1_137/B POR2X1_556/A 0.02fF
C17956 POR2X1_493/B POR2X1_493/CTRL 0.04fF
C17957 POR2X1_365/Y POR2X1_191/Y 0.05fF
C17958 PAND2X1_23/Y POR2X1_508/A 0.01fF
C17959 PAND2X1_824/B POR2X1_447/CTRL 0.07fF
C17960 PAND2X1_23/Y POR2X1_359/O 0.01fF
C17961 POR2X1_853/A POR2X1_192/B 0.05fF
C17962 POR2X1_367/a_16_28# POR2X1_169/A 0.03fF
C17963 POR2X1_327/Y POR2X1_112/Y 0.00fF
C17964 POR2X1_78/B PAND2X1_166/a_76_28# 0.05fF
C17965 PAND2X1_211/CTRL2 POR2X1_20/B 0.00fF
C17966 PAND2X1_96/B POR2X1_186/B 0.13fF
C17967 PAND2X1_501/CTRL2 PAND2X1_862/B 0.01fF
C17968 POR2X1_347/A PAND2X1_60/B 0.01fF
C17969 POR2X1_352/O POR2X1_854/B 0.33fF
C17970 PAND2X1_455/Y POR2X1_77/Y 0.03fF
C17971 PAND2X1_93/B PAND2X1_86/O 0.03fF
C17972 INPUT_3 PAND2X1_33/m4_208_n4# 0.06fF
C17973 PAND2X1_775/CTRL2 POR2X1_77/Y 0.01fF
C17974 POR2X1_730/Y POR2X1_151/CTRL2 0.01fF
C17975 PAND2X1_212/CTRL2 POR2X1_20/B 0.00fF
C17976 POR2X1_431/O POR2X1_37/Y 0.01fF
C17977 PAND2X1_23/Y POR2X1_568/B 0.05fF
C17978 POR2X1_130/A PAND2X1_72/A 0.06fF
C17979 POR2X1_119/Y PAND2X1_661/B 0.05fF
C17980 PAND2X1_462/CTRL POR2X1_293/Y 0.01fF
C17981 PAND2X1_221/Y PAND2X1_354/A 0.03fF
C17982 POR2X1_539/A POR2X1_733/Y 0.01fF
C17983 POR2X1_16/A PAND2X1_737/B 0.05fF
C17984 POR2X1_20/B POR2X1_260/B 0.07fF
C17985 POR2X1_25/Y POR2X1_3/A 0.07fF
C17986 POR2X1_65/O D_INPUT_0 0.02fF
C17987 POR2X1_375/a_76_344# POR2X1_260/A 0.00fF
C17988 POR2X1_566/A PAND2X1_72/A 0.14fF
C17989 POR2X1_16/A PAND2X1_216/B 0.12fF
C17990 PAND2X1_93/B POR2X1_556/A 0.06fF
C17991 POR2X1_270/CTRL POR2X1_567/A 0.01fF
C17992 PAND2X1_111/B POR2X1_294/A 0.03fF
C17993 PAND2X1_849/B PAND2X1_358/A 0.07fF
C17994 PAND2X1_73/Y POR2X1_688/CTRL2 0.01fF
C17995 POR2X1_4/Y PAND2X1_60/B 0.12fF
C17996 POR2X1_813/CTRL POR2X1_263/Y 0.01fF
C17997 POR2X1_123/O PAND2X1_72/A -0.00fF
C17998 PAND2X1_723/A PAND2X1_716/B 0.01fF
C17999 POR2X1_83/Y POR2X1_229/Y 0.02fF
C18000 PAND2X1_110/O PAND2X1_52/B 0.06fF
C18001 POR2X1_168/CTRL2 POR2X1_566/B 0.17fF
C18002 PAND2X1_557/A POR2X1_250/Y 0.01fF
C18003 POR2X1_35/B POR2X1_621/CTRL 0.01fF
C18004 POR2X1_532/A PAND2X1_134/a_76_28# 0.06fF
C18005 POR2X1_186/CTRL POR2X1_326/A 0.05fF
C18006 POR2X1_834/Y PAND2X1_48/A 0.10fF
C18007 POR2X1_23/Y PAND2X1_407/a_16_344# 0.00fF
C18008 PAND2X1_862/B PAND2X1_860/A 0.20fF
C18009 POR2X1_78/A POR2X1_556/A 2.22fF
C18010 POR2X1_329/A PAND2X1_733/O 0.01fF
C18011 POR2X1_495/a_16_28# POR2X1_55/Y 0.03fF
C18012 POR2X1_466/A POR2X1_446/B 0.02fF
C18013 POR2X1_499/A POR2X1_474/CTRL2 0.01fF
C18014 PAND2X1_73/Y PAND2X1_9/Y 0.00fF
C18015 PAND2X1_111/O PAND2X1_72/A 0.15fF
C18016 D_INPUT_5 PAND2X1_752/CTRL2 0.04fF
C18017 POR2X1_65/A POR2X1_292/a_16_28# 0.03fF
C18018 POR2X1_416/B POR2X1_108/CTRL2 0.01fF
C18019 PAND2X1_417/CTRL POR2X1_750/B 0.14fF
C18020 POR2X1_846/Y POR2X1_752/Y 0.00fF
C18021 PAND2X1_437/a_76_28# POR2X1_192/Y 0.05fF
C18022 POR2X1_38/O POR2X1_37/Y 0.05fF
C18023 PAND2X1_282/CTRL POR2X1_260/B 0.01fF
C18024 POR2X1_500/O POR2X1_500/Y 0.00fF
C18025 POR2X1_227/B POR2X1_242/O 0.03fF
C18026 POR2X1_491/O POR2X1_150/Y 0.01fF
C18027 POR2X1_373/Y POR2X1_373/CTRL2 0.01fF
C18028 POR2X1_49/Y PAND2X1_201/O 0.02fF
C18029 POR2X1_602/CTRL POR2X1_296/B 0.04fF
C18030 PAND2X1_72/A POR2X1_573/A 0.03fF
C18031 POR2X1_32/CTRL POR2X1_29/Y 0.01fF
C18032 POR2X1_736/A POR2X1_128/B 0.25fF
C18033 PAND2X1_571/A PAND2X1_571/O 0.00fF
C18034 PAND2X1_418/m4_208_n4# PAND2X1_41/B 0.12fF
C18035 POR2X1_71/a_16_28# POR2X1_62/Y 0.03fF
C18036 PAND2X1_830/CTRL2 POR2X1_416/B 0.01fF
C18037 POR2X1_731/a_16_28# PAND2X1_52/B 0.03fF
C18038 POR2X1_270/Y POR2X1_269/CTRL 0.01fF
C18039 PAND2X1_269/a_16_344# INPUT_0 0.04fF
C18040 PAND2X1_221/Y PAND2X1_730/CTRL 0.00fF
C18041 POR2X1_378/O PAND2X1_9/Y 0.01fF
C18042 POR2X1_326/A POR2X1_324/Y 0.04fF
C18043 POR2X1_475/O POR2X1_734/A 0.03fF
C18044 POR2X1_54/Y POR2X1_750/B 0.06fF
C18045 POR2X1_812/A POR2X1_809/CTRL2 0.01fF
C18046 PAND2X1_48/B PAND2X1_234/a_16_344# 0.01fF
C18047 POR2X1_20/B PAND2X1_803/A 0.03fF
C18048 PAND2X1_657/O POR2X1_23/Y 0.07fF
C18049 PAND2X1_666/CTRL PAND2X1_73/Y 0.01fF
C18050 POR2X1_490/Y PAND2X1_557/A 0.01fF
C18051 POR2X1_274/A POR2X1_141/Y 0.03fF
C18052 PAND2X1_492/O POR2X1_556/A 0.02fF
C18053 POR2X1_568/A POR2X1_854/B 0.03fF
C18054 PAND2X1_96/B PAND2X1_628/O 0.01fF
C18055 POR2X1_864/A PAND2X1_760/CTRL 0.00fF
C18056 PAND2X1_73/CTRL2 POR2X1_66/A 0.02fF
C18057 PAND2X1_214/CTRL PAND2X1_214/A 0.00fF
C18058 PAND2X1_807/O PAND2X1_221/Y 0.02fF
C18059 POR2X1_452/O VDD 0.00fF
C18060 POR2X1_20/B PAND2X1_673/Y 0.20fF
C18061 POR2X1_66/B POR2X1_98/CTRL 0.00fF
C18062 POR2X1_48/A PAND2X1_540/CTRL2 0.01fF
C18063 POR2X1_753/Y PAND2X1_58/A 0.10fF
C18064 POR2X1_416/B PAND2X1_537/a_76_28# 0.02fF
C18065 POR2X1_260/B PAND2X1_381/CTRL2 0.03fF
C18066 D_INPUT_0 POR2X1_40/Y 3.67fF
C18067 PAND2X1_817/O POR2X1_29/A 0.02fF
C18068 POR2X1_497/O POR2X1_32/A 0.01fF
C18069 POR2X1_814/A POR2X1_562/B 0.03fF
C18070 POR2X1_862/A POR2X1_472/Y 0.04fF
C18071 POR2X1_559/A PAND2X1_52/B 0.07fF
C18072 POR2X1_35/B D_INPUT_0 0.03fF
C18073 POR2X1_260/B POR2X1_410/CTRL2 0.01fF
C18074 POR2X1_78/A POR2X1_474/O 0.02fF
C18075 POR2X1_436/B POR2X1_436/O 0.02fF
C18076 PAND2X1_61/CTRL PAND2X1_61/Y 0.01fF
C18077 PAND2X1_73/Y POR2X1_808/A 0.03fF
C18078 POR2X1_462/CTRL2 PAND2X1_69/A 0.02fF
C18079 POR2X1_23/Y POR2X1_697/O 0.01fF
C18080 POR2X1_433/CTRL2 POR2X1_72/B 0.03fF
C18081 POR2X1_62/Y POR2X1_522/a_56_344# 0.00fF
C18082 POR2X1_278/Y PAND2X1_205/CTRL 0.05fF
C18083 POR2X1_458/Y PAND2X1_60/B 1.20fF
C18084 PAND2X1_719/Y PAND2X1_718/Y 0.00fF
C18085 POR2X1_296/B POR2X1_788/O 0.04fF
C18086 PAND2X1_93/B POR2X1_400/A 0.01fF
C18087 POR2X1_286/B POR2X1_294/B 0.22fF
C18088 POR2X1_179/CTRL2 POR2X1_411/B 0.01fF
C18089 POR2X1_322/a_76_344# POR2X1_441/Y 0.00fF
C18090 PAND2X1_23/Y POR2X1_341/A 0.10fF
C18091 PAND2X1_846/a_76_28# POR2X1_816/Y 0.02fF
C18092 POR2X1_32/A POR2X1_226/Y 0.00fF
C18093 POR2X1_654/O POR2X1_121/B 0.02fF
C18094 POR2X1_661/A POR2X1_308/B 0.03fF
C18095 POR2X1_628/Y POR2X1_55/Y 0.04fF
C18096 PAND2X1_576/B PAND2X1_571/Y 0.03fF
C18097 POR2X1_49/Y POR2X1_820/CTRL2 0.00fF
C18098 PAND2X1_771/Y PAND2X1_580/B 0.17fF
C18099 POR2X1_333/A POR2X1_186/Y 0.02fF
C18100 POR2X1_66/B POR2X1_404/CTRL2 0.00fF
C18101 POR2X1_496/Y POR2X1_627/O 0.03fF
C18102 POR2X1_460/Y PAND2X1_69/A 0.03fF
C18103 POR2X1_633/A POR2X1_734/A 0.47fF
C18104 POR2X1_335/O POR2X1_66/A 0.01fF
C18105 POR2X1_590/A POR2X1_362/B 4.58fF
C18106 PAND2X1_255/CTRL2 POR2X1_260/A 0.01fF
C18107 PAND2X1_266/CTRL2 POR2X1_7/A 0.01fF
C18108 POR2X1_290/a_56_344# POR2X1_83/B 0.01fF
C18109 POR2X1_665/O POR2X1_665/A 0.03fF
C18110 POR2X1_104/CTRL POR2X1_5/Y 0.00fF
C18111 POR2X1_806/O POR2X1_807/A 0.01fF
C18112 PAND2X1_863/a_16_344# POR2X1_102/Y 0.01fF
C18113 PAND2X1_557/A PAND2X1_205/Y 0.02fF
C18114 PAND2X1_43/CTRL2 PAND2X1_69/A 0.01fF
C18115 POR2X1_329/A POR2X1_385/CTRL2 0.04fF
C18116 POR2X1_847/A POR2X1_847/B 0.01fF
C18117 PAND2X1_95/B PAND2X1_31/CTRL2 0.01fF
C18118 POR2X1_678/O PAND2X1_69/A 0.01fF
C18119 POR2X1_83/B POR2X1_48/CTRL 0.00fF
C18120 POR2X1_694/CTRL POR2X1_257/A 0.01fF
C18121 POR2X1_48/A POR2X1_232/CTRL 0.01fF
C18122 POR2X1_528/m4_208_n4# PAND2X1_447/m4_208_n4# 0.13fF
C18123 PAND2X1_793/Y POR2X1_37/Y 0.03fF
C18124 POR2X1_407/A POR2X1_676/O 0.01fF
C18125 POR2X1_60/A PAND2X1_473/B 0.03fF
C18126 POR2X1_264/Y POR2X1_260/B 0.04fF
C18127 POR2X1_257/A POR2X1_90/Y 0.07fF
C18128 POR2X1_673/A POR2X1_673/CTRL2 0.00fF
C18129 PAND2X1_860/A PAND2X1_716/B 0.03fF
C18130 PAND2X1_474/Y POR2X1_497/CTRL 0.00fF
C18131 POR2X1_490/a_16_28# POR2X1_73/Y 0.02fF
C18132 PAND2X1_213/CTRL2 PAND2X1_161/Y 0.03fF
C18133 PAND2X1_90/A PAND2X1_277/O 0.02fF
C18134 POR2X1_811/B POR2X1_596/Y 0.09fF
C18135 POR2X1_148/CTRL2 POR2X1_532/A 0.03fF
C18136 POR2X1_32/A PAND2X1_151/m4_208_n4# 0.08fF
C18137 PAND2X1_430/CTRL POR2X1_750/B 0.02fF
C18138 PAND2X1_73/Y POR2X1_445/O 0.02fF
C18139 POR2X1_476/O POR2X1_476/Y 0.00fF
C18140 POR2X1_667/Y POR2X1_293/Y 0.03fF
C18141 POR2X1_631/A PAND2X1_39/B 0.00fF
C18142 PAND2X1_282/CTRL PAND2X1_55/Y 0.03fF
C18143 POR2X1_251/Y POR2X1_102/Y 0.02fF
C18144 PAND2X1_195/O VDD 0.00fF
C18145 POR2X1_356/A POR2X1_241/B 0.01fF
C18146 POR2X1_54/Y POR2X1_750/O 0.03fF
C18147 PAND2X1_73/Y POR2X1_149/Y 0.03fF
C18148 POR2X1_68/A POR2X1_856/B 0.06fF
C18149 POR2X1_528/a_56_344# POR2X1_48/A 0.00fF
C18150 POR2X1_632/CTRL2 PAND2X1_88/Y 0.01fF
C18151 PAND2X1_46/CTRL INPUT_0 0.11fF
C18152 POR2X1_466/A POR2X1_732/CTRL 0.47fF
C18153 PAND2X1_736/Y POR2X1_32/A 0.01fF
C18154 POR2X1_174/B POR2X1_579/Y 0.01fF
C18155 PAND2X1_576/B POR2X1_52/Y 0.03fF
C18156 POR2X1_14/Y POR2X1_372/Y 0.03fF
C18157 PAND2X1_219/A POR2X1_7/B 1.61fF
C18158 POR2X1_693/a_16_28# POR2X1_83/B 0.03fF
C18159 PAND2X1_20/CTRL VDD -0.00fF
C18160 PAND2X1_296/O POR2X1_42/Y -0.00fF
C18161 POR2X1_61/Y VDD 1.70fF
C18162 POR2X1_5/Y POR2X1_372/O 0.02fF
C18163 PAND2X1_169/Y PAND2X1_714/CTRL2 0.00fF
C18164 PAND2X1_76/Y POR2X1_272/Y 3.80fF
C18165 POR2X1_264/Y PAND2X1_265/CTRL2 0.01fF
C18166 PAND2X1_58/A POR2X1_459/A 0.00fF
C18167 PAND2X1_6/A POR2X1_29/A 0.20fF
C18168 POR2X1_683/Y POR2X1_604/Y 0.31fF
C18169 PAND2X1_54/CTRL2 VDD -0.00fF
C18170 POR2X1_666/A VDD 0.03fF
C18171 D_INPUT_0 POR2X1_550/CTRL 0.01fF
C18172 POR2X1_177/Y VDD 0.21fF
C18173 PAND2X1_603/m4_208_n4# PAND2X1_604/m4_208_n4# 0.13fF
C18174 POR2X1_752/Y INPUT_5 0.09fF
C18175 POR2X1_20/B PAND2X1_722/CTRL2 0.01fF
C18176 PAND2X1_570/a_16_344# PAND2X1_577/Y 0.02fF
C18177 PAND2X1_360/O POR2X1_42/Y 0.03fF
C18178 POR2X1_730/CTRL2 POR2X1_330/Y 0.02fF
C18179 POR2X1_79/Y PAND2X1_363/Y 0.02fF
C18180 PAND2X1_641/Y POR2X1_63/Y 0.01fF
C18181 POR2X1_96/A PAND2X1_541/a_56_28# 0.00fF
C18182 PAND2X1_206/A PAND2X1_100/CTRL 0.01fF
C18183 POR2X1_355/A POR2X1_785/A 0.03fF
C18184 PAND2X1_811/a_76_28# PAND2X1_805/A 0.01fF
C18185 POR2X1_552/Y VDD 0.00fF
C18186 POR2X1_763/A POR2X1_46/Y 0.31fF
C18187 PAND2X1_655/Y PAND2X1_660/B 0.15fF
C18188 POR2X1_490/Y PAND2X1_723/A 0.01fF
C18189 PAND2X1_818/a_56_28# POR2X1_376/B 0.00fF
C18190 POR2X1_60/a_76_344# D_INPUT_0 0.02fF
C18191 POR2X1_66/A PAND2X1_305/CTRL2 0.00fF
C18192 PAND2X1_11/Y PAND2X1_69/A 0.03fF
C18193 PAND2X1_206/B POR2X1_4/Y 0.07fF
C18194 PAND2X1_96/B PAND2X1_39/CTRL 0.01fF
C18195 PAND2X1_675/A POR2X1_251/A 0.03fF
C18196 PAND2X1_20/A POR2X1_78/O 0.01fF
C18197 POR2X1_58/Y POR2X1_376/B 0.02fF
C18198 POR2X1_850/B POR2X1_804/A 0.03fF
C18199 POR2X1_29/Y POR2X1_14/Y 0.05fF
C18200 PAND2X1_63/m4_208_n4# POR2X1_66/A 0.08fF
C18201 PAND2X1_473/Y INPUT_0 0.07fF
C18202 PAND2X1_57/B POR2X1_770/A 0.00fF
C18203 POR2X1_590/A POR2X1_550/O 0.02fF
C18204 POR2X1_252/O POR2X1_5/Y 0.01fF
C18205 POR2X1_66/B POR2X1_712/A 0.03fF
C18206 POR2X1_567/B PAND2X1_315/CTRL 0.13fF
C18207 PAND2X1_675/A POR2X1_72/B 0.01fF
C18208 POR2X1_542/B PAND2X1_58/A 0.03fF
C18209 POR2X1_508/CTRL POR2X1_852/B 0.03fF
C18210 PAND2X1_23/Y PAND2X1_395/CTRL 0.00fF
C18211 PAND2X1_193/CTRL POR2X1_7/B 0.01fF
C18212 PAND2X1_469/B POR2X1_72/B 0.04fF
C18213 POR2X1_791/B PAND2X1_586/a_16_344# 0.03fF
C18214 PAND2X1_29/CTRL2 PAND2X1_41/B 0.01fF
C18215 POR2X1_486/B POR2X1_486/CTRL2 0.08fF
C18216 PAND2X1_95/B PAND2X1_588/CTRL 0.01fF
C18217 PAND2X1_41/B POR2X1_350/O 0.10fF
C18218 POR2X1_355/A PAND2X1_504/O 0.02fF
C18219 POR2X1_180/B POR2X1_856/B 0.03fF
C18220 POR2X1_566/A POR2X1_244/B 0.05fF
C18221 POR2X1_61/Y POR2X1_741/Y 0.15fF
C18222 PAND2X1_23/Y PAND2X1_58/CTRL2 0.00fF
C18223 PAND2X1_57/B POR2X1_76/Y 0.03fF
C18224 POR2X1_443/CTRL POR2X1_191/Y 0.11fF
C18225 POR2X1_443/O POR2X1_192/B 0.06fF
C18226 POR2X1_652/Y VDD 0.23fF
C18227 PAND2X1_65/B POR2X1_205/CTRL 0.01fF
C18228 PAND2X1_736/Y PAND2X1_741/B 0.01fF
C18229 PAND2X1_731/O PAND2X1_731/B 0.00fF
C18230 PAND2X1_65/B POR2X1_800/A 0.00fF
C18231 PAND2X1_661/O POR2X1_13/A 0.17fF
C18232 PAND2X1_644/CTRL2 POR2X1_236/Y 0.11fF
C18233 POR2X1_41/B PAND2X1_734/B 0.02fF
C18234 POR2X1_235/Y POR2X1_32/A 0.01fF
C18235 POR2X1_596/Y POR2X1_783/B 0.02fF
C18236 POR2X1_43/B POR2X1_278/O 0.04fF
C18237 PAND2X1_651/Y PAND2X1_456/CTRL 0.01fF
C18238 POR2X1_290/O PAND2X1_642/B 0.01fF
C18239 POR2X1_289/Y POR2X1_394/A 0.04fF
C18240 POR2X1_49/Y POR2X1_90/Y 0.30fF
C18241 POR2X1_433/Y POR2X1_432/Y 0.01fF
C18242 POR2X1_60/A POR2X1_239/Y 0.06fF
C18243 POR2X1_8/Y POR2X1_23/Y 0.03fF
C18244 POR2X1_20/B PAND2X1_338/CTRL 0.01fF
C18245 POR2X1_48/A POR2X1_764/CTRL 0.02fF
C18246 POR2X1_300/O POR2X1_272/Y 0.01fF
C18247 PAND2X1_137/CTRL POR2X1_96/A 0.01fF
C18248 POR2X1_110/Y POR2X1_257/A 0.06fF
C18249 PAND2X1_580/B POR2X1_42/Y 0.03fF
C18250 POR2X1_380/CTRL2 POR2X1_5/Y 0.01fF
C18251 POR2X1_515/CTRL2 POR2X1_68/A 0.16fF
C18252 POR2X1_122/Y POR2X1_43/B 0.00fF
C18253 POR2X1_548/a_16_28# PAND2X1_90/A 0.02fF
C18254 PAND2X1_552/B VDD 0.01fF
C18255 POR2X1_20/B PAND2X1_352/O 0.16fF
C18256 POR2X1_809/A POR2X1_676/a_76_344# 0.00fF
C18257 PAND2X1_41/B POR2X1_758/CTRL 0.01fF
C18258 PAND2X1_803/Y POR2X1_417/Y 0.02fF
C18259 POR2X1_687/A PAND2X1_73/Y 0.01fF
C18260 PAND2X1_793/Y POR2X1_293/Y 0.03fF
C18261 POR2X1_566/A POR2X1_562/CTRL 0.14fF
C18262 POR2X1_833/A POR2X1_499/a_76_344# 0.01fF
C18263 PAND2X1_470/CTRL PAND2X1_803/A 0.00fF
C18264 PAND2X1_57/B POR2X1_740/Y 0.11fF
C18265 PAND2X1_48/B PAND2X1_152/CTRL2 0.01fF
C18266 POR2X1_78/B POR2X1_407/A 0.18fF
C18267 PAND2X1_347/Y PAND2X1_357/Y 0.03fF
C18268 PAND2X1_673/CTRL2 POR2X1_38/B 0.01fF
C18269 POR2X1_218/Y POR2X1_244/Y 0.16fF
C18270 POR2X1_35/Y VDD 1.20fF
C18271 PAND2X1_262/a_16_344# POR2X1_38/B 0.02fF
C18272 POR2X1_614/A PAND2X1_129/O 0.01fF
C18273 POR2X1_71/Y POR2X1_72/Y 0.28fF
C18274 POR2X1_855/B POR2X1_783/CTRL 0.01fF
C18275 POR2X1_447/B POR2X1_629/CTRL2 0.05fF
C18276 POR2X1_119/Y PAND2X1_560/a_76_28# 0.05fF
C18277 POR2X1_668/a_16_28# PAND2X1_69/A 0.01fF
C18278 POR2X1_294/B PAND2X1_110/CTRL2 0.01fF
C18279 POR2X1_52/A PAND2X1_242/CTRL2 0.02fF
C18280 POR2X1_463/Y POR2X1_805/Y 0.03fF
C18281 PAND2X1_14/CTRL2 POR2X1_68/B 0.03fF
C18282 PAND2X1_862/Y POR2X1_23/Y 0.03fF
C18283 POR2X1_376/B POR2X1_9/CTRL 0.01fF
C18284 PAND2X1_65/B PAND2X1_26/O 0.02fF
C18285 POR2X1_156/B POR2X1_155/CTRL2 0.01fF
C18286 POR2X1_60/A POR2X1_534/Y 0.28fF
C18287 PAND2X1_80/CTRL2 POR2X1_68/B 0.00fF
C18288 PAND2X1_129/O POR2X1_38/B 0.05fF
C18289 POR2X1_68/A POR2X1_722/Y 0.03fF
C18290 POR2X1_334/Y POR2X1_97/A 0.12fF
C18291 POR2X1_23/Y POR2X1_385/Y 0.05fF
C18292 POR2X1_96/A POR2X1_255/Y 0.05fF
C18293 POR2X1_614/A POR2X1_724/a_56_344# 0.00fF
C18294 PAND2X1_73/Y POR2X1_558/Y 0.28fF
C18295 POR2X1_849/A POR2X1_550/B 0.04fF
C18296 PAND2X1_239/CTRL POR2X1_191/Y 0.10fF
C18297 PAND2X1_696/CTRL POR2X1_866/A 0.27fF
C18298 POR2X1_335/B VDD 0.21fF
C18299 POR2X1_245/Y POR2X1_5/Y 0.03fF
C18300 PAND2X1_6/Y POR2X1_247/CTRL2 -0.00fF
C18301 POR2X1_120/CTRL PAND2X1_60/B 0.01fF
C18302 POR2X1_387/Y POR2X1_236/Y 0.07fF
C18303 POR2X1_122/CTRL POR2X1_102/Y 0.01fF
C18304 POR2X1_800/A PAND2X1_599/O 0.00fF
C18305 POR2X1_516/Y POR2X1_129/Y 0.03fF
C18306 POR2X1_28/a_56_344# POR2X1_4/Y 0.00fF
C18307 POR2X1_7/B POR2X1_816/A 0.03fF
C18308 PAND2X1_6/Y POR2X1_783/B 0.02fF
C18309 POR2X1_819/m4_208_n4# POR2X1_523/m4_208_n4# 0.13fF
C18310 POR2X1_253/Y POR2X1_55/Y 0.18fF
C18311 POR2X1_530/Y VDD 0.04fF
C18312 POR2X1_327/Y POR2X1_830/CTRL 0.06fF
C18313 POR2X1_49/Y PAND2X1_732/A 0.03fF
C18314 POR2X1_65/A PAND2X1_714/Y 0.07fF
C18315 POR2X1_307/B POR2X1_796/A 4.68fF
C18316 POR2X1_35/Y POR2X1_741/Y 0.11fF
C18317 POR2X1_29/Y POR2X1_55/Y 0.04fF
C18318 POR2X1_78/B PAND2X1_315/CTRL 0.06fF
C18319 POR2X1_814/B POR2X1_463/Y 0.03fF
C18320 POR2X1_20/O POR2X1_38/B 0.00fF
C18321 POR2X1_123/A VDD 0.42fF
C18322 PAND2X1_865/Y POR2X1_487/CTRL 0.01fF
C18323 POR2X1_102/O POR2X1_37/Y 0.17fF
C18324 PAND2X1_212/CTRL POR2X1_77/Y 0.00fF
C18325 PAND2X1_649/A PAND2X1_400/O 0.02fF
C18326 POR2X1_599/A PAND2X1_717/a_56_28# 0.00fF
C18327 POR2X1_814/B POR2X1_756/Y 0.01fF
C18328 POR2X1_327/Y POR2X1_188/A 0.02fF
C18329 PAND2X1_480/B PAND2X1_175/B 0.05fF
C18330 POR2X1_689/A POR2X1_38/Y 0.01fF
C18331 PAND2X1_90/A POR2X1_68/B 3.94fF
C18332 PAND2X1_572/O PAND2X1_364/B 0.09fF
C18333 POR2X1_654/CTRL POR2X1_774/A 0.00fF
C18334 POR2X1_239/O POR2X1_55/Y 0.00fF
C18335 POR2X1_770/A POR2X1_707/Y 0.01fF
C18336 POR2X1_504/O POR2X1_504/Y 0.01fF
C18337 POR2X1_309/Y PAND2X1_337/A 0.03fF
C18338 POR2X1_343/Y POR2X1_260/B 0.03fF
C18339 POR2X1_856/B POR2X1_169/A 0.03fF
C18340 PAND2X1_658/B PAND2X1_174/m4_208_n4# 0.02fF
C18341 PAND2X1_368/O VDD -0.00fF
C18342 POR2X1_9/Y POR2X1_67/Y 0.03fF
C18343 POR2X1_389/A POR2X1_294/B 0.03fF
C18344 POR2X1_235/Y PAND2X1_35/Y 0.03fF
C18345 POR2X1_316/a_76_344# PAND2X1_390/Y -0.00fF
C18346 POR2X1_840/B PAND2X1_275/a_16_344# 0.02fF
C18347 POR2X1_55/Y POR2X1_9/O 0.04fF
C18348 PAND2X1_289/a_76_28# PAND2X1_52/B 0.02fF
C18349 POR2X1_771/A POR2X1_770/A 0.08fF
C18350 POR2X1_41/B PAND2X1_661/Y 0.00fF
C18351 PAND2X1_787/Y PAND2X1_348/A 0.10fF
C18352 PAND2X1_472/CTRL VDD 0.00fF
C18353 POR2X1_602/B POR2X1_722/O 0.01fF
C18354 PAND2X1_854/A POR2X1_7/B 0.04fF
C18355 POR2X1_335/B POR2X1_741/Y 0.03fF
C18356 POR2X1_532/A POR2X1_713/CTRL 0.06fF
C18357 POR2X1_518/Y POR2X1_73/Y 0.04fF
C18358 PAND2X1_96/B POR2X1_515/Y 0.01fF
C18359 POR2X1_252/Y POR2X1_482/Y 0.03fF
C18360 POR2X1_574/CTRL POR2X1_724/A 0.00fF
C18361 POR2X1_176/O POR2X1_312/Y 0.01fF
C18362 POR2X1_693/a_56_344# PAND2X1_550/B 0.00fF
C18363 POR2X1_158/Y POR2X1_48/A 0.00fF
C18364 PAND2X1_93/B POR2X1_325/B 0.05fF
C18365 PAND2X1_94/A POR2X1_121/Y 0.03fF
C18366 POR2X1_68/B PAND2X1_19/O 0.04fF
C18367 PAND2X1_784/O POR2X1_7/A 0.01fF
C18368 POR2X1_49/Y POR2X1_110/Y 0.07fF
C18369 POR2X1_445/CTRL2 POR2X1_456/B 0.00fF
C18370 PAND2X1_844/B POR2X1_56/Y 0.03fF
C18371 PAND2X1_653/CTRL2 POR2X1_83/B 0.01fF
C18372 PAND2X1_349/A POR2X1_42/Y 0.02fF
C18373 POR2X1_687/B POR2X1_687/A 0.02fF
C18374 POR2X1_840/O POR2X1_513/Y 0.00fF
C18375 PAND2X1_63/B POR2X1_42/Y 0.03fF
C18376 POR2X1_137/Y POR2X1_218/A 0.10fF
C18377 POR2X1_541/CTRL POR2X1_702/A 0.00fF
C18378 PAND2X1_615/CTRL D_INPUT_1 0.01fF
C18379 PAND2X1_696/CTRL2 POR2X1_602/B 0.01fF
C18380 POR2X1_542/B PAND2X1_96/B 0.14fF
C18381 POR2X1_724/O POR2X1_703/Y 0.02fF
C18382 PAND2X1_445/Y PAND2X1_308/Y 0.01fF
C18383 POR2X1_204/a_16_28# POR2X1_84/Y 0.05fF
C18384 POR2X1_140/A POR2X1_318/A 0.03fF
C18385 POR2X1_326/A POR2X1_480/A 0.07fF
C18386 PAND2X1_736/m4_208_n4# PAND2X1_853/B 0.15fF
C18387 PAND2X1_96/B PAND2X1_79/Y 0.06fF
C18388 POR2X1_383/A POR2X1_341/CTRL 0.03fF
C18389 POR2X1_357/a_16_28# POR2X1_353/Y -0.00fF
C18390 PAND2X1_56/Y POR2X1_274/B 0.03fF
C18391 PAND2X1_90/A POR2X1_561/O 0.01fF
C18392 PAND2X1_48/B POR2X1_151/O 0.03fF
C18393 PAND2X1_209/A PAND2X1_797/CTRL2 0.01fF
C18394 POR2X1_416/B POR2X1_487/a_16_28# 0.02fF
C18395 POR2X1_9/Y POR2X1_818/CTRL2 0.04fF
C18396 PAND2X1_96/B POR2X1_736/O 0.01fF
C18397 POR2X1_525/Y PAND2X1_726/B 0.06fF
C18398 POR2X1_65/A PAND2X1_865/Y 0.07fF
C18399 D_INPUT_1 PAND2X1_60/B 0.07fF
C18400 POR2X1_377/CTRL PAND2X1_94/A 0.00fF
C18401 POR2X1_861/O POR2X1_101/Y 0.03fF
C18402 POR2X1_255/Y POR2X1_7/A 0.03fF
C18403 POR2X1_686/B POR2X1_809/A 0.63fF
C18404 PAND2X1_20/A POR2X1_736/A 0.02fF
C18405 POR2X1_93/A POR2X1_382/Y 0.59fF
C18406 POR2X1_741/Y PAND2X1_368/O 0.04fF
C18407 PAND2X1_422/CTRL2 POR2X1_788/B 0.03fF
C18408 PAND2X1_57/B POR2X1_774/A 0.03fF
C18409 POR2X1_277/CTRL2 PAND2X1_560/B 0.03fF
C18410 POR2X1_760/Y POR2X1_595/Y 0.07fF
C18411 D_INPUT_3 POR2X1_9/CTRL2 0.14fF
C18412 PAND2X1_735/a_76_28# POR2X1_153/Y 0.02fF
C18413 POR2X1_78/A POR2X1_325/B 0.02fF
C18414 PAND2X1_593/CTRL POR2X1_385/Y 0.01fF
C18415 D_INPUT_3 PAND2X1_509/a_16_344# 0.00fF
C18416 POR2X1_13/A POR2X1_371/CTRL2 0.00fF
C18417 PAND2X1_625/CTRL2 POR2X1_260/A 0.10fF
C18418 POR2X1_537/Y POR2X1_130/A 0.05fF
C18419 POR2X1_123/A PAND2X1_32/B 0.03fF
C18420 POR2X1_245/a_16_28# POR2X1_90/Y 0.03fF
C18421 POR2X1_383/A POR2X1_649/CTRL 0.01fF
C18422 POR2X1_333/A POR2X1_168/A 0.06fF
C18423 POR2X1_241/B PAND2X1_72/A 0.06fF
C18424 PAND2X1_60/B POR2X1_724/A 0.03fF
C18425 D_GATE_662 POR2X1_353/A 0.03fF
C18426 POR2X1_32/A POR2X1_387/m4_208_n4# 0.01fF
C18427 POR2X1_49/a_16_28# POR2X1_37/Y 0.03fF
C18428 POR2X1_143/CTRL2 PAND2X1_341/B 0.02fF
C18429 PAND2X1_841/CTRL POR2X1_153/Y 0.01fF
C18430 PAND2X1_20/A POR2X1_500/O 0.01fF
C18431 POR2X1_88/CTRL POR2X1_9/Y 0.01fF
C18432 PAND2X1_57/B PAND2X1_328/CTRL 0.01fF
C18433 PAND2X1_737/O VDD 0.00fF
C18434 PAND2X1_473/B POR2X1_589/CTRL2 0.01fF
C18435 POR2X1_68/A POR2X1_799/a_16_28# 0.08fF
C18436 POR2X1_16/A POR2X1_234/O 0.01fF
C18437 POR2X1_334/Y POR2X1_294/B 0.07fF
C18438 POR2X1_719/A PAND2X1_72/A 0.00fF
C18439 POR2X1_355/B POR2X1_337/Y 0.23fF
C18440 POR2X1_101/Y POR2X1_500/Y 0.05fF
C18441 PAND2X1_69/A PAND2X1_133/O 0.03fF
C18442 POR2X1_416/B POR2X1_423/Y 0.03fF
C18443 POR2X1_101/Y PAND2X1_150/CTRL 0.13fF
C18444 POR2X1_96/B D_INPUT_3 0.03fF
C18445 POR2X1_394/A PAND2X1_188/a_76_28# 0.03fF
C18446 POR2X1_814/B POR2X1_736/A 0.05fF
C18447 PAND2X1_552/B PAND2X1_703/CTRL 0.01fF
C18448 POR2X1_862/CTRL2 POR2X1_480/A 0.03fF
C18449 POR2X1_13/Y PAND2X1_538/a_16_344# 0.02fF
C18450 POR2X1_119/Y POR2X1_406/O 0.26fF
C18451 PAND2X1_118/a_56_28# POR2X1_559/A 0.00fF
C18452 POR2X1_43/B PAND2X1_508/Y 0.03fF
C18453 POR2X1_130/CTRL2 POR2X1_318/A 0.01fF
C18454 PAND2X1_300/O PAND2X1_60/B 0.02fF
C18455 POR2X1_65/A PAND2X1_326/O 0.01fF
C18456 PAND2X1_850/Y POR2X1_46/Y 0.10fF
C18457 POR2X1_150/Y POR2X1_411/B 0.38fF
C18458 PAND2X1_140/A PAND2X1_346/Y 0.03fF
C18459 POR2X1_684/Y POR2X1_42/Y 0.01fF
C18460 POR2X1_96/A POR2X1_189/CTRL2 0.01fF
C18461 PAND2X1_525/O PAND2X1_52/B 0.02fF
C18462 POR2X1_549/O PAND2X1_52/B 0.04fF
C18463 PAND2X1_630/a_16_344# PAND2X1_156/A 0.06fF
C18464 PAND2X1_824/B POR2X1_98/B 0.53fF
C18465 POR2X1_105/Y PAND2X1_72/A 0.01fF
C18466 POR2X1_485/a_16_28# POR2X1_102/Y 0.03fF
C18467 POR2X1_407/A POR2X1_294/A 0.13fF
C18468 POR2X1_583/O POR2X1_583/Y 0.01fF
C18469 PAND2X1_610/O POR2X1_293/Y 0.02fF
C18470 POR2X1_343/Y POR2X1_723/O 0.02fF
C18471 POR2X1_669/B POR2X1_827/CTRL2 0.01fF
C18472 POR2X1_566/A POR2X1_555/CTRL 0.01fF
C18473 PAND2X1_734/B POR2X1_77/Y 0.01fF
C18474 PAND2X1_865/Y PAND2X1_190/Y 0.10fF
C18475 POR2X1_271/A POR2X1_387/Y 0.05fF
C18476 POR2X1_73/Y PAND2X1_325/O 0.02fF
C18477 POR2X1_137/Y POR2X1_557/B 0.01fF
C18478 POR2X1_373/Y POR2X1_142/Y 0.03fF
C18479 PAND2X1_335/CTRL2 POR2X1_77/Y 0.01fF
C18480 PAND2X1_652/O PAND2X1_652/A 0.06fF
C18481 POR2X1_391/m4_208_n4# POR2X1_260/A 0.15fF
C18482 POR2X1_493/CTRL2 PAND2X1_48/A 0.00fF
C18483 POR2X1_529/Y POR2X1_384/A 0.03fF
C18484 POR2X1_43/CTRL2 POR2X1_42/Y 0.01fF
C18485 POR2X1_540/A POR2X1_552/a_76_344# 0.01fF
C18486 POR2X1_249/Y POR2X1_734/O 0.01fF
C18487 POR2X1_778/a_16_28# POR2X1_717/B 0.02fF
C18488 PAND2X1_438/CTRL2 PAND2X1_72/A 0.00fF
C18489 POR2X1_190/CTRL POR2X1_188/Y 0.01fF
C18490 PAND2X1_476/A PAND2X1_734/O 0.00fF
C18491 POR2X1_333/Y POR2X1_351/O 0.06fF
C18492 POR2X1_698/Y POR2X1_763/A 0.01fF
C18493 POR2X1_260/A POR2X1_156/Y 0.00fF
C18494 PAND2X1_467/Y POR2X1_394/A 0.03fF
C18495 PAND2X1_813/O POR2X1_673/Y 0.02fF
C18496 POR2X1_647/B POR2X1_643/Y 0.02fF
C18497 POR2X1_164/Y POR2X1_165/Y 0.02fF
C18498 POR2X1_494/Y POR2X1_80/CTRL2 0.00fF
C18499 POR2X1_246/O POR2X1_39/B 0.01fF
C18500 POR2X1_416/B POR2X1_57/Y 0.06fF
C18501 PAND2X1_94/A POR2X1_54/CTRL2 0.00fF
C18502 POR2X1_783/B PAND2X1_52/B 0.06fF
C18503 POR2X1_260/B POR2X1_624/Y 0.11fF
C18504 POR2X1_130/CTRL2 POR2X1_574/Y 0.09fF
C18505 POR2X1_67/Y PAND2X1_225/CTRL2 0.12fF
C18506 POR2X1_458/Y POR2X1_750/B 0.17fF
C18507 POR2X1_192/B POR2X1_577/m4_208_n4# 0.06fF
C18508 PAND2X1_557/A POR2X1_329/A 0.12fF
C18509 POR2X1_613/Y POR2X1_408/Y 0.05fF
C18510 POR2X1_773/B POR2X1_768/Y 0.03fF
C18511 POR2X1_432/CTRL POR2X1_271/B 0.01fF
C18512 POR2X1_390/B PAND2X1_48/A 0.03fF
C18513 POR2X1_68/A PAND2X1_681/CTRL2 0.10fF
C18514 PAND2X1_826/CTRL2 POR2X1_294/Y 0.00fF
C18515 PAND2X1_575/A PAND2X1_332/Y 0.03fF
C18516 POR2X1_362/Y POR2X1_556/A 0.01fF
C18517 POR2X1_539/O POR2X1_537/Y 0.00fF
C18518 POR2X1_334/a_16_28# POR2X1_334/A 0.03fF
C18519 PAND2X1_479/CTRL POR2X1_329/A 0.01fF
C18520 POR2X1_416/B POR2X1_136/a_16_28# 0.03fF
C18521 POR2X1_119/Y PAND2X1_301/CTRL2 0.01fF
C18522 PAND2X1_301/a_16_344# PAND2X1_716/B 0.02fF
C18523 POR2X1_505/CTRL PAND2X1_631/A 0.01fF
C18524 PAND2X1_319/B POR2X1_416/B 0.17fF
C18525 POR2X1_333/Y POR2X1_502/Y 0.17fF
C18526 PAND2X1_425/Y PAND2X1_582/CTRL 0.01fF
C18527 PAND2X1_405/CTRL2 POR2X1_46/Y 0.01fF
C18528 POR2X1_813/a_16_28# POR2X1_32/A 0.02fF
C18529 POR2X1_861/A POR2X1_244/Y 0.10fF
C18530 POR2X1_505/Y POR2X1_20/B 0.01fF
C18531 POR2X1_647/CTRL POR2X1_296/B 0.44fF
C18532 POR2X1_820/a_76_344# POR2X1_411/B 0.01fF
C18533 POR2X1_141/Y POR2X1_276/B 0.02fF
C18534 PAND2X1_458/O POR2X1_372/Y 0.02fF
C18535 PAND2X1_661/Y POR2X1_77/Y 0.03fF
C18536 POR2X1_567/A POR2X1_334/Y 0.10fF
C18537 PAND2X1_479/A POR2X1_329/A 0.02fF
C18538 PAND2X1_419/CTRL POR2X1_296/B 0.01fF
C18539 PAND2X1_267/O POR2X1_102/Y 0.04fF
C18540 POR2X1_54/Y POR2X1_389/Y 0.03fF
C18541 POR2X1_333/A POR2X1_478/a_16_28# 0.05fF
C18542 POR2X1_799/CTRL2 PAND2X1_72/A 0.01fF
C18543 POR2X1_302/m4_208_n4# POR2X1_284/m4_208_n4# 0.13fF
C18544 POR2X1_431/Y POR2X1_236/Y 0.03fF
C18545 POR2X1_420/O POR2X1_102/Y 0.01fF
C18546 PAND2X1_613/O PAND2X1_41/B 0.03fF
C18547 PAND2X1_404/Y PAND2X1_500/O 0.05fF
C18548 POR2X1_566/A POR2X1_443/CTRL2 0.09fF
C18549 POR2X1_681/Y POR2X1_682/CTRL 0.01fF
C18550 PAND2X1_98/CTRL VDD -0.00fF
C18551 POR2X1_707/B PAND2X1_25/CTRL2 0.01fF
C18552 POR2X1_83/B POR2X1_496/Y 2.79fF
C18553 POR2X1_814/A POR2X1_800/A 0.05fF
C18554 POR2X1_603/Y POR2X1_669/B 0.03fF
C18555 POR2X1_12/A POR2X1_2/CTRL2 0.01fF
C18556 POR2X1_860/O PAND2X1_72/A 0.02fF
C18557 POR2X1_424/Y VDD 0.05fF
C18558 POR2X1_174/B POR2X1_590/A 0.03fF
C18559 POR2X1_91/a_16_28# POR2X1_91/Y 0.02fF
C18560 POR2X1_257/A INPUT_0 0.15fF
C18561 POR2X1_32/A PAND2X1_719/Y 0.24fF
C18562 PAND2X1_571/A PAND2X1_576/CTRL 0.01fF
C18563 POR2X1_52/A POR2X1_150/Y 0.18fF
C18564 POR2X1_830/CTRL2 POR2X1_590/A 0.03fF
C18565 POR2X1_270/Y POR2X1_814/B 0.03fF
C18566 POR2X1_24/O POR2X1_409/B 0.02fF
C18567 POR2X1_496/Y POR2X1_626/Y 0.02fF
C18568 POR2X1_411/B PAND2X1_364/B 0.08fF
C18569 POR2X1_78/B PAND2X1_601/a_16_344# 0.02fF
C18570 POR2X1_484/Y POR2X1_763/Y 0.16fF
C18571 POR2X1_703/a_16_28# POR2X1_169/A 0.05fF
C18572 POR2X1_814/A POR2X1_702/A 0.73fF
C18573 POR2X1_446/B POR2X1_724/CTRL 0.01fF
C18574 INPUT_3 POR2X1_7/B 0.27fF
C18575 POR2X1_150/Y POR2X1_152/A 0.04fF
C18576 POR2X1_809/A PAND2X1_681/CTRL 0.01fF
C18577 PAND2X1_586/O PAND2X1_72/A 0.03fF
C18578 POR2X1_496/Y POR2X1_752/Y 2.83fF
C18579 POR2X1_72/B POR2X1_498/Y 0.02fF
C18580 POR2X1_405/O POR2X1_296/B 0.04fF
C18581 POR2X1_850/A D_INPUT_0 0.03fF
C18582 POR2X1_850/B POR2X1_794/B 0.03fF
C18583 POR2X1_83/B PAND2X1_733/A 0.03fF
C18584 POR2X1_504/Y POR2X1_669/B 0.00fF
C18585 D_INPUT_0 POR2X1_5/Y 7.05fF
C18586 POR2X1_399/A POR2X1_20/B 0.01fF
C18587 POR2X1_634/A POR2X1_792/m4_208_n4# 0.06fF
C18588 POR2X1_347/B POR2X1_202/A 0.04fF
C18589 PAND2X1_268/O POR2X1_193/A 0.01fF
C18590 PAND2X1_464/B PAND2X1_785/CTRL 0.02fF
C18591 PAND2X1_793/Y POR2X1_67/CTRL 0.01fF
C18592 POR2X1_814/B POR2X1_288/O 0.01fF
C18593 POR2X1_496/O POR2X1_55/Y 0.01fF
C18594 POR2X1_55/CTRL POR2X1_5/Y 0.01fF
C18595 POR2X1_260/B INPUT_4 0.03fF
C18596 POR2X1_555/A POR2X1_590/A 0.03fF
C18597 PAND2X1_55/Y POR2X1_624/Y 0.03fF
C18598 POR2X1_20/B PAND2X1_546/CTRL 0.01fF
C18599 PAND2X1_58/A PAND2X1_395/CTRL2 0.01fF
C18600 PAND2X1_793/CTRL POR2X1_29/A 0.01fF
C18601 POR2X1_163/Y PAND2X1_725/B 0.02fF
C18602 POR2X1_705/B PAND2X1_69/A 0.05fF
C18603 POR2X1_446/B POR2X1_659/CTRL2 0.01fF
C18604 PAND2X1_73/Y POR2X1_455/CTRL 0.01fF
C18605 POR2X1_856/B POR2X1_435/Y 0.02fF
C18606 POR2X1_83/B PAND2X1_180/CTRL2 0.03fF
C18607 PAND2X1_217/B PAND2X1_476/CTRL 0.27fF
C18608 POR2X1_864/A POR2X1_532/A 0.00fF
C18609 POR2X1_260/B PAND2X1_536/CTRL2 0.01fF
C18610 POR2X1_138/O POR2X1_260/B 0.01fF
C18611 POR2X1_20/B PAND2X1_785/O 0.05fF
C18612 POR2X1_750/B PAND2X1_52/Y 0.05fF
C18613 PAND2X1_615/CTRL INPUT_3 0.06fF
C18614 PAND2X1_473/Y POR2X1_102/Y 0.03fF
C18615 POR2X1_68/A POR2X1_866/A 0.25fF
C18616 POR2X1_32/A POR2X1_817/A 0.03fF
C18617 PAND2X1_78/CTRL PAND2X1_580/B 0.00fF
C18618 PAND2X1_429/CTRL INPUT_5 0.01fF
C18619 POR2X1_682/Y POR2X1_60/A 0.02fF
C18620 POR2X1_35/B POR2X1_621/B 0.01fF
C18621 POR2X1_760/A POR2X1_385/O 0.00fF
C18622 POR2X1_71/Y POR2X1_32/A 0.07fF
C18623 PAND2X1_93/a_16_344# PAND2X1_93/B 0.02fF
C18624 POR2X1_814/A POR2X1_768/O 0.03fF
C18625 POR2X1_812/O POR2X1_121/B -0.02fF
C18626 POR2X1_428/Y PAND2X1_711/O 0.17fF
C18627 POR2X1_20/A POR2X1_38/B 0.00fF
C18628 POR2X1_748/A VDD 2.34fF
C18629 PAND2X1_58/A POR2X1_722/Y 0.08fF
C18630 PAND2X1_48/B POR2X1_269/O 0.01fF
C18631 POR2X1_861/CTRL POR2X1_218/Y 0.05fF
C18632 PAND2X1_613/CTRL POR2X1_68/B 0.00fF
C18633 POR2X1_477/O POR2X1_854/B 0.01fF
C18634 POR2X1_377/O D_INPUT_0 0.01fF
C18635 PAND2X1_6/Y PAND2X1_258/CTRL 0.01fF
C18636 PAND2X1_793/Y POR2X1_60/A 0.07fF
C18637 POR2X1_32/A POR2X1_42/Y 0.20fF
C18638 POR2X1_21/O D_INPUT_5 0.01fF
C18639 POR2X1_56/B POR2X1_420/Y 0.02fF
C18640 POR2X1_54/Y POR2X1_713/B 0.06fF
C18641 PAND2X1_668/a_76_28# POR2X1_83/B 0.02fF
C18642 POR2X1_62/CTRL2 PAND2X1_58/A 0.04fF
C18643 POR2X1_49/Y INPUT_0 2.18fF
C18644 PAND2X1_631/O POR2X1_48/A 0.04fF
C18645 POR2X1_556/A PAND2X1_368/a_16_344# 0.02fF
C18646 PAND2X1_632/B POR2X1_20/B 0.01fF
C18647 POR2X1_459/O POR2X1_750/B 0.01fF
C18648 POR2X1_28/a_56_344# D_INPUT_1 0.01fF
C18649 PAND2X1_308/B POR2X1_306/Y 0.05fF
C18650 PAND2X1_58/A POR2X1_791/O 0.17fF
C18651 PAND2X1_295/O PAND2X1_60/B 0.02fF
C18652 PAND2X1_649/A POR2X1_689/a_16_28# 0.02fF
C18653 POR2X1_376/B POR2X1_701/Y 0.03fF
C18654 POR2X1_302/B PAND2X1_322/CTRL 0.01fF
C18655 POR2X1_856/B PAND2X1_96/B 0.03fF
C18656 PAND2X1_513/a_16_344# PAND2X1_512/Y 0.02fF
C18657 PAND2X1_48/B POR2X1_634/A 0.12fF
C18658 PAND2X1_39/B POR2X1_101/Y 0.15fF
C18659 PAND2X1_90/CTRL2 POR2X1_814/A 0.01fF
C18660 POR2X1_356/A POR2X1_436/CTRL 0.01fF
C18661 POR2X1_290/a_16_28# POR2X1_236/Y 0.02fF
C18662 POR2X1_218/Y POR2X1_501/B 0.07fF
C18663 PAND2X1_159/a_56_28# POR2X1_7/B 0.00fF
C18664 PAND2X1_6/Y POR2X1_296/B 0.18fF
C18665 POR2X1_65/A POR2X1_424/CTRL2 0.11fF
C18666 POR2X1_66/A POR2X1_194/O 0.01fF
C18667 PAND2X1_90/A PAND2X1_73/O 0.01fF
C18668 POR2X1_655/A POR2X1_725/Y 0.01fF
C18669 PAND2X1_93/B PAND2X1_60/B 10.26fF
C18670 PAND2X1_740/a_56_28# PAND2X1_738/Y 0.00fF
C18671 PAND2X1_58/A POR2X1_565/O 0.01fF
C18672 PAND2X1_644/Y POR2X1_757/O 0.08fF
C18673 POR2X1_590/A POR2X1_705/O 0.02fF
C18674 PAND2X1_206/B PAND2X1_101/B 0.01fF
C18675 PAND2X1_20/A PAND2X1_6/A 0.45fF
C18676 POR2X1_49/Y POR2X1_617/O 0.03fF
C18677 POR2X1_48/A PAND2X1_348/Y 0.03fF
C18678 PAND2X1_621/Y POR2X1_847/B 0.61fF
C18679 POR2X1_840/B PAND2X1_73/Y 0.21fF
C18680 PAND2X1_575/B POR2X1_184/Y 0.00fF
C18681 PAND2X1_770/CTRL VDD -0.00fF
C18682 PAND2X1_689/a_16_344# PAND2X1_32/B 0.01fF
C18683 POR2X1_670/CTRL2 POR2X1_42/Y 0.01fF
C18684 PAND2X1_480/B POR2X1_272/Y 0.14fF
C18685 POR2X1_178/O POR2X1_60/A 0.01fF
C18686 POR2X1_41/B POR2X1_144/Y 0.12fF
C18687 POR2X1_79/A VDD 0.13fF
C18688 POR2X1_489/B PAND2X1_69/A 0.02fF
C18689 PAND2X1_860/A PAND2X1_862/CTRL 0.01fF
C18690 POR2X1_417/Y POR2X1_309/Y 0.03fF
C18691 POR2X1_219/B PAND2X1_394/CTRL 0.03fF
C18692 POR2X1_800/a_16_28# POR2X1_800/A 0.03fF
C18693 POR2X1_16/A PAND2X1_404/Y 0.01fF
C18694 POR2X1_573/O POR2X1_404/Y 0.02fF
C18695 PAND2X1_849/O PAND2X1_859/B 0.02fF
C18696 POR2X1_97/A POR2X1_212/CTRL2 0.03fF
C18697 POR2X1_60/A PAND2X1_711/A 0.02fF
C18698 POR2X1_460/B POR2X1_752/Y 0.25fF
C18699 POR2X1_511/Y POR2X1_372/Y 0.07fF
C18700 POR2X1_296/B POR2X1_575/CTRL2 0.01fF
C18701 PAND2X1_468/CTRL2 VDD 0.00fF
C18702 POR2X1_628/Y POR2X1_129/Y 0.27fF
C18703 POR2X1_614/A PAND2X1_582/CTRL 0.01fF
C18704 PAND2X1_659/B PAND2X1_735/Y 0.11fF
C18705 PAND2X1_58/A PAND2X1_757/CTRL2 0.00fF
C18706 PAND2X1_394/O PAND2X1_88/Y 0.02fF
C18707 POR2X1_750/B POR2X1_816/A 0.03fF
C18708 POR2X1_435/Y POR2X1_722/Y 0.06fF
C18709 PAND2X1_90/A PAND2X1_80/CTRL2 0.03fF
C18710 POR2X1_78/A PAND2X1_60/B 0.18fF
C18711 POR2X1_13/A PAND2X1_668/CTRL2 0.01fF
C18712 POR2X1_278/Y POR2X1_251/Y 0.06fF
C18713 POR2X1_537/O POR2X1_260/B 0.04fF
C18714 POR2X1_706/CTRL2 POR2X1_383/A 0.01fF
C18715 POR2X1_440/Y POR2X1_434/A 0.01fF
C18716 PAND2X1_90/Y PAND2X1_145/CTRL 0.01fF
C18717 POR2X1_219/B POR2X1_330/Y 0.07fF
C18718 POR2X1_750/B D_INPUT_1 0.11fF
C18719 POR2X1_96/A POR2X1_693/CTRL 0.00fF
C18720 POR2X1_322/a_76_344# POR2X1_376/B 0.01fF
C18721 POR2X1_356/A POR2X1_781/O 0.03fF
C18722 PAND2X1_93/B POR2X1_353/A 0.03fF
C18723 POR2X1_29/O POR2X1_55/Y 0.18fF
C18724 POR2X1_814/B PAND2X1_6/A 6.53fF
C18725 PAND2X1_41/B PAND2X1_518/CTRL2 0.00fF
C18726 POR2X1_13/O POR2X1_7/B 0.02fF
C18727 PAND2X1_94/A PAND2X1_282/CTRL2 0.02fF
C18728 POR2X1_96/A POR2X1_46/Y 0.03fF
C18729 PAND2X1_786/CTRL POR2X1_91/Y 0.06fF
C18730 POR2X1_186/Y POR2X1_556/Y 0.03fF
C18731 POR2X1_57/A PAND2X1_557/A 0.03fF
C18732 POR2X1_444/A POR2X1_545/CTRL 0.07fF
C18733 PAND2X1_48/B POR2X1_130/A 0.10fF
C18734 PAND2X1_56/Y POR2X1_483/A 0.03fF
C18735 POR2X1_260/B POR2X1_186/B 1.21fF
C18736 PAND2X1_423/O POR2X1_804/A 0.29fF
C18737 PAND2X1_467/Y POR2X1_669/B 0.07fF
C18738 POR2X1_631/A POR2X1_200/O 0.01fF
C18739 PAND2X1_90/A POR2X1_243/Y 0.00fF
C18740 D_INPUT_0 POR2X1_576/O 0.01fF
C18741 POR2X1_750/B POR2X1_724/A 0.10fF
C18742 PAND2X1_787/Y POR2X1_183/Y 0.05fF
C18743 POR2X1_368/Y PAND2X1_76/Y 0.06fF
C18744 PAND2X1_269/m4_208_n4# POR2X1_39/B 0.15fF
C18745 INPUT_1 PAND2X1_623/CTRL2 0.01fF
C18746 PAND2X1_48/B POR2X1_566/A 0.04fF
C18747 PAND2X1_644/Y POR2X1_394/A 0.19fF
C18748 POR2X1_52/A PAND2X1_364/B 0.02fF
C18749 POR2X1_253/Y POR2X1_511/Y 0.01fF
C18750 POR2X1_567/A POR2X1_854/CTRL 0.04fF
C18751 PAND2X1_162/O VDD 0.00fF
C18752 PAND2X1_61/Y POR2X1_38/Y 0.05fF
C18753 PAND2X1_865/CTRL POR2X1_102/Y 0.01fF
C18754 PAND2X1_381/Y POR2X1_391/B 0.01fF
C18755 PAND2X1_570/CTRL2 VDD 0.00fF
C18756 POR2X1_439/Y POR2X1_540/A 0.04fF
C18757 PAND2X1_6/Y POR2X1_464/CTRL 0.01fF
C18758 POR2X1_45/Y PAND2X1_274/CTRL 0.01fF
C18759 POR2X1_302/CTRL POR2X1_513/Y 0.00fF
C18760 PAND2X1_829/CTRL2 POR2X1_260/A 0.01fF
C18761 PAND2X1_803/A POR2X1_73/Y 0.03fF
C18762 PAND2X1_20/A POR2X1_101/Y 0.05fF
C18763 POR2X1_306/Y POR2X1_239/Y 0.00fF
C18764 POR2X1_330/Y POR2X1_366/A 0.05fF
C18765 PAND2X1_140/A PAND2X1_354/A 0.03fF
C18766 POR2X1_302/Y POR2X1_68/A 0.02fF
C18767 POR2X1_136/Y POR2X1_423/Y 0.38fF
C18768 PAND2X1_91/O POR2X1_192/B 0.16fF
C18769 PAND2X1_91/CTRL2 POR2X1_191/Y 0.00fF
C18770 POR2X1_685/CTRL2 POR2X1_685/B 0.03fF
C18771 PAND2X1_7/Y POR2X1_228/Y 0.12fF
C18772 POR2X1_111/CTRL POR2X1_5/Y 0.01fF
C18773 PAND2X1_627/CTRL PAND2X1_69/A 0.00fF
C18774 POR2X1_297/m4_208_n4# PAND2X1_359/m4_208_n4# 0.13fF
C18775 POR2X1_596/A PAND2X1_65/B 0.06fF
C18776 POR2X1_304/a_76_344# POR2X1_90/Y 0.00fF
C18777 POR2X1_809/A POR2X1_678/Y 0.02fF
C18778 PAND2X1_659/Y PAND2X1_267/Y 0.03fF
C18779 POR2X1_119/Y PAND2X1_444/CTRL 0.00fF
C18780 POR2X1_783/O POR2X1_796/A 0.01fF
C18781 POR2X1_78/A POR2X1_353/A 0.00fF
C18782 PAND2X1_848/A POR2X1_7/B 0.10fF
C18783 POR2X1_851/a_16_28# POR2X1_851/A 0.11fF
C18784 PAND2X1_855/a_16_344# POR2X1_236/Y 0.00fF
C18785 PAND2X1_460/O POR2X1_5/Y 0.09fF
C18786 POR2X1_265/Y POR2X1_23/Y 0.03fF
C18787 POR2X1_41/B PAND2X1_852/O 0.04fF
C18788 POR2X1_835/B PAND2X1_52/B 0.01fF
C18789 PAND2X1_569/B POR2X1_40/Y 0.11fF
C18790 POR2X1_40/Y POR2X1_158/B 0.06fF
C18791 PAND2X1_675/A POR2X1_7/B 0.03fF
C18792 POR2X1_254/Y POR2X1_804/A 0.02fF
C18793 PAND2X1_55/Y PAND2X1_536/CTRL2 -0.01fF
C18794 POR2X1_356/A D_GATE_741 0.03fF
C18795 PAND2X1_484/CTRL POR2X1_590/A 0.01fF
C18796 POR2X1_836/CTRL2 POR2X1_192/B 0.07fF
C18797 POR2X1_383/A POR2X1_287/B 0.03fF
C18798 PAND2X1_469/B POR2X1_7/B 0.05fF
C18799 POR2X1_174/CTRL2 POR2X1_175/A 0.01fF
C18800 POR2X1_41/B PAND2X1_546/O 0.04fF
C18801 D_INPUT_3 POR2X1_236/Y 0.10fF
C18802 POR2X1_260/Y POR2X1_205/CTRL 0.00fF
C18803 POR2X1_291/Y VDD 0.12fF
C18804 PAND2X1_217/CTRL2 INPUT_0 0.01fF
C18805 PAND2X1_499/O POR2X1_283/A 0.02fF
C18806 POR2X1_631/A VDD 0.06fF
C18807 POR2X1_51/A POR2X1_36/CTRL 0.01fF
C18808 PAND2X1_549/a_76_28# POR2X1_531/Y 0.05fF
C18809 POR2X1_814/B POR2X1_101/Y 0.34fF
C18810 POR2X1_71/Y PAND2X1_651/Y 0.05fF
C18811 PAND2X1_319/B PAND2X1_738/Y 0.10fF
C18812 PAND2X1_206/A PAND2X1_358/O 0.01fF
C18813 PAND2X1_492/O PAND2X1_60/B 0.02fF
C18814 PAND2X1_724/B PAND2X1_357/Y 0.02fF
C18815 POR2X1_184/Y POR2X1_42/Y 0.02fF
C18816 PAND2X1_674/O POR2X1_732/B 0.16fF
C18817 POR2X1_483/A POR2X1_383/A 0.04fF
C18818 POR2X1_752/Y PAND2X1_376/O 0.07fF
C18819 POR2X1_417/CTRL2 POR2X1_372/Y 0.05fF
C18820 POR2X1_667/A PAND2X1_123/Y 0.05fF
C18821 PAND2X1_860/A POR2X1_329/A 0.03fF
C18822 POR2X1_369/a_16_28# POR2X1_83/B 0.02fF
C18823 POR2X1_237/Y PAND2X1_445/CTRL 0.01fF
C18824 PAND2X1_657/O PAND2X1_657/B 0.00fF
C18825 POR2X1_43/B PAND2X1_228/a_56_28# 0.00fF
C18826 PAND2X1_11/Y PAND2X1_3/B 0.06fF
C18827 PAND2X1_651/Y POR2X1_42/Y 0.03fF
C18828 POR2X1_66/A PAND2X1_179/CTRL 0.00fF
C18829 POR2X1_675/A POR2X1_456/B 0.00fF
C18830 POR2X1_119/Y PAND2X1_446/O 0.01fF
C18831 POR2X1_614/A POR2X1_563/Y 0.03fF
C18832 POR2X1_383/A PAND2X1_8/Y 0.11fF
C18833 PAND2X1_308/O POR2X1_306/Y 0.10fF
C18834 POR2X1_795/O PAND2X1_32/B 0.01fF
C18835 POR2X1_729/CTRL POR2X1_614/A 0.01fF
C18836 PAND2X1_349/A PAND2X1_139/Y 0.01fF
C18837 PAND2X1_65/B POR2X1_598/O 0.01fF
C18838 POR2X1_614/A PAND2X1_599/a_16_344# 0.02fF
C18839 PAND2X1_252/O PAND2X1_55/Y 0.05fF
C18840 POR2X1_334/B PAND2X1_767/O 0.02fF
C18841 PAND2X1_48/B POR2X1_573/A 0.03fF
C18842 POR2X1_447/O POR2X1_294/B 0.01fF
C18843 POR2X1_102/Y POR2X1_7/Y 0.01fF
C18844 PAND2X1_803/A PAND2X1_727/O 0.00fF
C18845 PAND2X1_823/a_76_28# PAND2X1_41/B 0.02fF
C18846 POR2X1_685/A POR2X1_676/Y 0.01fF
C18847 PAND2X1_127/CTRL2 POR2X1_78/B 0.13fF
C18848 POR2X1_468/B POR2X1_319/Y 0.47fF
C18849 POR2X1_46/Y POR2X1_7/A 0.08fF
C18850 PAND2X1_61/Y POR2X1_153/Y 0.05fF
C18851 POR2X1_730/Y POR2X1_155/CTRL2 0.03fF
C18852 PAND2X1_857/A POR2X1_821/a_76_344# 0.01fF
C18853 POR2X1_55/Y PAND2X1_344/O 0.17fF
C18854 POR2X1_222/Y POR2X1_194/O 0.09fF
C18855 POR2X1_66/A D_INPUT_4 0.01fF
C18856 POR2X1_396/Y POR2X1_669/a_16_28# 0.03fF
C18857 POR2X1_502/A PAND2X1_373/O 0.04fF
C18858 PAND2X1_39/B POR2X1_579/O 0.07fF
C18859 POR2X1_463/Y VDD 0.11fF
C18860 POR2X1_365/Y POR2X1_212/CTRL 0.03fF
C18861 POR2X1_23/Y PAND2X1_327/CTRL 0.01fF
C18862 POR2X1_62/Y PAND2X1_41/B 1.18fF
C18863 POR2X1_465/B POR2X1_569/A 0.07fF
C18864 POR2X1_83/B POR2X1_373/a_16_28# 0.03fF
C18865 PAND2X1_550/CTRL POR2X1_394/A 0.01fF
C18866 PAND2X1_624/A POR2X1_283/A 0.07fF
C18867 POR2X1_110/Y POR2X1_110/a_16_28# 0.02fF
C18868 POR2X1_756/Y VDD 0.13fF
C18869 PAND2X1_88/Y POR2X1_562/B 0.04fF
C18870 POR2X1_220/Y POR2X1_456/B 0.06fF
C18871 PAND2X1_4/CTRL PAND2X1_6/A 0.01fF
C18872 POR2X1_678/Y POR2X1_728/A 0.00fF
C18873 POR2X1_65/A PAND2X1_800/a_76_28# 0.02fF
C18874 POR2X1_614/A POR2X1_809/Y 0.01fF
C18875 POR2X1_481/Y PAND2X1_854/A 0.02fF
C18876 PAND2X1_209/O POR2X1_394/A 0.02fF
C18877 POR2X1_63/CTRL2 PAND2X1_63/B 0.01fF
C18878 POR2X1_65/A PAND2X1_341/B 0.03fF
C18879 POR2X1_316/CTRL INPUT_0 0.03fF
C18880 POR2X1_569/A POR2X1_501/CTRL 0.02fF
C18881 POR2X1_416/B PAND2X1_34/O 0.09fF
C18882 POR2X1_68/A POR2X1_7/A 0.03fF
C18883 PAND2X1_73/Y PAND2X1_56/A 0.02fF
C18884 POR2X1_356/A POR2X1_338/m4_208_n4# 0.06fF
C18885 POR2X1_404/Y POR2X1_456/B 0.03fF
C18886 POR2X1_43/B POR2X1_283/A 0.88fF
C18887 POR2X1_76/B POR2X1_76/A 0.22fF
C18888 POR2X1_13/A PAND2X1_301/a_76_28# 0.02fF
C18889 POR2X1_379/Y PAND2X1_380/O 0.00fF
C18890 D_INPUT_1 POR2X1_750/O 0.02fF
C18891 POR2X1_174/B PAND2X1_109/a_16_344# 0.07fF
C18892 POR2X1_537/Y POR2X1_733/O 0.01fF
C18893 POR2X1_16/A POR2X1_683/a_16_28# 0.09fF
C18894 POR2X1_75/CTRL2 PAND2X1_349/A 0.01fF
C18895 PAND2X1_359/O PAND2X1_348/Y 0.06fF
C18896 PAND2X1_57/B POR2X1_398/CTRL 0.01fF
C18897 POR2X1_296/B PAND2X1_52/B 0.09fF
C18898 PAND2X1_560/a_16_344# POR2X1_73/Y 0.02fF
C18899 PAND2X1_730/A VDD 0.00fF
C18900 POR2X1_73/O PAND2X1_6/A 0.05fF
C18901 PAND2X1_565/a_16_344# PAND2X1_550/Y 0.03fF
C18902 POR2X1_729/a_16_28# POR2X1_855/B 0.03fF
C18903 POR2X1_245/CTRL2 POR2X1_245/Y 0.06fF
C18904 POR2X1_537/O PAND2X1_55/Y -0.02fF
C18905 POR2X1_855/B PAND2X1_69/A 0.03fF
C18906 PAND2X1_94/A POR2X1_391/Y 0.10fF
C18907 POR2X1_68/A POR2X1_703/A 0.07fF
C18908 PAND2X1_48/B POR2X1_344/Y 0.03fF
C18909 PAND2X1_314/CTRL2 POR2X1_854/B 0.16fF
C18910 PAND2X1_850/Y PAND2X1_787/Y 0.27fF
C18911 POR2X1_183/Y PAND2X1_114/O 0.00fF
C18912 POR2X1_197/O POR2X1_99/B 0.00fF
C18913 PAND2X1_177/O POR2X1_854/B 0.02fF
C18914 PAND2X1_862/B POR2X1_171/Y 0.44fF
C18915 PAND2X1_55/Y POR2X1_186/B 11.65fF
C18916 POR2X1_582/a_16_28# POR2X1_582/A 0.03fF
C18917 POR2X1_557/B POR2X1_294/B 0.29fF
C18918 PAND2X1_190/a_76_28# POR2X1_131/A 0.05fF
C18919 POR2X1_614/A POR2X1_675/Y 0.03fF
C18920 PAND2X1_117/CTRL PAND2X1_48/A 0.01fF
C18921 POR2X1_722/O POR2X1_513/B 0.02fF
C18922 INPUT_3 PAND2X1_206/B 0.10fF
C18923 POR2X1_550/A POR2X1_550/a_16_28# -0.00fF
C18924 PAND2X1_350/O POR2X1_7/A 0.04fF
C18925 POR2X1_599/A POR2X1_394/A 0.22fF
C18926 POR2X1_119/Y PAND2X1_659/a_56_28# 0.00fF
C18927 PAND2X1_48/B POR2X1_349/CTRL2 0.01fF
C18928 POR2X1_5/Y PAND2X1_198/CTRL 0.01fF
C18929 POR2X1_52/A POR2X1_150/O 0.18fF
C18930 POR2X1_203/Y POR2X1_260/A 0.02fF
C18931 POR2X1_339/O POR2X1_556/Y 0.16fF
C18932 POR2X1_416/B POR2X1_743/CTRL2 0.03fF
C18933 POR2X1_83/Y POR2X1_81/Y 0.01fF
C18934 PAND2X1_107/O POR2X1_532/A 0.18fF
C18935 PAND2X1_640/CTRL POR2X1_153/Y 0.06fF
C18936 PAND2X1_229/CTRL2 PAND2X1_72/A 0.00fF
C18937 PAND2X1_563/A POR2X1_90/Y 0.10fF
C18938 POR2X1_760/Y PAND2X1_863/B 0.02fF
C18939 POR2X1_566/A POR2X1_181/CTRL 0.15fF
C18940 POR2X1_707/a_56_344# POR2X1_407/Y -0.00fF
C18941 POR2X1_681/CTRL2 POR2X1_681/Y 0.01fF
C18942 POR2X1_112/a_16_28# POR2X1_332/B 0.08fF
C18943 PAND2X1_96/B POR2X1_244/Y 0.03fF
C18944 PAND2X1_221/Y PAND2X1_798/CTRL2 0.00fF
C18945 POR2X1_508/A POR2X1_508/CTRL 0.01fF
C18946 PAND2X1_352/CTRL POR2X1_55/Y 0.01fF
C18947 PAND2X1_673/O POR2X1_416/B 0.03fF
C18948 POR2X1_740/Y POR2X1_195/m4_208_n4# 0.06fF
C18949 POR2X1_312/Y POR2X1_167/Y 0.00fF
C18950 PAND2X1_476/A PAND2X1_197/Y 0.03fF
C18951 VDD POR2X1_736/A 2.27fF
C18952 POR2X1_293/Y PAND2X1_860/CTRL 0.02fF
C18953 PAND2X1_800/O POR2X1_761/Y 0.00fF
C18954 PAND2X1_6/Y POR2X1_342/CTRL 0.01fF
C18955 POR2X1_416/B POR2X1_13/CTRL 0.01fF
C18956 POR2X1_318/CTRL POR2X1_445/A 0.01fF
C18957 PAND2X1_271/O POR2X1_116/A 0.00fF
C18958 POR2X1_65/A POR2X1_166/Y 0.15fF
C18959 POR2X1_218/CTRL2 POR2X1_260/A 0.01fF
C18960 PAND2X1_650/a_16_344# PAND2X1_641/Y 0.02fF
C18961 POR2X1_180/B POR2X1_703/A 0.03fF
C18962 POR2X1_266/A POR2X1_68/B 0.03fF
C18963 POR2X1_547/B PAND2X1_52/B 0.05fF
C18964 POR2X1_456/B POR2X1_737/CTRL2 0.00fF
C18965 POR2X1_20/Y POR2X1_4/Y 0.01fF
C18966 POR2X1_477/A POR2X1_568/B 0.05fF
C18967 POR2X1_821/m4_208_n4# PAND2X1_659/Y 0.15fF
C18968 PAND2X1_23/Y POR2X1_343/O 0.03fF
C18969 POR2X1_388/O POR2X1_540/Y 0.03fF
C18970 INPUT_6 PAND2X1_18/B 0.20fF
C18971 POR2X1_520/B POR2X1_520/A 0.20fF
C18972 POR2X1_326/A POR2X1_319/Y 0.09fF
C18973 PAND2X1_795/B PAND2X1_332/Y 0.07fF
C18974 POR2X1_188/A POR2X1_643/O 0.01fF
C18975 PAND2X1_699/CTRL2 POR2X1_496/Y 0.05fF
C18976 PAND2X1_163/O POR2X1_210/A 0.01fF
C18977 PAND2X1_254/O POR2X1_77/Y 0.05fF
C18978 POR2X1_591/CTRL POR2X1_77/Y 0.01fF
C18979 POR2X1_157/O POR2X1_416/B 0.18fF
C18980 POR2X1_332/B PAND2X1_135/CTRL 0.01fF
C18981 PAND2X1_63/B PAND2X1_48/A 0.03fF
C18982 PAND2X1_372/O POR2X1_717/B 0.00fF
C18983 POR2X1_654/B POR2X1_643/a_76_344# 0.01fF
C18984 POR2X1_324/Y POR2X1_319/Y 0.04fF
C18985 POR2X1_416/B PAND2X1_798/B 0.07fF
C18986 POR2X1_630/B POR2X1_630/A 0.31fF
C18987 POR2X1_67/Y POR2X1_69/A 0.00fF
C18988 POR2X1_846/Y POR2X1_753/a_76_344# 0.00fF
C18989 PAND2X1_222/B PAND2X1_643/A 0.09fF
C18990 POR2X1_301/A POR2X1_76/A 0.02fF
C18991 POR2X1_156/O POR2X1_162/Y 0.01fF
C18992 POR2X1_77/CTRL2 POR2X1_48/A 0.03fF
C18993 POR2X1_296/Y POR2X1_296/CTRL 0.02fF
C18994 POR2X1_610/O POR2X1_862/A 0.01fF
C18995 POR2X1_394/A POR2X1_599/O 0.01fF
C18996 POR2X1_508/B PAND2X1_823/CTRL 0.00fF
C18997 PAND2X1_641/O PAND2X1_341/B 0.19fF
C18998 POR2X1_471/A POR2X1_454/B 0.03fF
C18999 POR2X1_600/Y POR2X1_601/O 0.01fF
C19000 PAND2X1_469/B POR2X1_173/a_16_28# 0.03fF
C19001 POR2X1_60/A POR2X1_253/CTRL 0.01fF
C19002 POR2X1_257/A POR2X1_102/Y 0.13fF
C19003 PAND2X1_312/O POR2X1_736/A 0.32fF
C19004 POR2X1_349/CTRL POR2X1_363/A 0.01fF
C19005 POR2X1_567/CTRL POR2X1_854/B 0.15fF
C19006 PAND2X1_349/A PAND2X1_840/Y 0.04fF
C19007 PAND2X1_240/CTRL2 POR2X1_411/B 0.01fF
C19008 POR2X1_501/B POR2X1_138/A 0.03fF
C19009 D_INPUT_5 POR2X1_634/A 0.03fF
C19010 PAND2X1_175/B PAND2X1_861/B 0.02fF
C19011 POR2X1_14/Y PAND2X1_35/A 0.01fF
C19012 POR2X1_303/B POR2X1_723/B 0.50fF
C19013 INPUT_3 POR2X1_750/B 0.07fF
C19014 POR2X1_703/A POR2X1_169/A 0.01fF
C19015 POR2X1_48/A PAND2X1_400/O 0.01fF
C19016 POR2X1_257/A PAND2X1_436/A 0.20fF
C19017 PAND2X1_294/a_56_28# POR2X1_60/A 0.00fF
C19018 POR2X1_527/CTRL POR2X1_39/B 0.01fF
C19019 PAND2X1_644/Y POR2X1_669/B 0.17fF
C19020 POR2X1_54/Y POR2X1_40/Y 0.06fF
C19021 POR2X1_579/a_16_28# POR2X1_576/Y 0.03fF
C19022 POR2X1_866/A PAND2X1_58/A 0.03fF
C19023 PAND2X1_659/A PAND2X1_203/O 0.03fF
C19024 POR2X1_88/CTRL POR2X1_69/A 0.01fF
C19025 PAND2X1_33/O POR2X1_5/Y 0.16fF
C19026 PAND2X1_73/Y POR2X1_266/a_16_28# 0.00fF
C19027 POR2X1_54/Y POR2X1_35/B 0.05fF
C19028 POR2X1_815/O VDD 0.00fF
C19029 POR2X1_602/B PAND2X1_601/CTRL 0.01fF
C19030 POR2X1_741/O POR2X1_186/B 0.02fF
C19031 D_INPUT_0 POR2X1_413/CTRL2 0.00fF
C19032 INPUT_1 PAND2X1_462/O 0.01fF
C19033 POR2X1_49/Y PAND2X1_340/B 3.53fF
C19034 D_INPUT_5 PAND2X1_588/CTRL2 0.00fF
C19035 PAND2X1_156/A PAND2X1_508/B 0.05fF
C19036 POR2X1_760/A POR2X1_46/Y 0.01fF
C19037 POR2X1_57/A PAND2X1_860/A 0.09fF
C19038 D_INPUT_7 PAND2X1_587/CTRL 0.01fF
C19039 PAND2X1_93/B POR2X1_750/B 0.05fF
C19040 PAND2X1_58/A PAND2X1_381/Y 0.02fF
C19041 POR2X1_502/A POR2X1_444/CTRL 0.01fF
C19042 POR2X1_482/O POR2X1_482/Y 0.01fF
C19043 POR2X1_661/A PAND2X1_306/CTRL 0.06fF
C19044 PAND2X1_576/B PAND2X1_576/CTRL2 0.01fF
C19045 PAND2X1_687/a_16_344# POR2X1_761/A 0.01fF
C19046 POR2X1_856/B POR2X1_355/A 0.02fF
C19047 POR2X1_376/B POR2X1_817/CTRL2 0.01fF
C19048 PAND2X1_61/a_56_28# POR2X1_60/A 0.00fF
C19049 POR2X1_777/B D_INPUT_0 0.05fF
C19050 POR2X1_78/B POR2X1_222/O 0.06fF
C19051 POR2X1_467/Y POR2X1_296/B 0.07fF
C19052 POR2X1_60/A POR2X1_516/Y 0.01fF
C19053 PAND2X1_746/O PAND2X1_52/B 0.05fF
C19054 POR2X1_660/A D_INPUT_0 3.71fF
C19055 INPUT_3 POR2X1_618/CTRL 0.06fF
C19056 POR2X1_150/Y PAND2X1_390/CTRL 0.00fF
C19057 POR2X1_555/A POR2X1_66/A 0.03fF
C19058 POR2X1_856/CTRL2 PAND2X1_73/Y 0.01fF
C19059 POR2X1_13/A POR2X1_672/Y 0.00fF
C19060 POR2X1_78/A POR2X1_750/B 0.10fF
C19061 POR2X1_16/A POR2X1_16/CTRL2 0.01fF
C19062 POR2X1_596/A POR2X1_814/A 0.05fF
C19063 POR2X1_628/Y POR2X1_293/Y 0.03fF
C19064 PAND2X1_65/B D_INPUT_0 16.51fF
C19065 PAND2X1_472/B PAND2X1_35/A 0.02fF
C19066 POR2X1_424/Y POR2X1_424/m4_208_n4# 0.02fF
C19067 PAND2X1_223/B PAND2X1_223/O 0.01fF
C19068 PAND2X1_611/CTRL POR2X1_68/B 0.01fF
C19069 POR2X1_270/Y VDD 0.19fF
C19070 POR2X1_609/Y PAND2X1_403/Y 0.00fF
C19071 POR2X1_49/Y POR2X1_102/Y 0.17fF
C19072 POR2X1_83/A POR2X1_20/B 0.02fF
C19073 PAND2X1_23/Y PAND2X1_39/B 0.05fF
C19074 POR2X1_13/A PAND2X1_124/Y 0.03fF
C19075 POR2X1_66/B PAND2X1_88/O 0.02fF
C19076 POR2X1_418/Y POR2X1_417/Y 0.00fF
C19077 POR2X1_334/B POR2X1_473/CTRL2 0.13fF
C19078 POR2X1_263/Y VDD 0.55fF
C19079 POR2X1_66/B POR2X1_476/O 0.07fF
C19080 POR2X1_806/a_16_28# POR2X1_330/Y 0.04fF
C19081 PAND2X1_85/Y PAND2X1_15/CTRL 0.06fF
C19082 POR2X1_102/Y PAND2X1_558/CTRL2 0.01fF
C19083 PAND2X1_612/B POR2X1_642/CTRL2 0.00fF
C19084 PAND2X1_90/A PAND2X1_613/CTRL 0.09fF
C19085 POR2X1_669/B PAND2X1_550/CTRL 0.04fF
C19086 PAND2X1_35/A POR2X1_55/Y 0.02fF
C19087 POR2X1_96/A PAND2X1_571/A 0.02fF
C19088 PAND2X1_625/O PAND2X1_39/B 0.03fF
C19089 POR2X1_774/Y POR2X1_812/A 0.03fF
C19090 POR2X1_20/B POR2X1_90/Y 0.22fF
C19091 POR2X1_695/Y PAND2X1_707/O 0.00fF
C19092 POR2X1_347/B POR2X1_68/CTRL2 0.10fF
C19093 POR2X1_567/B POR2X1_776/B 0.62fF
C19094 POR2X1_65/A POR2X1_295/O 0.02fF
C19095 POR2X1_669/B PAND2X1_556/B 0.19fF
C19096 PAND2X1_810/A PAND2X1_805/A 0.03fF
C19097 POR2X1_817/Y PAND2X1_340/B 0.01fF
C19098 PAND2X1_289/CTRL2 POR2X1_210/Y 0.01fF
C19099 POR2X1_260/B POR2X1_459/A 0.03fF
C19100 POR2X1_52/A POR2X1_626/O 0.01fF
C19101 POR2X1_355/O POR2X1_355/A 0.02fF
C19102 POR2X1_120/a_56_344# POR2X1_78/A 0.00fF
C19103 POR2X1_241/B POR2X1_483/B 0.02fF
C19104 POR2X1_437/O PAND2X1_794/B 0.01fF
C19105 PAND2X1_418/a_16_344# POR2X1_854/B 0.06fF
C19106 POR2X1_590/A PAND2X1_372/CTRL -0.00fF
C19107 PAND2X1_76/Y PAND2X1_390/Y 0.03fF
C19108 PAND2X1_254/Y POR2X1_669/B 0.07fF
C19109 POR2X1_631/m4_208_n4# POR2X1_193/Y 0.08fF
C19110 POR2X1_478/m4_208_n4# POR2X1_468/m4_208_n4# 0.13fF
C19111 POR2X1_270/Y POR2X1_741/Y 0.06fF
C19112 POR2X1_13/A POR2X1_83/B 0.54fF
C19113 POR2X1_376/B POR2X1_427/Y 0.19fF
C19114 PAND2X1_93/B PAND2X1_72/CTRL2 0.01fF
C19115 POR2X1_811/A PAND2X1_599/O 0.00fF
C19116 D_INPUT_2 D_INPUT_0 0.00fF
C19117 PAND2X1_58/A PAND2X1_754/CTRL 0.01fF
C19118 PAND2X1_859/A PAND2X1_859/a_76_28# 0.04fF
C19119 POR2X1_477/B VDD 0.00fF
C19120 POR2X1_66/B POR2X1_404/B 0.00fF
C19121 PAND2X1_261/CTRL POR2X1_330/Y 0.10fF
C19122 POR2X1_83/B PAND2X1_214/B 0.01fF
C19123 PAND2X1_674/O POR2X1_466/A 0.31fF
C19124 POR2X1_333/A POR2X1_468/B 0.18fF
C19125 POR2X1_102/Y PAND2X1_553/B 0.07fF
C19126 POR2X1_628/Y POR2X1_408/Y 0.05fF
C19127 POR2X1_60/O PAND2X1_404/Y 0.01fF
C19128 POR2X1_416/Y POR2X1_37/Y 0.08fF
C19129 POR2X1_857/a_16_28# POR2X1_192/Y 0.10fF
C19130 PAND2X1_661/B PAND2X1_124/Y 0.03fF
C19131 POR2X1_63/CTRL2 POR2X1_32/A 0.01fF
C19132 PAND2X1_65/B PAND2X1_90/Y 1.21fF
C19133 PAND2X1_96/B POR2X1_195/A 0.03fF
C19134 PAND2X1_23/Y POR2X1_805/Y 0.03fF
C19135 POR2X1_857/CTRL2 POR2X1_795/B 0.01fF
C19136 POR2X1_556/A POR2X1_773/B 0.05fF
C19137 PAND2X1_423/CTRL2 PAND2X1_57/B 0.01fF
C19138 POR2X1_329/A PAND2X1_156/A 0.10fF
C19139 POR2X1_102/Y PAND2X1_188/O 0.11fF
C19140 POR2X1_135/Y PAND2X1_332/O 0.03fF
C19141 PAND2X1_23/Y PAND2X1_20/A 0.47fF
C19142 POR2X1_23/Y PAND2X1_457/m4_208_n4# 0.06fF
C19143 PAND2X1_48/B POR2X1_719/A 0.00fF
C19144 PAND2X1_392/a_16_344# POR2X1_816/A 0.01fF
C19145 POR2X1_200/CTRL2 POR2X1_294/B 0.07fF
C19146 POR2X1_52/A PAND2X1_465/O 0.01fF
C19147 POR2X1_75/CTRL2 POR2X1_32/A 0.03fF
C19148 PAND2X1_604/CTRL2 POR2X1_750/B 0.07fF
C19149 POR2X1_63/O POR2X1_83/B 0.16fF
C19150 POR2X1_43/B POR2X1_14/Y 0.30fF
C19151 POR2X1_832/B POR2X1_330/Y 0.05fF
C19152 POR2X1_65/A POR2X1_683/O 0.02fF
C19153 POR2X1_476/m4_208_n4# POR2X1_121/Y 0.09fF
C19154 PAND2X1_65/B PAND2X1_760/O 0.03fF
C19155 POR2X1_441/Y POR2X1_394/A 0.17fF
C19156 PAND2X1_23/Y PAND2X1_96/CTRL 0.00fF
C19157 POR2X1_94/A POR2X1_42/Y 0.06fF
C19158 POR2X1_288/O PAND2X1_32/B 0.01fF
C19159 POR2X1_78/B POR2X1_194/B 0.01fF
C19160 PAND2X1_16/CTRL POR2X1_785/A 0.00fF
C19161 POR2X1_260/B POR2X1_375/CTRL2 0.03fF
C19162 PAND2X1_229/O POR2X1_231/B 0.02fF
C19163 PAND2X1_798/B POR2X1_487/Y 0.07fF
C19164 PAND2X1_23/Y PAND2X1_250/O 0.07fF
C19165 POR2X1_65/A POR2X1_517/Y 0.01fF
C19166 POR2X1_49/Y POR2X1_528/CTRL2 0.03fF
C19167 POR2X1_688/Y POR2X1_260/A 0.01fF
C19168 PAND2X1_474/Y PAND2X1_795/B 0.17fF
C19169 INPUT_0 PAND2X1_8/Y 0.16fF
C19170 POR2X1_13/A PAND2X1_140/Y 1.77fF
C19171 POR2X1_16/A POR2X1_88/CTRL 0.00fF
C19172 PAND2X1_220/CTRL2 PAND2X1_220/Y 0.00fF
C19173 PAND2X1_661/B POR2X1_83/B 0.03fF
C19174 POR2X1_693/Y POR2X1_72/B 0.11fF
C19175 PAND2X1_223/a_76_28# POR2X1_7/B 0.01fF
C19176 PAND2X1_23/Y POR2X1_814/B 0.20fF
C19177 POR2X1_657/CTRL2 POR2X1_724/A 0.03fF
C19178 PAND2X1_48/B POR2X1_105/Y 6.99fF
C19179 POR2X1_686/CTRL PAND2X1_73/Y 0.01fF
C19180 POR2X1_240/B PAND2X1_88/Y 0.00fF
C19181 POR2X1_827/CTRL2 POR2X1_39/B -0.00fF
C19182 PAND2X1_826/CTRL POR2X1_507/A 0.04fF
C19183 POR2X1_174/B POR2X1_532/A 0.03fF
C19184 POR2X1_14/Y POR2X1_38/B 0.58fF
C19185 POR2X1_78/A PAND2X1_424/O 0.03fF
C19186 POR2X1_150/Y PAND2X1_716/B 0.03fF
C19187 POR2X1_72/a_16_28# POR2X1_71/Y 0.06fF
C19188 POR2X1_13/A PAND2X1_795/B 0.00fF
C19189 POR2X1_813/Y POR2X1_263/Y 0.01fF
C19190 PAND2X1_675/A PAND2X1_220/Y 0.10fF
C19191 POR2X1_110/Y POR2X1_20/B 0.09fF
C19192 POR2X1_468/O VDD 0.00fF
C19193 PAND2X1_6/Y POR2X1_186/Y 0.10fF
C19194 POR2X1_809/A PAND2X1_39/B 0.02fF
C19195 PAND2X1_46/O D_INPUT_1 0.08fF
C19196 PAND2X1_198/Y PAND2X1_35/Y 0.04fF
C19197 PAND2X1_215/B VDD 0.02fF
C19198 POR2X1_649/a_16_28# POR2X1_294/A 0.07fF
C19199 PAND2X1_23/Y POR2X1_325/A 2.59fF
C19200 POR2X1_60/A POR2X1_534/O 0.01fF
C19201 POR2X1_614/Y PAND2X1_63/B 0.18fF
C19202 D_INPUT_1 POR2X1_389/Y 0.02fF
C19203 POR2X1_866/A POR2X1_596/a_76_344# 0.03fF
C19204 POR2X1_407/A POR2X1_475/A 0.03fF
C19205 PAND2X1_6/A PAND2X1_392/B 0.10fF
C19206 POR2X1_811/CTRL POR2X1_260/A 0.01fF
C19207 PAND2X1_644/a_16_344# POR2X1_761/A 0.02fF
C19208 POR2X1_860/CTRL POR2X1_218/Y 0.04fF
C19209 POR2X1_720/A POR2X1_816/A 0.04fF
C19210 POR2X1_653/O POR2X1_740/Y 0.00fF
C19211 POR2X1_315/O PAND2X1_803/A 0.00fF
C19212 POR2X1_32/A PAND2X1_550/B 0.34fF
C19213 PAND2X1_57/B POR2X1_404/Y 0.03fF
C19214 PAND2X1_58/A POR2X1_7/A 0.03fF
C19215 POR2X1_60/A PAND2X1_843/Y 0.03fF
C19216 POR2X1_73/a_76_344# POR2X1_37/Y 0.00fF
C19217 POR2X1_329/A PAND2X1_339/O 0.03fF
C19218 POR2X1_68/B POR2X1_734/A 0.09fF
C19219 PAND2X1_378/O PAND2X1_377/Y 0.00fF
C19220 PAND2X1_787/A POR2X1_40/Y 0.03fF
C19221 POR2X1_590/A PAND2X1_528/O 0.05fF
C19222 POR2X1_355/B POR2X1_579/Y 0.20fF
C19223 PAND2X1_94/A POR2X1_650/CTRL2 0.34fF
C19224 POR2X1_433/Y PAND2X1_499/Y 0.02fF
C19225 POR2X1_516/A POR2X1_516/Y 0.01fF
C19226 PAND2X1_731/a_76_28# PAND2X1_738/B 0.03fF
C19227 POR2X1_449/a_16_28# POR2X1_832/B -0.00fF
C19228 POR2X1_23/Y PAND2X1_853/B 0.09fF
C19229 POR2X1_333/O POR2X1_174/B 0.00fF
C19230 POR2X1_68/A POR2X1_206/A 0.01fF
C19231 PAND2X1_840/A PAND2X1_499/a_76_28# 0.05fF
C19232 PAND2X1_654/CTRL POR2X1_46/Y 0.01fF
C19233 POR2X1_293/Y POR2X1_372/Y 0.02fF
C19234 PAND2X1_798/B PAND2X1_738/Y 0.10fF
C19235 POR2X1_612/Y POR2X1_5/CTRL 0.04fF
C19236 POR2X1_43/B PAND2X1_735/O 0.06fF
C19237 POR2X1_252/CTRL POR2X1_55/Y 0.01fF
C19238 POR2X1_555/A POR2X1_532/A 0.00fF
C19239 PAND2X1_6/A VDD 5.62fF
C19240 POR2X1_567/B POR2X1_180/CTRL 0.01fF
C19241 POR2X1_184/Y PAND2X1_139/Y 0.00fF
C19242 POR2X1_401/CTRL2 PAND2X1_69/A 0.03fF
C19243 POR2X1_286/CTRL POR2X1_774/A 0.00fF
C19244 PAND2X1_93/O PAND2X1_57/B 0.01fF
C19245 POR2X1_307/a_56_344# POR2X1_796/A 0.00fF
C19246 POR2X1_355/B POR2X1_545/A 0.03fF
C19247 POR2X1_391/A POR2X1_391/CTRL2 0.00fF
C19248 PAND2X1_389/CTRL VDD 0.00fF
C19249 POR2X1_851/CTRL2 POR2X1_590/A 0.03fF
C19250 PAND2X1_65/B POR2X1_789/O 0.07fF
C19251 PAND2X1_516/CTRL2 POR2X1_513/Y 0.03fF
C19252 POR2X1_13/A POR2X1_494/O 0.16fF
C19253 PAND2X1_216/B PAND2X1_561/Y 0.71fF
C19254 POR2X1_270/CTRL2 POR2X1_78/B 0.16fF
C19255 PAND2X1_653/Y INPUT_0 0.02fF
C19256 PAND2X1_651/Y PAND2X1_455/Y 0.00fF
C19257 PAND2X1_652/A PAND2X1_592/Y 0.07fF
C19258 POR2X1_538/CTRL POR2X1_193/A 0.03fF
C19259 POR2X1_740/Y POR2X1_294/B 0.09fF
C19260 POR2X1_366/Y POR2X1_740/Y 0.03fF
C19261 PAND2X1_688/O POR2X1_38/Y 0.04fF
C19262 D_INPUT_3 POR2X1_58/CTRL 0.28fF
C19263 PAND2X1_90/Y POR2X1_712/O 0.10fF
C19264 PAND2X1_766/O POR2X1_707/Y 0.17fF
C19265 PAND2X1_335/CTRL POR2X1_309/Y 0.07fF
C19266 POR2X1_43/B PAND2X1_341/CTRL2 0.01fF
C19267 PAND2X1_124/Y PAND2X1_199/O 0.03fF
C19268 POR2X1_416/Y POR2X1_293/Y 1.68fF
C19269 POR2X1_441/Y PAND2X1_326/CTRL 0.01fF
C19270 POR2X1_763/Y PAND2X1_546/CTRL 0.08fF
C19271 PAND2X1_787/Y POR2X1_7/A 0.05fF
C19272 PAND2X1_243/CTRL2 PAND2X1_35/Y 0.01fF
C19273 POR2X1_43/B POR2X1_55/Y 0.11fF
C19274 POR2X1_124/CTRL2 POR2X1_556/A 0.01fF
C19275 POR2X1_480/A POR2X1_319/Y 0.07fF
C19276 POR2X1_253/Y POR2X1_293/Y 0.02fF
C19277 PAND2X1_39/B POR2X1_711/Y 0.07fF
C19278 POR2X1_334/B POR2X1_124/m4_208_n4# 0.06fF
C19279 PAND2X1_700/a_56_28# POR2X1_532/A 0.00fF
C19280 POR2X1_296/B POR2X1_722/CTRL2 0.03fF
C19281 PAND2X1_665/CTRL PAND2X1_93/B 0.02fF
C19282 PAND2X1_472/B POR2X1_38/B 0.07fF
C19283 POR2X1_257/A POR2X1_320/Y 0.01fF
C19284 PAND2X1_848/B POR2X1_382/CTRL2 0.01fF
C19285 PAND2X1_491/CTRL2 POR2X1_294/B 0.10fF
C19286 PAND2X1_631/A POR2X1_482/CTRL 0.01fF
C19287 GATE_741 PAND2X1_568/B 0.03fF
C19288 POR2X1_38/Y POR2X1_46/Y 0.09fF
C19289 VDD POR2X1_351/CTRL2 0.00fF
C19290 PAND2X1_206/O POR2X1_7/A 0.02fF
C19291 POR2X1_669/B POR2X1_320/O 0.01fF
C19292 POR2X1_316/CTRL PAND2X1_436/A 0.03fF
C19293 INPUT_1 POR2X1_710/A 0.01fF
C19294 D_GATE_222 POR2X1_775/CTRL2 0.03fF
C19295 POR2X1_66/B PAND2X1_481/a_16_344# 0.01fF
C19296 POR2X1_76/Y POR2X1_203/O 0.03fF
C19297 PAND2X1_755/a_16_344# PAND2X1_60/B 0.02fF
C19298 POR2X1_685/CTRL POR2X1_687/A 0.01fF
C19299 POR2X1_76/Y PAND2X1_111/B 0.02fF
C19300 POR2X1_588/Y VDD 0.25fF
C19301 PAND2X1_653/Y PAND2X1_218/CTRL 0.02fF
C19302 PAND2X1_830/Y PAND2X1_389/Y 0.12fF
C19303 POR2X1_542/B PAND2X1_55/Y 0.04fF
C19304 POR2X1_38/B POR2X1_55/Y 0.00fF
C19305 POR2X1_332/B POR2X1_366/A 0.10fF
C19306 POR2X1_804/A POR2X1_130/Y 0.26fF
C19307 POR2X1_116/CTRL POR2X1_260/A 0.00fF
C19308 PAND2X1_623/Y POR2X1_38/Y 0.03fF
C19309 POR2X1_75/CTRL2 POR2X1_184/Y 0.00fF
C19310 POR2X1_124/a_16_28# POR2X1_123/Y 0.04fF
C19311 PAND2X1_55/Y PAND2X1_79/Y 0.14fF
C19312 POR2X1_101/Y VDD 3.90fF
C19313 POR2X1_280/Y VDD 0.20fF
C19314 PAND2X1_716/CTRL POR2X1_52/Y 0.01fF
C19315 POR2X1_335/A PAND2X1_311/CTRL2 0.01fF
C19316 POR2X1_583/CTRL POR2X1_42/Y 0.04fF
C19317 POR2X1_333/A POR2X1_324/Y 0.33fF
C19318 PAND2X1_864/CTRL2 GATE_741 0.01fF
C19319 POR2X1_102/Y PAND2X1_865/A 0.06fF
C19320 VDD PAND2X1_112/O 0.00fF
C19321 POR2X1_719/CTRL PAND2X1_48/B 0.00fF
C19322 POR2X1_13/A PAND2X1_196/CTRL 0.01fF
C19323 PAND2X1_55/Y POR2X1_736/O 0.10fF
C19324 POR2X1_20/Y D_INPUT_1 -0.01fF
C19325 POR2X1_355/B POR2X1_440/Y 0.03fF
C19326 POR2X1_71/CTRL POR2X1_5/Y 0.01fF
C19327 POR2X1_65/A POR2X1_177/O 0.01fF
C19328 POR2X1_65/CTRL POR2X1_9/Y 0.08fF
C19329 POR2X1_740/Y PAND2X1_111/B 0.05fF
C19330 PAND2X1_798/B PAND2X1_575/O 0.03fF
C19331 PAND2X1_678/O PAND2X1_860/A 0.04fF
C19332 POR2X1_68/A POR2X1_140/O 0.02fF
C19333 PAND2X1_797/Y POR2X1_60/A 0.05fF
C19334 POR2X1_557/A PAND2X1_57/B 0.01fF
C19335 PAND2X1_636/O POR2X1_260/A 0.01fF
C19336 PAND2X1_693/CTRL2 POR2X1_383/A 0.01fF
C19337 POR2X1_83/O PAND2X1_35/Y 0.01fF
C19338 POR2X1_119/Y PAND2X1_217/B 0.19fF
C19339 POR2X1_605/A PAND2X1_69/A 0.01fF
C19340 POR2X1_583/Y VDD 0.00fF
C19341 POR2X1_502/A POR2X1_260/A 0.03fF
C19342 PAND2X1_237/CTRL PAND2X1_72/A 0.00fF
C19343 POR2X1_783/A POR2X1_260/A 0.01fF
C19344 PAND2X1_602/Y PAND2X1_648/a_76_28# 0.05fF
C19345 PAND2X1_484/CTRL2 INPUT_0 0.03fF
C19346 POR2X1_383/A POR2X1_264/Y 0.07fF
C19347 POR2X1_32/A PAND2X1_840/Y 4.89fF
C19348 POR2X1_99/B PAND2X1_7/Y 0.66fF
C19349 POR2X1_337/CTRL POR2X1_260/A 0.01fF
C19350 POR2X1_570/B POR2X1_341/Y 0.01fF
C19351 POR2X1_72/CTRL2 POR2X1_72/B 0.00fF
C19352 POR2X1_189/Y PAND2X1_728/CTRL2 0.01fF
C19353 POR2X1_63/a_16_28# POR2X1_38/Y 0.08fF
C19354 POR2X1_114/O POR2X1_113/Y 0.03fF
C19355 POR2X1_516/CTRL2 POR2X1_283/A 0.01fF
C19356 POR2X1_680/CTRL POR2X1_40/Y 0.01fF
C19357 PAND2X1_666/O PAND2X1_72/A 0.03fF
C19358 POR2X1_330/Y POR2X1_330/O 0.06fF
C19359 D_INPUT_1 POR2X1_318/A 0.07fF
C19360 PAND2X1_551/CTRL2 POR2X1_90/Y 0.01fF
C19361 POR2X1_78/B PAND2X1_48/A 0.07fF
C19362 POR2X1_804/A POR2X1_228/Y 0.07fF
C19363 POR2X1_257/A POR2X1_677/Y 3.09fF
C19364 POR2X1_55/Y PAND2X1_336/O 0.05fF
C19365 POR2X1_122/a_16_28# POR2X1_122/A 0.03fF
C19366 INPUT_1 PAND2X1_623/Y 0.01fF
C19367 POR2X1_462/B POR2X1_713/B 0.05fF
C19368 POR2X1_29/Y POR2X1_408/Y 0.00fF
C19369 PAND2X1_20/A POR2X1_711/Y 2.28fF
C19370 POR2X1_46/Y POR2X1_153/Y 0.32fF
C19371 POR2X1_132/O VDD 0.00fF
C19372 POR2X1_41/B PAND2X1_200/B 1.57fF
C19373 PAND2X1_342/O POR2X1_248/Y 0.02fF
C19374 POR2X1_687/A POR2X1_730/O 0.01fF
C19375 POR2X1_502/A PAND2X1_142/O 0.04fF
C19376 POR2X1_592/Y POR2X1_593/B 0.05fF
C19377 POR2X1_494/O PAND2X1_510/B 0.01fF
C19378 POR2X1_722/O VDD 0.00fF
C19379 POR2X1_724/A POR2X1_318/A 0.07fF
C19380 POR2X1_244/B POR2X1_228/O 0.01fF
C19381 POR2X1_49/Y POR2X1_761/A 1.93fF
C19382 POR2X1_814/O POR2X1_260/B 0.01fF
C19383 POR2X1_119/Y VDD 4.56fF
C19384 POR2X1_863/A POR2X1_466/A 0.07fF
C19385 POR2X1_68/A INPUT_1 5.67fF
C19386 POR2X1_523/Y POR2X1_546/CTRL2 0.03fF
C19387 POR2X1_762/O INPUT_4 0.01fF
C19388 POR2X1_633/A PAND2X1_52/B 0.03fF
C19389 POR2X1_101/Y PAND2X1_32/B 0.07fF
C19390 POR2X1_504/Y POR2X1_39/B 0.03fF
C19391 POR2X1_278/Y POR2X1_7/Y 0.05fF
C19392 PAND2X1_661/B PAND2X1_196/CTRL 0.01fF
C19393 POR2X1_673/Y PAND2X1_6/A 0.06fF
C19394 PAND2X1_824/B PAND2X1_93/CTRL 0.01fF
C19395 POR2X1_316/Y POR2X1_5/Y 0.03fF
C19396 POR2X1_447/B POR2X1_835/Y 0.02fF
C19397 POR2X1_774/A POR2X1_294/B 0.03fF
C19398 POR2X1_114/O POR2X1_260/A 0.16fF
C19399 POR2X1_383/A POR2X1_712/CTRL 0.01fF
C19400 POR2X1_8/Y POR2X1_672/A 0.01fF
C19401 PAND2X1_716/B PAND2X1_364/B 0.09fF
C19402 PAND2X1_690/CTRL2 PAND2X1_32/B 0.01fF
C19403 PAND2X1_843/O POR2X1_416/B 0.01fF
C19404 PAND2X1_96/B POR2X1_703/A 0.03fF
C19405 POR2X1_814/B POR2X1_711/Y 0.07fF
C19406 POR2X1_468/Y POR2X1_568/Y 0.36fF
C19407 POR2X1_68/A POR2X1_782/O 0.01fF
C19408 PAND2X1_23/Y POR2X1_332/Y 0.01fF
C19409 PAND2X1_48/B POR2X1_773/A 0.12fF
C19410 POR2X1_574/A POR2X1_366/A 0.01fF
C19411 PAND2X1_721/CTRL POR2X1_77/Y 0.01fF
C19412 POR2X1_174/O PAND2X1_32/B 0.02fF
C19413 POR2X1_727/CTRL2 POR2X1_854/B 0.04fF
C19414 POR2X1_186/Y PAND2X1_52/B 0.26fF
C19415 POR2X1_341/Y POR2X1_351/a_16_28# 0.03fF
C19416 POR2X1_536/CTRL PAND2X1_222/B 0.01fF
C19417 POR2X1_187/a_16_28# POR2X1_594/A 0.03fF
C19418 POR2X1_529/a_16_28# POR2X1_384/A 0.02fF
C19419 POR2X1_383/A POR2X1_351/O 0.03fF
C19420 POR2X1_16/A PAND2X1_568/B 0.03fF
C19421 POR2X1_567/A POR2X1_740/Y 0.03fF
C19422 POR2X1_345/CTRL2 POR2X1_197/Y 0.03fF
C19423 POR2X1_447/CTRL2 POR2X1_186/B 0.04fF
C19424 PAND2X1_439/O POR2X1_438/Y 0.09fF
C19425 POR2X1_190/Y POR2X1_568/B 0.21fF
C19426 POR2X1_13/A PAND2X1_841/Y 0.04fF
C19427 POR2X1_222/A POR2X1_456/B 0.03fF
C19428 POR2X1_326/A POR2X1_788/B 0.01fF
C19429 POR2X1_240/B PAND2X1_234/O 0.00fF
C19430 POR2X1_814/A D_INPUT_0 0.11fF
C19431 PAND2X1_216/B PAND2X1_717/Y 0.12fF
C19432 POR2X1_814/A POR2X1_811/A 0.05fF
C19433 POR2X1_57/A PAND2X1_156/A 0.03fF
C19434 PAND2X1_620/a_16_344# POR2X1_408/Y 0.07fF
C19435 POR2X1_164/Y POR2X1_16/A 0.03fF
C19436 PAND2X1_454/B PAND2X1_796/B 0.02fF
C19437 PAND2X1_323/CTRL2 PAND2X1_32/B 0.01fF
C19438 PAND2X1_6/Y POR2X1_542/Y 0.01fF
C19439 POR2X1_121/CTRL2 POR2X1_537/Y 0.01fF
C19440 POR2X1_814/B PAND2X1_233/CTRL 0.08fF
C19441 PAND2X1_222/O PAND2X1_222/A 0.02fF
C19442 POR2X1_257/A PAND2X1_469/a_16_344# 0.01fF
C19443 POR2X1_68/B PAND2X1_396/O 0.03fF
C19444 INPUT_1 POR2X1_376/O 0.18fF
C19445 POR2X1_329/A PAND2X1_215/CTRL 0.03fF
C19446 POR2X1_416/B PAND2X1_552/B 0.03fF
C19447 POR2X1_385/Y POR2X1_387/Y 0.04fF
C19448 POR2X1_49/Y POR2X1_9/Y 0.34fF
C19449 POR2X1_623/Y POR2X1_296/B 0.03fF
C19450 POR2X1_184/Y PAND2X1_840/Y 0.06fF
C19451 POR2X1_411/B POR2X1_616/a_16_28# 0.03fF
C19452 POR2X1_486/B PAND2X1_69/A 0.32fF
C19453 POR2X1_510/Y POR2X1_540/Y 0.43fF
C19454 POR2X1_441/Y POR2X1_669/B 0.05fF
C19455 POR2X1_193/A PAND2X1_135/CTRL 0.00fF
C19456 PAND2X1_663/O PAND2X1_662/Y 0.00fF
C19457 POR2X1_579/Y PAND2X1_135/CTRL 0.00fF
C19458 POR2X1_135/O POR2X1_7/A 0.01fF
C19459 PAND2X1_651/Y PAND2X1_840/Y 0.03fF
C19460 PAND2X1_480/B POR2X1_310/CTRL2 0.30fF
C19461 POR2X1_286/B PAND2X1_595/O 0.01fF
C19462 PAND2X1_865/Y POR2X1_283/A 0.07fF
C19463 POR2X1_23/CTRL2 POR2X1_20/B 0.01fF
C19464 POR2X1_48/A POR2X1_600/Y 0.01fF
C19465 PAND2X1_242/Y POR2X1_372/Y 0.12fF
C19466 POR2X1_539/A POR2X1_374/O 0.02fF
C19467 POR2X1_344/Y POR2X1_359/B 0.00fF
C19468 PAND2X1_274/O POR2X1_677/Y 0.00fF
C19469 POR2X1_860/CTRL POR2X1_861/A 0.04fF
C19470 POR2X1_514/CTRL POR2X1_138/A 0.00fF
C19471 POR2X1_188/Y POR2X1_260/A 0.00fF
C19472 PAND2X1_6/Y POR2X1_717/B 0.05fF
C19473 POR2X1_438/a_16_28# POR2X1_77/Y 0.03fF
C19474 POR2X1_814/A PAND2X1_90/Y 0.19fF
C19475 PAND2X1_65/B POR2X1_260/O 0.18fF
C19476 POR2X1_242/CTRL2 POR2X1_776/A 0.01fF
C19477 POR2X1_614/A PAND2X1_135/CTRL 0.01fF
C19478 PAND2X1_620/O POR2X1_613/Y -0.00fF
C19479 POR2X1_838/B PAND2X1_67/O 0.00fF
C19480 POR2X1_597/Y POR2X1_40/Y 0.18fF
C19481 POR2X1_431/CTRL POR2X1_236/Y 0.04fF
C19482 POR2X1_593/O POR2X1_802/A 0.05fF
C19483 PAND2X1_60/O PAND2X1_58/A 0.11fF
C19484 POR2X1_41/B POR2X1_846/A 0.19fF
C19485 POR2X1_67/CTRL2 POR2X1_83/B 0.02fF
C19486 POR2X1_383/A POR2X1_343/Y 0.21fF
C19487 POR2X1_150/Y PAND2X1_205/Y 2.29fF
C19488 POR2X1_416/B POR2X1_416/CTRL2 0.01fF
C19489 PAND2X1_467/Y POR2X1_39/B 0.03fF
C19490 POR2X1_579/O PAND2X1_32/B 0.01fF
C19491 POR2X1_411/B POR2X1_272/a_76_344# 0.01fF
C19492 POR2X1_253/Y PAND2X1_242/Y 0.02fF
C19493 PAND2X1_48/A POR2X1_294/A 0.23fF
C19494 POR2X1_486/CTRL PAND2X1_57/B 0.01fF
C19495 POR2X1_411/B POR2X1_432/Y 0.03fF
C19496 PAND2X1_175/B PAND2X1_862/O 0.02fF
C19497 POR2X1_54/Y POR2X1_654/B 0.03fF
C19498 POR2X1_417/Y PAND2X1_212/CTRL 0.01fF
C19499 POR2X1_635/CTRL2 VDD 0.00fF
C19500 POR2X1_139/Y POR2X1_814/A 0.10fF
C19501 PAND2X1_239/a_76_28# POR2X1_590/A 0.01fF
C19502 POR2X1_35/B POR2X1_34/O 0.02fF
C19503 POR2X1_150/Y PAND2X1_151/CTRL 0.03fF
C19504 POR2X1_12/A POR2X1_12/O 0.01fF
C19505 POR2X1_54/Y POR2X1_5/Y 0.16fF
C19506 POR2X1_664/CTRL2 PAND2X1_72/A 0.01fF
C19507 POR2X1_20/B INPUT_0 0.08fF
C19508 POR2X1_66/B POR2X1_294/Y 0.03fF
C19509 POR2X1_842/O POR2X1_794/B 0.01fF
C19510 POR2X1_566/A POR2X1_318/O 0.04fF
C19511 POR2X1_848/A POR2X1_734/A 0.13fF
C19512 POR2X1_45/Y PAND2X1_717/A 8.18fF
C19513 POR2X1_83/B POR2X1_29/A 0.15fF
C19514 POR2X1_14/Y POR2X1_590/A 0.03fF
C19515 POR2X1_383/A POR2X1_579/m4_208_n4# 0.09fF
C19516 POR2X1_427/CTRL POR2X1_40/Y 0.01fF
C19517 POR2X1_504/Y POR2X1_48/A 0.00fF
C19518 POR2X1_278/Y POR2X1_257/A 0.18fF
C19519 POR2X1_343/Y PAND2X1_71/Y 0.05fF
C19520 POR2X1_486/CTRL2 PAND2X1_69/A 0.03fF
C19521 POR2X1_287/B POR2X1_458/a_56_344# 0.00fF
C19522 POR2X1_856/B POR2X1_436/a_76_344# 0.09fF
C19523 PAND2X1_65/B PAND2X1_59/B 0.03fF
C19524 PAND2X1_454/CTRL2 PAND2X1_446/Y 0.01fF
C19525 POR2X1_342/a_16_28# POR2X1_342/B 0.07fF
C19526 POR2X1_45/O POR2X1_23/Y 0.01fF
C19527 POR2X1_637/a_16_28# POR2X1_637/A 0.03fF
C19528 PAND2X1_219/A POR2X1_40/Y 0.04fF
C19529 POR2X1_416/Y POR2X1_412/O 0.01fF
C19530 POR2X1_446/B POR2X1_276/CTRL2 0.01fF
C19531 POR2X1_416/B PAND2X1_737/O 0.04fF
C19532 PAND2X1_39/B POR2X1_733/A 0.05fF
C19533 POR2X1_348/CTRL2 POR2X1_814/A 0.05fF
C19534 PAND2X1_139/O POR2X1_102/Y 0.03fF
C19535 POR2X1_597/Y POR2X1_761/a_16_28# 0.03fF
C19536 PAND2X1_58/A PAND2X1_525/CTRL2 0.01fF
C19537 PAND2X1_499/a_16_344# POR2X1_496/Y 0.02fF
C19538 POR2X1_706/O POR2X1_706/B 0.01fF
C19539 POR2X1_96/A POR2X1_271/O 0.02fF
C19540 PAND2X1_449/a_16_344# POR2X1_90/Y 0.01fF
C19541 POR2X1_669/B PAND2X1_381/O 0.30fF
C19542 POR2X1_682/O POR2X1_60/A 0.01fF
C19543 PAND2X1_721/B PAND2X1_721/O 0.03fF
C19544 POR2X1_35/B PAND2X1_616/CTRL 0.01fF
C19545 PAND2X1_9/Y PAND2X1_6/A 0.04fF
C19546 POR2X1_377/O POR2X1_54/Y 0.01fF
C19547 POR2X1_20/B POR2X1_619/m4_208_n4# 0.12fF
C19548 POR2X1_801/a_16_28# POR2X1_121/B 0.08fF
C19549 POR2X1_19/O POR2X1_38/B 0.00fF
C19550 PAND2X1_56/Y POR2X1_624/Y 0.10fF
C19551 POR2X1_122/A POR2X1_102/Y 0.01fF
C19552 PAND2X1_443/Y POR2X1_236/Y 0.02fF
C19553 POR2X1_174/B POR2X1_852/O 0.03fF
C19554 PAND2X1_772/a_16_344# PAND2X1_768/Y 0.03fF
C19555 PAND2X1_677/CTRL POR2X1_718/A 0.01fF
C19556 POR2X1_341/A POR2X1_702/A 0.10fF
C19557 POR2X1_196/a_16_28# PAND2X1_48/Y 0.00fF
C19558 POR2X1_333/A POR2X1_480/A 0.10fF
C19559 PAND2X1_714/A POR2X1_40/Y 0.14fF
C19560 PAND2X1_58/A POR2X1_206/A 0.02fF
C19561 PAND2X1_734/B POR2X1_32/A 0.03fF
C19562 POR2X1_65/A POR2X1_423/Y 7.73fF
C19563 POR2X1_452/Y POR2X1_730/a_16_28# 0.03fF
C19564 PAND2X1_489/O POR2X1_42/Y 0.01fF
C19565 POR2X1_52/a_16_28# POR2X1_102/Y 0.02fF
C19566 POR2X1_841/a_16_28# PAND2X1_69/A 0.01fF
C19567 POR2X1_669/B POR2X1_625/Y 0.01fF
C19568 POR2X1_442/Y VDD -0.00fF
C19569 PAND2X1_776/Y POR2X1_238/Y 0.03fF
C19570 PAND2X1_441/m4_208_n4# POR2X1_854/B 0.04fF
C19571 POR2X1_355/B POR2X1_590/A 0.06fF
C19572 POR2X1_836/a_76_344# POR2X1_578/Y 0.01fF
C19573 POR2X1_92/O INPUT_3 0.37fF
C19574 POR2X1_66/A POR2X1_563/Y 0.01fF
C19575 POR2X1_72/B PAND2X1_778/O 0.01fF
C19576 PAND2X1_793/Y PAND2X1_794/CTRL 0.01fF
C19577 POR2X1_818/Y PAND2X1_6/A 1.20fF
C19578 POR2X1_323/O POR2X1_65/A 0.01fF
C19579 POR2X1_302/A D_INPUT_0 0.07fF
C19580 POR2X1_196/CTRL2 POR2X1_814/A 0.06fF
C19581 POR2X1_489/B POR2X1_489/A 0.02fF
C19582 POR2X1_130/A POR2X1_330/Y 0.05fF
C19583 POR2X1_673/A POR2X1_35/B 0.01fF
C19584 POR2X1_301/A PAND2X1_69/A 0.05fF
C19585 PAND2X1_416/m4_208_n4# POR2X1_816/A 0.15fF
C19586 PAND2X1_445/Y POR2X1_417/Y 0.03fF
C19587 POR2X1_60/A POR2X1_372/Y 0.39fF
C19588 POR2X1_801/CTRL VDD 0.00fF
C19589 PAND2X1_810/O PAND2X1_810/B 0.01fF
C19590 PAND2X1_63/Y POR2X1_493/A 0.26fF
C19591 POR2X1_149/B PAND2X1_603/CTRL2 0.01fF
C19592 POR2X1_556/A POR2X1_116/Y 0.00fF
C19593 POR2X1_475/CTRL2 POR2X1_101/Y 0.17fF
C19594 PAND2X1_480/B POR2X1_272/O 0.02fF
C19595 PAND2X1_480/B PAND2X1_390/Y 0.05fF
C19596 POR2X1_403/CTRL POR2X1_403/B 0.01fF
C19597 POR2X1_594/Y POR2X1_83/B 0.00fF
C19598 POR2X1_13/A PAND2X1_795/O 0.03fF
C19599 POR2X1_383/A POR2X1_624/Y 0.10fF
C19600 POR2X1_78/B POR2X1_193/Y 0.11fF
C19601 PAND2X1_641/CTRL2 POR2X1_63/Y 0.01fF
C19602 PAND2X1_843/O PAND2X1_738/Y 0.23fF
C19603 POR2X1_590/A PAND2X1_536/CTRL 0.01fF
C19604 POR2X1_66/B POR2X1_554/Y 0.05fF
C19605 PAND2X1_597/CTRL VDD 0.00fF
C19606 POR2X1_49/Y POR2X1_278/Y 0.05fF
C19607 PAND2X1_474/A PAND2X1_735/O 0.05fF
C19608 PAND2X1_494/CTRL2 POR2X1_78/A 0.03fF
C19609 PAND2X1_52/B POR2X1_717/B 0.06fF
C19610 POR2X1_334/B PAND2X1_20/A 0.15fF
C19611 POR2X1_630/A POR2X1_785/A 0.03fF
C19612 POR2X1_68/O PAND2X1_69/A 0.01fF
C19613 POR2X1_494/O POR2X1_29/A 0.01fF
C19614 POR2X1_52/A PAND2X1_455/CTRL 0.01fF
C19615 PAND2X1_93/B POR2X1_318/A 0.07fF
C19616 PAND2X1_725/B VDD 0.04fF
C19617 POR2X1_829/Y VDD 0.06fF
C19618 PAND2X1_808/O POR2X1_60/A 0.02fF
C19619 POR2X1_163/A PAND2X1_725/Y 0.02fF
C19620 POR2X1_147/A POR2X1_788/A 0.01fF
C19621 POR2X1_661/B POR2X1_750/B 0.03fF
C19622 POR2X1_502/A POR2X1_718/A 0.03fF
C19623 POR2X1_49/Y POR2X1_829/A 0.01fF
C19624 POR2X1_440/Y POR2X1_434/CTRL2 0.01fF
C19625 POR2X1_502/A PAND2X1_588/CTRL 0.01fF
C19626 INPUT_1 POR2X1_709/A 0.04fF
C19627 POR2X1_509/B POR2X1_340/CTRL2 0.01fF
C19628 POR2X1_260/B POR2X1_391/O 0.01fF
C19629 POR2X1_274/A POR2X1_274/B 0.09fF
C19630 PAND2X1_205/Y PAND2X1_364/B 0.02fF
C19631 PAND2X1_784/O POR2X1_72/B 0.01fF
C19632 POR2X1_407/Y POR2X1_770/B 0.01fF
C19633 POR2X1_262/Y PAND2X1_560/B 0.00fF
C19634 PAND2X1_222/A PAND2X1_537/CTRL 0.00fF
C19635 PAND2X1_452/A PAND2X1_452/O 0.01fF
C19636 POR2X1_411/B POR2X1_394/A 0.53fF
C19637 POR2X1_302/O POR2X1_302/Y 0.01fF
C19638 PAND2X1_282/a_16_344# POR2X1_532/A 0.05fF
C19639 POR2X1_60/A POR2X1_253/Y 0.01fF
C19640 POR2X1_788/A PAND2X1_69/A 0.03fF
C19641 PAND2X1_653/Y POR2X1_102/Y 0.03fF
C19642 PAND2X1_20/A POR2X1_204/a_16_28# 0.03fF
C19643 PAND2X1_626/CTRL2 PAND2X1_69/A 0.00fF
C19644 PAND2X1_864/B PAND2X1_286/a_16_344# 0.02fF
C19645 POR2X1_445/A POR2X1_543/O 0.08fF
C19646 POR2X1_814/B POR2X1_733/A 0.01fF
C19647 POR2X1_105/Y POR2X1_717/Y 0.43fF
C19648 POR2X1_563/O POR2X1_553/Y 0.00fF
C19649 POR2X1_116/A PAND2X1_48/A 4.05fF
C19650 POR2X1_334/B POR2X1_814/B 0.07fF
C19651 PAND2X1_453/a_16_344# POR2X1_376/B 0.02fF
C19652 POR2X1_52/A PAND2X1_84/CTRL 0.01fF
C19653 PAND2X1_652/A PAND2X1_192/CTRL2 0.03fF
C19654 POR2X1_678/A PAND2X1_69/A 0.05fF
C19655 POR2X1_40/Y POR2X1_816/A 0.07fF
C19656 POR2X1_496/Y POR2X1_245/Y 0.07fF
C19657 D_INPUT_1 POR2X1_40/Y 0.03fF
C19658 POR2X1_446/B POR2X1_186/B 0.03fF
C19659 POR2X1_510/B POR2X1_590/A 0.00fF
C19660 POR2X1_54/CTRL POR2X1_54/Y 0.05fF
C19661 POR2X1_260/B POR2X1_244/Y 0.03fF
C19662 POR2X1_493/A POR2X1_260/A 0.68fF
C19663 PAND2X1_35/Y PAND2X1_734/B 0.02fF
C19664 POR2X1_402/A PAND2X1_395/CTRL2 0.01fF
C19665 POR2X1_401/a_16_28# POR2X1_401/B 0.07fF
C19666 POR2X1_834/Y PAND2X1_591/CTRL 0.28fF
C19667 POR2X1_35/B D_INPUT_1 0.09fF
C19668 PAND2X1_7/Y POR2X1_193/a_16_28# 0.03fF
C19669 POR2X1_60/A POR2X1_9/O 0.01fF
C19670 PAND2X1_794/B PAND2X1_363/Y 0.02fF
C19671 PAND2X1_562/B PAND2X1_357/Y 0.07fF
C19672 PAND2X1_661/Y POR2X1_32/A 0.03fF
C19673 PAND2X1_65/B D_GATE_222 0.10fF
C19674 POR2X1_495/Y POR2X1_236/Y 0.01fF
C19675 POR2X1_624/Y PAND2X1_71/Y 0.46fF
C19676 PAND2X1_387/O POR2X1_712/Y 0.04fF
C19677 PAND2X1_641/a_16_344# POR2X1_23/Y 0.01fF
C19678 POR2X1_128/A PAND2X1_96/B 0.04fF
C19679 POR2X1_330/Y POR2X1_573/A 0.03fF
C19680 PAND2X1_115/a_76_28# POR2X1_106/Y 0.02fF
C19681 POR2X1_516/Y PAND2X1_175/B 0.03fF
C19682 POR2X1_755/CTRL VDD -0.00fF
C19683 PAND2X1_23/Y VDD 4.59fF
C19684 POR2X1_43/B PAND2X1_276/O 0.16fF
C19685 POR2X1_648/Y POR2X1_779/O 0.01fF
C19686 PAND2X1_736/A PAND2X1_730/B 0.02fF
C19687 POR2X1_254/Y POR2X1_795/CTRL 0.02fF
C19688 POR2X1_43/B POR2X1_511/Y 0.03fF
C19689 POR2X1_62/Y PAND2X1_613/CTRL2 0.00fF
C19690 PAND2X1_818/CTRL POR2X1_42/Y 0.01fF
C19691 POR2X1_355/B POR2X1_857/B 0.03fF
C19692 PAND2X1_93/B POR2X1_574/Y 0.03fF
C19693 POR2X1_174/A POR2X1_726/Y 0.02fF
C19694 POR2X1_88/Y PAND2X1_341/CTRL 0.01fF
C19695 POR2X1_311/Y POR2X1_103/Y 0.01fF
C19696 PAND2X1_738/Y PAND2X1_552/B 0.05fF
C19697 PAND2X1_232/CTRL POR2X1_590/A 0.00fF
C19698 POR2X1_264/Y INPUT_0 0.19fF
C19699 PAND2X1_837/O POR2X1_39/B 0.17fF
C19700 PAND2X1_55/Y PAND2X1_38/CTRL 0.08fF
C19701 POR2X1_123/B PAND2X1_41/B 0.22fF
C19702 POR2X1_237/CTRL2 POR2X1_90/Y 0.01fF
C19703 PAND2X1_436/a_16_344# PAND2X1_508/Y 0.02fF
C19704 PAND2X1_55/Y POR2X1_722/Y 0.08fF
C19705 PAND2X1_725/A PAND2X1_707/CTRL2 0.01fF
C19706 POR2X1_66/A POR2X1_544/B 0.09fF
C19707 PAND2X1_319/B POR2X1_65/A 0.24fF
C19708 POR2X1_325/CTRL POR2X1_750/B 0.03fF
C19709 POR2X1_68/A POR2X1_215/O 0.01fF
C19710 POR2X1_496/Y PAND2X1_507/CTRL 0.06fF
C19711 POR2X1_62/Y POR2X1_623/CTRL2 0.06fF
C19712 INPUT_1 PAND2X1_58/A 0.32fF
C19713 PAND2X1_267/CTRL POR2X1_7/Y 0.01fF
C19714 POR2X1_114/B PAND2X1_57/B 0.00fF
C19715 POR2X1_13/A PAND2X1_357/Y 0.03fF
C19716 PAND2X1_289/CTRL POR2X1_568/B 0.03fF
C19717 PAND2X1_659/B POR2X1_816/A 0.01fF
C19718 POR2X1_675/CTRL2 POR2X1_456/B 0.00fF
C19719 PAND2X1_57/B PAND2X1_744/a_16_344# 0.02fF
C19720 POR2X1_728/B POR2X1_467/CTRL 0.00fF
C19721 PAND2X1_96/B POR2X1_206/A 0.01fF
C19722 POR2X1_344/A PAND2X1_6/Y 0.03fF
C19723 POR2X1_96/A PAND2X1_472/A 0.32fF
C19724 PAND2X1_651/Y PAND2X1_734/B 0.05fF
C19725 PAND2X1_821/a_16_344# POR2X1_857/B 0.01fF
C19726 POR2X1_102/Y POR2X1_7/a_16_28# 0.02fF
C19727 PAND2X1_823/CTRL2 PAND2X1_41/B 0.02fF
C19728 INPUT_0 PAND2X1_548/a_16_344# 0.07fF
C19729 POR2X1_137/CTRL POR2X1_391/Y 0.02fF
C19730 POR2X1_685/A PAND2X1_679/CTRL 0.01fF
C19731 POR2X1_326/A POR2X1_436/B 0.15fF
C19732 POR2X1_795/B POR2X1_785/A 1.48fF
C19733 PAND2X1_23/Y POR2X1_741/Y 1.06fF
C19734 POR2X1_70/O POR2X1_90/Y 0.01fF
C19735 PAND2X1_243/CTRL PAND2X1_734/B 0.01fF
C19736 POR2X1_814/B POR2X1_218/O 0.01fF
C19737 PAND2X1_700/CTRL PAND2X1_60/B 0.01fF
C19738 POR2X1_186/Y PAND2X1_172/O 0.09fF
C19739 PAND2X1_803/Y POR2X1_481/A 0.02fF
C19740 POR2X1_406/Y PAND2X1_560/O 0.04fF
C19741 POR2X1_140/B POR2X1_740/Y 0.03fF
C19742 POR2X1_472/CTRL2 VDD -0.00fF
C19743 D_INPUT_3 POR2X1_88/Y 0.03fF
C19744 POR2X1_763/Y POR2X1_90/Y 0.12fF
C19745 POR2X1_271/Y POR2X1_394/A 0.05fF
C19746 PAND2X1_90/A POR2X1_786/Y 0.01fF
C19747 POR2X1_296/B PAND2X1_527/O 0.00fF
C19748 PAND2X1_625/O POR2X1_741/Y 0.11fF
C19749 PAND2X1_625/a_56_28# POR2X1_740/Y 0.00fF
C19750 PAND2X1_90/A PAND2X1_316/a_56_28# 0.00fF
C19751 PAND2X1_651/Y PAND2X1_506/CTRL2 0.00fF
C19752 POR2X1_13/A POR2X1_278/A 0.06fF
C19753 POR2X1_93/A POR2X1_618/CTRL2 0.01fF
C19754 POR2X1_638/Y POR2X1_638/O 0.01fF
C19755 POR2X1_356/A POR2X1_341/Y 0.05fF
C19756 PAND2X1_23/Y PAND2X1_32/B 0.17fF
C19757 PAND2X1_140/A POR2X1_13/A 0.05fF
C19758 PAND2X1_658/A POR2X1_90/Y 0.03fF
C19759 POR2X1_802/O POR2X1_435/Y 0.04fF
C19760 POR2X1_447/B POR2X1_836/B 0.01fF
C19761 POR2X1_137/Y POR2X1_404/Y 0.03fF
C19762 PAND2X1_370/CTRL PAND2X1_566/Y 0.00fF
C19763 POR2X1_502/A POR2X1_725/Y 0.07fF
C19764 PAND2X1_41/B PAND2X1_384/O 0.00fF
C19765 PAND2X1_744/CTRL POR2X1_644/A 0.02fF
C19766 POR2X1_96/A POR2X1_527/Y 0.03fF
C19767 PAND2X1_632/CTRL INPUT_0 0.01fF
C19768 POR2X1_376/B POR2X1_394/A 1.63fF
C19769 PAND2X1_633/O POR2X1_153/Y 0.08fF
C19770 POR2X1_242/CTRL2 POR2X1_191/Y 0.12fF
C19771 POR2X1_242/CTRL POR2X1_192/B 0.28fF
C19772 D_INPUT_0 PAND2X1_358/O 0.35fF
C19773 POR2X1_16/A PAND2X1_473/Y 0.05fF
C19774 POR2X1_579/Y POR2X1_366/A 0.03fF
C19775 POR2X1_119/Y PAND2X1_786/a_16_344# 0.04fF
C19776 PAND2X1_631/CTRL2 POR2X1_93/A 0.06fF
C19777 POR2X1_532/A POR2X1_710/CTRL 0.02fF
C19778 PAND2X1_600/CTRL2 PAND2X1_72/A 0.01fF
C19779 POR2X1_383/A POR2X1_785/A 0.07fF
C19780 POR2X1_109/a_16_28# POR2X1_77/Y 0.02fF
C19781 PAND2X1_90/Y POR2X1_151/Y 0.05fF
C19782 POR2X1_57/A POR2X1_396/O 0.01fF
C19783 POR2X1_719/B VDD 0.10fF
C19784 PAND2X1_40/a_16_344# POR2X1_407/Y 0.01fF
C19785 POR2X1_855/B PAND2X1_599/CTRL2 0.01fF
C19786 POR2X1_90/Y POR2X1_73/Y 0.29fF
C19787 POR2X1_68/A PAND2X1_312/CTRL 0.01fF
C19788 D_INPUT_1 POR2X1_550/CTRL 0.00fF
C19789 POR2X1_505/Y PAND2X1_631/A 0.01fF
C19790 PAND2X1_686/O POR2X1_13/A 0.17fF
C19791 PAND2X1_206/O POR2X1_153/Y 0.15fF
C19792 POR2X1_575/B POR2X1_569/A 0.12fF
C19793 POR2X1_623/A POR2X1_55/Y 0.23fF
C19794 PAND2X1_651/Y POR2X1_229/m4_208_n4# 0.07fF
C19795 POR2X1_596/A POR2X1_770/CTRL 0.01fF
C19796 POR2X1_119/Y POR2X1_609/a_16_28# 0.07fF
C19797 PAND2X1_55/Y POR2X1_151/CTRL2 0.00fF
C19798 POR2X1_110/Y POR2X1_237/CTRL2 0.04fF
C19799 PAND2X1_414/a_16_344# POR2X1_67/Y 0.01fF
C19800 POR2X1_502/A POR2X1_559/A 0.05fF
C19801 PAND2X1_661/B POR2X1_278/A 0.02fF
C19802 PAND2X1_200/Y PAND2X1_207/A 0.01fF
C19803 PAND2X1_598/O POR2X1_394/A 0.12fF
C19804 PAND2X1_732/A POR2X1_763/Y 0.15fF
C19805 POR2X1_833/A POR2X1_404/Y 0.07fF
C19806 POR2X1_809/A VDD 0.98fF
C19807 POR2X1_83/A PAND2X1_244/B 0.01fF
C19808 PAND2X1_430/a_16_344# PAND2X1_3/B 0.01fF
C19809 POR2X1_614/A POR2X1_366/A 0.03fF
C19810 PAND2X1_362/B PAND2X1_355/a_16_344# 0.02fF
C19811 PAND2X1_216/B PAND2X1_736/Y 0.15fF
C19812 POR2X1_5/Y POR2X1_4/Y 0.23fF
C19813 POR2X1_456/B POR2X1_732/B 0.09fF
C19814 POR2X1_52/A POR2X1_394/A 0.30fF
C19815 POR2X1_8/Y PAND2X1_341/CTRL 0.00fF
C19816 POR2X1_167/CTRL2 POR2X1_73/Y 0.05fF
C19817 POR2X1_134/Y PAND2X1_854/A 0.06fF
C19818 POR2X1_43/B PAND2X1_124/O 0.04fF
C19819 POR2X1_389/A POR2X1_537/B 0.04fF
C19820 POR2X1_416/B POR2X1_748/A 0.12fF
C19821 POR2X1_566/A POR2X1_337/Y 0.11fF
C19822 POR2X1_383/A POR2X1_493/CTRL 0.01fF
C19823 PAND2X1_55/Y PAND2X1_527/CTRL2 0.03fF
C19824 POR2X1_532/A PAND2X1_528/O 0.01fF
C19825 PAND2X1_48/B POR2X1_342/CTRL2 0.01fF
C19826 PAND2X1_56/Y POR2X1_186/B 0.03fF
C19827 POR2X1_546/B POR2X1_550/B 0.02fF
C19828 VDD PAND2X1_326/B 0.02fF
C19829 PAND2X1_6/A POR2X1_751/Y 0.03fF
C19830 POR2X1_795/B POR2X1_186/B 0.07fF
C19831 PAND2X1_727/O POR2X1_90/Y 0.15fF
C19832 INPUT_1 PAND2X1_96/B 0.06fF
C19833 POR2X1_43/B POR2X1_129/Y 9.19fF
C19834 PAND2X1_26/CTRL2 POR2X1_260/A 0.00fF
C19835 POR2X1_3/O POR2X1_260/A 0.04fF
C19836 PAND2X1_732/A POR2X1_73/Y 0.01fF
C19837 POR2X1_20/CTRL POR2X1_4/Y 0.07fF
C19838 PAND2X1_686/O PAND2X1_643/Y 0.07fF
C19839 POR2X1_73/Y PAND2X1_123/a_76_28# 0.01fF
C19840 POR2X1_760/A PAND2X1_217/a_16_344# 0.02fF
C19841 POR2X1_260/A PAND2X1_670/CTRL2 0.03fF
C19842 PAND2X1_551/CTRL PAND2X1_569/B 0.01fF
C19843 POR2X1_709/O POR2X1_713/B 0.02fF
C19844 POR2X1_447/B POR2X1_294/B 0.10fF
C19845 INPUT_0 POR2X1_372/CTRL2 0.09fF
C19846 POR2X1_16/Y POR2X1_73/Y 0.01fF
C19847 POR2X1_773/B PAND2X1_60/B 0.05fF
C19848 PAND2X1_423/O PAND2X1_72/A 0.03fF
C19849 POR2X1_438/CTRL POR2X1_373/Y 0.01fF
C19850 PAND2X1_549/CTRL POR2X1_39/B 0.01fF
C19851 INPUT_1 POR2X1_248/Y 0.01fF
C19852 POR2X1_8/Y D_INPUT_3 0.03fF
C19853 PAND2X1_659/Y POR2X1_43/B 0.03fF
C19854 PAND2X1_658/A PAND2X1_185/CTRL2 0.01fF
C19855 PAND2X1_94/A PAND2X1_63/B 0.03fF
C19856 POR2X1_510/Y POR2X1_260/A 0.03fF
C19857 POR2X1_859/A POR2X1_39/B 18.05fF
C19858 POR2X1_559/a_16_28# POR2X1_559/A 0.03fF
C19859 POR2X1_123/Y POR2X1_557/B 0.01fF
C19860 POR2X1_809/A PAND2X1_32/B 0.04fF
C19861 PAND2X1_860/A PAND2X1_795/CTRL2 0.01fF
C19862 POR2X1_96/Y POR2X1_43/B 0.03fF
C19863 PAND2X1_661/B POR2X1_117/Y 0.01fF
C19864 PAND2X1_490/CTRL2 POR2X1_4/Y 0.05fF
C19865 POR2X1_248/Y POR2X1_153/Y 0.05fF
C19866 POR2X1_416/B POR2X1_79/Y 0.03fF
C19867 POR2X1_110/Y POR2X1_73/Y 0.10fF
C19868 POR2X1_294/B POR2X1_510/O 0.01fF
C19869 POR2X1_728/O PAND2X1_52/B 0.01fF
C19870 POR2X1_276/Y POR2X1_260/A 0.03fF
C19871 POR2X1_119/Y PAND2X1_852/B 0.00fF
C19872 POR2X1_389/A PAND2X1_48/A 0.03fF
C19873 PAND2X1_185/CTRL2 POR2X1_73/Y 0.00fF
C19874 POR2X1_254/Y PAND2X1_72/A 0.03fF
C19875 POR2X1_383/A POR2X1_186/B 0.21fF
C19876 POR2X1_509/CTRL2 POR2X1_857/B 0.03fF
C19877 PAND2X1_253/CTRL2 POR2X1_186/B 0.04fF
C19878 PAND2X1_175/CTRL PAND2X1_853/B 0.01fF
C19879 PAND2X1_221/Y PAND2X1_363/Y 0.02fF
C19880 POR2X1_599/A POR2X1_39/B 0.17fF
C19881 PAND2X1_434/CTRL POR2X1_129/Y 0.01fF
C19882 PAND2X1_409/O PAND2X1_52/B 0.21fF
C19883 INPUT_1 POR2X1_4/O 0.00fF
C19884 POR2X1_681/CTRL POR2X1_60/A 0.01fF
C19885 PAND2X1_653/Y POR2X1_761/A 0.00fF
C19886 POR2X1_556/A POR2X1_218/Y 0.14fF
C19887 POR2X1_499/O POR2X1_341/A 0.06fF
C19888 POR2X1_52/A POR2X1_90/CTRL2 0.00fF
C19889 POR2X1_496/a_16_28# POR2X1_260/B 0.00fF
C19890 POR2X1_43/B PAND2X1_333/Y 0.00fF
C19891 POR2X1_864/A PAND2X1_73/Y 0.01fF
C19892 POR2X1_738/A POR2X1_726/O 0.16fF
C19893 POR2X1_866/A POR2X1_260/B 0.05fF
C19894 POR2X1_41/B PAND2X1_147/CTRL2 0.12fF
C19895 POR2X1_669/B POR2X1_411/B 0.05fF
C19896 POR2X1_850/A POR2X1_458/Y 0.01fF
C19897 POR2X1_711/Y PAND2X1_32/B 0.07fF
C19898 PAND2X1_498/a_56_28# PAND2X1_72/A 0.00fF
C19899 PAND2X1_844/O POR2X1_153/Y 0.02fF
C19900 POR2X1_14/Y PAND2X1_33/CTRL 0.01fF
C19901 POR2X1_52/A POR2X1_91/CTRL 0.01fF
C19902 POR2X1_20/B POR2X1_102/Y 0.15fF
C19903 POR2X1_16/A POR2X1_7/Y 0.05fF
C19904 POR2X1_351/Y PAND2X1_52/B 0.01fF
C19905 PAND2X1_632/B PAND2X1_631/A 1.25fF
C19906 POR2X1_416/B PAND2X1_785/A 0.00fF
C19907 POR2X1_48/A PAND2X1_644/Y 0.03fF
C19908 PAND2X1_29/a_76_28# PAND2X1_52/B 0.02fF
C19909 POR2X1_341/Y PAND2X1_72/A 0.03fF
C19910 POR2X1_260/B PAND2X1_381/Y 0.01fF
C19911 POR2X1_333/Y POR2X1_191/Y 0.05fF
C19912 POR2X1_859/CTRL PAND2X1_41/B 0.03fF
C19913 POR2X1_188/A POR2X1_841/O 0.01fF
C19914 POR2X1_124/CTRL2 PAND2X1_60/B 0.01fF
C19915 D_INPUT_5 PAND2X1_425/CTRL2 0.00fF
C19916 POR2X1_519/CTRL POR2X1_416/B 0.01fF
C19917 POR2X1_817/a_76_344# POR2X1_32/A 0.01fF
C19918 POR2X1_736/A POR2X1_737/O 0.02fF
C19919 POR2X1_113/O POR2X1_768/A 0.02fF
C19920 POR2X1_863/A POR2X1_209/A 0.01fF
C19921 POR2X1_327/Y POR2X1_532/CTRL 0.28fF
C19922 POR2X1_153/Y PAND2X1_860/a_16_344# 0.04fF
C19923 POR2X1_329/A PAND2X1_364/B 0.07fF
C19924 POR2X1_187/Y POR2X1_385/Y 0.20fF
C19925 POR2X1_88/m4_208_n4# POR2X1_14/Y 0.12fF
C19926 PAND2X1_860/A PAND2X1_858/Y 0.03fF
C19927 POR2X1_192/B POR2X1_551/A 0.05fF
C19928 PAND2X1_48/B PAND2X1_85/CTRL 0.11fF
C19929 POR2X1_447/B POR2X1_567/A 0.10fF
C19930 PAND2X1_253/a_76_28# POR2X1_78/A 0.02fF
C19931 PAND2X1_789/O POR2X1_39/B 0.17fF
C19932 POR2X1_337/Y PAND2X1_167/CTRL 0.00fF
C19933 POR2X1_54/Y PAND2X1_65/B 0.03fF
C19934 POR2X1_805/Y POR2X1_792/CTRL 0.01fF
C19935 PAND2X1_358/A POR2X1_39/B 0.10fF
C19936 PAND2X1_435/CTRL POR2X1_271/B 0.01fF
C19937 POR2X1_23/Y POR2X1_49/CTRL 0.01fF
C19938 PAND2X1_796/B POR2X1_372/A 0.00fF
C19939 PAND2X1_472/B PAND2X1_33/CTRL 0.03fF
C19940 POR2X1_52/A POR2X1_816/CTRL2 0.01fF
C19941 POR2X1_814/A D_GATE_222 0.07fF
C19942 PAND2X1_779/CTRL POR2X1_39/B -0.00fF
C19943 PAND2X1_413/O POR2X1_634/A 0.00fF
C19944 POR2X1_658/CTRL POR2X1_193/A 0.03fF
C19945 POR2X1_624/Y INPUT_0 0.03fF
C19946 POR2X1_133/O POR2X1_257/A 0.01fF
C19947 POR2X1_12/A VDD 0.26fF
C19948 POR2X1_333/A PAND2X1_745/a_76_28# 0.04fF
C19949 POR2X1_320/O POR2X1_39/B 0.00fF
C19950 POR2X1_390/B POR2X1_303/B 0.02fF
C19951 POR2X1_416/B PAND2X1_730/A 0.03fF
C19952 POR2X1_491/CTRL2 POR2X1_102/Y 0.01fF
C19953 PAND2X1_852/A VDD 0.00fF
C19954 POR2X1_854/CTRL POR2X1_776/B 0.01fF
C19955 POR2X1_475/A POR2X1_479/B 0.01fF
C19956 PAND2X1_793/Y POR2X1_679/A 0.03fF
C19957 INPUT_1 POR2X1_825/Y 0.03fF
C19958 PAND2X1_65/B POR2X1_644/B 0.06fF
C19959 PAND2X1_808/Y POR2X1_20/B 0.03fF
C19960 PAND2X1_773/Y VDD 0.04fF
C19961 POR2X1_260/B PAND2X1_378/O 0.10fF
C19962 POR2X1_644/O PAND2X1_57/B 0.23fF
C19963 PAND2X1_31/O VDD 0.00fF
C19964 PAND2X1_620/Y POR2X1_422/Y 0.05fF
C19965 POR2X1_68/A POR2X1_556/A 0.08fF
C19966 POR2X1_376/B POR2X1_669/B 0.79fF
C19967 POR2X1_130/A POR2X1_558/B 0.01fF
C19968 POR2X1_445/A POR2X1_445/a_16_28# -0.00fF
C19969 POR2X1_729/CTRL POR2X1_452/Y 0.01fF
C19970 POR2X1_225/O POR2X1_5/Y 0.02fF
C19971 POR2X1_436/B POR2X1_480/A 0.02fF
C19972 POR2X1_54/Y D_INPUT_2 0.03fF
C19973 POR2X1_669/B POR2X1_430/A 0.04fF
C19974 PAND2X1_848/B INPUT_3 0.05fF
C19975 PAND2X1_612/B POR2X1_294/B 0.03fF
C19976 POR2X1_49/Y POR2X1_69/A 0.01fF
C19977 POR2X1_499/A PAND2X1_69/A 0.21fF
C19978 POR2X1_841/CTRL2 POR2X1_804/A 0.14fF
C19979 PAND2X1_248/CTRL POR2X1_404/Y 0.01fF
C19980 PAND2X1_669/CTRL2 POR2X1_668/Y 0.01fF
C19981 POR2X1_566/A PAND2X1_258/O 0.27fF
C19982 POR2X1_49/Y PAND2X1_169/Y 0.03fF
C19983 POR2X1_268/O VDD 0.00fF
C19984 POR2X1_470/O VDD 0.00fF
C19985 PAND2X1_219/A POR2X1_5/Y 0.17fF
C19986 POR2X1_48/A PAND2X1_254/Y 0.04fF
C19987 POR2X1_78/A POR2X1_788/m4_208_n4# 0.09fF
C19988 D_INPUT_0 PAND2X1_206/m4_208_n4# 0.06fF
C19989 POR2X1_659/A POR2X1_222/Y 0.01fF
C19990 POR2X1_193/A POR2X1_222/a_16_28# 0.03fF
C19991 PAND2X1_286/B VDD 0.19fF
C19992 POR2X1_866/A PAND2X1_55/Y 0.07fF
C19993 POR2X1_411/CTRL POR2X1_37/Y 0.03fF
C19994 D_INPUT_0 PAND2X1_804/B 0.12fF
C19995 POR2X1_57/A POR2X1_150/Y 0.17fF
C19996 PAND2X1_211/O PAND2X1_357/Y 0.02fF
C19997 PAND2X1_93/B PAND2X1_275/CTRL2 0.03fF
C19998 POR2X1_121/A POR2X1_655/A 0.03fF
C19999 PAND2X1_96/B PAND2X1_43/O 0.33fF
C20000 PAND2X1_73/Y POR2X1_608/a_76_344# 0.00fF
C20001 POR2X1_820/a_16_28# POR2X1_820/A 0.09fF
C20002 POR2X1_83/B POR2X1_250/O 0.02fF
C20003 POR2X1_23/Y POR2X1_238/Y 0.05fF
C20004 POR2X1_41/B POR2X1_309/CTRL 0.01fF
C20005 POR2X1_809/Y POR2X1_452/Y 0.01fF
C20006 POR2X1_49/Y POR2X1_743/CTRL 0.02fF
C20007 POR2X1_23/Y PAND2X1_658/B 0.37fF
C20008 PAND2X1_803/A PAND2X1_211/A 0.02fF
C20009 POR2X1_678/Y POR2X1_800/A 0.02fF
C20010 POR2X1_52/A POR2X1_669/B 0.32fF
C20011 POR2X1_63/Y PAND2X1_338/B 0.03fF
C20012 POR2X1_836/A POR2X1_192/Y 0.03fF
C20013 POR2X1_614/A POR2X1_809/CTRL2 0.02fF
C20014 PAND2X1_390/Y PAND2X1_473/B 0.03fF
C20015 PAND2X1_58/A PAND2X1_56/O 0.02fF
C20016 POR2X1_13/A POR2X1_667/A 3.18fF
C20017 PAND2X1_20/A POR2X1_128/CTRL2 0.01fF
C20018 PAND2X1_820/B VDD 0.11fF
C20019 POR2X1_644/CTRL2 POR2X1_644/A 0.01fF
C20020 POR2X1_43/B PAND2X1_97/a_16_344# 0.02fF
C20021 POR2X1_502/A POR2X1_811/B 0.23fF
C20022 POR2X1_240/CTRL PAND2X1_88/Y 0.01fF
C20023 POR2X1_538/CTRL POR2X1_66/A 0.01fF
C20024 POR2X1_752/Y POR2X1_585/a_76_344# 0.01fF
C20025 POR2X1_63/Y POR2X1_235/CTRL 0.01fF
C20026 POR2X1_659/A POR2X1_532/A 0.01fF
C20027 POR2X1_110/Y PAND2X1_458/CTRL2 0.01fF
C20028 POR2X1_679/B POR2X1_679/O 0.00fF
C20029 PAND2X1_96/B PAND2X1_406/O 0.02fF
C20030 POR2X1_645/a_16_28# POR2X1_330/Y 0.02fF
C20031 POR2X1_260/B POR2X1_501/B 0.03fF
C20032 POR2X1_43/B POR2X1_37/Y 4.75fF
C20033 POR2X1_603/Y POR2X1_597/A 0.17fF
C20034 POR2X1_669/B POR2X1_152/A 0.03fF
C20035 POR2X1_866/A POR2X1_407/Y 0.05fF
C20036 POR2X1_78/B PAND2X1_16/O 0.04fF
C20037 POR2X1_65/A PAND2X1_687/Y 0.03fF
C20038 PAND2X1_93/B POR2X1_219/O 0.18fF
C20039 PAND2X1_798/B POR2X1_487/CTRL 0.05fF
C20040 PAND2X1_48/Y POR2X1_483/A 0.01fF
C20041 PAND2X1_792/B POR2X1_759/Y 0.01fF
C20042 POR2X1_46/O POR2X1_46/Y 0.01fF
C20043 POR2X1_299/Y POR2X1_90/Y 0.01fF
C20044 POR2X1_72/B POR2X1_46/Y 7.23fF
C20045 POR2X1_502/A PAND2X1_387/CTRL2 0.02fF
C20046 POR2X1_76/CTRL POR2X1_569/A 0.05fF
C20047 POR2X1_287/a_76_344# POR2X1_733/A 0.04fF
C20048 POR2X1_257/A POR2X1_766/O 0.09fF
C20049 POR2X1_674/Y POR2X1_331/a_16_28# 0.02fF
C20050 POR2X1_265/a_16_28# POR2X1_73/Y 0.01fF
C20051 POR2X1_820/CTRL POR2X1_42/Y 0.15fF
C20052 POR2X1_269/m4_208_n4# POR2X1_741/Y 0.12fF
C20053 POR2X1_77/Y PAND2X1_147/CTRL2 0.01fF
C20054 POR2X1_38/B POR2X1_37/Y 1.20fF
C20055 PAND2X1_792/O POR2X1_759/Y 0.02fF
C20056 PAND2X1_240/O POR2X1_234/Y 0.00fF
C20057 PAND2X1_619/O POR2X1_260/A 0.10fF
C20058 POR2X1_356/A POR2X1_856/CTRL 0.27fF
C20059 POR2X1_356/A PAND2X1_41/B 0.06fF
C20060 POR2X1_590/A POR2X1_513/Y 0.06fF
C20061 POR2X1_671/CTRL VDD -0.00fF
C20062 POR2X1_60/A PAND2X1_339/Y 0.02fF
C20063 POR2X1_16/A POR2X1_257/A 21.55fF
C20064 POR2X1_753/Y POR2X1_90/Y 0.01fF
C20065 POR2X1_96/A PAND2X1_803/A 0.03fF
C20066 POR2X1_509/B POR2X1_579/Y 0.01fF
C20067 POR2X1_319/A POR2X1_317/A 0.01fF
C20068 D_INPUT_1 POR2X1_390/CTRL2 0.01fF
C20069 POR2X1_188/A POR2X1_662/Y 0.81fF
C20070 POR2X1_590/A POR2X1_219/B 0.01fF
C20071 PAND2X1_20/A POR2X1_562/B 0.02fF
C20072 POR2X1_791/Y POR2X1_792/B 0.12fF
C20073 POR2X1_846/B POR2X1_750/B 0.05fF
C20074 PAND2X1_6/Y PAND2X1_230/O 0.00fF
C20075 POR2X1_49/Y PAND2X1_478/CTRL2 0.01fF
C20076 PAND2X1_217/B PAND2X1_575/A 0.03fF
C20077 POR2X1_820/Y VDD 0.01fF
C20078 POR2X1_13/A POR2X1_372/O 0.18fF
C20079 PAND2X1_675/A POR2X1_40/Y 0.03fF
C20080 POR2X1_260/B POR2X1_596/CTRL2 0.01fF
C20081 POR2X1_356/A POR2X1_781/A 0.15fF
C20082 POR2X1_634/A PAND2X1_47/CTRL2 0.04fF
C20083 PAND2X1_239/CTRL POR2X1_566/B 0.33fF
C20084 PAND2X1_499/O POR2X1_293/Y 0.06fF
C20085 PAND2X1_469/B POR2X1_40/Y 0.34fF
C20086 POR2X1_482/CTRL POR2X1_7/A 0.02fF
C20087 POR2X1_814/B POR2X1_477/A 0.07fF
C20088 PAND2X1_661/B POR2X1_667/A 0.03fF
C20089 POR2X1_41/B PAND2X1_192/a_56_28# 0.00fF
C20090 PAND2X1_428/CTRL2 PAND2X1_32/B 0.01fF
C20091 POR2X1_29/A PAND2X1_670/CTRL 0.00fF
C20092 POR2X1_467/CTRL POR2X1_330/Y 0.04fF
C20093 POR2X1_68/A POR2X1_202/O 0.02fF
C20094 POR2X1_760/CTRL POR2X1_7/B 0.01fF
C20095 POR2X1_376/B PAND2X1_174/CTRL 0.09fF
C20096 PAND2X1_164/O POR2X1_776/B 0.02fF
C20097 POR2X1_276/A POR2X1_218/Y 0.07fF
C20098 POR2X1_407/A POR2X1_780/O 0.02fF
C20099 POR2X1_852/B D_GATE_222 0.03fF
C20100 PAND2X1_658/B PAND2X1_513/CTRL 0.00fF
C20101 PAND2X1_55/Y POR2X1_207/A 0.03fF
C20102 POR2X1_65/A PAND2X1_798/B 0.07fF
C20103 POR2X1_96/A PAND2X1_673/Y 0.13fF
C20104 POR2X1_79/Y PAND2X1_738/Y 0.17fF
C20105 POR2X1_96/Y PAND2X1_201/CTRL2 0.02fF
C20106 PAND2X1_232/CTRL POR2X1_66/A 0.02fF
C20107 PAND2X1_97/CTRL2 POR2X1_153/Y 0.13fF
C20108 PAND2X1_832/CTRL PAND2X1_651/Y 0.00fF
C20109 PAND2X1_401/O POR2X1_5/Y 0.17fF
C20110 POR2X1_74/a_56_344# POR2X1_23/Y 0.03fF
C20111 POR2X1_74/Y POR2X1_20/B 0.76fF
C20112 POR2X1_569/a_16_28# POR2X1_853/A 0.03fF
C20113 POR2X1_466/A POR2X1_456/B 0.09fF
C20114 POR2X1_102/Y PAND2X1_121/CTRL2 0.01fF
C20115 POR2X1_733/A VDD 1.23fF
C20116 POR2X1_174/B POR2X1_854/B 0.10fF
C20117 POR2X1_333/A POR2X1_319/Y 0.03fF
C20118 POR2X1_612/CTRL2 POR2X1_4/Y 0.01fF
C20119 PAND2X1_488/CTRL POR2X1_532/A 0.01fF
C20120 D_INPUT_2 PAND2X1_14/O 0.01fF
C20121 POR2X1_334/B VDD 4.36fF
C20122 POR2X1_271/O POR2X1_153/Y 0.18fF
C20123 POR2X1_98/CTRL POR2X1_260/A 0.00fF
C20124 PAND2X1_73/Y POR2X1_553/A 0.01fF
C20125 PAND2X1_575/A VDD 0.09fF
C20126 PAND2X1_675/a_56_28# POR2X1_250/Y 0.00fF
C20127 PAND2X1_488/O POR2X1_68/B 0.01fF
C20128 POR2X1_5/Y POR2X1_816/A 0.08fF
C20129 PAND2X1_812/CTRL VDD 0.00fF
C20130 PAND2X1_661/B POR2X1_117/O 0.01fF
C20131 PAND2X1_658/A INPUT_0 0.05fF
C20132 POR2X1_220/Y POR2X1_294/B 0.13fF
C20133 POR2X1_366/Y POR2X1_220/Y 0.07fF
C20134 PAND2X1_94/A PAND2X1_77/CTRL2 0.01fF
C20135 POR2X1_379/O PAND2X1_20/A 0.00fF
C20136 POR2X1_634/A PAND2X1_764/O 0.16fF
C20137 D_INPUT_1 POR2X1_5/Y 0.39fF
C20138 POR2X1_614/A POR2X1_786/CTRL 0.05fF
C20139 PAND2X1_140/A PAND2X1_554/O 0.00fF
C20140 POR2X1_68/A POR2X1_400/A 0.04fF
C20141 POR2X1_43/B POR2X1_406/Y 0.05fF
C20142 POR2X1_853/A POR2X1_192/Y 0.01fF
C20143 PAND2X1_568/a_76_28# POR2X1_7/B 0.01fF
C20144 POR2X1_43/B PAND2X1_715/O 0.15fF
C20145 PAND2X1_794/B VDD 1.03fF
C20146 PAND2X1_801/B POR2X1_761/Y 0.36fF
C20147 PAND2X1_207/a_16_344# PAND2X1_123/Y 0.02fF
C20148 POR2X1_294/B POR2X1_404/Y 0.03fF
C20149 POR2X1_83/B PAND2X1_392/CTRL2 0.09fF
C20150 PAND2X1_95/B PAND2X1_409/O 0.00fF
C20151 POR2X1_332/B PAND2X1_111/O 0.02fF
C20152 POR2X1_41/B PAND2X1_546/Y 0.01fF
C20153 POR2X1_103/a_16_28# POR2X1_48/A 0.00fF
C20154 POR2X1_124/B VDD 0.19fF
C20155 POR2X1_853/CTRL POR2X1_795/B 0.01fF
C20156 POR2X1_23/Y PAND2X1_657/B 0.02fF
C20157 POR2X1_66/A POR2X1_195/CTRL2 0.01fF
C20158 INPUT_2 PAND2X1_8/Y 0.02fF
C20159 POR2X1_271/B POR2X1_77/Y 0.03fF
C20160 PAND2X1_842/a_16_344# PAND2X1_388/Y 0.01fF
C20161 PAND2X1_41/B POR2X1_569/A 0.07fF
C20162 POR2X1_96/A PAND2X1_365/B 0.03fF
C20163 INPUT_0 POR2X1_73/Y 0.33fF
C20164 POR2X1_804/A PAND2X1_131/a_16_344# 0.06fF
C20165 POR2X1_48/A POR2X1_320/O 0.01fF
C20166 POR2X1_43/B POR2X1_293/Y 18.41fF
C20167 POR2X1_280/CTRL VDD 0.00fF
C20168 PAND2X1_6/Y POR2X1_307/Y 0.03fF
C20169 PAND2X1_819/O POR2X1_750/B 0.03fF
C20170 POR2X1_686/B POR2X1_596/A 0.01fF
C20171 POR2X1_41/B PAND2X1_845/O 0.00fF
C20172 POR2X1_96/A POR2X1_759/A 0.01fF
C20173 POR2X1_741/Y POR2X1_733/A 0.00fF
C20174 POR2X1_548/B POR2X1_68/A 0.01fF
C20175 PAND2X1_245/CTRL2 PAND2X1_71/Y 0.01fF
C20176 POR2X1_599/A PAND2X1_197/Y 0.03fF
C20177 POR2X1_638/Y PAND2X1_386/Y 0.10fF
C20178 POR2X1_65/A PAND2X1_691/Y 2.27fF
C20179 POR2X1_20/CTRL D_INPUT_1 0.01fF
C20180 PAND2X1_6/CTRL POR2X1_35/B 0.01fF
C20181 POR2X1_166/O PAND2X1_738/Y 0.02fF
C20182 PAND2X1_41/B POR2X1_570/Y 0.07fF
C20183 POR2X1_49/Y POR2X1_16/A 0.20fF
C20184 POR2X1_322/Y VDD 0.00fF
C20185 POR2X1_416/Y POR2X1_411/a_16_28# 0.03fF
C20186 PAND2X1_663/CTRL PAND2X1_660/B 0.01fF
C20187 PAND2X1_848/A PAND2X1_848/B 0.00fF
C20188 POR2X1_724/O POR2X1_724/A 0.02fF
C20189 PAND2X1_296/CTRL PAND2X1_359/Y 0.01fF
C20190 POR2X1_725/a_16_28# POR2X1_713/Y 0.04fF
C20191 POR2X1_355/B POR2X1_532/A 0.04fF
C20192 POR2X1_186/Y POR2X1_151/a_76_344# 0.00fF
C20193 POR2X1_57/CTRL2 POR2X1_38/Y 0.00fF
C20194 POR2X1_500/a_16_28# POR2X1_844/B 0.05fF
C20195 POR2X1_614/A POR2X1_832/B 0.18fF
C20196 POR2X1_23/Y POR2X1_184/CTRL2 0.03fF
C20197 POR2X1_311/CTRL2 POR2X1_481/A 0.01fF
C20198 PAND2X1_803/a_16_344# POR2X1_60/A 0.05fF
C20199 POR2X1_477/a_76_344# PAND2X1_52/B 0.01fF
C20200 PAND2X1_798/B PAND2X1_190/Y 0.10fF
C20201 VDD POR2X1_107/Y 0.11fF
C20202 PAND2X1_604/O PAND2X1_69/A 0.03fF
C20203 POR2X1_57/A PAND2X1_364/B 0.07fF
C20204 PAND2X1_810/CTRL2 PAND2X1_366/Y 0.03fF
C20205 POR2X1_733/A PAND2X1_32/B 0.05fF
C20206 POR2X1_45/Y POR2X1_52/Y 0.07fF
C20207 POR2X1_219/B POR2X1_214/B 0.01fF
C20208 PAND2X1_79/O POR2X1_844/B 0.02fF
C20209 PAND2X1_137/Y POR2X1_387/Y 0.10fF
C20210 PAND2X1_367/A VDD 0.00fF
C20211 POR2X1_860/A POR2X1_244/Y 0.00fF
C20212 POR2X1_13/A POR2X1_245/Y 0.23fF
C20213 POR2X1_334/B PAND2X1_32/B 0.30fF
C20214 PAND2X1_202/O POR2X1_7/A 0.02fF
C20215 POR2X1_218/O VDD 0.00fF
C20216 POR2X1_41/B PAND2X1_270/O 0.16fF
C20217 POR2X1_562/CTRL POR2X1_341/Y 0.01fF
C20218 POR2X1_377/O D_INPUT_1 0.01fF
C20219 PAND2X1_394/CTRL2 POR2X1_330/Y 0.03fF
C20220 PAND2X1_645/B POR2X1_42/Y 0.01fF
C20221 POR2X1_86/O D_INPUT_0 0.02fF
C20222 POR2X1_78/B PAND2X1_94/A 0.12fF
C20223 POR2X1_27/CTRL POR2X1_9/Y 0.01fF
C20224 POR2X1_566/A POR2X1_538/A 0.44fF
C20225 POR2X1_102/Y PAND2X1_141/O 0.03fF
C20226 PAND2X1_318/O PAND2X1_787/A 0.01fF
C20227 POR2X1_404/Y PAND2X1_111/B 0.03fF
C20228 PAND2X1_56/Y POR2X1_542/B 0.03fF
C20229 POR2X1_378/CTRL2 POR2X1_62/Y 0.01fF
C20230 POR2X1_423/Y PAND2X1_508/Y 0.89fF
C20231 POR2X1_72/B POR2X1_371/CTRL 0.01fF
C20232 POR2X1_60/A PAND2X1_352/CTRL 0.26fF
C20233 POR2X1_315/O POR2X1_90/Y 0.16fF
C20234 POR2X1_130/A POR2X1_362/A 0.03fF
C20235 POR2X1_119/Y PAND2X1_403/B 1.05fF
C20236 PAND2X1_6/Y PAND2X1_72/O 0.01fF
C20237 POR2X1_558/CTRL2 POR2X1_558/A 0.00fF
C20238 POR2X1_29/Y POR2X1_409/CTRL2 0.01fF
C20239 POR2X1_407/A PAND2X1_153/CTRL2 0.00fF
C20240 POR2X1_234/A POR2X1_411/B 0.02fF
C20241 POR2X1_566/A POR2X1_507/O 0.29fF
C20242 PAND2X1_624/A POR2X1_408/Y 0.06fF
C20243 POR2X1_334/Y POR2X1_193/Y 0.04fF
C20244 POR2X1_66/A POR2X1_181/a_16_28# 0.03fF
C20245 POR2X1_41/B PAND2X1_830/O 0.08fF
C20246 PAND2X1_117/O POR2X1_383/A 0.03fF
C20247 POR2X1_501/a_16_28# POR2X1_500/Y 0.02fF
C20248 PAND2X1_90/O POR2X1_94/A 0.06fF
C20249 POR2X1_405/a_56_344# POR2X1_737/A 0.00fF
C20250 POR2X1_804/A POR2X1_112/Y 0.11fF
C20251 PAND2X1_491/CTRL PAND2X1_96/B 0.00fF
C20252 POR2X1_124/B PAND2X1_32/B 0.80fF
C20253 POR2X1_179/CTRL POR2X1_142/Y 0.00fF
C20254 PAND2X1_6/Y POR2X1_68/B 0.07fF
C20255 POR2X1_49/Y POR2X1_599/a_16_28# 0.03fF
C20256 PAND2X1_664/O PAND2X1_645/B 0.10fF
C20257 INPUT_5 POR2X1_158/B 0.76fF
C20258 PAND2X1_220/O PAND2X1_388/Y 0.02fF
C20259 POR2X1_219/a_56_344# POR2X1_631/B 0.00fF
C20260 POR2X1_42/Y PAND2X1_154/O 0.02fF
C20261 POR2X1_777/B POR2X1_4/Y 0.00fF
C20262 PAND2X1_844/CTRL VDD 0.00fF
C20263 POR2X1_677/Y POR2X1_20/B 0.04fF
C20264 PAND2X1_192/Y PAND2X1_730/A 0.00fF
C20265 POR2X1_43/B POR2X1_408/Y 0.05fF
C20266 PAND2X1_6/A POR2X1_384/CTRL2 0.09fF
C20267 POR2X1_32/Y POR2X1_38/Y 0.05fF
C20268 POR2X1_351/Y POR2X1_350/B 0.01fF
C20269 POR2X1_41/B PAND2X1_641/Y 0.02fF
C20270 INPUT_0 POR2X1_186/B 0.03fF
C20271 POR2X1_68/A PAND2X1_393/O 0.02fF
C20272 POR2X1_9/Y POR2X1_20/B 0.54fF
C20273 POR2X1_557/A POR2X1_294/B 0.01fF
C20274 PAND2X1_55/Y POR2X1_703/A 0.10fF
C20275 D_INPUT_0 PAND2X1_332/Y 0.05fF
C20276 POR2X1_468/O POR2X1_444/Y 0.02fF
C20277 POR2X1_415/Y POR2X1_750/Y 0.01fF
C20278 D_INPUT_3 POR2X1_68/B 0.03fF
C20279 PAND2X1_94/A POR2X1_247/m4_208_n4# 0.15fF
C20280 POR2X1_380/a_16_28# POR2X1_380/A 0.03fF
C20281 POR2X1_814/A PAND2X1_417/CTRL 0.01fF
C20282 POR2X1_68/A POR2X1_180/A 0.07fF
C20283 POR2X1_271/A PAND2X1_515/O 0.06fF
C20284 PAND2X1_65/B POR2X1_4/Y 0.01fF
C20285 PAND2X1_216/B POR2X1_42/Y 0.03fF
C20286 POR2X1_383/A PAND2X1_110/m4_208_n4# 0.07fF
C20287 POR2X1_51/A POR2X1_53/O 0.03fF
C20288 POR2X1_275/CTRL2 POR2X1_129/Y 0.01fF
C20289 POR2X1_229/O POR2X1_229/Y 0.01fF
C20290 POR2X1_38/B POR2X1_408/Y 0.05fF
C20291 PAND2X1_691/Y POR2X1_761/m4_208_n4# 0.12fF
C20292 POR2X1_539/A PAND2X1_69/A 0.01fF
C20293 PAND2X1_90/CTRL2 POR2X1_546/A 0.09fF
C20294 POR2X1_283/A POR2X1_248/O 0.01fF
C20295 POR2X1_383/A POR2X1_542/B 0.03fF
C20296 PAND2X1_603/a_76_28# PAND2X1_72/A 0.02fF
C20297 PAND2X1_738/Y PAND2X1_730/A 0.05fF
C20298 POR2X1_465/B POR2X1_553/CTRL 0.01fF
C20299 PAND2X1_94/A PAND2X1_767/CTRL 0.05fF
C20300 POR2X1_365/Y POR2X1_357/CTRL 0.00fF
C20301 PAND2X1_566/Y POR2X1_176/Y 0.00fF
C20302 POR2X1_110/Y PAND2X1_785/Y 0.02fF
C20303 POR2X1_66/A PAND2X1_125/O 0.05fF
C20304 POR2X1_593/CTRL POR2X1_832/B 0.01fF
C20305 POR2X1_327/CTRL PAND2X1_48/A 0.01fF
C20306 PAND2X1_90/A PAND2X1_384/CTRL 0.12fF
C20307 PAND2X1_270/CTRL2 POR2X1_283/A 0.01fF
C20308 INPUT_1 PAND2X1_472/A 11.02fF
C20309 POR2X1_712/A POR2X1_260/A 0.59fF
C20310 PAND2X1_382/m4_208_n4# POR2X1_816/A 0.08fF
C20311 POR2X1_407/Y POR2X1_596/CTRL2 0.01fF
C20312 PAND2X1_90/Y POR2X1_568/B 0.07fF
C20313 D_INPUT_1 POR2X1_6/CTRL2 0.03fF
C20314 POR2X1_54/Y POR2X1_814/A 0.15fF
C20315 POR2X1_313/CTRL POR2X1_313/Y 0.01fF
C20316 PAND2X1_359/Y POR2X1_42/Y 0.34fF
C20317 POR2X1_569/A POR2X1_228/Y 0.10fF
C20318 PAND2X1_96/B POR2X1_758/Y 0.01fF
C20319 PAND2X1_472/A POR2X1_153/Y 0.23fF
C20320 POR2X1_81/A PAND2X1_735/a_16_344# 0.04fF
C20321 PAND2X1_348/A POR2X1_90/Y 0.07fF
C20322 POR2X1_509/O PAND2X1_41/B 0.01fF
C20323 PAND2X1_341/B POR2X1_55/Y 0.03fF
C20324 POR2X1_52/A POR2X1_41/Y 0.01fF
C20325 PAND2X1_41/B PAND2X1_72/A 0.23fF
C20326 POR2X1_54/Y POR2X1_846/Y 0.10fF
C20327 POR2X1_557/A PAND2X1_111/B 0.03fF
C20328 PAND2X1_824/B POR2X1_206/CTRL 0.06fF
C20329 POR2X1_218/A PAND2X1_48/A 0.07fF
C20330 POR2X1_730/Y PAND2X1_60/B 0.06fF
C20331 POR2X1_327/Y PAND2X1_63/Y 0.16fF
C20332 INPUT_1 POR2X1_380/Y 0.02fF
C20333 POR2X1_41/B POR2X1_680/O 0.08fF
C20334 PAND2X1_736/A PAND2X1_330/CTRL 0.02fF
C20335 POR2X1_528/Y POR2X1_744/CTRL2 0.03fF
C20336 PAND2X1_96/B POR2X1_741/A 0.04fF
C20337 POR2X1_54/CTRL D_INPUT_1 0.01fF
C20338 POR2X1_283/A POR2X1_310/Y 0.03fF
C20339 POR2X1_55/Y PAND2X1_352/Y 0.01fF
C20340 PAND2X1_714/O PAND2X1_326/B 0.02fF
C20341 D_INPUT_2 POR2X1_4/Y 0.66fF
C20342 POR2X1_625/Y POR2X1_39/B 4.12fF
C20343 PAND2X1_271/CTRL POR2X1_556/A 0.01fF
C20344 POR2X1_360/CTRL POR2X1_244/Y 0.01fF
C20345 POR2X1_274/B POR2X1_456/B 0.04fF
C20346 POR2X1_110/CTRL2 POR2X1_73/Y 0.04fF
C20347 POR2X1_294/A POR2X1_576/Y 0.03fF
C20348 POR2X1_388/CTRL POR2X1_337/Y 0.02fF
C20349 PAND2X1_213/Y PAND2X1_704/a_56_28# 0.00fF
C20350 PAND2X1_79/Y PAND2X1_71/Y 0.03fF
C20351 POR2X1_387/Y PAND2X1_853/B 0.07fF
C20352 PAND2X1_687/B POR2X1_683/Y 0.02fF
C20353 PAND2X1_81/CTRL POR2X1_4/Y 0.01fF
C20354 POR2X1_598/CTRL POR2X1_260/A 0.01fF
C20355 POR2X1_441/O POR2X1_669/B 0.03fF
C20356 POR2X1_652/a_16_28# POR2X1_652/A 0.02fF
C20357 PAND2X1_631/A POR2X1_90/Y 0.03fF
C20358 POR2X1_560/a_16_28# POR2X1_844/B 0.02fF
C20359 POR2X1_343/Y PAND2X1_498/O 0.03fF
C20360 POR2X1_119/Y PAND2X1_711/a_16_344# 0.01fF
C20361 POR2X1_730/Y POR2X1_353/A 1.86fF
C20362 POR2X1_468/B PAND2X1_52/B 0.03fF
C20363 POR2X1_520/O POR2X1_559/A 0.03fF
C20364 POR2X1_527/m4_208_n4# POR2X1_511/m4_208_n4# 0.13fF
C20365 PAND2X1_475/CTRL2 POR2X1_329/A 0.01fF
C20366 POR2X1_416/B POR2X1_628/O 0.01fF
C20367 POR2X1_212/CTRL2 POR2X1_192/B 0.09fF
C20368 POR2X1_394/A PAND2X1_124/a_16_344# 0.02fF
C20369 POR2X1_809/A POR2X1_687/A 0.04fF
C20370 POR2X1_327/Y POR2X1_260/A 0.20fF
C20371 PAND2X1_696/CTRL PAND2X1_60/B 0.01fF
C20372 POR2X1_341/A D_INPUT_0 0.03fF
C20373 POR2X1_416/B PAND2X1_6/A 0.03fF
C20374 PAND2X1_644/CTRL POR2X1_40/Y 0.01fF
C20375 PAND2X1_94/A POR2X1_294/A 0.14fF
C20376 PAND2X1_221/Y VDD 0.16fF
C20377 POR2X1_130/Y PAND2X1_72/A 0.23fF
C20378 PAND2X1_20/A POR2X1_554/B 0.02fF
C20379 POR2X1_41/B POR2X1_846/CTRL2 0.06fF
C20380 PAND2X1_23/Y POR2X1_568/A 0.06fF
C20381 PAND2X1_592/Y PAND2X1_850/CTRL2 0.00fF
C20382 POR2X1_856/B POR2X1_446/B 0.03fF
C20383 POR2X1_431/O PAND2X1_390/Y 0.01fF
C20384 PAND2X1_804/B POR2X1_173/Y 0.06fF
C20385 PAND2X1_411/O PAND2X1_52/B 0.02fF
C20386 POR2X1_510/B POR2X1_510/CTRL2 0.00fF
C20387 POR2X1_443/A POR2X1_97/A 0.03fF
C20388 POR2X1_52/A POR2X1_234/A 1.94fF
C20389 POR2X1_245/CTRL POR2X1_39/B 0.01fF
C20390 POR2X1_556/A PAND2X1_58/A 0.03fF
C20391 PAND2X1_611/CTRL POR2X1_734/A 0.06fF
C20392 PAND2X1_61/Y PAND2X1_206/B 0.00fF
C20393 PAND2X1_72/CTRL PAND2X1_72/A 0.00fF
C20394 POR2X1_509/CTRL2 POR2X1_532/A 0.01fF
C20395 POR2X1_652/O PAND2X1_72/A 0.01fF
C20396 PAND2X1_586/CTRL2 PAND2X1_48/A 0.34fF
C20397 POR2X1_651/Y POR2X1_294/B 0.03fF
C20398 POR2X1_394/A PAND2X1_716/B 0.10fF
C20399 POR2X1_62/Y PAND2X1_358/A 0.20fF
C20400 POR2X1_68/B PAND2X1_52/B 0.37fF
C20401 POR2X1_262/Y POR2X1_40/Y 0.03fF
C20402 POR2X1_557/B PAND2X1_48/A 0.03fF
C20403 POR2X1_477/B POR2X1_477/O 0.00fF
C20404 POR2X1_866/A POR2X1_807/a_16_28# 0.04fF
C20405 POR2X1_220/a_16_28# POR2X1_220/B -0.00fF
C20406 POR2X1_476/A POR2X1_66/A 0.03fF
C20407 PAND2X1_177/a_16_344# PAND2X1_72/A 0.01fF
C20408 GATE_479 POR2X1_485/Y 0.03fF
C20409 POR2X1_714/CTRL PAND2X1_72/A 0.00fF
C20410 POR2X1_166/CTRL POR2X1_167/Y 0.01fF
C20411 PAND2X1_366/a_76_28# PAND2X1_354/Y 0.01fF
C20412 POR2X1_471/A POR2X1_750/B 0.03fF
C20413 PAND2X1_217/B PAND2X1_217/O 0.02fF
C20414 POR2X1_228/Y PAND2X1_72/A 0.03fF
C20415 POR2X1_257/A POR2X1_495/O 0.03fF
C20416 POR2X1_411/B PAND2X1_340/CTRL 0.00fF
C20417 POR2X1_554/B POR2X1_325/A 0.03fF
C20418 POR2X1_499/A POR2X1_778/CTRL2 0.01fF
C20419 PAND2X1_221/Y PAND2X1_365/O 0.02fF
C20420 POR2X1_65/Y PAND2X1_61/Y 0.00fF
C20421 PAND2X1_810/B PAND2X1_366/Y 0.12fF
C20422 PAND2X1_72/A POR2X1_704/O 0.01fF
C20423 POR2X1_127/Y POR2X1_257/A 0.07fF
C20424 POR2X1_54/Y PAND2X1_55/CTRL2 0.04fF
C20425 PAND2X1_245/O POR2X1_66/A 0.02fF
C20426 POR2X1_135/a_16_28# POR2X1_394/A 0.01fF
C20427 POR2X1_68/A PAND2X1_94/Y 0.06fF
C20428 POR2X1_411/B PAND2X1_499/Y 0.03fF
C20429 INPUT_3 POR2X1_5/Y 0.45fF
C20430 PAND2X1_466/B PAND2X1_803/A 0.00fF
C20431 POR2X1_150/Y PAND2X1_84/Y 0.01fF
C20432 POR2X1_486/CTRL POR2X1_294/B 0.04fF
C20433 PAND2X1_48/B PAND2X1_53/CTRL2 0.03fF
C20434 PAND2X1_58/A PAND2X1_591/O 0.02fF
C20435 PAND2X1_820/B POR2X1_818/Y 0.01fF
C20436 PAND2X1_809/A PAND2X1_809/a_76_28# 0.02fF
C20437 POR2X1_202/B POR2X1_296/B 0.09fF
C20438 PAND2X1_217/B PAND2X1_124/Y 0.01fF
C20439 PAND2X1_299/O POR2X1_260/B 0.09fF
C20440 POR2X1_278/Y POR2X1_20/B 0.03fF
C20441 PAND2X1_571/A POR2X1_72/B 0.03fF
C20442 PAND2X1_214/CTRL POR2X1_40/Y 0.01fF
C20443 POR2X1_646/A POR2X1_294/B 0.01fF
C20444 PAND2X1_217/O VDD -0.00fF
C20445 POR2X1_174/B PAND2X1_73/Y 0.18fF
C20446 PAND2X1_309/CTRL2 POR2X1_556/A 0.08fF
C20447 POR2X1_500/A D_INPUT_0 0.02fF
C20448 POR2X1_98/B PAND2X1_234/CTRL2 0.00fF
C20449 POR2X1_641/CTRL2 POR2X1_267/A 0.00fF
C20450 POR2X1_41/B POR2X1_63/Y 0.02fF
C20451 POR2X1_54/Y POR2X1_401/B 0.04fF
C20452 POR2X1_711/Y PAND2X1_692/CTRL 0.01fF
C20453 POR2X1_470/CTRL2 POR2X1_186/Y 0.37fF
C20454 POR2X1_672/Y VDD 0.08fF
C20455 POR2X1_37/Y PAND2X1_474/A 0.07fF
C20456 POR2X1_188/A POR2X1_646/Y 0.03fF
C20457 PAND2X1_39/B POR2X1_646/CTRL -0.00fF
C20458 PAND2X1_443/O VDD 0.00fF
C20459 PAND2X1_717/A POR2X1_498/A 0.01fF
C20460 POR2X1_326/A PAND2X1_52/B 0.03fF
C20461 PAND2X1_255/O PAND2X1_60/B 0.01fF
C20462 POR2X1_460/O POR2X1_460/Y 0.02fF
C20463 POR2X1_119/Y POR2X1_416/B 0.30fF
C20464 PAND2X1_124/Y VDD 0.16fF
C20465 POR2X1_866/A POR2X1_779/a_16_28# 0.09fF
C20466 POR2X1_654/B POR2X1_78/A 11.31fF
C20467 POR2X1_334/B PAND2X1_9/Y 0.13fF
C20468 POR2X1_43/B POR2X1_275/A 0.59fF
C20469 POR2X1_65/A POR2X1_423/CTRL 0.01fF
C20470 POR2X1_452/Y POR2X1_730/CTRL2 0.01fF
C20471 POR2X1_142/CTRL2 POR2X1_49/Y 0.01fF
C20472 POR2X1_814/B POR2X1_240/B 0.02fF
C20473 PAND2X1_59/B PAND2X1_587/Y 0.06fF
C20474 PAND2X1_474/Y D_INPUT_0 0.05fF
C20475 POR2X1_257/A PAND2X1_324/Y 0.01fF
C20476 PAND2X1_39/B POR2X1_800/A -0.01fF
C20477 POR2X1_117/CTRL POR2X1_60/A 0.03fF
C20478 POR2X1_188/A POR2X1_830/a_56_344# 0.00fF
C20479 POR2X1_78/A POR2X1_5/Y 0.03fF
C20480 POR2X1_276/a_16_28# POR2X1_276/B 0.02fF
C20481 POR2X1_48/A POR2X1_625/Y 0.23fF
C20482 POR2X1_102/Y POR2X1_237/CTRL2 0.01fF
C20483 PAND2X1_104/CTRL POR2X1_814/B 0.00fF
C20484 POR2X1_13/A D_INPUT_0 0.14fF
C20485 PAND2X1_96/B POR2X1_556/A 0.11fF
C20486 POR2X1_831/CTRL2 PAND2X1_69/A 0.01fF
C20487 PAND2X1_416/CTRL2 POR2X1_816/A 0.12fF
C20488 PAND2X1_224/a_76_28# POR2X1_566/B 0.05fF
C20489 POR2X1_43/B PAND2X1_211/a_16_344# 0.01fF
C20490 PAND2X1_90/Y PAND2X1_585/CTRL2 0.01fF
C20491 PAND2X1_48/B PAND2X1_485/CTRL2 0.00fF
C20492 PAND2X1_219/A PAND2X1_723/Y 0.03fF
C20493 POR2X1_56/CTRL POR2X1_516/B 0.00fF
C20494 POR2X1_556/A POR2X1_216/CTRL2 0.01fF
C20495 PAND2X1_39/B POR2X1_702/A 0.03fF
C20496 D_INPUT_3 POR2X1_263/O 0.10fF
C20497 POR2X1_78/B POR2X1_606/Y 0.04fF
C20498 PAND2X1_659/B POR2X1_498/Y 0.12fF
C20499 POR2X1_83/B VDD 3.98fF
C20500 PAND2X1_423/CTRL2 POR2X1_807/A 0.01fF
C20501 POR2X1_502/A POR2X1_296/B 0.07fF
C20502 POR2X1_96/A PAND2X1_577/Y 0.01fF
C20503 POR2X1_102/Y PAND2X1_579/B 0.03fF
C20504 POR2X1_332/B POR2X1_241/B 0.03fF
C20505 POR2X1_13/A PAND2X1_435/Y 0.04fF
C20506 PAND2X1_394/O VDD 0.00fF
C20507 POR2X1_78/A POR2X1_724/O 0.04fF
C20508 POR2X1_709/A POR2X1_410/Y 0.01fF
C20509 PAND2X1_404/Y POR2X1_56/Y 0.03fF
C20510 POR2X1_862/CTRL2 PAND2X1_52/B 0.01fF
C20511 POR2X1_590/A PAND2X1_152/CTRL2 0.02fF
C20512 PAND2X1_478/Y PAND2X1_803/A 0.00fF
C20513 POR2X1_144/Y PAND2X1_731/B 0.02fF
C20514 POR2X1_523/Y POR2X1_849/B 0.01fF
C20515 POR2X1_23/Y PAND2X1_705/CTRL 0.01fF
C20516 POR2X1_829/O VDD 0.00fF
C20517 POR2X1_646/CTRL POR2X1_805/Y 0.02fF
C20518 PAND2X1_73/Y POR2X1_828/CTRL2 0.01fF
C20519 POR2X1_856/B POR2X1_795/B 0.19fF
C20520 POR2X1_49/Y PAND2X1_828/O 0.03fF
C20521 POR2X1_626/Y VDD 0.00fF
C20522 POR2X1_653/CTRL POR2X1_750/B 0.00fF
C20523 PAND2X1_263/a_76_28# POR2X1_94/A 0.05fF
C20524 POR2X1_270/O POR2X1_446/B 0.01fF
C20525 POR2X1_851/A POR2X1_513/Y 0.06fF
C20526 POR2X1_702/B PAND2X1_65/B 0.02fF
C20527 PAND2X1_796/B POR2X1_387/Y 0.04fF
C20528 POR2X1_65/A POR2X1_666/A 0.01fF
C20529 PAND2X1_244/CTRL2 POR2X1_293/Y 0.01fF
C20530 POR2X1_331/Y PAND2X1_730/B 0.02fF
C20531 PAND2X1_852/A PAND2X1_852/B 0.00fF
C20532 POR2X1_60/A POR2X1_252/CTRL 0.01fF
C20533 POR2X1_443/O POR2X1_568/Y 0.04fF
C20534 POR2X1_849/B PAND2X1_69/A 0.01fF
C20535 PAND2X1_476/O PAND2X1_473/Y 0.04fF
C20536 GATE_741 POR2X1_331/Y 0.01fF
C20537 POR2X1_593/B VDD 0.49fF
C20538 POR2X1_752/Y VDD 0.53fF
C20539 POR2X1_448/B POR2X1_448/A 0.00fF
C20540 POR2X1_257/A PAND2X1_549/B 0.10fF
C20541 POR2X1_467/Y POR2X1_468/B 0.06fF
C20542 POR2X1_260/B POR2X1_140/O 0.01fF
C20543 PAND2X1_217/B PAND2X1_795/B 0.03fF
C20544 POR2X1_43/B PAND2X1_61/O 0.01fF
C20545 POR2X1_334/B PAND2X1_15/O 0.03fF
C20546 POR2X1_23/O POR2X1_42/Y 0.01fF
C20547 POR2X1_298/m4_208_n4# PAND2X1_302/m4_208_n4# 0.05fF
C20548 POR2X1_505/Y POR2X1_96/A 0.35fF
C20549 POR2X1_407/A POR2X1_858/O 0.08fF
C20550 POR2X1_78/A PAND2X1_145/CTRL 0.01fF
C20551 POR2X1_681/O POR2X1_153/Y 0.05fF
C20552 POR2X1_830/Y POR2X1_733/A 0.13fF
C20553 PAND2X1_20/A PAND2X1_95/CTRL2 0.00fF
C20554 POR2X1_244/B PAND2X1_41/B 0.03fF
C20555 POR2X1_814/B POR2X1_723/CTRL 0.01fF
C20556 POR2X1_105/CTRL POR2X1_717/Y 0.01fF
C20557 POR2X1_315/m4_208_n4# PAND2X1_469/m4_208_n4# 0.13fF
C20558 POR2X1_29/Y POR2X1_409/B 0.02fF
C20559 POR2X1_519/CTRL PAND2X1_838/B 0.01fF
C20560 POR2X1_322/O POR2X1_83/B 0.01fF
C20561 POR2X1_334/B POR2X1_267/A 0.03fF
C20562 PAND2X1_793/Y PAND2X1_390/Y 0.35fF
C20563 PAND2X1_658/A POR2X1_102/Y 0.12fF
C20564 POR2X1_596/A POR2X1_678/Y 0.01fF
C20565 POR2X1_809/Y POR2X1_636/B 0.09fF
C20566 POR2X1_849/A POR2X1_550/CTRL2 0.03fF
C20567 POR2X1_60/A PAND2X1_714/m4_208_n4# 0.08fF
C20568 POR2X1_623/B PAND2X1_6/A 0.02fF
C20569 PAND2X1_20/A PAND2X1_79/a_16_344# 0.02fF
C20570 PAND2X1_417/O POR2X1_186/B 0.05fF
C20571 POR2X1_655/Y PAND2X1_55/Y 0.33fF
C20572 POR2X1_43/B POR2X1_60/A 0.13fF
C20573 POR2X1_23/Y POR2X1_387/Y 0.10fF
C20574 POR2X1_119/Y PAND2X1_608/CTRL 0.08fF
C20575 POR2X1_454/A POR2X1_569/A 0.07fF
C20576 POR2X1_695/CTRL POR2X1_23/Y 0.01fF
C20577 POR2X1_695/CTRL2 POR2X1_48/A 0.01fF
C20578 POR2X1_122/CTRL2 POR2X1_20/B 0.01fF
C20579 POR2X1_33/O D_INPUT_1 0.01fF
C20580 POR2X1_66/A POR2X1_205/A 0.01fF
C20581 PAND2X1_40/O PAND2X1_11/Y 0.01fF
C20582 POR2X1_128/A PAND2X1_55/Y 0.18fF
C20583 POR2X1_814/A POR2X1_4/Y 0.05fF
C20584 POR2X1_624/Y PAND2X1_184/CTRL2 0.01fF
C20585 PAND2X1_140/Y VDD 0.20fF
C20586 POR2X1_65/A PAND2X1_564/a_76_28# 0.01fF
C20587 POR2X1_97/CTRL POR2X1_454/A 0.01fF
C20588 POR2X1_218/Y PAND2X1_60/B 0.07fF
C20589 POR2X1_333/A POR2X1_775/O 0.05fF
C20590 POR2X1_305/Y POR2X1_748/A 0.10fF
C20591 POR2X1_383/A POR2X1_856/B 0.10fF
C20592 POR2X1_65/A POR2X1_761/CTRL2 0.03fF
C20593 PAND2X1_795/B VDD 0.28fF
C20594 POR2X1_614/A POR2X1_634/A 0.02fF
C20595 POR2X1_102/Y POR2X1_73/Y 0.16fF
C20596 PAND2X1_430/CTRL INPUT_5 0.01fF
C20597 POR2X1_451/A PAND2X1_52/B 0.00fF
C20598 POR2X1_502/A POR2X1_547/B 0.04fF
C20599 POR2X1_566/A POR2X1_471/CTRL 0.16fF
C20600 POR2X1_20/B PAND2X1_357/O 0.15fF
C20601 POR2X1_65/A PAND2X1_552/B 0.03fF
C20602 POR2X1_66/B POR2X1_804/A 0.05fF
C20603 INPUT_1 POR2X1_260/B 0.02fF
C20604 PAND2X1_785/Y INPUT_0 2.96fF
C20605 POR2X1_338/a_76_344# POR2X1_567/B 0.04fF
C20606 POR2X1_810/a_16_28# POR2X1_750/B 0.02fF
C20607 PAND2X1_84/O POR2X1_293/Y 0.03fF
C20608 POR2X1_188/A POR2X1_804/A 0.05fF
C20609 PAND2X1_436/A POR2X1_73/Y 0.07fF
C20610 POR2X1_283/A POR2X1_225/CTRL 0.01fF
C20611 POR2X1_68/A POR2X1_797/A 0.01fF
C20612 POR2X1_13/A PAND2X1_351/CTRL2 0.01fF
C20613 PAND2X1_65/B PAND2X1_744/CTRL2 0.01fF
C20614 PAND2X1_485/O POR2X1_260/A 0.01fF
C20615 POR2X1_67/A PAND2X1_154/O 0.01fF
C20616 POR2X1_47/CTRL VDD 0.00fF
C20617 POR2X1_149/B POR2X1_448/B 0.02fF
C20618 PAND2X1_55/Y POR2X1_206/A 0.01fF
C20619 POR2X1_213/B PAND2X1_146/O 0.15fF
C20620 POR2X1_490/Y POR2X1_394/A 0.03fF
C20621 PAND2X1_96/B POR2X1_202/O 0.01fF
C20622 POR2X1_752/Y PAND2X1_32/B 0.02fF
C20623 POR2X1_362/Y PAND2X1_106/O 0.14fF
C20624 POR2X1_477/A VDD 0.26fF
C20625 POR2X1_72/B POR2X1_511/CTRL2 0.01fF
C20626 POR2X1_734/A POR2X1_705/a_76_344# 0.03fF
C20627 VDD PAND2X1_709/O 0.00fF
C20628 POR2X1_566/A POR2X1_193/A 0.00fF
C20629 POR2X1_566/A POR2X1_579/Y 0.05fF
C20630 POR2X1_254/Y PAND2X1_48/B 0.28fF
C20631 POR2X1_717/CTRL POR2X1_777/B 0.01fF
C20632 POR2X1_860/A POR2X1_501/B 0.03fF
C20633 POR2X1_130/A POR2X1_572/B 0.03fF
C20634 POR2X1_508/CTRL VDD -0.00fF
C20635 POR2X1_46/Y POR2X1_7/B 0.05fF
C20636 PAND2X1_389/Y POR2X1_40/Y 0.03fF
C20637 POR2X1_23/Y PAND2X1_713/CTRL 0.01fF
C20638 POR2X1_763/A POR2X1_90/Y 0.12fF
C20639 POR2X1_785/CTRL POR2X1_785/A 0.00fF
C20640 PAND2X1_127/O POR2X1_66/A 0.05fF
C20641 POR2X1_813/Y POR2X1_83/B 0.07fF
C20642 PAND2X1_65/B POR2X1_462/B 0.03fF
C20643 PAND2X1_406/CTRL PAND2X1_48/A 0.01fF
C20644 POR2X1_59/CTRL2 POR2X1_32/A 0.03fF
C20645 PAND2X1_244/B POR2X1_102/Y 0.03fF
C20646 POR2X1_277/O POR2X1_46/Y 0.01fF
C20647 PAND2X1_65/B D_INPUT_1 0.91fF
C20648 PAND2X1_6/Y POR2X1_480/A 0.10fF
C20649 POR2X1_345/A POR2X1_197/Y 0.00fF
C20650 POR2X1_281/CTRL2 POR2X1_102/Y 0.03fF
C20651 PAND2X1_795/CTRL PAND2X1_175/B 0.01fF
C20652 POR2X1_505/Y POR2X1_7/A 0.28fF
C20653 VDD POR2X1_562/B 0.40fF
C20654 POR2X1_566/A POR2X1_545/A 0.04fF
C20655 POR2X1_102/Y PAND2X1_508/CTRL 0.02fF
C20656 PAND2X1_56/Y POR2X1_722/Y 0.03fF
C20657 POR2X1_614/A POR2X1_130/A 0.03fF
C20658 POR2X1_119/Y POR2X1_265/CTRL 0.11fF
C20659 POR2X1_423/Y POR2X1_283/A 0.06fF
C20660 POR2X1_140/B POR2X1_220/Y 0.01fF
C20661 POR2X1_479/B POR2X1_774/A 0.14fF
C20662 PAND2X1_51/O PAND2X1_47/B -0.00fF
C20663 PAND2X1_6/Y POR2X1_243/Y 0.15fF
C20664 POR2X1_49/Y PAND2X1_549/B 0.07fF
C20665 PAND2X1_651/A POR2X1_750/B 0.01fF
C20666 POR2X1_407/A POR2X1_220/Y 0.07fF
C20667 POR2X1_522/Y VDD 0.02fF
C20668 POR2X1_411/B POR2X1_39/B 0.24fF
C20669 POR2X1_83/B POR2X1_59/O 0.18fF
C20670 POR2X1_32/A PAND2X1_200/B 0.02fF
C20671 POR2X1_614/A POR2X1_566/A 0.29fF
C20672 POR2X1_186/Y POR2X1_738/A 0.05fF
C20673 POR2X1_383/A PAND2X1_386/O 0.02fF
C20674 POR2X1_231/B D_GATE_222 0.03fF
C20675 PAND2X1_372/CTRL POR2X1_778/B 0.00fF
C20676 PAND2X1_661/Y POR2X1_39/O 0.01fF
C20677 PAND2X1_94/A POR2X1_94/A 0.65fF
C20678 PAND2X1_191/a_16_344# PAND2X1_190/Y 0.07fF
C20679 POR2X1_673/O POR2X1_260/A 0.01fF
C20680 POR2X1_579/Y PAND2X1_111/O 0.00fF
C20681 PAND2X1_57/B POR2X1_644/A 0.34fF
C20682 POR2X1_730/Y POR2X1_750/B 0.03fF
C20683 POR2X1_260/B PAND2X1_136/CTRL 0.01fF
C20684 POR2X1_368/CTRL2 POR2X1_387/Y 0.05fF
C20685 POR2X1_108/Y PAND2X1_562/B 0.11fF
C20686 VDD PAND2X1_168/CTRL2 -0.00fF
C20687 PAND2X1_55/Y POR2X1_455/A 0.03fF
C20688 POR2X1_85/Y POR2X1_63/Y 0.58fF
C20689 POR2X1_313/Y POR2X1_72/B 0.03fF
C20690 PAND2X1_845/CTRL2 POR2X1_55/Y 0.01fF
C20691 POR2X1_555/B POR2X1_228/O 0.02fF
C20692 POR2X1_259/O PAND2X1_52/Y 0.01fF
C20693 POR2X1_508/a_16_28# POR2X1_857/B 0.03fF
C20694 POR2X1_471/A PAND2X1_179/m4_208_n4# 0.09fF
C20695 POR2X1_696/CTRL POR2X1_394/A 0.01fF
C20696 PAND2X1_350/CTRL2 POR2X1_88/Y 0.00fF
C20697 PAND2X1_371/CTRL PAND2X1_69/A -0.03fF
C20698 POR2X1_96/A PAND2X1_785/O 0.02fF
C20699 PAND2X1_6/Y PAND2X1_90/A 0.03fF
C20700 POR2X1_65/A POR2X1_41/CTRL2 0.03fF
C20701 PAND2X1_347/Y PAND2X1_854/A 0.02fF
C20702 POR2X1_786/a_76_344# PAND2X1_60/B 0.00fF
C20703 PAND2X1_6/A POR2X1_619/CTRL2 0.01fF
C20704 PAND2X1_319/B PAND2X1_182/A 0.17fF
C20705 PAND2X1_597/a_76_28# POR2X1_796/A 0.01fF
C20706 POR2X1_143/CTRL D_INPUT_3 0.14fF
C20707 GATE_479 PAND2X1_726/B 0.07fF
C20708 POR2X1_244/B POR2X1_228/Y 0.01fF
C20709 POR2X1_368/CTRL POR2X1_283/A 0.03fF
C20710 PAND2X1_55/Y POR2X1_435/O 0.10fF
C20711 PAND2X1_47/B PAND2X1_3/B 0.04fF
C20712 INPUT_0 PAND2X1_656/A 0.00fF
C20713 POR2X1_137/O PAND2X1_96/B 0.01fF
C20714 PAND2X1_90/Y POR2X1_151/CTRL 0.01fF
C20715 POR2X1_518/CTRL2 POR2X1_669/B 0.02fF
C20716 INPUT_1 POR2X1_381/CTRL2 0.01fF
C20717 POR2X1_193/A POR2X1_573/A 0.03fF
C20718 POR2X1_326/A POR2X1_467/Y 0.02fF
C20719 POR2X1_606/Y POR2X1_294/A 0.06fF
C20720 PAND2X1_23/Y POR2X1_840/B 0.05fF
C20721 POR2X1_90/Y PAND2X1_302/O 0.01fF
C20722 D_INPUT_2 D_INPUT_1 0.07fF
C20723 PAND2X1_737/B PAND2X1_733/Y 0.00fF
C20724 POR2X1_341/A POR2X1_715/O 0.05fF
C20725 POR2X1_516/O POR2X1_184/Y 0.01fF
C20726 POR2X1_614/A PAND2X1_111/O 0.01fF
C20727 PAND2X1_388/Y PAND2X1_553/B 0.07fF
C20728 POR2X1_775/A POR2X1_570/B 0.03fF
C20729 POR2X1_22/A POR2X1_3/CTRL2 0.01fF
C20730 PAND2X1_61/Y PAND2X1_560/B 0.00fF
C20731 POR2X1_192/Y PAND2X1_315/O 0.05fF
C20732 POR2X1_523/Y PAND2X1_69/A 0.03fF
C20733 POR2X1_700/a_16_28# PAND2X1_711/A 0.02fF
C20734 PAND2X1_762/CTRL PAND2X1_52/B 0.01fF
C20735 PAND2X1_787/A PAND2X1_724/B 0.02fF
C20736 POR2X1_614/A POR2X1_844/B 0.03fF
C20737 POR2X1_516/O PAND2X1_651/Y 0.04fF
C20738 POR2X1_481/Y PAND2X1_555/Y 0.01fF
C20739 PAND2X1_572/O PAND2X1_197/Y 0.00fF
C20740 POR2X1_814/A POR2X1_458/Y 0.03fF
C20741 PAND2X1_557/A POR2X1_385/Y 0.03fF
C20742 POR2X1_83/A PAND2X1_243/O 0.19fF
C20743 PAND2X1_152/a_16_344# PAND2X1_60/B 0.01fF
C20744 POR2X1_197/Y PAND2X1_55/Y 0.03fF
C20745 POR2X1_46/Y PAND2X1_123/CTRL 0.03fF
C20746 POR2X1_805/Y PAND2X1_759/O 0.04fF
C20747 POR2X1_454/A PAND2X1_72/A 0.03fF
C20748 D_GATE_222 PAND2X1_88/Y 0.03fF
C20749 POR2X1_57/A POR2X1_312/CTRL 0.01fF
C20750 PAND2X1_278/CTRL POR2X1_294/A 0.07fF
C20751 PAND2X1_675/A PAND2X1_388/O 0.07fF
C20752 PAND2X1_20/A POR2X1_558/m4_208_n4# 0.10fF
C20753 PAND2X1_760/CTRL2 POR2X1_260/A 0.01fF
C20754 PAND2X1_216/B PAND2X1_139/Y 0.00fF
C20755 POR2X1_96/A PAND2X1_632/B 0.07fF
C20756 POR2X1_378/A POR2X1_55/Y 0.00fF
C20757 INPUT_1 PAND2X1_673/Y 0.03fF
C20758 PAND2X1_198/Y PAND2X1_737/B 0.07fF
C20759 POR2X1_222/A POR2X1_294/B 0.03fF
C20760 POR2X1_38/B POR2X1_844/B 0.03fF
C20761 POR2X1_729/CTRL POR2X1_687/Y 0.01fF
C20762 POR2X1_489/O POR2X1_113/B 0.09fF
C20763 PAND2X1_23/Y POR2X1_544/a_16_28# 0.03fF
C20764 POR2X1_614/A PAND2X1_150/O 0.02fF
C20765 PAND2X1_737/a_16_344# POR2X1_40/Y 0.02fF
C20766 POR2X1_68/A PAND2X1_60/B 7.15fF
C20767 PAND2X1_94/A PAND2X1_110/CTRL2 0.03fF
C20768 POR2X1_51/B POR2X1_47/O 0.03fF
C20769 POR2X1_45/Y PAND2X1_349/A 0.02fF
C20770 POR2X1_219/B POR2X1_532/A 0.25fF
C20771 POR2X1_821/Y POR2X1_73/Y 0.07fF
C20772 PAND2X1_673/Y POR2X1_153/Y 1.99fF
C20773 POR2X1_464/Y POR2X1_543/CTRL 0.01fF
C20774 POR2X1_354/a_56_344# POR2X1_319/Y 0.00fF
C20775 POR2X1_7/B POR2X1_376/O 0.01fF
C20776 POR2X1_36/B POR2X1_36/CTRL 0.03fF
C20777 POR2X1_546/B POR2X1_546/CTRL 0.04fF
C20778 PAND2X1_57/B PAND2X1_701/a_16_344# 0.01fF
C20779 POR2X1_532/A POR2X1_205/A 0.07fF
C20780 INPUT_1 PAND2X1_55/Y 0.15fF
C20781 POR2X1_399/CTRL POR2X1_119/Y 0.01fF
C20782 PAND2X1_41/B PAND2X1_165/a_76_28# 0.02fF
C20783 POR2X1_271/Y POR2X1_39/B 0.01fF
C20784 POR2X1_617/Y VDD 0.09fF
C20785 POR2X1_178/Y PAND2X1_675/A 0.05fF
C20786 PAND2X1_84/Y POR2X1_150/O 0.10fF
C20787 POR2X1_78/B POR2X1_370/a_16_28# 0.00fF
C20788 POR2X1_37/Y POR2X1_90/CTRL 0.01fF
C20789 PAND2X1_23/Y POR2X1_444/Y 0.06fF
C20790 PAND2X1_48/B POR2X1_731/A 0.04fF
C20791 PAND2X1_481/CTRL POR2X1_294/B 0.01fF
C20792 POR2X1_20/B PAND2X1_269/CTRL 0.00fF
C20793 POR2X1_456/B PAND2X1_316/CTRL2 0.01fF
C20794 POR2X1_335/A POR2X1_260/A 0.87fF
C20795 POR2X1_276/A PAND2X1_96/B 0.18fF
C20796 POR2X1_643/O POR2X1_643/Y 0.00fF
C20797 PAND2X1_65/B PAND2X1_134/O 0.05fF
C20798 VDD POR2X1_357/B 0.09fF
C20799 POR2X1_532/A POR2X1_366/A 0.03fF
C20800 POR2X1_41/B PAND2X1_357/a_16_344# 0.02fF
C20801 POR2X1_346/B PAND2X1_6/Y 0.02fF
C20802 POR2X1_16/A PAND2X1_398/a_56_28# 0.00fF
C20803 PAND2X1_171/O POR2X1_776/B 0.01fF
C20804 POR2X1_68/A POR2X1_546/O 0.17fF
C20805 PAND2X1_631/A INPUT_0 0.03fF
C20806 PAND2X1_482/O POR2X1_294/B 0.03fF
C20807 POR2X1_514/Y POR2X1_574/Y 0.00fF
C20808 INPUT_6 POR2X1_1/O 0.00fF
C20809 POR2X1_376/B POR2X1_39/B 0.12fF
C20810 POR2X1_13/A PAND2X1_643/A 0.12fF
C20811 PAND2X1_551/CTRL PAND2X1_854/A 0.00fF
C20812 POR2X1_655/a_16_28# POR2X1_655/A 0.02fF
C20813 POR2X1_394/A PAND2X1_302/a_56_28# 0.00fF
C20814 PAND2X1_674/O POR2X1_186/B 0.04fF
C20815 POR2X1_68/A POR2X1_370/CTRL2 0.01fF
C20816 PAND2X1_659/Y POR2X1_494/Y 0.02fF
C20817 PAND2X1_768/Y POR2X1_77/Y 0.03fF
C20818 PAND2X1_824/B PAND2X1_69/A 0.03fF
C20819 POR2X1_81/A PAND2X1_862/B 0.01fF
C20820 PAND2X1_69/A PAND2X1_528/m4_208_n4# 0.07fF
C20821 PAND2X1_725/A PAND2X1_725/O 0.01fF
C20822 POR2X1_717/a_76_344# POR2X1_101/Y 0.02fF
C20823 POR2X1_119/Y PAND2X1_839/CTRL 0.01fF
C20824 PAND2X1_127/O POR2X1_532/A 0.04fF
C20825 POR2X1_569/O PAND2X1_52/B 0.01fF
C20826 VDD PAND2X1_841/Y 0.04fF
C20827 POR2X1_809/A PAND2X1_583/CTRL2 0.01fF
C20828 POR2X1_165/Y POR2X1_73/Y 0.01fF
C20829 PAND2X1_854/A PAND2X1_346/Y 0.02fF
C20830 POR2X1_376/B POR2X1_80/a_56_344# 0.03fF
C20831 PAND2X1_632/B POR2X1_7/A 0.03fF
C20832 POR2X1_489/O POR2X1_768/A 0.02fF
C20833 POR2X1_294/B PAND2X1_122/CTRL2 0.05fF
C20834 PAND2X1_850/Y POR2X1_275/CTRL 0.04fF
C20835 POR2X1_802/B POR2X1_532/CTRL2 0.02fF
C20836 PAND2X1_251/O POR2X1_814/A 0.19fF
C20837 PAND2X1_440/CTRL PAND2X1_580/B 0.00fF
C20838 PAND2X1_797/Y PAND2X1_714/a_16_344# 0.01fF
C20839 POR2X1_360/A PAND2X1_290/CTRL 0.05fF
C20840 POR2X1_570/B POR2X1_339/Y 0.01fF
C20841 POR2X1_16/A POR2X1_235/O 0.01fF
C20842 POR2X1_57/A PAND2X1_170/CTRL2 0.01fF
C20843 POR2X1_96/B POR2X1_96/CTRL 0.00fF
C20844 POR2X1_480/A PAND2X1_52/B 0.25fF
C20845 POR2X1_78/CTRL POR2X1_571/Y 0.01fF
C20846 PAND2X1_94/Y PAND2X1_58/A 0.01fF
C20847 PAND2X1_224/O POR2X1_590/A 0.02fF
C20848 POR2X1_52/A POR2X1_39/B 0.53fF
C20849 INPUT_1 PAND2X1_28/O -0.00fF
C20850 POR2X1_383/A POR2X1_244/Y 0.41fF
C20851 PAND2X1_69/A POR2X1_512/CTRL 0.00fF
C20852 POR2X1_669/B PAND2X1_87/CTRL 0.31fF
C20853 POR2X1_78/B POR2X1_147/a_76_344# 0.00fF
C20854 POR2X1_140/B POR2X1_554/CTRL 0.01fF
C20855 POR2X1_334/Y POR2X1_360/O 0.01fF
C20856 POR2X1_98/B POR2X1_294/A 0.00fF
C20857 POR2X1_353/a_16_28# POR2X1_353/A 0.02fF
C20858 POR2X1_109/Y POR2X1_91/Y 0.05fF
C20859 PAND2X1_348/A PAND2X1_348/CTRL 0.08fF
C20860 POR2X1_763/Y POR2X1_320/Y 0.19fF
C20861 POR2X1_327/Y POR2X1_725/Y 0.10fF
C20862 PAND2X1_726/CTRL POR2X1_39/B 0.01fF
C20863 D_GATE_222 POR2X1_568/B 0.07fF
C20864 PAND2X1_735/Y PAND2X1_332/Y 0.07fF
C20865 POR2X1_41/CTRL POR2X1_41/O -0.00fF
C20866 POR2X1_579/B POR2X1_569/A 0.02fF
C20867 PAND2X1_39/B PAND2X1_609/O 0.15fF
C20868 PAND2X1_657/a_16_344# POR2X1_329/A 0.01fF
C20869 POR2X1_361/a_16_28# PAND2X1_48/A 0.00fF
C20870 POR2X1_274/A POR2X1_624/Y 0.07fF
C20871 POR2X1_48/A POR2X1_411/B 0.32fF
C20872 PAND2X1_687/A PAND2X1_687/O -0.00fF
C20873 POR2X1_119/Y POR2X1_823/Y 0.01fF
C20874 POR2X1_278/Y PAND2X1_349/O 0.17fF
C20875 POR2X1_532/A POR2X1_532/CTRL2 0.01fF
C20876 PAND2X1_90/A PAND2X1_52/B 0.12fF
C20877 PAND2X1_93/B PAND2X1_268/CTRL 0.01fF
C20878 POR2X1_416/B POR2X1_57/a_16_28# 0.06fF
C20879 POR2X1_349/a_16_28# POR2X1_532/A 0.02fF
C20880 POR2X1_112/O PAND2X1_60/B 0.01fF
C20881 POR2X1_332/CTRL2 POR2X1_186/B 0.03fF
C20882 POR2X1_101/Y POR2X1_737/A 0.06fF
C20883 POR2X1_569/A POR2X1_571/Y 0.02fF
C20884 PAND2X1_6/Y POR2X1_716/CTRL 0.00fF
C20885 POR2X1_616/Y PAND2X1_154/O 0.02fF
C20886 POR2X1_129/O POR2X1_411/B 0.01fF
C20887 PAND2X1_213/Y PAND2X1_326/B 0.03fF
C20888 POR2X1_260/B PAND2X1_406/O 0.03fF
C20889 PAND2X1_717/A PAND2X1_168/Y 0.12fF
C20890 PAND2X1_813/CTRL2 POR2X1_266/A 0.01fF
C20891 POR2X1_326/A PAND2X1_533/CTRL2 0.00fF
C20892 PAND2X1_132/a_76_28# PAND2X1_52/B 0.01fF
C20893 PAND2X1_604/a_76_28# PAND2X1_72/A 0.02fF
C20894 POR2X1_99/A PAND2X1_86/O 0.03fF
C20895 POR2X1_651/Y PAND2X1_386/Y 0.01fF
C20896 POR2X1_68/A POR2X1_716/a_16_28# 0.02fF
C20897 PAND2X1_71/Y POR2X1_244/Y 0.03fF
C20898 POR2X1_863/A POR2X1_785/A 0.01fF
C20899 POR2X1_702/B POR2X1_814/A 0.02fF
C20900 POR2X1_191/CTRL2 POR2X1_568/Y 0.34fF
C20901 POR2X1_83/B PAND2X1_9/Y 0.03fF
C20902 POR2X1_635/CTRL POR2X1_750/B 0.01fF
C20903 PAND2X1_71/Y PAND2X1_527/CTRL2 0.01fF
C20904 POR2X1_774/A PAND2X1_48/A 0.03fF
C20905 POR2X1_97/A POR2X1_212/a_16_28# 0.03fF
C20906 PAND2X1_449/a_76_28# POR2X1_423/Y 0.01fF
C20907 PAND2X1_337/CTRL PAND2X1_336/Y 0.01fF
C20908 PAND2X1_609/O POR2X1_805/Y 0.16fF
C20909 POR2X1_614/O POR2X1_614/Y 0.11fF
C20910 POR2X1_119/Y POR2X1_122/O 0.10fF
C20911 PAND2X1_699/CTRL2 VDD -0.00fF
C20912 PAND2X1_20/A PAND2X1_609/O 0.02fF
C20913 POR2X1_83/A POR2X1_826/a_16_28# 0.02fF
C20914 POR2X1_60/A PAND2X1_407/a_76_28# 0.02fF
C20915 POR2X1_262/Y POR2X1_5/Y 0.02fF
C20916 POR2X1_137/B PAND2X1_65/B 0.13fF
C20917 POR2X1_65/A POR2X1_424/Y 3.56fF
C20918 PAND2X1_658/A POR2X1_9/Y 0.02fF
C20919 POR2X1_34/O POR2X1_34/Y 0.19fF
C20920 D_INPUT_0 POR2X1_29/A 0.11fF
C20921 POR2X1_554/B VDD 0.34fF
C20922 PAND2X1_52/B POR2X1_727/O 0.07fF
C20923 PAND2X1_208/CTRL2 PAND2X1_124/Y 0.03fF
C20924 POR2X1_153/CTRL2 POR2X1_416/B 0.06fF
C20925 POR2X1_408/Y POR2X1_90/CTRL 0.01fF
C20926 POR2X1_356/A POR2X1_466/a_16_28# 0.13fF
C20927 POR2X1_319/A PAND2X1_41/B 0.03fF
C20928 POR2X1_45/a_56_344# POR2X1_411/B 0.00fF
C20929 PAND2X1_341/B POR2X1_96/Y 0.03fF
C20930 POR2X1_677/Y POR2X1_73/Y 0.03fF
C20931 PAND2X1_48/B POR2X1_486/a_76_344# 0.01fF
C20932 POR2X1_24/CTRL POR2X1_23/Y 0.01fF
C20933 PAND2X1_96/B PAND2X1_94/Y 0.00fF
C20934 PAND2X1_620/Y POR2X1_422/O 0.02fF
C20935 PAND2X1_666/a_76_28# PAND2X1_20/A 0.02fF
C20936 POR2X1_37/Y POR2X1_609/CTRL 0.01fF
C20937 POR2X1_666/CTRL2 PAND2X1_719/Y 0.00fF
C20938 POR2X1_602/B D_INPUT_0 0.03fF
C20939 PAND2X1_19/Y POR2X1_68/B 0.01fF
C20940 POR2X1_275/CTRL2 POR2X1_275/A 0.01fF
C20941 POR2X1_696/CTRL POR2X1_669/B 0.04fF
C20942 PAND2X1_341/B POR2X1_86/a_56_344# 0.00fF
C20943 POR2X1_644/Y POR2X1_718/A 0.00fF
C20944 POR2X1_634/A POR2X1_590/A 0.03fF
C20945 POR2X1_434/O POR2X1_480/A -0.00fF
C20946 POR2X1_848/A POR2X1_625/O 0.03fF
C20947 POR2X1_462/B POR2X1_814/A 0.03fF
C20948 POR2X1_814/B POR2X1_499/O 0.01fF
C20949 POR2X1_49/Y PAND2X1_68/O 0.03fF
C20950 PAND2X1_93/B PAND2X1_65/B 0.17fF
C20951 PAND2X1_633/O PAND2X1_640/B 0.09fF
C20952 POR2X1_814/A D_INPUT_1 0.04fF
C20953 POR2X1_48/A POR2X1_376/B 0.71fF
C20954 POR2X1_718/CTRL D_INPUT_0 0.10fF
C20955 POR2X1_23/Y POR2X1_696/Y 0.02fF
C20956 POR2X1_554/B POR2X1_741/Y 0.03fF
C20957 POR2X1_692/O POR2X1_692/Y 0.00fF
C20958 POR2X1_83/B PAND2X1_208/CTRL2 0.01fF
C20959 PAND2X1_285/CTRL VDD 0.00fF
C20960 POR2X1_78/A POR2X1_777/B 0.03fF
C20961 POR2X1_244/B POR2X1_454/A 0.02fF
C20962 POR2X1_850/B POR2X1_330/Y 0.05fF
C20963 POR2X1_41/B PAND2X1_222/A 0.03fF
C20964 POR2X1_862/B POR2X1_296/B 0.02fF
C20965 PAND2X1_390/Y POR2X1_516/Y 0.03fF
C20966 POR2X1_695/Y PAND2X1_712/CTRL 0.02fF
C20967 POR2X1_48/A PAND2X1_712/O 0.04fF
C20968 PAND2X1_43/O PAND2X1_55/Y 0.01fF
C20969 POR2X1_846/Y POR2X1_816/A 0.03fF
C20970 POR2X1_3/A POR2X1_18/CTRL 0.06fF
C20971 PAND2X1_41/O POR2X1_294/B 0.01fF
C20972 POR2X1_818/Y POR2X1_415/CTRL2 0.01fF
C20973 POR2X1_462/B POR2X1_846/Y 1.23fF
C20974 PAND2X1_75/CTRL POR2X1_724/A 0.00fF
C20975 POR2X1_640/a_16_28# PAND2X1_73/Y 0.01fF
C20976 POR2X1_14/Y POR2X1_423/Y 0.03fF
C20977 POR2X1_654/B POR2X1_285/Y 0.03fF
C20978 PAND2X1_600/O POR2X1_130/A 0.04fF
C20979 POR2X1_29/O POR2X1_409/B 0.04fF
C20980 D_INPUT_2 INPUT_3 0.20fF
C20981 PAND2X1_93/B POR2X1_653/a_16_28# 0.01fF
C20982 POR2X1_863/A POR2X1_186/B 0.06fF
C20983 PAND2X1_206/A PAND2X1_101/CTRL2 0.01fF
C20984 POR2X1_341/A D_GATE_222 0.06fF
C20985 POR2X1_60/A PAND2X1_474/A 0.11fF
C20986 POR2X1_188/A POR2X1_794/B 0.03fF
C20987 POR2X1_439/CTRL2 PAND2X1_41/B 0.00fF
C20988 PAND2X1_206/B PAND2X1_350/O 0.00fF
C20989 PAND2X1_65/B POR2X1_78/A 6.60fF
C20990 POR2X1_423/O POR2X1_5/Y 0.02fF
C20991 POR2X1_855/A PAND2X1_73/Y 0.01fF
C20992 POR2X1_478/Y POR2X1_480/A 0.04fF
C20993 POR2X1_66/CTRL2 PAND2X1_39/B 0.07fF
C20994 POR2X1_658/CTRL POR2X1_532/A 0.01fF
C20995 POR2X1_558/CTRL2 POR2X1_260/B 0.01fF
C20996 D_GATE_662 POR2X1_444/B 0.06fF
C20997 PAND2X1_404/Y POR2X1_42/Y 0.02fF
C20998 PAND2X1_585/a_56_28# PAND2X1_41/B 0.00fF
C20999 POR2X1_864/O POR2X1_774/Y 0.03fF
C21000 PAND2X1_217/B PAND2X1_795/O 0.04fF
C21001 POR2X1_621/A PAND2X1_49/O 0.00fF
C21002 POR2X1_54/Y POR2X1_790/A 0.03fF
C21003 PAND2X1_23/Y POR2X1_610/O -0.00fF
C21004 POR2X1_65/A POR2X1_748/A 0.21fF
C21005 POR2X1_52/A POR2X1_48/A 0.60fF
C21006 POR2X1_163/A POR2X1_23/Y 0.11fF
C21007 POR2X1_49/Y PAND2X1_476/O 0.17fF
C21008 POR2X1_400/A POR2X1_400/B 0.06fF
C21009 POR2X1_105/a_16_28# POR2X1_814/B 0.01fF
C21010 POR2X1_240/B VDD 0.00fF
C21011 POR2X1_130/A POR2X1_590/A 0.09fF
C21012 PAND2X1_862/Y PAND2X1_860/A 0.60fF
C21013 POR2X1_344/CTRL2 PAND2X1_65/B 0.00fF
C21014 PAND2X1_6/Y POR2X1_84/B 0.02fF
C21015 PAND2X1_84/O POR2X1_60/A 0.02fF
C21016 POR2X1_302/Y POR2X1_121/B 0.02fF
C21017 POR2X1_566/A POR2X1_590/A 0.05fF
C21018 PAND2X1_317/Y POR2X1_48/A 4.55fF
C21019 POR2X1_43/B PAND2X1_444/O 0.01fF
C21020 POR2X1_48/A POR2X1_152/A 0.16fF
C21021 POR2X1_777/B POR2X1_573/CTRL 0.21fF
C21022 PAND2X1_473/Y PAND2X1_561/Y 0.04fF
C21023 POR2X1_596/A PAND2X1_39/B 0.03fF
C21024 POR2X1_48/A PAND2X1_726/CTRL 0.01fF
C21025 POR2X1_23/Y PAND2X1_726/O 0.01fF
C21026 PAND2X1_205/A POR2X1_599/A 0.00fF
C21027 POR2X1_102/Y PAND2X1_785/Y 0.00fF
C21028 POR2X1_77/Y PAND2X1_169/m4_208_n4# 0.09fF
C21029 PAND2X1_444/Y VDD 0.00fF
C21030 POR2X1_760/A PAND2X1_593/Y 0.70fF
C21031 PAND2X1_491/CTRL POR2X1_260/B 0.01fF
C21032 PAND2X1_243/B POR2X1_669/B 0.07fF
C21033 POR2X1_376/B PAND2X1_513/O 0.15fF
C21034 POR2X1_378/Y PAND2X1_58/A 0.03fF
C21035 POR2X1_65/A POR2X1_107/CTRL 0.01fF
C21036 POR2X1_241/B POR2X1_193/A 0.01fF
C21037 POR2X1_814/A POR2X1_734/m4_208_n4# 0.06fF
C21038 POR2X1_329/A POR2X1_394/A 0.10fF
C21039 POR2X1_241/B POR2X1_579/Y 0.17fF
C21040 POR2X1_188/O PAND2X1_39/B 0.01fF
C21041 POR2X1_188/A PAND2X1_108/O 0.02fF
C21042 POR2X1_307/B POR2X1_807/A 0.03fF
C21043 POR2X1_319/A PAND2X1_314/CTRL 0.01fF
C21044 PAND2X1_56/Y POR2X1_269/CTRL2 0.05fF
C21045 PAND2X1_58/A POR2X1_7/B 0.03fF
C21046 POR2X1_774/Y D_GATE_865 0.01fF
C21047 PAND2X1_66/CTRL POR2X1_38/Y 0.01fF
C21048 POR2X1_83/B PAND2X1_714/O 0.06fF
C21049 POR2X1_447/B POR2X1_837/B 0.01fF
C21050 PAND2X1_90/Y POR2X1_213/B 0.01fF
C21051 POR2X1_319/A POR2X1_714/CTRL 0.01fF
C21052 POR2X1_45/Y POR2X1_32/A 0.05fF
C21053 POR2X1_730/Y POR2X1_467/a_16_28# 0.02fF
C21054 PAND2X1_601/O PAND2X1_60/B 0.02fF
C21055 POR2X1_502/A POR2X1_186/Y 0.03fF
C21056 POR2X1_68/A PAND2X1_603/a_16_344# 0.01fF
C21057 POR2X1_16/A POR2X1_20/B 0.22fF
C21058 POR2X1_25/Y POR2X1_18/CTRL 0.00fF
C21059 POR2X1_52/A PAND2X1_512/O 0.01fF
C21060 POR2X1_309/m4_208_n4# PAND2X1_335/m4_208_n4# 0.13fF
C21061 POR2X1_309/O POR2X1_309/Y 0.01fF
C21062 POR2X1_660/Y POR2X1_513/Y 0.03fF
C21063 POR2X1_174/B POR2X1_35/Y 3.05fF
C21064 D_INPUT_3 POR2X1_23/Y 0.03fF
C21065 POR2X1_96/A PAND2X1_721/CTRL2 0.00fF
C21066 D_INPUT_0 POR2X1_500/Y 0.01fF
C21067 POR2X1_79/Y PAND2X1_740/CTRL2 0.01fF
C21068 POR2X1_287/B PAND2X1_57/B 0.06fF
C21069 POR2X1_422/a_16_28# POR2X1_93/A 0.03fF
C21070 POR2X1_72/B POR2X1_531/O 0.01fF
C21071 POR2X1_65/A POR2X1_79/Y 0.03fF
C21072 PAND2X1_39/B POR2X1_598/O 0.33fF
C21073 POR2X1_590/A POR2X1_844/B 0.04fF
C21074 POR2X1_516/CTRL2 POR2X1_60/A 0.00fF
C21075 POR2X1_840/B POR2X1_656/O 0.02fF
C21076 POR2X1_383/A POR2X1_866/A 0.01fF
C21077 POR2X1_614/A POR2X1_241/B 2.06fF
C21078 PAND2X1_266/CTRL POR2X1_7/Y 0.01fF
C21079 POR2X1_43/B PAND2X1_556/O 0.02fF
C21080 POR2X1_464/Y POR2X1_186/Y 0.03fF
C21081 PAND2X1_91/O POR2X1_568/Y 0.38fF
C21082 POR2X1_41/B PAND2X1_842/O 0.06fF
C21083 POR2X1_661/A POR2X1_711/Y 3.01fF
C21084 POR2X1_423/Y POR2X1_55/Y 0.03fF
C21085 POR2X1_74/a_16_28# POR2X1_20/B 0.03fF
C21086 POR2X1_435/Y POR2X1_794/CTRL2 0.03fF
C21087 POR2X1_264/Y POR2X1_264/O 0.01fF
C21088 PAND2X1_69/A POR2X1_720/O 0.03fF
C21089 PAND2X1_48/B PAND2X1_41/B 0.16fF
C21090 PAND2X1_862/B PAND2X1_499/Y 0.05fF
C21091 POR2X1_483/A PAND2X1_57/B 0.03fF
C21092 PAND2X1_254/Y PAND2X1_76/Y 0.01fF
C21093 PAND2X1_89/O POR2X1_61/Y 0.04fF
C21094 POR2X1_723/CTRL VDD 0.00fF
C21095 POR2X1_197/CTRL POR2X1_244/B 0.01fF
C21096 POR2X1_41/B POR2X1_692/Y 0.01fF
C21097 POR2X1_693/Y POR2X1_40/Y 0.02fF
C21098 PAND2X1_209/A PAND2X1_161/CTRL2 0.01fF
C21099 PAND2X1_73/Y POR2X1_541/O 0.02fF
C21100 PAND2X1_658/B PAND2X1_185/CTRL 0.09fF
C21101 POR2X1_702/B POR2X1_260/Y 0.16fF
C21102 POR2X1_390/B POR2X1_301/A 0.00fF
C21103 PAND2X1_787/Y POR2X1_7/B 0.01fF
C21104 POR2X1_278/Y PAND2X1_579/B 0.07fF
C21105 POR2X1_68/A POR2X1_750/B 0.35fF
C21106 POR2X1_306/Y POR2X1_43/B 0.01fF
C21107 PAND2X1_48/B POR2X1_781/A 0.20fF
C21108 POR2X1_43/B PAND2X1_639/O 0.01fF
C21109 D_INPUT_5 POR2X1_752/a_16_28# -0.00fF
C21110 POR2X1_383/A POR2X1_269/CTRL2 0.03fF
C21111 POR2X1_646/CTRL VDD -0.00fF
C21112 POR2X1_62/Y POR2X1_411/B 0.03fF
C21113 PAND2X1_61/Y POR2X1_521/CTRL2 0.01fF
C21114 POR2X1_19/CTRL POR2X1_4/Y 0.07fF
C21115 PAND2X1_736/Y PAND2X1_736/O 0.00fF
C21116 POR2X1_389/A POR2X1_606/Y 0.03fF
C21117 GATE_479 POR2X1_43/B 0.01fF
C21118 POR2X1_83/B PAND2X1_370/m4_208_n4# 0.08fF
C21119 PAND2X1_857/A POR2X1_669/B 0.03fF
C21120 POR2X1_564/Y POR2X1_566/A 0.02fF
C21121 POR2X1_38/B POR2X1_750/A 0.12fF
C21122 PAND2X1_58/A PAND2X1_60/B 6.04fF
C21123 POR2X1_555/A POR2X1_35/Y 0.00fF
C21124 POR2X1_641/CTRL PAND2X1_60/B 0.09fF
C21125 PAND2X1_340/m4_208_n4# POR2X1_42/Y 0.04fF
C21126 PAND2X1_90/Y POR2X1_805/A 0.07fF
C21127 PAND2X1_211/A POR2X1_90/Y 0.02fF
C21128 POR2X1_102/Y PAND2X1_656/A 0.10fF
C21129 POR2X1_614/A POR2X1_774/Y 0.18fF
C21130 PAND2X1_262/CTRL PAND2X1_69/A 0.01fF
C21131 POR2X1_697/Y VDD 0.43fF
C21132 POR2X1_186/Y PAND2X1_747/CTRL2 0.30fF
C21133 POR2X1_29/A PAND2X1_133/CTRL 0.01fF
C21134 POR2X1_96/A PAND2X1_191/Y 0.60fF
C21135 PAND2X1_90/Y POR2X1_712/Y 0.11fF
C21136 POR2X1_663/B POR2X1_540/Y 0.05fF
C21137 POR2X1_119/Y PAND2X1_838/B 0.05fF
C21138 POR2X1_215/O POR2X1_205/Y 0.04fF
C21139 PAND2X1_662/O PAND2X1_660/B 0.02fF
C21140 POR2X1_788/O POR2X1_788/B 0.04fF
C21141 POR2X1_39/CTRL POR2X1_38/Y 0.01fF
C21142 POR2X1_855/Y POR2X1_863/B 0.04fF
C21143 PAND2X1_859/B POR2X1_13/A 0.03fF
C21144 PAND2X1_675/A PAND2X1_347/Y 0.03fF
C21145 POR2X1_532/A POR2X1_509/B 0.02fF
C21146 POR2X1_800/A VDD 0.53fF
C21147 PAND2X1_793/Y PAND2X1_592/Y 0.03fF
C21148 POR2X1_296/B POR2X1_276/Y 0.05fF
C21149 POR2X1_96/A PAND2X1_758/O 0.04fF
C21150 PAND2X1_46/CTRL PAND2X1_111/B 0.01fF
C21151 POR2X1_496/Y PAND2X1_748/O 0.04fF
C21152 PAND2X1_56/O PAND2X1_55/Y 0.03fF
C21153 POR2X1_72/B PAND2X1_168/CTRL 0.01fF
C21154 POR2X1_102/Y PAND2X1_861/CTRL2 0.01fF
C21155 POR2X1_438/Y POR2X1_373/Y 0.08fF
C21156 POR2X1_43/B PAND2X1_636/CTRL2 0.03fF
C21157 PAND2X1_30/CTRL POR2X1_451/A 0.01fF
C21158 POR2X1_539/O POR2X1_590/A 0.01fF
C21159 POR2X1_529/Y POR2X1_40/Y 0.01fF
C21160 PAND2X1_69/A POR2X1_778/CTRL2 0.02fF
C21161 PAND2X1_357/Y VDD 1.22fF
C21162 POR2X1_65/A POR2X1_166/O 0.01fF
C21163 POR2X1_567/B POR2X1_564/B 0.37fF
C21164 POR2X1_311/Y PAND2X1_593/Y 0.03fF
C21165 POR2X1_334/B PAND2X1_80/a_76_28# 0.03fF
C21166 POR2X1_494/Y POR2X1_293/Y 0.03fF
C21167 POR2X1_185/CTRL PAND2X1_57/B 0.00fF
C21168 PAND2X1_354/A PAND2X1_854/A 0.01fF
C21169 POR2X1_52/A PAND2X1_197/Y 0.00fF
C21170 POR2X1_45/Y PAND2X1_35/Y 0.03fF
C21171 POR2X1_614/A POR2X1_155/CTRL 0.01fF
C21172 POR2X1_143/CTRL2 PAND2X1_6/A 0.03fF
C21173 POR2X1_83/A POR2X1_96/A 2.48fF
C21174 PAND2X1_380/O PAND2X1_32/B 0.03fF
C21175 POR2X1_614/A POR2X1_645/a_16_28# 0.02fF
C21176 POR2X1_708/O POR2X1_407/A 0.16fF
C21177 POR2X1_617/Y POR2X1_818/Y 0.00fF
C21178 VDD POR2X1_702/A 0.96fF
C21179 POR2X1_72/B POR2X1_527/Y 0.19fF
C21180 POR2X1_567/A POR2X1_629/CTRL -0.01fF
C21181 PAND2X1_57/B POR2X1_705/CTRL2 0.01fF
C21182 POR2X1_356/A POR2X1_775/A 0.03fF
C21183 POR2X1_180/B POR2X1_750/B 0.06fF
C21184 POR2X1_614/A PAND2X1_257/CTRL 0.01fF
C21185 POR2X1_136/O PAND2X1_480/B 0.02fF
C21186 PAND2X1_104/CTRL POR2X1_673/Y 0.03fF
C21187 POR2X1_16/A POR2X1_491/CTRL2 0.11fF
C21188 POR2X1_366/Y POR2X1_732/B 0.03fF
C21189 POR2X1_102/Y PAND2X1_348/A 0.07fF
C21190 POR2X1_670/Y POR2X1_42/Y 0.01fF
C21191 POR2X1_128/a_16_28# POR2X1_222/Y 0.01fF
C21192 PAND2X1_470/A PAND2X1_803/A 0.00fF
C21193 POR2X1_83/Y POR2X1_23/Y 0.01fF
C21194 PAND2X1_48/B POR2X1_130/Y 0.03fF
C21195 POR2X1_566/A POR2X1_336/CTRL2 0.01fF
C21196 POR2X1_278/Y POR2X1_73/Y 0.12fF
C21197 POR2X1_96/A POR2X1_90/Y 0.13fF
C21198 POR2X1_101/O POR2X1_814/B 0.01fF
C21199 PAND2X1_824/B PAND2X1_420/O 0.05fF
C21200 POR2X1_368/Y POR2X1_372/Y 0.01fF
C21201 POR2X1_707/CTRL2 PAND2X1_41/B 0.01fF
C21202 POR2X1_65/A PAND2X1_264/CTRL 0.01fF
C21203 PAND2X1_88/O POR2X1_260/A 0.01fF
C21204 PAND2X1_341/B POR2X1_37/Y 0.11fF
C21205 POR2X1_372/A POR2X1_387/Y 0.08fF
C21206 POR2X1_97/B POR2X1_97/A 0.01fF
C21207 POR2X1_278/A VDD 0.23fF
C21208 POR2X1_78/B PAND2X1_393/CTRL 0.01fF
C21209 POR2X1_646/CTRL PAND2X1_32/B 0.03fF
C21210 POR2X1_391/Y PAND2X1_132/O 0.05fF
C21211 POR2X1_130/A POR2X1_361/CTRL 0.10fF
C21212 POR2X1_188/A PAND2X1_701/CTRL2 0.09fF
C21213 POR2X1_102/Y POR2X1_300/Y 0.04fF
C21214 PAND2X1_140/A VDD 0.55fF
C21215 POR2X1_45/Y POR2X1_184/Y 0.02fF
C21216 POR2X1_856/O POR2X1_260/A 0.03fF
C21217 POR2X1_435/Y PAND2X1_60/B 0.07fF
C21218 POR2X1_483/B POR2X1_228/Y 0.12fF
C21219 POR2X1_596/A POR2X1_513/B 0.05fF
C21220 POR2X1_809/A POR2X1_866/CTRL2 0.01fF
C21221 POR2X1_582/O INPUT_5 0.01fF
C21222 PAND2X1_445/CTRL2 POR2X1_90/Y 0.01fF
C21223 POR2X1_416/B POR2X1_12/A 8.06fF
C21224 POR2X1_528/Y VDD 0.72fF
C21225 POR2X1_115/a_16_28# POR2X1_112/Y 0.01fF
C21226 POR2X1_113/A POR2X1_640/Y 0.01fF
C21227 POR2X1_489/B POR2X1_294/A 0.01fF
C21228 POR2X1_302/Y POR2X1_383/A 0.04fF
C21229 POR2X1_68/A PAND2X1_72/CTRL2 0.38fF
C21230 POR2X1_407/A POR2X1_114/B 0.03fF
C21231 PAND2X1_832/CTRL2 POR2X1_153/Y 0.00fF
C21232 POR2X1_315/Y PAND2X1_556/B 0.07fF
C21233 POR2X1_840/B POR2X1_733/A 0.10fF
C21234 PAND2X1_221/CTRL2 PAND2X1_730/A 0.00fF
C21235 POR2X1_740/Y POR2X1_731/O 0.00fF
C21236 PAND2X1_470/m4_208_n4# POR2X1_418/m4_208_n4# 0.05fF
C21237 PAND2X1_473/Y PAND2X1_717/Y 0.03fF
C21238 POR2X1_62/Y PAND2X1_459/CTRL2 0.01fF
C21239 POR2X1_154/CTRL POR2X1_855/B 0.01fF
C21240 POR2X1_741/Y POR2X1_702/A 0.06fF
C21241 PAND2X1_212/B PAND2X1_352/B 0.00fF
C21242 POR2X1_800/A PAND2X1_32/B 0.03fF
C21243 PAND2X1_90/a_76_28# POR2X1_590/A 0.02fF
C21244 POR2X1_96/CTRL POR2X1_236/Y 0.02fF
C21245 PAND2X1_663/CTRL VDD 0.00fF
C21246 PAND2X1_319/B POR2X1_55/Y 0.00fF
C21247 PAND2X1_566/a_16_344# PAND2X1_211/A 0.03fF
C21248 PAND2X1_613/CTRL PAND2X1_52/B 0.11fF
C21249 PAND2X1_96/B POR2X1_574/CTRL 0.01fF
C21250 PAND2X1_735/Y PAND2X1_510/B 0.02fF
C21251 PAND2X1_631/A POR2X1_102/Y 0.03fF
C21252 PAND2X1_90/Y POR2X1_520/B 0.00fF
C21253 PAND2X1_55/Y PAND2X1_312/CTRL 0.11fF
C21254 POR2X1_780/CTRL POR2X1_294/A 0.04fF
C21255 PAND2X1_48/B POR2X1_228/Y 0.03fF
C21256 POR2X1_536/CTRL POR2X1_13/A 0.03fF
C21257 POR2X1_415/O POR2X1_750/Y 0.01fF
C21258 INPUT_1 POR2X1_58/a_76_344# 0.01fF
C21259 PAND2X1_865/Y POR2X1_60/A 0.07fF
C21260 PAND2X1_48/Y POR2X1_186/B 0.01fF
C21261 POR2X1_804/A PAND2X1_311/CTRL2 0.31fF
C21262 POR2X1_68/A PAND2X1_424/O 0.09fF
C21263 PAND2X1_47/CTRL PAND2X1_32/B 0.01fF
C21264 POR2X1_702/A PAND2X1_32/B 0.19fF
C21265 POR2X1_538/a_16_28# PAND2X1_69/A 0.02fF
C21266 POR2X1_389/CTRL POR2X1_725/Y 0.04fF
C21267 PAND2X1_531/CTRL2 POR2X1_547/B 0.00fF
C21268 PAND2X1_90/Y POR2X1_543/m4_208_n4# 0.03fF
C21269 POR2X1_22/CTRL POR2X1_260/A 0.03fF
C21270 PAND2X1_6/A POR2X1_376/A 0.01fF
C21271 INPUT_2 POR2X1_73/Y 0.00fF
C21272 POR2X1_65/A PAND2X1_730/A 0.03fF
C21273 POR2X1_186/Y POR2X1_188/Y 0.03fF
C21274 POR2X1_62/Y POR2X1_376/B 0.05fF
C21275 POR2X1_112/O POR2X1_750/B 0.02fF
C21276 POR2X1_383/A POR2X1_861/CTRL 0.01fF
C21277 PAND2X1_830/Y PAND2X1_114/O 0.03fF
C21278 PAND2X1_859/B PAND2X1_510/B 0.04fF
C21279 POR2X1_458/CTRL POR2X1_343/B 0.01fF
C21280 PAND2X1_594/O POR2X1_711/Y 0.05fF
C21281 POR2X1_432/CTRL POR2X1_77/Y 0.03fF
C21282 PAND2X1_275/CTRL POR2X1_569/A 0.06fF
C21283 POR2X1_43/B PAND2X1_175/B 0.03fF
C21284 PAND2X1_798/B POR2X1_283/A 0.07fF
C21285 POR2X1_38/B POR2X1_380/m4_208_n4# 0.09fF
C21286 PAND2X1_484/CTRL2 PAND2X1_57/B 0.02fF
C21287 POR2X1_140/B POR2X1_222/A 0.01fF
C21288 PAND2X1_451/O VDD 0.00fF
C21289 PAND2X1_810/a_16_344# POR2X1_7/B 0.02fF
C21290 POR2X1_516/CTRL2 POR2X1_516/A 0.01fF
C21291 PAND2X1_547/CTRL2 POR2X1_527/Y 0.01fF
C21292 PAND2X1_4/O POR2X1_38/B 0.04fF
C21293 POR2X1_56/B PAND2X1_308/Y 0.02fF
C21294 POR2X1_46/Y PAND2X1_560/B 0.03fF
C21295 PAND2X1_855/CTRL PAND2X1_854/A 0.01fF
C21296 PAND2X1_96/B PAND2X1_60/B 3.22fF
C21297 PAND2X1_390/Y POR2X1_589/O 0.01fF
C21298 PAND2X1_48/B PAND2X1_103/a_76_28# 0.02fF
C21299 POR2X1_567/A POR2X1_741/a_16_28# 0.03fF
C21300 PAND2X1_341/A PAND2X1_338/B 0.03fF
C21301 POR2X1_7/A POR2X1_90/Y 0.06fF
C21302 POR2X1_507/O D_GATE_741 0.33fF
C21303 POR2X1_860/CTRL2 POR2X1_218/A 0.00fF
C21304 POR2X1_860/O POR2X1_572/B 0.01fF
C21305 POR2X1_750/B POR2X1_169/A 0.05fF
C21306 POR2X1_45/Y PAND2X1_196/a_16_344# 0.02fF
C21307 POR2X1_532/A PAND2X1_534/CTRL2 0.01fF
C21308 PAND2X1_56/Y POR2X1_703/A 0.34fF
C21309 PAND2X1_96/B POR2X1_758/a_16_28# 0.05fF
C21310 PAND2X1_545/Y PAND2X1_551/A 0.02fF
C21311 PAND2X1_90/A POR2X1_216/Y 0.08fF
C21312 POR2X1_137/B POR2X1_814/A 0.07fF
C21313 POR2X1_383/A POR2X1_501/B 0.06fF
C21314 POR2X1_569/A POR2X1_112/Y 0.07fF
C21315 POR2X1_267/Y POR2X1_276/Y 0.00fF
C21316 D_INPUT_5 D_INPUT_7 0.03fF
C21317 PAND2X1_812/A GATE_741 0.04fF
C21318 POR2X1_580/O POR2X1_191/Y 0.06fF
C21319 POR2X1_356/A POR2X1_339/Y 0.05fF
C21320 PAND2X1_23/Y PAND2X1_481/O 0.02fF
C21321 POR2X1_220/A POR2X1_162/Y 0.04fF
C21322 PAND2X1_542/CTRL2 PAND2X1_552/B -0.00fF
C21323 POR2X1_201/Y PAND2X1_88/Y 0.01fF
C21324 POR2X1_110/Y POR2X1_96/A 0.11fF
C21325 PAND2X1_793/Y POR2X1_767/CTRL2 0.01fF
C21326 POR2X1_52/A POR2X1_62/Y 0.00fF
C21327 POR2X1_283/A POR2X1_310/a_16_28# 0.11fF
C21328 POR2X1_55/Y PAND2X1_357/CTRL2 0.02fF
C21329 POR2X1_99/B POR2X1_244/B 1.19fF
C21330 PAND2X1_382/a_76_28# PAND2X1_69/A 0.02fF
C21331 POR2X1_569/a_76_344# POR2X1_568/B 0.02fF
C21332 POR2X1_72/CTRL2 PAND2X1_659/B 0.00fF
C21333 POR2X1_625/CTRL POR2X1_39/B 0.01fF
C21334 POR2X1_336/m4_208_n4# POR2X1_538/A 0.03fF
C21335 POR2X1_541/CTRL2 POR2X1_456/B 0.01fF
C21336 PAND2X1_850/Y INPUT_0 0.01fF
C21337 POR2X1_447/B POR2X1_776/B 0.03fF
C21338 POR2X1_567/B POR2X1_440/O 0.02fF
C21339 POR2X1_323/Y PAND2X1_325/O 0.00fF
C21340 PAND2X1_31/CTRL D_INPUT_7 0.01fF
C21341 PAND2X1_341/B POR2X1_293/Y 0.03fF
C21342 PAND2X1_738/Y PAND2X1_326/B 0.05fF
C21343 PAND2X1_96/B POR2X1_353/A 0.03fF
C21344 POR2X1_554/Y POR2X1_540/Y 0.63fF
C21345 PAND2X1_96/B POR2X1_332/O 0.01fF
C21346 POR2X1_845/a_16_28# POR2X1_7/A 0.03fF
C21347 POR2X1_319/O POR2X1_191/Y 0.06fF
C21348 POR2X1_316/Y POR2X1_13/A 0.04fF
C21349 POR2X1_652/CTRL2 POR2X1_652/A 0.00fF
C21350 POR2X1_493/B PAND2X1_60/B 0.04fF
C21351 PAND2X1_858/O POR2X1_43/B 0.17fF
C21352 INPUT_0 PAND2X1_102/O 0.17fF
C21353 POR2X1_866/A POR2X1_648/Y 4.11fF
C21354 POR2X1_834/Y POR2X1_513/O 0.04fF
C21355 PAND2X1_531/CTRL PAND2X1_32/B 0.00fF
C21356 PAND2X1_190/Y PAND2X1_730/A 0.00fF
C21357 POR2X1_108/O PAND2X1_348/A 0.02fF
C21358 PAND2X1_93/B POR2X1_814/A 1.32fF
C21359 POR2X1_508/B POR2X1_508/O 0.01fF
C21360 POR2X1_57/A POR2X1_394/A 0.64fF
C21361 POR2X1_9/Y POR2X1_753/Y 0.18fF
C21362 PAND2X1_48/B PAND2X1_122/O 0.15fF
C21363 PAND2X1_48/B PAND2X1_665/O 0.01fF
C21364 POR2X1_638/Y PAND2X1_48/A 0.10fF
C21365 PAND2X1_763/CTRL PAND2X1_52/B 0.01fF
C21366 POR2X1_43/B PAND2X1_500/CTRL 0.01fF
C21367 PAND2X1_643/O PAND2X1_643/A 0.03fF
C21368 POR2X1_829/A PAND2X1_207/A 0.00fF
C21369 POR2X1_741/CTRL POR2X1_741/Y 0.00fF
C21370 POR2X1_416/B PAND2X1_668/CTRL2 0.04fF
C21371 POR2X1_130/CTRL POR2X1_141/A 0.01fF
C21372 GATE_222 POR2X1_283/Y 0.63fF
C21373 POR2X1_68/B PAND2X1_527/O 0.15fF
C21374 PAND2X1_6/Y POR2X1_691/A 0.00fF
C21375 POR2X1_76/B POR2X1_274/Y 0.23fF
C21376 POR2X1_260/B POR2X1_556/A 0.15fF
C21377 POR2X1_348/CTRL POR2X1_334/Y 0.03fF
C21378 POR2X1_407/Y PAND2X1_328/O 0.02fF
C21379 POR2X1_56/B POR2X1_77/Y 0.10fF
C21380 POR2X1_669/B POR2X1_329/A 0.07fF
C21381 PAND2X1_119/a_16_344# POR2X1_294/A 0.04fF
C21382 POR2X1_78/A POR2X1_814/A 0.38fF
C21383 PAND2X1_804/B POR2X1_173/CTRL 0.08fF
C21384 POR2X1_502/A POR2X1_717/B 0.01fF
C21385 POR2X1_609/Y POR2X1_411/A 0.02fF
C21386 PAND2X1_393/CTRL POR2X1_294/A 0.01fF
C21387 PAND2X1_366/A PAND2X1_354/Y 0.05fF
C21388 POR2X1_180/CTRL2 POR2X1_180/A 0.01fF
C21389 POR2X1_188/CTRL2 POR2X1_188/Y 0.03fF
C21390 PAND2X1_831/Y POR2X1_119/Y 0.03fF
C21391 POR2X1_84/Y POR2X1_4/Y 0.02fF
C21392 PAND2X1_138/CTRL POR2X1_7/A 0.01fF
C21393 PAND2X1_632/A PAND2X1_508/Y 0.01fF
C21394 PAND2X1_632/B POR2X1_153/Y 0.05fF
C21395 POR2X1_452/Y POR2X1_809/CTRL2 0.01fF
C21396 PAND2X1_206/B PAND2X1_58/A 0.03fF
C21397 POR2X1_394/A POR2X1_744/O 0.02fF
C21398 PAND2X1_835/CTRL POR2X1_77/Y 0.00fF
C21399 PAND2X1_96/B POR2X1_554/O 0.01fF
C21400 POR2X1_110/Y POR2X1_7/A 0.03fF
C21401 PAND2X1_94/A POR2X1_557/B 0.05fF
C21402 POR2X1_146/O POR2X1_146/Y 0.01fF
C21403 POR2X1_305/CTRL2 PAND2X1_651/Y 0.00fF
C21404 POR2X1_664/Y PAND2X1_72/A 0.02fF
C21405 PAND2X1_64/CTRL2 PAND2X1_26/A 0.01fF
C21406 POR2X1_416/B PAND2X1_794/B 0.06fF
C21407 PAND2X1_450/CTRL POR2X1_158/Y 0.00fF
C21408 PAND2X1_450/O POR2X1_416/B 0.17fF
C21409 PAND2X1_621/CTRL2 POR2X1_617/Y 0.01fF
C21410 POR2X1_271/B POR2X1_32/A 0.03fF
C21411 PAND2X1_717/Y POR2X1_7/Y 0.00fF
C21412 PAND2X1_39/B D_INPUT_0 0.33fF
C21413 POR2X1_775/A PAND2X1_72/A 0.05fF
C21414 PAND2X1_39/B POR2X1_811/A 0.01fF
C21415 POR2X1_116/A POR2X1_474/CTRL2 0.00fF
C21416 POR2X1_813/O POR2X1_669/B 0.01fF
C21417 PAND2X1_35/A POR2X1_409/B 0.06fF
C21418 PAND2X1_39/B POR2X1_287/CTRL2 0.01fF
C21419 POR2X1_196/CTRL POR2X1_334/Y 0.08fF
C21420 POR2X1_825/Y POR2X1_7/B 0.00fF
C21421 POR2X1_339/a_16_28# POR2X1_332/Y 0.03fF
C21422 POR2X1_677/Y PAND2X1_785/Y 0.03fF
C21423 POR2X1_568/B POR2X1_148/B 0.02fF
C21424 POR2X1_567/B POR2X1_446/a_76_344# 0.04fF
C21425 POR2X1_169/A POR2X1_704/CTRL 0.02fF
C21426 PAND2X1_60/B POR2X1_342/B 0.03fF
C21427 PAND2X1_48/B POR2X1_635/B 0.01fF
C21428 PAND2X1_72/A POR2X1_112/Y 0.04fF
C21429 POR2X1_169/O POR2X1_169/B 0.00fF
C21430 POR2X1_16/CTRL2 POR2X1_42/Y 0.01fF
C21431 POR2X1_744/Y POR2X1_40/Y 0.01fF
C21432 POR2X1_859/CTRL2 POR2X1_734/A 0.05fF
C21433 POR2X1_48/A POR2X1_484/CTRL2 0.11fF
C21434 PAND2X1_48/A PAND2X1_692/CTRL2 0.01fF
C21435 POR2X1_612/Y POR2X1_414/CTRL2 0.05fF
C21436 POR2X1_545/a_16_28# POR2X1_551/A 0.02fF
C21437 POR2X1_13/A POR2X1_667/O 0.01fF
C21438 PAND2X1_497/CTRL2 PAND2X1_58/A 0.01fF
C21439 PAND2X1_72/A POR2X1_162/Y 0.02fF
C21440 POR2X1_447/B POR2X1_192/B 0.03fF
C21441 POR2X1_343/Y POR2X1_456/B 0.05fF
C21442 POR2X1_567/A POR2X1_97/B 0.02fF
C21443 POR2X1_657/CTRL2 POR2X1_218/Y 0.10fF
C21444 POR2X1_54/Y PAND2X1_395/CTRL 0.05fF
C21445 POR2X1_23/Y PAND2X1_76/CTRL 0.01fF
C21446 POR2X1_754/a_76_344# POR2X1_39/B 0.01fF
C21447 PAND2X1_796/B PAND2X1_778/CTRL2 0.00fF
C21448 POR2X1_814/B POR2X1_240/CTRL 0.03fF
C21449 POR2X1_16/A POR2X1_86/Y 0.00fF
C21450 PAND2X1_39/B PAND2X1_90/Y 0.07fF
C21451 PAND2X1_20/A D_INPUT_0 3.82fF
C21452 POR2X1_67/Y POR2X1_42/Y 0.05fF
C21453 POR2X1_835/B POR2X1_578/Y 0.03fF
C21454 POR2X1_558/B POR2X1_474/a_76_344# 0.03fF
C21455 POR2X1_624/Y POR2X1_573/O 0.01fF
C21456 POR2X1_634/A POR2X1_66/A 10.36fF
C21457 POR2X1_13/A POR2X1_603/O 0.02fF
C21458 POR2X1_16/A POR2X1_43/Y 0.11fF
C21459 PAND2X1_58/CTRL2 POR2X1_202/A 0.05fF
C21460 POR2X1_14/Y POR2X1_422/Y 0.00fF
C21461 PAND2X1_716/B POR2X1_39/B 0.03fF
C21462 POR2X1_655/A POR2X1_480/A 0.03fF
C21463 PAND2X1_279/CTRL2 PAND2X1_58/A 0.01fF
C21464 POR2X1_15/O POR2X1_9/Y 0.02fF
C21465 POR2X1_567/B POR2X1_439/Y 0.05fF
C21466 PAND2X1_39/B PAND2X1_760/O 0.16fF
C21467 PAND2X1_224/O POR2X1_532/A 0.06fF
C21468 POR2X1_106/a_16_28# POR2X1_60/A 0.00fF
C21469 POR2X1_54/Y POR2X1_13/A 0.12fF
C21470 POR2X1_168/m4_208_n4# POR2X1_191/Y 0.03fF
C21471 POR2X1_816/Y VDD 0.00fF
C21472 POR2X1_65/A POR2X1_263/Y 0.03fF
C21473 POR2X1_117/CTRL POR2X1_409/B 0.01fF
C21474 PAND2X1_115/O POR2X1_150/Y 0.09fF
C21475 PAND2X1_431/CTRL2 POR2X1_480/A 0.05fF
C21476 D_INPUT_0 PAND2X1_525/CTRL 0.01fF
C21477 POR2X1_814/B D_INPUT_0 0.08fF
C21478 PAND2X1_220/Y PAND2X1_352/A 0.01fF
C21479 PAND2X1_212/B POR2X1_40/Y 0.09fF
C21480 POR2X1_49/Y PAND2X1_623/CTRL 0.00fF
C21481 POR2X1_556/A PAND2X1_55/Y 0.07fF
C21482 POR2X1_814/A POR2X1_784/CTRL 0.01fF
C21483 POR2X1_69/m4_208_n4# POR2X1_29/A 0.15fF
C21484 POR2X1_119/O POR2X1_411/B 0.01fF
C21485 PAND2X1_811/A PAND2X1_805/A 0.12fF
C21486 POR2X1_634/A POR2X1_634/CTRL2 0.01fF
C21487 POR2X1_266/A PAND2X1_52/B 0.03fF
C21488 POR2X1_139/Y PAND2X1_39/B 0.01fF
C21489 PAND2X1_287/Y PAND2X1_580/B 0.03fF
C21490 PAND2X1_68/CTRL POR2X1_5/Y 0.03fF
C21491 POR2X1_66/B POR2X1_650/a_16_28# 0.03fF
C21492 PAND2X1_219/A PAND2X1_733/A 0.00fF
C21493 POR2X1_220/Y POR2X1_222/O 0.01fF
C21494 POR2X1_420/Y POR2X1_419/Y 0.01fF
C21495 POR2X1_115/O POR2X1_76/A 0.01fF
C21496 POR2X1_353/Y POR2X1_97/A 0.15fF
C21497 PAND2X1_58/A POR2X1_750/B 0.07fF
C21498 POR2X1_294/Y PAND2X1_58/CTRL 0.01fF
C21499 PAND2X1_717/A POR2X1_91/Y 0.03fF
C21500 POR2X1_37/Y POR2X1_497/Y 0.02fF
C21501 PAND2X1_299/O POR2X1_121/B 0.18fF
C21502 POR2X1_105/Y POR2X1_590/A 4.61fF
C21503 POR2X1_19/CTRL D_INPUT_1 0.01fF
C21504 PAND2X1_475/CTRL PAND2X1_217/B 0.29fF
C21505 PAND2X1_832/m4_208_n4# PAND2X1_436/m4_208_n4# 0.13fF
C21506 POR2X1_407/A PAND2X1_761/CTRL2 0.01fF
C21507 PAND2X1_57/B PAND2X1_248/a_16_344# 0.02fF
C21508 PAND2X1_695/CTRL2 PAND2X1_11/Y 0.02fF
C21509 POR2X1_130/A POR2X1_66/A 0.10fF
C21510 POR2X1_567/B POR2X1_192/Y 0.13fF
C21511 PAND2X1_651/Y POR2X1_271/B 0.05fF
C21512 POR2X1_63/Y POR2X1_406/A 0.05fF
C21513 POR2X1_717/B POR2X1_188/Y 0.03fF
C21514 POR2X1_590/A POR2X1_733/O 0.01fF
C21515 PAND2X1_52/B POR2X1_691/A 0.00fF
C21516 POR2X1_805/Y PAND2X1_90/Y 0.04fF
C21517 POR2X1_357/B POR2X1_568/A 0.01fF
C21518 POR2X1_66/Y PAND2X1_625/O 0.08fF
C21519 POR2X1_260/B PAND2X1_385/CTRL 0.09fF
C21520 POR2X1_566/A POR2X1_66/A 0.20fF
C21521 POR2X1_83/B POR2X1_697/CTRL2 0.03fF
C21522 PAND2X1_20/A PAND2X1_90/Y 0.10fF
C21523 POR2X1_423/Y PAND2X1_541/CTRL 0.01fF
C21524 POR2X1_428/Y POR2X1_426/O 0.01fF
C21525 PAND2X1_423/O POR2X1_330/Y 0.02fF
C21526 PAND2X1_673/O POR2X1_14/Y 0.08fF
C21527 D_INPUT_0 POR2X1_513/B 0.17fF
C21528 PAND2X1_459/O POR2X1_376/Y 0.08fF
C21529 POR2X1_201/a_76_344# PAND2X1_65/Y 0.01fF
C21530 POR2X1_259/A PAND2X1_52/Y 0.01fF
C21531 POR2X1_677/Y POR2X1_300/Y 0.00fF
C21532 PAND2X1_803/A POR2X1_72/B 0.03fF
C21533 POR2X1_667/A VDD 0.22fF
C21534 POR2X1_355/B PAND2X1_73/Y 0.03fF
C21535 POR2X1_20/B PAND2X1_388/Y 0.03fF
C21536 POR2X1_366/Y POR2X1_466/A 0.10fF
C21537 POR2X1_343/A POR2X1_287/B 0.07fF
C21538 PAND2X1_9/Y POR2X1_278/A 0.23fF
C21539 PAND2X1_55/Y PAND2X1_591/O 0.01fF
C21540 POR2X1_596/A POR2X1_678/a_16_28# 0.01fF
C21541 POR2X1_810/CTRL2 POR2X1_636/B 0.01fF
C21542 POR2X1_293/CTRL POR2X1_5/Y 0.01fF
C21543 PAND2X1_849/O PAND2X1_61/Y 0.02fF
C21544 PAND2X1_471/O POR2X1_14/Y 0.17fF
C21545 POR2X1_234/Y POR2X1_102/Y 0.01fF
C21546 POR2X1_314/a_16_28# POR2X1_48/A 0.01fF
C21547 POR2X1_20/B PAND2X1_549/B 0.03fF
C21548 POR2X1_376/B PAND2X1_333/O 0.09fF
C21549 POR2X1_814/B PAND2X1_90/Y 2.67fF
C21550 POR2X1_857/B POR2X1_241/B 0.03fF
C21551 PAND2X1_20/A POR2X1_401/a_16_28# 0.03fF
C21552 POR2X1_41/B POR2X1_142/CTRL 0.05fF
C21553 POR2X1_337/A POR2X1_556/A 0.07fF
C21554 POR2X1_66/A POR2X1_204/CTRL 0.01fF
C21555 POR2X1_13/A PAND2X1_784/A 0.01fF
C21556 POR2X1_43/B POR2X1_409/B 0.03fF
C21557 POR2X1_601/Y VDD 0.01fF
C21558 PAND2X1_65/B PAND2X1_65/Y 0.01fF
C21559 POR2X1_63/Y PAND2X1_63/B 0.04fF
C21560 POR2X1_254/Y POR2X1_330/Y 0.07fF
C21561 PAND2X1_845/CTRL2 POR2X1_37/Y 0.01fF
C21562 POR2X1_635/Y POR2X1_750/B 0.01fF
C21563 POR2X1_118/CTRL2 POR2X1_37/Y 0.12fF
C21564 POR2X1_410/Y POR2X1_260/B 0.01fF
C21565 POR2X1_427/Y POR2X1_236/Y 0.01fF
C21566 POR2X1_435/Y POR2X1_750/B 0.07fF
C21567 POR2X1_390/B POR2X1_499/A 0.03fF
C21568 POR2X1_614/A POR2X1_614/a_16_28# -0.00fF
C21569 POR2X1_139/Y PAND2X1_20/A 0.01fF
C21570 PAND2X1_465/B POR2X1_14/Y 0.34fF
C21571 PAND2X1_859/A INPUT_0 0.31fF
C21572 PAND2X1_546/Y POR2X1_32/A 0.00fF
C21573 POR2X1_66/A POR2X1_844/B 0.03fF
C21574 POR2X1_60/A POR2X1_494/Y 0.03fF
C21575 POR2X1_653/B VDD 0.04fF
C21576 PAND2X1_787/O PAND2X1_556/B 0.00fF
C21577 POR2X1_855/B POR2X1_803/a_56_344# 0.00fF
C21578 POR2X1_48/A PAND2X1_324/a_16_344# 0.05fF
C21579 PAND2X1_193/Y POR2X1_761/A 0.03fF
C21580 PAND2X1_590/O POR2X1_38/Y 0.03fF
C21581 PAND2X1_795/a_56_28# INPUT_0 0.00fF
C21582 PAND2X1_282/CTRL2 PAND2X1_69/A 0.03fF
C21583 POR2X1_655/A PAND2X1_305/O 0.15fF
C21584 POR2X1_830/A VDD 0.38fF
C21585 PAND2X1_717/A POR2X1_109/Y 0.01fF
C21586 POR2X1_58/O POR2X1_236/Y 0.03fF
C21587 POR2X1_260/B POR2X1_702/O 0.04fF
C21588 POR2X1_409/B POR2X1_38/B 0.06fF
C21589 PAND2X1_32/O POR2X1_294/A 0.17fF
C21590 PAND2X1_712/B VDD 0.17fF
C21591 PAND2X1_229/CTRL2 POR2X1_579/Y 0.00fF
C21592 PAND2X1_479/B PAND2X1_479/O 0.00fF
C21593 POR2X1_276/A POR2X1_260/B 0.02fF
C21594 POR2X1_150/Y PAND2X1_182/B 0.01fF
C21595 POR2X1_102/Y POR2X1_183/Y 0.03fF
C21596 PAND2X1_771/Y PAND2X1_568/B 0.05fF
C21597 PAND2X1_4/CTRL D_INPUT_0 0.00fF
C21598 POR2X1_624/Y POR2X1_456/B 0.04fF
C21599 PAND2X1_55/Y POR2X1_202/O 0.01fF
C21600 POR2X1_376/B PAND2X1_99/CTRL 0.03fF
C21601 POR2X1_87/Y VDD 0.12fF
C21602 POR2X1_179/a_76_344# POR2X1_102/Y 0.01fF
C21603 PAND2X1_41/B POR2X1_717/Y 0.03fF
C21604 PAND2X1_467/B POR2X1_694/CTRL 0.01fF
C21605 POR2X1_378/O POR2X1_55/Y 0.17fF
C21606 POR2X1_390/B POR2X1_76/A 0.03fF
C21607 POR2X1_46/Y PAND2X1_332/O 0.18fF
C21608 POR2X1_65/A PAND2X1_215/B 0.06fF
C21609 POR2X1_177/Y PAND2X1_182/A 0.00fF
C21610 POR2X1_78/B POR2X1_192/Y 0.10fF
C21611 POR2X1_808/A POR2X1_800/A 0.08fF
C21612 POR2X1_57/A POR2X1_669/B 0.23fF
C21613 POR2X1_487/Y PAND2X1_794/B 0.01fF
C21614 PAND2X1_90/Y POR2X1_513/B 0.19fF
C21615 POR2X1_96/A POR2X1_230/a_16_28# 0.03fF
C21616 POR2X1_693/Y PAND2X1_706/O 0.00fF
C21617 POR2X1_376/Y PAND2X1_375/CTRL 0.01fF
C21618 POR2X1_3/A POR2X1_32/A 0.06fF
C21619 POR2X1_407/A POR2X1_783/O 0.01fF
C21620 PAND2X1_558/Y POR2X1_599/A 0.12fF
C21621 POR2X1_763/A POR2X1_700/CTRL 0.05fF
C21622 POR2X1_94/O POR2X1_94/A 0.06fF
C21623 PAND2X1_283/CTRL2 POR2X1_734/A 0.02fF
C21624 POR2X1_389/O POR2X1_814/B 0.06fF
C21625 POR2X1_502/A POR2X1_794/O 0.01fF
C21626 POR2X1_782/A POR2X1_750/B 0.06fF
C21627 POR2X1_290/a_16_28# POR2X1_290/Y 0.02fF
C21628 POR2X1_188/A PAND2X1_536/a_16_344# 0.01fF
C21629 PAND2X1_805/O POR2X1_7/B 0.01fF
C21630 PAND2X1_626/O PAND2X1_96/B 0.04fF
C21631 POR2X1_608/Y PAND2X1_60/B 0.04fF
C21632 POR2X1_719/CTRL2 POR2X1_121/B 0.08fF
C21633 POR2X1_96/A INPUT_0 0.10fF
C21634 POR2X1_537/Y POR2X1_841/CTRL2 0.01fF
C21635 PAND2X1_422/CTRL POR2X1_296/B 0.06fF
C21636 POR2X1_809/A PAND2X1_761/CTRL 0.01fF
C21637 POR2X1_497/Y POR2X1_293/Y 0.07fF
C21638 POR2X1_186/Y POR2X1_731/CTRL2 0.16fF
C21639 POR2X1_448/A POR2X1_294/B 0.09fF
C21640 POR2X1_78/B PAND2X1_322/a_56_28# 0.00fF
C21641 POR2X1_254/A PAND2X1_96/B 0.03fF
C21642 PAND2X1_213/Y POR2X1_83/B 0.06fF
C21643 POR2X1_634/A POR2X1_532/A 0.27fF
C21644 POR2X1_478/Y POR2X1_319/Y 0.01fF
C21645 PAND2X1_620/Y PAND2X1_6/A 0.07fF
C21646 POR2X1_130/O POR2X1_260/B 0.01fF
C21647 POR2X1_566/A PAND2X1_524/CTRL 0.05fF
C21648 POR2X1_20/B POR2X1_397/CTRL 0.01fF
C21649 POR2X1_208/A POR2X1_590/A 0.00fF
C21650 POR2X1_73/O D_INPUT_0 0.02fF
C21651 PAND2X1_169/Y POR2X1_73/Y 0.01fF
C21652 POR2X1_49/Y PAND2X1_470/CTRL2 0.01fF
C21653 POR2X1_65/A PAND2X1_6/A 0.26fF
C21654 PAND2X1_64/O POR2X1_260/A 0.02fF
C21655 POR2X1_483/A POR2X1_795/a_76_344# 0.02fF
C21656 PAND2X1_244/CTRL2 PAND2X1_175/B 0.01fF
C21657 POR2X1_251/m4_208_n4# PAND2X1_190/Y 0.10fF
C21658 PAND2X1_96/B POR2X1_750/B 0.38fF
C21659 POR2X1_110/Y PAND2X1_466/B 0.03fF
C21660 PAND2X1_641/O POR2X1_263/Y 0.02fF
C21661 POR2X1_653/a_16_28# POR2X1_661/B 0.03fF
C21662 POR2X1_284/B POR2X1_740/Y 0.05fF
C21663 POR2X1_294/Y POR2X1_260/A 0.04fF
C21664 POR2X1_774/Y PAND2X1_583/O 0.08fF
C21665 PAND2X1_852/CTRL VDD 0.00fF
C21666 PAND2X1_512/CTRL POR2X1_239/Y 0.01fF
C21667 PAND2X1_297/CTRL POR2X1_296/B 0.01fF
C21668 POR2X1_336/CTRL POR2X1_814/B 0.00fF
C21669 PAND2X1_76/m4_208_n4# POR2X1_91/Y 0.12fF
C21670 POR2X1_285/a_16_28# POR2X1_285/A 0.05fF
C21671 POR2X1_13/A POR2X1_13/Y 0.02fF
C21672 POR2X1_99/A PAND2X1_60/B 0.03fF
C21673 POR2X1_640/A PAND2X1_32/B 0.00fF
C21674 POR2X1_108/CTRL PAND2X1_562/B 0.05fF
C21675 VDD PAND2X1_146/O 0.00fF
C21676 POR2X1_465/B POR2X1_193/A 0.03fF
C21677 PAND2X1_55/Y POR2X1_445/CTRL 0.11fF
C21678 POR2X1_313/a_16_28# POR2X1_72/B 0.01fF
C21679 POR2X1_251/Y POR2X1_42/Y 0.05fF
C21680 PAND2X1_52/Y PAND2X1_88/Y 0.51fF
C21681 PAND2X1_90/A PAND2X1_92/O 0.01fF
C21682 POR2X1_66/B POR2X1_569/A 0.07fF
C21683 PAND2X1_48/B POR2X1_360/A 0.07fF
C21684 POR2X1_495/CTRL2 POR2X1_283/A 0.01fF
C21685 PAND2X1_641/Y POR2X1_32/A 0.07fF
C21686 PAND2X1_347/Y PAND2X1_578/A 0.00fF
C21687 PAND2X1_738/Y PAND2X1_794/B 0.05fF
C21688 POR2X1_186/Y POR2X1_510/Y 0.03fF
C21689 POR2X1_348/CTRL2 POR2X1_814/B 0.01fF
C21690 POR2X1_814/B POR2X1_361/O 0.28fF
C21691 PAND2X1_465/B POR2X1_55/Y 0.01fF
C21692 PAND2X1_478/O POR2X1_46/Y 0.04fF
C21693 POR2X1_355/B POR2X1_509/A 0.15fF
C21694 PAND2X1_823/O POR2X1_836/A 0.02fF
C21695 PAND2X1_231/CTRL POR2X1_229/Y 0.01fF
C21696 POR2X1_43/B PAND2X1_351/Y 0.05fF
C21697 POR2X1_826/CTRL PAND2X1_338/B 0.00fF
C21698 POR2X1_347/B POR2X1_68/A 0.00fF
C21699 POR2X1_52/A PAND2X1_652/A 0.05fF
C21700 PAND2X1_673/CTRL D_INPUT_3 0.12fF
C21701 POR2X1_549/CTRL2 POR2X1_383/A 0.03fF
C21702 POR2X1_383/A PAND2X1_299/O 0.04fF
C21703 POR2X1_710/A POR2X1_713/B 0.00fF
C21704 POR2X1_48/A PAND2X1_716/B 0.03fF
C21705 PAND2X1_242/O POR2X1_7/B 0.15fF
C21706 POR2X1_225/CTRL POR2X1_129/Y 0.01fF
C21707 PAND2X1_41/B POR2X1_218/CTRL 0.01fF
C21708 PAND2X1_620/Y POR2X1_588/Y 0.04fF
C21709 POR2X1_416/Y POR2X1_232/CTRL 0.01fF
C21710 PAND2X1_340/O POR2X1_408/Y 0.10fF
C21711 POR2X1_327/Y POR2X1_296/B 0.69fF
C21712 PAND2X1_845/O PAND2X1_35/Y 0.02fF
C21713 POR2X1_579/Y D_GATE_741 0.22fF
C21714 PAND2X1_830/CTRL PAND2X1_562/B 0.04fF
C21715 POR2X1_596/A VDD 0.01fF
C21716 POR2X1_529/Y POR2X1_5/Y 0.02fF
C21717 POR2X1_188/A PAND2X1_698/CTRL 0.01fF
C21718 POR2X1_130/A POR2X1_532/A 0.07fF
C21719 POR2X1_656/O POR2X1_737/A 0.01fF
C21720 PAND2X1_41/B PAND2X1_503/CTRL2 0.01fF
C21721 POR2X1_862/CTRL2 POR2X1_647/B 0.01fF
C21722 POR2X1_49/Y POR2X1_419/CTRL 0.07fF
C21723 PAND2X1_472/A POR2X1_7/B 0.01fF
C21724 PAND2X1_244/CTRL POR2X1_153/Y 0.07fF
C21725 POR2X1_445/O POR2X1_702/A 0.00fF
C21726 POR2X1_149/B POR2X1_294/B 0.03fF
C21727 POR2X1_566/A POR2X1_532/A 0.05fF
C21728 PAND2X1_661/B POR2X1_277/CTRL2 0.03fF
C21729 PAND2X1_200/Y POR2X1_153/Y 0.04fF
C21730 POR2X1_795/CTRL2 POR2X1_786/Y 0.03fF
C21731 PAND2X1_477/B PAND2X1_241/CTRL 0.01fF
C21732 POR2X1_559/Y POR2X1_294/B 0.06fF
C21733 POR2X1_654/B POR2X1_773/B 0.32fF
C21734 PAND2X1_137/CTRL POR2X1_134/Y 0.01fF
C21735 POR2X1_311/Y PAND2X1_360/Y 0.03fF
C21736 POR2X1_563/CTRL POR2X1_569/A 0.05fF
C21737 POR2X1_25/Y POR2X1_32/A 0.04fF
C21738 POR2X1_85/CTRL2 POR2X1_23/Y 0.01fF
C21739 POR2X1_548/O PAND2X1_63/B 0.02fF
C21740 POR2X1_176/CTRL POR2X1_83/B 0.01fF
C21741 POR2X1_68/A PAND2X1_604/a_16_344# 0.02fF
C21742 POR2X1_32/A POR2X1_701/CTRL 0.01fF
C21743 POR2X1_541/B PAND2X1_72/A 0.03fF
C21744 PAND2X1_69/A POR2X1_208/O 0.09fF
C21745 POR2X1_13/A PAND2X1_787/A 0.03fF
C21746 POR2X1_362/B POR2X1_101/Y 0.05fF
C21747 INPUT_1 PAND2X1_721/CTRL2 0.11fF
C21748 POR2X1_245/Y VDD 0.14fF
C21749 POR2X1_41/B POR2X1_93/A 0.07fF
C21750 PAND2X1_821/O POR2X1_510/A 0.00fF
C21751 POR2X1_219/CTRL POR2X1_294/B 0.03fF
C21752 PAND2X1_139/B PAND2X1_349/A 0.00fF
C21753 PAND2X1_599/CTRL POR2X1_828/A 0.02fF
C21754 INPUT_0 POR2X1_7/A 1.00fF
C21755 POR2X1_750/A POR2X1_749/O 0.02fF
C21756 POR2X1_41/B POR2X1_91/Y 0.10fF
C21757 POR2X1_649/CTRL POR2X1_294/B 0.00fF
C21758 POR2X1_52/A POR2X1_152/Y 0.27fF
C21759 POR2X1_416/B POR2X1_672/Y 0.05fF
C21760 POR2X1_278/Y PAND2X1_656/A 0.05fF
C21761 POR2X1_389/A PAND2X1_385/CTRL2 0.00fF
C21762 PAND2X1_318/CTRL POR2X1_91/Y 0.09fF
C21763 POR2X1_207/B PAND2X1_55/Y 0.03fF
C21764 POR2X1_416/B POR2X1_699/CTRL2 0.01fF
C21765 POR2X1_423/Y POR2X1_129/Y 0.01fF
C21766 POR2X1_13/Y PAND2X1_643/Y 0.01fF
C21767 POR2X1_56/B PAND2X1_241/Y 0.03fF
C21768 PAND2X1_228/O PAND2X1_341/A 0.05fF
C21769 POR2X1_708/B PAND2X1_60/B 0.01fF
C21770 PAND2X1_341/B POR2X1_60/A 0.03fF
C21771 POR2X1_591/CTRL2 POR2X1_591/Y 0.01fF
C21772 PAND2X1_462/CTRL2 POR2X1_48/A 0.03fF
C21773 POR2X1_380/Y POR2X1_7/B 0.03fF
C21774 POR2X1_68/B PAND2X1_110/a_16_344# 0.01fF
C21775 POR2X1_462/B POR2X1_790/A 0.07fF
C21776 POR2X1_829/A PAND2X1_656/A 0.01fF
C21777 POR2X1_118/Y POR2X1_77/Y 0.85fF
C21778 PAND2X1_652/A PAND2X1_186/O 0.27fF
C21779 POR2X1_416/B PAND2X1_124/Y 0.07fF
C21780 PAND2X1_6/Y POR2X1_786/Y 0.21fF
C21781 POR2X1_790/A D_INPUT_1 0.02fF
C21782 POR2X1_483/A POR2X1_833/A 0.01fF
C21783 PAND2X1_715/O POR2X1_310/Y 0.02fF
C21784 PAND2X1_592/Y PAND2X1_843/Y 0.02fF
C21785 PAND2X1_726/CTRL POR2X1_152/Y 0.01fF
C21786 PAND2X1_850/Y POR2X1_102/Y 0.07fF
C21787 POR2X1_717/a_16_28# POR2X1_717/Y 0.03fF
C21788 VDD POR2X1_703/Y 0.17fF
C21789 PAND2X1_579/A VDD 0.00fF
C21790 PAND2X1_551/CTRL2 PAND2X1_324/Y 0.00fF
C21791 PAND2X1_6/Y POR2X1_788/B 0.06fF
C21792 POR2X1_614/A POR2X1_685/B 0.01fF
C21793 POR2X1_532/A POR2X1_844/B 0.03fF
C21794 POR2X1_131/Y PAND2X1_137/Y 0.20fF
C21795 POR2X1_68/A POR2X1_318/A 0.10fF
C21796 PAND2X1_126/O PAND2X1_90/A 0.03fF
C21797 PAND2X1_84/Y POR2X1_394/A 0.29fF
C21798 POR2X1_100/CTRL PAND2X1_69/A 0.00fF
C21799 PAND2X1_812/O PAND2X1_568/B 0.02fF
C21800 POR2X1_725/Y POR2X1_777/O 0.04fF
C21801 PAND2X1_270/O POR2X1_184/Y 0.01fF
C21802 POR2X1_618/a_16_28# POR2X1_7/A 0.02fF
C21803 POR2X1_293/Y POR2X1_310/Y 0.01fF
C21804 POR2X1_596/A PAND2X1_32/B 0.03fF
C21805 POR2X1_65/A POR2X1_119/Y 0.08fF
C21806 PAND2X1_498/CTRL2 POR2X1_260/A 0.00fF
C21807 PAND2X1_641/Y PAND2X1_35/Y 0.02fF
C21808 D_GATE_662 PAND2X1_373/CTRL2 0.08fF
C21809 POR2X1_110/Y POR2X1_485/CTRL2 0.00fF
C21810 POR2X1_224/O POR2X1_394/A 0.12fF
C21811 PAND2X1_6/Y PAND2X1_27/CTRL2 0.01fF
C21812 POR2X1_404/m4_208_n4# PAND2X1_399/m4_208_n4# 0.05fF
C21813 POR2X1_60/A POR2X1_533/Y 0.20fF
C21814 POR2X1_254/Y POR2X1_715/A 0.01fF
C21815 POR2X1_532/A POR2X1_573/A 0.05fF
C21816 POR2X1_383/A PAND2X1_519/O 0.03fF
C21817 POR2X1_94/A PAND2X1_379/CTRL 0.00fF
C21818 PAND2X1_651/Y PAND2X1_270/O 0.12fF
C21819 POR2X1_717/CTRL POR2X1_865/B 0.00fF
C21820 POR2X1_416/B POR2X1_83/B 0.52fF
C21821 POR2X1_438/a_56_344# POR2X1_142/Y 0.00fF
C21822 PAND2X1_824/B POR2X1_208/O 0.03fF
C21823 PAND2X1_308/Y PAND2X1_303/CTRL 0.01fF
C21824 POR2X1_346/B PAND2X1_625/CTRL2 0.00fF
C21825 POR2X1_192/Y POR2X1_180/O 0.06fF
C21826 PAND2X1_351/CTRL POR2X1_153/Y 0.30fF
C21827 PAND2X1_772/a_16_344# POR2X1_77/Y 0.01fF
C21828 POR2X1_96/A PAND2X1_355/CTRL 0.01fF
C21829 PAND2X1_511/O PAND2X1_48/A 0.07fF
C21830 POR2X1_856/B POR2X1_863/A 16.63fF
C21831 PAND2X1_548/a_76_28# POR2X1_530/Y 0.04fF
C21832 PAND2X1_550/B PAND2X1_565/A 0.04fF
C21833 POR2X1_83/A INPUT_1 0.22fF
C21834 PAND2X1_29/CTRL2 POR2X1_260/A 0.03fF
C21835 POR2X1_416/B POR2X1_626/Y 0.00fF
C21836 POR2X1_333/A PAND2X1_52/B 0.05fF
C21837 POR2X1_165/a_16_28# POR2X1_73/Y 0.05fF
C21838 POR2X1_333/A POR2X1_212/B 0.17fF
C21839 PAND2X1_358/A PAND2X1_341/O 0.07fF
C21840 PAND2X1_341/A PAND2X1_100/CTRL2 0.01fF
C21841 POR2X1_565/B POR2X1_6/a_16_28# 0.09fF
C21842 POR2X1_593/B PAND2X1_56/A 0.01fF
C21843 PAND2X1_25/m4_208_n4# PAND2X1_72/A 0.12fF
C21844 POR2X1_404/Y PAND2X1_48/A 0.01fF
C21845 POR2X1_66/B PAND2X1_72/A 0.13fF
C21846 POR2X1_785/CTRL POR2X1_191/Y 0.24fF
C21847 POR2X1_63/Y POR2X1_262/a_16_28# 0.03fF
C21848 POR2X1_13/A POR2X1_4/Y 0.03fF
C21849 POR2X1_562/CTRL POR2X1_339/Y 0.01fF
C21850 POR2X1_96/CTRL2 POR2X1_38/B 0.01fF
C21851 INPUT_1 POR2X1_90/Y 0.51fF
C21852 POR2X1_83/A POR2X1_153/Y 0.19fF
C21853 PAND2X1_38/O POR2X1_4/Y 0.16fF
C21854 POR2X1_220/Y POR2X1_330/CTRL2 0.00fF
C21855 POR2X1_68/A POR2X1_574/Y 0.05fF
C21856 POR2X1_16/A POR2X1_73/Y 5.52fF
C21857 POR2X1_733/A POR2X1_737/A 0.05fF
C21858 PAND2X1_90/A PAND2X1_527/O 0.01fF
C21859 POR2X1_52/A PAND2X1_506/Y 0.01fF
C21860 POR2X1_712/CTRL POR2X1_707/Y 0.01fF
C21861 POR2X1_49/Y PAND2X1_847/O 0.17fF
C21862 POR2X1_734/A PAND2X1_52/B 0.07fF
C21863 PAND2X1_149/CTRL PAND2X1_797/Y 0.04fF
C21864 PAND2X1_716/B PAND2X1_197/Y 0.00fF
C21865 POR2X1_265/Y POR2X1_406/a_16_28# 0.07fF
C21866 POR2X1_327/Y POR2X1_267/Y 0.00fF
C21867 PAND2X1_834/O POR2X1_236/Y 0.06fF
C21868 PAND2X1_48/B POR2X1_99/B 0.03fF
C21869 POR2X1_90/Y POR2X1_153/Y 0.03fF
C21870 GATE_662 POR2X1_413/A 0.01fF
C21871 PAND2X1_802/a_16_344# POR2X1_42/Y 0.02fF
C21872 PAND2X1_172/CTRL2 POR2X1_854/B 0.02fF
C21873 POR2X1_763/Y POR2X1_320/a_16_28# 0.09fF
C21874 POR2X1_862/CTRL POR2X1_130/A 0.29fF
C21875 POR2X1_203/O PAND2X1_72/Y 0.02fF
C21876 POR2X1_860/CTRL POR2X1_383/A 0.00fF
C21877 PAND2X1_308/Y POR2X1_91/Y 0.07fF
C21878 POR2X1_390/B POR2X1_539/A 0.02fF
C21879 PAND2X1_72/Y PAND2X1_111/B 0.60fF
C21880 INPUT_1 POR2X1_383/A 0.06fF
C21881 PAND2X1_59/CTRL2 PAND2X1_18/B 0.01fF
C21882 POR2X1_119/Y PAND2X1_836/CTRL2 0.01fF
C21883 POR2X1_343/Y PAND2X1_57/B 0.00fF
C21884 POR2X1_132/Y POR2X1_132/O 0.01fF
C21885 POR2X1_394/A PAND2X1_149/A 0.03fF
C21886 POR2X1_347/CTRL2 POR2X1_402/A 0.01fF
C21887 POR2X1_349/CTRL2 POR2X1_532/A 0.01fF
C21888 POR2X1_325/CTRL2 POR2X1_544/B 0.01fF
C21889 PAND2X1_612/B PAND2X1_612/a_76_28# 0.01fF
C21890 PAND2X1_173/O POR2X1_186/B -0.00fF
C21891 PAND2X1_243/B POR2X1_39/B 0.03fF
C21892 POR2X1_858/A POR2X1_733/A 0.20fF
C21893 POR2X1_614/A POR2X1_560/O 0.03fF
C21894 POR2X1_732/B POR2X1_181/a_56_344# 0.03fF
C21895 POR2X1_96/B POR2X1_394/A 0.03fF
C21896 D_GATE_662 POR2X1_568/B 0.10fF
C21897 POR2X1_333/Y POR2X1_566/B 0.03fF
C21898 POR2X1_16/A PAND2X1_727/O 0.04fF
C21899 POR2X1_38/B POR2X1_560/O 0.10fF
C21900 POR2X1_110/CTRL2 POR2X1_7/A 0.03fF
C21901 POR2X1_411/B PAND2X1_205/A 0.03fF
C21902 PAND2X1_96/B PAND2X1_122/CTRL 0.00fF
C21903 PAND2X1_192/Y PAND2X1_221/Y 0.01fF
C21904 POR2X1_659/CTRL POR2X1_736/A 0.11fF
C21905 POR2X1_416/B PAND2X1_709/O 0.04fF
C21906 POR2X1_190/Y POR2X1_568/A 0.03fF
C21907 POR2X1_567/A POR2X1_540/a_76_344# 0.01fF
C21908 POR2X1_713/CTRL POR2X1_711/Y 0.01fF
C21909 PAND2X1_724/O PAND2X1_326/B 0.02fF
C21910 POR2X1_456/B POR2X1_186/B 0.06fF
C21911 PAND2X1_221/a_16_344# POR2X1_250/Y 0.02fF
C21912 POR2X1_721/O POR2X1_559/A 0.08fF
C21913 POR2X1_102/Y POR2X1_412/CTRL2 0.00fF
C21914 PAND2X1_865/Y PAND2X1_175/B 0.04fF
C21915 POR2X1_181/B POR2X1_540/Y 0.10fF
C21916 PAND2X1_32/O POR2X1_94/A 0.04fF
C21917 POR2X1_678/Y POR2X1_808/CTRL 0.00fF
C21918 POR2X1_63/Y POR2X1_32/A 3.29fF
C21919 PAND2X1_587/CTRL2 PAND2X1_52/B 0.21fF
C21920 PAND2X1_51/O PAND2X1_3/B 0.04fF
C21921 PAND2X1_510/a_56_28# PAND2X1_508/Y 0.00fF
C21922 POR2X1_824/CTRL POR2X1_16/A 0.00fF
C21923 POR2X1_768/CTRL POR2X1_113/B 0.01fF
C21924 POR2X1_814/A PAND2X1_65/Y 0.07fF
C21925 POR2X1_829/A PAND2X1_193/Y 0.03fF
C21926 POR2X1_54/Y POR2X1_29/A 0.11fF
C21927 POR2X1_93/A POR2X1_77/Y 0.04fF
C21928 POR2X1_816/A PAND2X1_332/Y 0.03fF
C21929 POR2X1_77/Y POR2X1_91/Y 1.26fF
C21930 PAND2X1_549/B POR2X1_372/CTRL2 0.11fF
C21931 PAND2X1_508/a_16_344# PAND2X1_506/Y 0.02fF
C21932 POR2X1_711/Y PAND2X1_305/CTRL2 0.01fF
C21933 POR2X1_158/Y POR2X1_526/Y 0.00fF
C21934 PAND2X1_857/A POR2X1_39/B 0.03fF
C21935 PAND2X1_629/CTRL2 POR2X1_20/B 0.03fF
C21936 POR2X1_804/A PAND2X1_135/O 0.00fF
C21937 POR2X1_528/Y POR2X1_305/O 0.03fF
C21938 PAND2X1_58/A POR2X1_606/CTRL2 0.01fF
C21939 POR2X1_711/Y POR2X1_513/a_16_28# 0.06fF
C21940 PAND2X1_39/B POR2X1_780/CTRL2 0.01fF
C21941 POR2X1_78/B POR2X1_646/B -0.00fF
C21942 PAND2X1_374/O POR2X1_39/B 0.04fF
C21943 POR2X1_260/B POR2X1_267/CTRL 0.01fF
C21944 POR2X1_860/A POR2X1_556/A 0.03fF
C21945 PAND2X1_406/O POR2X1_121/B 0.17fF
C21946 PAND2X1_108/a_16_344# POR2X1_814/A 0.04fF
C21947 PAND2X1_163/CTRL PAND2X1_52/B 0.01fF
C21948 PAND2X1_94/Y PAND2X1_55/Y 0.05fF
C21949 POR2X1_676/CTRL2 POR2X1_750/B 0.01fF
C21950 POR2X1_16/A PAND2X1_207/A 0.01fF
C21951 POR2X1_39/B POR2X1_260/A 0.06fF
C21952 POR2X1_318/A POR2X1_138/A 0.04fF
C21953 POR2X1_841/B POR2X1_806/CTRL 0.00fF
C21954 POR2X1_760/A INPUT_0 1.07fF
C21955 POR2X1_459/Y VDD 0.14fF
C21956 PAND2X1_457/Y POR2X1_417/Y 0.24fF
C21957 PAND2X1_76/Y POR2X1_411/B 0.03fF
C21958 POR2X1_241/B POR2X1_66/A 0.03fF
C21959 PAND2X1_63/a_56_28# POR2X1_296/B 0.00fF
C21960 POR2X1_57/A POR2X1_234/A 0.03fF
C21961 PAND2X1_859/A PAND2X1_340/B 0.01fF
C21962 PAND2X1_94/Y POR2X1_402/A 0.02fF
C21963 POR2X1_102/Y PAND2X1_722/CTRL 0.08fF
C21964 POR2X1_719/A POR2X1_66/A 0.07fF
C21965 PAND2X1_313/CTRL PAND2X1_72/A 0.01fF
C21966 POR2X1_647/B POR2X1_480/A 0.02fF
C21967 POR2X1_624/Y PAND2X1_131/CTRL2 0.09fF
C21968 PAND2X1_340/B POR2X1_381/a_56_344# 0.00fF
C21969 POR2X1_760/A PAND2X1_218/CTRL 0.03fF
C21970 PAND2X1_472/A PAND2X1_608/CTRL2 0.06fF
C21971 PAND2X1_217/B D_INPUT_0 0.17fF
C21972 POR2X1_423/Y POR2X1_37/Y 0.03fF
C21973 POR2X1_63/Y PAND2X1_35/Y 0.16fF
C21974 POR2X1_471/A POR2X1_724/O 0.01fF
C21975 POR2X1_23/Y POR2X1_238/CTRL2 0.03fF
C21976 GATE_222 PAND2X1_568/B 0.03fF
C21977 POR2X1_483/m4_208_n4# POR2X1_556/A 0.09fF
C21978 POR2X1_77/Y POR2X1_109/Y 0.03fF
C21979 PAND2X1_57/B POR2X1_624/Y 0.07fF
C21980 POR2X1_792/CTRL2 PAND2X1_41/B 0.02fF
C21981 POR2X1_857/A POR2X1_785/A 0.01fF
C21982 PAND2X1_805/a_16_344# PAND2X1_287/Y 0.02fF
C21983 POR2X1_866/A PAND2X1_511/CTRL2 0.06fF
C21984 PAND2X1_473/O POR2X1_329/A 0.03fF
C21985 PAND2X1_307/O POR2X1_102/Y 0.03fF
C21986 POR2X1_60/A POR2X1_295/O 0.00fF
C21987 POR2X1_826/Y POR2X1_42/Y 0.00fF
C21988 PAND2X1_404/Y PAND2X1_734/B 0.03fF
C21989 PAND2X1_42/CTRL2 POR2X1_267/A 0.03fF
C21990 D_INPUT_5 PAND2X1_17/CTRL2 0.00fF
C21991 PAND2X1_404/Y PAND2X1_573/a_16_344# 0.01fF
C21992 PAND2X1_557/A PAND2X1_221/O 0.01fF
C21993 PAND2X1_796/O PAND2X1_783/Y 0.03fF
C21994 POR2X1_287/A POR2X1_249/O 0.01fF
C21995 POR2X1_32/A PAND2X1_736/CTRL 0.01fF
C21996 PAND2X1_473/Y PAND2X1_571/CTRL2 0.03fF
C21997 POR2X1_554/B POR2X1_840/B 0.03fF
C21998 PAND2X1_5/m4_208_n4# POR2X1_612/A 0.01fF
C21999 POR2X1_411/B PAND2X1_566/Y 0.14fF
C22000 D_INPUT_0 VDD 5.05fF
C22001 POR2X1_848/A POR2X1_790/CTRL 0.08fF
C22002 POR2X1_260/B POR2X1_7/B 0.77fF
C22003 POR2X1_67/Y POR2X1_391/CTRL2 0.00fF
C22004 POR2X1_77/Y PAND2X1_169/CTRL2 0.09fF
C22005 POR2X1_68/A POR2X1_831/O 0.02fF
C22006 PAND2X1_23/Y PAND2X1_487/CTRL 0.06fF
C22007 POR2X1_474/O POR2X1_860/A 0.01fF
C22008 POR2X1_830/Y POR2X1_830/A 0.14fF
C22009 PAND2X1_860/A PAND2X1_853/B 0.04fF
C22010 GATE_479 PAND2X1_478/B 0.12fF
C22011 POR2X1_605/CTRL2 PAND2X1_90/Y 0.06fF
C22012 POR2X1_547/O POR2X1_624/Y 0.09fF
C22013 POR2X1_491/O PAND2X1_558/Y 0.00fF
C22014 POR2X1_149/A PAND2X1_90/Y 0.00fF
C22015 PAND2X1_651/Y POR2X1_63/Y 0.05fF
C22016 PAND2X1_41/B POR2X1_330/Y 0.03fF
C22017 POR2X1_55/CTRL VDD 0.00fF
C22018 POR2X1_566/A POR2X1_220/B 0.07fF
C22019 POR2X1_257/A POR2X1_56/Y 0.02fF
C22020 POR2X1_39/CTRL POR2X1_72/B 0.01fF
C22021 POR2X1_597/Y PAND2X1_643/Y 4.66fF
C22022 POR2X1_490/Y PAND2X1_197/Y 0.16fF
C22023 POR2X1_341/A D_INPUT_1 0.07fF
C22024 PAND2X1_435/Y VDD 0.04fF
C22025 PAND2X1_557/A PAND2X1_740/O 0.02fF
C22026 POR2X1_78/B POR2X1_788/A 0.05fF
C22027 POR2X1_651/Y PAND2X1_48/A 0.03fF
C22028 POR2X1_60/A POR2X1_497/Y 0.03fF
C22029 POR2X1_677/a_56_344# PAND2X1_390/Y 0.00fF
C22030 POR2X1_260/B PAND2X1_753/m4_208_n4# 0.01fF
C22031 PAND2X1_362/B POR2X1_594/O 0.01fF
C22032 PAND2X1_793/Y POR2X1_487/O 0.01fF
C22033 POR2X1_311/Y INPUT_0 0.06fF
C22034 POR2X1_268/Y POR2X1_5/Y 0.07fF
C22035 POR2X1_682/Y POR2X1_603/Y 0.01fF
C22036 POR2X1_83/B PAND2X1_738/Y 0.05fF
C22037 POR2X1_341/A POR2X1_724/A 0.03fF
C22038 POR2X1_270/Y POR2X1_659/CTRL 0.01fF
C22039 POR2X1_56/O PAND2X1_254/Y 0.00fF
C22040 PAND2X1_630/B PAND2X1_156/A 0.22fF
C22041 PAND2X1_432/CTRL2 VDD -0.00fF
C22042 D_INPUT_0 PAND2X1_351/a_76_28# 0.04fF
C22043 POR2X1_96/A POR2X1_102/Y 0.31fF
C22044 PAND2X1_45/CTRL2 POR2X1_260/A 0.00fF
C22045 D_INPUT_0 POR2X1_501/CTRL2 0.01fF
C22046 POR2X1_225/CTRL POR2X1_293/Y 0.00fF
C22047 POR2X1_853/O POR2X1_78/A 0.07fF
C22048 POR2X1_188/A POR2X1_285/O 0.01fF
C22049 PAND2X1_61/Y POR2X1_5/Y 0.02fF
C22050 POR2X1_586/Y POR2X1_293/Y 0.03fF
C22051 POR2X1_448/Y POR2X1_449/Y 0.00fF
C22052 POR2X1_68/A POR2X1_855/CTRL 0.01fF
C22053 POR2X1_66/B POR2X1_244/B 0.06fF
C22054 POR2X1_814/B POR2X1_621/B 0.05fF
C22055 POR2X1_502/A PAND2X1_279/O 0.04fF
C22056 PAND2X1_787/A PAND2X1_211/O 0.00fF
C22057 POR2X1_70/CTRL2 POR2X1_40/Y 0.01fF
C22058 PAND2X1_362/B POR2X1_331/Y 0.13fF
C22059 PAND2X1_475/a_16_344# INPUT_0 0.01fF
C22060 PAND2X1_659/O POR2X1_72/B 0.01fF
C22061 POR2X1_315/Y POR2X1_411/B 0.16fF
C22062 POR2X1_198/B POR2X1_590/A 0.01fF
C22063 POR2X1_686/m4_208_n4# PAND2X1_39/B 0.01fF
C22064 PAND2X1_58/A POR2X1_756/CTRL2 0.00fF
C22065 POR2X1_498/CTRL2 POR2X1_72/B 0.03fF
C22066 POR2X1_78/B POR2X1_456/O 0.03fF
C22067 POR2X1_57/O PAND2X1_219/A 0.10fF
C22068 PAND2X1_738/B VDD 0.05fF
C22069 POR2X1_388/CTRL POR2X1_66/A 0.01fF
C22070 POR2X1_432/Y POR2X1_236/Y 0.03fF
C22071 POR2X1_128/CTRL POR2X1_750/B 0.14fF
C22072 POR2X1_335/A POR2X1_296/B 0.02fF
C22073 POR2X1_46/Y POR2X1_40/Y 0.10fF
C22074 PAND2X1_850/Y POR2X1_677/Y 0.07fF
C22075 PAND2X1_93/B PAND2X1_88/Y 0.07fF
C22076 POR2X1_241/B POR2X1_222/Y 0.03fF
C22077 PAND2X1_340/B POR2X1_7/A 0.03fF
C22078 INPUT_1 PAND2X1_33/a_16_344# 0.02fF
C22079 POR2X1_260/B PAND2X1_60/B 0.49fF
C22080 PAND2X1_118/O POR2X1_78/A 0.05fF
C22081 D_INPUT_0 PAND2X1_32/B 1.26fF
C22082 POR2X1_445/A POR2X1_181/B 0.03fF
C22083 POR2X1_48/A PAND2X1_655/B 0.01fF
C22084 POR2X1_222/O POR2X1_222/A 0.02fF
C22085 POR2X1_65/A POR2X1_693/CTRL2 0.03fF
C22086 PAND2X1_90/Y VDD 10.65fF
C22087 POR2X1_13/A PAND2X1_714/A 0.24fF
C22088 PAND2X1_685/a_16_344# POR2X1_603/Y 0.01fF
C22089 POR2X1_41/B POR2X1_278/CTRL2 0.00fF
C22090 POR2X1_840/CTRL2 POR2X1_660/Y 0.01fF
C22091 PAND2X1_20/A D_GATE_222 0.19fF
C22092 POR2X1_646/A PAND2X1_48/A 0.01fF
C22093 POR2X1_423/Y POR2X1_293/Y 4.66fF
C22094 POR2X1_646/B POR2X1_294/A -0.06fF
C22095 PAND2X1_808/B PAND2X1_592/Y 0.01fF
C22096 POR2X1_567/B POR2X1_704/CTRL2 0.03fF
C22097 PAND2X1_845/CTRL2 POR2X1_60/A 0.03fF
C22098 PAND2X1_496/O POR2X1_777/B 0.02fF
C22099 PAND2X1_90/Y POR2X1_793/a_16_28# 0.13fF
C22100 POR2X1_719/CTRL POR2X1_66/A 0.01fF
C22101 PAND2X1_7/CTRL POR2X1_750/B 0.11fF
C22102 POR2X1_52/A POR2X1_847/B 0.03fF
C22103 POR2X1_614/A POR2X1_850/B 0.03fF
C22104 POR2X1_330/Y POR2X1_130/Y 0.03fF
C22105 POR2X1_441/Y POR2X1_373/Y 0.04fF
C22106 POR2X1_66/B POR2X1_793/A 0.06fF
C22107 PAND2X1_771/Y POR2X1_765/Y 0.06fF
C22108 POR2X1_809/A POR2X1_864/A 0.05fF
C22109 PAND2X1_859/A POR2X1_382/CTRL 0.01fF
C22110 POR2X1_52/A PAND2X1_76/Y 0.00fF
C22111 D_INPUT_2 POR2X1_293/CTRL 0.01fF
C22112 POR2X1_121/CTRL2 POR2X1_590/A 0.01fF
C22113 POR2X1_856/a_16_28# POR2X1_855/Y 0.01fF
C22114 POR2X1_287/B POR2X1_294/B 0.03fF
C22115 POR2X1_679/B PAND2X1_205/A 0.02fF
C22116 POR2X1_669/B POR2X1_320/m4_208_n4# 0.17fF
C22117 POR2X1_865/B POR2X1_78/A 0.03fF
C22118 POR2X1_68/A POR2X1_35/B 0.03fF
C22119 POR2X1_108/CTRL2 POR2X1_60/A 0.04fF
C22120 POR2X1_254/Y POR2X1_332/B 0.07fF
C22121 PAND2X1_96/B POR2X1_675/CTRL 0.01fF
C22122 POR2X1_669/B PAND2X1_149/A 0.03fF
C22123 POR2X1_263/Y POR2X1_235/a_76_344# 0.00fF
C22124 PAND2X1_433/CTRL2 POR2X1_480/A -0.01fF
C22125 PAND2X1_11/Y INPUT_6 0.20fF
C22126 PAND2X1_23/Y POR2X1_362/B 0.07fF
C22127 POR2X1_150/Y POR2X1_385/Y 0.03fF
C22128 POR2X1_121/B PAND2X1_583/a_76_28# 0.04fF
C22129 POR2X1_555/B POR2X1_228/Y 0.01fF
C22130 POR2X1_649/CTRL POR2X1_643/A 0.03fF
C22131 PAND2X1_570/B PAND2X1_577/Y 0.07fF
C22132 POR2X1_49/Y POR2X1_56/Y 0.03fF
C22133 POR2X1_483/A POR2X1_294/B 0.04fF
C22134 POR2X1_467/Y POR2X1_788/B 0.05fF
C22135 POR2X1_260/B POR2X1_332/O 0.01fF
C22136 PAND2X1_354/A PAND2X1_354/a_16_344# 0.02fF
C22137 POR2X1_641/CTRL POR2X1_318/A 0.05fF
C22138 POR2X1_139/Y VDD 0.10fF
C22139 POR2X1_368/CTRL POR2X1_293/Y 0.02fF
C22140 PAND2X1_73/Y POR2X1_366/A 0.03fF
C22141 POR2X1_329/A POR2X1_39/B 0.10fF
C22142 PAND2X1_90/Y POR2X1_741/Y 0.05fF
C22143 POR2X1_840/B PAND2X1_74/a_56_28# 0.00fF
C22144 POR2X1_15/O POR2X1_69/A 0.01fF
C22145 POR2X1_502/A POR2X1_307/Y 0.03fF
C22146 PAND2X1_673/Y POR2X1_7/B 0.03fF
C22147 POR2X1_625/Y POR2X1_754/A 0.06fF
C22148 POR2X1_43/B POR2X1_58/CTRL2 0.03fF
C22149 POR2X1_102/Y POR2X1_7/A 2.21fF
C22150 POR2X1_294/B PAND2X1_8/Y 0.05fF
C22151 POR2X1_814/B PAND2X1_411/a_76_28# 0.01fF
C22152 PAND2X1_96/B POR2X1_389/Y 0.03fF
C22153 POR2X1_483/CTRL POR2X1_193/A 0.00fF
C22154 POR2X1_443/A POR2X1_192/B 0.36fF
C22155 POR2X1_596/A POR2X1_808/A 0.17fF
C22156 POR2X1_16/A PAND2X1_571/O -0.01fF
C22157 POR2X1_388/a_76_344# POR2X1_750/B 0.01fF
C22158 POR2X1_673/Y D_INPUT_0 0.03fF
C22159 PAND2X1_425/m4_208_n4# POR2X1_17/m4_208_n4# 0.13fF
C22160 POR2X1_215/CTRL2 POR2X1_740/Y 0.28fF
C22161 PAND2X1_809/B POR2X1_760/A 0.07fF
C22162 POR2X1_174/A POR2X1_180/A 10.02fF
C22163 POR2X1_433/O PAND2X1_349/A 0.01fF
C22164 POR2X1_83/a_16_28# POR2X1_23/Y 0.02fF
C22165 PAND2X1_94/A PAND2X1_15/CTRL 0.01fF
C22166 PAND2X1_830/CTRL2 POR2X1_60/A 0.06fF
C22167 PAND2X1_477/B PAND2X1_803/A 0.00fF
C22168 POR2X1_164/O POR2X1_376/B 0.19fF
C22169 PAND2X1_48/B PAND2X1_131/a_16_344# 0.02fF
C22170 POR2X1_249/Y POR2X1_296/B 0.03fF
C22171 POR2X1_174/CTRL2 PAND2X1_73/Y 0.01fF
C22172 POR2X1_333/O POR2X1_241/B 0.01fF
C22173 POR2X1_330/Y POR2X1_228/Y 0.05fF
C22174 PAND2X1_115/Y PAND2X1_553/B 0.07fF
C22175 POR2X1_83/B POR2X1_172/CTRL2 0.09fF
C22176 POR2X1_368/a_16_28# POR2X1_372/Y 0.06fF
C22177 POR2X1_55/CTRL POR2X1_673/Y 0.02fF
C22178 POR2X1_455/CTRL POR2X1_702/A 0.00fF
C22179 PAND2X1_139/B POR2X1_184/Y 0.61fF
C22180 POR2X1_325/A POR2X1_140/A 0.00fF
C22181 PAND2X1_90/Y PAND2X1_32/B 3.17fF
C22182 PAND2X1_578/a_76_28# PAND2X1_577/Y 0.01fF
C22183 POR2X1_748/A POR2X1_283/A 0.03fF
C22184 PAND2X1_808/Y POR2X1_96/A 0.03fF
C22185 PAND2X1_257/CTRL POR2X1_222/Y 0.03fF
C22186 POR2X1_61/CTRL PAND2X1_58/A 0.02fF
C22187 PAND2X1_218/A INPUT_0 0.01fF
C22188 POR2X1_38/B POR2X1_236/CTRL 0.03fF
C22189 PAND2X1_865/a_16_344# POR2X1_516/Y 0.02fF
C22190 PAND2X1_614/O POR2X1_245/Y 0.04fF
C22191 PAND2X1_643/CTRL2 POR2X1_7/B 0.01fF
C22192 POR2X1_174/B POR2X1_174/O 0.05fF
C22193 POR2X1_502/A PAND2X1_411/O 0.05fF
C22194 POR2X1_859/A POR2X1_793/A 0.03fF
C22195 PAND2X1_48/B POR2X1_664/Y 0.04fF
C22196 PAND2X1_469/B PAND2X1_804/B 0.30fF
C22197 POR2X1_421/O POR2X1_90/Y 0.00fF
C22198 POR2X1_355/B POR2X1_35/Y 0.03fF
C22199 PAND2X1_617/a_16_344# PAND2X1_52/B 0.04fF
C22200 POR2X1_614/A POR2X1_483/CTRL 0.03fF
C22201 POR2X1_115/CTRL2 POR2X1_112/Y 0.01fF
C22202 POR2X1_230/a_16_28# POR2X1_38/Y 0.06fF
C22203 POR2X1_336/CTRL VDD 0.00fF
C22204 POR2X1_96/A POR2X1_531/Y 0.02fF
C22205 POR2X1_763/Y PAND2X1_324/Y 0.01fF
C22206 POR2X1_13/A POR2X1_816/A 0.03fF
C22207 POR2X1_785/A POR2X1_341/CTRL2 0.03fF
C22208 POR2X1_66/A POR2X1_773/A 0.54fF
C22209 PAND2X1_562/B PAND2X1_854/A 0.05fF
C22210 POR2X1_158/Y POR2X1_485/Y 0.00fF
C22211 POR2X1_393/Y POR2X1_394/CTRL 0.01fF
C22212 POR2X1_394/Y POR2X1_394/O 0.01fF
C22213 PAND2X1_856/O POR2X1_102/Y 0.01fF
C22214 POR2X1_111/CTRL VDD 0.00fF
C22215 POR2X1_213/B POR2X1_148/B 0.02fF
C22216 POR2X1_813/O POR2X1_39/B 0.04fF
C22217 POR2X1_41/B POR2X1_310/CTRL 0.05fF
C22218 POR2X1_38/Y INPUT_0 9.87fF
C22219 PAND2X1_65/CTRL2 POR2X1_4/Y 0.01fF
C22220 PAND2X1_319/B PAND2X1_151/CTRL2 0.01fF
C22221 PAND2X1_671/CTRL POR2X1_35/B 0.01fF
C22222 POR2X1_68/A PAND2X1_275/CTRL2 0.07fF
C22223 POR2X1_62/Y PAND2X1_10/O 0.17fF
C22224 POR2X1_502/A POR2X1_68/B 0.08fF
C22225 PAND2X1_469/Y POR2X1_236/Y 0.16fF
C22226 POR2X1_348/CTRL2 VDD 0.00fF
C22227 POR2X1_606/Y POR2X1_774/A 0.06fF
C22228 PAND2X1_317/Y PAND2X1_566/Y 0.07fF
C22229 POR2X1_759/A POR2X1_7/B 0.13fF
C22230 PAND2X1_643/O POR2X1_13/Y 0.02fF
C22231 PAND2X1_7/Y POR2X1_260/A 0.04fF
C22232 POR2X1_262/CTRL POR2X1_73/Y 0.01fF
C22233 POR2X1_51/A POR2X1_3/A 0.00fF
C22234 PAND2X1_610/CTRL POR2X1_48/A 0.01fF
C22235 PAND2X1_65/B POR2X1_576/CTRL2 0.01fF
C22236 PAND2X1_352/A PAND2X1_352/B 0.00fF
C22237 POR2X1_67/O POR2X1_39/B 0.19fF
C22238 PAND2X1_473/B PAND2X1_175/CTRL2 0.03fF
C22239 PAND2X1_48/B POR2X1_112/Y 0.03fF
C22240 POR2X1_48/A PAND2X1_508/B 0.03fF
C22241 POR2X1_539/A POR2X1_370/Y 0.07fF
C22242 PAND2X1_65/B POR2X1_773/B 0.05fF
C22243 GATE_741 PAND2X1_366/A 0.01fF
C22244 POR2X1_29/A POR2X1_4/Y 0.26fF
C22245 POR2X1_41/B PAND2X1_338/B 0.03fF
C22246 POR2X1_13/A PAND2X1_854/A 0.16fF
C22247 POR2X1_673/Y PAND2X1_90/Y 0.15fF
C22248 POR2X1_108/Y VDD -0.00fF
C22249 POR2X1_294/B POR2X1_209/A 0.19fF
C22250 PAND2X1_803/Y PAND2X1_553/B 0.07fF
C22251 POR2X1_327/Y POR2X1_186/Y 0.17fF
C22252 POR2X1_750/B POR2X1_735/CTRL2 0.30fF
C22253 POR2X1_537/Y POR2X1_830/CTRL 0.01fF
C22254 POR2X1_66/B POR2X1_537/Y 0.03fF
C22255 POR2X1_79/Y POR2X1_283/A 0.03fF
C22256 PAND2X1_865/Y PAND2X1_794/CTRL -0.01fF
C22257 PAND2X1_90/A PAND2X1_150/a_56_28# 0.00fF
C22258 POR2X1_16/A PAND2X1_804/A 0.02fF
C22259 POR2X1_65/A POR2X1_83/m4_208_n4# 0.09fF
C22260 POR2X1_68/A POR2X1_219/O 0.01fF
C22261 PAND2X1_231/a_16_344# POR2X1_153/Y 0.05fF
C22262 PAND2X1_279/O POR2X1_188/Y 0.02fF
C22263 PAND2X1_449/Y POR2X1_90/Y 0.01fF
C22264 POR2X1_407/A POR2X1_644/A 0.27fF
C22265 PAND2X1_849/B POR2X1_88/Y 0.02fF
C22266 POR2X1_370/CTRL POR2X1_543/A 0.01fF
C22267 PAND2X1_55/Y PAND2X1_60/B 3.66fF
C22268 POR2X1_55/Y POR2X1_530/Y 0.02fF
C22269 INPUT_1 INPUT_0 1.53fF
C22270 POR2X1_188/A POR2X1_537/Y 0.03fF
C22271 POR2X1_52/A POR2X1_315/Y 0.01fF
C22272 POR2X1_71/CTRL2 PAND2X1_84/Y 0.01fF
C22273 POR2X1_672/CTRL POR2X1_38/B 0.01fF
C22274 POR2X1_114/O POR2X1_68/B 0.01fF
C22275 POR2X1_313/CTRL POR2X1_90/Y 0.00fF
C22276 PAND2X1_341/A POR2X1_52/Y 1.27fF
C22277 POR2X1_208/Y POR2X1_206/CTRL2 0.03fF
C22278 PAND2X1_61/a_16_344# POR2X1_39/B 0.04fF
C22279 POR2X1_394/A POR2X1_236/Y 1.04fF
C22280 POR2X1_502/A POR2X1_502/O 0.15fF
C22281 POR2X1_840/B POR2X1_702/A 0.03fF
C22282 POR2X1_78/A POR2X1_568/B 0.08fF
C22283 PAND2X1_632/A POR2X1_55/Y 0.03fF
C22284 PAND2X1_41/B POR2X1_337/Y 0.18fF
C22285 POR2X1_859/A POR2X1_753/CTRL2 0.02fF
C22286 POR2X1_267/Y POR2X1_361/CTRL2 0.03fF
C22287 POR2X1_788/Y PAND2X1_60/B 0.01fF
C22288 PAND2X1_583/a_16_344# PAND2X1_32/B 0.02fF
C22289 PAND2X1_658/A PAND2X1_549/B 0.01fF
C22290 POR2X1_315/Y POR2X1_152/A 0.07fF
C22291 INPUT_0 POR2X1_153/Y 0.19fF
C22292 POR2X1_402/A PAND2X1_60/B 0.04fF
C22293 PAND2X1_23/Y POR2X1_553/A 0.03fF
C22294 POR2X1_190/Y POR2X1_444/Y 0.03fF
C22295 POR2X1_307/B PAND2X1_48/A 0.02fF
C22296 POR2X1_384/A INPUT_0 0.05fF
C22297 POR2X1_574/O POR2X1_574/A 0.03fF
C22298 PAND2X1_480/B PAND2X1_112/m4_208_n4# 0.04fF
C22299 POR2X1_528/O POR2X1_528/Y 0.02fF
C22300 POR2X1_102/a_56_344# POR2X1_40/Y 0.00fF
C22301 PAND2X1_96/B POR2X1_318/A 0.15fF
C22302 PAND2X1_57/B POR2X1_186/B 0.03fF
C22303 PAND2X1_610/a_16_344# POR2X1_40/Y 0.02fF
C22304 PAND2X1_858/CTRL2 INPUT_0 0.10fF
C22305 POR2X1_119/Y POR2X1_122/Y 0.02fF
C22306 POR2X1_81/Y POR2X1_394/A 0.10fF
C22307 PAND2X1_55/Y POR2X1_353/A 0.01fF
C22308 PAND2X1_6/Y PAND2X1_368/CTRL2 0.01fF
C22309 POR2X1_326/A POR2X1_502/A 0.00fF
C22310 POR2X1_65/A PAND2X1_326/B 0.09fF
C22311 PAND2X1_659/Y POR2X1_393/CTRL 0.00fF
C22312 POR2X1_96/A PAND2X1_354/Y 0.16fF
C22313 POR2X1_379/CTRL2 POR2X1_532/A 0.07fF
C22314 POR2X1_816/A PAND2X1_510/B 0.02fF
C22315 POR2X1_29/A POR2X1_80/a_16_28# 0.03fF
C22316 PAND2X1_720/CTRL2 POR2X1_73/Y -0.01fF
C22317 INPUT_1 POR2X1_618/a_16_28# 0.00fF
C22318 PAND2X1_484/CTRL2 POR2X1_294/B 0.03fF
C22319 POR2X1_167/O POR2X1_90/Y 0.01fF
C22320 POR2X1_208/A POR2X1_532/A 0.01fF
C22321 POR2X1_61/A VDD -0.00fF
C22322 POR2X1_23/Y PAND2X1_860/A 0.03fF
C22323 PAND2X1_728/O POR2X1_816/A 0.02fF
C22324 PAND2X1_6/Y PAND2X1_528/a_16_344# 0.01fF
C22325 PAND2X1_798/Y PAND2X1_363/Y 0.75fF
C22326 POR2X1_188/A POR2X1_285/B 0.00fF
C22327 POR2X1_16/A POR2X1_315/O 0.01fF
C22328 POR2X1_701/a_16_28# POR2X1_236/Y -0.00fF
C22329 PAND2X1_643/A VDD 0.13fF
C22330 POR2X1_333/A POR2X1_161/O 0.05fF
C22331 POR2X1_196/CTRL POR2X1_740/Y 0.29fF
C22332 POR2X1_612/A POR2X1_612/a_16_28# 0.02fF
C22333 PAND2X1_39/B PAND2X1_32/CTRL2 0.05fF
C22334 POR2X1_390/B PAND2X1_69/A 0.04fF
C22335 PAND2X1_738/CTRL POR2X1_39/B 0.01fF
C22336 PAND2X1_863/B PAND2X1_729/CTRL2 0.01fF
C22337 POR2X1_275/a_16_28# POR2X1_394/A 0.02fF
C22338 POR2X1_326/A POR2X1_532/Y 0.07fF
C22339 POR2X1_96/A POR2X1_74/Y 0.08fF
C22340 POR2X1_385/Y PAND2X1_364/B 0.12fF
C22341 PAND2X1_798/B POR2X1_129/Y 0.01fF
C22342 POR2X1_826/CTRL POR2X1_77/Y 0.01fF
C22343 POR2X1_41/CTRL POR2X1_73/Y 0.02fF
C22344 PAND2X1_330/CTRL POR2X1_331/A 0.05fF
C22345 PAND2X1_79/Y POR2X1_456/B 0.03fF
C22346 POR2X1_777/Y POR2X1_725/Y 0.02fF
C22347 POR2X1_57/A POR2X1_527/O 0.02fF
C22348 PAND2X1_803/CTRL2 POR2X1_90/Y 0.00fF
C22349 POR2X1_299/CTRL PAND2X1_308/Y 0.01fF
C22350 POR2X1_332/Y D_GATE_222 0.02fF
C22351 POR2X1_456/B POR2X1_736/O 0.15fF
C22352 PAND2X1_862/B POR2X1_184/CTRL 0.03fF
C22353 PAND2X1_6/A PAND2X1_508/Y 0.07fF
C22354 PAND2X1_799/CTRL PAND2X1_539/Y 0.01fF
C22355 POR2X1_71/a_16_28# POR2X1_43/B 0.02fF
C22356 POR2X1_822/CTRL POR2X1_77/Y 0.01fF
C22357 PAND2X1_801/O PAND2X1_863/B 0.02fF
C22358 POR2X1_114/B PAND2X1_48/A 0.10fF
C22359 POR2X1_63/Y POR2X1_813/CTRL2 0.04fF
C22360 PAND2X1_96/B POR2X1_574/Y 0.04fF
C22361 PAND2X1_744/O POR2X1_294/A 0.06fF
C22362 POR2X1_16/A PAND2X1_656/A 0.07fF
C22363 PAND2X1_797/Y PAND2X1_213/A 0.07fF
C22364 POR2X1_51/B POR2X1_31/a_56_344# 0.00fF
C22365 D_INPUT_7 PAND2X1_429/CTRL2 0.00fF
C22366 POR2X1_204/CTRL2 POR2X1_4/Y 0.01fF
C22367 POR2X1_48/A POR2X1_329/A 0.10fF
C22368 PAND2X1_639/Y POR2X1_43/B 0.04fF
C22369 POR2X1_162/Y POR2X1_210/B 0.04fF
C22370 POR2X1_383/A POR2X1_758/Y 0.10fF
C22371 POR2X1_556/A POR2X1_446/B 0.02fF
C22372 POR2X1_532/A PAND2X1_394/CTRL2 0.03fF
C22373 PAND2X1_242/Y POR2X1_423/Y 0.16fF
C22374 PAND2X1_632/A PAND2X1_508/O 0.02fF
C22375 POR2X1_16/A PAND2X1_124/CTRL2 0.01fF
C22376 POR2X1_410/O PAND2X1_52/B 0.01fF
C22377 PAND2X1_20/A PAND2X1_607/O 0.04fF
C22378 PAND2X1_23/Y D_INPUT_4 0.03fF
C22379 PAND2X1_127/CTRL POR2X1_456/B 0.00fF
C22380 POR2X1_688/CTRL2 D_INPUT_0 0.00fF
C22381 POR2X1_304/O POR2X1_43/B 0.01fF
C22382 POR2X1_168/A POR2X1_578/Y 0.03fF
C22383 POR2X1_540/A POR2X1_552/A 0.01fF
C22384 POR2X1_510/A POR2X1_568/B 0.03fF
C22385 POR2X1_54/Y PAND2X1_618/Y 0.00fF
C22386 POR2X1_23/Y POR2X1_253/CTRL2 0.03fF
C22387 PAND2X1_859/A POR2X1_9/Y 0.05fF
C22388 PAND2X1_93/B POR2X1_341/A 0.07fF
C22389 POR2X1_394/A POR2X1_757/Y 0.06fF
C22390 POR2X1_283/A PAND2X1_730/A 0.03fF
C22391 POR2X1_760/A POR2X1_102/Y 0.05fF
C22392 POR2X1_257/A PAND2X1_771/Y 0.02fF
C22393 VDD POR2X1_173/Y 0.00fF
C22394 PAND2X1_9/Y D_INPUT_0 0.06fF
C22395 POR2X1_270/Y PAND2X1_268/O 0.08fF
C22396 POR2X1_311/CTRL PAND2X1_336/Y 0.01fF
C22397 POR2X1_814/B PAND2X1_607/O 0.04fF
C22398 PAND2X1_341/A PAND2X1_358/CTRL2 0.00fF
C22399 POR2X1_69/Y POR2X1_94/A 0.05fF
C22400 POR2X1_556/Y POR2X1_632/Y 0.01fF
C22401 POR2X1_416/B PAND2X1_357/Y 0.03fF
C22402 POR2X1_509/CTRL2 POR2X1_35/Y 0.01fF
C22403 POR2X1_193/A POR2X1_556/CTRL2 0.04fF
C22404 POR2X1_848/O POR2X1_734/A 0.05fF
C22405 POR2X1_294/A PAND2X1_103/CTRL 0.03fF
C22406 POR2X1_568/Y POR2X1_551/A 0.05fF
C22407 POR2X1_741/Y POR2X1_715/O 0.01fF
C22408 POR2X1_475/CTRL POR2X1_590/A 0.00fF
C22409 POR2X1_57/A POR2X1_39/B 4.84fF
C22410 POR2X1_137/a_16_28# POR2X1_768/A 0.05fF
C22411 PAND2X1_3/A PAND2X1_26/A 0.03fF
C22412 POR2X1_38/Y POR2X1_522/CTRL2 0.06fF
C22413 PAND2X1_699/CTRL POR2X1_750/B 0.02fF
C22414 PAND2X1_846/O POR2X1_38/B 0.01fF
C22415 POR2X1_96/A POR2X1_677/Y 0.03fF
C22416 PAND2X1_826/CTRL POR2X1_202/B 0.01fF
C22417 PAND2X1_838/B POR2X1_83/B 0.03fF
C22418 PAND2X1_222/A POR2X1_32/A 0.03fF
C22419 PAND2X1_338/B POR2X1_77/Y 0.12fF
C22420 POR2X1_8/Y POR2X1_749/Y 0.00fF
C22421 POR2X1_685/O POR2X1_814/A 0.29fF
C22422 POR2X1_614/A POR2X1_556/CTRL2 0.09fF
C22423 POR2X1_715/O PAND2X1_32/B 0.02fF
C22424 POR2X1_54/Y PAND2X1_20/A 0.19fF
C22425 POR2X1_85/Y PAND2X1_338/B 0.03fF
C22426 PAND2X1_140/A POR2X1_416/B 0.03fF
C22427 POR2X1_454/A POR2X1_555/B 0.09fF
C22428 POR2X1_444/Y POR2X1_738/CTRL 0.03fF
C22429 POR2X1_411/B PAND2X1_558/Y 0.03fF
C22430 POR2X1_343/Y POR2X1_575/O 0.28fF
C22431 POR2X1_85/Y POR2X1_235/CTRL 0.01fF
C22432 POR2X1_528/Y POR2X1_416/B 0.10fF
C22433 POR2X1_78/B PAND2X1_418/CTRL2 0.05fF
C22434 PAND2X1_20/A POR2X1_202/A 0.07fF
C22435 POR2X1_707/CTRL D_INPUT_4 0.03fF
C22436 POR2X1_326/A POR2X1_188/Y 0.16fF
C22437 D_INPUT_0 PAND2X1_591/a_16_344# 0.01fF
C22438 POR2X1_744/O POR2X1_39/B 0.16fF
C22439 POR2X1_554/B POR2X1_217/CTRL 0.01fF
C22440 POR2X1_832/A PAND2X1_72/A 0.80fF
C22441 POR2X1_376/B PAND2X1_98/CTRL2 0.01fF
C22442 POR2X1_807/CTRL2 POR2X1_590/A 0.01fF
C22443 PAND2X1_737/B PAND2X1_198/O 0.02fF
C22444 POR2X1_78/B POR2X1_659/a_16_28# 0.11fF
C22445 POR2X1_41/B PAND2X1_717/A 0.07fF
C22446 PAND2X1_65/B POR2X1_227/B 0.03fF
C22447 POR2X1_65/A POR2X1_253/O 0.02fF
C22448 POR2X1_736/A POR2X1_675/Y 0.39fF
C22449 PAND2X1_96/CTRL POR2X1_202/A 0.03fF
C22450 POR2X1_54/Y POR2X1_814/B 0.18fF
C22451 POR2X1_341/A POR2X1_573/CTRL 0.07fF
C22452 POR2X1_620/A POR2X1_296/B 0.01fF
C22453 PAND2X1_65/B POR2X1_471/A 0.03fF
C22454 PAND2X1_255/CTRL2 POR2X1_786/Y 0.02fF
C22455 POR2X1_343/Y POR2X1_833/A 0.03fF
C22456 POR2X1_260/B POR2X1_750/B 0.46fF
C22457 D_INPUT_0 POR2X1_267/A 0.03fF
C22458 PAND2X1_341/Y POR2X1_77/Y 0.10fF
C22459 POR2X1_78/B PAND2X1_41/CTRL 0.01fF
C22460 PAND2X1_435/CTRL2 POR2X1_20/B 0.01fF
C22461 POR2X1_544/B POR2X1_736/A 0.05fF
C22462 POR2X1_519/O POR2X1_43/Y 0.00fF
C22463 POR2X1_77/Y PAND2X1_337/CTRL2 0.01fF
C22464 POR2X1_514/Y POR2X1_814/A 0.03fF
C22465 POR2X1_65/A PAND2X1_852/A 0.01fF
C22466 POR2X1_260/B PAND2X1_13/O 0.17fF
C22467 POR2X1_669/B POR2X1_819/a_76_344# 0.10fF
C22468 PAND2X1_480/B POR2X1_411/B 0.18fF
C22469 PAND2X1_848/a_56_28# POR2X1_669/B 0.00fF
C22470 POR2X1_525/CTRL2 POR2X1_23/Y 0.03fF
C22471 POR2X1_260/O POR2X1_741/Y 0.01fF
C22472 POR2X1_558/B PAND2X1_41/B 0.09fF
C22473 POR2X1_808/A POR2X1_811/A 0.06fF
C22474 POR2X1_854/CTRL POR2X1_192/Y 0.01fF
C22475 POR2X1_78/B POR2X1_644/CTRL 0.03fF
C22476 POR2X1_48/A PAND2X1_738/CTRL 0.01fF
C22477 POR2X1_63/Y POR2X1_406/CTRL2 0.01fF
C22478 POR2X1_474/a_76_344# POR2X1_590/A 0.01fF
C22479 PAND2X1_841/CTRL2 POR2X1_411/B 0.01fF
C22480 POR2X1_32/A PAND2X1_168/Y 0.02fF
C22481 POR2X1_49/Y POR2X1_754/Y 0.07fF
C22482 PAND2X1_48/B POR2X1_541/B 0.02fF
C22483 POR2X1_327/Y POR2X1_717/B 0.03fF
C22484 POR2X1_302/Y POR2X1_274/A 0.56fF
C22485 POR2X1_9/Y POR2X1_7/A 0.24fF
C22486 POR2X1_14/Y POR2X1_748/A 0.05fF
C22487 POR2X1_102/Y PAND2X1_140/CTRL2 0.01fF
C22488 PAND2X1_56/Y POR2X1_556/A 0.05fF
C22489 POR2X1_748/A PAND2X1_453/A 0.05fF
C22490 POR2X1_411/B PAND2X1_398/CTRL 0.01fF
C22491 POR2X1_820/B POR2X1_48/A -0.00fF
C22492 PAND2X1_59/B VDD 0.35fF
C22493 PAND2X1_326/B PAND2X1_169/O 0.02fF
C22494 PAND2X1_244/CTRL POR2X1_72/B 0.01fF
C22495 POR2X1_460/Y POR2X1_459/B 0.01fF
C22496 POR2X1_35/B PAND2X1_58/A 0.03fF
C22497 PAND2X1_200/Y POR2X1_72/B 0.04fF
C22498 POR2X1_13/A POR2X1_93/Y 0.03fF
C22499 POR2X1_656/O POR2X1_362/B 0.18fF
C22500 POR2X1_629/B POR2X1_186/Y 0.03fF
C22501 PAND2X1_473/Y PAND2X1_576/B 0.40fF
C22502 POR2X1_60/A POR2X1_423/Y 0.03fF
C22503 POR2X1_502/A POR2X1_848/A 0.05fF
C22504 POR2X1_274/A PAND2X1_516/a_16_344# 0.01fF
C22505 POR2X1_843/a_56_344# POR2X1_287/B 0.00fF
C22506 POR2X1_32/A POR2X1_692/Y 0.00fF
C22507 POR2X1_48/A POR2X1_256/O 0.02fF
C22508 POR2X1_669/B POR2X1_236/Y 19.98fF
C22509 POR2X1_23/Y PAND2X1_515/O 0.02fF
C22510 POR2X1_673/A POR2X1_29/A 0.02fF
C22511 PAND2X1_39/B PAND2X1_29/CTRL 0.07fF
C22512 POR2X1_60/A PAND2X1_513/a_16_344# 0.02fF
C22513 POR2X1_41/B POR2X1_692/O 0.02fF
C22514 POR2X1_197/CTRL POR2X1_555/B 0.01fF
C22515 PAND2X1_236/O POR2X1_590/A 0.00fF
C22516 POR2X1_336/O POR2X1_556/A 0.10fF
C22517 PAND2X1_76/CTRL2 PAND2X1_76/Y 0.00fF
C22518 POR2X1_141/a_56_344# PAND2X1_20/A 0.00fF
C22519 POR2X1_644/B POR2X1_513/B 0.01fF
C22520 POR2X1_465/B POR2X1_66/A 0.03fF
C22521 PAND2X1_70/CTRL2 POR2X1_750/B 0.01fF
C22522 POR2X1_102/Y PAND2X1_719/CTRL 0.01fF
C22523 POR2X1_674/Y PAND2X1_740/Y 0.02fF
C22524 POR2X1_814/A POR2X1_773/B 0.03fF
C22525 POR2X1_97/O POR2X1_814/A 0.05fF
C22526 PAND2X1_580/O PAND2X1_578/Y 0.09fF
C22527 PAND2X1_787/Y POR2X1_40/Y 0.03fF
C22528 PAND2X1_10/a_76_28# PAND2X1_8/Y 0.02fF
C22529 POR2X1_41/B PAND2X1_623/O 0.08fF
C22530 POR2X1_808/A PAND2X1_90/Y 0.02fF
C22531 POR2X1_102/Y POR2X1_609/A 0.57fF
C22532 POR2X1_81/O PAND2X1_862/B 0.01fF
C22533 POR2X1_383/A POR2X1_556/A 0.14fF
C22534 POR2X1_48/A PAND2X1_506/a_16_344# 0.01fF
C22535 D_INPUT_5 D_INPUT_6 0.29fF
C22536 PAND2X1_717/A PAND2X1_308/Y 0.03fF
C22537 PAND2X1_206/O POR2X1_40/Y 0.01fF
C22538 PAND2X1_805/A PAND2X1_367/a_76_28# 0.01fF
C22539 PAND2X1_340/B POR2X1_38/Y 6.13fF
C22540 PAND2X1_620/Y POR2X1_627/O 0.11fF
C22541 POR2X1_150/Y PAND2X1_181/O 0.03fF
C22542 POR2X1_422/Y POR2X1_293/Y 0.03fF
C22543 POR2X1_137/Y POR2X1_624/Y 0.08fF
C22544 POR2X1_842/a_16_28# POR2X1_741/Y 0.00fF
C22545 POR2X1_464/a_16_28# POR2X1_750/B 0.01fF
C22546 PAND2X1_128/O PAND2X1_577/Y 0.06fF
C22547 POR2X1_65/A PAND2X1_206/CTRL 0.01fF
C22548 PAND2X1_59/B PAND2X1_32/B 0.19fF
C22549 POR2X1_375/Y POR2X1_7/B 0.01fF
C22550 POR2X1_174/B PAND2X1_23/Y 0.03fF
C22551 D_INPUT_2 POR2X1_414/CTRL 0.01fF
C22552 POR2X1_487/CTRL PAND2X1_794/B 0.01fF
C22553 PAND2X1_217/B PAND2X1_735/Y 0.10fF
C22554 POR2X1_814/B POR2X1_572/CTRL2 0.16fF
C22555 POR2X1_84/A PAND2X1_88/Y 0.03fF
C22556 POR2X1_291/CTRL POR2X1_20/B 0.01fF
C22557 PAND2X1_832/a_56_28# PAND2X1_499/Y 0.00fF
C22558 PAND2X1_420/CTRL POR2X1_785/A 0.01fF
C22559 POR2X1_48/A PAND2X1_702/CTRL 0.01fF
C22560 POR2X1_46/Y PAND2X1_706/O 0.01fF
C22561 PAND2X1_71/a_76_28# POR2X1_296/B 0.02fF
C22562 POR2X1_152/CTRL POR2X1_669/B 0.08fF
C22563 POR2X1_358/a_56_344# PAND2X1_20/A 0.00fF
C22564 PAND2X1_805/A VDD 0.39fF
C22565 POR2X1_805/CTRL2 PAND2X1_60/B 0.01fF
C22566 POR2X1_276/A POR2X1_446/B 0.03fF
C22567 POR2X1_475/O POR2X1_249/Y 0.01fF
C22568 POR2X1_62/Y POR2X1_329/A 0.03fF
C22569 POR2X1_783/A POR2X1_783/m4_208_n4# 0.01fF
C22570 POR2X1_311/Y PAND2X1_808/Y 0.03fF
C22571 POR2X1_56/B POR2X1_419/Y 0.56fF
C22572 POR2X1_66/B PAND2X1_48/B 0.70fF
C22573 PAND2X1_609/a_16_344# PAND2X1_60/B 0.01fF
C22574 POR2X1_436/CTRL POR2X1_802/B 0.01fF
C22575 POR2X1_505/Y POR2X1_7/B 0.03fF
C22576 PAND2X1_272/CTRL2 PAND2X1_32/B 0.01fF
C22577 POR2X1_57/A POR2X1_48/A 9.15fF
C22578 POR2X1_52/A PAND2X1_558/Y 0.03fF
C22579 POR2X1_322/CTRL2 POR2X1_72/B 0.01fF
C22580 POR2X1_621/B VDD 0.01fF
C22581 PAND2X1_675/A POR2X1_674/Y 0.02fF
C22582 POR2X1_866/CTRL2 POR2X1_800/A 0.08fF
C22583 POR2X1_477/A POR2X1_675/O 0.02fF
C22584 POR2X1_254/A PAND2X1_55/Y 0.03fF
C22585 POR2X1_748/A POR2X1_55/Y 0.03fF
C22586 POR2X1_29/A POR2X1_816/A 0.06fF
C22587 POR2X1_388/m4_208_n4# PAND2X1_93/B 0.08fF
C22588 POR2X1_96/A POR2X1_297/a_16_28# 0.00fF
C22589 POR2X1_49/Y PAND2X1_454/CTRL2 0.01fF
C22590 POR2X1_43/B POR2X1_309/a_16_28# 0.02fF
C22591 POR2X1_188/A PAND2X1_48/B 0.03fF
C22592 POR2X1_29/A D_INPUT_1 0.36fF
C22593 PAND2X1_807/B PAND2X1_354/O 0.02fF
C22594 PAND2X1_39/CTRL2 PAND2X1_69/A 0.00fF
C22595 POR2X1_66/B PAND2X1_625/CTRL 0.01fF
C22596 PAND2X1_55/Y POR2X1_750/B 0.17fF
C22597 POR2X1_251/CTRL2 PAND2X1_190/Y 0.01fF
C22598 PAND2X1_217/B PAND2X1_493/Y 0.05fF
C22599 POR2X1_567/B PAND2X1_173/a_16_344# 0.06fF
C22600 POR2X1_856/B PAND2X1_173/O 0.02fF
C22601 PAND2X1_659/A POR2X1_494/Y 0.12fF
C22602 POR2X1_121/B POR2X1_777/a_16_28# 0.03fF
C22603 POR2X1_65/A POR2X1_314/CTRL 0.01fF
C22604 PAND2X1_94/A PAND2X1_612/B 0.03fF
C22605 POR2X1_46/Y POR2X1_5/Y 0.08fF
C22606 POR2X1_502/A POR2X1_480/A 0.07fF
C22607 POR2X1_717/a_16_28# POR2X1_558/B -0.00fF
C22608 POR2X1_119/Y PAND2X1_464/B 0.07fF
C22609 POR2X1_49/Y POR2X1_42/Y 0.95fF
C22610 POR2X1_93/Y PAND2X1_510/B 0.02fF
C22611 POR2X1_833/A POR2X1_624/Y 0.11fF
C22612 INPUT_1 PAND2X1_340/B 0.03fF
C22613 PAND2X1_214/O PAND2X1_656/A 0.05fF
C22614 POR2X1_487/Y PAND2X1_357/Y 0.00fF
C22615 PAND2X1_735/Y VDD 0.08fF
C22616 POR2X1_43/B PAND2X1_390/Y 0.03fF
C22617 PAND2X1_55/Y PAND2X1_13/O 0.04fF
C22618 POR2X1_458/Y POR2X1_343/O 0.01fF
C22619 PAND2X1_180/a_76_28# PAND2X1_182/A 0.01fF
C22620 PAND2X1_660/O POR2X1_413/A 0.02fF
C22621 PAND2X1_58/A POR2X1_550/CTRL 0.01fF
C22622 POR2X1_93/A POR2X1_268/a_16_28# 0.05fF
C22623 POR2X1_102/Y POR2X1_38/Y 4.82fF
C22624 POR2X1_499/A POR2X1_294/A 0.05fF
C22625 POR2X1_417/Y PAND2X1_457/CTRL 0.01fF
C22626 PAND2X1_90/Y POR2X1_149/Y 0.01fF
C22627 PAND2X1_23/Y POR2X1_555/A 0.01fF
C22628 POR2X1_13/A POR2X1_13/O 0.12fF
C22629 POR2X1_634/CTRL PAND2X1_32/B 0.01fF
C22630 POR2X1_455/O POR2X1_193/A 0.07fF
C22631 POR2X1_24/Y POR2X1_394/A 0.27fF
C22632 POR2X1_509/A POR2X1_509/B 0.00fF
C22633 POR2X1_114/B POR2X1_288/A 0.03fF
C22634 POR2X1_264/Y POR2X1_650/A 0.02fF
C22635 POR2X1_362/B POR2X1_733/A 0.05fF
C22636 PAND2X1_675/A PAND2X1_562/B 0.07fF
C22637 PAND2X1_230/a_76_28# PAND2X1_32/B 0.07fF
C22638 POR2X1_278/Y POR2X1_96/A 0.18fF
C22639 POR2X1_673/CTRL POR2X1_38/B 0.01fF
C22640 PAND2X1_319/B POR2X1_60/A 0.10fF
C22641 PAND2X1_479/O POR2X1_599/A 0.31fF
C22642 POR2X1_422/Y POR2X1_408/Y 0.05fF
C22643 POR2X1_65/A PAND2X1_794/B 0.03fF
C22644 POR2X1_116/A POR2X1_362/CTRL 0.00fF
C22645 POR2X1_72/B POR2X1_90/Y 1.81fF
C22646 PAND2X1_41/CTRL POR2X1_294/A 0.01fF
C22647 PAND2X1_825/CTRL POR2X1_296/B 0.00fF
C22648 POR2X1_612/Y POR2X1_4/CTRL 0.04fF
C22649 POR2X1_447/B PAND2X1_43/CTRL2 0.04fF
C22650 POR2X1_423/Y PAND2X1_702/CTRL2 0.01fF
C22651 POR2X1_856/B POR2X1_456/B 0.06fF
C22652 PAND2X1_192/Y PAND2X1_357/Y 0.03fF
C22653 POR2X1_407/A POR2X1_287/B 0.03fF
C22654 PAND2X1_859/B VDD 0.96fF
C22655 POR2X1_52/A PAND2X1_480/B 0.03fF
C22656 POR2X1_16/A PAND2X1_561/CTRL2 0.12fF
C22657 PAND2X1_493/Y VDD 0.03fF
C22658 POR2X1_40/Y POR2X1_511/CTRL2 0.01fF
C22659 POR2X1_68/A POR2X1_5/Y 11.06fF
C22660 POR2X1_254/Y POR2X1_193/A 0.09fF
C22661 POR2X1_96/A POR2X1_829/A 0.03fF
C22662 POR2X1_254/Y POR2X1_579/Y 0.03fF
C22663 PAND2X1_218/CTRL2 VDD 0.00fF
C22664 POR2X1_558/CTRL2 INPUT_0 0.06fF
C22665 POR2X1_111/Y POR2X1_48/A 0.02fF
C22666 PAND2X1_854/O VDD 0.00fF
C22667 PAND2X1_717/A POR2X1_77/Y 0.03fF
C22668 PAND2X1_23/Y POR2X1_544/A 0.01fF
C22669 PAND2X1_180/O PAND2X1_566/Y 0.00fF
C22670 PAND2X1_48/B POR2X1_859/A 0.05fF
C22671 POR2X1_52/A POR2X1_754/A 0.03fF
C22672 PAND2X1_174/O VDD 0.00fF
C22673 POR2X1_580/CTRL2 D_GATE_741 0.02fF
C22674 POR2X1_252/Y POR2X1_257/A 0.12fF
C22675 PAND2X1_90/A POR2X1_502/A 0.05fF
C22676 PAND2X1_89/CTRL2 POR2X1_785/A 0.10fF
C22677 POR2X1_120/CTRL POR2X1_712/Y 0.03fF
C22678 POR2X1_61/Y POR2X1_219/B 0.77fF
C22679 PAND2X1_39/B POR2X1_4/Y 0.03fF
C22680 D_GATE_222 VDD 0.61fF
C22681 POR2X1_502/A POR2X1_756/a_56_344# 0.00fF
C22682 PAND2X1_793/Y POR2X1_488/Y 0.02fF
C22683 POR2X1_650/O POR2X1_773/B 0.29fF
C22684 POR2X1_49/Y PAND2X1_99/Y 0.02fF
C22685 POR2X1_159/O PAND2X1_63/B 0.01fF
C22686 PAND2X1_865/Y POR2X1_679/A 0.07fF
C22687 PAND2X1_675/A POR2X1_13/A 0.03fF
C22688 PAND2X1_65/Y PAND2X1_88/Y 0.03fF
C22689 POR2X1_23/Y PAND2X1_156/A 0.23fF
C22690 POR2X1_146/m4_208_n4# POR2X1_669/B 0.01fF
C22691 POR2X1_140/A VDD 0.00fF
C22692 PAND2X1_553/B POR2X1_42/Y 0.03fF
C22693 PAND2X1_41/B POR2X1_711/m4_208_n4# 0.07fF
C22694 POR2X1_13/A PAND2X1_469/B 0.03fF
C22695 PAND2X1_738/Y PAND2X1_357/Y 0.05fF
C22696 POR2X1_8/Y POR2X1_104/CTRL2 0.01fF
C22697 POR2X1_174/A POR2X1_353/A 0.12fF
C22698 INPUT_1 POR2X1_102/Y 0.06fF
C22699 POR2X1_79/Y PAND2X1_730/O 0.02fF
C22700 POR2X1_322/Y POR2X1_65/A 0.00fF
C22701 PAND2X1_205/A PAND2X1_716/B 0.00fF
C22702 POR2X1_130/A POR2X1_778/B 0.23fF
C22703 POR2X1_655/Y POR2X1_796/A 0.01fF
C22704 PAND2X1_491/CTRL INPUT_0 0.05fF
C22705 POR2X1_817/Y POR2X1_817/A 0.04fF
C22706 PAND2X1_682/O POR2X1_220/Y 0.01fF
C22707 POR2X1_254/Y POR2X1_614/A 0.08fF
C22708 PAND2X1_764/O PAND2X1_41/B 0.03fF
C22709 POR2X1_465/B POR2X1_222/Y 0.03fF
C22710 POR2X1_546/A POR2X1_816/A 0.03fF
C22711 POR2X1_516/A POR2X1_423/Y 0.61fF
C22712 POR2X1_23/Y POR2X1_373/CTRL 0.01fF
C22713 PAND2X1_28/O POR2X1_750/B 0.03fF
C22714 D_INPUT_1 POR2X1_546/A 3.56fF
C22715 PAND2X1_778/CTRL2 POR2X1_387/Y 0.06fF
C22716 POR2X1_65/A POR2X1_107/Y 0.04fF
C22717 POR2X1_347/A PAND2X1_20/A 0.03fF
C22718 POR2X1_198/CTRL POR2X1_198/B 0.01fF
C22719 POR2X1_16/A PAND2X1_78/O 0.06fF
C22720 PAND2X1_434/CTRL PAND2X1_390/Y 0.01fF
C22721 POR2X1_264/Y POR2X1_294/B 0.09fF
C22722 POR2X1_627/a_16_28# POR2X1_93/A 0.03fF
C22723 POR2X1_78/A PAND2X1_142/CTRL 0.01fF
C22724 POR2X1_193/Y POR2X1_222/A 0.02fF
C22725 PAND2X1_770/a_16_344# POR2X1_73/Y 0.02fF
C22726 PAND2X1_665/CTRL POR2X1_260/B 0.01fF
C22727 POR2X1_542/B PAND2X1_57/B 0.03fF
C22728 PAND2X1_777/CTRL2 PAND2X1_784/A 0.01fF
C22729 POR2X1_102/Y POR2X1_153/Y 0.39fF
C22730 INPUT_0 POR2X1_591/Y 0.03fF
C22731 PAND2X1_6/Y PAND2X1_183/O 0.02fF
C22732 POR2X1_495/Y PAND2X1_658/B 0.03fF
C22733 POR2X1_43/B POR2X1_277/a_56_344# 0.03fF
C22734 PAND2X1_73/Y PAND2X1_527/CTRL 0.02fF
C22735 POR2X1_557/A PAND2X1_42/CTRL 0.00fF
C22736 POR2X1_72/B PAND2X1_732/A 0.03fF
C22737 POR2X1_56/B PAND2X1_651/Y 0.03fF
C22738 POR2X1_334/CTRL2 POR2X1_814/B 0.01fF
C22739 POR2X1_96/A POR2X1_761/Y 0.03fF
C22740 POR2X1_404/Y POR2X1_576/Y 0.03fF
C22741 POR2X1_96/A PAND2X1_359/a_76_28# 0.02fF
C22742 INPUT_1 PAND2X1_23/O 0.16fF
C22743 POR2X1_29/A POR2X1_620/B 0.03fF
C22744 PAND2X1_661/a_16_344# PAND2X1_653/Y 0.01fF
C22745 POR2X1_347/A PAND2X1_96/CTRL 0.01fF
C22746 POR2X1_222/Y D_GATE_741 0.07fF
C22747 POR2X1_271/CTRL2 POR2X1_39/B 0.03fF
C22748 POR2X1_308/CTRL POR2X1_725/Y 0.04fF
C22749 POR2X1_592/Y PAND2X1_93/B 0.00fF
C22750 POR2X1_480/A POR2X1_799/CTRL 0.02fF
C22751 PAND2X1_436/A POR2X1_153/Y 0.09fF
C22752 PAND2X1_140/A PAND2X1_738/Y 0.05fF
C22753 POR2X1_332/B POR2X1_228/Y 0.03fF
C22754 POR2X1_356/A POR2X1_210/Y 0.07fF
C22755 PAND2X1_785/O POR2X1_7/B 0.17fF
C22756 POR2X1_131/a_16_28# PAND2X1_137/Y 0.11fF
C22757 POR2X1_722/Y POR2X1_513/CTRL 0.01fF
C22758 PAND2X1_794/B PAND2X1_190/Y 0.05fF
C22759 POR2X1_579/Y POR2X1_341/Y 0.03fF
C22760 POR2X1_368/O POR2X1_7/A 0.03fF
C22761 POR2X1_327/Y POR2X1_453/a_76_344# 0.03fF
C22762 POR2X1_730/Y PAND2X1_65/B 0.03fF
C22763 POR2X1_619/A POR2X1_7/B 0.03fF
C22764 POR2X1_514/Y POR2X1_139/O 0.16fF
C22765 POR2X1_278/Y POR2X1_7/A 0.05fF
C22766 POR2X1_99/B POR2X1_555/B 0.00fF
C22767 PAND2X1_48/B PAND2X1_59/O 0.01fF
C22768 PAND2X1_309/a_16_344# POR2X1_335/B 0.01fF
C22769 POR2X1_713/A INPUT_1 0.01fF
C22770 POR2X1_481/Y PAND2X1_555/O 0.01fF
C22771 POR2X1_198/B POR2X1_532/A 0.21fF
C22772 PAND2X1_569/B VDD 0.00fF
C22773 POR2X1_566/A POR2X1_854/B 0.10fF
C22774 POR2X1_110/Y PAND2X1_465/CTRL2 0.09fF
C22775 VDD POR2X1_158/B 0.55fF
C22776 POR2X1_346/B POR2X1_403/Y 0.03fF
C22777 PAND2X1_784/CTRL2 POR2X1_387/Y 0.05fF
C22778 POR2X1_346/O PAND2X1_23/Y 0.00fF
C22779 D_GATE_222 PAND2X1_32/B 0.12fF
C22780 PAND2X1_46/CTRL2 POR2X1_294/A 0.00fF
C22781 PAND2X1_20/A POR2X1_4/Y 0.03fF
C22782 POR2X1_219/B POR2X1_35/Y 0.00fF
C22783 POR2X1_8/Y POR2X1_58/O 0.01fF
C22784 POR2X1_647/CTRL PAND2X1_52/B 0.01fF
C22785 POR2X1_687/A PAND2X1_760/O 0.04fF
C22786 POR2X1_426/CTRL2 POR2X1_425/Y 0.01fF
C22787 POR2X1_741/Y POR2X1_702/CTRL2 0.01fF
C22788 POR2X1_376/B POR2X1_373/Y 0.03fF
C22789 PAND2X1_676/a_16_344# POR2X1_599/A 0.02fF
C22790 POR2X1_99/B POR2X1_330/Y 0.03fF
C22791 POR2X1_614/A POR2X1_341/Y 0.01fF
C22792 PAND2X1_602/Y POR2X1_757/O 0.01fF
C22793 POR2X1_315/CTRL POR2X1_91/Y 0.01fF
C22794 INPUT_7 PAND2X1_18/B 0.03fF
C22795 D_INPUT_1 POR2X1_500/Y 0.03fF
C22796 POR2X1_82/a_16_28# INPUT_1 0.03fF
C22797 POR2X1_16/A POR2X1_234/Y 0.01fF
C22798 POR2X1_662/Y POR2X1_725/Y 0.03fF
C22799 PAND2X1_632/B POR2X1_7/B 0.05fF
C22800 POR2X1_294/B PAND2X1_528/CTRL 0.08fF
C22801 PAND2X1_56/Y POR2X1_702/O 0.02fF
C22802 POR2X1_41/B POR2X1_385/a_56_344# 0.00fF
C22803 POR2X1_371/CTRL POR2X1_5/Y 0.01fF
C22804 POR2X1_379/m4_208_n4# PAND2X1_18/m4_208_n4# 0.13fF
C22805 D_INPUT_0 POR2X1_522/O 0.06fF
C22806 POR2X1_544/Y VDD 0.13fF
C22807 PAND2X1_385/a_76_28# PAND2X1_60/B 0.01fF
C22808 POR2X1_20/Y POR2X1_380/Y 0.95fF
C22809 PAND2X1_76/Y PAND2X1_716/B 0.15fF
C22810 POR2X1_702/CTRL2 PAND2X1_32/B 0.03fF
C22811 POR2X1_322/Y PAND2X1_565/O 0.00fF
C22812 POR2X1_322/O PAND2X1_569/B 0.01fF
C22813 POR2X1_814/B POR2X1_4/Y 0.07fF
C22814 PAND2X1_288/O PAND2X1_221/Y 0.09fF
C22815 PAND2X1_25/CTRL2 PAND2X1_72/A 0.10fF
C22816 D_INPUT_7 PAND2X1_425/Y 0.03fF
C22817 POR2X1_300/a_76_344# PAND2X1_349/A 0.00fF
C22818 PAND2X1_41/B PAND2X1_759/CTRL 0.01fF
C22819 PAND2X1_6/A POR2X1_283/A 0.17fF
C22820 POR2X1_855/B POR2X1_796/CTRL 0.01fF
C22821 POR2X1_210/CTRL PAND2X1_52/B 0.01fF
C22822 POR2X1_210/Y POR2X1_220/A 1.04fF
C22823 POR2X1_108/CTRL2 POR2X1_142/Y 0.06fF
C22824 POR2X1_356/A POR2X1_782/B 0.04fF
C22825 POR2X1_552/O VDD 0.00fF
C22826 POR2X1_416/B POR2X1_667/A 0.09fF
C22827 POR2X1_417/O POR2X1_387/Y 0.06fF
C22828 POR2X1_45/Y PAND2X1_737/B 0.03fF
C22829 POR2X1_41/O POR2X1_42/Y 0.01fF
C22830 POR2X1_416/B POR2X1_607/A 0.01fF
C22831 PAND2X1_69/A PAND2X1_63/B 0.10fF
C22832 PAND2X1_39/B POR2X1_458/Y 0.02fF
C22833 POR2X1_390/B POR2X1_723/B 0.00fF
C22834 POR2X1_134/Y POR2X1_103/Y 0.00fF
C22835 PAND2X1_500/CTRL POR2X1_497/Y 0.01fF
C22836 POR2X1_498/Y PAND2X1_332/Y 0.03fF
C22837 POR2X1_41/Y POR2X1_236/Y 0.03fF
C22838 INPUT_4 PAND2X1_18/B 0.07fF
C22839 POR2X1_405/Y PAND2X1_48/A 0.04fF
C22840 POR2X1_416/B POR2X1_255/O 0.03fF
C22841 PAND2X1_48/B PAND2X1_484/O 0.17fF
C22842 POR2X1_532/A POR2X1_520/CTRL2 0.01fF
C22843 POR2X1_567/A POR2X1_653/a_76_344# 0.01fF
C22844 PAND2X1_727/a_76_28# POR2X1_152/A 0.01fF
C22845 POR2X1_784/A PAND2X1_48/A 3.69fF
C22846 PAND2X1_349/A POR2X1_91/Y 0.03fF
C22847 POR2X1_334/B POR2X1_334/A 0.02fF
C22848 POR2X1_68/B POR2X1_520/O 0.02fF
C22849 PAND2X1_602/Y POR2X1_394/A 0.07fF
C22850 PAND2X1_264/O POR2X1_73/Y 0.05fF
C22851 POR2X1_92/m4_208_n4# POR2X1_38/Y 0.01fF
C22852 POR2X1_661/CTRL2 POR2X1_711/Y 0.05fF
C22853 POR2X1_541/m4_208_n4# POR2X1_366/A 0.12fF
C22854 POR2X1_804/A POR2X1_260/A 0.05fF
C22855 POR2X1_538/A POR2X1_228/Y 0.00fF
C22856 PAND2X1_555/Y PAND2X1_346/Y 0.10fF
C22857 POR2X1_405/O PAND2X1_52/B 0.09fF
C22858 POR2X1_316/Y VDD 0.49fF
C22859 POR2X1_499/A POR2X1_116/A 0.03fF
C22860 POR2X1_68/B POR2X1_768/CTRL2 0.03fF
C22861 POR2X1_394/A PAND2X1_547/O 0.02fF
C22862 PAND2X1_798/Y VDD 0.72fF
C22863 POR2X1_118/CTRL POR2X1_153/Y 0.06fF
C22864 POR2X1_270/O POR2X1_456/B 0.01fF
C22865 POR2X1_851/a_16_28# POR2X1_733/A 0.09fF
C22866 PAND2X1_7/CTRL2 POR2X1_99/B 0.00fF
C22867 POR2X1_493/O POR2X1_773/B 0.01fF
C22868 PAND2X1_23/Y PAND2X1_396/CTRL 0.00fF
C22869 POR2X1_614/A POR2X1_370/CTRL 0.01fF
C22870 POR2X1_68/B PAND2X1_531/CTRL2 0.01fF
C22871 PAND2X1_730/O PAND2X1_730/A 0.02fF
C22872 POR2X1_540/Y PAND2X1_178/O 0.02fF
C22873 PAND2X1_788/O POR2X1_533/Y -0.00fF
C22874 PAND2X1_33/CTRL2 POR2X1_24/Y 0.01fF
C22875 POR2X1_383/A PAND2X1_298/CTRL 0.05fF
C22876 POR2X1_707/B POR2X1_451/A 0.02fF
C22877 POR2X1_513/B PAND2X1_304/a_76_28# 0.04fF
C22878 POR2X1_679/a_56_344# POR2X1_679/A 0.00fF
C22879 PAND2X1_838/B PAND2X1_838/O 0.02fF
C22880 PAND2X1_388/Y PAND2X1_348/A 0.07fF
C22881 POR2X1_98/A POR2X1_590/A 0.03fF
C22882 PAND2X1_687/CTRL2 PAND2X1_643/Y 0.03fF
C22883 PAND2X1_90/Y POR2X1_568/A 4.86fF
C22884 POR2X1_38/Y PAND2X1_120/a_16_344# 0.02fF
C22885 POR2X1_116/A POR2X1_76/A 0.03fF
C22886 POR2X1_532/A POR2X1_342/CTRL2 0.01fF
C22887 POR2X1_557/A PAND2X1_94/A 0.03fF
C22888 POR2X1_41/B POR2X1_77/Y 0.63fF
C22889 POR2X1_735/CTRL2 POR2X1_318/A 0.05fF
C22890 PAND2X1_678/a_76_28# POR2X1_257/A 0.02fF
C22891 POR2X1_41/B POR2X1_85/Y 0.02fF
C22892 PAND2X1_94/A PAND2X1_184/O 0.04fF
C22893 POR2X1_376/B POR2X1_386/Y 0.01fF
C22894 POR2X1_343/Y POR2X1_294/B 0.05fF
C22895 POR2X1_65/A PAND2X1_221/Y 0.01fF
C22896 POR2X1_333/Y POR2X1_502/CTRL2 0.00fF
C22897 POR2X1_244/Y POR2X1_456/B 0.03fF
C22898 POR2X1_234/A POR2X1_236/Y 0.01fF
C22899 PAND2X1_832/O POR2X1_677/Y 0.00fF
C22900 POR2X1_356/A POR2X1_181/Y 0.03fF
C22901 POR2X1_304/CTRL POR2X1_90/Y 0.01fF
C22902 POR2X1_661/A POR2X1_830/A 0.07fF
C22903 POR2X1_396/CTRL POR2X1_39/B 0.01fF
C22904 PAND2X1_6/Y POR2X1_632/Y 0.03fF
C22905 PAND2X1_272/CTRL POR2X1_556/A 0.00fF
C22906 POR2X1_315/Y PAND2X1_716/B 0.97fF
C22907 POR2X1_119/Y POR2X1_283/A 0.07fF
C22908 POR2X1_65/A POR2X1_250/a_16_28# 0.03fF
C22909 POR2X1_554/B POR2X1_657/CTRL 0.01fF
C22910 POR2X1_119/Y PAND2X1_121/CTRL 0.02fF
C22911 POR2X1_508/B POR2X1_383/A 0.00fF
C22912 POR2X1_329/A POR2X1_594/a_16_28# 0.03fF
C22913 POR2X1_38/Y POR2X1_761/A 0.02fF
C22914 POR2X1_833/A POR2X1_186/B 0.01fF
C22915 PAND2X1_189/O POR2X1_353/A 0.00fF
C22916 PAND2X1_631/A PAND2X1_549/B 0.12fF
C22917 PAND2X1_640/O POR2X1_77/Y 0.15fF
C22918 PAND2X1_65/B PAND2X1_255/O 0.01fF
C22919 POR2X1_270/Y POR2X1_659/A 0.00fF
C22920 POR2X1_440/CTRL2 VDD -0.00fF
C22921 PAND2X1_20/A POR2X1_296/O 0.01fF
C22922 POR2X1_537/Y POR2X1_858/B 0.02fF
C22923 INPUT_3 POR2X1_29/A 0.09fF
C22924 POR2X1_20/B PAND2X1_721/B 0.08fF
C22925 POR2X1_364/A POR2X1_168/A 0.01fF
C22926 PAND2X1_157/CTRL2 PAND2X1_3/B 0.00fF
C22927 PAND2X1_20/A POR2X1_78/Y 0.04fF
C22928 PAND2X1_6/Y PAND2X1_52/B 5.10fF
C22929 PAND2X1_404/CTRL POR2X1_411/B 0.11fF
C22930 POR2X1_257/A POR2X1_67/A 0.03fF
C22931 PAND2X1_6/O POR2X1_294/A 0.03fF
C22932 POR2X1_52/A POR2X1_386/Y 0.08fF
C22933 PAND2X1_258/O POR2X1_454/A 0.03fF
C22934 POR2X1_458/Y POR2X1_325/A 0.03fF
C22935 POR2X1_39/B PAND2X1_149/A 0.05fF
C22936 POR2X1_87/O POR2X1_38/B 0.02fF
C22937 POR2X1_456/B POR2X1_703/a_16_28# 0.03fF
C22938 POR2X1_492/Y PAND2X1_717/Y 0.01fF
C22939 POR2X1_750/Y PAND2X1_526/CTRL2 0.14fF
C22940 PAND2X1_826/O POR2X1_296/B 0.32fF
C22941 PAND2X1_464/CTRL POR2X1_417/Y 0.01fF
C22942 POR2X1_841/CTRL2 POR2X1_330/Y 0.32fF
C22943 POR2X1_343/Y PAND2X1_111/B 0.05fF
C22944 PAND2X1_1/CTRL D_INPUT_4 0.01fF
C22945 PAND2X1_859/A PAND2X1_227/O 0.02fF
C22946 POR2X1_287/B POR2X1_287/A 0.00fF
C22947 PAND2X1_39/B POR2X1_400/O 0.01fF
C22948 PAND2X1_93/B POR2X1_269/CTRL 0.01fF
C22949 POR2X1_416/B POR2X1_245/Y 0.00fF
C22950 POR2X1_66/B D_INPUT_5 0.03fF
C22951 POR2X1_118/Y POR2X1_32/A 0.02fF
C22952 PAND2X1_485/CTRL2 POR2X1_590/A 0.01fF
C22953 POR2X1_102/Y POR2X1_248/A 0.02fF
C22954 POR2X1_707/B PAND2X1_762/CTRL 0.01fF
C22955 POR2X1_265/CTRL POR2X1_667/A 0.01fF
C22956 PAND2X1_86/O INPUT_0 0.02fF
C22957 PAND2X1_20/A POR2X1_34/O 0.01fF
C22958 PAND2X1_175/B POR2X1_173/CTRL2 0.01fF
C22959 POR2X1_383/A POR2X1_325/B 0.03fF
C22960 POR2X1_110/Y POR2X1_110/O 0.01fF
C22961 POR2X1_669/B POR2X1_626/CTRL 0.04fF
C22962 POR2X1_634/A POR2X1_862/A 0.10fF
C22963 POR2X1_257/A PAND2X1_161/a_76_28# 0.01fF
C22964 POR2X1_504/Y POR2X1_628/Y 0.06fF
C22965 POR2X1_294/Y POR2X1_296/B 0.09fF
C22966 POR2X1_54/Y PAND2X1_526/CTRL 0.29fF
C22967 POR2X1_411/B PAND2X1_473/B 0.09fF
C22968 PAND2X1_58/A PAND2X1_3/A 0.01fF
C22969 PAND2X1_659/Y PAND2X1_737/O 0.03fF
C22970 PAND2X1_698/CTRL2 PAND2X1_52/B 0.16fF
C22971 POR2X1_441/Y PAND2X1_544/a_16_344# 0.01fF
C22972 PAND2X1_308/Y POR2X1_77/Y 0.03fF
C22973 POR2X1_260/B POR2X1_389/Y 0.03fF
C22974 POR2X1_842/a_16_28# POR2X1_830/Y 0.02fF
C22975 POR2X1_602/B PAND2X1_93/B 0.03fF
C22976 POR2X1_416/B PAND2X1_507/CTRL 0.00fF
C22977 POR2X1_120/CTRL PAND2X1_39/B 0.01fF
C22978 POR2X1_78/A POR2X1_29/A 0.15fF
C22979 PAND2X1_652/A POR2X1_329/A 0.28fF
C22980 POR2X1_32/A PAND2X1_573/B 0.01fF
C22981 PAND2X1_65/B PAND2X1_26/A 0.07fF
C22982 PAND2X1_694/O PAND2X1_425/Y 0.01fF
C22983 POR2X1_292/O POR2X1_90/Y 0.01fF
C22984 PAND2X1_508/B PAND2X1_506/Y 0.14fF
C22985 POR2X1_648/CTRL VDD 0.00fF
C22986 POR2X1_49/Y PAND2X1_576/B 0.03fF
C22987 POR2X1_9/Y POR2X1_38/Y 0.13fF
C22988 POR2X1_54/Y VDD 5.90fF
C22989 POR2X1_68/A PAND2X1_617/CTRL2 0.03fF
C22990 PAND2X1_73/Y POR2X1_634/A 0.13fF
C22991 POR2X1_777/B POR2X1_218/Y 0.10fF
C22992 POR2X1_774/Y POR2X1_636/B 0.00fF
C22993 PAND2X1_5/CTRL POR2X1_612/A 0.01fF
C22994 POR2X1_159/O POR2X1_32/A 0.01fF
C22995 POR2X1_119/Y POR2X1_518/a_16_28# 0.07fF
C22996 POR2X1_655/CTRL POR2X1_307/A 0.00fF
C22997 POR2X1_122/Y PAND2X1_852/A 0.04fF
C22998 POR2X1_98/O PAND2X1_41/B 0.01fF
C22999 PAND2X1_860/A PAND2X1_175/CTRL 0.01fF
C23000 POR2X1_834/a_76_344# POR2X1_330/Y 0.03fF
C23001 POR2X1_298/O VDD -0.00fF
C23002 PAND2X1_266/CTRL POR2X1_73/Y 0.02fF
C23003 PAND2X1_404/Y PAND2X1_84/a_76_28# 0.01fF
C23004 PAND2X1_48/B PAND2X1_416/CTRL 0.01fF
C23005 POR2X1_750/B POR2X1_375/Y 0.01fF
C23006 POR2X1_624/Y POR2X1_294/B 0.05fF
C23007 POR2X1_65/A POR2X1_83/B 1.45fF
C23008 POR2X1_20/B POR2X1_56/Y 0.48fF
C23009 POR2X1_94/CTRL2 POR2X1_24/Y 0.01fF
C23010 POR2X1_644/B VDD 0.10fF
C23011 PAND2X1_39/B PAND2X1_744/CTRL2 0.02fF
C23012 POR2X1_688/CTRL POR2X1_532/A 0.01fF
C23013 POR2X1_78/A POR2X1_213/B 0.01fF
C23014 POR2X1_96/A POR2X1_420/CTRL2 0.01fF
C23015 POR2X1_346/A VDD 0.00fF
C23016 PAND2X1_770/a_76_28# PAND2X1_771/Y 0.02fF
C23017 INPUT_1 POR2X1_9/Y 0.23fF
C23018 PAND2X1_408/O D_INPUT_6 -0.00fF
C23019 PAND2X1_80/CTRL POR2X1_296/B 0.00fF
C23020 POR2X1_648/Y POR2X1_407/CTRL2 0.01fF
C23021 PAND2X1_58/A POR2X1_5/Y 0.03fF
C23022 PAND2X1_169/Y PAND2X1_211/A 0.03fF
C23023 POR2X1_65/A POR2X1_829/O 0.01fF
C23024 POR2X1_814/B PAND2X1_616/CTRL 0.01fF
C23025 POR2X1_120/CTRL POR2X1_805/Y 0.03fF
C23026 POR2X1_60/A PAND2X1_333/a_16_344# 0.02fF
C23027 POR2X1_306/Y PAND2X1_512/a_16_344# 0.05fF
C23028 PAND2X1_824/B PAND2X1_234/CTRL2 0.01fF
C23029 POR2X1_677/Y POR2X1_153/Y 0.03fF
C23030 PAND2X1_57/O POR2X1_590/A 0.15fF
C23031 POR2X1_686/A POR2X1_750/B 0.05fF
C23032 POR2X1_114/B POR2X1_475/a_16_28# 0.00fF
C23033 POR2X1_130/A PAND2X1_73/Y 0.38fF
C23034 D_INPUT_0 POR2X1_232/CTRL2 0.03fF
C23035 PAND2X1_57/B POR2X1_770/B 0.03fF
C23036 PAND2X1_494/CTRL2 POR2X1_260/B 0.01fF
C23037 POR2X1_60/A PAND2X1_687/Y 0.01fF
C23038 PAND2X1_675/A POR2X1_437/O 0.18fF
C23039 POR2X1_432/a_16_28# POR2X1_236/Y 0.02fF
C23040 POR2X1_669/Y PAND2X1_720/CTRL2 0.01fF
C23041 POR2X1_566/A PAND2X1_73/Y 0.05fF
C23042 POR2X1_54/Y PAND2X1_32/B 0.03fF
C23043 POR2X1_452/Y POR2X1_685/B 0.16fF
C23044 POR2X1_730/Y POR2X1_814/A 0.03fF
C23045 POR2X1_52/A POR2X1_484/O 0.16fF
C23046 PAND2X1_803/Y POR2X1_20/B 0.02fF
C23047 POR2X1_13/A POR2X1_423/O 0.18fF
C23048 POR2X1_676/O PAND2X1_69/A 0.04fF
C23049 PAND2X1_832/a_16_344# POR2X1_423/Y 0.02fF
C23050 POR2X1_263/Y POR2X1_55/Y 0.03fF
C23051 POR2X1_538/CTRL POR2X1_270/Y 0.00fF
C23052 POR2X1_311/Y POR2X1_278/Y 0.03fF
C23053 PAND2X1_402/O POR2X1_5/Y 0.05fF
C23054 PAND2X1_276/a_76_28# POR2X1_271/Y 0.00fF
C23055 POR2X1_48/A PAND2X1_649/CTRL 0.01fF
C23056 POR2X1_66/A PAND2X1_385/O 0.04fF
C23057 POR2X1_97/A POR2X1_785/A 0.03fF
C23058 PAND2X1_93/B POR2X1_712/Y 0.07fF
C23059 POR2X1_423/CTRL POR2X1_293/Y 0.01fF
C23060 POR2X1_484/a_16_28# POR2X1_763/Y 0.07fF
C23061 POR2X1_636/a_56_344# POR2X1_636/A 0.00fF
C23062 POR2X1_753/Y POR2X1_615/Y 0.02fF
C23063 POR2X1_862/B POR2X1_480/A 0.03fF
C23064 POR2X1_72/B INPUT_0 10.38fF
C23065 POR2X1_78/B POR2X1_403/CTRL2 0.01fF
C23066 POR2X1_624/Y PAND2X1_111/B 0.01fF
C23067 POR2X1_644/a_56_344# POR2X1_407/Y 0.00fF
C23068 PAND2X1_570/a_16_344# PAND2X1_771/Y 0.04fF
C23069 POR2X1_673/A POR2X1_814/B 0.03fF
C23070 POR2X1_446/B PAND2X1_60/B 0.03fF
C23071 POR2X1_634/A PAND2X1_132/CTRL2 0.01fF
C23072 POR2X1_846/Y POR2X1_753/CTRL 0.01fF
C23073 PAND2X1_52/B POR2X1_212/B 0.03fF
C23074 PAND2X1_449/O PAND2X1_308/Y 0.02fF
C23075 POR2X1_260/B POR2X1_318/A 0.51fF
C23076 PAND2X1_676/CTRL PAND2X1_205/A 0.00fF
C23077 POR2X1_283/O PAND2X1_365/B 0.01fF
C23078 POR2X1_257/A PAND2X1_550/B 5.88fF
C23079 POR2X1_99/m4_208_n4# POR2X1_360/m4_208_n4# 0.05fF
C23080 PAND2X1_97/CTRL POR2X1_91/Y 0.01fF
C23081 PAND2X1_217/CTRL2 PAND2X1_576/B 0.01fF
C23082 POR2X1_275/CTRL2 PAND2X1_390/Y 0.01fF
C23083 POR2X1_830/CTRL2 POR2X1_733/A 0.03fF
C23084 POR2X1_706/A VDD -0.00fF
C23085 POR2X1_40/Y POR2X1_531/O 0.02fF
C23086 POR2X1_288/A POR2X1_405/Y 0.42fF
C23087 POR2X1_119/Y POR2X1_399/Y 0.17fF
C23088 POR2X1_840/B D_INPUT_0 0.23fF
C23089 POR2X1_260/B POR2X1_713/B 0.05fF
C23090 POR2X1_78/A POR2X1_712/Y 8.03fF
C23091 PAND2X1_73/Y POR2X1_844/B 0.05fF
C23092 POR2X1_98/CTRL POR2X1_68/B 0.07fF
C23093 PAND2X1_267/CTRL POR2X1_7/A 0.01fF
C23094 POR2X1_51/a_56_344# PAND2X1_635/Y 0.00fF
C23095 POR2X1_288/A POR2X1_784/A 0.03fF
C23096 PAND2X1_80/CTRL POR2X1_547/B 0.01fF
C23097 POR2X1_499/a_16_28# D_INPUT_1 0.02fF
C23098 PAND2X1_84/Y PAND2X1_558/a_16_344# 0.01fF
C23099 POR2X1_60/A PAND2X1_798/B 0.07fF
C23100 POR2X1_78/B POR2X1_608/CTRL 0.01fF
C23101 PAND2X1_615/O D_INPUT_0 0.05fF
C23102 PAND2X1_236/CTRL2 INPUT_0 0.00fF
C23103 PAND2X1_72/A PAND2X1_135/O 0.16fF
C23104 POR2X1_29/A POR2X1_748/CTRL2 0.01fF
C23105 PAND2X1_652/A PAND2X1_361/O 0.20fF
C23106 POR2X1_72/B PAND2X1_717/CTRL2 0.01fF
C23107 PAND2X1_449/Y POR2X1_102/Y 0.01fF
C23108 POR2X1_13/A PAND2X1_828/CTRL 0.01fF
C23109 PAND2X1_512/Y POR2X1_372/O 0.01fF
C23110 POR2X1_14/Y PAND2X1_6/A 0.10fF
C23111 POR2X1_48/A PAND2X1_149/A 0.76fF
C23112 POR2X1_230/O POR2X1_230/Y 0.01fF
C23113 PAND2X1_41/B POR2X1_579/Y 0.03fF
C23114 POR2X1_54/Y POR2X1_673/Y 0.03fF
C23115 PAND2X1_501/B VDD 0.17fF
C23116 POR2X1_150/Y PAND2X1_853/B 0.43fF
C23117 PAND2X1_721/CTRL2 POR2X1_7/B 0.03fF
C23118 POR2X1_625/CTRL POR2X1_754/A 0.01fF
C23119 POR2X1_83/B PAND2X1_565/O 0.01fF
C23120 POR2X1_614/A PAND2X1_427/CTRL2 0.03fF
C23121 PAND2X1_55/Y POR2X1_389/Y 0.07fF
C23122 PAND2X1_651/Y PAND2X1_573/B 0.03fF
C23123 PAND2X1_20/A POR2X1_462/B 0.03fF
C23124 PAND2X1_802/CTRL POR2X1_760/A 0.01fF
C23125 PAND2X1_41/B POR2X1_572/B 0.01fF
C23126 PAND2X1_73/Y POR2X1_573/A 0.00fF
C23127 PAND2X1_20/A D_INPUT_1 6.76fF
C23128 PAND2X1_466/CTRL2 PAND2X1_803/A 0.00fF
C23129 POR2X1_683/CTRL POR2X1_236/Y 0.03fF
C23130 POR2X1_221/Y POR2X1_186/Y 0.01fF
C23131 POR2X1_669/B POR2X1_619/Y 0.05fF
C23132 POR2X1_96/B POR2X1_48/A 0.03fF
C23133 POR2X1_16/A POR2X1_437/CTRL 0.02fF
C23134 POR2X1_179/O POR2X1_40/Y 0.18fF
C23135 PAND2X1_809/B PAND2X1_809/CTRL2 0.01fF
C23136 POR2X1_806/O PAND2X1_69/A 0.01fF
C23137 POR2X1_32/A POR2X1_91/Y 0.10fF
C23138 POR2X1_81/Y PAND2X1_499/Y 0.23fF
C23139 POR2X1_96/A PAND2X1_730/B 0.03fF
C23140 POR2X1_52/A PAND2X1_473/B 0.03fF
C23141 POR2X1_502/A POR2X1_459/CTRL2 0.01fF
C23142 POR2X1_114/B PAND2X1_299/CTRL2 0.01fF
C23143 PAND2X1_41/B POR2X1_545/A 0.03fF
C23144 POR2X1_814/B D_GATE_662 0.19fF
C23145 POR2X1_102/Y POR2X1_591/Y 0.03fF
C23146 POR2X1_334/B PAND2X1_262/a_16_344# 0.04fF
C23147 POR2X1_509/B POR2X1_35/Y 0.02fF
C23148 POR2X1_253/O PAND2X1_508/Y 0.00fF
C23149 PAND2X1_20/A POR2X1_724/A 0.03fF
C23150 PAND2X1_216/CTRL INPUT_0 0.01fF
C23151 POR2X1_330/Y POR2X1_112/Y 0.31fF
C23152 POR2X1_407/A POR2X1_647/Y 0.06fF
C23153 PAND2X1_724/CTRL2 PAND2X1_731/B 0.01fF
C23154 PAND2X1_88/CTRL POR2X1_38/B 0.01fF
C23155 PAND2X1_57/B POR2X1_722/Y 0.03fF
C23156 POR2X1_812/B POR2X1_812/A 0.02fF
C23157 PAND2X1_478/O PAND2X1_803/A 0.00fF
C23158 POR2X1_614/A PAND2X1_41/B 0.31fF
C23159 POR2X1_121/B PAND2X1_60/B 0.24fF
C23160 PAND2X1_23/Y POR2X1_663/O 0.01fF
C23161 POR2X1_646/Y POR2X1_725/Y 0.07fF
C23162 POR2X1_273/O POR2X1_129/Y 0.01fF
C23163 POR2X1_859/A POR2X1_790/O 0.35fF
C23164 POR2X1_260/B POR2X1_574/Y 0.03fF
C23165 PAND2X1_854/a_76_28# PAND2X1_805/A 0.01fF
C23166 POR2X1_241/B POR2X1_854/B 0.03fF
C23167 POR2X1_391/A PAND2X1_69/A 0.03fF
C23168 POR2X1_356/A POR2X1_570/CTRL 0.00fF
C23169 POR2X1_68/A PAND2X1_65/B 0.31fF
C23170 POR2X1_654/B PAND2X1_96/B 3.27fF
C23171 POR2X1_814/B D_INPUT_1 0.11fF
C23172 POR2X1_13/Y VDD 0.37fF
C23173 POR2X1_52/A POR2X1_627/Y 0.00fF
C23174 POR2X1_417/Y POR2X1_91/Y 0.03fF
C23175 POR2X1_812/A POR2X1_780/B 0.03fF
C23176 POR2X1_38/B PAND2X1_41/B 2.34fF
C23177 POR2X1_57/A PAND2X1_349/B 0.01fF
C23178 POR2X1_16/A PAND2X1_722/CTRL 0.00fF
C23179 POR2X1_78/B POR2X1_147/A 0.02fF
C23180 POR2X1_41/B PAND2X1_486/O 0.04fF
C23181 POR2X1_588/Y POR2X1_14/Y 0.05fF
C23182 PAND2X1_451/a_76_28# POR2X1_428/Y 0.01fF
C23183 POR2X1_40/Y PAND2X1_168/CTRL 0.01fF
C23184 POR2X1_37/Y PAND2X1_100/a_56_28# 0.00fF
C23185 POR2X1_69/A POR2X1_7/A 2.24fF
C23186 POR2X1_312/Y PAND2X1_182/a_76_28# 0.01fF
C23187 POR2X1_333/A POR2X1_738/A 0.13fF
C23188 POR2X1_14/Y POR2X1_419/CTRL2 0.00fF
C23189 POR2X1_231/CTRL2 POR2X1_785/A 0.00fF
C23190 POR2X1_717/CTRL POR2X1_814/B 0.01fF
C23191 PAND2X1_80/O PAND2X1_81/B 0.01fF
C23192 POR2X1_81/a_56_344# PAND2X1_510/B 0.00fF
C23193 POR2X1_330/Y POR2X1_162/Y 0.02fF
C23194 POR2X1_814/B POR2X1_724/A 0.12fF
C23195 PAND2X1_661/B PAND2X1_828/CTRL 0.01fF
C23196 PAND2X1_453/A POR2X1_419/CTRL2 0.01fF
C23197 PAND2X1_213/Y PAND2X1_738/B 0.03fF
C23198 POR2X1_41/B PAND2X1_742/B 0.03fF
C23199 PAND2X1_691/Y POR2X1_60/A 0.03fF
C23200 POR2X1_823/a_16_28# POR2X1_236/Y 0.03fF
C23201 INPUT_1 PAND2X1_638/B 0.01fF
C23202 PAND2X1_456/CTRL2 POR2X1_283/A 0.01fF
C23203 PAND2X1_449/O POR2X1_77/Y 0.08fF
C23204 PAND2X1_738/Y PAND2X1_182/CTRL2 0.06fF
C23205 POR2X1_688/Y POR2X1_691/A 0.02fF
C23206 POR2X1_78/B PAND2X1_69/A 0.29fF
C23207 POR2X1_650/A POR2X1_493/CTRL 0.02fF
C23208 POR2X1_353/Y POR2X1_353/CTRL2 0.01fF
C23209 POR2X1_57/A PAND2X1_139/a_76_28# 0.01fF
C23210 POR2X1_65/A PAND2X1_509/m4_208_n4# 0.08fF
C23211 POR2X1_294/B POR2X1_785/A 8.72fF
C23212 POR2X1_97/A POR2X1_186/B 0.06fF
C23213 POR2X1_202/B POR2X1_507/A 0.04fF
C23214 POR2X1_572/CTRL2 PAND2X1_32/B 0.01fF
C23215 POR2X1_376/B POR2X1_239/Y 0.05fF
C23216 POR2X1_628/O POR2X1_55/Y 0.01fF
C23217 POR2X1_347/B POR2X1_402/A 0.01fF
C23218 GATE_741 PAND2X1_362/O 0.05fF
C23219 POR2X1_822/Y VDD 0.01fF
C23220 POR2X1_280/Y POR2X1_279/Y 0.02fF
C23221 INPUT_2 POR2X1_609/A 0.01fF
C23222 POR2X1_23/Y POR2X1_171/Y 0.03fF
C23223 PAND2X1_40/a_16_344# PAND2X1_57/B 0.04fF
C23224 POR2X1_87/B PAND2X1_32/O 0.01fF
C23225 POR2X1_189/a_16_28# POR2X1_498/A 0.05fF
C23226 POR2X1_307/B POR2X1_307/A 0.00fF
C23227 POR2X1_440/Y PAND2X1_41/B 0.07fF
C23228 POR2X1_248/Y POR2X1_5/Y 0.03fF
C23229 PAND2X1_694/O POR2X1_614/A 0.17fF
C23230 POR2X1_673/A PAND2X1_4/CTRL 0.00fF
C23231 PAND2X1_693/O PAND2X1_48/B 0.04fF
C23232 POR2X1_14/Y POR2X1_583/Y 0.00fF
C23233 POR2X1_785/CTRL2 PAND2X1_32/B 0.04fF
C23234 POR2X1_740/Y POR2X1_574/CTRL2 0.04fF
C23235 PAND2X1_65/B POR2X1_577/a_16_28# 0.02fF
C23236 PAND2X1_717/O PAND2X1_493/Y 0.02fF
C23237 POR2X1_278/Y POR2X1_38/Y 0.21fF
C23238 PAND2X1_787/A VDD 0.18fF
C23239 PAND2X1_386/O POR2X1_707/Y 0.02fF
C23240 POR2X1_294/B PAND2X1_504/O 0.04fF
C23241 POR2X1_32/A POR2X1_109/Y 0.04fF
C23242 PAND2X1_322/O PAND2X1_32/B 0.03fF
C23243 PAND2X1_72/CTRL POR2X1_579/Y 0.00fF
C23244 PAND2X1_6/A POR2X1_55/Y 0.51fF
C23245 POR2X1_16/A PAND2X1_211/A 0.02fF
C23246 POR2X1_7/B POR2X1_90/Y 0.41fF
C23247 POR2X1_57/A PAND2X1_549/O 0.04fF
C23248 POR2X1_54/CTRL PAND2X1_58/A 0.01fF
C23249 PAND2X1_731/O POR2X1_763/Y 0.09fF
C23250 PAND2X1_621/a_56_28# POR2X1_750/B 0.00fF
C23251 POR2X1_327/Y PAND2X1_279/O 0.04fF
C23252 VDD POR2X1_148/B 0.13fF
C23253 POR2X1_247/Y POR2X1_294/A 0.10fF
C23254 POR2X1_180/B PAND2X1_65/B 0.04fF
C23255 PAND2X1_90/A POR2X1_243/CTRL2 0.03fF
C23256 PAND2X1_799/O INPUT_0 0.05fF
C23257 POR2X1_829/A POR2X1_38/Y 0.02fF
C23258 POR2X1_174/B PAND2X1_165/CTRL2 0.06fF
C23259 PAND2X1_341/A PAND2X1_197/CTRL2 0.01fF
C23260 PAND2X1_228/O POR2X1_52/Y 0.15fF
C23261 POR2X1_748/A POR2X1_129/Y 0.03fF
C23262 PAND2X1_725/Y POR2X1_394/A 0.03fF
C23263 POR2X1_201/Y VDD 0.02fF
C23264 POR2X1_618/O POR2X1_38/B 0.03fF
C23265 PAND2X1_421/CTRL POR2X1_596/A 0.01fF
C23266 POR2X1_502/A POR2X1_319/Y 13.91fF
C23267 POR2X1_580/O POR2X1_566/B 0.02fF
C23268 PAND2X1_658/A PAND2X1_548/CTRL 0.01fF
C23269 PAND2X1_44/CTRL2 PAND2X1_18/B -0.00fF
C23270 POR2X1_593/O POR2X1_750/B 0.01fF
C23271 POR2X1_119/Y POR2X1_14/Y 0.03fF
C23272 POR2X1_517/CTRL2 POR2X1_669/B 0.01fF
C23273 POR2X1_52/A POR2X1_239/Y 0.01fF
C23274 POR2X1_570/CTRL POR2X1_569/A 0.08fF
C23275 PAND2X1_592/O POR2X1_283/A 0.09fF
C23276 PAND2X1_255/O POR2X1_814/A 0.02fF
C23277 POR2X1_193/A POR2X1_228/Y 0.12fF
C23278 POR2X1_493/CTRL POR2X1_294/B 0.14fF
C23279 POR2X1_579/Y POR2X1_228/Y 0.03fF
C23280 POR2X1_632/a_16_28# POR2X1_632/Y 0.03fF
C23281 POR2X1_175/B VDD 0.11fF
C23282 PAND2X1_55/Y POR2X1_318/A 0.19fF
C23283 POR2X1_614/A PAND2X1_72/CTRL 0.01fF
C23284 PAND2X1_96/B PAND2X1_316/CTRL 0.01fF
C23285 PAND2X1_748/O VDD -0.00fF
C23286 POR2X1_57/A PAND2X1_652/A 0.03fF
C23287 POR2X1_16/A POR2X1_821/CTRL 0.02fF
C23288 POR2X1_416/CTRL2 POR2X1_293/Y 0.01fF
C23289 PAND2X1_477/B POR2X1_90/Y 0.02fF
C23290 POR2X1_78/B PAND2X1_824/B 0.10fF
C23291 POR2X1_203/Y POR2X1_786/Y 0.03fF
C23292 POR2X1_333/CTRL POR2X1_578/Y 0.03fF
C23293 PAND2X1_84/CTRL2 POR2X1_394/A 0.05fF
C23294 PAND2X1_495/CTRL2 PAND2X1_69/A 0.00fF
C23295 PAND2X1_793/Y PAND2X1_489/CTRL 0.01fF
C23296 POR2X1_65/A PAND2X1_325/CTRL 0.00fF
C23297 D_INPUT_0 PAND2X1_56/A 0.03fF
C23298 POR2X1_403/CTRL2 POR2X1_294/A 0.00fF
C23299 POR2X1_96/A PAND2X1_356/a_56_28# 0.00fF
C23300 PAND2X1_651/Y PAND2X1_341/A 0.05fF
C23301 POR2X1_83/Y POR2X1_60/Y 0.90fF
C23302 POR2X1_416/B D_INPUT_0 0.15fF
C23303 POR2X1_49/Y POR2X1_616/Y 0.03fF
C23304 POR2X1_795/B PAND2X1_60/B 0.02fF
C23305 PAND2X1_56/Y PAND2X1_60/B 0.03fF
C23306 POR2X1_184/Y POR2X1_91/Y 0.03fF
C23307 POR2X1_16/A POR2X1_96/A 1.05fF
C23308 PAND2X1_215/B POR2X1_7/CTRL2 0.03fF
C23309 POR2X1_177/CTRL POR2X1_236/Y 0.01fF
C23310 POR2X1_680/Y PAND2X1_728/CTRL 0.01fF
C23311 PAND2X1_522/O INPUT_0 0.04fF
C23312 POR2X1_327/Y POR2X1_217/O 0.01fF
C23313 PAND2X1_388/Y POR2X1_183/Y 0.03fF
C23314 POR2X1_740/Y POR2X1_568/Y 0.05fF
C23315 PAND2X1_4/CTRL D_INPUT_1 0.01fF
C23316 PAND2X1_57/B POR2X1_244/Y 0.03fF
C23317 POR2X1_353/Y POR2X1_192/B 0.85fF
C23318 PAND2X1_651/Y POR2X1_91/Y 0.10fF
C23319 PAND2X1_90/A POR2X1_276/Y 0.03fF
C23320 POR2X1_745/Y POR2X1_73/Y 0.00fF
C23321 POR2X1_88/Y POR2X1_394/A 0.05fF
C23322 POR2X1_614/A POR2X1_228/Y 0.32fF
C23323 POR2X1_388/a_16_28# PAND2X1_69/A 0.03fF
C23324 POR2X1_730/B POR2X1_729/Y 0.23fF
C23325 POR2X1_574/Y PAND2X1_516/CTRL 0.01fF
C23326 POR2X1_333/A POR2X1_731/Y 0.09fF
C23327 POR2X1_528/Y POR2X1_305/Y 0.12fF
C23328 POR2X1_62/Y PAND2X1_84/Y 0.29fF
C23329 POR2X1_87/O POR2X1_590/A 0.05fF
C23330 POR2X1_550/A POR2X1_614/A 0.23fF
C23331 POR2X1_608/CTRL POR2X1_294/A 0.03fF
C23332 PAND2X1_447/O POR2X1_329/A 0.06fF
C23333 POR2X1_829/A POR2X1_153/Y 0.00fF
C23334 POR2X1_447/B PAND2X1_627/CTRL 0.06fF
C23335 POR2X1_3/A INPUT_6 0.04fF
C23336 POR2X1_804/A POR2X1_725/Y 0.10fF
C23337 PAND2X1_853/B PAND2X1_364/B 0.07fF
C23338 PAND2X1_319/B POR2X1_142/Y 0.07fF
C23339 POR2X1_502/A POR2X1_266/A 0.03fF
C23340 POR2X1_46/Y PAND2X1_123/Y 0.09fF
C23341 POR2X1_624/B POR2X1_623/Y 0.00fF
C23342 PAND2X1_201/O PAND2X1_206/B 0.00fF
C23343 POR2X1_740/Y POR2X1_787/a_76_344# 0.03fF
C23344 POR2X1_110/O INPUT_0 0.06fF
C23345 D_INPUT_6 POR2X1_1/CTRL2 0.01fF
C23346 PAND2X1_90/A PAND2X1_531/CTRL2 0.07fF
C23347 PAND2X1_65/B PAND2X1_517/O 0.02fF
C23348 PAND2X1_305/a_76_28# PAND2X1_32/B 0.02fF
C23349 INPUT_1 PAND2X1_401/a_16_344# 0.02fF
C23350 PAND2X1_23/Y POR2X1_544/B 1.32fF
C23351 VDD POR2X1_4/Y 4.56fF
C23352 POR2X1_383/A PAND2X1_494/m4_208_n4# 0.07fF
C23353 POR2X1_325/A POR2X1_374/CTRL 0.01fF
C23354 POR2X1_732/CTRL POR2X1_353/A 0.01fF
C23355 POR2X1_327/Y PAND2X1_421/O 0.17fF
C23356 POR2X1_814/B PAND2X1_179/a_56_28# 0.00fF
C23357 POR2X1_294/B POR2X1_186/B 0.03fF
C23358 POR2X1_366/Y POR2X1_186/B 0.07fF
C23359 PAND2X1_392/CTRL2 POR2X1_816/A 0.01fF
C23360 POR2X1_145/Y POR2X1_146/CTRL2 0.00fF
C23361 PAND2X1_659/Y POR2X1_79/Y 0.00fF
C23362 POR2X1_467/Y PAND2X1_52/B 0.01fF
C23363 PAND2X1_493/a_76_28# PAND2X1_480/B 0.01fF
C23364 POR2X1_20/B PAND2X1_97/Y 0.42fF
C23365 PAND2X1_797/Y PAND2X1_209/O 0.02fF
C23366 PAND2X1_7/a_16_344# POR2X1_259/B 0.01fF
C23367 PAND2X1_65/B POR2X1_169/A 0.04fF
C23368 PAND2X1_297/CTRL POR2X1_68/B 0.01fF
C23369 POR2X1_175/B PAND2X1_32/B 0.01fF
C23370 PAND2X1_94/A POR2X1_649/B 0.09fF
C23371 POR2X1_383/A PAND2X1_60/B 3.99fF
C23372 INPUT_1 INPUT_2 0.03fF
C23373 POR2X1_110/Y POR2X1_7/B 0.03fF
C23374 PAND2X1_642/O PAND2X1_642/B 0.00fF
C23375 POR2X1_661/A D_INPUT_0 0.07fF
C23376 POR2X1_162/Y PAND2X1_158/CTRL 0.01fF
C23377 PAND2X1_242/Y POR2X1_423/CTRL 0.06fF
C23378 POR2X1_289/O POR2X1_394/A 0.06fF
C23379 PAND2X1_44/O PAND2X1_72/A 0.01fF
C23380 POR2X1_72/B PAND2X1_327/a_76_28# 0.01fF
C23381 PAND2X1_311/O POR2X1_260/A 0.17fF
C23382 POR2X1_236/Y POR2X1_39/B 2.56fF
C23383 POR2X1_814/A POR2X1_220/O 0.25fF
C23384 PAND2X1_90/Y PAND2X1_56/A 0.03fF
C23385 POR2X1_16/A POR2X1_689/Y 0.01fF
C23386 POR2X1_123/B POR2X1_260/A 0.01fF
C23387 POR2X1_119/Y POR2X1_55/Y 0.03fF
C23388 POR2X1_621/a_16_28# POR2X1_621/A 0.03fF
C23389 POR2X1_567/A POR2X1_785/A 0.05fF
C23390 POR2X1_131/Y POR2X1_387/Y 0.01fF
C23391 POR2X1_98/A POR2X1_66/A 2.34fF
C23392 POR2X1_777/B POR2X1_138/A 0.05fF
C23393 POR2X1_715/A POR2X1_112/Y 0.07fF
C23394 PAND2X1_79/O POR2X1_571/Y 0.04fF
C23395 POR2X1_65/Y PAND2X1_201/O 0.04fF
C23396 POR2X1_643/CTRL2 POR2X1_590/A 0.01fF
C23397 PAND2X1_846/CTRL2 INPUT_0 0.32fF
C23398 PAND2X1_241/Y PAND2X1_308/Y 0.01fF
C23399 POR2X1_16/A POR2X1_7/A 0.10fF
C23400 POR2X1_66/m4_208_n4# PAND2X1_39/B 0.07fF
C23401 POR2X1_96/A POR2X1_184/a_76_344# 0.03fF
C23402 POR2X1_416/B POR2X1_697/a_16_28# 0.02fF
C23403 PAND2X1_53/CTRL2 POR2X1_66/A 0.01fF
C23404 PAND2X1_765/CTRL POR2X1_260/A 0.02fF
C23405 POR2X1_383/A POR2X1_353/A 0.03fF
C23406 PAND2X1_476/A POR2X1_43/B 0.05fF
C23407 PAND2X1_81/B POR2X1_4/Y 0.00fF
C23408 PAND2X1_69/A POR2X1_294/A 0.97fF
C23409 POR2X1_394/A POR2X1_757/CTRL 0.05fF
C23410 POR2X1_567/A PAND2X1_504/O -0.01fF
C23411 POR2X1_54/Y PAND2X1_9/Y 0.03fF
C23412 POR2X1_814/A POR2X1_218/Y 0.07fF
C23413 POR2X1_856/B PAND2X1_52/O 0.27fF
C23414 POR2X1_614/A POR2X1_156/CTRL 0.01fF
C23415 POR2X1_809/A POR2X1_809/Y 0.27fF
C23416 POR2X1_262/Y PAND2X1_560/a_76_28# 0.01fF
C23417 POR2X1_383/A POR2X1_571/O 0.07fF
C23418 POR2X1_241/Y PAND2X1_52/B 0.00fF
C23419 VDD POR2X1_173/CTRL -0.00fF
C23420 POR2X1_703/A POR2X1_456/B 0.07fF
C23421 POR2X1_103/O PAND2X1_349/A 0.01fF
C23422 POR2X1_57/A PAND2X1_779/O 0.04fF
C23423 POR2X1_532/A PAND2X1_692/O 0.16fF
C23424 POR2X1_25/Y INPUT_6 0.03fF
C23425 POR2X1_4/Y PAND2X1_32/B 0.07fF
C23426 PAND2X1_71/Y PAND2X1_60/B 0.03fF
C23427 POR2X1_38/O POR2X1_411/B 0.02fF
C23428 POR2X1_411/B PAND2X1_218/B 0.02fF
C23429 POR2X1_8/Y POR2X1_10/CTRL2 0.01fF
C23430 POR2X1_23/Y POR2X1_150/Y 0.03fF
C23431 POR2X1_188/O POR2X1_737/A 0.01fF
C23432 POR2X1_136/Y POR2X1_183/O 0.03fF
C23433 PAND2X1_854/A PAND2X1_345/Y 0.82fF
C23434 PAND2X1_716/B PAND2X1_303/B 0.13fF
C23435 POR2X1_20/B PAND2X1_771/Y 0.05fF
C23436 POR2X1_152/CTRL POR2X1_39/B 0.00fF
C23437 POR2X1_101/A POR2X1_101/a_16_28# 0.05fF
C23438 PAND2X1_691/Y PAND2X1_686/a_76_28# 0.02fF
C23439 PAND2X1_93/B PAND2X1_39/B 0.10fF
C23440 POR2X1_788/CTRL PAND2X1_60/B 0.01fF
C23441 POR2X1_407/A POR2X1_779/O 0.16fF
C23442 PAND2X1_95/B PAND2X1_52/B 0.05fF
C23443 POR2X1_54/Y POR2X1_818/Y 0.05fF
C23444 PAND2X1_655/Y PAND2X1_691/O 0.03fF
C23445 POR2X1_730/Y POR2X1_151/Y 0.03fF
C23446 POR2X1_8/Y POR2X1_394/A 4.21fF
C23447 POR2X1_561/a_16_28# POR2X1_558/Y 0.10fF
C23448 POR2X1_407/A POR2X1_343/Y 0.05fF
C23449 POR2X1_234/A PAND2X1_520/O 0.02fF
C23450 POR2X1_8/Y POR2X1_749/CTRL 0.01fF
C23451 POR2X1_754/Y POR2X1_20/B 0.07fF
C23452 POR2X1_591/Y POR2X1_761/A 0.03fF
C23453 POR2X1_86/CTRL2 PAND2X1_338/B 0.01fF
C23454 POR2X1_540/Y POR2X1_569/A 0.01fF
C23455 POR2X1_250/Y PAND2X1_742/a_16_344# 0.04fF
C23456 POR2X1_546/CTRL2 POR2X1_550/B 0.00fF
C23457 PAND2X1_72/Y PAND2X1_48/A 0.01fF
C23458 PAND2X1_184/a_16_344# PAND2X1_71/Y 0.02fF
C23459 PAND2X1_20/A POR2X1_137/B 0.50fF
C23460 D_GATE_222 POR2X1_568/A 0.07fF
C23461 POR2X1_274/A POR2X1_274/CTRL2 0.01fF
C23462 POR2X1_621/A POR2X1_296/B 0.03fF
C23463 PAND2X1_824/B POR2X1_294/A 0.03fF
C23464 POR2X1_456/B PAND2X1_167/CTRL2 0.11fF
C23465 PAND2X1_94/A PAND2X1_122/CTRL2 0.13fF
C23466 PAND2X1_108/CTRL2 PAND2X1_60/B 0.01fF
C23467 POR2X1_327/Y POR2X1_326/A 0.12fF
C23468 POR2X1_20/B PAND2X1_719/Y 0.01fF
C23469 POR2X1_571/O POR2X1_560/Y 0.00fF
C23470 POR2X1_78/A PAND2X1_39/B 0.34fF
C23471 PAND2X1_76/Y POR2X1_329/A 0.07fF
C23472 POR2X1_66/B POR2X1_649/O 0.17fF
C23473 POR2X1_673/Y POR2X1_4/Y 0.07fF
C23474 POR2X1_1/CTRL D_INPUT_4 0.03fF
C23475 PAND2X1_241/Y POR2X1_77/Y 0.03fF
C23476 PAND2X1_838/B POR2X1_667/A 0.05fF
C23477 PAND2X1_91/a_16_344# POR2X1_97/A 0.01fF
C23478 POR2X1_834/O POR2X1_260/B 0.01fF
C23479 PAND2X1_613/O POR2X1_296/B 0.04fF
C23480 POR2X1_220/A POR2X1_161/CTRL 0.01fF
C23481 PAND2X1_63/O POR2X1_66/A 0.10fF
C23482 POR2X1_567/A POR2X1_186/B 0.11fF
C23483 POR2X1_350/B PAND2X1_52/B 0.03fF
C23484 PAND2X1_497/O POR2X1_590/A 0.10fF
C23485 POR2X1_846/Y POR2X1_615/a_16_28# 0.01fF
C23486 POR2X1_648/Y PAND2X1_511/a_16_344# 0.01fF
C23487 POR2X1_65/A PAND2X1_838/O 0.01fF
C23488 POR2X1_503/CTRL2 POR2X1_77/Y 0.01fF
C23489 POR2X1_416/B POR2X1_108/Y 0.33fF
C23490 POR2X1_760/A PAND2X1_730/B 0.01fF
C23491 POR2X1_623/O POR2X1_296/B 0.02fF
C23492 POR2X1_722/A PAND2X1_696/O 0.03fF
C23493 POR2X1_446/B POR2X1_750/B 0.05fF
C23494 PAND2X1_434/O POR2X1_83/B 0.15fF
C23495 POR2X1_453/Y VDD 0.10fF
C23496 PAND2X1_20/A PAND2X1_93/B 0.27fF
C23497 POR2X1_150/Y PAND2X1_558/O 0.02fF
C23498 POR2X1_808/A POR2X1_808/CTRL 0.07fF
C23499 POR2X1_23/Y PAND2X1_794/O 0.01fF
C23500 PAND2X1_86/CTRL POR2X1_404/Y 0.00fF
C23501 POR2X1_294/a_16_28# POR2X1_355/A 0.03fF
C23502 POR2X1_709/A PAND2X1_65/B 0.03fF
C23503 POR2X1_458/Y POR2X1_741/Y 0.07fF
C23504 PAND2X1_373/O PAND2X1_72/A 0.18fF
C23505 POR2X1_65/A PAND2X1_206/A 0.01fF
C23506 POR2X1_78/Y VDD 0.27fF
C23507 POR2X1_271/A POR2X1_39/B 0.03fF
C23508 POR2X1_597/Y VDD 0.08fF
C23509 PAND2X1_571/O PAND2X1_561/Y 0.00fF
C23510 POR2X1_849/B POR2X1_94/A 0.02fF
C23511 POR2X1_56/a_56_344# POR2X1_496/Y 0.00fF
C23512 POR2X1_270/Y POR2X1_269/Y 0.08fF
C23513 PAND2X1_9/CTRL2 POR2X1_29/A 0.09fF
C23514 PAND2X1_73/Y POR2X1_241/B 0.12fF
C23515 POR2X1_748/A POR2X1_37/Y 5.14fF
C23516 PAND2X1_352/O PAND2X1_352/B 0.00fF
C23517 PAND2X1_469/CTRL2 POR2X1_236/Y 0.01fF
C23518 PAND2X1_689/O POR2X1_812/A 0.04fF
C23519 POR2X1_89/CTRL2 POR2X1_5/Y 0.00fF
C23520 POR2X1_78/A POR2X1_805/Y 0.51fF
C23521 POR2X1_20/B POR2X1_233/CTRL 0.00fF
C23522 PAND2X1_258/CTRL2 PAND2X1_52/Y 0.01fF
C23523 POR2X1_465/CTRL2 POR2X1_563/Y 0.01fF
C23524 PAND2X1_97/CTRL2 POR2X1_5/Y 0.00fF
C23525 POR2X1_68/A POR2X1_814/A 0.25fF
C23526 POR2X1_13/A PAND2X1_98/O 0.06fF
C23527 POR2X1_814/B PAND2X1_93/B 0.10fF
C23528 POR2X1_458/Y PAND2X1_32/B 0.01fF
C23529 POR2X1_49/Y PAND2X1_61/CTRL2 0.00fF
C23530 PAND2X1_20/A POR2X1_78/A 2.19fF
C23531 POR2X1_719/A PAND2X1_73/Y 0.00fF
C23532 PAND2X1_793/Y POR2X1_411/B 0.03fF
C23533 PAND2X1_862/B PAND2X1_203/O 0.08fF
C23534 PAND2X1_477/O PAND2X1_803/A 0.00fF
C23535 POR2X1_72/O POR2X1_23/Y 0.02fF
C23536 POR2X1_32/A PAND2X1_706/CTRL2 0.02fF
C23537 POR2X1_66/B POR2X1_555/B 0.03fF
C23538 PAND2X1_45/O POR2X1_741/Y 0.01fF
C23539 PAND2X1_88/CTRL POR2X1_590/A 0.01fF
C23540 PAND2X1_561/O PAND2X1_558/Y 0.02fF
C23541 PAND2X1_841/B POR2X1_411/B 0.51fF
C23542 POR2X1_193/A POR2X1_657/Y 0.05fF
C23543 POR2X1_20/B POR2X1_42/Y 0.17fF
C23544 POR2X1_864/A POR2X1_800/A 0.05fF
C23545 POR2X1_23/Y POR2X1_29/CTRL 0.00fF
C23546 PAND2X1_93/B POR2X1_325/A 0.10fF
C23547 POR2X1_251/A POR2X1_102/Y 1.25fF
C23548 POR2X1_83/B POR2X1_698/CTRL2 0.00fF
C23549 POR2X1_260/B PAND2X1_131/O 0.02fF
C23550 POR2X1_121/B POR2X1_750/B 0.05fF
C23551 POR2X1_590/A PAND2X1_41/B 9.87fF
C23552 POR2X1_383/A POR2X1_655/O 0.01fF
C23553 POR2X1_102/Y POR2X1_72/B 0.23fF
C23554 POR2X1_48/A POR2X1_236/Y 0.08fF
C23555 POR2X1_807/O POR2X1_480/A 0.03fF
C23556 POR2X1_499/A POR2X1_218/A 0.07fF
C23557 POR2X1_866/A PAND2X1_57/B 0.05fF
C23558 POR2X1_416/B PAND2X1_643/A 0.06fF
C23559 POR2X1_565/B POR2X1_624/Y 0.03fF
C23560 POR2X1_66/B POR2X1_330/Y 0.06fF
C23561 POR2X1_549/CTRL POR2X1_78/A 0.01fF
C23562 POR2X1_138/CTRL2 POR2X1_624/Y 0.09fF
C23563 POR2X1_814/B POR2X1_78/A 10.94fF
C23564 POR2X1_20/B POR2X1_309/Y 0.03fF
C23565 POR2X1_411/B POR2X1_665/Y 0.37fF
C23566 PAND2X1_217/CTRL POR2X1_599/A 0.01fF
C23567 PAND2X1_594/O PAND2X1_90/Y 0.21fF
C23568 POR2X1_648/Y PAND2X1_60/B 0.03fF
C23569 POR2X1_60/A PAND2X1_185/O 0.05fF
C23570 POR2X1_695/Y VDD 0.09fF
C23571 PAND2X1_673/CTRL2 POR2X1_83/B 0.00fF
C23572 POR2X1_496/Y PAND2X1_778/O 0.02fF
C23573 POR2X1_454/A POR2X1_579/Y 0.03fF
C23574 POR2X1_188/A POR2X1_330/Y 0.05fF
C23575 PAND2X1_829/O PAND2X1_65/B 0.03fF
C23576 POR2X1_52/A PAND2X1_218/B 0.06fF
C23577 PAND2X1_93/B POR2X1_513/B 0.07fF
C23578 PAND2X1_717/A PAND2X1_349/A 0.03fF
C23579 PAND2X1_630/B PAND2X1_507/CTRL2 0.01fF
C23580 POR2X1_126/CTRL D_INPUT_2 0.00fF
C23581 PAND2X1_65/B PAND2X1_58/A 0.08fF
C23582 POR2X1_422/O POR2X1_293/Y 0.26fF
C23583 POR2X1_23/Y PAND2X1_364/B 0.07fF
C23584 POR2X1_140/B POR2X1_624/Y 0.03fF
C23585 PAND2X1_296/CTRL2 PAND2X1_347/Y 0.01fF
C23586 POR2X1_78/A POR2X1_325/A 0.03fF
C23587 PAND2X1_781/O POR2X1_745/Y 0.04fF
C23588 PAND2X1_629/O POR2X1_626/Y 0.01fF
C23589 POR2X1_416/B PAND2X1_198/CTRL 0.06fF
C23590 POR2X1_32/A PAND2X1_596/m4_208_n4# 0.09fF
C23591 POR2X1_102/Y PAND2X1_756/O 0.02fF
C23592 POR2X1_43/B PAND2X1_436/CTRL 0.01fF
C23593 POR2X1_114/B PAND2X1_406/CTRL2 0.06fF
C23594 INPUT_3 POR2X1_380/a_16_28# 0.06fF
C23595 POR2X1_97/A POR2X1_853/CTRL 0.00fF
C23596 POR2X1_119/Y PAND2X1_862/m4_208_n4# 0.04fF
C23597 PAND2X1_803/A POR2X1_40/Y 0.03fF
C23598 POR2X1_311/Y PAND2X1_730/B 5.11fF
C23599 PAND2X1_39/B POR2X1_784/CTRL 0.00fF
C23600 POR2X1_591/A POR2X1_666/A 0.02fF
C23601 PAND2X1_219/A VDD 0.22fF
C23602 POR2X1_78/B PAND2X1_420/O 0.01fF
C23603 PAND2X1_267/Y POR2X1_599/A 0.03fF
C23604 PAND2X1_71/CTRL2 POR2X1_296/B 0.03fF
C23605 POR2X1_311/Y GATE_741 0.05fF
C23606 PAND2X1_360/CTRL PAND2X1_347/Y 0.01fF
C23607 POR2X1_20/B PAND2X1_99/Y 0.02fF
C23608 PAND2X1_210/CTRL PAND2X1_725/Y 0.00fF
C23609 PAND2X1_106/CTRL POR2X1_116/A 0.00fF
C23610 POR2X1_614/A POR2X1_454/A 0.03fF
C23611 PAND2X1_220/Y PAND2X1_540/a_76_28# 0.03fF
C23612 PAND2X1_651/Y POR2X1_613/CTRL2 0.00fF
C23613 PAND2X1_616/CTRL VDD 0.00fF
C23614 POR2X1_186/Y POR2X1_742/CTRL2 0.01fF
C23615 POR2X1_78/A POR2X1_513/B 0.03fF
C23616 POR2X1_450/A VDD 0.00fF
C23617 POR2X1_333/A POR2X1_502/A 0.14fF
C23618 POR2X1_220/CTRL POR2X1_210/Y 0.01fF
C23619 POR2X1_220/CTRL2 POR2X1_220/A 0.01fF
C23620 POR2X1_446/B POR2X1_714/CTRL2 0.01fF
C23621 POR2X1_366/CTRL2 POR2X1_556/A 0.01fF
C23622 POR2X1_16/A POR2X1_760/A 0.10fF
C23623 POR2X1_67/A PAND2X1_790/Y 0.07fF
C23624 POR2X1_272/Y POR2X1_423/Y 0.00fF
C23625 POR2X1_188/A POR2X1_733/a_76_344# 0.00fF
C23626 POR2X1_221/a_16_28# POR2X1_186/Y 0.02fF
C23627 POR2X1_273/Y D_INPUT_0 0.03fF
C23628 POR2X1_605/B POR2X1_220/Y 0.01fF
C23629 POR2X1_48/A POR2X1_232/Y 0.01fF
C23630 POR2X1_41/B POR2X1_482/Y 0.02fF
C23631 POR2X1_23/Y POR2X1_229/O 0.01fF
C23632 PAND2X1_458/a_76_28# PAND2X1_716/B 0.02fF
C23633 PAND2X1_52/Y VDD 0.46fF
C23634 PAND2X1_275/O POR2X1_296/B 0.01fF
C23635 POR2X1_702/B VDD 0.38fF
C23636 PAND2X1_714/A VDD 0.08fF
C23637 POR2X1_829/A PAND2X1_214/A 0.25fF
C23638 POR2X1_609/Y POR2X1_234/O 0.00fF
C23639 POR2X1_502/A POR2X1_734/A 0.07fF
C23640 PAND2X1_782/O POR2X1_747/Y 0.00fF
C23641 POR2X1_516/a_16_28# POR2X1_48/A 0.02fF
C23642 POR2X1_748/A POR2X1_293/Y 0.10fF
C23643 POR2X1_63/Y PAND2X1_737/B 0.03fF
C23644 PAND2X1_667/O PAND2X1_65/B 0.00fF
C23645 POR2X1_445/A POR2X1_569/A 0.07fF
C23646 POR2X1_278/CTRL2 PAND2X1_35/Y 0.01fF
C23647 POR2X1_66/A POR2X1_341/Y 0.04fF
C23648 POR2X1_672/CTRL2 POR2X1_102/Y 0.07fF
C23649 PAND2X1_65/B POR2X1_435/Y 0.03fF
C23650 POR2X1_135/Y VDD 0.12fF
C23651 POR2X1_857/B PAND2X1_41/B 15.74fF
C23652 D_INPUT_0 PAND2X1_575/O 0.02fF
C23653 PAND2X1_456/CTRL2 POR2X1_55/Y 0.00fF
C23654 POR2X1_855/B POR2X1_808/a_76_344# 0.00fF
C23655 POR2X1_861/A POR2X1_814/A 0.07fF
C23656 POR2X1_673/A VDD 0.11fF
C23657 POR2X1_834/O POR2X1_407/Y 0.01fF
C23658 POR2X1_237/Y POR2X1_14/Y 0.03fF
C23659 PAND2X1_793/Y POR2X1_376/B 0.03fF
C23660 POR2X1_57/CTRL2 POR2X1_5/Y 0.01fF
C23661 POR2X1_41/B POR2X1_106/Y 0.03fF
C23662 POR2X1_35/B PAND2X1_55/Y 0.03fF
C23663 PAND2X1_835/Y POR2X1_102/Y 0.02fF
C23664 POR2X1_750/B POR2X1_795/B 0.10fF
C23665 PAND2X1_721/B POR2X1_73/Y 0.03fF
C23666 POR2X1_136/Y D_INPUT_0 0.01fF
C23667 POR2X1_67/Y PAND2X1_526/CTRL2 0.01fF
C23668 PAND2X1_272/CTRL PAND2X1_60/B 0.02fF
C23669 POR2X1_65/A POR2X1_697/Y 0.04fF
C23670 PAND2X1_23/Y PAND2X1_55/CTRL 0.00fF
C23671 POR2X1_849/A POR2X1_7/A 0.01fF
C23672 POR2X1_130/A PAND2X1_755/O 0.05fF
C23673 POR2X1_523/Y POR2X1_94/A 0.03fF
C23674 POR2X1_459/O VDD 0.00fF
C23675 PAND2X1_480/B PAND2X1_151/CTRL 0.25fF
C23676 PAND2X1_245/CTRL2 PAND2X1_111/B 0.01fF
C23677 POR2X1_54/Y PAND2X1_522/a_16_344# 0.06fF
C23678 POR2X1_32/A PAND2X1_338/B 0.03fF
C23679 INPUT_0 POR2X1_572/O 0.08fF
C23680 POR2X1_72/B POR2X1_531/Y 0.04fF
C23681 POR2X1_41/B PAND2X1_580/B 0.03fF
C23682 PAND2X1_849/B POR2X1_23/Y 0.01fF
C23683 PAND2X1_52/Y POR2X1_741/Y 0.02fF
C23684 PAND2X1_593/CTRL PAND2X1_364/B 0.07fF
C23685 POR2X1_422/CTRL POR2X1_260/A 0.02fF
C23686 POR2X1_814/A POR2X1_169/A 0.29fF
C23687 POR2X1_235/CTRL POR2X1_32/A 0.01fF
C23688 POR2X1_68/A PAND2X1_55/CTRL2 0.03fF
C23689 PAND2X1_13/O POR2X1_795/B 0.05fF
C23690 POR2X1_201/CTRL2 PAND2X1_88/Y 0.01fF
C23691 PAND2X1_598/CTRL2 POR2X1_46/Y 0.01fF
C23692 PAND2X1_217/B POR2X1_816/A 0.07fF
C23693 POR2X1_594/a_16_28# POR2X1_594/A 0.02fF
C23694 POR2X1_69/A POR2X1_38/Y 0.03fF
C23695 POR2X1_94/A PAND2X1_69/A 0.37fF
C23696 INPUT_0 POR2X1_7/B 0.24fF
C23697 POR2X1_65/A PAND2X1_357/Y 0.03fF
C23698 POR2X1_717/a_16_28# POR2X1_590/A 0.00fF
C23699 PAND2X1_105/O PAND2X1_562/B 0.11fF
C23700 PAND2X1_483/O POR2X1_23/Y 0.03fF
C23701 POR2X1_550/A POR2X1_590/A 1.11fF
C23702 POR2X1_655/Y POR2X1_784/O 0.00fF
C23703 PAND2X1_13/CTRL2 PAND2X1_32/B 0.03fF
C23704 POR2X1_89/Y PAND2X1_244/B 0.01fF
C23705 POR2X1_13/A PAND2X1_735/a_76_28# 0.02fF
C23706 PAND2X1_401/CTRL POR2X1_236/Y 0.01fF
C23707 PAND2X1_96/B POR2X1_777/B 0.09fF
C23708 POR2X1_614/A POR2X1_264/a_16_28# 0.01fF
C23709 POR2X1_106/m4_208_n4# POR2X1_108/m4_208_n4# 0.13fF
C23710 POR2X1_556/A POR2X1_554/CTRL2 0.06fF
C23711 POR2X1_383/A PAND2X1_279/CTRL2 0.08fF
C23712 D_INPUT_1 PAND2X1_526/CTRL 0.02fF
C23713 PAND2X1_392/B POR2X1_816/A 0.01fF
C23714 PAND2X1_9/Y POR2X1_4/Y 0.18fF
C23715 POR2X1_274/a_16_28# POR2X1_274/B 0.07fF
C23716 PAND2X1_797/Y POR2X1_441/Y 0.03fF
C23717 PAND2X1_96/B POR2X1_194/A 0.03fF
C23718 POR2X1_367/a_16_28# POR2X1_366/Y 0.03fF
C23719 POR2X1_52/A PAND2X1_793/Y 0.03fF
C23720 PAND2X1_472/A POR2X1_5/Y 0.03fF
C23721 POR2X1_294/a_56_344# POR2X1_294/A 0.00fF
C23722 POR2X1_566/A PAND2X1_292/a_76_28# 0.04fF
C23723 POR2X1_490/Y PAND2X1_557/a_16_344# 0.05fF
C23724 POR2X1_308/a_16_28# POR2X1_740/Y 0.01fF
C23725 D_GATE_662 VDD 1.38fF
C23726 POR2X1_40/CTRL2 POR2X1_83/B 0.00fF
C23727 POR2X1_690/Y VDD 0.03fF
C23728 POR2X1_96/A PAND2X1_188/CTRL2 0.01fF
C23729 POR2X1_96/A POR2X1_680/Y 0.00fF
C23730 PAND2X1_6/A POR2X1_511/Y 0.07fF
C23731 PAND2X1_731/B POR2X1_91/Y 0.01fF
C23732 POR2X1_102/O POR2X1_411/B 0.01fF
C23733 POR2X1_271/A POR2X1_48/A 0.03fF
C23734 POR2X1_123/A POR2X1_634/A 0.03fF
C23735 PAND2X1_779/a_16_344# PAND2X1_549/B 0.01fF
C23736 POR2X1_848/O PAND2X1_52/B 0.01fF
C23737 POR2X1_41/B POR2X1_256/a_16_28# 0.05fF
C23738 PAND2X1_486/CTRL POR2X1_763/Y 0.03fF
C23739 POR2X1_355/B PAND2X1_23/Y 0.03fF
C23740 POR2X1_97/A PAND2X1_503/a_16_344# 0.02fF
C23741 POR2X1_358/CTRL2 POR2X1_578/Y 0.03fF
C23742 POR2X1_254/Y POR2X1_222/Y 0.07fF
C23743 PAND2X1_205/Y PAND2X1_186/a_56_28# 0.00fF
C23744 POR2X1_383/A POR2X1_254/A 0.03fF
C23745 POR2X1_210/CTRL2 POR2X1_210/B 0.01fF
C23746 POR2X1_32/Y POR2X1_5/Y 0.11fF
C23747 POR2X1_332/B POR2X1_775/A 0.85fF
C23748 PAND2X1_65/B PAND2X1_96/B 0.18fF
C23749 POR2X1_725/Y POR2X1_794/B 0.07fF
C23750 PAND2X1_213/B PAND2X1_213/A 0.02fF
C23751 POR2X1_8/Y POR2X1_669/B 0.08fF
C23752 POR2X1_32/A PAND2X1_341/Y 0.03fF
C23753 POR2X1_383/A POR2X1_750/B 0.17fF
C23754 POR2X1_409/a_16_28# POR2X1_5/Y 0.02fF
C23755 VDD POR2X1_816/A 1.60fF
C23756 POR2X1_566/A POR2X1_35/Y 0.05fF
C23757 POR2X1_462/B VDD 0.65fF
C23758 PAND2X1_569/A VDD 0.00fF
C23759 POR2X1_311/Y POR2X1_16/A 0.07fF
C23760 POR2X1_78/B POR2X1_538/a_16_28# 0.00fF
C23761 PAND2X1_620/O POR2X1_422/Y 0.05fF
C23762 PAND2X1_472/CTRL POR2X1_60/A 0.03fF
C23763 D_INPUT_1 VDD 2.35fF
C23764 PAND2X1_6/CTRL PAND2X1_20/A 0.01fF
C23765 PAND2X1_23/Y POR2X1_276/CTRL 0.03fF
C23766 POR2X1_65/A PAND2X1_140/A 0.03fF
C23767 POR2X1_49/Y PAND2X1_661/Y 0.01fF
C23768 POR2X1_57/A POR2X1_297/A 0.01fF
C23769 POR2X1_13/A POR2X1_299/CTRL2 0.03fF
C23770 D_INPUT_0 POR2X1_737/A 0.03fF
C23771 POR2X1_380/Y POR2X1_5/Y 0.04fF
C23772 POR2X1_502/A POR2X1_775/O 0.31fF
C23773 POR2X1_532/A POR2X1_794/CTRL 0.01fF
C23774 PAND2X1_710/CTRL2 POR2X1_763/A 0.04fF
C23775 POR2X1_65/A POR2X1_528/Y 0.07fF
C23776 POR2X1_332/B POR2X1_112/Y 0.07fF
C23777 PAND2X1_254/Y POR2X1_253/Y 0.03fF
C23778 POR2X1_628/CTRL2 PAND2X1_6/A 0.04fF
C23779 POR2X1_582/O VDD -0.00fF
C23780 POR2X1_840/B POR2X1_217/a_76_344# 0.04fF
C23781 VDD POR2X1_724/A 0.14fF
C23782 POR2X1_170/B POR2X1_577/CTRL2 0.09fF
C23783 PAND2X1_754/CTRL2 PAND2X1_69/A 0.01fF
C23784 POR2X1_433/CTRL POR2X1_153/Y 0.06fF
C23785 POR2X1_43/B PAND2X1_466/CTRL 0.01fF
C23786 POR2X1_709/O POR2X1_814/B 0.01fF
C23787 PAND2X1_676/CTRL PAND2X1_480/B 0.07fF
C23788 POR2X1_693/O POR2X1_73/Y 0.01fF
C23789 POR2X1_691/CTRL POR2X1_800/A 0.00fF
C23790 POR2X1_62/Y POR2X1_296/B 0.06fF
C23791 POR2X1_83/B PAND2X1_337/a_16_344# 0.02fF
C23792 POR2X1_83/B PAND2X1_508/Y 0.03fF
C23793 INPUT_0 PAND2X1_60/B 0.10fF
C23794 POR2X1_96/Y POR2X1_263/Y 0.03fF
C23795 POR2X1_360/A POR2X1_38/B 0.04fF
C23796 POR2X1_460/A INPUT_5 0.91fF
C23797 PAND2X1_319/m4_208_n4# POR2X1_258/m4_208_n4# 0.13fF
C23798 PAND2X1_854/A VDD 2.08fF
C23799 POR2X1_829/A POR2X1_591/Y 0.03fF
C23800 POR2X1_165/Y POR2X1_72/B 0.02fF
C23801 PAND2X1_658/A POR2X1_56/Y 0.03fF
C23802 PAND2X1_557/A PAND2X1_557/O 0.00fF
C23803 POR2X1_376/B POR2X1_376/CTRL 0.01fF
C23804 PAND2X1_35/Y PAND2X1_338/B 0.03fF
C23805 VDD POR2X1_356/B 0.44fF
C23806 POR2X1_293/Y POR2X1_291/Y 0.00fF
C23807 POR2X1_246/CTRL POR2X1_90/Y 0.01fF
C23808 POR2X1_532/Y POR2X1_788/B 0.03fF
C23809 PAND2X1_48/B POR2X1_210/Y 4.54fF
C23810 POR2X1_43/B PAND2X1_734/CTRL 0.01fF
C23811 POR2X1_311/Y PAND2X1_336/Y 0.08fF
C23812 POR2X1_712/A PAND2X1_697/CTRL 0.01fF
C23813 POR2X1_655/A POR2X1_725/CTRL 0.01fF
C23814 POR2X1_96/A PAND2X1_549/B 0.00fF
C23815 POR2X1_858/A D_INPUT_0 0.01fF
C23816 POR2X1_855/B POR2X1_220/Y 0.03fF
C23817 PAND2X1_81/B D_INPUT_1 0.03fF
C23818 POR2X1_564/Y POR2X1_704/O 0.01fF
C23819 POR2X1_41/B PAND2X1_349/A 0.03fF
C23820 POR2X1_192/Y POR2X1_714/a_16_28# 0.04fF
C23821 PAND2X1_591/CTRL2 PAND2X1_56/A 0.01fF
C23822 POR2X1_785/CTRL POR2X1_566/B 0.07fF
C23823 POR2X1_262/CTRL POR2X1_7/A 0.01fF
C23824 POR2X1_23/a_76_344# POR2X1_4/Y 0.01fF
C23825 POR2X1_41/B PAND2X1_63/B 0.01fF
C23826 POR2X1_673/A POR2X1_673/Y 0.01fF
C23827 PAND2X1_553/a_16_344# POR2X1_55/Y 0.02fF
C23828 POR2X1_655/A PAND2X1_52/B 0.01fF
C23829 PAND2X1_170/a_76_28# PAND2X1_168/Y 0.02fF
C23830 PAND2X1_691/Y PAND2X1_719/O 0.04fF
C23831 POR2X1_804/B PAND2X1_69/A 0.01fF
C23832 PAND2X1_220/Y PAND2X1_360/Y 0.03fF
C23833 POR2X1_743/CTRL POR2X1_153/Y 0.01fF
C23834 POR2X1_741/Y POR2X1_724/A 8.76fF
C23835 POR2X1_21/a_16_28# INPUT_5 0.00fF
C23836 PAND2X1_139/B PAND2X1_216/B 0.01fF
C23837 PAND2X1_741/B POR2X1_7/a_76_344# 0.03fF
C23838 PAND2X1_57/B POR2X1_596/CTRL2 0.00fF
C23839 POR2X1_771/CTRL2 PAND2X1_32/B 0.01fF
C23840 POR2X1_228/CTRL PAND2X1_52/Y 0.01fF
C23841 POR2X1_56/Y POR2X1_73/Y 11.38fF
C23842 POR2X1_816/A PAND2X1_32/B 0.03fF
C23843 PAND2X1_57/B POR2X1_703/A 0.07fF
C23844 POR2X1_334/O INPUT_0 0.10fF
C23845 PAND2X1_228/CTRL PAND2X1_656/A 0.01fF
C23846 D_INPUT_1 PAND2X1_32/B 0.13fF
C23847 POR2X1_123/A POR2X1_123/O 0.03fF
C23848 POR2X1_304/CTRL POR2X1_102/Y 0.01fF
C23849 POR2X1_57/A PAND2X1_566/Y 0.06fF
C23850 POR2X1_383/A PAND2X1_71/a_16_344# 0.02fF
C23851 POR2X1_327/Y POR2X1_480/A 0.10fF
C23852 POR2X1_287/B PAND2X1_48/A 0.03fF
C23853 PAND2X1_768/Y PAND2X1_359/Y 0.02fF
C23854 POR2X1_52/O POR2X1_102/Y 0.01fF
C23855 PAND2X1_220/A POR2X1_77/Y 0.14fF
C23856 POR2X1_116/Y POR2X1_392/O 0.02fF
C23857 POR2X1_96/A PAND2X1_472/O 0.03fF
C23858 POR2X1_153/CTRL2 PAND2X1_472/B 0.05fF
C23859 PAND2X1_812/O PAND2X1_811/Y 0.03fF
C23860 PAND2X1_793/Y PAND2X1_510/CTRL 0.01fF
C23861 PAND2X1_798/B PAND2X1_175/B 0.02fF
C23862 POR2X1_754/A POR2X1_260/A 0.03fF
C23863 PAND2X1_140/A PAND2X1_190/Y 0.17fF
C23864 POR2X1_857/B POR2X1_502/CTRL 0.03fF
C23865 PAND2X1_472/a_56_28# PAND2X1_673/Y 0.00fF
C23866 POR2X1_103/CTRL2 POR2X1_13/A 0.00fF
C23867 POR2X1_357/Y POR2X1_319/Y 0.01fF
C23868 POR2X1_724/A PAND2X1_32/B 0.06fF
C23869 D_GATE_741 POR2X1_854/B 0.10fF
C23870 POR2X1_305/Y POR2X1_245/Y 0.02fF
C23871 POR2X1_356/A POR2X1_260/A 0.12fF
C23872 POR2X1_483/A PAND2X1_48/A 0.00fF
C23873 POR2X1_306/a_56_344# POR2X1_90/Y 0.00fF
C23874 POR2X1_62/Y POR2X1_236/Y 0.05fF
C23875 PAND2X1_357/CTRL VDD 0.00fF
C23876 POR2X1_283/A PAND2X1_794/B 0.03fF
C23877 PAND2X1_81/CTRL2 PAND2X1_63/B 0.01fF
C23878 POR2X1_133/O POR2X1_384/A 0.01fF
C23879 POR2X1_336/CTRL2 POR2X1_228/Y 0.01fF
C23880 POR2X1_486/CTRL POR2X1_705/B 0.00fF
C23881 PAND2X1_243/CTRL PAND2X1_338/B 0.03fF
C23882 PAND2X1_653/O PAND2X1_557/A 0.02fF
C23883 POR2X1_96/A POR2X1_533/CTRL2 0.02fF
C23884 POR2X1_51/B POR2X1_587/a_56_344# 0.00fF
C23885 VDD POR2X1_620/B 0.23fF
C23886 PAND2X1_79/Y PAND2X1_111/B 0.03fF
C23887 POR2X1_132/Y PAND2X1_140/A 0.01fF
C23888 POR2X1_323/a_16_28# POR2X1_110/Y 0.02fF
C23889 PAND2X1_718/Y POR2X1_77/Y 0.01fF
C23890 POR2X1_845/CTRL2 POR2X1_532/A 0.03fF
C23891 POR2X1_565/a_16_28# POR2X1_550/Y 0.03fF
C23892 POR2X1_851/CTRL2 POR2X1_733/A 0.05fF
C23893 POR2X1_396/Y POR2X1_395/Y 0.16fF
C23894 POR2X1_482/Y POR2X1_77/Y 0.08fF
C23895 VDD PAND2X1_101/B 0.13fF
C23896 POR2X1_41/B POR2X1_144/O 0.05fF
C23897 PAND2X1_63/Y POR2X1_569/A 0.10fF
C23898 POR2X1_455/A POR2X1_456/B 0.01fF
C23899 PAND2X1_589/m4_208_n4# PAND2X1_142/m4_208_n4# 0.13fF
C23900 POR2X1_327/Y PAND2X1_90/A 0.03fF
C23901 POR2X1_294/A POR2X1_121/Y 0.03fF
C23902 D_INPUT_2 POR2X1_4/O 0.02fF
C23903 POR2X1_416/B POR2X1_609/O 0.03fF
C23904 POR2X1_447/B POR2X1_192/Y 0.05fF
C23905 PAND2X1_115/a_16_344# PAND2X1_853/B 0.01fF
C23906 PAND2X1_96/B POR2X1_259/O 0.02fF
C23907 POR2X1_170/B POR2X1_192/B 0.38fF
C23908 POR2X1_57/A POR2X1_315/Y 0.07fF
C23909 PAND2X1_499/CTRL POR2X1_39/B 0.01fF
C23910 POR2X1_390/B POR2X1_335/Y 0.00fF
C23911 POR2X1_673/Y D_INPUT_1 0.10fF
C23912 POR2X1_790/A POR2X1_753/CTRL 0.04fF
C23913 POR2X1_68/B POR2X1_249/Y 0.02fF
C23914 PAND2X1_843/CTRL2 POR2X1_251/Y 0.01fF
C23915 PAND2X1_71/a_16_344# PAND2X1_71/Y 0.01fF
C23916 POR2X1_205/A POR2X1_101/Y 0.10fF
C23917 PAND2X1_659/Y PAND2X1_215/B 0.07fF
C23918 PAND2X1_213/Y PAND2X1_569/B 0.07fF
C23919 PAND2X1_226/CTRL2 POR2X1_191/Y 0.00fF
C23920 PAND2X1_226/O POR2X1_192/B 0.21fF
C23921 POR2X1_7/A PAND2X1_549/B 0.07fF
C23922 PAND2X1_148/a_76_28# POR2X1_145/Y 0.04fF
C23923 POR2X1_60/Y PAND2X1_351/A 0.01fF
C23924 POR2X1_16/A POR2X1_38/Y 0.27fF
C23925 POR2X1_416/B PAND2X1_805/A 0.03fF
C23926 POR2X1_540/O POR2X1_703/A 0.01fF
C23927 POR2X1_106/Y POR2X1_77/Y 0.02fF
C23928 POR2X1_52/A POR2X1_613/Y 0.04fF
C23929 POR2X1_616/Y PAND2X1_790/Y 0.03fF
C23930 PAND2X1_6/A POR2X1_129/Y 0.09fF
C23931 POR2X1_41/B PAND2X1_857/O 0.06fF
C23932 PAND2X1_717/Y PAND2X1_656/A 0.06fF
C23933 PAND2X1_8/Y PAND2X1_102/CTRL2 0.03fF
C23934 PAND2X1_496/a_16_344# POR2X1_294/A 0.02fF
C23935 POR2X1_529/Y PAND2X1_510/B 0.02fF
C23936 POR2X1_285/B POR2X1_285/CTRL 0.00fF
C23937 POR2X1_7/B POR2X1_767/a_16_28# 0.01fF
C23938 POR2X1_648/A POR2X1_644/Y 0.02fF
C23939 PAND2X1_865/Y PAND2X1_592/Y 0.07fF
C23940 PAND2X1_218/a_76_28# PAND2X1_853/B 0.02fF
C23941 POR2X1_216/a_16_28# POR2X1_101/Y -0.00fF
C23942 POR2X1_216/a_76_344# POR2X1_116/Y 0.00fF
C23943 POR2X1_334/Y PAND2X1_69/A 0.03fF
C23944 POR2X1_158/Y PAND2X1_210/O 0.02fF
C23945 PAND2X1_61/Y PAND2X1_332/Y 0.02fF
C23946 POR2X1_83/Y PAND2X1_197/a_76_28# 0.03fF
C23947 PAND2X1_580/B POR2X1_77/Y 0.03fF
C23948 PAND2X1_812/A PAND2X1_812/O 0.05fF
C23949 PAND2X1_40/O PAND2X1_3/B 0.03fF
C23950 POR2X1_68/B POR2X1_571/m4_208_n4# 0.07fF
C23951 POR2X1_7/B PAND2X1_539/a_76_28# 0.01fF
C23952 POR2X1_126/CTRL2 POR2X1_411/B 0.01fF
C23953 PAND2X1_575/a_16_344# POR2X1_394/A 0.04fF
C23954 PAND2X1_809/B POR2X1_7/B 0.03fF
C23955 POR2X1_569/A POR2X1_260/A 0.07fF
C23956 POR2X1_620/B PAND2X1_32/B 0.03fF
C23957 POR2X1_244/Y POR2X1_575/O 0.01fF
C23958 PAND2X1_819/CTRL POR2X1_260/A 0.00fF
C23959 POR2X1_96/Y PAND2X1_6/A 0.07fF
C23960 PAND2X1_467/Y PAND2X1_726/B 0.07fF
C23961 POR2X1_274/A POR2X1_556/A 0.03fF
C23962 PAND2X1_246/CTRL POR2X1_66/A 0.03fF
C23963 POR2X1_711/B POR2X1_532/A 0.02fF
C23964 PAND2X1_593/Y PAND2X1_537/O 0.04fF
C23965 PAND2X1_550/Y POR2X1_394/A 0.05fF
C23966 PAND2X1_454/CTRL POR2X1_77/Y 0.00fF
C23967 POR2X1_387/Y PAND2X1_156/A 0.10fF
C23968 POR2X1_677/Y POR2X1_72/B 0.00fF
C23969 PAND2X1_437/CTRL POR2X1_186/Y 0.03fF
C23970 PAND2X1_717/A POR2X1_32/A 0.36fF
C23971 POR2X1_16/A INPUT_1 0.06fF
C23972 PAND2X1_109/CTRL D_GATE_222 0.06fF
C23973 POR2X1_57/A PAND2X1_737/CTRL 0.01fF
C23974 PAND2X1_779/CTRL2 POR2X1_527/Y 0.01fF
C23975 PAND2X1_134/O PAND2X1_32/B 0.17fF
C23976 POR2X1_814/A PAND2X1_58/A 0.07fF
C23977 PAND2X1_23/Y POR2X1_509/CTRL2 0.04fF
C23978 POR2X1_567/A POR2X1_736/O 0.03fF
C23979 POR2X1_166/CTRL2 PAND2X1_326/B 0.01fF
C23980 POR2X1_84/A PAND2X1_39/B 0.07fF
C23981 POR2X1_833/A POR2X1_244/Y 0.46fF
C23982 POR2X1_16/A POR2X1_153/Y 0.17fF
C23983 PAND2X1_69/A POR2X1_343/CTRL 0.02fF
C23984 PAND2X1_547/O POR2X1_39/B 0.15fF
C23985 PAND2X1_349/A PAND2X1_141/CTRL 0.01fF
C23986 POR2X1_815/Y POR2X1_816/Y 0.19fF
C23987 POR2X1_417/Y PAND2X1_717/A 0.03fF
C23988 PAND2X1_761/CTRL D_INPUT_0 0.00fF
C23989 POR2X1_564/O POR2X1_180/A 0.02fF
C23990 POR2X1_411/B POR2X1_268/CTRL 0.01fF
C23991 PAND2X1_337/A POR2X1_77/Y 0.03fF
C23992 POR2X1_846/Y PAND2X1_58/A 0.03fF
C23993 POR2X1_556/A POR2X1_269/A 0.21fF
C23994 POR2X1_48/A POR2X1_24/Y 0.06fF
C23995 POR2X1_43/Y POR2X1_42/Y 0.03fF
C23996 POR2X1_20/B POR2X1_67/A 0.14fF
C23997 PAND2X1_23/Y PAND2X1_135/CTRL 0.01fF
C23998 PAND2X1_26/O D_INPUT_4 0.17fF
C23999 POR2X1_42/Y POR2X1_589/Y 0.02fF
C24000 POR2X1_78/Y POR2X1_267/A 0.13fF
C24001 POR2X1_411/B POR2X1_516/Y 0.03fF
C24002 INPUT_3 POR2X1_819/O 0.06fF
C24003 PAND2X1_848/O INPUT_3 0.04fF
C24004 POR2X1_270/Y POR2X1_222/a_16_28# 0.02fF
C24005 POR2X1_836/B POR2X1_776/A 0.01fF
C24006 PAND2X1_88/Y POR2X1_555/O 0.01fF
C24007 POR2X1_554/a_16_28# POR2X1_228/Y 0.08fF
C24008 POR2X1_634/A POR2X1_859/O 0.01fF
C24009 POR2X1_440/a_56_344# POR2X1_192/Y 0.00fF
C24010 POR2X1_362/Y PAND2X1_39/B 0.06fF
C24011 PAND2X1_404/Y POR2X1_609/Y 0.02fF
C24012 PAND2X1_295/CTRL2 POR2X1_296/B 0.00fF
C24013 PAND2X1_63/Y PAND2X1_72/A 0.32fF
C24014 POR2X1_657/CTRL2 POR2X1_446/B 0.01fF
C24015 POR2X1_644/a_76_344# D_INPUT_0 0.01fF
C24016 PAND2X1_628/CTRL2 POR2X1_785/A 0.01fF
C24017 PAND2X1_639/B POR2X1_386/Y 0.01fF
C24018 POR2X1_48/A POR2X1_626/CTRL 0.01fF
C24019 POR2X1_606/CTRL2 POR2X1_121/B 0.03fF
C24020 POR2X1_751/Y POR2X1_4/Y 0.03fF
C24021 PAND2X1_434/CTRL2 POR2X1_39/B 0.11fF
C24022 POR2X1_590/A POR2X1_454/A 0.01fF
C24023 POR2X1_86/Y PAND2X1_99/Y 0.57fF
C24024 POR2X1_119/Y POR2X1_129/Y 0.03fF
C24025 PAND2X1_349/A POR2X1_77/Y 0.03fF
C24026 PAND2X1_63/B POR2X1_77/Y 0.14fF
C24027 POR2X1_263/Y POR2X1_37/Y 0.04fF
C24028 POR2X1_730/Y POR2X1_568/B 0.05fF
C24029 POR2X1_97/A POR2X1_856/B 0.03fF
C24030 PAND2X1_480/B POR2X1_329/A 0.01fF
C24031 PAND2X1_309/CTRL2 POR2X1_814/A 0.00fF
C24032 POR2X1_18/CTRL2 INPUT_4 0.01fF
C24033 POR2X1_416/B PAND2X1_569/B 0.07fF
C24034 POR2X1_864/A POR2X1_780/m4_208_n4# 0.12fF
C24035 POR2X1_416/B POR2X1_158/B 7.70fF
C24036 PAND2X1_415/O POR2X1_414/Y 0.18fF
C24037 PAND2X1_20/A POR2X1_84/A 0.01fF
C24038 PAND2X1_319/CTRL POR2X1_20/B 0.01fF
C24039 POR2X1_119/Y PAND2X1_659/Y 0.07fF
C24040 POR2X1_607/A POR2X1_612/Y 0.10fF
C24041 PAND2X1_640/B POR2X1_102/Y 0.01fF
C24042 PAND2X1_865/Y POR2X1_767/CTRL2 0.00fF
C24043 PAND2X1_39/B PAND2X1_65/Y 0.10fF
C24044 POR2X1_43/B POR2X1_827/CTRL2 0.01fF
C24045 POR2X1_66/B POR2X1_558/B 0.03fF
C24046 POR2X1_137/B VDD 0.07fF
C24047 PAND2X1_436/a_16_344# PAND2X1_390/Y 0.01fF
C24048 PAND2X1_493/O POR2X1_492/Y 0.00fF
C24049 POR2X1_654/B POR2X1_260/B 0.03fF
C24050 PAND2X1_797/Y PAND2X1_714/B 0.04fF
C24051 PAND2X1_200/CTRL2 POR2X1_32/A 0.01fF
C24052 PAND2X1_88/CTRL POR2X1_66/A 0.01fF
C24053 INPUT_3 VDD 4.38fF
C24054 POR2X1_666/CTRL POR2X1_102/Y 0.01fF
C24055 PAND2X1_72/A POR2X1_260/A 2.07fF
C24056 PAND2X1_87/CTRL2 PAND2X1_6/A 0.06fF
C24057 POR2X1_846/Y POR2X1_790/a_56_344# 0.00fF
C24058 POR2X1_814/B POR2X1_84/A 0.07fF
C24059 POR2X1_78/A POR2X1_605/CTRL2 0.03fF
C24060 POR2X1_850/A POR2X1_260/B 0.03fF
C24061 POR2X1_383/CTRL POR2X1_383/Y 0.01fF
C24062 POR2X1_149/A POR2X1_78/A 0.00fF
C24063 PAND2X1_717/A POR2X1_184/Y 0.03fF
C24064 POR2X1_66/B PAND2X1_413/O 0.15fF
C24065 POR2X1_3/A PAND2X1_635/Y 0.01fF
C24066 PAND2X1_73/Y PAND2X1_74/CTRL2 0.01fF
C24067 PAND2X1_108/a_16_344# PAND2X1_39/B 0.01fF
C24068 POR2X1_428/Y VDD 0.43fF
C24069 POR2X1_446/A POR2X1_192/Y 0.03fF
C24070 POR2X1_66/A PAND2X1_41/B 1.87fF
C24071 PAND2X1_26/A PAND2X1_587/Y 0.03fF
C24072 PAND2X1_96/B POR2X1_814/A 0.19fF
C24073 PAND2X1_142/O PAND2X1_72/A 0.03fF
C24074 POR2X1_88/O INPUT_0 0.06fF
C24075 POR2X1_102/Y POR2X1_272/CTRL2 0.01fF
C24076 POR2X1_681/Y POR2X1_682/Y 0.09fF
C24077 POR2X1_93/Y VDD 0.09fF
C24078 PAND2X1_205/A PAND2X1_84/Y 0.00fF
C24079 POR2X1_502/A POR2X1_602/CTRL 0.01fF
C24080 PAND2X1_93/B VDD 1.69fF
C24081 POR2X1_456/m4_208_n4# POR2X1_66/A 0.08fF
C24082 D_INPUT_0 PAND2X1_332/a_16_344# 0.02fF
C24083 PAND2X1_402/CTRL POR2X1_14/Y 0.01fF
C24084 POR2X1_257/A PAND2X1_254/O 0.02fF
C24085 POR2X1_121/B POR2X1_389/Y 0.01fF
C24086 POR2X1_852/B PAND2X1_58/A 0.00fF
C24087 PAND2X1_58/A PAND2X1_55/CTRL2 0.00fF
C24088 PAND2X1_571/CTRL PAND2X1_571/Y 0.01fF
C24089 POR2X1_634/CTRL2 PAND2X1_41/B 0.01fF
C24090 POR2X1_406/Y POR2X1_263/Y 0.00fF
C24091 POR2X1_20/B PAND2X1_642/B 0.03fF
C24092 POR2X1_402/B POR2X1_66/A 0.01fF
C24093 POR2X1_65/A POR2X1_667/A 0.06fF
C24094 POR2X1_262/Y PAND2X1_716/a_16_344# 0.02fF
C24095 POR2X1_440/CTRL POR2X1_353/A 0.02fF
C24096 POR2X1_23/Y POR2X1_252/CTRL2 -0.00fF
C24097 POR2X1_143/CTRL2 D_INPUT_0 0.01fF
C24098 POR2X1_137/B PAND2X1_32/B 0.31fF
C24099 POR2X1_316/Y POR2X1_416/B 0.03fF
C24100 POR2X1_39/CTRL POR2X1_40/Y 0.01fF
C24101 PAND2X1_9/Y D_INPUT_1 0.03fF
C24102 POR2X1_43/CTRL2 POR2X1_77/Y 0.07fF
C24103 POR2X1_669/B POR2X1_516/B 0.03fF
C24104 POR2X1_78/A VDD 3.85fF
C24105 POR2X1_614/A POR2X1_266/CTRL2 0.05fF
C24106 PAND2X1_209/A POR2X1_257/A 1.92fF
C24107 PAND2X1_60/a_56_28# POR2X1_35/Y 0.00fF
C24108 POR2X1_263/Y POR2X1_293/Y 0.03fF
C24109 POR2X1_671/m4_208_n4# POR2X1_37/Y 0.01fF
C24110 PAND2X1_438/O POR2X1_544/B 0.01fF
C24111 POR2X1_725/CTRL2 POR2X1_711/Y 0.01fF
C24112 POR2X1_72/B PAND2X1_736/CTRL2 0.01fF
C24113 PAND2X1_244/B PAND2X1_97/Y 0.03fF
C24114 POR2X1_814/A PAND2X1_503/CTRL 0.06fF
C24115 PAND2X1_52/B POR2X1_182/a_16_28# 0.00fF
C24116 POR2X1_185/O POR2X1_260/B 0.02fF
C24117 POR2X1_856/B POR2X1_294/B 0.12fF
C24118 POR2X1_366/Y POR2X1_856/B 0.10fF
C24119 PAND2X1_60/CTRL PAND2X1_69/A 0.01fF
C24120 PAND2X1_23/Y POR2X1_476/A 0.07fF
C24121 PAND2X1_149/O POR2X1_669/B 0.03fF
C24122 PAND2X1_93/B POR2X1_741/Y 0.11fF
C24123 POR2X1_41/B POR2X1_32/A 0.22fF
C24124 POR2X1_614/A POR2X1_450/Y 0.04fF
C24125 POR2X1_853/A POR2X1_567/B 0.05fF
C24126 POR2X1_72/B PAND2X1_513/a_76_28# 0.02fF
C24127 PAND2X1_58/A POR2X1_401/B 0.01fF
C24128 POR2X1_337/a_16_28# POR2X1_270/Y 0.01fF
C24129 PAND2X1_602/Y POR2X1_48/A 0.51fF
C24130 POR2X1_119/Y PAND2X1_403/CTRL2 0.01fF
C24131 POR2X1_360/A POR2X1_590/A 0.03fF
C24132 POR2X1_814/B PAND2X1_65/Y 0.03fF
C24133 PAND2X1_73/Y POR2X1_465/B 0.01fF
C24134 POR2X1_477/A POR2X1_434/A 0.59fF
C24135 POR2X1_49/Y POR2X1_144/Y 0.01fF
C24136 POR2X1_83/B PAND2X1_435/a_16_344# 0.01fF
C24137 POR2X1_83/B PAND2X1_182/A 0.01fF
C24138 POR2X1_25/Y PAND2X1_635/Y 0.02fF
C24139 PAND2X1_104/O PAND2X1_8/Y 0.13fF
C24140 POR2X1_60/A POR2X1_79/Y 0.03fF
C24141 POR2X1_66/B POR2X1_332/B 0.15fF
C24142 PAND2X1_830/Y POR2X1_102/Y 0.03fF
C24143 PAND2X1_793/CTRL PAND2X1_793/A 0.01fF
C24144 POR2X1_29/A PAND2X1_375/O 0.01fF
C24145 PAND2X1_205/Y PAND2X1_473/B 0.12fF
C24146 PAND2X1_58/A INPUT_5 0.02fF
C24147 PAND2X1_13/m4_208_n4# POR2X1_750/B 0.03fF
C24148 POR2X1_818/Y POR2X1_816/A 0.03fF
C24149 POR2X1_102/Y POR2X1_7/B 2.62fF
C24150 POR2X1_150/Y PAND2X1_175/CTRL 0.00fF
C24151 POR2X1_750/B INPUT_0 0.02fF
C24152 POR2X1_814/B PAND2X1_54/CTRL 0.08fF
C24153 POR2X1_307/O POR2X1_513/B 0.00fF
C24154 POR2X1_20/B PAND2X1_550/B 0.03fF
C24155 PAND2X1_93/B PAND2X1_32/B 0.13fF
C24156 PAND2X1_6/A POR2X1_37/Y 0.01fF
C24157 POR2X1_864/A POR2X1_598/O 0.00fF
C24158 POR2X1_278/Y POR2X1_72/B 0.12fF
C24159 PAND2X1_840/A POR2X1_496/Y 0.00fF
C24160 POR2X1_41/B POR2X1_417/Y 0.20fF
C24161 POR2X1_94/m4_208_n4# POR2X1_23/Y 0.07fF
C24162 POR2X1_223/CTRL2 POR2X1_186/Y 0.01fF
C24163 PAND2X1_56/Y POR2X1_657/CTRL2 0.13fF
C24164 PAND2X1_771/Y POR2X1_73/Y 1.69fF
C24165 PAND2X1_572/O PAND2X1_267/Y -0.00fF
C24166 POR2X1_78/A POR2X1_741/Y 0.03fF
C24167 PAND2X1_318/CTRL POR2X1_417/Y 0.01fF
C24168 POR2X1_420/a_56_344# POR2X1_90/Y 0.00fF
C24169 POR2X1_13/A PAND2X1_61/Y 0.02fF
C24170 POR2X1_573/CTRL VDD 0.00fF
C24171 PAND2X1_798/B PAND2X1_794/CTRL 0.01fF
C24172 POR2X1_241/B POR2X1_35/Y 0.03fF
C24173 D_INPUT_2 POR2X1_37/CTRL2 0.03fF
C24174 PAND2X1_834/CTRL2 POR2X1_677/Y 0.03fF
C24175 PAND2X1_340/CTRL POR2X1_88/Y 0.01fF
C24176 POR2X1_673/Y INPUT_3 0.15fF
C24177 PAND2X1_93/B PAND2X1_312/O 0.05fF
C24178 POR2X1_407/A POR2X1_656/a_76_344# 0.01fF
C24179 POR2X1_97/A POR2X1_577/CTRL 0.00fF
C24180 POR2X1_502/A POR2X1_640/m4_208_n4# 0.06fF
C24181 POR2X1_164/CTRL2 POR2X1_83/B 0.03fF
C24182 PAND2X1_41/B POR2X1_792/B 0.05fF
C24183 POR2X1_804/A POR2X1_296/B 0.05fF
C24184 POR2X1_865/B POR2X1_218/Y 0.09fF
C24185 POR2X1_250/A PAND2X1_364/B 0.07fF
C24186 PAND2X1_612/B POR2X1_773/CTRL2 0.00fF
C24187 POR2X1_859/CTRL POR2X1_559/A 0.03fF
C24188 PAND2X1_69/O POR2X1_296/B 0.17fF
C24189 POR2X1_707/B PAND2X1_587/CTRL2 0.02fF
C24190 PAND2X1_477/B POR2X1_102/Y 0.88fF
C24191 POR2X1_377/CTRL POR2X1_94/A 0.01fF
C24192 PAND2X1_740/Y VDD 0.35fF
C24193 POR2X1_78/A PAND2X1_32/B 1.06fF
C24194 POR2X1_13/A PAND2X1_778/O 0.15fF
C24195 POR2X1_654/B PAND2X1_55/Y 0.07fF
C24196 POR2X1_393/O VDD 0.00fF
C24197 PAND2X1_714/A PAND2X1_714/O -0.00fF
C24198 POR2X1_811/O POR2X1_780/B 0.04fF
C24199 PAND2X1_741/a_76_28# PAND2X1_473/B 0.02fF
C24200 PAND2X1_114/Y POR2X1_106/Y 0.15fF
C24201 POR2X1_38/B PAND2X1_531/O 0.24fF
C24202 PAND2X1_659/B PAND2X1_659/O 0.01fF
C24203 POR2X1_550/A POR2X1_66/A 0.03fF
C24204 POR2X1_222/Y PAND2X1_41/B 0.03fF
C24205 PAND2X1_217/B PAND2X1_469/B 0.02fF
C24206 PAND2X1_852/CTRL POR2X1_65/A 0.01fF
C24207 D_INPUT_0 POR2X1_513/a_16_28# 0.01fF
C24208 PAND2X1_778/CTRL POR2X1_293/Y 0.01fF
C24209 POR2X1_78/B POR2X1_231/CTRL 0.01fF
C24210 PAND2X1_243/B POR2X1_397/Y 0.03fF
C24211 POR2X1_504/Y POR2X1_43/B 0.03fF
C24212 PAND2X1_641/Y PAND2X1_404/Y 0.12fF
C24213 PAND2X1_787/Y PAND2X1_724/B 0.02fF
C24214 PAND2X1_575/B POR2X1_73/Y 0.01fF
C24215 POR2X1_677/O PAND2X1_658/B 0.21fF
C24216 PAND2X1_650/a_76_28# D_INPUT_0 0.01fF
C24217 POR2X1_446/B POR2X1_574/Y 0.00fF
C24218 POR2X1_389/CTRL POR2X1_480/A 0.00fF
C24219 PAND2X1_607/O PAND2X1_56/A 0.02fF
C24220 PAND2X1_47/B INPUT_6 0.04fF
C24221 POR2X1_192/Y POR2X1_220/Y 0.07fF
C24222 PAND2X1_94/A PAND2X1_94/O 0.05fF
C24223 POR2X1_529/Y POR2X1_29/A 0.01fF
C24224 POR2X1_236/Y POR2X1_395/O 0.01fF
C24225 POR2X1_330/Y PAND2X1_311/CTRL2 0.13fF
C24226 INPUT_1 PAND2X1_637/O 0.03fF
C24227 POR2X1_48/A PAND2X1_155/O 0.01fF
C24228 PAND2X1_9/Y POR2X1_620/B 0.03fF
C24229 PAND2X1_250/CTRL2 PAND2X1_69/A 0.02fF
C24230 POR2X1_616/Y POR2X1_20/B 0.04fF
C24231 POR2X1_108/a_16_28# POR2X1_102/Y 0.02fF
C24232 POR2X1_669/B PAND2X1_550/Y 0.03fF
C24233 D_INPUT_5 POR2X1_3/B 0.04fF
C24234 PAND2X1_862/B PAND2X1_793/Y 0.03fF
C24235 POR2X1_406/Y PAND2X1_215/B 0.03fF
C24236 POR2X1_615/O PAND2X1_6/A 0.09fF
C24237 PAND2X1_804/B POR2X1_46/Y 0.02fF
C24238 PAND2X1_88/O POR2X1_68/B 0.05fF
C24239 POR2X1_41/B PAND2X1_35/Y 6.76fF
C24240 POR2X1_283/A POR2X1_226/CTRL2 0.05fF
C24241 POR2X1_49/Y PAND2X1_209/A 0.01fF
C24242 POR2X1_83/B POR2X1_283/A 0.06fF
C24243 POR2X1_66/A POR2X1_721/CTRL 0.09fF
C24244 PAND2X1_96/B POR2X1_852/B 0.01fF
C24245 POR2X1_100/O POR2X1_99/A 0.01fF
C24246 POR2X1_567/A POR2X1_776/A 0.32fF
C24247 POR2X1_267/a_16_28# POR2X1_318/A 0.08fF
C24248 POR2X1_853/CTRL2 POR2X1_785/A 0.00fF
C24249 POR2X1_341/A PAND2X1_323/CTRL 0.07fF
C24250 POR2X1_532/A PAND2X1_41/B 0.58fF
C24251 POR2X1_475/A PAND2X1_69/A 0.12fF
C24252 POR2X1_13/A PAND2X1_784/O 0.15fF
C24253 POR2X1_722/B POR2X1_722/Y 0.37fF
C24254 POR2X1_556/A PAND2X1_134/a_16_344# 0.03fF
C24255 PAND2X1_803/Y PAND2X1_360/a_16_344# 0.02fF
C24256 POR2X1_708/CTRL2 POR2X1_779/A 0.01fF
C24257 POR2X1_78/B PAND2X1_81/CTRL2 0.04fF
C24258 PAND2X1_675/A VDD 0.77fF
C24259 POR2X1_294/B POR2X1_722/Y 0.01fF
C24260 POR2X1_16/A PAND2X1_794/CTRL2 0.01fF
C24261 PAND2X1_469/B VDD 2.29fF
C24262 PAND2X1_253/O POR2X1_78/A 0.02fF
C24263 POR2X1_510/A VDD 0.00fF
C24264 POR2X1_14/Y POR2X1_754/CTRL2 0.03fF
C24265 POR2X1_73/CTRL2 POR2X1_40/Y 0.02fF
C24266 POR2X1_673/Y POR2X1_78/A 0.03fF
C24267 PAND2X1_23/O PAND2X1_60/B 0.02fF
C24268 POR2X1_41/B POR2X1_189/Y 0.06fF
C24269 PAND2X1_629/CTRL2 POR2X1_7/A 0.03fF
C24270 POR2X1_32/A PAND2X1_308/Y 0.03fF
C24271 POR2X1_13/A POR2X1_669/A 0.01fF
C24272 POR2X1_95/O POR2X1_12/A 0.01fF
C24273 PAND2X1_808/Y POR2X1_7/B 0.03fF
C24274 POR2X1_383/A POR2X1_389/Y 0.03fF
C24275 POR2X1_344/O POR2X1_383/A 0.07fF
C24276 POR2X1_278/A POR2X1_278/O 0.12fF
C24277 POR2X1_857/B POR2X1_350/CTRL2 0.04fF
C24278 POR2X1_357/O POR2X1_220/B 0.00fF
C24279 POR2X1_41/B POR2X1_184/Y 0.08fF
C24280 POR2X1_186/Y POR2X1_181/B 0.06fF
C24281 POR2X1_43/B POR2X1_586/O 0.01fF
C24282 POR2X1_83/B POR2X1_385/a_16_28# 0.03fF
C24283 POR2X1_23/Y PAND2X1_851/O 0.08fF
C24284 POR2X1_463/Y POR2X1_634/A 0.03fF
C24285 POR2X1_208/A POR2X1_61/Y 0.06fF
C24286 POR2X1_775/A POR2X1_579/Y 0.03fF
C24287 PAND2X1_293/CTRL POR2X1_68/B 0.04fF
C24288 POR2X1_163/Y PAND2X1_725/CTRL 0.01fF
C24289 PAND2X1_309/O POR2X1_68/A 0.05fF
C24290 POR2X1_66/B POR2X1_768/CTRL 0.00fF
C24291 PAND2X1_658/A POR2X1_42/Y 0.05fF
C24292 POR2X1_227/A PAND2X1_52/B 0.00fF
C24293 PAND2X1_480/B PAND2X1_702/CTRL 0.25fF
C24294 POR2X1_842/a_16_28# POR2X1_737/A 0.02fF
C24295 POR2X1_333/A PAND2X1_745/O 0.06fF
C24296 POR2X1_41/B PAND2X1_651/Y 0.14fF
C24297 POR2X1_605/A POR2X1_220/Y 0.00fF
C24298 PAND2X1_6/A POR2X1_293/Y 0.21fF
C24299 PAND2X1_116/O POR2X1_283/A 0.01fF
C24300 POR2X1_567/A POR2X1_856/B 0.02fF
C24301 POR2X1_119/Y POR2X1_37/Y 0.12fF
C24302 POR2X1_119/Y POR2X1_271/a_16_28# 0.04fF
C24303 INPUT_1 POR2X1_495/O 0.02fF
C24304 POR2X1_185/O PAND2X1_55/Y 0.04fF
C24305 POR2X1_66/A PAND2X1_143/CTRL 0.03fF
C24306 POR2X1_294/B POR2X1_565/O 0.18fF
C24307 INPUT_7 PAND2X1_1/O 0.00fF
C24308 POR2X1_417/Y PAND2X1_308/Y 0.02fF
C24309 POR2X1_13/A PAND2X1_555/Y 0.02fF
C24310 POR2X1_358/O POR2X1_350/Y 0.00fF
C24311 POR2X1_8/Y PAND2X1_35/B 0.05fF
C24312 POR2X1_41/B PAND2X1_243/CTRL 0.00fF
C24313 POR2X1_81/a_76_344# POR2X1_153/Y 0.03fF
C24314 POR2X1_62/CTRL PAND2X1_6/A 0.01fF
C24315 PAND2X1_407/a_16_344# POR2X1_39/B 0.04fF
C24316 POR2X1_193/A POR2X1_112/Y 0.03fF
C24317 POR2X1_97/A POR2X1_191/Y 0.05fF
C24318 PAND2X1_8/Y PAND2X1_670/O 0.04fF
C24319 PAND2X1_132/CTRL PAND2X1_32/B 0.01fF
C24320 POR2X1_416/B POR2X1_54/Y 0.07fF
C24321 POR2X1_579/Y POR2X1_112/Y 0.05fF
C24322 POR2X1_71/Y POR2X1_73/Y 0.00fF
C24323 POR2X1_480/A POR2X1_590/O 0.04fF
C24324 POR2X1_590/A POR2X1_571/Y 0.03fF
C24325 POR2X1_283/A PAND2X1_140/Y 0.03fF
C24326 POR2X1_629/A PAND2X1_69/A 0.01fF
C24327 PAND2X1_23/Y POR2X1_513/Y 0.03fF
C24328 POR2X1_865/O POR2X1_784/A 0.01fF
C24329 PAND2X1_73/Y POR2X1_557/O 0.34fF
C24330 POR2X1_614/A POR2X1_775/A 0.03fF
C24331 PAND2X1_496/O POR2X1_500/Y 0.15fF
C24332 POR2X1_140/B POR2X1_515/Y 0.00fF
C24333 POR2X1_42/Y POR2X1_73/Y 0.42fF
C24334 POR2X1_68/A POR2X1_790/A 0.02fF
C24335 PAND2X1_549/B POR2X1_372/m4_208_n4# 0.15fF
C24336 PAND2X1_665/O POR2X1_66/A 0.03fF
C24337 POR2X1_351/Y POR2X1_350/O 0.01fF
C24338 PAND2X1_220/Y PAND2X1_343/a_16_344# 0.04fF
C24339 POR2X1_647/B PAND2X1_52/B 0.00fF
C24340 POR2X1_89/O POR2X1_77/Y 0.00fF
C24341 PAND2X1_478/O POR2X1_90/Y 0.01fF
C24342 POR2X1_447/B PAND2X1_626/CTRL2 0.04fF
C24343 POR2X1_52/A PAND2X1_843/Y 0.03fF
C24344 PAND2X1_856/B VDD 0.01fF
C24345 POR2X1_78/B POR2X1_834/Y 0.10fF
C24346 PAND2X1_738/Y PAND2X1_569/B 0.10fF
C24347 INPUT_1 PAND2X1_54/O 0.01fF
C24348 PAND2X1_46/O PAND2X1_71/Y 0.02fF
C24349 POR2X1_606/a_76_344# PAND2X1_56/A 0.00fF
C24350 POR2X1_460/A POR2X1_460/B 0.16fF
C24351 POR2X1_57/A PAND2X1_398/CTRL 0.01fF
C24352 POR2X1_78/O POR2X1_844/B 0.01fF
C24353 POR2X1_532/A POR2X1_130/Y 1.24fF
C24354 PAND2X1_319/B POR2X1_312/CTRL2 0.05fF
C24355 PAND2X1_273/CTRL2 PAND2X1_60/B 0.03fF
C24356 POR2X1_341/A POR2X1_579/a_56_344# 0.01fF
C24357 POR2X1_65/A PAND2X1_170/O 0.01fF
C24358 POR2X1_547/a_16_28# POR2X1_614/A 0.06fF
C24359 POR2X1_652/Y POR2X1_799/CTRL2 0.03fF
C24360 POR2X1_376/B PAND2X1_708/CTRL 0.01fF
C24361 POR2X1_425/CTRL POR2X1_158/B 0.01fF
C24362 POR2X1_614/A POR2X1_112/Y 0.07fF
C24363 PAND2X1_69/A PAND2X1_146/a_76_28# 0.01fF
C24364 PAND2X1_556/B PAND2X1_726/B 0.03fF
C24365 POR2X1_68/A PAND2X1_88/Y 0.03fF
C24366 POR2X1_61/Y PAND2X1_394/CTRL2 0.05fF
C24367 PAND2X1_56/Y POR2X1_318/A 0.10fF
C24368 POR2X1_179/CTRL2 POR2X1_387/Y 0.32fF
C24369 POR2X1_244/B POR2X1_260/A 0.03fF
C24370 POR2X1_55/Y POR2X1_107/Y 0.00fF
C24371 PAND2X1_23/Y POR2X1_366/A 0.11fF
C24372 INPUT_1 PAND2X1_57/B 0.54fF
C24373 POR2X1_222/Y POR2X1_228/Y 0.07fF
C24374 PAND2X1_96/B POR2X1_190/CTRL2 0.01fF
C24375 PAND2X1_90/A PAND2X1_133/CTRL2 0.01fF
C24376 PAND2X1_674/O PAND2X1_60/B 0.20fF
C24377 POR2X1_145/m4_208_n4# PAND2X1_213/Y 0.01fF
C24378 PAND2X1_23/Y PAND2X1_373/CTRL 0.01fF
C24379 POR2X1_32/A POR2X1_77/Y 0.15fF
C24380 POR2X1_334/CTRL POR2X1_404/Y 0.17fF
C24381 POR2X1_208/A POR2X1_35/Y 0.01fF
C24382 PAND2X1_631/A PAND2X1_456/CTRL 0.02fF
C24383 PAND2X1_6/A POR2X1_408/Y 0.22fF
C24384 PAND2X1_659/Y PAND2X1_204/CTRL2 0.00fF
C24385 POR2X1_848/A POR2X1_90/CTRL2 0.05fF
C24386 PAND2X1_56/Y PAND2X1_306/m4_208_n4# 0.06fF
C24387 POR2X1_470/CTRL2 PAND2X1_52/B 0.04fF
C24388 POR2X1_85/Y POR2X1_32/A 0.02fF
C24389 PAND2X1_126/CTRL PAND2X1_6/A 0.00fF
C24390 POR2X1_56/Y PAND2X1_656/A 0.00fF
C24391 PAND2X1_173/CTRL PAND2X1_32/B 0.01fF
C24392 POR2X1_137/Y POR2X1_501/B 0.03fF
C24393 POR2X1_614/A POR2X1_162/Y 0.00fF
C24394 PAND2X1_467/CTRL PAND2X1_725/A 0.00fF
C24395 PAND2X1_115/Y PAND2X1_348/A 0.03fF
C24396 PAND2X1_55/Y POR2X1_576/O 0.02fF
C24397 PAND2X1_467/Y POR2X1_43/B 0.03fF
C24398 POR2X1_3/A POR2X1_36/B 0.28fF
C24399 POR2X1_532/A POR2X1_228/Y 0.03fF
C24400 POR2X1_575/CTRL POR2X1_573/A 0.01fF
C24401 POR2X1_294/B POR2X1_244/Y 0.03fF
C24402 POR2X1_416/B PAND2X1_784/A 0.03fF
C24403 POR2X1_287/B POR2X1_343/CTRL2 0.01fF
C24404 PAND2X1_308/Y PAND2X1_302/CTRL 0.01fF
C24405 POR2X1_119/Y POR2X1_406/Y 0.31fF
C24406 POR2X1_13/A PAND2X1_141/CTRL2 0.01fF
C24407 POR2X1_417/Y POR2X1_77/Y 0.08fF
C24408 POR2X1_550/A POR2X1_532/A 0.03fF
C24409 POR2X1_477/A POR2X1_544/B 0.13fF
C24410 PAND2X1_281/O POR2X1_121/Y 0.04fF
C24411 POR2X1_674/Y POR2X1_331/O 0.01fF
C24412 PAND2X1_793/Y PAND2X1_716/B 0.03fF
C24413 POR2X1_113/O POR2X1_113/Y 0.00fF
C24414 POR2X1_489/A POR2X1_294/A 0.03fF
C24415 POR2X1_383/A POR2X1_318/A 0.07fF
C24416 POR2X1_670/CTRL2 POR2X1_77/Y 0.03fF
C24417 POR2X1_576/CTRL2 POR2X1_500/Y 0.00fF
C24418 PAND2X1_661/O PAND2X1_659/Y 0.01fF
C24419 POR2X1_816/A POR2X1_171/a_76_344# 0.00fF
C24420 POR2X1_461/A PAND2X1_52/B 0.00fF
C24421 POR2X1_502/Y POR2X1_776/B 3.86fF
C24422 POR2X1_235/CTRL2 POR2X1_7/A 0.02fF
C24423 POR2X1_366/CTRL2 PAND2X1_60/B 0.03fF
C24424 POR2X1_796/A PAND2X1_60/B 0.03fF
C24425 POR2X1_119/Y POR2X1_293/Y 0.80fF
C24426 POR2X1_751/Y POR2X1_816/A 0.95fF
C24427 VDD POR2X1_365/O 0.00fF
C24428 POR2X1_316/a_56_344# POR2X1_43/B 0.00fF
C24429 POR2X1_16/A POR2X1_591/Y 0.22fF
C24430 POR2X1_833/A PAND2X1_150/CTRL2 0.03fF
C24431 POR2X1_264/Y PAND2X1_48/A 0.02fF
C24432 PAND2X1_206/B PAND2X1_340/B 0.00fF
C24433 PAND2X1_394/CTRL2 POR2X1_35/Y 0.01fF
C24434 POR2X1_493/B POR2X1_493/O 0.09fF
C24435 PAND2X1_48/B POR2X1_540/Y 0.08fF
C24436 POR2X1_661/Y POR2X1_661/A 0.02fF
C24437 PAND2X1_93/B PAND2X1_85/CTRL2 0.01fF
C24438 PAND2X1_824/B POR2X1_447/O 0.06fF
C24439 POR2X1_52/A PAND2X1_797/Y 0.03fF
C24440 POR2X1_556/A POR2X1_276/B 0.03fF
C24441 POR2X1_88/Y POR2X1_39/B 0.03fF
C24442 PAND2X1_55/Y PAND2X1_41/Y 0.00fF
C24443 POR2X1_568/Y POR2X1_577/Y 0.00fF
C24444 PAND2X1_96/B POR2X1_151/Y 0.05fF
C24445 POR2X1_228/O POR2X1_631/B 0.01fF
C24446 POR2X1_184/Y PAND2X1_141/CTRL 0.00fF
C24447 PAND2X1_6/Y POR2X1_349/CTRL 0.01fF
C24448 PAND2X1_803/Y PAND2X1_348/A 0.02fF
C24449 INPUT_3 PAND2X1_9/Y 0.05fF
C24450 POR2X1_244/Y PAND2X1_111/B 0.03fF
C24451 POR2X1_566/A POR2X1_736/A 0.05fF
C24452 POR2X1_16/A POR2X1_167/O 0.02fF
C24453 POR2X1_57/A POR2X1_373/Y 0.03fF
C24454 POR2X1_762/CTRL D_INPUT_6 0.02fF
C24455 PAND2X1_864/a_76_28# PAND2X1_568/B 0.02fF
C24456 POR2X1_592/a_16_28# POR2X1_592/A 0.05fF
C24457 PAND2X1_631/A POR2X1_56/Y 0.01fF
C24458 POR2X1_730/Y POR2X1_151/CTRL 0.01fF
C24459 PAND2X1_212/CTRL POR2X1_20/B 0.01fF
C24460 POR2X1_85/Y PAND2X1_35/Y 0.03fF
C24461 PAND2X1_527/CTRL2 PAND2X1_111/B 0.01fF
C24462 POR2X1_676/Y PAND2X1_52/B 0.02fF
C24463 PAND2X1_549/B POR2X1_153/Y 0.07fF
C24464 POR2X1_271/CTRL POR2X1_411/B 0.01fF
C24465 POR2X1_63/Y PAND2X1_404/Y 0.03fF
C24466 POR2X1_25/Y POR2X1_36/B 0.16fF
C24467 POR2X1_411/B PAND2X1_267/Y 0.06fF
C24468 PAND2X1_862/B PAND2X1_862/O 0.05fF
C24469 POR2X1_375/a_16_28# POR2X1_260/A 0.03fF
C24470 PAND2X1_608/CTRL2 POR2X1_102/Y 0.01fF
C24471 POR2X1_68/A POR2X1_568/B 0.07fF
C24472 POR2X1_270/O POR2X1_567/A 0.23fF
C24473 POR2X1_16/A PAND2X1_803/CTRL2 0.01fF
C24474 POR2X1_864/A D_INPUT_0 0.03fF
C24475 POR2X1_416/B POR2X1_13/Y 0.08fF
C24476 INPUT_1 PAND2X1_701/O 0.03fF
C24477 POR2X1_864/A POR2X1_811/A 2.06fF
C24478 POR2X1_445/A POR2X1_319/A 0.04fF
C24479 POR2X1_463/CTRL2 POR2X1_750/B 0.01fF
C24480 PAND2X1_73/Y POR2X1_688/CTRL 0.01fF
C24481 POR2X1_456/B POR2X1_741/A 0.01fF
C24482 PAND2X1_472/O POR2X1_153/Y 0.01fF
C24483 POR2X1_669/Y PAND2X1_721/B 0.03fF
C24484 PAND2X1_338/B PAND2X1_338/O 0.26fF
C24485 PAND2X1_269/CTRL POR2X1_72/B 0.00fF
C24486 PAND2X1_110/a_16_344# PAND2X1_52/B 0.06fF
C24487 POR2X1_513/Y POR2X1_711/Y 0.03fF
C24488 PAND2X1_651/Y POR2X1_77/Y 0.03fF
C24489 POR2X1_841/CTRL2 POR2X1_590/A 0.03fF
C24490 PAND2X1_634/CTRL2 POR2X1_607/A 0.00fF
C24491 POR2X1_23/Y PAND2X1_407/a_56_28# 0.00fF
C24492 POR2X1_490/Y PAND2X1_218/B 0.05fF
C24493 POR2X1_814/Y POR2X1_752/Y 0.01fF
C24494 POR2X1_709/A POR2X1_496/Y 0.08fF
C24495 D_GATE_662 POR2X1_568/A 0.07fF
C24496 POR2X1_499/A POR2X1_474/CTRL 0.00fF
C24497 POR2X1_78/A PAND2X1_9/Y 0.03fF
C24498 D_INPUT_5 PAND2X1_752/CTRL 0.01fF
C24499 POR2X1_416/B POR2X1_108/CTRL 0.01fF
C24500 POR2X1_66/A POR2X1_454/A 0.03fF
C24501 PAND2X1_417/O POR2X1_750/B 0.01fF
C24502 POR2X1_416/B PAND2X1_787/A 0.03fF
C24503 POR2X1_612/Y D_INPUT_0 0.07fF
C24504 PAND2X1_282/O POR2X1_260/B 0.04fF
C24505 POR2X1_49/Y PAND2X1_201/a_16_344# 0.02fF
C24506 PAND2X1_63/B PAND2X1_529/O 0.03fF
C24507 POR2X1_602/O POR2X1_296/B 0.03fF
C24508 PAND2X1_270/a_76_28# POR2X1_39/B 0.02fF
C24509 POR2X1_9/Y POR2X1_7/B 2.76fF
C24510 PAND2X1_866/O PAND2X1_865/Y 0.00fF
C24511 POR2X1_77/Y POR2X1_503/Y 0.01fF
C24512 PAND2X1_242/Y PAND2X1_6/A 0.10fF
C24513 POR2X1_672/Y POR2X1_14/Y 0.03fF
C24514 POR2X1_848/A POR2X1_669/B 0.10fF
C24515 POR2X1_270/Y POR2X1_269/O 0.18fF
C24516 PAND2X1_830/CTRL POR2X1_416/B 0.01fF
C24517 PAND2X1_606/O POR2X1_102/Y 0.17fF
C24518 PAND2X1_269/a_56_28# INPUT_0 0.00fF
C24519 PAND2X1_221/Y PAND2X1_730/O 0.00fF
C24520 POR2X1_66/B PAND2X1_609/CTRL 0.11fF
C24521 PAND2X1_96/B PAND2X1_125/CTRL 0.06fF
C24522 POR2X1_812/A POR2X1_809/CTRL 0.01fF
C24523 POR2X1_57/A PAND2X1_850/CTRL2 0.03fF
C24524 PAND2X1_666/O PAND2X1_73/Y 0.01fF
C24525 POR2X1_738/A PAND2X1_52/B 0.03fF
C24526 PAND2X1_793/Y POR2X1_250/Y 0.03fF
C24527 POR2X1_725/Y PAND2X1_72/A 0.07fF
C24528 PAND2X1_466/A VDD 0.15fF
C24529 POR2X1_754/Y POR2X1_753/Y 1.27fF
C24530 POR2X1_227/A POR2X1_241/Y 0.37fF
C24531 POR2X1_669/B PAND2X1_711/B 0.03fF
C24532 POR2X1_777/B POR2X1_260/B 0.06fF
C24533 POR2X1_863/A PAND2X1_60/B 0.03fF
C24534 PAND2X1_341/B PAND2X1_476/A 0.02fF
C24535 POR2X1_262/Y VDD 0.14fF
C24536 POR2X1_60/A POR2X1_263/Y 0.03fF
C24537 POR2X1_497/CTRL POR2X1_37/Y 0.03fF
C24538 PAND2X1_93/B POR2X1_808/A 0.02fF
C24539 POR2X1_864/A PAND2X1_760/O 0.00fF
C24540 PAND2X1_73/CTRL POR2X1_66/A 0.03fF
C24541 PAND2X1_214/O PAND2X1_214/A 0.04fF
C24542 PAND2X1_678/O PAND2X1_480/B 0.02fF
C24543 POR2X1_567/B POR2X1_439/O 0.02fF
C24544 POR2X1_48/A PAND2X1_725/Y 0.03fF
C24545 POR2X1_66/B POR2X1_98/O 0.02fF
C24546 POR2X1_48/A PAND2X1_540/CTRL 0.02fF
C24547 POR2X1_260/B PAND2X1_381/CTRL 0.00fF
C24548 POR2X1_78/A POR2X1_267/A 7.01fF
C24549 PAND2X1_65/B POR2X1_260/B 0.26fF
C24550 POR2X1_840/B POR2X1_458/Y 0.05fF
C24551 POR2X1_83/B POR2X1_14/Y 1.10fF
C24552 POR2X1_669/B POR2X1_27/Y 0.17fF
C24553 POR2X1_72/B PAND2X1_777/O 0.01fF
C24554 POR2X1_343/Y PAND2X1_48/A 0.05fF
C24555 POR2X1_559/A PAND2X1_72/A 0.15fF
C24556 PAND2X1_436/CTRL2 INPUT_0 0.10fF
C24557 POR2X1_220/B PAND2X1_41/B 0.03fF
C24558 POR2X1_541/B POR2X1_579/Y 0.03fF
C24559 PAND2X1_412/a_76_28# POR2X1_260/B 0.02fF
C24560 POR2X1_129/a_56_344# PAND2X1_390/Y 0.01fF
C24561 PAND2X1_23/Y POR2X1_444/CTRL2 0.01fF
C24562 PAND2X1_222/a_16_344# INPUT_0 0.01fF
C24563 POR2X1_65/A D_INPUT_0 0.04fF
C24564 POR2X1_52/A POR2X1_628/Y 0.03fF
C24565 POR2X1_863/A POR2X1_353/A 0.03fF
C24566 POR2X1_84/A VDD 0.20fF
C24567 POR2X1_462/CTRL PAND2X1_69/A 0.03fF
C24568 POR2X1_326/a_16_28# POR2X1_568/A 0.03fF
C24569 POR2X1_220/B POR2X1_781/A 0.03fF
C24570 D_INPUT_0 POR2X1_362/B 0.03fF
C24571 POR2X1_433/CTRL POR2X1_72/B 0.01fF
C24572 POR2X1_476/Y POR2X1_66/A 0.46fF
C24573 POR2X1_278/Y PAND2X1_205/O 0.08fF
C24574 PAND2X1_860/A PAND2X1_861/O 0.07fF
C24575 POR2X1_657/Y POR2X1_222/Y 0.01fF
C24576 POR2X1_416/B POR2X1_4/Y 0.07fF
C24577 POR2X1_179/CTRL POR2X1_411/B 0.01fF
C24578 POR2X1_620/CTRL2 PAND2X1_9/Y 0.01fF
C24579 PAND2X1_214/CTRL VDD 0.00fF
C24580 POR2X1_169/A POR2X1_568/B 0.03fF
C24581 PAND2X1_220/Y POR2X1_102/Y 0.03fF
C24582 POR2X1_20/Y PAND2X1_33/a_16_344# 0.04fF
C24583 POR2X1_66/B POR2X1_404/CTRL 0.01fF
C24584 PAND2X1_48/B POR2X1_445/A 0.00fF
C24585 POR2X1_514/Y PAND2X1_39/B 0.03fF
C24586 POR2X1_48/A POR2X1_88/Y 0.03fF
C24587 POR2X1_566/A POR2X1_270/Y 0.03fF
C24588 POR2X1_496/Y POR2X1_627/a_56_344# 0.01fF
C24589 POR2X1_614/A POR2X1_541/B 0.08fF
C24590 POR2X1_52/A PAND2X1_267/Y 0.02fF
C24591 POR2X1_68/A POR2X1_341/A 0.10fF
C24592 PAND2X1_266/CTRL POR2X1_7/A 0.01fF
C24593 POR2X1_29/Y POR2X1_411/B 0.03fF
C24594 POR2X1_624/Y POR2X1_565/CTRL 0.01fF
C24595 PAND2X1_798/B POR2X1_679/A 0.03fF
C24596 POR2X1_60/A POR2X1_251/m4_208_n4# 0.12fF
C24597 POR2X1_866/A POR2X1_294/B 0.03fF
C24598 PAND2X1_863/a_56_28# POR2X1_102/Y 0.00fF
C24599 POR2X1_830/CTRL2 POR2X1_830/A 0.01fF
C24600 POR2X1_67/Y POR2X1_748/Y 0.00fF
C24601 POR2X1_516/O POR2X1_257/A 0.01fF
C24602 POR2X1_83/B POR2X1_237/CTRL 0.01fF
C24603 PAND2X1_43/CTRL PAND2X1_69/A 0.01fF
C24604 POR2X1_158/a_16_28# POR2X1_416/B 0.01fF
C24605 POR2X1_83/B POR2X1_48/O 0.10fF
C24606 POR2X1_694/O POR2X1_257/A 0.18fF
C24607 POR2X1_195/A POR2X1_294/B 0.03fF
C24608 POR2X1_48/A POR2X1_232/O 0.01fF
C24609 POR2X1_130/A POR2X1_288/O 0.10fF
C24610 POR2X1_360/A POR2X1_66/A 0.03fF
C24611 POR2X1_362/Y VDD 0.00fF
C24612 PAND2X1_6/Y POR2X1_688/Y 0.04fF
C24613 POR2X1_683/CTRL2 POR2X1_669/B 0.01fF
C24614 POR2X1_285/Y VDD -0.00fF
C24615 POR2X1_199/CTRL2 POR2X1_590/A 0.00fF
C24616 POR2X1_150/Y POR2X1_387/Y 0.07fF
C24617 PAND2X1_213/CTRL PAND2X1_161/Y 0.01fF
C24618 POR2X1_334/B POR2X1_476/A 0.02fF
C24619 POR2X1_366/Y POR2X1_269/CTRL2 0.01fF
C24620 PAND2X1_430/O POR2X1_750/B 0.07fF
C24621 PAND2X1_650/O PAND2X1_9/Y 0.02fF
C24622 POR2X1_413/A PAND2X1_656/CTRL2 0.01fF
C24623 PAND2X1_472/B POR2X1_83/B 0.98fF
C24624 PAND2X1_240/O POR2X1_5/Y 0.03fF
C24625 PAND2X1_282/O PAND2X1_55/Y 0.07fF
C24626 PAND2X1_661/Y POR2X1_20/B 0.03fF
C24627 PAND2X1_84/Y PAND2X1_558/Y 0.01fF
C24628 POR2X1_691/CTRL POR2X1_811/A 0.00fF
C24629 POR2X1_276/A POR2X1_276/B 0.08fF
C24630 PAND2X1_630/CTRL2 POR2X1_496/Y 0.06fF
C24631 POR2X1_78/A POR2X1_149/Y 0.04fF
C24632 PAND2X1_46/O INPUT_0 0.01fF
C24633 PAND2X1_742/B POR2X1_32/A 0.03fF
C24634 POR2X1_454/A POR2X1_532/A 0.02fF
C24635 PAND2X1_440/m4_208_n4# PAND2X1_804/m4_208_n4# 0.05fF
C24636 PAND2X1_309/O PAND2X1_58/A 0.02fF
C24637 POR2X1_634/A POR2X1_638/CTRL2 0.17fF
C24638 PAND2X1_658/A POR2X1_67/A 0.02fF
C24639 PAND2X1_839/CTRL2 POR2X1_102/Y 0.01fF
C24640 POR2X1_60/A PAND2X1_215/B 0.03fF
C24641 POR2X1_83/B POR2X1_55/Y 2.08fF
C24642 POR2X1_129/CTRL2 POR2X1_90/Y 0.01fF
C24643 POR2X1_96/A PAND2X1_76/a_76_28# 0.01fF
C24644 PAND2X1_20/A PAND2X1_496/O 0.03fF
C24645 POR2X1_556/A POR2X1_456/B 0.03fF
C24646 POR2X1_257/A PAND2X1_467/CTRL2 0.00fF
C24647 POR2X1_66/B POR2X1_193/A 0.03fF
C24648 PAND2X1_296/a_16_344# POR2X1_42/Y 0.02fF
C24649 POR2X1_66/B POR2X1_579/Y 0.03fF
C24650 POR2X1_523/Y POR2X1_819/CTRL2 0.01fF
C24651 PAND2X1_48/B POR2X1_792/a_16_28# 0.01fF
C24652 PAND2X1_307/a_76_28# POR2X1_304/Y 0.07fF
C24653 POR2X1_300/m4_208_n4# D_INPUT_0 0.09fF
C24654 POR2X1_41/B PAND2X1_731/B 0.04fF
C24655 POR2X1_274/A PAND2X1_60/B 0.03fF
C24656 PAND2X1_65/Y VDD 0.18fF
C24657 PAND2X1_169/Y PAND2X1_714/CTRL 0.01fF
C24658 POR2X1_66/B POR2X1_445/m4_208_n4# 0.15fF
C24659 POR2X1_264/Y PAND2X1_265/CTRL 0.01fF
C24660 POR2X1_779/A PAND2X1_73/Y 0.01fF
C24661 POR2X1_427/O PAND2X1_565/A 0.00fF
C24662 PAND2X1_58/A POR2X1_460/B 0.02fF
C24663 PAND2X1_362/A PAND2X1_794/B 0.00fF
C24664 PAND2X1_82/O POR2X1_84/A 0.03fF
C24665 POR2X1_115/a_76_344# POR2X1_330/Y 0.04fF
C24666 POR2X1_514/Y PAND2X1_20/A 0.01fF
C24667 PAND2X1_833/a_56_28# POR2X1_376/B 0.00fF
C24668 POR2X1_415/A POR2X1_750/Y -0.00fF
C24669 POR2X1_626/Y POR2X1_55/Y 0.00fF
C24670 POR2X1_52/A PAND2X1_808/B 0.01fF
C24671 PAND2X1_657/CTRL2 POR2X1_816/A 0.03fF
C24672 POR2X1_683/Y POR2X1_603/Y 0.01fF
C24673 POR2X1_807/A POR2X1_722/Y 0.04fF
C24674 PAND2X1_54/CTRL VDD -0.00fF
C24675 D_INPUT_0 POR2X1_550/O 0.01fF
C24676 POR2X1_786/A PAND2X1_41/B 0.42fF
C24677 PAND2X1_454/a_76_28# POR2X1_60/A 0.02fF
C24678 POR2X1_65/A PAND2X1_364/CTRL2 0.03fF
C24679 PAND2X1_58/A POR2X1_790/A 6.75fF
C24680 POR2X1_66/B POR2X1_43/B 0.01fF
C24681 PAND2X1_206/A PAND2X1_100/O 0.05fF
C24682 POR2X1_60/A PAND2X1_6/A 0.24fF
C24683 POR2X1_777/B PAND2X1_55/Y 0.10fF
C24684 PAND2X1_787/Y PAND2X1_804/B 0.10fF
C24685 POR2X1_477/Y POR2X1_478/B 0.04fF
C24686 POR2X1_752/Y POR2X1_55/Y 0.03fF
C24687 POR2X1_66/B POR2X1_789/A 0.03fF
C24688 POR2X1_555/A POR2X1_555/a_16_28# 0.05fF
C24689 POR2X1_376/B POR2X1_372/Y 0.76fF
C24690 POR2X1_66/A PAND2X1_305/CTRL 0.01fF
C24691 PAND2X1_246/CTRL2 POR2X1_4/Y 0.01fF
C24692 PAND2X1_96/B PAND2X1_39/O 0.11fF
C24693 PAND2X1_863/B POR2X1_236/Y 0.03fF
C24694 PAND2X1_480/B PAND2X1_84/Y 0.03fF
C24695 POR2X1_660/A PAND2X1_55/Y 0.02fF
C24696 POR2X1_66/B POR2X1_614/A 0.04fF
C24697 POR2X1_623/A POR2X1_623/CTRL2 0.01fF
C24698 POR2X1_567/B PAND2X1_315/O 0.30fF
C24699 POR2X1_198/B POR2X1_61/Y 0.05fF
C24700 POR2X1_508/O POR2X1_852/B 0.07fF
C24701 PAND2X1_808/Y PAND2X1_220/Y 0.03fF
C24702 POR2X1_96/A PAND2X1_362/B 0.03fF
C24703 POR2X1_102/Y PAND2X1_575/CTRL 0.00fF
C24704 PAND2X1_65/B POR2X1_205/Y 0.00fF
C24705 PAND2X1_208/O POR2X1_599/A 0.25fF
C24706 POR2X1_486/B POR2X1_486/CTRL 0.02fF
C24707 PAND2X1_95/B PAND2X1_588/O 0.03fF
C24708 PAND2X1_65/B PAND2X1_55/Y 0.25fF
C24709 POR2X1_207/A POR2X1_294/B 0.01fF
C24710 POR2X1_188/A POR2X1_614/A 0.03fF
C24711 POR2X1_418/Y POR2X1_73/Y 0.01fF
C24712 POR2X1_66/B POR2X1_38/B 0.03fF
C24713 POR2X1_40/Y POR2X1_90/Y 0.15fF
C24714 POR2X1_824/Y POR2X1_102/Y 0.12fF
C24715 POR2X1_602/A PAND2X1_60/B 0.01fF
C24716 POR2X1_13/A POR2X1_46/Y 0.14fF
C24717 POR2X1_443/a_56_344# POR2X1_192/B 0.00fF
C24718 POR2X1_661/B VDD 0.00fF
C24719 PAND2X1_65/B POR2X1_205/O 0.18fF
C24720 POR2X1_278/Y POR2X1_7/B 0.03fF
C24721 POR2X1_624/Y PAND2X1_48/A 0.02fF
C24722 PAND2X1_96/B POR2X1_259/A 0.09fF
C24723 PAND2X1_73/Y POR2X1_598/CTRL2 0.01fF
C24724 POR2X1_416/B POR2X1_827/a_76_344# 0.01fF
C24725 POR2X1_8/Y POR2X1_48/A 18.39fF
C24726 POR2X1_68/A PAND2X1_58/CTRL2 0.01fF
C24727 POR2X1_61/O POR2X1_66/A 0.01fF
C24728 POR2X1_376/B POR2X1_253/Y 0.01fF
C24729 PAND2X1_287/O VDD 0.00fF
C24730 POR2X1_153/CTRL2 POR2X1_37/Y 0.01fF
C24731 POR2X1_380/CTRL POR2X1_5/Y 0.00fF
C24732 PAND2X1_48/B PAND2X1_48/O 0.05fF
C24733 POR2X1_706/CTRL2 PAND2X1_94/A 0.03fF
C24734 PAND2X1_241/Y POR2X1_417/Y 0.54fF
C24735 POR2X1_29/Y POR2X1_376/B 0.03fF
C24736 POR2X1_302/CTRL2 PAND2X1_6/Y 0.03fF
C24737 POR2X1_23/Y POR2X1_394/A 3.01fF
C24738 PAND2X1_41/B POR2X1_758/O 0.04fF
C24739 POR2X1_664/CTRL2 PAND2X1_73/Y 0.03fF
C24740 POR2X1_45/Y PAND2X1_473/Y 0.03fF
C24741 PAND2X1_494/CTRL2 INPUT_0 0.06fF
C24742 POR2X1_753/Y POR2X1_754/CTRL 0.02fF
C24743 POR2X1_754/Y POR2X1_754/O 0.01fF
C24744 POR2X1_566/A POR2X1_562/O 0.30fF
C24745 POR2X1_43/B PAND2X1_556/B 0.05fF
C24746 POR2X1_355/B POR2X1_477/A 0.03fF
C24747 PAND2X1_470/O PAND2X1_803/A 0.00fF
C24748 PAND2X1_48/B PAND2X1_152/CTRL 0.01fF
C24749 PAND2X1_20/A POR2X1_576/CTRL2 0.01fF
C24750 POR2X1_785/A POR2X1_776/B 0.03fF
C24751 POR2X1_614/A PAND2X1_129/a_16_344# 0.02fF
C24752 PAND2X1_65/B POR2X1_407/Y 0.04fF
C24753 POR2X1_855/B POR2X1_783/O 0.01fF
C24754 PAND2X1_213/Y PAND2X1_714/A 0.07fF
C24755 PAND2X1_578/A VDD 0.00fF
C24756 POR2X1_256/CTRL POR2X1_255/Y 0.01fF
C24757 POR2X1_859/A POR2X1_789/A 0.07fF
C24758 POR2X1_97/O PAND2X1_20/A 0.18fF
C24759 POR2X1_78/B POR2X1_335/Y 0.01fF
C24760 POR2X1_376/B POR2X1_9/O 0.02fF
C24761 POR2X1_154/O POR2X1_68/A 0.02fF
C24762 POR2X1_50/a_56_344# INPUT_6 0.00fF
C24763 PAND2X1_80/CTRL POR2X1_68/B 0.01fF
C24764 POR2X1_57/A PAND2X1_473/B 0.03fF
C24765 PAND2X1_129/a_16_344# POR2X1_38/B 0.01fF
C24766 POR2X1_52/A POR2X1_22/A 0.02fF
C24767 PAND2X1_6/Y POR2X1_502/A 0.06fF
C24768 POR2X1_400/A POR2X1_206/CTRL2 0.11fF
C24769 POR2X1_407/A POR2X1_722/Y 0.15fF
C24770 POR2X1_812/A POR2X1_260/A 0.01fF
C24771 POR2X1_614/A POR2X1_155/Y 0.01fF
C24772 POR2X1_351/B POR2X1_97/A 0.01fF
C24773 POR2X1_57/A POR2X1_397/Y 0.01fF
C24774 POR2X1_52/A POR2X1_519/Y 0.02fF
C24775 PAND2X1_182/A PAND2X1_357/Y 0.01fF
C24776 PAND2X1_6/Y POR2X1_783/A 0.00fF
C24777 PAND2X1_455/Y POR2X1_73/Y 0.00fF
C24778 POR2X1_78/A POR2X1_558/Y 0.03fF
C24779 PAND2X1_115/Y POR2X1_183/Y 0.00fF
C24780 POR2X1_684/a_16_28# POR2X1_42/Y 0.02fF
C24781 PAND2X1_239/O POR2X1_191/Y 0.05fF
C24782 PAND2X1_239/a_16_344# POR2X1_192/B 0.03fF
C24783 POR2X1_859/A POR2X1_38/B 0.07fF
C24784 PAND2X1_6/Y POR2X1_247/CTRL 0.01fF
C24785 POR2X1_16/A POR2X1_72/B 1.53fF
C24786 PAND2X1_371/CTRL2 PAND2X1_32/B 0.03fF
C24787 PAND2X1_389/Y VDD 0.18fF
C24788 PAND2X1_732/A POR2X1_40/Y 0.09fF
C24789 PAND2X1_197/CTRL2 POR2X1_52/Y 0.00fF
C24790 PAND2X1_661/B POR2X1_46/Y 0.69fF
C24791 POR2X1_198/B POR2X1_35/Y 0.03fF
C24792 POR2X1_718/CTRL2 POR2X1_834/Y 0.15fF
C24793 POR2X1_578/Y POR2X1_775/O 0.01fF
C24794 PAND2X1_6/Y POR2X1_464/Y 0.01fF
C24795 INPUT_0 POR2X1_318/A 0.07fF
C24796 POR2X1_28/a_76_344# POR2X1_4/Y 0.02fF
C24797 PAND2X1_662/CTRL2 POR2X1_413/A 0.01fF
C24798 POR2X1_403/B PAND2X1_60/B 0.03fF
C24799 POR2X1_81/CTRL PAND2X1_573/B 0.01fF
C24800 POR2X1_21/CTRL2 INPUT_4 0.05fF
C24801 POR2X1_106/Y PAND2X1_114/B 0.01fF
C24802 PAND2X1_94/A POR2X1_287/B 0.05fF
C24803 PAND2X1_213/B PAND2X1_161/Y 0.04fF
C24804 PAND2X1_844/CTRL2 POR2X1_60/Y 0.01fF
C24805 POR2X1_52/A POR2X1_239/O 0.01fF
C24806 POR2X1_327/Y POR2X1_830/O 0.33fF
C24807 POR2X1_48/A PAND2X1_346/CTRL 0.00fF
C24808 POR2X1_733/A POR2X1_513/Y 0.07fF
C24809 PAND2X1_632/B POR2X1_5/Y 0.03fF
C24810 POR2X1_315/Y POR2X1_236/Y 0.45fF
C24811 POR2X1_761/Y POR2X1_7/B 0.03fF
C24812 POR2X1_78/B PAND2X1_315/O 0.07fF
C24813 POR2X1_83/B PAND2X1_199/B 0.03fF
C24814 PAND2X1_865/Y POR2X1_487/O 0.00fF
C24815 POR2X1_748/A PAND2X1_156/B 1.11fF
C24816 PAND2X1_69/A POR2X1_740/Y 0.07fF
C24817 PAND2X1_212/O POR2X1_77/Y 0.08fF
C24818 POR2X1_312/Y POR2X1_394/A 0.03fF
C24819 POR2X1_640/Y POR2X1_557/B 0.03fF
C24820 POR2X1_390/B POR2X1_78/B 0.03fF
C24821 POR2X1_688/Y PAND2X1_52/B 0.02fF
C24822 POR2X1_130/A POR2X1_101/Y 0.19fF
C24823 POR2X1_119/Y POR2X1_60/A 0.55fF
C24824 PAND2X1_823/CTRL VDD -0.00fF
C24825 POR2X1_651/O PAND2X1_60/B 0.00fF
C24826 PAND2X1_94/A PAND2X1_8/Y 0.16fF
C24827 POR2X1_9/Y PAND2X1_206/B 0.14fF
C24828 POR2X1_16/A PAND2X1_520/CTRL2 0.00fF
C24829 POR2X1_644/A POR2X1_796/CTRL2 0.02fF
C24830 PAND2X1_29/CTRL2 POR2X1_68/B 0.04fF
C24831 POR2X1_158/O POR2X1_669/B 0.06fF
C24832 PAND2X1_651/Y POR2X1_52/Y 0.05fF
C24833 POR2X1_333/Y PAND2X1_65/B 0.02fF
C24834 PAND2X1_672/O POR2X1_35/B 0.04fF
C24835 POR2X1_502/A PAND2X1_698/CTRL2 0.02fF
C24836 POR2X1_532/A POR2X1_713/O 0.34fF
C24837 PAND2X1_642/B POR2X1_73/Y 0.02fF
C24838 INPUT_0 PAND2X1_537/O 0.02fF
C24839 PAND2X1_702/a_76_28# POR2X1_42/Y 0.00fF
C24840 POR2X1_96/A POR2X1_419/CTRL 0.02fF
C24841 POR2X1_346/B POR2X1_404/B 0.07fF
C24842 POR2X1_42/Y PAND2X1_656/A 0.03fF
C24843 POR2X1_394/A PAND2X1_558/O 0.07fF
C24844 POR2X1_514/CTRL POR2X1_137/Y 0.01fF
C24845 POR2X1_693/a_76_344# PAND2X1_550/B 0.00fF
C24846 POR2X1_303/O POR2X1_330/Y 0.04fF
C24847 PAND2X1_48/B PAND2X1_747/a_76_28# 0.01fF
C24848 PAND2X1_490/CTRL POR2X1_38/B 0.00fF
C24849 PAND2X1_111/B PAND2X1_111/CTRL 0.01fF
C24850 PAND2X1_366/A POR2X1_42/Y 0.03fF
C24851 POR2X1_69/Y POR2X1_67/Y 0.10fF
C24852 POR2X1_445/CTRL POR2X1_456/B 0.01fF
C24853 PAND2X1_242/a_16_344# PAND2X1_241/Y 0.03fF
C24854 PAND2X1_653/CTRL POR2X1_83/B 0.01fF
C24855 POR2X1_541/O POR2X1_702/A 0.00fF
C24856 PAND2X1_803/Y POR2X1_183/Y 0.03fF
C24857 PAND2X1_615/O D_INPUT_1 0.06fF
C24858 POR2X1_16/A PAND2X1_216/CTRL -0.01fF
C24859 PAND2X1_696/CTRL POR2X1_602/B 0.01fF
C24860 PAND2X1_96/B PAND2X1_88/Y 0.03fF
C24861 POR2X1_865/B PAND2X1_96/B 0.02fF
C24862 PAND2X1_651/Y PAND2X1_241/Y 0.00fF
C24863 POR2X1_383/A POR2X1_341/O 0.03fF
C24864 INPUT_1 POR2X1_615/Y 0.00fF
C24865 POR2X1_65/A PAND2X1_643/A 0.02fF
C24866 POR2X1_366/Y POR2X1_703/A 0.08fF
C24867 POR2X1_283/A PAND2X1_357/Y 0.23fF
C24868 POR2X1_646/B POR2X1_646/A 0.06fF
C24869 POR2X1_364/A POR2X1_319/Y 4.31fF
C24870 PAND2X1_209/A PAND2X1_797/CTRL 0.01fF
C24871 PAND2X1_48/B POR2X1_260/A 4.12fF
C24872 POR2X1_9/Y POR2X1_818/CTRL 0.08fF
C24873 POR2X1_556/Y POR2X1_510/Y 0.01fF
C24874 POR2X1_516/A PAND2X1_6/A 0.01fF
C24875 PAND2X1_638/O POR2X1_588/Y 0.08fF
C24876 POR2X1_635/B PAND2X1_762/O 0.01fF
C24877 POR2X1_416/B PAND2X1_219/A 0.03fF
C24878 POR2X1_65/Y POR2X1_9/Y 0.02fF
C24879 POR2X1_740/Y PAND2X1_368/a_76_28# 0.03fF
C24880 POR2X1_741/Y PAND2X1_368/a_16_344# 0.02fF
C24881 POR2X1_185/CTRL PAND2X1_94/A 0.06fF
C24882 PAND2X1_422/CTRL POR2X1_788/B 0.01fF
C24883 POR2X1_52/A PAND2X1_620/a_16_344# 0.01fF
C24884 POR2X1_38/Y POR2X1_235/CTRL2 0.03fF
C24885 PAND2X1_723/a_16_344# PAND2X1_656/A 0.01fF
C24886 POR2X1_62/Y POR2X1_88/Y 0.05fF
C24887 PAND2X1_593/O POR2X1_385/Y 0.04fF
C24888 POR2X1_13/A POR2X1_371/CTRL 0.01fF
C24889 PAND2X1_348/A POR2X1_42/Y 0.07fF
C24890 PAND2X1_824/B POR2X1_740/Y 0.10fF
C24891 PAND2X1_854/a_76_28# PAND2X1_856/B 0.04fF
C24892 D_GATE_662 POR2X1_444/Y 0.04fF
C24893 PAND2X1_48/B POR2X1_363/A 0.46fF
C24894 POR2X1_811/B PAND2X1_72/A 0.03fF
C24895 PAND2X1_784/CTRL2 PAND2X1_156/A 0.28fF
C24896 PAND2X1_550/B POR2X1_73/Y 0.06fF
C24897 PAND2X1_731/B POR2X1_77/Y 0.02fF
C24898 POR2X1_760/Y PAND2X1_687/Y 0.17fF
C24899 POR2X1_49/Y PAND2X1_198/O 0.02fF
C24900 POR2X1_614/A PAND2X1_313/CTRL 0.08fF
C24901 POR2X1_416/B PAND2X1_221/a_76_28# 0.02fF
C24902 PAND2X1_841/O POR2X1_153/Y 0.17fF
C24903 PAND2X1_254/CTRL2 PAND2X1_508/Y 0.00fF
C24904 PAND2X1_57/B PAND2X1_328/O 0.17fF
C24905 POR2X1_88/O POR2X1_9/Y 0.02fF
C24906 POR2X1_293/Y POR2X1_371/CTRL2 0.01fF
C24907 PAND2X1_473/B POR2X1_589/CTRL 0.01fF
C24908 POR2X1_862/O POR2X1_389/Y 0.09fF
C24909 POR2X1_25/CTRL2 D_INPUT_4 0.01fF
C24910 POR2X1_101/Y PAND2X1_150/O 0.10fF
C24911 POR2X1_68/A PAND2X1_142/CTRL 0.04fF
C24912 PAND2X1_551/Y POR2X1_394/A 0.01fF
C24913 POR2X1_43/B PAND2X1_358/A 0.15fF
C24914 POR2X1_775/A POR2X1_332/a_16_28# 0.02fF
C24915 POR2X1_785/A POR2X1_192/B 0.03fF
C24916 PAND2X1_552/B PAND2X1_703/O 0.17fF
C24917 PAND2X1_106/O POR2X1_383/A 0.01fF
C24918 POR2X1_22/A POR2X1_3/B 0.73fF
C24919 PAND2X1_717/Y POR2X1_7/A 0.03fF
C24920 POR2X1_118/CTRL PAND2X1_560/B 0.03fF
C24921 POR2X1_38/B POR2X1_6/CTRL 0.06fF
C24922 POR2X1_544/m4_208_n4# POR2X1_854/B 0.08fF
C24923 PAND2X1_202/a_16_344# POR2X1_66/A 0.02fF
C24924 POR2X1_416/B PAND2X1_193/CTRL 0.08fF
C24925 POR2X1_814/A POR2X1_260/B 0.16fF
C24926 PAND2X1_75/CTRL POR2X1_260/B 0.01fF
C24927 POR2X1_567/A PAND2X1_280/a_76_28# -0.00fF
C24928 POR2X1_523/Y POR2X1_550/B 0.01fF
C24929 POR2X1_45/Y POR2X1_7/Y 0.03fF
C24930 PAND2X1_631/A POR2X1_42/Y 0.23fF
C24931 POR2X1_16/A PAND2X1_570/B 0.01fF
C24932 POR2X1_327/Y POR2X1_788/B 0.03fF
C24933 POR2X1_294/B POR2X1_342/a_16_28# 0.02fF
C24934 POR2X1_99/B POR2X1_222/Y 0.03fF
C24935 POR2X1_863/A POR2X1_750/B 0.06fF
C24936 POR2X1_383/A POR2X1_734/CTRL2 0.02fF
C24937 POR2X1_537/O POR2X1_537/B 0.02fF
C24938 POR2X1_846/Y POR2X1_260/B 0.03fF
C24939 POR2X1_669/B POR2X1_827/CTRL 0.01fF
C24940 PAND2X1_6/Y POR2X1_188/Y 0.03fF
C24941 POR2X1_456/B POR2X1_180/A 0.03fF
C24942 POR2X1_49/Y POR2X1_90/a_76_344# 0.01fF
C24943 POR2X1_265/Y PAND2X1_734/O 0.02fF
C24944 PAND2X1_152/CTRL2 POR2X1_711/Y 0.05fF
C24945 POR2X1_57/A POR2X1_131/A 0.12fF
C24946 PAND2X1_675/CTRL PAND2X1_736/A 0.02fF
C24947 PAND2X1_335/CTRL POR2X1_77/Y 0.01fF
C24948 PAND2X1_849/B PAND2X1_100/a_16_344# 0.01fF
C24949 POR2X1_493/CTRL PAND2X1_48/A 0.00fF
C24950 POR2X1_502/A PAND2X1_52/B 0.24fF
C24951 POR2X1_43/CTRL POR2X1_42/Y 0.01fF
C24952 POR2X1_540/A POR2X1_552/a_16_28# 0.02fF
C24953 PAND2X1_286/CTRL2 GATE_222 0.01fF
C24954 POR2X1_783/A PAND2X1_52/B 0.00fF
C24955 POR2X1_1/m4_208_n4# POR2X1_260/A 0.09fF
C24956 POR2X1_99/B POR2X1_532/A 0.03fF
C24957 POR2X1_9/Y POR2X1_750/B 0.07fF
C24958 POR2X1_782/A POR2X1_568/B 0.05fF
C24959 POR2X1_845/A POR2X1_845/CTRL2 0.04fF
C24960 POR2X1_494/Y POR2X1_80/CTRL 0.00fF
C24961 POR2X1_647/B POR2X1_655/A 0.01fF
C24962 POR2X1_57/A POR2X1_518/CTRL 0.01fF
C24963 POR2X1_67/Y PAND2X1_225/CTRL 0.00fF
C24964 POR2X1_711/B POR2X1_710/B -0.02fF
C24965 POR2X1_120/O POR2X1_651/Y 0.07fF
C24966 PAND2X1_96/B POR2X1_568/B 0.03fF
C24967 PAND2X1_196/CTRL PAND2X1_199/B 0.00fF
C24968 PAND2X1_440/O POR2X1_437/Y -0.00fF
C24969 POR2X1_554/a_16_28# POR2X1_112/Y 0.01fF
C24970 POR2X1_432/O POR2X1_271/B 0.01fF
C24971 POR2X1_345/A POR2X1_814/A 0.04fF
C24972 POR2X1_390/B POR2X1_294/A 0.03fF
C24973 POR2X1_68/A PAND2X1_681/CTRL 0.03fF
C24974 POR2X1_407/A PAND2X1_681/CTRL2 0.01fF
C24975 PAND2X1_55/Y PAND2X1_178/CTRL2 0.13fF
C24976 POR2X1_588/a_16_28# POR2X1_587/Y 0.10fF
C24977 PAND2X1_826/CTRL POR2X1_294/Y 0.02fF
C24978 POR2X1_8/Y POR2X1_62/Y 1.20fF
C24979 POR2X1_815/O POR2X1_750/A 0.02fF
C24980 POR2X1_539/CTRL POR2X1_567/A 0.01fF
C24981 PAND2X1_479/O POR2X1_329/A 0.03fF
C24982 POR2X1_147/a_16_28# POR2X1_147/A 0.03fF
C24983 POR2X1_119/Y PAND2X1_301/CTRL 0.01fF
C24984 POR2X1_864/A POR2X1_780/CTRL2 0.01fF
C24985 POR2X1_760/Y PAND2X1_691/Y 0.00fF
C24986 POR2X1_505/a_16_28# PAND2X1_156/A 0.04fF
C24987 POR2X1_804/A POR2X1_717/B 0.05fF
C24988 PAND2X1_48/A POR2X1_186/B 0.06fF
C24989 POR2X1_262/Y PAND2X1_786/a_16_344# 0.02fF
C24990 PAND2X1_213/Y PAND2X1_169/a_76_28# 0.01fF
C24991 PAND2X1_425/Y PAND2X1_582/O 0.02fF
C24992 PAND2X1_109/O POR2X1_854/B 0.04fF
C24993 POR2X1_228/Y POR2X1_716/O 0.02fF
C24994 PAND2X1_831/CTRL2 POR2X1_411/B 0.01fF
C24995 POR2X1_9/Y POR2X1_618/CTRL 0.15fF
C24996 POR2X1_647/O POR2X1_296/B 0.02fF
C24997 POR2X1_416/B PAND2X1_854/A 0.11fF
C24998 POR2X1_540/A POR2X1_181/A 0.12fF
C24999 POR2X1_485/Y POR2X1_376/B 0.03fF
C25000 POR2X1_23/Y POR2X1_669/B 1.93fF
C25001 POR2X1_344/Y POR2X1_359/a_16_28# 0.00fF
C25002 POR2X1_760/A PAND2X1_362/B 0.01fF
C25003 POR2X1_379/CTRL PAND2X1_52/B 0.13fF
C25004 PAND2X1_793/Y POR2X1_329/A 0.03fF
C25005 PAND2X1_86/O PAND2X1_57/B 0.05fF
C25006 PAND2X1_96/O PAND2X1_60/B 0.03fF
C25007 POR2X1_814/B POR2X1_471/A 0.01fF
C25008 POR2X1_76/A POR2X1_141/Y 0.03fF
C25009 POR2X1_260/B POR2X1_405/CTRL2 0.01fF
C25010 PAND2X1_841/B POR2X1_329/A 0.03fF
C25011 PAND2X1_771/Y PAND2X1_564/B 0.36fF
C25012 POR2X1_79/a_56_344# PAND2X1_354/A 0.00fF
C25013 POR2X1_16/A PAND2X1_440/O 0.26fF
C25014 POR2X1_814/A POR2X1_205/Y 0.07fF
C25015 POR2X1_442/CTRL2 POR2X1_236/Y 0.01fF
C25016 POR2X1_814/A PAND2X1_55/Y 0.20fF
C25017 POR2X1_753/Y POR2X1_67/A 0.04fF
C25018 PAND2X1_404/Y PAND2X1_500/a_16_344# 0.01fF
C25019 PAND2X1_23/Y POR2X1_284/a_16_28# 0.02fF
C25020 POR2X1_252/Y PAND2X1_631/A 0.04fF
C25021 POR2X1_681/Y POR2X1_682/O 0.01fF
C25022 PAND2X1_98/O VDD 0.00fF
C25023 POR2X1_556/A PAND2X1_57/B 0.13fF
C25024 POR2X1_866/A POR2X1_807/A 0.03fF
C25025 POR2X1_115/O POR2X1_116/A 0.01fF
C25026 POR2X1_12/A POR2X1_2/CTRL 0.01fF
C25027 POR2X1_265/a_16_28# POR2X1_40/Y 0.02fF
C25028 POR2X1_52/CTRL POR2X1_7/Y 0.01fF
C25029 PAND2X1_844/CTRL2 PAND2X1_351/A 0.00fF
C25030 POR2X1_554/B POR2X1_276/CTRL 0.01fF
C25031 POR2X1_48/A PAND2X1_62/CTRL2 0.02fF
C25032 PAND2X1_571/A PAND2X1_576/O 0.03fF
C25033 PAND2X1_603/CTRL2 POR2X1_750/B 0.10fF
C25034 POR2X1_417/Y PAND2X1_220/A 0.03fF
C25035 POR2X1_830/CTRL POR2X1_590/A 0.01fF
C25036 POR2X1_66/B POR2X1_590/A 0.13fF
C25037 POR2X1_490/CTRL2 PAND2X1_215/B 0.00fF
C25038 PAND2X1_58/A PAND2X1_585/CTRL2 0.00fF
C25039 INPUT_2 PAND2X1_608/CTRL2 0.01fF
C25040 POR2X1_43/B PAND2X1_447/CTRL2 0.03fF
C25041 PAND2X1_307/CTRL2 POR2X1_14/Y 0.00fF
C25042 POR2X1_27/CTRL2 POR2X1_38/Y 0.03fF
C25043 POR2X1_446/B POR2X1_724/O 0.01fF
C25044 POR2X1_754/Y POR2X1_615/CTRL 0.00fF
C25045 POR2X1_753/Y POR2X1_615/CTRL2 0.07fF
C25046 POR2X1_450/B PAND2X1_427/CTRL2 0.01fF
C25047 PAND2X1_307/CTRL2 PAND2X1_453/A 0.01fF
C25048 POR2X1_814/A POR2X1_407/Y 0.05fF
C25049 POR2X1_188/A POR2X1_590/A 0.06fF
C25050 POR2X1_253/O POR2X1_293/Y 0.07fF
C25051 PAND2X1_48/B POR2X1_610/Y 0.21fF
C25052 PAND2X1_792/O PAND2X1_805/A 0.02fF
C25053 PAND2X1_423/CTRL POR2X1_78/A 0.01fF
C25054 POR2X1_671/CTRL POR2X1_37/Y 0.04fF
C25055 POR2X1_654/B POR2X1_121/B 0.01fF
C25056 PAND2X1_225/CTRL2 POR2X1_750/B 0.01fF
C25057 PAND2X1_793/Y POR2X1_67/O 0.01fF
C25058 PAND2X1_52/B POR2X1_188/Y 0.01fF
C25059 POR2X1_55/O POR2X1_5/Y 0.01fF
C25060 POR2X1_260/B INPUT_5 0.02fF
C25061 POR2X1_296/CTRL2 POR2X1_68/B 0.01fF
C25062 POR2X1_48/A POR2X1_516/B 0.00fF
C25063 PAND2X1_58/A PAND2X1_395/CTRL 0.01fF
C25064 POR2X1_45/Y POR2X1_257/A 1.81fF
C25065 POR2X1_20/B PAND2X1_546/O 0.02fF
C25066 PAND2X1_65/B POR2X1_174/A 0.03fF
C25067 POR2X1_294/CTRL2 D_GATE_741 0.01fF
C25068 POR2X1_850/A POR2X1_121/B 0.03fF
C25069 POR2X1_20/B PAND2X1_182/CTRL 0.01fF
C25070 PAND2X1_73/Y POR2X1_455/O 0.02fF
C25071 POR2X1_477/A POR2X1_434/CTRL2 0.00fF
C25072 POR2X1_83/B PAND2X1_180/CTRL 0.01fF
C25073 PAND2X1_57/B PAND2X1_591/O 0.01fF
C25074 POR2X1_337/A POR2X1_814/A 0.03fF
C25075 PAND2X1_75/m4_208_n4# POR2X1_574/m4_208_n4# 0.13fF
C25076 PAND2X1_644/Y PAND2X1_758/CTRL2 0.00fF
C25077 POR2X1_150/Y PAND2X1_186/a_16_344# 0.02fF
C25078 PAND2X1_11/Y PAND2X1_18/a_16_344# 0.02fF
C25079 POR2X1_860/A POR2X1_777/B 0.03fF
C25080 POR2X1_302/A POR2X1_260/B 0.12fF
C25081 POR2X1_20/B PAND2X1_785/a_16_344# 0.01fF
C25082 PAND2X1_96/B POR2X1_341/A 2.33fF
C25083 POR2X1_254/Y PAND2X1_73/Y 0.05fF
C25084 POR2X1_94/CTRL2 POR2X1_23/Y 0.07fF
C25085 POR2X1_311/Y PAND2X1_362/B 2.02fF
C25086 POR2X1_760/A PAND2X1_717/Y 0.07fF
C25087 PAND2X1_859/A POR2X1_226/Y 0.99fF
C25088 PAND2X1_615/O INPUT_3 0.06fF
C25089 POR2X1_487/m4_208_n4# PAND2X1_738/Y 0.04fF
C25090 POR2X1_66/A POR2X1_664/Y 0.02fF
C25091 PAND2X1_106/CTRL2 POR2X1_556/A 0.01fF
C25092 PAND2X1_611/CTRL POR2X1_249/Y 0.01fF
C25093 PAND2X1_777/O POR2X1_7/B 0.05fF
C25094 POR2X1_407/A POR2X1_866/A 0.03fF
C25095 POR2X1_65/A PAND2X1_231/O 0.07fF
C25096 PAND2X1_429/O INPUT_5 0.01fF
C25097 POR2X1_72/Y POR2X1_32/A 0.05fF
C25098 PAND2X1_65/B POR2X1_860/A 0.03fF
C25099 POR2X1_640/a_16_28# POR2X1_640/A 0.09fF
C25100 POR2X1_686/A PAND2X1_65/B 0.16fF
C25101 POR2X1_68/A POR2X1_678/Y 0.07fF
C25102 POR2X1_155/O POR2X1_467/Y 0.02fF
C25103 POR2X1_775/A POR2X1_66/A 0.03fF
C25104 POR2X1_376/B POR2X1_677/a_56_344# 0.03fF
C25105 POR2X1_861/O POR2X1_218/Y 0.04fF
C25106 POR2X1_333/Y POR2X1_814/A 0.03fF
C25107 PAND2X1_787/Y PAND2X1_562/B 0.10fF
C25108 PAND2X1_613/O POR2X1_68/B 0.07fF
C25109 INPUT_0 POR2X1_40/Y 0.21fF
C25110 POR2X1_472/O POR2X1_472/B 0.01fF
C25111 PAND2X1_460/Y POR2X1_94/A 0.01fF
C25112 PAND2X1_73/Y POR2X1_575/B 0.01fF
C25113 PAND2X1_808/m4_208_n4# POR2X1_437/m4_208_n4# 0.05fF
C25114 POR2X1_69/A POR2X1_7/B 0.03fF
C25115 POR2X1_68/A POR2X1_29/A 0.14fF
C25116 POR2X1_302/B PAND2X1_322/O 0.02fF
C25117 PAND2X1_738/Y PAND2X1_714/A 0.10fF
C25118 PAND2X1_23/Y POR2X1_634/A 0.03fF
C25119 PAND2X1_287/Y PAND2X1_568/B 0.84fF
C25120 PAND2X1_90/CTRL POR2X1_814/A 0.01fF
C25121 POR2X1_356/A POR2X1_436/O 0.02fF
C25122 POR2X1_801/A VDD 0.00fF
C25123 PAND2X1_201/CTRL2 PAND2X1_358/A 0.02fF
C25124 POR2X1_529/a_16_28# POR2X1_29/A 0.09fF
C25125 POR2X1_65/A POR2X1_424/CTRL 0.00fF
C25126 PAND2X1_90/A PAND2X1_73/a_16_344# 0.01fF
C25127 POR2X1_78/B POR2X1_370/Y 0.03fF
C25128 POR2X1_13/A PAND2X1_787/Y 0.05fF
C25129 POR2X1_623/B D_INPUT_1 0.01fF
C25130 PAND2X1_740/a_76_28# PAND2X1_738/Y 0.04fF
C25131 PAND2X1_576/B PAND2X1_656/A 1.07fF
C25132 PAND2X1_859/a_76_28# POR2X1_13/A 0.02fF
C25133 D_INPUT_5 POR2X1_260/A 0.11fF
C25134 PAND2X1_630/B POR2X1_39/B 0.03fF
C25135 PAND2X1_467/Y PAND2X1_452/O 0.02fF
C25136 PAND2X1_480/B POR2X1_236/Y 0.00fF
C25137 POR2X1_305/Y PAND2X1_784/A 0.02fF
C25138 POR2X1_852/B PAND2X1_55/Y 0.13fF
C25139 PAND2X1_770/O VDD 0.00fF
C25140 POR2X1_809/B VDD 0.10fF
C25141 POR2X1_23/Y POR2X1_171/CTRL2 0.01fF
C25142 POR2X1_41/B PAND2X1_833/CTRL 0.07fF
C25143 POR2X1_743/CTRL POR2X1_7/B 0.01fF
C25144 POR2X1_149/B POR2X1_605/B 0.04fF
C25145 PAND2X1_55/CTRL2 PAND2X1_55/Y 0.01fF
C25146 PAND2X1_6/Y POR2X1_457/CTRL 0.01fF
C25147 PAND2X1_798/B PAND2X1_390/Y 0.03fF
C25148 POR2X1_49/Y POR2X1_45/Y 0.03fF
C25149 POR2X1_219/B PAND2X1_394/O 0.03fF
C25150 PAND2X1_341/B POR2X1_65/a_56_344# 0.00fF
C25151 POR2X1_121/B PAND2X1_536/m4_208_n4# 0.15fF
C25152 PAND2X1_803/A PAND2X1_724/B 0.03fF
C25153 POR2X1_525/Y PAND2X1_712/B 0.02fF
C25154 POR2X1_97/A POR2X1_212/CTRL 0.03fF
C25155 POR2X1_366/O PAND2X1_93/B 0.02fF
C25156 PAND2X1_558/CTRL PAND2X1_493/Y 0.02fF
C25157 PAND2X1_468/CTRL VDD 0.00fF
C25158 POR2X1_614/A PAND2X1_582/O 0.18fF
C25159 PAND2X1_205/B VDD 0.02fF
C25160 POR2X1_862/B PAND2X1_536/O 0.00fF
C25161 POR2X1_231/A POR2X1_231/a_16_28# 0.03fF
C25162 POR2X1_805/A POR2X1_710/A 0.03fF
C25163 POR2X1_274/O POR2X1_569/A 0.04fF
C25164 POR2X1_7/B PAND2X1_730/B 0.02fF
C25165 PAND2X1_394/a_16_344# PAND2X1_88/Y 0.01fF
C25166 PAND2X1_272/CTRL2 POR2X1_553/A 0.01fF
C25167 PAND2X1_90/A PAND2X1_80/CTRL 0.01fF
C25168 POR2X1_32/A PAND2X1_349/A 0.03fF
C25169 POR2X1_188/A PAND2X1_752/Y 0.01fF
C25170 POR2X1_13/A PAND2X1_668/CTRL 0.01fF
C25171 POR2X1_706/CTRL POR2X1_383/A 0.01fF
C25172 PAND2X1_90/Y PAND2X1_145/O 0.04fF
C25173 POR2X1_32/A PAND2X1_63/B 0.03fF
C25174 POR2X1_16/A PAND2X1_640/B 0.03fF
C25175 GATE_741 POR2X1_7/B 0.03fF
C25176 POR2X1_355/B POR2X1_190/Y 0.01fF
C25177 PAND2X1_96/B POR2X1_500/A 0.01fF
C25178 POR2X1_96/A POR2X1_693/O 0.00fF
C25179 PAND2X1_242/CTRL POR2X1_511/Y 0.03fF
C25180 PAND2X1_41/B PAND2X1_518/CTRL 0.01fF
C25181 PAND2X1_94/A PAND2X1_282/CTRL 0.03fF
C25182 POR2X1_296/B POR2X1_569/A 0.07fF
C25183 POR2X1_444/A POR2X1_545/O 0.05fF
C25184 POR2X1_99/A PAND2X1_88/Y 0.05fF
C25185 PAND2X1_23/Y POR2X1_130/A 0.10fF
C25186 POR2X1_846/B VDD 0.01fF
C25187 PAND2X1_725/Y POR2X1_152/Y 0.11fF
C25188 POR2X1_528/Y POR2X1_14/Y 0.04fF
C25189 INPUT_0 PAND2X1_188/a_16_344# 0.02fF
C25190 PAND2X1_377/O POR2X1_42/Y 0.07fF
C25191 POR2X1_514/Y VDD 0.00fF
C25192 INPUT_1 PAND2X1_623/CTRL 0.01fF
C25193 PAND2X1_23/Y POR2X1_566/A 0.05fF
C25194 POR2X1_497/Y POR2X1_521/CTRL 0.00fF
C25195 POR2X1_528/Y PAND2X1_453/A 0.75fF
C25196 POR2X1_379/Y POR2X1_260/B 0.05fF
C25197 POR2X1_502/A PAND2X1_95/B 2.79fF
C25198 POR2X1_693/Y VDD 0.26fF
C25199 POR2X1_553/Y POR2X1_554/Y 0.09fF
C25200 POR2X1_90/Y POR2X1_5/Y 0.15fF
C25201 POR2X1_567/A POR2X1_854/O 0.03fF
C25202 POR2X1_29/A POR2X1_391/B 0.01fF
C25203 PAND2X1_570/CTRL VDD 0.00fF
C25204 POR2X1_675/A POR2X1_540/A 0.00fF
C25205 POR2X1_45/Y PAND2X1_274/O 0.00fF
C25206 PAND2X1_829/CTRL POR2X1_260/A 0.01fF
C25207 PAND2X1_6/Y POR2X1_464/O 0.01fF
C25208 PAND2X1_96/B PAND2X1_58/CTRL2 0.03fF
C25209 PAND2X1_550/a_76_28# PAND2X1_546/Y 0.02fF
C25210 POR2X1_41/B PAND2X1_35/CTRL 0.00fF
C25211 POR2X1_68/A POR2X1_546/A 0.03fF
C25212 POR2X1_72/B PAND2X1_549/B 0.13fF
C25213 PAND2X1_6/A POR2X1_224/CTRL 0.10fF
C25214 PAND2X1_91/CTRL POR2X1_191/Y -0.01fF
C25215 PAND2X1_91/a_16_344# POR2X1_192/B 0.02fF
C25216 POR2X1_685/CTRL POR2X1_685/B 0.00fF
C25217 POR2X1_111/O POR2X1_5/Y 0.02fF
C25218 PAND2X1_627/O PAND2X1_69/A 0.15fF
C25219 POR2X1_402/A POR2X1_401/B 0.02fF
C25220 PAND2X1_42/O PAND2X1_111/B 0.02fF
C25221 POR2X1_66/A POR2X1_339/Y 0.03fF
C25222 POR2X1_119/Y PAND2X1_444/O 0.15fF
C25223 PAND2X1_439/O POR2X1_167/Y 0.02fF
C25224 PAND2X1_281/a_76_28# POR2X1_643/Y 0.03fF
C25225 POR2X1_260/Y POR2X1_205/Y 0.17fF
C25226 POR2X1_383/A POR2X1_654/B 0.03fF
C25227 PAND2X1_41/B POR2X1_854/B 0.06fF
C25228 POR2X1_45/Y PAND2X1_553/B 0.00fF
C25229 POR2X1_528/CTRL POR2X1_56/B 0.01fF
C25230 POR2X1_156/B VDD 0.18fF
C25231 POR2X1_226/Y POR2X1_7/A 0.03fF
C25232 POR2X1_174/a_16_28# POR2X1_174/A 0.05fF
C25233 PAND2X1_484/O POR2X1_590/A 0.04fF
C25234 POR2X1_836/CTRL POR2X1_192/B 0.07fF
C25235 POR2X1_383/A POR2X1_850/A 0.07fF
C25236 POR2X1_525/Y PAND2X1_546/CTRL2 0.01fF
C25237 POR2X1_260/Y POR2X1_205/O 0.00fF
C25238 PAND2X1_446/Y POR2X1_77/Y 0.05fF
C25239 POR2X1_249/Y POR2X1_734/A 0.04fF
C25240 POR2X1_65/A PAND2X1_569/B 0.14fF
C25241 POR2X1_83/B POR2X1_129/Y 0.04fF
C25242 POR2X1_65/A POR2X1_158/B 0.02fF
C25243 POR2X1_416/B INPUT_3 0.05fF
C25244 PAND2X1_245/CTRL2 PAND2X1_48/A 0.01fF
C25245 POR2X1_135/Y POR2X1_136/Y 0.00fF
C25246 POR2X1_51/A POR2X1_36/O 0.01fF
C25247 PAND2X1_357/Y POR2X1_55/Y 3.08fF
C25248 POR2X1_775/A POR2X1_222/Y 0.03fF
C25249 PAND2X1_773/B PAND2X1_854/A 0.25fF
C25250 PAND2X1_461/CTRL POR2X1_612/Y 0.06fF
C25251 PAND2X1_442/CTRL POR2X1_568/Y 0.01fF
C25252 POR2X1_178/Y PAND2X1_540/a_76_28# 0.02fF
C25253 PAND2X1_674/a_16_344# POR2X1_732/B 0.05fF
C25254 POR2X1_81/A POR2X1_23/Y 0.03fF
C25255 POR2X1_417/CTRL POR2X1_372/Y 0.08fF
C25256 POR2X1_529/Y VDD 0.15fF
C25257 POR2X1_78/B PAND2X1_63/B 0.03fF
C25258 POR2X1_57/A PAND2X1_793/Y 0.03fF
C25259 POR2X1_416/B POR2X1_428/Y 0.06fF
C25260 PAND2X1_23/Y POR2X1_363/a_16_28# 0.03fF
C25261 PAND2X1_48/B POR2X1_205/m4_208_n4# 0.17fF
C25262 PAND2X1_657/a_16_344# PAND2X1_657/B 0.03fF
C25263 POR2X1_43/B PAND2X1_228/a_76_28# 0.04fF
C25264 PAND2X1_90/Y PAND2X1_313/CTRL2 0.02fF
C25265 POR2X1_258/Y VDD 0.01fF
C25266 POR2X1_698/O POR2X1_394/A 0.02fF
C25267 POR2X1_455/CTRL2 POR2X1_456/B 0.00fF
C25268 PAND2X1_94/A POR2X1_410/CTRL2 0.02fF
C25269 PAND2X1_659/Y POR2X1_83/B 0.03fF
C25270 POR2X1_664/Y POR2X1_532/A 0.03fF
C25271 POR2X1_848/A POR2X1_39/B 0.13fF
C25272 PAND2X1_59/B D_INPUT_4 0.79fF
C25273 POR2X1_222/Y POR2X1_112/Y 0.12fF
C25274 PAND2X1_23/Y POR2X1_573/A 0.03fF
C25275 POR2X1_383/A PAND2X1_52/m4_208_n4# 0.14fF
C25276 POR2X1_514/Y PAND2X1_32/B 0.21fF
C25277 POR2X1_13/A POR2X1_103/Y 0.00fF
C25278 POR2X1_539/A POR2X1_220/Y 0.03fF
C25279 POR2X1_685/A POR2X1_728/B 0.12fF
C25280 POR2X1_96/A POR2X1_235/Y 0.04fF
C25281 PAND2X1_428/O PAND2X1_48/A 0.04fF
C25282 PAND2X1_371/a_76_28# POR2X1_68/B 0.07fF
C25283 PAND2X1_244/B PAND2X1_734/B 0.01fF
C25284 PAND2X1_8/Y PAND2X1_133/O 0.04fF
C25285 PAND2X1_857/A POR2X1_821/a_16_28# 0.03fF
C25286 INPUT_1 POR2X1_625/m4_208_n4# 0.01fF
C25287 POR2X1_96/Y POR2X1_83/B 15.86fF
C25288 POR2X1_57/A PAND2X1_334/CTRL2 0.03fF
C25289 POR2X1_590/A POR2X1_199/B 0.00fF
C25290 POR2X1_773/B VDD 1.26fF
C25291 PAND2X1_96/B PAND2X1_176/m4_208_n4# 0.15fF
C25292 POR2X1_281/a_16_28# POR2X1_236/Y 0.04fF
C25293 POR2X1_459/B PAND2X1_69/A 0.00fF
C25294 POR2X1_407/A POR2X1_501/B 0.89fF
C25295 PAND2X1_835/a_16_344# POR2X1_821/Y 0.02fF
C25296 POR2X1_398/Y POR2X1_398/O 0.00fF
C25297 PAND2X1_140/A POR2X1_55/Y 0.03fF
C25298 POR2X1_365/Y POR2X1_212/O 0.10fF
C25299 POR2X1_732/m4_208_n4# PAND2X1_152/m4_208_n4# 0.05fF
C25300 POR2X1_23/Y PAND2X1_327/O 0.03fF
C25301 POR2X1_57/A POR2X1_665/Y 0.31fF
C25302 POR2X1_122/a_16_28# POR2X1_40/Y 0.00fF
C25303 POR2X1_508/A POR2X1_355/A 0.01fF
C25304 POR2X1_391/B POR2X1_546/A 0.09fF
C25305 POR2X1_313/Y POR2X1_13/A 0.02fF
C25306 PAND2X1_99/O PAND2X1_97/Y 0.08fF
C25307 POR2X1_60/A PAND2X1_326/B 0.03fF
C25308 PAND2X1_48/B POR2X1_725/Y 0.07fF
C25309 POR2X1_68/B PAND2X1_518/CTRL2 0.01fF
C25310 POR2X1_528/Y POR2X1_55/Y 0.10fF
C25311 PAND2X1_96/B PAND2X1_767/O 0.11fF
C25312 POR2X1_72/B PAND2X1_330/CTRL 0.01fF
C25313 PAND2X1_636/CTRL2 POR2X1_583/Y 0.01fF
C25314 PAND2X1_144/O PAND2X1_60/B 0.17fF
C25315 PAND2X1_109/CTRL POR2X1_78/A 0.01fF
C25316 POR2X1_691/CTRL2 POR2X1_855/B 0.02fF
C25317 POR2X1_691/O POR2X1_691/B 0.04fF
C25318 PAND2X1_4/O PAND2X1_6/A 0.02fF
C25319 PAND2X1_866/A PAND2X1_865/Y 0.01fF
C25320 POR2X1_614/A POR2X1_812/B 0.05fF
C25321 POR2X1_299/O POR2X1_90/Y 0.01fF
C25322 POR2X1_532/A POR2X1_112/Y 0.03fF
C25323 PAND2X1_383/CTRL2 POR2X1_816/A 0.01fF
C25324 POR2X1_96/O PAND2X1_472/B 0.01fF
C25325 PAND2X1_79/CTRL2 POR2X1_569/A 0.02fF
C25326 POR2X1_63/CTRL PAND2X1_63/B 0.01fF
C25327 PAND2X1_435/CTRL2 POR2X1_153/Y 0.03fF
C25328 GATE_479 POR2X1_119/Y 0.01fF
C25329 POR2X1_16/A POR2X1_7/B 0.07fF
C25330 POR2X1_518/a_16_28# POR2X1_667/A 0.02fF
C25331 POR2X1_52/A PAND2X1_726/B 0.13fF
C25332 PAND2X1_693/CTRL2 PAND2X1_94/A 0.03fF
C25333 POR2X1_110/Y POR2X1_5/Y 0.01fF
C25334 POR2X1_184/Y PAND2X1_349/A 5.12fF
C25335 POR2X1_569/A POR2X1_501/O 0.04fF
C25336 POR2X1_78/A PAND2X1_56/A 0.03fF
C25337 POR2X1_48/A POR2X1_167/Y 0.00fF
C25338 POR2X1_25/O PAND2X1_18/B 0.05fF
C25339 PAND2X1_6/Y POR2X1_510/Y 0.05fF
C25340 POR2X1_278/Y PAND2X1_560/B 0.42fF
C25341 POR2X1_239/CTRL POR2X1_239/Y 0.01fF
C25342 INPUT_1 POR2X1_294/B 1.63fF
C25343 POR2X1_712/A POR2X1_712/a_16_28# 0.07fF
C25344 POR2X1_341/a_16_28# POR2X1_228/Y -0.00fF
C25345 PAND2X1_94/A POR2X1_264/Y 0.05fF
C25346 POR2X1_75/CTRL PAND2X1_349/A 0.01fF
C25347 POR2X1_326/a_76_344# POR2X1_468/B 0.03fF
C25348 PAND2X1_533/CTRL2 POR2X1_532/Y 0.01fF
C25349 PAND2X1_651/Y PAND2X1_349/A 0.03fF
C25350 POR2X1_114/CTRL2 POR2X1_101/Y 0.12fF
C25351 PAND2X1_359/a_16_344# PAND2X1_348/Y 0.03fF
C25352 PAND2X1_57/B POR2X1_398/O 0.01fF
C25353 PAND2X1_836/a_76_28# POR2X1_823/Y 0.07fF
C25354 POR2X1_25/a_16_28# POR2X1_3/B 0.04fF
C25355 POR2X1_548/a_76_344# POR2X1_620/B 0.01fF
C25356 POR2X1_110/Y PAND2X1_549/CTRL2 0.01fF
C25357 POR2X1_452/A POR2X1_450/Y 0.03fF
C25358 POR2X1_514/O POR2X1_101/Y 0.04fF
C25359 POR2X1_296/B PAND2X1_72/A 0.16fF
C25360 PAND2X1_844/CTRL POR2X1_293/Y 0.02fF
C25361 PAND2X1_483/a_16_344# POR2X1_55/Y 0.01fF
C25362 POR2X1_502/A POR2X1_722/CTRL2 0.01fF
C25363 PAND2X1_6/Y POR2X1_348/a_76_344# 0.01fF
C25364 POR2X1_855/B POR2X1_644/A 0.04fF
C25365 PAND2X1_48/B POR2X1_559/A 0.08fF
C25366 PAND2X1_661/Y POR2X1_73/Y 0.07fF
C25367 PAND2X1_6/Y POR2X1_276/Y 0.50fF
C25368 POR2X1_367/a_16_28# POR2X1_192/B 0.07fF
C25369 POR2X1_367/a_76_344# POR2X1_191/Y 0.02fF
C25370 POR2X1_65/A PAND2X1_798/Y 0.03fF
C25371 POR2X1_730/Y POR2X1_467/CTRL2 0.01fF
C25372 PAND2X1_659/Y PAND2X1_795/B 0.03fF
C25373 PAND2X1_23/Y POR2X1_344/Y 0.03fF
C25374 PAND2X1_314/CTRL POR2X1_854/B 0.14fF
C25375 POR2X1_707/B PAND2X1_52/B 0.64fF
C25376 POR2X1_750/Y PAND2X1_69/A 0.01fF
C25377 POR2X1_95/CTRL2 POR2X1_51/A 0.01fF
C25378 PAND2X1_55/Y POR2X1_151/Y 0.01fF
C25379 POR2X1_137/Y POR2X1_361/m4_208_n4# 0.15fF
C25380 POR2X1_768/Y POR2X1_294/B 0.03fF
C25381 POR2X1_773/B PAND2X1_32/B 0.11fF
C25382 POR2X1_347/CTRL2 PAND2X1_57/B 0.01fF
C25383 PAND2X1_117/O PAND2X1_48/A 0.15fF
C25384 PAND2X1_716/B POR2X1_372/Y 0.08fF
C25385 POR2X1_326/A POR2X1_662/Y 0.03fF
C25386 POR2X1_415/A POR2X1_67/Y 0.01fF
C25387 POR2X1_408/Y POR2X1_583/a_16_28# 0.08fF
C25388 POR2X1_322/Y PAND2X1_374/CTRL 0.00fF
C25389 PAND2X1_801/a_16_344# POR2X1_236/Y 0.00fF
C25390 POR2X1_7/B PAND2X1_336/Y 0.01fF
C25391 POR2X1_245/Y POR2X1_283/A 0.04fF
C25392 POR2X1_235/Y POR2X1_7/A 0.01fF
C25393 POR2X1_196/Y PAND2X1_824/B 0.02fF
C25394 POR2X1_862/B PAND2X1_52/B 0.02fF
C25395 POR2X1_557/B POR2X1_391/Y 0.07fF
C25396 D_INPUT_3 POR2X1_96/CTRL 0.12fF
C25397 POR2X1_464/CTRL2 POR2X1_736/A 0.34fF
C25398 POR2X1_707/a_76_344# POR2X1_407/Y 0.00fF
C25399 POR2X1_681/CTRL POR2X1_681/Y 0.01fF
C25400 PAND2X1_221/Y PAND2X1_798/CTRL 0.00fF
C25401 POR2X1_456/B PAND2X1_60/B 0.07fF
C25402 POR2X1_78/A POR2X1_661/A 0.07fF
C25403 POR2X1_508/A POR2X1_508/O 0.02fF
C25404 INPUT_1 PAND2X1_111/B 0.00fF
C25405 PAND2X1_73/Y POR2X1_643/CTRL2 0.05fF
C25406 PAND2X1_652/A POR2X1_385/Y 0.07fF
C25407 PAND2X1_779/CTRL2 POR2X1_90/Y 0.03fF
C25408 PAND2X1_865/Y POR2X1_488/Y 0.01fF
C25409 POR2X1_188/O POR2X1_675/Y 0.01fF
C25410 POR2X1_130/A POR2X1_711/Y 0.10fF
C25411 POR2X1_257/A POR2X1_271/B 0.03fF
C25412 POR2X1_293/Y PAND2X1_860/O 0.04fF
C25413 POR2X1_502/CTRL POR2X1_854/B 0.31fF
C25414 POR2X1_416/B PAND2X1_740/Y 0.06fF
C25415 POR2X1_518/CTRL2 POR2X1_519/Y 0.06fF
C25416 PAND2X1_850/Y POR2X1_42/Y 0.70fF
C25417 POR2X1_416/B POR2X1_13/O 0.01fF
C25418 POR2X1_318/O POR2X1_445/A 0.01fF
C25419 POR2X1_218/CTRL POR2X1_260/A 0.00fF
C25420 POR2X1_49/Y PAND2X1_147/CTRL2 0.01fF
C25421 POR2X1_62/Y POR2X1_68/B 0.03fF
C25422 POR2X1_456/B POR2X1_737/CTRL 0.01fF
C25423 PAND2X1_632/B PAND2X1_632/O 0.00fF
C25424 PAND2X1_555/Y PAND2X1_345/Y 0.02fF
C25425 PAND2X1_620/O POR2X1_588/Y 0.00fF
C25426 POR2X1_42/CTRL2 POR2X1_4/Y 0.06fF
C25427 POR2X1_411/B PAND2X1_35/A 0.12fF
C25428 POR2X1_447/B PAND2X1_69/A 0.05fF
C25429 PAND2X1_683/O POR2X1_596/A 0.02fF
C25430 INPUT_6 PAND2X1_3/B 3.03fF
C25431 POR2X1_508/O POR2X1_568/B 0.07fF
C25432 POR2X1_490/Y PAND2X1_217/CTRL 0.01fF
C25433 POR2X1_411/Y POR2X1_416/B 0.01fF
C25434 POR2X1_188/A POR2X1_643/a_56_344# -0.00fF
C25435 PAND2X1_699/CTRL POR2X1_496/Y 0.05fF
C25436 POR2X1_329/A POR2X1_516/Y 14.95fF
C25437 PAND2X1_254/a_16_344# POR2X1_77/Y 0.01fF
C25438 POR2X1_191/B POR2X1_568/Y 0.05fF
C25439 PAND2X1_462/CTRL2 POR2X1_416/Y 0.01fF
C25440 POR2X1_591/O POR2X1_77/Y 0.18fF
C25441 POR2X1_332/B PAND2X1_135/O 0.02fF
C25442 POR2X1_54/Y POR2X1_815/Y 0.44fF
C25443 POR2X1_158/Y PAND2X1_707/Y 0.66fF
C25444 PAND2X1_63/B POR2X1_294/A 0.03fF
C25445 POR2X1_654/B POR2X1_643/a_16_28# 0.07fF
C25446 POR2X1_119/Y PAND2X1_175/B 0.05fF
C25447 PAND2X1_675/A POR2X1_416/B 9.89fF
C25448 POR2X1_437/CTRL2 POR2X1_385/Y 0.14fF
C25449 PAND2X1_206/B POR2X1_69/A 0.88fF
C25450 POR2X1_416/B PAND2X1_469/B 0.03fF
C25451 POR2X1_832/O POR2X1_661/A 0.05fF
C25452 POR2X1_633/A POR2X1_633/CTRL2 0.01fF
C25453 PAND2X1_39/B POR2X1_218/Y 0.07fF
C25454 POR2X1_77/CTRL POR2X1_48/A 0.03fF
C25455 POR2X1_296/Y POR2X1_296/O 0.06fF
C25456 POR2X1_490/Y PAND2X1_267/Y 0.06fF
C25457 INPUT_3 POR2X1_623/B 0.04fF
C25458 POR2X1_267/Y PAND2X1_72/A 0.22fF
C25459 POR2X1_447/B PAND2X1_823/O 0.15fF
C25460 POR2X1_359/B POR2X1_363/A -0.02fF
C25461 POR2X1_804/A POR2X1_715/CTRL2 0.01fF
C25462 POR2X1_659/a_76_344# POR2X1_750/B 0.04fF
C25463 POR2X1_48/A POR2X1_848/A 0.07fF
C25464 PAND2X1_94/Y PAND2X1_57/B 0.02fF
C25465 POR2X1_510/Y POR2X1_632/Y 25.11fF
C25466 POR2X1_454/CTRL2 POR2X1_454/B 0.01fF
C25467 POR2X1_447/B PAND2X1_824/B 0.09fF
C25468 POR2X1_60/A POR2X1_253/O 0.18fF
C25469 POR2X1_101/Y PAND2X1_136/O 0.04fF
C25470 POR2X1_416/A POR2X1_416/a_16_28# 0.05fF
C25471 PAND2X1_86/O PAND2X1_85/Y 0.00fF
C25472 POR2X1_567/O POR2X1_854/B 0.04fF
C25473 PAND2X1_240/CTRL POR2X1_411/B 0.01fF
C25474 POR2X1_287/B POR2X1_705/B 0.05fF
C25475 POR2X1_14/Y POR2X1_816/Y 0.03fF
C25476 POR2X1_65/A POR2X1_603/O 0.02fF
C25477 POR2X1_600/O VDD 0.00fF
C25478 PAND2X1_404/Y PAND2X1_573/B 0.20fF
C25479 POR2X1_559/A PAND2X1_517/CTRL 0.02fF
C25480 PAND2X1_294/a_76_28# POR2X1_60/A 0.05fF
C25481 POR2X1_119/Y PAND2X1_858/O 0.13fF
C25482 PAND2X1_477/O POR2X1_102/Y 0.04fF
C25483 POR2X1_88/O POR2X1_69/A 0.01fF
C25484 PAND2X1_340/B POR2X1_40/Y 0.03fF
C25485 PAND2X1_771/Y PAND2X1_542/O 0.06fF
C25486 POR2X1_602/B PAND2X1_601/O 0.02fF
C25487 PAND2X1_824/B POR2X1_510/O 0.02fF
C25488 D_INPUT_0 POR2X1_413/CTRL 0.01fF
C25489 POR2X1_302/Y POR2X1_287/A 0.02fF
C25490 POR2X1_540/Y POR2X1_337/Y 0.40fF
C25491 POR2X1_126/O POR2X1_94/A 0.01fF
C25492 POR2X1_520/O PAND2X1_52/B 0.01fF
C25493 POR2X1_83/B POR2X1_37/Y 0.25fF
C25494 POR2X1_98/A POR2X1_35/Y 0.02fF
C25495 D_INPUT_5 PAND2X1_588/CTRL 0.01fF
C25496 POR2X1_227/B VDD 0.13fF
C25497 POR2X1_862/A PAND2X1_41/B 0.10fF
C25498 PAND2X1_853/B POR2X1_39/B 0.03fF
C25499 POR2X1_129/Y PAND2X1_841/Y 0.02fF
C25500 POR2X1_188/A POR2X1_851/A 0.01fF
C25501 POR2X1_744/Y VDD 0.17fF
C25502 D_INPUT_7 PAND2X1_587/O 0.03fF
C25503 POR2X1_66/B POR2X1_66/A 2.27fF
C25504 PAND2X1_205/Y PAND2X1_267/Y 0.02fF
C25505 POR2X1_661/A POR2X1_513/CTRL2 0.02fF
C25506 POR2X1_448/CTRL POR2X1_296/B 0.08fF
C25507 PAND2X1_58/A POR2X1_29/A 0.14fF
C25508 POR2X1_471/A VDD 0.46fF
C25509 POR2X1_502/A POR2X1_444/O 0.02fF
C25510 PAND2X1_230/CTRL2 POR2X1_78/A 0.03fF
C25511 POR2X1_260/B POR2X1_285/CTRL2 0.01fF
C25512 POR2X1_661/A PAND2X1_306/O 0.11fF
C25513 POR2X1_188/A POR2X1_66/A 0.03fF
C25514 PAND2X1_576/B PAND2X1_576/CTRL 0.01fF
C25515 PAND2X1_687/a_56_28# POR2X1_761/A 0.00fF
C25516 POR2X1_559/CTRL POR2X1_814/A 0.01fF
C25517 POR2X1_590/Y PAND2X1_72/A 0.01fF
C25518 POR2X1_355/CTRL POR2X1_567/B 0.00fF
C25519 POR2X1_376/B POR2X1_817/CTRL 0.01fF
C25520 POR2X1_417/Y POR2X1_32/A 0.03fF
C25521 POR2X1_49/Y PAND2X1_796/CTRL2 0.01fF
C25522 POR2X1_776/A POR2X1_776/B 15.73fF
C25523 POR2X1_60/A POR2X1_251/CTRL2 0.11fF
C25524 POR2X1_634/A PAND2X1_428/CTRL2 0.06fF
C25525 POR2X1_23/Y PAND2X1_499/Y 0.05fF
C25526 PAND2X1_57/B POR2X1_648/a_16_28# 0.01fF
C25527 POR2X1_856/CTRL PAND2X1_73/Y 0.01fF
C25528 POR2X1_102/Y POR2X1_40/Y 4.73fF
C25529 PAND2X1_73/Y PAND2X1_41/B 1.59fF
C25530 POR2X1_16/A POR2X1_16/CTRL 0.01fF
C25531 POR2X1_78/B POR2X1_567/B 0.10fF
C25532 POR2X1_777/B POR2X1_121/B 0.18fF
C25533 POR2X1_786/A POR2X1_266/CTRL2 0.01fF
C25534 POR2X1_114/B POR2X1_499/A 0.02fF
C25535 POR2X1_154/a_16_28# PAND2X1_39/B 0.03fF
C25536 POR2X1_554/B POR2X1_513/Y 0.03fF
C25537 INPUT_3 POR2X1_619/CTRL2 0.01fF
C25538 POR2X1_705/B POR2X1_705/CTRL2 0.00fF
C25539 PAND2X1_611/O POR2X1_68/B 0.16fF
C25540 POR2X1_43/B POR2X1_411/B 0.10fF
C25541 POR2X1_829/A PAND2X1_207/CTRL2 0.00fF
C25542 POR2X1_218/Y POR2X1_325/A 0.07fF
C25543 POR2X1_69/A POR2X1_750/B 0.03fF
C25544 POR2X1_814/A POR2X1_360/CTRL 0.07fF
C25545 PAND2X1_258/CTRL POR2X1_244/B 0.01fF
C25546 PAND2X1_618/a_76_28# PAND2X1_6/A 0.02fF
C25547 POR2X1_334/B POR2X1_473/CTRL 0.04fF
C25548 PAND2X1_215/O PAND2X1_205/Y -0.00fF
C25549 POR2X1_489/B POR2X1_287/B 0.01fF
C25550 POR2X1_260/B POR2X1_231/B 0.00fF
C25551 PAND2X1_612/B POR2X1_642/CTRL 0.00fF
C25552 POR2X1_96/A PAND2X1_771/Y 0.02fF
C25553 PAND2X1_90/A PAND2X1_613/O 0.01fF
C25554 PAND2X1_65/B POR2X1_121/B 0.03fF
C25555 POR2X1_68/A PAND2X1_39/B 0.11fF
C25556 PAND2X1_137/Y POR2X1_48/A 0.03fF
C25557 POR2X1_441/Y POR2X1_438/a_56_344# 0.00fF
C25558 POR2X1_499/A POR2X1_458/B 0.01fF
C25559 PAND2X1_37/CTRL VDD 0.00fF
C25560 PAND2X1_462/B PAND2X1_606/O 0.15fF
C25561 POR2X1_356/A PAND2X1_237/O 0.05fF
C25562 POR2X1_814/B POR2X1_439/CTRL 0.02fF
C25563 POR2X1_347/B POR2X1_68/CTRL 0.03fF
C25564 PAND2X1_212/B VDD 0.04fF
C25565 POR2X1_856/B POR2X1_776/B 0.01fF
C25566 POR2X1_411/B POR2X1_38/B 0.08fF
C25567 POR2X1_541/B POR2X1_532/A 0.07fF
C25568 PAND2X1_848/B PAND2X1_340/B 0.02fF
C25569 POR2X1_20/B POR2X1_382/Y 0.89fF
C25570 POR2X1_260/B POR2X1_460/B 0.04fF
C25571 POR2X1_124/B POR2X1_473/CTRL 0.15fF
C25572 POR2X1_624/Y POR2X1_576/Y 0.03fF
C25573 POR2X1_137/Y POR2X1_556/A 2.10fF
C25574 PAND2X1_65/B POR2X1_267/a_16_28# 0.03fF
C25575 POR2X1_130/A POR2X1_641/CTRL2 0.02fF
C25576 POR2X1_554/B POR2X1_366/A 0.03fF
C25577 POR2X1_120/a_76_344# POR2X1_78/A 0.00fF
C25578 PAND2X1_35/Y POR2X1_32/A 0.03fF
C25579 POR2X1_300/CTRL2 D_INPUT_0 0.09fF
C25580 POR2X1_593/B PAND2X1_589/CTRL2 0.01fF
C25581 POR2X1_260/B POR2X1_790/A 0.06fF
C25582 POR2X1_201/CTRL2 VDD 0.00fF
C25583 POR2X1_624/Y POR2X1_140/CTRL2 0.08fF
C25584 POR2X1_16/A PAND2X1_206/B 0.47fF
C25585 PAND2X1_58/A POR2X1_546/A 0.03fF
C25586 POR2X1_290/Y POR2X1_669/B 0.07fF
C25587 POR2X1_3/A POR2X1_257/A 0.04fF
C25588 POR2X1_515/a_76_344# PAND2X1_20/A 0.00fF
C25589 POR2X1_813/CTRL2 PAND2X1_63/B 0.01fF
C25590 PAND2X1_668/CTRL2 POR2X1_60/A 0.03fF
C25591 PAND2X1_658/CTRL VDD 0.00fF
C25592 PAND2X1_262/a_76_28# PAND2X1_41/B 0.01fF
C25593 POR2X1_492/CTRL2 VDD -0.00fF
C25594 POR2X1_268/Y VDD 0.10fF
C25595 PAND2X1_404/Y PAND2X1_341/A 0.03fF
C25596 PAND2X1_58/A PAND2X1_754/O 0.02fF
C25597 PAND2X1_492/CTRL PAND2X1_41/B 0.01fF
C25598 PAND2X1_860/A PAND2X1_860/CTRL2 0.01fF
C25599 POR2X1_96/A PAND2X1_575/B 0.02fF
C25600 PAND2X1_261/O POR2X1_330/Y 0.01fF
C25601 PAND2X1_48/O POR2X1_330/Y 0.03fF
C25602 POR2X1_83/B POR2X1_293/Y 0.13fF
C25603 POR2X1_118/O POR2X1_118/Y 0.01fF
C25604 PAND2X1_23/Y POR2X1_241/B 0.03fF
C25605 POR2X1_63/CTRL POR2X1_32/A 0.01fF
C25606 PAND2X1_391/CTRL2 POR2X1_816/A 0.01fF
C25607 PAND2X1_58/A PAND2X1_110/CTRL 0.01fF
C25608 PAND2X1_404/Y POR2X1_91/Y 0.07fF
C25609 PAND2X1_61/Y VDD 0.16fF
C25610 POR2X1_669/B PAND2X1_658/B 0.18fF
C25611 POR2X1_441/Y PAND2X1_714/Y 0.07fF
C25612 POR2X1_254/O POR2X1_483/B 0.00fF
C25613 PAND2X1_48/B POR2X1_811/B 0.03fF
C25614 POR2X1_274/A POR2X1_318/A 0.07fF
C25615 PAND2X1_288/A POR2X1_283/Y 0.01fF
C25616 POR2X1_616/CTRL2 POR2X1_93/A 0.00fF
C25617 PAND2X1_476/a_56_28# INPUT_0 0.00fF
C25618 POR2X1_663/O PAND2X1_90/Y 0.02fF
C25619 PAND2X1_699/CTRL2 POR2X1_129/Y 0.05fF
C25620 PAND2X1_831/O PAND2X1_785/Y 0.01fF
C25621 POR2X1_32/A POR2X1_184/Y 0.03fF
C25622 POR2X1_718/CTRL POR2X1_435/Y 0.01fF
C25623 PAND2X1_795/a_16_344# PAND2X1_785/Y 0.02fF
C25624 POR2X1_135/Y PAND2X1_332/a_16_344# 0.01fF
C25625 PAND2X1_859/A POR2X1_817/A 0.00fF
C25626 POR2X1_707/B PAND2X1_95/B 0.02fF
C25627 POR2X1_174/B D_GATE_222 0.10fF
C25628 PAND2X1_484/CTRL2 POR2X1_705/B 0.00fF
C25629 POR2X1_397/Y POR2X1_236/Y 0.00fF
C25630 POR2X1_200/CTRL POR2X1_294/B 0.08fF
C25631 POR2X1_75/CTRL POR2X1_32/A 0.01fF
C25632 INPUT_0 POR2X1_5/Y 0.28fF
C25633 PAND2X1_94/CTRL2 PAND2X1_60/B 0.01fF
C25634 PAND2X1_651/Y POR2X1_32/A 0.02fF
C25635 POR2X1_356/A POR2X1_186/Y 0.19fF
C25636 PAND2X1_857/CTRL2 POR2X1_329/A 0.03fF
C25637 POR2X1_16/A POR2X1_65/Y 0.11fF
C25638 PAND2X1_94/A POR2X1_624/Y 0.05fF
C25639 PAND2X1_604/CTRL POR2X1_750/B 0.00fF
C25640 PAND2X1_119/CTRL2 PAND2X1_73/Y 0.09fF
C25641 POR2X1_68/A PAND2X1_20/A 2.53fF
C25642 PAND2X1_58/A POR2X1_712/Y 0.03fF
C25643 POR2X1_66/B POR2X1_222/Y 18.75fF
C25644 POR2X1_628/Y POR2X1_260/A 0.03fF
C25645 POR2X1_752/Y POR2X1_293/Y 0.17fF
C25646 POR2X1_526/O POR2X1_669/B 0.06fF
C25647 PAND2X1_741/O PAND2X1_741/B 0.06fF
C25648 POR2X1_60/A PAND2X1_794/B 2.11fF
C25649 POR2X1_502/A PAND2X1_589/O 0.05fF
C25650 POR2X1_55/a_16_28# PAND2X1_6/A 0.00fF
C25651 PAND2X1_48/B PAND2X1_387/CTRL2 0.03fF
C25652 PAND2X1_597/O POR2X1_513/B 0.05fF
C25653 POR2X1_37/Y POR2X1_380/A 0.01fF
C25654 POR2X1_43/B POR2X1_271/Y 0.14fF
C25655 POR2X1_593/B POR2X1_832/B 0.00fF
C25656 PAND2X1_859/A POR2X1_42/Y 0.05fF
C25657 PAND2X1_16/O POR2X1_785/A 0.01fF
C25658 POR2X1_260/B POR2X1_375/CTRL 0.01fF
C25659 POR2X1_632/a_16_28# POR2X1_510/Y 0.01fF
C25660 PAND2X1_752/a_16_344# PAND2X1_32/B 0.01fF
C25661 PAND2X1_667/O POR2X1_546/A 0.03fF
C25662 POR2X1_362/Y POR2X1_840/B 0.19fF
C25663 POR2X1_16/A POR2X1_88/O 0.00fF
C25664 PAND2X1_128/O POR2X1_127/Y 0.02fF
C25665 PAND2X1_140/A POR2X1_127/CTRL 0.01fF
C25666 PAND2X1_220/CTRL PAND2X1_220/Y 0.00fF
C25667 POR2X1_220/B POR2X1_162/Y 0.03fF
C25668 POR2X1_68/A PAND2X1_96/CTRL 0.07fF
C25669 POR2X1_657/CTRL POR2X1_724/A 0.04fF
C25670 POR2X1_40/Y POR2X1_531/Y 0.01fF
C25671 POR2X1_686/O PAND2X1_73/Y 0.01fF
C25672 PAND2X1_862/B PAND2X1_573/CTRL2 0.01fF
C25673 PAND2X1_454/O PAND2X1_803/A 0.00fF
C25674 POR2X1_827/CTRL POR2X1_39/B 0.01fF
C25675 PAND2X1_826/O POR2X1_507/A 0.05fF
C25676 POR2X1_43/B POR2X1_497/a_16_28# 0.03fF
C25677 PAND2X1_55/Y POR2X1_285/CTRL2 0.03fF
C25678 PAND2X1_651/Y POR2X1_419/Y 0.00fF
C25679 POR2X1_57/A PAND2X1_360/CTRL2 0.03fF
C25680 PAND2X1_73/Y POR2X1_228/Y 0.03fF
C25681 POR2X1_842/CTRL2 POR2X1_456/B 0.00fF
C25682 PAND2X1_675/A PAND2X1_192/Y 0.03fF
C25683 PAND2X1_695/O PAND2X1_48/B 0.01fF
C25684 POR2X1_66/B POR2X1_532/A 0.10fF
C25685 POR2X1_68/A POR2X1_814/B 0.18fF
C25686 POR2X1_697/Y POR2X1_511/Y 0.10fF
C25687 POR2X1_555/A D_GATE_222 8.40fF
C25688 POR2X1_52/A PAND2X1_190/CTRL 0.05fF
C25689 POR2X1_43/B POR2X1_376/B 0.12fF
C25690 PAND2X1_65/B POR2X1_795/B 0.05fF
C25691 PAND2X1_56/Y PAND2X1_65/B 0.03fF
C25692 POR2X1_680/Y PAND2X1_192/a_76_28# 0.02fF
C25693 POR2X1_365/Y VDD 0.08fF
C25694 POR2X1_274/A POR2X1_574/Y 0.03fF
C25695 POR2X1_776/A POR2X1_192/B 0.05fF
C25696 POR2X1_821/Y POR2X1_40/Y 0.03fF
C25697 PAND2X1_795/B POR2X1_293/Y 0.02fF
C25698 D_INPUT_1 POR2X1_392/B 0.05fF
C25699 POR2X1_866/A POR2X1_596/a_16_28# 0.06fF
C25700 PAND2X1_20/A POR2X1_472/CTRL 0.10fF
C25701 POR2X1_811/O POR2X1_260/A 0.02fF
C25702 POR2X1_188/A POR2X1_532/A 0.05fF
C25703 POR2X1_484/CTRL2 PAND2X1_726/B 0.03fF
C25704 POR2X1_476/A POR2X1_768/O 0.02fF
C25705 POR2X1_334/B POR2X1_130/A 0.10fF
C25706 POR2X1_445/A POR2X1_703/O -0.00fF
C25707 POR2X1_78/A POR2X1_592/a_16_28# 0.01fF
C25708 PAND2X1_23/Y PAND2X1_438/CTRL2 0.01fF
C25709 POR2X1_83/B PAND2X1_374/CTRL 0.01fF
C25710 POR2X1_68/A POR2X1_325/A 0.06fF
C25711 POR2X1_861/A PAND2X1_39/B 0.17fF
C25712 PAND2X1_94/A POR2X1_650/CTRL 0.01fF
C25713 POR2X1_186/Y POR2X1_220/A 0.16fF
C25714 POR2X1_445/A POR2X1_337/Y 0.10fF
C25715 POR2X1_294/Y POR2X1_507/A 0.03fF
C25716 POR2X1_858/B POR2X1_590/A 0.04fF
C25717 POR2X1_96/A POR2X1_42/Y 20.99fF
C25718 POR2X1_48/A PAND2X1_853/B 0.03fF
C25719 POR2X1_669/A VDD 0.00fF
C25720 POR2X1_376/B POR2X1_38/B 1.08fF
C25721 PAND2X1_654/O POR2X1_46/Y 0.02fF
C25722 PAND2X1_48/B POR2X1_247/CTRL2 0.08fF
C25723 POR2X1_52/A PAND2X1_624/A 0.05fF
C25724 POR2X1_555/B POR2X1_260/A 2.40fF
C25725 PAND2X1_640/CTRL VDD 0.00fF
C25726 POR2X1_43/B PAND2X1_735/a_16_344# 0.01fF
C25727 POR2X1_252/O POR2X1_55/Y 0.01fF
C25728 PAND2X1_93/B POR2X1_737/A 0.03fF
C25729 INPUT_1 PAND2X1_721/B 0.03fF
C25730 POR2X1_567/B POR2X1_180/O 0.04fF
C25731 PAND2X1_484/O POR2X1_66/A 0.01fF
C25732 POR2X1_255/Y VDD 0.16fF
C25733 POR2X1_267/A POR2X1_773/B 0.01fF
C25734 POR2X1_286/O POR2X1_774/A 0.01fF
C25735 POR2X1_685/A POR2X1_330/Y 0.05fF
C25736 PAND2X1_254/CTRL2 POR2X1_55/Y 0.02fF
C25737 POR2X1_94/A PAND2X1_63/B 0.05fF
C25738 POR2X1_383/A POR2X1_777/B 0.07fF
C25739 PAND2X1_50/CTRL2 INPUT_6 0.00fF
C25740 POR2X1_186/Y PAND2X1_187/O -0.00fF
C25741 POR2X1_628/Y PAND2X1_508/B 0.06fF
C25742 POR2X1_558/CTRL2 POR2X1_294/B 0.13fF
C25743 POR2X1_391/A POR2X1_391/CTRL 0.00fF
C25744 PAND2X1_389/O VDD 0.00fF
C25745 PAND2X1_472/A POR2X1_13/A 0.03fF
C25746 PAND2X1_516/O POR2X1_515/Y -0.00fF
C25747 POR2X1_186/Y POR2X1_569/A 0.07fF
C25748 POR2X1_270/CTRL POR2X1_78/B 0.06fF
C25749 POR2X1_448/B PAND2X1_60/B 0.00fF
C25750 POR2X1_52/A POR2X1_43/B 0.14fF
C25751 POR2X1_612/Y POR2X1_4/Y 0.21fF
C25752 PAND2X1_798/B PAND2X1_592/Y 0.07fF
C25753 PAND2X1_642/a_16_344# POR2X1_102/Y 0.02fF
C25754 POR2X1_231/O POR2X1_795/B 0.05fF
C25755 D_INPUT_3 POR2X1_58/O 0.02fF
C25756 POR2X1_394/A POR2X1_764/a_16_28# 0.01fF
C25757 POR2X1_407/Y PAND2X1_587/Y 0.03fF
C25758 POR2X1_483/A POR2X1_702/CTRL 0.01fF
C25759 PAND2X1_651/Y PAND2X1_35/Y 0.05fF
C25760 PAND2X1_849/B POR2X1_60/Y 0.02fF
C25761 PAND2X1_555/Y VDD 0.13fF
C25762 PAND2X1_335/O POR2X1_309/Y 0.02fF
C25763 POR2X1_719/B POR2X1_719/A 0.17fF
C25764 POR2X1_220/Y PAND2X1_69/A 3.89fF
C25765 POR2X1_330/Y POR2X1_260/A 0.12fF
C25766 PAND2X1_124/Y PAND2X1_199/a_16_344# 0.02fF
C25767 PAND2X1_658/B PAND2X1_174/CTRL 0.23fF
C25768 POR2X1_750/B POR2X1_456/B 0.08fF
C25769 POR2X1_383/A PAND2X1_65/B 0.30fF
C25770 POR2X1_119/Y POR2X1_409/B 0.05fF
C25771 POR2X1_307/Y POR2X1_804/A 0.05fF
C25772 PAND2X1_131/CTRL2 PAND2X1_60/B 0.00fF
C25773 POR2X1_180/B POR2X1_814/B 0.04fF
C25774 POR2X1_441/Y PAND2X1_326/O 0.02fF
C25775 POR2X1_763/Y PAND2X1_546/O 0.08fF
C25776 POR2X1_43/B POR2X1_152/A 0.03fF
C25777 POR2X1_353/Y POR2X1_568/Y 0.05fF
C25778 PAND2X1_243/CTRL PAND2X1_35/Y 0.01fF
C25779 PAND2X1_182/CTRL2 POR2X1_55/Y 0.03fF
C25780 PAND2X1_65/B PAND2X1_253/CTRL2 0.00fF
C25781 POR2X1_296/B POR2X1_722/CTRL 0.04fF
C25782 PAND2X1_584/a_56_28# POR2X1_774/B 0.00fF
C25783 PAND2X1_69/A POR2X1_404/Y 0.03fF
C25784 POR2X1_78/A POR2X1_737/A 0.03fF
C25785 PAND2X1_493/CTRL POR2X1_60/A 0.01fF
C25786 PAND2X1_848/B POR2X1_382/CTRL 0.01fF
C25787 POR2X1_16/A PAND2X1_220/Y 0.10fF
C25788 POR2X1_537/Y POR2X1_296/B 0.05fF
C25789 POR2X1_390/B POR2X1_475/A 0.03fF
C25790 PAND2X1_491/CTRL POR2X1_294/B 0.03fF
C25791 PAND2X1_631/A POR2X1_482/O 0.05fF
C25792 POR2X1_102/Y POR2X1_533/O 0.06fF
C25793 POR2X1_236/Y POR2X1_511/a_16_28# 0.01fF
C25794 POR2X1_52/A POR2X1_38/B 0.02fF
C25795 POR2X1_165/Y POR2X1_40/Y 0.00fF
C25796 PAND2X1_6/Y POR2X1_803/A 0.02fF
C25797 INPUT_1 POR2X1_226/Y 0.03fF
C25798 POR2X1_334/B POR2X1_844/B 0.03fF
C25799 POR2X1_57/A POR2X1_821/a_16_28# 0.01fF
C25800 POR2X1_416/B POR2X1_695/O 0.15fF
C25801 POR2X1_32/A PAND2X1_199/CTRL2 0.01fF
C25802 PAND2X1_57/B PAND2X1_60/B 0.16fF
C25803 POR2X1_66/A POR2X1_199/B 0.01fF
C25804 D_GATE_222 POR2X1_775/CTRL 0.06fF
C25805 POR2X1_685/O POR2X1_687/A 0.01fF
C25806 PAND2X1_273/CTRL PAND2X1_69/A 0.01fF
C25807 POR2X1_350/Y POR2X1_35/Y 0.01fF
C25808 POR2X1_112/CTRL POR2X1_241/B 0.00fF
C25809 PAND2X1_830/Y PAND2X1_388/Y 4.09fF
C25810 POR2X1_327/Y POR2X1_405/O 0.09fF
C25811 PAND2X1_90/Y POR2X1_675/Y 0.03fF
C25812 POR2X1_205/Y PAND2X1_88/Y 0.03fF
C25813 POR2X1_96/A POR2X1_534/a_16_28# 0.03fF
C25814 PAND2X1_644/Y POR2X1_533/Y 0.05fF
C25815 POR2X1_23/Y POR2X1_39/B 4.30fF
C25816 POR2X1_116/O POR2X1_260/A 0.01fF
C25817 POR2X1_75/CTRL POR2X1_184/Y 0.00fF
C25818 PAND2X1_388/Y POR2X1_7/B 0.03fF
C25819 PAND2X1_55/Y PAND2X1_88/Y 0.03fF
C25820 POR2X1_7/A POR2X1_817/A 0.03fF
C25821 PAND2X1_480/CTRL PAND2X1_803/A 0.00fF
C25822 PAND2X1_55/Y POR2X1_84/Y 0.07fF
C25823 POR2X1_116/Y VDD 0.27fF
C25824 POR2X1_447/B POR2X1_506/B 0.01fF
C25825 PAND2X1_716/O POR2X1_52/Y 0.17fF
C25826 POR2X1_335/A PAND2X1_311/CTRL 0.01fF
C25827 POR2X1_60/A POR2X1_373/O 0.02fF
C25828 PAND2X1_852/O POR2X1_73/Y 0.04fF
C25829 POR2X1_777/B PAND2X1_71/Y 0.04fF
C25830 PAND2X1_355/O POR2X1_331/Y 0.00fF
C25831 POR2X1_283/A PAND2X1_364/CTRL2 0.01fF
C25832 PAND2X1_831/O POR2X1_300/Y 0.09fF
C25833 POR2X1_730/Y VDD 0.46fF
C25834 POR2X1_13/A PAND2X1_196/O 0.15fF
C25835 POR2X1_16/A PAND2X1_645/O 0.04fF
C25836 POR2X1_7/B PAND2X1_549/B 0.03fF
C25837 PAND2X1_90/Y POR2X1_544/B 0.10fF
C25838 PAND2X1_291/O POR2X1_198/B 0.01fF
C25839 POR2X1_65/A PAND2X1_120/O 0.01fF
C25840 PAND2X1_364/B POR2X1_385/CTRL2 0.04fF
C25841 POR2X1_71/O POR2X1_5/Y 0.18fF
C25842 POR2X1_65/O POR2X1_9/Y 0.31fF
C25843 POR2X1_809/A POR2X1_774/Y 0.16fF
C25844 POR2X1_208/A PAND2X1_23/Y 0.09fF
C25845 POR2X1_368/Y PAND2X1_785/A 0.02fF
C25846 POR2X1_170/B POR2X1_169/CTRL2 0.03fF
C25847 POR2X1_62/Y PAND2X1_340/CTRL2 0.01fF
C25848 PAND2X1_735/CTRL2 POR2X1_153/Y 0.06fF
C25849 POR2X1_7/A POR2X1_42/Y 1.34fF
C25850 PAND2X1_386/O PAND2X1_48/A 0.21fF
C25851 POR2X1_157/CTRL2 POR2X1_158/B 0.01fF
C25852 POR2X1_614/A POR2X1_210/Y 0.07fF
C25853 PAND2X1_490/CTRL POR2X1_532/A 0.01fF
C25854 POR2X1_119/Y PAND2X1_659/A 0.16fF
C25855 POR2X1_245/CTRL2 POR2X1_90/Y 0.01fF
C25856 POR2X1_334/O PAND2X1_57/B 0.01fF
C25857 POR2X1_110/CTRL2 POR2X1_5/Y 0.01fF
C25858 POR2X1_407/Y POR2X1_770/CTRL 0.01fF
C25859 PAND2X1_237/O PAND2X1_72/A 0.01fF
C25860 PAND2X1_65/B PAND2X1_71/Y 0.03fF
C25861 PAND2X1_57/B POR2X1_353/A 0.09fF
C25862 PAND2X1_651/Y PAND2X1_844/B 0.05fF
C25863 PAND2X1_862/Y PAND2X1_76/Y 0.01fF
C25864 PAND2X1_220/Y PAND2X1_336/Y 0.01fF
C25865 POR2X1_136/Y PAND2X1_469/B 0.05fF
C25866 POR2X1_32/A POR2X1_387/CTRL 0.01fF
C25867 PAND2X1_347/Y PAND2X1_360/Y 0.03fF
C25868 PAND2X1_824/B POR2X1_220/Y 0.07fF
C25869 POR2X1_516/CTRL POR2X1_283/A 0.00fF
C25870 PAND2X1_570/O PAND2X1_570/B 0.00fF
C25871 POR2X1_247/O POR2X1_260/A 0.02fF
C25872 POR2X1_360/A POR2X1_101/A 0.08fF
C25873 PAND2X1_472/O POR2X1_7/B 0.01fF
C25874 POR2X1_355/B POR2X1_352/a_16_28# 0.02fF
C25875 POR2X1_228/Y POR2X1_631/B 0.04fF
C25876 POR2X1_846/A POR2X1_20/B 1.33fF
C25877 VDD PAND2X1_2/CTRL 0.00fF
C25878 PAND2X1_7/CTRL2 POR2X1_260/A 0.03fF
C25879 PAND2X1_551/CTRL POR2X1_90/Y 0.01fF
C25880 POR2X1_614/A POR2X1_550/Y 0.00fF
C25881 POR2X1_78/B POR2X1_294/A 0.31fF
C25882 POR2X1_111/CTRL2 POR2X1_387/Y 0.02fF
C25883 POR2X1_55/Y PAND2X1_336/a_16_344# 0.01fF
C25884 PAND2X1_824/B POR2X1_404/Y 0.03fF
C25885 POR2X1_174/A POR2X1_180/Y 0.00fF
C25886 PAND2X1_193/O POR2X1_7/Y 0.03fF
C25887 POR2X1_366/A POR2X1_702/A 0.03fF
C25888 POR2X1_502/A PAND2X1_142/a_16_344# 0.02fF
C25889 POR2X1_119/Y POR2X1_272/Y 3.87fF
C25890 POR2X1_409/a_76_344# POR2X1_408/Y 0.02fF
C25891 POR2X1_740/A POR2X1_740/Y 0.02fF
C25892 POR2X1_494/a_56_344# PAND2X1_510/B 0.00fF
C25893 PAND2X1_798/Y PAND2X1_356/B 0.14fF
C25894 PAND2X1_96/B POR2X1_128/B 0.05fF
C25895 POR2X1_15/CTRL2 POR2X1_7/A 0.01fF
C25896 POR2X1_22/A POR2X1_260/A 0.10fF
C25897 POR2X1_38/B POR2X1_550/Y 0.00fF
C25898 POR2X1_143/CTRL POR2X1_62/Y 0.00fF
C25899 POR2X1_57/A PAND2X1_843/Y 0.03fF
C25900 PAND2X1_483/CTRL PAND2X1_6/A 0.03fF
C25901 POR2X1_111/CTRL POR2X1_283/A 0.08fF
C25902 POR2X1_722/Y PAND2X1_48/A 0.02fF
C25903 POR2X1_369/Y VDD 0.23fF
C25904 POR2X1_555/m4_208_n4# POR2X1_186/B 0.09fF
C25905 POR2X1_814/B POR2X1_169/A 0.10fF
C25906 POR2X1_840/O POR2X1_725/Y 0.05fF
C25907 PAND2X1_6/Y POR2X1_774/B 0.05fF
C25908 POR2X1_235/Y POR2X1_38/Y 0.03fF
C25909 POR2X1_731/O POR2X1_726/Y 0.00fF
C25910 POR2X1_523/Y POR2X1_546/CTRL 0.01fF
C25911 POR2X1_564/a_16_28# POR2X1_552/Y 0.04fF
C25912 PAND2X1_213/Y PAND2X1_738/A 0.11fF
C25913 PAND2X1_6/A POR2X1_384/m4_208_n4# 0.07fF
C25914 PAND2X1_661/B PAND2X1_196/O 0.01fF
C25915 POR2X1_116/Y PAND2X1_32/B 0.02fF
C25916 POR2X1_327/Y POR2X1_276/O 0.01fF
C25917 PAND2X1_824/B PAND2X1_93/O 0.03fF
C25918 POR2X1_228/CTRL2 POR2X1_294/B 0.03fF
C25919 POR2X1_508/B POR2X1_835/Y 0.02fF
C25920 POR2X1_447/B POR2X1_836/Y 0.01fF
C25921 POR2X1_557/A PAND2X1_69/A 0.02fF
C25922 PAND2X1_113/O PAND2X1_114/B 0.00fF
C25923 POR2X1_383/A POR2X1_712/O 0.01fF
C25924 POR2X1_42/Y POR2X1_384/Y 0.41fF
C25925 POR2X1_394/A PAND2X1_705/CTRL 0.01fF
C25926 PAND2X1_6/CTRL2 POR2X1_68/B 0.05fF
C25927 PAND2X1_20/A POR2X1_138/A 0.00fF
C25928 PAND2X1_611/CTRL2 POR2X1_54/Y 0.03fF
C25929 PAND2X1_690/CTRL PAND2X1_32/B 0.01fF
C25930 PAND2X1_90/A POR2X1_62/Y 0.13fF
C25931 POR2X1_478/B POR2X1_568/Y 0.05fF
C25932 POR2X1_791/O PAND2X1_48/A 0.02fF
C25933 PAND2X1_519/a_76_28# POR2X1_260/A 0.02fF
C25934 POR2X1_814/A POR2X1_446/B 0.01fF
C25935 PAND2X1_23/Y POR2X1_773/A 0.14fF
C25936 PAND2X1_191/O POR2X1_385/Y 0.17fF
C25937 POR2X1_776/B POR2X1_191/Y 0.05fF
C25938 PAND2X1_721/O POR2X1_77/Y 0.15fF
C25939 POR2X1_56/Y POR2X1_153/Y 0.03fF
C25940 POR2X1_327/Y PAND2X1_6/Y 0.12fF
C25941 POR2X1_186/Y PAND2X1_72/A 0.20fF
C25942 POR2X1_727/CTRL POR2X1_854/B 0.03fF
C25943 POR2X1_83/B PAND2X1_242/Y 0.05fF
C25944 VDD POR2X1_746/Y 0.01fF
C25945 PAND2X1_48/B POR2X1_726/O 0.01fF
C25946 POR2X1_329/A PAND2X1_267/Y 0.12fF
C25947 POR2X1_832/m4_208_n4# POR2X1_512/m4_208_n4# 0.13fF
C25948 POR2X1_176/O PAND2X1_566/Y 0.01fF
C25949 POR2X1_447/CTRL POR2X1_186/B 0.03fF
C25950 POR2X1_353/Y POR2X1_356/Y 0.04fF
C25951 POR2X1_481/A POR2X1_77/Y 0.51fF
C25952 POR2X1_709/B PAND2X1_69/A 0.02fF
C25953 PAND2X1_462/O VDD 0.00fF
C25954 POR2X1_307/O POR2X1_661/A 0.05fF
C25955 PAND2X1_158/CTRL2 POR2X1_156/Y 0.01fF
C25956 POR2X1_553/O POR2X1_573/A 0.02fF
C25957 POR2X1_155/CTRL POR2X1_728/A 0.00fF
C25958 POR2X1_394/A POR2X1_387/Y 0.10fF
C25959 POR2X1_81/A PAND2X1_658/B 0.30fF
C25960 POR2X1_192/B POR2X1_577/CTRL 0.01fF
C25961 POR2X1_622/B D_INPUT_0 0.01fF
C25962 PAND2X1_323/CTRL PAND2X1_32/B 0.01fF
C25963 INPUT_6 PAND2X1_2/O 0.02fF
C25964 PAND2X1_824/B POR2X1_215/A 0.04fF
C25965 POR2X1_119/Y PAND2X1_560/CTRL2 0.15fF
C25966 POR2X1_761/a_16_28# POR2X1_761/A 0.08fF
C25967 POR2X1_394/A PAND2X1_121/O 0.02fF
C25968 POR2X1_9/Y POR2X1_40/Y 0.10fF
C25969 POR2X1_216/Y POR2X1_276/Y 0.01fF
C25970 POR2X1_814/A POR2X1_121/B 0.05fF
C25971 POR2X1_260/B POR2X1_341/A 0.13fF
C25972 POR2X1_814/B PAND2X1_233/O 0.09fF
C25973 POR2X1_257/A PAND2X1_469/a_56_28# 0.00fF
C25974 POR2X1_578/Y PAND2X1_52/B 0.12fF
C25975 POR2X1_329/A PAND2X1_215/O 0.02fF
C25976 PAND2X1_22/O PAND2X1_26/A -0.00fF
C25977 POR2X1_252/Y POR2X1_7/A 0.03fF
C25978 POR2X1_93/CTRL2 POR2X1_77/Y 0.01fF
C25979 PAND2X1_99/Y PAND2X1_338/a_16_344# 0.03fF
C25980 POR2X1_158/Y PAND2X1_705/O 0.00fF
C25981 POR2X1_813/CTRL2 POR2X1_32/A 0.01fF
C25982 PAND2X1_326/B POR2X1_142/Y 0.10fF
C25983 POR2X1_193/A PAND2X1_135/O 0.03fF
C25984 PAND2X1_663/CTRL PAND2X1_659/Y 0.00fF
C25985 POR2X1_579/Y PAND2X1_135/O 0.00fF
C25986 PAND2X1_713/CTRL POR2X1_394/A 0.01fF
C25987 POR2X1_23/CTRL POR2X1_20/B 0.01fF
C25988 POR2X1_694/Y POR2X1_695/Y 0.06fF
C25989 PAND2X1_206/A POR2X1_37/Y 0.03fF
C25990 POR2X1_458/Y POR2X1_362/B 0.03fF
C25991 POR2X1_673/O POR2X1_624/B 0.09fF
C25992 POR2X1_290/Y POR2X1_234/A 0.04fF
C25993 POR2X1_651/Y PAND2X1_755/a_76_28# 0.03fF
C25994 POR2X1_160/O POR2X1_356/B 0.06fF
C25995 PAND2X1_645/B POR2X1_77/Y 0.06fF
C25996 POR2X1_602/CTRL2 POR2X1_66/A 0.01fF
C25997 PAND2X1_865/Y PAND2X1_489/CTRL 0.01fF
C25998 POR2X1_337/Y POR2X1_260/A 0.00fF
C25999 POR2X1_244/Y PAND2X1_48/A 0.03fF
C26000 POR2X1_760/A PAND2X1_361/a_76_28# 0.01fF
C26001 PAND2X1_65/B POR2X1_648/Y 1.45fF
C26002 POR2X1_23/Y POR2X1_48/A 0.56fF
C26003 PAND2X1_39/B PAND2X1_58/A 0.26fF
C26004 POR2X1_661/B POR2X1_661/A 0.07fF
C26005 POR2X1_96/O POR2X1_96/Y 0.01fF
C26006 POR2X1_614/A PAND2X1_135/O 0.05fF
C26007 PAND2X1_73/Y POR2X1_454/A 0.03fF
C26008 POR2X1_431/O POR2X1_236/Y 0.05fF
C26009 PAND2X1_341/B PAND2X1_358/A 0.07fF
C26010 POR2X1_738/A POR2X1_731/Y 0.02fF
C26011 PAND2X1_60/a_16_344# PAND2X1_58/A 0.02fF
C26012 POR2X1_67/CTRL POR2X1_83/B 0.00fF
C26013 POR2X1_417/Y PAND2X1_211/CTRL 0.01fF
C26014 POR2X1_567/A POR2X1_741/A 0.02fF
C26015 PAND2X1_618/Y PAND2X1_58/A 0.00fF
C26016 POR2X1_49/Y POR2X1_63/Y 0.15fF
C26017 POR2X1_411/B POR2X1_272/a_16_28# 0.02fF
C26018 POR2X1_65/A POR2X1_597/Y 0.00fF
C26019 POR2X1_486/O PAND2X1_57/B 0.01fF
C26020 POR2X1_650/A POR2X1_556/A 0.03fF
C26021 PAND2X1_449/CTRL2 VDD 0.00fF
C26022 POR2X1_119/Y POR2X1_150/CTRL 0.13fF
C26023 POR2X1_60/A PAND2X1_124/Y 0.03fF
C26024 POR2X1_709/A POR2X1_814/B 0.00fF
C26025 PAND2X1_496/m4_208_n4# POR2X1_573/m4_208_n4# 0.04fF
C26026 POR2X1_192/B POR2X1_191/Y 0.04fF
C26027 POR2X1_417/Y PAND2X1_212/O 0.02fF
C26028 POR2X1_329/A POR2X1_372/Y 0.07fF
C26029 POR2X1_333/Y POR2X1_568/B 0.03fF
C26030 POR2X1_635/CTRL VDD 0.00fF
C26031 PAND2X1_848/B POR2X1_9/Y 0.05fF
C26032 POR2X1_260/B POR2X1_500/A 0.03fF
C26033 POR2X1_445/A POR2X1_543/A 0.01fF
C26034 PAND2X1_75/CTRL2 POR2X1_740/Y 0.37fF
C26035 POR2X1_116/A POR2X1_116/a_16_28# -0.00fF
C26036 POR2X1_703/CTRL2 POR2X1_169/A 0.01fF
C26037 POR2X1_316/Y PAND2X1_508/Y 10.28fF
C26038 POR2X1_14/Y D_INPUT_0 0.07fF
C26039 POR2X1_774/B PAND2X1_52/B 0.43fF
C26040 POR2X1_150/Y PAND2X1_151/O 0.09fF
C26041 POR2X1_10/a_16_28# POR2X1_77/Y 0.01fF
C26042 PAND2X1_61/O POR2X1_83/B 0.07fF
C26043 POR2X1_150/Y PAND2X1_592/CTRL2 0.10fF
C26044 POR2X1_664/CTRL PAND2X1_72/A 0.01fF
C26045 PAND2X1_340/B POR2X1_5/Y 0.03fF
C26046 PAND2X1_56/Y POR2X1_814/A 0.12fF
C26047 POR2X1_188/A POR2X1_858/CTRL2 0.01fF
C26048 PAND2X1_56/Y PAND2X1_75/CTRL 0.01fF
C26049 POR2X1_634/A POR2X1_792/CTRL 0.01fF
C26050 POR2X1_760/A POR2X1_42/Y 0.03fF
C26051 POR2X1_523/Y POR2X1_67/Y 0.03fF
C26052 POR2X1_48/A POR2X1_312/Y 0.98fF
C26053 POR2X1_669/B PAND2X1_195/CTRL2 0.01fF
C26054 POR2X1_76/B POR2X1_274/B 0.02fF
C26055 POR2X1_499/A POR2X1_784/A 0.01fF
C26056 POR2X1_158/Y PAND2X1_713/O 0.00fF
C26057 PAND2X1_359/Y POR2X1_77/Y 0.03fF
C26058 PAND2X1_201/CTRL POR2X1_55/Y 0.29fF
C26059 PAND2X1_52/B POR2X1_317/B 0.03fF
C26060 PAND2X1_661/Y PAND2X1_193/Y 0.00fF
C26061 POR2X1_83/B POR2X1_60/A 4.04fF
C26062 PAND2X1_20/A PAND2X1_58/A 0.16fF
C26063 POR2X1_327/Y PAND2X1_52/B 0.05fF
C26064 POR2X1_486/CTRL PAND2X1_69/A 0.01fF
C26065 POR2X1_505/Y POR2X1_496/Y 0.02fF
C26066 PAND2X1_26/A VDD 0.36fF
C26067 PAND2X1_251/O POR2X1_362/B 0.01fF
C26068 POR2X1_287/B POR2X1_458/a_76_344# 0.00fF
C26069 POR2X1_856/B POR2X1_436/a_16_28# 0.11fF
C26070 POR2X1_220/O VDD 0.00fF
C26071 POR2X1_366/Y POR2X1_556/A 0.04fF
C26072 POR2X1_556/A POR2X1_294/B 5.19fF
C26073 POR2X1_67/Y PAND2X1_69/A 0.06fF
C26074 POR2X1_121/B POR2X1_405/CTRL2 0.00fF
C26075 PAND2X1_454/CTRL PAND2X1_446/Y 0.01fF
C26076 POR2X1_450/a_16_28# POR2X1_450/A 0.05fF
C26077 POR2X1_78/A POR2X1_302/B 0.03fF
C26078 POR2X1_274/A PAND2X1_131/O 0.01fF
C26079 POR2X1_812/a_16_28# POR2X1_452/Y 0.03fF
C26080 POR2X1_864/A PAND2X1_744/CTRL2 0.00fF
C26081 PAND2X1_612/B POR2X1_121/Y 0.03fF
C26082 POR2X1_661/CTRL2 POR2X1_661/Y 0.02fF
C26083 PAND2X1_96/CTRL PAND2X1_58/A 0.01fF
C26084 PAND2X1_55/Y POR2X1_341/A 0.14fF
C26085 PAND2X1_810/B PAND2X1_794/B 6.35fF
C26086 POR2X1_67/Y POR2X1_93/A 0.13fF
C26087 POR2X1_176/a_16_28# POR2X1_77/Y 0.01fF
C26088 PAND2X1_489/O PAND2X1_580/B 0.00fF
C26089 PAND2X1_206/A POR2X1_293/Y 0.04fF
C26090 PAND2X1_309/m4_208_n4# POR2X1_556/A 0.12fF
C26091 POR2X1_612/Y POR2X1_607/Y 0.23fF
C26092 POR2X1_833/a_16_28# POR2X1_541/B 0.11fF
C26093 PAND2X1_58/A PAND2X1_525/CTRL 0.01fF
C26094 POR2X1_814/B PAND2X1_58/A 0.07fF
C26095 PAND2X1_11/Y INPUT_7 0.03fF
C26096 INPUT_3 PAND2X1_19/CTRL2 0.03fF
C26097 POR2X1_218/Y VDD 1.41fF
C26098 POR2X1_646/Y POR2X1_480/A 0.01fF
C26099 POR2X1_35/B PAND2X1_616/O 0.04fF
C26100 POR2X1_383/A POR2X1_814/A 23.44fF
C26101 POR2X1_852/B POR2X1_630/A 0.04fF
C26102 POR2X1_102/Y POR2X1_5/Y 0.30fF
C26103 POR2X1_542/Y PAND2X1_72/A 0.04fF
C26104 PAND2X1_677/O POR2X1_718/A 0.04fF
C26105 POR2X1_718/A POR2X1_330/Y 0.05fF
C26106 PAND2X1_58/A POR2X1_325/A 0.03fF
C26107 POR2X1_383/A PAND2X1_256/CTRL2 0.06fF
C26108 PAND2X1_814/O INPUT_3 0.18fF
C26109 POR2X1_51/A POR2X1_32/A 0.02fF
C26110 POR2X1_257/A POR2X1_498/A 0.01fF
C26111 POR2X1_23/Y PAND2X1_197/Y 0.00fF
C26112 PAND2X1_96/B PAND2X1_39/B 0.07fF
C26113 POR2X1_567/B POR2X1_340/O 0.04fF
C26114 PAND2X1_69/O POR2X1_68/Y 0.00fF
C26115 PAND2X1_489/a_16_344# POR2X1_42/Y 0.02fF
C26116 POR2X1_61/Y PAND2X1_41/B 0.02fF
C26117 POR2X1_669/B POR2X1_669/CTRL2 -0.03fF
C26118 POR2X1_396/Y POR2X1_20/B 0.01fF
C26119 INPUT_3 POR2X1_376/A 0.02fF
C26120 PAND2X1_279/CTRL2 PAND2X1_57/B 0.00fF
C26121 D_INPUT_0 POR2X1_55/Y 0.13fF
C26122 POR2X1_257/A PAND2X1_284/Y 0.10fF
C26123 POR2X1_836/a_16_28# POR2X1_578/Y 0.03fF
C26124 POR2X1_65/A PAND2X1_714/A 0.16fF
C26125 POR2X1_376/B PAND2X1_474/A 0.03fF
C26126 POR2X1_60/A PAND2X1_795/B 0.05fF
C26127 PAND2X1_11/Y INPUT_4 0.03fF
C26128 PAND2X1_10/CTRL PAND2X1_55/Y 0.01fF
C26129 PAND2X1_652/Y POR2X1_32/A 0.01fF
C26130 POR2X1_815/Y D_INPUT_1 0.13fF
C26131 POR2X1_460/A PAND2X1_22/O 0.03fF
C26132 POR2X1_218/Y POR2X1_741/Y 0.07fF
C26133 POR2X1_813/a_16_28# POR2X1_38/Y 0.07fF
C26134 PAND2X1_58/A POR2X1_513/B 0.04fF
C26135 POR2X1_791/Y PAND2X1_90/Y 0.00fF
C26136 PAND2X1_48/B POR2X1_296/B 0.13fF
C26137 POR2X1_626/CTRL2 PAND2X1_6/A 0.09fF
C26138 PAND2X1_644/CTRL2 POR2X1_669/B 0.01fF
C26139 POR2X1_841/B PAND2X1_69/A 0.10fF
C26140 PAND2X1_224/CTRL POR2X1_192/B 0.28fF
C26141 POR2X1_346/O POR2X1_202/A 0.03fF
C26142 POR2X1_278/Y POR2X1_40/Y 0.12fF
C26143 POR2X1_777/B INPUT_0 7.49fF
C26144 POR2X1_502/A POR2X1_461/A 0.01fF
C26145 POR2X1_102/Y POR2X1_522/a_16_28# 0.06fF
C26146 POR2X1_130/A POR2X1_593/B 0.88fF
C26147 POR2X1_271/Y POR2X1_275/CTRL2 0.00fF
C26148 POR2X1_121/CTRL POR2X1_655/A 0.00fF
C26149 POR2X1_801/O VDD 0.00fF
C26150 PAND2X1_63/Y POR2X1_558/B 0.03fF
C26151 POR2X1_475/CTRL POR2X1_101/Y 0.01fF
C26152 PAND2X1_57/B POR2X1_750/B 0.18fF
C26153 POR2X1_149/B PAND2X1_603/CTRL 0.01fF
C26154 POR2X1_57/A PAND2X1_267/Y 0.03fF
C26155 POR2X1_710/A VDD -0.00fF
C26156 PAND2X1_97/Y POR2X1_153/Y 0.05fF
C26157 POR2X1_244/B POR2X1_186/Y 0.03fF
C26158 POR2X1_41/B PAND2X1_614/CTRL2 0.03fF
C26159 PAND2X1_755/O PAND2X1_41/B 0.05fF
C26160 POR2X1_814/A PAND2X1_71/Y 0.05fF
C26161 POR2X1_96/A POR2X1_533/A 0.00fF
C26162 POR2X1_403/O POR2X1_403/B 0.01fF
C26163 POR2X1_311/Y POR2X1_42/Y 0.09fF
C26164 PAND2X1_641/CTRL POR2X1_63/Y 0.01fF
C26165 PAND2X1_81/O POR2X1_66/A 0.07fF
C26166 PAND2X1_597/O VDD 0.00fF
C26167 POR2X1_829/A POR2X1_40/Y 0.03fF
C26168 POR2X1_66/A PAND2X1_311/CTRL2 0.01fF
C26169 POR2X1_135/Y POR2X1_45/CTRL 0.01fF
C26170 POR2X1_708/B POR2X1_602/B 0.01fF
C26171 PAND2X1_217/B POR2X1_46/Y 0.21fF
C26172 PAND2X1_474/A PAND2X1_735/a_16_344# 0.01fF
C26173 POR2X1_302/A POR2X1_121/B 0.36fF
C26174 PAND2X1_494/CTRL POR2X1_78/A 0.04fF
C26175 PAND2X1_204/CTRL VDD 0.00fF
C26176 PAND2X1_65/B INPUT_0 0.23fF
C26177 POR2X1_467/Y POR2X1_803/A 0.03fF
C26178 PAND2X1_61/Y PAND2X1_523/CTRL2 0.01fF
C26179 POR2X1_482/Y PAND2X1_254/a_16_344# 0.03fF
C26180 POR2X1_328/O POR2X1_329/A 0.01fF
C26181 POR2X1_149/B POR2X1_788/A 0.45fF
C26182 PAND2X1_682/CTRL2 POR2X1_467/Y 0.05fF
C26183 POR2X1_14/Y POR2X1_584/CTRL 0.01fF
C26184 POR2X1_624/Y PAND2X1_133/O 0.04fF
C26185 PAND2X1_722/m4_208_n4# POR2X1_591/m4_208_n4# 0.13fF
C26186 POR2X1_254/A POR2X1_341/CTRL2 0.01fF
C26187 PAND2X1_20/A PAND2X1_83/CTRL2 0.01fF
C26188 POR2X1_440/Y POR2X1_434/CTRL 0.01fF
C26189 POR2X1_502/A PAND2X1_588/O 0.10fF
C26190 POR2X1_376/B PAND2X1_350/A 0.00fF
C26191 PAND2X1_55/Y POR2X1_500/A 0.03fF
C26192 POR2X1_278/A POR2X1_37/Y 0.02fF
C26193 POR2X1_411/B PAND2X1_566/O 0.06fF
C26194 POR2X1_355/B PAND2X1_90/Y 0.06fF
C26195 PAND2X1_403/B PAND2X1_398/O 0.03fF
C26196 POR2X1_346/O POR2X1_346/A 0.02fF
C26197 PAND2X1_6/Y POR2X1_629/B 0.01fF
C26198 PAND2X1_725/Y PAND2X1_162/CTRL 0.00fF
C26199 POR2X1_29/A POR2X1_409/a_16_28# 0.03fF
C26200 PAND2X1_96/B POR2X1_805/Y 0.04fF
C26201 PAND2X1_862/B PAND2X1_659/CTRL 0.00fF
C26202 POR2X1_750/B PAND2X1_178/a_76_28# 0.02fF
C26203 POR2X1_66/B PAND2X1_697/O 0.01fF
C26204 POR2X1_16/A PAND2X1_207/CTRL2 0.01fF
C26205 PAND2X1_626/CTRL PAND2X1_69/A 0.01fF
C26206 PAND2X1_793/Y POR2X1_236/Y 0.03fF
C26207 PAND2X1_20/A PAND2X1_96/B 0.23fF
C26208 POR2X1_278/Y PAND2X1_659/B 0.07fF
C26209 POR2X1_116/A POR2X1_294/A 0.03fF
C26210 POR2X1_669/B POR2X1_387/Y 0.07fF
C26211 POR2X1_46/Y VDD 4.47fF
C26212 POR2X1_13/A PAND2X1_673/Y 0.21fF
C26213 PAND2X1_82/Y POR2X1_66/A 0.05fF
C26214 POR2X1_433/Y POR2X1_423/Y 0.06fF
C26215 PAND2X1_41/B POR2X1_35/Y 0.06fF
C26216 POR2X1_52/A PAND2X1_84/O 0.01fF
C26217 POR2X1_675/CTRL2 POR2X1_540/A 0.03fF
C26218 PAND2X1_55/Y PAND2X1_58/CTRL2 0.01fF
C26219 PAND2X1_652/A PAND2X1_192/CTRL 0.02fF
C26220 POR2X1_646/Y PAND2X1_305/O 0.05fF
C26221 POR2X1_750/B POR2X1_828/A 0.19fF
C26222 PAND2X1_638/O POR2X1_752/Y 0.05fF
C26223 INPUT_2 POR2X1_40/Y 0.03fF
C26224 POR2X1_67/A POR2X1_7/A 0.08fF
C26225 POR2X1_106/a_76_344# POR2X1_387/Y 0.02fF
C26226 PAND2X1_724/CTRL PAND2X1_169/Y 0.01fF
C26227 PAND2X1_108/CTRL2 POR2X1_814/A 0.13fF
C26228 POR2X1_102/Y PAND2X1_222/B 0.57fF
C26229 POR2X1_590/A POR2X1_550/Y 0.12fF
C26230 POR2X1_402/A PAND2X1_395/CTRL 0.01fF
C26231 POR2X1_558/B POR2X1_260/A 0.07fF
C26232 POR2X1_316/Y PAND2X1_464/B 0.75fF
C26233 INPUT_2 POR2X1_35/B 0.54fF
C26234 PAND2X1_821/CTRL2 VDD 0.00fF
C26235 PAND2X1_96/B PAND2X1_96/CTRL 0.01fF
C26236 POR2X1_558/A PAND2X1_20/A 0.03fF
C26237 POR2X1_693/Y POR2X1_697/CTRL2 0.01fF
C26238 POR2X1_507/m4_208_n4# POR2X1_854/m4_208_n4# 0.13fF
C26239 PAND2X1_623/Y VDD 0.24fF
C26240 PAND2X1_641/a_56_28# POR2X1_23/Y 0.00fF
C26241 PAND2X1_258/O POR2X1_260/A 0.01fF
C26242 POR2X1_755/O VDD 0.00fF
C26243 PAND2X1_20/CTRL2 POR2X1_68/B 0.01fF
C26244 PAND2X1_6/Y PAND2X1_423/a_16_344# 0.02fF
C26245 PAND2X1_865/Y POR2X1_411/B 0.19fF
C26246 POR2X1_814/B POR2X1_204/m4_208_n4# 0.15fF
C26247 PAND2X1_632/B POR2X1_496/Y 0.02fF
C26248 POR2X1_254/Y POR2X1_795/O 0.02fF
C26249 PAND2X1_284/CTRL VDD -0.00fF
C26250 POR2X1_62/Y PAND2X1_613/CTRL 0.00fF
C26251 INPUT_1 POR2X1_754/Y 2.75fF
C26252 POR2X1_814/B PAND2X1_96/B 0.11fF
C26253 POR2X1_109/CTRL2 POR2X1_109/Y 0.03fF
C26254 POR2X1_66/B PAND2X1_397/CTRL 0.00fF
C26255 POR2X1_88/Y PAND2X1_341/O 0.17fF
C26256 POR2X1_842/a_16_28# POR2X1_675/Y 0.02fF
C26257 POR2X1_566/A POR2X1_477/A 0.02fF
C26258 POR2X1_865/B POR2X1_860/A 0.03fF
C26259 PAND2X1_232/O POR2X1_590/A 0.15fF
C26260 PAND2X1_274/CTRL2 POR2X1_273/Y 0.01fF
C26261 PAND2X1_55/Y PAND2X1_38/O 0.01fF
C26262 POR2X1_84/O PAND2X1_57/B 0.01fF
C26263 POR2X1_68/A VDD 10.30fF
C26264 POR2X1_304/Y POR2X1_43/B 0.01fF
C26265 POR2X1_866/A PAND2X1_48/A 7.23fF
C26266 POR2X1_334/Y POR2X1_567/B 0.49fF
C26267 POR2X1_383/A POR2X1_405/CTRL2 0.12fF
C26268 POR2X1_402/B POR2X1_35/Y 0.01fF
C26269 POR2X1_480/A POR2X1_804/A 0.10fF
C26270 POR2X1_12/A POR2X1_762/a_16_28# 0.08fF
C26271 PAND2X1_725/A PAND2X1_707/CTRL 0.00fF
C26272 POR2X1_66/A PAND2X1_384/CTRL2 0.03fF
C26273 PAND2X1_779/a_16_344# PAND2X1_550/B 0.01fF
C26274 POR2X1_330/Y POR2X1_725/Y 0.10fF
C26275 PAND2X1_862/B POR2X1_43/B 0.03fF
C26276 POR2X1_343/A PAND2X1_60/B 0.02fF
C26277 POR2X1_122/Y POR2X1_822/Y 0.00fF
C26278 PAND2X1_220/Y PAND2X1_388/Y 0.00fF
C26279 POR2X1_62/Y POR2X1_23/Y 0.03fF
C26280 PAND2X1_857/B POR2X1_40/Y 0.02fF
C26281 POR2X1_62/Y POR2X1_623/CTRL 0.06fF
C26282 PAND2X1_20/A PAND2X1_503/CTRL 0.01fF
C26283 POR2X1_42/a_16_28# POR2X1_5/Y 0.01fF
C26284 PAND2X1_96/B POR2X1_325/A 0.03fF
C26285 POR2X1_66/B POR2X1_752/CTRL 0.12fF
C26286 PAND2X1_48/B POR2X1_363/CTRL2 0.01fF
C26287 PAND2X1_496/CTRL POR2X1_575/B 0.06fF
C26288 POR2X1_255/a_56_344# PAND2X1_349/A 0.00fF
C26289 POR2X1_72/B PAND2X1_717/Y 0.01fF
C26290 POR2X1_123/A PAND2X1_41/B 0.06fF
C26291 POR2X1_186/Y POR2X1_736/a_16_28# 0.00fF
C26292 POR2X1_566/A POR2X1_562/B 0.05fF
C26293 POR2X1_542/B POR2X1_284/B 0.30fF
C26294 POR2X1_439/Y POR2X1_190/a_16_28# 0.02fF
C26295 POR2X1_675/CTRL POR2X1_456/B 0.01fF
C26296 PAND2X1_376/O POR2X1_375/Y -0.00fF
C26297 PAND2X1_23/Y POR2X1_198/B 0.03fF
C26298 POR2X1_65/A PAND2X1_854/A 2.88fF
C26299 PAND2X1_738/O PAND2X1_149/A 0.04fF
C26300 POR2X1_460/A VDD 0.24fF
C26301 POR2X1_389/A POR2X1_78/B 0.03fF
C26302 PAND2X1_621/Y PAND2X1_6/A 0.04fF
C26303 PAND2X1_553/A PAND2X1_553/O -0.00fF
C26304 PAND2X1_73/Y POR2X1_579/B 0.00fF
C26305 PAND2X1_572/CTRL2 INPUT_0 0.01fF
C26306 POR2X1_685/A PAND2X1_679/O 0.01fF
C26307 PAND2X1_23/Y D_GATE_741 0.18fF
C26308 PAND2X1_243/O PAND2X1_734/B 0.02fF
C26309 PAND2X1_421/CTRL2 PAND2X1_69/A 0.01fF
C26310 POR2X1_186/Y PAND2X1_172/a_16_344# 0.06fF
C26311 D_GATE_741 PAND2X1_504/CTRL2 0.02fF
C26312 PAND2X1_424/O PAND2X1_57/B -0.00fF
C26313 POR2X1_472/CTRL VDD 0.00fF
C26314 POR2X1_327/Y POR2X1_467/Y 0.14fF
C26315 POR2X1_68/A POR2X1_741/Y 0.08fF
C26316 PAND2X1_73/Y POR2X1_571/Y 0.05fF
C26317 POR2X1_259/B POR2X1_750/B 0.05fF
C26318 PAND2X1_460/O PAND2X1_472/B 0.02fF
C26319 PAND2X1_625/a_76_28# POR2X1_740/Y 0.05fF
C26320 PAND2X1_90/A PAND2X1_316/a_76_28# 0.01fF
C26321 PAND2X1_724/B POR2X1_90/Y 0.03fF
C26322 POR2X1_507/a_16_28# POR2X1_355/A 0.02fF
C26323 POR2X1_227/B POR2X1_568/A 0.07fF
C26324 POR2X1_335/A PAND2X1_6/Y 0.03fF
C26325 PAND2X1_188/O POR2X1_498/A 0.01fF
C26326 POR2X1_180/B VDD 0.02fF
C26327 PAND2X1_41/B POR2X1_227/CTRL2 0.01fF
C26328 POR2X1_38/Y POR2X1_42/Y 10.88fF
C26329 POR2X1_82/CTRL POR2X1_16/A 0.00fF
C26330 POR2X1_447/B POR2X1_836/A 0.01fF
C26331 POR2X1_508/B POR2X1_836/B 0.00fF
C26332 POR2X1_514/Y POR2X1_840/B 0.05fF
C26333 POR2X1_540/A POR2X1_732/B 0.07fF
C26334 POR2X1_96/A PAND2X1_728/CTRL2 0.01fF
C26335 PAND2X1_556/B POR2X1_310/Y 0.06fF
C26336 POR2X1_114/B PAND2X1_69/A 0.10fF
C26337 POR2X1_356/A POR2X1_338/CTRL 0.26fF
C26338 POR2X1_68/A PAND2X1_32/B 0.26fF
C26339 POR2X1_356/A PAND2X1_824/O 0.05fF
C26340 PAND2X1_632/O INPUT_0 0.05fF
C26341 POR2X1_96/A PAND2X1_550/B 0.15fF
C26342 PAND2X1_744/O POR2X1_644/A 0.05fF
C26343 POR2X1_150/Y PAND2X1_860/A 0.03fF
C26344 POR2X1_94/A POR2X1_294/A 0.03fF
C26345 POR2X1_170/B POR2X1_568/Y 0.03fF
C26346 POR2X1_242/O POR2X1_192/B 0.02fF
C26347 POR2X1_57/A POR2X1_757/A 0.01fF
C26348 PAND2X1_219/a_16_344# POR2X1_591/Y 0.01fF
C26349 POR2X1_696/Y POR2X1_394/A 0.01fF
C26350 PAND2X1_216/B PAND2X1_571/Y 0.02fF
C26351 POR2X1_391/B VDD 0.04fF
C26352 POR2X1_57/A POR2X1_519/Y 1.72fF
C26353 POR2X1_294/B POR2X1_702/O 0.01fF
C26354 POR2X1_575/B POR2X1_575/CTRL 0.03fF
C26355 PAND2X1_810/B PAND2X1_221/Y 4.66fF
C26356 PAND2X1_723/A PAND2X1_364/B 0.04fF
C26357 INPUT_0 POR2X1_385/a_76_344# 0.00fF
C26358 PAND2X1_859/B POR2X1_283/A 0.03fF
C26359 POR2X1_383/A POR2X1_260/Y 0.04fF
C26360 POR2X1_228/Y POR2X1_715/a_16_28# 0.10fF
C26361 PAND2X1_600/CTRL PAND2X1_72/A 0.01fF
C26362 PAND2X1_90/Y POR2X1_209/O 0.02fF
C26363 POR2X1_174/A POR2X1_568/B 11.02fF
C26364 POR2X1_596/A PAND2X1_743/CTRL2 0.01fF
C26365 D_INPUT_0 POR2X1_500/CTRL2 0.01fF
C26366 POR2X1_63/CTRL2 POR2X1_7/A 0.03fF
C26367 PAND2X1_388/Y PAND2X1_370/CTRL2 0.01fF
C26368 POR2X1_855/B PAND2X1_599/CTRL 0.01fF
C26369 POR2X1_814/A POR2X1_648/Y 0.05fF
C26370 INPUT_1 POR2X1_817/A 0.05fF
C26371 POR2X1_301/CTRL PAND2X1_60/B 0.09fF
C26372 POR2X1_68/A PAND2X1_312/O 0.04fF
C26373 PAND2X1_23/Y POR2X1_507/CTRL2 0.01fF
C26374 D_INPUT_1 POR2X1_550/O 0.01fF
C26375 POR2X1_458/B PAND2X1_69/A 0.05fF
C26376 POR2X1_78/B POR2X1_334/Y 0.10fF
C26377 POR2X1_488/Y PAND2X1_363/O 0.03fF
C26378 POR2X1_302/A POR2X1_383/A 0.47fF
C26379 POR2X1_460/A PAND2X1_32/B 0.06fF
C26380 PAND2X1_206/a_16_344# POR2X1_153/Y 0.05fF
C26381 POR2X1_775/A POR2X1_854/B 0.05fF
C26382 POR2X1_5/Y POR2X1_5/O 0.00fF
C26383 POR2X1_596/A POR2X1_770/O 0.01fF
C26384 PAND2X1_716/CTRL PAND2X1_656/A 0.01fF
C26385 POR2X1_362/B POR2X1_362/CTRL2 0.01fF
C26386 PAND2X1_55/Y POR2X1_151/CTRL 0.01fF
C26387 POR2X1_16/A PAND2X1_776/CTRL 0.01fF
C26388 POR2X1_390/B POR2X1_740/Y 0.03fF
C26389 PAND2X1_48/B POR2X1_543/CTRL 0.01fF
C26390 INPUT_1 POR2X1_42/Y 0.15fF
C26391 PAND2X1_329/CTRL PAND2X1_69/A 0.01fF
C26392 PAND2X1_802/B POR2X1_42/Y 0.01fF
C26393 POR2X1_164/Y PAND2X1_565/CTRL2 0.01fF
C26394 PAND2X1_649/A POR2X1_689/CTRL2 0.01fF
C26395 PAND2X1_841/B POR2X1_271/A 1.26fF
C26396 POR2X1_131/O PAND2X1_349/A 0.01fF
C26397 POR2X1_163/A POR2X1_394/A 0.21fF
C26398 POR2X1_8/Y PAND2X1_341/O 0.07fF
C26399 POR2X1_68/A POR2X1_543/CTRL2 0.01fF
C26400 POR2X1_167/CTRL POR2X1_73/Y 0.07fF
C26401 POR2X1_780/B POR2X1_532/A 0.03fF
C26402 POR2X1_41/B POR2X1_595/CTRL2 0.04fF
C26403 POR2X1_137/Y PAND2X1_60/B 0.05fF
C26404 POR2X1_68/A POR2X1_673/Y 0.06fF
C26405 PAND2X1_117/CTRL POR2X1_557/B 0.00fF
C26406 POR2X1_486/B POR2X1_287/B 0.01fF
C26407 POR2X1_42/Y POR2X1_153/Y 0.02fF
C26408 PAND2X1_714/A PAND2X1_169/O 0.31fF
C26409 POR2X1_366/a_76_344# PAND2X1_6/Y 0.03fF
C26410 POR2X1_383/A POR2X1_493/O 0.01fF
C26411 PAND2X1_480/O POR2X1_43/B 0.01fF
C26412 PAND2X1_652/A PAND2X1_853/B 0.03fF
C26413 POR2X1_553/A POR2X1_724/A 0.11fF
C26414 VDD PAND2X1_517/O 0.00fF
C26415 PAND2X1_94/A PAND2X1_79/Y 0.06fF
C26416 POR2X1_391/B PAND2X1_32/B 0.02fF
C26417 PAND2X1_48/B POR2X1_342/CTRL 0.01fF
C26418 POR2X1_528/Y POR2X1_408/Y 0.19fF
C26419 VDD POR2X1_181/O 0.00fF
C26420 POR2X1_164/Y POR2X1_91/Y 0.01fF
C26421 PAND2X1_26/CTRL POR2X1_260/A 0.01fF
C26422 PAND2X1_55/Y POR2X1_735/O 0.00fF
C26423 POR2X1_20/O POR2X1_4/Y 0.05fF
C26424 VDD POR2X1_169/A 0.37fF
C26425 POR2X1_52/A PAND2X1_865/Y 0.07fF
C26426 PAND2X1_284/a_76_28# POR2X1_394/A 0.02fF
C26427 PAND2X1_551/O PAND2X1_569/B 0.00fF
C26428 POR2X1_20/B POR2X1_271/B 0.03fF
C26429 POR2X1_456/B POR2X1_318/A 0.11fF
C26430 INPUT_6 PAND2X1_157/CTRL2 0.01fF
C26431 INPUT_0 POR2X1_372/CTRL 0.01fF
C26432 POR2X1_43/B PAND2X1_716/B 0.03fF
C26433 PAND2X1_200/B POR2X1_73/Y 0.03fF
C26434 POR2X1_121/A POR2X1_537/Y 0.00fF
C26435 POR2X1_438/O POR2X1_373/Y 0.18fF
C26436 POR2X1_38/B POR2X1_673/B 0.01fF
C26437 PAND2X1_612/a_76_28# POR2X1_472/B 0.01fF
C26438 POR2X1_833/A PAND2X1_60/B 0.10fF
C26439 POR2X1_793/CTRL PAND2X1_52/B 0.01fF
C26440 POR2X1_538/A POR2X1_260/A 0.01fF
C26441 POR2X1_332/Y PAND2X1_96/B 0.15fF
C26442 D_INPUT_3 POR2X1_394/A 0.07fF
C26443 POR2X1_809/A POR2X1_685/B 0.01fF
C26444 POR2X1_290/Y POR2X1_39/B 0.09fF
C26445 POR2X1_57/A PAND2X1_325/CTRL2 0.01fF
C26446 POR2X1_730/Y POR2X1_687/A 0.02fF
C26447 POR2X1_760/A PAND2X1_576/B 0.10fF
C26448 PAND2X1_187/a_16_344# POR2X1_444/Y 0.02fF
C26449 PAND2X1_659/Y POR2X1_7/m4_208_n4# 0.12fF
C26450 POR2X1_99/B POR2X1_631/B 0.03fF
C26451 POR2X1_245/Y POR2X1_129/Y 0.10fF
C26452 POR2X1_389/A POR2X1_294/A 0.07fF
C26453 PAND2X1_69/A PAND2X1_122/CTRL2 0.01fF
C26454 POR2X1_383/A POR2X1_151/Y 0.01fF
C26455 VDD POR2X1_138/A -0.00fF
C26456 PAND2X1_60/B PAND2X1_18/B 0.01fF
C26457 POR2X1_88/a_16_28# POR2X1_88/A 0.03fF
C26458 POR2X1_564/Y POR2X1_181/Y 0.02fF
C26459 PAND2X1_634/CTRL POR2X1_48/A 0.01fF
C26460 POR2X1_416/B PAND2X1_375/O 0.01fF
C26461 POR2X1_571/a_16_28# POR2X1_569/A 0.07fF
C26462 POR2X1_509/CTRL POR2X1_857/B 0.09fF
C26463 PAND2X1_658/B POR2X1_39/B 0.03fF
C26464 PAND2X1_267/B PAND2X1_267/O 0.00fF
C26465 PAND2X1_350/m4_208_n4# POR2X1_394/A 0.06fF
C26466 PAND2X1_175/O PAND2X1_853/B 0.08fF
C26467 POR2X1_112/CTRL2 POR2X1_510/Y 0.03fF
C26468 PAND2X1_73/Y PAND2X1_79/a_76_28# 0.04fF
C26469 POR2X1_616/Y POR2X1_7/A 0.06fF
C26470 POR2X1_43/a_76_344# POR2X1_43/B 0.01fF
C26471 POR2X1_416/B POR2X1_693/Y 0.03fF
C26472 POR2X1_609/Y POR2X1_20/B 0.06fF
C26473 POR2X1_854/CTRL POR2X1_567/B 0.03fF
C26474 POR2X1_698/Y VDD -0.00fF
C26475 POR2X1_499/a_56_344# POR2X1_341/A 0.01fF
C26476 POR2X1_52/A POR2X1_90/CTRL 0.00fF
C26477 POR2X1_416/B POR2X1_765/a_56_344# 0.00fF
C26478 POR2X1_9/Y POR2X1_5/Y 1.10fF
C26479 PAND2X1_797/Y PAND2X1_149/A 0.00fF
C26480 PAND2X1_639/Y POR2X1_588/Y 0.02fF
C26481 POR2X1_567/A POR2X1_566/B 0.45fF
C26482 POR2X1_287/B POR2X1_486/CTRL2 0.01fF
C26483 PAND2X1_498/a_76_28# PAND2X1_72/A 0.01fF
C26484 POR2X1_8/Y POR2X1_153/a_16_28# 0.02fF
C26485 POR2X1_711/B POR2X1_463/Y 0.10fF
C26486 POR2X1_14/Y PAND2X1_33/O 0.17fF
C26487 POR2X1_257/A POR2X1_432/CTRL 0.02fF
C26488 POR2X1_826/a_16_28# PAND2X1_734/B 0.03fF
C26489 POR2X1_703/A POR2X1_703/a_76_344# 0.03fF
C26490 PAND2X1_39/B POR2X1_608/Y 0.02fF
C26491 POR2X1_52/A POR2X1_91/O 0.01fF
C26492 POR2X1_865/CTRL2 PAND2X1_52/B 0.01fF
C26493 INPUT_1 POR2X1_252/Y 0.03fF
C26494 POR2X1_316/Y POR2X1_283/A 0.03fF
C26495 PAND2X1_39/B POR2X1_400/B 0.01fF
C26496 PAND2X1_798/Y POR2X1_283/A 0.03fF
C26497 PAND2X1_601/CTRL2 POR2X1_296/B 0.03fF
C26498 PAND2X1_39/B POR2X1_806/CTRL2 0.03fF
C26499 PAND2X1_862/O PAND2X1_858/Y 0.03fF
C26500 POR2X1_411/B POR2X1_609/CTRL 0.01fF
C26501 PAND2X1_639/Y POR2X1_583/Y 0.37fF
C26502 POR2X1_673/Y PAND2X1_517/O 0.03fF
C26503 POR2X1_260/B POR2X1_29/A 0.03fF
C26504 POR2X1_266/A POR2X1_62/Y 0.18fF
C26505 POR2X1_138/A PAND2X1_32/B 0.07fF
C26506 POR2X1_60/A PAND2X1_206/A 0.09fF
C26507 POR2X1_814/A INPUT_0 0.19fF
C26508 POR2X1_859/O PAND2X1_41/B 0.09fF
C26509 POR2X1_99/A PAND2X1_39/B 0.03fF
C26510 POR2X1_421/a_16_28# POR2X1_329/A 0.06fF
C26511 POR2X1_49/Y POR2X1_415/A 0.07fF
C26512 POR2X1_817/a_16_28# POR2X1_32/A 0.02fF
C26513 POR2X1_704/Y POR2X1_568/B 0.55fF
C26514 POR2X1_647/B POR2X1_862/B 0.00fF
C26515 POR2X1_153/Y PAND2X1_860/a_56_28# 0.00fF
C26516 POR2X1_130/CTRL POR2X1_343/Y -0.00fF
C26517 POR2X1_482/CTRL2 POR2X1_60/A 0.01fF
C26518 POR2X1_249/Y PAND2X1_52/B 0.03fF
C26519 PAND2X1_48/B PAND2X1_85/O 0.01fF
C26520 POR2X1_667/A POR2X1_37/Y 0.05fF
C26521 PAND2X1_336/Y PAND2X1_352/B 0.01fF
C26522 POR2X1_607/A POR2X1_37/Y 0.03fF
C26523 POR2X1_608/Y POR2X1_805/Y 0.18fF
C26524 PAND2X1_73/Y PAND2X1_531/O 0.13fF
C26525 PAND2X1_217/B PAND2X1_571/A 0.05fF
C26526 PAND2X1_472/B PAND2X1_33/O 0.06fF
C26527 POR2X1_709/A VDD 0.46fF
C26528 PAND2X1_20/A POR2X1_608/Y 0.01fF
C26529 POR2X1_411/a_56_344# POR2X1_411/A 0.00fF
C26530 POR2X1_329/A PAND2X1_339/Y 0.68fF
C26531 POR2X1_65/A POR2X1_93/Y 0.01fF
C26532 POR2X1_52/A POR2X1_816/CTRL 0.01fF
C26533 POR2X1_730/Y POR2X1_568/A 0.03fF
C26534 POR2X1_257/A PAND2X1_707/CTRL2 0.00fF
C26535 POR2X1_41/B PAND2X1_247/CTRL2 0.03fF
C26536 POR2X1_66/B POR2X1_586/Y 0.03fF
C26537 POR2X1_658/O POR2X1_193/A 0.03fF
C26538 PAND2X1_9/Y POR2X1_46/Y 0.01fF
C26539 D_INPUT_5 POR2X1_25/a_76_344# 0.01fF
C26540 POR2X1_460/Y POR2X1_459/A 0.00fF
C26541 PAND2X1_205/a_76_28# PAND2X1_473/B 0.02fF
C26542 POR2X1_491/CTRL POR2X1_102/Y 0.01fF
C26543 POR2X1_854/O POR2X1_776/B 0.01fF
C26544 POR2X1_260/B POR2X1_546/A 0.07fF
C26545 POR2X1_20/B PAND2X1_546/Y 0.03fF
C26546 POR2X1_814/B POR2X1_608/Y 0.01fF
C26547 POR2X1_140/B POR2X1_556/A 0.03fF
C26548 PAND2X1_75/O POR2X1_532/A 0.04fF
C26549 POR2X1_41/B PAND2X1_404/Y 0.03fF
C26550 POR2X1_696/Y POR2X1_669/B 0.02fF
C26551 GATE_479 POR2X1_83/B 0.03fF
C26552 POR2X1_633/CTRL2 POR2X1_68/B 0.02fF
C26553 POR2X1_68/A PAND2X1_9/Y 0.03fF
C26554 PAND2X1_169/Y POR2X1_40/Y 0.96fF
C26555 POR2X1_285/CTRL POR2X1_590/A 0.01fF
C26556 PAND2X1_787/A PAND2X1_464/B 0.01fF
C26557 POR2X1_78/A POR2X1_362/B 0.10fF
C26558 POR2X1_257/A PAND2X1_725/A 0.00fF
C26559 POR2X1_841/CTRL POR2X1_804/A 0.07fF
C26560 PAND2X1_248/O POR2X1_404/Y 0.03fF
C26561 PAND2X1_669/CTRL POR2X1_668/Y 0.01fF
C26562 POR2X1_730/Y POR2X1_440/a_16_28# 0.02fF
C26563 POR2X1_95/a_16_28# POR2X1_416/B 0.01fF
C26564 POR2X1_411/Y POR2X1_612/Y 0.09fF
C26565 POR2X1_57/A POR2X1_485/Y 0.00fF
C26566 POR2X1_856/B POR2X1_855/Y 0.01fF
C26567 POR2X1_102/Y PAND2X1_723/Y 0.01fF
C26568 POR2X1_48/A POR2X1_290/Y 0.03fF
C26569 PAND2X1_673/Y POR2X1_29/A 0.03fF
C26570 POR2X1_40/Y POR2X1_743/CTRL 0.08fF
C26571 PAND2X1_65/B PAND2X1_766/CTRL2 0.01fF
C26572 POR2X1_3/A POR2X1_20/B 0.03fF
C26573 POR2X1_260/B POR2X1_805/A 0.03fF
C26574 POR2X1_454/A POR2X1_35/Y 0.02fF
C26575 PAND2X1_58/A VDD 4.80fF
C26576 POR2X1_614/A POR2X1_445/A 0.09fF
C26577 PAND2X1_73/Y POR2X1_608/a_16_28# 0.04fF
C26578 POR2X1_78/A POR2X1_608/a_76_344# 0.00fF
C26579 POR2X1_43/B POR2X1_490/Y 0.05fF
C26580 PAND2X1_827/CTRL2 POR2X1_741/Y 0.06fF
C26581 PAND2X1_827/O POR2X1_740/Y 0.02fF
C26582 POR2X1_102/Y PAND2X1_778/a_56_28# 0.00fF
C26583 POR2X1_480/A POR2X1_794/B 0.07fF
C26584 POR2X1_23/Y PAND2X1_652/A 1.22fF
C26585 PAND2X1_270/O POR2X1_20/B 0.02fF
C26586 PAND2X1_360/CTRL VDD 0.00fF
C26587 POR2X1_67/Y PAND2X1_789/CTRL2 0.01fF
C26588 POR2X1_41/B POR2X1_309/O 0.01fF
C26589 POR2X1_812/B POR2X1_452/Y 0.02fF
C26590 PAND2X1_402/CTRL2 POR2X1_236/Y 0.01fF
C26591 POR2X1_49/Y POR2X1_743/O 0.12fF
C26592 POR2X1_48/A PAND2X1_658/B 0.03fF
C26593 POR2X1_411/B PAND2X1_383/O 0.04fF
C26594 POR2X1_614/A POR2X1_809/CTRL 0.01fF
C26595 PAND2X1_20/A POR2X1_128/CTRL 0.01fF
C26596 PAND2X1_683/a_56_28# POR2X1_78/B 0.00fF
C26597 POR2X1_644/CTRL POR2X1_644/A 0.06fF
C26598 PAND2X1_691/Y PAND2X1_644/m4_208_n4# 0.12fF
C26599 POR2X1_629/CTRL PAND2X1_69/A 0.01fF
C26600 PAND2X1_627/CTRL2 POR2X1_852/B 0.06fF
C26601 POR2X1_240/O PAND2X1_88/Y 0.01fF
C26602 POR2X1_63/Y POR2X1_235/O 0.01fF
C26603 POR2X1_127/a_16_28# POR2X1_7/B 0.01fF
C26604 POR2X1_110/Y PAND2X1_458/CTRL 0.01fF
C26605 POR2X1_296/B POR2X1_717/Y 0.03fF
C26606 POR2X1_38/CTRL POR2X1_38/B 0.01fF
C26607 POR2X1_411/B PAND2X1_348/CTRL2 0.01fF
C26608 PAND2X1_73/Y POR2X1_664/Y 0.52fF
C26609 POR2X1_260/B POR2X1_500/Y 0.03fF
C26610 POR2X1_40/Y POR2X1_393/a_56_344# 0.01fF
C26611 POR2X1_460/Y PAND2X1_376/CTRL 0.01fF
C26612 POR2X1_133/O POR2X1_40/Y 0.01fF
C26613 PAND2X1_139/B PAND2X1_139/O 0.00fF
C26614 PAND2X1_798/B POR2X1_487/O 0.03fF
C26615 PAND2X1_48/B PAND2X1_15/a_16_344# 0.01fF
C26616 POR2X1_686/B POR2X1_686/A 0.00fF
C26617 D_INPUT_0 POR2X1_513/Y 0.03fF
C26618 PAND2X1_6/Y POR2X1_34/B 0.08fF
C26619 POR2X1_60/A POR2X1_697/Y 0.02fF
C26620 PAND2X1_425/Y POR2X1_260/A 0.04fF
C26621 POR2X1_33/A POR2X1_68/B 0.00fF
C26622 PAND2X1_862/B PAND2X1_474/A 0.03fF
C26623 PAND2X1_254/Y POR2X1_423/Y 0.03fF
C26624 POR2X1_502/A PAND2X1_387/CTRL 0.05fF
C26625 POR2X1_76/O POR2X1_569/A 0.04fF
C26626 POR2X1_287/a_16_28# POR2X1_733/A 0.08fF
C26627 POR2X1_23/Y POR2X1_152/Y 0.03fF
C26628 PAND2X1_58/A POR2X1_741/Y 0.03fF
C26629 POR2X1_94/CTRL POR2X1_14/Y 0.01fF
C26630 PAND2X1_790/a_16_344# POR2X1_7/A 0.01fF
C26631 POR2X1_566/A PAND2X1_229/O 0.03fF
C26632 PAND2X1_787/Y VDD 2.02fF
C26633 POR2X1_466/A POR2X1_540/A 0.05fF
C26634 POR2X1_76/A POR2X1_274/B 0.00fF
C26635 PAND2X1_794/CTRL PAND2X1_794/B 0.01fF
C26636 POR2X1_368/O POR2X1_5/Y 0.02fF
C26637 POR2X1_828/Y POR2X1_220/Y 0.03fF
C26638 POR2X1_496/Y POR2X1_90/Y 0.07fF
C26639 POR2X1_49/Y POR2X1_56/B 0.13fF
C26640 POR2X1_548/O PAND2X1_8/Y 0.18fF
C26641 POR2X1_278/Y POR2X1_5/Y 2.06fF
C26642 POR2X1_602/B PAND2X1_55/Y 0.03fF
C26643 POR2X1_457/B VDD 0.15fF
C26644 PAND2X1_736/Y POR2X1_72/B 0.01fF
C26645 PAND2X1_73/Y POR2X1_112/Y 0.05fF
C26646 POR2X1_473/a_56_344# POR2X1_276/Y 0.00fF
C26647 POR2X1_814/B POR2X1_791/CTRL2 0.01fF
C26648 POR2X1_60/A PAND2X1_357/Y 0.08fF
C26649 PAND2X1_667/O VDD 0.00fF
C26650 PAND2X1_48/B POR2X1_186/Y 4.70fF
C26651 D_INPUT_1 POR2X1_390/CTRL 0.04fF
C26652 POR2X1_130/CTRL POR2X1_624/Y 0.03fF
C26653 POR2X1_23/Y POR2X1_437/CTRL2 0.03fF
C26654 POR2X1_67/A POR2X1_38/Y 0.16fF
C26655 POR2X1_673/CTRL PAND2X1_6/A 0.04fF
C26656 POR2X1_315/Y PAND2X1_776/Y 0.18fF
C26657 PAND2X1_6/Y PAND2X1_230/a_16_344# 0.02fF
C26658 POR2X1_635/Y VDD 0.20fF
C26659 POR2X1_66/A POR2X1_548/A 0.00fF
C26660 PAND2X1_659/A PAND2X1_575/A 0.06fF
C26661 PAND2X1_58/A PAND2X1_32/B 0.79fF
C26662 POR2X1_435/Y VDD -0.00fF
C26663 POR2X1_37/Y POR2X1_245/Y 0.16fF
C26664 POR2X1_496/a_16_28# POR2X1_789/B 0.03fF
C26665 POR2X1_376/B POR2X1_494/Y 0.03fF
C26666 POR2X1_66/A POR2X1_550/Y 0.03fF
C26667 D_INPUT_3 POR2X1_669/B 0.05fF
C26668 PAND2X1_499/a_16_344# POR2X1_293/Y 0.01fF
C26669 POR2X1_482/O POR2X1_7/A 0.19fF
C26670 POR2X1_634/A PAND2X1_47/CTRL 0.17fF
C26671 PAND2X1_239/O POR2X1_566/B 0.04fF
C26672 POR2X1_514/a_16_28# PAND2X1_20/A 0.03fF
C26673 POR2X1_865/B POR2X1_121/B 0.02fF
C26674 POR2X1_102/Y PAND2X1_572/CTRL2 0.09fF
C26675 POR2X1_832/B POR2X1_830/A 0.02fF
C26676 POR2X1_72/B POR2X1_56/Y 0.03fF
C26677 PAND2X1_668/CTRL VDD 0.00fF
C26678 POR2X1_760/O POR2X1_7/B 0.02fF
C26679 PAND2X1_117/CTRL2 VDD 0.00fF
C26680 POR2X1_25/Y POR2X1_20/B 0.21fF
C26681 POR2X1_483/O POR2X1_483/B 0.04fF
C26682 POR2X1_625/m4_208_n4# POR2X1_7/B 0.07fF
C26683 POR2X1_293/Y POR2X1_372/O 0.13fF
C26684 POR2X1_96/A PAND2X1_734/B 0.08fF
C26685 POR2X1_83/B POR2X1_142/Y 0.03fF
C26686 POR2X1_614/Y POR2X1_7/A 0.02fF
C26687 POR2X1_347/B PAND2X1_57/B 0.01fF
C26688 POR2X1_96/Y PAND2X1_201/CTRL 0.03fF
C26689 POR2X1_814/A PAND2X1_122/a_76_28# 0.01fF
C26690 POR2X1_49/Y PAND2X1_724/CTRL2 0.03fF
C26691 PAND2X1_232/O POR2X1_66/A 0.01fF
C26692 PAND2X1_267/B POR2X1_7/Y 0.01fF
C26693 PAND2X1_377/Y VDD 0.13fF
C26694 POR2X1_370/Y POR2X1_740/Y 0.03fF
C26695 POR2X1_16/A POR2X1_487/CTRL2 0.02fF
C26696 PAND2X1_57/B POR2X1_756/CTRL2 0.01fF
C26697 PAND2X1_750/CTRL POR2X1_749/Y 0.00fF
C26698 POR2X1_411/B PAND2X1_352/Y 0.03fF
C26699 POR2X1_612/CTRL POR2X1_4/Y 0.01fF
C26700 POR2X1_745/CTRL2 VDD -0.00fF
C26701 POR2X1_79/Y PAND2X1_592/Y 0.03fF
C26702 PAND2X1_796/B PAND2X1_506/Y 0.02fF
C26703 POR2X1_334/A PAND2X1_93/B 0.01fF
C26704 POR2X1_98/O POR2X1_260/A 0.06fF
C26705 PAND2X1_205/A PAND2X1_853/B 0.03fF
C26706 POR2X1_92/CTRL POR2X1_49/Y 0.00fF
C26707 POR2X1_45/Y PAND2X1_579/B 8.95fF
C26708 POR2X1_406/Y PAND2X1_716/CTRL2 0.01fF
C26709 D_GATE_662 POR2X1_544/A 0.02fF
C26710 INPUT_2 POR2X1_5/Y 0.03fF
C26711 INPUT_1 POR2X1_67/A 0.07fF
C26712 POR2X1_631/A PAND2X1_41/B 0.03fF
C26713 PAND2X1_94/A PAND2X1_77/CTRL 0.01fF
C26714 POR2X1_614/A POR2X1_786/O 0.05fF
C26715 PAND2X1_140/A PAND2X1_554/a_16_344# 0.03fF
C26716 POR2X1_52/A POR2X1_494/Y 0.00fF
C26717 POR2X1_782/A VDD 0.00fF
C26718 POR2X1_334/B POR2X1_124/CTRL 0.25fF
C26719 POR2X1_270/Y POR2X1_370/CTRL 0.03fF
C26720 POR2X1_770/CTRL2 POR2X1_770/A 0.01fF
C26721 POR2X1_20/A POR2X1_4/Y 0.04fF
C26722 PAND2X1_309/CTRL2 POR2X1_741/Y 0.00fF
C26723 PAND2X1_309/CTRL POR2X1_740/Y 0.00fF
C26724 D_INPUT_0 POR2X1_129/Y 0.03fF
C26725 POR2X1_94/CTRL PAND2X1_472/B 0.06fF
C26726 POR2X1_383/A PAND2X1_428/a_16_344# 0.01fF
C26727 POR2X1_413/A POR2X1_290/Y 0.04fF
C26728 POR2X1_355/B D_GATE_222 0.07fF
C26729 POR2X1_567/B POR2X1_726/CTRL2 0.52fF
C26730 POR2X1_673/Y PAND2X1_58/A 0.03fF
C26731 POR2X1_65/A PAND2X1_650/O 0.07fF
C26732 POR2X1_38/Y PAND2X1_733/Y 0.15fF
C26733 POR2X1_853/O POR2X1_795/B 0.01fF
C26734 POR2X1_650/A PAND2X1_60/B 0.03fF
C26735 POR2X1_66/A POR2X1_195/CTRL 0.01fF
C26736 PAND2X1_96/B VDD 2.42fF
C26737 POR2X1_231/B POR2X1_795/B 0.03fF
C26738 POR2X1_131/CTRL POR2X1_13/A 0.01fF
C26739 PAND2X1_738/Y PAND2X1_388/CTRL2 0.15fF
C26740 POR2X1_360/A POR2X1_35/Y 0.11fF
C26741 PAND2X1_56/Y PAND2X1_309/O 0.07fF
C26742 PAND2X1_247/CTRL2 POR2X1_77/Y 0.01fF
C26743 PAND2X1_844/a_76_28# D_INPUT_0 0.04fF
C26744 PAND2X1_435/Y POR2X1_129/Y 0.02fF
C26745 PAND2X1_131/CTRL2 POR2X1_318/A 0.03fF
C26746 POR2X1_16/A POR2X1_40/Y 2.70fF
C26747 POR2X1_68/A POR2X1_149/Y 0.18fF
C26748 POR2X1_271/A POR2X1_516/Y 0.06fF
C26749 PAND2X1_659/Y D_INPUT_0 0.03fF
C26750 PAND2X1_319/B PAND2X1_556/B 0.03fF
C26751 PAND2X1_55/Y POR2X1_805/A 0.54fF
C26752 PAND2X1_51/CTRL POR2X1_750/B 0.01fF
C26753 PAND2X1_245/CTRL PAND2X1_71/Y 0.01fF
C26754 POR2X1_409/Y POR2X1_94/A 0.02fF
C26755 POR2X1_298/Y PAND2X1_716/B 0.12fF
C26756 POR2X1_649/B POR2X1_121/Y 0.07fF
C26757 PAND2X1_94/A PAND2X1_395/CTRL2 0.00fF
C26758 POR2X1_38/Y PAND2X1_198/Y 0.01fF
C26759 POR2X1_43/B PAND2X1_639/B 0.13fF
C26760 PAND2X1_69/A POR2X1_784/A 0.07fF
C26761 POR2X1_20/O D_INPUT_1 0.01fF
C26762 POR2X1_485/CTRL2 PAND2X1_550/B 0.01fF
C26763 POR2X1_463/Y PAND2X1_41/B 0.03fF
C26764 PAND2X1_65/B POR2X1_796/A 0.03fF
C26765 POR2X1_248/Y VDD 0.00fF
C26766 PAND2X1_663/O PAND2X1_660/B 0.02fF
C26767 PAND2X1_296/O PAND2X1_359/Y 0.02fF
C26768 POR2X1_186/Y POR2X1_151/a_16_28# 0.00fF
C26769 POR2X1_96/Y D_INPUT_0 0.03fF
C26770 PAND2X1_57/B POR2X1_318/A 0.07fF
C26771 PAND2X1_733/A POR2X1_16/Y 0.24fF
C26772 PAND2X1_675/A PAND2X1_190/Y 0.03fF
C26773 POR2X1_23/Y POR2X1_184/CTRL 0.01fF
C26774 POR2X1_477/a_16_28# PAND2X1_52/B 0.03fF
C26775 PAND2X1_795/B PAND2X1_175/B 0.11fF
C26776 POR2X1_719/O POR2X1_502/A 0.29fF
C26777 PAND2X1_404/Y POR2X1_77/Y 0.03fF
C26778 PAND2X1_57/B POR2X1_713/B 0.04fF
C26779 PAND2X1_491/O POR2X1_334/B 0.03fF
C26780 POR2X1_177/Y POR2X1_176/Y 0.54fF
C26781 PAND2X1_55/Y POR2X1_500/Y 0.56fF
C26782 POR2X1_96/A PAND2X1_344/a_56_28# 0.00fF
C26783 POR2X1_85/Y PAND2X1_404/Y 0.05fF
C26784 POR2X1_591/Y POR2X1_42/Y 0.03fF
C26785 POR2X1_562/O POR2X1_341/Y 0.01fF
C26786 POR2X1_27/O POR2X1_9/Y 0.01fF
C26787 PAND2X1_96/B POR2X1_741/Y 0.16fF
C26788 POR2X1_63/CTRL2 POR2X1_38/Y 0.03fF
C26789 POR2X1_348/A POR2X1_334/Y 0.02fF
C26790 POR2X1_192/Y POR2X1_351/O 0.06fF
C26791 POR2X1_750/B PAND2X1_18/B 0.07fF
C26792 POR2X1_722/B PAND2X1_60/B 0.77fF
C26793 POR2X1_378/CTRL POR2X1_62/Y 0.02fF
C26794 POR2X1_493/B VDD 0.11fF
C26795 POR2X1_728/CTRL POR2X1_730/Y 0.01fF
C26796 PAND2X1_81/B PAND2X1_96/B 0.37fF
C26797 POR2X1_78/A PAND2X1_179/CTRL 0.02fF
C26798 POR2X1_414/a_16_28# POR2X1_4/Y 0.02fF
C26799 POR2X1_659/CTRL POR2X1_724/A 0.02fF
C26800 POR2X1_245/Y POR2X1_293/Y 0.07fF
C26801 POR2X1_40/Y POR2X1_599/a_16_28# 0.03fF
C26802 POR2X1_294/B PAND2X1_60/B 0.35fF
C26803 POR2X1_193/a_16_28# POR2X1_631/B 0.00fF
C26804 PAND2X1_216/B PAND2X1_580/B 0.03fF
C26805 POR2X1_775/A PAND2X1_173/CTRL2 0.01fF
C26806 POR2X1_407/A PAND2X1_153/CTRL 0.00fF
C26807 POR2X1_29/Y POR2X1_409/CTRL 0.01fF
C26808 POR2X1_614/A PAND2X1_63/Y 0.08fF
C26809 POR2X1_119/Y PAND2X1_390/Y 0.03fF
C26810 PAND2X1_55/Y POR2X1_128/B 0.03fF
C26811 PAND2X1_111/a_76_28# PAND2X1_32/B 0.02fF
C26812 POR2X1_222/A POR2X1_556/O 0.12fF
C26813 POR2X1_219/a_76_344# POR2X1_631/B 0.00fF
C26814 PAND2X1_482/CTRL POR2X1_483/A 0.01fF
C26815 POR2X1_614/A PAND2X1_495/O 0.07fF
C26816 PAND2X1_96/B PAND2X1_32/B 2.64fF
C26817 POR2X1_491/Y POR2X1_102/Y 0.01fF
C26818 POR2X1_83/m4_208_n4# PAND2X1_231/m4_208_n4# 0.13fF
C26819 PAND2X1_63/Y POR2X1_38/B 0.15fF
C26820 PAND2X1_216/a_76_28# PAND2X1_723/A 0.01fF
C26821 POR2X1_573/A POR2X1_702/A 0.06fF
C26822 POR2X1_795/a_16_28# POR2X1_222/A 0.02fF
C26823 POR2X1_42/Y PAND2X1_154/a_16_344# 0.06fF
C26824 POR2X1_103/CTRL2 PAND2X1_738/Y 0.34fF
C26825 POR2X1_101/Y POR2X1_575/B 0.10fF
C26826 POR2X1_635/B POR2X1_635/A 0.02fF
C26827 PAND2X1_857/A POR2X1_43/B 0.03fF
C26828 PAND2X1_467/Y PAND2X1_707/Y 0.03fF
C26829 PAND2X1_341/B POR2X1_376/B 0.01fF
C26830 POR2X1_140/B POR2X1_276/A 0.68fF
C26831 POR2X1_210/Y POR2X1_532/A 0.35fF
C26832 POR2X1_99/B POR2X1_61/Y 0.03fF
C26833 POR2X1_853/A POR2X1_577/Y 0.01fF
C26834 PAND2X1_195/CTRL2 POR2X1_39/B -0.00fF
C26835 POR2X1_407/A POR2X1_407/CTRL2 0.00fF
C26836 POR2X1_558/A PAND2X1_32/B 0.57fF
C26837 POR2X1_302/CTRL2 POR2X1_188/Y 0.01fF
C26838 PAND2X1_552/B POR2X1_176/Y 0.00fF
C26839 POR2X1_814/A PAND2X1_417/O 0.01fF
C26840 POR2X1_731/CTRL2 POR2X1_738/A -0.00fF
C26841 POR2X1_572/B POR2X1_260/A 0.03fF
C26842 POR2X1_68/A POR2X1_687/A 0.23fF
C26843 POR2X1_685/A POR2X1_614/A 0.01fF
C26844 PAND2X1_779/Y POR2X1_527/Y 0.01fF
C26845 POR2X1_769/A PAND2X1_52/B 0.00fF
C26846 POR2X1_341/Y POR2X1_351/CTRL2 0.01fF
C26847 POR2X1_449/A POR2X1_832/B 0.76fF
C26848 POR2X1_532/A POR2X1_548/A 0.03fF
C26849 PAND2X1_90/CTRL POR2X1_546/A 0.00fF
C26850 POR2X1_43/B POR2X1_260/A 0.06fF
C26851 POR2X1_532/A POR2X1_550/Y 0.01fF
C26852 POR2X1_406/A PAND2X1_737/B 0.01fF
C26853 POR2X1_465/B POR2X1_553/O 0.18fF
C26854 POR2X1_590/A POR2X1_343/B 0.03fF
C26855 POR2X1_529/CTRL2 POR2X1_384/A 0.01fF
C26856 POR2X1_383/A POR2X1_865/B 0.09fF
C26857 POR2X1_356/A POR2X1_326/A 0.03fF
C26858 POR2X1_789/A POR2X1_260/A 0.03fF
C26859 POR2X1_68/B POR2X1_569/A 0.07fF
C26860 POR2X1_177/CTRL2 PAND2X1_552/B 0.00fF
C26861 PAND2X1_111/B PAND2X1_60/B 0.06fF
C26862 POR2X1_61/CTRL2 PAND2X1_69/A 0.01fF
C26863 PAND2X1_501/O POR2X1_72/B 0.01fF
C26864 PAND2X1_90/A PAND2X1_384/O 0.01fF
C26865 PAND2X1_270/CTRL POR2X1_283/A 0.00fF
C26866 POR2X1_614/A POR2X1_260/A 0.16fF
C26867 POR2X1_502/A POR2X1_188/Y 0.03fF
C26868 PAND2X1_620/CTRL2 PAND2X1_651/Y 0.00fF
C26869 POR2X1_493/B PAND2X1_32/B 0.01fF
C26870 PAND2X1_865/Y PAND2X1_862/B 0.03fF
C26871 PAND2X1_592/Y PAND2X1_730/A 0.03fF
C26872 PAND2X1_176/CTRL POR2X1_337/Y 0.01fF
C26873 POR2X1_38/B POR2X1_260/A 4.50fF
C26874 PAND2X1_82/Y PAND2X1_397/CTRL 0.01fF
C26875 D_INPUT_2 POR2X1_5/O 0.02fF
C26876 POR2X1_514/CTRL PAND2X1_48/A 0.03fF
C26877 POR2X1_527/CTRL2 PAND2X1_549/B 0.01fF
C26878 VDD POR2X1_342/B 0.00fF
C26879 POR2X1_416/B POR2X1_760/CTRL 0.01fF
C26880 PAND2X1_824/B POR2X1_206/O 0.06fF
C26881 PAND2X1_661/Y PAND2X1_660/Y 0.01fF
C26882 PAND2X1_6/Y POR2X1_552/CTRL2 0.01fF
C26883 POR2X1_63/Y POR2X1_20/B 0.03fF
C26884 POR2X1_218/A POR2X1_294/A 0.07fF
C26885 POR2X1_528/Y POR2X1_744/CTRL 0.03fF
C26886 POR2X1_218/CTRL2 POR2X1_276/Y 0.01fF
C26887 PAND2X1_87/CTRL2 D_INPUT_0 0.00fF
C26888 PAND2X1_216/B PAND2X1_349/A 0.03fF
C26889 POR2X1_502/Y POR2X1_502/m4_208_n4# 0.10fF
C26890 PAND2X1_271/O POR2X1_556/A 0.02fF
C26891 POR2X1_360/O POR2X1_244/Y 0.20fF
C26892 POR2X1_110/CTRL POR2X1_73/Y 0.03fF
C26893 POR2X1_316/Y POR2X1_55/Y 0.03fF
C26894 POR2X1_366/a_16_28# POR2X1_366/A 0.07fF
C26895 POR2X1_702/CTRL POR2X1_186/B 0.01fF
C26896 PAND2X1_213/Y PAND2X1_704/a_76_28# 0.01fF
C26897 POR2X1_217/O PAND2X1_72/A 0.10fF
C26898 PAND2X1_341/A POR2X1_7/Y 0.23fF
C26899 PAND2X1_65/B POR2X1_863/A 0.06fF
C26900 POR2X1_452/O POR2X1_450/Y 0.00fF
C26901 POR2X1_616/Y POR2X1_38/Y 0.00fF
C26902 POR2X1_860/CTRL2 POR2X1_244/Y 0.00fF
C26903 POR2X1_795/B POR2X1_568/B 0.03fF
C26904 POR2X1_319/a_16_28# POR2X1_169/A 0.03fF
C26905 POR2X1_730/Y POR2X1_444/Y 0.05fF
C26906 PAND2X1_385/O POR2X1_711/Y 0.06fF
C26907 POR2X1_57/A PAND2X1_352/CTRL 0.01fF
C26908 POR2X1_520/a_16_28# POR2X1_520/B 0.02fF
C26909 PAND2X1_39/B POR2X1_260/B 0.13fF
C26910 POR2X1_212/CTRL POR2X1_192/B 0.07fF
C26911 PAND2X1_94/A PAND2X1_527/CTRL2 0.01fF
C26912 PAND2X1_48/B POR2X1_717/B 0.07fF
C26913 POR2X1_730/Y POR2X1_210/A 0.01fF
C26914 POR2X1_283/A POR2X1_4/Y 0.07fF
C26915 PAND2X1_65/B POR2X1_9/Y 0.07fF
C26916 POR2X1_416/B POR2X1_255/Y 0.06fF
C26917 PAND2X1_644/O POR2X1_40/Y 0.02fF
C26918 PAND2X1_73/Y POR2X1_541/B 0.12fF
C26919 POR2X1_118/O POR2X1_77/Y 0.19fF
C26920 POR2X1_119/Y PAND2X1_123/O 0.19fF
C26921 POR2X1_41/B POR2X1_846/CTRL 0.06fF
C26922 PAND2X1_483/CTRL2 POR2X1_252/Y 0.01fF
C26923 POR2X1_431/a_56_344# PAND2X1_390/Y 0.00fF
C26924 PAND2X1_411/a_16_344# PAND2X1_52/B 0.02fF
C26925 POR2X1_4/Y PAND2X1_528/O 0.09fF
C26926 POR2X1_848/CTRL2 PAND2X1_90/Y 0.07fF
C26927 INPUT_1 POR2X1_616/Y 0.03fF
C26928 PAND2X1_562/Y PAND2X1_577/Y 0.47fF
C26929 PAND2X1_611/O POR2X1_734/A 0.11fF
C26930 PAND2X1_435/O POR2X1_677/Y 0.00fF
C26931 POR2X1_614/A PAND2X1_681/O 0.01fF
C26932 PAND2X1_9/Y PAND2X1_58/A 0.03fF
C26933 POR2X1_184/m4_208_n4# POR2X1_91/Y 0.12fF
C26934 POR2X1_416/B PAND2X1_555/Y 0.02fF
C26935 POR2X1_387/Y POR2X1_39/B 0.16fF
C26936 PAND2X1_72/O PAND2X1_72/A 0.15fF
C26937 PAND2X1_138/CTRL2 POR2X1_129/Y 0.03fF
C26938 POR2X1_383/A POR2X1_568/B 0.03fF
C26939 POR2X1_509/CTRL POR2X1_532/A 0.01fF
C26940 PAND2X1_586/CTRL PAND2X1_48/A 0.01fF
C26941 POR2X1_567/A POR2X1_353/A 0.03fF
C26942 POR2X1_409/B PAND2X1_124/Y 0.03fF
C26943 PAND2X1_73/Y POR2X1_848/Y 0.00fF
C26944 POR2X1_643/Y POR2X1_590/A 0.15fF
C26945 POR2X1_54/Y POR2X1_14/Y 0.27fF
C26946 POR2X1_557/B POR2X1_294/A 0.15fF
C26947 POR2X1_554/B POR2X1_105/Y 0.06fF
C26948 POR2X1_588/Y POR2X1_588/O 0.01fF
C26949 PAND2X1_177/a_76_28# PAND2X1_52/B 0.02fF
C26950 POR2X1_260/B POR2X1_805/Y 0.01fF
C26951 D_INPUT_0 POR2X1_37/Y 0.10fF
C26952 PAND2X1_116/CTRL POR2X1_150/Y 0.00fF
C26953 POR2X1_116/A POR2X1_475/A 0.58fF
C26954 PAND2X1_20/A POR2X1_260/B 0.19fF
C26955 PAND2X1_803/O PAND2X1_797/Y 0.01fF
C26956 POR2X1_411/B PAND2X1_340/O 0.01fF
C26957 POR2X1_66/B POR2X1_862/A 0.12fF
C26958 PAND2X1_58/A POR2X1_818/Y 0.03fF
C26959 POR2X1_499/A POR2X1_778/CTRL 0.01fF
C26960 PAND2X1_221/Y PAND2X1_365/a_16_344# 0.02fF
C26961 POR2X1_54/Y PAND2X1_55/CTRL 0.01fF
C26962 PAND2X1_865/Y PAND2X1_716/B 0.03fF
C26963 POR2X1_419/a_16_28# POR2X1_39/B 0.01fF
C26964 POR2X1_664/a_16_28# POR2X1_78/A -0.00fF
C26965 POR2X1_83/B POR2X1_409/B 0.10fF
C26966 POR2X1_188/A POR2X1_862/A 0.01fF
C26967 PAND2X1_273/CTRL2 POR2X1_814/A 0.00fF
C26968 POR2X1_486/O POR2X1_294/B 0.03fF
C26969 PAND2X1_48/A PAND2X1_136/CTRL 0.02fF
C26970 POR2X1_49/Y PAND2X1_477/CTRL 0.01fF
C26971 POR2X1_153/Y PAND2X1_840/Y 0.03fF
C26972 POR2X1_814/B POR2X1_260/B 0.16fF
C26973 POR2X1_176/CTRL2 POR2X1_77/Y 0.00fF
C26974 PAND2X1_214/O POR2X1_40/Y 0.01fF
C26975 POR2X1_174/B POR2X1_78/A 0.05fF
C26976 POR2X1_9/Y POR2X1_245/CTRL2 0.05fF
C26977 POR2X1_43/B POR2X1_329/A 0.14fF
C26978 POR2X1_227/A POR2X1_578/Y 0.03fF
C26979 PAND2X1_231/CTRL2 POR2X1_263/Y 0.01fF
C26980 PAND2X1_634/O POR2X1_290/Y 0.03fF
C26981 POR2X1_257/A PAND2X1_274/CTRL 0.08fF
C26982 POR2X1_98/B PAND2X1_234/CTRL 0.01fF
C26983 PAND2X1_58/A POR2X1_267/A 0.03fF
C26984 POR2X1_66/B PAND2X1_73/Y 0.13fF
C26985 POR2X1_641/CTRL POR2X1_267/A 0.01fF
C26986 POR2X1_260/B POR2X1_325/A 0.03fF
C26987 POR2X1_60/A POR2X1_667/A 0.06fF
C26988 POR2X1_711/Y PAND2X1_692/O 0.02fF
C26989 POR2X1_470/CTRL POR2X1_186/Y 0.01fF
C26990 POR2X1_296/B POR2X1_330/Y 0.16fF
C26991 POR2X1_23/Y PAND2X1_76/Y 0.16fF
C26992 POR2X1_177/Y POR2X1_438/Y 0.01fF
C26993 POR2X1_263/Y POR2X1_230/CTRL2 0.01fF
C26994 POR2X1_54/Y PAND2X1_472/B 0.07fF
C26995 POR2X1_48/A POR2X1_689/CTRL2 0.00fF
C26996 PAND2X1_487/CTRL2 PAND2X1_57/B 0.01fF
C26997 PAND2X1_39/B POR2X1_646/O 0.17fF
C26998 POR2X1_188/A PAND2X1_73/Y 0.13fF
C26999 POR2X1_179/CTRL2 POR2X1_150/Y 0.01fF
C27000 POR2X1_81/a_16_28# PAND2X1_573/B 0.02fF
C27001 POR2X1_326/A PAND2X1_72/A 0.03fF
C27002 POR2X1_329/Y PAND2X1_357/Y 0.03fF
C27003 POR2X1_119/Y POR2X1_158/Y 0.00fF
C27004 PAND2X1_39/B PAND2X1_55/Y 0.13fF
C27005 POR2X1_116/A POR2X1_218/A 0.53fF
C27006 POR2X1_83/B POR2X1_677/CTRL2 0.00fF
C27007 POR2X1_43/B POR2X1_275/Y 0.03fF
C27008 POR2X1_428/a_16_28# POR2X1_236/Y -0.00fF
C27009 POR2X1_54/Y POR2X1_55/Y 0.04fF
C27010 POR2X1_123/a_16_28# POR2X1_556/A 0.02fF
C27011 PAND2X1_631/CTRL2 POR2X1_20/B 0.03fF
C27012 POR2X1_65/A POR2X1_423/O 0.01fF
C27013 POR2X1_385/Y POR2X1_331/CTRL 0.45fF
C27014 POR2X1_142/CTRL POR2X1_49/Y 0.01fF
C27015 POR2X1_260/B POR2X1_513/B 0.05fF
C27016 PAND2X1_56/Y POR2X1_341/A 0.10fF
C27017 POR2X1_341/A POR2X1_795/B 0.03fF
C27018 POR2X1_406/Y D_INPUT_0 0.02fF
C27019 PAND2X1_863/B POR2X1_23/Y 0.21fF
C27020 POR2X1_848/A POR2X1_754/A 0.10fF
C27021 POR2X1_117/O POR2X1_60/A 0.09fF
C27022 POR2X1_640/CTRL PAND2X1_41/B 0.00fF
C27023 POR2X1_188/A POR2X1_830/a_76_344# 0.00fF
C27024 PAND2X1_193/Y PAND2X1_200/B 0.01fF
C27025 PAND2X1_6/Y POR2X1_663/B 0.03fF
C27026 POR2X1_362/Y POR2X1_362/B 0.01fF
C27027 POR2X1_271/B POR2X1_73/Y 0.03fF
C27028 POR2X1_123/Y POR2X1_556/A 0.01fF
C27029 PAND2X1_497/CTRL2 POR2X1_294/B 0.14fF
C27030 POR2X1_608/Y VDD 0.09fF
C27031 POR2X1_496/Y INPUT_0 0.07fF
C27032 PAND2X1_9/Y POR2X1_204/m4_208_n4# 0.15fF
C27033 POR2X1_831/CTRL PAND2X1_69/A 0.01fF
C27034 POR2X1_634/A POR2X1_640/A 0.00fF
C27035 PAND2X1_90/Y PAND2X1_585/CTRL 0.00fF
C27036 POR2X1_400/B VDD 0.13fF
C27037 PAND2X1_48/B PAND2X1_485/CTRL 0.01fF
C27038 PAND2X1_284/Y POR2X1_20/B 0.03fF
C27039 POR2X1_56/O POR2X1_516/B 0.00fF
C27040 POR2X1_805/CTRL2 POR2X1_805/A 0.01fF
C27041 POR2X1_164/Y PAND2X1_717/A 0.00fF
C27042 POR2X1_556/A POR2X1_216/CTRL 0.01fF
C27043 POR2X1_60/A POR2X1_372/O 0.01fF
C27044 POR2X1_49/Y PAND2X1_849/CTRL 0.01fF
C27045 PAND2X1_73/Y POR2X1_859/A 0.42fF
C27046 POR2X1_301/O POR2X1_76/A 0.00fF
C27047 D_INPUT_0 POR2X1_293/Y 0.10fF
C27048 PAND2X1_39/B POR2X1_407/Y 0.05fF
C27049 PAND2X1_246/CTRL POR2X1_101/Y 0.28fF
C27050 POR2X1_567/B POR2X1_740/Y 0.05fF
C27051 POR2X1_78/B POR2X1_200/CTRL2 0.01fF
C27052 POR2X1_20/A D_INPUT_1 0.01fF
C27053 PAND2X1_462/O POR2X1_416/B 0.04fF
C27054 PAND2X1_653/Y PAND2X1_222/A 0.01fF
C27055 PAND2X1_404/Y POR2X1_52/Y 0.03fF
C27056 POR2X1_257/A POR2X1_93/A 1.11fF
C27057 POR2X1_20/B POR2X1_751/a_76_344# 0.01fF
C27058 POR2X1_590/A PAND2X1_152/CTRL 0.00fF
C27059 POR2X1_169/A POR2X1_568/A 0.03fF
C27060 POR2X1_48/A PAND2X1_705/CTRL 0.01fF
C27061 POR2X1_533/Y POR2X1_759/CTRL 0.03fF
C27062 PAND2X1_20/A PAND2X1_516/CTRL 0.01fF
C27063 POR2X1_257/A POR2X1_91/Y 0.17fF
C27064 PAND2X1_864/B PAND2X1_286/B 0.12fF
C27065 PAND2X1_810/A GATE_741 0.04fF
C27066 POR2X1_646/O POR2X1_805/Y 0.07fF
C27067 POR2X1_186/Y PAND2X1_321/O 0.17fF
C27068 PAND2X1_469/B POR2X1_273/m4_208_n4# 0.03fF
C27069 PAND2X1_73/Y POR2X1_828/CTRL 0.01fF
C27070 POR2X1_653/O POR2X1_750/B 0.01fF
C27071 POR2X1_672/A POR2X1_48/A 0.00fF
C27072 POR2X1_78/A PAND2X1_89/O 0.01fF
C27073 PAND2X1_721/B POR2X1_7/B 0.25fF
C27074 POR2X1_99/A VDD 0.15fF
C27075 PAND2X1_48/Y PAND2X1_65/B 0.02fF
C27076 POR2X1_355/A VDD -0.00fF
C27077 POR2X1_277/a_16_28# POR2X1_37/Y 0.03fF
C27078 POR2X1_383/A POR2X1_341/A 0.09fF
C27079 POR2X1_829/A PAND2X1_200/CTRL 0.00fF
C27080 POR2X1_60/A POR2X1_252/O 0.01fF
C27081 POR2X1_808/A POR2X1_435/Y 0.03fF
C27082 POR2X1_60/A PAND2X1_254/CTRL2 0.00fF
C27083 POR2X1_411/B POR2X1_310/Y 0.82fF
C27084 POR2X1_115/O POR2X1_141/Y 0.18fF
C27085 POR2X1_78/A PAND2X1_145/O 0.01fF
C27086 PAND2X1_20/A PAND2X1_55/Y 15.45fF
C27087 POR2X1_262/CTRL POR2X1_40/Y 0.01fF
C27088 PAND2X1_20/A PAND2X1_95/CTRL 0.00fF
C27089 POR2X1_866/A POR2X1_307/A 0.03fF
C27090 POR2X1_814/B POR2X1_723/O 0.01fF
C27091 POR2X1_105/O POR2X1_717/Y 0.01fF
C27092 PAND2X1_784/A POR2X1_55/Y 0.03fF
C27093 POR2X1_751/A POR2X1_816/A 0.01fF
C27094 POR2X1_71/Y POR2X1_72/B 0.03fF
C27095 POR2X1_708/CTRL PAND2X1_65/B 0.01fF
C27096 POR2X1_840/B POR2X1_218/Y 0.10fF
C27097 POR2X1_812/B POR2X1_636/B 0.01fF
C27098 POR2X1_76/a_16_28# POR2X1_366/A 0.03fF
C27099 POR2X1_849/A POR2X1_550/CTRL 0.01fF
C27100 POR2X1_428/Y PAND2X1_710/O 0.03fF
C27101 POR2X1_343/Y POR2X1_76/B 0.58fF
C27102 PAND2X1_844/Y POR2X1_60/Y 0.01fF
C27103 POR2X1_680/Y POR2X1_40/Y 0.04fF
C27104 POR2X1_609/Y POR2X1_73/Y 0.03fF
C27105 PAND2X1_473/B PAND2X1_736/m4_208_n4# 0.15fF
C27106 POR2X1_330/Y POR2X1_363/CTRL2 0.01fF
C27107 POR2X1_220/B POR2X1_210/Y 0.03fF
C27108 POR2X1_270/Y POR2X1_228/Y 0.03fF
C27109 POR2X1_750/B POR2X1_294/B 0.10fF
C27110 POR2X1_366/Y POR2X1_750/B 0.07fF
C27111 PAND2X1_417/a_16_344# POR2X1_186/B 0.01fF
C27112 POR2X1_134/a_16_28# POR2X1_257/A 0.02fF
C27113 POR2X1_119/Y PAND2X1_608/O 0.01fF
C27114 PAND2X1_96/CTRL PAND2X1_55/Y 0.01fF
C27115 POR2X1_72/B POR2X1_42/Y 0.03fF
C27116 PAND2X1_20/A POR2X1_402/A 0.68fF
C27117 POR2X1_48/A POR2X1_387/Y 0.15fF
C27118 POR2X1_695/CTRL POR2X1_48/A 0.01fF
C27119 PAND2X1_94/A PAND2X1_27/O 0.02fF
C27120 POR2X1_143/O POR2X1_376/B 0.01fF
C27121 POR2X1_241/B POR2X1_702/A 0.03fF
C27122 PAND2X1_431/a_16_344# PAND2X1_60/B 0.01fF
C27123 POR2X1_40/Y PAND2X1_324/Y 0.02fF
C27124 POR2X1_624/Y PAND2X1_184/CTRL 0.01fF
C27125 PAND2X1_771/Y PAND2X1_570/B 0.16fF
C27126 PAND2X1_808/Y PAND2X1_354/A 0.03fF
C27127 POR2X1_278/Y PAND2X1_347/Y 0.04fF
C27128 PAND2X1_865/Y POR2X1_250/Y 0.07fF
C27129 POR2X1_355/A POR2X1_741/Y 0.03fF
C27130 D_INPUT_0 POR2X1_408/Y 0.05fF
C27131 POR2X1_814/B PAND2X1_55/Y 0.22fF
C27132 INPUT_6 POR2X1_32/A 0.05fF
C27133 PAND2X1_96/B POR2X1_267/A 0.03fF
C27134 PAND2X1_13/O POR2X1_294/B 0.03fF
C27135 POR2X1_65/A POR2X1_761/CTRL 0.01fF
C27136 PAND2X1_430/O INPUT_5 0.01fF
C27137 POR2X1_451/A PAND2X1_72/A 0.04fF
C27138 PAND2X1_9/O PAND2X1_69/A 0.02fF
C27139 POR2X1_236/Y POR2X1_531/CTRL 0.01fF
C27140 POR2X1_566/A POR2X1_471/O 0.01fF
C27141 POR2X1_356/A POR2X1_480/A 0.10fF
C27142 POR2X1_57/CTRL2 VDD 0.00fF
C27143 POR2X1_52/A POR2X1_497/Y 0.07fF
C27144 PAND2X1_462/B POR2X1_5/Y 0.07fF
C27145 POR2X1_236/Y POR2X1_372/Y 0.12fF
C27146 POR2X1_774/Y POR2X1_800/A 0.03fF
C27147 POR2X1_113/Y POR2X1_590/A 0.03fF
C27148 POR2X1_141/CTRL2 POR2X1_514/Y 0.00fF
C27149 POR2X1_312/Y PAND2X1_566/Y 0.10fF
C27150 PAND2X1_472/CTRL2 POR2X1_23/Y 0.09fF
C27151 POR2X1_409/B PAND2X1_196/CTRL 0.01fF
C27152 POR2X1_66/A PAND2X1_373/O 0.04fF
C27153 POR2X1_284/O POR2X1_325/A 0.01fF
C27154 POR2X1_708/B VDD 0.20fF
C27155 POR2X1_226/a_76_344# POR2X1_382/Y 0.02fF
C27156 POR2X1_814/B POR2X1_402/A 0.00fF
C27157 POR2X1_283/A POR2X1_225/O 0.01fF
C27158 POR2X1_257/A POR2X1_109/Y 0.09fF
C27159 PAND2X1_771/Y PAND2X1_578/a_76_28# 0.02fF
C27160 POR2X1_97/A POR2X1_502/CTRL2 0.02fF
C27161 POR2X1_13/A PAND2X1_351/CTRL 0.01fF
C27162 PAND2X1_65/B PAND2X1_744/CTRL 0.01fF
C27163 POR2X1_78/B POR2X1_740/Y 0.08fF
C27164 PAND2X1_198/a_16_344# PAND2X1_197/Y 0.02fF
C27165 POR2X1_149/B POR2X1_788/a_16_28# 0.07fF
C27166 POR2X1_614/A POR2X1_718/A 0.01fF
C27167 POR2X1_49/Y PAND2X1_341/A 0.03fF
C27168 PAND2X1_562/B POR2X1_90/Y 0.07fF
C27169 POR2X1_519/Y POR2X1_236/Y 0.00fF
C27170 PAND2X1_632/B POR2X1_482/a_16_28# 0.02fF
C27171 POR2X1_192/Y POR2X1_785/A 0.11fF
C27172 PAND2X1_862/B POR2X1_494/Y 0.13fF
C27173 POR2X1_734/A POR2X1_705/a_16_28# 0.03fF
C27174 POR2X1_254/Y PAND2X1_23/Y 0.10fF
C27175 POR2X1_717/O POR2X1_777/B 0.03fF
C27176 POR2X1_536/Y PAND2X1_222/B 0.06fF
C27177 POR2X1_332/Y POR2X1_260/B 0.03fF
C27178 PAND2X1_388/Y POR2X1_40/Y 0.06fF
C27179 POR2X1_48/A PAND2X1_713/CTRL 0.01fF
C27180 PAND2X1_127/a_16_344# POR2X1_66/A 0.02fF
C27181 PAND2X1_669/m4_208_n4# POR2X1_750/Y 0.01fF
C27182 PAND2X1_254/Y PAND2X1_465/B 0.01fF
C27183 POR2X1_49/Y POR2X1_93/A 0.08fF
C27184 POR2X1_785/O POR2X1_785/A 0.19fF
C27185 POR2X1_763/A POR2X1_700/Y 0.21fF
C27186 PAND2X1_406/O PAND2X1_48/A 0.01fF
C27187 POR2X1_253/Y POR2X1_236/Y 0.01fF
C27188 POR2X1_59/CTRL POR2X1_32/A 0.01fF
C27189 POR2X1_49/Y POR2X1_91/Y 0.10fF
C27190 PAND2X1_216/B POR2X1_32/A 0.03fF
C27191 PAND2X1_118/O INPUT_0 0.11fF
C27192 POR2X1_590/A POR2X1_260/A 13.83fF
C27193 POR2X1_518/Y VDD 0.05fF
C27194 PAND2X1_65/B PAND2X1_518/O 0.04fF
C27195 POR2X1_281/CTRL POR2X1_102/Y 0.01fF
C27196 POR2X1_537/Y POR2X1_832/Y 0.00fF
C27197 PAND2X1_55/Y POR2X1_513/B 0.15fF
C27198 PAND2X1_695/CTRL POR2X1_407/Y 0.01fF
C27199 POR2X1_790/A INPUT_0 0.03fF
C27200 PAND2X1_472/A VDD 0.38fF
C27201 PAND2X1_795/O PAND2X1_175/B 0.02fF
C27202 POR2X1_197/O PAND2X1_6/Y 0.16fF
C27203 POR2X1_3/A INPUT_7 0.15fF
C27204 PAND2X1_402/B PAND2X1_402/O 0.00fF
C27205 POR2X1_302/O PAND2X1_32/B 0.01fF
C27206 PAND2X1_812/A PAND2X1_287/Y 0.04fF
C27207 POR2X1_10/a_16_28# POR2X1_32/A 0.02fF
C27208 POR2X1_502/A POR2X1_357/Y 0.05fF
C27209 POR2X1_119/Y POR2X1_265/O 0.08fF
C27210 POR2X1_789/A POR2X1_790/CTRL2 0.03fF
C27211 PAND2X1_405/m4_208_n4# PAND2X1_327/m4_208_n4# 0.05fF
C27212 POR2X1_119/Y PAND2X1_606/a_16_344# 0.02fF
C27213 POR2X1_32/Y VDD 0.01fF
C27214 PAND2X1_546/Y POR2X1_763/Y 0.04fF
C27215 PAND2X1_769/a_76_28# POR2X1_73/Y 0.01fF
C27216 POR2X1_505/a_16_28# POR2X1_669/B 0.09fF
C27217 POR2X1_84/O POR2X1_294/B 0.01fF
C27218 POR2X1_13/A POR2X1_90/Y 0.07fF
C27219 POR2X1_526/a_56_344# PAND2X1_556/B 0.00fF
C27220 PAND2X1_484/O PAND2X1_73/Y 0.05fF
C27221 PAND2X1_41/B POR2X1_101/Y 0.23fF
C27222 PAND2X1_104/O INPUT_1 0.17fF
C27223 POR2X1_447/B POR2X1_836/CTRL2 0.00fF
C27224 PAND2X1_286/a_76_28# PAND2X1_568/B 0.02fF
C27225 POR2X1_337/A POR2X1_814/B 0.01fF
C27226 PAND2X1_798/B POR2X1_488/Y 0.02fF
C27227 POR2X1_333/Y PAND2X1_20/A 0.03fF
C27228 POR2X1_43/B PAND2X1_335/a_76_28# 0.02fF
C27229 POR2X1_38/Y PAND2X1_734/B 0.02fF
C27230 POR2X1_66/A POR2X1_540/Y 0.01fF
C27231 POR2X1_273/CTRL POR2X1_39/B 0.01fF
C27232 PAND2X1_480/O PAND2X1_478/B 0.02fF
C27233 VDD PAND2X1_168/CTRL 0.00fF
C27234 POR2X1_861/CTRL2 POR2X1_218/A 0.01fF
C27235 PAND2X1_222/B PAND2X1_730/B 0.12fF
C27236 POR2X1_833/A PAND2X1_46/O 0.04fF
C27237 POR2X1_696/O POR2X1_394/A 0.01fF
C27238 PAND2X1_476/A POR2X1_263/Y 3.85fF
C27239 POR2X1_380/Y VDD 0.21fF
C27240 POR2X1_57/A PAND2X1_520/a_16_344# 0.02fF
C27241 PAND2X1_371/O PAND2X1_69/A 0.11fF
C27242 POR2X1_96/A PAND2X1_785/a_16_344# 0.01fF
C27243 POR2X1_407/Y POR2X1_513/B 0.02fF
C27244 POR2X1_569/O POR2X1_570/Y 0.03fF
C27245 PAND2X1_65/B PAND2X1_103/CTRL2 0.09fF
C27246 POR2X1_70/O POR2X1_3/A 0.00fF
C27247 POR2X1_144/a_16_28# POR2X1_669/B 0.09fF
C27248 POR2X1_140/B POR2X1_574/CTRL 0.00fF
C27249 POR2X1_68/A PAND2X1_273/O 0.01fF
C27250 POR2X1_786/a_16_28# PAND2X1_60/B 0.01fF
C27251 POR2X1_3/A INPUT_4 0.14fF
C27252 PAND2X1_6/A POR2X1_619/CTRL 0.01fF
C27253 POR2X1_447/B PAND2X1_39/CTRL2 0.05fF
C27254 POR2X1_111/CTRL POR2X1_293/Y 0.02fF
C27255 POR2X1_109/CTRL2 POR2X1_77/Y 0.01fF
C27256 PAND2X1_90/Y POR2X1_151/O 0.02fF
C27257 POR2X1_523/Y POR2X1_559/Y 0.12fF
C27258 POR2X1_668/O POR2X1_260/A 0.08fF
C27259 POR2X1_16/A POR2X1_5/Y 0.14fF
C27260 INPUT_1 POR2X1_381/CTRL 0.01fF
C27261 POR2X1_527/Y VDD 0.00fF
C27262 PAND2X1_386/Y PAND2X1_60/B 0.00fF
C27263 PAND2X1_530/O PAND2X1_32/B 0.01fF
C27264 POR2X1_460/CTRL2 PAND2X1_32/B 0.00fF
C27265 INPUT_2 D_INPUT_2 0.09fF
C27266 PAND2X1_831/O POR2X1_153/Y 0.17fF
C27267 PAND2X1_770/a_56_28# POR2X1_765/Y 0.00fF
C27268 PAND2X1_803/Y POR2X1_7/B 0.02fF
C27269 PAND2X1_737/B PAND2X1_741/B 0.01fF
C27270 POR2X1_416/Y POR2X1_232/Y 0.01fF
C27271 POR2X1_383/A PAND2X1_38/O 0.01fF
C27272 POR2X1_22/A POR2X1_3/CTRL 0.01fF
C27273 PAND2X1_216/B PAND2X1_741/B 0.03fF
C27274 POR2X1_14/Y POR2X1_4/Y 0.16fF
C27275 POR2X1_192/Y PAND2X1_315/a_16_344# 0.02fF
C27276 PAND2X1_631/O PAND2X1_6/A 0.03fF
C27277 PAND2X1_787/A POR2X1_55/Y 0.10fF
C27278 POR2X1_439/Y POR2X1_186/B 0.03fF
C27279 PAND2X1_638/B POR2X1_585/CTRL2 0.05fF
C27280 POR2X1_198/O PAND2X1_88/Y 0.01fF
C27281 POR2X1_278/Y PAND2X1_346/Y 0.09fF
C27282 POR2X1_786/Y POR2X1_804/A 0.01fF
C27283 PAND2X1_107/a_76_28# PAND2X1_65/B 0.02fF
C27284 POR2X1_83/A PAND2X1_243/a_16_344# 0.01fF
C27285 POR2X1_57/A POR2X1_43/B 0.91fF
C27286 POR2X1_553/Y POR2X1_569/A 0.02fF
C27287 POR2X1_366/Y POR2X1_704/CTRL 0.07fF
C27288 PAND2X1_152/a_56_28# PAND2X1_60/B 0.00fF
C27289 POR2X1_567/A POR2X1_254/A 0.05fF
C27290 POR2X1_57/A POR2X1_312/O 0.01fF
C27291 POR2X1_390/B POR2X1_220/Y 0.09fF
C27292 PAND2X1_278/O POR2X1_294/A 0.12fF
C27293 PAND2X1_254/O POR2X1_7/A 0.06fF
C27294 PAND2X1_760/CTRL POR2X1_260/A 0.01fF
C27295 PAND2X1_798/Y PAND2X1_362/A 0.03fF
C27296 POR2X1_96/A PAND2X1_539/Y 0.03fF
C27297 POR2X1_252/Y POR2X1_72/B 0.03fF
C27298 INPUT_1 PAND2X1_734/B 0.02fF
C27299 POR2X1_52/A PAND2X1_160/CTRL2 0.03fF
C27300 POR2X1_567/A POR2X1_750/B 0.06fF
C27301 PAND2X1_90/A POR2X1_569/A 0.14fF
C27302 PAND2X1_64/O PAND2X1_52/B 0.23fF
C27303 PAND2X1_192/CTRL2 PAND2X1_730/A 0.00fF
C27304 POR2X1_45/Y PAND2X1_656/A 0.03fF
C27305 POR2X1_140/B PAND2X1_60/B 0.02fF
C27306 POR2X1_537/a_16_28# POR2X1_480/A 0.02fF
C27307 PAND2X1_357/Y POR2X1_142/Y 0.03fF
C27308 POR2X1_25/Y INPUT_7 0.05fF
C27309 POR2X1_566/A POR2X1_703/Y 0.05fF
C27310 POR2X1_57/CTRL PAND2X1_737/B 0.01fF
C27311 POR2X1_78/B POR2X1_774/A 0.03fF
C27312 PAND2X1_72/CTRL2 PAND2X1_111/B 0.01fF
C27313 PAND2X1_464/Y PAND2X1_241/Y 0.02fF
C27314 POR2X1_752/O INPUT_5 0.16fF
C27315 POR2X1_407/A PAND2X1_60/B 0.06fF
C27316 POR2X1_785/B POR2X1_785/A 0.00fF
C27317 POR2X1_180/CTRL2 VDD -0.00fF
C27318 PAND2X1_658/A POR2X1_748/Y 0.12fF
C27319 POR2X1_788/B POR2X1_535/A 0.04fF
C27320 POR2X1_68/A POR2X1_544/a_16_28# 0.00fF
C27321 POR2X1_356/CTRL2 POR2X1_356/B 0.05fF
C27322 PAND2X1_734/B POR2X1_153/Y 0.06fF
C27323 POR2X1_192/Y POR2X1_186/B 0.32fF
C27324 POR2X1_96/A PAND2X1_507/O 0.02fF
C27325 POR2X1_43/B POR2X1_584/Y 0.07fF
C27326 POR2X1_153/CTRL POR2X1_7/B 0.01fF
C27327 POR2X1_464/Y POR2X1_543/O 0.22fF
C27328 PAND2X1_654/A POR2X1_46/Y 0.01fF
C27329 POR2X1_283/A POR2X1_816/A 0.03fF
C27330 POR2X1_36/B POR2X1_36/O 0.05fF
C27331 POR2X1_546/B POR2X1_546/O 0.06fF
C27332 PAND2X1_270/O POR2X1_73/Y 0.03fF
C27333 POR2X1_614/A POR2X1_725/Y 0.07fF
C27334 PAND2X1_119/a_76_28# PAND2X1_96/B 0.01fF
C27335 POR2X1_189/Y PAND2X1_216/B 0.03fF
C27336 POR2X1_271/A POR2X1_372/Y 0.02fF
C27337 POR2X1_162/a_16_28# POR2X1_161/Y 0.02fF
C27338 POR2X1_468/Y POR2X1_478/B 0.00fF
C27339 POR2X1_835/B POR2X1_835/A 0.00fF
C27340 POR2X1_37/Y POR2X1_90/O 0.17fF
C27341 POR2X1_246/Y PAND2X1_342/O -0.00fF
C27342 POR2X1_829/A PAND2X1_123/Y 0.36fF
C27343 POR2X1_20/B PAND2X1_269/O 0.01fF
C27344 POR2X1_456/B PAND2X1_316/CTRL 0.01fF
C27345 PAND2X1_65/B PAND2X1_134/a_16_344# 0.01fF
C27346 POR2X1_110/Y POR2X1_13/A 0.04fF
C27347 PAND2X1_216/B POR2X1_184/Y 0.03fF
C27348 PAND2X1_659/Y PAND2X1_735/Y 0.02fF
C27349 PAND2X1_661/Y POR2X1_38/Y 0.06fF
C27350 POR2X1_25/Y INPUT_4 0.23fF
C27351 D_GATE_662 POR2X1_544/B 0.45fF
C27352 PAND2X1_793/Y POR2X1_385/Y 0.05fF
C27353 PAND2X1_844/B POR2X1_521/Y 0.07fF
C27354 PAND2X1_56/Y PAND2X1_142/CTRL 0.01fF
C27355 POR2X1_662/CTRL2 POR2X1_725/Y 0.05fF
C27356 POR2X1_332/Y PAND2X1_55/Y 0.05fF
C27357 PAND2X1_472/B POR2X1_4/Y 0.07fF
C27358 PAND2X1_551/O PAND2X1_854/A 0.00fF
C27359 POR2X1_494/Y PAND2X1_716/B 0.03fF
C27360 POR2X1_547/CTRL2 POR2X1_266/A 0.01fF
C27361 POR2X1_596/A POR2X1_596/CTRL 0.01fF
C27362 PAND2X1_534/a_56_28# PAND2X1_60/B 0.00fF
C27363 PAND2X1_23/Y POR2X1_711/B 0.05fF
C27364 PAND2X1_470/a_76_28# PAND2X1_467/Y 0.01fF
C27365 POR2X1_614/A POR2X1_559/A 0.17fF
C27366 POR2X1_740/Y POR2X1_294/A 0.19fF
C27367 PAND2X1_659/Y PAND2X1_218/CTRL2 0.09fF
C27368 PAND2X1_342/CTRL2 POR2X1_153/Y 0.13fF
C27369 POR2X1_274/A POR2X1_814/A 0.01fF
C27370 PAND2X1_476/A PAND2X1_215/B 0.03fF
C27371 POR2X1_717/a_16_28# POR2X1_101/Y 0.04fF
C27372 POR2X1_158/Y PAND2X1_725/B 0.16fF
C27373 POR2X1_119/Y PAND2X1_839/O 0.12fF
C27374 POR2X1_55/Y POR2X1_4/Y 0.03fF
C27375 POR2X1_96/Y PAND2X1_859/B 0.17fF
C27376 POR2X1_38/B POR2X1_559/A 0.00fF
C27377 POR2X1_537/CTRL PAND2X1_60/B 0.01fF
C27378 PAND2X1_850/Y POR2X1_275/O 0.03fF
C27379 POR2X1_294/B PAND2X1_122/CTRL 0.08fF
C27380 POR2X1_802/B POR2X1_532/CTRL 0.04fF
C27381 POR2X1_222/Y POR2X1_540/Y 0.30fF
C27382 POR2X1_163/a_16_28# POR2X1_158/Y 0.00fF
C27383 POR2X1_415/A POR2X1_20/B 0.03fF
C27384 POR2X1_57/A PAND2X1_170/CTRL 0.01fF
C27385 POR2X1_124/B POR2X1_113/B 0.03fF
C27386 POR2X1_78/O POR2X1_571/Y 0.02fF
C27387 POR2X1_480/A PAND2X1_72/A 0.61fF
C27388 POR2X1_558/A POR2X1_558/Y 0.01fF
C27389 POR2X1_554/Y POR2X1_632/Y 0.05fF
C27390 D_INPUT_3 POR2X1_5/CTRL2 0.01fF
C27391 POR2X1_416/B POR2X1_46/Y 0.26fF
C27392 PAND2X1_69/A POR2X1_512/O 0.10fF
C27393 POR2X1_575/O POR2X1_574/Y 0.02fF
C27394 POR2X1_7/A PAND2X1_507/O 0.01fF
C27395 POR2X1_669/B PAND2X1_87/O 0.02fF
C27396 POR2X1_814/A POR2X1_269/A 0.01fF
C27397 POR2X1_78/B POR2X1_147/a_16_28# 0.00fF
C27398 POR2X1_140/B POR2X1_554/O 0.01fF
C27399 INPUT_0 PAND2X1_332/Y 0.07fF
C27400 PAND2X1_661/Y POR2X1_153/Y 0.19fF
C27401 PAND2X1_82/CTRL2 POR2X1_294/A 0.00fF
C27402 POR2X1_343/Y PAND2X1_71/O 0.02fF
C27403 POR2X1_532/A POR2X1_540/Y 0.02fF
C27404 POR2X1_81/CTRL2 PAND2X1_510/B 0.01fF
C27405 PAND2X1_726/O POR2X1_39/B 0.02fF
C27406 POR2X1_270/Y POR2X1_657/Y 0.00fF
C27407 POR2X1_850/a_16_28# POR2X1_737/A 0.02fF
C27408 POR2X1_678/a_16_28# POR2X1_260/B 0.01fF
C27409 PAND2X1_844/Y PAND2X1_351/A 0.01fF
C27410 POR2X1_275/A D_INPUT_0 0.03fF
C27411 POR2X1_16/A POR2X1_599/CTRL 0.12fF
C27412 PAND2X1_618/CTRL2 POR2X1_29/A 0.03fF
C27413 POR2X1_119/Y PAND2X1_839/B 0.03fF
C27414 POR2X1_532/A POR2X1_532/CTRL 0.01fF
C27415 PAND2X1_90/A PAND2X1_72/A 0.03fF
C27416 PAND2X1_93/B PAND2X1_268/O 0.04fF
C27417 PAND2X1_674/CTRL2 PAND2X1_72/A 0.01fF
C27418 POR2X1_717/Y POR2X1_717/B 0.03fF
C27419 POR2X1_569/A POR2X1_572/Y 0.04fF
C27420 POR2X1_54/Y POR2X1_476/A 0.03fF
C27421 POR2X1_20/B POR2X1_432/CTRL 0.01fF
C27422 PAND2X1_29/CTRL2 PAND2X1_52/B 0.15fF
C27423 PAND2X1_813/CTRL POR2X1_266/A 0.01fF
C27424 POR2X1_334/B POR2X1_768/A 0.05fF
C27425 POR2X1_445/A POR2X1_66/A 0.04fF
C27426 POR2X1_150/Y PAND2X1_794/O 0.03fF
C27427 POR2X1_178/a_56_344# POR2X1_416/B 0.01fF
C27428 PAND2X1_48/Y POR2X1_814/A 0.09fF
C27429 POR2X1_610/Y POR2X1_590/A 0.03fF
C27430 POR2X1_191/CTRL POR2X1_568/Y 0.01fF
C27431 POR2X1_782/A POR2X1_568/A 0.01fF
C27432 POR2X1_635/O POR2X1_750/B 0.01fF
C27433 POR2X1_866/A POR2X1_801/B 0.00fF
C27434 POR2X1_774/A POR2X1_294/A 0.07fF
C27435 POR2X1_191/Y POR2X1_545/a_16_28# 0.03fF
C27436 PAND2X1_337/O PAND2X1_336/Y 0.03fF
C27437 POR2X1_411/B POR2X1_423/Y 0.06fF
C27438 POR2X1_673/A POR2X1_622/B 0.02fF
C27439 POR2X1_260/B POR2X1_605/CTRL2 0.01fF
C27440 POR2X1_442/a_56_344# POR2X1_40/Y 0.01fF
C27441 POR2X1_834/Y POR2X1_513/A 0.05fF
C27442 POR2X1_68/A POR2X1_661/A 0.10fF
C27443 PAND2X1_656/O PAND2X1_656/B 0.00fF
C27444 PAND2X1_699/CTRL VDD 0.00fF
C27445 PAND2X1_20/A PAND2X1_609/a_16_344# 0.02fF
C27446 POR2X1_20/B POR2X1_692/Y 0.01fF
C27447 POR2X1_316/Y POR2X1_129/Y 0.32fF
C27448 POR2X1_552/a_16_28# POR2X1_552/A 0.04fF
C27449 POR2X1_408/Y POR2X1_90/O 0.56fF
C27450 POR2X1_119/Y PAND2X1_476/A 0.05fF
C27451 POR2X1_484/Y VDD 0.00fF
C27452 POR2X1_60/A D_INPUT_0 0.19fF
C27453 POR2X1_326/A POR2X1_532/O 0.18fF
C27454 POR2X1_496/Y POR2X1_102/Y 1.55fF
C27455 POR2X1_634/A D_INPUT_0 0.01fF
C27456 PAND2X1_576/B POR2X1_72/B 0.03fF
C27457 POR2X1_260/B PAND2X1_526/CTRL 0.01fF
C27458 POR2X1_24/O POR2X1_23/Y 0.01fF
C27459 POR2X1_341/A INPUT_0 0.07fF
C27460 PAND2X1_620/Y POR2X1_422/a_56_344# 0.00fF
C27461 POR2X1_37/Y POR2X1_609/O 0.16fF
C27462 POR2X1_666/CTRL PAND2X1_719/Y 0.02fF
C27463 PAND2X1_341/B POR2X1_86/a_76_344# 0.00fF
C27464 POR2X1_696/O POR2X1_669/B 0.03fF
C27465 POR2X1_631/CTRL2 POR2X1_590/A 0.00fF
C27466 POR2X1_67/A POR2X1_72/B 0.11fF
C27467 POR2X1_260/B VDD 3.01fF
C27468 PAND2X1_416/a_16_344# POR2X1_859/A 0.07fF
C27469 POR2X1_622/B D_INPUT_1 0.01fF
C27470 PAND2X1_206/A PAND2X1_351/Y 0.00fF
C27471 POR2X1_102/Y PAND2X1_733/A 0.00fF
C27472 POR2X1_186/Y POR2X1_555/B 0.00fF
C27473 POR2X1_3/A POR2X1_18/O 0.37fF
C27474 POR2X1_571/Y POR2X1_500/O 0.02fF
C27475 POR2X1_818/Y POR2X1_415/CTRL 0.01fF
C27476 POR2X1_814/B POR2X1_174/A 0.07fF
C27477 POR2X1_218/Y POR2X1_217/CTRL 0.03fF
C27478 POR2X1_482/CTRL VDD 0.00fF
C27479 POR2X1_23/Y PAND2X1_480/B 0.09fF
C27480 PAND2X1_206/A PAND2X1_101/CTRL 0.01fF
C27481 POR2X1_466/A POR2X1_724/CTRL2 0.03fF
C27482 POR2X1_130/A D_INPUT_0 0.03fF
C27483 PAND2X1_860/A POR2X1_394/A 0.03fF
C27484 POR2X1_87/B POR2X1_294/A 0.02fF
C27485 PAND2X1_640/O POR2X1_826/Y 0.02fF
C27486 POR2X1_186/Y POR2X1_330/Y 0.10fF
C27487 POR2X1_445/A POR2X1_222/Y 0.03fF
C27488 POR2X1_66/B POR2X1_61/Y 0.08fF
C27489 POR2X1_663/O POR2X1_78/A 0.16fF
C27490 POR2X1_658/O POR2X1_532/A 0.02fF
C27491 PAND2X1_585/a_76_28# PAND2X1_41/B 0.01fF
C27492 PAND2X1_92/CTRL POR2X1_66/A 0.28fF
C27493 PAND2X1_841/CTRL2 POR2X1_23/Y 0.01fF
C27494 POR2X1_24/a_16_28# POR2X1_40/Y 0.01fF
C27495 POR2X1_63/Y POR2X1_73/Y 0.03fF
C27496 POR2X1_814/A PAND2X1_103/CTRL2 0.01fF
C27497 POR2X1_634/A PAND2X1_90/Y 0.79fF
C27498 POR2X1_260/B POR2X1_741/Y 0.03fF
C27499 POR2X1_647/B POR2X1_865/CTRL2 0.01fF
C27500 POR2X1_324/B POR2X1_324/A 0.00fF
C27501 PAND2X1_319/B POR2X1_411/B 0.07fF
C27502 PAND2X1_640/B POR2X1_42/Y 0.03fF
C27503 POR2X1_83/B PAND2X1_520/CTRL 0.00fF
C27504 PAND2X1_81/B POR2X1_260/B 0.00fF
C27505 PAND2X1_48/B PAND2X1_277/O 0.06fF
C27506 POR2X1_814/B POR2X1_860/A 0.03fF
C27507 PAND2X1_128/O PAND2X1_771/Y 0.18fF
C27508 PAND2X1_859/B POR2X1_37/Y 3.55fF
C27509 POR2X1_754/Y POR2X1_7/B 0.04fF
C27510 POR2X1_389/a_16_28# POR2X1_260/B 0.03fF
C27511 POR2X1_186/Y POR2X1_776/O 0.01fF
C27512 POR2X1_558/O POR2X1_558/B 0.01fF
C27513 POR2X1_257/A POR2X1_425/Y 0.15fF
C27514 POR2X1_777/B POR2X1_573/O 0.03fF
C27515 POR2X1_48/A PAND2X1_726/O 0.01fF
C27516 POR2X1_334/B PAND2X1_63/O 0.03fF
C27517 POR2X1_848/A POR2X1_793/A 0.03fF
C27518 POR2X1_250/Y PAND2X1_343/O 0.06fF
C27519 POR2X1_466/A PAND2X1_183/a_76_28# 0.03fF
C27520 POR2X1_760/A PAND2X1_539/Y 0.02fF
C27521 POR2X1_445/A POR2X1_532/A 0.06fF
C27522 POR2X1_362/B POR2X1_405/a_76_344# 0.01fF
C27523 POR2X1_260/B PAND2X1_32/B 10.39fF
C27524 GATE_479 PAND2X1_712/B 0.03fF
C27525 PAND2X1_561/A VDD -0.00fF
C27526 POR2X1_558/B POR2X1_267/Y 0.00fF
C27527 POR2X1_659/A POR2X1_724/A 0.09fF
C27528 INPUT_3 POR2X1_283/A 0.32fF
C27529 PAND2X1_786/CTRL2 POR2X1_293/Y 0.13fF
C27530 POR2X1_32/A PAND2X1_717/CTRL 0.01fF
C27531 POR2X1_319/A PAND2X1_314/O 0.15fF
C27532 PAND2X1_56/Y POR2X1_269/CTRL 0.01fF
C27533 POR2X1_695/a_16_28# POR2X1_425/Y 0.02fF
C27534 PAND2X1_786/a_76_28# PAND2X1_84/Y 0.02fF
C27535 POR2X1_865/O POR2X1_866/A 0.01fF
C27536 POR2X1_278/Y PAND2X1_354/A 0.03fF
C27537 POR2X1_590/A PAND2X1_110/O 0.04fF
C27538 PAND2X1_66/O POR2X1_38/Y 0.01fF
C27539 POR2X1_63/Y PAND2X1_244/B 0.03fF
C27540 POR2X1_78/A POR2X1_563/Y 0.03fF
C27541 D_INPUT_0 POR2X1_844/B 2.19fF
C27542 POR2X1_263/Y PAND2X1_734/CTRL 0.01fF
C27543 POR2X1_68/A POR2X1_68/a_16_28# 0.03fF
C27544 PAND2X1_63/Y POR2X1_66/A 0.08fF
C27545 POR2X1_840/CTRL2 D_INPUT_0 0.03fF
C27546 PAND2X1_803/A VDD 0.00fF
C27547 POR2X1_166/O POR2X1_438/Y 0.01fF
C27548 POR2X1_687/A POR2X1_676/CTRL2 0.03fF
C27549 POR2X1_607/A POR2X1_411/a_16_28# 0.04fF
C27550 PAND2X1_453/a_76_28# POR2X1_60/A 0.02fF
C27551 POR2X1_25/Y POR2X1_18/O 0.00fF
C27552 POR2X1_488/O PAND2X1_738/Y 0.04fF
C27553 POR2X1_130/A PAND2X1_90/Y 0.17fF
C27554 POR2X1_52/A POR2X1_423/Y 0.03fF
C27555 POR2X1_612/A POR2X1_4/Y 0.02fF
C27556 PAND2X1_863/B POR2X1_250/A 0.03fF
C27557 PAND2X1_401/O POR2X1_14/Y 0.02fF
C27558 POR2X1_272/CTRL2 POR2X1_42/Y 0.01fF
C27559 POR2X1_630/CTRL2 POR2X1_510/Y 0.01fF
C27560 POR2X1_96/A PAND2X1_721/CTRL 0.01fF
C27561 D_INPUT_3 POR2X1_48/A 0.93fF
C27562 D_INPUT_0 POR2X1_573/A 0.06fF
C27563 POR2X1_79/Y PAND2X1_740/CTRL 0.01fF
C27564 POR2X1_267/A PAND2X1_767/CTRL2 0.00fF
C27565 POR2X1_29/A POR2X1_90/Y 0.03fF
C27566 POR2X1_68/A POR2X1_866/CTRL2 0.12fF
C27567 POR2X1_516/CTRL POR2X1_60/A 0.01fF
C27568 POR2X1_93/Y POR2X1_283/A 0.26fF
C27569 POR2X1_566/A PAND2X1_90/Y 0.39fF
C27570 PAND2X1_266/O POR2X1_7/Y 0.02fF
C27571 POR2X1_43/B PAND2X1_556/a_16_344# 0.02fF
C27572 POR2X1_416/B POR2X1_698/Y 0.15fF
C27573 POR2X1_409/B POR2X1_278/A 0.04fF
C27574 GATE_366 VDD 0.00fF
C27575 POR2X1_287/B PAND2X1_371/CTRL 0.01fF
C27576 PAND2X1_231/O POR2X1_293/Y 0.02fF
C27577 POR2X1_66/B POR2X1_35/Y 0.07fF
C27578 POR2X1_41/B PAND2X1_842/a_16_344# 0.01fF
C27579 PAND2X1_474/Y INPUT_0 0.03fF
C27580 POR2X1_14/Y POR2X1_816/A 0.03fF
C27581 PAND2X1_23/Y PAND2X1_41/B 13.03fF
C27582 POR2X1_569/CTRL2 POR2X1_853/A 0.01fF
C27583 POR2X1_8/Y POR2X1_126/CTRL2 0.01fF
C27584 PAND2X1_265/CTRL2 PAND2X1_32/B 0.01fF
C27585 POR2X1_45/O PAND2X1_480/B 0.32fF
C27586 PAND2X1_90/A PAND2X1_412/O 0.07fF
C27587 POR2X1_14/Y D_INPUT_1 0.06fF
C27588 POR2X1_41/B PAND2X1_713/B 0.02fF
C27589 PAND2X1_673/Y VDD 0.67fF
C27590 POR2X1_614/A PAND2X1_677/CTRL2 0.01fF
C27591 PAND2X1_74/CTRL2 POR2X1_702/A 0.00fF
C27592 PAND2X1_202/O VDD 0.00fF
C27593 POR2X1_62/Y POR2X1_88/A 0.00fF
C27594 PAND2X1_48/Y POR2X1_260/Y 0.02fF
C27595 POR2X1_556/A PAND2X1_48/A 0.03fF
C27596 POR2X1_13/A INPUT_0 0.66fF
C27597 POR2X1_49/Y PAND2X1_551/A 0.01fF
C27598 POR2X1_407/A POR2X1_750/B 0.19fF
C27599 POR2X1_728/O POR2X1_728/B 0.00fF
C27600 POR2X1_58/O POR2X1_58/Y 0.01fF
C27601 PAND2X1_437/CTRL2 PAND2X1_72/A 0.01fF
C27602 POR2X1_383/A POR2X1_269/CTRL 0.01fF
C27603 POR2X1_48/A PAND2X1_350/m4_208_n4# 0.12fF
C27604 POR2X1_65/A POR2X1_693/Y 0.01fF
C27605 POR2X1_19/O POR2X1_4/Y 0.05fF
C27606 PAND2X1_93/B POR2X1_675/Y 0.03fF
C27607 PAND2X1_6/Y PAND2X1_7/Y 0.03fF
C27608 POR2X1_848/A POR2X1_753/CTRL2 0.05fF
C27609 POR2X1_257/A PAND2X1_725/O 0.16fF
C27610 POR2X1_614/A POR2X1_254/O 0.01fF
C27611 POR2X1_65/A PAND2X1_105/O 0.01fF
C27612 PAND2X1_828/CTRL2 POR2X1_599/A 0.01fF
C27613 VDD POR2X1_340/CTRL 0.00fF
C27614 PAND2X1_475/O POR2X1_38/Y 0.04fF
C27615 POR2X1_205/Y VDD 0.19fF
C27616 POR2X1_590/A POR2X1_725/Y 0.19fF
C27617 POR2X1_641/O PAND2X1_60/B 0.01fF
C27618 PAND2X1_55/Y VDD 4.54fF
C27619 POR2X1_502/A POR2X1_578/Y 0.10fF
C27620 POR2X1_66/A POR2X1_260/A 0.31fF
C27621 PAND2X1_23/Y POR2X1_402/B 0.00fF
C27622 PAND2X1_218/O PAND2X1_741/B 0.05fF
C27623 POR2X1_614/A POR2X1_549/O 0.03fF
C27624 POR2X1_389/O POR2X1_130/A 0.04fF
C27625 PAND2X1_93/B POR2X1_544/B 0.03fF
C27626 POR2X1_655/Y POR2X1_307/A 0.02fF
C27627 POR2X1_287/B PAND2X1_69/A 0.06fF
C27628 POR2X1_215/a_56_344# POR2X1_205/Y 0.00fF
C27629 PAND2X1_820/O POR2X1_669/B 0.52fF
C27630 POR2X1_311/O POR2X1_102/Y 0.02fF
C27631 POR2X1_166/CTRL2 PAND2X1_714/A 0.01fF
C27632 PAND2X1_859/A POR2X1_382/Y 0.13fF
C27633 PAND2X1_48/B PAND2X1_751/CTRL2 0.10fF
C27634 POR2X1_78/A PAND2X1_528/O 0.05fF
C27635 POR2X1_43/B PAND2X1_84/Y 0.03fF
C27636 POR2X1_496/Y PAND2X1_748/a_16_344# 0.05fF
C27637 PAND2X1_46/O PAND2X1_111/B 0.02fF
C27638 PAND2X1_48/B POR2X1_468/B 0.03fF
C27639 POR2X1_72/B PAND2X1_168/O 0.03fF
C27640 POR2X1_108/Y POR2X1_60/A 0.01fF
C27641 POR2X1_23/Y POR2X1_373/Y 0.01fF
C27642 PAND2X1_30/O POR2X1_451/A 0.06fF
C27643 POR2X1_43/B PAND2X1_636/CTRL 0.01fF
C27644 PAND2X1_520/O POR2X1_519/Y 0.00fF
C27645 PAND2X1_520/CTRL2 PAND2X1_642/B 0.01fF
C27646 POR2X1_402/A VDD 0.00fF
C27647 POR2X1_66/B PAND2X1_765/O 0.01fF
C27648 POR2X1_41/B PAND2X1_736/A 0.07fF
C27649 POR2X1_49/Y PAND2X1_338/B 0.00fF
C27650 PAND2X1_69/A POR2X1_778/CTRL 0.00fF
C27651 POR2X1_355/B D_GATE_662 0.07fF
C27652 PAND2X1_90/A PAND2X1_667/m4_208_n4# 0.15fF
C27653 POR2X1_78/A POR2X1_675/Y 0.03fF
C27654 PAND2X1_365/B VDD 0.11fF
C27655 PAND2X1_803/Y PAND2X1_220/Y 0.14fF
C27656 POR2X1_303/CTRL POR2X1_274/A 0.03fF
C27657 POR2X1_7/B POR2X1_42/Y 0.32fF
C27658 PAND2X1_473/CTRL PAND2X1_473/B 0.06fF
C27659 POR2X1_185/O PAND2X1_57/B 0.11fF
C27660 PAND2X1_594/CTRL2 POR2X1_151/Y 0.00fF
C27661 POR2X1_52/A POR2X1_57/Y 0.02fF
C27662 PAND2X1_675/A PAND2X1_182/A 0.03fF
C27663 POR2X1_814/B POR2X1_360/CTRL 0.01fF
C27664 PAND2X1_490/CTRL2 PAND2X1_57/B 0.03fF
C27665 POR2X1_759/A VDD 0.00fF
C27666 PAND2X1_735/O POR2X1_816/A 0.01fF
C27667 POR2X1_273/Y POR2X1_46/Y 0.05fF
C27668 POR2X1_833/CTRL2 POR2X1_294/B 0.01fF
C27669 PAND2X1_69/A PAND2X1_8/Y 0.20fF
C27670 POR2X1_72/B PAND2X1_550/B 0.06fF
C27671 POR2X1_343/Y POR2X1_499/A 0.05fF
C27672 PAND2X1_579/B POR2X1_498/A 0.01fF
C27673 POR2X1_590/A POR2X1_559/A 0.08fF
C27674 PAND2X1_57/B POR2X1_705/CTRL 0.01fF
C27675 PAND2X1_591/O PAND2X1_48/A 0.03fF
C27676 POR2X1_407/Y VDD 0.93fF
C27677 POR2X1_409/B POR2X1_117/Y 0.01fF
C27678 PAND2X1_107/CTRL POR2X1_640/Y 0.01fF
C27679 POR2X1_78/A POR2X1_544/B 1.49fF
C27680 POR2X1_447/B POR2X1_567/B 0.03fF
C27681 POR2X1_16/A POR2X1_491/CTRL 0.08fF
C27682 PAND2X1_494/CTRL2 POR2X1_294/B 0.13fF
C27683 POR2X1_7/B POR2X1_309/Y 0.03fF
C27684 POR2X1_826/Y POR2X1_77/Y 0.04fF
C27685 PAND2X1_55/Y POR2X1_741/Y 0.03fF
C27686 PAND2X1_23/Y POR2X1_130/Y 0.01fF
C27687 POR2X1_566/A POR2X1_336/CTRL 0.01fF
C27688 POR2X1_783/Y VDD 0.10fF
C27689 PAND2X1_549/B POR2X1_5/Y 0.03fF
C27690 PAND2X1_676/CTRL2 PAND2X1_735/Y 0.05fF
C27691 POR2X1_116/Y POR2X1_392/B 0.00fF
C27692 POR2X1_707/CTRL PAND2X1_41/B 0.01fF
C27693 POR2X1_777/B POR2X1_456/B 0.05fF
C27694 PAND2X1_562/B PAND2X1_348/CTRL 0.06fF
C27695 PAND2X1_521/CTRL INPUT_0 0.01fF
C27696 POR2X1_646/O PAND2X1_32/B 0.09fF
C27697 PAND2X1_94/A PAND2X1_42/O 0.03fF
C27698 POR2X1_130/A POR2X1_361/O 0.05fF
C27699 POR2X1_188/A PAND2X1_701/CTRL 0.00fF
C27700 POR2X1_51/A INPUT_6 0.00fF
C27701 POR2X1_55/Y POR2X1_816/A 0.03fF
C27702 PAND2X1_862/Y POR2X1_516/Y 0.03fF
C27703 PAND2X1_575/O POR2X1_46/Y 0.27fF
C27704 POR2X1_844/a_16_28# POR2X1_546/A 0.02fF
C27705 D_INPUT_1 POR2X1_55/Y 0.03fF
C27706 PAND2X1_740/Y POR2X1_283/A 0.70fF
C27707 PAND2X1_569/B PAND2X1_544/CTRL 0.03fF
C27708 PAND2X1_564/CTRL POR2X1_765/Y 0.01fF
C27709 POR2X1_809/A POR2X1_866/CTRL 0.01fF
C27710 POR2X1_49/Y POR2X1_599/CTRL2 0.01fF
C27711 INPUT_1 POR2X1_585/O 0.01fF
C27712 PAND2X1_55/Y PAND2X1_32/B 0.14fF
C27713 PAND2X1_445/CTRL POR2X1_90/Y 0.01fF
C27714 PAND2X1_6/Y PAND2X1_275/O 0.01fF
C27715 PAND2X1_65/B POR2X1_456/B 0.06fF
C27716 POR2X1_559/B INPUT_0 0.04fF
C27717 PAND2X1_48/B POR2X1_68/B 0.02fF
C27718 POR2X1_337/A VDD 0.00fF
C27719 POR2X1_188/A POR2X1_851/O 0.01fF
C27720 PAND2X1_832/CTRL POR2X1_153/Y 0.01fF
C27721 POR2X1_136/Y POR2X1_46/Y 0.12fF
C27722 POR2X1_316/Y POR2X1_37/Y 0.03fF
C27723 POR2X1_567/B POR2X1_510/O 0.26fF
C27724 PAND2X1_28/O VDD 0.00fF
C27725 PAND2X1_221/CTRL PAND2X1_730/A 0.00fF
C27726 PAND2X1_790/Y POR2X1_93/A 0.01fF
C27727 INPUT_0 PAND2X1_510/B 0.05fF
C27728 POR2X1_62/Y PAND2X1_459/CTRL 0.01fF
C27729 POR2X1_635/B POR2X1_635/CTRL2 0.02fF
C27730 POR2X1_813/Y PAND2X1_673/Y 0.18fF
C27731 PAND2X1_365/B PAND2X1_365/O 0.00fF
C27732 PAND2X1_499/Y PAND2X1_861/O 0.06fF
C27733 POR2X1_32/CTRL INPUT_3 0.49fF
C27734 PAND2X1_13/CTRL POR2X1_186/B 0.01fF
C27735 PAND2X1_319/B PAND2X1_317/Y 0.12fF
C27736 POR2X1_213/CTRL2 POR2X1_532/A 0.03fF
C27737 PAND2X1_319/B POR2X1_152/A 0.01fF
C27738 POR2X1_853/A POR2X1_578/CTRL2 0.01fF
C27739 PAND2X1_613/O PAND2X1_52/B 0.20fF
C27740 PAND2X1_93/CTRL2 PAND2X1_88/Y 0.01fF
C27741 POR2X1_311/CTRL2 POR2X1_7/B 0.00fF
C27742 PAND2X1_55/Y PAND2X1_312/O 0.04fF
C27743 PAND2X1_69/A POR2X1_705/CTRL2 0.03fF
C27744 D_INPUT_0 PAND2X1_339/CTRL2 0.06fF
C27745 PAND2X1_20/A PAND2X1_692/a_76_28# 0.01fF
C27746 POR2X1_780/O POR2X1_294/A 0.03fF
C27747 PAND2X1_23/Y POR2X1_228/Y 0.06fF
C27748 PAND2X1_63/B POR2X1_404/Y 0.03fF
C27749 INPUT_1 POR2X1_58/a_16_28# 0.03fF
C27750 POR2X1_186/Y POR2X1_703/O 0.06fF
C27751 POR2X1_776/B POR2X1_566/B 0.22fF
C27752 POR2X1_68/A PAND2X1_177/O 0.02fF
C27753 POR2X1_327/Y POR2X1_302/CTRL2 0.01fF
C27754 POR2X1_383/A PAND2X1_110/CTRL 0.00fF
C27755 POR2X1_360/A POR2X1_101/Y 0.09fF
C27756 PAND2X1_652/O POR2X1_83/B 0.04fF
C27757 PAND2X1_473/B PAND2X1_853/B 0.06fF
C27758 POR2X1_186/Y POR2X1_337/Y 0.07fF
C27759 POR2X1_804/A PAND2X1_311/CTRL 0.27fF
C27760 POR2X1_124/O POR2X1_276/Y 0.06fF
C27761 POR2X1_407/Y PAND2X1_32/B 0.03fF
C27762 POR2X1_22/O POR2X1_260/A 0.03fF
C27763 POR2X1_840/B PAND2X1_96/B 0.03fF
C27764 POR2X1_406/CTRL2 PAND2X1_737/B 0.01fF
C27765 POR2X1_333/Y VDD 0.14fF
C27766 POR2X1_78/B POR2X1_398/CTRL 0.01fF
C27767 POR2X1_123/a_16_28# PAND2X1_60/B 0.03fF
C27768 POR2X1_383/A POR2X1_861/O 0.01fF
C27769 POR2X1_52/A PAND2X1_477/A 0.02fF
C27770 POR2X1_458/O POR2X1_343/B 0.02fF
C27771 POR2X1_432/O POR2X1_77/Y 0.01fF
C27772 PAND2X1_675/A POR2X1_283/A 11.64fF
C27773 PAND2X1_148/Y PAND2X1_149/A 0.05fF
C27774 POR2X1_220/B POR2X1_161/CTRL 0.03fF
C27775 PAND2X1_469/B POR2X1_283/A 0.10fF
C27776 POR2X1_337/A POR2X1_741/Y 0.07fF
C27777 POR2X1_383/A POR2X1_712/Y 0.01fF
C27778 PAND2X1_382/CTRL POR2X1_816/A 0.00fF
C27779 POR2X1_516/CTRL POR2X1_516/A 0.01fF
C27780 PAND2X1_281/CTRL VDD 0.00fF
C27781 POR2X1_537/Y POR2X1_480/A 0.03fF
C27782 PAND2X1_733/A POR2X1_761/A 0.03fF
C27783 POR2X1_327/Y POR2X1_502/A 0.07fF
C27784 PAND2X1_58/A PAND2X1_56/A 1.26fF
C27785 POR2X1_814/A POR2X1_467/O 0.37fF
C27786 POR2X1_123/Y PAND2X1_60/B 0.01fF
C27787 PAND2X1_489/CTRL PAND2X1_798/B 0.03fF
C27788 POR2X1_832/B POR2X1_592/A 0.07fF
C27789 PAND2X1_363/a_76_28# POR2X1_42/Y 0.01fF
C27790 PAND2X1_855/O PAND2X1_854/A 0.03fF
C27791 POR2X1_110/CTRL2 POR2X1_13/A 0.00fF
C27792 POR2X1_71/CTRL POR2X1_293/Y 0.05fF
C27793 PAND2X1_6/Y PAND2X1_300/CTRL2 0.01fF
C27794 POR2X1_532/A PAND2X1_534/CTRL 0.00fF
C27795 POR2X1_222/Y POR2X1_260/A 0.06fF
C27796 PAND2X1_137/Y POR2X1_131/A 0.03fF
C27797 PAND2X1_615/CTRL2 PAND2X1_63/B 0.01fF
C27798 POR2X1_72/B POR2X1_387/CTRL2 0.03fF
C27799 POR2X1_96/B POR2X1_38/B 0.03fF
C27800 POR2X1_220/Y POR2X1_553/a_16_28# 0.03fF
C27801 POR2X1_7/A POR2X1_382/Y 0.03fF
C27802 VDD PAND2X1_338/CTRL 0.00fF
C27803 POR2X1_54/Y POR2X1_848/CTRL2 0.03fF
C27804 POR2X1_580/a_16_28# POR2X1_192/B 0.11fF
C27805 POR2X1_54/Y PAND2X1_87/CTRL2 0.13fF
C27806 POR2X1_102/Y PAND2X1_332/Y 0.03fF
C27807 D_INPUT_7 PAND2X1_581/CTRL 0.03fF
C27808 PAND2X1_793/Y POR2X1_767/CTRL 0.01fF
C27809 POR2X1_617/Y PAND2X1_621/Y 0.01fF
C27810 PAND2X1_48/B POR2X1_326/A 0.01fF
C27811 POR2X1_334/Y POR2X1_740/Y 0.10fF
C27812 POR2X1_55/Y PAND2X1_357/CTRL 0.01fF
C27813 PAND2X1_266/a_76_28# POR2X1_262/Y 0.05fF
C27814 POR2X1_257/A PAND2X1_717/A 21.06fF
C27815 POR2X1_41/B POR2X1_7/Y 0.03fF
C27816 PAND2X1_390/O PAND2X1_853/B 0.01fF
C27817 PAND2X1_385/CTRL PAND2X1_48/A 0.01fF
C27818 POR2X1_625/O POR2X1_39/B 0.05fF
C27819 PAND2X1_187/O POR2X1_319/Y 0.08fF
C27820 POR2X1_62/Y PAND2X1_341/CTRL 0.01fF
C27821 POR2X1_541/CTRL POR2X1_456/B 0.01fF
C27822 POR2X1_330/Y POR2X1_717/B 0.05fF
C27823 POR2X1_508/B POR2X1_776/B 0.03fF
C27824 PAND2X1_31/O D_INPUT_7 0.04fF
C27825 POR2X1_532/A POR2X1_260/A 3.71fF
C27826 POR2X1_57/A PAND2X1_714/Y 0.07fF
C27827 PAND2X1_484/CTRL2 PAND2X1_69/A 0.03fF
C27828 POR2X1_119/Y PAND2X1_466/CTRL 0.01fF
C27829 PAND2X1_96/B PAND2X1_184/a_56_28# 0.00fF
C27830 POR2X1_416/B PAND2X1_787/Y 0.01fF
C27831 POR2X1_333/Y PAND2X1_32/B 0.03fF
C27832 PAND2X1_228/O POR2X1_7/Y 0.02fF
C27833 POR2X1_313/Y PAND2X1_213/Y 0.06fF
C27834 POR2X1_68/A POR2X1_737/A 0.05fF
C27835 POR2X1_87/B POR2X1_94/A 0.04fF
C27836 PAND2X1_635/Y POR2X1_32/A 0.17fF
C27837 PAND2X1_569/B PAND2X1_374/CTRL -0.01fF
C27838 PAND2X1_6/Y POR2X1_62/Y 0.03fF
C27839 POR2X1_661/A PAND2X1_58/A 0.17fF
C27840 POR2X1_48/A POR2X1_600/CTRL2 0.00fF
C27841 POR2X1_739/a_76_344# POR2X1_444/Y 0.01fF
C27842 POR2X1_730/Y POR2X1_727/CTRL2 0.01fF
C27843 POR2X1_532/A POR2X1_363/A 0.07fF
C27844 POR2X1_557/A PAND2X1_63/B 0.16fF
C27845 POR2X1_499/A POR2X1_624/Y 0.00fF
C27846 POR2X1_23/Y POR2X1_441/a_76_344# 0.01fF
C27847 POR2X1_316/Y POR2X1_293/Y 0.07fF
C27848 PAND2X1_23/Y PAND2X1_122/O 0.12fF
C27849 POR2X1_16/A PAND2X1_489/CTRL2 0.02fF
C27850 POR2X1_389/A POR2X1_774/A 0.07fF
C27851 POR2X1_382/Y POR2X1_384/Y 0.00fF
C27852 PAND2X1_850/Y POR2X1_45/Y 0.07fF
C27853 PAND2X1_643/a_16_344# PAND2X1_643/A 0.01fF
C27854 POR2X1_741/O POR2X1_741/Y 0.02fF
C27855 POR2X1_416/B PAND2X1_668/CTRL 0.00fF
C27856 PAND2X1_94/A INPUT_1 1.29fF
C27857 POR2X1_16/A PAND2X1_100/CTRL 0.00fF
C27858 D_INPUT_3 POR2X1_62/Y 2.12fF
C27859 POR2X1_348/O POR2X1_334/Y 0.03fF
C27860 PAND2X1_830/O PAND2X1_348/A 0.04fF
C27861 POR2X1_407/Y PAND2X1_328/a_16_344# 0.01fF
C27862 PAND2X1_539/Y PAND2X1_802/B 0.01fF
C27863 PAND2X1_119/a_56_28# POR2X1_294/A 0.00fF
C27864 POR2X1_145/O POR2X1_77/Y 0.05fF
C27865 POR2X1_76/A POR2X1_624/Y -0.03fF
C27866 PAND2X1_804/B POR2X1_173/O 0.06fF
C27867 POR2X1_180/CTRL POR2X1_180/A 0.01fF
C27868 POR2X1_188/CTRL POR2X1_188/Y 0.02fF
C27869 POR2X1_57/A PAND2X1_865/Y 0.07fF
C27870 POR2X1_205/A POR2X1_4/Y 0.22fF
C27871 POR2X1_567/A POR2X1_318/A 0.10fF
C27872 POR2X1_416/B POR2X1_745/CTRL2 -0.00fF
C27873 POR2X1_452/Y POR2X1_809/CTRL 0.01fF
C27874 PAND2X1_220/O POR2X1_77/Y 0.17fF
C27875 POR2X1_387/Y PAND2X1_506/Y 0.07fF
C27876 POR2X1_385/Y PAND2X1_843/Y 0.05fF
C27877 PAND2X1_835/O POR2X1_77/Y 0.15fF
C27878 POR2X1_823/CTRL2 POR2X1_77/Y -0.00fF
C27879 POR2X1_567/B POR2X1_446/A 0.25fF
C27880 POR2X1_16/A PAND2X1_123/Y 0.04fF
C27881 POR2X1_566/B POR2X1_192/B 0.28fF
C27882 POR2X1_602/B POR2X1_648/Y 0.03fF
C27883 PAND2X1_450/O POR2X1_158/Y 0.00fF
C27884 PAND2X1_621/CTRL POR2X1_617/Y 0.01fF
C27885 POR2X1_750/Y POR2X1_294/A 0.22fF
C27886 POR2X1_54/Y POR2X1_37/Y 0.12fF
C27887 PAND2X1_493/CTRL2 POR2X1_394/A 0.05fF
C27888 POR2X1_394/A PAND2X1_708/CTRL2 0.01fF
C27889 POR2X1_49/Y PAND2X1_717/A 0.07fF
C27890 POR2X1_220/CTRL2 POR2X1_220/B 0.03fF
C27891 POR2X1_146/CTRL2 PAND2X1_797/Y 0.01fF
C27892 POR2X1_669/B PAND2X1_750/CTRL 0.01fF
C27893 POR2X1_260/B POR2X1_818/Y 0.03fF
C27894 POR2X1_169/CTRL2 POR2X1_191/Y 0.13fF
C27895 POR2X1_20/B PAND2X1_573/B 0.02fF
C27896 POR2X1_116/A POR2X1_474/CTRL 0.00fF
C27897 PAND2X1_632/a_76_28# PAND2X1_508/Y 0.04fF
C27898 PAND2X1_482/CTRL POR2X1_186/B 0.01fF
C27899 POR2X1_333/a_16_28# POR2X1_192/B 0.04fF
C27900 PAND2X1_39/B POR2X1_287/CTRL 0.01fF
C27901 POR2X1_677/Y PAND2X1_804/B 0.00fF
C27902 POR2X1_567/B POR2X1_446/a_16_28# 0.11fF
C27903 POR2X1_593/a_16_28# POR2X1_449/A 0.03fF
C27904 INPUT_3 POR2X1_14/Y 0.17fF
C27905 PAND2X1_39/B POR2X1_121/B 0.13fF
C27906 POR2X1_383/A POR2X1_343/O 0.02fF
C27907 POR2X1_16/CTRL POR2X1_42/Y 0.01fF
C27908 PAND2X1_404/Y POR2X1_32/A 0.15fF
C27909 POR2X1_294/A POR2X1_398/CTRL 0.01fF
C27910 POR2X1_859/CTRL POR2X1_734/A 0.03fF
C27911 POR2X1_327/Y POR2X1_188/Y 0.06fF
C27912 PAND2X1_20/A POR2X1_446/B 0.04fF
C27913 POR2X1_48/A POR2X1_484/CTRL 0.00fF
C27914 POR2X1_612/Y POR2X1_414/CTRL 0.08fF
C27915 POR2X1_847/O POR2X1_5/Y 0.07fF
C27916 PAND2X1_849/CTRL POR2X1_20/B 0.02fF
C27917 POR2X1_260/B POR2X1_267/A 0.03fF
C27918 PAND2X1_274/O PAND2X1_717/A 0.07fF
C27919 POR2X1_65/A POR2X1_744/Y 0.01fF
C27920 PAND2X1_497/CTRL PAND2X1_58/A 0.01fF
C27921 POR2X1_83/Y POR2X1_62/Y 0.02fF
C27922 POR2X1_74/Y POR2X1_75/Y 0.13fF
C27923 POR2X1_502/A PAND2X1_53/CTRL 0.06fF
C27924 POR2X1_447/B POR2X1_294/A 0.09fF
C27925 PAND2X1_403/Y POR2X1_20/B 0.06fF
C27926 POR2X1_508/B POR2X1_192/B 0.03fF
C27927 PAND2X1_717/A PAND2X1_553/B 0.03fF
C27928 POR2X1_667/O POR2X1_293/Y 0.08fF
C27929 POR2X1_657/CTRL POR2X1_218/Y 0.03fF
C27930 POR2X1_54/Y POR2X1_615/O 0.01fF
C27931 POR2X1_313/Y POR2X1_416/B 0.03fF
C27932 PAND2X1_106/a_16_344# PAND2X1_72/A 0.02fF
C27933 POR2X1_329/A POR2X1_494/Y 0.03fF
C27934 POR2X1_808/A POR2X1_260/B 0.03fF
C27935 POR2X1_54/Y PAND2X1_395/O 0.04fF
C27936 POR2X1_814/B POR2X1_446/B 0.03fF
C27937 POR2X1_9/Y POR2X1_790/A 0.07fF
C27938 POR2X1_852/B POR2X1_629/CTRL2 0.06fF
C27939 POR2X1_23/Y PAND2X1_76/O 0.01fF
C27940 PAND2X1_717/A PAND2X1_303/O 0.03fF
C27941 POR2X1_814/B POR2X1_240/O 0.02fF
C27942 POR2X1_409/B POR2X1_667/A 0.03fF
C27943 POR2X1_286/a_16_28# POR2X1_285/Y 0.04fF
C27944 PAND2X1_206/B POR2X1_42/Y 0.10fF
C27945 POR2X1_133/CTRL POR2X1_411/B 0.00fF
C27946 POR2X1_558/B POR2X1_474/a_16_28# 0.03fF
C27947 POR2X1_852/a_76_344# POR2X1_776/A 0.01fF
C27948 POR2X1_458/Y POR2X1_513/Y 0.15fF
C27949 PAND2X1_9/Y PAND2X1_673/Y 0.03fF
C27950 D_INPUT_0 POR2X1_750/A 0.01fF
C27951 POR2X1_805/Y POR2X1_121/B 0.01fF
C27952 POR2X1_446/B POR2X1_325/A 0.03fF
C27953 POR2X1_811/B POR2X1_590/A 0.01fF
C27954 POR2X1_776/A POR2X1_192/Y 0.03fF
C27955 POR2X1_48/A PAND2X1_541/O 0.04fF
C27956 POR2X1_416/B PAND2X1_708/O 0.01fF
C27957 PAND2X1_308/B PAND2X1_796/B 0.25fF
C27958 PAND2X1_20/A POR2X1_121/B 0.03fF
C27959 PAND2X1_472/B INPUT_3 0.10fF
C27960 PAND2X1_279/CTRL PAND2X1_58/A 0.00fF
C27961 PAND2X1_659/B PAND2X1_203/a_76_28# 0.02fF
C27962 POR2X1_294/A PAND2X1_122/m4_208_n4# 0.06fF
C27963 POR2X1_754/Y POR2X1_750/B 0.77fF
C27964 POR2X1_856/B POR2X1_439/Y 0.45fF
C27965 POR2X1_60/A PAND2X1_786/CTRL2 0.01fF
C27966 PAND2X1_838/B POR2X1_46/Y 0.00fF
C27967 POR2X1_837/B PAND2X1_60/B 0.00fF
C27968 POR2X1_69/CTRL PAND2X1_58/A 0.11fF
C27969 POR2X1_56/CTRL2 POR2X1_423/Y 0.03fF
C27970 POR2X1_41/B POR2X1_257/A 1.77fF
C27971 POR2X1_117/O POR2X1_409/B 0.01fF
C27972 PAND2X1_431/CTRL POR2X1_480/A 0.06fF
C27973 POR2X1_718/A POR2X1_66/A 0.03fF
C27974 POR2X1_13/A PAND2X1_340/B 0.00fF
C27975 POR2X1_23/Y PAND2X1_473/B 0.03fF
C27976 POR2X1_49/Y PAND2X1_623/O 0.01fF
C27977 POR2X1_814/A POR2X1_784/O 0.04fF
C27978 POR2X1_62/Y PAND2X1_52/B 0.05fF
C27979 POR2X1_634/A POR2X1_634/CTRL 0.01fF
C27980 PAND2X1_9/Y PAND2X1_55/Y 0.07fF
C27981 INPUT_3 POR2X1_55/Y 0.05fF
C27982 POR2X1_15/CTRL2 PAND2X1_206/B 0.00fF
C27983 PAND2X1_68/O POR2X1_5/Y 0.11fF
C27984 POR2X1_83/B PAND2X1_390/Y 0.03fF
C27985 POR2X1_106/CTRL2 POR2X1_106/Y 0.01fF
C27986 PAND2X1_219/A PAND2X1_733/CTRL2 0.03fF
C27987 POR2X1_130/A PAND2X1_591/CTRL2 0.01fF
C27988 PAND2X1_404/Y PAND2X1_35/Y 0.03fF
C27989 PAND2X1_798/B POR2X1_411/B 0.03fF
C27990 PAND2X1_23/Y PAND2X1_826/CTRL2 0.01fF
C27991 POR2X1_156/CTRL POR2X1_728/A 0.00fF
C27992 POR2X1_590/A PAND2X1_525/O 0.04fF
C27993 POR2X1_37/Y PAND2X1_501/B 0.01fF
C27994 POR2X1_814/B POR2X1_121/B 0.03fF
C27995 POR2X1_19/O D_INPUT_1 0.01fF
C27996 POR2X1_670/CTRL POR2X1_102/Y 0.00fF
C27997 PAND2X1_487/CTRL2 POR2X1_294/B 0.03fF
C27998 POR2X1_709/A PAND2X1_411/CTRL2 0.00fF
C27999 POR2X1_102/Y PAND2X1_562/B 0.27fF
C28000 POR2X1_68/A PAND2X1_761/CTRL 0.03fF
C28001 PAND2X1_206/B PAND2X1_99/Y 0.01fF
C28002 PAND2X1_404/Y PAND2X1_197/CTRL2 0.01fF
C28003 PAND2X1_658/A POR2X1_415/A 0.34fF
C28004 PAND2X1_56/Y PAND2X1_39/B 0.03fF
C28005 POR2X1_699/CTRL POR2X1_7/B 0.01fF
C28006 POR2X1_856/B POR2X1_192/Y 0.04fF
C28007 PAND2X1_55/Y PAND2X1_67/a_16_344# 0.01fF
C28008 POR2X1_688/m4_208_n4# PAND2X1_32/B 0.15fF
C28009 POR2X1_83/B POR2X1_697/CTRL 0.01fF
C28010 PAND2X1_577/Y VDD 0.14fF
C28011 POR2X1_20/B PAND2X1_341/A 0.03fF
C28012 POR2X1_121/B POR2X1_325/A 0.03fF
C28013 POR2X1_29/A INPUT_0 0.41fF
C28014 POR2X1_174/A VDD 0.80fF
C28015 POR2X1_609/Y POR2X1_234/Y 0.00fF
C28016 PAND2X1_72/A PAND2X1_179/O 0.08fF
C28017 POR2X1_257/A POR2X1_256/Y 0.01fF
C28018 PAND2X1_474/Y POR2X1_102/Y 0.00fF
C28019 POR2X1_20/B POR2X1_93/A 1.07fF
C28020 POR2X1_461/a_16_28# POR2X1_461/A 0.05fF
C28021 POR2X1_498/a_16_28# D_INPUT_0 0.01fF
C28022 POR2X1_20/B POR2X1_91/Y 0.06fF
C28023 POR2X1_814/A POR2X1_456/B 0.03fF
C28024 PAND2X1_459/a_16_344# POR2X1_376/Y 0.02fF
C28025 POR2X1_201/a_16_28# PAND2X1_65/Y 0.02fF
C28026 POR2X1_65/A PAND2X1_61/Y 0.03fF
C28027 POR2X1_375/Y VDD 0.28fF
C28028 POR2X1_610/Y POR2X1_532/A 0.03fF
C28029 POR2X1_355/B POR2X1_78/A 0.06fF
C28030 POR2X1_13/A POR2X1_102/Y 2.32fF
C28031 POR2X1_12/A POR2X1_587/m4_208_n4# 0.12fF
C28032 POR2X1_39/CTRL2 POR2X1_236/Y 0.09fF
C28033 POR2X1_67/A POR2X1_7/B 0.02fF
C28034 POR2X1_810/CTRL POR2X1_636/B 0.01fF
C28035 POR2X1_376/B POR2X1_743/CTRL2 0.00fF
C28036 POR2X1_60/A PAND2X1_735/Y 0.07fF
C28037 POR2X1_52/A POR2X1_422/Y 4.05fF
C28038 PAND2X1_824/B POR2X1_630/B 0.01fF
C28039 POR2X1_193/A POR2X1_296/B 0.03fF
C28040 PAND2X1_796/B POR2X1_239/Y 0.02fF
C28041 POR2X1_579/Y POR2X1_296/B 0.09fF
C28042 POR2X1_505/Y VDD 0.01fF
C28043 POR2X1_54/Y PAND2X1_521/O 0.07fF
C28044 POR2X1_660/CTRL2 PAND2X1_55/Y 0.00fF
C28045 POR2X1_65/A POR2X1_760/CTRL 0.01fF
C28046 POR2X1_41/B POR2X1_142/O 0.05fF
C28047 POR2X1_728/O POR2X1_330/Y 0.03fF
C28048 PAND2X1_640/B PAND2X1_642/B 3.01fF
C28049 POR2X1_66/A POR2X1_204/O 0.05fF
C28050 PAND2X1_65/B POR2X1_448/B 0.03fF
C28051 PAND2X1_404/Y PAND2X1_844/B 0.03fF
C28052 POR2X1_54/Y POR2X1_408/Y 0.10fF
C28053 POR2X1_13/A PAND2X1_436/A 0.00fF
C28054 POR2X1_572/B POR2X1_296/B 0.03fF
C28055 POR2X1_333/A POR2X1_356/A 0.10fF
C28056 PAND2X1_55/Y PAND2X1_15/O 0.03fF
C28057 POR2X1_383/A PAND2X1_39/B 18.58fF
C28058 PAND2X1_217/B POR2X1_498/CTRL2 0.05fF
C28059 POR2X1_730/Y POR2X1_864/A 0.03fF
C28060 PAND2X1_691/Y POR2X1_411/B 0.03fF
C28061 POR2X1_860/A VDD 0.29fF
C28062 POR2X1_686/A VDD 0.15fF
C28063 POR2X1_685/A POR2X1_452/Y 0.02fF
C28064 PAND2X1_859/B POR2X1_60/A 0.03fF
C28065 POR2X1_586/Y POR2X1_790/B 0.01fF
C28066 POR2X1_60/A PAND2X1_493/Y 0.01fF
C28067 PAND2X1_784/A POR2X1_293/Y 0.02fF
C28068 POR2X1_829/A PAND2X1_733/A 0.03fF
C28069 POR2X1_855/B POR2X1_803/a_76_344# 0.00fF
C28070 PAND2X1_714/CTRL2 PAND2X1_731/B 0.01fF
C28071 PAND2X1_795/a_76_28# INPUT_0 0.01fF
C28072 PAND2X1_282/CTRL PAND2X1_69/A 0.02fF
C28073 POR2X1_41/B POR2X1_49/Y 0.45fF
C28074 POR2X1_60/A PAND2X1_174/O 0.05fF
C28075 PAND2X1_56/Y PAND2X1_20/A 0.05fF
C28076 PAND2X1_20/A POR2X1_795/B 0.14fF
C28077 POR2X1_614/A POR2X1_296/B 1.53fF
C28078 POR2X1_341/A POR2X1_332/CTRL2 0.04fF
C28079 PAND2X1_169/Y PAND2X1_724/B 0.00fF
C28080 PAND2X1_3/O D_INPUT_5 0.04fF
C28081 PAND2X1_272/CTRL2 POR2X1_573/A 0.01fF
C28082 POR2X1_287/B POR2X1_121/Y 0.06fF
C28083 POR2X1_118/O POR2X1_32/A 0.02fF
C28084 PAND2X1_65/B PAND2X1_57/B 0.20fF
C28085 PAND2X1_711/B PAND2X1_711/A 0.12fF
C28086 PAND2X1_96/B PAND2X1_594/O 0.02fF
C28087 POR2X1_750/B POR2X1_42/Y 0.07fF
C28088 PAND2X1_4/O D_INPUT_0 0.03fF
C28089 POR2X1_174/A PAND2X1_32/B 0.03fF
C28090 POR2X1_20/B PAND2X1_100/m4_208_n4# 0.15fF
C28091 POR2X1_257/A PAND2X1_308/Y 0.06fF
C28092 POR2X1_38/B POR2X1_296/B 0.10fF
C28093 PAND2X1_473/Y PAND2X1_571/Y 0.87fF
C28094 POR2X1_46/Y PAND2X1_332/a_16_344# 0.03fF
C28095 PAND2X1_467/B POR2X1_694/O 0.01fF
C28096 PAND2X1_412/a_76_28# PAND2X1_57/B 0.06fF
C28097 POR2X1_504/Y POR2X1_628/O 0.01fF
C28098 POR2X1_687/CTRL2 POR2X1_729/Y 0.01fF
C28099 POR2X1_334/B PAND2X1_41/B 3.85fF
C28100 POR2X1_78/B POR2X1_220/Y 0.10fF
C28101 POR2X1_192/Y POR2X1_776/a_16_28# 0.02fF
C28102 PAND2X1_220/Y POR2X1_42/Y 0.03fF
C28103 D_INPUT_2 POR2X1_414/Y 0.01fF
C28104 PAND2X1_643/Y POR2X1_102/Y 0.04fF
C28105 INPUT_0 POR2X1_546/A 0.07fF
C28106 D_INPUT_0 PAND2X1_175/B 0.03fF
C28107 POR2X1_36/B POR2X1_32/A 0.02fF
C28108 POR2X1_68/A POR2X1_302/B 0.03fF
C28109 INPUT_3 POR2X1_376/a_16_28# 0.11fF
C28110 PAND2X1_733/Y POR2X1_7/B 0.01fF
C28111 PAND2X1_464/Y POR2X1_417/Y 0.16fF
C28112 POR2X1_763/A POR2X1_700/O 0.04fF
C28113 POR2X1_763/Y POR2X1_692/Y 0.03fF
C28114 POR2X1_66/A POR2X1_725/Y 0.42fF
C28115 PAND2X1_283/CTRL POR2X1_734/A 0.03fF
C28116 POR2X1_375/Y PAND2X1_32/B 0.00fF
C28117 POR2X1_20/B POR2X1_109/Y 0.03fF
C28118 POR2X1_423/CTRL2 POR2X1_387/Y 0.06fF
C28119 POR2X1_377/CTRL2 POR2X1_5/Y 0.03fF
C28120 POR2X1_792/O PAND2X1_60/B 0.01fF
C28121 PAND2X1_56/Y POR2X1_814/B 0.05fF
C28122 POR2X1_78/B POR2X1_404/Y 0.03fF
C28123 POR2X1_407/A POR2X1_389/Y 0.00fF
C28124 PAND2X1_48/B POR2X1_480/A 0.07fF
C28125 POR2X1_537/Y POR2X1_841/CTRL 0.01fF
C28126 PAND2X1_422/O POR2X1_296/B 0.07fF
C28127 PAND2X1_65/B POR2X1_341/CTRL2 0.00fF
C28128 POR2X1_333/A POR2X1_220/A 0.05fF
C28129 POR2X1_504/Y PAND2X1_6/A 0.03fF
C28130 PAND2X1_39/B PAND2X1_71/Y 0.03fF
C28131 POR2X1_78/B PAND2X1_322/a_76_28# 0.01fF
C28132 POR2X1_566/A PAND2X1_524/O 0.05fF
C28133 POR2X1_106/CTRL2 PAND2X1_114/B 0.03fF
C28134 POR2X1_677/Y PAND2X1_332/Y 0.03fF
C28135 GATE_479 POR2X1_694/CTRL2 0.03fF
C28136 POR2X1_20/B POR2X1_397/O 0.02fF
C28137 POR2X1_614/A PAND2X1_679/CTRL2 0.00fF
C28138 POR2X1_32/A PAND2X1_123/CTRL2 0.01fF
C28139 POR2X1_124/B PAND2X1_41/B 0.00fF
C28140 PAND2X1_168/Y POR2X1_73/Y 0.12fF
C28141 POR2X1_66/B POR2X1_631/A -0.00fF
C28142 POR2X1_96/A POR2X1_329/O 0.18fF
C28143 PAND2X1_362/A PAND2X1_854/A 0.05fF
C28144 PAND2X1_455/Y POR2X1_7/B 0.01fF
C28145 POR2X1_808/A POR2X1_407/Y 0.03fF
C28146 PAND2X1_712/O PAND2X1_707/Y 0.02fF
C28147 PAND2X1_139/CTRL POR2X1_150/Y 0.11fF
C28148 POR2X1_383/A POR2X1_805/Y 0.03fF
C28149 POR2X1_260/B POR2X1_558/Y 0.01fF
C28150 PAND2X1_48/B POR2X1_243/Y 0.07fF
C28151 PAND2X1_739/Y POR2X1_42/Y 0.07fF
C28152 PAND2X1_775/CTRL2 POR2X1_7/B 0.00fF
C28153 PAND2X1_56/Y POR2X1_325/A 0.03fF
C28154 POR2X1_41/B PAND2X1_553/B 0.07fF
C28155 POR2X1_383/A PAND2X1_20/A 0.29fF
C28156 POR2X1_43/B POR2X1_236/Y 0.12fF
C28157 PAND2X1_218/B PAND2X1_853/B 0.05fF
C28158 POR2X1_489/O POR2X1_68/B 0.01fF
C28159 PAND2X1_612/B POR2X1_294/A 0.03fF
C28160 PAND2X1_297/O POR2X1_296/B 0.17fF
C28161 POR2X1_336/O POR2X1_814/B 0.01fF
C28162 PAND2X1_65/B POR2X1_828/A 0.04fF
C28163 PAND2X1_711/CTRL POR2X1_763/A 0.07fF
C28164 PAND2X1_467/B PAND2X1_467/CTRL2 0.01fF
C28165 POR2X1_52/A PAND2X1_465/B 0.36fF
C28166 POR2X1_718/A POR2X1_532/A 0.03fF
C28167 POR2X1_60/A PAND2X1_569/B 0.07fF
C28168 POR2X1_66/A POR2X1_559/A 6.65fF
C28169 POR2X1_108/O PAND2X1_562/B 0.02fF
C28170 PAND2X1_480/B POR2X1_238/Y 0.01fF
C28171 PAND2X1_55/Y POR2X1_445/O 0.01fF
C28172 POR2X1_471/A PAND2X1_179/CTRL 0.01fF
C28173 POR2X1_614/A POR2X1_547/B 0.02fF
C28174 PAND2X1_23/Y POR2X1_360/A 0.02fF
C28175 POR2X1_96/A POR2X1_45/Y 0.03fF
C28176 POR2X1_566/A D_GATE_222 0.10fF
C28177 POR2X1_383/A POR2X1_254/CTRL 0.02fF
C28178 PAND2X1_489/m4_208_n4# PAND2X1_363/m4_208_n4# 0.13fF
C28179 POR2X1_495/CTRL POR2X1_283/A 0.01fF
C28180 POR2X1_3/A POR2X1_763/A 0.29fF
C28181 PAND2X1_773/CTRL VDD -0.00fF
C28182 POR2X1_459/m4_208_n4# PAND2X1_378/m4_208_n4# 0.13fF
C28183 PAND2X1_661/Y POR2X1_72/B 0.03fF
C28184 PAND2X1_48/B PAND2X1_90/A 0.00fF
C28185 POR2X1_38/B POR2X1_236/Y 6.15fF
C28186 POR2X1_355/B POR2X1_510/A 0.03fF
C28187 PAND2X1_3/A PAND2X1_18/B 0.03fF
C28188 POR2X1_750/B PAND2X1_1/O 0.02fF
C28189 POR2X1_669/B PAND2X1_708/CTRL2 0.03fF
C28190 POR2X1_52/A PAND2X1_798/B 0.07fF
C28191 POR2X1_38/B POR2X1_547/B 0.03fF
C28192 POR2X1_43/B POR2X1_81/Y 0.02fF
C28193 POR2X1_549/CTRL POR2X1_383/A 0.03fF
C28194 POR2X1_383/A POR2X1_814/B 0.26fF
C28195 POR2X1_750/B PAND2X1_376/CTRL2 0.01fF
C28196 PAND2X1_76/Y POR2X1_387/Y 0.07fF
C28197 POR2X1_364/A POR2X1_502/A 0.10fF
C28198 PAND2X1_41/B POR2X1_218/O 0.16fF
C28199 POR2X1_225/O POR2X1_129/Y 0.01fF
C28200 INPUT_0 POR2X1_500/Y 0.03fF
C28201 POR2X1_474/a_16_28# POR2X1_362/A 0.05fF
C28202 POR2X1_416/Y POR2X1_232/O 0.01fF
C28203 PAND2X1_340/a_16_344# POR2X1_408/Y 0.04fF
C28204 PAND2X1_592/Y PAND2X1_794/B 0.03fF
C28205 D_GATE_579 D_GATE_741 0.03fF
C28206 POR2X1_619/A VDD 0.06fF
C28207 PAND2X1_675/A POR2X1_55/Y 0.03fF
C28208 POR2X1_669/B PAND2X1_156/A 0.10fF
C28209 POR2X1_188/A PAND2X1_698/O 0.02fF
C28210 POR2X1_71/CTRL POR2X1_60/A 0.01fF
C28211 POR2X1_78/A POR2X1_209/O 0.01fF
C28212 POR2X1_16/A PAND2X1_354/A 0.03fF
C28213 PAND2X1_183/CTRL2 POR2X1_540/A 0.10fF
C28214 PAND2X1_469/B POR2X1_55/Y 0.05fF
C28215 POR2X1_188/A POR2X1_463/Y 3.05fF
C28216 POR2X1_49/Y POR2X1_419/O 0.06fF
C28217 PAND2X1_787/A PAND2X1_151/CTRL2 0.02fF
C28218 POR2X1_65/A POR2X1_291/CTRL2 0.10fF
C28219 POR2X1_257/A POR2X1_77/Y 10.69fF
C28220 POR2X1_37/Y POR2X1_4/Y 1.25fF
C28221 POR2X1_795/CTRL POR2X1_786/Y 0.03fF
C28222 PAND2X1_107/CTRL2 PAND2X1_65/B 0.01fF
C28223 PAND2X1_477/B PAND2X1_241/O 0.15fF
C28224 POR2X1_383/A POR2X1_325/A 0.03fF
C28225 POR2X1_563/O POR2X1_569/A 0.05fF
C28226 POR2X1_572/B POR2X1_267/Y 0.02fF
C28227 PAND2X1_65/B POR2X1_707/Y 1.55fF
C28228 POR2X1_32/A POR2X1_701/O 0.01fF
C28229 POR2X1_840/O POR2X1_307/Y 0.01fF
C28230 PAND2X1_20/A PAND2X1_71/Y 0.03fF
C28231 PAND2X1_58/A POR2X1_737/A 0.03fF
C28232 POR2X1_73/CTRL2 VDD 0.00fF
C28233 POR2X1_356/A POR2X1_788/B 0.08fF
C28234 POR2X1_49/Y PAND2X1_308/Y 0.07fF
C28235 INPUT_1 PAND2X1_721/CTRL 0.00fF
C28236 POR2X1_219/O POR2X1_294/B 0.02fF
C28237 POR2X1_66/B POR2X1_537/m4_208_n4# 0.08fF
C28238 PAND2X1_370/CTRL2 POR2X1_309/Y 0.01fF
C28239 PAND2X1_599/O POR2X1_828/A 0.02fF
C28240 PAND2X1_20/A POR2X1_560/Y 0.01fF
C28241 PAND2X1_23/Y POR2X1_544/CTRL2 0.01fF
C28242 PAND2X1_659/Y PAND2X1_219/A 0.03fF
C28243 POR2X1_141/a_16_28# POR2X1_141/A 0.12fF
C28244 POR2X1_390/B POR2X1_335/CTRL 0.00fF
C28245 POR2X1_251/Y PAND2X1_349/A 0.02fF
C28246 PAND2X1_632/B VDD 0.07fF
C28247 POR2X1_591/CTRL POR2X1_591/Y 0.01fF
C28248 PAND2X1_593/Y VDD 0.17fF
C28249 POR2X1_138/CTRL2 POR2X1_318/A 0.03fF
C28250 D_INPUT_3 POR2X1_119/O 0.02fF
C28251 POR2X1_43/B PAND2X1_858/Y 0.01fF
C28252 POR2X1_383/A POR2X1_513/B 0.09fF
C28253 PAND2X1_6/Y POR2X1_804/A 0.07fF
C28254 PAND2X1_592/Y PAND2X1_842/Y 0.00fF
C28255 PAND2X1_726/O POR2X1_152/Y 0.06fF
C28256 POR2X1_383/A POR2X1_327/O 0.01fF
C28257 PAND2X1_490/O PAND2X1_6/Y 0.17fF
C28258 PAND2X1_422/m4_208_n4# PAND2X1_72/A 0.15fF
C28259 POR2X1_423/Y PAND2X1_716/B 0.03fF
C28260 POR2X1_814/B PAND2X1_71/Y 0.03fF
C28261 POR2X1_313/Y PAND2X1_738/Y 0.05fF
C28262 POR2X1_178/m4_208_n4# PAND2X1_675/A 0.12fF
C28263 POR2X1_141/a_76_344# POR2X1_244/Y 0.01fF
C28264 PAND2X1_724/CTRL2 POR2X1_73/Y 0.01fF
C28265 PAND2X1_551/CTRL PAND2X1_324/Y 0.01fF
C28266 POR2X1_469/a_16_28# POR2X1_468/Y 0.04fF
C28267 POR2X1_532/A POR2X1_713/Y 0.09fF
C28268 POR2X1_78/B PAND2X1_399/CTRL 0.01fF
C28269 PAND2X1_330/a_16_344# POR2X1_385/Y 0.04fF
C28270 POR2X1_135/Y POR2X1_129/Y 0.03fF
C28271 POR2X1_316/Y POR2X1_60/A 0.03fF
C28272 POR2X1_90/Y POR2X1_321/a_16_28# 0.01fF
C28273 POR2X1_45/Y POR2X1_7/A 0.15fF
C28274 POR2X1_608/Y PAND2X1_56/A 0.01fF
C28275 POR2X1_558/B POR2X1_717/B 0.20fF
C28276 PAND2X1_23/Y POR2X1_787/CTRL2 0.01fF
C28277 POR2X1_639/Y POR2X1_407/Y 0.03fF
C28278 POR2X1_510/B POR2X1_510/A 0.01fF
C28279 POR2X1_41/B POR2X1_41/O 0.01fF
C28280 D_GATE_662 PAND2X1_373/CTRL 0.03fF
C28281 POR2X1_179/Y PAND2X1_675/A 0.05fF
C28282 POR2X1_110/Y POR2X1_485/CTRL 0.02fF
C28283 POR2X1_224/a_56_344# POR2X1_394/A 0.00fF
C28284 PAND2X1_440/CTRL2 POR2X1_60/A 0.01fF
C28285 PAND2X1_6/Y PAND2X1_27/CTRL 0.01fF
C28286 POR2X1_16/A PAND2X1_724/B 0.03fF
C28287 POR2X1_515/a_16_28# POR2X1_574/Y 0.02fF
C28288 POR2X1_94/A PAND2X1_379/O 0.09fF
C28289 PAND2X1_82/Y POR2X1_35/Y 0.04fF
C28290 POR2X1_717/O POR2X1_865/B 0.01fF
C28291 POR2X1_762/O VDD 0.00fF
C28292 POR2X1_646/Y PAND2X1_52/B 0.04fF
C28293 POR2X1_425/Y POR2X1_426/Y 0.01fF
C28294 POR2X1_65/A POR2X1_518/O 0.01fF
C28295 PAND2X1_793/Y PAND2X1_853/B 0.03fF
C28296 POR2X1_135/a_16_28# POR2X1_423/Y 0.02fF
C28297 PAND2X1_308/Y PAND2X1_303/O 0.04fF
C28298 POR2X1_66/B POR2X1_736/A 0.01fF
C28299 POR2X1_346/B PAND2X1_625/CTRL 0.00fF
C28300 PAND2X1_351/O POR2X1_153/Y 0.04fF
C28301 INPUT_3 POR2X1_612/A 0.00fF
C28302 POR2X1_96/A PAND2X1_355/O 0.17fF
C28303 PAND2X1_390/Y PAND2X1_841/Y 0.00fF
C28304 PAND2X1_69/A PAND2X1_528/CTRL 0.00fF
C28305 POR2X1_136/m4_208_n4# PAND2X1_702/m4_208_n4# 0.15fF
C28306 PAND2X1_491/CTRL PAND2X1_94/A 0.26fF
C28307 PAND2X1_560/B POR2X1_42/Y 0.11fF
C28308 POR2X1_30/O POR2X1_260/A 0.01fF
C28309 POR2X1_192/Y POR2X1_191/Y 0.05fF
C28310 PAND2X1_697/O POR2X1_260/A 0.01fF
C28311 POR2X1_49/Y POR2X1_77/Y 0.13fF
C28312 POR2X1_614/A POR2X1_543/CTRL 0.01fF
C28313 POR2X1_648/Y PAND2X1_39/B 0.03fF
C28314 POR2X1_404/Y POR2X1_294/A 0.03fF
C28315 POR2X1_785/O POR2X1_191/Y -0.01fF
C28316 POR2X1_562/O POR2X1_339/Y 0.01fF
C28317 POR2X1_140/B POR2X1_574/Y 0.86fF
C28318 POR2X1_616/Y POR2X1_7/B 0.33fF
C28319 PAND2X1_812/A PAND2X1_288/A 0.02fF
C28320 PAND2X1_38/a_16_344# POR2X1_4/Y 0.06fF
C28321 PAND2X1_777/CTRL2 POR2X1_90/Y 0.01fF
C28322 POR2X1_42/Y PAND2X1_538/a_16_344# 0.02fF
C28323 POR2X1_108/Y POR2X1_142/Y -0.00fF
C28324 POR2X1_740/Y POR2X1_726/CTRL2 0.00fF
C28325 POR2X1_712/O POR2X1_707/Y 0.18fF
C28326 INPUT_1 POR2X1_382/Y 0.07fF
C28327 POR2X1_332/Y POR2X1_795/B 0.02fF
C28328 POR2X1_96/A POR2X1_304/CTRL2 0.01fF
C28329 POR2X1_293/Y POR2X1_4/Y 0.03fF
C28330 PAND2X1_149/O PAND2X1_797/Y 0.02fF
C28331 POR2X1_43/Y PAND2X1_195/a_76_28# 0.02fF
C28332 POR2X1_57/A PAND2X1_343/O 0.01fF
C28333 POR2X1_13/A POR2X1_761/A 0.04fF
C28334 PAND2X1_23/Y POR2X1_99/B 0.03fF
C28335 PAND2X1_808/O POR2X1_385/Y 0.04fF
C28336 POR2X1_543/A POR2X1_717/B 0.12fF
C28337 POR2X1_465/CTRL2 POR2X1_454/A 0.04fF
C28338 PAND2X1_172/CTRL POR2X1_854/B 0.10fF
C28339 POR2X1_196/Y POR2X1_334/Y 0.04fF
C28340 POR2X1_532/A POR2X1_559/A 0.19fF
C28341 POR2X1_335/A POR2X1_188/Y 0.00fF
C28342 POR2X1_96/A POR2X1_305/CTRL2 0.02fF
C28343 POR2X1_40/Y POR2X1_321/CTRL2 0.01fF
C28344 PAND2X1_492/CTRL2 PAND2X1_72/A 0.03fF
C28345 POR2X1_567/A POR2X1_341/O 0.24fF
C28346 PAND2X1_683/CTRL PAND2X1_69/A 0.01fF
C28347 POR2X1_240/B POR2X1_98/A 0.08fF
C28348 POR2X1_119/Y PAND2X1_836/CTRL -0.02fF
C28349 POR2X1_52/Y POR2X1_7/Y 0.13fF
C28350 PAND2X1_631/CTRL2 PAND2X1_631/A 0.03fF
C28351 POR2X1_347/CTRL POR2X1_402/A 0.01fF
C28352 POR2X1_416/B POR2X1_57/CTRL2 0.05fF
C28353 POR2X1_186/O POR2X1_725/Y 0.05fF
C28354 POR2X1_832/a_16_28# POR2X1_711/Y 0.01fF
C28355 POR2X1_325/CTRL POR2X1_544/B 0.01fF
C28356 POR2X1_165/Y PAND2X1_168/a_76_28# 0.07fF
C28357 PAND2X1_503/a_76_28# POR2X1_854/B 0.04fF
C28358 PAND2X1_612/B POR2X1_286/B 0.02fF
C28359 PAND2X1_319/B PAND2X1_716/B 0.10fF
C28360 POR2X1_765/Y PAND2X1_569/a_76_28# 0.01fF
C28361 POR2X1_495/Y POR2X1_39/B 0.68fF
C28362 PAND2X1_48/A PAND2X1_60/B 0.26fF
C28363 POR2X1_278/Y PAND2X1_332/Y 0.07fF
C28364 PAND2X1_653/O PAND2X1_652/A 0.04fF
C28365 POR2X1_250/Y POR2X1_487/a_16_28# 0.01fF
C28366 POR2X1_124/B PAND2X1_122/O 0.01fF
C28367 POR2X1_24/Y PAND2X1_35/A 0.01fF
C28368 POR2X1_609/Y POR2X1_412/CTRL2 0.01fF
C28369 POR2X1_110/CTRL POR2X1_7/A 0.03fF
C28370 POR2X1_68/A POR2X1_716/CTRL2 0.15fF
C28371 POR2X1_542/B POR2X1_374/O 0.01fF
C28372 POR2X1_835/B POR2X1_590/A 0.18fF
C28373 POR2X1_327/Y POR2X1_276/Y 0.05fF
C28374 POR2X1_57/A PAND2X1_352/Y 0.04fF
C28375 PAND2X1_20/A POR2X1_648/Y 0.06fF
C28376 PAND2X1_860/A PAND2X1_499/Y 0.03fF
C28377 POR2X1_659/O POR2X1_736/A 0.06fF
C28378 POR2X1_858/B POR2X1_851/O 0.00fF
C28379 POR2X1_567/A POR2X1_540/a_16_28# 0.03fF
C28380 POR2X1_78/B POR2X1_651/Y 0.03fF
C28381 POR2X1_713/O POR2X1_711/Y 0.01fF
C28382 PAND2X1_341/B POR2X1_229/Y 0.17fF
C28383 PAND2X1_661/B POR2X1_761/A 0.01fF
C28384 PAND2X1_643/Y POR2X1_761/A 4.36fF
C28385 POR2X1_462/a_16_28# POR2X1_590/A 0.02fF
C28386 PAND2X1_569/B POR2X1_373/CTRL2 0.01fF
C28387 PAND2X1_472/A POR2X1_416/B 0.01fF
C28388 POR2X1_102/Y POR2X1_412/CTRL 0.00fF
C28389 POR2X1_191/Y POR2X1_568/Y 0.05fF
C28390 POR2X1_540/A POR2X1_181/a_76_344# 0.01fF
C28391 PAND2X1_466/A POR2X1_14/Y 0.01fF
C28392 PAND2X1_467/Y POR2X1_119/Y 0.02fF
C28393 PAND2X1_32/a_16_344# POR2X1_94/A 0.02fF
C28394 PAND2X1_200/B POR2X1_153/Y 0.00fF
C28395 POR2X1_343/Y PAND2X1_69/A 0.03fF
C28396 POR2X1_67/Y POR2X1_391/A 0.25fF
C28397 POR2X1_249/Y POR2X1_188/Y 0.03fF
C28398 POR2X1_678/Y POR2X1_808/O 0.23fF
C28399 PAND2X1_587/CTRL PAND2X1_52/B 0.06fF
C28400 POR2X1_174/B POR2X1_227/B 0.03fF
C28401 POR2X1_38/Y PAND2X1_198/O 0.15fF
C28402 POR2X1_416/B POR2X1_32/Y 0.01fF
C28403 PAND2X1_510/a_76_28# PAND2X1_508/Y 0.01fF
C28404 POR2X1_52/CTRL POR2X1_7/A 0.01fF
C28405 POR2X1_13/A POR2X1_677/Y 0.05fF
C28406 POR2X1_824/O POR2X1_16/A 0.07fF
C28407 POR2X1_768/O POR2X1_113/B 0.03fF
C28408 POR2X1_192/B POR2X1_353/A 0.01fF
C28409 POR2X1_86/Y PAND2X1_341/A 0.03fF
C28410 POR2X1_51/A PAND2X1_635/Y 0.03fF
C28411 PAND2X1_166/O POR2X1_854/B 0.04fF
C28412 POR2X1_13/A POR2X1_9/Y 0.01fF
C28413 PAND2X1_399/CTRL POR2X1_294/A 0.01fF
C28414 PAND2X1_549/B POR2X1_372/CTRL 0.00fF
C28415 POR2X1_66/Y PAND2X1_58/A 0.01fF
C28416 POR2X1_116/A POR2X1_141/Y 0.01fF
C28417 POR2X1_711/Y PAND2X1_305/CTRL 0.08fF
C28418 POR2X1_316/a_16_28# POR2X1_129/Y 0.02fF
C28419 PAND2X1_72/A POR2X1_788/B 0.03fF
C28420 POR2X1_329/A POR2X1_497/Y 0.13fF
C28421 POR2X1_357/CTRL2 POR2X1_191/Y 0.11fF
C28422 PAND2X1_106/CTRL POR2X1_343/Y 0.28fF
C28423 PAND2X1_22/CTRL PAND2X1_11/Y 0.01fF
C28424 PAND2X1_469/a_76_28# POR2X1_32/A 0.01fF
C28425 POR2X1_54/Y POR2X1_634/A 0.03fF
C28426 PAND2X1_58/A POR2X1_606/CTRL 0.01fF
C28427 POR2X1_409/B D_INPUT_0 0.03fF
C28428 POR2X1_357/O POR2X1_357/B 0.00fF
C28429 POR2X1_327/Y POR2X1_741/CTRL2 0.02fF
C28430 POR2X1_416/B POR2X1_527/Y 0.03fF
C28431 POR2X1_814/A PAND2X1_57/B 0.25fF
C28432 PAND2X1_163/CTRL PAND2X1_72/A 0.01fF
C28433 POR2X1_320/Y POR2X1_321/Y 0.07fF
C28434 POR2X1_676/CTRL POR2X1_750/B 0.01fF
C28435 POR2X1_353/Y POR2X1_443/O 0.03fF
C28436 POR2X1_416/B PAND2X1_196/O 0.02fF
C28437 POR2X1_841/B POR2X1_806/O 0.10fF
C28438 POR2X1_535/O POR2X1_788/B 0.00fF
C28439 POR2X1_648/Y POR2X1_513/B 0.10fF
C28440 POR2X1_648/CTRL2 POR2X1_718/A 0.02fF
C28441 POR2X1_411/B POR2X1_666/A 1.04fF
C28442 PAND2X1_340/B POR2X1_820/A 0.01fF
C28443 PAND2X1_63/a_76_28# POR2X1_296/B 0.01fF
C28444 POR2X1_329/O POR2X1_760/A 0.02fF
C28445 POR2X1_811/B POR2X1_66/A 0.05fF
C28446 PAND2X1_93/B POR2X1_269/Y 0.01fF
C28447 POR2X1_590/A POR2X1_296/B 2.60fF
C28448 POR2X1_102/Y PAND2X1_722/O 0.03fF
C28449 POR2X1_814/A POR2X1_193/O 0.07fF
C28450 PAND2X1_2/CTRL D_INPUT_4 0.01fF
C28451 PAND2X1_175/B POR2X1_173/Y 0.08fF
C28452 POR2X1_462/B POR2X1_848/CTRL2 0.01fF
C28453 PAND2X1_39/B INPUT_0 0.02fF
C28454 PAND2X1_340/B POR2X1_381/a_76_344# 0.00fF
C28455 POR2X1_54/Y POR2X1_130/A 0.24fF
C28456 PAND2X1_472/A PAND2X1_608/CTRL 0.04fF
C28457 POR2X1_446/B VDD 0.87fF
C28458 POR2X1_116/A POR2X1_404/Y 0.03fF
C28459 POR2X1_66/A PAND2X1_387/CTRL2 0.01fF
C28460 POR2X1_760/A POR2X1_45/Y 0.07fF
C28461 POR2X1_456/B PAND2X1_125/CTRL 0.00fF
C28462 POR2X1_502/A POR2X1_818/a_16_28# 0.02fF
C28463 POR2X1_792/CTRL PAND2X1_41/B 0.03fF
C28464 POR2X1_333/Y POR2X1_568/A 0.03fF
C28465 POR2X1_814/B PAND2X1_15/CTRL2 0.03fF
C28466 D_GATE_662 POR2X1_444/CTRL2 0.12fF
C28467 POR2X1_866/A PAND2X1_511/CTRL 0.04fF
C28468 POR2X1_302/B PAND2X1_58/A 0.03fF
C28469 PAND2X1_307/a_16_344# POR2X1_102/Y 0.02fF
C28470 POR2X1_68/A POR2X1_864/A 0.11fF
C28471 POR2X1_272/Y D_INPUT_0 0.03fF
C28472 PAND2X1_319/a_76_28# POR2X1_48/A 0.02fF
C28473 PAND2X1_790/a_16_344# POR2X1_7/B 0.02fF
C28474 POR2X1_32/A PAND2X1_736/O 0.01fF
C28475 POR2X1_257/A POR2X1_426/CTRL2 0.03fF
C28476 PAND2X1_473/Y PAND2X1_571/CTRL 0.01fF
C28477 PAND2X1_73/Y POR2X1_285/CTRL 0.07fF
C28478 POR2X1_848/A POR2X1_790/O 0.04fF
C28479 POR2X1_67/Y POR2X1_391/CTRL 0.00fF
C28480 PAND2X1_48/B PAND2X1_487/O 0.17fF
C28481 POR2X1_760/A PAND2X1_799/CTRL2 0.01fF
C28482 POR2X1_78/Y PAND2X1_767/a_16_344# 0.02fF
C28483 PAND2X1_793/Y POR2X1_23/Y 0.03fF
C28484 PAND2X1_48/B PAND2X1_251/CTRL2 0.01fF
C28485 POR2X1_446/B POR2X1_741/Y 0.03fF
C28486 POR2X1_159/CTRL2 POR2X1_376/B 0.03fF
C28487 POR2X1_605/CTRL PAND2X1_90/Y 0.06fF
C28488 POR2X1_376/B PAND2X1_502/a_76_28# 0.04fF
C28489 POR2X1_20/B POR2X1_299/CTRL 0.03fF
C28490 POR2X1_590/A POR2X1_547/B 0.03fF
C28491 PAND2X1_841/B POR2X1_23/Y 0.03fF
C28492 PAND2X1_809/CTRL2 PAND2X1_539/Y 0.01fF
C28493 POR2X1_226/Y POR2X1_40/Y 0.03fF
C28494 POR2X1_590/A POR2X1_214/CTRL2 0.00fF
C28495 PAND2X1_37/O PAND2X1_8/Y 0.03fF
C28496 POR2X1_66/A PAND2X1_176/CTRL 0.01fF
C28497 POR2X1_254/A POR2X1_254/a_16_28# 0.04fF
C28498 PAND2X1_557/A PAND2X1_740/a_16_344# 0.02fF
C28499 POR2X1_121/B VDD 1.32fF
C28500 POR2X1_651/Y POR2X1_294/A 0.07fF
C28501 POR2X1_624/Y PAND2X1_69/A 0.03fF
C28502 POR2X1_82/a_16_28# POR2X1_29/A 0.04fF
C28503 POR2X1_677/a_76_344# PAND2X1_390/Y 0.00fF
C28504 POR2X1_66/Y PAND2X1_96/B 0.04fF
C28505 PAND2X1_200/Y VDD 0.13fF
C28506 PAND2X1_20/A INPUT_0 0.39fF
C28507 POR2X1_20/B PAND2X1_338/B 0.03fF
C28508 POR2X1_376/B PAND2X1_185/O 0.12fF
C28509 POR2X1_270/Y POR2X1_659/O 0.01fF
C28510 POR2X1_630/A VDD 0.11fF
C28511 PAND2X1_39/B POR2X1_780/A 0.02fF
C28512 POR2X1_96/A POR2X1_420/Y 0.01fF
C28513 PAND2X1_45/CTRL POR2X1_260/A 0.00fF
C28514 POR2X1_814/A POR2X1_259/B 0.02fF
C28515 PAND2X1_39/B PAND2X1_393/CTRL2 0.01fF
C28516 D_INPUT_0 POR2X1_501/CTRL 0.01fF
C28517 PAND2X1_808/Y PAND2X1_811/A 0.01fF
C28518 POR2X1_225/O POR2X1_293/Y 0.01fF
C28519 POR2X1_188/A POR2X1_285/a_56_344# 0.00fF
C28520 POR2X1_68/A POR2X1_855/O 0.01fF
C28521 PAND2X1_93/B POR2X1_513/Y 0.03fF
C28522 POR2X1_840/B POR2X1_260/B 0.07fF
C28523 POR2X1_366/CTRL POR2X1_116/A 0.00fF
C28524 POR2X1_409/B POR2X1_277/a_16_28# 0.02fF
C28525 POR2X1_154/CTRL2 POR2X1_750/B 0.11fF
C28526 POR2X1_83/B PAND2X1_592/Y 0.03fF
C28527 PAND2X1_824/B POR2X1_240/A 0.01fF
C28528 POR2X1_70/CTRL POR2X1_40/Y 0.01fF
C28529 PAND2X1_93/B POR2X1_219/B 0.15fF
C28530 POR2X1_74/CTRL2 POR2X1_20/B 0.01fF
C28531 PAND2X1_94/A POR2X1_556/A 0.05fF
C28532 PAND2X1_58/A POR2X1_756/CTRL 0.01fF
C28533 POR2X1_118/Y POR2X1_73/Y 0.03fF
C28534 POR2X1_498/CTRL POR2X1_72/B 0.01fF
C28535 POR2X1_37/Y POR2X1_816/A 0.03fF
C28536 PAND2X1_721/CTRL2 VDD 0.00fF
C28537 POR2X1_52/A PAND2X1_195/O 0.01fF
C28538 PAND2X1_445/CTRL POR2X1_102/Y 0.01fF
C28539 POR2X1_307/Y POR2X1_330/Y 0.05fF
C28540 POR2X1_814/B INPUT_0 0.21fF
C28541 POR2X1_128/O POR2X1_750/B 0.34fF
C28542 POR2X1_37/Y D_INPUT_1 0.01fF
C28543 POR2X1_811/CTRL2 POR2X1_532/A 0.03fF
C28544 PAND2X1_115/Y POR2X1_40/Y 1.50fF
C28545 POR2X1_241/B D_GATE_222 0.03fF
C28546 PAND2X1_93/B POR2X1_205/A 0.07fF
C28547 POR2X1_669/B POR2X1_396/O 0.07fF
C28548 POR2X1_471/A PAND2X1_313/CTRL2 0.01fF
C28549 POR2X1_48/A PAND2X1_553/O 0.04fF
C28550 PAND2X1_118/a_16_344# PAND2X1_73/Y 0.02fF
C28551 POR2X1_65/A POR2X1_693/CTRL 0.01fF
C28552 PAND2X1_217/B POR2X1_275/CTRL 0.01fF
C28553 PAND2X1_643/O POR2X1_102/Y 0.01fF
C28554 POR2X1_65/A POR2X1_46/Y 0.06fF
C28555 POR2X1_41/B POR2X1_278/CTRL 0.00fF
C28556 POR2X1_150/Y POR2X1_394/A 0.03fF
C28557 POR2X1_502/A POR2X1_461/a_16_28# 0.01fF
C28558 PAND2X1_280/CTRL2 PAND2X1_90/Y 0.12fF
C28559 POR2X1_840/CTRL POR2X1_660/Y 0.01fF
C28560 POR2X1_83/B PAND2X1_370/CTRL 0.03fF
C28561 POR2X1_186/Y POR2X1_579/Y 0.03fF
C28562 POR2X1_62/Y POR2X1_623/Y 0.01fF
C28563 PAND2X1_659/B PAND2X1_735/CTRL2 0.00fF
C28564 PAND2X1_93/B POR2X1_366/A 0.00fF
C28565 POR2X1_654/B POR2X1_294/B 0.10fF
C28566 POR2X1_404/B POR2X1_403/Y 0.01fF
C28567 POR2X1_477/A PAND2X1_41/B 0.03fF
C28568 POR2X1_614/A POR2X1_864/CTRL2 0.01fF
C28569 POR2X1_66/B PAND2X1_6/A 0.05fF
C28570 POR2X1_121/B PAND2X1_32/B 7.63fF
C28571 POR2X1_278/Y PAND2X1_474/Y 0.05fF
C28572 POR2X1_801/B PAND2X1_583/a_76_28# 0.04fF
C28573 POR2X1_254/O POR2X1_222/Y 0.04fF
C28574 POR2X1_448/CTRL POR2X1_788/B 0.01fF
C28575 PAND2X1_39/B POR2X1_398/CTRL2 0.05fF
C28576 PAND2X1_859/A POR2X1_382/O 0.01fF
C28577 PAND2X1_6/Y POR2X1_794/B 0.03fF
C28578 POR2X1_368/O POR2X1_13/A 0.17fF
C28579 PAND2X1_758/CTRL2 POR2X1_236/Y 0.10fF
C28580 POR2X1_811/B POR2X1_532/A 0.03fF
C28581 POR2X1_278/Y POR2X1_13/A 0.01fF
C28582 POR2X1_108/CTRL POR2X1_60/A 0.07fF
C28583 PAND2X1_96/B POR2X1_675/O 0.01fF
C28584 PAND2X1_351/CTRL VDD 0.00fF
C28585 PAND2X1_90/A PAND2X1_667/CTRL 0.00fF
C28586 POR2X1_818/CTRL2 POR2X1_294/A 0.01fF
C28587 PAND2X1_191/Y VDD 0.15fF
C28588 POR2X1_614/A POR2X1_186/Y 0.15fF
C28589 POR2X1_467/Y POR2X1_535/A 0.01fF
C28590 PAND2X1_84/Y POR2X1_494/Y 0.02fF
C28591 POR2X1_660/Y POR2X1_725/Y 0.04fF
C28592 POR2X1_641/O POR2X1_318/A 0.10fF
C28593 POR2X1_13/A POR2X1_829/A 0.04fF
C28594 PAND2X1_758/O VDD 0.00fF
C28595 PAND2X1_615/CTRL2 POR2X1_94/A 0.16fF
C28596 POR2X1_840/B PAND2X1_74/a_76_28# 0.03fF
C28597 PAND2X1_445/Y POR2X1_7/B 0.00fF
C28598 POR2X1_498/a_16_28# PAND2X1_735/Y 0.04fF
C28599 POR2X1_344/CTRL2 POR2X1_205/A 0.03fF
C28600 POR2X1_43/B POR2X1_58/CTRL 0.01fF
C28601 POR2X1_376/Y PAND2X1_6/A 0.81fF
C28602 POR2X1_623/A POR2X1_296/B 0.07fF
C28603 POR2X1_614/A PAND2X1_263/CTRL2 0.00fF
C28604 POR2X1_590/a_56_344# POR2X1_296/B 0.03fF
C28605 POR2X1_483/O POR2X1_193/A 0.01fF
C28606 POR2X1_214/CTRL2 POR2X1_214/B 0.01fF
C28607 POR2X1_215/CTRL POR2X1_740/Y 0.01fF
C28608 PAND2X1_392/B POR2X1_90/Y 0.03fF
C28609 POR2X1_51/B PAND2X1_11/Y 0.10fF
C28610 POR2X1_433/a_56_344# PAND2X1_349/A 0.00fF
C28611 POR2X1_7/B PAND2X1_335/CTRL2 0.00fF
C28612 POR2X1_260/Y PAND2X1_57/B 0.03fF
C28613 PAND2X1_803/Y POR2X1_40/Y 0.02fF
C28614 POR2X1_683/Y POR2X1_236/Y 0.02fF
C28615 PAND2X1_830/CTRL POR2X1_60/A 0.17fF
C28616 POR2X1_795/B VDD 0.03fF
C28617 PAND2X1_56/Y VDD 5.30fF
C28618 POR2X1_137/Y POR2X1_777/B 0.05fF
C28619 POR2X1_732/CTRL VDD 0.00fF
C28620 POR2X1_83/A VDD 0.24fF
C28621 PAND2X1_114/Y PAND2X1_553/B 0.07fF
C28622 POR2X1_76/Y POR2X1_740/Y 0.03fF
C28623 POR2X1_55/O POR2X1_673/Y 0.01fF
C28624 POR2X1_83/B POR2X1_172/CTRL 0.00fF
C28625 POR2X1_66/B POR2X1_588/Y 0.03fF
C28626 POR2X1_302/a_56_344# POR2X1_114/B 0.00fF
C28627 POR2X1_455/O POR2X1_702/A 0.00fF
C28628 POR2X1_7/B PAND2X1_506/CTRL2 0.00fF
C28629 POR2X1_288/A PAND2X1_60/B 0.03fF
C28630 PAND2X1_685/CTRL POR2X1_829/A 0.00fF
C28631 PAND2X1_862/B PAND2X1_798/B 0.03fF
C28632 POR2X1_853/A POR2X1_170/B 0.16fF
C28633 POR2X1_66/B POR2X1_101/Y 0.03fF
C28634 POR2X1_333/a_56_344# PAND2X1_20/A 0.00fF
C28635 POR2X1_360/A POR2X1_334/B 0.06fF
C28636 POR2X1_38/B POR2X1_236/O 0.05fF
C28637 PAND2X1_659/B POR2X1_56/Y 0.03fF
C28638 POR2X1_861/CTRL2 POR2X1_404/Y 0.08fF
C28639 PAND2X1_614/a_16_344# POR2X1_245/Y 0.02fF
C28640 POR2X1_90/Y VDD 1.89fF
C28641 POR2X1_602/B POR2X1_796/A 0.03fF
C28642 POR2X1_66/A POR2X1_703/CTRL 0.00fF
C28643 POR2X1_502/A PAND2X1_411/a_16_344# 0.01fF
C28644 POR2X1_137/Y PAND2X1_65/B 0.03fF
C28645 PAND2X1_477/B PAND2X1_445/Y 0.15fF
C28646 POR2X1_614/A POR2X1_483/O 0.10fF
C28647 PAND2X1_783/O PAND2X1_779/Y 0.04fF
C28648 POR2X1_440/Y POR2X1_186/Y 0.05fF
C28649 POR2X1_254/Y POR2X1_702/A 0.05fF
C28650 POR2X1_43/B PAND2X1_523/CTRL 0.30fF
C28651 PAND2X1_254/Y PAND2X1_6/A 0.02fF
C28652 PAND2X1_317/Y PAND2X1_552/B 0.12fF
C28653 PAND2X1_215/B POR2X1_599/A 0.10fF
C28654 POR2X1_393/Y POR2X1_394/O 0.01fF
C28655 PAND2X1_565/O POR2X1_46/Y 0.01fF
C28656 POR2X1_96/Y POR2X1_93/Y 0.04fF
C28657 POR2X1_16/A PAND2X1_733/A 0.07fF
C28658 PAND2X1_845/a_16_344# PAND2X1_673/Y 0.02fF
C28659 PAND2X1_23/Y POR2X1_775/A 0.01fF
C28660 POR2X1_415/a_16_28# POR2X1_816/A 0.00fF
C28661 POR2X1_300/m4_208_n4# POR2X1_46/Y 0.06fF
C28662 PAND2X1_65/CTRL POR2X1_4/Y 0.01fF
C28663 POR2X1_808/A POR2X1_598/a_56_344# 0.00fF
C28664 PAND2X1_69/A INPUT_4 3.53fF
C28665 PAND2X1_4/CTRL INPUT_0 0.00fF
C28666 POR2X1_41/B PAND2X1_653/Y 0.02fF
C28667 PAND2X1_319/B PAND2X1_151/CTRL 0.01fF
C28668 PAND2X1_671/O POR2X1_35/B 0.03fF
C28669 POR2X1_572/a_16_28# POR2X1_267/Y 0.08fF
C28670 POR2X1_293/Y POR2X1_816/A 0.03fF
C28671 PAND2X1_490/CTRL2 POR2X1_294/B 0.01fF
C28672 PAND2X1_90/Y POR2X1_520/CTRL2 0.01fF
C28673 PAND2X1_409/O PAND2X1_408/Y 0.03fF
C28674 POR2X1_438/Y PAND2X1_326/B 0.03fF
C28675 PAND2X1_661/B POR2X1_829/A 0.01fF
C28676 PAND2X1_56/Y POR2X1_741/Y 9.54fF
C28677 PAND2X1_26/A D_INPUT_4 0.09fF
C28678 POR2X1_7/B POR2X1_386/CTRL2 0.01fF
C28679 POR2X1_833/A POR2X1_777/B 0.15fF
C28680 POR2X1_829/A PAND2X1_643/Y 0.03fF
C28681 POR2X1_376/B POR2X1_428/CTRL2 0.03fF
C28682 POR2X1_46/CTRL2 POR2X1_153/Y 0.13fF
C28683 POR2X1_51/A POR2X1_36/B 0.09fF
C28684 POR2X1_806/CTRL2 POR2X1_737/A 0.01fF
C28685 POR2X1_247/CTRL2 POR2X1_532/A 0.01fF
C28686 PAND2X1_69/A POR2X1_785/A 0.03fF
C28687 POR2X1_383/A VDD 7.11fF
C28688 POR2X1_164/CTRL2 POR2X1_693/Y 0.01fF
C28689 PAND2X1_480/B POR2X1_387/Y 0.10fF
C28690 PAND2X1_473/B PAND2X1_175/CTRL 0.02fF
C28691 POR2X1_296/B POR2X1_788/CTRL2 0.05fF
C28692 POR2X1_575/B POR2X1_702/A 0.03fF
C28693 PAND2X1_23/Y POR2X1_112/Y 0.13fF
C28694 POR2X1_532/A POR2X1_783/B 0.02fF
C28695 POR2X1_538/CTRL2 PAND2X1_69/A 0.01fF
C28696 PAND2X1_846/O POR2X1_816/Y 0.02fF
C28697 PAND2X1_481/O POR2X1_355/A 0.02fF
C28698 POR2X1_840/B PAND2X1_55/Y 0.00fF
C28699 POR2X1_260/B PAND2X1_56/A 0.03fF
C28700 POR2X1_833/A PAND2X1_65/B 0.10fF
C28701 PAND2X1_624/A POR2X1_619/Y 0.21fF
C28702 PAND2X1_56/Y PAND2X1_32/B 0.07fF
C28703 POR2X1_795/B PAND2X1_32/B 0.17fF
C28704 POR2X1_42/Y POR2X1_748/a_76_344# 0.04fF
C28705 POR2X1_364/A POR2X1_357/Y 0.06fF
C28706 POR2X1_537/Y POR2X1_830/O 0.01fF
C28707 PAND2X1_476/A POR2X1_83/B 0.02fF
C28708 PAND2X1_194/CTRL2 POR2X1_42/Y 0.01fF
C28709 POR2X1_336/O POR2X1_741/Y 0.02fF
C28710 PAND2X1_5/O D_INPUT_2 0.02fF
C28711 PAND2X1_284/a_76_28# PAND2X1_566/Y 0.02fF
C28712 PAND2X1_90/A PAND2X1_150/a_76_28# 0.01fF
C28713 POR2X1_45/Y POR2X1_38/Y 0.03fF
C28714 PAND2X1_658/A POR2X1_93/A 0.03fF
C28715 PAND2X1_472/A PAND2X1_401/a_76_28# 0.01fF
C28716 PAND2X1_58/A PAND2X1_304/CTRL2 0.01fF
C28717 POR2X1_812/A POR2X1_691/A 0.27fF
C28718 POR2X1_8/Y POR2X1_29/O 0.00fF
C28719 POR2X1_39/Y POR2X1_236/Y 0.02fF
C28720 POR2X1_268/CTRL2 POR2X1_39/B 0.01fF
C28721 PAND2X1_48/B POR2X1_319/Y 0.03fF
C28722 POR2X1_370/O POR2X1_543/A 0.01fF
C28723 POR2X1_832/B POR2X1_592/CTRL2 0.01fF
C28724 PAND2X1_6/Y POR2X1_570/B 2.04fF
C28725 PAND2X1_732/A VDD 0.05fF
C28726 POR2X1_62/a_16_28# PAND2X1_69/A 0.03fF
C28727 POR2X1_616/Y POR2X1_750/B 0.09fF
C28728 PAND2X1_56/Y POR2X1_336/a_16_28# 0.02fF
C28729 POR2X1_672/O POR2X1_38/B 0.02fF
C28730 PAND2X1_58/O POR2X1_507/A 0.05fF
C28731 POR2X1_208/Y POR2X1_206/CTRL 0.08fF
C28732 POR2X1_394/A POR2X1_701/Y 0.01fF
C28733 POR2X1_16/Y VDD -0.00fF
C28734 PAND2X1_65/B PAND2X1_18/B 0.04fF
C28735 PAND2X1_341/A POR2X1_73/Y 0.17fF
C28736 POR2X1_383/A POR2X1_741/Y 0.17fF
C28737 PAND2X1_723/A PAND2X1_197/Y 0.31fF
C28738 PAND2X1_50/CTRL PAND2X1_18/B 0.06fF
C28739 PAND2X1_641/Y POR2X1_96/A 0.01fF
C28740 POR2X1_777/a_16_28# POR2X1_307/A 0.02fF
C28741 POR2X1_220/A POR2X1_162/O 0.05fF
C28742 PAND2X1_360/Y VDD 0.20fF
C28743 POR2X1_408/Y POR2X1_816/A 0.03fF
C28744 PAND2X1_778/CTRL2 PAND2X1_506/Y 0.00fF
C28745 POR2X1_73/Y POR2X1_91/Y 0.07fF
C28746 PAND2X1_71/Y VDD 0.57fF
C28747 POR2X1_83/B PAND2X1_327/CTRL2 0.05fF
C28748 PAND2X1_630/B POR2X1_628/Y 0.22fF
C28749 PAND2X1_469/B PAND2X1_353/O 0.11fF
C28750 POR2X1_334/Y POR2X1_220/Y 0.07fF
C28751 PAND2X1_858/CTRL INPUT_0 0.03fF
C28752 POR2X1_560/Y VDD 0.10fF
C28753 PAND2X1_71/O POR2X1_244/Y 0.07fF
C28754 POR2X1_394/A PAND2X1_364/B 0.07fF
C28755 PAND2X1_824/B POR2X1_785/A 0.07fF
C28756 POR2X1_110/Y VDD 0.41fF
C28757 POR2X1_383/A PAND2X1_32/B 0.17fF
C28758 PAND2X1_6/Y PAND2X1_368/CTRL 0.01fF
C28759 POR2X1_661/A POR2X1_260/B 0.07fF
C28760 POR2X1_539/A POR2X1_542/B 0.03fF
C28761 PAND2X1_659/Y POR2X1_393/O 0.01fF
C28762 POR2X1_708/O POR2X1_294/A 0.12fF
C28763 POR2X1_119/Y PAND2X1_556/B 0.03fF
C28764 PAND2X1_559/CTRL2 POR2X1_73/Y 0.05fF
C28765 PAND2X1_720/CTRL POR2X1_73/Y 0.04fF
C28766 PAND2X1_717/A POR2X1_20/B 0.03fF
C28767 POR2X1_857/O PAND2X1_72/A 0.01fF
C28768 PAND2X1_832/a_16_344# POR2X1_316/Y 0.02fF
C28769 POR2X1_307/a_16_28# POR2X1_711/Y 0.09fF
C28770 PAND2X1_244/B PAND2X1_341/A 0.03fF
C28771 POR2X1_60/A POR2X1_80/a_16_28# 0.02fF
C28772 PAND2X1_191/CTRL2 PAND2X1_730/A 0.00fF
C28773 POR2X1_45/Y POR2X1_153/Y 0.03fF
C28774 PAND2X1_39/B PAND2X1_32/CTRL 0.07fF
C28775 POR2X1_119/Y PAND2X1_254/Y 0.01fF
C28776 PAND2X1_863/B PAND2X1_729/CTRL 0.01fF
C28777 POR2X1_316/a_16_28# POR2X1_293/Y 0.02fF
C28778 POR2X1_52/A PAND2X1_330/CTRL2 0.00fF
C28779 PAND2X1_94/A POR2X1_410/Y 0.05fF
C28780 POR2X1_862/O POR2X1_814/B 0.01fF
C28781 POR2X1_59/O POR2X1_90/Y 0.01fF
C28782 PAND2X1_469/B POR2X1_129/Y 2.23fF
C28783 PAND2X1_569/B POR2X1_142/Y 0.07fF
C28784 PAND2X1_6/A PAND2X1_358/A 0.01fF
C28785 POR2X1_416/B PAND2X1_803/A 0.03fF
C28786 POR2X1_447/B POR2X1_629/A 0.06fF
C28787 POR2X1_62/O POR2X1_62/Y 0.08fF
C28788 PAND2X1_127/CTRL2 POR2X1_318/A 0.04fF
C28789 POR2X1_334/B POR2X1_571/Y 0.03fF
C28790 POR2X1_343/Y POR2X1_778/CTRL2 0.04fF
C28791 POR2X1_56/B PAND2X1_631/A 0.00fF
C28792 PAND2X1_803/CTRL POR2X1_90/Y 0.01fF
C28793 POR2X1_730/Y PAND2X1_163/CTRL2 0.01fF
C28794 PAND2X1_81/B PAND2X1_71/Y 0.04fF
C28795 PAND2X1_798/B PAND2X1_716/B 0.03fF
C28796 PAND2X1_862/B POR2X1_184/O 0.09fF
C28797 PAND2X1_727/O POR2X1_91/Y 0.02fF
C28798 PAND2X1_69/A POR2X1_186/B 0.04fF
C28799 PAND2X1_799/O PAND2X1_539/Y 0.03fF
C28800 POR2X1_822/O POR2X1_77/Y 0.16fF
C28801 PAND2X1_72/CTRL2 PAND2X1_48/A 0.01fF
C28802 POR2X1_43/B PAND2X1_851/CTRL 0.01fF
C28803 POR2X1_294/B PAND2X1_41/Y 0.01fF
C28804 POR2X1_442/CTRL POR2X1_411/B 0.00fF
C28805 POR2X1_383/A PAND2X1_253/O 0.04fF
C28806 POR2X1_732/B POR2X1_552/A 0.03fF
C28807 POR2X1_112/CTRL POR2X1_775/A 0.01fF
C28808 D_INPUT_1 PAND2X1_527/CTRL 0.03fF
C28809 POR2X1_9/Y POR2X1_29/A 0.03fF
C28810 POR2X1_725/Y POR2X1_308/B 0.17fF
C28811 D_INPUT_7 PAND2X1_429/CTRL 0.01fF
C28812 POR2X1_204/CTRL POR2X1_4/Y 0.01fF
C28813 PAND2X1_410/O POR2X1_411/A 0.01fF
C28814 POR2X1_416/B PAND2X1_673/Y 0.01fF
C28815 PAND2X1_649/A PAND2X1_649/O 0.01fF
C28816 POR2X1_657/Y POR2X1_222/CTRL2 0.01fF
C28817 POR2X1_776/B POR2X1_567/CTRL2 0.03fF
C28818 POR2X1_649/B POR2X1_294/A 0.37fF
C28819 PAND2X1_755/CTRL2 PAND2X1_72/A 0.01fF
C28820 POR2X1_16/A PAND2X1_124/CTRL 0.00fF
C28821 POR2X1_62/Y PAND2X1_350/CTRL2 0.01fF
C28822 VDD POR2X1_162/B 0.24fF
C28823 POR2X1_112/CTRL POR2X1_112/Y 0.00fF
C28824 POR2X1_257/A POR2X1_253/a_16_28# 0.01fF
C28825 PAND2X1_20/A PAND2X1_607/a_16_344# 0.01fF
C28826 PAND2X1_206/B POR2X1_614/Y 0.02fF
C28827 POR2X1_688/CTRL D_INPUT_0 0.01fF
C28828 PAND2X1_55/Y PAND2X1_56/A 0.12fF
C28829 PAND2X1_643/CTRL2 POR2X1_416/B 0.01fF
C28830 POR2X1_692/O POR2X1_20/B 0.03fF
C28831 PAND2X1_182/B PAND2X1_336/O 0.02fF
C28832 POR2X1_48/A POR2X1_253/CTRL2 0.01fF
C28833 POR2X1_23/Y POR2X1_253/CTRL 0.04fF
C28834 PAND2X1_126/O POR2X1_62/Y 0.05fF
C28835 POR2X1_73/Y PAND2X1_169/CTRL2 0.01fF
C28836 POR2X1_38/Y PAND2X1_379/CTRL 0.10fF
C28837 POR2X1_862/A POR2X1_643/Y 0.00fF
C28838 POR2X1_688/CTRL2 POR2X1_121/B 0.15fF
C28839 POR2X1_343/Y POR2X1_723/B 0.05fF
C28840 INPUT_3 POR2X1_37/Y 1.10fF
C28841 PAND2X1_123/O POR2X1_117/Y 0.01fF
C28842 POR2X1_311/O PAND2X1_336/Y 0.02fF
C28843 PAND2X1_341/A PAND2X1_358/CTRL 0.01fF
C28844 POR2X1_67/Y POR2X1_94/A 0.12fF
C28845 POR2X1_509/CTRL POR2X1_35/Y 0.01fF
C28846 PAND2X1_824/B POR2X1_186/B 0.07fF
C28847 POR2X1_193/A POR2X1_556/CTRL 0.03fF
C28848 POR2X1_329/A POR2X1_423/Y 0.13fF
C28849 POR2X1_460/A D_INPUT_4 0.19fF
C28850 POR2X1_864/A PAND2X1_829/O 0.00fF
C28851 POR2X1_294/A PAND2X1_103/O 0.09fF
C28852 POR2X1_826/Y POR2X1_32/A 0.09fF
C28853 POR2X1_343/A POR2X1_814/A 0.01fF
C28854 POR2X1_73/a_56_344# PAND2X1_341/B 0.00fF
C28855 POR2X1_475/O POR2X1_590/A 0.01fF
C28856 PAND2X1_699/O POR2X1_750/B 0.01fF
C28857 POR2X1_597/Y POR2X1_60/A 0.03fF
C28858 POR2X1_672/m4_208_n4# POR2X1_102/Y 0.01fF
C28859 POR2X1_9/Y POR2X1_546/A 0.09fF
C28860 POR2X1_614/A POR2X1_717/B 0.03fF
C28861 POR2X1_93/Y POR2X1_37/Y 3.79fF
C28862 PAND2X1_826/O POR2X1_202/B 0.05fF
C28863 POR2X1_445/A PAND2X1_73/Y 0.00fF
C28864 POR2X1_646/Y POR2X1_655/A 0.37fF
C28865 PAND2X1_73/Y POR2X1_643/Y 0.01fF
C28866 POR2X1_77/CTRL2 POR2X1_83/B 0.00fF
C28867 POR2X1_21/a_16_28# D_INPUT_4 0.01fF
C28868 POR2X1_614/A POR2X1_556/CTRL 0.00fF
C28869 POR2X1_434/a_16_28# POR2X1_434/A 0.01fF
C28870 POR2X1_661/A PAND2X1_55/Y 0.07fF
C28871 PAND2X1_86/CTRL2 VDD -0.00fF
C28872 POR2X1_257/A POR2X1_482/Y 0.07fF
C28873 POR2X1_648/Y VDD 0.21fF
C28874 POR2X1_444/Y POR2X1_738/O 0.11fF
C28875 POR2X1_85/Y POR2X1_235/O 0.16fF
C28876 PAND2X1_832/O POR2X1_271/B 0.02fF
C28877 POR2X1_333/A POR2X1_319/A 0.03fF
C28878 POR2X1_54/Y POR2X1_750/A 0.07fF
C28879 POR2X1_78/B PAND2X1_418/CTRL 0.04fF
C28880 POR2X1_728/A POR2X1_162/Y 2.03fF
C28881 POR2X1_814/A PAND2X1_89/CTRL2 0.03fF
C28882 POR2X1_304/CTRL2 POR2X1_153/Y 0.03fF
C28883 POR2X1_67/Y PAND2X1_754/CTRL2 0.01fF
C28884 PAND2X1_41/m4_208_n4# POR2X1_330/Y 0.12fF
C28885 POR2X1_376/B PAND2X1_98/CTRL 0.01fF
C28886 POR2X1_456/B PAND2X1_167/m4_208_n4# 0.12fF
C28887 POR2X1_807/CTRL POR2X1_590/A 0.01fF
C28888 POR2X1_66/A POR2X1_296/B 0.10fF
C28889 POR2X1_23/Y POR2X1_516/Y 0.02fF
C28890 POR2X1_98/CTRL2 POR2X1_590/A 0.00fF
C28891 POR2X1_294/Y POR2X1_202/B 0.00fF
C28892 POR2X1_20/B PAND2X1_541/a_76_28# 0.02fF
C28893 POR2X1_433/CTRL2 POR2X1_37/Y 0.01fF
C28894 PAND2X1_318/CTRL2 PAND2X1_464/B 0.03fF
C28895 POR2X1_341/A POR2X1_573/O 0.06fF
C28896 POR2X1_168/CTRL POR2X1_191/Y 0.24fF
C28897 POR2X1_168/O POR2X1_192/B 0.34fF
C28898 PAND2X1_563/A POR2X1_77/Y 0.02fF
C28899 POR2X1_389/A POR2X1_651/Y 0.39fF
C28900 POR2X1_78/B PAND2X1_41/O 0.03fF
C28901 PAND2X1_435/CTRL POR2X1_20/B 0.01fF
C28902 POR2X1_77/Y PAND2X1_337/CTRL 0.01fF
C28903 PAND2X1_156/A POR2X1_39/B 0.03fF
C28904 POR2X1_669/B POR2X1_819/a_16_28# 0.13fF
C28905 PAND2X1_798/B POR2X1_250/Y 0.07fF
C28906 POR2X1_541/B PAND2X1_48/a_56_28# 0.00fF
C28907 PAND2X1_848/a_76_28# POR2X1_669/B 0.04fF
C28908 POR2X1_41/B POR2X1_20/B 1.55fF
C28909 POR2X1_96/A POR2X1_63/Y 0.05fF
C28910 POR2X1_502/A POR2X1_663/B 0.07fF
C28911 PAND2X1_458/CTRL2 POR2X1_91/Y 0.03fF
C28912 PAND2X1_318/CTRL POR2X1_20/B 0.01fF
C28913 POR2X1_479/B POR2X1_389/Y 0.03fF
C28914 POR2X1_854/O POR2X1_192/Y 0.01fF
C28915 PAND2X1_137/O POR2X1_20/B 0.04fF
C28916 POR2X1_78/B POR2X1_644/O 0.05fF
C28917 POR2X1_63/Y POR2X1_406/CTRL 0.01fF
C28918 POR2X1_376/B PAND2X1_68/CTRL2 0.02fF
C28919 POR2X1_614/Y POR2X1_750/B 0.12fF
C28920 POR2X1_663/B PAND2X1_176/O 0.02fF
C28921 POR2X1_841/CTRL2 POR2X1_733/A 0.05fF
C28922 PAND2X1_818/O PAND2X1_340/B 0.02fF
C28923 POR2X1_602/B POR2X1_602/A 0.01fF
C28924 POR2X1_464/Y POR2X1_663/B 0.11fF
C28925 POR2X1_267/A POR2X1_267/a_16_28# -0.00fF
C28926 POR2X1_590/A POR2X1_186/Y 0.45fF
C28927 POR2X1_302/Y POR2X1_301/A 1.04fF
C28928 PAND2X1_622/CTRL POR2X1_29/A 0.01fF
C28929 POR2X1_476/Y PAND2X1_595/CTRL2 0.00fF
C28930 POR2X1_240/B PAND2X1_41/B 0.01fF
C28931 POR2X1_102/Y PAND2X1_140/CTRL 0.01fF
C28932 POR2X1_97/A PAND2X1_65/B 0.06fF
C28933 POR2X1_366/Y PAND2X1_268/CTRL 0.01fF
C28934 POR2X1_89/Y POR2X1_5/Y 0.01fF
C28935 POR2X1_471/A POR2X1_563/Y 0.01fF
C28936 PAND2X1_20/A PAND2X1_23/O 0.01fF
C28937 PAND2X1_601/m4_208_n4# PAND2X1_57/B 0.07fF
C28938 POR2X1_83/A PAND2X1_9/Y 0.03fF
C28939 POR2X1_78/Y POR2X1_844/B 0.01fF
C28940 POR2X1_69/Y POR2X1_7/A 0.01fF
C28941 POR2X1_843/a_16_28# POR2X1_343/A 0.02fF
C28942 POR2X1_843/a_76_344# POR2X1_287/B 0.00fF
C28943 PAND2X1_750/CTRL2 POR2X1_816/A 0.01fF
C28944 POR2X1_12/A POR2X1_587/CTRL2 0.10fF
C28945 POR2X1_32/A PAND2X1_713/B 0.01fF
C28946 POR2X1_462/a_16_28# POR2X1_532/A 0.05fF
C28947 POR2X1_654/B POR2X1_643/A 2.77fF
C28948 PAND2X1_446/Y PAND2X1_466/a_76_28# 0.05fF
C28949 POR2X1_707/A PAND2X1_41/B 0.01fF
C28950 POR2X1_609/Y POR2X1_609/A 0.03fF
C28951 POR2X1_713/A PAND2X1_20/A 0.04fF
C28952 PAND2X1_76/CTRL PAND2X1_76/Y 0.00fF
C28953 POR2X1_13/A PAND2X1_777/O 0.16fF
C28954 POR2X1_554/B POR2X1_228/Y 0.40fF
C28955 POR2X1_376/B POR2X1_748/A 0.12fF
C28956 PAND2X1_93/B POR2X1_832/B 0.03fF
C28957 PAND2X1_411/CTRL2 POR2X1_260/B 0.01fF
C28958 POR2X1_430/Y VDD 0.13fF
C28959 PAND2X1_272/CTRL2 POR2X1_465/B 0.03fF
C28960 PAND2X1_478/B POR2X1_236/Y 1.35fF
C28961 POR2X1_411/Y POR2X1_37/Y 0.03fF
C28962 POR2X1_139/A POR2X1_624/Y 0.04fF
C28963 POR2X1_480/A POR2X1_330/Y 0.10fF
C28964 POR2X1_290/Y POR2X1_667/Y 0.01fF
C28965 POR2X1_833/A POR2X1_814/A 0.10fF
C28966 POR2X1_485/Y PAND2X1_550/Y 0.01fF
C28967 POR2X1_207/CTRL2 POR2X1_330/Y 0.04fF
C28968 PAND2X1_485/CTRL POR2X1_789/A 0.11fF
C28969 POR2X1_302/O POR2X1_302/B 0.01fF
C28970 POR2X1_12/A D_INPUT_6 0.01fF
C28971 POR2X1_226/Y POR2X1_5/Y 0.06fF
C28972 INPUT_3 POR2X1_408/Y 0.12fF
C28973 POR2X1_63/Y POR2X1_7/A 0.08fF
C28974 PAND2X1_404/A PAND2X1_404/a_76_28# 0.01fF
C28975 POR2X1_383/A PAND2X1_9/Y 0.03fF
C28976 PAND2X1_65/B POR2X1_650/A 0.04fF
C28977 POR2X1_114/Y POR2X1_390/a_16_28# 0.03fF
C28978 PAND2X1_474/Y PAND2X1_500/O 0.00fF
C28979 PAND2X1_736/A POR2X1_32/A 0.07fF
C28980 POR2X1_20/B PAND2X1_100/CTRL2 0.10fF
C28981 PAND2X1_217/B INPUT_0 0.51fF
C28982 POR2X1_849/A POR2X1_790/A 0.54fF
C28983 POR2X1_257/A PAND2X1_349/A 0.06fF
C28984 PAND2X1_473/Y PAND2X1_576/CTRL2 0.03fF
C28985 POR2X1_78/A POR2X1_832/B 0.09fF
C28986 POR2X1_65/A PAND2X1_206/O 0.15fF
C28987 POR2X1_177/Y PAND2X1_180/O -0.00fF
C28988 POR2X1_40/Y POR2X1_817/A 0.01fF
C28989 D_INPUT_2 POR2X1_414/O 0.02fF
C28990 POR2X1_487/O PAND2X1_794/B 0.02fF
C28991 POR2X1_423/Y POR2X1_256/O 0.01fF
C28992 PAND2X1_659/A PAND2X1_735/Y 0.13fF
C28993 POR2X1_52/A POR2X1_748/A 0.03fF
C28994 PAND2X1_39/B POR2X1_796/A 0.07fF
C28995 POR2X1_291/O POR2X1_20/B 0.01fF
C28996 POR2X1_121/A POR2X1_590/A 0.03fF
C28997 PAND2X1_420/O POR2X1_785/A 0.06fF
C28998 POR2X1_88/CTRL2 POR2X1_7/A 0.01fF
C28999 PAND2X1_456/CTRL2 PAND2X1_254/Y 0.01fF
C29000 POR2X1_805/CTRL PAND2X1_60/B 0.01fF
C29001 PAND2X1_798/B PAND2X1_798/O 0.07fF
C29002 POR2X1_846/B POR2X1_14/Y 0.11fF
C29003 PAND2X1_41/B POR2X1_190/Y 0.02fF
C29004 POR2X1_68/a_16_28# POR2X1_402/A 0.02fF
C29005 PAND2X1_831/Y POR2X1_271/O 0.01fF
C29006 POR2X1_856/B POR2X1_540/A 0.03fF
C29007 PAND2X1_56/Y POR2X1_830/Y 0.29fF
C29008 POR2X1_566/A PAND2X1_52/Y 0.05fF
C29009 POR2X1_66/B PAND2X1_23/Y 0.26fF
C29010 POR2X1_436/O POR2X1_802/B 0.01fF
C29011 PAND2X1_272/CTRL PAND2X1_32/B 0.01fF
C29012 POR2X1_407/A POR2X1_390/CTRL2 0.00fF
C29013 POR2X1_341/A POR2X1_456/B 0.03fF
C29014 POR2X1_20/B PAND2X1_308/Y 0.03fF
C29015 POR2X1_866/CTRL POR2X1_800/A 0.00fF
C29016 POR2X1_446/B POR2X1_714/m4_208_n4# 0.12fF
C29017 POR2X1_40/Y POR2X1_42/Y 0.17fF
C29018 POR2X1_399/A PAND2X1_403/B 0.03fF
C29019 POR2X1_49/Y PAND2X1_454/CTRL 0.06fF
C29020 INPUT_2 POR2X1_29/A 0.03fF
C29021 POR2X1_271/B POR2X1_153/Y 0.05fF
C29022 PAND2X1_63/Y PAND2X1_73/Y 0.07fF
C29023 POR2X1_188/A PAND2X1_23/Y 0.05fF
C29024 POR2X1_102/Y POR2X1_239/CTRL2 0.01fF
C29025 POR2X1_66/B PAND2X1_625/O 0.01fF
C29026 PAND2X1_557/A PAND2X1_652/A 0.24fF
C29027 PAND2X1_48/B POR2X1_734/A 0.12fF
C29028 PAND2X1_39/CTRL PAND2X1_69/A 0.01fF
C29029 POR2X1_251/CTRL PAND2X1_190/Y 0.02fF
C29030 POR2X1_567/B PAND2X1_173/a_56_28# 0.00fF
C29031 PAND2X1_742/B POR2X1_331/Y 0.05fF
C29032 POR2X1_65/A POR2X1_314/O 0.07fF
C29033 POR2X1_60/A POR2X1_816/A 0.06fF
C29034 INPUT_0 VDD 15.28fF
C29035 POR2X1_532/A POR2X1_296/B 0.13fF
C29036 PAND2X1_553/B POR2X1_106/Y 0.22fF
C29037 POR2X1_634/A POR2X1_771/CTRL2 0.06fF
C29038 PAND2X1_39/B PAND2X1_399/CTRL2 0.01fF
C29039 PAND2X1_460/Y PAND2X1_8/Y 0.01fF
C29040 POR2X1_753/Y POR2X1_93/A 0.19fF
C29041 PAND2X1_635/CTRL2 POR2X1_748/A 0.03fF
C29042 PAND2X1_214/a_16_344# PAND2X1_656/A 0.01fF
C29043 PAND2X1_229/CTRL2 D_GATE_222 0.03fF
C29044 POR2X1_462/B POR2X1_634/A 0.03fF
C29045 POR2X1_40/Y POR2X1_309/Y 0.08fF
C29046 POR2X1_8/Y PAND2X1_35/A 0.05fF
C29047 POR2X1_565/B POR2X1_5/Y 0.12fF
C29048 POR2X1_862/A POR2X1_260/A 0.07fF
C29049 PAND2X1_55/Y PAND2X1_13/a_16_344# 0.02fF
C29050 POR2X1_48/A PAND2X1_114/CTRL2 0.01fF
C29051 PAND2X1_58/A POR2X1_550/O 0.01fF
C29052 PAND2X1_57/B PAND2X1_587/Y 0.16fF
C29053 POR2X1_366/Y PAND2X1_65/B 0.07fF
C29054 POR2X1_417/Y PAND2X1_457/O 0.03fF
C29055 PAND2X1_65/B POR2X1_294/B 0.20fF
C29056 PAND2X1_808/Y PAND2X1_363/Y 0.04fF
C29057 POR2X1_634/O PAND2X1_32/B 0.18fF
C29058 POR2X1_496/Y PAND2X1_549/B 0.07fF
C29059 POR2X1_116/A POR2X1_362/O 0.00fF
C29060 POR2X1_71/Y PAND2X1_659/B 0.03fF
C29061 POR2X1_555/A POR2X1_68/A 0.17fF
C29062 PAND2X1_41/O POR2X1_294/A 0.15fF
C29063 POR2X1_150/Y PAND2X1_353/Y 0.13fF
C29064 PAND2X1_825/O POR2X1_296/B 0.15fF
C29065 POR2X1_612/Y POR2X1_4/O 0.03fF
C29066 POR2X1_447/B PAND2X1_43/CTRL 0.06fF
C29067 POR2X1_54/Y POR2X1_773/A 0.03fF
C29068 POR2X1_423/Y PAND2X1_702/CTRL 0.01fF
C29069 PAND2X1_842/a_16_344# POR2X1_184/Y 0.02fF
C29070 POR2X1_817/CTRL2 POR2X1_394/A 0.05fF
C29071 POR2X1_362/Y POR2X1_366/A 0.00fF
C29072 POR2X1_832/O POR2X1_832/B 0.01fF
C29073 POR2X1_779/A PAND2X1_90/Y 0.06fF
C29074 POR2X1_52/A POR2X1_79/Y 0.03fF
C29075 POR2X1_5/Y POR2X1_56/Y 0.03fF
C29076 PAND2X1_267/Y PAND2X1_853/B 0.03fF
C29077 POR2X1_56/B PAND2X1_471/B 0.29fF
C29078 POR2X1_606/CTRL2 PAND2X1_48/A 0.03fF
C29079 POR2X1_280/CTRL2 POR2X1_312/Y 0.03fF
C29080 INPUT_1 POR2X1_609/Y 0.03fF
C29081 PAND2X1_849/B POR2X1_669/B 0.02fF
C29082 POR2X1_57/A POR2X1_423/Y 0.03fF
C29083 D_INPUT_3 POR2X1_293/CTRL2 0.01fF
C29084 PAND2X1_6/A PAND2X1_381/O 0.04fF
C29085 POR2X1_438/a_16_28# POR2X1_72/B 0.03fF
C29086 POR2X1_198/O VDD 0.00fF
C29087 PAND2X1_20/A PAND2X1_397/O 0.02fF
C29088 POR2X1_580/CTRL D_GATE_741 0.06fF
C29089 POR2X1_443/A POR2X1_551/A 0.02fF
C29090 POR2X1_260/B POR2X1_737/A 0.02fF
C29091 POR2X1_777/B PAND2X1_111/B 0.04fF
C29092 PAND2X1_483/O POR2X1_669/B -0.01fF
C29093 PAND2X1_73/Y POR2X1_260/A 1.22fF
C29094 PAND2X1_96/B POR2X1_362/B 0.59fF
C29095 POR2X1_422/Y POR2X1_260/A 0.03fF
C29096 POR2X1_68/A POR2X1_544/A 0.07fF
C29097 POR2X1_43/B POR2X1_88/Y 0.03fF
C29098 POR2X1_857/A POR2X1_568/B 0.00fF
C29099 POR2X1_537/B POR2X1_389/Y 1.78fF
C29100 POR2X1_83/B POR2X1_176/Y 0.01fF
C29101 POR2X1_48/A PAND2X1_156/A 0.08fF
C29102 POR2X1_57/A POR2X1_323/O 0.02fF
C29103 PAND2X1_65/Y POR2X1_205/A 0.02fF
C29104 POR2X1_460/A PAND2X1_21/CTRL 0.00fF
C29105 PAND2X1_793/Y PAND2X1_658/B 0.05fF
C29106 POR2X1_96/A PAND2X1_631/CTRL2 0.00fF
C29107 POR2X1_279/Y POR2X1_258/Y 0.12fF
C29108 POR2X1_130/A D_INPUT_1 4.67fF
C29109 POR2X1_38/Y PAND2X1_340/a_76_28# 0.02fF
C29110 POR2X1_49/Y PAND2X1_63/B 0.03fF
C29111 POR2X1_66/B POR2X1_537/CTRL2 0.09fF
C29112 POR2X1_625/Y PAND2X1_6/A 0.39fF
C29113 POR2X1_539/CTRL2 POR2X1_750/B 0.01fF
C29114 PAND2X1_848/B POR2X1_817/A 0.66fF
C29115 PAND2X1_764/a_16_344# PAND2X1_41/B 0.02fF
C29116 INPUT_0 PAND2X1_32/B 0.16fF
C29117 PAND2X1_65/B PAND2X1_111/B 0.03fF
C29118 PAND2X1_857/CTRL2 POR2X1_23/Y 0.01fF
C29119 POR2X1_20/B POR2X1_77/Y 0.22fF
C29120 PAND2X1_738/Y PAND2X1_113/CTRL2 0.08fF
C29121 POR2X1_135/CTRL2 POR2X1_48/A 0.01fF
C29122 PAND2X1_748/CTRL2 POR2X1_752/Y 0.01fF
C29123 POR2X1_65/A POR2X1_103/Y 0.04fF
C29124 POR2X1_346/B POR2X1_330/Y 0.03fF
C29125 POR2X1_218/A POR2X1_404/Y 0.07fF
C29126 PAND2X1_469/B POR2X1_293/Y 0.05fF
C29127 POR2X1_324/A POR2X1_568/Y 0.38fF
C29128 PAND2X1_57/B POR2X1_770/CTRL 0.01fF
C29129 POR2X1_537/CTRL2 POR2X1_188/A 0.01fF
C29130 POR2X1_25/Y POR2X1_26/a_16_28# 0.02fF
C29131 POR2X1_500/A POR2X1_456/B 0.01fF
C29132 POR2X1_96/A POR2X1_498/A 0.02fF
C29133 PAND2X1_48/B PAND2X1_145/a_16_344# 0.01fF
C29134 POR2X1_570/O POR2X1_570/B 0.02fF
C29135 POR2X1_780/A VDD 0.00fF
C29136 PAND2X1_777/CTRL PAND2X1_784/A 0.01fF
C29137 POR2X1_193/Y POR2X1_200/A 0.00fF
C29138 POR2X1_364/A POR2X1_578/Y 0.03fF
C29139 POR2X1_351/Y POR2X1_579/Y 0.11fF
C29140 PAND2X1_393/CTRL2 VDD 0.00fF
C29141 PAND2X1_383/O POR2X1_236/Y 0.04fF
C29142 POR2X1_137/CTRL2 PAND2X1_32/B 0.00fF
C29143 PAND2X1_105/O POR2X1_55/Y 0.06fF
C29144 PAND2X1_95/B POR2X1_638/B 0.01fF
C29145 PAND2X1_57/B PAND2X1_88/Y 0.03fF
C29146 PAND2X1_848/B POR2X1_42/Y 0.05fF
C29147 PAND2X1_773/O POR2X1_7/B 0.04fF
C29148 POR2X1_502/A POR2X1_544/CTRL 0.01fF
C29149 PAND2X1_115/B POR2X1_310/CTRL 0.04fF
C29150 PAND2X1_797/Y POR2X1_23/Y 0.03fF
C29151 PAND2X1_57/B POR2X1_84/Y 0.01fF
C29152 POR2X1_566/A POR2X1_724/A 0.03fF
C29153 PAND2X1_90/Y POR2X1_407/CTRL 0.02fF
C29154 POR2X1_96/A PAND2X1_284/Y 0.01fF
C29155 PAND2X1_48/B POR2X1_786/Y 0.09fF
C29156 POR2X1_49/Y PAND2X1_480/CTRL2 0.01fF
C29157 PAND2X1_90/Y POR2X1_317/A 0.00fF
C29158 POR2X1_308/O POR2X1_725/Y 0.04fF
C29159 POR2X1_111/Y POR2X1_423/Y 0.02fF
C29160 D_GATE_222 D_GATE_741 0.02fF
C29161 POR2X1_65/A POR2X1_313/Y 0.03fF
C29162 POR2X1_32/A POR2X1_7/Y 0.03fF
C29163 PAND2X1_139/B POR2X1_7/A 0.01fF
C29164 PAND2X1_659/Y POR2X1_498/Y 0.32fF
C29165 POR2X1_480/A POR2X1_799/O 0.03fF
C29166 POR2X1_72/B PAND2X1_200/B 0.06fF
C29167 POR2X1_669/B POR2X1_749/Y 0.57fF
C29168 POR2X1_463/Y POR2X1_805/B 0.48fF
C29169 POR2X1_383/A POR2X1_483/CTRL2 0.06fF
C29170 PAND2X1_139/B PAND2X1_130/O 0.00fF
C29171 POR2X1_722/Y POR2X1_513/O 0.01fF
C29172 POR2X1_327/Y POR2X1_453/a_16_28# 0.07fF
C29173 PAND2X1_444/a_16_344# POR2X1_39/B 0.02fF
C29174 PAND2X1_745/a_16_344# PAND2X1_41/B 0.02fF
C29175 POR2X1_618/CTRL2 POR2X1_7/A 0.03fF
C29176 POR2X1_427/Y POR2X1_394/A 0.03fF
C29177 PAND2X1_784/CTRL POR2X1_387/Y 0.04fF
C29178 POR2X1_49/Y POR2X1_144/O 0.01fF
C29179 PAND2X1_46/CTRL POR2X1_294/A 0.00fF
C29180 POR2X1_401/A POR2X1_68/B 0.01fF
C29181 D_INPUT_3 PAND2X1_341/O 0.15fF
C29182 PAND2X1_20/A POR2X1_554/CTRL2 0.01fF
C29183 POR2X1_647/O PAND2X1_52/B 0.02fF
C29184 POR2X1_426/CTRL POR2X1_425/Y 0.01fF
C29185 POR2X1_673/Y INPUT_0 0.21fF
C29186 PAND2X1_496/CTRL2 POR2X1_569/A 0.01fF
C29187 POR2X1_796/A POR2X1_513/B 0.06fF
C29188 POR2X1_529/Y POR2X1_55/Y 0.23fF
C29189 PAND2X1_363/Y PAND2X1_354/Y 0.18fF
C29190 POR2X1_244/B POR2X1_259/a_16_28# 0.02fF
C29191 PAND2X1_291/CTRL2 POR2X1_35/Y 0.01fF
C29192 POR2X1_346/O POR2X1_68/A 0.02fF
C29193 POR2X1_16/A POR2X1_13/A 0.16fF
C29194 PAND2X1_63/Y PAND2X1_316/m4_208_n4# 0.06fF
C29195 POR2X1_542/B PAND2X1_69/A 0.03fF
C29196 PAND2X1_390/Y PAND2X1_851/a_16_344# 0.01fF
C29197 POR2X1_810/a_16_28# POR2X1_809/Y 0.07fF
C29198 POR2X1_315/O POR2X1_91/Y 0.01fF
C29199 INPUT_7 PAND2X1_3/B 0.01fF
C29200 PAND2X1_79/Y PAND2X1_69/A 0.22fF
C29201 PAND2X1_849/B PAND2X1_844/Y 0.01fF
C29202 PAND2X1_539/Y POR2X1_7/B 0.03fF
C29203 POR2X1_416/B POR2X1_626/a_16_28# 0.03fF
C29204 PAND2X1_566/Y PAND2X1_347/a_76_28# 0.02fF
C29205 POR2X1_165/CTRL2 POR2X1_73/Y 0.01fF
C29206 PAND2X1_58/A D_INPUT_4 0.02fF
C29207 D_INPUT_0 POR2X1_522/a_56_344# 0.00fF
C29208 POR2X1_16/A POR2X1_57/O -0.01fF
C29209 POR2X1_565/B POR2X1_6/CTRL2 0.00fF
C29210 POR2X1_41/B PAND2X1_303/Y 0.06fF
C29211 PAND2X1_442/O POR2X1_192/B 0.06fF
C29212 PAND2X1_442/CTRL2 POR2X1_191/Y 0.01fF
C29213 PAND2X1_25/CTRL PAND2X1_52/B 0.01fF
C29214 POR2X1_81/A PAND2X1_244/a_76_28# 0.03fF
C29215 POR2X1_186/CTRL2 PAND2X1_55/Y 0.00fF
C29216 PAND2X1_220/m4_208_n4# POR2X1_142/Y 0.09fF
C29217 POR2X1_228/Y POR2X1_702/A 0.03fF
C29218 POR2X1_724/A POR2X1_573/A 0.03fF
C29219 PAND2X1_41/B PAND2X1_759/O 0.01fF
C29220 POR2X1_855/B POR2X1_796/O 0.01fF
C29221 POR2X1_567/A PAND2X1_65/B 0.08fF
C29222 POR2X1_78/CTRL2 POR2X1_569/A 0.03fF
C29223 POR2X1_57/A PAND2X1_319/B 0.11fF
C29224 PAND2X1_338/B POR2X1_73/Y 0.03fF
C29225 POR2X1_210/O PAND2X1_52/B 0.01fF
C29226 PAND2X1_60/B POR2X1_140/CTRL2 0.01fF
C29227 POR2X1_463/a_16_28# POR2X1_459/Y -0.00fF
C29228 PAND2X1_6/Y POR2X1_569/A 0.07fF
C29229 PAND2X1_341/B POR2X1_236/Y 0.05fF
C29230 PAND2X1_741/B POR2X1_7/Y 0.02fF
C29231 POR2X1_108/CTRL POR2X1_142/Y 0.01fF
C29232 POR2X1_492/Y POR2X1_492/O 0.02fF
C29233 POR2X1_66/B POR2X1_711/Y 0.43fF
C29234 POR2X1_92/CTRL2 POR2X1_408/Y 0.41fF
C29235 POR2X1_7/B PAND2X1_507/O 0.05fF
C29236 PAND2X1_341/A PAND2X1_656/A 2.13fF
C29237 POR2X1_38/B POR2X1_384/CTRL 0.01fF
C29238 PAND2X1_658/A PAND2X1_789/CTRL2 0.01fF
C29239 PAND2X1_816/a_76_28# POR2X1_463/Y 0.02fF
C29240 POR2X1_349/a_16_28# PAND2X1_65/Y 0.01fF
C29241 POR2X1_590/A POR2X1_717/B 6.41fF
C29242 PAND2X1_785/Y POR2X1_109/Y -0.00fF
C29243 POR2X1_325/O POR2X1_542/B 0.01fF
C29244 PAND2X1_534/O POR2X1_788/B 0.01fF
C29245 POR2X1_383/A POR2X1_639/Y 0.03fF
C29246 POR2X1_390/B POR2X1_301/O -0.00fF
C29247 POR2X1_505/Y POR2X1_416/B 0.08fF
C29248 INPUT_5 PAND2X1_18/B 0.10fF
C29249 INPUT_4 PAND2X1_3/B 0.03fF
C29250 POR2X1_8/Y POR2X1_43/B 3.15fF
C29251 PAND2X1_793/Y PAND2X1_657/B 0.21fF
C29252 D_INPUT_6 PAND2X1_1/CTRL 0.02fF
C29253 POR2X1_356/A POR2X1_209/a_56_344# 0.03fF
C29254 POR2X1_359/O PAND2X1_57/B 0.01fF
C29255 POR2X1_417/a_16_28# POR2X1_283/A 0.09fF
C29256 POR2X1_532/A POR2X1_520/CTRL 0.00fF
C29257 POR2X1_567/A POR2X1_653/a_16_28# 0.03fF
C29258 PAND2X1_574/O POR2X1_73/Y 0.17fF
C29259 PAND2X1_322/CTRL2 POR2X1_188/Y 0.06fF
C29260 PAND2X1_140/A PAND2X1_348/Y 0.16fF
C29261 POR2X1_631/B POR2X1_260/A 0.03fF
C29262 PAND2X1_83/a_76_28# PAND2X1_82/Y 0.01fF
C29263 POR2X1_96/A PAND2X1_802/O 0.05fF
C29264 POR2X1_52/A PAND2X1_730/A 0.03fF
C29265 POR2X1_795/a_16_28# POR2X1_186/B 0.02fF
C29266 POR2X1_575/CTRL2 POR2X1_569/A 0.04fF
C29267 POR2X1_327/Y POR2X1_335/A 0.03fF
C29268 POR2X1_661/CTRL POR2X1_711/Y 0.06fF
C29269 PAND2X1_65/B POR2X1_779/CTRL2 0.01fF
C29270 POR2X1_16/A PAND2X1_661/B 0.03fF
C29271 PAND2X1_556/B PAND2X1_326/B 0.03fF
C29272 POR2X1_16/A PAND2X1_643/Y 0.11fF
C29273 PAND2X1_23/Y POR2X1_54/O 0.00fF
C29274 PAND2X1_824/B POR2X1_208/Y 0.03fF
C29275 POR2X1_554/B POR2X1_657/Y 0.03fF
C29276 POR2X1_705/B POR2X1_556/A 0.12fF
C29277 POR2X1_9/Y PAND2X1_66/a_76_28# 0.04fF
C29278 POR2X1_208/A POR2X1_201/Y 0.29fF
C29279 POR2X1_236/Y POR2X1_533/Y 0.03fF
C29280 POR2X1_68/B POR2X1_768/CTRL 0.01fF
C29281 POR2X1_832/CTRL2 POR2X1_711/Y 0.03fF
C29282 PAND2X1_809/B VDD 0.01fF
C29283 POR2X1_713/CTRL2 PAND2X1_48/A 0.01fF
C29284 POR2X1_567/A POR2X1_231/O 0.06fF
C29285 PAND2X1_99/B PAND2X1_99/O 0.01fF
C29286 POR2X1_8/Y POR2X1_38/B 1.13fF
C29287 PAND2X1_641/Y POR2X1_38/Y 0.00fF
C29288 PAND2X1_94/A PAND2X1_60/B 0.40fF
C29289 POR2X1_447/B POR2X1_740/Y 0.10fF
C29290 POR2X1_158/Y PAND2X1_712/B 0.00fF
C29291 PAND2X1_793/Y POR2X1_184/CTRL2 0.01fF
C29292 PAND2X1_18/CTRL2 PAND2X1_52/B 0.15fF
C29293 POR2X1_334/B PAND2X1_134/CTRL2 0.13fF
C29294 POR2X1_614/A POR2X1_370/O 0.01fF
C29295 POR2X1_527/CTRL2 PAND2X1_550/B 0.01fF
C29296 PAND2X1_700/CTRL2 PAND2X1_52/B 0.14fF
C29297 PAND2X1_33/CTRL POR2X1_24/Y 0.01fF
C29298 POR2X1_327/Y POR2X1_361/CTRL2 0.01fF
C29299 PAND2X1_687/CTRL PAND2X1_643/Y 0.02fF
C29300 POR2X1_814/B POR2X1_863/A 0.07fF
C29301 POR2X1_58/Y POR2X1_39/B 0.14fF
C29302 PAND2X1_281/O POR2X1_649/B 0.14fF
C29303 POR2X1_97/A POR2X1_814/A 0.07fF
C29304 POR2X1_532/A POR2X1_342/CTRL 0.01fF
C29305 POR2X1_569/Y POR2X1_570/Y -0.00fF
C29306 POR2X1_155/Y POR2X1_728/A 0.00fF
C29307 POR2X1_65/A POR2X1_825/Y 0.02fF
C29308 POR2X1_264/Y POR2X1_383/Y 0.11fF
C29309 POR2X1_99/Y PAND2X1_39/B 0.07fF
C29310 POR2X1_416/B POR2X1_411/O 0.02fF
C29311 POR2X1_383/A POR2X1_558/Y 0.03fF
C29312 PAND2X1_48/A POR2X1_318/A 0.07fF
C29313 POR2X1_334/Y POR2X1_222/A 0.03fF
C29314 PAND2X1_48/A POR2X1_713/B 0.01fF
C29315 POR2X1_416/B PAND2X1_35/CTRL2 0.01fF
C29316 POR2X1_610/Y POR2X1_862/A 0.07fF
C29317 POR2X1_416/B POR2X1_32/O 0.02fF
C29318 POR2X1_356/A PAND2X1_52/B 0.07fF
C29319 PAND2X1_631/A POR2X1_93/A 0.01fF
C29320 POR2X1_41/B POR2X1_43/Y 0.03fF
C29321 PAND2X1_631/A POR2X1_91/Y 0.07fF
C29322 POR2X1_396/O POR2X1_39/B 0.17fF
C29323 POR2X1_557/A POR2X1_557/B 0.41fF
C29324 PAND2X1_308/Y PAND2X1_303/Y 0.01fF
C29325 PAND2X1_272/O POR2X1_556/A 0.07fF
C29326 POR2X1_97/a_56_344# POR2X1_186/B 0.00fF
C29327 POR2X1_66/CTRL PAND2X1_58/A 0.03fF
C29328 POR2X1_554/B POR2X1_657/O 0.08fF
C29329 POR2X1_332/Y POR2X1_332/CTRL2 0.01fF
C29330 POR2X1_165/O PAND2X1_326/B 0.01fF
C29331 POR2X1_54/Y POR2X1_409/B 0.07fF
C29332 POR2X1_440/B POR2X1_186/Y 0.03fF
C29333 POR2X1_440/CTRL VDD 0.00fF
C29334 POR2X1_862/O PAND2X1_32/B 0.06fF
C29335 POR2X1_474/CTRL2 POR2X1_556/A 0.01fF
C29336 POR2X1_39/B POR2X1_9/CTRL 0.29fF
C29337 POR2X1_795/B POR2X1_568/A 0.01fF
C29338 PAND2X1_157/CTRL PAND2X1_3/B 0.01fF
C29339 POR2X1_257/A POR2X1_32/A 12.75fF
C29340 PAND2X1_6/Y PAND2X1_72/A 2.60fF
C29341 POR2X1_137/B POR2X1_634/A 0.04fF
C29342 POR2X1_537/Y POR2X1_851/CTRL 0.01fF
C29343 POR2X1_463/CTRL2 VDD 0.00fF
C29344 POR2X1_491/Y PAND2X1_717/Y 0.12fF
C29345 PAND2X1_464/O POR2X1_417/Y 0.03fF
C29346 POR2X1_841/CTRL POR2X1_330/Y 0.01fF
C29347 PAND2X1_97/Y POR2X1_5/Y 0.01fF
C29348 POR2X1_54/Y POR2X1_55/a_16_28# 0.03fF
C29349 PAND2X1_85/CTRL2 INPUT_0 0.00fF
C29350 POR2X1_99/A POR2X1_99/a_16_28# 0.01fF
C29351 POR2X1_632/Y POR2X1_569/A 0.07fF
C29352 POR2X1_220/A PAND2X1_52/B 0.88fF
C29353 POR2X1_428/Y POR2X1_60/A 0.00fF
C29354 PAND2X1_313/CTRL2 POR2X1_169/A 0.01fF
C29355 POR2X1_850/A POR2X1_287/A 0.03fF
C29356 PAND2X1_93/B POR2X1_269/O 0.02fF
C29357 PAND2X1_717/A PAND2X1_579/B 6.90fF
C29358 POR2X1_257/A POR2X1_417/Y 0.06fF
C29359 PAND2X1_20/A POR2X1_274/A 0.03fF
C29360 PAND2X1_485/CTRL POR2X1_590/A 0.01fF
C29361 POR2X1_313/a_76_344# POR2X1_167/Y 0.00fF
C29362 POR2X1_129/CTRL2 POR2X1_67/A 0.10fF
C29363 POR2X1_635/B PAND2X1_47/CTRL 0.00fF
C29364 POR2X1_265/O POR2X1_667/A 0.19fF
C29365 POR2X1_569/A POR2X1_500/CTRL 0.04fF
C29366 PAND2X1_175/B POR2X1_173/CTRL 0.01fF
C29367 POR2X1_661/A PAND2X1_385/a_76_28# 0.02fF
C29368 POR2X1_60/A POR2X1_93/Y 0.03fF
C29369 POR2X1_37/CTRL2 POR2X1_612/Y 0.05fF
C29370 POR2X1_86/Y PAND2X1_100/CTRL2 0.00fF
C29371 POR2X1_669/B POR2X1_626/O 0.02fF
C29372 PAND2X1_632/B POR2X1_416/B 0.18fF
C29373 POR2X1_416/B PAND2X1_593/Y 0.03fF
C29374 PAND2X1_611/a_16_344# POR2X1_130/A 0.07fF
C29375 POR2X1_569/A PAND2X1_52/B 0.03fF
C29376 PAND2X1_201/CTRL2 POR2X1_88/Y 0.00fF
C29377 POR2X1_54/Y PAND2X1_526/O 0.02fF
C29378 POR2X1_99/Y POR2X1_814/B 0.02fF
C29379 POR2X1_129/CTRL POR2X1_83/B 0.01fF
C29380 POR2X1_814/A POR2X1_294/B 0.35fF
C29381 PAND2X1_698/CTRL PAND2X1_52/B 0.02fF
C29382 POR2X1_570/Y PAND2X1_52/B 0.07fF
C29383 PAND2X1_64/m4_208_n4# PAND2X1_11/Y 0.09fF
C29384 POR2X1_52/A POR2X1_815/O 0.02fF
C29385 POR2X1_274/A POR2X1_814/B 0.03fF
C29386 POR2X1_454/A PAND2X1_229/O 0.04fF
C29387 POR2X1_567/B POR2X1_857/m4_208_n4# 0.06fF
C29388 PAND2X1_9/Y INPUT_0 0.05fF
C29389 PAND2X1_798/B POR2X1_329/A 0.03fF
C29390 PAND2X1_39/B POR2X1_403/B 0.01fF
C29391 PAND2X1_502/CTRL POR2X1_77/Y 0.01fF
C29392 D_INPUT_5 PAND2X1_21/O 0.02fF
C29393 D_INPUT_0 PAND2X1_390/Y 0.03fF
C29394 PAND2X1_635/Y INPUT_6 0.03fF
C29395 PAND2X1_57/B POR2X1_341/A 0.07fF
C29396 POR2X1_66/A POR2X1_186/Y 0.10fF
C29397 POR2X1_68/A PAND2X1_617/CTRL 0.02fF
C29398 POR2X1_105/Y PAND2X1_251/O 0.01fF
C29399 POR2X1_262/Y POR2X1_293/Y 0.16fF
C29400 PAND2X1_414/m4_208_n4# POR2X1_42/Y 0.04fF
C29401 PAND2X1_340/B VDD 0.38fF
C29402 PAND2X1_116/CTRL POR2X1_48/A 0.01fF
C29403 PAND2X1_865/Y POR2X1_767/Y 0.04fF
C29404 POR2X1_274/A POR2X1_325/A 0.05fF
C29405 PAND2X1_629/CTRL2 POR2X1_496/Y 0.06fF
C29406 POR2X1_655/O POR2X1_307/A 0.00fF
C29407 GATE_479 POR2X1_695/Y 0.03fF
C29408 POR2X1_66/B POR2X1_641/CTRL2 0.01fF
C29409 POR2X1_302/Y POR2X1_76/A 0.18fF
C29410 PAND2X1_860/A PAND2X1_175/O 0.04fF
C29411 POR2X1_861/CTRL POR2X1_499/A 0.02fF
C29412 POR2X1_834/a_16_28# POR2X1_330/Y 0.09fF
C29413 PAND2X1_717/A POR2X1_73/Y 0.03fF
C29414 PAND2X1_435/Y PAND2X1_390/Y 0.00fF
C29415 POR2X1_49/Y POR2X1_32/A 0.24fF
C29416 PAND2X1_644/O PAND2X1_643/Y 0.08fF
C29417 PAND2X1_20/A PAND2X1_616/O 0.04fF
C29418 PAND2X1_266/O POR2X1_73/Y 0.05fF
C29419 POR2X1_669/B POR2X1_427/Y 0.07fF
C29420 PAND2X1_217/B POR2X1_102/Y 0.44fF
C29421 POR2X1_666/Y POR2X1_102/Y 0.69fF
C29422 POR2X1_838/B POR2X1_852/B 0.05fF
C29423 POR2X1_32/A PAND2X1_558/CTRL2 0.03fF
C29424 POR2X1_754/Y POR2X1_5/Y 0.07fF
C29425 PAND2X1_52/O PAND2X1_88/Y 0.00fF
C29426 POR2X1_113/m4_208_n4# PAND2X1_96/B 0.17fF
C29427 PAND2X1_48/B PAND2X1_416/O 0.15fF
C29428 POR2X1_66/Y PAND2X1_55/Y 1.49fF
C29429 POR2X1_260/B PAND2X1_753/CTRL 0.00fF
C29430 POR2X1_814/A PAND2X1_111/B 0.05fF
C29431 POR2X1_66/CTRL PAND2X1_96/B 0.05fF
C29432 POR2X1_566/A PAND2X1_93/B 0.03fF
C29433 POR2X1_650/O POR2X1_650/A 0.01fF
C29434 POR2X1_411/B PAND2X1_6/A 0.10fF
C29435 POR2X1_356/A POR2X1_434/O 0.02fF
C29436 POR2X1_175/CTRL PAND2X1_73/Y 0.01fF
C29437 PAND2X1_39/B PAND2X1_744/CTRL 0.01fF
C29438 POR2X1_688/O POR2X1_532/A 0.01fF
C29439 PAND2X1_703/a_76_28# POR2X1_167/Y 0.02fF
C29440 POR2X1_257/A POR2X1_184/Y 0.06fF
C29441 POR2X1_864/a_16_28# POR2X1_750/B 0.03fF
C29442 POR2X1_96/A POR2X1_420/CTRL 0.01fF
C29443 POR2X1_49/Y POR2X1_419/Y 0.04fF
C29444 POR2X1_105/a_16_28# PAND2X1_41/B 0.00fF
C29445 POR2X1_504/Y POR2X1_626/Y 0.06fF
C29446 POR2X1_23/Y POR2X1_372/Y 0.10fF
C29447 PAND2X1_42/CTRL2 PAND2X1_41/B 0.01fF
C29448 POR2X1_65/A POR2X1_829/a_56_344# 0.00fF
C29449 POR2X1_814/B PAND2X1_616/O 0.04fF
C29450 POR2X1_409/B POR2X1_277/CTRL2 0.01fF
C29451 PAND2X1_824/B PAND2X1_234/CTRL 0.01fF
C29452 PAND2X1_16/CTRL2 PAND2X1_41/B 0.03fF
C29453 PAND2X1_651/Y POR2X1_257/A 0.01fF
C29454 PAND2X1_214/O PAND2X1_214/B 0.00fF
C29455 POR2X1_49/Y PAND2X1_576/CTRL2 0.03fF
C29456 PAND2X1_658/CTRL2 POR2X1_376/B 0.06fF
C29457 POR2X1_692/O POR2X1_763/Y 0.06fF
C29458 POR2X1_130/A POR2X1_78/A 0.18fF
C29459 PAND2X1_279/CTRL2 POR2X1_284/B 0.00fF
C29460 PAND2X1_90/A POR2X1_558/B 0.03fF
C29461 POR2X1_63/Y POR2X1_38/Y 1.87fF
C29462 POR2X1_133/O POR2X1_29/A 0.01fF
C29463 POR2X1_342/Y POR2X1_343/Y 0.01fF
C29464 POR2X1_102/Y VDD 2.11fF
C29465 D_INPUT_0 POR2X1_232/CTRL 0.03fF
C29466 PAND2X1_494/CTRL POR2X1_260/B 0.01fF
C29467 PAND2X1_404/A POR2X1_14/Y 0.01fF
C29468 POR2X1_669/Y PAND2X1_720/CTRL 0.01fF
C29469 POR2X1_566/A POR2X1_78/A 0.21fF
C29470 POR2X1_669/B POR2X1_252/CTRL2 0.02fF
C29471 PAND2X1_733/Y POR2X1_40/Y 0.03fF
C29472 PAND2X1_810/B PAND2X1_854/A 0.14fF
C29473 D_INPUT_0 POR2X1_575/B 0.11fF
C29474 POR2X1_632/Y PAND2X1_72/A 0.03fF
C29475 PAND2X1_409/CTRL2 PAND2X1_11/Y 0.01fF
C29476 POR2X1_32/A PAND2X1_553/B 0.03fF
C29477 POR2X1_614/A POR2X1_832/Y 0.16fF
C29478 POR2X1_48/A PAND2X1_649/O 0.15fF
C29479 POR2X1_549/A POR2X1_66/A 0.03fF
C29480 POR2X1_445/A POR2X1_540/CTRL2 0.14fF
C29481 POR2X1_461/Y POR2X1_713/B 0.03fF
C29482 POR2X1_786/A POR2X1_296/B 1.06fF
C29483 PAND2X1_644/Y PAND2X1_794/B 0.02fF
C29484 PAND2X1_436/A VDD 0.00fF
C29485 PAND2X1_65/B POR2X1_807/A 0.00fF
C29486 POR2X1_32/A PAND2X1_303/O 0.08fF
C29487 POR2X1_23/Y POR2X1_253/Y 0.02fF
C29488 POR2X1_423/O POR2X1_293/Y 0.14fF
C29489 POR2X1_451/CTRL POR2X1_635/Y 0.01fF
C29490 PAND2X1_212/B POR2X1_55/Y 0.01fF
C29491 POR2X1_123/O POR2X1_78/A 0.02fF
C29492 POR2X1_87/Y PAND2X1_41/B 0.01fF
C29493 POR2X1_78/B POR2X1_403/CTRL 0.01fF
C29494 POR2X1_644/a_76_344# POR2X1_407/Y 0.00fF
C29495 POR2X1_212/A POR2X1_319/Y 0.27fF
C29496 POR2X1_415/A POR2X1_7/A 0.12fF
C29497 POR2X1_404/B POR2X1_404/CTRL2 0.01fF
C29498 PAND2X1_198/Y POR2X1_40/Y 0.06fF
C29499 POR2X1_634/A PAND2X1_132/CTRL 0.01fF
C29500 PAND2X1_52/B PAND2X1_72/A 5.57fF
C29501 POR2X1_356/A POR2X1_467/Y 0.03fF
C29502 POR2X1_856/B PAND2X1_69/A 0.12fF
C29503 PAND2X1_93/B POR2X1_573/A 0.03fF
C29504 POR2X1_296/Y PAND2X1_55/Y 0.00fF
C29505 PAND2X1_676/O PAND2X1_205/A 0.00fF
C29506 POR2X1_49/Y PAND2X1_35/Y 0.06fF
C29507 POR2X1_671/O POR2X1_5/Y 0.01fF
C29508 PAND2X1_793/Y PAND2X1_185/CTRL 0.01fF
C29509 PAND2X1_307/O POR2X1_56/B 0.02fF
C29510 POR2X1_830/CTRL POR2X1_733/A 0.05fF
C29511 POR2X1_713/A VDD -0.00fF
C29512 POR2X1_66/B POR2X1_334/B 0.08fF
C29513 POR2X1_529/CTRL2 POR2X1_40/Y 0.03fF
C29514 PAND2X1_73/Y POR2X1_713/Y 0.00fF
C29515 PAND2X1_675/A POR2X1_60/A 0.07fF
C29516 POR2X1_83/B POR2X1_433/Y 0.03fF
C29517 POR2X1_16/A PAND2X1_562/Y 0.01fF
C29518 POR2X1_98/O POR2X1_68/B 0.03fF
C29519 POR2X1_78/A POR2X1_844/B 0.03fF
C29520 POR2X1_51/a_76_344# PAND2X1_635/Y 0.00fF
C29521 POR2X1_268/Y POR2X1_55/Y 0.08fF
C29522 POR2X1_78/B POR2X1_608/O 0.01fF
C29523 PAND2X1_236/CTRL INPUT_0 0.01fF
C29524 POR2X1_29/A POR2X1_748/CTRL 0.01fF
C29525 POR2X1_567/A POR2X1_814/A 0.10fF
C29526 POR2X1_296/Y POR2X1_402/A 0.00fF
C29527 PAND2X1_615/a_16_344# D_INPUT_0 0.02fF
C29528 POR2X1_647/CTRL2 POR2X1_101/Y 0.02fF
C29529 POR2X1_13/A PAND2X1_828/O 0.15fF
C29530 POR2X1_141/Y POR2X1_740/Y 0.32fF
C29531 POR2X1_188/A POR2X1_733/A 0.00fF
C29532 POR2X1_817/A POR2X1_5/Y 0.07fF
C29533 PAND2X1_65/B PAND2X1_386/Y 0.00fF
C29534 POR2X1_852/B POR2X1_294/B 0.09fF
C29535 POR2X1_614/A PAND2X1_427/CTRL 0.01fF
C29536 POR2X1_63/Y POR2X1_153/Y 0.05fF
C29537 POR2X1_614/A PAND2X1_230/O 0.03fF
C29538 POR2X1_646/CTRL2 POR2X1_480/A 0.05fF
C29539 POR2X1_45/Y POR2X1_72/B 0.06fF
C29540 PAND2X1_778/Y POR2X1_32/A 0.01fF
C29541 PAND2X1_61/Y POR2X1_55/Y 0.05fF
C29542 POR2X1_71/Y POR2X1_5/Y 0.01fF
C29543 POR2X1_840/B POR2X1_121/B 0.01fF
C29544 POR2X1_844/CTRL POR2X1_590/A 0.11fF
C29545 PAND2X1_658/A PAND2X1_658/a_16_344# 0.02fF
C29546 POR2X1_614/A PAND2X1_279/O 0.07fF
C29547 PAND2X1_802/O POR2X1_760/A 0.02fF
C29548 POR2X1_664/Y PAND2X1_387/O 0.02fF
C29549 POR2X1_222/Y POR2X1_186/Y 0.12fF
C29550 POR2X1_83/CTRL2 POR2X1_23/Y 0.01fF
C29551 POR2X1_683/O POR2X1_236/Y 0.03fF
C29552 POR2X1_16/A POR2X1_437/O 0.15fF
C29553 POR2X1_143/O POR2X1_236/Y 0.02fF
C29554 POR2X1_66/B POR2X1_124/B 6.48fF
C29555 PAND2X1_630/a_16_344# POR2X1_748/A 0.04fF
C29556 PAND2X1_682/O POR2X1_750/B 0.02fF
C29557 PAND2X1_809/B PAND2X1_809/CTRL 0.01fF
C29558 PAND2X1_95/B PAND2X1_18/CTRL2 0.01fF
C29559 POR2X1_502/A POR2X1_459/CTRL 0.01fF
C29560 POR2X1_407/A POR2X1_777/B 0.03fF
C29561 POR2X1_114/B PAND2X1_299/CTRL 0.01fF
C29562 POR2X1_368/CTRL2 POR2X1_372/Y 0.05fF
C29563 PAND2X1_391/a_76_28# POR2X1_382/Y 0.04fF
C29564 POR2X1_65/A PAND2X1_242/O 0.01fF
C29565 PAND2X1_3/A PAND2X1_1/O 0.01fF
C29566 POR2X1_5/Y POR2X1_42/Y 0.13fF
C29567 POR2X1_346/O PAND2X1_58/A 0.17fF
C29568 D_INPUT_1 POR2X1_750/A 0.06fF
C29569 PAND2X1_659/CTRL2 POR2X1_494/Y 0.00fF
C29570 POR2X1_88/Y PAND2X1_350/A 0.01fF
C29571 INPUT_1 POR2X1_28/O 0.18fF
C29572 POR2X1_378/A POR2X1_296/B 0.00fF
C29573 POR2X1_76/Y POR2X1_220/Y 0.07fF
C29574 PAND2X1_778/O POR2X1_55/Y 0.01fF
C29575 POR2X1_407/A POR2X1_660/A 0.03fF
C29576 PAND2X1_420/a_76_28# PAND2X1_96/B 0.02fF
C29577 PAND2X1_216/O INPUT_0 0.02fF
C29578 POR2X1_65/A POR2X1_518/Y 0.01fF
C29579 POR2X1_502/A POR2X1_651/CTRL2 0.01fF
C29580 POR2X1_49/Y PAND2X1_651/Y 0.08fF
C29581 PAND2X1_454/a_76_28# POR2X1_376/B 0.02fF
C29582 POR2X1_114/B POR2X1_475/A 0.03fF
C29583 POR2X1_681/CTRL2 POR2X1_39/B 0.03fF
C29584 POR2X1_119/Y POR2X1_411/B 0.76fF
C29585 PAND2X1_498/O VDD 0.00fF
C29586 POR2X1_700/CTRL VDD 0.00fF
C29587 PAND2X1_612/B POR2X1_774/A 0.29fF
C29588 POR2X1_862/A POR2X1_559/A 0.03fF
C29589 POR2X1_376/B PAND2X1_6/A 0.26fF
C29590 POR2X1_217/O POR2X1_572/B 0.01fF
C29591 POR2X1_356/A POR2X1_570/O 0.04fF
C29592 POR2X1_407/A PAND2X1_65/B 2.20fF
C29593 POR2X1_68/A POR2X1_855/A 0.00fF
C29594 POR2X1_96/A POR2X1_56/B 0.02fF
C29595 POR2X1_315/Y PAND2X1_443/Y 0.02fF
C29596 POR2X1_78/B POR2X1_341/CTRL 0.19fF
C29597 PAND2X1_808/Y VDD 0.14fF
C29598 POR2X1_186/Y POR2X1_532/A 0.08fF
C29599 POR2X1_742/O POR2X1_741/Y 0.04fF
C29600 PAND2X1_824/B POR2X1_856/B 0.20fF
C29601 POR2X1_96/Y PAND2X1_98/O 0.00fF
C29602 POR2X1_441/Y PAND2X1_326/B 0.03fF
C29603 POR2X1_41/B POR2X1_763/Y 0.03fF
C29604 POR2X1_16/A PAND2X1_722/O 0.03fF
C29605 POR2X1_49/Y PAND2X1_844/B 1.65fF
C29606 POR2X1_525/Y POR2X1_46/Y 0.12fF
C29607 PAND2X1_651/A POR2X1_14/Y 0.02fF
C29608 PAND2X1_69/A POR2X1_786/CTRL2 0.00fF
C29609 POR2X1_502/A POR2X1_662/Y 0.00fF
C29610 POR2X1_41/B PAND2X1_115/B 0.21fF
C29611 POR2X1_40/Y PAND2X1_168/O 0.04fF
C29612 PAND2X1_674/O VDD 0.00fF
C29613 POR2X1_555/A PAND2X1_96/B 0.10fF
C29614 PAND2X1_467/Y POR2X1_83/B 0.03fF
C29615 POR2X1_37/Y PAND2X1_100/a_76_28# 0.01fF
C29616 D_GATE_662 PAND2X1_438/CTRL2 0.00fF
C29617 POR2X1_220/Y POR2X1_740/Y 0.03fF
C29618 POR2X1_52/A PAND2X1_215/B 0.02fF
C29619 PAND2X1_96/B POR2X1_563/CTRL2 0.04fF
C29620 PAND2X1_48/B PAND2X1_372/O 0.08fF
C29621 POR2X1_231/CTRL POR2X1_785/A 0.07fF
C29622 POR2X1_717/O POR2X1_814/B 0.01fF
C29623 PAND2X1_218/a_16_344# INPUT_0 0.01fF
C29624 POR2X1_81/a_76_344# PAND2X1_510/B -0.00fF
C29625 PAND2X1_661/B PAND2X1_828/O 0.02fF
C29626 PAND2X1_845/CTRL VDD 0.00fF
C29627 POR2X1_573/CTRL POR2X1_573/A 0.01fF
C29628 POR2X1_150/Y POR2X1_39/B 0.10fF
C29629 PAND2X1_714/A POR2X1_142/Y 0.07fF
C29630 PAND2X1_388/Y PAND2X1_562/B 0.07fF
C29631 POR2X1_78/B POR2X1_194/CTRL2 0.01fF
C29632 POR2X1_78/B POR2X1_644/A 0.03fF
C29633 PAND2X1_6/Y POR2X1_244/B 0.06fF
C29634 POR2X1_650/A POR2X1_493/O 0.01fF
C29635 POR2X1_448/Y PAND2X1_60/B 0.01fF
C29636 POR2X1_40/Y PAND2X1_550/B 0.03fF
C29637 PAND2X1_139/O PAND2X1_349/A 0.02fF
C29638 PAND2X1_73/Y POR2X1_559/A 0.10fF
C29639 PAND2X1_564/CTRL POR2X1_73/Y 0.08fF
C29640 POR2X1_483/B POR2X1_556/Y 0.01fF
C29641 PAND2X1_149/O PAND2X1_148/Y 0.01fF
C29642 POR2X1_853/A POR2X1_785/A 0.00fF
C29643 POR2X1_3/A POR2X1_25/O 0.36fF
C29644 POR2X1_821/Y VDD 0.08fF
C29645 PAND2X1_94/A POR2X1_750/B 0.03fF
C29646 POR2X1_52/A PAND2X1_6/A 0.13fF
C29647 POR2X1_87/B PAND2X1_32/a_16_344# 0.03fF
C29648 POR2X1_673/A PAND2X1_4/O 0.04fF
C29649 POR2X1_65/A POR2X1_527/Y 0.03fF
C29650 POR2X1_614/A POR2X1_307/Y 0.03fF
C29651 POR2X1_785/CTRL PAND2X1_32/B 0.03fF
C29652 PAND2X1_69/A POR2X1_722/Y 0.03fF
C29653 POR2X1_257/A POR2X1_524/a_16_28# 0.03fF
C29654 PAND2X1_803/Y PAND2X1_347/Y 0.01fF
C29655 PAND2X1_472/a_76_28# POR2X1_83/B 0.02fF
C29656 POR2X1_351/Y POR2X1_857/B 0.03fF
C29657 POR2X1_60/O POR2X1_13/A 0.01fF
C29658 PAND2X1_90/Y POR2X1_758/m4_208_n4# 0.12fF
C29659 POR2X1_488/Y PAND2X1_794/B 0.00fF
C29660 INPUT_0 POR2X1_597/CTRL 0.06fF
C29661 POR2X1_65/A POR2X1_83/CTRL 0.02fF
C29662 POR2X1_41/B POR2X1_73/Y 0.23fF
C29663 POR2X1_322/Y PAND2X1_556/B 0.03fF
C29664 POR2X1_409/B POR2X1_4/Y 0.07fF
C29665 POR2X1_294/B PAND2X1_504/a_16_344# 0.01fF
C29666 POR2X1_330/Y POR2X1_507/A 0.07fF
C29667 PAND2X1_72/O POR2X1_579/Y 0.00fF
C29668 PAND2X1_820/O POR2X1_847/B 0.01fF
C29669 PAND2X1_96/B PAND2X1_89/O 0.04fF
C29670 POR2X1_55/Y PAND2X1_548/CTRL2 0.01fF
C29671 PAND2X1_834/a_16_344# PAND2X1_349/A 0.00fF
C29672 POR2X1_66/A POR2X1_542/Y 0.01fF
C29673 POR2X1_13/A PAND2X1_388/Y 0.03fF
C29674 PAND2X1_90/A POR2X1_243/CTRL 0.01fF
C29675 PAND2X1_799/a_16_344# INPUT_0 0.00fF
C29676 POR2X1_516/Y PAND2X1_657/B 0.04fF
C29677 POR2X1_61/Y POR2X1_260/A 0.10fF
C29678 PAND2X1_490/CTRL POR2X1_334/B 0.01fF
C29679 PAND2X1_687/CTRL2 POR2X1_60/A 0.01fF
C29680 POR2X1_48/A POR2X1_524/O 0.02fF
C29681 PAND2X1_341/A PAND2X1_197/CTRL 0.01fF
C29682 PAND2X1_63/B PAND2X1_8/Y 0.04fF
C29683 POR2X1_334/A POR2X1_99/A 0.02fF
C29684 POR2X1_32/A PAND2X1_865/A 0.01fF
C29685 POR2X1_618/a_56_344# POR2X1_38/B 0.01fF
C29686 PAND2X1_41/B POR2X1_352/a_16_28# 0.03fF
C29687 PAND2X1_775/CTRL POR2X1_91/Y 0.01fF
C29688 POR2X1_13/A PAND2X1_720/CTRL2 0.01fF
C29689 POR2X1_335/O POR2X1_337/A 0.03fF
C29690 POR2X1_796/A VDD 0.27fF
C29691 POR2X1_13/A PAND2X1_549/B 0.03fF
C29692 PAND2X1_658/A PAND2X1_548/O 0.02fF
C29693 PAND2X1_44/CTRL PAND2X1_18/B 0.01fF
C29694 POR2X1_483/a_16_28# POR2X1_228/Y 0.03fF
C29695 PAND2X1_569/Y VDD 0.38fF
C29696 POR2X1_237/CTRL2 PAND2X1_308/Y 0.01fF
C29697 PAND2X1_563/A POR2X1_106/Y 0.18fF
C29698 POR2X1_517/CTRL POR2X1_669/B 0.02fF
C29699 POR2X1_283/A POR2X1_46/Y 0.10fF
C29700 POR2X1_570/O POR2X1_569/A 0.04fF
C29701 POR2X1_554/Y POR2X1_510/Y 0.04fF
C29702 PAND2X1_480/B PAND2X1_112/CTRL 0.27fF
C29703 POR2X1_493/O POR2X1_294/B 0.23fF
C29704 POR2X1_619/A POR2X1_619/CTRL2 0.01fF
C29705 POR2X1_559/CTRL2 POR2X1_68/B 0.01fF
C29706 POR2X1_56/B POR2X1_7/A 0.10fF
C29707 POR2X1_614/A PAND2X1_72/O 0.01fF
C29708 PAND2X1_96/B PAND2X1_316/O 0.15fF
C29709 POR2X1_52/A POR2X1_588/Y 0.03fF
C29710 POR2X1_57/A PAND2X1_798/B 0.07fF
C29711 POR2X1_41/B PAND2X1_244/B 0.05fF
C29712 POR2X1_440/Y POR2X1_468/B 0.03fF
C29713 POR2X1_16/A POR2X1_821/O 0.06fF
C29714 POR2X1_523/Y PAND2X1_521/CTRL2 0.01fF
C29715 POR2X1_750/B PAND2X1_680/CTRL2 0.01fF
C29716 POR2X1_447/B POR2X1_202/CTRL 0.18fF
C29717 PAND2X1_17/a_56_28# INPUT_6 0.00fF
C29718 PAND2X1_623/Y POR2X1_283/A 0.03fF
C29719 POR2X1_614/A POR2X1_68/B 0.10fF
C29720 PAND2X1_84/CTRL POR2X1_394/A 0.08fF
C29721 POR2X1_65/A PAND2X1_325/O 0.01fF
C29722 POR2X1_730/Y POR2X1_355/B 0.03fF
C29723 POR2X1_403/CTRL POR2X1_294/A 0.01fF
C29724 POR2X1_96/A PAND2X1_356/a_76_28# 0.01fF
C29725 POR2X1_198/B POR2X1_201/Y 0.01fF
C29726 POR2X1_259/CTRL2 POR2X1_785/A 0.09fF
C29727 POR2X1_165/Y VDD 0.03fF
C29728 POR2X1_740/A POR2X1_738/Y 0.00fF
C29729 POR2X1_177/O POR2X1_236/Y 0.01fF
C29730 POR2X1_316/CTRL2 POR2X1_13/A 0.03fF
C29731 POR2X1_566/A PAND2X1_313/a_16_344# 0.05fF
C29732 POR2X1_680/Y PAND2X1_728/O 0.15fF
C29733 POR2X1_567/A POR2X1_852/B 0.10fF
C29734 POR2X1_71/Y PAND2X1_574/a_16_344# 0.01fF
C29735 POR2X1_38/B POR2X1_68/B 0.54fF
C29736 PAND2X1_4/O D_INPUT_1 0.08fF
C29737 INPUT_0 POR2X1_558/Y 0.04fF
C29738 PAND2X1_840/A POR2X1_283/A 0.24fF
C29739 PAND2X1_213/Y POR2X1_90/Y 0.04fF
C29740 PAND2X1_30/CTRL2 POR2X1_635/A 0.05fF
C29741 POR2X1_119/Y POR2X1_376/B 0.07fF
C29742 POR2X1_346/O PAND2X1_96/B 0.01fF
C29743 PAND2X1_354/Y VDD 0.06fF
C29744 PAND2X1_57/B PAND2X1_142/CTRL 0.01fF
C29745 POR2X1_121/B PAND2X1_56/A 0.03fF
C29746 POR2X1_574/Y PAND2X1_516/O 0.02fF
C29747 PAND2X1_126/CTRL2 PAND2X1_69/A 0.01fF
C29748 POR2X1_52/A POR2X1_583/Y 0.00fF
C29749 INPUT_0 PAND2X1_851/CTRL2 0.09fF
C29750 POR2X1_608/O POR2X1_294/A 0.02fF
C29751 PAND2X1_587/Y PAND2X1_18/B 0.06fF
C29752 PAND2X1_642/B PAND2X1_559/O 0.06fF
C29753 POR2X1_447/B PAND2X1_627/O 0.03fF
C29754 PAND2X1_69/A POR2X1_391/O 0.01fF
C29755 POR2X1_36/B INPUT_6 0.46fF
C29756 POR2X1_383/A POR2X1_840/B 0.14fF
C29757 POR2X1_784/CTRL2 POR2X1_725/Y 0.03fF
C29758 D_INPUT_6 POR2X1_1/CTRL 0.01fF
C29759 POR2X1_76/B POR2X1_274/CTRL2 0.00fF
C29760 POR2X1_35/Y POR2X1_260/A 0.03fF
C29761 POR2X1_68/A POR2X1_675/Y 0.05fF
C29762 PAND2X1_641/CTRL PAND2X1_651/Y 0.24fF
C29763 PAND2X1_775/CTRL POR2X1_109/Y 0.01fF
C29764 PAND2X1_605/CTRL2 POR2X1_73/Y 0.03fF
C29765 PAND2X1_658/A PAND2X1_861/a_76_28# 0.01fF
C29766 PAND2X1_659/Y PAND2X1_205/B 0.03fF
C29767 POR2X1_846/B POR2X1_129/Y 0.00fF
C29768 POR2X1_467/Y PAND2X1_72/A 0.03fF
C29769 PAND2X1_75/CTRL2 POR2X1_624/Y 0.10fF
C29770 POR2X1_383/A PAND2X1_824/CTRL 0.01fF
C29771 PAND2X1_297/O POR2X1_68/B 0.04fF
C29772 POR2X1_57/A PAND2X1_691/Y 0.03fF
C29773 PAND2X1_671/a_76_28# PAND2X1_6/A 0.01fF
C29774 POR2X1_52/A POR2X1_119/Y 0.11fF
C29775 PAND2X1_642/a_16_344# PAND2X1_642/B 0.03fF
C29776 PAND2X1_651/a_56_28# POR2X1_43/B 0.00fF
C29777 POR2X1_162/Y PAND2X1_158/O 0.02fF
C29778 POR2X1_632/A POR2X1_632/Y 0.01fF
C29779 PAND2X1_493/CTRL POR2X1_599/A 0.05fF
C29780 POR2X1_416/B PAND2X1_540/a_76_28# 0.02fF
C29781 POR2X1_149/A POR2X1_863/A 0.01fF
C29782 PAND2X1_242/Y POR2X1_423/O 0.01fF
C29783 VDD POR2X1_761/A 0.05fF
C29784 POR2X1_235/O PAND2X1_63/B 0.00fF
C29785 POR2X1_335/B POR2X1_260/A 0.00fF
C29786 PAND2X1_308/Y POR2X1_73/Y 0.03fF
C29787 POR2X1_119/Y PAND2X1_398/CTRL2 0.01fF
C29788 POR2X1_662/Y POR2X1_188/Y 0.03fF
C29789 POR2X1_119/Y POR2X1_152/A 0.03fF
C29790 POR2X1_760/A PAND2X1_222/A 0.03fF
C29791 POR2X1_265/Y POR2X1_43/B 0.05fF
C29792 POR2X1_579/B POR2X1_702/A 0.16fF
C29793 POR2X1_714/CTRL POR2X1_703/Y 0.01fF
C29794 POR2X1_366/O POR2X1_383/A 0.01fF
C29795 POR2X1_537/Y PAND2X1_536/O 0.02fF
C29796 POR2X1_643/CTRL POR2X1_590/A 0.01fF
C29797 POR2X1_661/A POR2X1_121/B 0.08fF
C29798 POR2X1_467/Y POR2X1_535/O 0.01fF
C29799 POR2X1_244/B POR2X1_632/Y 0.03fF
C29800 POR2X1_176/CTRL POR2X1_90/Y 0.07fF
C29801 POR2X1_668/Y POR2X1_39/B 0.03fF
C29802 PAND2X1_55/Y PAND2X1_304/CTRL2 0.03fF
C29803 PAND2X1_846/CTRL INPUT_0 0.30fF
C29804 POR2X1_539/A POR2X1_703/A 0.03fF
C29805 PAND2X1_6/Y POR2X1_537/Y 0.03fF
C29806 POR2X1_123/A POR2X1_260/A 0.03fF
C29807 POR2X1_96/A POR2X1_184/a_16_28# 0.02fF
C29808 POR2X1_145/Y POR2X1_394/A 0.00fF
C29809 POR2X1_840/B PAND2X1_71/Y 0.03fF
C29810 PAND2X1_765/O POR2X1_260/A 0.04fF
C29811 POR2X1_644/A POR2X1_294/A 0.07fF
C29812 POR2X1_394/A POR2X1_757/O 0.03fF
C29813 POR2X1_8/Y POR2X1_384/O 0.16fF
C29814 POR2X1_614/A PAND2X1_143/O 0.05fF
C29815 PAND2X1_472/A POR2X1_397/a_16_28# 0.03fF
C29816 VDD POR2X1_173/O 0.00fF
C29817 POR2X1_244/B PAND2X1_52/B 0.04fF
C29818 POR2X1_763/Y POR2X1_77/Y 0.07fF
C29819 POR2X1_458/Y POR2X1_457/CTRL2 0.04fF
C29820 PAND2X1_217/B POR2X1_677/Y 0.05fF
C29821 POR2X1_485/Y POR2X1_23/Y 0.06fF
C29822 POR2X1_66/B PAND2X1_257/a_16_344# 0.02fF
C29823 PAND2X1_115/B POR2X1_77/Y 0.01fF
C29824 POR2X1_48/A POR2X1_150/Y 0.03fF
C29825 PAND2X1_602/Y POR2X1_533/Y 0.00fF
C29826 POR2X1_8/Y POR2X1_10/CTRL 0.01fF
C29827 POR2X1_368/Y POR2X1_316/Y 0.16fF
C29828 PAND2X1_860/A PAND2X1_76/Y 0.03fF
C29829 POR2X1_568/Y POR2X1_545/m4_208_n4# 0.06fF
C29830 POR2X1_564/B POR2X1_180/A 0.03fF
C29831 POR2X1_863/A VDD 1.18fF
C29832 PAND2X1_658/A POR2X1_77/Y 0.03fF
C29833 POR2X1_416/B POR2X1_232/a_16_28# 0.01fF
C29834 PAND2X1_308/Y PAND2X1_727/O 0.01fF
C29835 POR2X1_25/Y POR2X1_51/B 0.33fF
C29836 PAND2X1_95/B PAND2X1_72/A 0.03fF
C29837 PAND2X1_850/Y POR2X1_91/Y 0.07fF
C29838 PAND2X1_220/A POR2X1_20/B 0.01fF
C29839 POR2X1_8/Y POR2X1_749/O 0.20fF
C29840 PAND2X1_117/a_56_28# PAND2X1_72/A 0.00fF
C29841 POR2X1_365/A POR2X1_365/a_16_28# 0.03fF
C29842 POR2X1_86/CTRL PAND2X1_338/B 0.00fF
C29843 POR2X1_677/Y VDD 0.34fF
C29844 POR2X1_416/B POR2X1_90/Y 0.20fF
C29845 POR2X1_294/B POR2X1_535/CTRL2 0.01fF
C29846 POR2X1_793/A PAND2X1_52/B 0.38fF
C29847 POR2X1_73/Y POR2X1_77/Y 0.44fF
C29848 POR2X1_546/CTRL POR2X1_550/B 0.00fF
C29849 POR2X1_814/A POR2X1_807/A 0.05fF
C29850 POR2X1_60/A POR2X1_262/Y 0.12fF
C29851 POR2X1_9/Y VDD 4.68fF
C29852 POR2X1_85/Y POR2X1_73/Y 1.20fF
C29853 PAND2X1_632/A PAND2X1_508/B 0.01fF
C29854 POR2X1_274/A POR2X1_274/CTRL 0.04fF
C29855 PAND2X1_484/a_16_344# POR2X1_559/A 0.12fF
C29856 PAND2X1_802/O PAND2X1_802/B 0.00fF
C29857 PAND2X1_94/A PAND2X1_122/CTRL 0.13fF
C29858 POR2X1_20/B PAND2X1_718/Y 0.00fF
C29859 POR2X1_571/O POR2X1_561/Y 0.12fF
C29860 POR2X1_41/B PAND2X1_458/CTRL2 0.02fF
C29861 POR2X1_832/A POR2X1_711/Y -0.02fF
C29862 POR2X1_67/Y POR2X1_668/m4_208_n4# 0.08fF
C29863 PAND2X1_91/a_56_28# POR2X1_97/A 0.00fF
C29864 POR2X1_334/Y POR2X1_97/B 0.04fF
C29865 POR2X1_311/Y PAND2X1_222/O 0.17fF
C29866 POR2X1_333/A POR2X1_212/A 0.50fF
C29867 POR2X1_54/Y POR2X1_23/a_16_28# 0.03fF
C29868 POR2X1_311/Y PAND2X1_222/A 1.23fF
C29869 POR2X1_832/Y POR2X1_590/A 0.03fF
C29870 POR2X1_383/A PAND2X1_56/A 0.26fF
C29871 POR2X1_220/A POR2X1_161/O 0.01fF
C29872 POR2X1_323/CTRL POR2X1_485/Y 0.01fF
C29873 PAND2X1_56/Y POR2X1_661/A 0.07fF
C29874 POR2X1_394/A POR2X1_701/a_16_28# 0.03fF
C29875 PAND2X1_717/A PAND2X1_785/Y 0.16fF
C29876 POR2X1_863/A PAND2X1_32/B 0.17fF
C29877 POR2X1_85/Y PAND2X1_244/B 0.03fF
C29878 POR2X1_811/CTRL2 PAND2X1_73/Y 0.01fF
C29879 PAND2X1_35/A POR2X1_27/Y 0.12fF
C29880 POR2X1_590/Y PAND2X1_304/a_56_28# 0.00fF
C29881 POR2X1_390/B POR2X1_343/Y 0.05fF
C29882 POR2X1_250/Y POR2X1_79/Y 0.03fF
C29883 POR2X1_849/A POR2X1_29/A 0.00fF
C29884 PAND2X1_862/Y PAND2X1_865/Y 0.01fF
C29885 POR2X1_532/A PAND2X1_146/CTRL 0.01fF
C29886 POR2X1_719/A PAND2X1_93/B 0.07fF
C29887 POR2X1_808/A POR2X1_808/O 0.07fF
C29888 POR2X1_836/O POR2X1_836/B 0.00fF
C29889 PAND2X1_865/Y POR2X1_385/Y 0.10fF
C29890 PAND2X1_373/a_16_344# PAND2X1_72/A 0.02fF
C29891 POR2X1_276/B POR2X1_325/A 0.07fF
C29892 POR2X1_20/B PAND2X1_580/B 0.03fF
C29893 PAND2X1_172/a_16_344# PAND2X1_52/B 0.01fF
C29894 PAND2X1_60/B POR2X1_303/B 0.03fF
C29895 POR2X1_153/O POR2X1_77/Y 0.07fF
C29896 POR2X1_174/CTRL PAND2X1_72/A 0.00fF
C29897 POR2X1_709/A POR2X1_410/CTRL 0.01fF
C29898 POR2X1_56/a_76_344# POR2X1_496/Y 0.03fF
C29899 PAND2X1_714/B PAND2X1_326/B 0.00fF
C29900 PAND2X1_23/Y PAND2X1_75/O 0.18fF
C29901 POR2X1_78/A POR2X1_241/B 0.26fF
C29902 PAND2X1_9/CTRL POR2X1_29/A 0.01fF
C29903 POR2X1_257/A POR2X1_256/CTRL2 0.01fF
C29904 POR2X1_337/Y PAND2X1_179/O 0.23fF
C29905 POR2X1_734/B POR2X1_734/A 0.03fF
C29906 PAND2X1_469/CTRL POR2X1_236/Y 0.01fF
C29907 PAND2X1_601/a_16_344# PAND2X1_65/B 0.01fF
C29908 POR2X1_89/CTRL POR2X1_5/Y 0.04fF
C29909 POR2X1_416/B PAND2X1_360/Y 0.03fF
C29910 POR2X1_20/B POR2X1_233/O 0.01fF
C29911 POR2X1_96/A PAND2X1_267/B 0.02fF
C29912 PAND2X1_231/CTRL2 D_INPUT_0 0.01fF
C29913 POR2X1_465/CTRL POR2X1_563/Y 0.01fF
C29914 POR2X1_407/A POR2X1_814/A 0.48fF
C29915 POR2X1_260/B POR2X1_362/B 0.03fF
C29916 POR2X1_13/A PAND2X1_98/a_16_344# 0.02fF
C29917 POR2X1_629/a_76_344# POR2X1_186/Y 0.01fF
C29918 POR2X1_315/O PAND2X1_717/A 0.07fF
C29919 POR2X1_243/B VDD 0.06fF
C29920 POR2X1_99/Y VDD 0.00fF
C29921 POR2X1_383/A POR2X1_661/A 0.07fF
C29922 D_INPUT_0 PAND2X1_41/B 0.03fF
C29923 POR2X1_220/B POR2X1_186/Y 0.03fF
C29924 POR2X1_801/B POR2X1_750/B 1.76fF
C29925 POR2X1_32/A PAND2X1_706/CTRL 0.01fF
C29926 POR2X1_467/Y POR2X1_448/CTRL 0.01fF
C29927 POR2X1_828/a_16_28# POR2X1_828/A 0.03fF
C29928 POR2X1_274/A VDD 0.51fF
C29929 POR2X1_110/Y POR2X1_416/B 0.06fF
C29930 POR2X1_540/Y POR2X1_736/A 0.05fF
C29931 PAND2X1_11/Y POR2X1_750/B 0.03fF
C29932 POR2X1_23/Y POR2X1_29/O 0.01fF
C29933 POR2X1_632/A POR2X1_632/a_16_28# 0.05fF
C29934 POR2X1_83/B POR2X1_698/CTRL 0.01fF
C29935 POR2X1_416/Y PAND2X1_634/CTRL 0.01fF
C29936 POR2X1_427/CTRL2 POR2X1_236/Y 0.00fF
C29937 POR2X1_644/CTRL2 POR2X1_513/B 0.01fF
C29938 PAND2X1_545/CTRL POR2X1_40/Y 0.01fF
C29939 POR2X1_48/A PAND2X1_553/A 0.01fF
C29940 PAND2X1_9/O POR2X1_94/A 0.07fF
C29941 POR2X1_554/B POR2X1_112/Y 0.05fF
C29942 POR2X1_138/CTRL POR2X1_624/Y 0.05fF
C29943 PAND2X1_307/CTRL POR2X1_40/Y 0.02fF
C29944 POR2X1_67/A POR2X1_5/Y 1.28fF
C29945 POR2X1_454/A POR2X1_555/a_16_28# 0.07fF
C29946 PAND2X1_213/O PAND2X1_213/A 0.01fF
C29947 PAND2X1_10/CTRL2 PAND2X1_8/Y 0.03fF
C29948 PAND2X1_217/O POR2X1_599/A 0.24fF
C29949 PAND2X1_594/a_16_344# PAND2X1_90/Y 0.07fF
C29950 POR2X1_485/Y PAND2X1_565/a_16_344# 0.02fF
C29951 POR2X1_66/B POR2X1_752/Y 0.03fF
C29952 PAND2X1_474/a_16_344# POR2X1_43/B 0.01fF
C29953 POR2X1_60/A PAND2X1_185/a_16_344# 0.01fF
C29954 POR2X1_27/CTRL PAND2X1_63/B 0.01fF
C29955 POR2X1_864/A POR2X1_407/Y 0.00fF
C29956 POR2X1_502/A POR2X1_444/A 0.03fF
C29957 POR2X1_226/O POR2X1_5/Y 0.07fF
C29958 INPUT_3 POR2X1_409/CTRL2 0.17fF
C29959 PAND2X1_39/B POR2X1_249/CTRL 0.01fF
C29960 POR2X1_504/CTRL2 POR2X1_846/A 0.00fF
C29961 POR2X1_49/Y PAND2X1_731/B 0.05fF
C29962 POR2X1_614/A PAND2X1_761/O 0.01fF
C29963 PAND2X1_296/CTRL PAND2X1_347/Y 0.01fF
C29964 PAND2X1_77/CTRL2 PAND2X1_8/Y 0.01fF
C29965 PAND2X1_318/m4_208_n4# POR2X1_299/m4_208_n4# 0.13fF
C29966 POR2X1_286/B POR2X1_649/CTRL 0.01fF
C29967 POR2X1_602/A VDD 0.00fF
C29968 PAND2X1_638/B VDD 0.05fF
C29969 POR2X1_114/B PAND2X1_406/CTRL 0.03fF
C29970 POR2X1_83/B PAND2X1_556/B 0.02fF
C29971 POR2X1_97/A POR2X1_853/O 0.01fF
C29972 POR2X1_555/A POR2X1_355/A 0.01fF
C29973 PAND2X1_751/CTRL2 POR2X1_590/A 0.03fF
C29974 PAND2X1_39/B POR2X1_784/O 0.01fF
C29975 PAND2X1_124/Y POR2X1_599/A 0.36fF
C29976 PAND2X1_467/B PAND2X1_707/CTRL2 0.01fF
C29977 POR2X1_276/CTRL POR2X1_218/Y 0.02fF
C29978 POR2X1_43/B POR2X1_848/A 0.07fF
C29979 POR2X1_415/A POR2X1_38/Y 0.89fF
C29980 POR2X1_43/B PAND2X1_776/Y 0.02fF
C29981 POR2X1_79/Y PAND2X1_798/O 0.00fF
C29982 PAND2X1_210/O PAND2X1_725/Y 0.00fF
C29983 POR2X1_23/Y PAND2X1_339/Y 0.03fF
C29984 POR2X1_848/A POR2X1_789/A 0.07fF
C29985 PAND2X1_90/Y PAND2X1_41/B 0.55fF
C29986 POR2X1_447/CTRL2 POR2X1_447/A 0.01fF
C29987 POR2X1_760/A PAND2X1_537/CTRL 0.01fF
C29988 POR2X1_285/B PAND2X1_52/B 0.01fF
C29989 POR2X1_65/A PAND2X1_803/A 0.03fF
C29990 PAND2X1_651/Y POR2X1_613/CTRL 0.00fF
C29991 POR2X1_20/B PAND2X1_349/A 0.03fF
C29992 PAND2X1_254/Y POR2X1_83/B 0.03fF
C29993 POR2X1_186/Y POR2X1_742/CTRL 0.01fF
C29994 PAND2X1_594/CTRL POR2X1_740/Y 0.00fF
C29995 POR2X1_423/Y POR2X1_236/Y 0.10fF
C29996 PAND2X1_717/A PAND2X1_348/A 0.07fF
C29997 PAND2X1_73/Y POR2X1_783/B 0.02fF
C29998 POR2X1_20/B PAND2X1_63/B 0.01fF
C29999 PAND2X1_267/B POR2X1_7/A 0.04fF
C30000 D_INPUT_0 POR2X1_130/Y 0.07fF
C30001 POR2X1_674/a_76_344# PAND2X1_652/A 0.03fF
C30002 POR2X1_388/CTRL PAND2X1_93/B 0.00fF
C30003 POR2X1_96/A PAND2X1_772/a_16_344# 0.02fF
C30004 POR2X1_195/A PAND2X1_69/A 0.01fF
C30005 POR2X1_52/A POR2X1_497/CTRL 0.01fF
C30006 PAND2X1_95/B PAND2X1_752/O 0.06fF
C30007 POR2X1_502/A POR2X1_830/a_56_344# 0.00fF
C30008 POR2X1_602/B PAND2X1_57/B 0.03fF
C30009 POR2X1_278/Y PAND2X1_217/B 0.10fF
C30010 POR2X1_456/CTRL VDD -0.00fF
C30011 POR2X1_596/A POR2X1_644/a_16_28# 0.02fF
C30012 POR2X1_859/A POR2X1_752/Y 0.02fF
C30013 PAND2X1_48/Y VDD 0.25fF
C30014 D_INPUT_0 PAND2X1_744/m4_208_n4# 0.12fF
C30015 GATE_741 PAND2X1_363/Y 0.02fF
C30016 POR2X1_483/A PAND2X1_48/CTRL2 0.01fF
C30017 PAND2X1_230/CTRL2 POR2X1_795/B 0.04fF
C30018 PAND2X1_479/CTRL PAND2X1_480/B 0.00fF
C30019 POR2X1_825/CTRL2 POR2X1_42/Y 0.01fF
C30020 POR2X1_102/Y PAND2X1_717/O 0.03fF
C30021 POR2X1_556/A POR2X1_787/a_76_344# 0.00fF
C30022 POR2X1_505/O POR2X1_20/B 0.01fF
C30023 POR2X1_83/B POR2X1_599/A 0.05fF
C30024 POR2X1_52/A POR2X1_290/CTRL2 0.01fF
C30025 POR2X1_719/CTRL PAND2X1_93/B -0.01fF
C30026 PAND2X1_205/Y POR2X1_79/Y 0.01fF
C30027 POR2X1_40/Y PAND2X1_506/CTRL2 0.01fF
C30028 POR2X1_250/Y PAND2X1_730/A 0.03fF
C30029 PAND2X1_467/B PAND2X1_725/A 0.00fF
C30030 POR2X1_278/CTRL PAND2X1_35/Y 0.01fF
C30031 PAND2X1_381/Y PAND2X1_69/A 0.03fF
C30032 POR2X1_68/A POR2X1_14/Y 0.03fF
C30033 PAND2X1_39/B POR2X1_456/B 1.26fF
C30034 POR2X1_294/CTRL2 POR2X1_260/A 0.03fF
C30035 PAND2X1_848/A POR2X1_750/A 0.00fF
C30036 PAND2X1_73/Y PAND2X1_519/a_56_28# 0.00fF
C30037 INPUT_1 POR2X1_415/A 0.13fF
C30038 PAND2X1_854/a_76_28# POR2X1_102/Y 0.01fF
C30039 POR2X1_833/A POR2X1_341/A 0.12fF
C30040 POR2X1_208/A PAND2X1_93/B 0.01fF
C30041 PAND2X1_198/Y POR2X1_5/Y 0.01fF
C30042 PAND2X1_469/B PAND2X1_556/O 0.17fF
C30043 PAND2X1_545/a_16_344# PAND2X1_324/Y 0.04fF
C30044 POR2X1_834/a_56_344# POR2X1_407/Y 0.00fF
C30045 POR2X1_403/B VDD 0.12fF
C30046 PAND2X1_192/Y PAND2X1_191/Y 0.05fF
C30047 POR2X1_567/B POR2X1_190/a_16_28# 0.02fF
C30048 PAND2X1_631/A PAND2X1_717/A 0.07fF
C30049 POR2X1_260/B POR2X1_553/A 0.03fF
C30050 PAND2X1_6/Y POR2X1_812/A 0.29fF
C30051 POR2X1_590/A POR2X1_68/B 0.23fF
C30052 D_INPUT_0 POR2X1_228/Y 0.10fF
C30053 POR2X1_52/A POR2X1_238/CTRL 0.08fF
C30054 PAND2X1_852/B POR2X1_102/Y 0.01fF
C30055 POR2X1_529/Y POR2X1_37/Y 0.20fF
C30056 POR2X1_489/a_16_28# POR2X1_489/A 0.03fF
C30057 PAND2X1_674/CTRL POR2X1_186/Y 0.03fF
C30058 POR2X1_278/Y VDD 2.97fF
C30059 POR2X1_716/a_16_28# POR2X1_303/B 0.07fF
C30060 POR2X1_145/Y POR2X1_669/B 0.02fF
C30061 PAND2X1_34/a_76_28# POR2X1_38/Y 0.02fF
C30062 PAND2X1_272/O PAND2X1_60/B 0.04fF
C30063 PAND2X1_23/Y PAND2X1_55/O 0.00fF
C30064 POR2X1_550/A D_INPUT_0 0.04fF
C30065 POR2X1_529/CTRL2 POR2X1_5/Y 0.02fF
C30066 POR2X1_41/B PAND2X1_804/A 0.06fF
C30067 PAND2X1_460/Y PAND2X1_459/Y 0.02fF
C30068 PAND2X1_23/Y POR2X1_805/B 0.14fF
C30069 POR2X1_786/Y POR2X1_330/Y 0.07fF
C30070 PAND2X1_90/A PAND2X1_263/O 0.00fF
C30071 PAND2X1_480/B PAND2X1_151/O 0.00fF
C30072 PAND2X1_245/CTRL PAND2X1_111/B 0.01fF
C30073 POR2X1_54/Y PAND2X1_522/a_56_28# 0.00fF
C30074 POR2X1_264/Y POR2X1_267/B 0.01fF
C30075 PAND2X1_57/B POR2X1_546/A 0.51fF
C30076 POR2X1_775/A PAND2X1_229/O 0.02fF
C30077 PAND2X1_139/O POR2X1_184/Y 0.00fF
C30078 PAND2X1_96/B POR2X1_288/a_16_28# 0.02fF
C30079 PAND2X1_593/O PAND2X1_364/B 0.09fF
C30080 PAND2X1_118/CTRL2 PAND2X1_65/B 0.01fF
C30081 POR2X1_422/O POR2X1_260/A 0.01fF
C30082 POR2X1_68/A POR2X1_849/CTRL2 0.00fF
C30083 POR2X1_68/A PAND2X1_55/CTRL 0.03fF
C30084 PAND2X1_433/O PAND2X1_65/B 0.03fF
C30085 PAND2X1_329/CTRL2 POR2X1_149/A 0.00fF
C30086 POR2X1_441/Y POR2X1_373/O 0.01fF
C30087 POR2X1_235/O POR2X1_32/A 0.01fF
C30088 POR2X1_201/CTRL PAND2X1_88/Y 0.01fF
C30089 PAND2X1_659/A POR2X1_816/A 0.01fF
C30090 POR2X1_481/a_16_28# POR2X1_295/Y 0.04fF
C30091 PAND2X1_598/CTRL POR2X1_46/Y 0.13fF
C30092 POR2X1_41/B PAND2X1_785/Y 0.03fF
C30093 POR2X1_23/Y PAND2X1_726/B 0.07fF
C30094 POR2X1_78/B POR2X1_659/CTRL2 0.03fF
C30095 POR2X1_72/CTRL POR2X1_816/A 0.01fF
C30096 POR2X1_65/A PAND2X1_365/B 0.01fF
C30097 PAND2X1_347/Y POR2X1_42/Y 0.03fF
C30098 PAND2X1_483/O POR2X1_48/A 0.03fF
C30099 PAND2X1_632/CTRL2 POR2X1_496/Y 0.06fF
C30100 POR2X1_516/a_16_28# POR2X1_423/Y 0.01fF
C30101 POR2X1_648/Y PAND2X1_56/A 0.03fF
C30102 POR2X1_66/A POR2X1_773/a_16_28# 0.03fF
C30103 POR2X1_383/A PAND2X1_279/CTRL 0.03fF
C30104 PAND2X1_3/CTRL2 PAND2X1_11/Y 0.01fF
C30105 POR2X1_671/O D_INPUT_2 0.01fF
C30106 D_INPUT_1 PAND2X1_526/O 0.01fF
C30107 POR2X1_130/a_16_28# POR2X1_141/A 0.04fF
C30108 POR2X1_299/Y PAND2X1_308/Y 0.01fF
C30109 POR2X1_49/Y POR2X1_583/CTRL 0.02fF
C30110 POR2X1_294/a_76_344# POR2X1_294/A 0.00fF
C30111 POR2X1_608/CTRL2 POR2X1_712/Y 0.03fF
C30112 POR2X1_10/CTRL2 POR2X1_669/B 0.01fF
C30113 POR2X1_193/Y POR2X1_219/O 0.07fF
C30114 POR2X1_96/A PAND2X1_188/CTRL 0.01fF
C30115 PAND2X1_637/CTRL2 PAND2X1_638/B 0.01fF
C30116 POR2X1_652/O PAND2X1_90/Y 0.12fF
C30117 PAND2X1_744/CTRL VDD 0.00fF
C30118 POR2X1_330/Y PAND2X1_163/CTRL 0.04fF
C30119 POR2X1_614/A POR2X1_480/A 0.07fF
C30120 POR2X1_542/B POR2X1_663/CTRL2 0.06fF
C30121 POR2X1_46/Y POR2X1_55/Y 0.09fF
C30122 PAND2X1_211/A POR2X1_91/Y 0.02fF
C30123 PAND2X1_93/B PAND2X1_394/CTRL2 0.00fF
C30124 PAND2X1_486/O POR2X1_763/Y 0.05fF
C30125 POR2X1_358/CTRL POR2X1_578/Y 0.03fF
C30126 POR2X1_66/A POR2X1_546/a_16_28# 0.01fF
C30127 PAND2X1_787/Y PAND2X1_390/m4_208_n4# 0.07fF
C30128 POR2X1_254/Y D_GATE_222 1.31fF
C30129 PAND2X1_205/Y PAND2X1_186/a_76_28# 0.01fF
C30130 POR2X1_486/B POR2X1_556/A 0.02fF
C30131 D_INPUT_5 PAND2X1_2/a_76_28# 0.01fF
C30132 POR2X1_210/CTRL POR2X1_210/B 0.05fF
C30133 PAND2X1_742/B POR2X1_331/A 0.02fF
C30134 PAND2X1_197/Y PAND2X1_364/B 0.03fF
C30135 PAND2X1_661/Y POR2X1_40/Y 0.03fF
C30136 PAND2X1_7/Y POR2X1_510/Y 0.09fF
C30137 PAND2X1_95/a_76_28# PAND2X1_57/B 0.03fF
C30138 POR2X1_65/A POR2X1_313/a_16_28# 0.01fF
C30139 PAND2X1_58/A POR2X1_675/Y 0.03fF
C30140 PAND2X1_20/A POR2X1_456/B 0.06fF
C30141 PAND2X1_623/CTRL2 POR2X1_129/Y 0.01fF
C30142 POR2X1_355/B POR2X1_68/A 0.03fF
C30143 POR2X1_57/A POR2X1_666/A 1.01fF
C30144 POR2X1_593/a_16_28# PAND2X1_93/B 0.03fF
C30145 INPUT_2 VDD 1.02fF
C30146 POR2X1_669/B POR2X1_394/A 1.21fF
C30147 POR2X1_753/Y POR2X1_753/O 0.06fF
C30148 POR2X1_708/CTRL PAND2X1_32/B 0.11fF
C30149 POR2X1_302/Y PAND2X1_69/A 0.02fF
C30150 PAND2X1_90/A POR2X1_572/B 0.03fF
C30151 POR2X1_131/CTRL2 PAND2X1_137/Y 0.05fF
C30152 PAND2X1_738/Y POR2X1_90/Y 0.05fF
C30153 POR2X1_761/Y VDD 0.20fF
C30154 POR2X1_94/O POR2X1_7/B 0.01fF
C30155 PAND2X1_398/O POR2X1_293/Y 0.17fF
C30156 POR2X1_416/Y POR2X1_290/Y 0.09fF
C30157 POR2X1_775/CTRL2 POR2X1_776/B 0.00fF
C30158 PAND2X1_649/A PAND2X1_590/CTRL2 0.01fF
C30159 PAND2X1_94/A PAND2X1_46/O 0.01fF
C30160 POR2X1_532/A POR2X1_794/O 0.01fF
C30161 POR2X1_780/a_56_344# POR2X1_796/A 0.00fF
C30162 POR2X1_270/Y POR2X1_540/Y 0.05fF
C30163 POR2X1_52/A POR2X1_237/Y 0.02fF
C30164 POR2X1_559/CTRL2 PAND2X1_90/A 0.01fF
C30165 VDD PAND2X1_156/O 0.00fF
C30166 POR2X1_48/A POR2X1_749/Y 0.06fF
C30167 POR2X1_433/O POR2X1_153/Y 0.05fF
C30168 POR2X1_83/B PAND2X1_358/A 0.07fF
C30169 PAND2X1_754/CTRL PAND2X1_69/A 0.12fF
C30170 POR2X1_326/A POR2X1_590/A 0.12fF
C30171 PAND2X1_787/Y POR2X1_283/A 0.10fF
C30172 PAND2X1_90/Y POR2X1_704/O 0.01fF
C30173 POR2X1_344/A POR2X1_532/A 0.11fF
C30174 POR2X1_197/a_16_28# POR2X1_196/Y 0.02fF
C30175 POR2X1_254/Y POR2X1_702/CTRL2 0.08fF
C30176 POR2X1_288/A POR2X1_734/CTRL2 0.00fF
C30177 PAND2X1_6/Y PAND2X1_48/B 3.09fF
C30178 PAND2X1_859/a_76_28# POR2X1_283/A 0.04fF
C30179 PAND2X1_676/O PAND2X1_480/B 0.01fF
C30180 PAND2X1_593/a_76_28# POR2X1_591/Y 0.02fF
C30181 POR2X1_691/O POR2X1_800/A 0.00fF
C30182 POR2X1_614/A PAND2X1_90/A 0.29fF
C30183 PAND2X1_476/A D_INPUT_0 0.03fF
C30184 POR2X1_96/A POR2X1_93/A 0.16fF
C30185 POR2X1_529/a_16_28# POR2X1_55/Y 0.06fF
C30186 POR2X1_814/B POR2X1_456/B 0.13fF
C30187 POR2X1_121/B POR2X1_737/A 0.02fF
C30188 POR2X1_244/B POR2X1_350/B 0.03fF
C30189 POR2X1_440/Y POR2X1_480/A 0.02fF
C30190 POR2X1_96/A POR2X1_91/Y 0.06fF
C30191 POR2X1_16/A PAND2X1_363/Y 0.03fF
C30192 POR2X1_196/a_16_28# POR2X1_334/Y 0.05fF
C30193 POR2X1_750/B POR2X1_733/Y 0.06fF
C30194 POR2X1_618/CTRL POR2X1_382/Y 0.01fF
C30195 POR2X1_119/Y PAND2X1_404/CTRL2 0.00fF
C30196 POR2X1_253/Y PAND2X1_658/B 0.02fF
C30197 PAND2X1_857/B VDD 0.01fF
C30198 POR2X1_271/A POR2X1_423/Y 0.03fF
C30199 PAND2X1_90/A POR2X1_38/B 0.94fF
C30200 PAND2X1_550/B PAND2X1_549/CTRL2 0.01fF
C30201 POR2X1_82/CTRL2 INPUT_1 0.01fF
C30202 POR2X1_775/A POR2X1_702/A 0.00fF
C30203 PAND2X1_90/Y POR2X1_721/CTRL 0.06fF
C30204 POR2X1_294/B PAND2X1_88/Y 0.03fF
C30205 POR2X1_76/Y POR2X1_222/A 0.03fF
C30206 POR2X1_669/B POR2X1_701/a_16_28# 0.05fF
C30207 PAND2X1_48/B POR2X1_791/A 0.01fF
C30208 POR2X1_220/CTRL PAND2X1_52/B 0.01fF
C30209 POR2X1_84/Y POR2X1_294/B 0.01fF
C30210 POR2X1_41/B PAND2X1_656/A 0.03fF
C30211 POR2X1_192/Y POR2X1_566/B 0.05fF
C30212 POR2X1_655/A POR2X1_725/O 0.12fF
C30213 POR2X1_333/A POR2X1_169/B 0.02fF
C30214 POR2X1_20/O POR2X1_380/Y 0.11fF
C30215 POR2X1_325/A POR2X1_456/B 0.01fF
C30216 PAND2X1_76/a_76_28# POR2X1_75/Y 0.04fF
C30217 POR2X1_281/Y POR2X1_282/Y 0.20fF
C30218 POR2X1_192/Y POR2X1_180/A 0.10fF
C30219 POR2X1_319/A PAND2X1_52/B 0.03fF
C30220 PAND2X1_824/B POR2X1_207/A 0.05fF
C30221 POR2X1_590/A POR2X1_362/a_76_344# 0.00fF
C30222 POR2X1_785/O POR2X1_566/B 0.18fF
C30223 PAND2X1_220/CTRL2 POR2X1_142/Y 0.10fF
C30224 POR2X1_97/A POR2X1_568/B 0.03fF
C30225 PAND2X1_691/Y PAND2X1_719/a_16_344# 0.01fF
C30226 POR2X1_743/O POR2X1_153/Y 0.10fF
C30227 POR2X1_82/CTRL2 POR2X1_153/Y 0.09fF
C30228 POR2X1_96/A PAND2X1_641/CTRL2 0.03fF
C30229 POR2X1_360/A POR2X1_101/O 0.02fF
C30230 PAND2X1_741/B POR2X1_7/a_16_28# 0.07fF
C30231 PAND2X1_433/CTRL POR2X1_832/A 0.01fF
C30232 POR2X1_771/CTRL PAND2X1_32/B 0.01fF
C30233 POR2X1_52/Y POR2X1_73/Y 0.03fF
C30234 POR2X1_228/O PAND2X1_52/Y 0.11fF
C30235 POR2X1_112/Y POR2X1_702/A 0.29fF
C30236 PAND2X1_228/O PAND2X1_656/A 0.02fF
C30237 POR2X1_258/Y PAND2X1_555/A 0.01fF
C30238 POR2X1_349/CTRL2 PAND2X1_65/Y 0.01fF
C30239 PAND2X1_69/A PAND2X1_150/CTRL2 0.00fF
C30240 POR2X1_287/B POR2X1_294/A 0.06fF
C30241 POR2X1_458/O POR2X1_717/B 0.00fF
C30242 POR2X1_567/A POR2X1_259/A 0.05fF
C30243 POR2X1_368/Y PAND2X1_787/A 0.02fF
C30244 PAND2X1_663/CTRL2 POR2X1_413/A 0.01fF
C30245 POR2X1_821/Y PAND2X1_852/B 0.10fF
C30246 POR2X1_116/Y POR2X1_392/a_56_344# 0.00fF
C30247 PAND2X1_793/Y PAND2X1_510/O 0.01fF
C30248 PAND2X1_469/B PAND2X1_175/B 0.05fF
C30249 POR2X1_750/B PAND2X1_526/CTRL2 0.07fF
C30250 PAND2X1_467/Y POR2X1_697/Y 0.03fF
C30251 POR2X1_748/A PAND2X1_508/B 0.03fF
C30252 D_INPUT_3 POR2X1_63/a_76_344# 0.02fF
C30253 POR2X1_502/A POR2X1_6/O 0.02fF
C30254 POR2X1_857/B POR2X1_502/O 0.01fF
C30255 POR2X1_103/CTRL POR2X1_13/A 0.01fF
C30256 POR2X1_49/Y PAND2X1_338/O 0.15fF
C30257 POR2X1_616/Y POR2X1_5/Y 0.05fF
C30258 POR2X1_306/a_76_344# POR2X1_90/Y 0.00fF
C30259 POR2X1_41/B PAND2X1_348/A 0.07fF
C30260 POR2X1_96/Y PAND2X1_61/Y 0.73fF
C30261 PAND2X1_738/Y PAND2X1_360/Y 0.05fF
C30262 POR2X1_858/B POR2X1_733/A 0.03fF
C30263 PAND2X1_241/Y POR2X1_73/Y 0.00fF
C30264 PAND2X1_605/CTRL POR2X1_42/Y 0.01fF
C30265 PAND2X1_691/Y PAND2X1_649/CTRL 0.17fF
C30266 POR2X1_318/A POR2X1_140/CTRL2 0.02fF
C30267 POR2X1_316/Y PAND2X1_390/Y 0.01fF
C30268 POR2X1_336/CTRL POR2X1_228/Y 0.01fF
C30269 POR2X1_419/a_56_344# POR2X1_42/Y 0.00fF
C30270 PAND2X1_69/A POR2X1_7/A 0.03fF
C30271 PAND2X1_243/O PAND2X1_338/B 0.08fF
C30272 POR2X1_486/O POR2X1_705/B 0.00fF
C30273 POR2X1_707/Y POR2X1_712/Y 0.01fF
C30274 POR2X1_96/A POR2X1_533/CTRL 0.01fF
C30275 PAND2X1_489/CTRL PAND2X1_794/B 0.01fF
C30276 POR2X1_56/B POR2X1_153/Y 2.25fF
C30277 PAND2X1_236/O POR2X1_4/Y 0.04fF
C30278 POR2X1_845/CTRL POR2X1_532/A 0.04fF
C30279 POR2X1_438/CTRL PAND2X1_569/B 0.03fF
C30280 POR2X1_96/A POR2X1_109/Y 0.03fF
C30281 POR2X1_93/A POR2X1_7/A 0.10fF
C30282 POR2X1_812/A PAND2X1_52/B 0.03fF
C30283 PAND2X1_341/B POR2X1_88/Y 0.05fF
C30284 POR2X1_7/A POR2X1_91/Y 0.03fF
C30285 POR2X1_62/Y PAND2X1_364/B 0.33fF
C30286 POR2X1_119/Y PAND2X1_862/B 0.05fF
C30287 POR2X1_98/A POR2X1_202/A 0.02fF
C30288 POR2X1_447/B POR2X1_220/Y 0.07fF
C30289 PAND2X1_69/A POR2X1_703/A 0.38fF
C30290 POR2X1_852/A POR2X1_192/B 0.02fF
C30291 PAND2X1_502/O POR2X1_42/Y 0.06fF
C30292 POR2X1_283/A POR2X1_248/Y 0.03fF
C30293 POR2X1_20/B POR2X1_411/A 0.07fF
C30294 POR2X1_9/Y POR2X1_818/Y 0.04fF
C30295 POR2X1_43/B PAND2X1_853/B 5.13fF
C30296 PAND2X1_96/B POR2X1_675/Y 0.83fF
C30297 POR2X1_41/B PAND2X1_631/A 0.10fF
C30298 POR2X1_736/CTRL2 POR2X1_675/Y 0.01fF
C30299 PAND2X1_226/a_16_344# POR2X1_192/B 0.02fF
C30300 PAND2X1_226/CTRL POR2X1_191/Y -0.01fF
C30301 PAND2X1_61/Y PAND2X1_333/Y 0.03fF
C30302 POR2X1_62/Y PAND2X1_101/O 0.02fF
C30303 PAND2X1_56/Y POR2X1_737/A 0.03fF
C30304 POR2X1_41/B PAND2X1_857/a_16_344# 0.01fF
C30305 POR2X1_786/Y POR2X1_715/A 0.01fF
C30306 POR2X1_637/A PAND2X1_72/A 0.04fF
C30307 PAND2X1_8/Y PAND2X1_102/CTRL 0.01fF
C30308 POR2X1_383/A POR2X1_561/CTRL2 0.03fF
C30309 PAND2X1_94/A POR2X1_713/B 0.10fF
C30310 PAND2X1_96/B POR2X1_544/B 0.03fF
C30311 POR2X1_216/a_16_28# POR2X1_116/Y -0.00fF
C30312 POR2X1_566/B POR2X1_568/Y 1.32fF
C30313 POR2X1_840/a_16_28# POR2X1_834/Y 0.03fF
C30314 POR2X1_52/A PAND2X1_326/B 0.03fF
C30315 POR2X1_483/B POR2X1_632/Y 0.01fF
C30316 PAND2X1_569/a_76_28# POR2X1_73/Y 0.01fF
C30317 POR2X1_355/B POR2X1_169/A 0.03fF
C30318 POR2X1_853/A PAND2X1_165/O 0.01fF
C30319 POR2X1_785/B POR2X1_566/B 0.29fF
C30320 POR2X1_775/CTRL2 POR2X1_192/B 0.12fF
C30321 POR2X1_416/B INPUT_0 0.06fF
C30322 PAND2X1_40/a_16_344# PAND2X1_3/B 0.01fF
C30323 PAND2X1_785/Y POR2X1_77/Y 0.00fF
C30324 POR2X1_152/A PAND2X1_326/B 0.03fF
C30325 POR2X1_305/CTRL2 POR2X1_7/B 0.00fF
C30326 POR2X1_169/CTRL POR2X1_568/Y 0.22fF
C30327 POR2X1_93/A POR2X1_384/Y 0.01fF
C30328 POR2X1_16/A POR2X1_73/O 0.01fF
C30329 POR2X1_366/Y POR2X1_568/B 0.10fF
C30330 POR2X1_294/B POR2X1_568/B 0.08fF
C30331 POR2X1_804/A POR2X1_188/Y 0.03fF
C30332 POR2X1_245/O PAND2X1_156/A 0.16fF
C30333 POR2X1_123/A POR2X1_559/A 0.05fF
C30334 POR2X1_27/CTRL POR2X1_32/A 0.01fF
C30335 PAND2X1_48/B POR2X1_632/Y 0.04fF
C30336 POR2X1_566/CTRL2 POR2X1_854/B 0.01fF
C30337 PAND2X1_246/O POR2X1_66/A 0.07fF
C30338 PAND2X1_631/A POR2X1_256/Y 0.02fF
C30339 POR2X1_463/Y POR2X1_260/A 0.03fF
C30340 PAND2X1_437/O POR2X1_186/Y 0.03fF
C30341 PAND2X1_319/B PAND2X1_352/CTRL2 0.02fF
C30342 PAND2X1_69/A POR2X1_342/a_16_28# 0.02fF
C30343 POR2X1_567/A PAND2X1_88/Y 0.05fF
C30344 POR2X1_447/B PAND2X1_824/CTRL2 0.00fF
C30345 PAND2X1_109/O D_GATE_222 0.06fF
C30346 POR2X1_754/Y POR2X1_846/Y 0.08fF
C30347 POR2X1_57/A PAND2X1_737/O 0.02fF
C30348 PAND2X1_779/CTRL2 PAND2X1_550/B 0.01fF
C30349 POR2X1_383/A POR2X1_737/A 0.03fF
C30350 POR2X1_846/A POR2X1_750/B 0.12fF
C30351 POR2X1_814/Y PAND2X1_58/A 0.36fF
C30352 POR2X1_745/Y POR2X1_746/a_16_28# 0.02fF
C30353 PAND2X1_467/Y PAND2X1_451/O 0.01fF
C30354 POR2X1_446/A POR2X1_446/a_16_28# 0.03fF
C30355 PAND2X1_23/Y POR2X1_509/CTRL 0.03fF
C30356 POR2X1_52/A POR2X1_387/a_16_28# 0.03fF
C30357 PAND2X1_48/B PAND2X1_52/B 0.20fF
C30358 POR2X1_318/A PAND2X1_136/CTRL2 0.03fF
C30359 POR2X1_456/B POR2X1_703/CTRL2 0.01fF
C30360 POR2X1_748/A POR2X1_329/A 0.10fF
C30361 PAND2X1_349/A PAND2X1_141/O 0.02fF
C30362 POR2X1_71/CTRL2 POR2X1_394/A 0.03fF
C30363 PAND2X1_849/B POR2X1_62/Y 0.73fF
C30364 POR2X1_411/B POR2X1_268/O 0.01fF
C30365 D_INPUT_3 PAND2X1_610/O 0.04fF
C30366 POR2X1_20/B POR2X1_32/A 0.68fF
C30367 POR2X1_407/Y D_INPUT_4 0.00fF
C30368 POR2X1_16/A PAND2X1_345/Y 0.03fF
C30369 PAND2X1_480/B PAND2X1_860/A 0.05fF
C30370 POR2X1_326/A POR2X1_737/m4_208_n4# 0.08fF
C30371 POR2X1_597/CTRL POR2X1_761/A 0.01fF
C30372 PAND2X1_23/Y PAND2X1_135/O 0.04fF
C30373 POR2X1_83/B POR2X1_441/Y 0.03fF
C30374 POR2X1_863/A POR2X1_149/Y 0.03fF
C30375 POR2X1_41/B PAND2X1_193/Y 1.82fF
C30376 POR2X1_48/A POR2X1_817/CTRL2 0.04fF
C30377 POR2X1_836/A POR2X1_776/A 0.03fF
C30378 POR2X1_669/B POR2X1_604/a_16_28# 0.05fF
C30379 PAND2X1_63/Y POR2X1_500/O 0.33fF
C30380 POR2X1_147/CTRL2 POR2X1_532/A 0.01fF
C30381 POR2X1_257/A PAND2X1_161/CTRL2 0.00fF
C30382 POR2X1_709/A POR2X1_14/Y 0.09fF
C30383 PAND2X1_295/CTRL POR2X1_296/B 0.00fF
C30384 POR2X1_657/CTRL POR2X1_446/B 0.01fF
C30385 POR2X1_417/Y POR2X1_20/B 5.16fF
C30386 POR2X1_87/a_16_28# POR2X1_68/B 0.11fF
C30387 PAND2X1_480/O POR2X1_119/Y 0.17fF
C30388 POR2X1_644/a_16_28# D_INPUT_0 0.02fF
C30389 POR2X1_329/A PAND2X1_596/a_16_344# 0.02fF
C30390 PAND2X1_628/CTRL POR2X1_785/A 0.00fF
C30391 PAND2X1_269/CTRL VDD -0.00fF
C30392 POR2X1_77/Y PAND2X1_656/A 0.03fF
C30393 POR2X1_48/A POR2X1_626/O 0.02fF
C30394 POR2X1_606/O POR2X1_590/A 0.00fF
C30395 POR2X1_606/CTRL POR2X1_121/B 0.01fF
C30396 POR2X1_406/Y PAND2X1_266/CTRL2 0.01fF
C30397 POR2X1_686/A POR2X1_864/A 0.00fF
C30398 POR2X1_63/Y POR2X1_72/B 0.06fF
C30399 POR2X1_590/A POR2X1_458/CTRL2 0.09fF
C30400 POR2X1_670/CTRL2 POR2X1_20/B 0.01fF
C30401 PAND2X1_640/B POR2X1_609/Y 0.03fF
C30402 POR2X1_311/CTRL POR2X1_77/Y 0.00fF
C30403 POR2X1_652/A POR2X1_802/A 0.56fF
C30404 PAND2X1_449/CTRL2 POR2X1_511/Y 0.09fF
C30405 PAND2X1_649/A POR2X1_394/A 0.00fF
C30406 POR2X1_49/Y PAND2X1_446/Y 0.00fF
C30407 POR2X1_18/CTRL INPUT_4 0.01fF
C30408 POR2X1_119/Y PAND2X1_716/B 0.13fF
C30409 PAND2X1_474/a_16_344# PAND2X1_474/A 0.01fF
C30410 PAND2X1_507/CTRL2 POR2X1_39/B 0.02fF
C30411 POR2X1_601/Y POR2X1_600/Y 1.46fF
C30412 PAND2X1_39/B POR2X1_398/Y 0.04fF
C30413 PAND2X1_319/O POR2X1_20/B 0.17fF
C30414 PAND2X1_747/m4_208_n4# PAND2X1_52/B 0.12fF
C30415 PAND2X1_865/Y POR2X1_767/CTRL 0.01fF
C30416 POR2X1_49/Y PAND2X1_444/CTRL2 0.01fF
C30417 D_INPUT_3 POR2X1_49/a_16_28# 0.03fF
C30418 POR2X1_119/Y POR2X1_518/CTRL2 0.08fF
C30419 PAND2X1_861/B PAND2X1_861/O 0.00fF
C30420 POR2X1_43/B POR2X1_827/CTRL 0.01fF
C30421 PAND2X1_20/A POR2X1_849/A 0.05fF
C30422 PAND2X1_348/A POR2X1_77/Y 0.05fF
C30423 PAND2X1_73/Y POR2X1_296/B 0.06fF
C30424 POR2X1_101/Y POR2X1_343/B 0.03fF
C30425 PAND2X1_493/O POR2X1_491/Y -0.00fF
C30426 POR2X1_416/B PAND2X1_343/a_16_344# 0.01fF
C30427 POR2X1_276/B VDD 0.00fF
C30428 PAND2X1_52/B POR2X1_210/B 0.02fF
C30429 POR2X1_666/O POR2X1_102/Y 0.01fF
C30430 PAND2X1_59/B PAND2X1_41/B 0.04fF
C30431 PAND2X1_410/CTRL2 POR2X1_236/Y 0.01fF
C30432 POR2X1_276/A POR2X1_76/B 0.01fF
C30433 PAND2X1_87/CTRL PAND2X1_6/A 0.07fF
C30434 POR2X1_846/Y POR2X1_790/a_76_344# 0.00fF
C30435 POR2X1_23/Y PAND2X1_208/O 0.03fF
C30436 POR2X1_20/B PAND2X1_35/Y 0.03fF
C30437 POR2X1_37/Y POR2X1_268/Y 0.00fF
C30438 POR2X1_78/A POR2X1_605/CTRL 0.05fF
C30439 POR2X1_117/CTRL2 POR2X1_48/A 0.01fF
C30440 POR2X1_383/O POR2X1_383/Y 0.01fF
C30441 POR2X1_728/O POR2X1_452/Y 0.01fF
C30442 POR2X1_491/CTRL2 POR2X1_32/A 0.03fF
C30443 POR2X1_36/B PAND2X1_635/Y 0.02fF
C30444 PAND2X1_73/Y PAND2X1_74/CTRL 0.01fF
C30445 POR2X1_14/Y PAND2X1_58/A 0.03fF
C30446 PAND2X1_39/B PAND2X1_57/B 0.50fF
C30447 POR2X1_427/O POR2X1_72/B 0.01fF
C30448 POR2X1_66/B POR2X1_240/B 0.01fF
C30449 POR2X1_567/A POR2X1_568/B 0.02fF
C30450 PAND2X1_61/Y POR2X1_37/Y 0.03fF
C30451 PAND2X1_73/O POR2X1_590/A 0.05fF
C30452 PAND2X1_403/B POR2X1_102/Y 0.07fF
C30453 POR2X1_808/A POR2X1_602/A 0.02fF
C30454 POR2X1_862/B POR2X1_646/Y 0.02fF
C30455 POR2X1_102/Y POR2X1_272/CTRL 0.01fF
C30456 PAND2X1_652/A POR2X1_150/Y 0.74fF
C30457 PAND2X1_631/A POR2X1_77/Y 0.03fF
C30458 PAND2X1_655/B POR2X1_600/CTRL 0.00fF
C30459 POR2X1_24/a_16_28# POR2X1_29/A 0.02fF
C30460 POR2X1_502/A POR2X1_602/O 0.02fF
C30461 PAND2X1_402/O POR2X1_14/Y 0.03fF
C30462 POR2X1_257/A PAND2X1_254/a_16_344# 0.02fF
C30463 POR2X1_20/B POR2X1_184/Y 0.03fF
C30464 POR2X1_112/CTRL2 PAND2X1_72/A 0.00fF
C30465 PAND2X1_621/CTRL2 POR2X1_9/Y 0.03fF
C30466 PAND2X1_406/CTRL POR2X1_784/A 0.02fF
C30467 POR2X1_662/CTRL PAND2X1_55/Y 0.01fF
C30468 PAND2X1_58/A PAND2X1_55/CTRL 0.01fF
C30469 PAND2X1_571/O PAND2X1_571/Y 0.19fF
C30470 POR2X1_634/CTRL PAND2X1_41/B 0.00fF
C30471 PAND2X1_58/A POR2X1_791/Y 0.01fF
C30472 POR2X1_52/A PAND2X1_852/A 0.05fF
C30473 PAND2X1_20/A PAND2X1_20/O 0.02fF
C30474 POR2X1_43/B PAND2X1_796/B 0.02fF
C30475 POR2X1_48/A POR2X1_411/CTRL2 0.03fF
C30476 PAND2X1_651/Y POR2X1_20/B 0.08fF
C30477 POR2X1_490/Y PAND2X1_215/B 0.01fF
C30478 POR2X1_480/A POR2X1_590/A 0.32fF
C30479 PAND2X1_58/A POR2X1_637/B 0.01fF
C30480 POR2X1_541/B POR2X1_702/A 0.03fF
C30481 POR2X1_440/O POR2X1_353/A 0.11fF
C30482 POR2X1_43/B PAND2X1_454/B 0.03fF
C30483 POR2X1_23/Y POR2X1_252/CTRL 0.04fF
C30484 POR2X1_48/A POR2X1_252/CTRL2 0.01fF
C30485 PAND2X1_570/O PAND2X1_562/Y 0.02fF
C30486 POR2X1_590/A POR2X1_207/CTRL2 0.00fF
C30487 PAND2X1_73/Y POR2X1_547/B 0.14fF
C30488 POR2X1_43/CTRL POR2X1_77/Y 0.00fF
C30489 POR2X1_347/A POR2X1_98/A 0.00fF
C30490 POR2X1_12/A PAND2X1_635/CTRL2 0.01fF
C30491 PAND2X1_39/B POR2X1_828/A 0.05fF
C30492 POR2X1_9/Y POR2X1_751/Y 0.03fF
C30493 PAND2X1_93/B POR2X1_198/B 2.24fF
C30494 POR2X1_20/B PAND2X1_844/B 0.02fF
C30495 POR2X1_679/A POR2X1_816/A 0.03fF
C30496 POR2X1_67/Y POR2X1_750/Y 0.05fF
C30497 POR2X1_416/B POR2X1_747/CTRL2 0.00fF
C30498 PAND2X1_60/a_76_28# POR2X1_35/Y 0.01fF
C30499 PAND2X1_564/B PAND2X1_564/CTRL 0.01fF
C30500 POR2X1_72/B PAND2X1_736/CTRL 0.01fF
C30501 POR2X1_814/A PAND2X1_503/O 0.09fF
C30502 PAND2X1_57/B POR2X1_805/Y 0.03fF
C30503 PAND2X1_60/O PAND2X1_69/A 0.06fF
C30504 POR2X1_260/B PAND2X1_316/O 0.02fF
C30505 POR2X1_124/CTRL POR2X1_78/A 0.01fF
C30506 PAND2X1_352/A POR2X1_55/Y 0.01fF
C30507 POR2X1_853/A POR2X1_856/B 0.03fF
C30508 PAND2X1_65/B PAND2X1_386/CTRL2 0.01fF
C30509 POR2X1_150/Y POR2X1_437/CTRL2 0.01fF
C30510 PAND2X1_96/B POR2X1_659/A 0.03fF
C30511 POR2X1_43/B POR2X1_23/Y 0.19fF
C30512 PAND2X1_6/Y POR2X1_796/Y 0.01fF
C30513 PAND2X1_556/B PAND2X1_444/Y 0.01fF
C30514 PAND2X1_20/A PAND2X1_57/B 0.38fF
C30515 POR2X1_119/Y PAND2X1_403/CTRL 0.01fF
C30516 POR2X1_536/Y VDD 0.00fF
C30517 POR2X1_341/A PAND2X1_111/B 0.08fF
C30518 POR2X1_257/A POR2X1_172/Y 0.03fF
C30519 POR2X1_860/A POR2X1_362/B 0.29fF
C30520 PAND2X1_169/Y VDD 0.00fF
C30521 PAND2X1_222/A POR2X1_591/Y 0.03fF
C30522 POR2X1_186/Y POR2X1_798/a_16_28# 0.09fF
C30523 POR2X1_855/a_16_28# POR2X1_803/A 0.01fF
C30524 POR2X1_846/Y POR2X1_754/CTRL 0.01fF
C30525 POR2X1_60/A PAND2X1_205/B 0.11fF
C30526 PAND2X1_90/A POR2X1_590/A 5.55fF
C30527 POR2X1_94/A PAND2X1_8/Y 2.98fF
C30528 PAND2X1_404/Y POR2X1_521/a_16_28# 0.00fF
C30529 PAND2X1_674/CTRL2 POR2X1_590/A 0.03fF
C30530 POR2X1_502/A POR2X1_794/B 0.72fF
C30531 POR2X1_150/Y PAND2X1_175/O 0.04fF
C30532 POR2X1_814/B POR2X1_608/CTRL2 0.01fF
C30533 POR2X1_72/B PAND2X1_558/a_76_28# 0.01fF
C30534 POR2X1_814/B PAND2X1_54/O 0.08fF
C30535 POR2X1_296/B PAND2X1_144/CTRL 0.08fF
C30536 PAND2X1_863/a_76_28# PAND2X1_805/A 0.01fF
C30537 PAND2X1_404/O POR2X1_293/Y 0.17fF
C30538 POR2X1_558/CTRL POR2X1_78/A 0.04fF
C30539 POR2X1_558/O PAND2X1_73/Y 0.28fF
C30540 PAND2X1_58/A POR2X1_55/Y 0.08fF
C30541 POR2X1_194/B POR2X1_194/A 0.05fF
C30542 POR2X1_406/Y PAND2X1_61/Y 0.81fF
C30543 POR2X1_624/Y PAND2X1_63/B 0.03fF
C30544 POR2X1_23/Y POR2X1_38/B 0.04fF
C30545 POR2X1_223/CTRL POR2X1_186/Y 0.01fF
C30546 POR2X1_218/Y POR2X1_513/Y 0.07fF
C30547 POR2X1_66/B POR2X1_124/a_56_344# 0.00fF
C30548 POR2X1_421/Y POR2X1_42/Y 0.03fF
C30549 PAND2X1_56/Y POR2X1_657/CTRL 0.14fF
C30550 PAND2X1_20/A POR2X1_285/A 0.01fF
C30551 PAND2X1_572/CTRL2 PAND2X1_576/B 0.01fF
C30552 PAND2X1_84/CTRL2 POR2X1_497/Y 0.01fF
C30553 PAND2X1_287/a_76_28# PAND2X1_577/Y 0.01fF
C30554 PAND2X1_673/O POR2X1_236/Y 0.01fF
C30555 POR2X1_820/Y POR2X1_376/B 0.07fF
C30556 POR2X1_814/A POR2X1_383/CTRL2 0.03fF
C30557 POR2X1_420/a_76_344# POR2X1_90/Y 0.00fF
C30558 POR2X1_689/A POR2X1_591/A 0.01fF
C30559 POR2X1_814/B PAND2X1_57/B 0.27fF
C30560 POR2X1_66/A POR2X1_68/B 0.42fF
C30561 PAND2X1_652/A PAND2X1_794/O 0.15fF
C30562 PAND2X1_340/O POR2X1_88/Y 0.15fF
C30563 POR2X1_161/m4_208_n4# POR2X1_568/m4_208_n4# 0.04fF
C30564 PAND2X1_853/O POR2X1_83/B 0.04fF
C30565 PAND2X1_93/B PAND2X1_312/a_16_344# 0.01fF
C30566 POR2X1_407/A POR2X1_656/a_16_28# 0.02fF
C30567 PAND2X1_480/B PAND2X1_579/m4_208_n4# 0.04fF
C30568 POR2X1_478/O POR2X1_568/Y 0.37fF
C30569 POR2X1_164/CTRL POR2X1_83/B 0.01fF
C30570 POR2X1_133/CTRL POR2X1_236/Y 0.00fF
C30571 PAND2X1_695/CTRL PAND2X1_57/B 0.01fF
C30572 PAND2X1_105/O POR2X1_60/A 0.05fF
C30573 PAND2X1_592/CTRL2 PAND2X1_473/B 0.03fF
C30574 PAND2X1_612/B POR2X1_773/CTRL 0.00fF
C30575 POR2X1_859/O POR2X1_559/A 0.28fF
C30576 PAND2X1_61/Y POR2X1_293/Y 0.03fF
C30577 PAND2X1_205/Y PAND2X1_215/B 0.04fF
C30578 PAND2X1_730/B VDD 2.59fF
C30579 POR2X1_403/A POR2X1_403/B 0.00fF
C30580 POR2X1_707/B PAND2X1_587/CTRL 0.01fF
C30581 INPUT_0 PAND2X1_512/Y 0.07fF
C30582 PAND2X1_650/O POR2X1_409/B 0.02fF
C30583 POR2X1_748/A PAND2X1_506/a_16_344# 0.02fF
C30584 POR2X1_124/B POR2X1_650/a_56_344# 0.00fF
C30585 PAND2X1_57/B POR2X1_325/A 0.03fF
C30586 PAND2X1_65/B POR2X1_776/B 0.07fF
C30587 PAND2X1_56/Y POR2X1_302/B 0.03fF
C30588 PAND2X1_852/O POR2X1_40/Y 0.15fF
C30589 POR2X1_65/A POR2X1_591/CTRL2 0.03fF
C30590 PAND2X1_850/Y PAND2X1_717/A 0.07fF
C30591 POR2X1_52/A PAND2X1_859/a_56_28# 0.00fF
C30592 POR2X1_830/m4_208_n4# POR2X1_741/Y 0.09fF
C30593 POR2X1_106/Y PAND2X1_115/B 0.02fF
C30594 POR2X1_218/Y POR2X1_366/A 0.07fF
C30595 POR2X1_567/B POR2X1_351/O 0.04fF
C30596 POR2X1_41/B PAND2X1_715/CTRL2 0.05fF
C30597 PAND2X1_58/A POR2X1_791/B 0.00fF
C30598 D_GATE_222 PAND2X1_41/B 0.10fF
C30599 POR2X1_66/B POR2X1_702/A 0.03fF
C30600 POR2X1_416/B POR2X1_292/CTRL2 0.03fF
C30601 PAND2X1_778/O POR2X1_293/Y 0.11fF
C30602 POR2X1_260/B POR2X1_576/a_56_344# 0.00fF
C30603 POR2X1_625/a_16_28# POR2X1_293/Y 0.00fF
C30604 PAND2X1_206/A PAND2X1_358/A 0.03fF
C30605 PAND2X1_607/a_16_344# PAND2X1_56/A 0.01fF
C30606 POR2X1_77/O POR2X1_394/A 0.04fF
C30607 PAND2X1_404/A POR2X1_293/Y 0.10fF
C30608 POR2X1_264/O PAND2X1_32/B 0.01fF
C30609 POR2X1_121/B PAND2X1_305/CTRL2 0.10fF
C30610 POR2X1_556/A POR2X1_362/CTRL 0.01fF
C30611 POR2X1_270/Y POR2X1_260/A 0.03fF
C30612 POR2X1_72/B POR2X1_498/A 0.16fF
C30613 POR2X1_330/Y PAND2X1_311/CTRL 0.13fF
C30614 PAND2X1_250/CTRL PAND2X1_69/A 0.05fF
C30615 POR2X1_312/a_56_344# POR2X1_65/A 0.00fF
C30616 PAND2X1_57/B POR2X1_513/B 0.37fF
C30617 POR2X1_12/A POR2X1_3/B 0.03fF
C30618 POR2X1_57/A POR2X1_748/A 1.57fF
C30619 POR2X1_335/CTRL2 POR2X1_741/Y 0.01fF
C30620 PAND2X1_674/m4_208_n4# POR2X1_675/m4_208_n4# 0.13fF
C30621 PAND2X1_697/CTRL2 PAND2X1_90/Y 0.03fF
C30622 POR2X1_729/m4_208_n4# POR2X1_864/m4_208_n4# 0.13fF
C30623 PAND2X1_462/B VDD 0.02fF
C30624 PAND2X1_48/CTRL POR2X1_294/B 0.01fF
C30625 POR2X1_283/A POR2X1_226/CTRL 0.03fF
C30626 POR2X1_496/Y PAND2X1_508/CTRL2 0.04fF
C30627 POR2X1_330/Y POR2X1_541/a_76_344# 0.01fF
C30628 POR2X1_118/Y POR2X1_153/Y 0.07fF
C30629 PAND2X1_622/CTRL2 POR2X1_619/Y 0.01fF
C30630 PAND2X1_342/CTRL2 POR2X1_5/Y 0.04fF
C30631 POR2X1_468/B POR2X1_802/B 0.22fF
C30632 PAND2X1_96/B POR2X1_791/Y 0.02fF
C30633 POR2X1_341/A PAND2X1_323/O 0.08fF
C30634 PAND2X1_65/B POR2X1_577/CTRL2 0.03fF
C30635 PAND2X1_56/Y POR2X1_335/O 0.02fF
C30636 POR2X1_467/Y PAND2X1_534/O 0.02fF
C30637 POR2X1_537/Y POR2X1_655/A 0.02fF
C30638 PAND2X1_478/Y POR2X1_91/Y 0.05fF
C30639 POR2X1_188/A POR2X1_121/O 0.01fF
C30640 PAND2X1_90/Y POR2X1_758/CTRL2 0.15fF
C30641 PAND2X1_653/m4_208_n4# PAND2X1_652/A 0.05fF
C30642 POR2X1_48/A POR2X1_183/CTRL2 0.01fF
C30643 POR2X1_383/A POR2X1_302/B 0.14fF
C30644 PAND2X1_784/O POR2X1_293/Y 0.09fF
C30645 POR2X1_855/B POR2X1_750/B 0.05fF
C30646 POR2X1_119/Y POR2X1_490/Y 0.05fF
C30647 D_INPUT_0 POR2X1_579/B 0.01fF
C30648 POR2X1_806/CTRL2 POR2X1_675/Y 0.01fF
C30649 POR2X1_32/A PAND2X1_303/Y 0.03fF
C30650 POR2X1_502/A POR2X1_638/B 0.01fF
C30651 POR2X1_26/O POR2X1_83/B 0.01fF
C30652 POR2X1_206/A PAND2X1_69/A 0.02fF
C30653 POR2X1_439/Y PAND2X1_60/B 0.03fF
C30654 POR2X1_335/A PAND2X1_498/CTRL2 0.01fF
C30655 POR2X1_186/Y POR2X1_854/B 0.03fF
C30656 PAND2X1_48/B PAND2X1_95/B 0.38fF
C30657 POR2X1_322/Y POR2X1_376/B 0.01fF
C30658 POR2X1_857/B POR2X1_350/CTRL 0.03fF
C30659 POR2X1_723/a_16_28# POR2X1_723/B 0.05fF
C30660 POR2X1_65/A POR2X1_73/CTRL2 -0.00fF
C30661 POR2X1_41/B POR2X1_183/Y 0.94fF
C30662 PAND2X1_298/CTRL2 POR2X1_750/B 0.03fF
C30663 PAND2X1_93/O POR2X1_404/Y 0.05fF
C30664 POR2X1_52/A PAND2X1_794/B 0.03fF
C30665 POR2X1_208/A PAND2X1_65/Y 0.00fF
C30666 POR2X1_174/B POR2X1_333/Y 0.03fF
C30667 INPUT_1 POR2X1_159/O 0.00fF
C30668 PAND2X1_55/Y POR2X1_659/CTRL 0.00fF
C30669 POR2X1_356/A POR2X1_340/a_16_28# 0.12fF
C30670 PAND2X1_293/O POR2X1_68/B 0.08fF
C30671 POR2X1_56/B PAND2X1_449/Y 0.02fF
C30672 PAND2X1_94/A POR2X1_35/B 0.06fF
C30673 D_INPUT_0 POR2X1_571/Y 0.01fF
C30674 PAND2X1_573/B POR2X1_153/Y 0.03fF
C30675 POR2X1_66/B POR2X1_768/O 0.10fF
C30676 POR2X1_284/CTRL2 POR2X1_804/A 0.03fF
C30677 POR2X1_355/B PAND2X1_96/B 0.03fF
C30678 POR2X1_488/Y PAND2X1_357/Y 0.00fF
C30679 PAND2X1_753/O PAND2X1_752/Y 0.00fF
C30680 POR2X1_49/Y PAND2X1_620/CTRL2 0.01fF
C30681 POR2X1_66/A PAND2X1_143/O 0.04fF
C30682 POR2X1_41/B PAND2X1_243/O 0.00fF
C30683 PAND2X1_3/a_76_28# POR2X1_750/B 0.01fF
C30684 POR2X1_57/A POR2X1_79/Y 0.03fF
C30685 POR2X1_732/O POR2X1_732/B 0.01fF
C30686 POR2X1_72/Y POR2X1_73/Y 0.03fF
C30687 PAND2X1_35/B POR2X1_394/A 0.12fF
C30688 POR2X1_192/Y PAND2X1_60/B 0.15fF
C30689 PAND2X1_498/O POR2X1_840/B 0.05fF
C30690 POR2X1_651/O POR2X1_639/Y 0.03fF
C30691 PAND2X1_91/a_76_28# POR2X1_169/A 0.02fF
C30692 POR2X1_96/A PAND2X1_338/B 0.03fF
C30693 POR2X1_130/Y POR2X1_140/A 0.01fF
C30694 POR2X1_439/Y POR2X1_353/A 0.49fF
C30695 POR2X1_186/a_76_344# POR2X1_750/B 0.01fF
C30696 PAND2X1_691/Y POR2X1_236/Y 0.07fF
C30697 POR2X1_198/CTRL2 POR2X1_532/A 0.03fF
C30698 POR2X1_115/CTRL POR2X1_366/A 0.08fF
C30699 POR2X1_41/Y POR2X1_669/B 0.02fF
C30700 PAND2X1_320/m4_208_n4# POR2X1_568/Y 0.06fF
C30701 D_INPUT_5 PAND2X1_52/B 0.05fF
C30702 POR2X1_766/O VDD 0.00fF
C30703 POR2X1_322/Y POR2X1_52/A 0.03fF
C30704 POR2X1_402/A PAND2X1_69/CTRL2 0.01fF
C30705 POR2X1_68/A POR2X1_513/Y 0.03fF
C30706 POR2X1_853/A POR2X1_577/CTRL 0.01fF
C30707 POR2X1_447/B PAND2X1_626/CTRL 0.04fF
C30708 POR2X1_387/Y POR2X1_372/Y 0.05fF
C30709 POR2X1_346/O PAND2X1_55/Y 0.01fF
C30710 POR2X1_305/Y POR2X1_90/Y 0.15fF
C30711 POR2X1_68/A POR2X1_219/B 0.05fF
C30712 POR2X1_388/CTRL2 PAND2X1_69/A 0.01fF
C30713 INPUT_1 PAND2X1_54/a_16_344# 0.02fF
C30714 PAND2X1_46/a_16_344# PAND2X1_71/Y 0.01fF
C30715 POR2X1_456/B VDD 0.46fF
C30716 POR2X1_16/A VDD 4.49fF
C30717 POR2X1_777/B PAND2X1_48/A 0.43fF
C30718 POR2X1_130/A POR2X1_773/B 0.02fF
C30719 PAND2X1_738/Y PAND2X1_181/m4_208_n4# 0.04fF
C30720 POR2X1_322/Y POR2X1_152/A 0.03fF
C30721 POR2X1_341/A POR2X1_579/a_76_344# -0.02fF
C30722 POR2X1_794/B POR2X1_188/Y 0.02fF
C30723 POR2X1_796/Y PAND2X1_52/B 1.11fF
C30724 PAND2X1_216/B PAND2X1_473/Y 0.03fF
C30725 POR2X1_425/O POR2X1_158/B 0.01fF
C30726 POR2X1_356/A POR2X1_738/A 0.05fF
C30727 PAND2X1_824/B POR2X1_206/A 0.09fF
C30728 POR2X1_407/A POR2X1_865/B 0.03fF
C30729 POR2X1_566/A POR2X1_97/O 0.29fF
C30730 POR2X1_68/A POR2X1_205/A 0.10fF
C30731 PAND2X1_462/O POR2X1_37/Y 0.09fF
C30732 POR2X1_179/CTRL POR2X1_387/Y 0.02fF
C30733 POR2X1_55/Y POR2X1_103/Y 0.01fF
C30734 POR2X1_834/Y POR2X1_722/Y 0.03fF
C30735 D_GATE_222 POR2X1_228/Y 0.72fF
C30736 PAND2X1_251/CTRL POR2X1_717/B 0.01fF
C30737 POR2X1_192/Y POR2X1_353/A 0.15fF
C30738 PAND2X1_72/O POR2X1_532/A 0.05fF
C30739 PAND2X1_639/B POR2X1_588/Y 0.03fF
C30740 PAND2X1_674/a_16_344# PAND2X1_60/B 0.01fF
C30741 POR2X1_632/B POR2X1_632/Y 0.17fF
C30742 PAND2X1_65/B PAND2X1_48/A 0.17fF
C30743 PAND2X1_23/Y PAND2X1_373/O 0.02fF
C30744 PAND2X1_274/CTRL POR2X1_153/Y 0.01fF
C30745 PAND2X1_341/A POR2X1_38/Y 0.03fF
C30746 POR2X1_68/A POR2X1_366/A 0.04fF
C30747 POR2X1_707/CTRL2 PAND2X1_95/B 0.01fF
C30748 PAND2X1_65/B POR2X1_192/B 0.05fF
C30749 POR2X1_532/A POR2X1_68/B 0.11fF
C30750 PAND2X1_659/Y PAND2X1_204/CTRL 0.01fF
C30751 POR2X1_848/A POR2X1_90/CTRL 0.08fF
C30752 PAND2X1_476/A PAND2X1_231/O 0.00fF
C30753 PAND2X1_493/CTRL2 PAND2X1_480/B 0.03fF
C30754 POR2X1_470/CTRL PAND2X1_52/B 0.03fF
C30755 PAND2X1_173/O PAND2X1_32/B 0.06fF
C30756 POR2X1_52/Y PAND2X1_656/A 0.02fF
C30757 POR2X1_364/A POR2X1_578/a_16_28# 0.01fF
C30758 POR2X1_730/Y POR2X1_832/B 0.01fF
C30759 POR2X1_57/A POR2X1_291/Y 0.04fF
C30760 POR2X1_416/B POR2X1_102/Y 0.52fF
C30761 POR2X1_628/O POR2X1_260/A 0.01fF
C30762 POR2X1_46/Y POR2X1_129/Y 0.05fF
C30763 POR2X1_741/Y POR2X1_456/B 0.06fF
C30764 POR2X1_334/Y PAND2X1_89/CTRL 0.07fF
C30765 PAND2X1_349/A POR2X1_73/Y 0.03fF
C30766 VDD PAND2X1_336/Y 0.21fF
C30767 PAND2X1_639/B POR2X1_583/Y 0.21fF
C30768 PAND2X1_284/Y PAND2X1_570/B 0.02fF
C30769 PAND2X1_308/Y PAND2X1_302/O 0.04fF
C30770 POR2X1_287/B POR2X1_343/CTRL 0.01fF
C30771 PAND2X1_371/CTRL2 POR2X1_773/A 0.10fF
C30772 PAND2X1_63/Y POR2X1_101/Y 0.03fF
C30773 PAND2X1_623/Y POR2X1_129/Y 0.01fF
C30774 PAND2X1_6/A POR2X1_260/A 0.07fF
C30775 POR2X1_326/A POR2X1_802/B 0.00fF
C30776 POR2X1_327/Y POR2X1_662/Y 0.19fF
C30777 POR2X1_715/A POR2X1_715/a_76_344# 0.03fF
C30778 PAND2X1_659/Y POR2X1_46/Y 0.03fF
C30779 POR2X1_7/A PAND2X1_338/B 0.03fF
C30780 POR2X1_101/a_76_344# PAND2X1_69/A 0.00fF
C30781 POR2X1_62/Y PAND2X1_523/O 0.07fF
C30782 POR2X1_538/a_16_28# POR2X1_703/A 0.04fF
C30783 PAND2X1_641/CTRL2 POR2X1_38/Y 0.05fF
C30784 PAND2X1_48/B POR2X1_722/CTRL2 0.02fF
C30785 INPUT_1 PAND2X1_69/A 3.01fF
C30786 POR2X1_456/B PAND2X1_32/B 3.36fF
C30787 POR2X1_145/a_16_28# POR2X1_394/A 0.03fF
C30788 POR2X1_235/CTRL POR2X1_7/A 0.01fF
C30789 POR2X1_119/Y PAND2X1_243/B 0.03fF
C30790 POR2X1_113/Y POR2X1_101/Y 0.03fF
C30791 POR2X1_499/A POR2X1_556/A 0.03fF
C30792 INPUT_1 POR2X1_93/A 0.29fF
C30793 POR2X1_833/A PAND2X1_150/CTRL 0.02fF
C30794 PAND2X1_437/CTRL2 POR2X1_590/A 0.02fF
C30795 PAND2X1_6/Y POR2X1_359/B 0.02fF
C30796 PAND2X1_93/B PAND2X1_85/CTRL 0.01fF
C30797 D_INPUT_3 POR2X1_4/CTRL2 0.01fF
C30798 POR2X1_356/A PAND2X1_167/O 0.16fF
C30799 PAND2X1_341/A POR2X1_153/Y 0.05fF
C30800 POR2X1_40/a_16_28# INPUT_6 0.03fF
C30801 POR2X1_853/A POR2X1_191/Y 0.05fF
C30802 POR2X1_614/A POR2X1_266/A 0.21fF
C30803 PAND2X1_511/CTRL2 PAND2X1_56/A 0.01fF
C30804 PAND2X1_211/CTRL POR2X1_20/B 0.01fF
C30805 POR2X1_228/a_56_344# POR2X1_631/B 0.00fF
C30806 PAND2X1_321/O PAND2X1_52/B 0.05fF
C30807 PAND2X1_501/CTRL PAND2X1_862/B 0.01fF
C30808 POR2X1_184/Y PAND2X1_141/O 0.00fF
C30809 POR2X1_93/A POR2X1_384/A 0.91fF
C30810 POR2X1_153/Y POR2X1_91/Y 0.13fF
C30811 POR2X1_588/Y POR2X1_260/A 0.03fF
C30812 PAND2X1_341/Y POR2X1_7/A 0.04fF
C30813 POR2X1_630/a_16_28# POR2X1_630/B 0.07fF
C30814 POR2X1_326/A POR2X1_532/A 0.00fF
C30815 POR2X1_609/Y PAND2X1_608/CTRL2 0.00fF
C30816 PAND2X1_471/B POR2X1_77/Y 0.01fF
C30817 POR2X1_76/A POR2X1_556/A 0.03fF
C30818 POR2X1_101/Y POR2X1_260/A 0.15fF
C30819 POR2X1_568/Y POR2X1_353/A 0.05fF
C30820 POR2X1_669/B POR2X1_667/CTRL2 0.01fF
C30821 PAND2X1_775/CTRL POR2X1_77/Y 0.01fF
C30822 POR2X1_730/Y POR2X1_151/O 0.01fF
C30823 PAND2X1_212/O POR2X1_20/B 0.17fF
C30824 POR2X1_57/A PAND2X1_730/A 0.00fF
C30825 POR2X1_728/B PAND2X1_52/B 0.44fF
C30826 PAND2X1_690/CTRL2 POR2X1_260/A 0.06fF
C30827 PAND2X1_462/O POR2X1_293/Y 0.03fF
C30828 PAND2X1_63/B POR2X1_186/B 0.03fF
C30829 POR2X1_553/CTRL2 POR2X1_569/A 0.05fF
C30830 POR2X1_357/CTRL POR2X1_568/Y 0.27fF
C30831 PAND2X1_608/CTRL POR2X1_102/Y 0.01fF
C30832 POR2X1_583/Y POR2X1_260/A 0.03fF
C30833 POR2X1_659/A POR2X1_222/CTRL 0.01fF
C30834 INPUT_1 PAND2X1_528/m4_208_n4# 0.07fF
C30835 POR2X1_86/CTRL2 POR2X1_73/Y 0.01fF
C30836 PAND2X1_860/A PAND2X1_473/B 0.03fF
C30837 PAND2X1_808/Y POR2X1_416/B 0.03fF
C30838 POR2X1_16/A PAND2X1_803/CTRL 0.01fF
C30839 POR2X1_394/A PAND2X1_514/O 0.02fF
C30840 PAND2X1_433/CTRL2 PAND2X1_72/A 0.01fF
C30841 POR2X1_463/CTRL POR2X1_750/B 0.01fF
C30842 PAND2X1_73/Y POR2X1_688/O 0.01fF
C30843 POR2X1_760/A POR2X1_594/CTRL 0.01fF
C30844 INPUT_1 PAND2X1_632/m4_208_n4# 0.15fF
C30845 POR2X1_813/O POR2X1_263/Y 0.09fF
C30846 PAND2X1_269/O POR2X1_72/B 0.01fF
C30847 POR2X1_168/CTRL POR2X1_566/B 0.14fF
C30848 PAND2X1_23/Y POR2X1_343/B 0.03fF
C30849 POR2X1_35/B POR2X1_621/O 0.01fF
C30850 POR2X1_841/CTRL POR2X1_590/A 0.01fF
C30851 POR2X1_383/A PAND2X1_304/CTRL2 0.00fF
C30852 POR2X1_23/Y PAND2X1_407/a_76_28# 0.01fF
C30853 POR2X1_411/B POR2X1_226/CTRL2 0.01fF
C30854 POR2X1_383/a_16_28# POR2X1_520/A 0.02fF
C30855 POR2X1_186/O POR2X1_326/A 0.01fF
C30856 POR2X1_83/B POR2X1_411/B 0.18fF
C30857 POR2X1_145/Y POR2X1_39/B 0.00fF
C30858 POR2X1_499/A POR2X1_474/O 0.11fF
C30859 POR2X1_48/A PAND2X1_590/CTRL2 0.00fF
C30860 POR2X1_846/Y POR2X1_615/CTRL2 0.01fF
C30861 PAND2X1_358/CTRL2 PAND2X1_656/A 0.01fF
C30862 PAND2X1_35/A PAND2X1_34/CTRL2 0.01fF
C30863 POR2X1_416/B POR2X1_108/O 0.01fF
C30864 PAND2X1_651/CTRL2 PAND2X1_639/Y 0.03fF
C30865 POR2X1_778/B POR2X1_717/B 0.03fF
C30866 POR2X1_203/Y PAND2X1_72/A 0.01fF
C30867 POR2X1_741/B POR2X1_188/Y 0.01fF
C30868 POR2X1_832/Y POR2X1_660/Y 0.03fF
C30869 POR2X1_20/B POR2X1_94/A 0.03fF
C30870 POR2X1_373/Y POR2X1_373/CTRL 0.01fF
C30871 POR2X1_89/Y PAND2X1_97/O -0.00fF
C30872 POR2X1_760/A PAND2X1_539/B 0.02fF
C30873 PAND2X1_865/Y PAND2X1_853/B 0.07fF
C30874 POR2X1_796/A PAND2X1_56/A 0.03fF
C30875 POR2X1_343/Y POR2X1_141/A 0.05fF
C30876 PAND2X1_269/a_76_28# INPUT_0 0.04fF
C30877 POR2X1_96/A PAND2X1_717/A 0.03fF
C30878 POR2X1_378/a_56_344# PAND2X1_9/Y 0.00fF
C30879 POR2X1_265/Y PAND2X1_341/B 0.01fF
C30880 POR2X1_78/A POR2X1_807/CTRL2 0.01fF
C30881 POR2X1_66/B PAND2X1_609/O 0.01fF
C30882 POR2X1_343/A PAND2X1_39/B 0.02fF
C30883 PAND2X1_96/B PAND2X1_125/O 0.05fF
C30884 POR2X1_54/Y PAND2X1_41/B 0.03fF
C30885 POR2X1_814/A POR2X1_776/B 0.07fF
C30886 POR2X1_812/A POR2X1_809/O 0.01fF
C30887 PAND2X1_65/B POR2X1_461/Y 0.03fF
C30888 POR2X1_99/CTRL VDD 0.00fF
C30889 POR2X1_632/B POR2X1_632/a_16_28# 0.03fF
C30890 PAND2X1_478/B PAND2X1_776/Y 0.02fF
C30891 POR2X1_650/A POR2X1_473/CTRL2 0.01fF
C30892 PAND2X1_806/a_76_28# PAND2X1_362/A 0.01fF
C30893 POR2X1_9/Y POR2X1_382/a_16_28# 0.08fF
C30894 POR2X1_227/A POR2X1_244/B 0.05fF
C30895 POR2X1_342/Y POR2X1_244/Y 0.00fF
C30896 POR2X1_394/A POR2X1_39/B 4.45fF
C30897 POR2X1_857/A VDD 0.00fF
C30898 PAND2X1_628/CTRL2 PAND2X1_88/Y 0.01fF
C30899 POR2X1_76/B PAND2X1_60/B 0.03fF
C30900 POR2X1_106/O POR2X1_102/Y 0.02fF
C30901 POR2X1_376/B POR2X1_699/CTRL2 0.00fF
C30902 POR2X1_51/A POR2X1_20/B 0.03fF
C30903 PAND2X1_73/O POR2X1_66/A 0.08fF
C30904 POR2X1_174/B POR2X1_174/A 0.01fF
C30905 PAND2X1_214/a_16_344# PAND2X1_214/A 0.02fF
C30906 PAND2X1_807/a_16_344# PAND2X1_221/Y 0.02fF
C30907 POR2X1_78/B POR2X1_624/Y 0.03fF
C30908 POR2X1_470/O POR2X1_466/Y 0.00fF
C30909 POR2X1_48/A PAND2X1_540/O 0.05fF
C30910 POR2X1_60/A PAND2X1_212/B 0.05fF
C30911 POR2X1_450/a_16_28# POR2X1_121/B 0.11fF
C30912 POR2X1_23/Y PAND2X1_474/A 0.03fF
C30913 POR2X1_329/A PAND2X1_6/A 0.19fF
C30914 PAND2X1_66/O POR2X1_5/Y 0.04fF
C30915 POR2X1_96/A PAND2X1_783/B 0.01fF
C30916 POR2X1_566/A POR2X1_471/A 0.31fF
C30917 POR2X1_648/A POR2X1_532/A 0.01fF
C30918 POR2X1_260/B POR2X1_410/CTRL 0.01fF
C30919 PAND2X1_23/Y POR2X1_444/CTRL 0.01fF
C30920 PAND2X1_222/a_56_28# INPUT_0 0.00fF
C30921 POR2X1_661/A POR2X1_796/A 0.07fF
C30922 PAND2X1_61/O PAND2X1_61/Y 0.01fF
C30923 POR2X1_846/A POR2X1_713/B 0.05fF
C30924 PAND2X1_73/Y POR2X1_186/Y 0.03fF
C30925 POR2X1_262/a_16_28# POR2X1_73/Y 0.02fF
C30926 PAND2X1_659/A POR2X1_498/Y 0.15fF
C30927 POR2X1_462/O PAND2X1_69/A 0.02fF
C30928 POR2X1_74/Y POR2X1_416/B 0.01fF
C30929 POR2X1_480/A POR2X1_66/A 0.10fF
C30930 POR2X1_433/O POR2X1_72/B 0.01fF
C30931 POR2X1_399/CTRL2 POR2X1_609/Y 0.03fF
C30932 POR2X1_492/CTRL2 POR2X1_60/A 0.01fF
C30933 POR2X1_32/A INPUT_7 0.05fF
C30934 POR2X1_322/a_16_28# POR2X1_441/Y 0.03fF
C30935 POR2X1_119/Y PAND2X1_862/CTRL 0.19fF
C30936 D_INPUT_5 PAND2X1_95/B 0.09fF
C30937 POR2X1_48/CTRL2 POR2X1_32/A 0.01fF
C30938 POR2X1_49/Y POR2X1_820/CTRL 0.01fF
C30939 POR2X1_66/B PAND2X1_16/CTRL2 0.01fF
C30940 POR2X1_849/A VDD 0.26fF
C30941 PAND2X1_61/Y POR2X1_60/A 0.03fF
C30942 POR2X1_66/B POR2X1_404/O 0.15fF
C30943 POR2X1_376/B POR2X1_83/B 3.98fF
C30944 PAND2X1_717/A POR2X1_7/A 0.03fF
C30945 POR2X1_496/Y POR2X1_627/a_76_344# 0.01fF
C30946 POR2X1_52/A PAND2X1_124/Y 0.03fF
C30947 POR2X1_72/B PAND2X1_168/Y 0.01fF
C30948 POR2X1_121/B POR2X1_362/B 0.03fF
C30949 PAND2X1_255/CTRL POR2X1_260/A 0.01fF
C30950 POR2X1_423/CTRL POR2X1_236/Y 0.12fF
C30951 PAND2X1_266/O POR2X1_7/A 0.03fF
C30952 PAND2X1_469/B POR2X1_679/A 0.13fF
C30953 POR2X1_104/O POR2X1_5/Y 0.09fF
C30954 PAND2X1_20/A PAND2X1_85/Y 0.07fF
C30955 POR2X1_830/CTRL POR2X1_830/A 0.08fF
C30956 POR2X1_32/A PAND2X1_579/B 0.03fF
C30957 POR2X1_777/B POR2X1_288/A 0.05fF
C30958 POR2X1_37/Y POR2X1_46/Y 0.02fF
C30959 PAND2X1_43/O PAND2X1_69/A 0.03fF
C30960 POR2X1_329/A POR2X1_385/CTRL 0.03fF
C30961 PAND2X1_95/B PAND2X1_31/CTRL 0.01fF
C30962 POR2X1_220/B POR2X1_468/B 0.03fF
C30963 PAND2X1_250/CTRL2 POR2X1_287/B 0.01fF
C30964 POR2X1_454/A D_GATE_222 0.07fF
C30965 POR2X1_567/B POR2X1_785/A 0.05fF
C30966 POR2X1_544/A POR2X1_174/A 0.07fF
C30967 POR2X1_683/CTRL POR2X1_669/B 0.01fF
C30968 POR2X1_188/A POR2X1_830/A 0.03fF
C30969 POR2X1_141/Y POR2X1_217/CTRL2 0.00fF
C30970 POR2X1_416/B POR2X1_320/Y 0.06fF
C30971 POR2X1_32/A INPUT_4 0.09fF
C30972 POR2X1_673/A POR2X1_673/CTRL 0.01fF
C30973 PAND2X1_90/A POR2X1_66/A 0.23fF
C30974 PAND2X1_623/Y POR2X1_37/Y 0.06fF
C30975 PAND2X1_195/O POR2X1_236/Y 0.02fF
C30976 POR2X1_13/A PAND2X1_721/B 0.01fF
C30977 POR2X1_411/B POR2X1_380/A 0.11fF
C30978 POR2X1_307/Y POR2X1_660/Y 0.01fF
C30979 PAND2X1_474/Y POR2X1_497/O 0.00fF
C30980 POR2X1_66/B POR2X1_87/Y 0.01fF
C30981 POR2X1_516/CTRL2 POR2X1_23/Y 0.01fF
C30982 POR2X1_466/A POR2X1_740/Y 0.05fF
C30983 PAND2X1_213/O PAND2X1_161/Y 0.01fF
C30984 POR2X1_148/CTRL POR2X1_532/A 0.01fF
C30985 POR2X1_287/B POR2X1_475/A 0.02fF
C30986 PAND2X1_20/A PAND2X1_89/CTRL2 0.00fF
C30987 POR2X1_366/Y POR2X1_269/CTRL 0.01fF
C30988 PAND2X1_23/Y POR2X1_843/CTRL2 0.01fF
C30989 PAND2X1_612/B POR2X1_649/B 0.02fF
C30990 PAND2X1_430/a_16_344# POR2X1_750/B 0.02fF
C30991 POR2X1_413/A PAND2X1_656/CTRL 0.01fF
C30992 POR2X1_52/A POR2X1_226/CTRL2 0.01fF
C30993 POR2X1_496/Y POR2X1_42/Y 0.10fF
C30994 POR2X1_814/B PAND2X1_85/Y 0.18fF
C30995 POR2X1_52/A POR2X1_83/B 1.41fF
C30996 PAND2X1_840/A POR2X1_37/Y 0.00fF
C30997 PAND2X1_20/A PAND2X1_226/CTRL2 0.03fF
C30998 POR2X1_39/B POR2X1_90/CTRL2 0.03fF
C30999 POR2X1_691/O POR2X1_811/A 0.00fF
C31000 POR2X1_414/Y VDD 0.01fF
C31001 POR2X1_632/CTRL PAND2X1_88/Y 0.01fF
C31002 PAND2X1_80/O PAND2X1_41/B 0.04fF
C31003 POR2X1_466/A POR2X1_732/O 0.04fF
C31004 POR2X1_254/Y PAND2X1_13/CTRL2 0.07fF
C31005 POR2X1_127/Y VDD 0.01fF
C31006 PAND2X1_108/O POR2X1_862/B 0.06fF
C31007 PAND2X1_222/A PAND2X1_799/O 0.00fF
C31008 PAND2X1_793/Y PAND2X1_557/A 0.75fF
C31009 POR2X1_634/A POR2X1_638/CTRL 0.14fF
C31010 PAND2X1_839/CTRL POR2X1_102/Y 0.01fF
C31011 POR2X1_398/Y VDD 0.01fF
C31012 POR2X1_83/B POR2X1_152/A 0.03fF
C31013 POR2X1_242/a_16_28# POR2X1_241/Y 0.09fF
C31014 PAND2X1_96/B POR2X1_476/A 0.04fF
C31015 POR2X1_121/A PAND2X1_73/Y 0.05fF
C31016 POR2X1_814/A PAND2X1_48/A 0.20fF
C31017 POR2X1_257/A PAND2X1_467/CTRL 0.01fF
C31018 POR2X1_177/Y POR2X1_236/Y 0.03fF
C31019 POR2X1_523/Y POR2X1_819/CTRL 0.01fF
C31020 POR2X1_123/B POR2X1_493/A 0.03fF
C31021 POR2X1_448/B VDD 0.16fF
C31022 POR2X1_254/Y POR2X1_702/B 0.10fF
C31023 POR2X1_624/Y POR2X1_141/A 0.02fF
C31024 PAND2X1_169/Y PAND2X1_714/O 0.16fF
C31025 POR2X1_16/A PAND2X1_9/Y 0.03fF
C31026 POR2X1_264/Y PAND2X1_265/O 0.03fF
C31027 POR2X1_56/B POR2X1_72/B 0.07fF
C31028 POR2X1_433/Y PAND2X1_435/Y 0.01fF
C31029 POR2X1_41/B PAND2X1_211/A 0.10fF
C31030 PAND2X1_96/B POR2X1_288/CTRL2 0.01fF
C31031 POR2X1_722/B POR2X1_602/B 0.00fF
C31032 PAND2X1_6/Y POR2X1_555/B 0.03fF
C31033 PAND2X1_807/B PAND2X1_794/B 0.00fF
C31034 POR2X1_333/A POR2X1_545/A 0.05fF
C31035 POR2X1_119/Y POR2X1_329/A 0.05fF
C31036 POR2X1_852/B POR2X1_776/B 0.07fF
C31037 POR2X1_602/B POR2X1_294/B 0.03fF
C31038 POR2X1_620/A POR2X1_620/a_16_28# 0.07fF
C31039 PAND2X1_733/A POR2X1_42/Y 0.03fF
C31040 PAND2X1_217/B PAND2X1_188/CTRL2 0.35fF
C31041 PAND2X1_657/CTRL POR2X1_816/A 0.01fF
C31042 PAND2X1_20/A PAND2X1_612/CTRL2 0.03fF
C31043 PAND2X1_54/O VDD 0.00fF
C31044 PAND2X1_453/O POR2X1_423/Y 0.06fF
C31045 PAND2X1_804/A PAND2X1_580/B 0.02fF
C31046 PAND2X1_570/a_76_28# PAND2X1_577/Y 0.04fF
C31047 POR2X1_65/A PAND2X1_364/CTRL 0.01fF
C31048 POR2X1_32/A POR2X1_73/Y 0.29fF
C31049 PAND2X1_115/Y PAND2X1_562/B 0.03fF
C31050 POR2X1_502/A PAND2X1_700/CTRL2 0.07fF
C31051 POR2X1_322/CTRL POR2X1_49/Y 0.08fF
C31052 POR2X1_730/CTRL POR2X1_330/Y 0.03fF
C31053 POR2X1_814/A POR2X1_330/CTRL2 0.02fF
C31054 PAND2X1_860/A PAND2X1_861/B 0.17fF
C31055 PAND2X1_472/A POR2X1_14/Y 0.03fF
C31056 POR2X1_833/A PAND2X1_39/B 0.07fF
C31057 PAND2X1_48/B POR2X1_637/A 0.00fF
C31058 POR2X1_96/A PAND2X1_541/a_76_28# 0.01fF
C31059 POR2X1_66/B POR2X1_66/CTRL2 0.03fF
C31060 POR2X1_66/A PAND2X1_397/CTRL2 0.01fF
C31061 POR2X1_60/A POR2X1_255/Y 0.02fF
C31062 POR2X1_167/Y POR2X1_166/Y 0.24fF
C31063 POR2X1_333/A POR2X1_317/Y 0.18fF
C31064 POR2X1_791/CTRL2 POR2X1_637/B 0.01fF
C31065 PAND2X1_818/a_76_28# POR2X1_376/B 0.01fF
C31066 POR2X1_66/A PAND2X1_305/O 0.06fF
C31067 PAND2X1_246/CTRL POR2X1_4/Y 0.01fF
C31068 PAND2X1_257/O POR2X1_632/Y 0.06fF
C31069 POR2X1_832/Y POR2X1_308/B 0.12fF
C31070 POR2X1_263/Y POR2X1_229/Y 0.00fF
C31071 PAND2X1_57/B VDD 2.95fF
C31072 POR2X1_623/A POR2X1_623/CTRL 0.01fF
C31073 POR2X1_79/Y PAND2X1_84/Y 0.01fF
C31074 PAND2X1_6/Y POR2X1_330/Y 0.17fF
C31075 POR2X1_198/B PAND2X1_65/Y 0.03fF
C31076 PAND2X1_193/O POR2X1_7/B 0.04fF
C31077 POR2X1_102/Y PAND2X1_575/O 0.11fF
C31078 POR2X1_52/A PAND2X1_140/Y 0.03fF
C31079 PAND2X1_467/B POR2X1_425/Y 0.02fF
C31080 GATE_479 POR2X1_693/Y 0.03fF
C31081 POR2X1_486/B POR2X1_486/O 0.05fF
C31082 PAND2X1_29/CTRL PAND2X1_41/B 0.01fF
C31083 PAND2X1_390/Y POR2X1_816/A 0.02fF
C31084 PAND2X1_688/O POR2X1_293/Y -0.01fF
C31085 PAND2X1_93/B PAND2X1_298/O 0.01fF
C31086 PAND2X1_456/O POR2X1_184/Y 0.02fF
C31087 POR2X1_66/B POR2X1_596/A 0.03fF
C31088 POR2X1_417/Y POR2X1_73/Y 0.16fF
C31089 POR2X1_78/B POR2X1_785/A 0.06fF
C31090 PAND2X1_245/CTRL2 PAND2X1_63/B 0.01fF
C31091 PAND2X1_20/A POR2X1_137/Y 0.03fF
C31092 PAND2X1_104/a_76_28# PAND2X1_6/A 0.07fF
C31093 POR2X1_823/Y POR2X1_102/Y 0.02fF
C31094 PAND2X1_23/Y PAND2X1_58/CTRL 0.00fF
C31095 POR2X1_788/A PAND2X1_60/B 0.03fF
C31096 POR2X1_52/A PAND2X1_795/B 0.03fF
C31097 POR2X1_680/Y VDD 0.01fF
C31098 POR2X1_443/O POR2X1_191/Y 0.26fF
C31099 POR2X1_41/B POR2X1_96/A 0.13fF
C31100 POR2X1_14/Y POR2X1_380/Y 0.16fF
C31101 POR2X1_78/B POR2X1_538/CTRL2 0.03fF
C31102 PAND2X1_552/B POR2X1_236/Y 0.01fF
C31103 POR2X1_346/B POR2X1_66/A 0.06fF
C31104 PAND2X1_808/Y PAND2X1_773/B 0.01fF
C31105 POR2X1_594/Y PAND2X1_362/B 0.00fF
C31106 PAND2X1_244/B POR2X1_32/A 0.03fF
C31107 POR2X1_356/A POR2X1_502/A 0.05fF
C31108 POR2X1_192/Y POR2X1_223/a_16_28# 0.02fF
C31109 PAND2X1_651/Y PAND2X1_456/O 0.02fF
C31110 POR2X1_624/Y POR2X1_294/A 0.03fF
C31111 POR2X1_66/B PAND2X1_60/CTRL2 0.00fF
C31112 POR2X1_673/Y POR2X1_849/A 0.09fF
C31113 POR2X1_283/Y PAND2X1_568/B 0.05fF
C31114 POR2X1_65/A POR2X1_90/Y 7.26fF
C31115 POR2X1_416/B POR2X1_827/a_16_28# 0.02fF
C31116 POR2X1_20/B PAND2X1_338/O 0.03fF
C31117 POR2X1_657/m4_208_n4# POR2X1_228/Y 0.08fF
C31118 POR2X1_48/A POR2X1_764/O 0.01fF
C31119 PAND2X1_137/O POR2X1_96/A 0.01fF
C31120 VDD PAND2X1_324/Y 0.15fF
C31121 POR2X1_380/O POR2X1_5/Y 0.11fF
C31122 POR2X1_515/CTRL POR2X1_68/A 0.14fF
C31123 POR2X1_46/Y POR2X1_293/Y 0.13fF
C31124 POR2X1_706/CTRL PAND2X1_94/A 0.01fF
C31125 POR2X1_302/CTRL PAND2X1_6/Y 0.02fF
C31126 PAND2X1_808/Y PAND2X1_738/Y 0.05fF
C31127 POR2X1_48/A POR2X1_394/A 0.31fF
C31128 POR2X1_102/Y POR2X1_172/CTRL2 0.01fF
C31129 POR2X1_48/A POR2X1_749/CTRL 0.09fF
C31130 POR2X1_333/A POR2X1_440/Y 0.15fF
C31131 POR2X1_664/CTRL2 POR2X1_78/A 0.03fF
C31132 POR2X1_664/CTRL PAND2X1_73/Y 0.01fF
C31133 POR2X1_567/B POR2X1_186/B 0.07fF
C31134 PAND2X1_494/CTRL INPUT_0 0.07fF
C31135 PAND2X1_862/B PAND2X1_575/A 0.04fF
C31136 POR2X1_188/A POR2X1_188/O 0.02fF
C31137 PAND2X1_474/Y POR2X1_56/Y 0.00fF
C31138 PAND2X1_57/B POR2X1_741/Y 0.10fF
C31139 PAND2X1_673/CTRL POR2X1_38/B 0.00fF
C31140 POR2X1_25/CTRL2 D_INPUT_6 0.01fF
C31141 POR2X1_814/B POR2X1_137/Y 0.08fF
C31142 POR2X1_855/B POR2X1_783/a_56_344# 0.00fF
C31143 POR2X1_830/Y POR2X1_456/B 0.00fF
C31144 PAND2X1_803/Y PAND2X1_562/B 0.03fF
C31145 POR2X1_244/B POR2X1_340/a_16_28# 0.02fF
C31146 POR2X1_447/B POR2X1_629/CTRL 0.08fF
C31147 POR2X1_376/B PAND2X1_168/CTRL2 0.00fF
C31148 POR2X1_828/A VDD 0.07fF
C31149 POR2X1_52/A PAND2X1_242/CTRL 0.01fF
C31150 PAND2X1_14/CTRL POR2X1_68/B 0.03fF
C31151 POR2X1_294/B PAND2X1_110/CTRL 0.06fF
C31152 POR2X1_13/A POR2X1_56/Y 0.06fF
C31153 POR2X1_222/Y POR2X1_553/Y 0.11fF
C31154 POR2X1_411/B PAND2X1_841/Y 0.01fF
C31155 POR2X1_65/A POR2X1_167/CTRL2 0.03fF
C31156 POR2X1_156/B POR2X1_155/CTRL 0.01fF
C31157 PAND2X1_41/B POR2X1_201/Y 0.03fF
C31158 PAND2X1_362/B PAND2X1_362/a_16_344# 0.02fF
C31159 POR2X1_542/B POR2X1_370/Y 0.03fF
C31160 POR2X1_326/A POR2X1_220/B 0.06fF
C31161 PAND2X1_223/B PAND2X1_538/CTRL2 0.01fF
C31162 POR2X1_40/Y POR2X1_384/a_76_344# 0.01fF
C31163 POR2X1_343/Y POR2X1_116/A 0.05fF
C31164 POR2X1_400/A POR2X1_206/CTRL 0.00fF
C31165 PAND2X1_472/A PAND2X1_472/B 0.01fF
C31166 PAND2X1_840/A POR2X1_293/Y 0.03fF
C31167 PAND2X1_4/CTRL2 PAND2X1_8/Y 0.03fF
C31168 POR2X1_60/O VDD 0.00fF
C31169 PAND2X1_408/O PAND2X1_52/B 0.02fF
C31170 POR2X1_49/Y POR2X1_521/Y 0.01fF
C31171 PAND2X1_57/B PAND2X1_32/B 1.03fF
C31172 POR2X1_614/A POR2X1_724/a_16_28# 0.01fF
C31173 PAND2X1_114/Y POR2X1_183/Y 0.00fF
C31174 POR2X1_243/Y POR2X1_532/A 0.07fF
C31175 PAND2X1_215/B PAND2X1_723/CTRL2 0.02fF
C31176 PAND2X1_239/a_56_28# POR2X1_192/B 0.00fF
C31177 PAND2X1_865/Y POR2X1_23/Y 0.00fF
C31178 PAND2X1_696/O POR2X1_866/A 0.02fF
C31179 POR2X1_383/A POR2X1_362/B 0.33fF
C31180 PAND2X1_35/Y POR2X1_73/Y 0.03fF
C31181 POR2X1_324/Y POR2X1_220/B 0.07fF
C31182 POR2X1_49/Y PAND2X1_737/B 0.03fF
C31183 POR2X1_68/A POR2X1_832/B 0.03fF
C31184 PAND2X1_6/Y POR2X1_247/O 0.16fF
C31185 POR2X1_193/A POR2X1_786/Y 0.05fF
C31186 POR2X1_294/B POR2X1_712/Y 0.03fF
C31187 POR2X1_120/O PAND2X1_60/B 0.01fF
C31188 PAND2X1_388/Y VDD 0.54fF
C31189 POR2X1_649/O PAND2X1_52/B 0.01fF
C31190 PAND2X1_6/Y PAND2X1_7/CTRL2 0.00fF
C31191 PAND2X1_197/CTRL POR2X1_52/Y 0.01fF
C31192 POR2X1_461/B POR2X1_713/B 0.29fF
C31193 POR2X1_122/O POR2X1_102/Y 0.01fF
C31194 POR2X1_285/B POR2X1_647/B 0.17fF
C31195 POR2X1_43/B POR2X1_238/Y 0.03fF
C31196 POR2X1_741/Y POR2X1_715/m4_208_n4# 0.12fF
C31197 POR2X1_41/B PAND2X1_850/m4_208_n4# 0.08fF
C31198 POR2X1_137/B POR2X1_768/A 0.02fF
C31199 POR2X1_78/A POR2X1_113/B 0.03fF
C31200 POR2X1_356/A PAND2X1_747/CTRL2 0.05fF
C31201 POR2X1_13/A PAND2X1_803/Y 0.03fF
C31202 PAND2X1_720/CTRL2 VDD 0.00fF
C31203 POR2X1_514/O POR2X1_514/Y 0.00fF
C31204 PAND2X1_94/A POR2X1_5/Y 1.29fF
C31205 PAND2X1_549/B VDD 0.67fF
C31206 PAND2X1_471/B PAND2X1_241/Y 0.16fF
C31207 PAND2X1_200/B POR2X1_40/Y 0.02fF
C31208 PAND2X1_653/O PAND2X1_267/Y 0.07fF
C31209 POR2X1_65/A PAND2X1_732/A 0.01fF
C31210 POR2X1_416/B PAND2X1_606/CTRL2 0.01fF
C31211 POR2X1_192/Y POR2X1_704/CTRL 0.45fF
C31212 POR2X1_428/CTRL2 POR2X1_236/Y 0.01fF
C31213 PAND2X1_472/B POR2X1_380/Y 0.02fF
C31214 POR2X1_57/A PAND2X1_215/B 0.07fF
C31215 PAND2X1_90/A POR2X1_532/A 0.07fF
C31216 PAND2X1_785/Y PAND2X1_349/A 0.03fF
C31217 POR2X1_60/CTRL2 PAND2X1_339/Y 0.00fF
C31218 POR2X1_599/A PAND2X1_717/a_76_28# 0.01fF
C31219 POR2X1_220/Y POR2X1_222/A 21.40fF
C31220 POR2X1_707/Y VDD 0.00fF
C31221 POR2X1_212/A POR2X1_212/B 0.00fF
C31222 POR2X1_654/O POR2X1_774/A 0.01fF
C31223 PAND2X1_866/O PAND2X1_805/A 0.02fF
C31224 POR2X1_41/B POR2X1_7/A 0.65fF
C31225 POR2X1_52/A POR2X1_131/m4_208_n4# 0.14fF
C31226 POR2X1_76/Y POR2X1_274/B 0.13fF
C31227 PAND2X1_857/A PAND2X1_661/O 0.05fF
C31228 PAND2X1_832/CTRL2 PAND2X1_508/Y 0.01fF
C31229 POR2X1_106/Y PAND2X1_348/A 0.08fF
C31230 PAND2X1_408/CTRL2 PAND2X1_32/B 0.01fF
C31231 POR2X1_614/A POR2X1_786/Y -0.00fF
C31232 POR2X1_184/Y POR2X1_73/Y 0.03fF
C31233 POR2X1_65/A PAND2X1_360/Y 0.03fF
C31234 POR2X1_644/A POR2X1_796/CTRL 0.06fF
C31235 PAND2X1_486/a_76_28# POR2X1_526/Y 0.00fF
C31236 PAND2X1_244/B PAND2X1_35/Y 0.03fF
C31237 POR2X1_771/A VDD 0.11fF
C31238 POR2X1_502/A PAND2X1_698/CTRL 0.00fF
C31239 PAND2X1_848/B POR2X1_382/Y 0.01fF
C31240 PAND2X1_787/Y POR2X1_129/Y 0.03fF
C31241 INPUT_0 PAND2X1_537/a_16_344# 0.00fF
C31242 POR2X1_460/a_16_28# POR2X1_460/A 0.03fF
C31243 PAND2X1_96/B POR2X1_513/Y 0.18fF
C31244 PAND2X1_631/A POR2X1_482/Y 0.02fF
C31245 POR2X1_96/A POR2X1_419/O 0.02fF
C31246 PAND2X1_651/Y POR2X1_73/Y 0.15fF
C31247 POR2X1_347/A POR2X1_402/B 0.00fF
C31248 POR2X1_574/O POR2X1_724/A 0.01fF
C31249 POR2X1_669/B POR2X1_39/B 0.39fF
C31250 POR2X1_158/Y POR2X1_695/Y 0.55fF
C31251 POR2X1_32/A PAND2X1_207/A 0.01fF
C31252 POR2X1_259/B VDD 0.12fF
C31253 POR2X1_508/O POR2X1_510/B 0.01fF
C31254 POR2X1_555/B POR2X1_632/Y 0.03fF
C31255 PAND2X1_48/CTRL2 POR2X1_186/B 0.01fF
C31256 POR2X1_69/Y PAND2X1_206/B 0.05fF
C31257 POR2X1_307/Y POR2X1_308/B 0.44fF
C31258 POR2X1_65/A POR2X1_110/Y 1.19fF
C31259 POR2X1_22/A POR2X1_36/m4_208_n4# 0.12fF
C31260 POR2X1_78/B POR2X1_186/B 0.10fF
C31261 POR2X1_445/O POR2X1_456/B 0.16fF
C31262 POR2X1_740/Y POR2X1_274/B 0.05fF
C31263 POR2X1_76/Y PAND2X1_72/Y 0.16fF
C31264 PAND2X1_41/B POR2X1_4/Y 0.19fF
C31265 POR2X1_16/A PAND2X1_216/O 0.01fF
C31266 POR2X1_96/A PAND2X1_308/Y 0.03fF
C31267 PAND2X1_844/B POR2X1_73/Y 0.01fF
C31268 PAND2X1_216/B PAND2X1_553/B 0.00fF
C31269 PAND2X1_56/Y POR2X1_553/A 0.05fF
C31270 POR2X1_283/A PAND2X1_365/B 0.01fF
C31271 POR2X1_845/CTRL2 D_INPUT_1 0.02fF
C31272 POR2X1_351/Y POR2X1_854/B 0.05fF
C31273 PAND2X1_23/Y POR2X1_260/A 0.36fF
C31274 PAND2X1_55/Y POR2X1_675/Y 0.06fF
C31275 POR2X1_9/Y POR2X1_818/O 0.06fF
C31276 POR2X1_377/O PAND2X1_94/A 0.20fF
C31277 POR2X1_21/O POR2X1_460/A 0.13fF
C31278 POR2X1_256/Y POR2X1_7/A 0.01fF
C31279 POR2X1_56/Y PAND2X1_510/B 0.03fF
C31280 POR2X1_38/Y PAND2X1_338/B 0.07fF
C31281 POR2X1_346/B POR2X1_222/Y 0.03fF
C31282 POR2X1_185/O PAND2X1_94/A 0.35fF
C31283 PAND2X1_422/O POR2X1_788/B 0.07fF
C31284 PAND2X1_467/Y POR2X1_694/CTRL2 0.01fF
C31285 POR2X1_277/CTRL PAND2X1_560/B 0.03fF
C31286 PAND2X1_445/CTRL2 PAND2X1_308/Y 0.01fF
C31287 PAND2X1_96/B POR2X1_366/A 0.03fF
C31288 D_INPUT_3 POR2X1_9/O 0.03fF
C31289 POR2X1_38/Y POR2X1_235/CTRL 0.02fF
C31290 D_INPUT_3 PAND2X1_509/a_76_28# 0.00fF
C31291 PAND2X1_625/O POR2X1_260/A 0.01fF
C31292 POR2X1_164/Y PAND2X1_565/A 0.05fF
C31293 PAND2X1_55/Y POR2X1_544/B 0.03fF
C31294 POR2X1_461/Y POR2X1_814/A 0.04fF
C31295 PAND2X1_79/Y PAND2X1_63/B 0.02fF
C31296 PAND2X1_23/Y POR2X1_363/A 0.07fF
C31297 POR2X1_93/a_16_28# POR2X1_283/A 0.03fF
C31298 PAND2X1_784/CTRL PAND2X1_156/A 0.26fF
C31299 POR2X1_143/CTRL PAND2X1_341/B 0.02fF
C31300 PAND2X1_859/A POR2X1_77/Y 0.23fF
C31301 PAND2X1_254/CTRL PAND2X1_508/Y 0.00fF
C31302 POR2X1_293/Y POR2X1_371/CTRL 0.02fF
C31303 PAND2X1_575/B PAND2X1_332/Y 0.03fF
C31304 POR2X1_330/Y PAND2X1_52/B 0.10fF
C31305 POR2X1_771/A PAND2X1_32/B 0.04fF
C31306 POR2X1_435/Y POR2X1_532/CTRL2 0.04fF
C31307 POR2X1_356/A POR2X1_188/Y 0.05fF
C31308 POR2X1_93/A POR2X1_384/a_16_28# 0.02fF
C31309 PAND2X1_190/Y PAND2X1_360/Y 0.55fF
C31310 POR2X1_356/A POR2X1_726/a_56_344# 0.03fF
C31311 PAND2X1_127/O PAND2X1_96/B 0.02fF
C31312 POR2X1_88/CTRL2 PAND2X1_206/B 0.00fF
C31313 PAND2X1_575/A PAND2X1_716/B 0.03fF
C31314 POR2X1_862/CTRL POR2X1_480/A 0.00fF
C31315 PAND2X1_118/a_76_28# POR2X1_559/A 0.04fF
C31316 POR2X1_327/Y POR2X1_804/A 0.06fF
C31317 PAND2X1_675/a_16_344# PAND2X1_740/Y -0.00fF
C31318 POR2X1_130/CTRL POR2X1_318/A 0.04fF
C31319 POR2X1_552/a_16_28# POR2X1_732/B 0.06fF
C31320 POR2X1_416/B PAND2X1_740/m4_208_n4# 0.12fF
C31321 PAND2X1_807/B PAND2X1_221/Y 0.04fF
C31322 POR2X1_96/A POR2X1_189/CTRL 0.01fF
C31323 POR2X1_192/Y POR2X1_567/CTRL2 0.01fF
C31324 POR2X1_99/B D_GATE_222 0.03fF
C31325 POR2X1_383/A POR2X1_734/CTRL 0.12fF
C31326 POR2X1_368/O POR2X1_416/B 0.01fF
C31327 POR2X1_278/Y POR2X1_416/B 0.07fF
C31328 PAND2X1_338/B POR2X1_153/Y 0.07fF
C31329 POR2X1_96/A POR2X1_77/Y 14.23fF
C31330 POR2X1_669/B POR2X1_827/O 0.01fF
C31331 POR2X1_566/A POR2X1_555/O 0.04fF
C31332 POR2X1_566/A PAND2X1_292/CTRL2 0.15fF
C31333 PAND2X1_152/CTRL POR2X1_711/Y 0.08fF
C31334 PAND2X1_474/CTRL2 PAND2X1_404/Y 0.03fF
C31335 PAND2X1_675/O PAND2X1_736/A 0.07fF
C31336 POR2X1_763/Y POR2X1_524/a_16_28# 0.03fF
C31337 POR2X1_583/Y POR2X1_584/Y 0.14fF
C31338 PAND2X1_335/O POR2X1_77/Y 0.01fF
C31339 PAND2X1_404/Y POR2X1_826/Y 0.03fF
C31340 POR2X1_493/O PAND2X1_48/A 0.16fF
C31341 POR2X1_43/O POR2X1_42/Y 0.01fF
C31342 POR2X1_502/A PAND2X1_72/A 0.18fF
C31343 POR2X1_111/Y PAND2X1_112/O 0.00fF
C31344 POR2X1_57/A POR2X1_119/Y 0.63fF
C31345 POR2X1_190/O POR2X1_188/Y 0.02fF
C31346 PAND2X1_349/A POR2X1_300/Y 0.80fF
C31347 PAND2X1_675/a_16_344# PAND2X1_675/A 0.01fF
C31348 PAND2X1_813/a_16_344# POR2X1_673/Y 0.02fF
C31349 POR2X1_845/A POR2X1_845/CTRL 0.01fF
C31350 POR2X1_685/A POR2X1_809/A 0.01fF
C31351 POR2X1_156/Y POR2X1_210/B 0.01fF
C31352 POR2X1_494/Y POR2X1_80/O 0.00fF
C31353 PAND2X1_313/O POR2X1_317/B 0.00fF
C31354 PAND2X1_94/A POR2X1_54/CTRL 0.01fF
C31355 POR2X1_67/Y PAND2X1_225/O 0.01fF
C31356 PAND2X1_632/B PAND2X1_508/Y 0.25fF
C31357 POR2X1_130/CTRL POR2X1_574/Y 0.00fF
C31358 POR2X1_532/A POR2X1_160/a_56_344# 0.00fF
C31359 POR2X1_180/B POR2X1_180/a_16_28# 0.03fF
C31360 PAND2X1_196/O PAND2X1_199/B 0.00fF
C31361 POR2X1_78/B PAND2X1_628/O 0.13fF
C31362 POR2X1_809/A POR2X1_260/A 0.02fF
C31363 PAND2X1_22/CTRL2 PAND2X1_3/A 0.01fF
C31364 POR2X1_814/A POR2X1_288/A 0.05fF
C31365 POR2X1_407/A PAND2X1_681/CTRL 0.01fF
C31366 POR2X1_86/Y PAND2X1_101/a_76_28# 0.02fF
C31367 PAND2X1_826/O POR2X1_294/Y 0.01fF
C31368 POR2X1_61/CTRL2 POR2X1_447/B 0.05fF
C31369 POR2X1_799/a_16_28# POR2X1_652/A 0.02fF
C31370 INPUT_2 POR2X1_416/B 0.05fF
C31371 POR2X1_84/B POR2X1_66/A 0.02fF
C31372 POR2X1_732/B POR2X1_181/A 0.21fF
C31373 PAND2X1_793/Y PAND2X1_860/A 0.02fF
C31374 POR2X1_205/A POR2X1_342/B 0.02fF
C31375 POR2X1_815/a_56_344# POR2X1_750/A 0.00fF
C31376 POR2X1_814/A POR2X1_193/Y 0.04fF
C31377 POR2X1_119/Y PAND2X1_301/O 0.11fF
C31378 POR2X1_62/Y POR2X1_394/A 0.05fF
C31379 PAND2X1_301/a_76_28# PAND2X1_716/B 0.02fF
C31380 POR2X1_383/A D_INPUT_4 0.07fF
C31381 PAND2X1_646/O POR2X1_609/Y 0.00fF
C31382 POR2X1_505/O PAND2X1_631/A 0.01fF
C31383 POR2X1_150/Y PAND2X1_558/Y 0.01fF
C31384 PAND2X1_840/A PAND2X1_242/Y 0.02fF
C31385 PAND2X1_405/CTRL POR2X1_46/Y 0.01fF
C31386 POR2X1_7/A POR2X1_77/Y 0.20fF
C31387 PAND2X1_831/CTRL POR2X1_411/B 0.01fF
C31388 PAND2X1_267/B POR2X1_72/B 0.03fF
C31389 POR2X1_85/Y POR2X1_7/A 1.85fF
C31390 POR2X1_820/a_16_28# POR2X1_411/B 0.03fF
C31391 PAND2X1_853/B PAND2X1_352/Y 0.03fF
C31392 POR2X1_14/Y POR2X1_260/B 0.03fF
C31393 POR2X1_48/A POR2X1_669/B 0.57fF
C31394 POR2X1_539/A POR2X1_325/B 0.09fF
C31395 POR2X1_685/A POR2X1_728/A 0.58fF
C31396 POR2X1_273/Y POR2X1_677/Y 0.42fF
C31397 PAND2X1_856/a_76_28# PAND2X1_854/Y 0.02fF
C31398 POR2X1_13/A PAND2X1_97/Y 0.03fF
C31399 PAND2X1_419/O POR2X1_296/B 0.21fF
C31400 PAND2X1_3/A PAND2X1_11/Y 0.13fF
C31401 POR2X1_260/B POR2X1_405/CTRL 0.01fF
C31402 POR2X1_799/CTRL PAND2X1_72/A 0.07fF
C31403 POR2X1_79/m4_208_n4# PAND2X1_798/m4_208_n4# 0.13fF
C31404 POR2X1_41/B POR2X1_760/A 6.89fF
C31405 POR2X1_442/CTRL POR2X1_236/Y 0.01fF
C31406 POR2X1_424/Y POR2X1_236/Y 0.00fF
C31407 POR2X1_728/A POR2X1_260/A 0.00fF
C31408 POR2X1_118/Y POR2X1_72/B 0.15fF
C31409 PAND2X1_404/Y PAND2X1_500/a_56_28# 0.00fF
C31410 POR2X1_566/A POR2X1_443/CTRL 0.05fF
C31411 PAND2X1_480/B POR2X1_150/Y 0.13fF
C31412 PAND2X1_20/A POR2X1_97/A 1.51fF
C31413 POR2X1_66/B D_INPUT_0 0.03fF
C31414 POR2X1_191/CTRL2 POR2X1_191/Y 0.03fF
C31415 POR2X1_707/B PAND2X1_25/CTRL 0.01fF
C31416 POR2X1_275/A POR2X1_46/Y 0.03fF
C31417 POR2X1_162/CTRL2 POR2X1_161/Y 0.01fF
C31418 PAND2X1_9/Y PAND2X1_57/B 0.03fF
C31419 POR2X1_12/A POR2X1_2/O 0.01fF
C31420 POR2X1_11/a_76_344# INPUT_4 0.00fF
C31421 POR2X1_188/A D_INPUT_0 0.03fF
C31422 POR2X1_250/Y PAND2X1_794/B 0.03fF
C31423 POR2X1_730/B POR2X1_814/A 0.09fF
C31424 POR2X1_237/Y POR2X1_329/A 0.09fF
C31425 PAND2X1_603/CTRL POR2X1_750/B 0.00fF
C31426 POR2X1_830/O POR2X1_590/A 0.01fF
C31427 PAND2X1_436/O PAND2X1_499/Y 0.01fF
C31428 POR2X1_490/CTRL PAND2X1_215/B 0.01fF
C31429 PAND2X1_58/A PAND2X1_585/CTRL 0.01fF
C31430 PAND2X1_259/O PAND2X1_555/A 0.02fF
C31431 INPUT_2 PAND2X1_608/CTRL 0.01fF
C31432 POR2X1_43/B PAND2X1_447/CTRL 0.01fF
C31433 POR2X1_119/Y PAND2X1_339/CTRL 0.29fF
C31434 PAND2X1_353/Y POR2X1_39/B 2.19fF
C31435 POR2X1_450/B PAND2X1_427/CTRL 0.01fF
C31436 POR2X1_41/Y POR2X1_39/B 0.00fF
C31437 POR2X1_815/Y INPUT_0 0.02fF
C31438 POR2X1_415/A POR2X1_7/B 0.02fF
C31439 PAND2X1_211/CTRL2 POR2X1_55/Y 0.01fF
C31440 POR2X1_809/A PAND2X1_681/O 0.02fF
C31441 POR2X1_590/A POR2X1_734/A 0.19fF
C31442 POR2X1_624/Y PAND2X1_110/CTRL2 0.01fF
C31443 POR2X1_159/a_16_28# POR2X1_669/B 0.02fF
C31444 POR2X1_679/CTRL2 POR2X1_816/A 0.01fF
C31445 PAND2X1_39/B POR2X1_294/B 8.03fF
C31446 POR2X1_480/A POR2X1_220/B 0.07fF
C31447 POR2X1_360/A POR2X1_202/A 0.02fF
C31448 PAND2X1_23/Y POR2X1_610/Y 0.08fF
C31449 PAND2X1_464/B PAND2X1_785/O 0.04fF
C31450 PAND2X1_423/O POR2X1_78/A 0.03fF
C31451 POR2X1_467/Y POR2X1_330/Y 0.05fF
C31452 PAND2X1_225/CTRL POR2X1_750/B 0.02fF
C31453 POR2X1_669/B PAND2X1_199/A 0.01fF
C31454 POR2X1_337/Y POR2X1_212/B 0.07fF
C31455 PAND2X1_57/B POR2X1_818/Y 0.03fF
C31456 POR2X1_411/B PAND2X1_357/Y 0.06fF
C31457 PAND2X1_72/A POR2X1_188/Y 0.02fF
C31458 POR2X1_614/A POR2X1_452/CTRL2 0.03fF
C31459 PAND2X1_212/CTRL2 POR2X1_55/Y 0.01fF
C31460 POR2X1_296/CTRL POR2X1_68/B 0.00fF
C31461 POR2X1_130/A POR2X1_218/Y 0.10fF
C31462 PAND2X1_58/A PAND2X1_395/O 0.02fF
C31463 PAND2X1_793/O POR2X1_29/A 0.03fF
C31464 PAND2X1_58/A PAND2X1_589/CTRL2 0.01fF
C31465 POR2X1_294/CTRL D_GATE_741 0.02fF
C31466 POR2X1_556/A PAND2X1_69/A 0.04fF
C31467 POR2X1_20/B PAND2X1_182/O 0.17fF
C31468 POR2X1_634/A POR2X1_710/A 0.39fF
C31469 POR2X1_14/Y PAND2X1_803/A 0.03fF
C31470 POR2X1_446/B POR2X1_659/CTRL 0.01fF
C31471 POR2X1_477/A POR2X1_434/CTRL 0.01fF
C31472 POR2X1_83/B PAND2X1_180/O 0.01fF
C31473 PAND2X1_217/B PAND2X1_476/O 0.02fF
C31474 POR2X1_260/B POR2X1_55/Y 0.05fF
C31475 PAND2X1_13/CTRL POR2X1_750/B 0.29fF
C31476 POR2X1_555/A POR2X1_630/A 0.03fF
C31477 PAND2X1_644/Y PAND2X1_758/CTRL 0.00fF
C31478 POR2X1_23/Y POR2X1_494/Y 0.03fF
C31479 POR2X1_66/B PAND2X1_90/Y 0.18fF
C31480 POR2X1_260/B PAND2X1_536/CTRL 0.01fF
C31481 PAND2X1_785/Y POR2X1_32/A 0.74fF
C31482 POR2X1_84/a_16_28# POR2X1_84/B 0.02fF
C31483 POR2X1_604/Y INPUT_0 0.78fF
C31484 PAND2X1_224/CTRL2 POR2X1_590/A 0.02fF
C31485 PAND2X1_448/CTRL2 POR2X1_42/Y 0.02fF
C31486 POR2X1_188/A PAND2X1_90/Y 0.05fF
C31487 PAND2X1_106/CTRL POR2X1_556/A 0.01fF
C31488 PAND2X1_611/O POR2X1_249/Y 0.02fF
C31489 POR2X1_14/Y PAND2X1_673/Y 0.03fF
C31490 POR2X1_114/B POR2X1_841/B 0.03fF
C31491 PAND2X1_777/a_16_344# POR2X1_7/B 0.01fF
C31492 PAND2X1_78/O PAND2X1_580/B 0.00fF
C31493 POR2X1_244/CTRL VDD 0.00fF
C31494 POR2X1_76/CTRL POR2X1_724/A 0.08fF
C31495 POR2X1_84/B POR2X1_532/A 0.44fF
C31496 POR2X1_760/A POR2X1_385/a_56_344# 0.00fF
C31497 POR2X1_376/B PAND2X1_783/Y 0.64fF
C31498 PAND2X1_39/B PAND2X1_111/B 0.03fF
C31499 POR2X1_60/A POR2X1_46/Y 0.12fF
C31500 PAND2X1_717/A POR2X1_153/Y 0.03fF
C31501 POR2X1_334/A PAND2X1_86/CTRL2 0.00fF
C31502 POR2X1_297/O POR2X1_297/Y 0.01fF
C31503 PAND2X1_6/Y PAND2X1_258/O 0.17fF
C31504 PAND2X1_221/m4_208_n4# PAND2X1_738/Y 0.04fF
C31505 POR2X1_805/Y POR2X1_294/B 0.19fF
C31506 PAND2X1_459/Y POR2X1_94/A 0.06fF
C31507 POR2X1_343/A VDD 0.05fF
C31508 POR2X1_423/Y POR2X1_516/B 0.05fF
C31509 POR2X1_76/A PAND2X1_60/B 0.00fF
C31510 POR2X1_673/a_16_28# PAND2X1_8/Y 0.06fF
C31511 PAND2X1_58/A POR2X1_832/B 1.06fF
C31512 POR2X1_804/CTRL2 POR2X1_532/A 0.01fF
C31513 PAND2X1_20/A POR2X1_294/B 0.27fF
C31514 POR2X1_62/CTRL PAND2X1_58/A 0.03fF
C31515 POR2X1_65/A INPUT_0 0.30fF
C31516 POR2X1_234/A POR2X1_39/B 0.07fF
C31517 POR2X1_435/B POR2X1_796/A 0.01fF
C31518 POR2X1_174/B POR2X1_795/B 0.05fF
C31519 POR2X1_315/O POR2X1_32/A 0.01fF
C31520 POR2X1_278/Y PAND2X1_192/Y 0.03fF
C31521 POR2X1_475/A PAND2X1_372/CTRL2 0.03fF
C31522 POR2X1_226/a_16_28# POR2X1_42/Y 0.06fF
C31523 PAND2X1_85/Y VDD 0.33fF
C31524 PAND2X1_90/O POR2X1_814/A 0.02fF
C31525 PAND2X1_444/Y POR2X1_152/A 0.04fF
C31526 POR2X1_51/A INPUT_7 0.00fF
C31527 POR2X1_763/Y PAND2X1_731/B 0.04fF
C31528 PAND2X1_201/CTRL PAND2X1_358/A 0.03fF
C31529 PAND2X1_56/Y POR2X1_830/CTRL2 0.28fF
C31530 PAND2X1_159/a_76_28# POR2X1_7/B 0.01fF
C31531 POR2X1_65/A POR2X1_424/O 0.01fF
C31532 POR2X1_859/A PAND2X1_90/Y 0.07fF
C31533 POR2X1_467/O POR2X1_210/A 0.01fF
C31534 POR2X1_43/B PAND2X1_195/CTRL2 0.01fF
C31535 POR2X1_45/Y POR2X1_40/Y 0.03fF
C31536 POR2X1_493/a_16_28# POR2X1_493/A 0.03fF
C31537 PAND2X1_63/Y POR2X1_641/CTRL2 0.16fF
C31538 POR2X1_514/CTRL2 POR2X1_777/B 0.33fF
C31539 POR2X1_63/Y PAND2X1_560/B 0.03fF
C31540 PAND2X1_675/A PAND2X1_540/CTRL2 0.03fF
C31541 POR2X1_814/B POR2X1_294/B 0.06fF
C31542 POR2X1_366/Y POR2X1_814/B 0.07fF
C31543 POR2X1_78/A POR2X1_341/Y 0.03fF
C31544 POR2X1_743/O POR2X1_7/B 0.01fF
C31545 D_GATE_662 PAND2X1_41/B 0.07fF
C31546 POR2X1_670/CTRL POR2X1_42/Y 0.01fF
C31547 PAND2X1_55/CTRL PAND2X1_55/Y 0.01fF
C31548 POR2X1_835/Y VDD 0.16fF
C31549 PAND2X1_6/Y POR2X1_457/O 0.01fF
C31550 POR2X1_438/Y PAND2X1_569/B 0.08fF
C31551 POR2X1_72/B PAND2X1_565/CTRL2 0.01fF
C31552 POR2X1_231/a_16_28# POR2X1_186/Y 0.03fF
C31553 POR2X1_14/Y POR2X1_583/CTRL2 0.00fF
C31554 PAND2X1_469/B PAND2X1_390/Y 0.03fF
C31555 POR2X1_407/A POR2X1_602/B 0.03fF
C31556 PAND2X1_787/Y POR2X1_293/Y 0.03fF
C31557 POR2X1_376/B POR2X1_697/Y 0.03fF
C31558 PAND2X1_341/B POR2X1_65/a_76_344# -0.00fF
C31559 POR2X1_278/Y PAND2X1_738/Y 0.31fF
C31560 PAND2X1_860/A PAND2X1_862/O 0.04fF
C31561 POR2X1_814/A POR2X1_343/CTRL2 0.03fF
C31562 POR2X1_186/Y POR2X1_35/Y 0.03fF
C31563 PAND2X1_643/Y PAND2X1_719/Y 0.06fF
C31564 PAND2X1_474/A PAND2X1_658/B 0.09fF
C31565 POR2X1_97/A POR2X1_212/O 0.02fF
C31566 POR2X1_296/B POR2X1_575/CTRL 0.00fF
C31567 PAND2X1_558/O POR2X1_494/Y 0.00fF
C31568 POR2X1_71/Y PAND2X1_474/Y 0.02fF
C31569 POR2X1_32/A PAND2X1_656/A 0.03fF
C31570 POR2X1_808/A POR2X1_828/A 0.20fF
C31571 PAND2X1_206/O POR2X1_293/Y 0.05fF
C31572 PAND2X1_58/A PAND2X1_757/CTRL 0.01fF
C31573 POR2X1_62/a_16_28# POR2X1_94/A 0.01fF
C31574 POR2X1_777/B POR2X1_576/Y 0.05fF
C31575 POR2X1_366/Y POR2X1_325/A 0.01fF
C31576 POR2X1_483/A POR2X1_740/Y 0.05fF
C31577 POR2X1_51/A INPUT_4 0.03fF
C31578 POR2X1_462/B PAND2X1_41/B 0.03fF
C31579 PAND2X1_272/CTRL POR2X1_553/A 0.01fF
C31580 D_INPUT_0 POR2X1_575/a_16_28# 0.03fF
C31581 POR2X1_615/Y VDD 0.00fF
C31582 POR2X1_13/A PAND2X1_668/O 0.02fF
C31583 PAND2X1_6/Y POR2X1_543/A 0.01fF
C31584 POR2X1_662/a_16_28# POR2X1_353/A 0.08fF
C31585 PAND2X1_20/A PAND2X1_111/B 0.03fF
C31586 POR2X1_440/Y POR2X1_436/B 0.06fF
C31587 PAND2X1_731/B POR2X1_73/Y 0.02fF
C31588 PAND2X1_41/B D_INPUT_1 0.33fF
C31589 POR2X1_78/A POR2X1_590/CTRL2 0.01fF
C31590 PAND2X1_242/O POR2X1_511/Y 0.08fF
C31591 POR2X1_120/m4_208_n4# POR2X1_608/m4_208_n4# 0.13fF
C31592 POR2X1_722/A POR2X1_866/A 0.10fF
C31593 POR2X1_546/B POR2X1_546/A 0.02fF
C31594 POR2X1_183/Y POR2X1_106/Y 0.00fF
C31595 PAND2X1_94/A PAND2X1_282/O 0.12fF
C31596 PAND2X1_786/O POR2X1_91/Y 0.37fF
C31597 POR2X1_93/A POR2X1_72/B 0.26fF
C31598 PAND2X1_673/Y POR2X1_55/Y 0.03fF
C31599 POR2X1_208/A POR2X1_201/CTRL2 0.00fF
C31600 POR2X1_72/B POR2X1_91/Y 0.03fF
C31601 POR2X1_123/A POR2X1_633/A 0.13fF
C31602 POR2X1_13/A POR2X1_42/Y 0.64fF
C31603 INPUT_1 PAND2X1_623/O 0.07fF
C31604 POR2X1_56/B POR2X1_7/B 0.05fF
C31605 POR2X1_722/B POR2X1_513/B 0.03fF
C31606 POR2X1_96/A PAND2X1_742/B 0.03fF
C31607 POR2X1_294/B POR2X1_513/B 0.13fF
C31608 POR2X1_548/CTRL2 POR2X1_68/B 0.05fF
C31609 PAND2X1_462/B POR2X1_232/CTRL2 0.02fF
C31610 PAND2X1_865/O POR2X1_102/Y 0.02fF
C31611 POR2X1_119/Y POR2X1_271/CTRL2 0.07fF
C31612 POR2X1_302/O POR2X1_513/Y 0.01fF
C31613 PAND2X1_90/A POR2X1_786/A 0.03fF
C31614 POR2X1_193/A POR2X1_193/CTRL2 0.01fF
C31615 POR2X1_52/A POR2X1_697/Y 0.01fF
C31616 PAND2X1_433/a_16_344# POR2X1_722/Y 0.03fF
C31617 POR2X1_5/Y POR2X1_382/Y 0.03fF
C31618 PAND2X1_785/Y POR2X1_184/Y 0.03fF
C31619 PAND2X1_6/A POR2X1_224/O 0.01fF
C31620 POR2X1_566/A POR2X1_68/A 0.23fF
C31621 POR2X1_32/A PAND2X1_348/A 0.03fF
C31622 POR2X1_814/B PAND2X1_111/B 0.03fF
C31623 PAND2X1_91/O POR2X1_191/Y 0.17fF
C31624 POR2X1_78/B POR2X1_542/B 0.03fF
C31625 POR2X1_685/O POR2X1_685/B 0.11fF
C31626 PAND2X1_52/Y POR2X1_228/Y 0.01fF
C31627 POR2X1_502/A POR2X1_793/A 0.03fF
C31628 POR2X1_266/A POR2X1_66/A 0.06fF
C31629 PAND2X1_439/a_16_344# POR2X1_167/Y 0.01fF
C31630 POR2X1_78/B PAND2X1_79/Y 0.03fF
C31631 POR2X1_544/B POR2X1_174/A 0.03fF
C31632 POR2X1_16/A PAND2X1_403/B 0.01fF
C31633 PAND2X1_341/B POR2X1_23/Y 0.05fF
C31634 POR2X1_96/A POR2X1_52/Y 0.02fF
C31635 PAND2X1_200/CTRL2 POR2X1_153/Y 0.05fF
C31636 PAND2X1_55/Y PAND2X1_536/CTRL 0.02fF
C31637 POR2X1_528/Y POR2X1_376/B 0.03fF
C31638 POR2X1_62/Y POR2X1_620/A 0.01fF
C31639 PAND2X1_833/CTRL2 POR2X1_283/A 0.01fF
C31640 POR2X1_32/A POR2X1_300/Y 0.05fF
C31641 POR2X1_836/O POR2X1_192/B 0.08fF
C31642 POR2X1_836/CTRL2 POR2X1_191/Y 0.00fF
C31643 POR2X1_525/Y PAND2X1_546/CTRL 0.01fF
C31644 POR2X1_416/B PAND2X1_634/a_16_344# 0.02fF
C31645 POR2X1_174/CTRL POR2X1_175/A 0.01fF
C31646 PAND2X1_6/Y PAND2X1_369/CTRL2 0.01fF
C31647 POR2X1_305/a_16_28# POR2X1_90/Y 0.03fF
C31648 POR2X1_639/Y PAND2X1_57/B 0.03fF
C31649 POR2X1_137/Y VDD 0.36fF
C31650 POR2X1_62/Y POR2X1_669/B 0.05fF
C31651 PAND2X1_814/CTRL2 POR2X1_7/B 0.03fF
C31652 PAND2X1_245/CTRL PAND2X1_48/A 0.01fF
C31653 POR2X1_57/A POR2X1_693/CTRL2 0.01fF
C31654 PAND2X1_649/A POR2X1_48/A 0.02fF
C31655 POR2X1_775/A D_GATE_222 0.22fF
C31656 PAND2X1_206/A PAND2X1_358/a_56_28# 0.00fF
C31657 POR2X1_250/CTRL2 POR2X1_283/A 0.01fF
C31658 POR2X1_41/B POR2X1_38/Y 0.08fF
C31659 PAND2X1_442/O POR2X1_568/Y 0.04fF
C31660 POR2X1_511/Y POR2X1_527/Y 0.22fF
C31661 POR2X1_707/a_16_28# POR2X1_707/A 0.05fF
C31662 POR2X1_57/A PAND2X1_661/O 0.04fF
C31663 POR2X1_417/O POR2X1_372/Y 0.06fF
C31664 POR2X1_327/Y POR2X1_794/B 0.07fF
C31665 POR2X1_13/A PAND2X1_99/Y 0.01fF
C31666 PAND2X1_94/A PAND2X1_65/B 0.17fF
C31667 PAND2X1_621/O POR2X1_847/B 0.03fF
C31668 POR2X1_237/Y PAND2X1_445/O 0.02fF
C31669 POR2X1_158/Y POR2X1_428/Y 0.03fF
C31670 PAND2X1_90/Y PAND2X1_313/CTRL 0.01fF
C31671 POR2X1_334/B PAND2X1_63/Y 0.19fF
C31672 PAND2X1_96/B POR2X1_832/B 0.01fF
C31673 PAND2X1_631/A POR2X1_32/A 0.07fF
C31674 PAND2X1_643/Y POR2X1_42/Y 0.03fF
C31675 POR2X1_66/A PAND2X1_179/O 0.06fF
C31676 PAND2X1_308/a_16_344# POR2X1_306/Y 0.05fF
C31677 POR2X1_698/a_56_344# POR2X1_394/A 0.00fF
C31678 POR2X1_455/CTRL POR2X1_456/B 0.01fF
C31679 POR2X1_335/A POR2X1_804/A 0.05fF
C31680 POR2X1_729/O POR2X1_614/A 0.01fF
C31681 PAND2X1_207/O POR2X1_39/B 0.01fF
C31682 POR2X1_614/A PAND2X1_599/a_76_28# 0.02fF
C31683 POR2X1_68/A POR2X1_844/B 0.05fF
C31684 PAND2X1_35/Y PAND2X1_656/A 0.03fF
C31685 POR2X1_89/CTRL2 PAND2X1_333/Y 0.01fF
C31686 POR2X1_856/B PAND2X1_167/a_76_28# 0.02fF
C31687 POR2X1_519/O VDD 0.00fF
C31688 POR2X1_740/Y POR2X1_209/A 0.00fF
C31689 POR2X1_135/a_56_344# POR2X1_32/A 0.00fF
C31690 POR2X1_567/A PAND2X1_20/A 0.07fF
C31691 PAND2X1_127/CTRL POR2X1_78/B 0.09fF
C31692 POR2X1_301/a_16_28# POR2X1_335/A 0.03fF
C31693 POR2X1_468/B POR2X1_854/B 0.03fF
C31694 POR2X1_390/B POR2X1_302/Y 0.02fF
C31695 POR2X1_66/B POR2X1_61/A 0.01fF
C31696 POR2X1_180/B POR2X1_566/A 0.08fF
C31697 POR2X1_730/Y POR2X1_155/CTRL 0.03fF
C31698 PAND2X1_8/Y PAND2X1_133/a_16_344# 0.01fF
C31699 PAND2X1_197/CTRL2 PAND2X1_656/A 0.01fF
C31700 POR2X1_57/A PAND2X1_334/CTRL 0.01fF
C31701 POR2X1_52/A POR2X1_528/Y 0.20fF
C31702 POR2X1_57/A POR2X1_57/a_16_28# 0.03fF
C31703 POR2X1_114/B POR2X1_458/B 0.33fF
C31704 POR2X1_672/A POR2X1_38/B 0.01fF
C31705 POR2X1_68/A POR2X1_573/A 0.03fF
C31706 POR2X1_65/A POR2X1_110/CTRL2 0.03fF
C31707 POR2X1_833/A VDD 0.07fF
C31708 PAND2X1_41/B POR2X1_620/B 0.01fF
C31709 PAND2X1_824/B POR2X1_400/A 0.07fF
C31710 POR2X1_334/CTRL2 POR2X1_360/A 0.04fF
C31711 PAND2X1_631/A POR2X1_417/Y 0.19fF
C31712 PAND2X1_48/B POR2X1_738/A 1.41fF
C31713 POR2X1_493/A PAND2X1_72/A 0.06fF
C31714 POR2X1_68/B PAND2X1_518/CTRL 0.00fF
C31715 PAND2X1_550/O POR2X1_394/A 0.02fF
C31716 PAND2X1_732/CTRL2 POR2X1_39/B 0.01fF
C31717 POR2X1_43/B POR2X1_387/Y 0.08fF
C31718 PAND2X1_636/CTRL POR2X1_583/Y 0.01fF
C31719 PAND2X1_109/O POR2X1_78/A 0.10fF
C31720 POR2X1_41/B INPUT_1 0.61fF
C31721 POR2X1_567/A POR2X1_776/CTRL2 0.11fF
C31722 PAND2X1_810/A GATE_865 0.12fF
C31723 POR2X1_299/a_56_344# POR2X1_90/Y 0.00fF
C31724 POR2X1_777/B PAND2X1_136/CTRL2 0.33fF
C31725 PAND2X1_79/CTRL POR2X1_569/A 0.03fF
C31726 POR2X1_334/A INPUT_0 0.03fF
C31727 PAND2X1_435/CTRL POR2X1_153/Y 0.04fF
C31728 POR2X1_567/A POR2X1_814/B 4.18fF
C31729 POR2X1_316/O INPUT_0 0.02fF
C31730 POR2X1_124/B POR2X1_113/Y 0.03fF
C31731 POR2X1_347/A POR2X1_360/A 0.02fF
C31732 POR2X1_137/Y PAND2X1_32/B 0.04fF
C31733 POR2X1_355/B POR2X1_333/Y 0.03fF
C31734 POR2X1_7/A POR2X1_52/Y 0.01fF
C31735 PAND2X1_651/Y PAND2X1_656/A 0.05fF
C31736 VDD PAND2X1_18/B 0.63fF
C31737 POR2X1_41/B POR2X1_153/Y 0.21fF
C31738 POR2X1_733/A POR2X1_260/A 0.03fF
C31739 PAND2X1_73/Y POR2X1_715/CTRL2 0.01fF
C31740 POR2X1_75/O PAND2X1_349/A 0.01fF
C31741 POR2X1_305/CTRL2 POR2X1_40/Y 0.01fF
C31742 POR2X1_334/B POR2X1_260/A 0.19fF
C31743 PAND2X1_659/Y PAND2X1_741/CTRL2 0.03fF
C31744 POR2X1_114/CTRL POR2X1_101/Y 0.15fF
C31745 POR2X1_183/Y PAND2X1_114/B 0.04fF
C31746 POR2X1_119/Y PAND2X1_84/Y 0.27fF
C31747 PAND2X1_844/O POR2X1_293/Y 0.01fF
C31748 POR2X1_228/Y POR2X1_724/A 0.07fF
C31749 PAND2X1_795/B PAND2X1_716/B 11.10fF
C31750 POR2X1_48/A POR2X1_234/A 0.04fF
C31751 POR2X1_502/A POR2X1_722/CTRL 0.01fF
C31752 POR2X1_53/O INPUT_5 0.00fF
C31753 PAND2X1_651/Y PAND2X1_861/CTRL2 0.49fF
C31754 POR2X1_596/A POR2X1_780/B 0.01fF
C31755 PAND2X1_6/Y POR2X1_348/a_16_28# 0.02fF
C31756 POR2X1_245/CTRL POR2X1_245/Y 0.02fF
C31757 POR2X1_687/A POR2X1_828/A 0.91fF
C31758 PAND2X1_23/Y POR2X1_559/A 0.10fF
C31759 POR2X1_537/Y POR2X1_502/A 0.03fF
C31760 POR2X1_65/A PAND2X1_809/B 0.02fF
C31761 POR2X1_730/Y POR2X1_467/CTRL 0.01fF
C31762 POR2X1_334/Y POR2X1_785/A 0.07fF
C31763 PAND2X1_314/O POR2X1_854/B 0.29fF
C31764 POR2X1_222/Y POR2X1_507/A 0.07fF
C31765 POR2X1_824/a_16_28# POR2X1_236/Y 0.03fF
C31766 POR2X1_614/A PAND2X1_813/CTRL2 0.00fF
C31767 POR2X1_366/Y POR2X1_703/CTRL2 0.03fF
C31768 POR2X1_707/B PAND2X1_72/A 0.03fF
C31769 PAND2X1_838/B POR2X1_827/a_16_28# 0.01fF
C31770 PAND2X1_653/Y PAND2X1_737/B 0.03fF
C31771 POR2X1_639/Y POR2X1_707/Y 0.03fF
C31772 POR2X1_390/B POR2X1_501/B 0.03fF
C31773 PAND2X1_74/O PAND2X1_72/A 0.04fF
C31774 POR2X1_206/a_16_28# POR2X1_201/Y 0.03fF
C31775 POR2X1_537/A PAND2X1_60/B 0.05fF
C31776 POR2X1_264/Y POR2X1_557/B 0.03fF
C31777 POR2X1_68/A POR2X1_344/Y 0.49fF
C31778 POR2X1_347/CTRL PAND2X1_57/B 0.01fF
C31779 POR2X1_840/B POR2X1_456/B 0.03fF
C31780 PAND2X1_350/a_16_344# POR2X1_7/A 0.01fF
C31781 POR2X1_119/Y PAND2X1_659/a_76_28# 0.03fF
C31782 POR2X1_5/Y PAND2X1_198/O 0.03fF
C31783 PAND2X1_48/B POR2X1_349/CTRL 0.01fF
C31784 POR2X1_322/Y PAND2X1_374/O 0.00fF
C31785 POR2X1_510/Y POR2X1_569/A 0.07fF
C31786 PAND2X1_499/Y POR2X1_39/B 0.04fF
C31787 PAND2X1_193/Y POR2X1_32/A 0.03fF
C31788 POR2X1_416/B POR2X1_743/CTRL 0.01fF
C31789 PAND2X1_107/a_16_344# POR2X1_532/A 0.06fF
C31790 PAND2X1_640/O POR2X1_153/Y 0.04fF
C31791 PAND2X1_229/CTRL PAND2X1_72/A 0.01fF
C31792 PAND2X1_793/Y PAND2X1_860/CTRL2 0.01fF
C31793 POR2X1_184/Y POR2X1_300/Y 0.03fF
C31794 POR2X1_207/B PAND2X1_824/B 0.01fF
C31795 POR2X1_16/A PAND2X1_213/Y 0.03fF
C31796 POR2X1_566/A POR2X1_181/O 0.32fF
C31797 POR2X1_464/CTRL POR2X1_736/A 0.29fF
C31798 PAND2X1_860/A POR2X1_516/Y 0.03fF
C31799 PAND2X1_221/Y PAND2X1_798/O 0.00fF
C31800 POR2X1_566/A POR2X1_169/A 0.05fF
C31801 PAND2X1_73/Y POR2X1_643/CTRL 0.08fF
C31802 POR2X1_451/a_16_28# POR2X1_750/B 0.03fF
C31803 PAND2X1_798/B POR2X1_385/Y 0.10fF
C31804 PAND2X1_352/O POR2X1_55/Y 0.04fF
C31805 POR2X1_332/B POR2X1_632/Y 0.09fF
C31806 PAND2X1_162/A PAND2X1_161/Y 0.00fF
C31807 POR2X1_416/B PAND2X1_730/B 0.02fF
C31808 POR2X1_83/Y PAND2X1_339/Y 0.02fF
C31809 POR2X1_394/A POR2X1_152/Y 0.00fF
C31810 POR2X1_293/Y PAND2X1_860/a_16_344# 0.01fF
C31811 POR2X1_257/A PAND2X1_247/CTRL2 0.13fF
C31812 POR2X1_502/O POR2X1_854/B 0.02fF
C31813 POR2X1_776/B POR2X1_568/B 0.01fF
C31814 PAND2X1_6/Y POR2X1_342/O 0.17fF
C31815 INPUT_1 PAND2X1_528/CTRL2 0.07fF
C31816 PAND2X1_18/B PAND2X1_32/B 1.82fF
C31817 POR2X1_779/CTRL2 POR2X1_513/B 0.01fF
C31818 POR2X1_266/A POR2X1_532/A 0.02fF
C31819 PAND2X1_631/A POR2X1_184/Y 0.35fF
C31820 POR2X1_218/O POR2X1_260/A 0.11fF
C31821 POR2X1_771/A POR2X1_769/Y 0.04fF
C31822 POR2X1_390/B POR2X1_703/A -0.03fF
C31823 POR2X1_456/B POR2X1_737/O 0.16fF
C31824 POR2X1_865/B PAND2X1_48/A 0.02fF
C31825 POR2X1_42/CTRL POR2X1_4/Y 0.05fF
C31826 POR2X1_131/a_16_28# POR2X1_131/A 0.03fF
C31827 PAND2X1_631/A PAND2X1_651/Y 0.03fF
C31828 PAND2X1_48/B POR2X1_731/Y 0.05fF
C31829 POR2X1_559/A POR2X1_520/A 0.01fF
C31830 POR2X1_130/A POR2X1_138/A 0.07fF
C31831 POR2X1_490/Y PAND2X1_217/O 0.01fF
C31832 POR2X1_83/B POR2X1_431/CTRL2 0.04fF
C31833 PAND2X1_462/B POR2X1_416/B 0.05fF
C31834 POR2X1_326/A POR2X1_854/B 0.05fF
C31835 POR2X1_532/A POR2X1_691/A 0.01fF
C31836 POR2X1_73/Y POR2X1_150/a_16_28# 0.01fF
C31837 POR2X1_188/A POR2X1_643/a_76_344# 0.00fF
C31838 PAND2X1_699/O POR2X1_496/Y 0.09fF
C31839 POR2X1_83/B POR2X1_250/Y 0.01fF
C31840 POR2X1_680/m4_208_n4# PAND2X1_652/A 0.08fF
C31841 PAND2X1_853/B POR2X1_310/Y 0.02fF
C31842 POR2X1_65/A POR2X1_292/CTRL2 0.02fF
C31843 POR2X1_567/B POR2X1_776/A 0.74fF
C31844 POR2X1_57/A PAND2X1_326/B 0.04fF
C31845 POR2X1_343/Y POR2X1_218/A 0.13fF
C31846 PAND2X1_562/Y PAND2X1_771/Y 0.32fF
C31847 POR2X1_324/Y POR2X1_854/B 0.02fF
C31848 POR2X1_691/B POR2X1_691/A 0.02fF
C31849 POR2X1_713/Y POR2X1_711/Y 0.01fF
C31850 POR2X1_327/Y POR2X1_741/B 0.08fF
C31851 POR2X1_633/A POR2X1_633/CTRL 0.01fF
C31852 POR2X1_77/O POR2X1_48/A 0.02fF
C31853 POR2X1_490/Y PAND2X1_124/Y 0.00fF
C31854 POR2X1_334/Y POR2X1_186/B 0.07fF
C31855 POR2X1_38/Y POR2X1_77/Y 0.11fF
C31856 PAND2X1_172/m4_208_n4# PAND2X1_189/m4_208_n4# 0.05fF
C31857 POR2X1_825/Y POR2X1_293/Y 0.03fF
C31858 POR2X1_508/B PAND2X1_823/O 0.00fF
C31859 POR2X1_85/Y POR2X1_38/Y 0.02fF
C31860 POR2X1_607/A POR2X1_411/B 0.00fF
C31861 POR2X1_143/CTRL2 POR2X1_9/Y 0.02fF
C31862 POR2X1_804/A POR2X1_715/CTRL 0.00fF
C31863 POR2X1_659/a_16_28# POR2X1_750/B 0.08fF
C31864 POR2X1_456/B POR2X1_564/a_76_344# 0.01fF
C31865 PAND2X1_640/B POR2X1_118/Y 0.03fF
C31866 POR2X1_454/CTRL POR2X1_454/B 0.01fF
C31867 POR2X1_567/B POR2X1_856/B 0.03fF
C31868 POR2X1_640/Y POR2X1_556/A 0.01fF
C31869 POR2X1_137/B PAND2X1_41/B 0.07fF
C31870 POR2X1_349/O POR2X1_363/A 0.07fF
C31871 POR2X1_335/B POR2X1_717/B 0.00fF
C31872 POR2X1_725/Y POR2X1_711/Y 0.00fF
C31873 POR2X1_49/Y POR2X1_603/a_16_28# 0.03fF
C31874 POR2X1_502/A POR2X1_848/a_56_344# 0.00fF
C31875 POR2X1_415/A POR2X1_750/B 0.07fF
C31876 PAND2X1_497/O POR2X1_78/A 0.05fF
C31877 POR2X1_496/m4_208_n4# PAND2X1_58/A 0.07fF
C31878 POR2X1_510/Y PAND2X1_72/A 0.03fF
C31879 POR2X1_527/O POR2X1_39/B 0.18fF
C31880 POR2X1_48/A PAND2X1_732/CTRL2 0.03fF
C31881 POR2X1_20/B PAND2X1_721/O 0.05fF
C31882 PAND2X1_488/a_76_28# POR2X1_556/A 0.02fF
C31883 PAND2X1_477/a_16_344# POR2X1_102/Y 0.02fF
C31884 POR2X1_119/Y PAND2X1_858/a_16_344# 0.03fF
C31885 POR2X1_150/Y PAND2X1_473/B 0.06fF
C31886 INPUT_1 POR2X1_77/Y 0.10fF
C31887 PAND2X1_39/B POR2X1_807/A 0.20fF
C31888 PAND2X1_771/Y PAND2X1_542/a_16_344# 0.07fF
C31889 POR2X1_16/A POR2X1_416/B 0.56fF
C31890 PAND2X1_557/A PAND2X1_267/Y 0.03fF
C31891 POR2X1_60/A PAND2X1_571/A 0.01fF
C31892 D_INPUT_0 POR2X1_413/O 0.18fF
C31893 PAND2X1_9/Y PAND2X1_85/Y 0.01fF
C31894 PAND2X1_412/CTRL2 POR2X1_260/B 0.03fF
C31895 POR2X1_49/Y PAND2X1_404/Y 0.05fF
C31896 POR2X1_276/Y PAND2X1_72/A 0.03fF
C31897 D_INPUT_5 PAND2X1_588/O 0.15fF
C31898 PAND2X1_601/CTRL POR2X1_718/A 0.10fF
C31899 POR2X1_816/O POR2X1_859/A 0.01fF
C31900 POR2X1_329/A PAND2X1_575/A 0.03fF
C31901 PAND2X1_282/a_76_28# POR2X1_590/A 0.02fF
C31902 POR2X1_454/A PAND2X1_52/Y 0.02fF
C31903 POR2X1_77/Y POR2X1_153/Y 0.12fF
C31904 POR2X1_102/Y PAND2X1_792/O 0.01fF
C31905 POR2X1_326/CTRL2 POR2X1_568/A 0.01fF
C31906 POR2X1_85/Y POR2X1_153/Y 0.05fF
C31907 PAND2X1_722/O PAND2X1_719/Y 0.00fF
C31908 PAND2X1_722/CTRL PAND2X1_718/Y 0.01fF
C31909 PAND2X1_860/A PAND2X1_843/Y 0.00fF
C31910 POR2X1_661/A POR2X1_513/CTRL 0.03fF
C31911 POR2X1_448/O POR2X1_296/B 0.04fF
C31912 POR2X1_760/A PAND2X1_742/B -0.00fF
C31913 PAND2X1_831/Y POR2X1_677/Y 0.00fF
C31914 PAND2X1_230/CTRL POR2X1_78/A 0.03fF
C31915 PAND2X1_576/B PAND2X1_576/O 0.03fF
C31916 PAND2X1_687/a_76_28# POR2X1_761/A 0.01fF
C31917 POR2X1_355/O POR2X1_567/B 0.01fF
C31918 PAND2X1_865/Y POR2X1_184/CTRL2 0.00fF
C31919 POR2X1_66/A POR2X1_734/A 0.42fF
C31920 POR2X1_376/B POR2X1_817/O 0.02fF
C31921 POR2X1_29/Y PAND2X1_87/O 0.10fF
C31922 PAND2X1_61/a_76_28# POR2X1_60/A 0.01fF
C31923 PAND2X1_281/CTRL2 PAND2X1_52/B 0.01fF
C31924 POR2X1_437/CTRL PAND2X1_580/B 0.00fF
C31925 POR2X1_634/A PAND2X1_58/A 0.05fF
C31926 POR2X1_675/A POR2X1_466/A 0.24fF
C31927 POR2X1_60/A POR2X1_251/CTRL 0.00fF
C31928 POR2X1_621/a_16_28# PAND2X1_6/A 0.01fF
C31929 INPUT_3 POR2X1_618/O 0.02fF
C31930 POR2X1_23/Y POR2X1_497/Y 0.03fF
C31931 POR2X1_760/A POR2X1_52/Y 0.03fF
C31932 POR2X1_150/Y PAND2X1_390/O 0.03fF
C31933 PAND2X1_47/B POR2X1_750/B 0.01fF
C31934 POR2X1_662/Y POR2X1_663/B 0.03fF
C31935 POR2X1_78/A PAND2X1_41/B 5.72fF
C31936 POR2X1_16/A POR2X1_16/O 0.05fF
C31937 POR2X1_78/B POR2X1_856/B 0.10fF
C31938 PAND2X1_434/O INPUT_0 0.05fF
C31939 POR2X1_814/A POR2X1_307/A 0.05fF
C31940 POR2X1_52/A POR2X1_816/Y 0.01fF
C31941 POR2X1_815/A POR2X1_7/B 0.02fF
C31942 POR2X1_705/B POR2X1_705/CTRL 0.00fF
C31943 POR2X1_624/B POR2X1_38/B 0.12fF
C31944 INPUT_3 POR2X1_619/CTRL 0.01fF
C31945 POR2X1_83/B PAND2X1_205/Y 0.15fF
C31946 POR2X1_65/A POR2X1_102/Y 0.71fF
C31947 POR2X1_76/B POR2X1_574/Y 0.18fF
C31948 POR2X1_41/B POR2X1_248/A 0.03fF
C31949 POR2X1_308/CTRL2 POR2X1_660/Y 0.01fF
C31950 POR2X1_814/A POR2X1_360/O 0.09fF
C31951 PAND2X1_97/CTRL2 POR2X1_293/Y 0.10fF
C31952 POR2X1_63/Y PAND2X1_734/CTRL2 0.01fF
C31953 POR2X1_334/B POR2X1_473/O 0.11fF
C31954 PAND2X1_65/B PAND2X1_11/Y 0.27fF
C31955 POR2X1_97/A VDD 0.69fF
C31956 PAND2X1_85/Y PAND2X1_15/O 0.06fF
C31957 POR2X1_102/Y PAND2X1_558/CTRL 0.01fF
C31958 PAND2X1_612/B POR2X1_642/O 0.00fF
C31959 POR2X1_669/B PAND2X1_550/O 0.05fF
C31960 POR2X1_407/A PAND2X1_39/B 0.15fF
C31961 PAND2X1_476/a_16_344# POR2X1_72/B 0.02fF
C31962 POR2X1_624/Y POR2X1_218/A 0.01fF
C31963 POR2X1_60/A PAND2X1_787/Y 0.00fF
C31964 POR2X1_356/A PAND2X1_237/a_16_344# 0.09fF
C31965 PAND2X1_806/CTRL2 POR2X1_42/Y 0.01fF
C31966 POR2X1_860/CTRL2 POR2X1_814/A 0.01fF
C31967 PAND2X1_794/O PAND2X1_473/B 0.03fF
C31968 POR2X1_257/A PAND2X1_565/A 0.03fF
C31969 POR2X1_347/B POR2X1_68/O 0.03fF
C31970 PAND2X1_790/a_76_28# POR2X1_42/Y 0.02fF
C31971 POR2X1_838/B VDD 0.00fF
C31972 PAND2X1_94/A POR2X1_814/A 0.03fF
C31973 PAND2X1_866/A PAND2X1_805/A 0.13fF
C31974 POR2X1_657/Y POR2X1_724/A 0.02fF
C31975 PAND2X1_289/CTRL POR2X1_210/Y 0.01fF
C31976 PAND2X1_289/CTRL2 POR2X1_220/A 0.03fF
C31977 POR2X1_836/B VDD 0.10fF
C31978 POR2X1_674/CTRL2 PAND2X1_742/B 0.01fF
C31979 POR2X1_20/B INPUT_6 0.03fF
C31980 POR2X1_124/B POR2X1_473/O 0.01fF
C31981 PAND2X1_561/Y VDD 0.04fF
C31982 POR2X1_130/A PAND2X1_58/A 0.06fF
C31983 POR2X1_130/A POR2X1_641/CTRL 0.03fF
C31984 PAND2X1_93/B POR2X1_130/Y 0.07fF
C31985 PAND2X1_96/B POR2X1_473/CTRL 0.01fF
C31986 POR2X1_66/A PAND2X1_144/CTRL2 0.01fF
C31987 POR2X1_355/B POR2X1_174/A 32.33fF
C31988 POR2X1_656/CTRL2 POR2X1_733/A 0.17fF
C31989 POR2X1_593/B PAND2X1_589/CTRL 0.01fF
C31990 POR2X1_448/m4_208_n4# PAND2X1_90/Y 0.03fF
C31991 PAND2X1_418/a_76_28# POR2X1_854/B 0.04fF
C31992 POR2X1_624/Y POR2X1_140/CTRL -0.03fF
C31993 POR2X1_260/B PAND2X1_743/CTRL2 0.01fF
C31994 POR2X1_590/A PAND2X1_372/O 0.21fF
C31995 POR2X1_36/B POR2X1_257/A 0.00fF
C31996 PAND2X1_845/CTRL2 POR2X1_23/Y 0.08fF
C31997 POR2X1_864/A POR2X1_796/A 0.03fF
C31998 PAND2X1_769/O POR2X1_764/Y 0.00fF
C31999 PAND2X1_65/B POR2X1_448/Y 0.01fF
C32000 PAND2X1_668/CTRL POR2X1_60/A 0.03fF
C32001 PAND2X1_93/B PAND2X1_72/CTRL 0.00fF
C32002 PAND2X1_658/O VDD 0.00fF
C32003 POR2X1_29/A POR2X1_42/Y 0.08fF
C32004 POR2X1_492/CTRL VDD 0.00fF
C32005 PAND2X1_492/O PAND2X1_41/B 0.17fF
C32006 PAND2X1_243/B POR2X1_83/B 0.13fF
C32007 PAND2X1_860/A PAND2X1_860/CTRL 0.10fF
C32008 POR2X1_376/B PAND2X1_712/B 0.01fF
C32009 PAND2X1_812/O PAND2X1_811/A 0.03fF
C32010 POR2X1_663/B POR2X1_181/B 0.01fF
C32011 PAND2X1_217/CTRL PAND2X1_723/A 0.01fF
C32012 PAND2X1_803/A POR2X1_511/Y 0.03fF
C32013 PAND2X1_472/A POR2X1_37/Y 0.03fF
C32014 PAND2X1_20/A POR2X1_546/B 0.12fF
C32015 POR2X1_66/A POR2X1_786/Y 0.07fF
C32016 POR2X1_224/CTRL2 POR2X1_226/Y 0.00fF
C32017 POR2X1_78/B POR2X1_786/CTRL2 0.04fF
C32018 POR2X1_857/CTRL POR2X1_795/B 0.01fF
C32019 POR2X1_650/A VDD 0.23fF
C32020 POR2X1_616/CTRL POR2X1_93/A 0.01fF
C32021 PAND2X1_699/CTRL POR2X1_129/Y 0.03fF
C32022 PAND2X1_423/CTRL PAND2X1_57/B 0.01fF
C32023 POR2X1_198/B POR2X1_201/CTRL2 0.03fF
C32024 INPUT_0 PAND2X1_729/m4_208_n4# 0.07fF
C32025 POR2X1_14/CTRL2 POR2X1_68/B 0.02fF
C32026 PAND2X1_6/A POR2X1_296/B 0.06fF
C32027 POR2X1_12/CTRL2 INPUT_4 0.05fF
C32028 PAND2X1_61/Y PAND2X1_351/Y 0.02fF
C32029 POR2X1_97/A PAND2X1_32/B 0.05fF
C32030 POR2X1_102/Y PAND2X1_190/Y 0.21fF
C32031 POR2X1_260/B POR2X1_366/A 0.03fF
C32032 POR2X1_200/O POR2X1_294/B 0.02fF
C32033 PAND2X1_93/B POR2X1_228/Y 0.03fF
C32034 GATE_479 POR2X1_46/Y 0.03fF
C32035 POR2X1_75/O POR2X1_32/A 0.01fF
C32036 PAND2X1_478/B POR2X1_238/Y 0.04fF
C32037 PAND2X1_94/CTRL PAND2X1_60/B 0.01fF
C32038 PAND2X1_20/A POR2X1_140/B 0.01fF
C32039 POR2X1_602/a_16_28# PAND2X1_60/B 0.02fF
C32040 PAND2X1_836/CTRL2 POR2X1_102/Y 0.01fF
C32041 PAND2X1_604/O POR2X1_750/B 0.06fF
C32042 PAND2X1_119/CTRL2 POR2X1_78/A 0.02fF
C32043 PAND2X1_119/CTRL PAND2X1_73/Y 0.00fF
C32044 POR2X1_66/B D_GATE_222 0.03fF
C32045 POR2X1_807/A POR2X1_513/B 0.03fF
C32046 POR2X1_110/Y PAND2X1_464/B 0.01fF
C32047 PAND2X1_58/A POR2X1_844/B 0.01fF
C32048 POR2X1_502/A PAND2X1_589/a_16_344# 0.01fF
C32049 PAND2X1_362/B VDD 0.26fF
C32050 PAND2X1_267/Y PAND2X1_723/A 0.02fF
C32051 PAND2X1_48/B PAND2X1_387/CTRL 0.01fF
C32052 PAND2X1_73/Y POR2X1_68/B 0.14fF
C32053 POR2X1_296/B PAND2X1_505/CTRL2 0.00fF
C32054 POR2X1_302/A PAND2X1_299/CTRL2 0.01fF
C32055 POR2X1_260/B POR2X1_375/O 0.01fF
C32056 POR2X1_832/A D_INPUT_0 0.03fF
C32057 POR2X1_66/B POR2X1_140/A 0.04fF
C32058 POR2X1_669/B POR2X1_152/Y 0.04fF
C32059 PAND2X1_640/B PAND2X1_559/CTRL2 0.03fF
C32060 POR2X1_220/B POR2X1_319/Y 0.03fF
C32061 POR2X1_78/B POR2X1_722/Y 0.03fF
C32062 POR2X1_49/Y POR2X1_528/CTRL 0.04fF
C32063 D_INPUT_0 POR2X1_780/B 0.00fF
C32064 POR2X1_60/Y PAND2X1_339/Y 0.01fF
C32065 POR2X1_548/CTRL2 PAND2X1_90/A 0.03fF
C32066 POR2X1_811/A POR2X1_780/B 0.00fF
C32067 POR2X1_13/A PAND2X1_139/Y 0.01fF
C32068 PAND2X1_140/A POR2X1_127/O 0.01fF
C32069 POR2X1_65/A PAND2X1_808/Y 0.03fF
C32070 POR2X1_809/Y POR2X1_121/B 0.03fF
C32071 POR2X1_96/A PAND2X1_580/B 0.03fF
C32072 POR2X1_657/O POR2X1_724/A 0.02fF
C32073 PAND2X1_862/B PAND2X1_573/CTRL 0.01fF
C32074 POR2X1_333/A POR2X1_532/A 0.03fF
C32075 POR2X1_827/O POR2X1_39/B 0.16fF
C32076 POR2X1_78/Y POR2X1_571/Y 0.63fF
C32077 PAND2X1_96/B POR2X1_634/A 0.40fF
C32078 POR2X1_510/A PAND2X1_41/B 0.03fF
C32079 POR2X1_78/A PAND2X1_424/a_16_344# 0.02fF
C32080 POR2X1_68/B POR2X1_390/a_16_28# 0.03fF
C32081 PAND2X1_736/A PAND2X1_736/O 0.00fF
C32082 POR2X1_341/A PAND2X1_48/A 0.03fF
C32083 POR2X1_68/A POR2X1_774/Y 0.14fF
C32084 POR2X1_842/CTRL POR2X1_456/B 0.01fF
C32085 PAND2X1_695/O PAND2X1_23/Y 0.02fF
C32086 POR2X1_45/Y POR2X1_5/Y 0.03fF
C32087 POR2X1_407/A POR2X1_814/B 0.03fF
C32088 POR2X1_722/B VDD 0.05fF
C32089 POR2X1_65/A POR2X1_531/Y 0.00fF
C32090 POR2X1_550/A POR2X1_78/A 0.01fF
C32091 POR2X1_858/B D_INPUT_0 0.03fF
C32092 POR2X1_294/B VDD 7.20fF
C32093 PAND2X1_857/A POR2X1_83/B 0.03fF
C32094 PAND2X1_495/a_76_28# PAND2X1_20/A 0.01fF
C32095 PAND2X1_20/A POR2X1_472/O 0.01fF
C32096 POR2X1_3/A POR2X1_40/Y 0.02fF
C32097 POR2X1_101/Y POR2X1_296/B 0.12fF
C32098 POR2X1_860/O POR2X1_218/Y 0.05fF
C32099 POR2X1_484/CTRL PAND2X1_726/B 0.08fF
C32100 PAND2X1_205/A POR2X1_394/A 0.03fF
C32101 POR2X1_498/a_16_28# POR2X1_46/Y 0.09fF
C32102 POR2X1_532/A POR2X1_734/A 0.10fF
C32103 POR2X1_43/B POR2X1_237/O -0.00fF
C32104 PAND2X1_48/B POR2X1_502/A 1.34fF
C32105 POR2X1_140/B POR2X1_325/A 0.03fF
C32106 POR2X1_865/B POR2X1_288/A 0.02fF
C32107 POR2X1_650/A PAND2X1_32/B 0.09fF
C32108 POR2X1_73/a_16_28# POR2X1_37/Y 0.04fF
C32109 PAND2X1_6/A POR2X1_236/Y 0.17fF
C32110 POR2X1_46/O PAND2X1_338/B 0.03fF
C32111 POR2X1_83/B PAND2X1_374/O 0.01fF
C32112 POR2X1_65/A POR2X1_821/Y 0.03fF
C32113 PAND2X1_61/Y PAND2X1_560/CTRL2 0.01fF
C32114 POR2X1_163/A PAND2X1_213/B 0.09fF
C32115 POR2X1_506/B POR2X1_566/B 0.03fF
C32116 PAND2X1_94/A POR2X1_650/O 0.02fF
C32117 POR2X1_482/Y POR2X1_7/A 0.03fF
C32118 PAND2X1_119/a_16_344# POR2X1_654/B 0.00fF
C32119 POR2X1_750/CTRL2 POR2X1_720/A 0.01fF
C32120 POR2X1_272/Y POR2X1_255/Y 0.00fF
C32121 POR2X1_326/a_56_344# POR2X1_220/B 0.00fF
C32122 POR2X1_193/A POR2X1_795/CTRL2 0.05fF
C32123 POR2X1_193/Y PAND2X1_88/Y 0.03fF
C32124 PAND2X1_48/B POR2X1_247/CTRL 0.01fF
C32125 POR2X1_599/A PAND2X1_735/Y 0.02fF
C32126 POR2X1_612/Y POR2X1_5/O 0.02fF
C32127 PAND2X1_48/B POR2X1_464/Y 0.72fF
C32128 POR2X1_401/CTRL PAND2X1_69/A 0.01fF
C32129 POR2X1_149/B POR2X1_220/Y 0.03fF
C32130 PAND2X1_213/B PAND2X1_162/CTRL2 0.01fF
C32131 PAND2X1_254/CTRL POR2X1_55/Y 0.00fF
C32132 PAND2X1_548/CTRL VDD 0.00fF
C32133 PAND2X1_94/A POR2X1_34/Y 0.01fF
C32134 POR2X1_96/A POR2X1_406/A 0.00fF
C32135 POR2X1_130/CTRL2 POR2X1_66/B 0.01fF
C32136 POR2X1_391/A POR2X1_391/O 0.00fF
C32137 POR2X1_114/B POR2X1_405/Y 0.01fF
C32138 POR2X1_851/CTRL POR2X1_590/A 0.01fF
C32139 POR2X1_396/Y POR2X1_5/Y 0.00fF
C32140 POR2X1_130/A PAND2X1_96/B 0.12fF
C32141 PAND2X1_516/CTRL POR2X1_513/Y 0.00fF
C32142 PAND2X1_675/A PAND2X1_592/Y 0.03fF
C32143 POR2X1_270/O POR2X1_78/B 0.05fF
C32144 POR2X1_523/Y POR2X1_7/B 0.03fF
C32145 POR2X1_114/B POR2X1_784/A 0.07fF
C32146 POR2X1_16/A POR2X1_487/Y 0.05fF
C32147 POR2X1_407/A POR2X1_513/B 10.15fF
C32148 PAND2X1_89/a_16_344# D_GATE_222 0.02fF
C32149 PAND2X1_36/CTRL PAND2X1_18/B 0.00fF
C32150 POR2X1_538/O POR2X1_193/A 0.02fF
C32151 POR2X1_745/Y VDD 0.00fF
C32152 POR2X1_366/Y POR2X1_741/Y 0.03fF
C32153 POR2X1_741/Y POR2X1_294/B 0.08fF
C32154 PAND2X1_688/a_16_344# POR2X1_38/Y 0.02fF
C32155 POR2X1_566/A PAND2X1_96/B 0.03fF
C32156 POR2X1_632/A POR2X1_510/Y 0.01fF
C32157 POR2X1_599/A PAND2X1_493/Y 1.26fF
C32158 POR2X1_76/Y POR2X1_541/CTRL2 0.01fF
C32159 POR2X1_43/B PAND2X1_341/CTRL 0.00fF
C32160 POR2X1_378/Y PAND2X1_69/A 0.03fF
C32161 PAND2X1_124/Y PAND2X1_199/a_56_28# 0.00fF
C32162 PAND2X1_224/CTRL2 POR2X1_532/A 0.01fF
C32163 PAND2X1_472/A POR2X1_293/Y 0.01fF
C32164 PAND2X1_6/Y POR2X1_579/Y 0.03fF
C32165 POR2X1_852/CTRL2 POR2X1_854/B 0.33fF
C32166 POR2X1_231/CTRL2 PAND2X1_32/B 0.03fF
C32167 POR2X1_614/A POR2X1_795/CTRL2 0.01fF
C32168 PAND2X1_94/A PAND2X1_55/CTRL2 0.01fF
C32169 POR2X1_441/Y PAND2X1_326/a_16_344# 0.01fF
C32170 PAND2X1_644/CTRL2 POR2X1_683/Y 0.00fF
C32171 POR2X1_60/m4_208_n4# POR2X1_497/Y 0.09fF
C32172 PAND2X1_111/B VDD 0.86fF
C32173 PAND2X1_243/O PAND2X1_35/Y 0.02fF
C32174 PAND2X1_69/A POR2X1_7/B 0.03fF
C32175 POR2X1_480/A POR2X1_854/B 0.07fF
C32176 PAND2X1_808/Y PAND2X1_190/Y 0.61fF
C32177 PAND2X1_700/a_76_28# POR2X1_532/A 0.01fF
C32178 POR2X1_296/B POR2X1_722/O 0.02fF
C32179 PAND2X1_665/O PAND2X1_93/B 0.06fF
C32180 POR2X1_41/B POR2X1_591/Y 0.07fF
C32181 POR2X1_68/B PAND2X1_132/CTRL2 0.08fF
C32182 PAND2X1_848/B POR2X1_382/O 0.02fF
C32183 PAND2X1_55/Y POR2X1_513/Y 0.97fF
C32184 POR2X1_219/B POR2X1_205/Y 0.19fF
C32185 PAND2X1_491/CTRL2 POR2X1_264/Y 0.01fF
C32186 POR2X1_802/B POR2X1_788/B 0.03fF
C32187 POR2X1_244/B POR2X1_510/Y 0.03fF
C32188 VDD POR2X1_351/CTRL 0.00fF
C32189 POR2X1_294/B PAND2X1_32/B 0.40fF
C32190 PAND2X1_55/Y POR2X1_219/B 0.07fF
C32191 POR2X1_158/Y POR2X1_695/O 0.00fF
C32192 POR2X1_32/A PAND2X1_199/CTRL 0.01fF
C32193 POR2X1_316/O PAND2X1_436/A 0.03fF
C32194 POR2X1_280/Y POR2X1_236/Y 0.00fF
C32195 POR2X1_93/A POR2X1_7/B 0.03fF
C32196 PAND2X1_717/Y VDD 0.20fF
C32197 POR2X1_308/CTRL2 POR2X1_308/B 0.01fF
C32198 POR2X1_456/a_16_28# POR2X1_456/B 0.07fF
C32199 POR2X1_189/m4_208_n4# PAND2X1_676/m4_208_n4# 0.15fF
C32200 POR2X1_184/Y POR2X1_183/Y 0.02fF
C32201 POR2X1_76/Y POR2X1_203/a_56_344# 0.01fF
C32202 POR2X1_7/B POR2X1_91/Y 0.03fF
C32203 PAND2X1_755/a_76_28# PAND2X1_60/B 0.01fF
C32204 POR2X1_423/Y PAND2X1_853/B 10.82fF
C32205 POR2X1_351/Y POR2X1_35/Y 0.03fF
C32206 PAND2X1_653/Y PAND2X1_218/O 0.07fF
C32207 POR2X1_112/O POR2X1_241/B 0.01fF
C32208 POR2X1_248/A POR2X1_77/Y 0.05fF
C32209 POR2X1_46/Y PAND2X1_175/B 0.03fF
C32210 POR2X1_96/A PAND2X1_349/A 0.03fF
C32211 PAND2X1_556/B PAND2X1_569/B 0.07fF
C32212 D_GATE_662 POR2X1_544/CTRL2 0.09fF
C32213 POR2X1_65/A POR2X1_165/Y 0.01fF
C32214 PAND2X1_65/m4_208_n4# POR2X1_342/m4_208_n4# 0.13fF
C32215 POR2X1_75/O POR2X1_184/Y 0.00fF
C32216 POR2X1_48/A POR2X1_39/B 1.40fF
C32217 POR2X1_614/A PAND2X1_6/Y 3.20fF
C32218 POR2X1_170/B POR2X1_169/Y 0.01fF
C32219 POR2X1_508/B POR2X1_506/B 0.00fF
C32220 POR2X1_583/O POR2X1_42/Y 0.01fF
C32221 POR2X1_60/A POR2X1_373/a_56_344# 0.00fF
C32222 POR2X1_335/A PAND2X1_311/O 0.03fF
C32223 POR2X1_25/Y POR2X1_40/Y 0.01fF
C32224 PAND2X1_864/CTRL GATE_741 0.01fF
C32225 POR2X1_283/A PAND2X1_364/CTRL 0.01fF
C32226 PAND2X1_94/A POR2X1_401/B 0.01fF
C32227 POR2X1_719/O PAND2X1_48/B 0.01fF
C32228 PAND2X1_55/Y POR2X1_736/a_56_344# 0.00fF
C32229 PAND2X1_716/O POR2X1_73/Y 0.04fF
C32230 POR2X1_16/A PAND2X1_738/Y 0.12fF
C32231 PAND2X1_96/B POR2X1_844/B 0.03fF
C32232 POR2X1_205/Y POR2X1_366/A 0.36fF
C32233 POR2X1_677/a_16_28# POR2X1_129/Y 0.06fF
C32234 POR2X1_407/Y PAND2X1_743/CTRL2 0.01fF
C32235 PAND2X1_6/Y POR2X1_38/B 0.06fF
C32236 POR2X1_57/A PAND2X1_794/B 0.03fF
C32237 POR2X1_60/Y PAND2X1_338/CTRL2 0.01fF
C32238 D_INPUT_3 POR2X1_43/B 0.05fF
C32239 PAND2X1_55/Y POR2X1_366/A 0.01fF
C32240 POR2X1_741/Y PAND2X1_111/B 0.01fF
C32241 POR2X1_537/Y POR2X1_862/B 1.90fF
C32242 POR2X1_38/Y POR2X1_52/Y 0.03fF
C32243 POR2X1_532/A POR2X1_786/Y 0.07fF
C32244 PAND2X1_386/a_16_344# PAND2X1_48/A 0.04fF
C32245 POR2X1_62/Y PAND2X1_340/CTRL 0.01fF
C32246 POR2X1_101/A POR2X1_243/Y 0.02fF
C32247 POR2X1_147/A PAND2X1_60/B 0.01fF
C32248 PAND2X1_693/CTRL POR2X1_383/A 0.01fF
C32249 PAND2X1_81/B PAND2X1_111/B 0.01fF
C32250 POR2X1_110/CTRL POR2X1_5/Y 0.01fF
C32251 POR2X1_407/Y POR2X1_770/O 0.01fF
C32252 POR2X1_205/O POR2X1_366/A 0.04fF
C32253 POR2X1_350/CTRL POR2X1_854/B 0.32fF
C32254 PAND2X1_96/B POR2X1_573/A 0.03fF
C32255 PAND2X1_484/CTRL INPUT_0 0.01fF
C32256 POR2X1_99/B PAND2X1_52/Y 0.00fF
C32257 PAND2X1_632/B POR2X1_55/Y 0.03fF
C32258 POR2X1_532/A POR2X1_788/B 0.04fF
C32259 POR2X1_337/O POR2X1_260/A 0.18fF
C32260 PAND2X1_6/Y PAND2X1_422/O 0.01fF
C32261 POR2X1_189/Y PAND2X1_728/CTRL 0.01fF
C32262 POR2X1_68/A POR2X1_799/CTRL2 0.05fF
C32263 POR2X1_680/O POR2X1_40/Y 0.01fF
C32264 POR2X1_760/A PAND2X1_405/a_76_28# 0.01fF
C32265 PAND2X1_69/A PAND2X1_60/B 2.66fF
C32266 PAND2X1_508/Y INPUT_0 0.12fF
C32267 D_INPUT_3 POR2X1_38/B 3.08fF
C32268 PAND2X1_111/B PAND2X1_32/B 0.16fF
C32269 PAND2X1_551/O POR2X1_90/Y 0.03fF
C32270 PAND2X1_57/B PAND2X1_399/O 0.04fF
C32271 POR2X1_55/Y PAND2X1_336/a_56_28# 0.00fF
C32272 POR2X1_119/Y POR2X1_236/Y 0.11fF
C32273 POR2X1_775/A POR2X1_175/B 0.01fF
C32274 POR2X1_466/a_16_28# POR2X1_453/Y -0.00fF
C32275 POR2X1_32/Y POR2X1_408/Y 0.52fF
C32276 PAND2X1_94/A PAND2X1_49/CTRL2 0.01fF
C32277 POR2X1_283/A POR2X1_90/Y 0.14fF
C32278 POR2X1_356/A POR2X1_317/B 0.07fF
C32279 POR2X1_57/A POR2X1_322/Y 0.00fF
C32280 PAND2X1_56/Y POR2X1_675/Y 0.03fF
C32281 POR2X1_494/a_76_344# PAND2X1_510/B 0.00fF
C32282 POR2X1_65/A POR2X1_761/A 0.03fF
C32283 PAND2X1_213/Y PAND2X1_388/Y 0.06fF
C32284 POR2X1_15/CTRL POR2X1_7/A 0.01fF
C32285 POR2X1_567/A VDD 4.13fF
C32286 POR2X1_57/A PAND2X1_842/Y 0.00fF
C32287 POR2X1_111/O POR2X1_283/A 0.06fF
C32288 PAND2X1_649/A POR2X1_393/CTRL2 0.01fF
C32289 POR2X1_327/Y POR2X1_115/a_16_28# 0.02fF
C32290 POR2X1_523/Y POR2X1_546/O 0.01fF
C32291 POR2X1_266/A POR2X1_786/A 0.01fF
C32292 POR2X1_186/Y POR2X1_736/A 0.46fF
C32293 POR2X1_7/B POR2X1_109/Y 2.11fF
C32294 POR2X1_228/CTRL POR2X1_294/B 0.03fF
C32295 POR2X1_257/A POR2X1_67/Y 0.06fF
C32296 PAND2X1_449/Y PAND2X1_308/Y 0.01fF
C32297 POR2X1_508/B POR2X1_836/Y 0.02fF
C32298 PAND2X1_113/a_76_28# POR2X1_103/Y 0.04fF
C32299 PAND2X1_793/Y POR2X1_171/Y 0.02fF
C32300 PAND2X1_199/A POR2X1_39/B 0.01fF
C32301 POR2X1_542/O VDD 0.00fF
C32302 POR2X1_394/A PAND2X1_566/Y 4.50fF
C32303 POR2X1_7/B POR2X1_397/O 0.00fF
C32304 PAND2X1_63/B POR2X1_7/A 1.68fF
C32305 PAND2X1_191/a_16_344# POR2X1_385/Y 0.07fF
C32306 POR2X1_315/Y PAND2X1_469/Y 0.04fF
C32307 PAND2X1_48/B POR2X1_188/Y 0.03fF
C32308 POR2X1_68/A PAND2X1_394/CTRL2 0.01fF
C32309 POR2X1_727/O POR2X1_854/B 0.09fF
C32310 PAND2X1_39/B POR2X1_287/A 0.64fF
C32311 POR2X1_536/O PAND2X1_222/B 0.01fF
C32312 POR2X1_60/A POR2X1_825/Y 0.03fF
C32313 POR2X1_608/CTRL2 PAND2X1_56/A 0.01fF
C32314 POR2X1_316/Y PAND2X1_254/Y 0.03fF
C32315 POR2X1_1/CTRL POR2X1_260/A 0.09fF
C32316 POR2X1_345/CTRL POR2X1_197/Y 0.01fF
C32317 POR2X1_447/O POR2X1_186/B 0.02fF
C32318 POR2X1_567/A POR2X1_741/Y 0.06fF
C32319 POR2X1_447/B POR2X1_61/B 0.07fF
C32320 POR2X1_13/A POR2X1_387/CTRL2 0.00fF
C32321 PAND2X1_824/B PAND2X1_60/B 0.03fF
C32322 POR2X1_383/A POR2X1_675/Y 0.00fF
C32323 POR2X1_13/A PAND2X1_840/Y 0.00fF
C32324 PAND2X1_158/O POR2X1_260/A 0.10fF
C32325 PAND2X1_158/CTRL POR2X1_156/Y 0.01fF
C32326 POR2X1_647/B POR2X1_649/O 0.03fF
C32327 POR2X1_153/CTRL2 POR2X1_96/B 0.01fF
C32328 PAND2X1_57/B PAND2X1_56/A 0.03fF
C32329 POR2X1_835/B PAND2X1_239/CTRL2 0.03fF
C32330 POR2X1_119/Y POR2X1_232/Y 0.01fF
C32331 POR2X1_471/CTRL2 PAND2X1_72/A 0.03fF
C32332 POR2X1_52/CTRL2 POR2X1_599/A 0.33fF
C32333 POR2X1_193/A POR2X1_632/Y 0.08fF
C32334 POR2X1_579/Y POR2X1_632/Y 0.03fF
C32335 POR2X1_814/A POR2X1_801/B 0.05fF
C32336 PAND2X1_808/B PAND2X1_860/A 0.01fF
C32337 PAND2X1_850/Y POR2X1_184/Y 0.02fF
C32338 POR2X1_132/CTRL2 PAND2X1_140/A 0.01fF
C32339 POR2X1_567/A PAND2X1_32/B 0.05fF
C32340 POR2X1_244/Y POR2X1_141/A 0.08fF
C32341 POR2X1_315/Y POR2X1_394/A 0.03fF
C32342 PAND2X1_323/O PAND2X1_32/B 0.02fF
C32343 POR2X1_66/B PAND2X1_607/O 0.02fF
C32344 POR2X1_54/Y POR2X1_848/Y 0.04fF
C32345 POR2X1_257/A POR2X1_109/CTRL2 0.06fF
C32346 POR2X1_121/CTRL POR2X1_537/Y 0.01fF
C32347 POR2X1_55/CTRL2 POR2X1_624/B 0.01fF
C32348 POR2X1_83/B POR2X1_329/A 0.13fF
C32349 POR2X1_446/B POR2X1_659/A 0.05fF
C32350 POR2X1_257/A PAND2X1_469/a_76_28# 0.01fF
C32351 POR2X1_579/Y PAND2X1_52/B 0.05fF
C32352 POR2X1_416/B PAND2X1_324/Y 0.03fF
C32353 POR2X1_110/Y POR2X1_283/A 0.32fF
C32354 POR2X1_65/A POR2X1_9/Y 7.26fF
C32355 POR2X1_411/B D_INPUT_0 0.74fF
C32356 POR2X1_614/A POR2X1_632/Y 0.06fF
C32357 PAND2X1_634/CTRL2 POR2X1_102/Y 0.00fF
C32358 POR2X1_803/A PAND2X1_72/A 0.03fF
C32359 PAND2X1_717/A POR2X1_72/B 0.15fF
C32360 PAND2X1_65/B POR2X1_846/A 0.03fF
C32361 POR2X1_545/A PAND2X1_52/B 0.03fF
C32362 POR2X1_456/B POR2X1_737/A 0.01fF
C32363 POR2X1_773/B POR2X1_113/B 0.05fF
C32364 PAND2X1_663/O PAND2X1_659/Y 0.04fF
C32365 PAND2X1_339/Y PAND2X1_351/A 0.04fF
C32366 POR2X1_49/Y POR2X1_67/Y 0.03fF
C32367 POR2X1_86/CTRL2 POR2X1_7/A 0.01fF
C32368 POR2X1_227/A POR2X1_227/a_16_28# 0.10fF
C32369 PAND2X1_435/Y POR2X1_411/B 0.10fF
C32370 POR2X1_23/O POR2X1_20/B 0.02fF
C32371 POR2X1_661/A PAND2X1_57/B 0.07fF
C32372 PAND2X1_441/a_16_344# PAND2X1_41/B 0.01fF
C32373 POR2X1_614/A PAND2X1_52/B 0.45fF
C32374 POR2X1_591/Y POR2X1_77/Y 1.26fF
C32375 POR2X1_602/CTRL POR2X1_66/A 0.01fF
C32376 PAND2X1_275/CTRL2 POR2X1_76/B 0.00fF
C32377 POR2X1_860/O POR2X1_861/A 0.02fF
C32378 POR2X1_514/O POR2X1_138/A 0.01fF
C32379 POR2X1_38/B PAND2X1_52/B 0.28fF
C32380 POR2X1_438/m4_208_n4# POR2X1_77/Y 0.12fF
C32381 PAND2X1_12/CTRL2 PAND2X1_11/Y 0.01fF
C32382 POR2X1_416/B PAND2X1_388/Y 0.03fF
C32383 POR2X1_23/Y PAND2X1_477/a_76_28# 0.02fF
C32384 POR2X1_866/A POR2X1_811/m4_208_n4# 0.05fF
C32385 POR2X1_242/CTRL POR2X1_776/A 0.01fF
C32386 PAND2X1_808/O PAND2X1_860/A 0.04fF
C32387 POR2X1_63/Y POR2X1_40/Y 0.15fF
C32388 POR2X1_66/B POR2X1_54/Y 0.06fF
C32389 POR2X1_78/A POR2X1_454/A 0.03fF
C32390 POR2X1_431/a_56_344# POR2X1_236/Y 0.00fF
C32391 PAND2X1_43/CTRL2 POR2X1_852/B 0.03fF
C32392 POR2X1_67/O POR2X1_83/B 0.01fF
C32393 POR2X1_89/CTRL2 POR2X1_60/A 0.01fF
C32394 PAND2X1_65/B POR2X1_705/B 0.03fF
C32395 POR2X1_416/B POR2X1_416/CTRL 0.01fF
C32396 POR2X1_60/A PAND2X1_97/CTRL2 0.01fF
C32397 PAND2X1_422/CTRL PAND2X1_72/A 0.12fF
C32398 POR2X1_287/A POR2X1_325/A 0.06fF
C32399 PAND2X1_449/CTRL VDD -0.00fF
C32400 PAND2X1_241/CTRL2 POR2X1_329/A 0.02fF
C32401 POR2X1_440/Y PAND2X1_52/B 0.03fF
C32402 PAND2X1_388/a_76_28# POR2X1_167/Y 0.01fF
C32403 PAND2X1_358/CTRL2 POR2X1_153/Y 0.30fF
C32404 POR2X1_353/Y POR2X1_443/A 0.14fF
C32405 PAND2X1_298/a_16_344# POR2X1_736/A 0.06fF
C32406 POR2X1_627/CTRL2 POR2X1_628/Y 0.00fF
C32407 POR2X1_67/A POR2X1_29/A 0.09fF
C32408 POR2X1_333/A POR2X1_220/B 0.51fF
C32409 POR2X1_84/A PAND2X1_41/B 0.03fF
C32410 POR2X1_150/Y PAND2X1_592/CTRL 0.00fF
C32411 POR2X1_664/O PAND2X1_72/A 0.01fF
C32412 PAND2X1_472/m4_208_n4# POR2X1_39/B 0.03fF
C32413 POR2X1_271/Y D_INPUT_0 0.03fF
C32414 POR2X1_23/Y POR2X1_423/Y 0.12fF
C32415 PAND2X1_645/CTRL2 POR2X1_600/Y 0.01fF
C32416 PAND2X1_793/Y POR2X1_150/Y 0.03fF
C32417 POR2X1_62/Y POR2X1_39/B 0.74fF
C32418 POR2X1_603/CTRL2 POR2X1_597/A 0.00fF
C32419 PAND2X1_623/a_76_28# POR2X1_669/B 0.10fF
C32420 POR2X1_438/Y PAND2X1_714/A 0.07fF
C32421 PAND2X1_235/O POR2X1_296/B 0.03fF
C32422 POR2X1_669/B PAND2X1_195/CTRL 0.01fF
C32423 POR2X1_142/a_16_28# POR2X1_669/B 0.07fF
C32424 POR2X1_427/O POR2X1_40/Y 0.02fF
C32425 PAND2X1_216/B POR2X1_589/Y 0.00fF
C32426 PAND2X1_34/O POR2X1_27/Y 0.02fF
C32427 POR2X1_862/A POR2X1_480/A 0.55fF
C32428 PAND2X1_201/O POR2X1_55/Y 0.02fF
C32429 PAND2X1_72/A POR2X1_317/B 0.26fF
C32430 POR2X1_54/Y POR2X1_859/A 0.07fF
C32431 POR2X1_327/Y PAND2X1_72/A 2.84fF
C32432 POR2X1_486/O PAND2X1_69/A 0.07fF
C32433 POR2X1_78/B POR2X1_866/A 0.05fF
C32434 PAND2X1_463/CTRL2 PAND2X1_58/A 0.03fF
C32435 POR2X1_502/A D_INPUT_5 0.30fF
C32436 POR2X1_329/A POR2X1_522/Y 0.08fF
C32437 POR2X1_502/A PAND2X1_601/CTRL2 0.01fF
C32438 PAND2X1_206/B PAND2X1_69/A 0.03fF
C32439 POR2X1_376/B D_INPUT_0 0.04fF
C32440 PAND2X1_859/A POR2X1_32/A 0.00fF
C32441 POR2X1_78/B POR2X1_195/A 0.00fF
C32442 POR2X1_121/B POR2X1_405/CTRL 0.01fF
C32443 PAND2X1_9/Y POR2X1_294/B 0.09fF
C32444 PAND2X1_200/CTRL2 POR2X1_72/B 0.03fF
C32445 PAND2X1_206/B PAND2X1_341/A 0.00fF
C32446 POR2X1_864/A PAND2X1_744/CTRL 0.00fF
C32447 POR2X1_609/Y POR2X1_5/Y 0.03fF
C32448 POR2X1_342/a_16_28# POR2X1_342/A 0.03fF
C32449 POR2X1_474/CTRL2 POR2X1_777/B 0.13fF
C32450 POR2X1_661/CTRL POR2X1_661/Y 0.01fF
C32451 POR2X1_847/B POR2X1_669/B 0.05fF
C32452 POR2X1_556/A POR2X1_391/Y 0.02fF
C32453 POR2X1_78/A POR2X1_264/a_16_28# 0.03fF
C32454 POR2X1_446/B POR2X1_276/CTRL 0.01fF
C32455 PAND2X1_850/Y PAND2X1_858/B 0.11fF
C32456 POR2X1_624/Y POR2X1_740/Y 0.10fF
C32457 POR2X1_348/CTRL POR2X1_814/A 0.06fF
C32458 POR2X1_20/B POR2X1_234/O 0.03fF
C32459 POR2X1_650/A POR2X1_267/A 0.01fF
C32460 INPUT_3 PAND2X1_19/CTRL 0.01fF
C32461 PAND2X1_218/B PAND2X1_364/B 0.03fF
C32462 POR2X1_78/A POR2X1_476/Y 0.03fF
C32463 POR2X1_37/Y PAND2X1_673/Y 0.06fF
C32464 PAND2X1_80/CTRL2 PAND2X1_73/Y 0.03fF
C32465 POR2X1_360/A PAND2X1_93/B 0.05fF
C32466 POR2X1_311/Y POR2X1_106/Y 0.03fF
C32467 POR2X1_477/B POR2X1_186/Y 0.05fF
C32468 PAND2X1_20/A POR2X1_489/a_76_344# 0.01fF
C32469 POR2X1_417/Y PAND2X1_211/A 0.23fF
C32470 POR2X1_263/Y POR2X1_230/Y 0.01fF
C32471 POR2X1_122/Y POR2X1_102/Y 0.10fF
C32472 D_INPUT_0 PAND2X1_598/O 0.02fF
C32473 POR2X1_409/B POR2X1_46/Y 2.79fF
C32474 POR2X1_41/B PAND2X1_804/O 0.05fF
C32475 POR2X1_442/Y POR2X1_236/Y 0.01fF
C32476 POR2X1_174/B POR2X1_852/a_56_344# 0.01fF
C32477 POR2X1_499/A POR2X1_318/A 0.07fF
C32478 PAND2X1_721/B VDD 0.18fF
C32479 POR2X1_52/A D_INPUT_0 0.03fF
C32480 POR2X1_383/A PAND2X1_256/CTRL 0.07fF
C32481 POR2X1_311/Y PAND2X1_580/B 0.03fF
C32482 POR2X1_96/A POR2X1_32/A 0.15fF
C32483 POR2X1_65/Y PAND2X1_341/A 0.12fF
C32484 POR2X1_106/CTRL2 PAND2X1_553/B 0.05fF
C32485 POR2X1_413/A POR2X1_48/A 0.04fF
C32486 POR2X1_142/CTRL2 PAND2X1_738/Y 0.08fF
C32487 POR2X1_445/A POR2X1_702/A 0.00fF
C32488 POR2X1_669/B POR2X1_669/CTRL 0.01fF
C32489 PAND2X1_136/O POR2X1_138/A 0.02fF
C32490 PAND2X1_279/CTRL PAND2X1_57/B 0.01fF
C32491 POR2X1_643/A VDD 0.11fF
C32492 POR2X1_800/O VDD 0.00fF
C32493 POR2X1_290/CTRL2 POR2X1_236/Y 0.01fF
C32494 PAND2X1_11/Y INPUT_5 0.08fF
C32495 PAND2X1_139/B POR2X1_40/Y 0.05fF
C32496 POR2X1_529/CTRL2 POR2X1_29/A 0.02fF
C32497 PAND2X1_793/Y PAND2X1_794/O 0.02fF
C32498 PAND2X1_90/A PAND2X1_73/Y 0.24fF
C32499 POR2X1_441/Y PAND2X1_569/B 0.07fF
C32500 INPUT_2 POR2X1_612/Y 0.02fF
C32501 POR2X1_805/B PAND2X1_90/Y 0.18fF
C32502 POR2X1_196/CTRL POR2X1_814/A 0.07fF
C32503 PAND2X1_23/Y POR2X1_296/B 1.45fF
C32504 POR2X1_626/CTRL PAND2X1_6/A 0.03fF
C32505 POR2X1_76/A POR2X1_318/A -0.02fF
C32506 PAND2X1_235/CTRL2 PAND2X1_55/Y 0.03fF
C32507 POR2X1_96/A POR2X1_417/Y 0.03fF
C32508 PAND2X1_833/CTRL2 POR2X1_511/Y 0.03fF
C32509 POR2X1_96/A POR2X1_419/Y 0.00fF
C32510 POR2X1_566/A POR2X1_355/A 0.05fF
C32511 POR2X1_226/Y VDD 0.01fF
C32512 POR2X1_475/O POR2X1_101/Y 0.03fF
C32513 POR2X1_149/B PAND2X1_603/O 0.04fF
C32514 POR2X1_96/A POR2X1_829/a_16_28# 0.03fF
C32515 POR2X1_807/A VDD 0.54fF
C32516 POR2X1_41/B POR2X1_72/B 4.70fF
C32517 POR2X1_41/B PAND2X1_614/CTRL 0.03fF
C32518 PAND2X1_755/a_16_344# PAND2X1_41/B 0.01fF
C32519 POR2X1_847/A PAND2X1_623/Y 0.02fF
C32520 POR2X1_78/B POR2X1_207/A 0.01fF
C32521 POR2X1_278/Y PAND2X1_740/CTRL2 0.05fF
C32522 PAND2X1_843/a_16_344# PAND2X1_738/Y 0.04fF
C32523 POR2X1_590/A PAND2X1_536/O 0.02fF
C32524 POR2X1_121/B PAND2X1_536/CTRL 0.10fF
C32525 POR2X1_65/A POR2X1_278/Y 12.61fF
C32526 POR2X1_66/A PAND2X1_311/CTRL 0.01fF
C32527 PAND2X1_6/Y POR2X1_590/A 0.11fF
C32528 PAND2X1_242/O POR2X1_60/A 0.05fF
C32529 POR2X1_83/A POR2X1_14/Y 0.03fF
C32530 POR2X1_16/A PAND2X1_838/B 0.03fF
C32531 POR2X1_52/A PAND2X1_455/O 0.01fF
C32532 POR2X1_832/A PAND2X1_591/CTRL2 0.03fF
C32533 POR2X1_65/A POR2X1_829/A 0.03fF
C32534 POR2X1_624/Y PAND2X1_133/a_16_344# 0.05fF
C32535 POR2X1_647/m4_208_n4# PAND2X1_60/B 0.12fF
C32536 POR2X1_440/Y POR2X1_434/O 0.01fF
C32537 POR2X1_509/B POR2X1_340/CTRL 0.01fF
C32538 PAND2X1_531/O D_INPUT_1 0.03fF
C32539 PAND2X1_472/A POR2X1_60/A 0.46fF
C32540 PAND2X1_352/A POR2X1_142/Y 0.03fF
C32541 PAND2X1_96/B POR2X1_241/B 0.03fF
C32542 PAND2X1_804/CTRL2 POR2X1_283/A 0.01fF
C32543 PAND2X1_222/A PAND2X1_537/O 0.00fF
C32544 POR2X1_14/Y POR2X1_90/Y 0.07fF
C32545 PAND2X1_282/a_76_28# POR2X1_532/A 0.03fF
C32546 PAND2X1_725/Y PAND2X1_162/O 0.00fF
C32547 POR2X1_198/CTRL2 POR2X1_61/Y 0.01fF
C32548 POR2X1_32/A POR2X1_689/Y 0.00fF
C32549 POR2X1_614/A POR2X1_467/Y 0.03fF
C32550 POR2X1_69/CTRL2 PAND2X1_69/A 0.01fF
C32551 PAND2X1_732/CTRL2 POR2X1_152/Y 0.02fF
C32552 POR2X1_272/Y POR2X1_46/Y 0.05fF
C32553 PAND2X1_453/A POR2X1_90/Y 0.06fF
C32554 POR2X1_523/Y POR2X1_750/B 0.03fF
C32555 POR2X1_43/B POR2X1_60/Y 0.03fF
C32556 PAND2X1_626/O PAND2X1_69/A 0.15fF
C32557 D_INPUT_0 POR2X1_550/Y 1.33fF
C32558 PAND2X1_363/Y POR2X1_42/Y 0.05fF
C32559 POR2X1_57/A POR2X1_83/B 0.22fF
C32560 PAND2X1_386/Y VDD 0.23fF
C32561 POR2X1_13/A PAND2X1_734/B 0.24fF
C32562 PAND2X1_9/a_16_344# D_INPUT_1 0.02fF
C32563 PAND2X1_453/a_76_28# POR2X1_376/B 0.02fF
C32564 POR2X1_675/CTRL POR2X1_540/A 0.06fF
C32565 PAND2X1_486/CTRL VDD 0.00fF
C32566 PAND2X1_115/Y VDD 0.05fF
C32567 POR2X1_646/Y POR2X1_777/Y 0.01fF
C32568 POR2X1_628/Y PAND2X1_156/A 0.05fF
C32569 PAND2X1_467/Y POR2X1_695/Y 0.02fF
C32570 POR2X1_32/A POR2X1_7/A 0.10fF
C32571 POR2X1_76/A POR2X1_574/Y 0.03fF
C32572 POR2X1_750/B PAND2X1_69/A 2.26fF
C32573 POR2X1_102/Y POR2X1_755/Y 0.06fF
C32574 POR2X1_267/A PAND2X1_111/B 0.04fF
C32575 POR2X1_96/A PAND2X1_35/Y 0.03fF
C32576 POR2X1_329/A PAND2X1_841/Y 0.01fF
C32577 POR2X1_106/a_16_28# POR2X1_387/Y 0.04fF
C32578 PAND2X1_724/O PAND2X1_169/Y 0.15fF
C32579 POR2X1_565/B VDD 0.23fF
C32580 POR2X1_546/B VDD 0.03fF
C32581 POR2X1_54/O POR2X1_54/Y 0.05fF
C32582 POR2X1_541/B POR2X1_4/Y 0.01fF
C32583 POR2X1_402/A PAND2X1_395/O 0.03fF
C32584 POR2X1_834/Y PAND2X1_591/O 0.04fF
C32585 POR2X1_693/Y POR2X1_697/CTRL 0.01fF
C32586 PAND2X1_387/a_16_344# POR2X1_712/Y 0.00fF
C32587 POR2X1_311/Y PAND2X1_349/A 0.00fF
C32588 POR2X1_94/A PAND2X1_521/CTRL2 0.05fF
C32589 PAND2X1_94/A POR2X1_496/Y 0.05fF
C32590 POR2X1_415/Y VDD 0.12fF
C32591 PAND2X1_20/CTRL POR2X1_68/B 0.01fF
C32592 PAND2X1_172/CTRL2 POR2X1_174/A 0.01fF
C32593 POR2X1_118/Y PAND2X1_560/B 0.03fF
C32594 PAND2X1_613/CTRL2 POR2X1_620/B 0.14fF
C32595 POR2X1_62/Y PAND2X1_613/O 0.15fF
C32596 PAND2X1_27/O POR2X1_294/A 0.17fF
C32597 POR2X1_174/CTRL2 POR2X1_174/A 0.01fF
C32598 PAND2X1_818/O POR2X1_42/Y 0.04fF
C32599 PAND2X1_319/B POR2X1_312/Y 0.10fF
C32600 POR2X1_60/A POR2X1_527/Y 0.09fF
C32601 POR2X1_65/A POR2X1_761/Y 0.04fF
C32602 POR2X1_134/Y PAND2X1_768/Y 0.01fF
C32603 PAND2X1_429/CTRL POR2X1_260/A 0.01fF
C32604 POR2X1_140/B VDD 0.04fF
C32605 POR2X1_738/Y POR2X1_740/Y 0.00fF
C32606 POR2X1_417/Y POR2X1_7/A -0.01fF
C32607 POR2X1_419/Y POR2X1_7/A 0.15fF
C32608 POR2X1_237/CTRL POR2X1_90/Y 0.01fF
C32609 POR2X1_407/A VDD 0.91fF
C32610 POR2X1_130/A PAND2X1_767/CTRL2 0.02fF
C32611 POR2X1_96/A POR2X1_189/Y 0.01fF
C32612 POR2X1_297/Y PAND2X1_566/Y 0.05fF
C32613 POR2X1_334/Y POR2X1_856/B 0.10fF
C32614 POR2X1_866/A POR2X1_294/A 0.10fF
C32615 POR2X1_383/A POR2X1_405/CTRL 0.05fF
C32616 POR2X1_57/A PAND2X1_319/CTRL2 0.03fF
C32617 POR2X1_240/B POR2X1_260/A 0.01fF
C32618 POR2X1_56/Y VDD 0.67fF
C32619 PAND2X1_725/A PAND2X1_707/O 0.00fF
C32620 PAND2X1_349/A PAND2X1_140/CTRL2 0.01fF
C32621 PAND2X1_81/B POR2X1_786/a_16_28# 0.00fF
C32622 POR2X1_66/A PAND2X1_384/CTRL 0.01fF
C32623 POR2X1_355/B POR2X1_795/B 0.03fF
C32624 POR2X1_195/A POR2X1_294/A 0.00fF
C32625 INPUT_6 INPUT_7 12.29fF
C32626 POR2X1_325/O POR2X1_750/B 0.01fF
C32627 PAND2X1_771/Y PAND2X1_345/Y 0.23fF
C32628 POR2X1_122/Y POR2X1_821/Y 0.03fF
C32629 POR2X1_701/Y PAND2X1_711/A 0.02fF
C32630 POR2X1_62/Y POR2X1_48/A 0.03fF
C32631 POR2X1_96/A POR2X1_184/Y 0.03fF
C32632 POR2X1_128/a_16_28# PAND2X1_55/Y 0.03fF
C32633 POR2X1_62/Y POR2X1_623/O 0.26fF
C32634 PAND2X1_20/A PAND2X1_503/O 0.15fF
C32635 POR2X1_496/Y PAND2X1_507/O 0.08fF
C32636 PAND2X1_859/A POR2X1_503/Y 0.02fF
C32637 POR2X1_389/Y POR2X1_537/A 0.01fF
C32638 PAND2X1_23/Y POR2X1_363/CTRL2 0.01fF
C32639 PAND2X1_267/O POR2X1_7/Y 0.02fF
C32640 PAND2X1_496/O POR2X1_575/B 0.03fF
C32641 POR2X1_405/a_16_28# PAND2X1_60/B 0.02fF
C32642 PAND2X1_55/Y POR2X1_832/B 0.03fF
C32643 POR2X1_66/B PAND2X1_748/O 0.05fF
C32644 PAND2X1_289/O POR2X1_568/B 0.03fF
C32645 POR2X1_675/O POR2X1_456/B 0.16fF
C32646 POR2X1_258/O VDD 0.00fF
C32647 POR2X1_57/A PAND2X1_140/Y 0.03fF
C32648 POR2X1_99/B PAND2X1_93/B 0.03fF
C32649 INPUT_1 POR2X1_482/Y 0.03fF
C32650 POR2X1_96/A PAND2X1_651/Y 0.08fF
C32651 POR2X1_383/A POR2X1_637/B 0.00fF
C32652 POR2X1_278/Y PAND2X1_359/B 0.01fF
C32653 POR2X1_83/A POR2X1_55/Y 1.13fF
C32654 POR2X1_198/CTRL2 POR2X1_35/Y 0.01fF
C32655 INPUT_0 PAND2X1_548/a_76_28# 0.04fF
C32656 PAND2X1_823/CTRL PAND2X1_41/B 0.03fF
C32657 PAND2X1_572/CTRL INPUT_0 0.03fF
C32658 POR2X1_137/O POR2X1_391/Y 0.03fF
C32659 POR2X1_809/A POR2X1_296/B 0.03fF
C32660 POR2X1_68/A POR2X1_198/B 0.34fF
C32661 PAND2X1_787/A PAND2X1_556/B 0.11fF
C32662 PAND2X1_803/Y VDD 0.73fF
C32663 PAND2X1_48/B POR2X1_731/CTRL2 0.01fF
C32664 PAND2X1_243/a_16_344# PAND2X1_734/B 0.03fF
C32665 PAND2X1_741/B POR2X1_7/A 0.09fF
C32666 PAND2X1_700/O PAND2X1_60/B 0.01fF
C32667 POR2X1_102/Y PAND2X1_508/Y 0.03fF
C32668 POR2X1_72/B PAND2X1_308/Y 0.03fF
C32669 POR2X1_482/Y POR2X1_153/Y 0.05fF
C32670 PAND2X1_65/B POR2X1_352/CTRL2 0.01fF
C32671 PAND2X1_824/B POR2X1_750/B 0.10fF
C32672 POR2X1_140/B POR2X1_741/Y 0.03fF
C32673 PAND2X1_512/Y PAND2X1_549/B 3.03fF
C32674 POR2X1_55/Y POR2X1_90/Y 0.29fF
C32675 POR2X1_78/A POR2X1_571/Y 0.03fF
C32676 POR2X1_483/B POR2X1_510/Y 0.06fF
C32677 INPUT_6 INPUT_4 0.13fF
C32678 PAND2X1_651/Y PAND2X1_506/CTRL 0.00fF
C32679 POR2X1_93/A POR2X1_618/CTRL 0.01fF
C32680 POR2X1_391/CTRL2 POR2X1_546/A 0.01fF
C32681 POR2X1_72/B PAND2X1_861/a_76_28# 0.01fF
C32682 POR2X1_324/CTRL2 POR2X1_324/A 0.01fF
C32683 PAND2X1_558/Y POR2X1_394/A 0.29fF
C32684 POR2X1_283/A INPUT_0 0.07fF
C32685 PAND2X1_469/Y PAND2X1_480/B 0.03fF
C32686 POR2X1_110/Y POR2X1_14/Y 0.06fF
C32687 POR2X1_99/B POR2X1_78/A 0.01fF
C32688 POR2X1_78/B POR2X1_596/CTRL2 0.03fF
C32689 POR2X1_222/Y POR2X1_556/Y 0.03fF
C32690 PAND2X1_436/A PAND2X1_508/Y 0.39fF
C32691 PAND2X1_661/Y POR2X1_13/A 0.01fF
C32692 POR2X1_355/B POR2X1_383/A 0.03fF
C32693 POR2X1_78/B POR2X1_703/A 0.07fF
C32694 POR2X1_579/Y POR2X1_350/B 0.03fF
C32695 PAND2X1_41/B POR2X1_227/CTRL 0.00fF
C32696 POR2X1_508/B POR2X1_836/A 0.00fF
C32697 POR2X1_602/B PAND2X1_48/A 0.03fF
C32698 POR2X1_518/CTRL2 POR2X1_667/A 0.01fF
C32699 PAND2X1_370/O PAND2X1_566/Y 0.00fF
C32700 POR2X1_557/A PAND2X1_8/Y 0.02fF
C32701 PAND2X1_727/CTRL VDD -0.00fF
C32702 POR2X1_68/A POR2X1_685/B 0.02fF
C32703 POR2X1_407/A PAND2X1_32/B 0.10fF
C32704 PAND2X1_356/B PAND2X1_354/Y 0.05fF
C32705 PAND2X1_744/a_16_344# POR2X1_644/A 0.02fF
C32706 POR2X1_809/A PAND2X1_679/CTRL2 0.01fF
C32707 PAND2X1_48/B POR2X1_510/Y 0.03fF
C32708 POR2X1_242/CTRL POR2X1_191/Y 0.13fF
C32709 POR2X1_38/Y POR2X1_406/A 0.01fF
C32710 POR2X1_751/CTRL2 POR2X1_816/A 0.01fF
C32711 POR2X1_119/Y PAND2X1_786/a_56_28# 0.00fF
C32712 PAND2X1_6/A POR2X1_619/Y 0.00fF
C32713 PAND2X1_631/CTRL POR2X1_93/A 0.00fF
C32714 POR2X1_532/A POR2X1_710/O 0.15fF
C32715 POR2X1_596/A PAND2X1_743/CTRL 0.01fF
C32716 POR2X1_63/CTRL POR2X1_7/A 0.01fF
C32717 PAND2X1_449/Y PAND2X1_241/Y 0.03fF
C32718 POR2X1_855/B PAND2X1_599/O 0.02fF
C32719 PAND2X1_23/Y POR2X1_507/CTRL 0.01fF
C32720 POR2X1_270/Y POR2X1_717/B 0.02fF
C32721 PAND2X1_60/B POR2X1_723/B 0.03fF
C32722 POR2X1_296/B POR2X1_711/Y 0.10fF
C32723 PAND2X1_645/B POR2X1_73/Y 0.21fF
C32724 POR2X1_112/Y POR2X1_724/A 0.17fF
C32725 PAND2X1_635/Y POR2X1_20/B 0.03fF
C32726 POR2X1_853/A POR2X1_566/B 0.08fF
C32727 PAND2X1_48/B POR2X1_276/Y 0.95fF
C32728 PAND2X1_480/B POR2X1_394/A 0.14fF
C32729 POR2X1_611/O POR2X1_4/Y 0.01fF
C32730 PAND2X1_716/O PAND2X1_656/A 0.02fF
C32731 POR2X1_337/A POR2X1_337/a_16_28# 0.04fF
C32732 POR2X1_673/Y POR2X1_546/B 1.31fF
C32733 PAND2X1_55/Y POR2X1_151/O 0.16fF
C32734 POR2X1_110/Y POR2X1_237/CTRL 0.02fF
C32735 PAND2X1_651/Y POR2X1_7/A 0.18fF
C32736 POR2X1_346/CTRL2 PAND2X1_60/B 0.01fF
C32737 PAND2X1_48/B POR2X1_543/O 0.01fF
C32738 POR2X1_824/CTRL2 VDD 0.00fF
C32739 PAND2X1_598/a_56_28# POR2X1_394/A 0.00fF
C32740 POR2X1_814/A POR2X1_705/B 0.03fF
C32741 POR2X1_590/A PAND2X1_52/B 1.08fF
C32742 PAND2X1_465/CTRL2 POR2X1_77/Y 0.01fF
C32743 PAND2X1_329/O PAND2X1_69/A 0.03fF
C32744 POR2X1_7/B PAND2X1_337/CTRL2 0.00fF
C32745 POR2X1_97/A POR2X1_568/A 9.31fF
C32746 POR2X1_164/Y PAND2X1_565/CTRL 0.01fF
C32747 POR2X1_94/A PAND2X1_102/O 0.05fF
C32748 POR2X1_800/A POR2X1_260/A 0.00fF
C32749 PAND2X1_57/B POR2X1_737/A 0.03fF
C32750 PAND2X1_649/A POR2X1_689/CTRL 0.01fF
C32751 POR2X1_52/A PAND2X1_162/A 0.01fF
C32752 PAND2X1_659/Y PAND2X1_659/O 0.02fF
C32753 POR2X1_131/a_56_344# PAND2X1_349/A 0.00fF
C32754 POR2X1_383/A POR2X1_791/B 0.05fF
C32755 POR2X1_123/A POR2X1_68/B 0.03fF
C32756 POR2X1_218/A POR2X1_218/a_16_28# 0.03fF
C32757 PAND2X1_90/A POR2X1_576/a_16_28# 0.03fF
C32758 PAND2X1_659/Y POR2X1_498/CTRL2 0.00fF
C32759 POR2X1_41/B POR2X1_595/CTRL 0.03fF
C32760 POR2X1_38/Y PAND2X1_63/B 0.03fF
C32761 POR2X1_112/CTRL2 POR2X1_332/B 0.01fF
C32762 POR2X1_326/A POR2X1_652/Y 0.03fF
C32763 POR2X1_558/Y POR2X1_294/B 0.04fF
C32764 POR2X1_72/B POR2X1_77/Y 0.97fF
C32765 PAND2X1_117/O POR2X1_557/B 0.03fF
C32766 POR2X1_20/B POR2X1_667/a_16_28# 0.00fF
C32767 POR2X1_79/Y POR2X1_385/Y 0.05fF
C32768 POR2X1_740/Y POR2X1_186/B 0.05fF
C32769 POR2X1_836/B POR2X1_568/A 0.01fF
C32770 PAND2X1_313/a_76_28# POR2X1_732/B 0.05fF
C32771 PAND2X1_737/B POR2X1_73/Y 0.03fF
C32772 POR2X1_702/A POR2X1_260/A 0.00fF
C32773 POR2X1_416/B PAND2X1_742/a_76_28# 0.02fF
C32774 PAND2X1_55/Y PAND2X1_527/CTRL 0.02fF
C32775 PAND2X1_798/B PAND2X1_853/B 0.03fF
C32776 POR2X1_383/A POR2X1_510/B 0.03fF
C32777 POR2X1_319/Y POR2X1_854/B 0.74fF
C32778 POR2X1_62/Y PAND2X1_197/Y 0.01fF
C32779 PAND2X1_679/CTRL2 POR2X1_728/A 0.00fF
C32780 POR2X1_388/a_16_28# POR2X1_703/A 0.04fF
C32781 PAND2X1_26/O POR2X1_260/A 0.00fF
C32782 POR2X1_20/a_56_344# POR2X1_4/Y 0.01fF
C32783 POR2X1_3/a_76_344# POR2X1_260/A 0.00fF
C32784 POR2X1_260/A PAND2X1_670/CTRL 0.01fF
C32785 PAND2X1_716/CTRL2 PAND2X1_716/B 0.01fF
C32786 PAND2X1_48/A POR2X1_712/Y 0.12fF
C32787 INPUT_6 PAND2X1_157/CTRL 0.01fF
C32788 PAND2X1_341/A PAND2X1_560/B 0.07fF
C32789 PAND2X1_549/O POR2X1_39/B 0.17fF
C32790 INPUT_1 PAND2X1_63/B 0.05fF
C32791 POR2X1_680/a_16_28# POR2X1_79/Y 0.03fF
C32792 PAND2X1_860/A PAND2X1_795/CTRL 0.01fF
C32793 POR2X1_854/CTRL POR2X1_776/A 0.01fF
C32794 POR2X1_610/m4_208_n4# POR2X1_814/A 0.12fF
C32795 PAND2X1_48/A POR2X1_500/Y 0.03fF
C32796 PAND2X1_20/A POR2X1_837/B 0.00fF
C32797 POR2X1_177/Y POR2X1_167/Y 0.01fF
C32798 POR2X1_57/A PAND2X1_325/CTRL 0.01fF
C32799 PAND2X1_490/CTRL POR2X1_4/Y 0.06fF
C32800 PAND2X1_404/Y POR2X1_20/B 0.08fF
C32801 PAND2X1_349/A POR2X1_153/Y 0.07fF
C32802 POR2X1_424/a_16_28# POR2X1_77/Y 0.09fF
C32803 POR2X1_20/B POR2X1_616/CTRL2 0.03fF
C32804 POR2X1_150/Y POR2X1_437/a_16_28# 0.01fF
C32805 PAND2X1_69/A PAND2X1_122/CTRL 0.01fF
C32806 PAND2X1_634/O POR2X1_48/A 0.01fF
C32807 POR2X1_489/B POR2X1_814/A 0.00fF
C32808 PAND2X1_253/CTRL POR2X1_186/B 0.02fF
C32809 POR2X1_760/A POR2X1_32/A 0.03fF
C32810 POR2X1_857/B PAND2X1_52/B 5.21fF
C32811 PAND2X1_175/a_16_344# PAND2X1_853/B 0.01fF
C32812 PAND2X1_409/a_16_344# PAND2X1_52/B 0.04fF
C32813 POR2X1_754/A POR2X1_90/CTRL2 0.00fF
C32814 POR2X1_681/O POR2X1_60/A 0.01fF
C32815 POR2X1_854/O POR2X1_567/B 0.03fF
C32816 POR2X1_366/Y POR2X1_568/A 0.07fF
C32817 POR2X1_52/A POR2X1_90/O 0.11fF
C32818 POR2X1_334/Y POR2X1_244/Y 0.64fF
C32819 POR2X1_335/A PAND2X1_72/A 0.12fF
C32820 PAND2X1_835/Y POR2X1_77/Y 0.01fF
C32821 POR2X1_43/B PAND2X1_351/A 0.04fF
C32822 PAND2X1_639/Y PAND2X1_651/A -0.00fF
C32823 PAND2X1_552/B POR2X1_167/Y 0.18fF
C32824 POR2X1_41/B PAND2X1_147/CTRL 0.05fF
C32825 POR2X1_287/B POR2X1_486/CTRL 0.01fF
C32826 POR2X1_152/Y POR2X1_39/B 0.05fF
C32827 POR2X1_716/a_16_28# POR2X1_723/B 0.02fF
C32828 POR2X1_257/A POR2X1_432/O 0.09fF
C32829 POR2X1_66/B POR2X1_78/Y 0.00fF
C32830 POR2X1_153/a_16_28# POR2X1_394/A 0.05fF
C32831 POR2X1_502/A PAND2X1_438/CTRL 0.01fF
C32832 POR2X1_78/A POR2X1_266/CTRL2 0.03fF
C32833 PAND2X1_601/CTRL POR2X1_296/B 0.02fF
C32834 PAND2X1_39/B POR2X1_806/CTRL 0.01fF
C32835 POR2X1_102/Y PAND2X1_791/O 0.05fF
C32836 POR2X1_327/Y POR2X1_537/Y 0.06fF
C32837 POR2X1_411/B POR2X1_609/O 0.02fF
C32838 POR2X1_825/Y POR2X1_396/CTRL2 0.00fF
C32839 POR2X1_266/A POR2X1_845/A 0.01fF
C32840 POR2X1_361/CTRL2 PAND2X1_72/A 0.01fF
C32841 POR2X1_760/A PAND2X1_741/B 0.07fF
C32842 POR2X1_188/A POR2X1_841/a_56_344# 0.00fF
C32843 PAND2X1_780/CTRL2 VDD 0.00fF
C32844 PAND2X1_66/a_76_28# POR2X1_67/A 0.04fF
C32845 PAND2X1_97/Y VDD 0.21fF
C32846 D_INPUT_5 PAND2X1_425/CTRL 0.01fF
C32847 PAND2X1_730/A POR2X1_385/Y 0.05fF
C32848 PAND2X1_222/A POR2X1_40/Y 0.01fF
C32849 POR2X1_634/A POR2X1_260/B 0.02fF
C32850 POR2X1_519/O POR2X1_416/B 0.01fF
C32851 PAND2X1_717/A POR2X1_7/B 0.05fF
C32852 POR2X1_327/Y POR2X1_532/O 0.02fF
C32853 POR2X1_153/Y PAND2X1_860/a_76_28# 0.03fF
C32854 POR2X1_760/A PAND2X1_35/Y 0.07fF
C32855 POR2X1_614/A PAND2X1_255/CTRL2 0.05fF
C32856 POR2X1_482/CTRL POR2X1_60/A 0.01fF
C32857 POR2X1_101/Y POR2X1_717/B 0.01fF
C32858 POR2X1_675/CTRL2 POR2X1_466/A 0.14fF
C32859 POR2X1_191/Y POR2X1_551/A 0.03fF
C32860 POR2X1_614/Y POR2X1_29/A 0.05fF
C32861 POR2X1_656/m4_208_n4# D_INPUT_0 0.07fF
C32862 POR2X1_337/Y PAND2X1_167/O 0.30fF
C32863 POR2X1_805/Y POR2X1_792/O 0.02fF
C32864 PAND2X1_435/O POR2X1_271/B 0.01fF
C32865 POR2X1_411/B PAND2X1_735/Y 0.07fF
C32866 PAND2X1_73/Y PAND2X1_531/a_16_344# 0.04fF
C32867 POR2X1_777/B POR2X1_458/a_76_344# 0.03fF
C32868 POR2X1_609/Y POR2X1_607/O 0.05fF
C32869 POR2X1_52/A POR2X1_816/O 0.01fF
C32870 PAND2X1_779/O POR2X1_39/B 0.15fF
C32871 POR2X1_257/A PAND2X1_707/CTRL 0.01fF
C32872 POR2X1_41/B PAND2X1_247/CTRL 0.03fF
C32873 PAND2X1_446/O POR2X1_418/Y -0.00fF
C32874 PAND2X1_852/A POR2X1_236/Y 0.01fF
C32875 POR2X1_502/A POR2X1_212/A 0.16fF
C32876 POR2X1_76/A PAND2X1_131/O 0.01fF
C32877 POR2X1_814/B POR2X1_479/B 0.03fF
C32878 POR2X1_130/A POR2X1_260/B 0.18fF
C32879 POR2X1_411/B PAND2X1_218/CTRL2 0.01fF
C32880 POR2X1_670/Y POR2X1_20/B 0.01fF
C32881 PAND2X1_496/a_76_28# D_INPUT_1 0.02fF
C32882 POR2X1_360/A PAND2X1_82/a_16_344# 0.02fF
C32883 POR2X1_48/A POR2X1_393/CTRL2 0.00fF
C32884 POR2X1_808/B VDD 0.08fF
C32885 PAND2X1_771/Y VDD 2.89fF
C32886 POR2X1_666/Y PAND2X1_719/Y 0.02fF
C32887 POR2X1_66/B PAND2X1_13/CTRL2 0.03fF
C32888 PAND2X1_206/B PAND2X1_338/B 0.07fF
C32889 POR2X1_633/CTRL POR2X1_68/B 0.00fF
C32890 POR2X1_360/A POR2X1_84/A 11.07fF
C32891 PAND2X1_168/Y POR2X1_40/Y 0.01fF
C32892 POR2X1_729/O POR2X1_452/Y 0.01fF
C32893 POR2X1_20/B PAND2X1_565/A 0.03fF
C32894 POR2X1_528/Y POR2X1_329/A 0.07fF
C32895 POR2X1_855/B POR2X1_814/A 0.05fF
C32896 POR2X1_754/Y VDD 0.16fF
C32897 POR2X1_116/A POR2X1_501/B 0.03fF
C32898 POR2X1_66/B PAND2X1_52/Y 0.03fF
C32899 POR2X1_60/A PAND2X1_803/A 0.03fF
C32900 POR2X1_841/O POR2X1_804/A 0.24fF
C32901 PAND2X1_669/O POR2X1_668/Y 0.02fF
C32902 POR2X1_60/A POR2X1_677/a_16_28# 0.02fF
C32903 PAND2X1_794/CTRL2 PAND2X1_580/B 0.00fF
C32904 PAND2X1_211/A PAND2X1_731/B 0.35fF
C32905 POR2X1_341/A POR2X1_576/Y 0.02fF
C32906 POR2X1_65/A PAND2X1_169/Y 2.23fF
C32907 PAND2X1_93/B POR2X1_664/Y 0.02fF
C32908 PAND2X1_462/B POR2X1_612/Y 0.03fF
C32909 POR2X1_411/O POR2X1_37/Y 0.05fF
C32910 POR2X1_490/Y PAND2X1_716/CTRL2 0.03fF
C32911 PAND2X1_93/B PAND2X1_275/CTRL 0.02fF
C32912 POR2X1_286/Y POR2X1_389/Y 0.03fF
C32913 POR2X1_446/B POR2X1_513/Y 0.03fF
C32914 PAND2X1_11/Y PAND2X1_587/Y 0.10fF
C32915 POR2X1_23/Y PAND2X1_707/Y 0.39fF
C32916 PAND2X1_65/B PAND2X1_766/CTRL 0.01fF
C32917 POR2X1_462/B POR2X1_848/Y 0.01fF
C32918 POR2X1_40/Y POR2X1_743/O 0.01fF
C32919 POR2X1_677/Y PAND2X1_508/Y 0.03fF
C32920 POR2X1_818/Y POR2X1_415/Y 0.03fF
C32921 POR2X1_78/A POR2X1_608/a_16_28# 0.00fF
C32922 POR2X1_14/Y INPUT_0 0.08fF
C32923 POR2X1_669/B POR2X1_754/A 0.05fF
C32924 PAND2X1_827/CTRL POR2X1_741/Y 0.01fF
C32925 PAND2X1_318/a_76_28# PAND2X1_776/Y 0.04fF
C32926 PAND2X1_719/Y VDD 0.13fF
C32927 POR2X1_102/Y PAND2X1_778/a_76_28# 0.01fF
C32928 POR2X1_614/Y PAND2X1_754/O 0.00fF
C32929 PAND2X1_575/B VDD 0.01fF
C32930 POR2X1_60/A PAND2X1_673/Y 1.71fF
C32931 POR2X1_23/Y PAND2X1_798/B 0.03fF
C32932 POR2X1_296/Y PAND2X1_57/B 0.00fF
C32933 POR2X1_813/CTRL2 POR2X1_7/A 0.02fF
C32934 PAND2X1_475/O PAND2X1_474/Y 0.00fF
C32935 PAND2X1_402/CTRL POR2X1_236/Y 0.01fF
C32936 PAND2X1_6/Y POR2X1_851/A 0.00fF
C32937 PAND2X1_206/B PAND2X1_341/Y 0.00fF
C32938 POR2X1_411/B PAND2X1_383/a_16_344# 0.01fF
C32939 PAND2X1_283/CTRL2 POR2X1_66/A 0.01fF
C32940 POR2X1_614/A POR2X1_809/O 0.01fF
C32941 PAND2X1_477/a_76_28# POR2X1_238/Y 0.02fF
C32942 PAND2X1_20/A POR2X1_128/O 0.01fF
C32943 POR2X1_644/O POR2X1_644/A 0.02fF
C32944 PAND2X1_627/CTRL POR2X1_852/B 0.07fF
C32945 POR2X1_538/O POR2X1_66/A 0.18fF
C32946 POR2X1_820/a_16_28# POR2X1_820/B 0.02fF
C32947 POR2X1_752/Y POR2X1_585/a_16_28# 0.03fF
C32948 POR2X1_110/Y PAND2X1_458/O 0.01fF
C32949 PAND2X1_20/A POR2X1_776/B 0.28fF
C32950 POR2X1_78/A POR2X1_664/Y 0.03fF
C32951 POR2X1_60/A PAND2X1_788/m4_208_n4# 0.09fF
C32952 POR2X1_260/B POR2X1_573/A 0.03fF
C32953 PAND2X1_640/O PAND2X1_640/B 0.01fF
C32954 POR2X1_334/B POR2X1_296/B 0.03fF
C32955 POR2X1_502/A POR2X1_330/Y 0.05fF
C32956 POR2X1_300/CTRL2 POR2X1_102/Y 0.01fF
C32957 POR2X1_460/Y PAND2X1_376/O 0.02fF
C32958 POR2X1_257/A POR2X1_765/Y 0.03fF
C32959 PAND2X1_6/Y POR2X1_66/A 0.13fF
C32960 POR2X1_49/Y PAND2X1_473/Y 1.17fF
C32961 POR2X1_390/B POR2X1_556/A 0.03fF
C32962 POR2X1_433/Y POR2X1_432/CTRL2 0.01fF
C32963 POR2X1_302/B PAND2X1_57/B 0.04fF
C32964 POR2X1_78/B PAND2X1_16/a_16_344# 0.02fF
C32965 POR2X1_65/A PAND2X1_730/B 0.03fF
C32966 POR2X1_150/Y PAND2X1_130/a_76_28# 0.02fF
C32967 PAND2X1_433/a_76_28# D_INPUT_0 0.02fF
C32968 POR2X1_446/B POR2X1_366/A 0.03fF
C32969 POR2X1_65/A GATE_741 0.01fF
C32970 POR2X1_775/A POR2X1_78/A 0.08fF
C32971 PAND2X1_6/Y POR2X1_34/A 0.01fF
C32972 POR2X1_407/A POR2X1_660/CTRL2 0.04fF
C32973 POR2X1_56/B POR2X1_40/Y 0.03fF
C32974 POR2X1_634/A PAND2X1_55/Y 0.10fF
C32975 POR2X1_43/B PAND2X1_443/Y 0.04fF
C32976 PAND2X1_679/O POR2X1_676/Y -0.00fF
C32977 POR2X1_43/B POR2X1_497/CTRL2 0.01fF
C32978 POR2X1_71/Y PAND2X1_217/B 0.17fF
C32979 POR2X1_48/A POR2X1_152/Y 1.07fF
C32980 POR2X1_820/O POR2X1_42/Y 0.25fF
C32981 POR2X1_77/Y PAND2X1_147/CTRL 0.00fF
C32982 POR2X1_78/B POR2X1_206/A 0.03fF
C32983 POR2X1_68/A POR2X1_850/B 0.05fF
C32984 PAND2X1_65/B POR2X1_192/Y 0.09fF
C32985 POR2X1_329/m4_208_n4# PAND2X1_557/A 0.07fF
C32986 POR2X1_121/B PAND2X1_743/CTRL2 0.07fF
C32987 POR2X1_356/A POR2X1_856/O 0.04fF
C32988 PAND2X1_742/B POR2X1_72/B 0.03fF
C32989 PAND2X1_482/CTRL2 POR2X1_541/B 0.05fF
C32990 POR2X1_121/B POR2X1_513/Y 0.03fF
C32991 POR2X1_671/O VDD 0.00fF
C32992 POR2X1_618/CTRL2 POR2X1_5/Y 0.01fF
C32993 PAND2X1_217/B POR2X1_42/Y 0.11fF
C32994 POR2X1_356/A POR2X1_781/B 0.04fF
C32995 PAND2X1_208/a_76_28# PAND2X1_198/Y 0.02fF
C32996 POR2X1_814/B POR2X1_791/CTRL 0.01fF
C32997 PAND2X1_23/Y POR2X1_186/Y 0.12fF
C32998 POR2X1_38/Y POR2X1_32/A 0.70fF
C32999 PAND2X1_431/CTRL2 POR2X1_440/Y 0.01fF
C33000 D_INPUT_1 POR2X1_390/O 0.14fF
C33001 PAND2X1_84/Y PAND2X1_795/B 0.03fF
C33002 POR2X1_834/Y POR2X1_648/a_16_28# 0.03fF
C33003 POR2X1_60/A POR2X1_759/A 0.02fF
C33004 POR2X1_49/Y PAND2X1_478/CTRL 0.01fF
C33005 POR2X1_66/B POR2X1_816/A 0.03fF
C33006 POR2X1_73/CTRL2 POR2X1_37/Y 0.00fF
C33007 PAND2X1_859/B POR2X1_376/B 0.01fF
C33008 POR2X1_260/B POR2X1_596/CTRL 0.01fF
C33009 POR2X1_66/B D_INPUT_1 0.03fF
C33010 POR2X1_652/Y POR2X1_480/A 0.00fF
C33011 PAND2X1_96/B PAND2X1_74/CTRL2 0.00fF
C33012 POR2X1_817/A VDD 0.33fF
C33013 POR2X1_102/Y PAND2X1_572/CTRL 0.00fF
C33014 POR2X1_41/B PAND2X1_192/a_76_28# 0.01fF
C33015 PAND2X1_428/CTRL PAND2X1_32/B 0.01fF
C33016 POR2X1_634/A POR2X1_407/Y 0.05fF
C33017 POR2X1_29/A PAND2X1_670/O 0.11fF
C33018 POR2X1_72/B POR2X1_52/Y 0.03fF
C33019 POR2X1_378/CTRL2 D_INPUT_1 0.01fF
C33020 POR2X1_376/B PAND2X1_174/O 0.18fF
C33021 POR2X1_292/O POR2X1_77/Y 0.08fF
C33022 PAND2X1_281/CTRL2 POR2X1_647/B 0.03fF
C33023 POR2X1_71/Y VDD 0.20fF
C33024 POR2X1_51/A POR2X1_96/A 0.01fF
C33025 POR2X1_114/B POR2X1_287/B 0.03fF
C33026 POR2X1_632/B POR2X1_510/Y 1.56fF
C33027 PAND2X1_718/Y POR2X1_591/Y 0.01fF
C33028 POR2X1_137/B PAND2X1_134/CTRL2 0.01fF
C33029 PAND2X1_48/B POR2X1_471/CTRL2 0.01fF
C33030 POR2X1_66/B POR2X1_724/A 0.03fF
C33031 POR2X1_96/Y PAND2X1_201/O 0.04fF
C33032 PAND2X1_39/B PAND2X1_48/A 0.18fF
C33033 PAND2X1_341/CTRL2 INPUT_0 0.05fF
C33034 PAND2X1_69/A POR2X1_389/Y 0.07fF
C33035 PAND2X1_264/CTRL2 POR2X1_669/B 0.02fF
C33036 PAND2X1_656/a_56_28# PAND2X1_656/A 0.00fF
C33037 POR2X1_499/O POR2X1_260/A 0.01fF
C33038 POR2X1_52/A PAND2X1_735/Y 0.00fF
C33039 POR2X1_96/A POR2X1_406/CTRL2 0.03fF
C33040 POR2X1_334/B POR2X1_547/B 0.03fF
C33041 POR2X1_42/Y VDD 5.55fF
C33042 PAND2X1_97/CTRL POR2X1_153/Y 0.09fF
C33043 PAND2X1_832/O PAND2X1_651/Y 0.02fF
C33044 INPUT_0 POR2X1_55/Y 0.22fF
C33045 POR2X1_102/Y POR2X1_283/A 0.06fF
C33046 POR2X1_74/a_76_344# POR2X1_23/Y 0.03fF
C33047 POR2X1_41/B PAND2X1_830/Y 0.03fF
C33048 POR2X1_130/A PAND2X1_55/Y 1.66fF
C33049 PAND2X1_69/A POR2X1_720/A 0.05fF
C33050 PAND2X1_793/A POR2X1_90/Y 0.18fF
C33051 POR2X1_102/Y PAND2X1_121/CTRL 0.01fF
C33052 POR2X1_16/A POR2X1_487/CTRL 0.06fF
C33053 POR2X1_625/CTRL2 POR2X1_90/Y 0.03fF
C33054 PAND2X1_57/B POR2X1_756/CTRL 0.01fF
C33055 POR2X1_41/B POR2X1_7/B 0.18fF
C33056 POR2X1_333/A POR2X1_854/B 0.03fF
C33057 POR2X1_612/O POR2X1_4/Y 0.01fF
C33058 PAND2X1_488/O POR2X1_532/A 0.04fF
C33059 POR2X1_745/CTRL VDD 0.00fF
C33060 PAND2X1_794/B POR2X1_236/Y 0.02fF
C33061 D_INPUT_2 PAND2X1_14/a_16_344# 0.02fF
C33062 POR2X1_566/A PAND2X1_55/Y 0.03fF
C33063 POR2X1_16/A PAND2X1_214/m4_208_n4# 0.04fF
C33064 PAND2X1_218/A PAND2X1_741/B 0.04fF
C33065 POR2X1_270/CTRL2 POR2X1_814/B 0.05fF
C33066 PAND2X1_241/Y POR2X1_72/B 0.04fF
C33067 PAND2X1_562/CTRL VDD -0.00fF
C33068 POR2X1_856/B POR2X1_724/B 0.02fF
C33069 INPUT_1 POR2X1_32/A 0.06fF
C33070 POR2X1_287/B POR2X1_458/B 0.00fF
C33071 POR2X1_309/Y VDD 0.10fF
C33072 PAND2X1_94/A PAND2X1_77/O 0.02fF
C33073 INPUT_1 PAND2X1_77/CTRL2 0.01fF
C33074 POR2X1_511/Y POR2X1_90/Y 0.03fF
C33075 POR2X1_60/CTRL2 POR2X1_497/Y 0.10fF
C33076 POR2X1_52/A PAND2X1_859/B 0.23fF
C33077 POR2X1_316/Y POR2X1_411/B 0.03fF
C33078 POR2X1_220/A POR2X1_781/B 0.70fF
C33079 POR2X1_52/A PAND2X1_493/Y 0.17fF
C33080 POR2X1_383/A POR2X1_269/Y 0.01fF
C33081 POR2X1_94/A POR2X1_7/A 0.05fF
C33082 POR2X1_270/Y POR2X1_370/O 0.03fF
C33083 PAND2X1_6/A POR2X1_88/Y 0.03fF
C33084 PAND2X1_483/CTRL2 POR2X1_482/Y 0.01fF
C33085 POR2X1_814/B POR2X1_537/B 0.01fF
C33086 POR2X1_420/m4_208_n4# POR2X1_419/m4_208_n4# 0.13fF
C33087 POR2X1_201/m4_208_n4# POR2X1_201/Y 0.09fF
C33088 POR2X1_399/A POR2X1_293/Y 0.01fF
C33089 POR2X1_38/Y PAND2X1_741/B 0.01fF
C33090 POR2X1_32/A POR2X1_153/Y 0.41fF
C33091 VDD PAND2X1_347/CTRL -0.00fF
C33092 POR2X1_439/O POR2X1_180/A 0.00fF
C33093 POR2X1_123/Y VDD 0.00fF
C33094 POR2X1_859/A POR2X1_816/A 0.05fF
C33095 POR2X1_48/A PAND2X1_554/CTRL2 0.01fF
C33096 POR2X1_66/A POR2X1_195/O 0.01fF
C33097 POR2X1_462/B POR2X1_859/A 0.00fF
C33098 POR2X1_859/A D_INPUT_1 0.03fF
C33099 D_INPUT_0 PAND2X1_716/B 0.07fF
C33100 PAND2X1_247/CTRL POR2X1_77/Y 0.01fF
C33101 POR2X1_215/CTRL2 PAND2X1_88/Y 0.01fF
C33102 PAND2X1_602/Y POR2X1_755/CTRL 0.02fF
C33103 PAND2X1_661/Y PAND2X1_660/B 0.03fF
C33104 POR2X1_347/B PAND2X1_69/A 0.18fF
C33105 POR2X1_42/Y PAND2X1_850/CTRL 0.01fF
C33106 POR2X1_839/CTRL2 POR2X1_566/B 0.37fF
C33107 POR2X1_78/A POR2X1_339/Y 0.03fF
C33108 POR2X1_506/a_16_28# POR2X1_506/B -0.00fF
C33109 POR2X1_266/A PAND2X1_73/Y 0.16fF
C33110 PAND2X1_41/B POR2X1_773/B 0.05fF
C33111 PAND2X1_51/O POR2X1_750/B 0.02fF
C33112 PAND2X1_245/O PAND2X1_71/Y 0.02fF
C33113 VDD PAND2X1_99/Y 0.10fF
C33114 POR2X1_376/B PAND2X1_569/B 0.02fF
C33115 POR2X1_257/O PAND2X1_569/Y 0.02fF
C33116 PAND2X1_714/CTRL2 POR2X1_73/Y 0.01fF
C33117 PAND2X1_94/A PAND2X1_395/CTRL 0.01fF
C33118 POR2X1_639/Y PAND2X1_386/Y 0.03fF
C33119 POR2X1_525/CTRL2 PAND2X1_726/B 0.03fF
C33120 PAND2X1_96/B POR2X1_465/B 0.03fF
C33121 POR2X1_485/CTRL PAND2X1_550/B 0.01fF
C33122 POR2X1_805/Y PAND2X1_48/A 0.03fF
C33123 PAND2X1_6/O POR2X1_35/B 0.03fF
C33124 POR2X1_256/CTRL2 POR2X1_7/A 0.05fF
C33125 POR2X1_65/A POR2X1_16/A 0.93fF
C33126 POR2X1_346/B POR2X1_61/Y 0.02fF
C33127 POR2X1_57/CTRL POR2X1_38/Y 0.01fF
C33128 POR2X1_840/CTRL2 PAND2X1_55/Y 0.00fF
C33129 POR2X1_809/A POR2X1_864/CTRL2 0.01fF
C33130 POR2X1_537/Y POR2X1_858/a_16_28# 0.02fF
C33131 PAND2X1_95/B PAND2X1_752/Y 0.01fF
C33132 PAND2X1_20/A PAND2X1_48/A 0.18fF
C33133 PAND2X1_6/Y POR2X1_222/Y 0.03fF
C33134 POR2X1_23/Y POR2X1_184/O 0.01fF
C33135 POR2X1_311/CTRL POR2X1_481/A 0.01fF
C33136 POR2X1_840/B POR2X1_294/B 0.01fF
C33137 POR2X1_734/A POR2X1_734/a_16_28# 0.00fF
C33138 PAND2X1_290/CTRL2 POR2X1_66/A 0.01fF
C33139 POR2X1_861/CTRL2 POR2X1_501/B 0.04fF
C33140 POR2X1_542/B POR2X1_740/Y 0.03fF
C33141 PAND2X1_810/CTRL PAND2X1_366/Y 0.01fF
C33142 PAND2X1_20/A POR2X1_192/B 3.02fF
C33143 POR2X1_198/a_16_28# POR2X1_68/A 0.03fF
C33144 POR2X1_57/A POR2X1_697/Y 0.02fF
C33145 POR2X1_566/A POR2X1_337/A 0.13fF
C33146 POR2X1_63/CTRL POR2X1_38/Y 0.04fF
C33147 POR2X1_128/A POR2X1_735/CTRL 0.05fF
C33148 POR2X1_679/B PAND2X1_735/Y 0.03fF
C33149 POR2X1_750/B PAND2X1_3/B 6.43fF
C33150 PAND2X1_640/B POR2X1_77/Y 0.09fF
C33151 POR2X1_87/Y POR2X1_260/A 0.04fF
C33152 POR2X1_659/O POR2X1_724/A 0.05fF
C33153 POR2X1_72/B POR2X1_371/O 0.01fF
C33154 POR2X1_60/A PAND2X1_352/O 0.02fF
C33155 POR2X1_558/CTRL POR2X1_558/A 0.01fF
C33156 POR2X1_330/Y POR2X1_188/Y 0.05fF
C33157 POR2X1_29/Y POR2X1_409/O 0.09fF
C33158 POR2X1_775/A PAND2X1_173/CTRL 0.01fF
C33159 POR2X1_369/CTRL2 POR2X1_236/Y 0.01fF
C33160 INPUT_1 PAND2X1_38/CTRL2 0.01fF
C33161 PAND2X1_142/O POR2X1_830/A 0.01fF
C33162 POR2X1_57/A PAND2X1_357/Y 0.06fF
C33163 POR2X1_52/A PAND2X1_569/B 0.07fF
C33164 PAND2X1_6/Y POR2X1_532/A 0.43fF
C33165 POR2X1_814/B PAND2X1_48/A 13.81fF
C33166 POR2X1_322/a_16_28# POR2X1_57/A 0.03fF
C33167 POR2X1_49/Y POR2X1_7/Y 0.03fF
C33168 PAND2X1_90/a_16_344# POR2X1_94/A 0.03fF
C33169 INPUT_1 PAND2X1_35/Y 0.06fF
C33170 PAND2X1_651/Y POR2X1_38/Y 0.10fF
C33171 POR2X1_123/Y PAND2X1_32/B 0.01fF
C33172 PAND2X1_605/CTRL2 POR2X1_7/B 0.03fF
C33173 PAND2X1_491/O PAND2X1_96/B 0.10fF
C33174 POR2X1_179/O POR2X1_142/Y 0.10fF
C33175 PAND2X1_684/a_76_28# PAND2X1_90/Y 0.02fF
C33176 PAND2X1_397/CTRL2 POR2X1_35/Y 0.01fF
C33177 PAND2X1_808/Y POR2X1_283/A 0.04fF
C33178 POR2X1_814/B POR2X1_192/B 0.49fF
C33179 PAND2X1_482/O POR2X1_483/A 0.02fF
C33180 POR2X1_219/a_16_28# POR2X1_631/B 0.01fF
C33181 POR2X1_66/A PAND2X1_52/B 0.16fF
C33182 POR2X1_103/CTRL PAND2X1_738/Y 0.01fF
C33183 POR2X1_327/Y POR2X1_115/CTRL2 0.01fF
C33184 PAND2X1_569/B POR2X1_152/A 0.07fF
C33185 POR2X1_740/Y POR2X1_726/Y 0.00fF
C33186 POR2X1_451/A POR2X1_635/A 0.04fF
C33187 PAND2X1_6/Y POR2X1_691/B 0.01fF
C33188 PAND2X1_6/A POR2X1_384/CTRL 0.00fF
C33189 PAND2X1_850/O PAND2X1_842/Y -0.00fF
C33190 PAND2X1_181/m4_208_n4# POR2X1_55/Y 0.07fF
C33191 POR2X1_38/Y PAND2X1_844/B 0.03fF
C33192 PAND2X1_35/Y POR2X1_153/Y 0.05fF
C33193 POR2X1_98/B PAND2X1_88/Y 0.01fF
C33194 POR2X1_287/B PAND2X1_122/CTRL2 0.01fF
C33195 PAND2X1_195/CTRL POR2X1_39/B 0.01fF
C33196 POR2X1_507/B VDD 0.14fF
C33197 POR2X1_840/B PAND2X1_111/B 0.03fF
C33198 POR2X1_206/A POR2X1_294/A 0.03fF
C33199 POR2X1_383/A POR2X1_513/Y 0.10fF
C33200 PAND2X1_69/A POR2X1_713/B 0.06fF
C33201 POR2X1_302/CTRL POR2X1_188/Y 0.01fF
C33202 POR2X1_108/CTRL2 POR2X1_387/Y 0.15fF
C33203 PAND2X1_477/A POR2X1_238/Y 0.07fF
C33204 POR2X1_407/A POR2X1_687/A 0.07fF
C33205 POR2X1_51/A POR2X1_53/a_56_344# 0.01fF
C33206 PAND2X1_779/Y PAND2X1_550/B 0.06fF
C33207 POR2X1_57/A PAND2X1_130/CTRL2 0.01fF
C33208 POR2X1_275/CTRL POR2X1_129/Y 0.01fF
C33209 POR2X1_16/A PAND2X1_190/Y 0.10fF
C33210 POR2X1_346/B POR2X1_35/Y 0.54fF
C33211 POR2X1_327/Y PAND2X1_152/O 0.07fF
C33212 POR2X1_252/Y VDD 0.00fF
C33213 POR2X1_20/B POR2X1_67/Y 0.03fF
C33214 POR2X1_814/B PAND2X1_102/CTRL2 0.05fF
C33215 PAND2X1_90/O POR2X1_546/A 0.01fF
C33216 POR2X1_863/A POR2X1_434/A 0.03fF
C33217 POR2X1_327/Y PAND2X1_48/B 0.20fF
C33218 POR2X1_529/CTRL POR2X1_384/A 0.01fF
C33219 POR2X1_57/A POR2X1_528/Y 9.36fF
C33220 POR2X1_513/B PAND2X1_48/A 0.13fF
C33221 POR2X1_186/Y POR2X1_711/Y 0.08fF
C33222 POR2X1_383/A POR2X1_205/A 0.02fF
C33223 PAND2X1_94/A PAND2X1_767/O 0.01fF
C33224 POR2X1_365/Y POR2X1_357/O 0.00fF
C33225 POR2X1_61/CTRL PAND2X1_69/A 0.01fF
C33226 POR2X1_66/A PAND2X1_125/a_16_344# 0.01fF
C33227 POR2X1_593/O POR2X1_832/B 0.01fF
C33228 POR2X1_8/Y PAND2X1_6/A 0.04fF
C33229 POR2X1_327/O PAND2X1_48/A 0.16fF
C33230 POR2X1_218/A POR2X1_244/Y 0.00fF
C33231 POR2X1_614/A POR2X1_156/Y 0.71fF
C33232 PAND2X1_698/CTRL2 POR2X1_532/A 0.01fF
C33233 PAND2X1_76/Y POR2X1_39/B 0.03fF
C33234 POR2X1_407/Y POR2X1_596/CTRL 0.01fF
C33235 PAND2X1_477/B PAND2X1_308/Y 0.21fF
C33236 POR2X1_184/Y POR2X1_153/Y 0.02fF
C33237 D_INPUT_1 POR2X1_6/CTRL 0.04fF
C33238 PAND2X1_176/O POR2X1_337/Y 0.14fF
C33239 POR2X1_112/CTRL2 POR2X1_579/Y 0.00fF
C33240 POR2X1_124/CTRL2 PAND2X1_41/B 0.05fF
C33241 POR2X1_313/O POR2X1_313/Y 0.01fF
C33242 PAND2X1_704/CTRL2 POR2X1_90/Y 0.00fF
C33243 POR2X1_262/O POR2X1_7/Y 0.01fF
C33244 POR2X1_383/A POR2X1_366/A 0.03fF
C33245 POR2X1_596/A POR2X1_260/A 0.03fF
C33246 POR2X1_447/B POR2X1_785/A 0.07fF
C33247 PAND2X1_651/Y POR2X1_153/Y 0.09fF
C33248 POR2X1_387/Y POR2X1_310/Y 0.04fF
C33249 POR2X1_129/Y POR2X1_90/Y 0.13fF
C33250 POR2X1_834/Y PAND2X1_60/B 0.03fF
C33251 POR2X1_494/a_16_28# POR2X1_384/A 0.03fF
C33252 POR2X1_416/B POR2X1_760/O 0.01fF
C33253 PAND2X1_737/B PAND2X1_656/A 0.03fF
C33254 PAND2X1_655/Y POR2X1_690/CTRL2 0.01fF
C33255 PAND2X1_6/Y POR2X1_552/CTRL 0.01fF
C33256 POR2X1_416/B PAND2X1_362/B 0.03fF
C33257 POR2X1_52/A POR2X1_316/Y 0.05fF
C33258 PAND2X1_736/A PAND2X1_330/O 0.12fF
C33259 POR2X1_218/CTRL2 POR2X1_362/A 0.01fF
C33260 POR2X1_218/CTRL POR2X1_276/Y 0.01fF
C33261 POR2X1_528/Y POR2X1_744/O 0.05fF
C33262 PAND2X1_216/B PAND2X1_656/A 0.02fF
C33263 INPUT_1 POR2X1_9/a_16_28# 0.04fF
C33264 POR2X1_732/B PAND2X1_179/CTRL2 0.21fF
C33265 POR2X1_846/A POR2X1_496/Y 0.01fF
C33266 POR2X1_54/O D_INPUT_1 0.01fF
C33267 PAND2X1_87/CTRL D_INPUT_0 0.01fF
C33268 POR2X1_54/Y POR2X1_411/B 1.13fF
C33269 PAND2X1_425/Y PAND2X1_581/CTRL2 0.01fF
C33270 POR2X1_110/Y POR2X1_417/CTRL2 0.01fF
C33271 POR2X1_553/A POR2X1_456/B 0.01fF
C33272 POR2X1_388/O POR2X1_337/Y 0.14fF
C33273 POR2X1_7/B POR2X1_77/Y 10.18fF
C33274 PAND2X1_81/O POR2X1_4/Y 0.02fF
C33275 POR2X1_327/Y PAND2X1_534/O 0.06fF
C33276 POR2X1_598/O POR2X1_260/A 0.01fF
C33277 PAND2X1_3/m4_208_n4# POR2X1_21/m4_208_n4# 0.05fF
C33278 POR2X1_782/CTRL2 POR2X1_260/A 0.11fF
C33279 PAND2X1_93/B POR2X1_541/B 0.07fF
C33280 POR2X1_294/B PAND2X1_56/A 0.03fF
C33281 POR2X1_222/Y POR2X1_632/Y 0.03fF
C33282 PAND2X1_341/B D_INPUT_3 0.06fF
C33283 POR2X1_119/Y PAND2X1_711/a_56_28# 0.00fF
C33284 POR2X1_730/Y POR2X1_731/A 0.03fF
C33285 PAND2X1_718/CTRL2 POR2X1_77/Y 0.00fF
C33286 PAND2X1_475/CTRL POR2X1_329/A 0.01fF
C33287 POR2X1_121/A POR2X1_711/Y 0.03fF
C33288 POR2X1_703/A POR2X1_543/a_16_28# 0.04fF
C33289 POR2X1_722/a_16_28# PAND2X1_60/B 0.03fF
C33290 POR2X1_212/CTRL2 POR2X1_191/Y 0.25fF
C33291 POR2X1_212/O POR2X1_192/B 0.17fF
C33292 PAND2X1_339/Y PAND2X1_339/O 0.00fF
C33293 PAND2X1_635/Y INPUT_7 0.03fF
C33294 POR2X1_394/A PAND2X1_124/a_76_28# 0.02fF
C33295 POR2X1_438/CTRL2 POR2X1_77/Y 0.11fF
C33296 PAND2X1_23/Y POR2X1_717/B 0.09fF
C33297 PAND2X1_830/m4_208_n4# PAND2X1_114/m4_208_n4# 0.15fF
C33298 POR2X1_25/Y POR2X1_26/CTRL2 0.01fF
C33299 POR2X1_65/CTRL2 POR2X1_40/Y 0.03fF
C33300 PAND2X1_422/a_76_28# PAND2X1_93/B 0.04fF
C33301 PAND2X1_696/O PAND2X1_60/B 0.02fF
C33302 POR2X1_532/A POR2X1_632/Y 0.08fF
C33303 GATE_222 VDD 0.00fF
C33304 INPUT_1 POR2X1_294/A 0.04fF
C33305 POR2X1_118/a_56_344# POR2X1_77/Y 0.00fF
C33306 POR2X1_41/B POR2X1_846/O 0.08fF
C33307 POR2X1_245/Y PAND2X1_508/B 0.03fF
C33308 POR2X1_431/a_76_344# PAND2X1_390/Y 0.00fF
C33309 POR2X1_837/B VDD 0.28fF
C33310 POR2X1_848/CTRL PAND2X1_90/Y 0.02fF
C33311 POR2X1_687/a_16_28# POR2X1_452/Y 0.02fF
C33312 POR2X1_245/O POR2X1_39/B 0.01fF
C33313 POR2X1_67/Y PAND2X1_381/CTRL2 0.01fF
C33314 POR2X1_416/B POR2X1_745/Y 0.01fF
C33315 POR2X1_334/Y POR2X1_351/B 0.04fF
C33316 POR2X1_23/Y PAND2X1_214/CTRL2 0.01fF
C33317 PAND2X1_138/CTRL POR2X1_129/Y 0.01fF
C33318 PAND2X1_635/Y INPUT_4 0.13fF
C33319 POR2X1_532/A PAND2X1_52/B 13.87fF
C33320 POR2X1_192/a_16_28# POR2X1_192/B 0.09fF
C33321 POR2X1_773/B PAND2X1_122/O -0.01fF
C33322 POR2X1_317/A POR2X1_169/A 0.02fF
C33323 POR2X1_655/A POR2X1_590/A 0.05fF
C33324 POR2X1_315/Y POR2X1_39/B 0.07fF
C33325 POR2X1_153/Y PAND2X1_199/CTRL2 0.05fF
C33326 PAND2X1_358/A PAND2X1_101/B -0.00fF
C33327 POR2X1_768/Y POR2X1_294/A 0.06fF
C33328 POR2X1_260/B POR2X1_241/B 0.03fF
C33329 POR2X1_43/B PAND2X1_860/A 0.08fF
C33330 PAND2X1_431/CTRL2 POR2X1_590/A 0.07fF
C33331 POR2X1_809/CTRL2 POR2X1_121/B 0.03fF
C33332 POR2X1_815/CTRL2 INPUT_0 0.21fF
C33333 POR2X1_691/B PAND2X1_52/B 0.02fF
C33334 POR2X1_814/A POR2X1_192/Y 0.10fF
C33335 PAND2X1_472/CTRL2 POR2X1_39/B 0.03fF
C33336 POR2X1_714/O PAND2X1_72/A 0.01fF
C33337 POR2X1_166/O POR2X1_167/Y 0.18fF
C33338 POR2X1_814/B POR2X1_461/Y 0.01fF
C33339 POR2X1_49/Y POR2X1_257/A 0.17fF
C33340 POR2X1_719/A POR2X1_260/B 0.10fF
C33341 PAND2X1_39/B POR2X1_288/A 0.03fF
C33342 POR2X1_499/A POR2X1_778/O 0.01fF
C33343 POR2X1_83/Y PAND2X1_341/B 0.35fF
C33344 PAND2X1_47/B PAND2X1_3/A 0.02fF
C33345 INPUT_3 POR2X1_376/Y 0.04fF
C33346 POR2X1_66/B PAND2X1_93/B 0.18fF
C33347 POR2X1_54/Y PAND2X1_55/O 0.03fF
C33348 POR2X1_54/Y POR2X1_376/B 0.07fF
C33349 POR2X1_68/A POR2X1_98/A 0.01fF
C33350 POR2X1_415/A POR2X1_5/Y 0.03fF
C33351 POR2X1_556/A POR2X1_370/Y 0.03fF
C33352 PAND2X1_443/CTRL2 PAND2X1_803/A 0.00fF
C33353 PAND2X1_605/a_76_28# POR2X1_604/Y 0.03fF
C33354 POR2X1_465/a_16_28# POR2X1_465/A 0.03fF
C33355 POR2X1_862/A POR2X1_734/A 0.02fF
C33356 PAND2X1_48/B PAND2X1_53/CTRL 0.01fF
C33357 POR2X1_188/A PAND2X1_93/B 0.01fF
C33358 POR2X1_864/A PAND2X1_57/B 0.00fF
C33359 POR2X1_612/Y POR2X1_414/Y 0.03fF
C33360 POR2X1_445/A PAND2X1_90/Y 0.10fF
C33361 PAND2X1_847/CTRL2 POR2X1_394/A 0.32fF
C33362 PAND2X1_217/B PAND2X1_576/B 0.00fF
C33363 POR2X1_326/A POR2X1_736/A 0.39fF
C33364 PAND2X1_309/CTRL POR2X1_556/A 0.00fF
C33365 POR2X1_676/CTRL VDD 0.00fF
C33366 POR2X1_14/Y POR2X1_102/Y 0.13fF
C33367 POR2X1_257/A PAND2X1_274/O 0.01fF
C33368 POR2X1_850/B PAND2X1_58/A 0.03fF
C33369 PAND2X1_214/A POR2X1_32/A 0.01fF
C33370 POR2X1_476/A POR2X1_476/a_16_28# 0.02fF
C33371 POR2X1_66/B POR2X1_78/A 0.10fF
C33372 PAND2X1_453/A POR2X1_102/Y 0.03fF
C33373 POR2X1_847/B POR2X1_48/A 0.03fF
C33374 POR2X1_641/O POR2X1_267/A 0.18fF
C33375 PAND2X1_217/CTRL PAND2X1_364/B 0.03fF
C33376 POR2X1_470/O POR2X1_186/Y 0.04fF
C33377 POR2X1_48/A PAND2X1_76/Y 0.03fF
C33378 PAND2X1_287/Y PAND2X1_347/Y 0.65fF
C33379 PAND2X1_124/Y POR2X1_236/Y 0.07fF
C33380 POR2X1_263/Y POR2X1_230/CTRL 0.01fF
C33381 PAND2X1_51/CTRL2 POR2X1_451/A 0.01fF
C33382 POR2X1_48/A POR2X1_689/CTRL 0.01fF
C33383 PAND2X1_487/CTRL PAND2X1_57/B 0.01fF
C33384 PAND2X1_257/O POR2X1_510/Y 0.01fF
C33385 POR2X1_257/A PAND2X1_553/B 0.91fF
C33386 POR2X1_188/A POR2X1_78/A 0.06fF
C33387 POR2X1_52/A POR2X1_54/Y 0.01fF
C33388 POR2X1_179/CTRL POR2X1_150/Y 0.01fF
C33389 PAND2X1_73/Y POR2X1_734/A 0.45fF
C33390 POR2X1_9/Y POR2X1_283/A 0.17fF
C33391 PAND2X1_9/Y POR2X1_42/Y 0.03fF
C33392 POR2X1_667/a_16_28# POR2X1_73/Y 0.07fF
C33393 POR2X1_624/Y POR2X1_404/Y 0.03fF
C33394 PAND2X1_410/CTRL2 POR2X1_290/Y 0.02fF
C33395 POR2X1_863/A POR2X1_544/B 0.03fF
C33396 PAND2X1_576/B VDD 0.12fF
C33397 PAND2X1_75/CTRL2 PAND2X1_60/B 0.00fF
C33398 POR2X1_41/B POR2X1_265/CTRL2 0.00fF
C33399 PAND2X1_810/B PAND2X1_365/B 0.01fF
C33400 POR2X1_661/CTRL POR2X1_78/A 0.08fF
C33401 POR2X1_83/B POR2X1_677/CTRL 0.01fF
C33402 POR2X1_142/O POR2X1_49/Y 0.01fF
C33403 POR2X1_452/Y POR2X1_730/CTRL 0.01fF
C33404 POR2X1_482/Y POR2X1_72/B 0.03fF
C33405 POR2X1_864/A POR2X1_828/A 0.40fF
C33406 POR2X1_479/B VDD 0.04fF
C33407 PAND2X1_267/Y PAND2X1_364/B 0.25fF
C33408 PAND2X1_492/CTRL2 PAND2X1_73/Y 0.13fF
C33409 POR2X1_770/B POR2X1_770/A 0.03fF
C33410 POR2X1_397/Y POR2X1_669/B 0.07fF
C33411 POR2X1_640/O PAND2X1_41/B 0.01fF
C33412 POR2X1_102/Y POR2X1_237/CTRL 0.01fF
C33413 POR2X1_67/A VDD 0.85fF
C33414 PAND2X1_497/CTRL POR2X1_294/B 0.20fF
C33415 POR2X1_813/CTRL2 POR2X1_38/Y 0.03fF
C33416 PAND2X1_104/O POR2X1_814/B 0.03fF
C33417 POR2X1_83/B POR2X1_236/Y 5.99fF
C33418 POR2X1_831/O PAND2X1_69/A 0.01fF
C33419 PAND2X1_416/CTRL POR2X1_816/A 0.00fF
C33420 POR2X1_796/Y POR2X1_803/A 0.02fF
C33421 PAND2X1_206/B PAND2X1_100/CTRL2 0.00fF
C33422 PAND2X1_90/Y PAND2X1_585/O 0.08fF
C33423 POR2X1_251/A POR2X1_106/Y 0.11fF
C33424 POR2X1_828/Y POR2X1_750/B 0.03fF
C33425 PAND2X1_48/B PAND2X1_485/O 0.19fF
C33426 PAND2X1_6/Y POR2X1_808/CTRL2 0.00fF
C33427 POR2X1_805/CTRL POR2X1_805/A 0.00fF
C33428 POR2X1_814/B POR2X1_288/A 0.03fF
C33429 POR2X1_556/A POR2X1_216/O 0.01fF
C33430 PAND2X1_787/A POR2X1_411/B 0.03fF
C33431 POR2X1_566/A POR2X1_174/A 0.07fF
C33432 PAND2X1_659/B PAND2X1_573/B 0.16fF
C33433 PAND2X1_487/CTRL2 PAND2X1_69/A 0.01fF
C33434 POR2X1_308/CTRL POR2X1_794/B 0.02fF
C33435 PAND2X1_706/O POR2X1_692/Y 0.01fF
C33436 POR2X1_856/B POR2X1_740/Y 0.03fF
C33437 POR2X1_623/A POR2X1_623/Y 0.04fF
C33438 PAND2X1_246/O POR2X1_101/Y 0.04fF
C33439 PAND2X1_423/CTRL POR2X1_807/A 0.01fF
C33440 POR2X1_78/B POR2X1_200/CTRL 0.01fF
C33441 PAND2X1_95/B POR2X1_66/A 0.05fF
C33442 POR2X1_78/A POR2X1_724/a_76_344# 0.01fF
C33443 POR2X1_441/Y PAND2X1_854/A 0.01fF
C33444 POR2X1_862/CTRL PAND2X1_52/B 0.01fF
C33445 POR2X1_418/Y VDD 0.12fF
C33446 GATE_479 PAND2X1_803/A 0.05fF
C33447 POR2X1_23/Y PAND2X1_705/O 0.03fF
C33448 POR2X1_533/Y POR2X1_759/O 0.02fF
C33449 PAND2X1_20/A PAND2X1_516/O 0.02fF
C33450 POR2X1_3/A PAND2X1_12/CTRL2 0.20fF
C33451 PAND2X1_404/Y POR2X1_73/Y 0.05fF
C33452 POR2X1_186/Y PAND2X1_321/a_16_344# 0.03fF
C33453 PAND2X1_73/Y POR2X1_828/O 0.01fF
C33454 POR2X1_48/A PAND2X1_566/Y 0.07fF
C33455 POR2X1_533/A VDD 0.15fF
C33456 PAND2X1_244/CTRL POR2X1_293/Y 0.00fF
C33457 PAND2X1_212/CTRL2 POR2X1_142/Y 0.00fF
C33458 PAND2X1_55/Y POR2X1_241/B 0.03fF
C33459 PAND2X1_214/A PAND2X1_35/Y 0.00fF
C33460 PAND2X1_222/A PAND2X1_222/B 0.10fF
C33461 POR2X1_102/Y POR2X1_55/Y 7.54fF
C33462 POR2X1_130/A POR2X1_860/A 0.03fF
C33463 POR2X1_60/A PAND2X1_254/CTRL 0.01fF
C33464 POR2X1_284/CTRL2 POR2X1_330/Y 0.51fF
C33465 PAND2X1_776/Y PAND2X1_785/A 0.00fF
C33466 POR2X1_467/Y POR2X1_802/B 0.32fF
C33467 PAND2X1_768/Y PAND2X1_347/Y 0.02fF
C33468 POR2X1_528/CTRL2 POR2X1_14/Y 0.00fF
C33469 PAND2X1_390/Y POR2X1_46/Y 0.05fF
C33470 POR2X1_852/B POR2X1_192/Y 0.10fF
C33471 POR2X1_37/Y POR2X1_90/Y 0.07fF
C33472 POR2X1_41/B POR2X1_750/B 1.09fF
C33473 PAND2X1_63/Y D_INPUT_0 0.05fF
C33474 POR2X1_528/CTRL2 PAND2X1_453/A 0.01fF
C33475 PAND2X1_20/A PAND2X1_95/O 0.00fF
C33476 POR2X1_379/CTRL2 POR2X1_260/B 0.03fF
C33477 POR2X1_315/Y PAND2X1_469/CTRL2 0.05fF
C33478 POR2X1_479/B PAND2X1_32/B 0.03fF
C33479 PAND2X1_6/Y POR2X1_660/Y 0.03fF
C33480 POR2X1_519/O PAND2X1_838/B 0.01fF
C33481 POR2X1_141/Y POR2X1_276/CTRL2 0.00fF
C33482 POR2X1_105/Y POR2X1_723/O 0.02fF
C33483 PAND2X1_319/CTRL VDD 0.00fF
C33484 PAND2X1_94/A POR2X1_473/CTRL2 0.05fF
C33485 PAND2X1_41/B POR2X1_208/CTRL2 0.01fF
C33486 POR2X1_72/Y POR2X1_72/B 0.04fF
C33487 PAND2X1_733/Y VDD 0.00fF
C33488 POR2X1_849/A POR2X1_550/O 0.01fF
C33489 POR2X1_511/Y INPUT_0 0.07fF
C33490 POR2X1_557/A POR2X1_624/Y 0.03fF
C33491 POR2X1_329/A PAND2X1_851/a_16_344# 0.01fF
C33492 POR2X1_401/CTRL2 POR2X1_401/B 0.01fF
C33493 POR2X1_287/B POR2X1_784/A 0.03fF
C33494 PAND2X1_614/O POR2X1_42/Y 0.14fF
C33495 POR2X1_122/CTRL POR2X1_20/B 0.01fF
C33496 PAND2X1_377/CTRL VDD -0.00fF
C33497 POR2X1_464/Y POR2X1_543/A 0.21fF
C33498 PAND2X1_431/a_56_28# PAND2X1_60/B 0.00fF
C33499 PAND2X1_139/Y VDD -0.00fF
C33500 POR2X1_624/Y PAND2X1_184/O 0.02fF
C33501 POR2X1_32/A POR2X1_591/Y 0.06fF
C33502 POR2X1_194/B VDD 0.02fF
C33503 PAND2X1_552/B POR2X1_312/Y 1.15fF
C33504 PAND2X1_455/Y VDD 0.00fF
C33505 PAND2X1_565/CTRL2 POR2X1_40/Y 0.01fF
C33506 POR2X1_56/B POR2X1_5/Y 0.01fF
C33507 POR2X1_97/O POR2X1_454/A 0.05fF
C33508 POR2X1_814/B POR2X1_789/Y 0.01fF
C33509 PAND2X1_198/Y VDD 0.00fF
C33510 POR2X1_355/A D_GATE_741 0.03fF
C33511 POR2X1_355/CTRL2 D_GATE_741 0.02fF
C33512 POR2X1_333/A POR2X1_775/a_56_344# 0.03fF
C33513 POR2X1_65/A POR2X1_761/O 0.01fF
C33514 POR2X1_72/B POR2X1_406/A 0.01fF
C33515 POR2X1_49/Y POR2X1_817/Y 0.00fF
C33516 POR2X1_65/A PAND2X1_324/Y 1.38fF
C33517 POR2X1_865/B POR2X1_474/CTRL2 0.10fF
C33518 POR2X1_57/A POR2X1_667/A 0.03fF
C33519 POR2X1_486/B POR2X1_814/A 1.24fF
C33520 PAND2X1_862/B PAND2X1_735/Y 0.07fF
C33521 POR2X1_338/a_16_28# POR2X1_567/B 0.10fF
C33522 POR2X1_16/A PAND2X1_645/Y 0.03fF
C33523 POR2X1_776/B VDD 0.74fF
C33524 POR2X1_776/A PAND2X1_171/O 0.07fF
C33525 PAND2X1_260/a_16_344# PAND2X1_566/Y 0.04fF
C33526 POR2X1_12/A POR2X1_762/CTRL2 0.01fF
C33527 POR2X1_555/B POR2X1_510/Y 0.03fF
C33528 PAND2X1_472/CTRL POR2X1_23/Y 0.00fF
C33529 PAND2X1_824/a_76_28# POR2X1_856/B 0.01fF
C33530 PAND2X1_824/m4_208_n4# POR2X1_567/B 0.06fF
C33531 POR2X1_409/B PAND2X1_196/O 0.02fF
C33532 POR2X1_467/Y POR2X1_532/A 0.03fF
C33533 PAND2X1_62/CTRL2 PAND2X1_6/A 0.03fF
C33534 POR2X1_66/A PAND2X1_373/a_16_344# 0.01fF
C33535 D_INPUT_3 POR2X1_14/m4_208_n4# 0.09fF
C33536 POR2X1_226/a_16_28# POR2X1_382/Y 0.07fF
C33537 POR2X1_226/Y POR2X1_382/a_16_28# 0.01fF
C33538 PAND2X1_241/O VDD 0.00fF
C33539 POR2X1_35/B PAND2X1_69/A 0.03fF
C33540 PAND2X1_460/Y POR2X1_7/B 0.01fF
C33541 POR2X1_529/CTRL2 VDD -0.00fF
C33542 PAND2X1_659/CTRL2 PAND2X1_575/A 0.01fF
C33543 POR2X1_669/B POR2X1_511/a_16_28# 0.03fF
C33544 PAND2X1_249/O POR2X1_38/Y 0.00fF
C33545 PAND2X1_414/CTRL2 POR2X1_39/B 0.00fF
C33546 POR2X1_51/B POR2X1_32/A 0.04fF
C33547 POR2X1_411/B POR2X1_4/Y 0.12fF
C33548 POR2X1_13/A PAND2X1_351/O 0.03fF
C33549 PAND2X1_65/B PAND2X1_744/O 0.07fF
C33550 POR2X1_94/A POR2X1_38/Y 0.03fF
C33551 PAND2X1_216/B PAND2X1_561/CTRL2 0.00fF
C33552 PAND2X1_218/B POR2X1_394/A 0.03fF
C33553 POR2X1_93/A POR2X1_40/Y 0.02fF
C33554 PAND2X1_808/Y POR2X1_488/a_16_28# 0.05fF
C33555 D_INPUT_0 POR2X1_260/A 0.13fF
C33556 POR2X1_811/A POR2X1_260/A 0.00fF
C33557 PAND2X1_206/B POR2X1_77/Y 0.07fF
C33558 POR2X1_403/O PAND2X1_69/A 0.01fF
C33559 PAND2X1_94/A POR2X1_29/A 0.03fF
C33560 POR2X1_72/B POR2X1_511/CTRL 0.01fF
C33561 PAND2X1_812/a_76_28# PAND2X1_805/A 0.01fF
C33562 PAND2X1_830/Y PAND2X1_114/Y 0.24fF
C33563 POR2X1_85/Y PAND2X1_206/B 0.03fF
C33564 POR2X1_102/Y POR2X1_7/CTRL2 0.01fF
C33565 PAND2X1_351/CTRL POR2X1_293/Y 0.02fF
C33566 POR2X1_697/Y POR2X1_531/CTRL2 0.01fF
C33567 PAND2X1_470/A POR2X1_417/Y 0.02fF
C33568 POR2X1_23/Y PAND2X1_713/O 0.02fF
C33569 PAND2X1_469/B PAND2X1_556/B 0.49fF
C33570 POR2X1_828/Y POR2X1_686/CTRL2 0.00fF
C33571 POR2X1_740/Y POR2X1_722/Y 0.02fF
C33572 POR2X1_423/Y POR2X1_387/Y 0.09fF
C33573 POR2X1_45/Y PAND2X1_804/B 0.01fF
C33574 POR2X1_348/A POR2X1_197/Y 0.01fF
C33575 POR2X1_671/CTRL2 POR2X1_38/B 0.01fF
C33576 PAND2X1_642/B VDD 0.30fF
C33577 POR2X1_281/O POR2X1_102/Y 0.01fF
C33578 PAND2X1_632/B POR2X1_60/A 0.01fF
C33579 POR2X1_72/B PAND2X1_349/A 0.03fF
C33580 INPUT_6 POR2X1_763/A 0.07fF
C33581 PAND2X1_6/A POR2X1_516/B 0.07fF
C33582 POR2X1_213/m4_208_n4# PAND2X1_320/m4_208_n4# 0.13fF
C33583 POR2X1_36/B INPUT_7 0.07fF
C33584 POR2X1_682/a_16_28# POR2X1_591/Y 0.03fF
C33585 POR2X1_251/A PAND2X1_114/B 0.05fF
C33586 PAND2X1_585/m4_208_n4# POR2X1_758/m4_208_n4# 0.13fF
C33587 POR2X1_102/Y PAND2X1_508/O 0.05fF
C33588 POR2X1_614/A POR2X1_676/Y 0.01fF
C33589 POR2X1_383/A POR2X1_509/B 0.03fF
C33590 POR2X1_507/CTRL2 POR2X1_355/A 0.01fF
C33591 POR2X1_66/A POR2X1_722/CTRL2 0.01fF
C33592 POR2X1_789/A POR2X1_790/CTRL 0.03fF
C33593 POR2X1_770/B POR2X1_774/A 0.01fF
C33594 POR2X1_800/A POR2X1_783/B 0.00fF
C33595 POR2X1_276/A POR2X1_274/Y 0.01fF
C33596 POR2X1_65/A PAND2X1_549/B 0.07fF
C33597 POR2X1_333/Y POR2X1_241/B 0.01fF
C33598 POR2X1_83/A POR2X1_293/Y 0.03fF
C33599 POR2X1_265/Y POR2X1_263/Y 0.92fF
C33600 PAND2X1_545/Y POR2X1_40/Y 0.01fF
C33601 PAND2X1_564/a_76_28# PAND2X1_551/Y 0.07fF
C33602 POR2X1_335/A PAND2X1_48/B 0.03fF
C33603 POR2X1_566/A POR2X1_447/CTRL2 0.15fF
C33604 PAND2X1_56/Y POR2X1_832/B 0.01fF
C33605 PAND2X1_41/B POR2X1_116/Y 0.02fF
C33606 PAND2X1_58/A POR2X1_720/CTRL2 0.09fF
C33607 POR2X1_32/A POR2X1_150/CTRL2 0.03fF
C33608 PAND2X1_372/O POR2X1_778/B 0.01fF
C33609 POR2X1_447/B POR2X1_836/CTRL 0.01fF
C33610 POR2X1_508/B POR2X1_836/CTRL2 0.00fF
C33611 POR2X1_13/A POR2X1_289/a_16_28# 0.03fF
C33612 INPUT_1 POR2X1_94/A 0.06fF
C33613 POR2X1_725/Y POR2X1_830/A 0.07fF
C33614 PAND2X1_183/m4_208_n4# POR2X1_732/B 0.05fF
C33615 PAND2X1_803/O POR2X1_83/B 0.05fF
C33616 POR2X1_205/A INPUT_0 0.07fF
C33617 POR2X1_730/Y PAND2X1_41/B 0.02fF
C33618 POR2X1_260/B PAND2X1_136/O 0.02fF
C33619 POR2X1_368/CTRL POR2X1_387/Y 0.07fF
C33620 POR2X1_776/B PAND2X1_32/B 0.03fF
C33621 VDD PAND2X1_168/O 0.00fF
C33622 POR2X1_90/Y POR2X1_293/Y 0.19fF
C33623 PAND2X1_845/CTRL POR2X1_55/Y 0.00fF
C33624 POR2X1_861/CTRL POR2X1_218/A 0.01fF
C33625 POR2X1_537/B VDD 0.04fF
C33626 POR2X1_833/A PAND2X1_46/a_16_344# 0.02fF
C33627 PAND2X1_350/CTRL POR2X1_88/Y 0.01fF
C33628 POR2X1_65/A POR2X1_41/CTRL 0.01fF
C33629 POR2X1_38/Y POR2X1_406/CTRL2 0.00fF
C33630 PAND2X1_773/Y POR2X1_767/Y 0.03fF
C33631 PAND2X1_65/B PAND2X1_103/CTRL 0.00fF
C33632 POR2X1_3/A INPUT_5 0.18fF
C33633 PAND2X1_6/A POR2X1_619/O 0.02fF
C33634 POR2X1_36/B INPUT_4 1.00fF
C33635 POR2X1_452/Y PAND2X1_52/B 0.70fF
C33636 POR2X1_447/B PAND2X1_39/CTRL 0.06fF
C33637 POR2X1_143/O D_INPUT_3 0.17fF
C33638 POR2X1_563/CTRL2 POR2X1_456/B 0.12fF
C33639 PAND2X1_728/CTRL2 VDD 0.00fF
C33640 POR2X1_111/O POR2X1_293/Y 0.12fF
C33641 PAND2X1_852/B POR2X1_42/Y 0.00fF
C33642 POR2X1_368/O POR2X1_283/A 0.02fF
C33643 POR2X1_516/Y PAND2X1_851/O 0.04fF
C33644 POR2X1_278/Y POR2X1_283/A 0.07fF
C33645 POR2X1_518/CTRL POR2X1_669/B 0.06fF
C33646 INPUT_1 POR2X1_381/O 0.01fF
C33647 PAND2X1_550/B VDD 0.52fF
C33648 PAND2X1_90/Y POR2X1_260/A 0.05fF
C33649 PAND2X1_241/Y POR2X1_7/B 0.00fF
C33650 POR2X1_460/CTRL PAND2X1_32/B 0.01fF
C33651 POR2X1_122/Y POR2X1_16/A 0.01fF
C33652 POR2X1_808/CTRL2 PAND2X1_52/B 0.17fF
C33653 POR2X1_90/Y PAND2X1_302/a_16_344# 0.01fF
C33654 PAND2X1_770/a_76_28# POR2X1_765/Y 0.01fF
C33655 POR2X1_341/A POR2X1_715/a_56_344# 0.01fF
C33656 PAND2X1_768/O POR2X1_103/Y -0.00fF
C33657 POR2X1_119/Y POR2X1_609/CTRL2 0.02fF
C33658 PAND2X1_57/B POR2X1_553/A 0.03fF
C33659 POR2X1_218/A POR2X1_501/B 0.07fF
C33660 POR2X1_22/A POR2X1_3/O 0.01fF
C33661 PAND2X1_787/A POR2X1_152/A 0.02fF
C33662 POR2X1_640/A POR2X1_559/A 0.05fF
C33663 POR2X1_675/A POR2X1_186/B 0.01fF
C33664 POR2X1_407/A POR2X1_840/B 0.05fF
C33665 POR2X1_99/B POR2X1_244/CTRL2 0.00fF
C33666 POR2X1_68/A POR2X1_844/CTRL2 0.00fF
C33667 PAND2X1_762/O PAND2X1_52/B 0.01fF
C33668 POR2X1_198/a_56_344# PAND2X1_88/Y 0.00fF
C33669 PAND2X1_464/Y POR2X1_73/Y 0.03fF
C33670 PAND2X1_6/A POR2X1_68/B 0.01fF
C33671 POR2X1_614/A POR2X1_203/Y 0.01fF
C33672 POR2X1_46/Y PAND2X1_123/O 0.10fF
C33673 POR2X1_554/Y POR2X1_569/A 0.09fF
C33674 POR2X1_548/B PAND2X1_63/B 0.76fF
C33675 POR2X1_57/A PAND2X1_182/CTRL2 0.03fF
C33676 POR2X1_73/Y PAND2X1_565/A 0.01fF
C33677 PAND2X1_865/Y PAND2X1_557/A 0.02fF
C33678 PAND2X1_760/O POR2X1_260/A 0.04fF
C33679 PAND2X1_798/Y PAND2X1_807/B 0.02fF
C33680 POR2X1_52/A PAND2X1_160/CTRL 0.01fF
C33681 POR2X1_163/A PAND2X1_160/CTRL2 0.03fF
C33682 POR2X1_500/Y POR2X1_576/Y 0.01fF
C33683 POR2X1_711/B POR2X1_710/A 0.56fF
C33684 POR2X1_376/B POR2X1_701/CTRL2 0.05fF
C33685 POR2X1_729/O POR2X1_687/Y 0.17fF
C33686 POR2X1_181/B PAND2X1_178/O 0.00fF
C33687 PAND2X1_192/CTRL PAND2X1_730/A 0.00fF
C33688 POR2X1_68/A POR2X1_845/CTRL2 0.09fF
C33689 PAND2X1_714/A PAND2X1_714/B 0.03fF
C33690 PAND2X1_737/a_76_28# POR2X1_40/Y 0.01fF
C33691 PAND2X1_48/B POR2X1_249/Y 0.00fF
C33692 PAND2X1_477/B PAND2X1_241/Y 0.35fF
C33693 PAND2X1_94/A PAND2X1_110/CTRL 0.12fF
C33694 INPUT_0 POR2X1_129/Y 0.05fF
C33695 POR2X1_220/B PAND2X1_52/B 0.00fF
C33696 POR2X1_180/CTRL VDD -0.00fF
C33697 PAND2X1_533/CTRL2 POR2X1_802/B 0.03fF
C33698 POR2X1_40/Y PAND2X1_169/CTRL2 0.01fF
C33699 POR2X1_334/Y PAND2X1_257/CTRL2 0.04fF
C33700 POR2X1_139/A POR2X1_318/A 0.02fF
C33701 POR2X1_863/CTRL2 POR2X1_260/A 0.01fF
C33702 POR2X1_334/A PAND2X1_57/B 0.03fF
C33703 POR2X1_376/B POR2X1_4/Y 0.13fF
C33704 PAND2X1_115/CTRL2 PAND2X1_348/A 0.00fF
C33705 POR2X1_220/Y POR2X1_186/B 0.03fF
C33706 POR2X1_79/Y PAND2X1_853/B 0.03fF
C33707 PAND2X1_793/Y POR2X1_394/A 0.05fF
C33708 VDD PAND2X1_48/A 3.49fF
C33709 POR2X1_41/B PAND2X1_560/B 0.03fF
C33710 POR2X1_391/CTRL2 PAND2X1_32/B 0.00fF
C33711 POR2X1_710/O POR2X1_710/B 0.00fF
C33712 PAND2X1_94/A POR2X1_805/A 0.07fF
C33713 POR2X1_83/Y POR2X1_497/Y 0.02fF
C33714 POR2X1_399/O POR2X1_119/Y 0.28fF
C33715 VDD POR2X1_192/B 5.00fF
C33716 PAND2X1_659/Y INPUT_0 0.06fF
C33717 POR2X1_81/CTRL2 POR2X1_293/Y 0.03fF
C33718 POR2X1_662/Y POR2X1_741/B 0.07fF
C33719 POR2X1_404/Y POR2X1_186/B 0.03fF
C33720 POR2X1_751/Y POR2X1_42/Y 0.05fF
C33721 PAND2X1_735/Y PAND2X1_716/B 0.07fF
C33722 PAND2X1_481/O POR2X1_294/B 0.15fF
C33723 POR2X1_456/B PAND2X1_316/O 0.02fF
C33724 PAND2X1_811/Y PAND2X1_568/B 0.06fF
C33725 PAND2X1_216/B POR2X1_183/Y 0.21fF
C33726 PAND2X1_787/O POR2X1_39/B 0.01fF
C33727 POR2X1_68/B POR2X1_101/Y 0.07fF
C33728 POR2X1_854/CTRL2 POR2X1_854/B 0.01fF
C33729 POR2X1_96/Y INPUT_0 0.01fF
C33730 POR2X1_16/A PAND2X1_398/a_76_28# 0.01fF
C33731 PAND2X1_220/Y POR2X1_77/Y 0.03fF
C33732 PAND2X1_292/CTRL2 PAND2X1_41/B 0.03fF
C33733 POR2X1_265/Y PAND2X1_215/B 0.20fF
C33734 POR2X1_394/A POR2X1_665/Y 0.00fF
C33735 POR2X1_110/Y POR2X1_293/Y 0.02fF
C33736 POR2X1_547/CTRL POR2X1_266/A 0.01fF
C33737 POR2X1_52/A POR2X1_4/Y 0.03fF
C33738 POR2X1_394/A PAND2X1_302/a_76_28# 0.01fF
C33739 POR2X1_596/A POR2X1_596/O 0.01fF
C33740 POR2X1_68/A POR2X1_370/CTRL 0.01fF
C33741 POR2X1_532/A PAND2X1_533/CTRL2 0.01fF
C33742 POR2X1_327/Y POR2X1_861/a_16_28# 0.02fF
C33743 POR2X1_43/B PAND2X1_156/A 0.05fF
C33744 POR2X1_346/B POR2X1_631/A 0.02fF
C33745 PAND2X1_675/A POR2X1_103/a_16_28# 0.02fF
C33746 PAND2X1_659/Y PAND2X1_218/CTRL 0.00fF
C33747 POR2X1_390/B PAND2X1_60/B 0.03fF
C33748 PAND2X1_342/CTRL POR2X1_153/Y 0.06fF
C33749 PAND2X1_798/B PAND2X1_657/B 0.27fF
C33750 POR2X1_301/A POR2X1_814/A 0.02fF
C33751 POR2X1_440/Y POR2X1_738/A 0.03fF
C33752 POR2X1_750/B POR2X1_161/a_16_28# 0.05fF
C33753 VDD PAND2X1_840/Y 0.14fF
C33754 POR2X1_809/A PAND2X1_583/CTRL 0.01fF
C33755 PAND2X1_57/B D_INPUT_4 0.10fF
C33756 PAND2X1_480/B POR2X1_39/B 0.05fF
C33757 POR2X1_376/B POR2X1_80/a_16_28# 0.02fF
C33758 PAND2X1_440/O PAND2X1_580/B 0.00fF
C33759 PAND2X1_797/Y PAND2X1_714/a_76_28# 0.02fF
C33760 PAND2X1_209/A POR2X1_146/Y 0.02fF
C33761 POR2X1_360/A PAND2X1_290/O 0.10fF
C33762 PAND2X1_446/Y PAND2X1_466/B 0.26fF
C33763 POR2X1_754/A POR2X1_39/B 0.06fF
C33764 PAND2X1_48/A PAND2X1_32/B 0.25fF
C33765 POR2X1_57/A PAND2X1_170/O 0.04fF
C33766 POR2X1_96/B POR2X1_96/O 0.02fF
C33767 POR2X1_329/A D_INPUT_0 0.07fF
C33768 POR2X1_348/O POR2X1_244/Y 0.05fF
C33769 PAND2X1_96/B POR2X1_113/B 0.03fF
C33770 POR2X1_722/A PAND2X1_60/B 0.24fF
C33771 POR2X1_192/B PAND2X1_32/B 0.05fF
C33772 POR2X1_14/Y POR2X1_9/Y 0.11fF
C33773 PAND2X1_653/Y POR2X1_7/Y 0.03fF
C33774 PAND2X1_841/CTRL2 POR2X1_39/B 0.03fF
C33775 POR2X1_98/A PAND2X1_58/A 0.01fF
C33776 POR2X1_456/B PAND2X1_313/CTRL2 0.01fF
C33777 D_INPUT_3 POR2X1_5/CTRL 0.01fF
C33778 PAND2X1_798/B POR2X1_184/CTRL2 0.01fF
C33779 PAND2X1_115/Y POR2X1_416/B 0.01fF
C33780 POR2X1_409/Y INPUT_1 0.04fF
C33781 PAND2X1_82/CTRL POR2X1_294/A 0.01fF
C33782 POR2X1_305/O POR2X1_42/Y 0.05fF
C33783 PAND2X1_348/A PAND2X1_348/O 0.10fF
C33784 POR2X1_661/A POR2X1_807/A 0.03fF
C33785 POR2X1_263/Y POR2X1_263/O 0.01fF
C33786 POR2X1_678/O POR2X1_678/Y 0.01fF
C33787 PAND2X1_187/a_76_28# POR2X1_191/B 0.01fF
C33788 PAND2X1_618/CTRL POR2X1_29/A 0.01fF
C33789 PAND2X1_23/Y POR2X1_715/CTRL2 0.01fF
C33790 PAND2X1_853/m4_208_n4# PAND2X1_737/m4_208_n4# 0.05fF
C33791 POR2X1_548/A POR2X1_4/Y 0.05fF
C33792 POR2X1_407/A PAND2X1_56/A 0.03fF
C33793 POR2X1_355/B POR2X1_863/A 0.03fF
C33794 PAND2X1_20/A PAND2X1_85/a_76_28# 0.01fF
C33795 POR2X1_332/CTRL POR2X1_186/B 0.01fF
C33796 POR2X1_733/A POR2X1_717/B 0.08fF
C33797 PAND2X1_6/Y POR2X1_716/O 0.03fF
C33798 PAND2X1_93/B POR2X1_602/CTRL2 0.03fF
C33799 POR2X1_20/B POR2X1_432/O 0.02fF
C33800 PAND2X1_813/O POR2X1_266/A 0.02fF
C33801 POR2X1_326/A PAND2X1_533/CTRL 0.01fF
C33802 POR2X1_532/A POR2X1_555/CTRL2 0.01fF
C33803 POR2X1_655/A POR2X1_66/A 1.28fF
C33804 PAND2X1_834/CTRL2 PAND2X1_349/A 0.01fF
C33805 POR2X1_647/B POR2X1_590/A 0.03fF
C33806 POR2X1_493/A POR2X1_558/B 1.27fF
C33807 POR2X1_191/O POR2X1_568/Y 0.04fF
C33808 POR2X1_824/Y POR2X1_77/Y 0.08fF
C33809 POR2X1_66/Y POR2X1_838/B 0.00fF
C33810 POR2X1_416/B PAND2X1_803/Y 0.02fF
C33811 POR2X1_499/A POR2X1_777/B 0.05fF
C33812 PAND2X1_71/Y PAND2X1_527/CTRL 0.01fF
C33813 PAND2X1_96/B POR2X1_768/A 0.09fF
C33814 PAND2X1_216/B PAND2X1_850/Y 0.07fF
C33815 POR2X1_519/CTRL2 POR2X1_39/B 0.00fF
C33816 POR2X1_191/CTRL2 POR2X1_353/A 0.01fF
C33817 POR2X1_689/A POR2X1_689/a_16_28# 0.03fF
C33818 POR2X1_707/Y D_INPUT_4 0.02fF
C33819 POR2X1_721/CTRL2 POR2X1_383/Y 0.02fF
C33820 PAND2X1_606/m4_208_n4# POR2X1_37/Y 0.01fF
C33821 POR2X1_408/Y POR2X1_588/a_16_28# 0.03fF
C33822 POR2X1_260/B POR2X1_605/CTRL 0.01fF
C33823 POR2X1_9/Y POR2X1_55/Y 0.10fF
C33824 POR2X1_407/A POR2X1_661/A 0.07fF
C33825 PAND2X1_699/O VDD 0.00fF
C33826 POR2X1_119/Y POR2X1_265/Y 0.05fF
C33827 POR2X1_23/CTRL2 POR2X1_37/Y 0.01fF
C33828 POR2X1_16/CTRL2 POR2X1_73/Y 0.03fF
C33829 POR2X1_66/B POR2X1_84/A 0.03fF
C33830 POR2X1_78/B POR2X1_556/A 0.06fF
C33831 POR2X1_135/Y POR2X1_411/B 0.03fF
C33832 PAND2X1_432/O POR2X1_866/A 0.13fF
C33833 POR2X1_669/B POR2X1_667/Y 0.02fF
C33834 INPUT_3 PAND2X1_381/O 0.03fF
C33835 POR2X1_23/Y POR2X1_748/A 0.10fF
C33836 POR2X1_564/B POR2X1_568/B 0.03fF
C33837 POR2X1_153/CTRL POR2X1_416/B 0.01fF
C33838 PAND2X1_208/CTRL PAND2X1_124/Y 0.03fF
C33839 PAND2X1_6/Y POR2X1_457/Y 0.01fF
C33840 PAND2X1_560/B POR2X1_77/Y 3.34fF
C33841 PAND2X1_658/A POR2X1_67/Y 0.01fF
C33842 POR2X1_260/B PAND2X1_526/O 0.01fF
C33843 POR2X1_24/O POR2X1_48/A 0.06fF
C33844 POR2X1_98/a_76_344# PAND2X1_20/A 0.01fF
C33845 PAND2X1_96/B POR2X1_98/A 0.00fF
C33846 PAND2X1_620/Y POR2X1_422/a_76_344# 0.00fF
C33847 POR2X1_666/O PAND2X1_719/Y 0.21fF
C33848 POR2X1_275/CTRL POR2X1_275/A 0.01fF
C33849 POR2X1_850/B POR2X1_806/CTRL2 0.01fF
C33850 POR2X1_631/CTRL POR2X1_590/A 0.01fF
C33851 POR2X1_218/Y PAND2X1_41/B 0.01fF
C33852 PAND2X1_457/CTRL2 PAND2X1_464/B 0.03fF
C33853 PAND2X1_480/B PAND2X1_469/CTRL2 0.04fF
C33854 POR2X1_60/A PAND2X1_200/Y 0.01fF
C33855 POR2X1_72/B POR2X1_32/A 7.94fF
C33856 POR2X1_66/B POR2X1_285/Y 0.00fF
C33857 POR2X1_566/A POR2X1_446/B 0.05fF
C33858 POR2X1_718/O D_INPUT_0 0.01fF
C33859 POR2X1_83/B PAND2X1_208/CTRL 0.01fF
C33860 POR2X1_188/A POR2X1_285/Y 0.01fF
C33861 POR2X1_435/B POR2X1_294/B 0.01fF
C33862 POR2X1_856/B PAND2X1_627/O 0.02fF
C33863 POR2X1_695/Y PAND2X1_712/O 0.02fF
C33864 PAND2X1_626/CTRL2 POR2X1_852/B 0.06fF
C33865 PAND2X1_75/O POR2X1_724/A 0.01fF
C33866 POR2X1_818/Y POR2X1_415/O 0.01fF
C33867 PAND2X1_286/CTRL2 POR2X1_283/Y 0.01fF
C33868 PAND2X1_405/CTRL2 PAND2X1_737/B 0.01fF
C33869 POR2X1_840/B POR2X1_287/A 0.02fF
C33870 POR2X1_48/A PAND2X1_480/B 0.05fF
C33871 POR2X1_37/Y INPUT_0 0.21fF
C33872 POR2X1_23/Y PAND2X1_468/CTRL2 0.02fF
C33873 POR2X1_417/Y POR2X1_72/B 0.03fF
C33874 POR2X1_668/a_16_28# POR2X1_29/A 0.03fF
C33875 POR2X1_411/B POR2X1_816/A 0.06fF
C33876 POR2X1_447/A POR2X1_294/B 0.54fF
C33877 POR2X1_466/A POR2X1_724/CTRL 0.02fF
C33878 POR2X1_409/B PAND2X1_673/Y 0.07fF
C33879 POR2X1_54/Y POR2X1_790/B 0.06fF
C33880 POR2X1_439/CTRL PAND2X1_41/B 0.01fF
C33881 POR2X1_411/B D_INPUT_1 0.01fF
C33882 POR2X1_48/A POR2X1_754/A 0.06fF
C33883 PAND2X1_108/O POR2X1_646/Y 0.03fF
C33884 POR2X1_102/Y POR2X1_511/Y 0.03fF
C33885 POR2X1_490/Y PAND2X1_218/CTRL2 0.02fF
C33886 POR2X1_614/Y VDD 0.40fF
C33887 POR2X1_44/O POR2X1_748/A 0.07fF
C33888 POR2X1_558/CTRL POR2X1_260/B 0.01fF
C33889 PAND2X1_831/O PAND2X1_217/B 0.15fF
C33890 PAND2X1_92/O POR2X1_66/A 0.02fF
C33891 POR2X1_814/A PAND2X1_103/CTRL 0.01fF
C33892 POR2X1_487/m4_208_n4# POR2X1_488/m4_208_n4# 0.13fF
C33893 PAND2X1_65/B PAND2X1_46/CTRL2 0.01fF
C33894 POR2X1_130/A POR2X1_121/B 0.12fF
C33895 POR2X1_344/CTRL PAND2X1_65/B 0.01fF
C33896 PAND2X1_444/Y POR2X1_236/Y 0.01fF
C33897 POR2X1_220/Y PAND2X1_39/CTRL 0.02fF
C33898 POR2X1_83/B PAND2X1_520/O 0.01fF
C33899 POR2X1_477/B POR2X1_480/A 0.03fF
C33900 PAND2X1_48/B PAND2X1_277/a_16_344# 0.01fF
C33901 POR2X1_257/A POR2X1_426/Y 0.01fF
C33902 POR2X1_623/a_16_28# POR2X1_55/Y 0.02fF
C33903 POR2X1_848/A PAND2X1_6/A 0.07fF
C33904 POR2X1_343/A POR2X1_362/B 0.00fF
C33905 POR2X1_60/Y POR2X1_497/Y 0.02fF
C33906 POR2X1_411/B PAND2X1_854/A 0.02fF
C33907 PAND2X1_39/B POR2X1_307/A 0.03fF
C33908 PAND2X1_865/Y PAND2X1_860/A 0.01fF
C33909 PAND2X1_491/O POR2X1_260/B 0.02fF
C33910 POR2X1_718/A PAND2X1_90/Y 0.08fF
C33911 POR2X1_65/A POR2X1_107/O 0.01fF
C33912 POR2X1_288/A VDD 0.00fF
C33913 PAND2X1_48/B PAND2X1_594/a_56_28# 0.00fF
C33914 POR2X1_49/Y POR2X1_52/a_16_28# 0.00fF
C33915 POR2X1_188/A PAND2X1_108/a_16_344# 0.01fF
C33916 POR2X1_121/CTRL2 POR2X1_260/B 0.01fF
C33917 PAND2X1_56/Y POR2X1_269/O 0.02fF
C33918 PAND2X1_807/O PAND2X1_287/Y 0.09fF
C33919 PAND2X1_35/Y POR2X1_72/B 0.03fF
C33920 PAND2X1_810/A PAND2X1_288/A 0.03fF
C33921 POR2X1_319/A POR2X1_714/O 0.16fF
C33922 PAND2X1_22/m4_208_n4# PAND2X1_32/B 0.15fF
C33923 PAND2X1_3/A PAND2X1_69/A 0.06fF
C33924 POR2X1_669/B POR2X1_665/Y 0.07fF
C33925 POR2X1_496/CTRL2 POR2X1_789/B 0.00fF
C33926 PAND2X1_223/B PAND2X1_794/B 0.03fF
C33927 POR2X1_193/Y VDD 0.17fF
C33928 PAND2X1_73/CTRL2 POR2X1_294/B 0.15fF
C33929 POR2X1_840/CTRL D_INPUT_0 0.01fF
C33930 PAND2X1_404/Y PAND2X1_656/A 0.03fF
C33931 POR2X1_514/CTRL2 PAND2X1_20/A 0.01fF
C33932 POR2X1_68/A PAND2X1_603/a_76_28# 0.02fF
C33933 PAND2X1_94/A PAND2X1_39/B 0.16fF
C33934 POR2X1_81/m4_208_n4# PAND2X1_735/m4_208_n4# 0.13fF
C33935 PAND2X1_492/a_16_344# PAND2X1_65/B 0.01fF
C33936 POR2X1_687/A POR2X1_676/CTRL 0.01fF
C33937 POR2X1_499/a_16_28# POR2X1_576/Y 0.02fF
C33938 PAND2X1_863/B POR2X1_595/Y 0.01fF
C33939 POR2X1_466/A POR2X1_209/A 0.64fF
C33940 POR2X1_57/A D_INPUT_0 0.03fF
C33941 POR2X1_78/B POR2X1_400/A 0.12fF
C33942 POR2X1_284/B POR2X1_325/A 0.02fF
C33943 POR2X1_272/CTRL POR2X1_42/Y 0.01fF
C33944 POR2X1_630/CTRL POR2X1_510/Y 0.01fF
C33945 POR2X1_96/A PAND2X1_721/O 0.03fF
C33946 POR2X1_296/B POR2X1_702/A 0.05fF
C33947 POR2X1_79/Y PAND2X1_740/O 0.02fF
C33948 POR2X1_669/B PAND2X1_711/A 0.03fF
C33949 POR2X1_68/A POR2X1_866/CTRL 0.05fF
C33950 PAND2X1_419/a_76_28# PAND2X1_69/A 0.08fF
C33951 PAND2X1_821/CTRL2 PAND2X1_41/B 0.03fF
C33952 PAND2X1_620/Y POR2X1_615/Y 0.02fF
C33953 POR2X1_628/Y PAND2X1_507/CTRL2 0.00fF
C33954 PAND2X1_830/Y POR2X1_106/Y 0.02fF
C33955 PAND2X1_378/CTRL2 VDD 0.00fF
C33956 POR2X1_154/m4_208_n4# POR2X1_750/B 0.15fF
C33957 POR2X1_477/A POR2X1_186/Y 0.07fF
C33958 POR2X1_458/CTRL2 POR2X1_101/Y 0.08fF
C33959 POR2X1_287/B PAND2X1_371/O 0.02fF
C33960 PAND2X1_231/a_16_344# POR2X1_293/Y 0.02fF
C33961 POR2X1_294/CTRL2 POR2X1_507/A 0.03fF
C33962 POR2X1_406/Y INPUT_0 0.05fF
C33963 POR2X1_218/Y POR2X1_228/Y 0.12fF
C33964 PAND2X1_551/A POR2X1_40/Y 0.02fF
C33965 PAND2X1_20/A POR2X1_576/Y 0.01fF
C33966 PAND2X1_69/A POR2X1_720/a_76_344# 0.01fF
C33967 POR2X1_106/Y POR2X1_7/B 0.05fF
C33968 POR2X1_435/Y POR2X1_794/CTRL 0.03fF
C33969 PAND2X1_63/CTRL2 PAND2X1_63/B 0.01fF
C33970 INPUT_2 POR2X1_14/Y 0.00fF
C33971 PAND2X1_265/CTRL PAND2X1_32/B 0.01fF
C33972 PAND2X1_862/B PAND2X1_501/B 0.06fF
C33973 POR2X1_23/Y PAND2X1_574/CTRL2 0.06fF
C33974 POR2X1_60/A POR2X1_90/Y 0.08fF
C33975 PAND2X1_651/Y PAND2X1_465/CTRL2 0.00fF
C33976 PAND2X1_445/Y VDD 0.10fF
C33977 POR2X1_197/O POR2X1_244/B 0.01fF
C33978 POR2X1_567/B POR2X1_566/B 0.18fF
C33979 PAND2X1_734/B VDD 0.43fF
C33980 PAND2X1_317/Y PAND2X1_714/A 0.17fF
C33981 D_INPUT_0 POR2X1_229/Y 0.03fF
C33982 POR2X1_106/O PAND2X1_803/Y 0.00fF
C33983 PAND2X1_242/a_16_344# POR2X1_72/B 0.02fF
C33984 POR2X1_614/A PAND2X1_677/CTRL 0.01fF
C33985 POR2X1_567/B POR2X1_180/A 0.05fF
C33986 PAND2X1_209/A PAND2X1_161/CTRL 0.01fF
C33987 POR2X1_355/B POR2X1_798/m4_208_n4# 0.12fF
C33988 PAND2X1_74/CTRL POR2X1_702/A 0.00fF
C33989 PAND2X1_65/B PAND2X1_132/O 0.07fF
C33990 PAND2X1_658/B PAND2X1_185/O 0.16fF
C33991 D_INPUT_0 POR2X1_725/Y 0.07fF
C33992 POR2X1_556/A POR2X1_294/A 0.10fF
C33993 PAND2X1_92/CTRL2 INPUT_0 0.00fF
C33994 POR2X1_40/Y POR2X1_310/CTRL 0.01fF
C33995 POR2X1_596/A POR2X1_811/B 0.03fF
C33996 POR2X1_68/A PAND2X1_41/B 1.25fF
C33997 PAND2X1_437/CTRL PAND2X1_72/A 0.01fF
C33998 PAND2X1_615/a_16_344# PAND2X1_58/A 0.02fF
C33999 POR2X1_558/B POR2X1_276/Y 0.05fF
C34000 PAND2X1_651/Y POR2X1_72/B 0.08fF
C34001 POR2X1_383/A POR2X1_269/O 0.02fF
C34002 POR2X1_207/A POR2X1_740/Y 0.05fF
C34003 POR2X1_464/CTRL2 PAND2X1_55/Y 0.01fF
C34004 POR2X1_655/a_16_28# POR2X1_711/Y 0.09fF
C34005 PAND2X1_61/Y POR2X1_521/CTRL 0.01fF
C34006 PAND2X1_580/B POR2X1_7/B 0.03fF
C34007 PAND2X1_59/B POR2X1_260/A 0.04fF
C34008 PAND2X1_252/CTRL POR2X1_750/B 0.32fF
C34009 POR2X1_19/a_56_344# POR2X1_4/Y 0.01fF
C34010 POR2X1_832/A POR2X1_78/A 0.04fF
C34011 POR2X1_697/Y POR2X1_236/Y 0.04fF
C34012 POR2X1_257/A POR2X1_320/CTRL2 0.00fF
C34013 INPUT_0 POR2X1_293/Y 1.52fF
C34014 PAND2X1_828/CTRL POR2X1_599/A 0.01fF
C34015 POR2X1_49/Y PAND2X1_653/Y 0.09fF
C34016 POR2X1_654/B POR2X1_649/CTRL2 0.04fF
C34017 PAND2X1_249/O POR2X1_591/Y 0.05fF
C34018 PAND2X1_23/Y PAND2X1_293/CTRL2 0.00fF
C34019 POR2X1_654/B PAND2X1_69/A 0.07fF
C34020 INPUT_1 POR2X1_817/a_16_28# 0.03fF
C34021 POR2X1_288/A PAND2X1_32/B 0.06fF
C34022 POR2X1_447/B POR2X1_776/A 0.03fF
C34023 POR2X1_41/B POR2X1_13/a_16_28# 0.01fF
C34024 POR2X1_566/A PAND2X1_441/CTRL2 0.06fF
C34025 PAND2X1_274/a_76_28# PAND2X1_480/B 0.03fF
C34026 POR2X1_814/B POR2X1_576/Y 0.57fF
C34027 POR2X1_789/Y VDD 0.10fF
C34028 POR2X1_376/B POR2X1_816/A 0.03fF
C34029 POR2X1_394/Y PAND2X1_656/A 0.00fF
C34030 PAND2X1_262/O PAND2X1_69/A 0.17fF
C34031 POR2X1_278/Y POR2X1_55/Y 0.03fF
C34032 PAND2X1_434/CTRL2 POR2X1_83/B -0.00fF
C34033 PAND2X1_280/CTRL2 PAND2X1_55/Y 0.01fF
C34034 POR2X1_186/Y PAND2X1_747/CTRL 0.28fF
C34035 POR2X1_29/A PAND2X1_133/O 0.02fF
C34036 POR2X1_40/Y PAND2X1_338/B 0.03fF
C34037 POR2X1_111/Y D_INPUT_0 0.01fF
C34038 POR2X1_383/A POR2X1_634/A 0.18fF
C34039 POR2X1_39/O POR2X1_38/Y 0.20fF
C34040 PAND2X1_48/B PAND2X1_751/CTRL 0.00fF
C34041 PAND2X1_56/Y POR2X1_130/A 0.04fF
C34042 POR2X1_416/B PAND2X1_780/CTRL2 0.04fF
C34043 PAND2X1_69/A POR2X1_5/Y 0.06fF
C34044 POR2X1_367/O POR2X1_364/A 0.08fF
C34045 POR2X1_272/CTRL2 PAND2X1_349/A 0.01fF
C34046 POR2X1_68/A POR2X1_402/B 0.02fF
C34047 POR2X1_13/A POR2X1_45/Y 0.07fF
C34048 PAND2X1_341/A POR2X1_5/Y 0.03fF
C34049 POR2X1_102/Y PAND2X1_861/CTRL 0.01fF
C34050 POR2X1_730/B VDD 0.04fF
C34051 POR2X1_43/B PAND2X1_636/O 0.03fF
C34052 POR2X1_566/A POR2X1_795/B 0.10fF
C34053 PAND2X1_56/Y POR2X1_566/A 0.03fF
C34054 PAND2X1_94/A PAND2X1_20/A 0.19fF
C34055 PAND2X1_55/Y POR2X1_465/B 0.03fF
C34056 PAND2X1_69/A POR2X1_778/O 0.02fF
C34057 POR2X1_567/A POR2X1_447/A 0.21fF
C34058 POR2X1_508/CTRL2 POR2X1_579/Y 0.01fF
C34059 PAND2X1_65/B POR2X1_775/a_16_28# 0.02fF
C34060 POR2X1_274/Y PAND2X1_60/B 0.03fF
C34061 POR2X1_93/A POR2X1_5/Y 3.30fF
C34062 POR2X1_153/a_16_28# POR2X1_48/A 0.00fF
C34063 POR2X1_416/Y POR2X1_411/CTRL2 0.01fF
C34064 PAND2X1_473/O PAND2X1_473/B 0.01fF
C34065 POR2X1_123/A POR2X1_734/A 1.50fF
C34066 POR2X1_614/A POR2X1_155/O 0.18fF
C34067 POR2X1_814/B POR2X1_360/O 0.01fF
C34068 POR2X1_5/Y POR2X1_91/Y 0.39fF
C34069 PAND2X1_57/B PAND2X1_69/CTRL2 0.01fF
C34070 POR2X1_143/CTRL PAND2X1_6/A 0.03fF
C34071 POR2X1_731/O VDD 0.00fF
C34072 POR2X1_330/Y POR2X1_598/CTRL 0.30fF
C34073 POR2X1_833/CTRL POR2X1_294/B 0.01fF
C34074 POR2X1_616/Y POR2X1_818/Y 0.59fF
C34075 POR2X1_119/Y PAND2X1_776/Y 0.32fF
C34076 POR2X1_614/A POR2X1_502/A 0.22fF
C34077 POR2X1_567/A POR2X1_629/O -0.01fF
C34078 POR2X1_43/B POR2X1_58/Y 0.01fF
C34079 POR2X1_779/A POR2X1_708/B 0.00fF
C34080 PAND2X1_57/B POR2X1_705/O 0.01fF
C34081 POR2X1_780/CTRL2 POR2X1_260/A 0.01fF
C34082 POR2X1_254/Y PAND2X1_96/B 0.07fF
C34083 POR2X1_234/CTRL2 POR2X1_293/Y 0.00fF
C34084 POR2X1_447/B POR2X1_856/B 0.03fF
C34085 PAND2X1_104/O POR2X1_673/Y 0.01fF
C34086 POR2X1_7/B PAND2X1_337/A 0.01fF
C34087 PAND2X1_494/CTRL POR2X1_294/B 0.05fF
C34088 POR2X1_542/B POR2X1_220/Y 0.03fF
C34089 POR2X1_102/Y POR2X1_129/Y 0.13fF
C34090 POR2X1_52/A POR2X1_816/A 0.07fF
C34091 POR2X1_566/A POR2X1_336/O 0.01fF
C34092 PAND2X1_707/Y PAND2X1_705/CTRL 0.01fF
C34093 POR2X1_502/A POR2X1_38/B 0.10fF
C34094 PAND2X1_676/CTRL PAND2X1_735/Y 0.03fF
C34095 PAND2X1_492/CTRL2 POR2X1_123/A 0.01fF
C34096 PAND2X1_90/Y POR2X1_725/Y 0.10fF
C34097 POR2X1_52/A D_INPUT_1 0.03fF
C34098 PAND2X1_90/A PAND2X1_6/A 0.21fF
C34099 PAND2X1_362/A PAND2X1_354/Y 0.01fF
C34100 PAND2X1_498/a_76_28# POR2X1_733/A 0.02fF
C34101 POR2X1_65/A PAND2X1_264/O 0.01fF
C34102 PAND2X1_94/A POR2X1_814/B 0.58fF
C34103 PAND2X1_521/O INPUT_0 0.04fF
C34104 POR2X1_614/A POR2X1_464/Y 0.73fF
C34105 POR2X1_498/O POR2X1_38/Y 0.01fF
C34106 POR2X1_78/B PAND2X1_393/O 0.04fF
C34107 POR2X1_193/CTRL2 POR2X1_631/B 0.04fF
C34108 POR2X1_68/A POR2X1_130/Y 0.10fF
C34109 POR2X1_408/Y INPUT_0 0.10fF
C34110 POR2X1_7/B PAND2X1_347/O 0.03fF
C34111 POR2X1_13/A POR2X1_396/Y 0.03fF
C34112 PAND2X1_278/CTRL2 POR2X1_559/A 0.48fF
C34113 POR2X1_283/A PAND2X1_730/B 0.03fF
C34114 POR2X1_327/Y POR2X1_330/Y 0.09fF
C34115 PAND2X1_436/A POR2X1_129/Y 0.32fF
C34116 POR2X1_383/A POR2X1_130/A 0.41fF
C34117 POR2X1_332/B POR2X1_510/Y 0.03fF
C34118 PAND2X1_661/Y VDD 0.20fF
C34119 POR2X1_596/A POR2X1_783/B 0.02fF
C34120 POR2X1_809/A POR2X1_866/O 0.01fF
C34121 PAND2X1_659/Y POR2X1_102/Y 0.10fF
C34122 PAND2X1_96/B POR2X1_575/B 0.01fF
C34123 POR2X1_832/Y POR2X1_711/Y 0.02fF
C34124 PAND2X1_23/Y POR2X1_68/B 0.13fF
C34125 POR2X1_566/A POR2X1_383/A 0.10fF
C34126 POR2X1_68/A PAND2X1_72/CTRL 0.00fF
C34127 POR2X1_121/CTRL2 PAND2X1_55/Y 0.03fF
C34128 POR2X1_856/B POR2X1_510/O 0.28fF
C34129 PAND2X1_221/O PAND2X1_730/A 0.00fF
C34130 PAND2X1_661/B POR2X1_45/Y 0.03fF
C34131 POR2X1_451/A POR2X1_635/CTRL2 0.01fF
C34132 POR2X1_635/B POR2X1_635/CTRL 0.01fF
C34133 POR2X1_62/Y PAND2X1_459/O 0.12fF
C34134 POR2X1_154/O POR2X1_855/B 0.01fF
C34135 POR2X1_566/A PAND2X1_253/CTRL2 0.32fF
C34136 PAND2X1_499/Y PAND2X1_861/a_16_344# 0.01fF
C34137 POR2X1_51/A POR2X1_51/B 0.11fF
C34138 POR2X1_750/B POR2X1_652/A 0.03fF
C34139 PAND2X1_465/B POR2X1_387/Y 0.03fF
C34140 PAND2X1_830/Y PAND2X1_349/A 0.04fF
C34141 POR2X1_96/O POR2X1_236/Y 0.02fF
C34142 POR2X1_808/A PAND2X1_48/A 0.14fF
C34143 POR2X1_213/CTRL POR2X1_532/A 0.01fF
C34144 PAND2X1_56/Y POR2X1_573/A 0.05fF
C34145 POR2X1_853/A POR2X1_578/CTRL 0.01fF
C34146 POR2X1_789/B VDD 0.00fF
C34147 PAND2X1_93/CTRL PAND2X1_88/Y 0.01fF
C34148 POR2X1_517/CTRL2 POR2X1_83/B 0.00fF
C34149 PAND2X1_96/B POR2X1_574/O 0.01fF
C34150 POR2X1_394/A PAND2X1_738/O 0.04fF
C34151 PAND2X1_63/B POR2X1_7/B 0.03fF
C34152 PAND2X1_90/Y POR2X1_559/A 0.04fF
C34153 PAND2X1_69/A POR2X1_705/CTRL 0.01fF
C34154 D_INPUT_0 PAND2X1_339/CTRL 0.07fF
C34155 POR2X1_394/O VDD 0.00fF
C34156 POR2X1_536/O POR2X1_13/A 0.02fF
C34157 POR2X1_334/A PAND2X1_85/Y 0.00fF
C34158 POR2X1_96/A PAND2X1_737/B 0.01fF
C34159 POR2X1_72/B PAND2X1_199/CTRL2 0.03fF
C34160 PAND2X1_831/m4_208_n4# POR2X1_394/A 0.06fF
C34161 POR2X1_327/Y POR2X1_302/CTRL 0.01fF
C34162 POR2X1_807/A POR2X1_737/A 0.03fF
C34163 POR2X1_804/A PAND2X1_311/O 0.02fF
C34164 POR2X1_96/A PAND2X1_216/B 0.03fF
C34165 POR2X1_389/O POR2X1_725/Y 0.02fF
C34166 POR2X1_68/A POR2X1_228/Y 0.05fF
C34167 PAND2X1_90/A POR2X1_101/Y 0.12fF
C34168 PAND2X1_531/CTRL POR2X1_547/B 0.00fF
C34169 POR2X1_406/CTRL PAND2X1_737/B 0.01fF
C34170 POR2X1_57/A POR2X1_528/a_16_28# 0.03fF
C34171 POR2X1_78/B POR2X1_398/O 0.02fF
C34172 POR2X1_550/A POR2X1_68/A 0.03fF
C34173 PAND2X1_275/O POR2X1_569/A 0.08fF
C34174 POR2X1_539/CTRL2 POR2X1_741/Y 0.00fF
C34175 POR2X1_220/B POR2X1_161/O 0.02fF
C34176 POR2X1_614/A PAND2X1_158/CTRL2 0.00fF
C34177 PAND2X1_484/CTRL PAND2X1_57/B 0.02fF
C34178 PAND2X1_810/a_56_28# POR2X1_7/B 0.00fF
C34179 POR2X1_383/A POR2X1_844/B 0.03fF
C34180 PAND2X1_547/CTRL POR2X1_527/Y 0.01fF
C34181 POR2X1_299/O POR2X1_91/Y 0.06fF
C34182 POR2X1_400/A POR2X1_294/A 0.11fF
C34183 D_INPUT_1 POR2X1_550/Y 0.03fF
C34184 POR2X1_156/B POR2X1_162/Y 0.00fF
C34185 INPUT_1 POR2X1_32/a_56_344# 0.00fF
C34186 POR2X1_499/A POR2X1_814/A 0.03fF
C34187 PAND2X1_390/Y POR2X1_589/a_56_344# 0.00fF
C34188 POR2X1_110/CTRL POR2X1_13/A 0.01fF
C34189 POR2X1_96/A PAND2X1_359/Y 0.03fF
C34190 PAND2X1_41/B POR2X1_169/A 0.03fF
C34191 POR2X1_71/O POR2X1_293/Y 0.05fF
C34192 POR2X1_860/CTRL POR2X1_218/A 0.02fF
C34193 PAND2X1_6/Y PAND2X1_300/CTRL 0.01fF
C34194 POR2X1_679/B POR2X1_816/A 0.00fF
C34195 D_GATE_222 POR2X1_260/A 0.05fF
C34196 PAND2X1_215/B PAND2X1_853/B 0.07fF
C34197 POR2X1_208/Y POR2X1_215/A 0.04fF
C34198 PAND2X1_649/A PAND2X1_688/CTRL2 0.01fF
C34199 PAND2X1_139/CTRL2 PAND2X1_140/Y 0.03fF
C34200 POR2X1_383/A POR2X1_573/A 0.03fF
C34201 PAND2X1_615/CTRL PAND2X1_63/B 0.01fF
C34202 POR2X1_832/A POR2X1_513/CTRL2 0.03fF
C34203 POR2X1_72/B POR2X1_387/CTRL 0.01fF
C34204 POR2X1_508/A POR2X1_192/Y 0.05fF
C34205 POR2X1_580/a_76_344# POR2X1_191/Y 0.02fF
C34206 POR2X1_54/Y POR2X1_848/CTRL 0.01fF
C34207 POR2X1_110/CTRL2 POR2X1_293/Y 0.01fF
C34208 POR2X1_54/Y PAND2X1_87/CTRL 0.05fF
C34209 POR2X1_164/Y POR2X1_73/Y 0.03fF
C34210 PAND2X1_542/CTRL PAND2X1_552/B 0.01fF
C34211 PAND2X1_793/Y POR2X1_767/O 0.02fF
C34212 D_INPUT_7 PAND2X1_581/O 0.05fF
C34213 POR2X1_55/Y PAND2X1_357/O 0.01fF
C34214 PAND2X1_23/Y POR2X1_326/A 0.00fF
C34215 PAND2X1_63/B PAND2X1_60/B 0.10fF
C34216 PAND2X1_724/B PAND2X1_357/a_16_344# 0.03fF
C34217 POR2X1_569/a_16_28# POR2X1_568/B 0.06fF
C34218 POR2X1_557/A PAND2X1_79/Y 0.03fF
C34219 POR2X1_62/Y PAND2X1_341/O 0.05fF
C34220 POR2X1_684/Y POR2X1_7/B 0.04fF
C34221 POR2X1_541/O POR2X1_456/B 0.01fF
C34222 PAND2X1_312/CTRL2 POR2X1_703/A 0.10fF
C34223 POR2X1_7/A PAND2X1_154/O 0.01fF
C34224 POR2X1_397/Y POR2X1_39/B 0.01fF
C34225 PAND2X1_671/a_56_28# INPUT_2 0.00fF
C34226 POR2X1_116/A POR2X1_556/A 3.77fF
C34227 PAND2X1_560/B POR2X1_52/Y 0.03fF
C34228 POR2X1_600/O POR2X1_600/Y 0.01fF
C34229 POR2X1_702/CTRL2 POR2X1_260/A 0.01fF
C34230 POR2X1_81/A PAND2X1_793/Y 0.03fF
C34231 PAND2X1_96/B PAND2X1_184/a_76_28# 0.01fF
C34232 POR2X1_192/Y POR2X1_568/B 0.12fF
C34233 POR2X1_407/A POR2X1_737/A 0.03fF
C34234 POR2X1_68/A PAND2X1_482/a_16_344# 0.05fF
C34235 POR2X1_548/CTRL2 PAND2X1_52/B 0.32fF
C34236 PAND2X1_499/Y PAND2X1_861/B 0.06fF
C34237 POR2X1_319/a_16_28# POR2X1_192/B 0.04fF
C34238 POR2X1_652/CTRL POR2X1_652/A 0.00fF
C34239 INPUT_3 POR2X1_411/B 0.18fF
C34240 POR2X1_569/Y POR2X1_854/B 0.03fF
C34241 PAND2X1_569/B PAND2X1_374/O 0.00fF
C34242 POR2X1_560/Y POR2X1_844/B 0.01fF
C34243 POR2X1_789/a_16_28# POR2X1_789/B 0.03fF
C34244 PAND2X1_794/B POR2X1_385/Y 0.05fF
C34245 POR2X1_16/A POR2X1_283/A 0.07fF
C34246 PAND2X1_216/B POR2X1_7/A 0.03fF
C34247 POR2X1_730/Y POR2X1_727/CTRL 0.01fF
C34248 POR2X1_257/A POR2X1_20/B 0.46fF
C34249 PAND2X1_39/B PAND2X1_43/CTRL2 0.01fF
C34250 PAND2X1_352/CTRL2 PAND2X1_357/Y 0.01fF
C34251 POR2X1_497/Y PAND2X1_351/A 0.00fF
C34252 POR2X1_23/Y POR2X1_441/a_16_28# 0.02fF
C34253 POR2X1_614/A POR2X1_188/Y 0.03fF
C34254 POR2X1_815/a_16_28# POR2X1_815/A 0.05fF
C34255 POR2X1_276/Y POR2X1_362/A 1.12fF
C34256 POR2X1_57/A PAND2X1_138/CTRL2 0.01fF
C34257 PAND2X1_763/O PAND2X1_52/B 0.01fF
C34258 PAND2X1_69/A PAND2X1_396/CTRL2 0.03fF
C34259 POR2X1_307/Y POR2X1_711/Y 0.04fF
C34260 PAND2X1_501/CTRL2 POR2X1_494/Y 0.00fF
C34261 POR2X1_344/Y POR2X1_383/A 0.04fF
C34262 POR2X1_416/B PAND2X1_668/O 0.04fF
C34263 POR2X1_16/A PAND2X1_100/O 0.00fF
C34264 POR2X1_130/O POR2X1_141/A 0.01fF
C34265 PAND2X1_23/Y POR2X1_374/a_16_28# 0.02fF
C34266 POR2X1_222/A POR2X1_186/B 0.03fF
C34267 POR2X1_456/B POR2X1_675/Y 0.03fF
C34268 PAND2X1_787/A PAND2X1_716/B 0.03fF
C34269 PAND2X1_508/Y PAND2X1_549/B 0.03fF
C34270 POR2X1_416/B POR2X1_42/Y 3.91fF
C34271 PAND2X1_653/Y PAND2X1_737/m4_208_n4# 0.21fF
C34272 POR2X1_548/A POR2X1_620/B 0.12fF
C34273 PAND2X1_393/O POR2X1_294/A 0.15fF
C34274 POR2X1_180/O POR2X1_180/A 0.03fF
C34275 POR2X1_544/B POR2X1_456/B 0.03fF
C34276 POR2X1_452/Y POR2X1_809/O 0.01fF
C34277 PAND2X1_138/O POR2X1_7/A 0.15fF
C34278 POR2X1_416/B POR2X1_745/CTRL 0.01fF
C34279 POR2X1_338/a_16_28# POR2X1_334/Y 0.08fF
C34280 POR2X1_863/A POR2X1_570/CTRL2 0.01fF
C34281 POR2X1_776/B POR2X1_568/A 0.03fF
C34282 PAND2X1_242/Y INPUT_0 0.17fF
C34283 POR2X1_657/Y POR2X1_218/Y 0.08fF
C34284 PAND2X1_635/Y POR2X1_763/A 0.06fF
C34285 POR2X1_9/Y POR2X1_625/CTRL2 0.01fF
C34286 POR2X1_823/CTRL POR2X1_77/Y 0.01fF
C34287 PAND2X1_276/O POR2X1_677/Y 0.04fF
C34288 POR2X1_145/Y PAND2X1_797/Y 0.83fF
C34289 POR2X1_411/B POR2X1_432/CTRL2 0.01fF
C34290 POR2X1_677/Y POR2X1_511/Y 0.00fF
C34291 POR2X1_305/CTRL PAND2X1_651/Y 0.00fF
C34292 PAND2X1_717/A POR2X1_40/Y 0.01fF
C34293 POR2X1_610/Y POR2X1_610/a_16_28# 0.03fF
C34294 PAND2X1_64/CTRL PAND2X1_26/A 0.01fF
C34295 PAND2X1_266/O POR2X1_40/Y 0.04fF
C34296 PAND2X1_621/CTRL2 POR2X1_616/Y 0.01fF
C34297 POR2X1_772/CTRL2 POR2X1_294/A 0.03fF
C34298 POR2X1_647/B POR2X1_66/A 0.03fF
C34299 POR2X1_394/A PAND2X1_708/CTRL 0.01fF
C34300 POR2X1_814/B POR2X1_621/O 0.03fF
C34301 POR2X1_116/A POR2X1_474/O 0.00fF
C34302 POR2X1_707/B PAND2X1_425/Y 0.01fF
C34303 PAND2X1_518/CTRL PAND2X1_52/B 0.02fF
C34304 PAND2X1_482/O POR2X1_186/B 0.01fF
C34305 PAND2X1_39/B POR2X1_287/O 0.01fF
C34306 POR2X1_169/A POR2X1_704/O 0.02fF
C34307 POR2X1_557/B POR2X1_768/Y 0.01fF
C34308 PAND2X1_60/B POR2X1_342/A 0.00fF
C34309 POR2X1_114/a_56_344# POR2X1_717/B 0.00fF
C34310 POR2X1_568/B POR2X1_568/Y 0.04fF
C34311 POR2X1_577/CTRL2 POR2X1_568/A 0.03fF
C34312 POR2X1_23/Y POR2X1_263/Y 0.03fF
C34313 POR2X1_16/O POR2X1_42/Y 0.01fF
C34314 POR2X1_827/Y POR2X1_669/B 0.01fF
C34315 POR2X1_294/A POR2X1_398/O 0.18fF
C34316 POR2X1_811/CTRL2 D_INPUT_0 0.00fF
C34317 POR2X1_422/CTRL2 POR2X1_422/Y 0.01fF
C34318 POR2X1_49/Y POR2X1_20/B 0.20fF
C34319 POR2X1_859/O POR2X1_734/A 0.02fF
C34320 POR2X1_130/A POR2X1_648/Y 2.23fF
C34321 POR2X1_475/CTRL2 POR2X1_288/A 0.00fF
C34322 POR2X1_48/A POR2X1_484/O 0.02fF
C34323 PAND2X1_48/A PAND2X1_692/CTRL 0.01fF
C34324 POR2X1_612/Y POR2X1_414/O 0.05fF
C34325 POR2X1_329/A PAND2X1_735/Y 0.07fF
C34326 PAND2X1_797/Y POR2X1_394/A 1.29fF
C34327 PAND2X1_640/B POR2X1_32/A 0.20fF
C34328 PAND2X1_52/B POR2X1_854/B 0.34fF
C34329 PAND2X1_497/O PAND2X1_58/A 0.02fF
C34330 POR2X1_612/Y POR2X1_607/CTRL2 0.05fF
C34331 POR2X1_212/B POR2X1_854/B 0.05fF
C34332 POR2X1_376/B INPUT_3 0.03fF
C34333 POR2X1_447/B POR2X1_191/Y 0.05fF
C34334 PAND2X1_269/CTRL POR2X1_55/Y 0.00fF
C34335 POR2X1_846/A POR2X1_805/A 0.01fF
C34336 POR2X1_102/Y POR2X1_37/Y 1.79fF
C34337 POR2X1_657/O POR2X1_218/Y 0.01fF
C34338 POR2X1_485/a_16_28# POR2X1_73/Y 0.03fF
C34339 POR2X1_632/O POR2X1_750/B 0.02fF
C34340 PAND2X1_20/A POR2X1_637/CTRL2 0.00fF
C34341 POR2X1_705/B POR2X1_546/A 0.45fF
C34342 PAND2X1_96/B POR2X1_643/CTRL2 0.01fF
C34343 POR2X1_811/B D_INPUT_0 0.00fF
C34344 POR2X1_23/Y PAND2X1_658/CTRL2 0.01fF
C34345 PAND2X1_796/B PAND2X1_778/CTRL 0.00fF
C34346 PAND2X1_717/A PAND2X1_303/a_16_344# 0.02fF
C34347 POR2X1_428/Y POR2X1_376/B 0.02fF
C34348 POR2X1_811/B POR2X1_811/A 0.03fF
C34349 PAND2X1_415/CTRL2 VDD 0.00fF
C34350 PAND2X1_18/B D_INPUT_4 0.17fF
C34351 POR2X1_852/a_16_28# POR2X1_776/A 0.03fF
C34352 PAND2X1_659/Y POR2X1_761/A 0.03fF
C34353 PAND2X1_9/Y PAND2X1_734/B 0.25fF
C34354 POR2X1_326/A POR2X1_711/Y 0.07fF
C34355 POR2X1_376/B POR2X1_93/Y 0.11fF
C34356 POR2X1_123/CTRL2 POR2X1_556/A 0.01fF
C34357 PAND2X1_58/CTRL POR2X1_202/A 0.05fF
C34358 PAND2X1_20/A PAND2X1_11/Y 0.02fF
C34359 POR2X1_272/CTRL2 POR2X1_32/A 0.02fF
C34360 POR2X1_855/m4_208_n4# PAND2X1_829/m4_208_n4# 0.13fF
C34361 PAND2X1_20/A POR2X1_606/Y 0.06fF
C34362 POR2X1_52/A INPUT_3 0.15fF
C34363 POR2X1_33/O POR2X1_33/B 0.04fF
C34364 PAND2X1_600/a_16_344# POR2X1_814/B 0.01fF
C34365 POR2X1_69/O PAND2X1_58/A 0.01fF
C34366 POR2X1_56/CTRL POR2X1_423/Y 0.02fF
C34367 POR2X1_14/Y POR2X1_69/A 0.74fF
C34368 PAND2X1_431/O POR2X1_480/A 0.12fF
C34369 D_INPUT_0 PAND2X1_525/O 0.03fF
C34370 POR2X1_124/a_16_28# POR2X1_556/A 0.02fF
C34371 PAND2X1_220/Y PAND2X1_220/A 0.02fF
C34372 PAND2X1_48/B POR2X1_663/B 6.39fF
C34373 POR2X1_376/B POR2X1_432/CTRL2 0.08fF
C34374 POR2X1_634/A POR2X1_634/O 0.02fF
C34375 PAND2X1_75/CTRL2 POR2X1_318/A 0.01fF
C34376 POR2X1_43/B POR2X1_150/Y 0.07fF
C34377 POR2X1_15/CTRL PAND2X1_206/B 0.00fF
C34378 POR2X1_77/Y PAND2X1_352/B 0.01fF
C34379 POR2X1_106/CTRL POR2X1_106/Y 0.01fF
C34380 PAND2X1_219/A PAND2X1_733/CTRL 0.01fF
C34381 PAND2X1_675/A POR2X1_411/B 0.03fF
C34382 POR2X1_77/a_16_28# POR2X1_13/A 0.03fF
C34383 PAND2X1_240/a_76_28# D_INPUT_0 0.02fF
C34384 PAND2X1_58/A PAND2X1_41/B 0.10fF
C34385 PAND2X1_469/B POR2X1_411/B 0.03fF
C34386 PAND2X1_23/Y PAND2X1_826/CTRL 0.01fF
C34387 POR2X1_774/Y POR2X1_121/B 0.03fF
C34388 D_INPUT_0 PAND2X1_84/Y 0.03fF
C34389 POR2X1_294/Y PAND2X1_58/O 0.01fF
C34390 POR2X1_814/B POR2X1_606/Y 0.01fF
C34391 POR2X1_670/O POR2X1_102/Y 0.01fF
C34392 PAND2X1_487/CTRL POR2X1_294/B 0.04fF
C34393 PAND2X1_475/O PAND2X1_217/B 0.04fF
C34394 POR2X1_709/A PAND2X1_411/CTRL 0.02fF
C34395 PAND2X1_404/Y PAND2X1_197/CTRL 0.00fF
C34396 POR2X1_192/B POR2X1_568/A 0.10fF
C34397 POR2X1_407/A PAND2X1_761/CTRL 0.01fF
C34398 POR2X1_52/A POR2X1_93/Y 1.95fF
C34399 PAND2X1_203/CTRL2 POR2X1_816/A 0.03fF
C34400 POR2X1_72/B PAND2X1_731/B 0.02fF
C34401 POR2X1_68/A PAND2X1_826/CTRL2 0.05fF
C34402 POR2X1_811/B PAND2X1_90/Y 0.07fF
C34403 PAND2X1_23/Y POR2X1_458/CTRL2 0.01fF
C34404 POR2X1_260/B PAND2X1_385/O 0.01fF
C34405 POR2X1_83/B POR2X1_697/O 0.01fF
C34406 POR2X1_23/Y PAND2X1_215/B 0.03fF
C34407 POR2X1_677/Y POR2X1_129/Y 0.18fF
C34408 PAND2X1_677/CTRL2 PAND2X1_90/Y 0.03fF
C34409 POR2X1_423/Y PAND2X1_541/O 0.02fF
C34410 POR2X1_16/A POR2X1_399/Y 0.00fF
C34411 PAND2X1_16/a_76_28# POR2X1_630/A 0.04fF
C34412 POR2X1_164/a_16_28# POR2X1_20/B 0.02fF
C34413 POR2X1_364/A POR2X1_212/A 0.03fF
C34414 PAND2X1_673/a_16_344# POR2X1_14/Y 0.05fF
C34415 POR2X1_68/A POR2X1_454/A 0.02fF
C34416 POR2X1_493/A POR2X1_572/B 0.18fF
C34417 POR2X1_406/Y POR2X1_102/Y 0.15fF
C34418 PAND2X1_443/CTRL2 POR2X1_90/Y 0.00fF
C34419 POR2X1_311/Y POR2X1_481/A 1.16fF
C34420 PAND2X1_326/B POR2X1_167/Y 0.00fF
C34421 POR2X1_502/A POR2X1_590/A 0.09fF
C34422 D_INPUT_0 POR2X1_783/B 0.02fF
C34423 PAND2X1_58/A POR2X1_402/B 0.00fF
C34424 POR2X1_9/Y POR2X1_129/Y 0.07fF
C34425 PAND2X1_392/CTRL POR2X1_55/Y 0.00fF
C34426 POR2X1_811/A POR2X1_783/B 0.02fF
C34427 POR2X1_60/A INPUT_0 0.35fF
C34428 POR2X1_83/B POR2X1_88/Y 0.03fF
C34429 POR2X1_821/a_16_28# POR2X1_669/B 0.02fF
C34430 PAND2X1_236/CTRL2 POR2X1_94/A 0.03fF
C34431 POR2X1_274/A POR2X1_513/Y 11.88fF
C34432 POR2X1_634/A INPUT_0 0.05fF
C34433 POR2X1_309/CTRL2 POR2X1_293/Y 0.01fF
C34434 POR2X1_32/A POR2X1_7/B 0.14fF
C34435 PAND2X1_220/Y POR2X1_106/Y 0.03fF
C34436 PAND2X1_777/O POR2X1_55/Y 0.01fF
C34437 POR2X1_810/O POR2X1_636/B 0.01fF
C34438 POR2X1_760/A PAND2X1_737/B 0.03fF
C34439 POR2X1_293/O POR2X1_5/Y 0.05fF
C34440 POR2X1_666/Y PAND2X1_719/CTRL2 0.01fF
C34441 PAND2X1_42/CTRL2 POR2X1_547/B 0.00fF
C34442 POR2X1_23/Y PAND2X1_6/A 0.00fF
C34443 PAND2X1_216/B POR2X1_760/A 0.01fF
C34444 POR2X1_54/Y PAND2X1_521/a_16_344# 0.06fF
C34445 PAND2X1_299/CTRL2 VDD 0.00fF
C34446 POR2X1_660/CTRL PAND2X1_55/Y 0.01fF
C34447 POR2X1_102/Y POR2X1_293/Y 0.34fF
C34448 POR2X1_324/B VDD 0.14fF
C34449 POR2X1_66/A POR2X1_340/a_16_28# 0.03fF
C34450 POR2X1_65/A POR2X1_760/O 0.17fF
C34451 PAND2X1_42/CTRL VDD 0.00fF
C34452 POR2X1_566/A PAND2X1_230/m4_208_n4# 0.05fF
C34453 PAND2X1_659/A PAND2X1_659/O 0.01fF
C34454 PAND2X1_845/CTRL POR2X1_37/Y 0.01fF
C34455 POR2X1_8/Y PAND2X1_35/a_76_28# 0.01fF
C34456 POR2X1_118/CTRL POR2X1_37/Y 0.06fF
C34457 POR2X1_65/A PAND2X1_362/B 0.03fF
C34458 PAND2X1_220/Y PAND2X1_580/B 0.01fF
C34459 PAND2X1_217/B POR2X1_498/CTRL 0.01fF
C34460 POR2X1_244/B PAND2X1_7/Y 0.67fF
C34461 POR2X1_41/B POR2X1_40/Y 1.07fF
C34462 PAND2X1_340/B POR2X1_408/Y 2.12fF
C34463 POR2X1_585/Y POR2X1_790/B 0.00fF
C34464 POR2X1_96/Y POR2X1_9/Y 0.10fF
C34465 POR2X1_241/B POR2X1_795/B 0.07fF
C34466 POR2X1_417/Y POR2X1_7/B 0.02fF
C34467 POR2X1_419/Y POR2X1_7/B 0.00fF
C34468 POR2X1_654/B POR2X1_121/Y 0.03fF
C34469 PAND2X1_436/A POR2X1_293/Y 0.07fF
C34470 POR2X1_687/A POR2X1_803/O 0.08fF
C34471 PAND2X1_714/CTRL PAND2X1_731/B 0.01fF
C34472 POR2X1_119/a_16_28# POR2X1_14/Y 0.02fF
C34473 POR2X1_144/Y VDD 0.04fF
C34474 PAND2X1_282/O PAND2X1_69/A 0.04fF
C34475 POR2X1_389/A PAND2X1_666/CTRL2 0.10fF
C34476 POR2X1_274/A POR2X1_366/A 0.03fF
C34477 PAND2X1_6/Y PAND2X1_73/Y 0.15fF
C34478 POR2X1_114/O POR2X1_590/A 0.02fF
C34479 POR2X1_487/Y POR2X1_42/Y 0.01fF
C34480 POR2X1_236/a_16_28# POR2X1_236/Y 0.03fF
C34481 POR2X1_42/a_16_28# POR2X1_37/Y 0.08fF
C34482 D_INPUT_3 POR2X1_14/CTRL2 0.04fF
C34483 POR2X1_567/B PAND2X1_60/B 0.05fF
C34484 PAND2X1_272/CTRL POR2X1_573/A 0.01fF
C34485 POR2X1_48/A POR2X1_239/Y 0.05fF
C34486 POR2X1_54/Y POR2X1_260/A 0.10fF
C34487 PAND2X1_229/CTRL POR2X1_579/Y 0.00fF
C34488 POR2X1_284/B VDD 0.01fF
C34489 POR2X1_335/A POR2X1_330/Y 0.05fF
C34490 POR2X1_272/CTRL2 POR2X1_184/Y 0.00fF
C34491 POR2X1_130/A INPUT_0 0.17fF
C34492 POR2X1_855/B POR2X1_678/Y 0.02fF
C34493 PAND2X1_473/Y PAND2X1_579/B 0.01fF
C34494 POR2X1_179/a_16_28# POR2X1_102/Y 0.08fF
C34495 POR2X1_257/A PAND2X1_303/Y 0.09fF
C34496 POR2X1_707/B POR2X1_614/A 0.01fF
C34497 PAND2X1_39/B POR2X1_733/Y 0.02fF
C34498 PAND2X1_793/Y PAND2X1_499/Y 0.03fF
C34499 PAND2X1_403/B PAND2X1_642/B 0.07fF
C34500 POR2X1_687/CTRL POR2X1_729/Y 0.01fF
C34501 PAND2X1_192/Y POR2X1_42/Y 0.03fF
C34502 PAND2X1_90/Y POR2X1_783/B 0.03fF
C34503 POR2X1_376/Y PAND2X1_375/O 0.01fF
C34504 PAND2X1_477/B POR2X1_417/Y 0.02fF
C34505 POR2X1_763/Y PAND2X1_713/B 0.03fF
C34506 PAND2X1_741/B POR2X1_7/B 0.62fF
C34507 POR2X1_316/Y POR2X1_329/A 0.03fF
C34508 PAND2X1_283/O POR2X1_734/A 0.05fF
C34509 POR2X1_855/Y VDD -0.00fF
C34510 POR2X1_734/B POR2X1_249/Y 0.02fF
C34511 POR2X1_423/CTRL POR2X1_387/Y 0.05fF
C34512 PAND2X1_20/A POR2X1_98/B 0.03fF
C34513 POR2X1_377/CTRL POR2X1_5/Y 0.01fF
C34514 PAND2X1_626/a_56_28# PAND2X1_96/B 0.00fF
C34515 POR2X1_719/CTRL POR2X1_121/B 0.08fF
C34516 POR2X1_407/A POR2X1_392/B 0.17fF
C34517 POR2X1_537/Y POR2X1_841/O 0.01fF
C34518 PAND2X1_23/Y POR2X1_480/A 0.50fF
C34519 PAND2X1_864/B GATE_366 0.12fF
C34520 POR2X1_809/A PAND2X1_761/O 0.02fF
C34521 POR2X1_186/Y POR2X1_731/CTRL 0.15fF
C34522 POR2X1_777/B PAND2X1_69/A 0.27fF
C34523 POR2X1_306/Y POR2X1_90/Y 0.01fF
C34524 PAND2X1_299/CTRL2 PAND2X1_32/B 0.01fF
C34525 PAND2X1_236/O PAND2X1_55/Y 0.07fF
C34526 POR2X1_106/CTRL PAND2X1_114/B 0.01fF
C34527 GATE_479 POR2X1_694/CTRL 0.03fF
C34528 POR2X1_383/A POR2X1_241/B 0.47fF
C34529 POR2X1_614/A PAND2X1_679/CTRL 0.01fF
C34530 POR2X1_567/B POR2X1_353/A 0.05fF
C34531 POR2X1_32/A PAND2X1_123/CTRL 0.01fF
C34532 POR2X1_49/Y PAND2X1_470/CTRL 0.01fF
C34533 PAND2X1_267/Y POR2X1_394/A 0.03fF
C34534 POR2X1_194/A PAND2X1_69/A 0.01fF
C34535 PAND2X1_807/B PAND2X1_854/A 0.73fF
C34536 POR2X1_782/A POR2X1_781/A 0.03fF
C34537 PAND2X1_244/CTRL PAND2X1_175/B 0.01fF
C34538 POR2X1_502/A POR2X1_857/B 0.03fF
C34539 PAND2X1_96/B PAND2X1_41/B 1.14fF
C34540 PAND2X1_253/CTRL2 POR2X1_241/B 0.01fF
C34541 PAND2X1_381/Y POR2X1_750/Y 0.03fF
C34542 POR2X1_333/Y PAND2X1_237/CTRL 0.01fF
C34543 POR2X1_97/CTRL2 POR2X1_78/A 0.03fF
C34544 PAND2X1_641/a_16_344# POR2X1_263/Y 0.01fF
C34545 POR2X1_505/CTRL2 POR2X1_669/B 0.02fF
C34546 PAND2X1_738/Y POR2X1_42/Y 0.05fF
C34547 POR2X1_61/Y POR2X1_556/Y 0.03fF
C34548 PAND2X1_23/Y POR2X1_243/Y 0.07fF
C34549 POR2X1_284/B POR2X1_741/Y 0.03fF
C34550 PAND2X1_41/B POR2X1_216/CTRL2 0.00fF
C34551 PAND2X1_512/O POR2X1_239/Y 0.02fF
C34552 POR2X1_327/Y POR2X1_558/B 1.58fF
C34553 PAND2X1_65/B PAND2X1_69/A 1.84fF
C34554 PAND2X1_467/B PAND2X1_467/CTRL 0.01fF
C34555 POR2X1_458/Y POR2X1_343/B 0.01fF
C34556 POR2X1_428/a_16_28# POR2X1_394/A 0.03fF
C34557 POR2X1_435/CTRL2 VDD -0.00fF
C34558 PAND2X1_736/A POR2X1_331/A 0.03fF
C34559 PAND2X1_738/B PAND2X1_149/A 0.34fF
C34560 POR2X1_750/B PAND2X1_63/B 0.05fF
C34561 POR2X1_76/Y POR2X1_455/A 0.02fF
C34562 POR2X1_495/O POR2X1_283/A 0.01fF
C34563 POR2X1_16/A POR2X1_14/Y 0.10fF
C34564 PAND2X1_773/O VDD 0.00fF
C34565 POR2X1_348/CTRL POR2X1_814/B 0.01fF
C34566 POR2X1_284/B PAND2X1_32/B 0.01fF
C34567 POR2X1_3/A POR2X1_2/CTRL2 0.00fF
C34568 PAND2X1_209/A VDD 0.00fF
C34569 POR2X1_8/Y POR2X1_83/B 0.07fF
C34570 POR2X1_66/B POR2X1_773/B 0.01fF
C34571 PAND2X1_478/a_16_344# POR2X1_46/Y 0.01fF
C34572 POR2X1_686/B POR2X1_605/A 0.02fF
C34573 POR2X1_447/B POR2X1_195/A 0.08fF
C34574 POR2X1_52/A PAND2X1_675/A 0.08fF
C34575 PAND2X1_220/Y PAND2X1_349/A 0.03fF
C34576 PAND2X1_862/B POR2X1_816/A 0.03fF
C34577 POR2X1_43/B PAND2X1_364/B 0.10fF
C34578 PAND2X1_3/A PAND2X1_3/B 0.03fF
C34579 PAND2X1_231/O POR2X1_229/Y 0.17fF
C34580 PAND2X1_830/Y POR2X1_184/Y 1.45fF
C34581 PAND2X1_464/Y PAND2X1_471/B 0.00fF
C34582 POR2X1_360/A POR2X1_68/A 0.03fF
C34583 POR2X1_826/O PAND2X1_338/B 0.16fF
C34584 PAND2X1_96/B POR2X1_402/B 0.03fF
C34585 POR2X1_750/B PAND2X1_1/a_16_344# 0.02fF
C34586 POR2X1_669/B PAND2X1_708/CTRL 0.04fF
C34587 POR2X1_119/Y POR2X1_23/Y 0.15fF
C34588 PAND2X1_673/O D_INPUT_3 0.15fF
C34589 POR2X1_383/A POR2X1_105/Y 0.54fF
C34590 POR2X1_502/A PAND2X1_752/Y 0.02fF
C34591 POR2X1_280/Y POR2X1_312/Y 0.09fF
C34592 POR2X1_156/B POR2X1_155/Y 0.01fF
C34593 POR2X1_225/a_56_344# POR2X1_129/Y 0.00fF
C34594 PAND2X1_535/Y VDD 0.36fF
C34595 INPUT_0 PAND2X1_150/O 0.01fF
C34596 PAND2X1_220/Y PAND2X1_114/B 0.03fF
C34597 POR2X1_390/B POR2X1_389/Y 0.32fF
C34598 PAND2X1_830/O PAND2X1_562/B 0.10fF
C34599 PAND2X1_476/A PAND2X1_571/A 0.27fF
C34600 POR2X1_78/B PAND2X1_60/B 7.77fF
C34601 POR2X1_273/Y POR2X1_42/Y 0.02fF
C34602 POR2X1_71/O POR2X1_60/A 0.02fF
C34603 POR2X1_493/B PAND2X1_41/B 0.01fF
C34604 PAND2X1_651/Y POR2X1_7/B 0.03fF
C34605 POR2X1_307/A VDD 0.00fF
C34606 PAND2X1_469/B POR2X1_152/A 0.07fF
C34607 PAND2X1_41/B PAND2X1_503/CTRL 0.00fF
C34608 PAND2X1_787/A PAND2X1_151/CTRL 0.03fF
C34609 POR2X1_862/CTRL POR2X1_647/B 0.01fF
C34610 POR2X1_634/CTRL POR2X1_559/A 0.29fF
C34611 PAND2X1_244/O POR2X1_153/Y 0.24fF
C34612 POR2X1_65/A POR2X1_291/CTRL 0.04fF
C34613 PAND2X1_568/B PAND2X1_568/CTRL2 0.03fF
C34614 PAND2X1_661/B POR2X1_277/CTRL 0.01fF
C34615 POR2X1_360/O VDD 0.00fF
C34616 POR2X1_795/O POR2X1_786/Y 0.04fF
C34617 POR2X1_311/Y PAND2X1_359/Y 0.04fF
C34618 POR2X1_52/A POR2X1_92/CTRL2 0.11fF
C34619 PAND2X1_137/O POR2X1_134/Y 0.03fF
C34620 POR2X1_85/CTRL POR2X1_23/Y 0.01fF
C34621 POR2X1_176/O POR2X1_83/B 0.01fF
C34622 POR2X1_427/Y PAND2X1_726/B 0.07fF
C34623 POR2X1_52/A POR2X1_526/a_76_344# 0.01fF
C34624 POR2X1_356/A POR2X1_535/A 0.03fF
C34625 INPUT_1 PAND2X1_721/O 0.01fF
C34626 POR2X1_290/Y POR2X1_291/Y 0.00fF
C34627 POR2X1_590/A POR2X1_188/Y 0.07fF
C34628 PAND2X1_821/m4_208_n4# POR2X1_509/m4_208_n4# 0.15fF
C34629 PAND2X1_388/Y PAND2X1_182/A 0.08fF
C34630 PAND2X1_599/O PAND2X1_69/A 0.04fF
C34631 PAND2X1_599/a_16_344# POR2X1_828/A 0.01fF
C34632 PAND2X1_20/A POR2X1_561/Y 0.04fF
C34633 POR2X1_83/B POR2X1_385/Y 0.03fF
C34634 POR2X1_514/CTRL2 PAND2X1_32/B 0.01fF
C34635 POR2X1_750/A POR2X1_749/a_76_344# 0.01fF
C34636 POR2X1_462/B POR2X1_790/B 0.00fF
C34637 POR2X1_40/a_16_28# INPUT_7 0.01fF
C34638 POR2X1_334/B POR2X1_68/B 0.19fF
C34639 POR2X1_389/A PAND2X1_385/CTRL 0.00fF
C34640 PAND2X1_797/Y POR2X1_669/B 0.95fF
C34641 PAND2X1_318/O POR2X1_91/Y 0.01fF
C34642 POR2X1_416/B POR2X1_699/CTRL 0.01fF
C34643 PAND2X1_96/B POR2X1_130/Y 0.03fF
C34644 PAND2X1_94/A VDD 3.92fF
C34645 POR2X1_327/Y POR2X1_543/A 0.10fF
C34646 POR2X1_591/O POR2X1_591/Y 0.03fF
C34647 PAND2X1_462/CTRL POR2X1_48/A 0.00fF
C34648 PAND2X1_539/Y VDD 0.12fF
C34649 POR2X1_138/CTRL POR2X1_318/A 0.04fF
C34650 POR2X1_193/A POR2X1_510/Y 0.04fF
C34651 PAND2X1_6/Y POR2X1_631/B 0.03fF
C34652 POR2X1_579/Y POR2X1_510/Y 0.03fF
C34653 POR2X1_78/B POR2X1_353/A 0.01fF
C34654 POR2X1_572/CTRL2 POR2X1_260/A 0.10fF
C34655 POR2X1_862/A PAND2X1_52/B 0.05fF
C34656 POR2X1_113/A PAND2X1_65/B 0.04fF
C34657 POR2X1_699/a_16_28# POR2X1_39/B 0.03fF
C34658 PAND2X1_847/CTRL2 POR2X1_48/A 0.03fF
C34659 POR2X1_136/Y POR2X1_42/Y 0.00fF
C34660 POR2X1_576/Y PAND2X1_32/B 0.14fF
C34661 POR2X1_76/B POR2X1_341/A 0.04fF
C34662 POR2X1_628/a_16_28# POR2X1_93/A 0.01fF
C34663 PAND2X1_57/B POR2X1_675/Y 0.03fF
C34664 POR2X1_124/B POR2X1_68/B 0.03fF
C34665 POR2X1_141/a_16_28# POR2X1_244/Y 0.02fF
C34666 PAND2X1_551/O PAND2X1_324/Y 0.16fF
C34667 POR2X1_673/A POR2X1_673/B 0.03fF
C34668 POR2X1_209/A POR2X1_535/a_16_28# 0.01fF
C34669 PAND2X1_73/Y POR2X1_632/Y 0.03fF
C34670 GATE_479 POR2X1_110/Y 0.03fF
C34671 PAND2X1_90/Y POR2X1_703/CTRL 0.05fF
C34672 POR2X1_121/A POR2X1_121/O 0.03fF
C34673 POR2X1_312/m4_208_n4# POR2X1_90/Y 0.01fF
C34674 PAND2X1_474/A POR2X1_171/Y 0.04fF
C34675 POR2X1_100/O PAND2X1_69/A 0.01fF
C34676 PAND2X1_659/Y PAND2X1_736/CTRL2 0.00fF
C34677 POR2X1_16/A PAND2X1_341/CTRL2 0.00fF
C34678 PAND2X1_23/Y POR2X1_787/CTRL 0.01fF
C34679 PAND2X1_498/CTRL POR2X1_260/A 0.01fF
C34680 PAND2X1_553/B PAND2X1_715/B 0.02fF
C34681 POR2X1_90/Y POR2X1_142/Y 0.03fF
C34682 POR2X1_38/B PAND2X1_670/CTRL2 0.01fF
C34683 D_GATE_662 PAND2X1_373/O 0.03fF
C34684 POR2X1_614/A POR2X1_510/Y 0.06fF
C34685 POR2X1_572/B POR2X1_276/Y 0.03fF
C34686 POR2X1_110/Y POR2X1_485/O 0.22fF
C34687 PAND2X1_495/CTRL2 PAND2X1_60/B 0.03fF
C34688 POR2X1_16/A POR2X1_55/Y 0.06fF
C34689 POR2X1_346/B PAND2X1_23/Y 0.03fF
C34690 PAND2X1_592/O PAND2X1_853/B 0.05fF
C34691 PAND2X1_651/Y PAND2X1_270/a_16_344# 0.12fF
C34692 PAND2X1_96/B POR2X1_228/Y 0.70fF
C34693 PAND2X1_297/CTRL2 POR2X1_402/A 0.01fF
C34694 PAND2X1_298/O PAND2X1_55/Y 0.00fF
C34695 PAND2X1_73/Y PAND2X1_52/B 0.14fF
C34696 PAND2X1_849/B POR2X1_43/B 0.04fF
C34697 PAND2X1_94/A PAND2X1_81/B 0.01fF
C34698 POR2X1_102/Y PAND2X1_862/CTRL2 0.01fF
C34699 POR2X1_804/A POR2X1_569/A 0.10fF
C34700 PAND2X1_291/m4_208_n4# POR2X1_35/Y 0.08fF
C34701 POR2X1_292/a_16_28# POR2X1_150/Y 0.02fF
C34702 POR2X1_346/B PAND2X1_625/O 0.00fF
C34703 POR2X1_730/B POR2X1_687/A 0.00fF
C34704 POR2X1_765/Y POR2X1_73/Y 1.24fF
C34705 PAND2X1_772/a_56_28# POR2X1_77/Y 0.00fF
C34706 POR2X1_215/Y PAND2X1_88/Y 0.01fF
C34707 PAND2X1_511/a_56_28# PAND2X1_48/A 0.00fF
C34708 POR2X1_40/Y POR2X1_77/Y 25.77fF
C34709 PAND2X1_798/B PAND2X1_510/O 0.00fF
C34710 POR2X1_831/CTRL2 POR2X1_814/A 0.00fF
C34711 POR2X1_278/Y PAND2X1_659/Y 0.01fF
C34712 PAND2X1_29/CTRL POR2X1_260/A 0.01fF
C34713 POR2X1_85/Y POR2X1_40/Y 0.02fF
C34714 POR2X1_129/Y POR2X1_586/a_16_28# 0.00fF
C34715 PAND2X1_94/A PAND2X1_32/B 0.17fF
C34716 POR2X1_732/B POR2X1_186/B 0.03fF
C34717 POR2X1_757/A POR2X1_394/A 0.03fF
C34718 POR2X1_54/a_16_28# POR2X1_401/B 0.05fF
C34719 POR2X1_614/A POR2X1_543/O 0.01fF
C34720 PAND2X1_659/Y POR2X1_829/A 0.03fF
C34721 PAND2X1_341/A PAND2X1_100/CTRL 0.01fF
C34722 POR2X1_57/A PAND2X1_569/B 0.08fF
C34723 POR2X1_57/A POR2X1_158/B 0.02fF
C34724 POR2X1_163/CTRL2 POR2X1_158/Y 0.00fF
C34725 POR2X1_39/a_16_28# POR2X1_669/B 0.03fF
C34726 POR2X1_96/CTRL POR2X1_38/B 0.00fF
C34727 PAND2X1_182/B PAND2X1_357/Y 0.13fF
C34728 POR2X1_38/Y PAND2X1_737/B 0.04fF
C34729 POR2X1_677/Y POR2X1_37/Y 0.33fF
C34730 POR2X1_283/A PAND2X1_549/B 0.03fF
C34731 PAND2X1_777/CTRL POR2X1_90/Y 0.00fF
C34732 POR2X1_220/Y POR2X1_330/CTRL 0.00fF
C34733 POR2X1_719/a_16_28# PAND2X1_60/B 0.03fF
C34734 POR2X1_537/Y POR2X1_662/Y 0.16fF
C34735 PAND2X1_242/Y POR2X1_102/Y 0.08fF
C34736 PAND2X1_185/a_76_28# POR2X1_77/Y 0.02fF
C34737 POR2X1_480/A POR2X1_711/Y 0.07fF
C34738 PAND2X1_687/B POR2X1_829/A 0.00fF
C34739 POR2X1_9/Y POR2X1_37/Y 0.42fF
C34740 POR2X1_416/B PAND2X1_733/Y 0.04fF
C34741 POR2X1_38/B PAND2X1_531/CTRL2 0.02fF
C34742 POR2X1_10/a_16_28# POR2X1_38/Y 0.04fF
C34743 POR2X1_730/Y POR2X1_162/Y 0.05fF
C34744 POR2X1_465/CTRL POR2X1_454/A 0.03fF
C34745 PAND2X1_172/O POR2X1_854/B 0.01fF
C34746 PAND2X1_436/A PAND2X1_242/Y 0.10fF
C34747 POR2X1_843/CTRL2 POR2X1_458/Y 0.01fF
C34748 POR2X1_394/A POR2X1_526/Y 0.06fF
C34749 POR2X1_862/O POR2X1_130/A 0.04fF
C34750 PAND2X1_716/B POR2X1_816/A 0.03fF
C34751 PAND2X1_285/CTRL2 POR2X1_282/Y 0.01fF
C34752 POR2X1_860/O POR2X1_383/A 0.02fF
C34753 POR2X1_68/A POR2X1_99/B 0.05fF
C34754 PAND2X1_793/Y POR2X1_39/B 0.03fF
C34755 POR2X1_840/B PAND2X1_48/A 0.03fF
C34756 PAND2X1_59/CTRL PAND2X1_18/B 0.01fF
C34757 POR2X1_416/B PAND2X1_198/Y 0.04fF
C34758 POR2X1_119/Y PAND2X1_836/O 0.12fF
C34759 PAND2X1_809/A PAND2X1_809/B 0.26fF
C34760 PAND2X1_841/B POR2X1_39/B 0.22fF
C34761 PAND2X1_94/A POR2X1_673/Y 0.03fF
C34762 POR2X1_349/CTRL POR2X1_532/A 0.01fF
C34763 POR2X1_814/B POR2X1_303/B 0.04fF
C34764 POR2X1_73/Y POR2X1_7/Y 0.06fF
C34765 PAND2X1_48/B POR2X1_39/B 0.03fF
C34766 PAND2X1_63/Y POR2X1_4/Y 2.49fF
C34767 POR2X1_327/Y POR2X1_538/A 0.01fF
C34768 POR2X1_614/A POR2X1_560/a_76_344# 0.01fF
C34769 PAND2X1_612/B POR2X1_472/B 1.80fF
C34770 POR2X1_636/A PAND2X1_52/B 0.01fF
C34771 PAND2X1_206/B POR2X1_32/A 0.07fF
C34772 POR2X1_732/B POR2X1_181/a_76_344# 0.03fF
C34773 PAND2X1_334/CTRL2 POR2X1_39/B 0.00fF
C34774 PAND2X1_69/A POR2X1_585/CTRL2 0.04fF
C34775 POR2X1_294/A PAND2X1_60/B 0.59fF
C34776 POR2X1_540/Y POR2X1_724/A 0.10fF
C34777 POR2X1_113/a_16_28# POR2X1_113/A 0.05fF
C34778 POR2X1_294/A POR2X1_758/a_16_28# 0.10fF
C34779 POR2X1_609/Y POR2X1_412/CTRL 0.00fF
C34780 POR2X1_325/A POR2X1_303/B 0.03fF
C34781 PAND2X1_96/B PAND2X1_122/O 0.01fF
C34782 POR2X1_327/Y POR2X1_362/A 0.03fF
C34783 PAND2X1_63/B PAND2X1_143/CTRL2 0.01fF
C34784 POR2X1_36/B POR2X1_328/m4_208_n4# 0.01fF
C34785 POR2X1_814/B POR2X1_846/A 0.03fF
C34786 POR2X1_635/B POR2X1_635/Y 0.24fF
C34787 PAND2X1_728/a_76_28# PAND2X1_853/B 0.02fF
C34788 POR2X1_75/CTRL2 POR2X1_416/B 0.01fF
C34789 POR2X1_416/B PAND2X1_642/B 0.03fF
C34790 POR2X1_187/CTRL POR2X1_385/Y 0.47fF
C34791 PAND2X1_221/a_76_28# POR2X1_250/Y 0.03fF
C34792 POR2X1_509/A PAND2X1_52/B 4.64fF
C34793 POR2X1_102/Y POR2X1_412/O 0.16fF
C34794 PAND2X1_55/Y POR2X1_556/CTRL2 0.01fF
C34795 POR2X1_134/Y POR2X1_77/Y 0.03fF
C34796 POR2X1_102/Y POR2X1_275/A 0.03fF
C34797 PAND2X1_606/CTRL2 POR2X1_37/Y 0.03fF
C34798 PAND2X1_587/O PAND2X1_52/B 0.13fF
C34799 POR2X1_192/B POR2X1_444/Y 1.21fF
C34800 PAND2X1_678/CTRL2 POR2X1_72/B 0.00fF
C34801 POR2X1_865/a_16_28# POR2X1_590/A 0.01fF
C34802 POR2X1_804/A PAND2X1_72/A 0.42fF
C34803 POR2X1_345/CTRL2 POR2X1_99/B 0.00fF
C34804 PAND2X1_717/A POR2X1_5/Y 0.03fF
C34805 POR2X1_4/Y POR2X1_260/A 0.03fF
C34806 POR2X1_122/CTRL2 PAND2X1_659/Y 0.00fF
C34807 POR2X1_677/Y POR2X1_293/Y 0.03fF
C34808 POR2X1_97/B POR2X1_186/B 0.03fF
C34809 POR2X1_711/Y PAND2X1_305/O 0.09fF
C34810 POR2X1_329/A PAND2X1_501/B 0.03fF
C34811 POR2X1_9/Y POR2X1_415/a_16_28# 0.04fF
C34812 PAND2X1_22/O PAND2X1_11/Y 0.02fF
C34813 PAND2X1_629/CTRL POR2X1_20/B 0.03fF
C34814 POR2X1_630/CTRL2 POR2X1_590/A 0.00fF
C34815 PAND2X1_39/B POR2X1_780/CTRL 0.02fF
C34816 PAND2X1_374/a_16_344# POR2X1_39/B 0.02fF
C34817 POR2X1_260/B POR2X1_267/O 0.01fF
C34818 POR2X1_475/A POR2X1_556/A 0.01fF
C34819 POR2X1_416/B PAND2X1_550/B 0.03fF
C34820 PAND2X1_163/O PAND2X1_52/B 0.03fF
C34821 POR2X1_210/A POR2X1_330/CTRL2 0.03fF
C34822 POR2X1_98/A PAND2X1_55/Y 0.00fF
C34823 POR2X1_676/O POR2X1_750/B 0.01fF
C34824 POR2X1_122/A POR2X1_20/B 0.01fF
C34825 POR2X1_353/Y POR2X1_443/a_56_344# 0.01fF
C34826 POR2X1_669/B POR2X1_428/a_16_28# 0.09fF
C34827 D_INPUT_0 POR2X1_296/B 0.20fF
C34828 POR2X1_460/Y VDD 0.24fF
C34829 POR2X1_445/A POR2X1_456/CTRL2 0.01fF
C34830 POR2X1_257/A INPUT_7 0.01fF
C34831 POR2X1_33/a_16_28# POR2X1_33/A 0.02fF
C34832 POR2X1_43/CTRL2 PAND2X1_560/B 0.12fF
C34833 POR2X1_760/A PAND2X1_216/CTRL2 0.03fF
C34834 POR2X1_66/B POR2X1_286/CTRL2 0.00fF
C34835 POR2X1_174/B POR2X1_97/A 0.07fF
C34836 PAND2X1_274/CTRL2 POR2X1_411/B 0.01fF
C34837 PAND2X1_313/O PAND2X1_72/A 0.03fF
C34838 POR2X1_355/B POR2X1_857/A 0.00fF
C34839 POR2X1_63/Y POR2X1_13/A 0.11fF
C34840 POR2X1_257/A PAND2X1_579/B 0.03fF
C34841 POR2X1_174/B POR2X1_836/B 0.01fF
C34842 POR2X1_462/B POR2X1_848/CTRL 0.01fF
C34843 POR2X1_624/Y PAND2X1_131/CTRL 0.03fF
C34844 POR2X1_661/A POR2X1_537/B 0.02fF
C34845 POR2X1_20/CTRL2 POR2X1_20/B 0.01fF
C34846 POR2X1_467/Y PAND2X1_73/Y 0.03fF
C34847 PAND2X1_20/A POR2X1_489/B 0.01fF
C34848 POR2X1_760/A PAND2X1_218/O 0.04fF
C34849 POR2X1_60/A POR2X1_102/Y 7.51fF
C34850 PAND2X1_48/A PAND2X1_56/A 0.08fF
C34851 PAND2X1_472/A PAND2X1_608/O 0.06fF
C34852 POR2X1_66/A PAND2X1_387/CTRL 0.01fF
C34853 POR2X1_23/Y POR2X1_238/CTRL 0.09fF
C34854 POR2X1_257/A INPUT_4 0.03fF
C34855 PAND2X1_206/A POR2X1_88/Y 0.03fF
C34856 POR2X1_814/A PAND2X1_69/A 2.45fF
C34857 POR2X1_54/Y POR2X1_790/CTRL2 0.03fF
C34858 POR2X1_23/Y PAND2X1_725/B 0.01fF
C34859 POR2X1_186/Y PAND2X1_331/CTRL2 0.01fF
C34860 POR2X1_9/Y POR2X1_408/Y 0.26fF
C34861 POR2X1_456/B PAND2X1_125/O 0.09fF
C34862 POR2X1_102/Y POR2X1_591/A 0.02fF
C34863 PAND2X1_695/O PAND2X1_59/B 0.05fF
C34864 PAND2X1_688/CTRL2 POR2X1_48/A 0.00fF
C34865 D_GATE_662 POR2X1_444/CTRL 0.05fF
C34866 POR2X1_257/A POR2X1_763/Y 0.10fF
C34867 POR2X1_254/Y POR2X1_260/B 0.17fF
C34868 POR2X1_389/A PAND2X1_607/m4_208_n4# 0.15fF
C34869 PAND2X1_436/A POR2X1_60/A 0.19fF
C34870 POR2X1_400/B PAND2X1_41/B 0.02fF
C34871 PAND2X1_805/a_76_28# PAND2X1_287/Y 0.02fF
C34872 POR2X1_862/B POR2X1_590/A 0.05fF
C34873 POR2X1_257/A PAND2X1_115/B 0.03fF
C34874 POR2X1_866/A PAND2X1_511/O 0.11fF
C34875 POR2X1_96/A PAND2X1_404/Y 0.03fF
C34876 POR2X1_265/CTRL2 PAND2X1_35/Y 0.01fF
C34877 PAND2X1_838/B POR2X1_42/Y 0.99fF
C34878 POR2X1_407/A POR2X1_864/A 0.03fF
C34879 POR2X1_66/A POR2X1_403/Y 0.02fF
C34880 POR2X1_556/A POR2X1_218/A 0.06fF
C34881 D_INPUT_0 POR2X1_236/Y 0.06fF
C34882 PAND2X1_42/CTRL POR2X1_267/A 0.02fF
C34883 D_INPUT_5 PAND2X1_17/CTRL 0.01fF
C34884 PAND2X1_480/B PAND2X1_205/A 0.05fF
C34885 POR2X1_63/O POR2X1_63/Y 0.01fF
C34886 POR2X1_257/A PAND2X1_658/A 0.02fF
C34887 POR2X1_477/Y VDD -0.00fF
C34888 POR2X1_460/Y PAND2X1_32/B 0.01fF
C34889 PAND2X1_90/Y POR2X1_296/B 0.12fF
C34890 POR2X1_257/A POR2X1_426/CTRL 0.01fF
C34891 PAND2X1_479/B PAND2X1_571/A 0.00fF
C34892 PAND2X1_473/Y PAND2X1_571/O 0.01fF
C34893 POR2X1_278/Y POR2X1_37/Y 0.17fF
C34894 POR2X1_801/B VDD 0.05fF
C34895 POR2X1_67/Y POR2X1_391/O 0.01fF
C34896 POR2X1_502/A POR2X1_66/A 0.30fF
C34897 POR2X1_276/B POR2X1_513/Y 0.06fF
C34898 PAND2X1_23/Y PAND2X1_487/O 0.12fF
C34899 POR2X1_760/A PAND2X1_799/CTRL 0.01fF
C34900 PAND2X1_808/Y PAND2X1_774/a_76_28# 0.01fF
C34901 PAND2X1_65/B POR2X1_506/B 0.02fF
C34902 POR2X1_99/A PAND2X1_41/B 0.01fF
C34903 POR2X1_605/O PAND2X1_90/Y 0.09fF
C34904 POR2X1_865/B POR2X1_499/A 0.09fF
C34905 POR2X1_417/Y PAND2X1_220/Y 0.03fF
C34906 PAND2X1_661/B POR2X1_63/Y 0.03fF
C34907 PAND2X1_809/CTRL PAND2X1_539/Y 0.01fF
C34908 PAND2X1_805/Y POR2X1_7/B 0.06fF
C34909 POR2X1_39/O POR2X1_72/B 0.01fF
C34910 PAND2X1_11/Y VDD 0.84fF
C34911 PAND2X1_362/A GATE_741 0.06fF
C34912 POR2X1_66/A PAND2X1_176/O 0.18fF
C34913 POR2X1_416/B PAND2X1_840/Y 0.00fF
C34914 POR2X1_257/A POR2X1_73/Y 0.13fF
C34915 POR2X1_606/Y VDD 0.04fF
C34916 POR2X1_661/A PAND2X1_48/A 0.07fF
C34917 PAND2X1_826/CTRL2 PAND2X1_96/B 0.03fF
C34918 POR2X1_116/A PAND2X1_60/B 0.03fF
C34919 POR2X1_847/O POR2X1_283/A 0.03fF
C34920 PAND2X1_47/B PAND2X1_587/Y 0.01fF
C34921 POR2X1_640/Y PAND2X1_65/B 0.00fF
C34922 POR2X1_23/Y PAND2X1_775/a_76_28# 0.02fF
C34923 POR2X1_83/B POR2X1_516/B 0.03fF
C34924 PAND2X1_391/CTRL2 POR2X1_42/Y 0.10fF
C34925 POR2X1_117/a_16_28# POR2X1_72/B 0.05fF
C34926 POR2X1_78/B POR2X1_254/A 0.05fF
C34927 POR2X1_56/B POR2X1_496/Y 0.12fF
C34928 PAND2X1_406/CTRL2 PAND2X1_32/B 0.02fF
C34929 POR2X1_669/B POR2X1_372/Y 0.07fF
C34930 PAND2X1_79/CTRL2 D_INPUT_0 0.01fF
C34931 POR2X1_376/B PAND2X1_185/a_16_344# 0.04fF
C34932 PAND2X1_865/a_76_28# POR2X1_329/A 0.02fF
C34933 POR2X1_139/Y POR2X1_296/B 0.01fF
C34934 PAND2X1_432/CTRL VDD 0.00fF
C34935 POR2X1_78/B POR2X1_750/B 0.14fF
C34936 POR2X1_688/Y POR2X1_532/A 0.01fF
C34937 POR2X1_611/m4_208_n4# POR2X1_4/Y 0.07fF
C34938 POR2X1_502/A POR2X1_634/CTRL2 0.14fF
C34939 POR2X1_23/Y POR2X1_237/Y 0.05fF
C34940 POR2X1_276/B POR2X1_366/A 0.02fF
C34941 POR2X1_445/A POR2X1_724/A 0.07fF
C34942 INPUT_0 POR2X1_750/A 0.03fF
C34943 PAND2X1_45/O POR2X1_260/A 0.04fF
C34944 D_INPUT_0 POR2X1_501/O 0.01fF
C34945 PAND2X1_39/B PAND2X1_393/CTRL 0.01fF
C34946 POR2X1_360/A PAND2X1_58/A 0.02fF
C34947 POR2X1_83/A POR2X1_409/B 0.04fF
C34948 PAND2X1_26/A D_INPUT_6 0.00fF
C34949 POR2X1_306/Y INPUT_0 0.01fF
C34950 POR2X1_333/A POR2X1_468/O 0.07fF
C34951 POR2X1_315/Y POR2X1_442/CTRL2 0.05fF
C34952 POR2X1_154/CTRL POR2X1_750/B 0.00fF
C34953 PAND2X1_809/A POR2X1_102/Y 0.03fF
C34954 POR2X1_814/B POR2X1_461/B 0.01fF
C34955 POR2X1_49/Y PAND2X1_579/B 0.01fF
C34956 PAND2X1_475/a_56_28# INPUT_0 0.00fF
C34957 POR2X1_855/B PAND2X1_39/B 0.00fF
C34958 POR2X1_106/CTRL2 POR2X1_183/Y 0.00fF
C34959 PAND2X1_58/A POR2X1_756/O 0.17fF
C34960 POR2X1_669/B POR2X1_519/Y 0.07fF
C34961 POR2X1_498/O POR2X1_72/B 0.06fF
C34962 POR2X1_709/A PAND2X1_748/CTRL2 0.01fF
C34963 POR2X1_448/Y VDD 0.10fF
C34964 PAND2X1_721/CTRL VDD 0.00fF
C34965 POR2X1_57/m4_208_n4# PAND2X1_214/m4_208_n4# 0.05fF
C34966 PAND2X1_94/A PAND2X1_9/Y 0.19fF
C34967 POR2X1_388/O POR2X1_66/A 0.18fF
C34968 POR2X1_52/A PAND2X1_195/a_16_344# 0.02fF
C34969 PAND2X1_291/CTRL2 PAND2X1_93/B 0.00fF
C34970 INPUT_2 POR2X1_37/Y 0.05fF
C34971 D_INPUT_0 POR2X1_796/a_16_28# 0.02fF
C34972 POR2X1_567/B POR2X1_714/CTRL2 0.31fF
C34973 POR2X1_218/Y POR2X1_112/Y 0.07fF
C34974 PAND2X1_114/Y POR2X1_40/Y 0.18fF
C34975 POR2X1_811/CTRL POR2X1_532/A 0.01fF
C34976 POR2X1_253/Y POR2X1_669/B 0.01fF
C34977 PAND2X1_404/Y POR2X1_7/A 0.03fF
C34978 INPUT_1 PAND2X1_33/a_76_28# 0.01fF
C34979 POR2X1_94/A POR2X1_7/B 1.66fF
C34980 PAND2X1_577/B PAND2X1_569/Y 0.01fF
C34981 POR2X1_558/B POR2X1_361/CTRL2 0.00fF
C34982 POR2X1_471/A PAND2X1_313/CTRL 0.00fF
C34983 POR2X1_801/B PAND2X1_32/B 0.01fF
C34984 POR2X1_20/B PAND2X1_563/A 0.03fF
C34985 POR2X1_29/Y POR2X1_669/B 0.04fF
C34986 POR2X1_485/Y POR2X1_394/A 6.92fF
C34987 POR2X1_559/a_16_28# POR2X1_66/A 0.02fF
C34988 POR2X1_65/A POR2X1_693/O 0.01fF
C34989 PAND2X1_217/B POR2X1_275/O 0.02fF
C34990 POR2X1_13/A PAND2X1_768/Y 0.01fF
C34991 POR2X1_697/a_16_28# POR2X1_236/Y 0.01fF
C34992 POR2X1_49/Y POR2X1_763/Y 0.07fF
C34993 PAND2X1_742/B POR2X1_40/Y 0.01fF
C34994 POR2X1_814/B PAND2X1_385/CTRL2 0.03fF
C34995 POR2X1_567/B POR2X1_704/CTRL 0.01fF
C34996 PAND2X1_658/CTRL2 PAND2X1_658/B 0.17fF
C34997 POR2X1_41/B POR2X1_5/Y 0.20fF
C34998 PAND2X1_845/CTRL POR2X1_60/A 0.02fF
C34999 POR2X1_130/A PAND2X1_511/CTRL2 0.01fF
C35000 POR2X1_556/A POR2X1_557/B 0.03fF
C35001 PAND2X1_11/Y PAND2X1_32/B 0.06fF
C35002 D_INPUT_2 POR2X1_611/CTRL2 0.01fF
C35003 POR2X1_719/O POR2X1_66/A 0.01fF
C35004 PAND2X1_7/O POR2X1_750/B 0.25fF
C35005 PAND2X1_615/O POR2X1_614/Y -0.00fF
C35006 POR2X1_614/A POR2X1_864/CTRL 0.00fF
C35007 PAND2X1_23/Y POR2X1_402/CTRL2 0.00fF
C35008 PAND2X1_84/Y PAND2X1_735/Y 0.01fF
C35009 PAND2X1_423/O PAND2X1_55/Y 0.04fF
C35010 POR2X1_669/B POR2X1_526/Y 0.04fF
C35011 POR2X1_278/Y POR2X1_406/Y 0.08fF
C35012 PAND2X1_860/A POR2X1_173/CTRL2 0.01fF
C35013 PAND2X1_139/B POR2X1_13/A 0.00fF
C35014 POR2X1_848/A POR2X1_754/CTRL2 0.03fF
C35015 POR2X1_555/A POR2X1_294/B 0.01fF
C35016 POR2X1_448/O POR2X1_788/B 0.02fF
C35017 D_INPUT_2 POR2X1_293/O 0.01fF
C35018 POR2X1_54/Y POR2X1_559/A 0.97fF
C35019 POR2X1_121/CTRL POR2X1_590/A 0.01fF
C35020 POR2X1_186/Y PAND2X1_146/O 0.02fF
C35021 PAND2X1_758/CTRL POR2X1_236/Y 0.03fF
C35022 POR2X1_220/B POR2X1_738/A 0.03fF
C35023 POR2X1_108/O POR2X1_60/A 0.13fF
C35024 POR2X1_590/A POR2X1_510/Y 0.01fF
C35025 PAND2X1_796/B POR2X1_371/CTRL2 0.00fF
C35026 PAND2X1_351/O VDD 0.00fF
C35027 PAND2X1_433/CTRL POR2X1_480/A 0.03fF
C35028 POR2X1_818/CTRL POR2X1_294/A 0.01fF
C35029 POR2X1_65/A POR2X1_56/Y 0.01fF
C35030 PAND2X1_205/Y POR2X1_816/A 0.03fF
C35031 PAND2X1_84/Y PAND2X1_493/Y 0.01fF
C35032 POR2X1_661/Y POR2X1_725/Y 0.09fF
C35033 POR2X1_258/CTRL2 POR2X1_312/Y 0.02fF
C35034 PAND2X1_265/O PAND2X1_60/B 0.02fF
C35035 PAND2X1_865/Y POR2X1_150/Y 0.07fF
C35036 POR2X1_29/A POR2X1_748/Y 0.01fF
C35037 POR2X1_368/O POR2X1_293/Y 0.12fF
C35038 PAND2X1_675/A PAND2X1_180/O 0.07fF
C35039 PAND2X1_50/m4_208_n4# INPUT_5 0.21fF
C35040 POR2X1_51/A POR2X1_7/B 0.02fF
C35041 PAND2X1_652/A PAND2X1_473/B 0.03fF
C35042 PAND2X1_6/Y POR2X1_61/Y 0.05fF
C35043 POR2X1_278/Y POR2X1_293/Y 0.10fF
C35044 PAND2X1_615/CTRL POR2X1_94/A 0.09fF
C35045 POR2X1_852/B PAND2X1_69/A 0.01fF
C35046 POR2X1_49/Y POR2X1_73/Y 0.17fF
C35047 POR2X1_407/A POR2X1_362/B 0.06fF
C35048 POR2X1_83/B PAND2X1_550/Y 0.04fF
C35049 POR2X1_14/Y PAND2X1_549/B 0.03fF
C35050 POR2X1_43/B POR2X1_58/O 0.02fF
C35051 POR2X1_614/A PAND2X1_263/CTRL 0.01fF
C35052 POR2X1_254/Y PAND2X1_55/Y 1.59fF
C35053 POR2X1_388/a_16_28# POR2X1_750/B 0.02fF
C35054 PAND2X1_453/A PAND2X1_549/B 0.03fF
C35055 POR2X1_748/A POR2X1_387/Y 0.10fF
C35056 POR2X1_215/O POR2X1_740/Y 0.02fF
C35057 POR2X1_72/B POR2X1_172/Y 0.90fF
C35058 POR2X1_7/B PAND2X1_335/CTRL 0.01fF
C35059 POR2X1_433/a_76_344# PAND2X1_349/A 0.00fF
C35060 POR2X1_855/Y POR2X1_149/Y 0.03fF
C35061 PAND2X1_94/A PAND2X1_15/O 0.17fF
C35062 PAND2X1_48/B POR2X1_651/CTRL2 0.03fF
C35063 D_INPUT_0 POR2X1_590/Y 0.05fF
C35064 POR2X1_174/CTRL PAND2X1_73/Y 0.01fF
C35065 PAND2X1_242/Y POR2X1_677/Y 0.05fF
C35066 PAND2X1_809/B PAND2X1_810/B 0.01fF
C35067 POR2X1_578/Y POR2X1_579/Y 0.08fF
C35068 POR2X1_83/B POR2X1_172/O 0.01fF
C35069 PAND2X1_94/A POR2X1_267/A 0.05fF
C35070 POR2X1_614/A POR2X1_471/CTRL2 0.03fF
C35071 POR2X1_302/a_76_344# POR2X1_114/B 0.00fF
C35072 PAND2X1_96/B POR2X1_476/Y 0.01fF
C35073 POR2X1_514/O INPUT_0 0.03fF
C35074 POR2X1_466/A POR2X1_186/B 0.03fF
C35075 POR2X1_802/B POR2X1_532/Y 0.10fF
C35076 POR2X1_779/A POR2X1_779/a_16_28# 0.03fF
C35077 POR2X1_445/CTRL2 POR2X1_455/A 0.01fF
C35078 POR2X1_267/B POR2X1_318/A 0.03fF
C35079 POR2X1_61/O PAND2X1_58/A 0.13fF
C35080 POR2X1_861/CTRL POR2X1_404/Y 0.00fF
C35081 PAND2X1_643/CTRL POR2X1_7/B 0.01fF
C35082 POR2X1_700/Y VDD 0.00fF
C35083 PAND2X1_742/a_76_28# POR2X1_283/A 0.02fF
C35084 POR2X1_32/A PAND2X1_560/B 0.03fF
C35085 PAND2X1_90/A POR2X1_334/B 0.03fF
C35086 PAND2X1_93/B POR2X1_540/Y 0.08fF
C35087 POR2X1_115/CTRL POR2X1_112/Y 0.01fF
C35088 POR2X1_49/Y PAND2X1_244/B 0.03fF
C35089 POR2X1_401/B PAND2X1_69/A 0.04fF
C35090 POR2X1_96/A PAND2X1_565/A 1.55fF
C35091 POR2X1_43/B PAND2X1_523/O 0.02fF
C35092 POR2X1_101/Y POR2X1_734/A 0.10fF
C35093 POR2X1_114/Y D_INPUT_1 0.01fF
C35094 POR2X1_785/A POR2X1_341/CTRL 0.03fF
C35095 POR2X1_382/Y VDD 0.11fF
C35096 POR2X1_98/B VDD 0.04fF
C35097 INPUT_1 PAND2X1_614/CTRL2 0.01fF
C35098 POR2X1_278/Y PAND2X1_676/CTRL2 0.05fF
C35099 POR2X1_41/B POR2X1_310/O 0.05fF
C35100 PAND2X1_65/O POR2X1_4/Y 0.02fF
C35101 POR2X1_502/A POR2X1_532/A 0.33fF
C35102 PAND2X1_69/A INPUT_5 0.03fF
C35103 PAND2X1_4/O INPUT_0 0.10fF
C35104 PAND2X1_319/B PAND2X1_151/O 0.02fF
C35105 POR2X1_305/Y POR2X1_42/Y 0.36fF
C35106 POR2X1_783/A POR2X1_532/A 0.01fF
C35107 POR2X1_68/A PAND2X1_275/CTRL 0.07fF
C35108 POR2X1_537/Y POR2X1_646/Y 0.16fF
C35109 PAND2X1_90/Y POR2X1_520/CTRL 0.01fF
C35110 INPUT_2 POR2X1_293/Y 0.02fF
C35111 POR2X1_7/B POR2X1_386/CTRL 0.01fF
C35112 POR2X1_376/B POR2X1_428/CTRL 0.04fF
C35113 POR2X1_46/CTRL POR2X1_153/Y 0.05fF
C35114 PAND2X1_150/CTRL2 POR2X1_404/Y 0.01fF
C35115 POR2X1_186/Y POR2X1_703/Y 0.10fF
C35116 INPUT_0 PAND2X1_175/B 0.03fF
C35117 PAND2X1_52/Y POR2X1_260/A 0.10fF
C35118 POR2X1_262/O POR2X1_73/Y 0.01fF
C35119 POR2X1_827/Y POR2X1_39/B 0.01fF
C35120 PAND2X1_610/O POR2X1_48/A 0.01fF
C35121 PAND2X1_682/CTRL2 POR2X1_614/A 0.00fF
C35122 PAND2X1_6/A PAND2X1_658/B 0.10fF
C35123 POR2X1_247/CTRL POR2X1_532/A 0.01fF
C35124 POR2X1_78/B POR2X1_200/A 0.01fF
C35125 POR2X1_702/B POR2X1_260/A 0.02fF
C35126 POR2X1_806/CTRL POR2X1_737/A 0.01fF
C35127 PAND2X1_65/B POR2X1_576/CTRL 0.00fF
C35128 POR2X1_164/CTRL POR2X1_693/Y 0.01fF
C35129 POR2X1_67/a_76_344# POR2X1_39/B 0.03fF
C35130 PAND2X1_473/B PAND2X1_175/O 0.04fF
C35131 POR2X1_532/A PAND2X1_530/CTRL2 0.01fF
C35132 POR2X1_383/A PAND2X1_280/CTRL2 0.03fF
C35133 POR2X1_52/A PAND2X1_389/Y 0.01fF
C35134 PAND2X1_6/Y POR2X1_35/Y 0.02fF
C35135 PAND2X1_853/CTRL2 PAND2X1_653/Y 0.03fF
C35136 PAND2X1_90/Y POR2X1_543/CTRL 0.19fF
C35137 POR2X1_532/A POR2X1_532/Y 0.83fF
C35138 POR2X1_130/A POR2X1_796/A 0.03fF
C35139 POR2X1_590/A POR2X1_741/CTRL2 0.03fF
C35140 POR2X1_123/CTRL2 PAND2X1_60/B 0.01fF
C35141 PAND2X1_698/a_56_28# PAND2X1_65/B 0.00fF
C35142 POR2X1_315/Y PAND2X1_480/B 0.07fF
C35143 PAND2X1_724/B POR2X1_91/Y 0.03fF
C35144 PAND2X1_852/O PAND2X1_852/B 0.00fF
C35145 PAND2X1_61/Y PAND2X1_358/A 0.01fF
C35146 POR2X1_42/Y POR2X1_748/a_16_28# 0.09fF
C35147 POR2X1_750/B POR2X1_735/CTRL 0.26fF
C35148 POR2X1_673/A POR2X1_260/A 0.84fF
C35149 PAND2X1_96/B POR2X1_713/O 0.02fF
C35150 PAND2X1_388/Y POR2X1_55/Y 0.03fF
C35151 PAND2X1_865/Y PAND2X1_794/O 0.00fF
C35152 PAND2X1_231/a_56_28# POR2X1_153/Y 0.00fF
C35153 POR2X1_220/B POR2X1_731/Y 0.01fF
C35154 POR2X1_517/CTRL2 POR2X1_667/A 0.01fF
C35155 PAND2X1_58/A PAND2X1_304/CTRL 0.01fF
C35156 PAND2X1_467/Y POR2X1_46/Y 5.39fF
C35157 POR2X1_268/CTRL POR2X1_39/B 0.01fF
C35158 PAND2X1_23/Y POR2X1_319/Y 0.03fF
C35159 POR2X1_124/a_16_28# PAND2X1_60/B 0.03fF
C35160 POR2X1_832/B POR2X1_592/CTRL 0.01fF
C35161 POR2X1_95/CTRL2 POR2X1_40/Y 0.01fF
C35162 PAND2X1_63/Y D_INPUT_1 0.07fF
C35163 POR2X1_220/Y POR2X1_703/A 0.07fF
C35164 POR2X1_55/Y PAND2X1_549/B 0.04fF
C35165 PAND2X1_48/B POR2X1_181/B 0.11fF
C35166 PAND2X1_803/Y PAND2X1_190/Y 0.01fF
C35167 POR2X1_677/Y POR2X1_275/A 0.25fF
C35168 POR2X1_71/CTRL PAND2X1_84/Y 0.01fF
C35169 PAND2X1_96/B POR2X1_758/CTRL2 0.01fF
C35170 POR2X1_313/O POR2X1_90/Y 0.04fF
C35171 VDD POR2X1_733/Y 0.02fF
C35172 POR2X1_208/Y POR2X1_206/O 0.06fF
C35173 PAND2X1_61/a_56_28# POR2X1_39/B 0.00fF
C35174 POR2X1_60/A POR2X1_761/A 0.03fF
C35175 PAND2X1_200/B VDD 0.23fF
C35176 POR2X1_859/A POR2X1_753/CTRL 0.05fF
C35177 PAND2X1_472/O PAND2X1_472/B 0.01fF
C35178 POR2X1_267/Y POR2X1_361/O 0.20fF
C35179 POR2X1_335/A POR2X1_538/A 0.01fF
C35180 POR2X1_140/A POR2X1_140/a_16_28# 0.03fF
C35181 GATE_741 PAND2X1_366/CTRL2 0.01fF
C35182 POR2X1_516/Y POR2X1_39/B 0.03fF
C35183 POR2X1_102/Y PAND2X1_339/CTRL2 0.01fF
C35184 POR2X1_356/A POR2X1_351/a_16_28# 0.10fF
C35185 POR2X1_409/Y POR2X1_7/B 0.06fF
C35186 POR2X1_366/Y PAND2X1_313/CTRL2 -0.01fF
C35187 PAND2X1_645/B POR2X1_591/Y 0.07fF
C35188 POR2X1_113/Y D_INPUT_1 0.81fF
C35189 POR2X1_846/A POR2X1_496/CTRL2 0.00fF
C35190 POR2X1_555/A POR2X1_567/A 0.10fF
C35191 PAND2X1_23/Y POR2X1_325/a_16_28# 0.02fF
C35192 PAND2X1_35/Y PAND2X1_560/B 0.04fF
C35193 POR2X1_559/m4_208_n4# POR2X1_68/B 0.09fF
C35194 POR2X1_102/a_16_28# POR2X1_40/Y 0.01fF
C35195 POR2X1_83/B PAND2X1_327/CTRL 0.01fF
C35196 POR2X1_57/A PAND2X1_787/A 0.06fF
C35197 PAND2X1_90/Y PAND2X1_759/CTRL2 0.10fF
C35198 PAND2X1_469/B PAND2X1_353/a_16_344# 0.03fF
C35199 POR2X1_122/CTRL2 POR2X1_293/Y 0.00fF
C35200 POR2X1_561/Y VDD 0.06fF
C35201 PAND2X1_858/O INPUT_0 0.02fF
C35202 PAND2X1_744/CTRL2 POR2X1_260/A 0.01fF
C35203 POR2X1_101/Y POR2X1_786/Y 0.10fF
C35204 PAND2X1_23/Y POR2X1_507/A 0.16fF
C35205 PAND2X1_6/Y PAND2X1_368/O 0.02fF
C35206 POR2X1_389/A PAND2X1_60/B 0.01fF
C35207 PAND2X1_771/B PAND2X1_771/O 0.00fF
C35208 POR2X1_643/CTRL2 POR2X1_260/B 0.01fF
C35209 POR2X1_379/CTRL POR2X1_532/A 0.01fF
C35210 POR2X1_570/B POR2X1_569/A 0.07fF
C35211 PAND2X1_720/O POR2X1_73/Y 0.05fF
C35212 PAND2X1_559/CTRL POR2X1_73/Y 0.07fF
C35213 PAND2X1_504/CTRL2 POR2X1_507/A 0.03fF
C35214 PAND2X1_73/Y POR2X1_579/CTRL2 0.01fF
C35215 PAND2X1_484/CTRL POR2X1_294/B 0.03fF
C35216 POR2X1_192/Y POR2X1_566/a_16_28# 0.02fF
C35217 PAND2X1_373/CTRL2 POR2X1_540/A 0.01fF
C35218 PAND2X1_763/a_76_28# PAND2X1_48/A 0.04fF
C35219 POR2X1_741/Y POR2X1_733/Y 0.02fF
C35220 POR2X1_327/Y POR2X1_572/B 3.59fF
C35221 POR2X1_816/A POR2X1_260/A 0.03fF
C35222 POR2X1_61/Y POR2X1_632/Y 0.08fF
C35223 POR2X1_462/B POR2X1_260/A 0.04fF
C35224 PAND2X1_191/CTRL PAND2X1_730/A 0.00fF
C35225 D_INPUT_1 POR2X1_260/A 0.19fF
C35226 PAND2X1_39/B PAND2X1_32/O 0.05fF
C35227 POR2X1_51/B INPUT_6 0.07fF
C35228 POR2X1_794/B PAND2X1_72/A 0.03fF
C35229 GATE_865 VDD 0.00fF
C35230 PAND2X1_738/O POR2X1_39/B 0.06fF
C35231 POR2X1_119/Y POR2X1_290/Y 0.07fF
C35232 POR2X1_827/Y POR2X1_827/O 0.01fF
C35233 POR2X1_343/Y POR2X1_287/B 0.01fF
C35234 POR2X1_315/Y PAND2X1_303/B 0.04fF
C35235 PAND2X1_171/CTRL2 D_GATE_741 0.01fF
C35236 POR2X1_494/Y POR2X1_171/Y 0.16fF
C35237 INPUT_0 PAND2X1_136/O 0.04fF
C35238 POR2X1_5/Y POR2X1_77/Y 6.11fF
C35239 POR2X1_826/O POR2X1_77/Y 0.15fF
C35240 POR2X1_41/O POR2X1_73/Y 0.03fF
C35241 PAND2X1_330/O POR2X1_331/A 0.01fF
C35242 POR2X1_327/Y POR2X1_614/A 8.25fF
C35243 POR2X1_483/A POR2X1_343/Y 0.05fF
C35244 POR2X1_343/Y POR2X1_778/CTRL 0.07fF
C35245 POR2X1_299/O PAND2X1_308/Y 0.02fF
C35246 POR2X1_499/A POR2X1_341/A 0.00fF
C35247 POR2X1_119/Y POR2X1_238/Y 1.67fF
C35248 POR2X1_333/Y POR2X1_341/Y 0.05fF
C35249 PAND2X1_61/O POR2X1_9/Y 0.01fF
C35250 POR2X1_43/B PAND2X1_851/O 0.17fF
C35251 POR2X1_63/Y POR2X1_813/CTRL 0.02fF
C35252 PAND2X1_96/B POR2X1_579/B 0.02fF
C35253 POR2X1_107/a_76_344# POR2X1_77/Y 0.02fF
C35254 POR2X1_722/Y POR2X1_513/A 0.02fF
C35255 POR2X1_456/B POR2X1_366/A 0.03fF
C35256 PAND2X1_844/B PAND2X1_560/B 0.01fF
C35257 POR2X1_442/O POR2X1_411/B 0.02fF
C35258 POR2X1_63/a_76_344# POR2X1_62/Y 0.01fF
C35259 POR2X1_112/O POR2X1_775/A 0.01fF
C35260 POR2X1_51/B POR2X1_31/a_16_28# 0.03fF
C35261 D_INPUT_7 PAND2X1_429/O 0.17fF
C35262 POR2X1_537/Y POR2X1_804/A 0.03fF
C35263 POR2X1_204/O POR2X1_4/Y 0.01fF
C35264 POR2X1_776/B POR2X1_567/CTRL 0.01fF
C35265 POR2X1_657/Y POR2X1_222/CTRL 0.01fF
C35266 PAND2X1_96/B POR2X1_571/Y 0.03fF
C35267 POR2X1_60/A POR2X1_9/Y 6.16fF
C35268 POR2X1_145/a_16_28# PAND2X1_797/Y 0.02fF
C35269 PAND2X1_476/A PAND2X1_472/A 0.02fF
C35270 POR2X1_334/Y PAND2X1_60/B 0.04fF
C35271 POR2X1_67/Y PAND2X1_381/Y 0.01fF
C35272 PAND2X1_755/CTRL PAND2X1_72/A 0.01fF
C35273 POR2X1_16/A PAND2X1_124/O 0.07fF
C35274 POR2X1_112/O POR2X1_112/Y 0.00fF
C35275 POR2X1_99/B PAND2X1_96/B 0.03fF
C35276 POR2X1_102/CTRL2 D_INPUT_1 0.01fF
C35277 PAND2X1_20/A PAND2X1_607/a_56_28# 0.00fF
C35278 POR2X1_736/A PAND2X1_178/CTRL 0.02fF
C35279 POR2X1_327/Y POR2X1_440/Y 0.03fF
C35280 POR2X1_688/O D_INPUT_0 0.17fF
C35281 PAND2X1_127/O POR2X1_456/B 0.01fF
C35282 POR2X1_16/A PAND2X1_704/CTRL2 0.01fF
C35283 PAND2X1_526/CTRL2 PAND2X1_32/B 0.00fF
C35284 POR2X1_329/A PAND2X1_219/A 0.03fF
C35285 PAND2X1_773/CTRL2 POR2X1_767/Y 0.01fF
C35286 POR2X1_35/Y POR2X1_632/Y 0.04fF
C35287 POR2X1_273/CTRL POR2X1_273/O -0.00fF
C35288 POR2X1_239/Y PAND2X1_506/Y 0.10fF
C35289 PAND2X1_182/B PAND2X1_336/a_16_344# 0.02fF
C35290 PAND2X1_482/CTRL2 POR2X1_260/A 0.01fF
C35291 POR2X1_7/Y PAND2X1_656/A 0.15fF
C35292 VDD POR2X1_303/B 0.04fF
C35293 POR2X1_23/Y POR2X1_253/O 0.02fF
C35294 POR2X1_48/A POR2X1_253/CTRL 0.01fF
C35295 PAND2X1_726/B POR2X1_394/A 0.07fF
C35296 POR2X1_444/A POR2X1_444/a_56_344# 0.00fF
C35297 PAND2X1_126/a_16_344# POR2X1_62/Y 0.01fF
C35298 POR2X1_73/Y PAND2X1_169/CTRL 0.01fF
C35299 POR2X1_566/A POR2X1_863/A 0.07fF
C35300 POR2X1_38/Y PAND2X1_379/O 0.01fF
C35301 POR2X1_485/Y POR2X1_669/B 0.07fF
C35302 POR2X1_688/CTRL POR2X1_121/B 0.25fF
C35303 POR2X1_640/Y POR2X1_814/A 0.01fF
C35304 PAND2X1_206/B POR2X1_94/A 0.16fF
C35305 PAND2X1_341/A PAND2X1_358/O 0.03fF
C35306 POR2X1_35/Y PAND2X1_52/B 0.05fF
C35307 PAND2X1_432/a_16_344# POR2X1_648/Y 0.01fF
C35308 POR2X1_638/B PAND2X1_72/A 0.11fF
C35309 POR2X1_16/A PAND2X1_659/Y 0.12fF
C35310 POR2X1_715/CTRL2 POR2X1_702/A 0.00fF
C35311 POR2X1_846/A VDD 0.15fF
C35312 POR2X1_38/Y POR2X1_522/CTRL 0.07fF
C35313 POR2X1_814/A POR2X1_778/CTRL2 0.01fF
C35314 POR2X1_16/A POR2X1_96/Y 0.03fF
C35315 POR2X1_570/B PAND2X1_72/A 0.03fF
C35316 PAND2X1_811/A PAND2X1_287/Y 0.03fF
C35317 POR2X1_445/A POR2X1_78/A 0.03fF
C35318 PAND2X1_207/CTRL2 POR2X1_32/A 0.01fF
C35319 PAND2X1_652/O PAND2X1_593/Y 0.05fF
C35320 POR2X1_234/A POR2X1_519/Y 0.02fF
C35321 POR2X1_77/CTRL POR2X1_83/B 0.01fF
C35322 POR2X1_123/B PAND2X1_72/A 0.02fF
C35323 POR2X1_643/CTRL2 PAND2X1_55/Y 0.03fF
C35324 POR2X1_737/A PAND2X1_48/A 0.12fF
C35325 PAND2X1_86/CTRL VDD 0.00fF
C35326 POR2X1_431/m4_208_n4# POR2X1_5/Y 0.05fF
C35327 POR2X1_250/Y PAND2X1_740/Y 0.15fF
C35328 POR2X1_423/Y POR2X1_253/CTRL2 0.01fF
C35329 POR2X1_257/A PAND2X1_541/CTRL2 0.01fF
C35330 POR2X1_78/B PAND2X1_418/O 0.11fF
C35331 POR2X1_54/Y POR2X1_104/a_16_28# 0.03fF
C35332 POR2X1_707/O D_INPUT_4 0.01fF
C35333 POR2X1_814/A POR2X1_121/Y 1.70fF
C35334 POR2X1_123/A PAND2X1_52/B 0.04fF
C35335 POR2X1_67/Y PAND2X1_754/CTRL 0.00fF
C35336 POR2X1_554/B POR2X1_217/O 0.01fF
C35337 POR2X1_376/B PAND2X1_98/O 0.03fF
C35338 POR2X1_807/O POR2X1_590/A 0.01fF
C35339 PAND2X1_272/CTRL2 POR2X1_296/B 0.03fF
C35340 POR2X1_48/A POR2X1_516/Y 0.01fF
C35341 POR2X1_98/CTRL POR2X1_590/A 0.01fF
C35342 POR2X1_660/O D_INPUT_0 0.03fF
C35343 PAND2X1_639/a_16_344# POR2X1_408/Y 0.08fF
C35344 POR2X1_705/B VDD 0.00fF
C35345 POR2X1_294/A PAND2X1_122/CTRL 0.24fF
C35346 POR2X1_433/CTRL POR2X1_37/Y 0.01fF
C35347 POR2X1_341/A POR2X1_573/a_56_344# 0.01fF
C35348 PAND2X1_255/CTRL POR2X1_786/Y 0.05fF
C35349 POR2X1_260/B PAND2X1_41/B 0.13fF
C35350 POR2X1_62/Y PAND2X1_529/CTRL2 0.03fF
C35351 POR2X1_848/A POR2X1_752/Y 0.06fF
C35352 POR2X1_556/A POR2X1_76/Y 0.03fF
C35353 POR2X1_77/Y PAND2X1_337/O 0.03fF
C35354 POR2X1_294/Y POR2X1_330/Y 0.07fF
C35355 PAND2X1_675/A POR2X1_250/Y 0.15fF
C35356 POR2X1_624/Y PAND2X1_8/Y 0.03fF
C35357 POR2X1_525/CTRL POR2X1_23/Y 0.03fF
C35358 POR2X1_66/A POR2X1_200/a_16_28# 0.03fF
C35359 POR2X1_37/Y PAND2X1_500/O 0.00fF
C35360 PAND2X1_458/CTRL POR2X1_91/Y 0.03fF
C35361 POR2X1_257/A PAND2X1_785/Y 2.48fF
C35362 POR2X1_329/A POR2X1_816/A 0.03fF
C35363 POR2X1_227/CTRL2 PAND2X1_52/B 0.03fF
C35364 POR2X1_150/Y POR2X1_494/Y 0.00fF
C35365 PAND2X1_137/a_16_344# POR2X1_20/B 0.01fF
C35366 POR2X1_48/A PAND2X1_738/O 0.01fF
C35367 POR2X1_63/Y POR2X1_406/O 0.01fF
C35368 PAND2X1_205/A PAND2X1_473/B 0.05fF
C35369 POR2X1_306/CTRL2 POR2X1_329/A 0.03fF
C35370 POR2X1_556/A POR2X1_740/Y 4.29fF
C35371 POR2X1_636/CTRL2 POR2X1_750/B 0.01fF
C35372 POR2X1_376/B PAND2X1_68/CTRL 0.02fF
C35373 PAND2X1_841/CTRL POR2X1_411/B 0.01fF
C35374 POR2X1_68/A POR2X1_66/O 0.02fF
C35375 POR2X1_841/CTRL POR2X1_733/A 0.07fF
C35376 POR2X1_49/Y POR2X1_753/Y 0.07fF
C35377 PAND2X1_818/a_16_344# PAND2X1_340/B 0.01fF
C35378 POR2X1_515/O PAND2X1_93/B 0.03fF
C35379 PAND2X1_797/Y POR2X1_39/B 0.03fF
C35380 POR2X1_16/A PAND2X1_403/CTRL2 0.01fF
C35381 POR2X1_476/Y PAND2X1_595/CTRL 0.01fF
C35382 POR2X1_306/Y POR2X1_102/Y 0.01fF
C35383 POR2X1_102/Y PAND2X1_140/O 0.07fF
C35384 PAND2X1_742/CTRL2 POR2X1_331/Y 0.03fF
C35385 POR2X1_411/B PAND2X1_398/O 0.02fF
C35386 POR2X1_68/A POR2X1_541/B 0.10fF
C35387 POR2X1_366/Y PAND2X1_268/O 0.03fF
C35388 PAND2X1_244/O POR2X1_72/B 0.01fF
C35389 PAND2X1_105/O POR2X1_411/B 0.02fF
C35390 POR2X1_13/A PAND2X1_99/B 0.61fF
C35391 POR2X1_621/B POR2X1_296/B 0.01fF
C35392 POR2X1_487/CTRL2 PAND2X1_580/B 0.00fF
C35393 POR2X1_274/A PAND2X1_516/a_56_28# 0.00fF
C35394 POR2X1_476/A PAND2X1_57/B 0.03fF
C35395 POR2X1_67/Y POR2X1_7/A 0.03fF
C35396 POR2X1_12/A POR2X1_587/CTRL 0.00fF
C35397 POR2X1_94/A POR2X1_750/B 0.07fF
C35398 PAND2X1_66/a_16_344# POR2X1_7/B 0.02fF
C35399 POR2X1_624/Y PAND2X1_316/CTRL2 0.01fF
C35400 POR2X1_502/A POR2X1_220/B 0.03fF
C35401 POR2X1_60/A PAND2X1_513/a_76_28# 0.02fF
C35402 POR2X1_257/A PAND2X1_324/CTRL2 0.00fF
C35403 POR2X1_633/A PAND2X1_90/Y 0.03fF
C35404 PAND2X1_39/B PAND2X1_29/O 0.01fF
C35405 POR2X1_149/CTRL2 POR2X1_532/A 0.01fF
C35406 POR2X1_197/O POR2X1_555/B 0.02fF
C35407 PAND2X1_20/A POR2X1_401/CTRL2 0.01fF
C35408 PAND2X1_76/O PAND2X1_76/Y 0.00fF
C35409 POR2X1_188/A POR2X1_710/A 0.05fF
C35410 POR2X1_260/B POR2X1_130/Y 0.02fF
C35411 POR2X1_313/Y PAND2X1_439/CTRL2 0.01fF
C35412 POR2X1_502/A POR2X1_660/Y 0.03fF
C35413 POR2X1_106/Y POR2X1_40/Y 0.03fF
C35414 POR2X1_489/B VDD 0.02fF
C35415 PAND2X1_411/CTRL POR2X1_260/B 0.01fF
C35416 POR2X1_141/a_76_344# PAND2X1_20/A 0.00fF
C35417 POR2X1_630/CTRL2 POR2X1_222/Y 0.10fF
C35418 PAND2X1_644/Y POR2X1_755/O 0.09fF
C35419 PAND2X1_651/Y PAND2X1_436/CTRL2 0.05fF
C35420 PAND2X1_272/CTRL POR2X1_465/B 0.04fF
C35421 POR2X1_23/Y PAND2X1_575/A 0.62fF
C35422 PAND2X1_862/B POR2X1_498/Y 0.03fF
C35423 POR2X1_114/B POR2X1_866/A 0.59fF
C35424 PAND2X1_70/CTRL POR2X1_750/B 0.01fF
C35425 POR2X1_102/Y PAND2X1_719/O 0.02fF
C35426 POR2X1_227/A POR2X1_854/B 0.31fF
C35427 PAND2X1_777/O POR2X1_293/Y 0.16fF
C35428 PAND2X1_462/B POR2X1_37/Y 0.08fF
C35429 PAND2X1_284/Y PAND2X1_562/Y 0.68fF
C35430 POR2X1_814/B POR2X1_439/Y 0.02fF
C35431 PAND2X1_58/A POR2X1_608/a_16_28# 0.02fF
C35432 POR2X1_186/Y PAND2X1_90/Y 0.11fF
C35433 POR2X1_278/Y POR2X1_60/A 0.12fF
C35434 POR2X1_318/a_16_28# POR2X1_318/A 0.03fF
C35435 PAND2X1_20/A POR2X1_192/Y 0.05fF
C35436 POR2X1_849/B POR2X1_790/A 0.02fF
C35437 POR2X1_20/B PAND2X1_121/CTRL2 0.01fF
C35438 PAND2X1_413/CTRL2 POR2X1_814/A 0.01fF
C35439 POR2X1_605/B VDD 0.02fF
C35440 POR2X1_590/A POR2X1_578/Y 0.95fF
C35441 POR2X1_23/Y PAND2X1_794/B 0.34fF
C35442 PAND2X1_717/A PAND2X1_112/a_76_28# 0.02fF
C35443 POR2X1_207/CTRL POR2X1_330/Y 0.03fF
C35444 POR2X1_202/CTRL2 VDD 0.00fF
C35445 POR2X1_40/Y PAND2X1_580/B 0.03fF
C35446 PAND2X1_20/A POR2X1_785/O 0.07fF
C35447 PAND2X1_340/B PAND2X1_509/O -0.00fF
C35448 PAND2X1_485/O POR2X1_789/A 0.01fF
C35449 POR2X1_780/CTRL VDD 0.00fF
C35450 PAND2X1_287/a_76_28# PAND2X1_771/Y 0.02fF
C35451 POR2X1_828/Y PAND2X1_65/B 1.63fF
C35452 POR2X1_48/A PAND2X1_506/a_56_28# 0.00fF
C35453 PAND2X1_404/Y POR2X1_38/Y 0.07fF
C35454 POR2X1_274/A POR2X1_573/A 0.03fF
C35455 POR2X1_51/A POR2X1_750/B 0.03fF
C35456 POR2X1_604/Y POR2X1_42/Y 0.01fF
C35457 PAND2X1_669/CTRL2 POR2X1_816/A 0.01fF
C35458 POR2X1_677/CTRL2 INPUT_0 0.09fF
C35459 PAND2X1_480/B PAND2X1_558/Y 0.03fF
C35460 PAND2X1_473/Y PAND2X1_576/CTRL 0.01fF
C35461 POR2X1_96/B POR2X1_54/Y 0.05fF
C35462 POR2X1_192/Y POR2X1_776/CTRL2 0.01fF
C35463 POR2X1_333/A PAND2X1_23/Y 0.05fF
C35464 POR2X1_137/B POR2X1_260/A 0.07fF
C35465 POR2X1_814/B POR2X1_572/CTRL 0.14fF
C35466 INPUT_1 PAND2X1_247/CTRL2 0.01fF
C35467 POR2X1_48/A POR2X1_280/CTRL2 0.01fF
C35468 POR2X1_66/B PAND2X1_376/m4_208_n4# 0.22fF
C35469 PAND2X1_420/a_16_344# POR2X1_785/A 0.02fF
C35470 POR2X1_88/CTRL POR2X1_7/A 0.01fF
C35471 PAND2X1_20/A POR2X1_574/CTRL2 0.01fF
C35472 PAND2X1_832/a_76_28# PAND2X1_499/Y 0.01fF
C35473 POR2X1_260/B POR2X1_228/Y 0.01fF
C35474 INPUT_3 POR2X1_376/CTRL2 0.05fF
C35475 POR2X1_48/A PAND2X1_702/O 0.04fF
C35476 PAND2X1_840/B POR2X1_83/B 0.01fF
C35477 POR2X1_814/B POR2X1_192/Y 0.10fF
C35478 POR2X1_152/O POR2X1_669/B 0.06fF
C35479 POR2X1_358/a_16_28# PAND2X1_20/A 0.01fF
C35480 POR2X1_832/m4_208_n4# POR2X1_330/Y 0.06fF
C35481 POR2X1_805/O PAND2X1_60/B 0.01fF
C35482 PAND2X1_56/Y POR2X1_850/B 0.03fF
C35483 POR2X1_290/CTRL2 POR2X1_290/Y 0.02fF
C35484 POR2X1_779/A POR2X1_121/B 0.03fF
C35485 PAND2X1_460/Y POR2X1_5/Y 0.39fF
C35486 POR2X1_549/B VDD 0.04fF
C35487 PAND2X1_272/O PAND2X1_32/B 0.03fF
C35488 POR2X1_407/A POR2X1_390/CTRL 0.00fF
C35489 PAND2X1_638/B PAND2X1_638/O 0.00fF
C35490 PAND2X1_627/CTRL VDD 0.00fF
C35491 POR2X1_322/CTRL POR2X1_72/B 0.01fF
C35492 POR2X1_866/O POR2X1_800/A 0.01fF
C35493 POR2X1_477/A POR2X1_675/a_76_344# 0.01fF
C35494 POR2X1_461/B VDD 0.17fF
C35495 POR2X1_66/B POR2X1_68/A 0.11fF
C35496 PAND2X1_39/O PAND2X1_69/A 0.15fF
C35497 PAND2X1_557/A PAND2X1_798/B 0.09fF
C35498 PAND2X1_23/Y POR2X1_734/A 0.10fF
C35499 PAND2X1_55/Y PAND2X1_41/B 0.23fF
C35500 POR2X1_567/B PAND2X1_173/a_76_28# 0.05fF
C35501 POR2X1_496/Y POR2X1_93/A 0.07fF
C35502 PAND2X1_275/CTRL2 POR2X1_274/Y 0.01fF
C35503 POR2X1_257/A PAND2X1_348/A 0.03fF
C35504 POR2X1_240/B POR2X1_68/B 0.02fF
C35505 POR2X1_66/A POR2X1_510/Y 0.13fF
C35506 POR2X1_45/Y PAND2X1_217/B 0.20fF
C35507 POR2X1_465/A VDD -0.00fF
C35508 POR2X1_41/B PAND2X1_723/Y 0.03fF
C35509 POR2X1_65/A POR2X1_42/Y 0.23fF
C35510 POR2X1_634/A POR2X1_771/CTRL 0.07fF
C35511 INPUT_2 POR2X1_60/A 0.00fF
C35512 PAND2X1_279/m4_208_n4# POR2X1_740/Y 0.06fF
C35513 POR2X1_270/Y PAND2X1_368/CTRL2 0.00fF
C35514 PAND2X1_635/CTRL POR2X1_748/A 0.01fF
C35515 POR2X1_188/A POR2X1_68/A 0.05fF
C35516 PAND2X1_137/Y PAND2X1_140/Y 0.03fF
C35517 PAND2X1_214/a_56_28# PAND2X1_656/A 0.00fF
C35518 POR2X1_40/Y PAND2X1_337/A 0.08fF
C35519 POR2X1_262/Y PAND2X1_716/B 0.03fF
C35520 PAND2X1_831/O POR2X1_273/Y 0.02fF
C35521 POR2X1_57/A PAND2X1_219/A 0.24fF
C35522 POR2X1_48/A PAND2X1_114/CTRL 0.01fF
C35523 PAND2X1_776/m4_208_n4# POR2X1_20/B 0.10fF
C35524 PAND2X1_781/Y POR2X1_747/Y 0.00fF
C35525 POR2X1_231/A POR2X1_795/B 0.08fF
C35526 POR2X1_505/CTRL2 POR2X1_48/A 0.01fF
C35527 POR2X1_113/Y POR2X1_78/A 0.03fF
C35528 POR2X1_66/B POR2X1_460/A 2.68fF
C35529 POR2X1_313/Y POR2X1_438/Y 0.00fF
C35530 PAND2X1_93/B POR2X1_260/A 0.13fF
C35531 PAND2X1_35/A POR2X1_394/A 0.08fF
C35532 POR2X1_102/Y POR2X1_142/Y 3.27fF
C35533 POR2X1_853/A PAND2X1_65/B 0.03fF
C35534 POR2X1_477/A POR2X1_480/A 0.08fF
C35535 POR2X1_693/Y POR2X1_376/B 0.02fF
C35536 PAND2X1_74/O POR2X1_532/A 0.04fF
C35537 POR2X1_673/O POR2X1_38/B 0.02fF
C35538 PAND2X1_404/Y POR2X1_153/Y 0.12fF
C35539 POR2X1_663/B POR2X1_337/Y 0.07fF
C35540 POR2X1_81/Y PAND2X1_735/Y 0.06fF
C35541 POR2X1_72/Y PAND2X1_659/B 0.25fF
C35542 POR2X1_121/A PAND2X1_90/Y 0.02fF
C35543 PAND2X1_785/Y PAND2X1_553/B 0.05fF
C35544 POR2X1_102/Y PAND2X1_175/B 3.56fF
C35545 POR2X1_150/Y PAND2X1_352/Y 0.00fF
C35546 POR2X1_56/B POR2X1_13/A 0.01fF
C35547 POR2X1_16/A POR2X1_37/Y 0.10fF
C35548 POR2X1_524/Y PAND2X1_324/Y 0.02fF
C35549 POR2X1_447/B PAND2X1_43/O 0.09fF
C35550 POR2X1_110/a_16_28# POR2X1_73/Y 0.00fF
C35551 PAND2X1_65/B POR2X1_391/Y 0.14fF
C35552 POR2X1_817/CTRL POR2X1_394/A 0.07fF
C35553 POR2X1_407/Y PAND2X1_41/B 0.04fF
C35554 POR2X1_16/A PAND2X1_561/CTRL 0.10fF
C35555 PAND2X1_564/B POR2X1_765/Y 0.00fF
C35556 POR2X1_40/Y POR2X1_511/CTRL 0.01fF
C35557 POR2X1_558/CTRL INPUT_0 0.07fF
C35558 POR2X1_606/CTRL2 POR2X1_294/A 0.09fF
C35559 POR2X1_606/CTRL PAND2X1_48/A 0.01fF
C35560 POR2X1_280/CTRL POR2X1_312/Y 0.01fF
C35561 POR2X1_5/Y POR2X1_52/Y 0.02fF
C35562 POR2X1_69/A POR2X1_408/Y 0.05fF
C35563 PAND2X1_96/CTRL2 PAND2X1_60/B 0.01fF
C35564 PAND2X1_93/B POR2X1_363/A 0.07fF
C35565 POR2X1_45/Y VDD 1.00fF
C35566 PAND2X1_762/Y VDD 0.12fF
C35567 POR2X1_517/O POR2X1_73/Y 0.03fF
C35568 PAND2X1_631/A POR2X1_257/A 0.07fF
C35569 POR2X1_580/O D_GATE_741 0.34fF
C35570 PAND2X1_89/CTRL POR2X1_785/A 0.00fF
C35571 POR2X1_529/m4_208_n4# POR2X1_5/Y 0.03fF
C35572 POR2X1_120/O POR2X1_712/Y 0.02fF
C35573 POR2X1_66/B POR2X1_21/a_16_28# 0.04fF
C35574 PAND2X1_20/A POR2X1_785/B 0.01fF
C35575 PAND2X1_349/A POR2X1_40/Y 0.03fF
C35576 POR2X1_302/Y POR2X1_114/B 0.01fF
C35577 POR2X1_78/A POR2X1_260/A 0.07fF
C35578 PAND2X1_63/B POR2X1_40/Y 0.11fF
C35579 PAND2X1_462/B POR2X1_293/Y 0.16fF
C35580 POR2X1_68/A POR2X1_859/A 0.01fF
C35581 POR2X1_455/A POR2X1_220/Y 0.06fF
C35582 POR2X1_49/Y PAND2X1_656/A 0.06fF
C35583 PAND2X1_793/Y PAND2X1_652/A 0.01fF
C35584 POR2X1_599/A POR2X1_46/Y 0.09fF
C35585 PAND2X1_65/B POR2X1_712/CTRL2 0.01fF
C35586 PAND2X1_20/A POR2X1_546/CTRL2 0.01fF
C35587 POR2X1_115/CTRL2 POR2X1_804/A 0.12fF
C35588 POR2X1_8/Y POR2X1_104/CTRL 0.01fF
C35589 PAND2X1_57/B PAND2X1_743/CTRL2 0.00fF
C35590 POR2X1_52/A POR2X1_693/Y 0.03fF
C35591 PAND2X1_491/O INPUT_0 0.12fF
C35592 POR2X1_57/A POR2X1_135/Y 0.46fF
C35593 PAND2X1_20/A POR2X1_571/CTRL2 0.01fF
C35594 POR2X1_633/CTRL PAND2X1_52/B 0.09fF
C35595 POR2X1_462/B POR2X1_790/CTRL2 0.01fF
C35596 POR2X1_327/Y POR2X1_590/A 0.16fF
C35597 POR2X1_196/Y POR2X1_215/O 0.06fF
C35598 POR2X1_23/Y POR2X1_373/O 0.02fF
C35599 POR2X1_390/m4_208_n4# POR2X1_260/A 0.01fF
C35600 PAND2X1_738/Y PAND2X1_113/CTRL 0.01fF
C35601 POR2X1_628/Y POR2X1_39/B 0.07fF
C35602 POR2X1_135/CTRL POR2X1_48/A 0.01fF
C35603 PAND2X1_778/CTRL POR2X1_387/Y 0.07fF
C35604 POR2X1_72/B PAND2X1_737/B 0.03fF
C35605 POR2X1_198/O POR2X1_198/B 0.01fF
C35606 POR2X1_78/B POR2X1_318/A 0.36fF
C35607 PAND2X1_57/B POR2X1_770/O 0.18fF
C35608 POR2X1_86/Y POR2X1_20/B 0.03fF
C35609 POR2X1_83/B PAND2X1_853/B 0.00fF
C35610 POR2X1_78/A PAND2X1_142/O 0.03fF
C35611 PAND2X1_665/O POR2X1_260/B 0.02fF
C35612 PAND2X1_770/a_76_28# POR2X1_73/Y 0.01fF
C35613 PAND2X1_216/B POR2X1_72/B 0.03fF
C35614 PAND2X1_190/Y POR2X1_42/Y 0.05fF
C35615 POR2X1_511/Y PAND2X1_549/B 0.03fF
C35616 POR2X1_396/Y VDD 0.10fF
C35617 POR2X1_137/CTRL PAND2X1_32/B 0.01fF
C35618 PAND2X1_773/a_16_344# POR2X1_7/B 0.02fF
C35619 PAND2X1_797/Y POR2X1_48/A 0.03fF
C35620 POR2X1_43/B POR2X1_277/a_76_344# 0.03fF
C35621 PAND2X1_73/Y PAND2X1_527/O 0.07fF
C35622 POR2X1_557/A PAND2X1_42/O 0.01fF
C35623 POR2X1_498/Y PAND2X1_716/B 0.03fF
C35624 POR2X1_334/CTRL POR2X1_814/B 0.00fF
C35625 PAND2X1_48/B POR2X1_804/A 0.03fF
C35626 PAND2X1_23/Y POR2X1_786/Y 0.07fF
C35627 POR2X1_271/CTRL POR2X1_39/B 0.01fF
C35628 POR2X1_237/Y POR2X1_238/Y 0.01fF
C35629 POR2X1_283/A PAND2X1_362/B 0.03fF
C35630 POR2X1_178/CTRL PAND2X1_675/A 0.09fF
C35631 POR2X1_855/B VDD 0.70fF
C35632 POR2X1_717/CTRL2 POR2X1_717/Y 0.01fF
C35633 POR2X1_834/Y PAND2X1_65/B 0.05fF
C35634 POR2X1_523/Y POR2X1_790/A 0.02fF
C35635 POR2X1_356/A POR2X1_220/A 0.03fF
C35636 POR2X1_333/Y PAND2X1_41/B 0.03fF
C35637 POR2X1_334/Y POR2X1_750/B 0.10fF
C35638 POR2X1_383/A POR2X1_483/CTRL 0.05fF
C35639 PAND2X1_57/B POR2X1_366/A 0.01fF
C35640 PAND2X1_651/Y POR2X1_521/CTRL2 0.06fF
C35641 POR2X1_635/A PAND2X1_52/B 0.01fF
C35642 POR2X1_460/B PAND2X1_69/A 0.00fF
C35643 POR2X1_802/O POR2X1_220/Y 0.06fF
C35644 POR2X1_775/A PAND2X1_96/B 0.03fF
C35645 VDD POR2X1_171/O 0.00fF
C35646 PAND2X1_532/CTRL2 VDD 0.00fF
C35647 POR2X1_236/Y POR2X1_172/a_16_28# 0.03fF
C35648 PAND2X1_793/Y POR2X1_437/CTRL2 0.01fF
C35649 POR2X1_188/a_76_344# POR2X1_220/Y 0.01fF
C35650 POR2X1_110/Y PAND2X1_465/CTRL 0.00fF
C35651 POR2X1_537/Y POR2X1_794/B 0.04fF
C35652 POR2X1_572/B POR2X1_361/CTRL2 0.01fF
C35653 POR2X1_790/A PAND2X1_69/A 0.03fF
C35654 PAND2X1_46/O POR2X1_294/A 0.02fF
C35655 PAND2X1_844/B POR2X1_521/CTRL2 0.01fF
C35656 POR2X1_135/Y POR2X1_111/Y 0.28fF
C35657 POR2X1_288/A POR2X1_737/A 0.02fF
C35658 PAND2X1_55/Y POR2X1_228/Y 0.10fF
C35659 PAND2X1_514/Y POR2X1_91/Y 0.03fF
C35660 POR2X1_130/CTRL VDD 0.00fF
C35661 PAND2X1_116/O PAND2X1_853/B 0.02fF
C35662 POR2X1_389/Y POR2X1_294/A 0.02fF
C35663 POR2X1_356/A POR2X1_569/A 0.10fF
C35664 POR2X1_426/O POR2X1_425/Y 0.01fF
C35665 POR2X1_502/A POR2X1_308/B 0.03fF
C35666 PAND2X1_372/O POR2X1_101/Y 0.02fF
C35667 POR2X1_741/Y POR2X1_702/CTRL 0.00fF
C35668 POR2X1_740/Y POR2X1_702/O 0.06fF
C35669 POR2X1_135/CTRL2 POR2X1_423/Y 0.01fF
C35670 POR2X1_859/A POR2X1_391/B 0.02fF
C35671 PAND2X1_291/CTRL POR2X1_35/Y 0.03fF
C35672 POR2X1_483/A POR2X1_186/B 0.01fF
C35673 PAND2X1_96/B POR2X1_112/Y 0.03fF
C35674 POR2X1_765/a_16_28# POR2X1_73/Y 0.09fF
C35675 POR2X1_222/Y POR2X1_510/Y 0.03fF
C35676 POR2X1_57/A POR2X1_816/A 5.35fF
C35677 POR2X1_219/CTRL2 PAND2X1_88/Y 0.01fF
C35678 PAND2X1_140/Y PAND2X1_853/B 0.03fF
C35679 POR2X1_43/B PAND2X1_469/Y 0.01fF
C35680 POR2X1_865/B PAND2X1_69/A 0.07fF
C35681 PAND2X1_69/A PAND2X1_88/Y 0.03fF
C35682 POR2X1_294/B PAND2X1_528/O 0.03fF
C35683 POR2X1_84/Y PAND2X1_69/A 0.00fF
C35684 POR2X1_86/CTRL2 POR2X1_40/Y 0.02fF
C35685 POR2X1_16/A POR2X1_293/Y 0.17fF
C35686 POR2X1_371/O POR2X1_5/Y 0.02fF
C35687 POR2X1_371/CTRL2 POR2X1_372/A 0.01fF
C35688 POR2X1_564/B VDD 0.02fF
C35689 PAND2X1_209/A PAND2X1_213/Y 0.01fF
C35690 POR2X1_192/Y POR2X1_192/a_16_28# 0.01fF
C35691 POR2X1_16/A PAND2X1_555/A 0.03fF
C35692 D_INPUT_0 POR2X1_717/B 0.03fF
C35693 POR2X1_702/CTRL PAND2X1_32/B 0.01fF
C35694 POR2X1_564/Y POR2X1_317/B 0.03fF
C35695 PAND2X1_800/O POR2X1_96/A 0.05fF
C35696 PAND2X1_442/CTRL POR2X1_191/Y 0.00fF
C35697 PAND2X1_725/B PAND2X1_725/a_76_28# 0.04fF
C35698 PAND2X1_25/CTRL PAND2X1_72/A 0.00fF
C35699 POR2X1_857/a_16_28# POR2X1_568/B 0.03fF
C35700 POR2X1_477/Y POR2X1_568/A 0.00fF
C35701 POR2X1_855/B POR2X1_796/a_56_344# 0.00fF
C35702 POR2X1_78/CTRL POR2X1_569/A 0.04fF
C35703 PAND2X1_60/B POR2X1_140/CTRL 0.01fF
C35704 POR2X1_537/Y PAND2X1_108/O 0.02fF
C35705 POR2X1_108/O POR2X1_142/Y 0.00fF
C35706 POR2X1_567/A POR2X1_663/O 0.30fF
C35707 POR2X1_41/B PAND2X1_123/Y 0.04fF
C35708 POR2X1_855/B PAND2X1_32/B 0.02fF
C35709 POR2X1_532/A POR2X1_510/Y 0.06fF
C35710 POR2X1_7/B PAND2X1_507/a_16_344# 0.02fF
C35711 POR2X1_96/A PAND2X1_538/O 0.05fF
C35712 PAND2X1_217/CTRL2 PAND2X1_656/A 0.01fF
C35713 POR2X1_57/A PAND2X1_854/A 0.02fF
C35714 POR2X1_814/A PAND2X1_268/CTRL2 0.03fF
C35715 PAND2X1_298/CTRL2 PAND2X1_32/B 0.01fF
C35716 INPUT_5 PAND2X1_3/B 0.82fF
C35717 PAND2X1_65/B POR2X1_383/Y 0.03fF
C35718 PAND2X1_349/A PAND2X1_840/CTRL2 0.01fF
C35719 POR2X1_763/Y POR2X1_320/CTRL2 0.05fF
C35720 POR2X1_187/Y POR2X1_79/Y 0.01fF
C35721 PAND2X1_476/A PAND2X1_673/Y 0.04fF
C35722 POR2X1_532/A POR2X1_520/O 0.01fF
C35723 POR2X1_43/B POR2X1_394/A 0.22fF
C35724 POR2X1_96/A PAND2X1_802/a_16_344# 0.01fF
C35725 PAND2X1_322/CTRL POR2X1_188/Y 0.00fF
C35726 PAND2X1_39/B POR2X1_646/B 0.02fF
C35727 POR2X1_318/A POR2X1_141/A 0.03fF
C35728 POR2X1_661/O POR2X1_711/Y 0.04fF
C35729 PAND2X1_65/B POR2X1_779/CTRL 0.01fF
C35730 PAND2X1_844/Y PAND2X1_338/CTRL2 0.01fF
C35731 POR2X1_66/B POR2X1_138/A 0.04fF
C35732 POR2X1_337/A POR2X1_228/Y 0.01fF
C35733 POR2X1_197/Y POR2X1_215/A 0.07fF
C35734 PAND2X1_863/A PAND2X1_863/B 0.15fF
C35735 POR2X1_462/B POR2X1_559/A 0.06fF
C35736 POR2X1_68/B POR2X1_768/O 0.01fF
C35737 POR2X1_738/A POR2X1_854/B 0.03fF
C35738 POR2X1_713/CTRL PAND2X1_48/A 0.01fF
C35739 POR2X1_118/O POR2X1_153/Y 0.05fF
C35740 PAND2X1_508/Y POR2X1_56/Y 0.02fF
C35741 PAND2X1_824/B PAND2X1_88/Y 0.07fF
C35742 PAND2X1_347/Y POR2X1_77/Y 0.03fF
C35743 POR2X1_38/B POR2X1_394/A 0.02fF
C35744 PAND2X1_7/CTRL POR2X1_99/B 0.00fF
C35745 POR2X1_567/A POR2X1_563/Y 0.01fF
C35746 POR2X1_16/A POR2X1_408/Y 0.03fF
C35747 PAND2X1_23/Y PAND2X1_396/O 0.10fF
C35748 POR2X1_751/Y POR2X1_382/Y 0.00fF
C35749 PAND2X1_793/Y POR2X1_184/CTRL 0.01fF
C35750 PAND2X1_18/CTRL PAND2X1_52/B 0.13fF
C35751 POR2X1_42/Y POR2X1_397/a_16_28# 0.02fF
C35752 POR2X1_68/B PAND2X1_531/CTRL 0.01fF
C35753 POR2X1_110/Y POR2X1_368/Y 0.01fF
C35754 POR2X1_648/Y POR2X1_807/CTRL2 0.03fF
C35755 PAND2X1_33/O POR2X1_24/Y 0.12fF
C35756 POR2X1_383/A PAND2X1_298/O 0.05fF
C35757 POR2X1_569/A POR2X1_570/Y 0.36fF
C35758 POR2X1_41/O PAND2X1_656/A 0.01fF
C35759 POR2X1_809/A POR2X1_788/B 0.02fF
C35760 POR2X1_327/Y POR2X1_361/CTRL 0.01fF
C35761 PAND2X1_586/CTRL2 PAND2X1_60/B 0.01fF
C35762 PAND2X1_687/O PAND2X1_643/Y 0.05fF
C35763 POR2X1_508/A PAND2X1_69/A 0.03fF
C35764 PAND2X1_90/CTRL2 POR2X1_68/B 0.01fF
C35765 POR2X1_557/B PAND2X1_60/B 0.03fF
C35766 POR2X1_75/Y POR2X1_91/Y 0.03fF
C35767 POR2X1_49/Y PAND2X1_193/Y 0.03fF
C35768 POR2X1_48/A PAND2X1_35/a_56_28# 0.00fF
C35769 POR2X1_283/A PAND2X1_502/CTRL2 0.03fF
C35770 POR2X1_490/Y POR2X1_262/Y 0.03fF
C35771 POR2X1_333/CTRL2 POR2X1_333/Y 0.00fF
C35772 POR2X1_735/CTRL POR2X1_318/A 0.06fF
C35773 POR2X1_129/Y PAND2X1_549/B 0.03fF
C35774 PAND2X1_96/B PAND2X1_134/CTRL2 0.01fF
C35775 POR2X1_153/Y PAND2X1_123/CTRL2 0.05fF
C35776 POR2X1_294/A POR2X1_318/A 0.07fF
C35777 POR2X1_9/Y POR2X1_750/A 0.02fF
C35778 POR2X1_574/Y POR2X1_141/A 0.03fF
C35779 PAND2X1_148/O POR2X1_146/Y 0.00fF
C35780 POR2X1_555/A PAND2X1_628/CTRL2 0.02fF
C35781 POR2X1_22/A POR2X1_39/B 0.10fF
C35782 POR2X1_519/Y POR2X1_39/B 0.01fF
C35783 POR2X1_646/B POR2X1_805/Y 0.27fF
C35784 POR2X1_76/B POR2X1_325/A 0.12fF
C35785 POR2X1_333/Y POR2X1_502/CTRL 0.00fF
C35786 POR2X1_647/B POR2X1_862/A 0.05fF
C35787 POR2X1_119/Y POR2X1_387/Y 0.07fF
C35788 PAND2X1_812/A PAND2X1_811/Y 0.32fF
C35789 POR2X1_356/A PAND2X1_72/A 0.19fF
C35790 POR2X1_35/Y POR2X1_555/CTRL2 0.01fF
C35791 POR2X1_304/O POR2X1_90/Y 0.00fF
C35792 PAND2X1_69/A POR2X1_568/B 0.05fF
C35793 POR2X1_576/m4_208_n4# POR2X1_260/A 0.15fF
C35794 PAND2X1_251/a_16_344# PAND2X1_39/B 0.04fF
C35795 PAND2X1_6/Y POR2X1_736/A 0.05fF
C35796 POR2X1_709/B INPUT_1 0.02fF
C35797 POR2X1_66/O PAND2X1_58/A 0.27fF
C35798 POR2X1_730/Y PAND2X1_533/a_76_28# 0.02fF
C35799 POR2X1_96/B POR2X1_4/Y 0.00fF
C35800 POR2X1_316/CTRL2 POR2X1_129/Y 0.01fF
C35801 POR2X1_119/Y PAND2X1_121/O 0.18fF
C35802 PAND2X1_341/B PAND2X1_849/B 0.03fF
C35803 POR2X1_644/a_16_28# POR2X1_260/B 0.03fF
C35804 PAND2X1_65/B PAND2X1_255/a_16_344# 0.02fF
C35805 POR2X1_241/CTRL2 POR2X1_776/A 0.01fF
C35806 POR2X1_39/B POR2X1_9/O 0.03fF
C35807 POR2X1_474/CTRL POR2X1_556/A 0.01fF
C35808 POR2X1_415/A POR2X1_29/A 0.02fF
C35809 POR2X1_23/Y PAND2X1_124/Y 0.03fF
C35810 POR2X1_416/B PAND2X1_547/a_76_28# 0.00fF
C35811 PAND2X1_157/O PAND2X1_3/B 0.15fF
C35812 POR2X1_54/Y POR2X1_296/B 0.07fF
C35813 POR2X1_814/B POR2X1_646/B 0.06fF
C35814 PAND2X1_404/O POR2X1_411/B 0.03fF
C35815 POR2X1_567/A POR2X1_675/Y 0.03fF
C35816 PAND2X1_535/Y POR2X1_416/B 0.02fF
C35817 POR2X1_257/A PAND2X1_564/B 0.03fF
C35818 POR2X1_46/CTRL2 PAND2X1_9/Y 0.01fF
C35819 POR2X1_202/A POR2X1_296/B 0.32fF
C35820 POR2X1_362/A POR2X1_362/a_16_28# 0.05fF
C35821 POR2X1_66/B POR2X1_709/A 0.06fF
C35822 POR2X1_841/O POR2X1_330/Y 0.04fF
C35823 POR2X1_411/B POR2X1_268/Y 0.01fF
C35824 POR2X1_536/a_16_28# PAND2X1_643/A 0.07fF
C35825 PAND2X1_1/O D_INPUT_4 0.04fF
C35826 POR2X1_285/Y POR2X1_643/Y 0.02fF
C35827 POR2X1_567/A POR2X1_544/B 0.10fF
C35828 POR2X1_856/B POR2X1_466/A 0.12fF
C35829 PAND2X1_85/CTRL INPUT_0 0.00fF
C35830 PAND2X1_798/B PAND2X1_860/A 0.02fF
C35831 POR2X1_191/B POR2X1_191/Y 0.18fF
C35832 PAND2X1_313/CTRL POR2X1_169/A 0.01fF
C35833 PAND2X1_332/Y POR2X1_91/Y 21.92fF
C35834 PAND2X1_600/CTRL2 POR2X1_121/B 0.07fF
C35835 PAND2X1_93/B POR2X1_243/A 0.07fF
C35836 POR2X1_20/B INPUT_7 0.03fF
C35837 POR2X1_831/m4_208_n4# POR2X1_330/Y 0.06fF
C35838 PAND2X1_485/O POR2X1_590/A 0.03fF
C35839 POR2X1_663/B POR2X1_543/A 0.03fF
C35840 POR2X1_814/A POR2X1_489/A 0.01fF
C35841 POR2X1_707/B PAND2X1_762/O 0.02fF
C35842 POR2X1_187/Y PAND2X1_730/A 0.02fF
C35843 POR2X1_23/Y POR2X1_83/B 0.84fF
C35844 PAND2X1_175/B POR2X1_173/O 0.01fF
C35845 POR2X1_12/A POR2X1_698/O 0.07fF
C35846 POR2X1_37/CTRL POR2X1_612/Y 0.08fF
C35847 POR2X1_569/A PAND2X1_72/A 0.14fF
C35848 POR2X1_49/Y PAND2X1_217/m4_208_n4# 0.08fF
C35849 PAND2X1_48/A PAND2X1_304/CTRL2 0.06fF
C35850 POR2X1_346/A POR2X1_296/B 0.01fF
C35851 PAND2X1_201/CTRL POR2X1_88/Y 0.01fF
C35852 POR2X1_271/B VDD 0.04fF
C35853 PAND2X1_829/CTRL2 PAND2X1_73/Y 0.01fF
C35854 PAND2X1_404/A POR2X1_411/B 0.03fF
C35855 POR2X1_41/B POR2X1_846/Y 0.03fF
C35856 PAND2X1_698/O PAND2X1_52/B 0.07fF
C35857 POR2X1_463/Y PAND2X1_52/B 0.46fF
C35858 POR2X1_570/Y PAND2X1_72/A 0.01fF
C35859 POR2X1_120/O PAND2X1_39/B 0.20fF
C35860 POR2X1_416/B PAND2X1_507/O 0.06fF
C35861 POR2X1_661/A POR2X1_307/A 0.09fF
C35862 PAND2X1_837/CTRL POR2X1_42/Y 0.01fF
C35863 PAND2X1_792/B POR2X1_533/A 0.28fF
C35864 POR2X1_66/A POR2X1_404/CTRL2 0.01fF
C35865 PAND2X1_859/O POR2X1_93/Y 0.01fF
C35866 PAND2X1_502/O POR2X1_77/Y 0.03fF
C35867 POR2X1_20/B INPUT_4 0.07fF
C35868 POR2X1_814/A POR2X1_391/Y 0.07fF
C35869 POR2X1_779/A POR2X1_648/Y 0.01fF
C35870 D_INPUT_5 PAND2X1_21/a_16_344# 0.02fF
C35871 PAND2X1_93/B POR2X1_718/A 0.03fF
C35872 POR2X1_68/A PAND2X1_617/O 0.06fF
C35873 POR2X1_20/B POR2X1_763/Y 0.07fF
C35874 POR2X1_677/Y PAND2X1_175/B 0.00fF
C35875 POR2X1_32/A POR2X1_40/Y 0.18fF
C35876 POR2X1_301/A POR2X1_325/A 0.08fF
C35877 POR2X1_39/CTRL2 POR2X1_669/B 0.01fF
C35878 POR2X1_66/B PAND2X1_58/A 0.80fF
C35879 POR2X1_624/B PAND2X1_6/A 1.65fF
C35880 POR2X1_66/B POR2X1_641/CTRL 0.01fF
C35881 POR2X1_861/O POR2X1_499/A 0.03fF
C35882 PAND2X1_71/O PAND2X1_39/B 0.05fF
C35883 POR2X1_67/Y POR2X1_38/Y 0.02fF
C35884 POR2X1_555/B PAND2X1_7/Y 0.01fF
C35885 POR2X1_60/A PAND2X1_169/Y 0.03fF
C35886 PAND2X1_41/B POR2X1_174/A 0.03fF
C35887 PAND2X1_658/A POR2X1_20/B 0.02fF
C35888 PAND2X1_217/CTRL PAND2X1_197/Y 0.00fF
C35889 POR2X1_188/A PAND2X1_58/A 0.03fF
C35890 PAND2X1_20/A PAND2X1_616/a_16_344# 0.01fF
C35891 PAND2X1_266/a_16_344# POR2X1_73/Y 0.02fF
C35892 POR2X1_51/B PAND2X1_635/Y 0.06fF
C35893 POR2X1_83/B POR2X1_312/Y -0.00fF
C35894 POR2X1_254/A POR2X1_254/CTRL2 0.01fF
C35895 PAND2X1_826/CTRL2 PAND2X1_55/Y 0.01fF
C35896 POR2X1_88/A PAND2X1_6/A 0.04fF
C35897 POR2X1_471/CTRL2 POR2X1_66/A 0.03fF
C35898 PAND2X1_594/a_76_28# POR2X1_186/Y 0.01fF
C35899 POR2X1_13/A POR2X1_118/Y 0.03fF
C35900 POR2X1_23/Y PAND2X1_795/B 0.03fF
C35901 POR2X1_650/CTRL2 PAND2X1_65/B 0.01fF
C35902 POR2X1_254/CTRL2 POR2X1_750/B 0.05fF
C35903 POR2X1_66/O PAND2X1_96/B 0.06fF
C35904 POR2X1_417/Y POR2X1_40/Y 0.03fF
C35905 PAND2X1_95/B POR2X1_635/A 0.01fF
C35906 POR2X1_419/Y POR2X1_40/Y 0.02fF
C35907 POR2X1_866/A POR2X1_784/A 0.08fF
C35908 PAND2X1_20/A POR2X1_456/O 0.01fF
C35909 POR2X1_609/Y VDD 0.16fF
C35910 POR2X1_94/CTRL POR2X1_24/Y 0.01fF
C35911 POR2X1_175/O PAND2X1_73/Y 0.01fF
C35912 PAND2X1_39/B PAND2X1_744/O 0.21fF
C35913 POR2X1_499/A POR2X1_500/Y 0.01fF
C35914 PAND2X1_436/A POR2X1_677/CTRL2 0.03fF
C35915 POR2X1_670/CTRL2 POR2X1_40/Y 0.02fF
C35916 POR2X1_96/A POR2X1_420/O 0.02fF
C35917 POR2X1_20/B POR2X1_73/Y 1.27fF
C35918 POR2X1_648/Y POR2X1_407/CTRL 0.01fF
C35919 PAND2X1_80/O POR2X1_296/B 0.00fF
C35920 PAND2X1_267/Y PAND2X1_197/Y 0.02fF
C35921 POR2X1_48/A POR2X1_372/Y 0.02fF
C35922 PAND2X1_659/B POR2X1_32/A 0.03fF
C35923 POR2X1_60/A PAND2X1_333/a_76_28# 0.02fF
C35924 POR2X1_102/Y POR2X1_272/Y 0.04fF
C35925 POR2X1_120/O POR2X1_805/Y 0.06fF
C35926 POR2X1_355/B POR2X1_97/A 0.03fF
C35927 PAND2X1_824/B PAND2X1_234/O 0.02fF
C35928 PAND2X1_16/CTRL PAND2X1_41/B 0.01fF
C35929 POR2X1_482/Y POR2X1_5/Y 0.03fF
C35930 POR2X1_49/Y PAND2X1_576/CTRL 0.01fF
C35931 POR2X1_411/B PAND2X1_555/Y 0.03fF
C35932 PAND2X1_658/CTRL POR2X1_376/B 0.05fF
C35933 POR2X1_860/A PAND2X1_41/B 0.03fF
C35934 PAND2X1_279/CTRL POR2X1_284/B 0.00fF
C35935 PAND2X1_697/CTRL2 POR2X1_260/B 0.01fF
C35936 D_INPUT_0 POR2X1_232/O 0.01fF
C35937 POR2X1_420/Y VDD 0.10fF
C35938 INPUT_1 POR2X1_67/Y 0.03fF
C35939 POR2X1_669/Y PAND2X1_720/O 0.02fF
C35940 POR2X1_174/B POR2X1_853/CTRL2 0.32fF
C35941 POR2X1_669/B POR2X1_252/CTRL 0.08fF
C35942 POR2X1_13/A PAND2X1_573/B 0.05fF
C35943 POR2X1_859/A PAND2X1_58/A 0.10fF
C35944 POR2X1_676/a_16_28# POR2X1_828/A 0.05fF
C35945 POR2X1_676/a_76_344# PAND2X1_69/A 0.01fF
C35946 PAND2X1_61/Y POR2X1_376/B 0.14fF
C35947 PAND2X1_571/A POR2X1_599/A 0.05fF
C35948 PAND2X1_409/CTRL PAND2X1_11/Y 0.01fF
C35949 POR2X1_48/A POR2X1_519/Y 0.14fF
C35950 POR2X1_538/O POR2X1_270/Y 0.01fF
C35951 POR2X1_445/A POR2X1_540/CTRL 0.13fF
C35952 POR2X1_416/Y POR2X1_48/A 0.01fF
C35953 POR2X1_857/CTRL2 POR2X1_785/A -0.00fF
C35954 PAND2X1_6/Y POR2X1_270/Y 0.08fF
C35955 POR2X1_389/CTRL2 POR2X1_121/B 0.01fF
C35956 POR2X1_636/a_16_28# POR2X1_636/A -0.00fF
C35957 POR2X1_48/A POR2X1_253/Y 0.01fF
C35958 PAND2X1_244/B POR2X1_20/B 0.03fF
C35959 PAND2X1_48/B PAND2X1_282/m4_208_n4# 0.07fF
C35960 PAND2X1_273/a_16_344# D_INPUT_0 0.01fF
C35961 POR2X1_78/B POR2X1_403/O 0.01fF
C35962 POR2X1_616/a_56_344# POR2X1_90/Y 0.00fF
C35963 POR2X1_295/a_16_28# POR2X1_481/A 0.08fF
C35964 POR2X1_678/A POR2X1_513/B 0.00fF
C35965 POR2X1_404/B POR2X1_404/CTRL 0.01fF
C35966 PAND2X1_35/Y POR2X1_40/Y 0.15fF
C35967 POR2X1_32/A POR2X1_587/Y 0.14fF
C35968 POR2X1_801/B PAND2X1_583/CTRL2 0.00fF
C35969 POR2X1_81/a_76_344# POR2X1_293/Y 0.01fF
C35970 POR2X1_439/Y VDD 0.30fF
C35971 PAND2X1_570/a_76_28# PAND2X1_771/Y 0.02fF
C35972 POR2X1_43/B POR2X1_669/B 0.08fF
C35973 POR2X1_335/A POR2X1_590/A 0.05fF
C35974 POR2X1_163/Y PAND2X1_725/A 0.06fF
C35975 POR2X1_846/Y POR2X1_753/O 0.01fF
C35976 POR2X1_856/CTRL2 POR2X1_855/Y 0.01fF
C35977 PAND2X1_148/Y POR2X1_669/B 0.03fF
C35978 PAND2X1_97/O POR2X1_91/Y 0.11fF
C35979 PAND2X1_774/O PAND2X1_773/Y 0.00fF
C35980 POR2X1_275/CTRL PAND2X1_390/Y 0.01fF
C35981 POR2X1_48/A POR2X1_526/Y 0.02fF
C35982 POR2X1_790/A POR2X1_720/O 0.06fF
C35983 PAND2X1_137/O PAND2X1_354/A 0.01fF
C35984 POR2X1_830/O POR2X1_733/A 0.03fF
C35985 POR2X1_529/CTRL POR2X1_40/Y 0.01fF
C35986 POR2X1_414/Y POR2X1_293/Y 0.53fF
C35987 POR2X1_137/Y POR2X1_476/A 0.05fF
C35988 POR2X1_437/Y POR2X1_60/A 0.01fF
C35989 POR2X1_78/A POR2X1_713/Y 0.01fF
C35990 POR2X1_137/B POR2X1_559/A 0.10fF
C35991 POR2X1_455/CTRL2 POR2X1_76/Y 0.03fF
C35992 PAND2X1_267/O POR2X1_7/A 0.03fF
C35993 PAND2X1_80/O POR2X1_547/B 0.02fF
C35994 POR2X1_189/Y POR2X1_40/Y 0.03fF
C35995 PAND2X1_236/O INPUT_0 0.16fF
C35996 POR2X1_29/A POR2X1_748/O 0.01fF
C35997 POR2X1_647/CTRL POR2X1_101/Y 0.01fF
C35998 PAND2X1_652/A PAND2X1_361/a_16_344# 0.05fF
C35999 POR2X1_72/B PAND2X1_717/CTRL 0.01fF
C36000 PAND2X1_659/CTRL2 PAND2X1_735/Y 0.05fF
C36001 POR2X1_669/B POR2X1_38/B 0.05fF
C36002 PAND2X1_841/m4_208_n4# POR2X1_516/Y 0.12fF
C36003 PAND2X1_93/B POR2X1_725/Y 0.07fF
C36004 PAND2X1_793/Y PAND2X1_76/Y 0.03fF
C36005 PAND2X1_511/CTRL VDD 0.00fF
C36006 PAND2X1_721/O POR2X1_7/B 0.08fF
C36007 PAND2X1_356/B POR2X1_42/Y 0.01fF
C36008 POR2X1_614/A PAND2X1_230/a_16_344# 0.02fF
C36009 POR2X1_41/B POR2X1_48/CTRL 0.09fF
C36010 POR2X1_646/CTRL POR2X1_480/A 0.01fF
C36011 PAND2X1_651/Y PAND2X1_512/CTRL2 0.00fF
C36012 POR2X1_184/Y POR2X1_40/Y 0.03fF
C36013 POR2X1_192/Y VDD 9.49fF
C36014 D_INPUT_3 POR2X1_414/CTRL2 0.03fF
C36015 POR2X1_864/A PAND2X1_48/A 0.00fF
C36016 POR2X1_844/O POR2X1_590/A 0.01fF
C36017 POR2X1_37/Y PAND2X1_549/B 0.03fF
C36018 D_GATE_222 POR2X1_186/Y 0.08fF
C36019 PAND2X1_466/CTRL PAND2X1_803/A 0.00fF
C36020 POR2X1_20/Y POR2X1_94/A 0.19fF
C36021 POR2X1_37/Y POR2X1_416/CTRL 0.01fF
C36022 PAND2X1_809/B PAND2X1_809/O 0.08fF
C36023 PAND2X1_95/B PAND2X1_18/CTRL 0.01fF
C36024 POR2X1_66/B PAND2X1_96/B 9.82fF
C36025 POR2X1_84/A POR2X1_260/A 0.03fF
C36026 POR2X1_814/A POR2X1_383/Y 3.27fF
C36027 POR2X1_114/B PAND2X1_299/O 0.02fF
C36028 PAND2X1_651/Y POR2X1_40/Y 0.05fF
C36029 PAND2X1_3/A PAND2X1_1/a_16_344# 0.03fF
C36030 POR2X1_334/B PAND2X1_262/a_56_28# 0.00fF
C36031 POR2X1_64/m4_208_n4# POR2X1_44/m4_208_n4# 0.18fF
C36032 POR2X1_122/Y POR2X1_42/Y 0.03fF
C36033 POR2X1_422/Y POR2X1_583/a_76_344# 0.01fF
C36034 POR2X1_481/A POR2X1_7/B 0.03fF
C36035 PAND2X1_216/a_16_344# INPUT_0 0.01fF
C36036 POR2X1_188/A PAND2X1_96/B 0.03fF
C36037 POR2X1_65/A PAND2X1_642/B 0.11fF
C36038 PAND2X1_88/O POR2X1_38/B 0.04fF
C36039 POR2X1_502/A POR2X1_651/CTRL 0.06fF
C36040 PAND2X1_724/CTRL PAND2X1_731/B 0.01fF
C36041 POR2X1_356/A POR2X1_244/B 0.05fF
C36042 POR2X1_681/CTRL POR2X1_39/B 0.02fF
C36043 PAND2X1_42/CTRL2 POR2X1_68/B 0.01fF
C36044 POR2X1_700/O VDD 0.00fF
C36045 POR2X1_78/A POR2X1_725/Y 0.07fF
C36046 PAND2X1_250/a_76_28# POR2X1_778/B 0.04fF
C36047 POR2X1_29/Y POR2X1_159/a_16_28# 0.01fF
C36048 POR2X1_406/A POR2X1_5/Y 0.01fF
C36049 POR2X1_657/a_16_28# POR2X1_510/Y -0.00fF
C36050 POR2X1_113/CTRL2 POR2X1_640/Y 0.01fF
C36051 POR2X1_13/A POR2X1_669/a_16_28# 0.03fF
C36052 POR2X1_78/B POR2X1_341/O 0.02fF
C36053 POR2X1_8/Y D_INPUT_0 0.02fF
C36054 POR2X1_590/A POR2X1_249/Y 0.03fF
C36055 PAND2X1_573/B PAND2X1_510/B 0.02fF
C36056 PAND2X1_57/B POR2X1_832/B 0.01fF
C36057 POR2X1_355/B POR2X1_366/Y 0.07fF
C36058 POR2X1_355/B POR2X1_294/B 0.06fF
C36059 POR2X1_41/B PAND2X1_724/B 0.01fF
C36060 POR2X1_96/A PAND2X1_736/A 0.07fF
C36061 PAND2X1_58/CTRL2 PAND2X1_69/A 0.06fF
C36062 POR2X1_254/Y PAND2X1_56/Y 0.10fF
C36063 POR2X1_254/Y POR2X1_795/B 0.17fF
C36064 POR2X1_305/a_16_28# POR2X1_42/Y 0.03fF
C36065 PAND2X1_96/B POR2X1_563/CTRL 0.03fF
C36066 POR2X1_832/a_16_28# PAND2X1_55/Y 0.01fF
C36067 POR2X1_14/Y POR2X1_419/CTRL 0.01fF
C36068 POR2X1_260/B POR2X1_571/Y 0.02fF
C36069 POR2X1_360/A PAND2X1_55/Y 0.02fF
C36070 POR2X1_327/Y POR2X1_66/A 0.03fF
C36071 PAND2X1_850/Y POR2X1_257/A 0.07fF
C36072 POR2X1_569/a_16_28# PAND2X1_32/B 0.02fF
C36073 POR2X1_347/A POR2X1_296/B 0.00fF
C36074 PAND2X1_453/A POR2X1_419/CTRL 0.01fF
C36075 POR2X1_573/O POR2X1_573/A 0.03fF
C36076 POR2X1_855/B POR2X1_808/A 0.00fF
C36077 POR2X1_298/Y POR2X1_394/A 0.96fF
C36078 POR2X1_16/A POR2X1_60/A 0.23fF
C36079 POR2X1_78/B POR2X1_194/CTRL 0.01fF
C36080 PAND2X1_456/CTRL POR2X1_283/A 0.00fF
C36081 PAND2X1_738/Y PAND2X1_182/CTRL 0.01fF
C36082 PAND2X1_651/Y PAND2X1_659/B 0.05fF
C36083 POR2X1_686/B PAND2X1_69/A 0.01fF
C36084 POR2X1_353/Y POR2X1_353/CTRL 0.01fF
C36085 PAND2X1_137/Y PAND2X1_357/Y 0.03fF
C36086 POR2X1_87/Y POR2X1_68/B 0.04fF
C36087 POR2X1_572/CTRL PAND2X1_32/B 0.01fF
C36088 POR2X1_283/A POR2X1_226/Y 0.02fF
C36089 POR2X1_78/A POR2X1_559/A 0.23fF
C36090 POR2X1_43/B PAND2X1_844/Y 0.02fF
C36091 PAND2X1_6/A PAND2X1_375/CTRL2 0.00fF
C36092 POR2X1_360/A POR2X1_402/A 0.04fF
C36093 POR2X1_16/A POR2X1_591/A 0.01fF
C36094 POR2X1_192/Y PAND2X1_32/B 2.56fF
C36095 PAND2X1_553/B POR2X1_183/Y 0.00fF
C36096 POR2X1_390/B POR2X1_777/B 0.03fF
C36097 POR2X1_3/A VDD 1.12fF
C36098 PAND2X1_86/Y POR2X1_99/A 0.01fF
C36099 POR2X1_13/A PAND2X1_341/A 0.06fF
C36100 PAND2X1_474/Y POR2X1_91/Y 0.03fF
C36101 PAND2X1_236/m4_208_n4# POR2X1_68/B 0.07fF
C36102 PAND2X1_693/a_16_344# PAND2X1_48/B 0.01fF
C36103 POR2X1_65/A PAND2X1_550/B 0.08fF
C36104 POR2X1_785/O PAND2X1_32/B 0.09fF
C36105 POR2X1_305/Y PAND2X1_506/CTRL2 0.01fF
C36106 POR2X1_83/Y POR2X1_263/Y 0.02fF
C36107 PAND2X1_63/B POR2X1_5/Y 0.54fF
C36108 POR2X1_740/Y POR2X1_574/CTRL 0.01fF
C36109 POR2X1_741/Y POR2X1_574/CTRL2 0.01fF
C36110 POR2X1_41/B PAND2X1_186/CTRL2 0.03fF
C36111 PAND2X1_672/a_76_28# POR2X1_260/A 0.02fF
C36112 POR2X1_150/Y POR2X1_173/CTRL2 0.01fF
C36113 POR2X1_413/A POR2X1_416/Y 0.03fF
C36114 POR2X1_13/A POR2X1_93/A 0.13fF
C36115 POR2X1_65/A POR2X1_83/O 0.01fF
C36116 POR2X1_343/Y POR2X1_624/Y 0.10fF
C36117 POR2X1_13/A POR2X1_91/Y 0.10fF
C36118 POR2X1_178/Y POR2X1_106/Y 0.12fF
C36119 POR2X1_7/B PAND2X1_645/B 0.01fF
C36120 POR2X1_54/O PAND2X1_58/A 0.01fF
C36121 POR2X1_55/Y PAND2X1_548/CTRL 0.01fF
C36122 PAND2X1_96/B PAND2X1_89/a_16_344# 0.02fF
C36123 PAND2X1_56/Y POR2X1_574/O 0.11fF
C36124 PAND2X1_621/a_76_28# POR2X1_750/B 0.01fF
C36125 POR2X1_327/Y PAND2X1_279/a_16_344# 0.01fF
C36126 POR2X1_532/A POR2X1_578/Y 0.03fF
C36127 PAND2X1_572/O POR2X1_46/Y 0.01fF
C36128 POR2X1_807/A POR2X1_675/Y 0.01fF
C36129 POR2X1_76/Y PAND2X1_60/B 0.03fF
C36130 PAND2X1_799/a_56_28# INPUT_0 0.00fF
C36131 PAND2X1_90/A POR2X1_243/O 0.01fF
C36132 POR2X1_174/B PAND2X1_165/CTRL 0.14fF
C36133 PAND2X1_687/CTRL POR2X1_60/A 0.01fF
C36134 POR2X1_265/Y POR2X1_667/A 0.01fF
C36135 PAND2X1_837/O POR2X1_825/Y 0.01fF
C36136 PAND2X1_341/A PAND2X1_197/O 0.02fF
C36137 POR2X1_296/B POR2X1_4/Y 0.15fF
C36138 POR2X1_254/Y POR2X1_383/A 0.15fF
C36139 PAND2X1_223/B PAND2X1_643/A 0.01fF
C36140 VDD POR2X1_568/Y 5.86fF
C36141 PAND2X1_725/Y PAND2X1_162/A 0.01fF
C36142 PAND2X1_830/O VDD 0.00fF
C36143 PAND2X1_775/O POR2X1_91/Y 0.02fF
C36144 PAND2X1_137/Y PAND2X1_140/A 0.34fF
C36145 PAND2X1_421/O POR2X1_596/A 0.02fF
C36146 POR2X1_13/A PAND2X1_720/CTRL 0.01fF
C36147 POR2X1_68/B POR2X1_8/a_16_28# 0.00fF
C36148 POR2X1_502/A POR2X1_854/B 0.14fF
C36149 PAND2X1_810/CTRL2 GATE_741 0.01fF
C36150 POR2X1_60/A PAND2X1_336/Y 0.05fF
C36151 POR2X1_785/B VDD 0.03fF
C36152 POR2X1_700/a_16_28# POR2X1_90/Y 0.05fF
C36153 PAND2X1_388/Y POR2X1_293/Y 0.00fF
C36154 PAND2X1_643/Y POR2X1_761/a_56_344# 0.00fF
C36155 PAND2X1_563/A PAND2X1_563/B 0.13fF
C36156 POR2X1_334/CTRL VDD 0.00fF
C36157 PAND2X1_79/Y PAND2X1_316/CTRL2 0.03fF
C36158 POR2X1_619/A POR2X1_619/CTRL 0.03fF
C36159 POR2X1_293/Y PAND2X1_549/B 0.07fF
C36160 PAND2X1_713/CTRL PAND2X1_725/B 0.02fF
C36161 PAND2X1_184/CTRL VDD -0.00fF
C36162 POR2X1_57/A PAND2X1_675/A 0.06fF
C36163 POR2X1_35/B POR2X1_294/A 0.02fF
C36164 POR2X1_740/Y PAND2X1_60/B 0.04fF
C36165 POR2X1_57/A PAND2X1_469/B 0.03fF
C36166 POR2X1_326/A POR2X1_653/B 0.03fF
C36167 PAND2X1_641/Y VDD 0.05fF
C36168 POR2X1_416/CTRL POR2X1_293/Y 0.01fF
C36169 POR2X1_566/A POR2X1_456/B 0.12fF
C36170 POR2X1_523/Y PAND2X1_521/CTRL 0.01fF
C36171 POR2X1_447/B POR2X1_202/O 0.01fF
C36172 POR2X1_383/A POR2X1_575/B 0.15fF
C36173 PAND2X1_17/a_76_28# INPUT_6 0.01fF
C36174 PAND2X1_572/CTRL2 POR2X1_52/Y 0.00fF
C36175 POR2X1_333/O POR2X1_578/Y 0.02fF
C36176 PAND2X1_23/Y PAND2X1_505/a_76_28# 0.04fF
C36177 PAND2X1_84/O POR2X1_394/A 0.07fF
C36178 POR2X1_345/A POR2X1_99/B 0.02fF
C36179 PAND2X1_495/CTRL PAND2X1_69/A 0.00fF
C36180 D_INPUT_3 PAND2X1_6/A 0.10fF
C36181 POR2X1_403/O POR2X1_294/A 0.17fF
C36182 POR2X1_259/CTRL POR2X1_785/A 0.00fF
C36183 POR2X1_549/O POR2X1_620/B 0.06fF
C36184 PAND2X1_737/B POR2X1_7/B 0.20fF
C36185 PAND2X1_215/B POR2X1_7/CTRL 0.08fF
C36186 POR2X1_362/B PAND2X1_48/A 0.00fF
C36187 POR2X1_455/A POR2X1_222/A 0.06fF
C36188 POR2X1_307/CTRL2 POR2X1_711/Y 0.05fF
C36189 POR2X1_353/Y POR2X1_191/Y 0.05fF
C36190 PAND2X1_95/B PAND2X1_51/CTRL2 0.03fF
C36191 PAND2X1_30/CTRL POR2X1_635/A 0.01fF
C36192 POR2X1_283/A POR2X1_56/Y 0.02fF
C36193 PAND2X1_659/Y POR2X1_822/CTRL2 0.01fF
C36194 PAND2X1_715/B PAND2X1_115/B 0.07fF
C36195 POR2X1_606/Y PAND2X1_56/A 0.01fF
C36196 POR2X1_316/CTRL2 POR2X1_293/Y 0.03fF
C36197 POR2X1_345/a_16_28# POR2X1_244/B 0.02fF
C36198 PAND2X1_466/A POR2X1_329/A 0.02fF
C36199 PAND2X1_94/A PAND2X1_411/CTRL2 0.01fF
C36200 POR2X1_754/A POR2X1_754/a_16_28# 0.04fF
C36201 POR2X1_25/Y VDD 0.00fF
C36202 PAND2X1_587/Y PAND2X1_3/B 4.32fF
C36203 PAND2X1_831/CTRL2 POR2X1_39/B 0.03fF
C36204 PAND2X1_6/Y POR2X1_101/Y 0.03fF
C36205 POR2X1_74/Y POR2X1_272/Y 0.05fF
C36206 POR2X1_262/Y POR2X1_329/A 0.03fF
C36207 POR2X1_327/Y POR2X1_802/B 0.10fF
C36208 POR2X1_13/A POR2X1_109/Y 0.03fF
C36209 PAND2X1_642/B PAND2X1_559/a_16_344# 0.02fF
C36210 POR2X1_784/CTRL POR2X1_725/Y 0.05fF
C36211 POR2X1_383/A POR2X1_341/Y 0.06fF
C36212 POR2X1_547/B POR2X1_4/Y 0.03fF
C36213 POR2X1_615/Y POR2X1_129/Y 0.00fF
C36214 POR2X1_740/Y POR2X1_787/a_16_28# 0.06fF
C36215 POR2X1_76/B POR2X1_274/CTRL 0.01fF
C36216 PAND2X1_90/A PAND2X1_531/CTRL 0.03fF
C36217 POR2X1_785/B PAND2X1_32/B 0.02fF
C36218 POR2X1_325/A POR2X1_374/O 0.01fF
C36219 POR2X1_732/O POR2X1_353/A 0.01fF
C36220 POR2X1_96/A POR2X1_7/Y 0.02fF
C36221 POR2X1_814/B PAND2X1_179/a_76_28# 0.01fF
C36222 PAND2X1_775/O POR2X1_109/Y 0.01fF
C36223 POR2X1_294/B POR2X1_195/CTRL2 0.01fF
C36224 PAND2X1_803/Y POR2X1_283/A 0.03fF
C36225 POR2X1_145/Y POR2X1_146/CTRL 0.00fF
C36226 POR2X1_383/A POR2X1_338/CTRL2 0.01fF
C36227 POR2X1_477/B PAND2X1_52/B 0.03fF
C36228 POR2X1_502/A POR2X1_374/CTRL2 0.01fF
C36229 POR2X1_51/B POR2X1_36/B 0.83fF
C36230 PAND2X1_90/A PAND2X1_90/CTRL2 0.01fF
C36231 POR2X1_532/A POR2X1_774/B 0.01fF
C36232 POR2X1_456/B POR2X1_573/A 0.04fF
C36233 PAND2X1_357/Y PAND2X1_853/B 0.03fF
C36234 POR2X1_486/B VDD 0.19fF
C36235 POR2X1_710/Y POR2X1_713/B 0.01fF
C36236 POR2X1_83/Y PAND2X1_215/B 0.02fF
C36237 POR2X1_99/B POR2X1_205/Y 0.03fF
C36238 POR2X1_169/Y POR2X1_566/B 0.04fF
C36239 POR2X1_99/B PAND2X1_55/Y 0.03fF
C36240 POR2X1_49/Y POR2X1_49/O 0.01fF
C36241 POR2X1_855/B POR2X1_687/A 0.02fF
C36242 POR2X1_643/O POR2X1_590/A 0.01fF
C36243 POR2X1_327/Y POR2X1_532/A 0.03fF
C36244 PAND2X1_55/Y PAND2X1_304/CTRL 0.00fF
C36245 PAND2X1_846/O INPUT_0 0.04fF
C36246 POR2X1_178/Y PAND2X1_114/B 0.00fF
C36247 POR2X1_687/CTRL2 POR2X1_814/A 0.02fF
C36248 POR2X1_83/Y PAND2X1_6/A 0.03fF
C36249 PAND2X1_156/B PAND2X1_156/O 0.00fF
C36250 POR2X1_41/Y POR2X1_43/B 0.00fF
C36251 POR2X1_458/Y POR2X1_296/B 0.01fF
C36252 PAND2X1_53/CTRL POR2X1_66/A 0.01fF
C36253 POR2X1_704/Y POR2X1_704/O 0.00fF
C36254 PAND2X1_830/a_76_28# POR2X1_108/Y 0.07fF
C36255 PAND2X1_284/Y PAND2X1_345/Y 0.09fF
C36256 POR2X1_774/A PAND2X1_60/B 0.06fF
C36257 POR2X1_614/A POR2X1_156/O 0.18fF
C36258 VDD POR2X1_356/Y 0.89fF
C36259 POR2X1_81/A POR2X1_43/B 0.09fF
C36260 PAND2X1_6/Y POR2X1_542/CTRL2 0.01fF
C36261 POR2X1_244/B PAND2X1_72/A 0.03fF
C36262 POR2X1_54/Y POR2X1_24/Y 0.00fF
C36263 POR2X1_371/CTRL2 POR2X1_387/Y 0.06fF
C36264 PAND2X1_6/Y POR2X1_359/a_16_28# 0.00fF
C36265 POR2X1_673/Y POR2X1_546/CTRL2 0.03fF
C36266 POR2X1_103/a_56_344# PAND2X1_349/A 0.00fF
C36267 PAND2X1_724/B POR2X1_77/Y 0.02fF
C36268 POR2X1_485/Y POR2X1_48/A 0.03fF
C36269 POR2X1_8/Y POR2X1_10/O 0.06fF
C36270 POR2X1_136/Y POR2X1_183/a_76_344# 0.01fF
C36271 POR2X1_76/B VDD 0.02fF
C36272 POR2X1_152/O POR2X1_39/B 0.01fF
C36273 PAND2X1_289/CTRL2 POR2X1_220/B 0.02fF
C36274 POR2X1_7/A POR2X1_7/Y 0.03fF
C36275 POR2X1_296/O POR2X1_296/B 0.01fF
C36276 POR2X1_499/A POR2X1_499/a_16_28# 0.03fF
C36277 POR2X1_447/B POR2X1_566/B 0.05fF
C36278 POR2X1_753/Y POR2X1_20/B 0.07fF
C36279 PAND2X1_117/a_76_28# PAND2X1_72/A 0.01fF
C36280 POR2X1_86/O PAND2X1_338/B 0.01fF
C36281 POR2X1_250/Y PAND2X1_742/a_56_28# 0.00fF
C36282 POR2X1_326/A POR2X1_449/A 0.03fF
C36283 PAND2X1_20/A POR2X1_499/A 0.03fF
C36284 POR2X1_546/O POR2X1_550/B 0.00fF
C36285 POR2X1_394/A POR2X1_314/Y 0.10fF
C36286 POR2X1_464/O POR2X1_457/Y 0.00fF
C36287 POR2X1_86/Y POR2X1_73/Y 0.11fF
C36288 POR2X1_832/Y D_INPUT_0 0.03fF
C36289 POR2X1_456/B PAND2X1_167/CTRL 0.00fF
C36290 PAND2X1_108/CTRL PAND2X1_60/B 0.01fF
C36291 PAND2X1_73/Y POR2X1_688/Y 0.09fF
C36292 POR2X1_23/Y POR2X1_482/CTRL2 0.03fF
C36293 POR2X1_20/B PAND2X1_541/CTRL2 0.02fF
C36294 POR2X1_41/B PAND2X1_458/CTRL 0.03fF
C36295 POR2X1_1/O D_INPUT_4 0.08fF
C36296 POR2X1_43/Y POR2X1_73/Y 0.03fF
C36297 POR2X1_69/Y VDD 0.06fF
C36298 POR2X1_203/CTRL2 PAND2X1_72/A 0.00fF
C36299 PAND2X1_91/a_76_28# POR2X1_97/A 0.03fF
C36300 POR2X1_537/a_16_28# POR2X1_537/Y 0.02fF
C36301 POR2X1_678/A POR2X1_678/a_16_28# 0.15fF
C36302 POR2X1_499/A POR2X1_814/B 0.03fF
C36303 PAND2X1_20/A POR2X1_76/A 0.03fF
C36304 POR2X1_849/B POR2X1_29/A 0.01fF
C36305 PAND2X1_865/Y POR2X1_394/A 0.05fF
C36306 POR2X1_646/B VDD 0.11fF
C36307 POR2X1_41/B POR2X1_441/CTRL2 0.10fF
C36308 PAND2X1_251/O POR2X1_296/B 0.02fF
C36309 POR2X1_84/A POR2X1_243/A 0.01fF
C36310 POR2X1_252/Y PAND2X1_508/Y 0.01fF
C36311 POR2X1_610/a_76_344# POR2X1_590/A 0.01fF
C36312 PAND2X1_717/A PAND2X1_804/B 0.05fF
C36313 POR2X1_76/B PAND2X1_32/B 0.01fF
C36314 POR2X1_811/CTRL PAND2X1_73/Y 0.01fF
C36315 PAND2X1_726/B POR2X1_39/B 0.24fF
C36316 POR2X1_68/CTRL2 POR2X1_296/B 0.00fF
C36317 POR2X1_648/Y PAND2X1_511/a_76_28# 0.01fF
C36318 PAND2X1_35/A PAND2X1_35/B 0.14fF
C36319 POR2X1_503/CTRL POR2X1_77/Y 0.01fF
C36320 POR2X1_590/Y PAND2X1_304/a_76_28# 0.03fF
C36321 POR2X1_20/B PAND2X1_563/B 0.00fF
C36322 PAND2X1_93/B POR2X1_811/B 0.08fF
C36323 POR2X1_329/Y PAND2X1_730/B 0.03fF
C36324 PAND2X1_796/B PAND2X1_783/Y 0.00fF
C36325 POR2X1_101/Y PAND2X1_52/B 0.03fF
C36326 POR2X1_597/Y POR2X1_236/Y 0.07fF
C36327 POR2X1_447/B POR2X1_508/B 0.00fF
C36328 POR2X1_552/O POR2X1_542/Y 0.04fF
C36329 PAND2X1_810/B GATE_741 0.00fF
C36330 PAND2X1_86/O POR2X1_404/Y 0.01fF
C36331 POR2X1_814/B POR2X1_76/A 0.03fF
C36332 POR2X1_202/A POR2X1_202/a_16_28# 0.02fF
C36333 POR2X1_614/O POR2X1_750/B 0.01fF
C36334 POR2X1_63/Y VDD 0.40fF
C36335 POR2X1_866/CTRL2 POR2X1_801/B 0.01fF
C36336 POR2X1_303/a_16_28# POR2X1_274/A 0.03fF
C36337 PAND2X1_93/B PAND2X1_387/CTRL2 0.02fF
C36338 POR2X1_56/a_16_28# POR2X1_496/Y 0.04fF
C36339 POR2X1_343/Y POR2X1_186/B 0.05fF
C36340 PAND2X1_23/Y PAND2X1_75/a_16_344# 0.01fF
C36341 PAND2X1_464/a_16_344# PAND2X1_445/Y 0.02fF
C36342 PAND2X1_48/A D_INPUT_4 0.99fF
C36343 POR2X1_411/B POR2X1_46/Y 0.05fF
C36344 POR2X1_78/A POR2X1_811/B 0.01fF
C36345 PAND2X1_469/O POR2X1_236/Y 0.02fF
C36346 PAND2X1_427/CTRL2 POR2X1_121/B 0.05fF
C36347 POR2X1_89/O POR2X1_5/Y 0.19fF
C36348 PAND2X1_97/CTRL POR2X1_5/Y 0.01fF
C36349 PAND2X1_258/CTRL PAND2X1_52/Y 0.01fF
C36350 POR2X1_465/O POR2X1_563/Y 0.01fF
C36351 POR2X1_556/A POR2X1_404/Y 0.12fF
C36352 POR2X1_88/CTRL2 VDD 0.00fF
C36353 POR2X1_49/Y PAND2X1_61/CTRL 0.01fF
C36354 POR2X1_96/A POR2X1_257/A 0.17fF
C36355 PAND2X1_62/CTRL2 D_INPUT_0 0.01fF
C36356 POR2X1_32/A PAND2X1_706/O 0.01fF
C36357 PAND2X1_630/B POR2X1_245/Y 0.03fF
C36358 PAND2X1_88/O POR2X1_590/A 0.17fF
C36359 PAND2X1_561/a_16_344# PAND2X1_558/Y 0.02fF
C36360 POR2X1_467/Y POR2X1_448/O 0.01fF
C36361 PAND2X1_79/CTRL2 POR2X1_78/Y 0.03fF
C36362 POR2X1_301/A VDD 0.15fF
C36363 POR2X1_824/O POR2X1_77/Y 0.00fF
C36364 PAND2X1_287/Y VDD 0.20fF
C36365 POR2X1_227/A POR2X1_35/Y 0.03fF
C36366 INPUT_1 PAND2X1_42/a_76_28# 0.01fF
C36367 POR2X1_83/B POR2X1_698/O 0.16fF
C36368 POR2X1_416/Y PAND2X1_634/O 0.02fF
C36369 POR2X1_427/CTRL POR2X1_236/Y 0.01fF
C36370 POR2X1_69/A POR2X1_750/A 0.02fF
C36371 POR2X1_644/CTRL POR2X1_513/B 0.02fF
C36372 POR2X1_83/B POR2X1_250/A 0.07fF
C36373 POR2X1_32/A POR2X1_5/Y 0.28fF
C36374 POR2X1_356/A POR2X1_319/A 0.05fF
C36375 POR2X1_66/B POR2X1_355/A 0.00fF
C36376 POR2X1_549/O POR2X1_78/A 0.01fF
C36377 POR2X1_138/O POR2X1_624/Y 0.11fF
C36378 POR2X1_13/A POR2X1_422/a_16_28# 0.01fF
C36379 POR2X1_40/Y PAND2X1_731/B 0.05fF
C36380 POR2X1_630/A PAND2X1_41/B 0.03fF
C36381 PAND2X1_235/CTRL2 PAND2X1_85/Y 0.01fF
C36382 PAND2X1_673/CTRL POR2X1_83/B 0.01fF
C36383 POR2X1_27/O PAND2X1_63/B 0.01fF
C36384 POR2X1_496/Y PAND2X1_778/a_16_344# 0.02fF
C36385 POR2X1_614/A POR2X1_663/B 0.03fF
C36386 POR2X1_673/A POR2X1_296/B 0.01fF
C36387 POR2X1_35/B POR2X1_94/A 0.03fF
C36388 PAND2X1_829/a_16_344# PAND2X1_65/B 0.02fF
C36389 INPUT_3 POR2X1_409/CTRL 0.13fF
C36390 D_INPUT_5 POR2X1_638/B 0.01fF
C36391 PAND2X1_630/B PAND2X1_507/CTRL 0.01fF
C36392 POR2X1_126/O D_INPUT_2 0.01fF
C36393 POR2X1_140/B POR2X1_659/A 0.11fF
C36394 PAND2X1_319/B POR2X1_150/Y 0.00fF
C36395 PAND2X1_296/O PAND2X1_347/Y 0.04fF
C36396 POR2X1_416/B PAND2X1_346/a_56_28# 0.00fF
C36397 POR2X1_307/Y D_INPUT_0 0.03fF
C36398 POR2X1_49/Y PAND2X1_211/A 0.02fF
C36399 PAND2X1_77/CTRL PAND2X1_8/Y 0.01fF
C36400 POR2X1_775/A POR2X1_260/B 0.84fF
C36401 POR2X1_390/B POR2X1_814/A 0.06fF
C36402 POR2X1_416/B PAND2X1_198/O 0.09fF
C36403 POR2X1_788/A VDD 0.27fF
C36404 POR2X1_23/Y POR2X1_697/Y 0.05fF
C36405 POR2X1_417/Y POR2X1_5/Y 0.04fF
C36406 POR2X1_43/B PAND2X1_436/O 0.17fF
C36407 POR2X1_114/B PAND2X1_406/O 0.03fF
C36408 POR2X1_476/A POR2X1_294/B 0.07fF
C36409 POR2X1_502/A PAND2X1_73/Y 0.20fF
C36410 POR2X1_673/Y POR2X1_69/Y 0.05fF
C36411 POR2X1_41/B POR2X1_496/Y 0.04fF
C36412 PAND2X1_73/Y POR2X1_783/A 0.01fF
C36413 POR2X1_66/B PAND2X1_377/CTRL2 0.13fF
C36414 PAND2X1_467/B PAND2X1_707/CTRL 0.01fF
C36415 PAND2X1_751/CTRL POR2X1_590/A 0.02fF
C36416 PAND2X1_225/CTRL VDD 0.00fF
C36417 PAND2X1_71/CTRL POR2X1_296/B 0.02fF
C36418 PAND2X1_360/O PAND2X1_347/Y 0.09fF
C36419 POR2X1_832/CTRL POR2X1_330/Y 0.01fF
C36420 POR2X1_678/A VDD -0.00fF
C36421 POR2X1_288/A POR2X1_362/B 0.03fF
C36422 POR2X1_20/B PAND2X1_656/A 0.03fF
C36423 PAND2X1_106/O POR2X1_116/A 0.00fF
C36424 POR2X1_66/B POR2X1_415/CTRL 0.02fF
C36425 PAND2X1_56/Y POR2X1_842/O 0.03fF
C36426 POR2X1_447/CTRL POR2X1_447/A 0.01fF
C36427 POR2X1_821/CTRL2 POR2X1_40/Y 0.00fF
C36428 POR2X1_174/B POR2X1_776/B 0.07fF
C36429 POR2X1_335/A POR2X1_66/A 0.88fF
C36430 PAND2X1_651/Y POR2X1_613/O 0.00fF
C36431 POR2X1_302/B POR2X1_284/B 0.61fF
C36432 POR2X1_634/A PAND2X1_57/B 0.11fF
C36433 POR2X1_220/CTRL POR2X1_220/A 0.01fF
C36434 POR2X1_220/O POR2X1_210/Y 0.01fF
C36435 POR2X1_290/Y POR2X1_83/B 0.03fF
C36436 POR2X1_674/a_16_28# PAND2X1_652/A 0.07fF
C36437 POR2X1_446/B POR2X1_714/CTRL 0.09fF
C36438 POR2X1_722/A POR2X1_814/A 0.31fF
C36439 POR2X1_13/A POR2X1_595/a_16_28# 0.07fF
C36440 POR2X1_366/CTRL POR2X1_556/A 0.01fF
C36441 PAND2X1_390/Y INPUT_0 0.08fF
C36442 POR2X1_813/Y POR2X1_63/Y 0.01fF
C36443 POR2X1_257/A POR2X1_7/A 0.24fF
C36444 PAND2X1_557/A POR2X1_79/Y 0.03fF
C36445 POR2X1_567/B POR2X1_535/m4_208_n4# 0.17fF
C36446 PAND2X1_714/A POR2X1_236/Y 0.01fF
C36447 POR2X1_51/A POR2X1_40/Y 0.01fF
C36448 POR2X1_446/B POR2X1_228/Y 0.03fF
C36449 POR2X1_271/Y POR2X1_46/Y 0.05fF
C36450 PAND2X1_65/CTRL2 PAND2X1_69/A 0.03fF
C36451 POR2X1_539/A PAND2X1_39/B 0.03fF
C36452 POR2X1_678/Y PAND2X1_69/A 0.01fF
C36453 POR2X1_480/A POR2X1_830/A 0.02fF
C36454 PAND2X1_220/Y POR2X1_481/A 0.03fF
C36455 POR2X1_644/Y POR2X1_532/A 0.04fF
C36456 POR2X1_278/Y PAND2X1_659/A 0.05fF
C36457 POR2X1_41/B PAND2X1_733/A 0.07fF
C36458 PAND2X1_209/A PAND2X1_782/Y 0.00fF
C36459 POR2X1_311/Y PAND2X1_736/A 0.01fF
C36460 POR2X1_523/Y POR2X1_29/A 0.03fF
C36461 POR2X1_683/Y POR2X1_669/B 0.01fF
C36462 POR2X1_49/Y POR2X1_96/A 0.31fF
C36463 POR2X1_13/A POR2X1_278/CTRL2 0.01fF
C36464 POR2X1_14/Y POR2X1_415/Y 0.11fF
C36465 PAND2X1_768/Y VDD 0.35fF
C36466 POR2X1_65/A PAND2X1_734/B 0.03fF
C36467 POR2X1_83/B PAND2X1_658/B 0.05fF
C36468 POR2X1_555/A POR2X1_194/B 0.10fF
C36469 POR2X1_526/CTRL2 POR2X1_32/A 0.03fF
C36470 POR2X1_856/B POR2X1_209/A 0.02fF
C36471 PAND2X1_479/O PAND2X1_480/B 0.00fF
C36472 PAND2X1_230/CTRL POR2X1_795/B 0.06fF
C36473 POR2X1_23/Y POR2X1_278/A 0.04fF
C36474 POR2X1_825/CTRL POR2X1_42/Y 0.01fF
C36475 D_INPUT_0 POR2X1_68/B 1.77fF
C36476 POR2X1_720/B PAND2X1_58/A 0.07fF
C36477 POR2X1_366/Y POR2X1_269/Y 0.04fF
C36478 PAND2X1_641/Y PAND2X1_9/Y 0.03fF
C36479 PAND2X1_90/A PAND2X1_42/CTRL2 0.02fF
C36480 POR2X1_29/A PAND2X1_69/A 24.66fF
C36481 PAND2X1_645/CTRL VDD -0.00fF
C36482 D_INPUT_1 POR2X1_296/B 0.02fF
C36483 POR2X1_376/B POR2X1_46/Y 0.10fF
C36484 INPUT_7 INPUT_4 0.93fF
C36485 POR2X1_672/CTRL POR2X1_102/Y 0.04fF
C36486 POR2X1_294/CTRL POR2X1_260/A 0.01fF
C36487 PAND2X1_474/CTRL2 POR2X1_153/Y 0.08fF
C36488 POR2X1_16/A PAND2X1_443/CTRL2 0.01fF
C36489 PAND2X1_469/B PAND2X1_556/a_16_344# 0.04fF
C36490 POR2X1_750/B POR2X1_740/Y 0.03fF
C36491 PAND2X1_139/B VDD 0.04fF
C36492 POR2X1_150/Y PAND2X1_357/CTRL2 0.06fF
C36493 POR2X1_66/B PAND2X1_767/CTRL2 0.01fF
C36494 PAND2X1_456/CTRL POR2X1_55/Y 0.01fF
C36495 POR2X1_834/a_76_344# POR2X1_407/Y 0.00fF
C36496 POR2X1_826/Y POR2X1_153/Y 0.20fF
C36497 POR2X1_615/O POR2X1_615/Y 0.01fF
C36498 POR2X1_760/A POR2X1_7/Y 0.03fF
C36499 POR2X1_57/CTRL POR2X1_5/Y 0.01fF
C36500 POR2X1_93/A POR2X1_29/A 0.16fF
C36501 POR2X1_296/B POR2X1_724/A 0.03fF
C36502 POR2X1_130/A PAND2X1_57/B 0.03fF
C36503 PAND2X1_41/B POR2X1_795/B 0.03fF
C36504 POR2X1_859/A POR2X1_415/CTRL 0.14fF
C36505 POR2X1_529/CTRL POR2X1_5/Y 0.17fF
C36506 PAND2X1_421/O PAND2X1_90/Y 0.01fF
C36507 POR2X1_312/Y PAND2X1_357/Y 1.49fF
C36508 POR2X1_804/A POR2X1_330/Y 0.29fF
C36509 POR2X1_834/Y PAND2X1_601/m4_208_n4# 0.04fF
C36510 POR2X1_754/Y POR2X1_283/A 0.07fF
C36511 POR2X1_566/A PAND2X1_57/B 0.03fF
C36512 PAND2X1_245/O PAND2X1_111/B 0.02fF
C36513 POR2X1_54/Y PAND2X1_522/a_76_28# 0.05fF
C36514 POR2X1_416/B POR2X1_846/A 0.00fF
C36515 POR2X1_72/B PAND2X1_565/A 0.70fF
C36516 POR2X1_163/a_16_28# POR2X1_163/A 0.03fF
C36517 PAND2X1_118/CTRL PAND2X1_65/B 0.01fF
C36518 PAND2X1_71/O VDD 0.00fF
C36519 POR2X1_68/A POR2X1_849/CTRL 0.01fF
C36520 POR2X1_66/A POR2X1_249/Y 0.06fF
C36521 PAND2X1_793/Y PAND2X1_480/B 0.05fF
C36522 POR2X1_68/A PAND2X1_55/O 0.09fF
C36523 POR2X1_441/Y POR2X1_373/a_56_344# 0.00fF
C36524 POR2X1_201/O PAND2X1_88/Y 0.01fF
C36525 PAND2X1_598/O POR2X1_46/Y 0.10fF
C36526 PAND2X1_278/CTRL2 POR2X1_68/B 0.03fF
C36527 POR2X1_60/A PAND2X1_388/Y 0.05fF
C36528 PAND2X1_217/B PAND2X1_575/CTRL2 0.32fF
C36529 POR2X1_48/A PAND2X1_726/B 0.13fF
C36530 POR2X1_146/CTRL POR2X1_669/B 0.03fF
C36531 POR2X1_832/A PAND2X1_58/A 0.03fF
C36532 POR2X1_84/CTRL VDD 0.00fF
C36533 POR2X1_251/CTRL2 POR2X1_387/Y 0.04fF
C36534 PAND2X1_631/A POR2X1_20/B 0.07fF
C36535 PAND2X1_411/O PAND2X1_90/Y 0.02fF
C36536 PAND2X1_13/CTRL PAND2X1_32/B 0.01fF
C36537 POR2X1_43/B PAND2X1_499/Y 0.08fF
C36538 PAND2X1_401/O POR2X1_236/Y 0.01fF
C36539 POR2X1_52/A POR2X1_46/Y 0.11fF
C36540 PAND2X1_478/B PAND2X1_469/Y 0.01fF
C36541 POR2X1_60/A PAND2X1_549/B 0.05fF
C36542 POR2X1_750/B PAND2X1_312/CTRL2 0.01fF
C36543 POR2X1_556/A POR2X1_554/CTRL 0.05fF
C36544 PAND2X1_169/Y POR2X1_142/Y 0.03fF
C36545 INPUT_6 POR2X1_750/B 0.03fF
C36546 PAND2X1_3/CTRL PAND2X1_11/Y 0.01fF
C36547 PAND2X1_651/Y POR2X1_5/Y 0.04fF
C36548 PAND2X1_425/a_16_344# D_INPUT_6 0.03fF
C36549 POR2X1_814/B POR2X1_540/A 0.21fF
C36550 POR2X1_608/CTRL POR2X1_712/Y 0.03fF
C36551 PAND2X1_69/A POR2X1_213/B 0.83fF
C36552 POR2X1_40/CTRL POR2X1_83/B 0.01fF
C36553 PAND2X1_592/Y PAND2X1_191/Y 0.01fF
C36554 POR2X1_10/CTRL POR2X1_669/B 0.01fF
C36555 POR2X1_96/A PAND2X1_188/O 0.04fF
C36556 PAND2X1_841/CTRL2 PAND2X1_841/B 0.02fF
C36557 POR2X1_24/Y POR2X1_4/Y 0.09fF
C36558 POR2X1_236/Y POR2X1_816/A 0.03fF
C36559 PAND2X1_280/O POR2X1_662/Y 0.02fF
C36560 POR2X1_241/B POR2X1_456/B 0.09fF
C36561 POR2X1_358/O POR2X1_578/Y 0.02fF
C36562 POR2X1_356/A PAND2X1_48/B 0.35fF
C36563 POR2X1_654/CTRL2 POR2X1_725/Y 0.01fF
C36564 PAND2X1_95/B POR2X1_638/CTRL2 0.01fF
C36565 POR2X1_51/A POR2X1_587/Y 0.03fF
C36566 PAND2X1_691/Y POR2X1_829/CTRL2 0.01fF
C36567 POR2X1_523/Y POR2X1_546/A 0.16fF
C36568 PAND2X1_90/Y POR2X1_68/B 0.11fF
C36569 POR2X1_669/B POR2X1_39/Y 0.01fF
C36570 POR2X1_276/A POR2X1_141/Y 0.29fF
C36571 POR2X1_210/O POR2X1_210/B 0.01fF
C36572 PAND2X1_844/B POR2X1_5/Y 0.06fF
C36573 D_INPUT_1 POR2X1_547/B 0.02fF
C36574 POR2X1_306/CTRL2 POR2X1_236/Y 0.01fF
C36575 POR2X1_49/Y POR2X1_7/A 0.16fF
C36576 POR2X1_72/B PAND2X1_123/CTRL2 0.03fF
C36577 POR2X1_777/B PAND2X1_63/B 0.12fF
C36578 POR2X1_383/A PAND2X1_41/B 0.81fF
C36579 VDD POR2X1_498/A 0.00fF
C36580 PAND2X1_623/CTRL POR2X1_129/Y 0.01fF
C36581 POR2X1_102/Y PAND2X1_532/O 0.01fF
C36582 POR2X1_130/a_16_28# POR2X1_244/Y 0.02fF
C36583 POR2X1_658/a_16_28# POR2X1_632/Y 0.03fF
C36584 PAND2X1_472/O POR2X1_60/A 0.04fF
C36585 POR2X1_259/A POR2X1_259/CTRL2 0.01fF
C36586 PAND2X1_6/O PAND2X1_20/A 0.02fF
C36587 PAND2X1_23/Y POR2X1_276/O 0.08fF
C36588 POR2X1_634/A POR2X1_771/A 0.05fF
C36589 PAND2X1_474/A POR2X1_171/CTRL2 0.00fF
C36590 PAND2X1_69/A POR2X1_546/A 0.03fF
C36591 POR2X1_814/B POR2X1_537/A 0.00fF
C36592 PAND2X1_645/O PAND2X1_645/B 0.01fF
C36593 POR2X1_539/A POR2X1_814/B 0.01fF
C36594 POR2X1_65/A PAND2X1_661/Y 0.03fF
C36595 POR2X1_16/A POR2X1_750/A 0.02fF
C36596 POR2X1_775/CTRL POR2X1_776/B 0.00fF
C36597 PAND2X1_284/Y VDD 0.41fF
C36598 POR2X1_13/A POR2X1_299/CTRL 0.01fF
C36599 POR2X1_775/A PAND2X1_55/Y 0.03fF
C36600 PAND2X1_710/CTRL POR2X1_763/A 0.08fF
C36601 POR2X1_628/CTRL PAND2X1_6/A 0.03fF
C36602 PAND2X1_65/B PAND2X1_63/B 0.03fF
C36603 POR2X1_840/B POR2X1_217/a_16_28# 0.07fF
C36604 POR2X1_539/A POR2X1_733/CTRL 0.02fF
C36605 PAND2X1_57/B POR2X1_573/A 0.03fF
C36606 POR2X1_170/B POR2X1_577/CTRL 0.11fF
C36607 PAND2X1_754/O PAND2X1_69/A 0.03fF
C36608 POR2X1_43/B PAND2X1_466/O 0.05fF
C36609 POR2X1_207/B POR2X1_207/a_16_28# 0.01fF
C36610 PAND2X1_478/B POR2X1_394/A 0.03fF
C36611 PAND2X1_854/A POR2X1_236/Y 0.05fF
C36612 POR2X1_55/Y POR2X1_56/Y 0.01fF
C36613 POR2X1_288/A POR2X1_734/CTRL 0.00fF
C36614 PAND2X1_467/Y PAND2X1_803/A 0.03fF
C36615 PAND2X1_6/Y PAND2X1_23/Y 0.16fF
C36616 POR2X1_296/B POR2X1_620/B 0.55fF
C36617 POR2X1_539/A POR2X1_325/A 0.03fF
C36618 POR2X1_366/Y POR2X1_513/Y 0.03fF
C36619 GATE_479 POR2X1_16/A 0.03fF
C36620 POR2X1_763/Y POR2X1_73/Y 0.03fF
C36621 POR2X1_66/B POR2X1_735/CTRL2 0.01fF
C36622 POR2X1_832/A POR2X1_435/Y 0.01fF
C36623 POR2X1_174/B POR2X1_192/B 0.17fF
C36624 PAND2X1_489/CTRL2 PAND2X1_580/B 0.00fF
C36625 PAND2X1_687/A POR2X1_13/A 0.00fF
C36626 POR2X1_68/A PAND2X1_49/O 0.01fF
C36627 POR2X1_256/Y PAND2X1_514/Y 0.05fF
C36628 POR2X1_790/A POR2X1_391/Y 0.01fF
C36629 POR2X1_400/A POR2X1_215/A 0.05fF
C36630 POR2X1_376/B POR2X1_376/O 0.01fF
C36631 PAND2X1_69/A PAND2X1_369/m4_208_n4# 0.12fF
C36632 POR2X1_805/A PAND2X1_69/A 0.03fF
C36633 PAND2X1_658/A POR2X1_73/Y 0.03fF
C36634 POR2X1_246/O POR2X1_90/Y 0.10fF
C36635 POR2X1_333/A POR2X1_357/B 0.03fF
C36636 POR2X1_205/A POR2X1_294/B 0.07fF
C36637 POR2X1_504/a_16_28# POR2X1_750/B 0.00fF
C36638 POR2X1_712/A PAND2X1_697/O 0.02fF
C36639 PAND2X1_557/A PAND2X1_730/A 0.03fF
C36640 POR2X1_43/B PAND2X1_734/O 0.02fF
C36641 POR2X1_38/B PAND2X1_29/CTRL2 0.01fF
C36642 D_INPUT_1 POR2X1_267/Y 0.03fF
C36643 PAND2X1_803/Y POR2X1_55/Y 0.02fF
C36644 PAND2X1_553/B POR2X1_7/A 0.01fF
C36645 POR2X1_319/A PAND2X1_72/A 0.03fF
C36646 PAND2X1_41/B PAND2X1_71/Y 0.03fF
C36647 PAND2X1_591/CTRL PAND2X1_56/A 0.01fF
C36648 POR2X1_760/Y POR2X1_102/Y 0.01fF
C36649 POR2X1_262/O POR2X1_7/A 0.01fF
C36650 POR2X1_449/A POR2X1_480/A 0.02fF
C36651 PAND2X1_631/O POR2X1_90/Y 0.01fF
C36652 POR2X1_96/A PAND2X1_641/CTRL 0.01fF
C36653 PAND2X1_438/CTRL2 POR2X1_456/B 0.03fF
C36654 POR2X1_654/B POR2X1_294/A 0.02fF
C36655 POR2X1_294/B POR2X1_366/A 0.03fF
C36656 PAND2X1_57/B POR2X1_596/CTRL 0.01fF
C36657 POR2X1_228/a_16_28# PAND2X1_7/Y 0.05fF
C36658 POR2X1_283/A POR2X1_42/Y 0.26fF
C36659 PAND2X1_56/Y POR2X1_228/Y 0.05fF
C36660 PAND2X1_48/B POR2X1_569/A 0.07fF
C36661 POR2X1_326/A PAND2X1_90/Y 0.05fF
C36662 POR2X1_304/O POR2X1_102/Y 0.01fF
C36663 PAND2X1_69/A PAND2X1_150/CTRL 0.01fF
C36664 POR2X1_119/Y PAND2X1_541/O 0.01fF
C36665 POR2X1_7/B PAND2X1_348/O 0.02fF
C36666 POR2X1_496/Y POR2X1_77/Y 0.07fF
C36667 POR2X1_48/m4_208_n4# PAND2X1_196/m4_208_n4# 0.05fF
C36668 POR2X1_836/A POR2X1_568/B 0.01fF
C36669 POR2X1_13/A POR2X1_599/CTRL2 0.00fF
C36670 PAND2X1_308/B PAND2X1_308/O 0.00fF
C36671 POR2X1_116/Y POR2X1_392/a_76_344# 0.01fF
C36672 POR2X1_68/A POR2X1_550/Y 0.05fF
C36673 POR2X1_153/CTRL PAND2X1_472/B 0.08fF
C36674 POR2X1_55/Y PAND2X1_508/CTRL2 0.03fF
C36675 PAND2X1_658/A PAND2X1_244/B 0.03fF
C36676 POR2X1_840/B PAND2X1_72/a_76_28# 0.01fF
C36677 POR2X1_344/Y PAND2X1_57/B 0.03fF
C36678 POR2X1_187/a_16_28# POR2X1_79/Y 0.02fF
C36679 PAND2X1_472/a_76_28# PAND2X1_673/Y 0.01fF
C36680 PAND2X1_333/a_16_344# POR2X1_171/Y 0.03fF
C36681 POR2X1_103/O POR2X1_13/A 0.18fF
C36682 PAND2X1_460/O POR2X1_68/B 0.01fF
C36683 POR2X1_638/Y PAND2X1_60/B 0.02fF
C36684 POR2X1_90/Y PAND2X1_348/Y 0.03fF
C36685 POR2X1_318/A POR2X1_140/CTRL 0.00fF
C36686 POR2X1_669/B PAND2X1_326/O 0.06fF
C36687 PAND2X1_691/Y PAND2X1_649/O 0.01fF
C36688 PAND2X1_81/CTRL PAND2X1_63/B 0.01fF
C36689 POR2X1_547/B POR2X1_620/B 0.06fF
C36690 POR2X1_16/A PAND2X1_649/CTRL2 0.01fF
C36691 POR2X1_81/A PAND2X1_474/A 0.10fF
C36692 POR2X1_336/O POR2X1_228/Y 0.02fF
C36693 POR2X1_57/A PAND2X1_389/Y 0.03fF
C36694 POR2X1_291/a_16_28# POR2X1_42/Y 0.02fF
C36695 POR2X1_349/CTRL2 PAND2X1_57/B 0.03fF
C36696 POR2X1_369/Y PAND2X1_543/O 0.00fF
C36697 POR2X1_301/CTRL2 POR2X1_260/A 0.00fF
C36698 PAND2X1_384/m4_208_n4# POR2X1_546/A 0.15fF
C36699 POR2X1_346/B POR2X1_66/CTRL2 0.00fF
C36700 PAND2X1_733/A POR2X1_77/Y 0.02fF
C36701 POR2X1_851/CTRL POR2X1_733/A 0.08fF
C36702 PAND2X1_778/Y POR2X1_7/A 0.03fF
C36703 PAND2X1_236/a_16_344# POR2X1_4/Y 0.08fF
C36704 POR2X1_845/O POR2X1_532/A 0.05fF
C36705 POR2X1_438/O PAND2X1_569/B 0.01fF
C36706 POR2X1_785/A POR2X1_186/B 0.03fF
C36707 PAND2X1_291/a_16_344# PAND2X1_88/Y 0.01fF
C36708 POR2X1_78/B PAND2X1_41/Y 0.01fF
C36709 PAND2X1_244/B POR2X1_73/Y 0.06fF
C36710 POR2X1_532/A PAND2X1_133/CTRL2 0.01fF
C36711 POR2X1_345/a_16_28# PAND2X1_48/B 0.02fF
C36712 PAND2X1_63/Y POR2X1_773/B 0.07fF
C36713 PAND2X1_111/B POR2X1_366/A 0.03fF
C36714 POR2X1_68/A POR2X1_782/B 0.04fF
C36715 POR2X1_110/Y POR2X1_368/a_16_28# 0.03fF
C36716 POR2X1_170/B POR2X1_191/Y 0.05fF
C36717 POR2X1_383/A POR2X1_228/Y 1.06fF
C36718 PAND2X1_96/B POR2X1_259/a_76_344# 0.01fF
C36719 POR2X1_840/Y VDD 0.18fF
C36720 PAND2X1_499/O POR2X1_39/B 0.01fF
C36721 POR2X1_790/A POR2X1_753/O 0.02fF
C36722 POR2X1_407/A PAND2X1_310/CTRL2 0.00fF
C36723 PAND2X1_180/CTRL2 POR2X1_77/Y 0.00fF
C36724 PAND2X1_865/CTRL2 PAND2X1_175/B 0.01fF
C36725 PAND2X1_226/O POR2X1_191/Y 0.17fF
C36726 POR2X1_736/CTRL POR2X1_675/Y 0.01fF
C36727 PAND2X1_661/B POR2X1_599/CTRL2 0.01fF
C36728 PAND2X1_543/CTRL2 POR2X1_77/Y 0.11fF
C36729 PAND2X1_301/CTRL2 POR2X1_91/Y 0.03fF
C36730 POR2X1_804/A POR2X1_715/A 0.03fF
C36731 POR2X1_113/Y POR2X1_773/B 0.05fF
C36732 POR2X1_16/A POR2X1_142/Y 0.03fF
C36733 POR2X1_62/Y PAND2X1_339/Y 0.03fF
C36734 PAND2X1_8/Y PAND2X1_102/O 0.05fF
C36735 POR2X1_346/B PAND2X1_60/CTRL2 0.00fF
C36736 POR2X1_285/B POR2X1_285/O 0.01fF
C36737 PAND2X1_6/Y POR2X1_809/A 0.02fF
C36738 POR2X1_383/A POR2X1_561/CTRL 0.00fF
C36739 POR2X1_566/B POR2X1_577/Y 0.03fF
C36740 POR2X1_775/CTRL POR2X1_192/B 0.15fF
C36741 POR2X1_825/O POR2X1_825/Y 0.01fF
C36742 POR2X1_800/A POR2X1_691/A 0.00fF
C36743 POR2X1_66/Y PAND2X1_43/CTRL2 0.01fF
C36744 POR2X1_446/B POR2X1_657/Y 0.92fF
C36745 POR2X1_126/CTRL POR2X1_411/B 0.01fF
C36746 PAND2X1_575/a_56_28# POR2X1_394/A 0.00fF
C36747 PAND2X1_353/CTRL2 PAND2X1_303/Y 0.01fF
C36748 POR2X1_751/Y POR2X1_748/Y 0.00fF
C36749 PAND2X1_819/O POR2X1_260/A 0.02fF
C36750 POR2X1_445/A POR2X1_471/A 0.03fF
C36751 POR2X1_220/Y POR2X1_325/B 0.00fF
C36752 POR2X1_27/O POR2X1_32/A 0.01fF
C36753 POR2X1_773/B POR2X1_260/A 0.03fF
C36754 PAND2X1_23/Y POR2X1_632/Y 0.03fF
C36755 POR2X1_853/A POR2X1_568/B 0.01fF
C36756 POR2X1_57/A POR2X1_397/CTRL2 0.03fF
C36757 POR2X1_101/Y POR2X1_216/Y 0.08fF
C36758 PAND2X1_771/a_76_28# PAND2X1_769/Y 0.02fF
C36759 PAND2X1_454/O POR2X1_77/Y 0.01fF
C36760 PAND2X1_223/O PAND2X1_221/Y 0.02fF
C36761 POR2X1_192/Y POR2X1_568/A 0.22fF
C36762 PAND2X1_336/Y POR2X1_142/Y 0.03fF
C36763 POR2X1_43/B POR2X1_39/B 1.06fF
C36764 POR2X1_411/B PAND2X1_571/A 0.03fF
C36765 PAND2X1_779/CTRL POR2X1_527/Y 0.01fF
C36766 POR2X1_364/A POR2X1_168/a_16_28# 0.01fF
C36767 PAND2X1_715/B PAND2X1_348/A 0.02fF
C36768 PAND2X1_152/O PAND2X1_72/A 0.02fF
C36769 POR2X1_416/B POR2X1_45/Y 0.07fF
C36770 POR2X1_166/CTRL PAND2X1_326/B 0.01fF
C36771 PAND2X1_360/Y PAND2X1_343/CTRL2 0.00fF
C36772 PAND2X1_23/Y PAND2X1_52/B 2.06fF
C36773 PAND2X1_48/B PAND2X1_72/A 0.18fF
C36774 PAND2X1_69/A POR2X1_343/O 0.10fF
C36775 PAND2X1_6/Y POR2X1_711/Y 0.07fF
C36776 PAND2X1_761/O D_INPUT_0 0.04fF
C36777 POR2X1_38/B POR2X1_39/B 0.07fF
C36778 POR2X1_48/A PAND2X1_35/A 0.06fF
C36779 PAND2X1_404/Y PAND2X1_640/B 0.07fF
C36780 POR2X1_648/A PAND2X1_90/Y 0.05fF
C36781 POR2X1_138/a_16_28# POR2X1_138/A 0.02fF
C36782 POR2X1_737/A POR2X1_733/Y 0.08fF
C36783 POR2X1_49/Y POR2X1_760/A 0.07fF
C36784 POR2X1_48/A POR2X1_817/CTRL 0.00fF
C36785 POR2X1_661/A PAND2X1_385/CTRL2 0.02fF
C36786 PAND2X1_631/A PAND2X1_715/B 0.03fF
C36787 PAND2X1_467/B POR2X1_257/A 0.05fF
C36788 PAND2X1_88/Y POR2X1_555/a_56_344# 0.00fF
C36789 PAND2X1_127/O POR2X1_567/A -0.02fF
C36790 POR2X1_147/CTRL POR2X1_532/A 0.01fF
C36791 PAND2X1_295/O POR2X1_296/B 0.15fF
C36792 POR2X1_657/O POR2X1_446/B 0.01fF
C36793 PAND2X1_635/Y POR2X1_7/B 0.03fF
C36794 PAND2X1_628/O POR2X1_785/A 0.07fF
C36795 PAND2X1_269/O VDD 0.00fF
C36796 PAND2X1_621/Y POR2X1_9/Y 0.02fF
C36797 POR2X1_604/CTRL2 POR2X1_72/B 0.03fF
C36798 POR2X1_347/A POR2X1_347/O 0.01fF
C36799 POR2X1_406/Y PAND2X1_266/CTRL 0.00fF
C36800 PAND2X1_434/CTRL POR2X1_39/B 0.00fF
C36801 POR2X1_590/A POR2X1_458/CTRL 0.00fF
C36802 POR2X1_472/CTRL2 PAND2X1_52/B 0.01fF
C36803 POR2X1_311/O POR2X1_77/Y 0.02fF
C36804 PAND2X1_449/CTRL POR2X1_511/Y 0.00fF
C36805 PAND2X1_93/B POR2X1_296/B 0.07fF
C36806 POR2X1_88/m4_208_n4# POR2X1_669/B 0.06fF
C36807 POR2X1_493/A PAND2X1_73/Y 0.07fF
C36808 POR2X1_13/A PAND2X1_717/A 0.17fF
C36809 POR2X1_49/Y PAND2X1_466/B 0.08fF
C36810 PAND2X1_39/B POR2X1_403/CTRL2 0.01fF
C36811 POR2X1_34/B POR2X1_34/A 0.60fF
C36812 PAND2X1_20/A POR2X1_849/B 0.01fF
C36813 POR2X1_66/B POR2X1_260/B 21.92fF
C36814 PAND2X1_309/CTRL POR2X1_814/A 0.01fF
C36815 PAND2X1_569/B PAND2X1_326/CTRL2 0.01fF
C36816 POR2X1_18/O INPUT_4 0.02fF
C36817 POR2X1_411/B PAND2X1_787/Y 0.01fF
C36818 PAND2X1_124/Y PAND2X1_195/CTRL2 0.01fF
C36819 POR2X1_23/Y POR2X1_667/A 0.73fF
C36820 POR2X1_536/O POR2X1_416/B 0.07fF
C36821 POR2X1_602/O POR2X1_330/Y 0.02fF
C36822 POR2X1_180/B POR2X1_181/Y 0.03fF
C36823 POR2X1_294/A PAND2X1_41/Y 0.01fF
C36824 POR2X1_499/A VDD 0.45fF
C36825 POR2X1_262/Y PAND2X1_84/Y 0.00fF
C36826 PAND2X1_73/Y PAND2X1_413/CTRL 0.00fF
C36827 POR2X1_188/A POR2X1_260/B 0.08fF
C36828 PAND2X1_865/Y POR2X1_767/O 0.01fF
C36829 D_INPUT_5 PAND2X1_18/CTRL2 0.00fF
C36830 POR2X1_484/Y PAND2X1_556/B 0.01fF
C36831 POR2X1_568/A POR2X1_568/Y 0.01fF
C36832 POR2X1_43/B POR2X1_827/O 0.02fF
C36833 POR2X1_862/B POR2X1_862/A 0.32fF
C36834 POR2X1_29/A POR2X1_720/O 0.10fF
C36835 POR2X1_78/A POR2X1_296/B 0.16fF
C36836 PAND2X1_624/a_76_28# POR2X1_20/B 0.02fF
C36837 POR2X1_479/B POR2X1_288/a_16_28# 0.01fF
C36838 POR2X1_609/Y PAND2X1_403/B 0.07fF
C36839 POR2X1_864/A POR2X1_855/Y 0.03fF
C36840 POR2X1_428/Y POR2X1_236/Y 0.01fF
C36841 PAND2X1_200/CTRL POR2X1_32/A 0.01fF
C36842 PAND2X1_88/O POR2X1_66/A 0.02fF
C36843 POR2X1_415/A VDD 0.15fF
C36844 PAND2X1_87/O PAND2X1_6/A 0.15fF
C36845 PAND2X1_508/Y PAND2X1_840/Y 0.03fF
C36846 POR2X1_106/CTRL2 POR2X1_251/A 0.11fF
C36847 POR2X1_78/A POR2X1_605/O 0.01fF
C36848 POR2X1_383/a_56_344# POR2X1_383/Y 0.00fF
C36849 POR2X1_117/CTRL POR2X1_48/A 0.01fF
C36850 PAND2X1_222/A VDD 0.00fF
C36851 POR2X1_491/CTRL POR2X1_32/A 0.01fF
C36852 PAND2X1_73/Y PAND2X1_74/O 0.09fF
C36853 POR2X1_76/A VDD 0.51fF
C36854 PAND2X1_108/a_56_28# PAND2X1_39/B 0.00fF
C36855 POR2X1_510/A POR2X1_835/B 0.00fF
C36856 PAND2X1_73/a_16_344# POR2X1_590/A 0.01fF
C36857 POR2X1_567/B PAND2X1_65/B 0.10fF
C36858 POR2X1_394/Y POR2X1_393/Y 0.01fF
C36859 POR2X1_809/A PAND2X1_52/B 0.02fF
C36860 POR2X1_504/Y POR2X1_626/a_16_28# 0.02fF
C36861 POR2X1_735/a_16_28# POR2X1_632/Y -0.00fF
C36862 POR2X1_852/B PAND2X1_39/CTRL2 0.06fF
C36863 POR2X1_88/a_56_344# INPUT_0 0.01fF
C36864 POR2X1_102/Y POR2X1_272/O 0.01fF
C36865 POR2X1_102/Y PAND2X1_390/Y 0.06fF
C36866 PAND2X1_20/A POR2X1_33/B 0.01fF
C36867 PAND2X1_798/B POR2X1_150/Y 0.54fF
C36868 POR2X1_260/B POR2X1_859/A 0.10fF
C36869 POR2X1_411/B PAND2X1_562/CTRL2 0.01fF
C36870 POR2X1_360/A POR2X1_240/O 0.08fF
C36871 PAND2X1_99/B VDD 0.00fF
C36872 D_INPUT_0 POR2X1_480/A 0.07fF
C36873 PAND2X1_406/O POR2X1_405/Y 0.00fF
C36874 POR2X1_486/m4_208_n4# POR2X1_532/A 0.06fF
C36875 POR2X1_432/CTRL2 POR2X1_236/Y 0.01fF
C36876 POR2X1_760/A PAND2X1_217/CTRL2 0.03fF
C36877 POR2X1_373/a_16_28# POR2X1_77/Y 0.03fF
C36878 PAND2X1_621/CTRL POR2X1_9/Y 0.04fF
C36879 PAND2X1_406/O POR2X1_784/A 0.01fF
C36880 PAND2X1_58/A PAND2X1_55/O 0.17fF
C36881 POR2X1_32/A PAND2X1_723/Y 0.07fF
C36882 PAND2X1_436/A PAND2X1_390/Y 0.01fF
C36883 POR2X1_499/A PAND2X1_32/B 0.03fF
C36884 POR2X1_634/O PAND2X1_41/B 0.01fF
C36885 POR2X1_614/A POR2X1_841/O 0.02fF
C36886 POR2X1_814/A PAND2X1_63/B 0.05fF
C36887 POR2X1_48/A POR2X1_411/CTRL 0.01fF
C36888 POR2X1_490/Y PAND2X1_228/CTRL2 0.03fF
C36889 POR2X1_79/CTRL PAND2X1_798/B 0.00fF
C36890 POR2X1_432/CTRL VDD 0.00fF
C36891 POR2X1_43/B PAND2X1_469/CTRL2 0.03fF
C36892 POR2X1_23/Y POR2X1_252/O 0.03fF
C36893 POR2X1_48/A POR2X1_252/CTRL 0.01fF
C36894 POR2X1_52/A PAND2X1_571/A 0.02fF
C36895 POR2X1_143/CTRL D_INPUT_0 0.01fF
C36896 POR2X1_504/Y POR2X1_505/Y 0.00fF
C36897 POR2X1_590/A POR2X1_207/CTRL 0.01fF
C36898 POR2X1_23/Y PAND2X1_254/CTRL2 0.01fF
C36899 POR2X1_39/O POR2X1_40/Y 0.01fF
C36900 POR2X1_78/A POR2X1_547/B 0.07fF
C36901 POR2X1_43/O POR2X1_77/Y 0.01fF
C36902 POR2X1_49/Y PAND2X1_478/Y 0.02fF
C36903 POR2X1_454/A POR2X1_795/B 0.07fF
C36904 PAND2X1_39/B PAND2X1_69/A 0.22fF
C36905 POR2X1_12/A PAND2X1_635/CTRL 0.01fF
C36906 POR2X1_834/CTRL2 POR2X1_513/B 0.03fF
C36907 PAND2X1_47/B VDD 0.42fF
C36908 POR2X1_186/Y PAND2X1_52/Y 0.03fF
C36909 POR2X1_679/Y POR2X1_816/A 0.01fF
C36910 POR2X1_614/A POR2X1_266/CTRL 0.06fF
C36911 POR2X1_94/A POR2X1_5/Y 1.11fF
C36912 POR2X1_725/CTRL POR2X1_711/Y 0.01fF
C36913 PAND2X1_90/A D_INPUT_0 0.13fF
C36914 POR2X1_72/B PAND2X1_736/O 0.03fF
C36915 POR2X1_613/Y POR2X1_386/Y 0.01fF
C36916 POR2X1_624/Y PAND2X1_79/Y 0.03fF
C36917 PAND2X1_498/CTRL2 POR2X1_590/A 0.03fF
C36918 POR2X1_423/CTRL2 POR2X1_372/Y 0.05fF
C36919 PAND2X1_65/B PAND2X1_386/CTRL 0.01fF
C36920 POR2X1_43/B POR2X1_48/A 0.45fF
C36921 POR2X1_83/B POR2X1_669/CTRL2 -0.00fF
C36922 PAND2X1_618/Y PAND2X1_69/A 0.01fF
C36923 POR2X1_333/A POR2X1_190/Y 0.05fF
C36924 POR2X1_119/Y PAND2X1_403/O 0.15fF
C36925 POR2X1_477/A POR2X1_436/B 0.01fF
C36926 PAND2X1_168/Y VDD 0.00fF
C36927 PAND2X1_354/A PAND2X1_580/B 0.03fF
C36928 POR2X1_311/Y PAND2X1_553/B 0.03fF
C36929 POR2X1_78/B POR2X1_194/A 0.00fF
C36930 POR2X1_817/Y POR2X1_817/m4_208_n4# 0.12fF
C36931 POR2X1_60/A PAND2X1_468/O 0.04fF
C36932 PAND2X1_793/O PAND2X1_793/A 0.02fF
C36933 POR2X1_13/Y PAND2X1_223/B 0.00fF
C36934 PAND2X1_23/Y POR2X1_478/Y 0.01fF
C36935 PAND2X1_52/B POR2X1_728/A 0.04fF
C36936 PAND2X1_644/Y POR2X1_759/A 0.00fF
C36937 POR2X1_308/CTRL2 POR2X1_830/A 0.09fF
C36938 POR2X1_814/B POR2X1_608/CTRL 0.01fF
C36939 PAND2X1_41/B INPUT_0 0.14fF
C36940 PAND2X1_640/B POR2X1_118/O 0.03fF
C36941 POR2X1_620/CTRL2 POR2X1_296/B 0.01fF
C36942 POR2X1_445/CTRL2 POR2X1_750/B 0.12fF
C36943 POR2X1_241/B POR2X1_341/CTRL2 0.01fF
C36944 POR2X1_480/A PAND2X1_90/Y 0.17fF
C36945 POR2X1_283/Y POR2X1_7/B 0.03fF
C36946 POR2X1_558/O POR2X1_78/A 0.03fF
C36947 POR2X1_96/A POR2X1_331/Y 0.03fF
C36948 POR2X1_14/Y POR2X1_42/Y 0.30fF
C36949 POR2X1_78/B PAND2X1_65/B 0.21fF
C36950 POR2X1_686/B POR2X1_828/Y 0.64fF
C36951 POR2X1_610/a_76_344# POR2X1_532/A 0.02fF
C36952 POR2X1_48/A POR2X1_38/B 0.06fF
C36953 POR2X1_223/O POR2X1_186/Y 0.01fF
C36954 PAND2X1_803/A PAND2X1_556/B 0.03fF
C36955 PAND2X1_56/Y POR2X1_657/O 0.31fF
C36956 POR2X1_431/a_16_28# POR2X1_129/Y 0.06fF
C36957 PAND2X1_453/A POR2X1_42/Y 0.02fF
C36958 PAND2X1_723/Y PAND2X1_741/B 0.02fF
C36959 POR2X1_66/B PAND2X1_55/Y 0.40fF
C36960 PAND2X1_572/CTRL PAND2X1_576/B 0.01fF
C36961 PAND2X1_84/CTRL POR2X1_497/Y 0.00fF
C36962 PAND2X1_318/O POR2X1_417/Y 0.03fF
C36963 POR2X1_814/A POR2X1_383/CTRL 0.02fF
C36964 POR2X1_383/A POR2X1_454/A 0.07fF
C36965 PAND2X1_798/B PAND2X1_794/O -0.02fF
C36966 D_INPUT_2 POR2X1_37/O 0.02fF
C36967 PAND2X1_834/CTRL POR2X1_677/Y 0.04fF
C36968 POR2X1_41/B PAND2X1_562/B 0.07fF
C36969 POR2X1_523/Y PAND2X1_20/A 0.04fF
C36970 INPUT_1 POR2X1_257/A 0.14fF
C36971 POR2X1_193/A PAND2X1_7/Y 0.08fF
C36972 PAND2X1_93/B PAND2X1_312/a_56_28# 0.00fF
C36973 POR2X1_188/A PAND2X1_55/Y 0.15fF
C36974 POR2X1_97/A POR2X1_577/O 0.01fF
C36975 PAND2X1_192/CTRL2 PAND2X1_191/Y 0.03fF
C36976 PAND2X1_592/CTRL PAND2X1_473/B 0.01fF
C36977 PAND2X1_612/B POR2X1_773/O 0.00fF
C36978 PAND2X1_824/B PAND2X1_39/B 0.07fF
C36979 POR2X1_8/Y POR2X1_54/Y 15.71fF
C36980 POR2X1_406/CTRL2 POR2X1_5/Y 0.01fF
C36981 POR2X1_707/B PAND2X1_587/O 0.04fF
C36982 PAND2X1_47/B PAND2X1_32/B 0.02fF
C36983 POR2X1_377/O POR2X1_94/A 0.04fF
C36984 PAND2X1_793/Y PAND2X1_473/B 0.03fF
C36985 PAND2X1_76/Y POR2X1_372/Y 0.03fF
C36986 PAND2X1_20/A PAND2X1_69/A 0.17fF
C36987 D_GATE_662 POR2X1_186/Y 0.12fF
C36988 POR2X1_814/B PAND2X1_372/a_76_28# 0.02fF
C36989 POR2X1_596/A POR2X1_834/a_16_28# 0.02fF
C36990 POR2X1_257/A POR2X1_153/Y 0.20fF
C36991 POR2X1_478/CTRL2 POR2X1_444/Y 0.04fF
C36992 POR2X1_65/A POR2X1_591/CTRL 0.01fF
C36993 POR2X1_52/A PAND2X1_859/a_76_28# 0.01fF
C36994 POR2X1_15/CTRL2 POR2X1_14/Y 0.01fF
C36995 POR2X1_257/A POR2X1_384/A 0.03fF
C36996 POR2X1_459/B POR2X1_750/B 0.01fF
C36997 PAND2X1_90/A PAND2X1_90/Y 0.01fF
C36998 POR2X1_41/B PAND2X1_715/CTRL 0.04fF
C36999 POR2X1_12/CTRL2 POR2X1_587/Y 0.01fF
C37000 POR2X1_416/B POR2X1_292/CTRL 0.01fF
C37001 PAND2X1_48/B POR2X1_632/A 0.05fF
C37002 PAND2X1_57/CTRL2 POR2X1_404/Y 0.03fF
C37003 POR2X1_8/Y POR2X1_77/a_56_344# 0.00fF
C37004 POR2X1_66/B POR2X1_407/Y 0.00fF
C37005 PAND2X1_852/O POR2X1_65/A 0.01fF
C37006 POR2X1_102/Y POR2X1_757/CTRL2 0.01fF
C37007 POR2X1_78/B POR2X1_231/O 0.02fF
C37008 PAND2X1_73/Y POR2X1_510/Y 0.03fF
C37009 POR2X1_56/B VDD 1.30fF
C37010 POR2X1_96/A POR2X1_305/a_76_344# 0.01fF
C37011 POR2X1_67/A POR2X1_283/A 0.03fF
C37012 POR2X1_197/CTRL2 POR2X1_740/Y 0.06fF
C37013 POR2X1_41/B POR2X1_13/A 0.58fF
C37014 PAND2X1_127/a_76_28# POR2X1_445/A 0.01fF
C37015 POR2X1_389/O POR2X1_480/A 0.01fF
C37016 POR2X1_83/B POR2X1_387/Y 0.07fF
C37017 PAND2X1_94/A PAND2X1_94/a_16_344# 0.02fF
C37018 PAND2X1_435/CTRL2 POR2X1_293/Y 0.01fF
C37019 POR2X1_121/B PAND2X1_305/CTRL 0.00fF
C37020 PAND2X1_592/Y INPUT_0 0.03fF
C37021 POR2X1_556/A POR2X1_362/O 0.01fF
C37022 POR2X1_330/Y PAND2X1_311/O 0.07fF
C37023 POR2X1_175/A POR2X1_570/B 0.03fF
C37024 PAND2X1_645/CTRL2 PAND2X1_602/Y 0.01fF
C37025 POR2X1_43/B PAND2X1_199/A 0.01fF
C37026 POR2X1_23/Y PAND2X1_579/A 0.01fF
C37027 PAND2X1_250/O PAND2X1_69/A 0.24fF
C37028 POR2X1_51/a_16_28# POR2X1_22/A 0.01fF
C37029 PAND2X1_90/Y PAND2X1_132/a_76_28# 0.02fF
C37030 POR2X1_453/CTRL2 PAND2X1_60/B 0.03fF
C37031 POR2X1_16/A POR2X1_409/B 0.03fF
C37032 PAND2X1_697/CTRL PAND2X1_90/Y 0.05fF
C37033 PAND2X1_58/A POR2X1_550/Y 0.06fF
C37034 PAND2X1_48/B POR2X1_244/B 0.03fF
C37035 PAND2X1_675/A POR2X1_236/Y 0.03fF
C37036 PAND2X1_23/Y POR2X1_241/Y 0.00fF
C37037 POR2X1_814/B PAND2X1_69/A 0.26fF
C37038 PAND2X1_411/CTRL2 POR2X1_461/B 0.00fF
C37039 POR2X1_283/A POR2X1_226/O 0.01fF
C37040 POR2X1_197/CTRL PAND2X1_56/Y 0.02fF
C37041 POR2X1_49/Y POR2X1_38/Y 0.22fF
C37042 PAND2X1_71/CTRL2 POR2X1_579/Y 0.00fF
C37043 POR2X1_330/Y POR2X1_541/a_16_28# 0.02fF
C37044 POR2X1_48/A PAND2X1_348/m4_208_n4# 0.12fF
C37045 PAND2X1_469/B POR2X1_236/Y 0.00fF
C37046 POR2X1_403/Y POR2X1_35/Y 0.02fF
C37047 POR2X1_66/A POR2X1_721/O 0.01fF
C37048 PAND2X1_382/a_76_28# POR2X1_29/A 0.02fF
C37049 POR2X1_26/CTRL2 POR2X1_32/A 0.03fF
C37050 POR2X1_186/Y POR2X1_724/A 0.07fF
C37051 D_GATE_811 VDD 0.04fF
C37052 POR2X1_458/Y POR2X1_717/B 0.03fF
C37053 PAND2X1_342/CTRL POR2X1_5/Y 0.02fF
C37054 PAND2X1_725/A VDD 0.00fF
C37055 POR2X1_141/Y PAND2X1_60/B 0.03fF
C37056 POR2X1_853/CTRL POR2X1_785/A 0.01fF
C37057 POR2X1_341/A PAND2X1_323/a_16_344# 0.04fF
C37058 PAND2X1_96/B POR2X1_805/B 0.17fF
C37059 PAND2X1_472/B POR2X1_42/Y 0.07fF
C37060 POR2X1_38/Y PAND2X1_558/CTRL2 0.01fF
C37061 POR2X1_471/A POR2X1_181/CTRL2 0.02fF
C37062 POR2X1_708/CTRL POR2X1_779/A 0.01fF
C37063 POR2X1_78/B PAND2X1_81/CTRL 0.02fF
C37064 PAND2X1_393/CTRL2 PAND2X1_41/B 0.02fF
C37065 POR2X1_188/A POR2X1_121/a_56_344# 0.00fF
C37066 POR2X1_16/A PAND2X1_794/CTRL -0.01fF
C37067 PAND2X1_69/A POR2X1_325/A 0.06fF
C37068 POR2X1_14/Y POR2X1_754/CTRL 0.03fF
C37069 POR2X1_73/CTRL POR2X1_40/Y 0.01fF
C37070 POR2X1_48/A POR2X1_183/CTRL 0.01fF
C37071 PAND2X1_629/CTRL POR2X1_7/A 0.01fF
C37072 PAND2X1_106/CTRL2 POR2X1_105/Y 0.01fF
C37073 POR2X1_806/CTRL POR2X1_675/Y 0.01fF
C37074 PAND2X1_74/CTRL2 POR2X1_456/B 0.01fF
C37075 POR2X1_675/A PAND2X1_60/B 0.01fF
C37076 POR2X1_52/A POR2X1_315/CTRL2 0.01fF
C37077 POR2X1_95/a_56_344# POR2X1_12/A 0.00fF
C37078 POR2X1_55/Y POR2X1_42/Y 0.65fF
C37079 POR2X1_78/A POR2X1_590/Y 0.01fF
C37080 PAND2X1_23/Y PAND2X1_95/B 0.03fF
C37081 POR2X1_332/B POR2X1_804/A 0.38fF
C37082 POR2X1_857/B POR2X1_350/O 0.01fF
C37083 POR2X1_614/A PAND2X1_71/CTRL2 0.05fF
C37084 POR2X1_164/Y POR2X1_72/B 0.98fF
C37085 POR2X1_540/A VDD 0.23fF
C37086 POR2X1_43/B POR2X1_586/a_56_344# 0.00fF
C37087 POR2X1_750/B POR2X1_750/Y 3.55fF
C37088 PAND2X1_824/B PAND2X1_20/A 0.03fF
C37089 PAND2X1_370/m4_208_n4# PAND2X1_352/m4_208_n4# 0.13fF
C37090 POR2X1_32/A PAND2X1_123/Y 0.04fF
C37091 PAND2X1_93/a_16_344# POR2X1_404/Y 0.02fF
C37092 PAND2X1_55/Y POR2X1_659/O 0.01fF
C37093 PAND2X1_69/A PAND2X1_176/CTRL2 0.01fF
C37094 POR2X1_113/A PAND2X1_20/A 0.00fF
C37095 POR2X1_163/Y PAND2X1_725/O 0.03fF
C37096 PAND2X1_730/O POR2X1_42/Y 0.05fF
C37097 PAND2X1_563/A PAND2X1_554/CTRL 0.01fF
C37098 POR2X1_221/Y POR2X1_222/Y 0.00fF
C37099 POR2X1_284/CTRL POR2X1_804/A 0.01fF
C37100 POR2X1_43/B PAND2X1_197/Y 0.05fF
C37101 POR2X1_55/Y POR2X1_309/Y 0.03fF
C37102 PAND2X1_480/B PAND2X1_702/O 0.04fF
C37103 POR2X1_333/A PAND2X1_745/a_16_344# 0.04fF
C37104 POR2X1_130/A POR2X1_137/Y 0.01fF
C37105 POR2X1_41/B PAND2X1_661/B 0.03fF
C37106 POR2X1_763/Y PAND2X1_324/CTRL2 0.01fF
C37107 POR2X1_49/Y INPUT_1 0.09fF
C37108 POR2X1_804/A PAND2X1_369/CTRL2 0.05fF
C37109 POR2X1_632/CTRL2 POR2X1_632/Y 0.01fF
C37110 POR2X1_65/A PAND2X1_539/Y 0.02fF
C37111 PAND2X1_6/Y POR2X1_733/A 0.07fF
C37112 POR2X1_45/Y POR2X1_273/Y 0.03fF
C37113 PAND2X1_6/Y POR2X1_334/B 0.05fF
C37114 POR2X1_81/a_16_28# POR2X1_153/Y 0.03fF
C37115 PAND2X1_407/a_76_28# POR2X1_39/B 0.04fF
C37116 POR2X1_62/O PAND2X1_6/A 0.16fF
C37117 PAND2X1_132/O PAND2X1_32/B 0.15fF
C37118 PAND2X1_864/O PAND2X1_805/A 0.06fF
C37119 POR2X1_539/A VDD 0.19fF
C37120 POR2X1_537/A VDD 0.00fF
C37121 POR2X1_220/Y PAND2X1_60/B 0.06fF
C37122 POR2X1_325/CTRL2 POR2X1_502/A 0.01fF
C37123 POR2X1_119/Y PAND2X1_443/Y 0.02fF
C37124 POR2X1_634/A PAND2X1_18/B 0.05fF
C37125 POR2X1_199/a_16_28# POR2X1_196/Y 0.07fF
C37126 POR2X1_78/B POR2X1_259/O 0.03fF
C37127 PAND2X1_824/B POR2X1_814/B 0.21fF
C37128 POR2X1_748/A PAND2X1_156/A 0.61fF
C37129 POR2X1_409/Y POR2X1_5/Y 0.04fF
C37130 POR2X1_36/B POR2X1_7/B 0.00fF
C37131 POR2X1_49/Y POR2X1_153/Y 0.07fF
C37132 POR2X1_123/A POR2X1_502/A 0.05fF
C37133 D_INPUT_5 PAND2X1_72/A 0.03fF
C37134 POR2X1_140/B POR2X1_513/Y -0.00fF
C37135 POR2X1_38/Y PAND2X1_188/O 0.01fF
C37136 POR2X1_404/Y PAND2X1_60/B 0.03fF
C37137 POR2X1_447/B PAND2X1_626/O 0.09fF
C37138 POR2X1_423/Y POR2X1_183/CTRL2 0.01fF
C37139 PAND2X1_464/Y PAND2X1_477/B 0.01fF
C37140 PAND2X1_534/CTRL2 POR2X1_294/B 0.05fF
C37141 POR2X1_260/Y POR2X1_359/Y 0.00fF
C37142 POR2X1_740/Y POR2X1_318/A 0.10fF
C37143 POR2X1_556/Y POR2X1_562/B 0.05fF
C37144 POR2X1_786/Y POR2X1_702/A 0.02fF
C37145 POR2X1_57/A POR2X1_693/Y 0.01fF
C37146 POR2X1_57/A PAND2X1_398/O 0.01fF
C37147 POR2X1_491/Y POR2X1_32/A 0.01fF
C37148 POR2X1_40/Y POR2X1_183/a_16_28# -0.00fF
C37149 PAND2X1_319/B POR2X1_312/CTRL 0.06fF
C37150 POR2X1_210/Y POR2X1_782/A 0.03fF
C37151 PAND2X1_790/Y POR2X1_7/A 0.04fF
C37152 POR2X1_62/Y PAND2X1_786/a_76_28# 0.04fF
C37153 PAND2X1_273/CTRL PAND2X1_60/B 0.03fF
C37154 POR2X1_254/Y POR2X1_332/CTRL2 0.03fF
C37155 POR2X1_741/a_16_28# POR2X1_741/A 0.11fF
C37156 POR2X1_652/Y POR2X1_799/CTRL 0.01fF
C37157 POR2X1_376/B PAND2X1_708/O 0.03fF
C37158 POR2X1_350/a_16_28# POR2X1_341/Y 0.03fF
C37159 POR2X1_447/B POR2X1_750/B 0.11fF
C37160 INPUT_1 POR2X1_586/CTRL2 0.01fF
C37161 POR2X1_497/Y POR2X1_394/A 0.07fF
C37162 PAND2X1_664/a_16_344# POR2X1_73/Y 0.02fF
C37163 PAND2X1_215/B PAND2X1_723/A 0.10fF
C37164 POR2X1_590/A POR2X1_39/B 0.03fF
C37165 POR2X1_416/B POR2X1_609/Y 0.03fF
C37166 POR2X1_785/a_16_28# POR2X1_785/B 0.05fF
C37167 POR2X1_220/Y POR2X1_353/A 0.03fF
C37168 PAND2X1_251/O POR2X1_717/B 0.02fF
C37169 PAND2X1_96/B POR2X1_190/CTRL 0.01fF
C37170 POR2X1_192/Y POR2X1_444/Y 0.01fF
C37171 PAND2X1_90/A PAND2X1_133/CTRL 0.01fF
C37172 POR2X1_13/A PAND2X1_308/Y 0.64fF
C37173 POR2X1_465/B POR2X1_456/B 0.18fF
C37174 POR2X1_539/A POR2X1_741/Y 0.03fF
C37175 PAND2X1_65/B POR2X1_294/A 0.42fF
C37176 POR2X1_140/B POR2X1_366/A 0.03fF
C37177 POR2X1_383/A POR2X1_713/O 0.03fF
C37178 POR2X1_89/Y PAND2X1_333/Y 0.04fF
C37179 PAND2X1_274/O POR2X1_153/Y 0.17fF
C37180 POR2X1_619/A POR2X1_751/CTRL2 0.10fF
C37181 POR2X1_707/CTRL PAND2X1_95/B 0.01fF
C37182 PAND2X1_70/O PAND2X1_3/B 0.05fF
C37183 POR2X1_334/O POR2X1_404/Y 0.01fF
C37184 POR2X1_8/Y POR2X1_143/a_56_344# 0.00fF
C37185 PAND2X1_631/A PAND2X1_456/O 0.07fF
C37186 POR2X1_848/A POR2X1_90/O 0.04fF
C37187 PAND2X1_659/Y PAND2X1_204/O 0.15fF
C37188 PAND2X1_56/Y POR2X1_787/CTRL2 0.16fF
C37189 POR2X1_470/O PAND2X1_52/B 0.10fF
C37190 PAND2X1_317/Y POR2X1_313/Y 0.01fF
C37191 PAND2X1_126/O PAND2X1_6/A 0.11fF
C37192 INPUT_1 POR2X1_669/m4_208_n4# 0.15fF
C37193 PAND2X1_467/O PAND2X1_725/A 0.00fF
C37194 PAND2X1_115/B PAND2X1_348/A 0.00fF
C37195 POR2X1_73/Y PAND2X1_656/A 0.10fF
C37196 POR2X1_711/CTRL2 POR2X1_713/B 0.00fF
C37197 POR2X1_539/A PAND2X1_32/B 0.03fF
C37198 POR2X1_537/A PAND2X1_32/B 0.10fF
C37199 INPUT_1 POR2X1_817/Y 0.01fF
C37200 POR2X1_575/O POR2X1_573/A 0.02fF
C37201 POR2X1_170/a_16_28# POR2X1_169/Y 0.03fF
C37202 PAND2X1_388/Y POR2X1_142/Y 0.03fF
C37203 PAND2X1_177/CTRL2 POR2X1_180/A 0.01fF
C37204 POR2X1_13/A PAND2X1_141/CTRL 0.01fF
C37205 POR2X1_46/Y PAND2X1_716/B 0.03fF
C37206 POR2X1_467/Y POR2X1_728/A 0.66fF
C37207 PAND2X1_476/A INPUT_0 0.05fF
C37208 PAND2X1_281/a_16_344# POR2X1_121/Y 0.01fF
C37209 POR2X1_7/B PAND2X1_365/A 0.06fF
C37210 POR2X1_88/Y POR2X1_4/Y 0.03fF
C37211 PAND2X1_738/A PAND2X1_149/A 0.02fF
C37212 POR2X1_782/A POR2X1_782/B 0.02fF
C37213 PAND2X1_641/CTRL POR2X1_38/Y 0.07fF
C37214 POR2X1_670/CTRL POR2X1_77/Y 0.03fF
C37215 POR2X1_576/CTRL POR2X1_500/Y 0.01fF
C37216 POR2X1_837/B PAND2X1_419/CTRL2 0.03fF
C37217 PAND2X1_562/B POR2X1_77/Y 0.20fF
C37218 PAND2X1_48/B POR2X1_722/CTRL 0.01fF
C37219 POR2X1_68/A POR2X1_673/B 0.20fF
C37220 POR2X1_390/B POR2X1_865/B 0.03fF
C37221 PAND2X1_481/a_16_344# POR2X1_222/Y 0.02fF
C37222 POR2X1_235/O POR2X1_7/A 0.01fF
C37223 POR2X1_366/CTRL PAND2X1_60/B 0.01fF
C37224 POR2X1_129/Y POR2X1_56/Y 0.03fF
C37225 POR2X1_750/O POR2X1_750/Y 0.02fF
C37226 PAND2X1_244/B PAND2X1_656/A 0.05fF
C37227 POR2X1_316/Y POR2X1_516/B 0.07fF
C37228 POR2X1_38/Y PAND2X1_121/m4_208_n4# 0.08fF
C37229 POR2X1_590/CTRL2 POR2X1_796/A 0.01fF
C37230 PAND2X1_726/B POR2X1_152/Y 0.36fF
C37231 POR2X1_833/A PAND2X1_150/O 0.09fF
C37232 POR2X1_252/Y POR2X1_55/Y 0.01fF
C37233 POR2X1_62/Y POR2X1_43/B 3.39fF
C37234 POR2X1_750/B POR2X1_181/A 0.01fF
C37235 PAND2X1_437/CTRL POR2X1_590/A 0.01fF
C37236 POR2X1_542/B POR2X1_186/B 0.03fF
C37237 PAND2X1_93/B PAND2X1_85/O 0.02fF
C37238 D_INPUT_3 POR2X1_4/CTRL 0.01fF
C37239 POR2X1_356/A PAND2X1_167/a_16_344# 0.12fF
C37240 POR2X1_614/A POR2X1_62/Y 0.12fF
C37241 PAND2X1_60/B POR2X1_332/CTRL 0.11fF
C37242 POR2X1_567/B POR2X1_814/A 0.10fF
C37243 PAND2X1_56/Y POR2X1_99/B 0.03fF
C37244 POR2X1_81/A POR2X1_494/Y 0.12fF
C37245 PAND2X1_511/CTRL PAND2X1_56/A 0.01fF
C37246 POR2X1_228/a_76_344# POR2X1_631/B 0.00fF
C37247 PAND2X1_321/a_16_344# PAND2X1_52/B 0.01fF
C37248 POR2X1_13/A POR2X1_77/Y 2.59fF
C37249 POR2X1_20/B POR2X1_299/a_16_28# 0.03fF
C37250 PAND2X1_6/Y POR2X1_349/O 0.18fF
C37251 POR2X1_7/B POR2X1_588/CTRL2 0.01fF
C37252 PAND2X1_290/CTRL2 POR2X1_334/B 0.09fF
C37253 POR2X1_7/A POR2X1_7/a_16_28# 0.03fF
C37254 POR2X1_609/Y PAND2X1_608/CTRL 0.00fF
C37255 POR2X1_762/O D_INPUT_6 0.01fF
C37256 INPUT_3 POR2X1_24/Y 0.05fF
C37257 POR2X1_568/Y POR2X1_444/Y 0.05fF
C37258 POR2X1_669/B POR2X1_667/CTRL -0.04fF
C37259 PAND2X1_793/Y PAND2X1_861/B 0.03fF
C37260 PAND2X1_775/O POR2X1_77/Y 0.03fF
C37261 POR2X1_730/Y POR2X1_260/A 0.03fF
C37262 PAND2X1_527/CTRL PAND2X1_111/B 0.01fF
C37263 POR2X1_677/Y PAND2X1_390/Y 0.04fF
C37264 POR2X1_431/a_16_28# POR2X1_37/Y 0.02fF
C37265 PAND2X1_690/CTRL POR2X1_260/A 0.01fF
C37266 POR2X1_383/A POR2X1_579/B 0.01fF
C37267 POR2X1_591/Y POR2X1_7/Y 0.03fF
C37268 PAND2X1_631/A POR2X1_73/Y 0.03fF
C37269 POR2X1_271/O POR2X1_411/B 0.01fF
C37270 PAND2X1_160/CTRL2 POR2X1_394/A 0.01fF
C37271 POR2X1_553/CTRL POR2X1_569/A 0.08fF
C37272 PAND2X1_608/O POR2X1_102/Y 0.02fF
C37273 PAND2X1_79/Y PAND2X1_527/m4_208_n4# 0.09fF
C37274 POR2X1_257/A POR2X1_248/A 0.05fF
C37275 POR2X1_270/a_76_344# POR2X1_567/A 0.00fF
C37276 POR2X1_86/CTRL POR2X1_73/Y 0.01fF
C37277 POR2X1_659/A POR2X1_222/O 0.06fF
C37278 POR2X1_383/A POR2X1_571/Y 0.06fF
C37279 POR2X1_864/A POR2X1_801/B 0.00fF
C37280 POR2X1_415/A POR2X1_818/Y 0.00fF
C37281 POR2X1_616/Y POR2X1_283/A 0.03fF
C37282 POR2X1_663/B POR2X1_66/A 0.03fF
C37283 POR2X1_20/B PAND2X1_722/CTRL 0.01fF
C37284 POR2X1_760/A POR2X1_594/O 0.01fF
C37285 POR2X1_463/O POR2X1_750/B 0.01fF
C37286 POR2X1_813/a_56_344# POR2X1_263/Y 0.00fF
C37287 POR2X1_180/B POR2X1_540/Y 0.09fF
C37288 POR2X1_841/O POR2X1_590/A 0.01fF
C37289 POR2X1_383/A PAND2X1_304/CTRL 0.01fF
C37290 PAND2X1_643/Y POR2X1_77/Y 0.03fF
C37291 PAND2X1_61/Y POR2X1_329/A 0.09fF
C37292 PAND2X1_634/CTRL POR2X1_607/A 0.00fF
C37293 POR2X1_411/B POR2X1_226/CTRL 0.01fF
C37294 POR2X1_83/B POR2X1_431/Y 0.03fF
C37295 POR2X1_646/a_76_344# PAND2X1_90/Y 0.01fF
C37296 POR2X1_346/B POR2X1_61/A 0.00fF
C37297 INPUT_1 POR2X1_397/a_56_344# 0.00fF
C37298 POR2X1_250/Y POR2X1_488/O 0.03fF
C37299 POR2X1_3/A POR2X1_416/B 0.05fF
C37300 PAND2X1_358/CTRL PAND2X1_656/A 0.01fF
C37301 D_INPUT_5 PAND2X1_752/O 0.17fF
C37302 PAND2X1_35/A PAND2X1_34/CTRL 0.01fF
C37303 PAND2X1_207/A PAND2X1_656/A 0.03fF
C37304 POR2X1_8/Y POR2X1_4/Y 0.24fF
C37305 POR2X1_78/B POR2X1_814/A 0.17fF
C37306 PAND2X1_644/CTRL POR2X1_236/Y 0.04fF
C37307 POR2X1_116/A POR2X1_777/B 0.03fF
C37308 POR2X1_506/a_16_28# POR2X1_447/B -0.00fF
C37309 POR2X1_23/Y D_INPUT_0 0.17fF
C37310 POR2X1_38/a_76_344# POR2X1_37/Y 0.01fF
C37311 POR2X1_450/Y POR2X1_121/B 0.04fF
C37312 POR2X1_49/Y PAND2X1_201/a_76_28# 0.02fF
C37313 POR2X1_20/B PAND2X1_211/A 0.00fF
C37314 PAND2X1_199/CTRL2 PAND2X1_123/Y 0.01fF
C37315 POR2X1_77/Y PAND2X1_510/B 0.05fF
C37316 PAND2X1_830/O POR2X1_416/B 0.02fF
C37317 POR2X1_441/Y PAND2X1_803/A 0.00fF
C37318 PAND2X1_466/A POR2X1_236/Y 0.02fF
C37319 POR2X1_378/a_76_344# PAND2X1_9/Y 0.00fF
C37320 POR2X1_840/B POR2X1_76/B 0.03fF
C37321 PAND2X1_445/Y PAND2X1_464/B 0.05fF
C37322 PAND2X1_797/Y POR2X1_373/Y 0.03fF
C37323 POR2X1_78/A POR2X1_807/CTRL 0.01fF
C37324 POR2X1_67/Y POR2X1_7/B 0.03fF
C37325 POR2X1_82/CTRL2 PAND2X1_9/Y 0.01fF
C37326 POR2X1_466/A POR2X1_454/B 0.01fF
C37327 PAND2X1_39/B POR2X1_405/a_16_28# 0.10fF
C37328 POR2X1_862/Y POR2X1_777/B 0.02fF
C37329 POR2X1_650/A POR2X1_473/CTRL 0.09fF
C37330 POR2X1_416/B PAND2X1_317/O 0.02fF
C37331 PAND2X1_267/O POR2X1_72/B 0.05fF
C37332 PAND2X1_628/CTRL PAND2X1_88/Y 0.01fF
C37333 PAND2X1_267/B VDD 0.05fF
C37334 POR2X1_497/O POR2X1_37/Y 0.05fF
C37335 PAND2X1_353/Y PAND2X1_352/Y 0.03fF
C37336 POR2X1_651/Y PAND2X1_60/B 0.12fF
C37337 POR2X1_362/Y POR2X1_296/B 0.11fF
C37338 PAND2X1_406/CTRL2 POR2X1_362/B 0.01fF
C37339 POR2X1_96/A POR2X1_20/B 26.96fF
C37340 POR2X1_54/Y PAND2X1_293/CTRL2 0.07fF
C37341 POR2X1_567/B POR2X1_852/B 0.07fF
C37342 PAND2X1_443/Y POR2X1_442/Y 0.06fF
C37343 PAND2X1_439/CTRL2 POR2X1_90/Y 0.00fF
C37344 POR2X1_260/B PAND2X1_381/O 0.04fF
C37345 POR2X1_329/A POR2X1_255/Y 0.19fF
C37346 PAND2X1_66/a_16_344# POR2X1_5/Y 0.01fF
C37347 POR2X1_828/Y POR2X1_678/Y 0.13fF
C37348 POR2X1_290/CTRL POR2X1_37/Y 0.28fF
C37349 POR2X1_815/A VDD 0.00fF
C37350 POR2X1_25/Y POR2X1_416/B 0.03fF
C37351 PAND2X1_436/CTRL INPUT_0 0.03fF
C37352 PAND2X1_23/Y POR2X1_444/O 0.01fF
C37353 POR2X1_418/Y POR2X1_14/Y 0.01fF
C37354 POR2X1_754/Y POR2X1_625/CTRL2 0.06fF
C37355 POR2X1_849/B VDD 0.10fF
C37356 POR2X1_78/A POR2X1_186/Y 0.11fF
C37357 POR2X1_168/CTRL2 POR2X1_168/A 0.01fF
C37358 POR2X1_118/Y VDD 0.11fF
C37359 PAND2X1_286/B PAND2X1_286/O 0.00fF
C37360 POR2X1_311/Y POR2X1_331/Y 0.01fF
C37361 PAND2X1_20/A POR2X1_640/Y 0.03fF
C37362 PAND2X1_203/CTRL PAND2X1_575/A 0.09fF
C37363 PAND2X1_658/O POR2X1_60/A 0.04fF
C37364 POR2X1_287/A POR2X1_513/Y 0.11fF
C37365 POR2X1_399/CTRL POR2X1_609/Y 0.03fF
C37366 POR2X1_492/CTRL POR2X1_60/A 0.01fF
C37367 POR2X1_109/CTRL2 POR2X1_7/B 0.00fF
C37368 POR2X1_490/Y POR2X1_46/Y 0.03fF
C37369 POR2X1_812/A POR2X1_801/CTRL2 0.01fF
C37370 POR2X1_52/A POR2X1_89/CTRL2 0.02fF
C37371 POR2X1_179/O POR2X1_411/B 0.02fF
C37372 PAND2X1_73/Y POR2X1_780/a_16_28# 0.03fF
C37373 POR2X1_52/A PAND2X1_97/CTRL2 0.03fF
C37374 POR2X1_669/Y POR2X1_73/Y 0.10fF
C37375 PAND2X1_263/CTRL2 POR2X1_78/A 0.03fF
C37376 POR2X1_620/CTRL PAND2X1_9/Y 0.01fF
C37377 POR2X1_709/A POR2X1_790/B 0.03fF
C37378 POR2X1_253/CTRL2 PAND2X1_6/A 0.13fF
C37379 PAND2X1_472/A POR2X1_411/B 0.03fF
C37380 POR2X1_48/CTRL POR2X1_32/A 0.01fF
C37381 POR2X1_66/B PAND2X1_16/CTRL 0.01fF
C37382 POR2X1_288/A POR2X1_288/a_16_28# 0.09fF
C37383 PAND2X1_853/B POR2X1_173/Y 0.04fF
C37384 POR2X1_49/Y PAND2X1_214/A 0.02fF
C37385 POR2X1_632/B POR2X1_632/A 0.01fF
C37386 PAND2X1_766/CTRL2 PAND2X1_41/B 0.10fF
C37387 PAND2X1_39/B POR2X1_723/B 0.33fF
C37388 POR2X1_473/CTRL2 POR2X1_391/Y 0.05fF
C37389 PAND2X1_255/O POR2X1_260/A 0.03fF
C37390 POR2X1_423/O POR2X1_236/Y 0.01fF
C37391 POR2X1_450/O VDD 0.00fF
C37392 POR2X1_290/a_16_28# POR2X1_83/B -0.00fF
C37393 POR2X1_624/Y POR2X1_565/O 0.00fF
C37394 POR2X1_665/a_16_28# POR2X1_665/A 0.10fF
C37395 PAND2X1_60/O POR2X1_61/B 0.08fF
C37396 POR2X1_247/Y VDD 0.01fF
C37397 POR2X1_566/A POR2X1_97/A 0.16fF
C37398 POR2X1_68/A POR2X1_445/A 0.16fF
C37399 PAND2X1_863/a_76_28# POR2X1_102/Y 0.01fF
C37400 POR2X1_830/O POR2X1_830/A 0.03fF
C37401 POR2X1_83/B POR2X1_237/O 0.01fF
C37402 POR2X1_329/A POR2X1_385/O 0.09fF
C37403 PAND2X1_73/m4_208_n4# PAND2X1_41/B 0.07fF
C37404 PAND2X1_95/B PAND2X1_31/O 0.02fF
C37405 POR2X1_57/A POR2X1_744/Y 0.01fF
C37406 PAND2X1_271/O POR2X1_513/Y 0.07fF
C37407 PAND2X1_573/B VDD 0.00fF
C37408 PAND2X1_250/CTRL POR2X1_287/B 0.01fF
C37409 POR2X1_856/B POR2X1_785/A 0.05fF
C37410 POR2X1_360/A PAND2X1_15/CTRL2 0.04fF
C37411 PAND2X1_850/Y POR2X1_589/Y 0.02fF
C37412 POR2X1_683/O POR2X1_669/B 0.01fF
C37413 POR2X1_446/B POR2X1_112/Y 0.03fF
C37414 INPUT_3 POR2X1_619/Y 0.00fF
C37415 POR2X1_119/Y PAND2X1_860/A 0.03fF
C37416 POR2X1_54/Y POR2X1_68/B 1.52fF
C37417 POR2X1_32/A INPUT_5 0.02fF
C37418 PAND2X1_455/Y POR2X1_14/Y 0.02fF
C37419 POR2X1_199/CTRL POR2X1_590/A 0.01fF
C37420 POR2X1_14/Y POR2X1_415/O 0.06fF
C37421 PAND2X1_319/O PAND2X1_354/A 0.01fF
C37422 POR2X1_89/Y POR2X1_293/Y 0.02fF
C37423 POR2X1_516/CTRL2 POR2X1_48/A 0.01fF
C37424 POR2X1_516/CTRL POR2X1_23/Y 0.04fF
C37425 POR2X1_20/B POR2X1_7/A 0.17fF
C37426 PAND2X1_90/A PAND2X1_277/a_76_28# 0.02fF
C37427 POR2X1_517/Y POR2X1_669/B 0.02fF
C37428 PAND2X1_863/B PAND2X1_249/CTRL2 0.01fF
C37429 POR2X1_33/B VDD 0.17fF
C37430 POR2X1_366/Y POR2X1_269/O 0.01fF
C37431 PAND2X1_23/Y POR2X1_843/CTRL 0.04fF
C37432 INPUT_7 POR2X1_763/A 0.07fF
C37433 POR2X1_20/B PAND2X1_344/a_76_28# 0.02fF
C37434 POR2X1_481/A POR2X1_40/Y 0.01fF
C37435 POR2X1_52/A POR2X1_226/CTRL 0.01fF
C37436 POR2X1_67/A POR2X1_55/Y 0.01fF
C37437 PAND2X1_473/Y POR2X1_72/B 0.01fF
C37438 POR2X1_438/Y POR2X1_90/Y 0.00fF
C37439 POR2X1_662/Y POR2X1_590/A 0.94fF
C37440 POR2X1_102/Y PAND2X1_174/CTRL2 0.01fF
C37441 POR2X1_39/B POR2X1_90/CTRL 0.01fF
C37442 PAND2X1_20/A PAND2X1_226/CTRL 0.00fF
C37443 PAND2X1_630/CTRL POR2X1_496/Y 0.07fF
C37444 POR2X1_37/Y POR2X1_56/Y 0.10fF
C37445 PAND2X1_362/A POR2X1_42/Y 0.04fF
C37446 POR2X1_567/B POR2X1_190/CTRL2 0.16fF
C37447 POR2X1_290/Y POR2X1_607/A 0.00fF
C37448 POR2X1_632/O PAND2X1_88/Y 0.01fF
C37449 POR2X1_220/Y POR2X1_750/B 0.06fF
C37450 POR2X1_549/A POR2X1_78/A 0.02fF
C37451 POR2X1_286/Y VDD 0.18fF
C37452 PAND2X1_289/m4_208_n4# POR2X1_220/A 0.07fF
C37453 POR2X1_674/Y PAND2X1_742/B 0.87fF
C37454 POR2X1_634/A POR2X1_638/O 0.24fF
C37455 PAND2X1_839/O POR2X1_102/Y 0.02fF
C37456 POR2X1_716/CTRL2 POR2X1_303/B 0.01fF
C37457 POR2X1_744/Y POR2X1_744/O 0.01fF
C37458 POR2X1_129/CTRL POR2X1_90/Y 0.00fF
C37459 POR2X1_130/A POR2X1_650/A 0.02fF
C37460 POR2X1_634/A POR2X1_294/B 0.01fF
C37461 POR2X1_29/A POR2X1_391/Y 0.10fF
C37462 PAND2X1_20/A PAND2X1_496/a_16_344# 0.02fF
C37463 PAND2X1_848/B PAND2X1_848/CTRL2 0.01fF
C37464 POR2X1_121/A POR2X1_78/A 0.00fF
C37465 POR2X1_814/A POR2X1_294/A 0.60fF
C37466 PAND2X1_621/CTRL2 POR2X1_415/A 0.05fF
C37467 POR2X1_523/Y POR2X1_819/O 0.01fF
C37468 POR2X1_123/B POR2X1_558/B 0.10fF
C37469 PAND2X1_403/Y VDD 0.12fF
C37470 POR2X1_647/B POR2X1_101/Y 0.07fF
C37471 POR2X1_356/A POR2X1_175/A 0.05fF
C37472 POR2X1_254/Y PAND2X1_48/Y 0.04fF
C37473 POR2X1_638/A POR2X1_638/a_16_28# 0.05fF
C37474 POR2X1_260/B POR2X1_780/B 0.01fF
C37475 PAND2X1_465/O PAND2X1_465/B 0.01fF
C37476 POR2X1_417/Y PAND2X1_724/B 0.02fF
C37477 POR2X1_712/A PAND2X1_73/Y 0.01fF
C37478 POR2X1_322/CTRL POR2X1_40/Y 0.12fF
C37479 POR2X1_180/B POR2X1_445/A 0.03fF
C37480 POR2X1_458/m4_208_n4# POR2X1_458/B 0.01fF
C37481 POR2X1_115/a_16_28# POR2X1_330/Y 0.08fF
C37482 POR2X1_196/m4_208_n4# POR2X1_740/Y 0.06fF
C37483 POR2X1_32/A PAND2X1_186/CTRL2 0.03fF
C37484 PAND2X1_833/a_76_28# POR2X1_376/B 0.03fF
C37485 PAND2X1_657/O POR2X1_816/A 0.01fF
C37486 PAND2X1_217/B PAND2X1_188/CTRL 0.01fF
C37487 POR2X1_633/Y VDD 0.09fF
C37488 PAND2X1_20/A PAND2X1_612/CTRL 0.03fF
C37489 POR2X1_763/A INPUT_4 0.08fF
C37490 PAND2X1_736/A POR2X1_72/B 0.07fF
C37491 POR2X1_62/Y PAND2X1_201/CTRL2 0.01fF
C37492 POR2X1_65/A PAND2X1_364/O 0.01fF
C37493 POR2X1_123/A POR2X1_493/A 0.01fF
C37494 PAND2X1_288/A PAND2X1_367/a_76_28# 0.04fF
C37495 D_INPUT_2 POR2X1_94/A 0.03fF
C37496 POR2X1_149/A PAND2X1_69/A 0.01fF
C37497 POR2X1_791/CTRL POR2X1_637/B 0.01fF
C37498 POR2X1_57/A PAND2X1_212/B 0.05fF
C37499 PAND2X1_26/A POR2X1_260/A 1.24fF
C37500 POR2X1_624/Y POR2X1_244/Y 0.07fF
C37501 PAND2X1_20/A POR2X1_139/A 0.00fF
C37502 POR2X1_807/A POR2X1_832/B 0.03fF
C37503 PAND2X1_564/B POR2X1_73/Y 0.02fF
C37504 PAND2X1_246/O POR2X1_4/Y 0.02fF
C37505 POR2X1_224/Y POR2X1_226/Y 0.13fF
C37506 PAND2X1_454/CTRL2 POR2X1_511/Y 0.03fF
C37507 POR2X1_60/A PAND2X1_389/a_16_344# 0.02fF
C37508 POR2X1_623/A POR2X1_623/O 0.01fF
C37509 POR2X1_300/a_76_344# PAND2X1_217/B 0.03fF
C37510 PAND2X1_735/CTRL2 POR2X1_293/Y 0.03fF
C37511 PAND2X1_499/Y POR2X1_494/Y 0.05fF
C37512 D_INPUT_3 POR2X1_83/B 0.13fF
C37513 PAND2X1_371/CTRL VDD 0.00fF
C37514 PAND2X1_787/Y PAND2X1_390/CTRL 0.02fF
C37515 POR2X1_376/B PAND2X1_242/O 0.04fF
C37516 PAND2X1_6/Y POR2X1_593/B 0.04fF
C37517 PAND2X1_223/B PAND2X1_854/A 0.02fF
C37518 POR2X1_360/A INPUT_0 0.10fF
C37519 PAND2X1_288/A VDD 0.15fF
C37520 PAND2X1_715/CTRL2 PAND2X1_115/B 0.03fF
C37521 POR2X1_814/B POR2X1_723/B 0.04fF
C37522 PAND2X1_245/CTRL PAND2X1_63/B 0.01fF
C37523 PAND2X1_839/B POR2X1_102/Y 0.01fF
C37524 PAND2X1_864/B GATE_741 0.00fF
C37525 PAND2X1_438/CTRL PAND2X1_72/A 0.01fF
C37526 PAND2X1_119/m4_208_n4# POR2X1_78/A 0.08fF
C37527 PAND2X1_48/B POR2X1_115/CTRL2 0.01fF
C37528 POR2X1_668/CTRL2 POR2X1_816/A 0.05fF
C37529 POR2X1_504/Y POR2X1_90/Y 0.07fF
C37530 POR2X1_383/A PAND2X1_531/O 0.07fF
C37531 POR2X1_130/A POR2X1_294/B 0.06fF
C37532 PAND2X1_852/O POR2X1_122/Y 0.04fF
C37533 PAND2X1_73/Y POR2X1_598/CTRL 0.01fF
C37534 POR2X1_566/A POR2X1_294/B 0.05fF
C37535 POR2X1_49/Y POR2X1_591/Y 0.03fF
C37536 POR2X1_68/A PAND2X1_58/CTRL 0.01fF
C37537 POR2X1_366/Y POR2X1_566/A 0.10fF
C37538 POR2X1_153/CTRL POR2X1_37/Y 0.01fF
C37539 POR2X1_646/B PAND2X1_56/A 0.00fF
C37540 PAND2X1_217/B POR2X1_91/Y 0.03fF
C37541 POR2X1_61/B POR2X1_206/A 0.02fF
C37542 POR2X1_515/O POR2X1_68/A 0.34fF
C37543 POR2X1_706/CTRL2 INPUT_1 0.01fF
C37544 POR2X1_60/A PAND2X1_717/Y 0.03fF
C37545 POR2X1_197/Y POR2X1_244/O 0.01fF
C37546 POR2X1_14/Y PAND2X1_550/B 0.06fF
C37547 POR2X1_523/Y VDD 0.09fF
C37548 POR2X1_102/Y POR2X1_172/CTRL 0.01fF
C37549 POR2X1_706/B POR2X1_532/A 0.02fF
C37550 POR2X1_48/A POR2X1_749/O 0.01fF
C37551 POR2X1_664/O PAND2X1_73/Y 0.05fF
C37552 POR2X1_664/CTRL POR2X1_78/A 0.00fF
C37553 PAND2X1_408/CTRL VDD 0.00fF
C37554 POR2X1_856/B POR2X1_186/B 0.04fF
C37555 POR2X1_753/Y POR2X1_754/O 0.01fF
C37556 POR2X1_93/A PAND2X1_392/B 0.03fF
C37557 PAND2X1_48/B PAND2X1_152/O 0.03fF
C37558 PAND2X1_20/A POR2X1_576/CTRL 0.01fF
C37559 POR2X1_49/Y PAND2X1_470/A 0.02fF
C37560 POR2X1_330/Y POR2X1_569/A 0.07fF
C37561 POR2X1_391/Y POR2X1_546/A 0.04fF
C37562 POR2X1_855/B POR2X1_783/a_76_344# 0.00fF
C37563 POR2X1_850/B POR2X1_456/B 0.54fF
C37564 PAND2X1_69/A VDD 3.20fF
C37565 POR2X1_376/B PAND2X1_168/CTRL 0.01fF
C37566 PAND2X1_571/A PAND2X1_716/B 0.00fF
C37567 POR2X1_172/Y POR2X1_5/Y 0.21fF
C37568 POR2X1_52/A PAND2X1_242/O 0.01fF
C37569 PAND2X1_14/O POR2X1_68/B 0.05fF
C37570 POR2X1_256/O POR2X1_255/Y 0.13fF
C37571 POR2X1_61/Y POR2X1_510/Y 0.07fF
C37572 POR2X1_222/Y POR2X1_554/Y 0.03fF
C37573 POR2X1_13/A POR2X1_52/Y 0.02fF
C37574 POR2X1_661/A POR2X1_655/CTRL2 0.05fF
C37575 POR2X1_65/A POR2X1_167/CTRL 0.01fF
C37576 PAND2X1_341/A VDD 0.00fF
C37577 PAND2X1_80/O POR2X1_68/B 0.15fF
C37578 POR2X1_327/Y PAND2X1_73/Y 0.00fF
C37579 POR2X1_400/A POR2X1_206/O 0.01fF
C37580 PAND2X1_737/B POR2X1_40/Y 0.10fF
C37581 POR2X1_52/A POR2X1_518/Y 0.03fF
C37582 POR2X1_834/Y POR2X1_602/B 0.05fF
C37583 POR2X1_93/A VDD 0.63fF
C37584 POR2X1_445/A POR2X1_169/A 0.03fF
C37585 POR2X1_468/Y VDD 0.00fF
C37586 POR2X1_293/Y POR2X1_56/Y 0.07fF
C37587 PAND2X1_216/B POR2X1_40/Y 0.01fF
C37588 POR2X1_376/B POR2X1_527/Y 0.16fF
C37589 VDD POR2X1_91/Y 0.55fF
C37590 PAND2X1_239/a_76_28# POR2X1_192/B 0.03fF
C37591 PAND2X1_41/B PAND2X1_184/CTRL2 0.10fF
C37592 POR2X1_790/a_16_28# POR2X1_790/A 0.01fF
C37593 POR2X1_62/Y POR2X1_590/A 0.03fF
C37594 PAND2X1_371/CTRL PAND2X1_32/B 0.01fF
C37595 POR2X1_579/Y POR2X1_804/A 0.03fF
C37596 PAND2X1_197/O POR2X1_52/Y 0.15fF
C37597 POR2X1_294/B POR2X1_844/B 0.06fF
C37598 POR2X1_718/CTRL POR2X1_834/Y 0.14fF
C37599 PAND2X1_6/Y POR2X1_477/A 5.32fF
C37600 D_INPUT_0 POR2X1_691/A 0.01fF
C37601 POR2X1_10/a_16_28# POR2X1_40/Y 0.02fF
C37602 PAND2X1_662/CTRL POR2X1_413/A 0.01fF
C37603 POR2X1_640/O POR2X1_559/A 0.11fF
C37604 POR2X1_316/Y PAND2X1_776/Y 0.23fF
C37605 POR2X1_21/CTRL INPUT_4 0.07fF
C37606 POR2X1_532/A POR2X1_554/Y 0.38fF
C37607 POR2X1_655/A POR2X1_711/Y 0.03fF
C37608 PAND2X1_720/CTRL VDD 0.00fF
C37609 PAND2X1_844/CTRL POR2X1_60/Y 0.01fF
C37610 PAND2X1_341/A PAND2X1_101/CTRL2 0.01fF
C37611 POR2X1_48/A PAND2X1_346/O 0.04fF
C37612 PAND2X1_211/A PAND2X1_303/Y 0.03fF
C37613 POR2X1_416/B PAND2X1_606/CTRL 0.01fF
C37614 POR2X1_423/Y POR2X1_394/A 0.03fF
C37615 POR2X1_78/B PAND2X1_232/CTRL2 0.01fF
C37616 POR2X1_96/A POR2X1_134/CTRL2 0.02fF
C37617 POR2X1_428/CTRL POR2X1_236/Y 0.01fF
C37618 PAND2X1_69/A POR2X1_741/Y 0.08fF
C37619 PAND2X1_56/Y POR2X1_112/Y 0.03fF
C37620 PAND2X1_568/B POR2X1_7/B 0.03fF
C37621 PAND2X1_6/Y POR2X1_562/B 0.02fF
C37622 POR2X1_654/B POR2X1_557/B 0.16fF
C37623 PAND2X1_81/B PAND2X1_69/A 0.17fF
C37624 POR2X1_78/A POR2X1_542/Y 0.01fF
C37625 POR2X1_187/CTRL2 POR2X1_79/Y 0.01fF
C37626 POR2X1_220/Y POR2X1_200/A 0.09fF
C37627 PAND2X1_545/Y VDD 0.17fF
C37628 POR2X1_326/CTRL VDD -0.00fF
C37629 PAND2X1_488/CTRL2 POR2X1_294/A 0.03fF
C37630 PAND2X1_832/CTRL PAND2X1_508/Y 0.00fF
C37631 PAND2X1_408/CTRL PAND2X1_32/B 0.01fF
C37632 PAND2X1_823/O VDD 0.00fF
C37633 POR2X1_614/A POR2X1_804/A 0.03fF
C37634 INPUT_1 PAND2X1_8/Y 0.31fF
C37635 POR2X1_16/A PAND2X1_520/CTRL 0.00fF
C37636 PAND2X1_23/Y PAND2X1_757/O 0.05fF
C37637 POR2X1_644/A POR2X1_796/O 0.01fF
C37638 PAND2X1_29/CTRL POR2X1_68/B 0.06fF
C37639 POR2X1_832/A PAND2X1_55/Y 0.13fF
C37640 PAND2X1_798/Y POR2X1_283/a_16_28# 0.04fF
C37641 POR2X1_72/B POR2X1_7/Y 0.03fF
C37642 INPUT_6 POR2X1_587/Y 0.01fF
C37643 POR2X1_852/B POR2X1_294/A 0.02fF
C37644 POR2X1_502/A PAND2X1_698/O 0.07fF
C37645 PAND2X1_69/A PAND2X1_32/B 0.23fF
C37646 PAND2X1_824/B VDD 3.21fF
C37647 POR2X1_502/A POR2X1_463/Y 0.01fF
C37648 POR2X1_304/a_76_344# POR2X1_153/Y 0.01fF
C37649 POR2X1_514/O POR2X1_137/Y 0.02fF
C37650 POR2X1_637/B PAND2X1_48/A 0.05fF
C37651 PAND2X1_111/B PAND2X1_111/O 0.07fF
C37652 POR2X1_114/B PAND2X1_60/B 0.04fF
C37653 PAND2X1_653/Y POR2X1_38/Y 0.03fF
C37654 PAND2X1_490/O POR2X1_38/B 0.04fF
C37655 INPUT_1 POR2X1_20/CTRL2 0.00fF
C37656 POR2X1_67/Y PAND2X1_206/B 0.01fF
C37657 PAND2X1_11/Y D_INPUT_4 0.23fF
C37658 POR2X1_35/Y POR2X1_510/Y 0.03fF
C37659 PAND2X1_653/O POR2X1_83/B 0.03fF
C37660 POR2X1_29/A POR2X1_77/Y 0.09fF
C37661 PAND2X1_785/Y PAND2X1_348/A 0.05fF
C37662 PAND2X1_696/O POR2X1_602/B 0.02fF
C37663 POR2X1_203/CTRL POR2X1_203/Y 0.00fF
C37664 PAND2X1_449/CTRL2 POR2X1_329/A -0.02fF
C37665 POR2X1_336/a_16_28# PAND2X1_69/A 0.03fF
C37666 PAND2X1_735/Y PAND2X1_853/B 0.07fF
C37667 POR2X1_685/A POR2X1_68/A 0.04fF
C37668 POR2X1_113/CTRL PAND2X1_96/B 0.09fF
C37669 POR2X1_567/B POR2X1_535/CTRL2 0.01fF
C37670 POR2X1_845/CTRL D_INPUT_1 0.04fF
C37671 VDD POR2X1_109/Y 0.15fF
C37672 POR2X1_252/Y POR2X1_511/Y 0.04fF
C37673 PAND2X1_785/Y POR2X1_300/Y 0.05fF
C37674 PAND2X1_209/A PAND2X1_797/O 0.03fF
C37675 POR2X1_407/Y POR2X1_780/B 0.03fF
C37676 PAND2X1_57/B POR2X1_342/CTRL2 0.03fF
C37677 PAND2X1_823/a_76_28# POR2X1_857/B 0.02fF
C37678 POR2X1_116/A POR2X1_814/A 0.03fF
C37679 POR2X1_346/B D_GATE_222 0.03fF
C37680 POR2X1_741/Y PAND2X1_368/a_76_28# 0.02fF
C37681 PAND2X1_467/Y POR2X1_694/CTRL 0.01fF
C37682 PAND2X1_445/CTRL PAND2X1_308/Y 0.01fF
C37683 POR2X1_52/A PAND2X1_620/a_56_28# 0.00fF
C37684 POR2X1_523/Y POR2X1_673/Y 0.03fF
C37685 PAND2X1_723/a_56_28# PAND2X1_656/A 0.00fF
C37686 POR2X1_78/A POR2X1_717/B 0.04fF
C37687 POR2X1_38/Y POR2X1_235/O 0.03fF
C37688 POR2X1_68/A POR2X1_260/A 1.92fF
C37689 POR2X1_62/Y PAND2X1_350/A 0.01fF
C37690 POR2X1_13/A POR2X1_371/O 0.18fF
C37691 PAND2X1_637/CTRL2 PAND2X1_69/A 0.00fF
C37692 PAND2X1_824/B POR2X1_741/Y 0.10fF
C37693 PAND2X1_6/Y POR2X1_802/m4_208_n4# 0.08fF
C37694 POR2X1_84/Y PAND2X1_63/B 0.29fF
C37695 POR2X1_129/Y POR2X1_42/Y 0.39fF
C37696 POR2X1_548/a_16_28# POR2X1_4/Y 0.04fF
C37697 POR2X1_614/A PAND2X1_313/O 0.01fF
C37698 PAND2X1_563/O POR2X1_394/A 0.02fF
C37699 POR2X1_567/A POR2X1_566/A 0.13fF
C37700 PAND2X1_859/CTRL2 POR2X1_77/Y 0.01fF
C37701 PAND2X1_254/O PAND2X1_508/Y 0.00fF
C37702 POR2X1_222/A PAND2X1_60/B 0.03fF
C37703 PAND2X1_473/B POR2X1_589/O 0.01fF
C37704 PAND2X1_631/A PAND2X1_785/Y 0.07fF
C37705 POR2X1_673/Y PAND2X1_69/A 0.03fF
C37706 POR2X1_16/A POR2X1_234/a_16_28# 0.03fF
C37707 POR2X1_57/A POR2X1_291/CTRL2 0.03fF
C37708 POR2X1_330/Y PAND2X1_72/A 0.15fF
C37709 POR2X1_356/A POR2X1_337/Y 0.10fF
C37710 POR2X1_25/CTRL D_INPUT_4 0.01fF
C37711 POR2X1_8/Y D_INPUT_1 0.01fF
C37712 POR2X1_68/A POR2X1_363/A 0.10fF
C37713 POR2X1_460/A POR2X1_260/A 0.03fF
C37714 POR2X1_175/A PAND2X1_72/A 0.03fF
C37715 POR2X1_435/Y POR2X1_532/CTRL 0.07fF
C37716 POR2X1_68/A PAND2X1_142/O 0.12fF
C37717 PAND2X1_659/Y POR2X1_42/Y 0.03fF
C37718 D_INPUT_1 POR2X1_749/CTRL2 0.01fF
C37719 POR2X1_328/m4_208_n4# INPUT_4 0.07fF
C37720 PAND2X1_23/Y POR2X1_112/CTRL2 0.01fF
C37721 POR2X1_88/CTRL PAND2X1_206/B 0.01fF
C37722 POR2X1_785/A POR2X1_191/Y 0.05fF
C37723 POR2X1_534/O POR2X1_534/Y 0.01fF
C37724 POR2X1_118/O PAND2X1_560/B 0.01fF
C37725 PAND2X1_6/A PAND2X1_156/A 0.10fF
C37726 POR2X1_38/B POR2X1_6/O 0.34fF
C37727 POR2X1_101/Y POR2X1_218/CTRL2 0.10fF
C37728 POR2X1_416/B PAND2X1_193/O 0.09fF
C37729 PAND2X1_202/a_76_28# POR2X1_66/A 0.01fF
C37730 PAND2X1_300/a_76_28# PAND2X1_60/B 0.02fF
C37731 PAND2X1_75/O POR2X1_260/B 0.02fF
C37732 PAND2X1_687/B POR2X1_42/Y 0.01fF
C37733 POR2X1_96/A POR2X1_189/O 0.02fF
C37734 PAND2X1_319/B POR2X1_394/A 0.05fF
C37735 POR2X1_192/Y POR2X1_567/CTRL 0.01fF
C37736 PAND2X1_630/a_76_28# PAND2X1_156/A 0.03fF
C37737 PAND2X1_715/B POR2X1_7/A 0.01fF
C37738 POR2X1_730/Y POR2X1_725/Y 0.00fF
C37739 POR2X1_863/A PAND2X1_41/B 0.03fF
C37740 POR2X1_502/A POR2X1_736/A 0.05fF
C37741 POR2X1_383/A POR2X1_734/O 0.01fF
C37742 POR2X1_21/a_16_28# POR2X1_260/A 0.01fF
C37743 POR2X1_391/a_16_28# POR2X1_391/B 0.09fF
C37744 POR2X1_51/A POR2X1_64/CTRL2 0.01fF
C37745 PAND2X1_474/CTRL PAND2X1_404/Y 0.01fF
C37746 POR2X1_218/O POR2X1_216/Y 0.00fF
C37747 PAND2X1_96/B POR2X1_540/Y 0.05fF
C37748 INPUT_2 POR2X1_5/a_16_28# 0.02fF
C37749 POR2X1_713/B PAND2X1_692/CTRL2 0.00fF
C37750 POR2X1_68/B POR2X1_4/Y 0.26fF
C37751 POR2X1_383/A POR2X1_339/Y 0.01fF
C37752 POR2X1_249/Y POR2X1_734/a_16_28# 0.01fF
C37753 PAND2X1_286/CTRL GATE_222 0.01fF
C37754 PAND2X1_349/A POR2X1_75/Y 0.01fF
C37755 POR2X1_305/CTRL2 POR2X1_305/Y 0.01fF
C37756 POR2X1_151/CTRL2 POR2X1_186/B 0.03fF
C37757 POR2X1_69/CTRL2 POR2X1_67/Y 0.01fF
C37758 POR2X1_826/Y PAND2X1_640/B 0.07fF
C37759 POR2X1_845/A POR2X1_845/O 0.03fF
C37760 POR2X1_54/Y POR2X1_848/A 0.37fF
C37761 POR2X1_62/Y POR2X1_623/A 0.01fF
C37762 POR2X1_57/A POR2X1_518/O 0.01fF
C37763 PAND2X1_530/CTRL PAND2X1_52/B 0.30fF
C37764 POR2X1_477/A PAND2X1_52/B 0.06fF
C37765 PAND2X1_631/CTRL2 POR2X1_416/B 0.01fF
C37766 POR2X1_565/CTRL2 PAND2X1_52/B 0.03fF
C37767 PAND2X1_665/CTRL2 PAND2X1_60/B 0.01fF
C37768 POR2X1_814/A POR2X1_94/A 0.00fF
C37769 POR2X1_110/Y PAND2X1_467/Y 0.07fF
C37770 POR2X1_67/Y POR2X1_750/B 0.03fF
C37771 POR2X1_78/B PAND2X1_628/a_16_344# 0.04fF
C37772 POR2X1_244/Y POR2X1_186/B 0.03fF
C37773 POR2X1_348/A POR2X1_814/A 0.02fF
C37774 POR2X1_68/A PAND2X1_681/O 0.03fF
C37775 POR2X1_61/CTRL POR2X1_447/B 0.08fF
C37776 POR2X1_180/B POR2X1_181/CTRL2 0.00fF
C37777 POR2X1_539/O POR2X1_567/A 0.01fF
C37778 POR2X1_864/A POR2X1_780/CTRL 0.00fF
C37779 PAND2X1_602/O POR2X1_600/Y 0.02fF
C37780 PAND2X1_747/CTRL PAND2X1_52/B 0.09fF
C37781 PAND2X1_631/A PAND2X1_348/A 0.90fF
C37782 POR2X1_707/B POR2X1_635/A 0.02fF
C37783 POR2X1_9/Y POR2X1_618/O 0.30fF
C37784 POR2X1_775/a_16_28# POR2X1_568/A 0.00fF
C37785 POR2X1_257/A POR2X1_72/B 1.08fF
C37786 POR2X1_479/B POR2X1_288/CTRL2 0.01fF
C37787 POR2X1_754/Y POR2X1_37/Y 0.17fF
C37788 POR2X1_760/A POR2X1_760/a_56_344# 0.00fF
C37789 POR2X1_329/A POR2X1_46/Y 0.03fF
C37790 POR2X1_520/B POR2X1_383/Y 0.02fF
C37791 POR2X1_379/O PAND2X1_52/B 0.32fF
C37792 POR2X1_329/Y PAND2X1_362/B 0.01fF
C37793 POR2X1_267/B POR2X1_341/A 0.05fF
C37794 PAND2X1_349/A PAND2X1_332/Y 0.03fF
C37795 POR2X1_828/Y PAND2X1_39/B 0.19fF
C37796 PAND2X1_86/a_16_344# PAND2X1_57/B 0.02fF
C37797 POR2X1_496/Y POR2X1_32/A 0.00fF
C37798 POR2X1_799/O PAND2X1_72/A 0.01fF
C37799 POR2X1_97/A POR2X1_241/B 0.03fF
C37800 POR2X1_646/Y POR2X1_590/A 0.14fF
C37801 PAND2X1_97/Y POR2X1_293/Y 0.05fF
C37802 POR2X1_442/O POR2X1_236/Y 0.01fF
C37803 POR2X1_266/a_56_344# PAND2X1_41/B 0.00fF
C37804 POR2X1_728/A POR2X1_156/Y 0.00fF
C37805 PAND2X1_404/Y PAND2X1_500/a_76_28# 0.01fF
C37806 PAND2X1_20/A POR2X1_33/CTRL2 0.01fF
C37807 POR2X1_150/Y POR2X1_79/Y 0.03fF
C37808 POR2X1_89/Y POR2X1_60/A 0.01fF
C37809 POR2X1_191/CTRL POR2X1_191/Y 0.01fF
C37810 POR2X1_283/O POR2X1_283/Y 0.01fF
C37811 PAND2X1_234/CTRL2 PAND2X1_88/Y 0.01fF
C37812 PAND2X1_317/CTRL2 POR2X1_167/Y 0.01fF
C37813 INPUT_3 POR2X1_88/Y 0.05fF
C37814 POR2X1_275/Y POR2X1_46/Y 0.32fF
C37815 POR2X1_162/CTRL POR2X1_161/Y 0.01fF
C37816 POR2X1_52/O POR2X1_7/Y 0.01fF
C37817 PAND2X1_844/CTRL PAND2X1_351/A 0.00fF
C37818 POR2X1_52/A POR2X1_484/Y 0.04fF
C37819 POR2X1_554/B POR2X1_276/O 0.01fF
C37820 PAND2X1_23/Y POR2X1_227/A 0.00fF
C37821 PAND2X1_341/B POR2X1_39/B 0.05fF
C37822 PAND2X1_48/A POR2X1_725/CTRL2 0.01fF
C37823 POR2X1_32/A PAND2X1_733/A 0.08fF
C37824 POR2X1_48/A PAND2X1_62/CTRL 0.02fF
C37825 PAND2X1_603/O POR2X1_750/B 0.01fF
C37826 POR2X1_715/A PAND2X1_72/A 0.02fF
C37827 POR2X1_180/CTRL2 POR2X1_181/Y 0.01fF
C37828 PAND2X1_436/a_16_344# PAND2X1_499/Y 0.02fF
C37829 POR2X1_66/B POR2X1_121/B 0.03fF
C37830 POR2X1_627/Y POR2X1_628/Y 0.00fF
C37831 POR2X1_490/O PAND2X1_215/B 0.18fF
C37832 PAND2X1_58/A PAND2X1_585/O 0.17fF
C37833 POR2X1_669/B POR2X1_423/Y 0.03fF
C37834 INPUT_2 PAND2X1_608/O 0.01fF
C37835 PAND2X1_622/CTRL2 POR2X1_669/B 0.51fF
C37836 POR2X1_43/B PAND2X1_447/O 0.01fF
C37837 PAND2X1_307/CTRL POR2X1_14/Y 0.01fF
C37838 POR2X1_736/A POR2X1_188/Y 0.05fF
C37839 POR2X1_119/Y PAND2X1_339/O 0.04fF
C37840 POR2X1_27/CTRL POR2X1_38/Y 0.04fF
C37841 PAND2X1_352/Y POR2X1_39/B 0.02fF
C37842 POR2X1_754/Y POR2X1_615/O 0.29fF
C37843 POR2X1_753/Y POR2X1_615/CTRL -0.02fF
C37844 PAND2X1_307/CTRL PAND2X1_453/A 0.01fF
C37845 POR2X1_188/A POR2X1_121/B 0.07fF
C37846 PAND2X1_6/Y POR2X1_554/B 0.01fF
C37847 POR2X1_66/B POR2X1_630/A 0.09fF
C37848 POR2X1_405/a_76_344# POR2X1_296/B 0.08fF
C37849 PAND2X1_622/a_76_28# POR2X1_48/A 0.01fF
C37850 PAND2X1_90/A POR2X1_54/Y 0.03fF
C37851 POR2X1_679/CTRL POR2X1_816/A 0.01fF
C37852 PAND2X1_48/B D_INPUT_5 0.34fF
C37853 POR2X1_337/Y PAND2X1_72/A 0.07fF
C37854 POR2X1_344/A PAND2X1_93/B 0.01fF
C37855 PAND2X1_464/B PAND2X1_785/a_16_344# 0.02fF
C37856 POR2X1_671/O POR2X1_37/Y 0.01fF
C37857 POR2X1_34/Y POR2X1_94/A 0.10fF
C37858 PAND2X1_225/O POR2X1_750/B 0.05fF
C37859 POR2X1_23/Y PAND2X1_735/Y 0.08fF
C37860 POR2X1_357/B POR2X1_212/B 0.09fF
C37861 PAND2X1_48/B PAND2X1_59/m4_208_n4# 0.07fF
C37862 POR2X1_614/A POR2X1_452/CTRL 0.01fF
C37863 POR2X1_296/O POR2X1_68/B 0.01fF
C37864 POR2X1_182/O POR2X1_180/Y 0.00fF
C37865 PAND2X1_212/CTRL POR2X1_55/Y 0.01fF
C37866 PAND2X1_41/B PAND2X1_531/a_76_28# 0.01fF
C37867 PAND2X1_58/A PAND2X1_589/CTRL 0.01fF
C37868 PAND2X1_659/CTRL2 POR2X1_498/Y 0.01fF
C37869 PAND2X1_793/Y POR2X1_437/a_16_28# 0.02fF
C37870 PAND2X1_6/Y POR2X1_803/CTRL2 0.00fF
C37871 POR2X1_294/O D_GATE_741 0.16fF
C37872 POR2X1_446/B POR2X1_659/O 0.01fF
C37873 PAND2X1_783/B PAND2X1_779/Y 0.02fF
C37874 POR2X1_477/A POR2X1_434/O 0.15fF
C37875 POR2X1_186/Y POR2X1_798/CTRL2 0.15fF
C37876 POR2X1_333/A PAND2X1_90/Y 1.76fF
C37877 POR2X1_49/Y POR2X1_72/B 0.20fF
C37878 PAND2X1_9/Y PAND2X1_69/A 0.20fF
C37879 POR2X1_651/CTRL2 POR2X1_66/A 0.01fF
C37880 POR2X1_20/B POR2X1_38/Y 0.17fF
C37881 PAND2X1_73/Y PAND2X1_760/CTRL2 0.01fF
C37882 PAND2X1_52/B PAND2X1_680/a_76_28# 0.02fF
C37883 POR2X1_274/A POR2X1_130/Y 0.03fF
C37884 PAND2X1_644/Y PAND2X1_758/O 0.00fF
C37885 PAND2X1_630/a_56_28# POR2X1_628/Y 0.00fF
C37886 PAND2X1_65/B POR2X1_254/CTRL2 0.00fF
C37887 POR2X1_71/Y POR2X1_37/Y 0.08fF
C37888 POR2X1_72/B PAND2X1_558/CTRL2 0.01fF
C37889 PAND2X1_771/Y PAND2X1_555/A 1.52fF
C37890 POR2X1_290/Y D_INPUT_0 0.05fF
C37891 POR2X1_244/B POR2X1_555/B 0.01fF
C37892 PAND2X1_831/Y POR2X1_271/B 0.22fF
C37893 POR2X1_138/a_16_28# POR2X1_260/B 0.02fF
C37894 POR2X1_475/A POR2X1_777/B 0.03fF
C37895 POR2X1_603/Y INPUT_0 6.66fF
C37896 PAND2X1_61/CTRL2 POR2X1_55/Y 0.12fF
C37897 POR2X1_20/B PAND2X1_785/a_56_28# 0.00fF
C37898 POR2X1_506/B VDD 0.45fF
C37899 POR2X1_94/CTRL POR2X1_23/Y 0.04fF
C37900 POR2X1_754/Y POR2X1_293/Y 0.00fF
C37901 PAND2X1_448/CTRL POR2X1_42/Y 0.03fF
C37902 POR2X1_37/Y POR2X1_42/Y 1.04fF
C37903 POR2X1_445/A PAND2X1_96/B 0.42fF
C37904 POR2X1_14/Y PAND2X1_734/B 0.02fF
C37905 POR2X1_855/B POR2X1_864/A 0.03fF
C37906 PAND2X1_90/Y POR2X1_734/A 0.09fF
C37907 POR2X1_850/B PAND2X1_57/B 0.05fF
C37908 PAND2X1_777/a_56_28# POR2X1_7/B 0.00fF
C37909 POR2X1_299/Y PAND2X1_302/O 0.00fF
C37910 POR2X1_244/B POR2X1_227/a_16_28# 0.01fF
C37911 PAND2X1_96/B POR2X1_643/Y 0.01fF
C37912 POR2X1_383/A POR2X1_541/B 0.05fF
C37913 POR2X1_106/Y PAND2X1_562/B 0.25fF
C37914 PAND2X1_793/Y POR2X1_516/Y 0.03fF
C37915 POR2X1_76/O POR2X1_724/A 0.01fF
C37916 POR2X1_376/B POR2X1_381/CTRL2 0.01fF
C37917 POR2X1_843/CTRL POR2X1_733/A 0.47fF
C37918 POR2X1_78/B POR2X1_259/A 0.05fF
C37919 POR2X1_376/B PAND2X1_803/A 0.04fF
C37920 POR2X1_640/Y VDD 0.29fF
C37921 POR2X1_812/a_16_28# POR2X1_121/B 0.09fF
C37922 PAND2X1_841/B POR2X1_516/Y 0.03fF
C37923 POR2X1_344/CTRL2 POR2X1_344/A 0.01fF
C37924 POR2X1_502/A POR2X1_640/CTRL 0.02fF
C37925 POR2X1_376/B POR2X1_677/a_16_28# 0.01fF
C37926 POR2X1_244/B POR2X1_330/Y 0.03fF
C37927 POR2X1_257/A PAND2X1_570/B 0.10fF
C37928 PAND2X1_48/B POR2X1_632/B 0.03fF
C37929 PAND2X1_48/B POR2X1_269/a_16_28# 0.02fF
C37930 POR2X1_241/B POR2X1_294/B 0.03fF
C37931 POR2X1_818/Y PAND2X1_69/A 0.03fF
C37932 POR2X1_334/Y POR2X1_814/A 0.02fF
C37933 POR2X1_334/A PAND2X1_86/CTRL 0.00fF
C37934 POR2X1_857/a_56_344# POR2X1_579/Y 0.00fF
C37935 POR2X1_293/O VDD -0.00fF
C37936 POR2X1_514/Y POR2X1_296/B 0.03fF
C37937 POR2X1_66/A PAND2X1_518/CTRL2 0.03fF
C37938 PAND2X1_579/B PAND2X1_579/O 0.01fF
C37939 POR2X1_692/CTRL2 POR2X1_526/Y 0.01fF
C37940 POR2X1_673/m4_208_n4# PAND2X1_8/Y 0.02fF
C37941 PAND2X1_714/CTRL2 POR2X1_40/Y 0.01fF
C37942 INPUT_1 POR2X1_20/B 0.19fF
C37943 POR2X1_251/A PAND2X1_553/B 0.18fF
C37944 POR2X1_274/A POR2X1_228/Y 0.03fF
C37945 POR2X1_28/a_16_28# D_INPUT_1 0.03fF
C37946 PAND2X1_499/Y POR2X1_497/Y 0.01fF
C37947 PAND2X1_787/A PAND2X1_776/Y 0.02fF
C37948 PAND2X1_272/CTRL POR2X1_112/Y 0.08fF
C37949 POR2X1_81/O POR2X1_43/B 0.02fF
C37950 PAND2X1_807/O PAND2X1_805/Y -0.00fF
C37951 POR2X1_251/Y PAND2X1_220/Y 0.16fF
C37952 POR2X1_114/B PAND2X1_279/CTRL2 0.00fF
C37953 PAND2X1_287/Y PAND2X1_578/CTRL2 -0.00fF
C37954 POR2X1_411/B PAND2X1_722/CTRL2 0.01fF
C37955 PAND2X1_539/B VDD 0.03fF
C37956 POR2X1_13/A POR2X1_106/Y 0.03fF
C37957 PAND2X1_201/O PAND2X1_358/A 0.05fF
C37958 PAND2X1_66/O POR2X1_283/A 0.06fF
C37959 PAND2X1_3/A INPUT_6 0.09fF
C37960 POR2X1_590/A POR2X1_804/A 0.05fF
C37961 PAND2X1_56/Y POR2X1_830/CTRL 0.01fF
C37962 POR2X1_651/O PAND2X1_41/B 0.02fF
C37963 POR2X1_66/B PAND2X1_56/Y 0.05fF
C37964 PAND2X1_724/B PAND2X1_731/B 0.13fF
C37965 POR2X1_66/B POR2X1_795/B 0.07fF
C37966 PAND2X1_20/A POR2X1_391/Y 0.07fF
C37967 POR2X1_221/CTRL POR2X1_220/Y 0.01fF
C37968 POR2X1_8/Y INPUT_3 0.93fF
C37969 PAND2X1_593/CTRL2 INPUT_0 0.01fF
C37970 POR2X1_66/A POR2X1_194/a_16_28# 0.03fF
C37971 POR2X1_417/Y PAND2X1_514/Y 0.08fF
C37972 POR2X1_20/B POR2X1_153/Y 0.17fF
C37973 POR2X1_43/B PAND2X1_195/CTRL 0.01fF
C37974 POR2X1_60/A POR2X1_56/Y 0.05fF
C37975 POR2X1_121/A POR2X1_654/CTRL2 0.01fF
C37976 POR2X1_52/A PAND2X1_803/A 0.02fF
C37977 PAND2X1_557/A PAND2X1_794/B 0.04fF
C37978 POR2X1_855/A POR2X1_855/Y 0.24fF
C37979 POR2X1_267/A PAND2X1_69/A 0.01fF
C37980 PAND2X1_63/Y POR2X1_641/CTRL 0.12fF
C37981 POR2X1_188/A PAND2X1_56/Y 0.05fF
C37982 PAND2X1_675/A PAND2X1_540/CTRL 0.02fF
C37983 POR2X1_48/A PAND2X1_348/CTRL2 0.11fF
C37984 POR2X1_855/B POR2X1_855/O 0.00fF
C37985 POR2X1_404/CTRL2 POR2X1_35/Y 0.01fF
C37986 PAND2X1_382/CTRL2 PAND2X1_381/Y 0.00fF
C37987 POR2X1_506/B PAND2X1_32/B 0.00fF
C37988 POR2X1_23/Y POR2X1_171/CTRL 0.01fF
C37989 POR2X1_41/B PAND2X1_833/O 0.09fF
C37990 PAND2X1_689/a_76_28# PAND2X1_32/B 0.02fF
C37991 POR2X1_670/O POR2X1_42/Y 0.01fF
C37992 PAND2X1_55/O PAND2X1_55/Y 0.02fF
C37993 POR2X1_23/Y PAND2X1_569/B 0.01fF
C37994 POR2X1_72/B PAND2X1_565/CTRL 0.01fF
C37995 POR2X1_777/B POR2X1_218/A 0.10fF
C37996 POR2X1_754/Y POR2X1_408/Y 0.10fF
C37997 POR2X1_267/CTRL2 POR2X1_318/A 0.02fF
C37998 POR2X1_66/A POR2X1_181/B 0.08fF
C37999 VDD POR2X1_121/Y 0.15fF
C38000 PAND2X1_96/B POR2X1_792/a_16_28# 0.02fF
C38001 POR2X1_96/A PAND2X1_579/B 0.03fF
C38002 POR2X1_150/Y PAND2X1_730/A 0.03fF
C38003 PAND2X1_803/A POR2X1_152/A 0.03fF
C38004 POR2X1_269/A POR2X1_228/Y 0.05fF
C38005 POR2X1_814/A POR2X1_343/CTRL 0.03fF
C38006 POR2X1_696/Y POR2X1_697/Y 0.00fF
C38007 PAND2X1_48/B PAND2X1_321/O 0.01fF
C38008 POR2X1_790/A POR2X1_391/A 0.03fF
C38009 PAND2X1_558/O PAND2X1_493/Y 0.06fF
C38010 PAND2X1_558/a_16_344# POR2X1_494/Y 0.03fF
C38011 POR2X1_808/A PAND2X1_69/A 0.09fF
C38012 PAND2X1_20/A PAND2X1_505/O 0.01fF
C38013 PAND2X1_206/a_16_344# POR2X1_293/Y 0.01fF
C38014 POR2X1_436/CTRL2 POR2X1_209/A 0.01fF
C38015 PAND2X1_803/Y POR2X1_60/A 0.03fF
C38016 POR2X1_51/A INPUT_5 2.47fF
C38017 POR2X1_43/B PAND2X1_76/Y 0.03fF
C38018 PAND2X1_90/A PAND2X1_80/O 0.01fF
C38019 PAND2X1_272/O POR2X1_553/A 0.02fF
C38020 POR2X1_502/A POR2X1_638/CTRL2 0.01fF
C38021 POR2X1_138/CTRL2 POR2X1_130/A 0.03fF
C38022 POR2X1_706/O POR2X1_383/A 0.02fF
C38023 POR2X1_278/Y PAND2X1_592/Y 0.07fF
C38024 PAND2X1_65/B POR2X1_218/A 0.91fF
C38025 POR2X1_713/A POR2X1_713/O 0.01fF
C38026 POR2X1_78/A POR2X1_590/CTRL 0.01fF
C38027 POR2X1_377/CTRL VDD 0.00fF
C38028 PAND2X1_41/B PAND2X1_518/O 0.17fF
C38029 PAND2X1_778/Y POR2X1_72/B 0.63fF
C38030 PAND2X1_211/A POR2X1_73/Y 0.01fF
C38031 PAND2X1_7/CTRL2 POR2X1_244/B 0.01fF
C38032 POR2X1_693/Y POR2X1_236/Y 0.03fF
C38033 POR2X1_260/B POR2X1_3/B 0.63fF
C38034 PAND2X1_734/B POR2X1_55/Y 0.63fF
C38035 POR2X1_208/A POR2X1_201/CTRL 0.00fF
C38036 PAND2X1_725/Y PAND2X1_731/A 0.00fF
C38037 POR2X1_66/B POR2X1_383/A 0.84fF
C38038 PAND2X1_553/CTRL2 POR2X1_106/Y 0.01fF
C38039 POR2X1_56/B PAND2X1_453/CTRL2 0.02fF
C38040 POR2X1_71/Y POR2X1_293/Y 0.02fF
C38041 POR2X1_497/Y POR2X1_521/O 0.01fF
C38042 VDD POR2X1_723/B 0.01fF
C38043 POR2X1_407/A POR2X1_130/A 0.06fF
C38044 POR2X1_548/CTRL POR2X1_68/B 0.10fF
C38045 PAND2X1_462/B POR2X1_232/CTRL 0.06fF
C38046 PAND2X1_90/Y POR2X1_788/B 0.36fF
C38047 PAND2X1_388/CTRL2 POR2X1_236/Y 0.01fF
C38048 POR2X1_356/A POR2X1_466/O 0.06fF
C38049 POR2X1_188/A POR2X1_383/A 0.10fF
C38050 PAND2X1_829/O POR2X1_260/A 0.04fF
C38051 POR2X1_293/Y POR2X1_42/Y 0.13fF
C38052 PAND2X1_96/B PAND2X1_58/CTRL 0.01fF
C38053 PAND2X1_58/A POR2X1_260/A 0.05fF
C38054 POR2X1_55/Y PAND2X1_506/CTRL2 0.01fF
C38055 PAND2X1_40/O PAND2X1_587/Y 0.01fF
C38056 POR2X1_41/B PAND2X1_35/O -0.00fF
C38057 PAND2X1_556/B POR2X1_90/Y 0.03fF
C38058 PAND2X1_91/a_76_28# POR2X1_192/B 0.02fF
C38059 POR2X1_403/A PAND2X1_69/A 0.06fF
C38060 PAND2X1_820/O PAND2X1_820/B 0.00fF
C38061 PAND2X1_48/B PAND2X1_516/m4_208_n4# 0.12fF
C38062 POR2X1_62/Y POR2X1_66/A 0.07fF
C38063 POR2X1_78/B PAND2X1_88/Y 0.08fF
C38064 POR2X1_67/A POR2X1_129/Y 0.04fF
C38065 POR2X1_508/A POR2X1_567/B 0.03fF
C38066 POR2X1_78/B POR2X1_84/Y 0.03fF
C38067 PAND2X1_258/a_76_28# POR2X1_186/B 0.00fF
C38068 POR2X1_134/Y PAND2X1_768/CTRL2 0.01fF
C38069 PAND2X1_855/a_76_28# POR2X1_236/Y 0.00fF
C38070 POR2X1_528/O POR2X1_56/B 0.01fF
C38071 POR2X1_288/CTRL2 PAND2X1_48/A 0.04fF
C38072 PAND2X1_182/A PAND2X1_182/CTRL 0.02fF
C38073 POR2X1_293/Y POR2X1_309/Y 0.01fF
C38074 POR2X1_32/A POR2X1_75/Y 0.01fF
C38075 POR2X1_709/CTRL2 PAND2X1_90/Y 0.06fF
C38076 POR2X1_96/A POR2X1_73/Y 0.10fF
C38077 POR2X1_836/CTRL POR2X1_191/Y -0.01fF
C38078 POR2X1_387/Y POR2X1_372/O 0.06fF
C38079 POR2X1_525/Y PAND2X1_546/O 0.02fF
C38080 POR2X1_466/A POR2X1_552/m4_208_n4# 0.06fF
C38081 PAND2X1_6/Y PAND2X1_369/CTRL 0.01fF
C38082 POR2X1_562/CTRL2 POR2X1_562/B 0.01fF
C38083 PAND2X1_338/B VDD 0.28fF
C38084 POR2X1_546/B POR2X1_844/B 0.11fF
C38085 PAND2X1_58/A PAND2X1_142/O 0.03fF
C38086 POR2X1_730/B POR2X1_730/CTRL2 0.01fF
C38087 PAND2X1_245/O PAND2X1_48/A 0.02fF
C38088 INPUT_4 POR2X1_386/O 0.01fF
C38089 POR2X1_57/A POR2X1_693/CTRL 0.01fF
C38090 POR2X1_52/A POR2X1_583/CTRL2 0.01fF
C38091 POR2X1_53/m4_208_n4# POR2X1_699/m4_208_n4# 0.13fF
C38092 POR2X1_57/A POR2X1_46/Y 0.08fF
C38093 PAND2X1_69/A POR2X1_149/Y 0.03fF
C38094 PAND2X1_461/O POR2X1_612/Y 0.12fF
C38095 PAND2X1_206/A PAND2X1_358/a_76_28# 0.01fF
C38096 POR2X1_579/Y POR2X1_570/B 0.03fF
C38097 POR2X1_220/Y POR2X1_318/A 0.07fF
C38098 POR2X1_278/m4_208_n4# PAND2X1_734/m4_208_n4# 0.13fF
C38099 POR2X1_547/CTRL2 POR2X1_614/A 0.03fF
C38100 POR2X1_511/Y PAND2X1_550/B 0.03fF
C38101 POR2X1_416/B PAND2X1_222/A 0.03fF
C38102 POR2X1_316/Y POR2X1_23/Y 0.12fF
C38103 POR2X1_124/CTRL POR2X1_137/Y 0.00fF
C38104 PAND2X1_6/Y POR2X1_800/A 0.02fF
C38105 POR2X1_141/Y POR2X1_574/Y 0.01fF
C38106 POR2X1_278/Y PAND2X1_348/Y 0.12fF
C38107 POR2X1_722/A POR2X1_602/B 0.04fF
C38108 PAND2X1_737/B POR2X1_5/Y 0.10fF
C38109 POR2X1_489/a_56_344# POR2X1_260/A 0.00fF
C38110 POR2X1_405/Y PAND2X1_60/B 0.03fF
C38111 POR2X1_567/B POR2X1_568/B 0.01fF
C38112 POR2X1_192/Y POR2X1_727/CTRL2 0.10fF
C38113 POR2X1_13/A PAND2X1_349/A 0.03fF
C38114 POR2X1_567/A POR2X1_241/B 0.03fF
C38115 POR2X1_404/Y POR2X1_318/A 0.07fF
C38116 PAND2X1_425/CTRL2 PAND2X1_18/B 0.03fF
C38117 POR2X1_455/O POR2X1_456/B 0.18fF
C38118 PAND2X1_94/A POR2X1_410/CTRL 0.05fF
C38119 PAND2X1_440/CTRL2 POR2X1_23/Y 0.03fF
C38120 POR2X1_784/A PAND2X1_60/B 0.02fF
C38121 POR2X1_145/CTRL PAND2X1_213/Y 0.00fF
C38122 PAND2X1_252/a_76_28# PAND2X1_55/Y 0.02fF
C38123 PAND2X1_661/Y PAND2X1_688/m4_208_n4# 0.09fF
C38124 PAND2X1_297/CTRL2 PAND2X1_57/B 0.01fF
C38125 POR2X1_89/CTRL PAND2X1_333/Y 0.01fF
C38126 POR2X1_567/B PAND2X1_167/m4_208_n4# 0.06fF
C38127 POR2X1_447/a_16_28# POR2X1_294/B 0.02fF
C38128 POR2X1_537/Y POR2X1_330/Y 0.05fF
C38129 POR2X1_96/A PAND2X1_244/B 0.03fF
C38130 PAND2X1_6/Y POR2X1_702/A 0.03fF
C38131 POR2X1_30/CTRL2 POR2X1_3/A 0.32fF
C38132 PAND2X1_197/CTRL PAND2X1_656/A 0.01fF
C38133 POR2X1_57/A PAND2X1_334/O 0.01fF
C38134 POR2X1_85/CTRL2 POR2X1_83/B 0.02fF
C38135 PAND2X1_632/B POR2X1_625/Y 0.03fF
C38136 POR2X1_408/Y POR2X1_42/Y 0.10fF
C38137 POR2X1_254/Y POR2X1_456/B 0.32fF
C38138 POR2X1_614/A POR2X1_570/B 0.05fF
C38139 POR2X1_732/B PAND2X1_60/B 0.42fF
C38140 PAND2X1_341/Y VDD 0.15fF
C38141 POR2X1_65/A POR2X1_110/CTRL 0.04fF
C38142 PAND2X1_65/B POR2X1_557/B 0.03fF
C38143 PAND2X1_413/CTRL2 VDD 0.00fF
C38144 PAND2X1_63/Y PAND2X1_96/B 1.23fF
C38145 POR2X1_139/A PAND2X1_32/B 0.06fF
C38146 POR2X1_68/B D_INPUT_1 0.33fF
C38147 PAND2X1_857/a_76_28# POR2X1_83/B 0.02fF
C38148 PAND2X1_808/Y PAND2X1_363/CTRL2 0.01fF
C38149 PAND2X1_658/A POR2X1_7/A 0.07fF
C38150 POR2X1_558/B PAND2X1_72/A 0.04fF
C38151 PAND2X1_732/CTRL POR2X1_39/B 0.01fF
C38152 PAND2X1_117/CTRL2 POR2X1_260/A 0.03fF
C38153 PAND2X1_636/O POR2X1_583/Y 0.02fF
C38154 POR2X1_834/Y POR2X1_513/B 0.01fF
C38155 POR2X1_72/B PAND2X1_330/O 0.09fF
C38156 POR2X1_691/CTRL POR2X1_855/B 0.01fF
C38157 POR2X1_327/m4_208_n4# POR2X1_216/m4_208_n4# 0.18fF
C38158 PAND2X1_392/m4_208_n4# POR2X1_39/B 0.05fF
C38159 PAND2X1_383/CTRL POR2X1_816/A 0.01fF
C38160 POR2X1_111/Y POR2X1_46/Y 0.26fF
C38161 PAND2X1_79/O POR2X1_569/A 0.05fF
C38162 POR2X1_694/a_16_28# POR2X1_425/Y 0.11fF
C38163 POR2X1_63/O PAND2X1_63/B 0.02fF
C38164 PAND2X1_731/m4_208_n4# PAND2X1_147/m4_208_n4# 0.13fF
C38165 POR2X1_865/B POR2X1_114/m4_208_n4# 0.15fF
C38166 POR2X1_68/A POR2X1_725/Y 0.10fF
C38167 POR2X1_315/Y POR2X1_43/B 0.01fF
C38168 POR2X1_55/Y POR2X1_789/B 0.14fF
C38169 POR2X1_538/CTRL2 POR2X1_703/A 0.02fF
C38170 PAND2X1_725/O VDD 0.00fF
C38171 PAND2X1_693/CTRL PAND2X1_94/A 0.01fF
C38172 PAND2X1_693/CTRL2 INPUT_1 0.01fF
C38173 POR2X1_575/B POR2X1_456/B 0.01fF
C38174 POR2X1_665/A PAND2X1_645/B 0.16fF
C38175 POR2X1_239/O POR2X1_239/Y 0.01fF
C38176 POR2X1_147/CTRL2 POR2X1_78/A 0.04fF
C38177 VDD PAND2X1_3/B 0.82fF
C38178 PAND2X1_551/Y PAND2X1_569/B 0.03fF
C38179 POR2X1_809/A POR2X1_676/Y 0.01fF
C38180 POR2X1_174/B PAND2X1_109/a_76_28# 0.06fF
C38181 PAND2X1_73/Y POR2X1_715/CTRL 0.01fF
C38182 POR2X1_75/a_56_344# PAND2X1_349/A 0.00fF
C38183 POR2X1_110/Y PAND2X1_471/CTRL2 0.02fF
C38184 PAND2X1_533/CTRL POR2X1_532/Y 0.01fF
C38185 POR2X1_7/A POR2X1_73/Y 0.10fF
C38186 PAND2X1_659/Y PAND2X1_741/CTRL 0.03fF
C38187 POR2X1_49/Y POR2X1_52/O 0.02fF
C38188 POR2X1_114/O POR2X1_101/Y 0.15fF
C38189 PAND2X1_850/Y PAND2X1_276/CTRL2 0.05fF
C38190 POR2X1_32/A PAND2X1_332/Y 0.22fF
C38191 POR2X1_188/A PAND2X1_108/CTRL2 0.01fF
C38192 POR2X1_548/a_16_28# POR2X1_620/B 0.02fF
C38193 POR2X1_110/Y PAND2X1_549/CTRL 0.01fF
C38194 PAND2X1_723/O PAND2X1_723/A 0.02fF
C38195 POR2X1_502/A POR2X1_722/O 0.02fF
C38196 POR2X1_596/A PAND2X1_765/CTRL2 0.01fF
C38197 POR2X1_687/A PAND2X1_69/A 0.03fF
C38198 PAND2X1_707/Y POR2X1_394/A 0.36fF
C38199 POR2X1_367/a_16_28# POR2X1_191/Y 0.03fF
C38200 POR2X1_334/Y POR2X1_260/Y 0.02fF
C38201 PAND2X1_48/B POR2X1_359/B -0.00fF
C38202 D_GATE_222 POR2X1_507/A 0.02fF
C38203 POR2X1_684/Y POR2X1_13/A 0.01fF
C38204 POR2X1_614/A PAND2X1_813/CTRL 0.01fF
C38205 POR2X1_493/B PAND2X1_63/Y 0.01fF
C38206 POR2X1_245/Y POR2X1_387/Y 0.08fF
C38207 POR2X1_278/Y PAND2X1_476/A 0.05fF
C38208 PAND2X1_798/B POR2X1_394/A 0.05fF
C38209 POR2X1_95/CTRL POR2X1_51/A 0.01fF
C38210 PAND2X1_74/a_16_344# PAND2X1_72/A 0.02fF
C38211 PAND2X1_696/CTRL2 POR2X1_502/A 0.02fF
C38212 PAND2X1_96/B POR2X1_260/A 0.20fF
C38213 POR2X1_7/B POR2X1_7/Y 0.05fF
C38214 POR2X1_78/B POR2X1_568/B 0.10fF
C38215 PAND2X1_850/Y PAND2X1_785/Y 0.15fF
C38216 POR2X1_92/CTRL2 POR2X1_8/Y 0.00fF
C38217 POR2X1_416/B POR2X1_743/O 0.03fF
C38218 PAND2X1_244/B POR2X1_7/A 0.03fF
C38219 PAND2X1_793/Y PAND2X1_860/CTRL 0.01fF
C38220 POR2X1_184/Y POR2X1_75/Y 0.00fF
C38221 PAND2X1_90/A POR2X1_4/Y 0.39fF
C38222 POR2X1_464/O POR2X1_736/A 0.04fF
C38223 PAND2X1_833/O POR2X1_77/Y 0.04fF
C38224 D_INPUT_3 POR2X1_96/O 0.15fF
C38225 POR2X1_463/Y POR2X1_711/a_16_28# 0.01fF
C38226 POR2X1_681/O POR2X1_681/Y 0.01fF
C38227 PAND2X1_675/A POR2X1_385/Y 0.03fF
C38228 PAND2X1_150/CTRL2 POR2X1_186/B 0.01fF
C38229 POR2X1_790/A POR2X1_294/A 0.03fF
C38230 PAND2X1_73/Y POR2X1_643/O 0.04fF
C38231 PAND2X1_779/CTRL POR2X1_90/Y 0.02fF
C38232 PAND2X1_714/A POR2X1_167/Y 0.17fF
C38233 PAND2X1_865/Y PAND2X1_652/A 0.00fF
C38234 POR2X1_257/A PAND2X1_247/CTRL 0.05fF
C38235 INPUT_1 PAND2X1_528/CTRL 0.00fF
C38236 PAND2X1_3/B PAND2X1_32/B 0.03fF
C38237 PAND2X1_787/A PAND2X1_853/B 0.00fF
C38238 POR2X1_518/CTRL POR2X1_519/Y 0.01fF
C38239 POR2X1_518/CTRL2 POR2X1_518/Y 0.02fF
C38240 POR2X1_779/CTRL POR2X1_513/B 0.01fF
C38241 PAND2X1_630/CTRL2 PAND2X1_508/B 0.01fF
C38242 POR2X1_406/Y PAND2X1_339/m4_208_n4# 0.01fF
C38243 POR2X1_49/Y PAND2X1_147/CTRL 0.01fF
C38244 POR2X1_68/B POR2X1_620/B 1.46fF
C38245 POR2X1_692/CTRL2 POR2X1_485/Y 0.00fF
C38246 POR2X1_676/Y POR2X1_728/A 0.00fF
C38247 INPUT_1 PAND2X1_632/CTRL 0.12fF
C38248 PAND2X1_704/m4_208_n4# POR2X1_142/Y 0.09fF
C38249 POR2X1_294/A PAND2X1_88/Y 0.03fF
C38250 POR2X1_42/O POR2X1_4/Y 0.06fF
C38251 POR2X1_493/B POR2X1_260/A 0.05fF
C38252 POR2X1_56/B POR2X1_416/B 0.02fF
C38253 POR2X1_332/B PAND2X1_72/A 0.06fF
C38254 POR2X1_190/Y PAND2X1_52/B 0.05fF
C38255 PAND2X1_501/CTRL2 PAND2X1_575/A 0.01fF
C38256 PAND2X1_557/A POR2X1_250/a_16_28# 0.03fF
C38257 PAND2X1_691/Y POR2X1_394/A 0.07fF
C38258 POR2X1_83/B POR2X1_431/CTRL 0.01fF
C38259 PAND2X1_319/B PAND2X1_353/Y 0.03fF
C38260 PAND2X1_845/CTRL2 POR2X1_39/B 0.18fF
C38261 PAND2X1_254/a_76_28# POR2X1_77/Y 0.02fF
C38262 PAND2X1_699/a_16_344# POR2X1_496/Y 0.05fF
C38263 POR2X1_703/A POR2X1_186/B 0.03fF
C38264 PAND2X1_35/O POR2X1_77/Y 0.08fF
C38265 PAND2X1_462/CTRL POR2X1_416/Y 0.01fF
C38266 POR2X1_65/A POR2X1_292/CTRL 0.03fF
C38267 POR2X1_856/B POR2X1_776/A 0.01fF
C38268 POR2X1_54/Y POR2X1_23/Y 0.03fF
C38269 POR2X1_60/A PAND2X1_97/Y 0.01fF
C38270 POR2X1_632/Y POR2X1_702/A 0.03fF
C38271 PAND2X1_63/Y POR2X1_342/B 0.01fF
C38272 POR2X1_800/A PAND2X1_52/B 0.02fF
C38273 POR2X1_191/B POR2X1_353/A 0.03fF
C38274 PAND2X1_217/B PAND2X1_717/A 0.07fF
C38275 PAND2X1_865/Y POR2X1_437/CTRL2 0.00fF
C38276 POR2X1_411/B PAND2X1_577/Y 4.29fF
C38277 PAND2X1_218/B PAND2X1_267/Y 0.01fF
C38278 PAND2X1_774/a_76_28# PAND2X1_771/Y 0.02fF
C38279 POR2X1_633/A POR2X1_633/O 0.09fF
C38280 POR2X1_67/Y POR2X1_720/A 0.03fF
C38281 POR2X1_814/A POR2X1_475/A 0.03fF
C38282 POR2X1_184/Y PAND2X1_332/Y 0.03fF
C38283 PAND2X1_243/B POR2X1_825/Y 0.03fF
C38284 POR2X1_326/A POR2X1_326/a_16_28# 0.03fF
C38285 POR2X1_456/B POR2X1_564/a_16_28# 0.03fF
C38286 POR2X1_454/O POR2X1_454/B 0.01fF
C38287 POR2X1_609/Y POR2X1_612/Y 0.07fF
C38288 PAND2X1_69/A POR2X1_568/A 0.03fF
C38289 PAND2X1_761/CTRL2 POR2X1_750/B 0.01fF
C38290 PAND2X1_3/A PAND2X1_36/CTRL2 0.01fF
C38291 PAND2X1_717/A VDD 0.80fF
C38292 POR2X1_326/a_16_28# POR2X1_324/Y 0.04fF
C38293 PAND2X1_832/CTRL2 POR2X1_411/B 0.01fF
C38294 POR2X1_738/A POR2X1_711/Y 0.04fF
C38295 PAND2X1_69/A PAND2X1_146/CTRL2 0.00fF
C38296 PAND2X1_41/CTRL2 PAND2X1_41/B 0.03fF
C38297 POR2X1_39/B POR2X1_310/Y 0.03fF
C38298 PAND2X1_240/O POR2X1_411/B 0.02fF
C38299 POR2X1_287/B POR2X1_556/A 0.01fF
C38300 PAND2X1_341/B POR2X1_62/Y 3.27fF
C38301 POR2X1_559/A PAND2X1_517/O 0.01fF
C38302 PAND2X1_497/a_16_344# POR2X1_78/A 0.02fF
C38303 POR2X1_646/Y POR2X1_66/A 0.03fF
C38304 POR2X1_48/A PAND2X1_732/CTRL 0.01fF
C38305 POR2X1_20/B PAND2X1_721/a_16_344# 0.01fF
C38306 POR2X1_67/A POR2X1_37/Y 0.01fF
C38307 PAND2X1_635/Y POR2X1_587/Y 0.04fF
C38308 PAND2X1_659/A PAND2X1_203/a_76_28# 0.05fF
C38309 POR2X1_483/A POR2X1_556/A 0.03fF
C38310 POR2X1_119/Y PAND2X1_858/a_56_28# 0.00fF
C38311 PAND2X1_404/Y POR2X1_40/Y 0.03fF
C38312 PAND2X1_58/A PAND2X1_28/m4_208_n4# 0.15fF
C38313 POR2X1_566/A POR2X1_465/O 0.36fF
C38314 POR2X1_202/A POR2X1_402/CTRL2 0.02fF
C38315 PAND2X1_412/CTRL POR2X1_260/B 0.01fF
C38316 PAND2X1_671/Y POR2X1_54/Y 0.04fF
C38317 POR2X1_362/A PAND2X1_72/A 0.01fF
C38318 PAND2X1_601/O POR2X1_718/A 0.01fF
C38319 POR2X1_776/A POR2X1_776/a_16_28# -0.00fF
C38320 POR2X1_129/Y PAND2X1_840/Y 0.23fF
C38321 POR2X1_674/Y POR2X1_32/A 0.14fF
C38322 PAND2X1_783/B VDD 0.04fF
C38323 POR2X1_805/CTRL2 POR2X1_805/B 0.01fF
C38324 POR2X1_326/CTRL POR2X1_568/A 0.03fF
C38325 POR2X1_814/A POR2X1_218/A 0.15fF
C38326 POR2X1_661/A POR2X1_513/O 0.04fF
C38327 PAND2X1_722/O PAND2X1_718/Y 0.06fF
C38328 POR2X1_322/CTRL2 POR2X1_441/Y 0.01fF
C38329 PAND2X1_230/O POR2X1_78/A 0.04fF
C38330 POR2X1_260/B POR2X1_285/CTRL 0.01fF
C38331 POR2X1_559/O POR2X1_814/A 0.01fF
C38332 PAND2X1_865/Y POR2X1_184/CTRL 0.00fF
C38333 POR2X1_590/A POR2X1_794/B 0.03fF
C38334 POR2X1_29/Y PAND2X1_87/a_16_344# 0.01fF
C38335 POR2X1_437/O PAND2X1_580/B 0.00fF
C38336 POR2X1_309/O POR2X1_40/Y 0.05fF
C38337 POR2X1_49/Y PAND2X1_796/CTRL -0.03fF
C38338 POR2X1_257/A POR2X1_7/B 0.03fF
C38339 PAND2X1_468/O POR2X1_679/A 0.05fF
C38340 POR2X1_634/A PAND2X1_428/CTRL 0.07fF
C38341 POR2X1_360/A POR2X1_243/B 0.03fF
C38342 POR2X1_360/A POR2X1_99/Y 0.02fF
C38343 POR2X1_23/Y PAND2X1_501/B 0.11fF
C38344 POR2X1_399/A POR2X1_411/B 0.01fF
C38345 PAND2X1_447/CTRL2 POR2X1_90/Y 0.01fF
C38346 POR2X1_591/A PAND2X1_719/Y 0.02fF
C38347 POR2X1_856/O PAND2X1_73/Y 0.01fF
C38348 POR2X1_692/O VDD -0.00fF
C38349 POR2X1_786/A POR2X1_266/CTRL 0.01fF
C38350 PAND2X1_485/CTRL2 PAND2X1_57/B 0.01fF
C38351 POR2X1_43/B POR2X1_442/CTRL2 0.03fF
C38352 INPUT_3 POR2X1_619/O 0.01fF
C38353 POR2X1_705/B POR2X1_705/O 0.00fF
C38354 PAND2X1_249/O PAND2X1_733/A 0.01fF
C38355 POR2X1_829/A PAND2X1_207/CTRL 0.00fF
C38356 POR2X1_308/CTRL POR2X1_660/Y 0.01fF
C38357 PAND2X1_58/A POR2X1_718/A 0.01fF
C38358 POR2X1_441/Y POR2X1_90/Y 0.03fF
C38359 PAND2X1_258/O POR2X1_244/B 0.02fF
C38360 POR2X1_137/B POR2X1_68/B 0.03fF
C38361 POR2X1_666/a_16_28# POR2X1_666/A 0.03fF
C38362 POR2X1_865/B POR2X1_116/A 0.03fF
C38363 POR2X1_198/CTRL2 PAND2X1_93/B 0.00fF
C38364 PAND2X1_108/O POR2X1_590/A 0.01fF
C38365 POR2X1_441/Y POR2X1_438/a_76_344# 0.00fF
C38366 PAND2X1_794/a_16_344# PAND2X1_473/B 0.01fF
C38367 POR2X1_814/B POR2X1_439/O 0.06fF
C38368 PAND2X1_806/CTRL POR2X1_42/Y 0.01fF
C38369 POR2X1_13/A POR2X1_32/A 1.75fF
C38370 POR2X1_260/B POR2X1_790/B 0.08fF
C38371 INPUT_3 POR2X1_68/B 0.91fF
C38372 PAND2X1_614/CTRL2 POR2X1_5/Y 0.00fF
C38373 POR2X1_836/A VDD 0.00fF
C38374 POR2X1_674/CTRL PAND2X1_742/B 0.01fF
C38375 POR2X1_717/a_76_344# POR2X1_499/A 0.01fF
C38376 POR2X1_16/A PAND2X1_608/O 0.01fF
C38377 POR2X1_130/A POR2X1_641/O 0.02fF
C38378 PAND2X1_96/B POR2X1_473/O 0.02fF
C38379 POR2X1_120/a_16_28# POR2X1_78/A 0.01fF
C38380 PAND2X1_9/Y PAND2X1_338/B 0.03fF
C38381 POR2X1_593/B PAND2X1_589/O 0.02fF
C38382 POR2X1_201/O VDD 0.00fF
C38383 POR2X1_66/B INPUT_0 0.24fF
C38384 POR2X1_624/Y POR2X1_140/O 0.02fF
C38385 POR2X1_268/Y POR2X1_236/Y 0.01fF
C38386 POR2X1_260/B PAND2X1_743/CTRL 0.01fF
C38387 POR2X1_78/B POR2X1_500/A 0.03fF
C38388 POR2X1_423/Y PAND2X1_499/Y 3.82fF
C38389 POR2X1_67/A POR2X1_293/Y 0.02fF
C38390 POR2X1_462/B POR2X1_848/A 0.00fF
C38391 PAND2X1_48/B POR2X1_555/B 0.03fF
C38392 POR2X1_813/CTRL PAND2X1_63/B 0.01fF
C38393 POR2X1_51/B POR2X1_20/B 0.03fF
C38394 PAND2X1_668/O POR2X1_60/A 0.04fF
C38395 PAND2X1_93/B PAND2X1_72/O 0.07fF
C38396 POR2X1_16/A POR2X1_679/CTRL2 0.21fF
C38397 PAND2X1_815/a_16_344# POR2X1_752/Y 0.02fF
C38398 PAND2X1_23/Y POR2X1_202/B 0.24fF
C38399 POR2X1_13/A POR2X1_417/Y 0.60fF
C38400 PAND2X1_319/B POR2X1_298/CTRL2 0.01fF
C38401 POR2X1_71/Y POR2X1_60/A 0.01fF
C38402 POR2X1_865/B POR2X1_862/Y 0.00fF
C38403 PAND2X1_860/A PAND2X1_860/O 0.01fF
C38404 POR2X1_814/A POR2X1_557/B 0.08fF
C38405 POR2X1_37/Y PAND2X1_642/B 0.05fF
C38406 POR2X1_478/O POR2X1_478/B 0.00fF
C38407 PAND2X1_217/O PAND2X1_723/A 0.00fF
C38408 POR2X1_685/A POR2X1_676/CTRL2 0.01fF
C38409 POR2X1_66/A POR2X1_804/A 0.05fF
C38410 POR2X1_60/CTRL2 D_INPUT_0 0.05fF
C38411 POR2X1_828/Y VDD 0.01fF
C38412 POR2X1_495/Y POR2X1_83/B 0.01fF
C38413 POR2X1_63/O POR2X1_32/A 0.01fF
C38414 PAND2X1_391/CTRL POR2X1_816/A 0.01fF
C38415 PAND2X1_58/A PAND2X1_110/O 0.02fF
C38416 POR2X1_224/CTRL POR2X1_226/Y 0.00fF
C38417 PAND2X1_65/B POR2X1_770/A 0.01fF
C38418 POR2X1_60/A POR2X1_42/Y 0.10fF
C38419 POR2X1_441/Y PAND2X1_732/A 0.13fF
C38420 PAND2X1_490/O POR2X1_66/A 0.02fF
C38421 PAND2X1_476/a_76_28# INPUT_0 0.01fF
C38422 POR2X1_616/O POR2X1_93/A 0.18fF
C38423 PAND2X1_699/O POR2X1_129/Y 0.06fF
C38424 POR2X1_198/B POR2X1_201/CTRL 0.01fF
C38425 PAND2X1_423/O PAND2X1_57/B 0.02fF
C38426 POR2X1_718/A POR2X1_435/Y 0.09fF
C38427 POR2X1_14/CTRL POR2X1_68/B 0.00fF
C38428 POR2X1_718/O POR2X1_435/Y 0.01fF
C38429 PAND2X1_755/CTRL2 PAND2X1_90/Y 0.01fF
C38430 POR2X1_390/B PAND2X1_39/B 0.02fF
C38431 PAND2X1_48/B POR2X1_330/Y 11.65fF
C38432 POR2X1_333/A D_GATE_222 0.10fF
C38433 PAND2X1_236/CTRL2 PAND2X1_8/Y 0.02fF
C38434 PAND2X1_484/CTRL POR2X1_705/B 0.00fF
C38435 POR2X1_707/A PAND2X1_95/B 0.00fF
C38436 POR2X1_12/CTRL INPUT_4 0.08fF
C38437 PAND2X1_404/A POR2X1_236/Y 0.01fF
C38438 POR2X1_49/Y POR2X1_7/B 0.14fF
C38439 POR2X1_57/A PAND2X1_352/A 0.01fF
C38440 POR2X1_60/A POR2X1_309/Y 0.05fF
C38441 PAND2X1_94/O PAND2X1_60/B 0.03fF
C38442 PAND2X1_20/A POR2X1_139/CTRL2 0.01fF
C38443 PAND2X1_857/CTRL POR2X1_329/A 0.03fF
C38444 INPUT_1 POR2X1_624/Y 0.01fF
C38445 PAND2X1_836/CTRL POR2X1_102/Y 0.01fF
C38446 PAND2X1_643/Y POR2X1_32/A 0.03fF
C38447 PAND2X1_119/CTRL POR2X1_78/A 0.11fF
C38448 POR2X1_629/A POR2X1_852/B 0.06fF
C38449 POR2X1_750/B POR2X1_732/B 0.03fF
C38450 PAND2X1_564/CTRL VDD 0.00fF
C38451 POR2X1_466/A PAND2X1_60/B 0.05fF
C38452 PAND2X1_741/a_16_344# PAND2X1_741/B 0.01fF
C38453 POR2X1_502/A PAND2X1_589/a_56_28# 0.00fF
C38454 PAND2X1_124/Y PAND2X1_723/A 0.02fF
C38455 POR2X1_78/A POR2X1_68/B 0.10fF
C38456 POR2X1_296/B PAND2X1_505/CTRL 0.01fF
C38457 POR2X1_302/A PAND2X1_299/CTRL 0.01fF
C38458 POR2X1_57/A PAND2X1_296/CTRL2 0.03fF
C38459 PAND2X1_640/B PAND2X1_559/CTRL 0.02fF
C38460 PAND2X1_57/B PAND2X1_57/O 0.04fF
C38461 POR2X1_43/B POR2X1_24/O 0.05fF
C38462 POR2X1_859/A INPUT_0 0.22fF
C38463 POR2X1_722/A PAND2X1_39/B 0.52fF
C38464 PAND2X1_84/Y POR2X1_46/Y 0.05fF
C38465 POR2X1_548/CTRL PAND2X1_90/A 0.01fF
C38466 POR2X1_94/A POR2X1_790/A 0.02fF
C38467 PAND2X1_220/O PAND2X1_220/Y 0.01fF
C38468 POR2X1_254/Y PAND2X1_57/B 0.07fF
C38469 POR2X1_812/B POR2X1_121/B 0.02fF
C38470 POR2X1_41/B VDD 7.15fF
C38471 POR2X1_692/CTRL2 PAND2X1_726/B 0.03fF
C38472 PAND2X1_862/B PAND2X1_573/O 0.01fF
C38473 POR2X1_40/Y PAND2X1_565/A 0.00fF
C38474 PAND2X1_65/B POR2X1_740/Y 0.05fF
C38475 POR2X1_202/A POR2X1_507/A 1.03fF
C38476 PAND2X1_55/Y POR2X1_285/CTRL 0.03fF
C38477 PAND2X1_238/CTRL VDD 0.00fF
C38478 POR2X1_13/A PAND2X1_35/Y 0.02fF
C38479 POR2X1_57/A PAND2X1_360/CTRL 0.01fF
C38480 PAND2X1_849/B POR2X1_263/Y 0.20fF
C38481 POR2X1_49/Y PAND2X1_477/B 0.01fF
C38482 POR2X1_341/A POR2X1_294/A 0.07fF
C38483 POR2X1_29/A PAND2X1_63/B 0.01fF
C38484 POR2X1_842/O POR2X1_456/B 0.16fF
C38485 POR2X1_315/Y POR2X1_298/Y 0.00fF
C38486 POR2X1_68/A PAND2X1_525/O 0.03fF
C38487 POR2X1_46/Y POR2X1_531/CTRL2 0.05fF
C38488 POR2X1_407/A POR2X1_105/Y 0.03fF
C38489 POR2X1_244/B POR2X1_340/CTRL2 0.01fF
C38490 POR2X1_548/B PAND2X1_8/Y 0.82fF
C38491 POR2X1_52/A PAND2X1_190/O 0.05fF
C38492 PAND2X1_360/CTRL2 PAND2X1_843/Y 0.01fF
C38493 POR2X1_776/A POR2X1_191/Y 0.05fF
C38494 PAND2X1_35/Y PAND2X1_214/B 0.01fF
C38495 PAND2X1_228/O VDD 0.00fF
C38496 PAND2X1_41/B POR2X1_206/CTRL2 0.01fF
C38497 PAND2X1_691/Y POR2X1_669/B 0.03fF
C38498 PAND2X1_6/Y POR2X1_830/A 0.01fF
C38499 POR2X1_466/A POR2X1_353/A 0.05fF
C38500 PAND2X1_612/CTRL POR2X1_472/Y 0.13fF
C38501 PAND2X1_58/A POR2X1_725/Y 0.07fF
C38502 POR2X1_853/A VDD 0.25fF
C38503 POR2X1_48/A POR2X1_766/m4_208_n4# 0.08fF
C38504 PAND2X1_830/Y PAND2X1_553/B 0.03fF
C38505 POR2X1_484/O PAND2X1_726/B 0.05fF
C38506 POR2X1_476/A POR2X1_768/a_76_344# 0.01fF
C38507 PAND2X1_23/Y POR2X1_502/A 0.09fF
C38508 POR2X1_43/B POR2X1_237/a_56_344# 0.00fF
C38509 PAND2X1_95/m4_208_n4# PAND2X1_588/m4_208_n4# 0.13fF
C38510 POR2X1_730/Y POR2X1_296/B 0.07fF
C38511 PAND2X1_14/CTRL2 D_INPUT_1 0.03fF
C38512 POR2X1_599/A INPUT_0 0.03fF
C38513 POR2X1_102/Y POR2X1_530/CTRL2 0.01fF
C38514 POR2X1_485/CTRL2 POR2X1_73/Y 0.01fF
C38515 POR2X1_356/A POR2X1_579/Y 0.05fF
C38516 POR2X1_684/CTRL2 POR2X1_42/Y 0.01fF
C38517 PAND2X1_541/CTRL2 POR2X1_7/A 0.03fF
C38518 PAND2X1_80/CTRL2 D_INPUT_1 0.05fF
C38519 POR2X1_391/Y VDD -0.00fF
C38520 POR2X1_654/O PAND2X1_60/B 0.02fF
C38521 POR2X1_346/A POR2X1_507/A 0.02fF
C38522 POR2X1_750/CTRL POR2X1_720/A 0.04fF
C38523 POR2X1_78/A POR2X1_502/O 0.02fF
C38524 PAND2X1_6/Y POR2X1_87/Y 0.00fF
C38525 PAND2X1_94/A POR2X1_14/Y 0.03fF
C38526 POR2X1_193/A POR2X1_795/CTRL 0.08fF
C38527 POR2X1_84/B POR2X1_4/Y 0.01fF
C38528 POR2X1_43/B PAND2X1_480/B 0.17fF
C38529 PAND2X1_651/Y PAND2X1_474/Y 0.03fF
C38530 PAND2X1_390/Y PAND2X1_549/B 0.03fF
C38531 PAND2X1_48/B POR2X1_247/O 0.01fF
C38532 PAND2X1_613/CTRL POR2X1_4/Y -0.00fF
C38533 POR2X1_13/A POR2X1_184/Y 0.23fF
C38534 POR2X1_403/CTRL PAND2X1_60/B 0.02fF
C38535 POR2X1_57/A PAND2X1_787/Y 0.05fF
C38536 POR2X1_41/B PAND2X1_850/CTRL 0.02fF
C38537 POR2X1_590/A POR2X1_741/B 0.13fF
C38538 POR2X1_256/Y VDD 0.08fF
C38539 PAND2X1_213/B PAND2X1_162/CTRL 0.01fF
C38540 POR2X1_401/O PAND2X1_69/A 0.01fF
C38541 PAND2X1_254/O POR2X1_55/Y -0.00fF
C38542 POR2X1_43/B POR2X1_754/A 0.03fF
C38543 PAND2X1_50/CTRL INPUT_6 0.01fF
C38544 POR2X1_260/B POR2X1_383/a_16_28# 0.02fF
C38545 POR2X1_307/a_16_28# POR2X1_796/A 0.01fF
C38546 PAND2X1_651/Y POR2X1_13/A 0.12fF
C38547 PAND2X1_495/m4_208_n4# POR2X1_814/B 0.15fF
C38548 POR2X1_558/CTRL POR2X1_294/B 0.05fF
C38549 POR2X1_391/A POR2X1_391/a_56_344# 0.01fF
C38550 POR2X1_558/CTRL2 POR2X1_264/Y 0.01fF
C38551 PAND2X1_516/O POR2X1_513/Y 0.04fF
C38552 POR2X1_437/Y PAND2X1_592/Y 0.00fF
C38553 POR2X1_448/A PAND2X1_60/B 0.01fF
C38554 POR2X1_625/Y POR2X1_90/Y 0.11fF
C38555 POR2X1_596/A POR2X1_596/Y 0.01fF
C38556 POR2X1_23/Y POR2X1_4/Y 0.10fF
C38557 D_GATE_741 POR2X1_294/B 0.36fF
C38558 POR2X1_616/Y POR2X1_37/Y 0.19fF
C38559 POR2X1_483/A POR2X1_702/O 0.01fF
C38560 POR2X1_536/CTRL POR2X1_250/A 0.09fF
C38561 PAND2X1_642/B POR2X1_293/Y 0.06fF
C38562 POR2X1_356/A POR2X1_614/A 0.18fF
C38563 POR2X1_52/A POR2X1_131/CTRL 0.08fF
C38564 PAND2X1_219/A PAND2X1_853/B 0.03fF
C38565 POR2X1_76/Y POR2X1_541/CTRL 0.01fF
C38566 POR2X1_43/B PAND2X1_341/O 0.03fF
C38567 POR2X1_863/A POR2X1_466/a_16_28# 0.01fF
C38568 PAND2X1_124/Y PAND2X1_199/a_76_28# 0.01fF
C38569 PAND2X1_658/B PAND2X1_174/O 0.01fF
C38570 POR2X1_326/A POR2X1_78/A 0.00fF
C38571 POR2X1_369/O POR2X1_60/A 0.08fF
C38572 POR2X1_13/A PAND2X1_844/B 0.02fF
C38573 POR2X1_355/A POR2X1_260/A 0.01fF
C38574 PAND2X1_41/B POR2X1_456/B 0.03fF
C38575 POR2X1_852/CTRL POR2X1_854/B 0.30fF
C38576 POR2X1_231/CTRL PAND2X1_32/B 0.01fF
C38577 POR2X1_96/Y PAND2X1_61/CTRL2 0.00fF
C38578 POR2X1_614/A POR2X1_795/CTRL 0.00fF
C38579 PAND2X1_131/CTRL PAND2X1_60/B 0.01fF
C38580 PAND2X1_94/A PAND2X1_55/CTRL 0.01fF
C38581 POR2X1_390/B POR2X1_814/B 0.03fF
C38582 PAND2X1_713/A PAND2X1_713/B 0.00fF
C38583 POR2X1_316/CTRL2 PAND2X1_390/Y 0.01fF
C38584 PAND2X1_182/CTRL POR2X1_55/Y 0.01fF
C38585 PAND2X1_65/B PAND2X1_253/CTRL 0.01fF
C38586 PAND2X1_651/Y PAND2X1_197/O 0.02fF
C38587 PAND2X1_858/m4_208_n4# POR2X1_271/m4_208_n4# 0.13fF
C38588 PAND2X1_90/A D_INPUT_1 0.77fF
C38589 PAND2X1_584/a_76_28# POR2X1_774/B 0.01fF
C38590 PAND2X1_493/O POR2X1_60/A 0.03fF
C38591 POR2X1_68/B PAND2X1_132/CTRL 0.00fF
C38592 PAND2X1_212/B PAND2X1_352/CTRL2 0.01fF
C38593 PAND2X1_491/O POR2X1_294/B 0.03fF
C38594 PAND2X1_702/CTRL2 POR2X1_42/Y 0.03fF
C38595 POR2X1_347/A POR2X1_402/CTRL2 0.01fF
C38596 PAND2X1_491/CTRL POR2X1_264/Y 0.01fF
C38597 POR2X1_65/A PAND2X1_641/Y 0.03fF
C38598 POR2X1_407/A POR2X1_114/CTRL2 0.00fF
C38599 POR2X1_32/A PAND2X1_199/O 0.04fF
C38600 POR2X1_128/A POR2X1_186/B 0.01fF
C38601 POR2X1_353/Y POR2X1_353/A 0.04fF
C38602 PAND2X1_108/a_76_28# PAND2X1_60/B 0.02fF
C38603 PAND2X1_785/Y POR2X1_7/A 0.03fF
C38604 POR2X1_308/CTRL POR2X1_308/B 0.04fF
C38605 POR2X1_96/A PAND2X1_656/A 0.02fF
C38606 POR2X1_853/A PAND2X1_32/B 0.06fF
C38607 D_GATE_222 POR2X1_775/O 0.06fF
C38608 POR2X1_390/B POR2X1_325/A 0.03fF
C38609 PAND2X1_273/O PAND2X1_69/A 0.01fF
C38610 POR2X1_131/Y PAND2X1_140/Y 0.05fF
C38611 POR2X1_252/Y POR2X1_60/A 1.05fF
C38612 POR2X1_16/A POR2X1_261/A 0.09fF
C38613 POR2X1_502/A POR2X1_520/A 0.05fF
C38614 PAND2X1_480/O PAND2X1_803/A 0.00fF
C38615 POR2X1_170/B POR2X1_566/B 0.03fF
C38616 PAND2X1_20/A PAND2X1_527/a_76_28# 0.01fF
C38617 POR2X1_391/Y PAND2X1_32/B 0.95fF
C38618 POR2X1_834/Y VDD 1.15fF
C38619 POR2X1_41/B POR2X1_813/Y 0.02fF
C38620 POR2X1_335/A POR2X1_335/B 0.00fF
C38621 POR2X1_283/A PAND2X1_364/O 0.03fF
C38622 POR2X1_48/CTRL2 POR2X1_153/Y 0.05fF
C38623 POR2X1_394/A POR2X1_666/A 0.05fF
C38624 PAND2X1_831/a_16_344# POR2X1_300/Y 0.01fF
C38625 POR2X1_37/Y PAND2X1_840/Y 0.30fF
C38626 POR2X1_210/Y PAND2X1_146/a_16_344# 0.02fF
C38627 PAND2X1_55/Y POR2X1_736/a_76_344# 0.00fF
C38628 POR2X1_42/O D_INPUT_1 0.00fF
C38629 POR2X1_193/A POR2X1_569/A 0.07fF
C38630 PAND2X1_65/B POR2X1_774/A 0.03fF
C38631 POR2X1_356/A POR2X1_440/Y 0.28fF
C38632 PAND2X1_308/Y VDD 0.60fF
C38633 POR2X1_407/Y PAND2X1_743/CTRL 0.01fF
C38634 PAND2X1_6/Y POR2X1_596/A 0.03fF
C38635 PAND2X1_226/O POR2X1_566/B 0.19fF
C38636 PAND2X1_364/B POR2X1_385/CTRL 0.06fF
C38637 POR2X1_840/B PAND2X1_69/A 0.05fF
C38638 POR2X1_303/CTRL2 POR2X1_814/B 0.03fF
C38639 POR2X1_809/A POR2X1_866/B 0.01fF
C38640 POR2X1_603/Y POR2X1_761/A 0.15fF
C38641 POR2X1_532/A POR2X1_804/A 0.08fF
C38642 POR2X1_170/B POR2X1_169/CTRL 0.01fF
C38643 POR2X1_493/a_16_28# POR2X1_572/B 0.02fF
C38644 POR2X1_786/Y POR2X1_702/CTRL2 0.02fF
C38645 PAND2X1_735/CTRL POR2X1_153/Y 0.03fF
C38646 PAND2X1_386/a_56_28# PAND2X1_48/A 0.00fF
C38647 POR2X1_149/B PAND2X1_60/B 0.02fF
C38648 POR2X1_62/Y PAND2X1_340/O 0.01fF
C38649 POR2X1_157/CTRL POR2X1_158/B 0.01fF
C38650 PAND2X1_410/CTRL2 POR2X1_234/A 0.01fF
C38651 POR2X1_614/A POR2X1_220/A 0.32fF
C38652 PAND2X1_693/O POR2X1_383/A 0.04fF
C38653 PAND2X1_490/O POR2X1_532/A 0.02fF
C38654 POR2X1_245/CTRL POR2X1_90/Y 0.01fF
C38655 PAND2X1_630/O POR2X1_7/A 0.05fF
C38656 PAND2X1_6/Y POR2X1_802/CTRL2 0.10fF
C38657 POR2X1_719/B POR2X1_502/A 0.04fF
C38658 POR2X1_38/Y POR2X1_73/Y 0.21fF
C38659 POR2X1_204/CTRL2 PAND2X1_63/B 0.01fF
C38660 POR2X1_350/O POR2X1_854/B 0.04fF
C38661 POR2X1_16/A PAND2X1_592/Y 0.07fF
C38662 PAND2X1_358/A INPUT_0 0.04fF
C38663 PAND2X1_94/A POR2X1_55/Y 0.01fF
C38664 PAND2X1_484/O INPUT_0 0.42fF
C38665 POR2X1_32/A POR2X1_387/O 0.00fF
C38666 PAND2X1_347/Y PAND2X1_359/Y 0.02fF
C38667 PAND2X1_175/B POR2X1_56/Y 0.03fF
C38668 PAND2X1_675/A PAND2X1_181/O 0.05fF
C38669 POR2X1_519/CTRL2 POR2X1_43/B 0.01fF
C38670 PAND2X1_6/Y PAND2X1_422/a_16_344# 0.02fF
C38671 POR2X1_189/Y PAND2X1_728/O 0.02fF
C38672 POR2X1_516/O POR2X1_283/A 0.09fF
C38673 POR2X1_247/a_76_344# POR2X1_260/A 0.01fF
C38674 VDD PAND2X1_2/O 0.00fF
C38675 PAND2X1_7/CTRL POR2X1_260/A 0.01fF
C38676 POR2X1_614/A POR2X1_569/A 0.07fF
C38677 POR2X1_111/CTRL POR2X1_387/Y 0.07fF
C38678 POR2X1_55/Y PAND2X1_336/a_76_28# 0.01fF
C38679 PAND2X1_865/Y PAND2X1_76/Y 0.03fF
C38680 PAND2X1_57/B PAND2X1_399/a_16_344# 0.01fF
C38681 POR2X1_461/Y POR2X1_848/CTRL2 0.01fF
C38682 INPUT_1 PAND2X1_658/A 0.03fF
C38683 PAND2X1_564/a_76_28# POR2X1_394/A 0.02fF
C38684 POR2X1_174/A POR2X1_181/Y 0.03fF
C38685 POR2X1_369/Y POR2X1_236/Y 0.01fF
C38686 PAND2X1_94/A PAND2X1_49/CTRL 0.01fF
C38687 POR2X1_775/A POR2X1_332/CTRL2 0.01fF
C38688 POR2X1_93/A POR2X1_384/CTRL2 0.01fF
C38689 PAND2X1_193/a_16_344# POR2X1_7/Y 0.02fF
C38690 PAND2X1_141/CTRL VDD 0.00fF
C38691 PAND2X1_849/B PAND2X1_6/A 0.07fF
C38692 POR2X1_289/a_16_28# POR2X1_283/A 0.02fF
C38693 PAND2X1_96/B POR2X1_725/Y 0.07fF
C38694 POR2X1_423/Y POR2X1_39/B 0.06fF
C38695 PAND2X1_803/Y POR2X1_142/Y 0.02fF
C38696 POR2X1_711/B PAND2X1_57/B 0.03fF
C38697 POR2X1_244/B POR2X1_228/a_16_28# 0.02fF
C38698 POR2X1_15/O POR2X1_7/A 0.01fF
C38699 POR2X1_283/A POR2X1_382/Y 0.13fF
C38700 POR2X1_544/CTRL POR2X1_854/B 0.01fF
C38701 POR2X1_143/O POR2X1_62/Y 0.11fF
C38702 PAND2X1_552/B POR2X1_394/A 0.03fF
C38703 PAND2X1_483/O PAND2X1_6/A 0.03fF
C38704 PAND2X1_244/B POR2X1_38/Y 0.07fF
C38705 POR2X1_222/A POR2X1_318/A 0.07fF
C38706 PAND2X1_649/A POR2X1_393/CTRL 0.01fF
C38707 PAND2X1_658/A POR2X1_153/Y 0.03fF
C38708 POR2X1_542/B POR2X1_703/A 0.02fF
C38709 POR2X1_228/O POR2X1_294/B 0.02fF
C38710 POR2X1_294/B POR2X1_342/CTRL2 0.01fF
C38711 POR2X1_7/A PAND2X1_656/A 0.03fF
C38712 PAND2X1_6/Y POR2X1_449/A 0.04fF
C38713 POR2X1_119/Y PAND2X1_364/B 0.10fF
C38714 POR2X1_96/A PAND2X1_631/A 0.46fF
C38715 POR2X1_455/A POR2X1_186/B 0.03fF
C38716 POR2X1_394/A PAND2X1_705/O 0.02fF
C38717 PAND2X1_90/A POR2X1_620/B 0.06fF
C38718 PAND2X1_20/A PAND2X1_125/CTRL2 0.01fF
C38719 PAND2X1_690/O PAND2X1_32/B 0.03fF
C38720 PAND2X1_6/CTRL POR2X1_68/B 0.03fF
C38721 PAND2X1_611/CTRL POR2X1_54/Y 0.01fF
C38722 POR2X1_567/A POR2X1_465/B 0.03fF
C38723 POR2X1_568/Y POR2X1_161/Y 0.19fF
C38724 POR2X1_271/A POR2X1_255/Y 0.19fF
C38725 PAND2X1_48/B POR2X1_337/Y 0.07fF
C38726 POR2X1_383/Y VDD 0.13fF
C38727 PAND2X1_853/B POR2X1_816/A 0.03fF
C38728 PAND2X1_23/Y POR2X1_188/Y 0.03fF
C38729 PAND2X1_55/Y POR2X1_540/Y 0.03fF
C38730 PAND2X1_96/B POR2X1_559/A 0.03fF
C38731 POR2X1_73/Y POR2X1_153/Y 0.18fF
C38732 POR2X1_456/B POR2X1_228/Y 0.03fF
C38733 POR2X1_468/Y POR2X1_444/Y 0.01fF
C38734 POR2X1_608/CTRL PAND2X1_56/A 0.01fF
C38735 POR2X1_342/Y VDD 0.10fF
C38736 POR2X1_383/A POR2X1_351/a_76_344# 0.01fF
C38737 VDD POR2X1_77/Y 1.61fF
C38738 PAND2X1_349/A PAND2X1_301/CTRL2 0.01fF
C38739 POR2X1_456/B POR2X1_704/O 0.01fF
C38740 POR2X1_85/Y VDD 0.18fF
C38741 POR2X1_567/A D_GATE_741 0.10fF
C38742 POR2X1_345/O POR2X1_197/Y 0.01fF
C38743 POR2X1_42/Y POR2X1_589/CTRL2 0.01fF
C38744 POR2X1_101/Y POR2X1_276/Y 0.03fF
C38745 POR2X1_13/A POR2X1_387/CTRL 0.01fF
C38746 POR2X1_719/O POR2X1_719/B 0.00fF
C38747 POR2X1_502/A POR2X1_711/Y 0.07fF
C38748 POR2X1_13/A PAND2X1_858/B 0.05fF
C38749 PAND2X1_158/a_16_344# POR2X1_260/A 0.01fF
C38750 PAND2X1_158/O POR2X1_156/Y 0.03fF
C38751 POR2X1_835/B PAND2X1_239/CTRL 0.01fF
C38752 PAND2X1_714/B POR2X1_90/Y 0.00fF
C38753 POR2X1_553/a_76_344# POR2X1_573/A 0.03fF
C38754 POR2X1_471/CTRL PAND2X1_72/A 0.03fF
C38755 POR2X1_155/O POR2X1_728/A 0.00fF
C38756 POR2X1_293/Y POR2X1_387/CTRL2 0.01fF
C38757 PAND2X1_236/m4_208_n4# PAND2X1_52/B 0.04fF
C38758 POR2X1_192/B POR2X1_577/O 0.04fF
C38759 PAND2X1_620/a_76_28# POR2X1_408/Y 0.03fF
C38760 POR2X1_119/Y PAND2X1_560/CTRL 0.10fF
C38761 POR2X1_428/CTRL2 POR2X1_394/A 0.01fF
C38762 POR2X1_378/A POR2X1_62/Y 0.01fF
C38763 POR2X1_539/A POR2X1_737/A 0.03fF
C38764 POR2X1_27/a_16_28# POR2X1_669/B 0.02fF
C38765 POR2X1_88/A D_INPUT_0 0.01fF
C38766 POR2X1_616/Y POR2X1_408/Y 0.01fF
C38767 POR2X1_193/A PAND2X1_72/A 0.03fF
C38768 POR2X1_675/Y POR2X1_733/Y 0.33fF
C38769 POR2X1_579/Y PAND2X1_72/A 0.10fF
C38770 POR2X1_260/B POR2X1_643/Y 0.01fF
C38771 PAND2X1_22/a_16_344# PAND2X1_26/A 0.05fF
C38772 POR2X1_572/B PAND2X1_72/A 0.06fF
C38773 PAND2X1_631/A POR2X1_7/A 0.55fF
C38774 PAND2X1_860/A PAND2X1_795/B 0.00fF
C38775 POR2X1_93/CTRL POR2X1_77/Y 0.01fF
C38776 PAND2X1_52/B PAND2X1_146/O 0.07fF
C38777 POR2X1_813/CTRL POR2X1_32/A 0.01fF
C38778 POR2X1_16/A POR2X1_767/CTRL2 0.01fF
C38779 PAND2X1_663/O GATE_662 0.00fF
C38780 POR2X1_49/Y PAND2X1_206/B 0.14fF
C38781 PAND2X1_319/B POR2X1_39/B 0.03fF
C38782 PAND2X1_713/O POR2X1_394/A 0.02fF
C38783 POR2X1_86/CTRL POR2X1_7/A 0.08fF
C38784 POR2X1_614/A PAND2X1_72/A 3.26fF
C38785 POR2X1_602/O POR2X1_66/A 0.01fF
C38786 POR2X1_428/Y PAND2X1_711/B 0.01fF
C38787 POR2X1_416/B POR2X1_93/A 0.03fF
C38788 POR2X1_16/A PAND2X1_476/A 0.03fF
C38789 POR2X1_344/Y POR2X1_359/CTRL2 0.10fF
C38790 POR2X1_539/A POR2X1_374/a_76_344# 0.01fF
C38791 POR2X1_775/A POR2X1_863/A 0.16fF
C38792 POR2X1_416/B POR2X1_91/Y 0.06fF
C38793 PAND2X1_798/Y PAND2X1_356/O 0.11fF
C38794 POR2X1_408/Y POR2X1_387/CTRL2 0.03fF
C38795 PAND2X1_12/CTRL PAND2X1_11/Y 0.01fF
C38796 POR2X1_23/Y POR2X1_695/Y 0.01fF
C38797 POR2X1_702/A POR2X1_579/CTRL2 0.02fF
C38798 PAND2X1_560/B POR2X1_7/Y 0.03fF
C38799 POR2X1_20/B POR2X1_72/B 0.14fF
C38800 POR2X1_604/CTRL2 POR2X1_40/Y 0.01fF
C38801 POR2X1_242/O POR2X1_776/A 0.01fF
C38802 PAND2X1_808/a_16_344# PAND2X1_860/A 0.01fF
C38803 POR2X1_43/B POR2X1_386/Y 0.03fF
C38804 POR2X1_431/a_76_344# POR2X1_236/Y 0.00fF
C38805 PAND2X1_449/CTRL2 POR2X1_236/Y 0.01fF
C38806 POR2X1_728/A PAND2X1_158/CTRL2 0.00fF
C38807 PAND2X1_43/CTRL POR2X1_852/B 0.02fF
C38808 POR2X1_417/Y PAND2X1_211/O 0.01fF
C38809 POR2X1_89/CTRL POR2X1_60/A 0.01fF
C38810 PAND2X1_422/O PAND2X1_72/A 0.01fF
C38811 POR2X1_416/B POR2X1_416/O 0.02fF
C38812 POR2X1_65/A POR2X1_63/Y 0.08fF
C38813 POR2X1_49/Y POR2X1_65/Y 0.08fF
C38814 POR2X1_579/a_16_28# PAND2X1_32/B 0.02fF
C38815 POR2X1_266/A POR2X1_4/Y 0.03fF
C38816 POR2X1_54/Y POR2X1_734/A 0.05fF
C38817 PAND2X1_247/CTRL2 POR2X1_5/Y 0.00fF
C38818 PAND2X1_644/Y POR2X1_102/Y 0.03fF
C38819 POR2X1_433/Y POR2X1_677/Y 0.02fF
C38820 PAND2X1_449/O VDD 0.00fF
C38821 POR2X1_416/B PAND2X1_545/Y 0.02fF
C38822 POR2X1_23/Y PAND2X1_219/A 0.01fF
C38823 POR2X1_119/Y POR2X1_150/O 0.09fF
C38824 POR2X1_218/Y POR2X1_296/B 0.07fF
C38825 PAND2X1_241/CTRL POR2X1_329/A 0.03fF
C38826 POR2X1_440/Y PAND2X1_72/A 0.03fF
C38827 POR2X1_661/A PAND2X1_69/A 0.07fF
C38828 PAND2X1_612/B POR2X1_654/B 0.03fF
C38829 POR2X1_796/Y POR2X1_330/Y 0.05fF
C38830 POR2X1_57/A POR2X1_825/Y 0.01fF
C38831 PAND2X1_358/CTRL POR2X1_153/Y 0.01fF
C38832 POR2X1_627/CTRL POR2X1_628/Y 0.00fF
C38833 POR2X1_153/Y PAND2X1_207/A 0.17fF
C38834 PAND2X1_678/CTRL2 PAND2X1_804/B 0.01fF
C38835 POR2X1_814/A POR2X1_740/Y 0.12fF
C38836 PAND2X1_75/CTRL POR2X1_740/Y 0.00fF
C38837 PAND2X1_75/CTRL2 POR2X1_741/Y 0.01fF
C38838 POR2X1_703/CTRL POR2X1_169/A 0.01fF
C38839 PAND2X1_689/O POR2X1_121/B 0.10fF
C38840 POR2X1_150/Y PAND2X1_592/O 0.01fF
C38841 PAND2X1_717/A PAND2X1_717/O 0.12fF
C38842 POR2X1_48/A POR2X1_423/Y 0.10fF
C38843 PAND2X1_404/Y POR2X1_5/Y 0.03fF
C38844 POR2X1_159/CTRL2 POR2X1_669/B 0.01fF
C38845 POR2X1_466/A POR2X1_750/B 0.05fF
C38846 POR2X1_188/A POR2X1_858/CTRL 0.01fF
C38847 POR2X1_25/Y D_INPUT_4 0.01fF
C38848 PAND2X1_56/Y PAND2X1_75/O 0.11fF
C38849 POR2X1_603/CTRL POR2X1_597/A 0.00fF
C38850 POR2X1_634/A POR2X1_792/O 0.04fF
C38851 POR2X1_257/A POR2X1_425/CTRL2 0.03fF
C38852 POR2X1_41/B PAND2X1_9/Y 0.00fF
C38853 POR2X1_669/B PAND2X1_195/O 0.02fF
C38854 PAND2X1_58/A POR2X1_811/B 0.02fF
C38855 POR2X1_593/CTRL PAND2X1_72/A 0.11fF
C38856 POR2X1_416/B POR2X1_109/Y 0.03fF
C38857 PAND2X1_93/B POR2X1_480/A 0.07fF
C38858 PAND2X1_251/a_16_344# POR2X1_362/B 0.02fF
C38859 POR2X1_502/A PAND2X1_601/CTRL 0.01fF
C38860 POR2X1_29/A POR2X1_391/A 0.03fF
C38861 POR2X1_135/Y POR2X1_23/Y 0.42fF
C38862 PAND2X1_90/A INPUT_3 0.03fF
C38863 PAND2X1_454/O PAND2X1_446/Y 0.01fF
C38864 POR2X1_864/A PAND2X1_744/O 0.00fF
C38865 PAND2X1_93/B POR2X1_243/Y 0.23fF
C38866 POR2X1_474/CTRL POR2X1_777/B 0.22fF
C38867 POR2X1_661/O POR2X1_661/Y 0.00fF
C38868 POR2X1_84/CTRL2 POR2X1_84/B 0.00fF
C38869 POR2X1_12/A PAND2X1_709/CTRL2 0.09fF
C38870 POR2X1_416/Y POR2X1_412/a_16_28# 0.03fF
C38871 POR2X1_257/A POR2X1_481/Y 0.06fF
C38872 POR2X1_491/CTRL2 POR2X1_72/B 0.01fF
C38873 POR2X1_445/A PAND2X1_55/Y 0.03fF
C38874 PAND2X1_81/CTRL2 PAND2X1_9/Y 0.00fF
C38875 POR2X1_348/O POR2X1_814/A 0.08fF
C38876 POR2X1_130/A POR2X1_479/B 0.05fF
C38877 POR2X1_842/O PAND2X1_57/B 0.07fF
C38878 PAND2X1_55/Y POR2X1_643/Y 0.01fF
C38879 PAND2X1_58/A PAND2X1_525/O 0.02fF
C38880 POR2X1_96/A POR2X1_271/a_76_344# 0.01fF
C38881 PAND2X1_835/Y POR2X1_20/B 0.00fF
C38882 INPUT_3 PAND2X1_19/O 0.01fF
C38883 POR2X1_22/A D_INPUT_5 0.02fF
C38884 POR2X1_78/A POR2X1_480/A 0.10fF
C38885 PAND2X1_80/CTRL PAND2X1_73/Y 0.03fF
C38886 POR2X1_411/B POR2X1_90/Y 9.63fF
C38887 PAND2X1_412/m4_208_n4# PAND2X1_277/m4_208_n4# 0.13fF
C38888 POR2X1_42/O INPUT_3 0.09fF
C38889 POR2X1_278/Y POR2X1_487/O 0.01fF
C38890 PAND2X1_90/A PAND2X1_93/B 0.01fF
C38891 POR2X1_760/A PAND2X1_656/A 0.04fF
C38892 PAND2X1_496/CTRL2 D_INPUT_0 0.01fF
C38893 POR2X1_807/CTRL2 POR2X1_294/B 0.03fF
C38894 POR2X1_383/A PAND2X1_256/O 0.14fF
C38895 POR2X1_306/CTRL2 PAND2X1_454/B 0.01fF
C38896 POR2X1_673/CTRL2 PAND2X1_8/Y 0.03fF
C38897 POR2X1_822/a_16_28# POR2X1_102/Y 0.03fF
C38898 POR2X1_174/B POR2X1_192/Y 0.10fF
C38899 POR2X1_106/CTRL PAND2X1_553/B 0.07fF
C38900 PAND2X1_833/O POR2X1_482/Y 0.06fF
C38901 POR2X1_142/CTRL PAND2X1_738/Y 0.02fF
C38902 POR2X1_669/B POR2X1_669/O 0.08fF
C38903 POR2X1_78/B POR2X1_602/B 0.06fF
C38904 POR2X1_356/A POR2X1_590/A 0.08fF
C38905 PAND2X1_63/Y POR2X1_260/B 0.05fF
C38906 POR2X1_829/A POR2X1_603/Y 0.03fF
C38907 PAND2X1_10/O PAND2X1_55/Y 0.01fF
C38908 POR2X1_594/Y POR2X1_32/A 0.01fF
C38909 POR2X1_529/CTRL POR2X1_29/A 0.03fF
C38910 INPUT_1 POR2X1_19/CTRL2 0.00fF
C38911 POR2X1_638/B POR2X1_66/A 0.02fF
C38912 POR2X1_23/Y POR2X1_816/A 2.08fF
C38913 POR2X1_96/A PAND2X1_78/O 0.05fF
C38914 PAND2X1_90/A POR2X1_78/A 5.57fF
C38915 POR2X1_119/CTRL2 POR2X1_102/Y 0.01fF
C38916 POR2X1_728/B POR2X1_330/Y 0.02fF
C38917 POR2X1_81/O POR2X1_494/Y 0.00fF
C38918 PAND2X1_23/Y POR2X1_637/m4_208_n4# 0.12fF
C38919 D_INPUT_5 POR2X1_1/CTRL2 0.06fF
C38920 POR2X1_78/CTRL2 D_INPUT_0 0.01fF
C38921 POR2X1_626/O PAND2X1_6/A 0.03fF
C38922 POR2X1_84/A POR2X1_68/B 0.07fF
C38923 POR2X1_750/B POR2X1_586/CTRL2 0.01fF
C38924 PAND2X1_6/Y D_INPUT_0 0.10fF
C38925 PAND2X1_224/O POR2X1_192/B 0.04fF
C38926 PAND2X1_224/CTRL POR2X1_191/Y -0.01fF
C38927 POR2X1_218/Y POR2X1_267/Y 0.11fF
C38928 POR2X1_49/Y PAND2X1_149/CTRL2 0.01fF
C38929 PAND2X1_6/Y POR2X1_811/A 0.01fF
C38930 POR2X1_391/A POR2X1_546/A 0.00fF
C38931 POR2X1_271/Y POR2X1_275/CTRL 0.00fF
C38932 POR2X1_121/O POR2X1_655/A 0.01fF
C38933 PAND2X1_580/B PAND2X1_363/Y 0.02fF
C38934 PAND2X1_57/B PAND2X1_41/B 6.20fF
C38935 POR2X1_798/CTRL2 POR2X1_468/B 0.01fF
C38936 POR2X1_68/A POR2X1_296/B 0.78fF
C38937 POR2X1_66/A POR2X1_570/B 0.02fF
C38938 POR2X1_41/B PAND2X1_614/O 0.07fF
C38939 PAND2X1_755/a_56_28# PAND2X1_41/B 0.00fF
C38940 PAND2X1_641/O POR2X1_63/Y 0.03fF
C38941 POR2X1_278/Y PAND2X1_740/CTRL 0.04fF
C38942 POR2X1_102/Y POR2X1_599/A 0.08fF
C38943 PAND2X1_474/A PAND2X1_735/a_56_28# 0.00fF
C38944 POR2X1_66/A PAND2X1_311/O 0.02fF
C38945 POR2X1_41/B PAND2X1_499/CTRL2 0.06fF
C38946 POR2X1_135/Y POR2X1_45/O 0.01fF
C38947 PAND2X1_494/O POR2X1_78/A 0.05fF
C38948 POR2X1_660/Y POR2X1_804/A 0.05fF
C38949 POR2X1_808/A PAND2X1_599/CTRL2 0.05fF
C38950 POR2X1_494/a_16_28# POR2X1_29/A 0.02fF
C38951 POR2X1_370/Y POR2X1_325/A 0.00fF
C38952 POR2X1_52/A PAND2X1_455/a_16_344# 0.03fF
C38953 POR2X1_330/Y PAND2X1_516/m4_208_n4# 0.06fF
C38954 PAND2X1_433/m4_208_n4# PAND2X1_591/m4_208_n4# 0.13fF
C38955 PAND2X1_61/Y PAND2X1_523/CTRL 0.01fF
C38956 PAND2X1_220/Y PAND2X1_553/B 0.10fF
C38957 PAND2X1_682/CTRL POR2X1_467/Y 0.00fF
C38958 POR2X1_623/B PAND2X1_69/A 0.02fF
C38959 POR2X1_419/Y PAND2X1_506/O 0.00fF
C38960 POR2X1_14/Y POR2X1_584/O 0.15fF
C38961 D_INPUT_3 D_INPUT_0 1.00fF
C38962 D_INPUT_0 POR2X1_575/CTRL2 0.01fF
C38963 POR2X1_254/A POR2X1_341/CTRL 0.01fF
C38964 PAND2X1_20/A PAND2X1_83/CTRL 0.01fF
C38965 PAND2X1_571/Y VDD 0.00fF
C38966 POR2X1_75/CTRL2 POR2X1_60/A 0.00fF
C38967 PAND2X1_63/Y PAND2X1_265/CTRL2 0.15fF
C38968 PAND2X1_425/Y PAND2X1_2/CTRL2 0.01fF
C38969 POR2X1_322/CTRL2 POR2X1_376/B 0.00fF
C38970 PAND2X1_801/B POR2X1_7/B 0.01fF
C38971 PAND2X1_48/B POR2X1_543/A 0.23fF
C38972 PAND2X1_460/Y VDD 0.15fF
C38973 POR2X1_852/B POR2X1_740/Y 0.10fF
C38974 PAND2X1_557/A PAND2X1_357/Y 0.03fF
C38975 POR2X1_271/B PAND2X1_508/Y 0.03fF
C38976 POR2X1_46/Y POR2X1_236/Y 0.26fF
C38977 POR2X1_13/Y POR2X1_250/A 0.03fF
C38978 POR2X1_149/B POR2X1_750/B 0.03fF
C38979 POR2X1_406/Y PAND2X1_734/B 0.01fF
C38980 POR2X1_550/A POR2X1_849/A 0.04fF
C38981 POR2X1_69/CTRL PAND2X1_69/A 0.00fF
C38982 POR2X1_192/Y POR2X1_544/A 0.05fF
C38983 PAND2X1_862/B PAND2X1_659/O 0.08fF
C38984 POR2X1_260/B POR2X1_260/A 1.80fF
C38985 POR2X1_16/A PAND2X1_207/CTRL -0.02fF
C38986 POR2X1_51/A POR2X1_13/A 0.03fF
C38987 POR2X1_68/A PAND2X1_679/CTRL2 0.07fF
C38988 PAND2X1_254/O POR2X1_511/Y 0.04fF
C38989 POR2X1_675/O POR2X1_540/A 0.01fF
C38990 PAND2X1_486/O VDD 0.00fF
C38991 POR2X1_7/B PAND2X1_8/Y 0.03fF
C38992 POR2X1_852/a_16_28# POR2X1_852/A 0.03fF
C38993 POR2X1_596/A POR2X1_467/Y 0.03fF
C38994 PAND2X1_114/Y VDD -0.00fF
C38995 PAND2X1_55/Y PAND2X1_58/CTRL 0.01fF
C38996 PAND2X1_652/A PAND2X1_192/O 0.05fF
C38997 PAND2X1_638/a_16_344# POR2X1_752/Y 0.02fF
C38998 POR2X1_750/B POR2X1_644/A 0.00fF
C38999 POR2X1_5/Y POR2X1_382/a_56_344# 0.00fF
C39000 PAND2X1_48/B POR2X1_723/CTRL2 0.00fF
C39001 POR2X1_566/A POR2X1_776/B 0.00fF
C39002 PAND2X1_108/CTRL POR2X1_814/A 0.09fF
C39003 POR2X1_590/A POR2X1_569/A 0.08fF
C39004 POR2X1_244/B POR2X1_579/Y 0.03fF
C39005 PAND2X1_734/B POR2X1_293/Y 0.03fF
C39006 PAND2X1_742/B VDD 0.02fF
C39007 PAND2X1_821/CTRL VDD 0.00fF
C39008 PAND2X1_131/CTRL2 POR2X1_130/Y 0.03fF
C39009 POR2X1_43/B PAND2X1_473/B 0.04fF
C39010 POR2X1_693/Y POR2X1_697/O 0.01fF
C39011 POR2X1_669/B POR2X1_428/CTRL2 0.03fF
C39012 PAND2X1_840/A POR2X1_236/Y 0.00fF
C39013 PAND2X1_6/Y PAND2X1_90/Y 0.12fF
C39014 PAND2X1_641/a_76_28# POR2X1_23/Y 0.01fF
C39015 PAND2X1_20/A PAND2X1_63/B 0.03fF
C39016 POR2X1_94/A PAND2X1_521/CTRL 0.04fF
C39017 POR2X1_376/B POR2X1_90/Y 0.07fF
C39018 PAND2X1_613/CTRL POR2X1_620/B 0.05fF
C39019 PAND2X1_172/CTRL POR2X1_174/A 0.01fF
C39020 PAND2X1_284/O VDD 0.00fF
C39021 POR2X1_78/B POR2X1_712/Y 0.03fF
C39022 POR2X1_52/A PAND2X1_191/Y 0.05fF
C39023 POR2X1_502/A POR2X1_733/A 0.07fF
C39024 POR2X1_327/Y POR2X1_270/Y 0.01fF
C39025 POR2X1_465/A POR2X1_563/Y 0.06fF
C39026 POR2X1_32/A PAND2X1_301/CTRL2 0.03fF
C39027 INPUT_1 POR2X1_753/Y 3.05fF
C39028 PAND2X1_48/B PAND2X1_280/O 0.05fF
C39029 POR2X1_109/CTRL POR2X1_109/Y 0.00fF
C39030 POR2X1_60/A PAND2X1_550/B 0.02fF
C39031 POR2X1_66/B PAND2X1_397/O 0.09fF
C39032 PAND2X1_65/B PAND2X1_153/CTRL2 0.01fF
C39033 PAND2X1_23/Y POR2X1_284/CTRL2 0.01fF
C39034 PAND2X1_768/Y PAND2X1_359/B 0.02fF
C39035 PAND2X1_429/O POR2X1_260/A 0.01fF
C39036 POR2X1_68/A POR2X1_214/CTRL2 0.04fF
C39037 POR2X1_139/CTRL2 VDD -0.00fF
C39038 POR2X1_865/B POR2X1_475/A 0.06fF
C39039 POR2X1_720/B INPUT_0 0.04fF
C39040 PAND2X1_274/CTRL POR2X1_273/Y 0.01fF
C39041 POR2X1_206/A POR2X1_208/Y 0.31fF
C39042 POR2X1_351/B POR2X1_856/B 0.02fF
C39043 POR2X1_52/Y VDD 0.00fF
C39044 POR2X1_404/B POR2X1_35/Y 0.00fF
C39045 POR2X1_539/A POR2X1_302/B 0.03fF
C39046 PAND2X1_349/A PAND2X1_140/CTRL 0.01fF
C39047 PAND2X1_137/Y PAND2X1_675/A 0.03fF
C39048 PAND2X1_62/m4_208_n4# PAND2X1_6/A 0.12fF
C39049 POR2X1_312/Y PAND2X1_854/A 0.02fF
C39050 POR2X1_66/A PAND2X1_384/O 0.01fF
C39051 POR2X1_423/Y PAND2X1_840/O 0.08fF
C39052 POR2X1_5/Y POR2X1_395/Y 0.19fF
C39053 POR2X1_287/B PAND2X1_60/B 0.05fF
C39054 POR2X1_278/Y PAND2X1_359/CTRL2 0.00fF
C39055 POR2X1_68/A POR2X1_215/a_16_28# 0.02fF
C39056 POR2X1_335/Y VDD 0.15fF
C39057 POR2X1_496/Y PAND2X1_507/a_16_344# -0.01fF
C39058 POR2X1_252/CTRL2 PAND2X1_6/A 0.04fF
C39059 POR2X1_66/B POR2X1_752/O 0.01fF
C39060 POR2X1_164/Y POR2X1_40/Y 0.01fF
C39061 POR2X1_343/Y POR2X1_556/A 0.05fF
C39062 PAND2X1_48/B POR2X1_363/CTRL 0.11fF
C39063 POR2X1_255/a_76_344# PAND2X1_349/A 0.00fF
C39064 POR2X1_567/B POR2X1_566/a_16_28# 0.08fF
C39065 PAND2X1_556/CTRL2 PAND2X1_348/A 0.03fF
C39066 POR2X1_66/B PAND2X1_748/a_16_344# 0.01fF
C39067 POR2X1_814/B PAND2X1_63/B 0.03fF
C39068 POR2X1_311/Y PAND2X1_348/A 0.07fF
C39069 PAND2X1_808/Y POR2X1_488/Y 0.04fF
C39070 PAND2X1_197/Y POR2X1_57/Y 0.00fF
C39071 POR2X1_56/B POR2X1_305/Y 0.00fF
C39072 PAND2X1_41/B POR2X1_707/Y 0.04fF
C39073 PAND2X1_9/Y POR2X1_77/Y 0.03fF
C39074 POR2X1_483/A PAND2X1_60/B 0.03fF
C39075 POR2X1_537/a_16_28# POR2X1_590/A 0.03fF
C39076 POR2X1_834/Y POR2X1_808/A 0.14fF
C39077 POR2X1_326/CTRL2 PAND2X1_41/B 0.03fF
C39078 POR2X1_42/Y POR2X1_396/CTRL2 0.01fF
C39079 PAND2X1_241/Y VDD 0.30fF
C39080 POR2X1_51/B INPUT_7 1.58fF
C39081 POR2X1_41/B PAND2X1_852/B 0.16fF
C39082 PAND2X1_572/O INPUT_0 0.02fF
C39083 POR2X1_83/Y D_INPUT_0 0.03fF
C39084 POR2X1_730/Y POR2X1_186/Y 0.08fF
C39085 POR2X1_52/A POR2X1_90/Y 1.40fF
C39086 POR2X1_96/A PAND2X1_243/O 0.04fF
C39087 POR2X1_537/CTRL2 POR2X1_862/B 0.00fF
C39088 POR2X1_828/Y POR2X1_687/A 0.01fF
C39089 PAND2X1_653/Y POR2X1_7/B 0.03fF
C39090 PAND2X1_421/CTRL PAND2X1_69/A 0.01fF
C39091 PAND2X1_96/B PAND2X1_176/CTRL 0.10fF
C39092 POR2X1_83/B PAND2X1_156/A 0.52fF
C39093 POR2X1_210/a_16_28# POR2X1_210/A 0.04fF
C39094 D_GATE_741 PAND2X1_504/CTRL 0.03fF
C39095 PAND2X1_65/B POR2X1_352/CTRL 0.01fF
C39096 PAND2X1_63/Y PAND2X1_55/Y 0.03fF
C39097 PAND2X1_57/B POR2X1_228/Y 10.51fF
C39098 POR2X1_152/A POR2X1_90/Y 0.03fF
C39099 POR2X1_138/CTRL PAND2X1_32/B 0.02fF
C39100 PAND2X1_651/Y PAND2X1_506/O -0.00fF
C39101 INPUT_6 INPUT_5 0.10fF
C39102 POR2X1_861/A POR2X1_296/B 0.19fF
C39103 POR2X1_391/CTRL POR2X1_546/A 0.01fF
C39104 POR2X1_376/B PAND2X1_732/A 0.03fF
C39105 POR2X1_203/CTRL2 POR2X1_579/Y 0.00fF
C39106 POR2X1_634/A PAND2X1_48/A 0.10fF
C39107 POR2X1_49/Y PAND2X1_560/B 0.00fF
C39108 POR2X1_192/Y POR2X1_190/m4_208_n4# 0.04fF
C39109 D_GATE_222 POR2X1_556/Y 0.03fF
C39110 PAND2X1_495/O PAND2X1_55/Y 0.00fF
C39111 POR2X1_326/A POR2X1_798/CTRL2 0.00fF
C39112 POR2X1_390/B VDD 0.02fF
C39113 POR2X1_25/Y POR2X1_698/CTRL2 0.01fF
C39114 PAND2X1_41/B POR2X1_227/O 0.01fF
C39115 POR2X1_82/O POR2X1_16/A 0.01fF
C39116 POR2X1_564/Y POR2X1_569/A 0.13fF
C39117 PAND2X1_784/CTRL2 POR2X1_245/Y 0.02fF
C39118 POR2X1_347/A POR2X1_347/a_16_28# 0.10fF
C39119 INPUT_1 POR2X1_627/m4_208_n4# 0.12fF
C39120 POR2X1_840/B POR2X1_723/B 0.05fF
C39121 POR2X1_51/B INPUT_4 0.03fF
C39122 POR2X1_356/A POR2X1_338/O 0.02fF
C39123 POR2X1_96/A PAND2X1_728/CTRL 0.01fF
C39124 PAND2X1_48/B POR2X1_711/m4_208_n4# 0.07fF
C39125 PAND2X1_23/Y POR2X1_711/a_16_28# 0.03fF
C39126 POR2X1_407/A POR2X1_685/B 0.01fF
C39127 PAND2X1_636/a_76_28# POR2X1_584/Y 0.05fF
C39128 VDD PAND2X1_157/CTRL2 -0.00fF
C39129 POR2X1_356/A PAND2X1_824/a_16_344# 0.02fF
C39130 POR2X1_809/A PAND2X1_679/CTRL 0.01fF
C39131 POR2X1_865/B POR2X1_218/A 0.07fF
C39132 PAND2X1_23/Y POR2X1_510/Y 0.03fF
C39133 POR2X1_242/O POR2X1_191/Y 0.17fF
C39134 PAND2X1_605/O INPUT_0 0.05fF
C39135 PAND2X1_219/a_56_28# POR2X1_591/Y 0.00fF
C39136 POR2X1_57/A POR2X1_518/Y 2.49fF
C39137 POR2X1_119/Y PAND2X1_240/CTRL2 0.02fF
C39138 POR2X1_575/B POR2X1_575/O 0.55fF
C39139 D_GATE_662 POR2X1_319/Y 0.07fF
C39140 POR2X1_57/A PAND2X1_472/A 0.03fF
C39141 POR2X1_751/CTRL POR2X1_816/A 0.01fF
C39142 POR2X1_614/A POR2X1_203/CTRL2 0.02fF
C39143 POR2X1_447/B POR2X1_194/A 0.08fF
C39144 PAND2X1_600/O PAND2X1_72/A 0.03fF
C39145 POR2X1_750/B PAND2X1_179/CTRL2 0.01fF
C39146 POR2X1_596/A PAND2X1_743/O 0.02fF
C39147 D_INPUT_0 POR2X1_500/CTRL 0.01fF
C39148 POR2X1_366/Y POR2X1_317/A 0.09fF
C39149 POR2X1_722/A VDD 0.00fF
C39150 PAND2X1_6/Y POR2X1_348/CTRL2 0.03fF
C39151 PAND2X1_388/Y PAND2X1_370/CTRL 0.01fF
C39152 POR2X1_855/B PAND2X1_599/a_16_344# 0.01fF
C39153 POR2X1_301/O PAND2X1_60/B 0.01fF
C39154 POR2X1_334/Y PAND2X1_261/CTRL2 0.05fF
C39155 POR2X1_547/O POR2X1_550/A 0.01fF
C39156 D_INPUT_0 PAND2X1_52/B 0.18fF
C39157 POR2X1_591/Y POR2X1_73/Y 0.07fF
C39158 PAND2X1_551/Y PAND2X1_854/A 0.42fF
C39159 PAND2X1_206/a_76_28# POR2X1_153/Y 0.05fF
C39160 POR2X1_811/A PAND2X1_52/B 0.01fF
C39161 POR2X1_567/A POR2X1_231/A 0.01fF
C39162 PAND2X1_785/Y POR2X1_153/Y 0.03fF
C39163 POR2X1_814/B POR2X1_552/A 0.03fF
C39164 PAND2X1_563/A POR2X1_7/B 0.03fF
C39165 POR2X1_362/B POR2X1_362/CTRL 0.01fF
C39166 POR2X1_16/A PAND2X1_776/O 0.04fF
C39167 PAND2X1_55/Y POR2X1_260/A 0.10fF
C39168 POR2X1_130/A PAND2X1_48/A 0.28fF
C39169 POR2X1_390/B POR2X1_741/Y 0.03fF
C39170 POR2X1_346/CTRL PAND2X1_60/B 0.01fF
C39171 PAND2X1_470/A POR2X1_73/Y 0.00fF
C39172 PAND2X1_214/A PAND2X1_207/A 0.01fF
C39173 PAND2X1_598/a_76_28# POR2X1_394/A 0.03fF
C39174 POR2X1_72/B POR2X1_372/CTRL2 0.03fF
C39175 POR2X1_590/A PAND2X1_72/A 0.46fF
C39176 POR2X1_7/B PAND2X1_337/CTRL 0.01fF
C39177 PAND2X1_770/O POR2X1_766/Y 0.00fF
C39178 POR2X1_546/A POR2X1_294/A 0.03fF
C39179 D_GATE_222 POR2X1_259/a_16_28# 0.02fF
C39180 POR2X1_38/Y PAND2X1_656/A 0.06fF
C39181 POR2X1_94/A PAND2X1_102/a_16_344# 0.01fF
C39182 POR2X1_8/Y PAND2X1_341/a_16_344# 0.02fF
C39183 POR2X1_184/Y PAND2X1_301/CTRL2 0.00fF
C39184 POR2X1_68/A POR2X1_543/CTRL 0.01fF
C39185 POR2X1_167/O POR2X1_73/Y 0.04fF
C39186 POR2X1_566/A POR2X1_192/B 0.10fF
C39187 POR2X1_296/B POR2X1_138/A 0.01fF
C39188 POR2X1_41/B POR2X1_595/O 0.10fF
C39189 PAND2X1_659/Y POR2X1_498/CTRL 0.01fF
C39190 POR2X1_311/CTRL2 POR2X1_142/Y 0.01fF
C39191 POR2X1_57/A POR2X1_527/Y 0.01fF
C39192 POR2X1_836/A POR2X1_568/A 0.03fF
C39193 POR2X1_740/Y POR2X1_151/Y 0.02fF
C39194 POR2X1_52/A POR2X1_110/Y 0.10fF
C39195 PAND2X1_162/A PAND2X1_162/CTRL2 0.00fF
C39196 PAND2X1_865/Y PAND2X1_480/B 0.05fF
C39197 POR2X1_366/a_16_28# PAND2X1_6/Y 0.02fF
C39198 POR2X1_294/B POR2X1_113/B 0.03fF
C39199 POR2X1_407/Y POR2X1_260/A 0.05fF
C39200 PAND2X1_94/A POR2X1_205/A 0.78fF
C39201 POR2X1_416/B POR2X1_24/m4_208_n4# 0.04fF
C39202 PAND2X1_48/B POR2X1_342/O 0.01fF
C39203 POR2X1_96/A PAND2X1_850/Y 0.27fF
C39204 PAND2X1_679/CTRL POR2X1_728/A 0.00fF
C39205 POR2X1_20/a_76_344# POR2X1_4/Y 0.02fF
C39206 POR2X1_3/a_16_28# POR2X1_260/A 0.01fF
C39207 POR2X1_131/Y PAND2X1_140/A 0.07fF
C39208 PAND2X1_852/O PAND2X1_659/Y 0.01fF
C39209 POR2X1_294/A POR2X1_712/Y 0.07fF
C39210 INPUT_6 PAND2X1_157/O 0.02fF
C39211 PAND2X1_90/Y PAND2X1_52/B 12.84fF
C39212 POR2X1_520/O POR2X1_520/A 0.01fF
C39213 POR2X1_556/A POR2X1_624/Y 0.12fF
C39214 PAND2X1_69/A POR2X1_737/A 0.04fF
C39215 POR2X1_614/A POR2X1_537/Y 0.03fF
C39216 POR2X1_793/O PAND2X1_52/B 0.04fF
C39217 PAND2X1_20/A PAND2X1_234/CTRL2 0.03fF
C39218 POR2X1_337/A POR2X1_260/A 0.00fF
C39219 PAND2X1_65/B POR2X1_181/A 0.01fF
C39220 PAND2X1_860/A PAND2X1_795/O 0.04fF
C39221 POR2X1_294/A POR2X1_500/Y 0.03fF
C39222 POR2X1_854/O POR2X1_776/A 0.01fF
C39223 POR2X1_153/Y PAND2X1_656/A 0.12fF
C39224 POR2X1_846/A POR2X1_14/Y 0.03fF
C39225 POR2X1_57/A PAND2X1_325/O 0.04fF
C39226 POR2X1_66/B POR2X1_9/Y 0.19fF
C39227 PAND2X1_270/O PAND2X1_508/Y 0.01fF
C39228 POR2X1_725/a_16_28# POR2X1_711/Y 0.03fF
C39229 POR2X1_20/B POR2X1_616/CTRL 0.01fF
C39230 PAND2X1_217/CTRL PAND2X1_267/Y 0.01fF
C39231 POR2X1_327/Y POR2X1_101/Y 0.03fF
C39232 PAND2X1_640/B POR2X1_20/B 0.03fF
C39233 PAND2X1_93/B POR2X1_243/a_16_28# 0.03fF
C39234 POR2X1_509/O POR2X1_857/B 0.05fF
C39235 PAND2X1_94/A POR2X1_129/Y 0.03fF
C39236 POR2X1_859/CTRL POR2X1_66/A 0.05fF
C39237 POR2X1_857/B PAND2X1_72/A 0.05fF
C39238 POR2X1_814/B PAND2X1_234/CTRL2 0.02fF
C39239 POR2X1_40/CTRL2 POR2X1_25/Y 0.01fF
C39240 INPUT_1 POR2X1_4/a_16_28# 0.08fF
C39241 POR2X1_112/CTRL POR2X1_510/Y 0.02fF
C39242 PAND2X1_447/CTRL2 POR2X1_102/Y 0.01fF
C39243 POR2X1_416/B PAND2X1_551/A 0.07fF
C39244 POR2X1_456/B POR2X1_579/B 0.02fF
C39245 POR2X1_754/A POR2X1_90/CTRL 0.00fF
C39246 POR2X1_510/Y POR2X1_735/a_16_28# 0.03fF
C39247 POR2X1_329/A PAND2X1_561/A 0.34fF
C39248 PAND2X1_646/CTRL2 POR2X1_612/Y 0.01fF
C39249 POR2X1_499/a_76_344# POR2X1_341/A 0.01fF
C39250 POR2X1_287/A POR2X1_287/a_16_28# 0.03fF
C39251 PAND2X1_852/B POR2X1_77/Y 0.03fF
C39252 POR2X1_316/Y POR2X1_387/Y 0.07fF
C39253 POR2X1_853/A POR2X1_568/A 0.03fF
C39254 POR2X1_741/A POR2X1_186/B 0.00fF
C39255 POR2X1_287/B POR2X1_486/O 0.01fF
C39256 POR2X1_96/A POR2X1_826/a_16_28# 0.08fF
C39257 POR2X1_300/Y POR2X1_153/Y 0.00fF
C39258 POR2X1_703/A POR2X1_703/a_16_28# 0.01fF
C39259 POR2X1_416/B POR2X1_425/Y 0.91fF
C39260 POR2X1_67/Y POR2X1_5/Y 0.03fF
C39261 POR2X1_567/A POR2X1_339/CTRL 0.25fF
C39262 POR2X1_865/CTRL PAND2X1_52/B 0.01fF
C39263 INPUT_1 PAND2X1_631/A 0.03fF
C39264 POR2X1_9/Y POR2X1_859/A 0.12fF
C39265 POR2X1_634/A POR2X1_461/Y 0.17fF
C39266 POR2X1_502/A PAND2X1_438/O 0.04fF
C39267 PAND2X1_39/B POR2X1_806/O 0.01fF
C39268 PAND2X1_601/O POR2X1_296/B 0.04fF
C39269 POR2X1_102/Y PAND2X1_791/a_16_344# 0.01fF
C39270 PAND2X1_862/a_16_344# PAND2X1_858/Y 0.01fF
C39271 POR2X1_266/A POR2X1_620/B 0.36fF
C39272 POR2X1_825/Y POR2X1_396/CTRL 0.00fF
C39273 POR2X1_361/CTRL PAND2X1_72/A 0.01fF
C39274 PAND2X1_631/A POR2X1_153/Y 0.03fF
C39275 PAND2X1_827/CTRL2 POR2X1_296/B 0.00fF
C39276 POR2X1_188/A POR2X1_841/a_76_344# 0.00fF
C39277 POR2X1_846/A POR2X1_55/Y 1.25fF
C39278 POR2X1_479/CTRL2 POR2X1_66/A 0.02fF
C39279 POR2X1_66/B POR2X1_274/A 0.03fF
C39280 D_INPUT_5 PAND2X1_425/O 0.17fF
C39281 POR2X1_673/Y PAND2X1_529/O 0.03fF
C39282 POR2X1_356/A POR2X1_440/B 0.68fF
C39283 PAND2X1_20/A POR2X1_567/B 0.05fF
C39284 POR2X1_99/CTRL2 POR2X1_243/Y 0.03fF
C39285 POR2X1_852/B PAND2X1_67/O 0.08fF
C39286 PAND2X1_97/Y PAND2X1_351/Y 0.01fF
C39287 PAND2X1_193/Y POR2X1_38/Y 0.02fF
C39288 POR2X1_130/O POR2X1_343/Y 0.02fF
C39289 POR2X1_482/O POR2X1_60/A 0.02fF
C39290 POR2X1_675/CTRL POR2X1_466/A 0.13fF
C39291 POR2X1_411/B INPUT_0 0.18fF
C39292 POR2X1_78/B PAND2X1_39/B 0.10fF
C39293 PAND2X1_57/B POR2X1_657/Y 0.02fF
C39294 POR2X1_260/B POR2X1_718/A 0.63fF
C39295 PAND2X1_58/A POR2X1_296/B 0.16fF
C39296 POR2X1_23/Y PAND2X1_332/CTRL2 0.03fF
C39297 POR2X1_777/B POR2X1_458/a_16_28# 0.07fF
C39298 POR2X1_60/Y D_INPUT_0 0.09fF
C39299 POR2X1_814/B POR2X1_567/B 0.10fF
C39300 POR2X1_660/Y POR2X1_794/B 0.03fF
C39301 POR2X1_257/A PAND2X1_707/O 0.17fF
C39302 POR2X1_807/A POR2X1_807/CTRL2 0.01fF
C39303 POR2X1_748/A POR2X1_669/B 0.10fF
C39304 POR2X1_20/B POR2X1_7/B 0.21fF
C39305 POR2X1_41/B PAND2X1_247/O 0.12fF
C39306 POR2X1_195/A POR2X1_207/A 0.00fF
C39307 POR2X1_65/A POR2X1_283/CTRL2 0.03fF
C39308 POR2X1_196/Y POR2X1_814/A 0.04fF
C39309 POR2X1_94/A POR2X1_29/A 0.85fF
C39310 POR2X1_96/A POR2X1_299/a_16_28# 0.01fF
C39311 PAND2X1_415/CTRL2 POR2X1_293/Y 0.01fF
C39312 POR2X1_744/Y POR2X1_743/Y 0.00fF
C39313 POR2X1_67/m4_208_n4# POR2X1_236/Y 0.09fF
C39314 PAND2X1_394/CTRL POR2X1_330/Y 0.02fF
C39315 POR2X1_411/B PAND2X1_218/CTRL 0.01fF
C39316 POR2X1_491/O POR2X1_102/Y 0.01fF
C39317 POR2X1_150/Y PAND2X1_794/B 0.03fF
C39318 POR2X1_548/B POR2X1_624/Y 0.03fF
C39319 POR2X1_48/A POR2X1_393/CTRL 0.01fF
C39320 POR2X1_411/B POR2X1_234/CTRL2 0.01fF
C39321 POR2X1_451/CTRL2 POR2X1_750/B 0.01fF
C39322 PAND2X1_571/CTRL VDD 0.00fF
C39323 POR2X1_850/B POR2X1_807/A 0.01fF
C39324 POR2X1_632/A POR2X1_590/A 0.01fF
C39325 POR2X1_633/O POR2X1_68/B 0.01fF
C39326 PAND2X1_193/Y POR2X1_153/Y 0.16fF
C39327 POR2X1_225/a_16_28# POR2X1_5/Y 0.03fF
C39328 POR2X1_285/O POR2X1_590/A 0.01fF
C39329 POR2X1_16/A POR2X1_827/CTRL2 0.04fF
C39330 POR2X1_54/Y POR2X1_672/A 0.06fF
C39331 PAND2X1_90/A POR2X1_84/A 0.03fF
C39332 POR2X1_65/A PAND2X1_168/Y 0.00fF
C39333 POR2X1_467/Y PAND2X1_90/Y 0.12fF
C39334 POR2X1_16/A PAND2X1_439/CTRL2 0.01fF
C39335 POR2X1_356/A POR2X1_66/A 0.05fF
C39336 POR2X1_78/B PAND2X1_20/A 0.30fF
C39337 POR2X1_148/CTRL2 PAND2X1_69/A 0.01fF
C39338 PAND2X1_660/CTRL2 PAND2X1_660/B 0.01fF
C39339 POR2X1_66/Y PAND2X1_69/A 0.04fF
C39340 POR2X1_334/B POR2X1_493/A 0.05fF
C39341 POR2X1_9/Y PAND2X1_358/A 0.07fF
C39342 POR2X1_48/A PAND2X1_707/Y 0.00fF
C39343 PAND2X1_65/B PAND2X1_766/O 0.03fF
C39344 POR2X1_441/O PAND2X1_732/A 0.06fF
C39345 POR2X1_614/A POR2X1_319/A 0.12fF
C39346 POR2X1_48/CTRL2 POR2X1_72/B 0.03fF
C39347 PAND2X1_65/B PAND2X1_423/CTRL2 0.03fF
C39348 POR2X1_319/A POR2X1_317/Y 0.02fF
C39349 PAND2X1_57/B POR2X1_657/O 0.05fF
C39350 PAND2X1_827/O POR2X1_741/Y 0.46fF
C39351 POR2X1_409/B POR2X1_42/Y 0.07fF
C39352 PAND2X1_675/A POR2X1_23/Y 1.04fF
C39353 POR2X1_482/Y VDD 0.35fF
C39354 POR2X1_614/Y PAND2X1_754/a_16_344# 0.05fF
C39355 POR2X1_23/Y PAND2X1_469/B 0.01fF
C39356 PAND2X1_667/m4_208_n4# POR2X1_590/A 0.15fF
C39357 POR2X1_67/Y PAND2X1_789/CTRL 0.01fF
C39358 POR2X1_271/Y INPUT_0 0.00fF
C39359 POR2X1_241/B POR2X1_776/B 0.03fF
C39360 PAND2X1_402/O POR2X1_236/Y 0.02fF
C39361 PAND2X1_478/B PAND2X1_480/B 0.14fF
C39362 PAND2X1_283/CTRL POR2X1_66/A 0.01fF
C39363 POR2X1_57/A PAND2X1_212/CTRL2 0.03fF
C39364 D_INPUT_7 PAND2X1_18/B 0.05fF
C39365 POR2X1_750/B PAND2X1_8/Y 0.01fF
C39366 PAND2X1_7/CTRL2 POR2X1_555/B 0.01fF
C39367 PAND2X1_683/a_76_28# POR2X1_78/B 0.01fF
C39368 POR2X1_58/Y POR2X1_83/B 0.03fF
C39369 POR2X1_72/B PAND2X1_579/B 0.03fF
C39370 POR2X1_629/O PAND2X1_69/A 0.16fF
C39371 PAND2X1_627/O POR2X1_852/B 0.16fF
C39372 POR2X1_240/a_56_344# PAND2X1_88/Y 0.00fF
C39373 PAND2X1_90/A PAND2X1_9/CTRL2 0.01fF
C39374 POR2X1_38/O POR2X1_38/B 0.02fF
C39375 POR2X1_78/B POR2X1_814/B 1.57fF
C39376 POR2X1_411/B PAND2X1_348/CTRL 0.01fF
C39377 POR2X1_130/A POR2X1_288/A 0.50fF
C39378 POR2X1_37/Y POR2X1_380/O 0.03fF
C39379 POR2X1_274/Y VDD 0.01fF
C39380 POR2X1_276/A POR2X1_624/Y 0.02fF
C39381 POR2X1_267/B VDD 0.10fF
C39382 POR2X1_32/a_16_28# POR2X1_32/A 0.14fF
C39383 POR2X1_502/A POR2X1_593/B 0.03fF
C39384 POR2X1_502/A POR2X1_752/Y 0.03fF
C39385 PAND2X1_61/Y POR2X1_88/Y 0.12fF
C39386 POR2X1_72/B POR2X1_331/A 0.01fF
C39387 POR2X1_106/Y VDD -0.00fF
C39388 POR2X1_376/B INPUT_0 0.54fF
C39389 POR2X1_504/CTRL2 POR2X1_20/B 0.03fF
C39390 POR2X1_407/A POR2X1_660/CTRL 0.03fF
C39391 POR2X1_333/A D_GATE_662 0.10fF
C39392 POR2X1_243/Y PAND2X1_65/Y 0.07fF
C39393 PAND2X1_581/a_56_28# INPUT_6 0.00fF
C39394 POR2X1_78/B POR2X1_325/A 0.03fF
C39395 POR2X1_502/A PAND2X1_387/O 0.34fF
C39396 POR2X1_777/B POR2X1_404/Y 0.01fF
C39397 POR2X1_72/Y PAND2X1_217/B 0.73fF
C39398 POR2X1_94/O POR2X1_14/Y 0.18fF
C39399 PAND2X1_73/Y PAND2X1_518/CTRL2 0.09fF
C39400 POR2X1_49/Y PAND2X1_466/CTRL2 0.01fF
C39401 POR2X1_260/B POR2X1_725/Y 0.07fF
C39402 POR2X1_72/CTRL POR2X1_71/Y 0.01fF
C39403 PAND2X1_794/O PAND2X1_794/B 0.08fF
C39404 POR2X1_68/A POR2X1_864/CTRL2 0.10fF
C39405 PAND2X1_65/B POR2X1_220/Y 0.06fF
C39406 PAND2X1_736/A POR2X1_40/Y 0.07fF
C39407 POR2X1_65/A POR2X1_56/B 0.10fF
C39408 PAND2X1_96/B POR2X1_296/B 0.10fF
C39409 POR2X1_121/B PAND2X1_743/CTRL 0.07fF
C39410 POR2X1_556/A POR2X1_186/B 0.03fF
C39411 PAND2X1_580/B VDD 0.04fF
C39412 POR2X1_370/Y VDD 0.23fF
C39413 POR2X1_233/CTRL2 POR2X1_236/Y 0.01fF
C39414 PAND2X1_658/A POR2X1_72/B 1.76fF
C39415 POR2X1_16/A POR2X1_600/Y 0.01fF
C39416 POR2X1_614/A POR2X1_812/A 0.00fF
C39417 PAND2X1_431/CTRL POR2X1_440/Y 0.01fF
C39418 POR2X1_296/Y PAND2X1_69/A 0.04fF
C39419 POR2X1_866/A POR2X1_596/CTRL2 0.13fF
C39420 POR2X1_130/O POR2X1_624/Y 0.02fF
C39421 PAND2X1_808/B PAND2X1_808/O 0.00fF
C39422 PAND2X1_65/B POR2X1_404/Y 0.03fF
C39423 POR2X1_338/CTRL2 POR2X1_97/A 0.01fF
C39424 POR2X1_48/A POR2X1_766/CTRL 0.02fF
C39425 POR2X1_673/O PAND2X1_6/A 0.05fF
C39426 POR2X1_49/Y PAND2X1_478/O 0.12fF
C39427 POR2X1_49/Y POR2X1_521/CTRL2 0.00fF
C39428 PAND2X1_73/CTRL2 PAND2X1_69/A 0.09fF
C39429 POR2X1_78/B POR2X1_513/B 0.07fF
C39430 POR2X1_260/B POR2X1_596/O 0.01fF
C39431 POR2X1_68/A POR2X1_186/Y 0.11fF
C39432 POR2X1_66/A POR2X1_569/A 0.07fF
C39433 PAND2X1_691/Y POR2X1_48/A 0.06fF
C39434 PAND2X1_824/B POR2X1_447/A 0.06fF
C39435 PAND2X1_96/B PAND2X1_74/CTRL 0.01fF
C39436 POR2X1_325/a_16_28# PAND2X1_93/B 0.01fF
C39437 PAND2X1_499/a_56_28# POR2X1_293/Y 0.00fF
C39438 POR2X1_626/m4_208_n4# POR2X1_408/Y 0.06fF
C39439 POR2X1_102/Y PAND2X1_572/O 0.01fF
C39440 POR2X1_16/A POR2X1_438/Y 0.22fF
C39441 POR2X1_614/A POR2X1_801/CTRL2 0.02fF
C39442 POR2X1_378/CTRL D_INPUT_1 0.00fF
C39443 PAND2X1_840/A PAND2X1_499/CTRL 0.00fF
C39444 PAND2X1_117/CTRL VDD 0.00fF
C39445 POR2X1_255/a_76_344# POR2X1_184/Y 0.01fF
C39446 POR2X1_302/B PAND2X1_69/A 0.03fF
C39447 POR2X1_52/A INPUT_0 1.22fF
C39448 POR2X1_462/B POR2X1_734/A 0.05fF
C39449 PAND2X1_7/Y POR2X1_631/B 0.03fF
C39450 POR2X1_272/Y POR2X1_42/Y 0.36fF
C39451 POR2X1_114/B POR2X1_850/A 0.03fF
C39452 PAND2X1_48/B POR2X1_471/CTRL 0.01fF
C39453 POR2X1_72/B POR2X1_73/Y 2.94fF
C39454 POR2X1_260/B POR2X1_559/A 0.05fF
C39455 PAND2X1_39/B POR2X1_294/A 16.64fF
C39456 POR2X1_360/A PAND2X1_57/B 0.08fF
C39457 POR2X1_857/B POR2X1_244/B 0.03fF
C39458 PAND2X1_264/CTRL POR2X1_669/B 0.05fF
C39459 PAND2X1_94/A POR2X1_35/O 0.03fF
C39460 POR2X1_702/B POR2X1_786/Y 0.02fF
C39461 POR2X1_65/A PAND2X1_724/CTRL2 0.03fF
C39462 POR2X1_49/Y PAND2X1_724/CTRL 0.01fF
C39463 PAND2X1_495/CTRL2 POR2X1_814/B 0.11fF
C39464 POR2X1_96/A POR2X1_406/CTRL 0.01fF
C39465 POR2X1_254/Y POR2X1_294/B 0.05fF
C39466 PAND2X1_810/A PAND2X1_568/B 8.74fF
C39467 PAND2X1_784/A POR2X1_387/Y 0.06fF
C39468 POR2X1_416/B PAND2X1_717/A 0.03fF
C39469 POR2X1_278/Y POR2X1_488/Y 0.07fF
C39470 POR2X1_370/Y POR2X1_741/Y 0.03fF
C39471 POR2X1_267/B PAND2X1_32/B 0.01fF
C39472 POR2X1_625/CTRL POR2X1_90/Y 0.01fF
C39473 PAND2X1_57/B POR2X1_756/O 0.01fF
C39474 POR2X1_16/A POR2X1_487/O 0.32fF
C39475 PAND2X1_661/Y POR2X1_60/A 0.03fF
C39476 PAND2X1_750/O POR2X1_749/Y 0.07fF
C39477 POR2X1_275/a_56_344# PAND2X1_785/Y 0.00fF
C39478 POR2X1_327/Y PAND2X1_431/O 0.09fF
C39479 POR2X1_502/A POR2X1_477/A 0.03fF
C39480 POR2X1_270/CTRL POR2X1_814/B 0.03fF
C39481 POR2X1_356/A POR2X1_802/B 0.03fF
C39482 PAND2X1_214/A PAND2X1_656/A 1.74fF
C39483 PAND2X1_94/A PAND2X1_235/CTRL2 0.00fF
C39484 PAND2X1_20/A POR2X1_141/A 0.00fF
C39485 PAND2X1_562/O VDD 0.00fF
C39486 POR2X1_137/Y PAND2X1_41/B 0.05fF
C39487 POR2X1_409/Y POR2X1_29/A 0.01fF
C39488 POR2X1_92/O POR2X1_49/Y 0.01fF
C39489 POR2X1_446/B POR2X1_540/Y 0.05fF
C39490 POR2X1_406/Y PAND2X1_716/CTRL 0.00fF
C39491 POR2X1_264/Y POR2X1_572/O 0.00fF
C39492 POR2X1_433/m4_208_n4# PAND2X1_549/B 0.15fF
C39493 POR2X1_52/A PAND2X1_717/CTRL2 0.00fF
C39494 INPUT_1 PAND2X1_77/CTRL 0.05fF
C39495 POR2X1_390/B POR2X1_105/CTRL2 0.00fF
C39496 POR2X1_440/B PAND2X1_72/A 0.01fF
C39497 POR2X1_32/A PAND2X1_777/CTRL2 0.01fF
C39498 PAND2X1_48/B POR2X1_193/A 0.03fF
C39499 POR2X1_57/A PAND2X1_803/A 0.03fF
C39500 PAND2X1_23/Y POR2X1_578/Y 0.03fF
C39501 PAND2X1_48/B POR2X1_579/Y 0.03fF
C39502 PAND2X1_652/Y POR2X1_594/Y 0.13fF
C39503 POR2X1_334/B POR2X1_124/O 0.02fF
C39504 PAND2X1_217/B PAND2X1_349/A 0.06fF
C39505 POR2X1_770/CTRL POR2X1_770/A 0.01fF
C39506 PAND2X1_864/CTRL2 PAND2X1_810/A 0.01fF
C39507 PAND2X1_211/m4_208_n4# PAND2X1_566/m4_208_n4# 0.13fF
C39508 PAND2X1_859/A POR2X1_7/A 0.03fF
C39509 PAND2X1_309/O POR2X1_740/Y 0.02fF
C39510 PAND2X1_309/CTRL POR2X1_741/Y 0.00fF
C39511 POR2X1_614/A POR2X1_483/B 0.05fF
C39512 POR2X1_94/O PAND2X1_472/B 0.04fF
C39513 POR2X1_304/Y POR2X1_90/Y 0.01fF
C39514 POR2X1_43/B PAND2X1_793/Y 0.03fF
C39515 POR2X1_829/A POR2X1_599/A 0.01fF
C39516 POR2X1_219/B POR2X1_215/CTRL2 0.13fF
C39517 PAND2X1_244/B POR2X1_72/B 0.18fF
C39518 POR2X1_567/B POR2X1_726/CTRL 0.00fF
C39519 POR2X1_525/Y PAND2X1_546/Y 0.03fF
C39520 VDD PAND2X1_347/O 0.00fF
C39521 PAND2X1_58/A POR2X1_590/Y 0.03fF
C39522 POR2X1_180/B POR2X1_186/Y 0.03fF
C39523 POR2X1_327/CTRL2 PAND2X1_63/Y 0.03fF
C39524 POR2X1_131/O POR2X1_13/A 0.18fF
C39525 PAND2X1_738/Y PAND2X1_388/CTRL 0.14fF
C39526 PAND2X1_247/O POR2X1_77/Y 0.03fF
C39527 GATE_479 PAND2X1_550/B 5.87fF
C39528 POR2X1_215/CTRL PAND2X1_88/Y 0.01fF
C39529 PAND2X1_602/Y POR2X1_755/O 0.01fF
C39530 POR2X1_804/A PAND2X1_131/a_76_28# 0.03fF
C39531 PAND2X1_131/CTRL POR2X1_318/A 0.01fF
C39532 POR2X1_57/A PAND2X1_673/Y 0.03fF
C39533 PAND2X1_48/B POR2X1_789/A 0.03fF
C39534 POR2X1_124/O POR2X1_124/B 0.01fF
C39535 POR2X1_216/O VDD 0.00fF
C39536 VDD POR2X1_359/Y 0.09fF
C39537 POR2X1_839/CTRL POR2X1_566/B 0.01fF
C39538 POR2X1_499/a_16_28# POR2X1_294/A 0.00fF
C39539 INPUT_6 PAND2X1_587/Y 0.01fF
C39540 POR2X1_266/A POR2X1_78/A 0.06fF
C39541 PAND2X1_245/a_16_344# PAND2X1_71/Y 0.01fF
C39542 POR2X1_614/A PAND2X1_48/B 0.06fF
C39543 PAND2X1_94/A PAND2X1_395/O 0.15fF
C39544 INPUT_2 POR2X1_119/CTRL2 0.01fF
C39545 PAND2X1_714/CTRL POR2X1_73/Y 0.01fF
C39546 POR2X1_860/A POR2X1_260/A 0.03fF
C39547 POR2X1_686/A POR2X1_260/A 0.02fF
C39548 POR2X1_537/Y POR2X1_590/A 2.36fF
C39549 POR2X1_485/O PAND2X1_550/B 0.01fF
C39550 POR2X1_805/Y POR2X1_294/A 0.03fF
C39551 PAND2X1_349/A VDD 1.02fF
C39552 POR2X1_356/A POR2X1_532/A 0.09fF
C39553 POR2X1_241/B POR2X1_192/B 0.03fF
C39554 POR2X1_724/a_16_28# POR2X1_724/A 0.01fF
C39555 PAND2X1_63/B VDD 1.47fF
C39556 POR2X1_41/B PAND2X1_213/Y 0.07fF
C39557 POR2X1_840/CTRL PAND2X1_55/Y 0.01fF
C39558 POR2X1_809/A POR2X1_864/CTRL 0.01fF
C39559 POR2X1_323/Y POR2X1_73/Y 0.01fF
C39560 PAND2X1_6/Y D_GATE_222 0.06fF
C39561 PAND2X1_20/A POR2X1_294/A 0.29fF
C39562 PAND2X1_658/B POR2X1_816/A 0.19fF
C39563 PAND2X1_803/a_76_28# POR2X1_60/A 0.05fF
C39564 POR2X1_779/A POR2X1_407/A 0.04fF
C39565 POR2X1_311/O POR2X1_481/A 0.01fF
C39566 PAND2X1_290/CTRL POR2X1_66/A 0.01fF
C39567 POR2X1_861/CTRL POR2X1_501/B 0.03fF
C39568 VDD PAND2X1_114/B 0.14fF
C39569 POR2X1_96/A POR2X1_7/A 0.26fF
C39570 PAND2X1_810/O PAND2X1_366/Y 0.01fF
C39571 POR2X1_740/Y PAND2X1_88/Y 0.05fF
C39572 POR2X1_96/A PAND2X1_344/a_76_28# 0.01fF
C39573 PAND2X1_631/m4_208_n4# POR2X1_55/Y 0.07fF
C39574 PAND2X1_651/Y POR2X1_239/CTRL2 0.00fF
C39575 POR2X1_276/A POR2X1_276/CTRL2 0.01fF
C39576 POR2X1_51/A POR2X1_744/CTRL2 0.01fF
C39577 POR2X1_378/O POR2X1_62/Y 0.12fF
C39578 PAND2X1_109/O POR2X1_97/A 0.01fF
C39579 POR2X1_728/O POR2X1_730/Y 0.01fF
C39580 POR2X1_40/Y POR2X1_7/Y 0.10fF
C39581 POR2X1_78/A PAND2X1_179/O 0.04fF
C39582 POR2X1_590/A POR2X1_532/O 0.03fF
C39583 POR2X1_264/Y PAND2X1_60/B 0.08fF
C39584 POR2X1_558/O POR2X1_558/A 0.21fF
C39585 POR2X1_793/A POR2X1_789/CTRL 0.08fF
C39586 POR2X1_775/A PAND2X1_173/O 0.02fF
C39587 POR2X1_407/A PAND2X1_153/O 0.00fF
C39588 POR2X1_369/CTRL POR2X1_236/Y 0.01fF
C39589 INPUT_1 PAND2X1_38/CTRL 0.01fF
C39590 PAND2X1_59/B PAND2X1_52/B 0.01fF
C39591 POR2X1_327/CTRL2 POR2X1_260/A 0.03fF
C39592 POR2X1_814/B POR2X1_294/A 0.22fF
C39593 POR2X1_785/A POR2X1_566/B 0.03fF
C39594 PAND2X1_55/Y POR2X1_725/Y 0.08fF
C39595 PAND2X1_48/B POR2X1_440/Y 0.09fF
C39596 PAND2X1_216/B PAND2X1_804/B 0.07fF
C39597 POR2X1_405/a_16_28# POR2X1_737/A 0.03fF
C39598 PAND2X1_96/B PAND2X1_125/m4_208_n4# 0.15fF
C39599 POR2X1_38/B POR2X1_565/a_16_28# 0.03fF
C39600 POR2X1_285/B POR2X1_590/A 0.33fF
C39601 POR2X1_292/CTRL2 POR2X1_411/B 0.05fF
C39602 POR2X1_693/Y PAND2X1_550/Y 0.75fF
C39603 POR2X1_222/Y POR2X1_569/A 0.07fF
C39604 D_INPUT_0 PAND2X1_351/A 0.07fF
C39605 POR2X1_66/A PAND2X1_72/A 10.69fF
C39606 POR2X1_103/O PAND2X1_738/Y 0.02fF
C39607 POR2X1_192/Y POR2X1_544/B 0.03fF
C39608 PAND2X1_686/CTRL2 POR2X1_42/Y 0.01fF
C39609 PAND2X1_81/B PAND2X1_63/B 0.12fF
C39610 POR2X1_81/CTRL2 PAND2X1_862/B 0.01fF
C39611 POR2X1_16/A PAND2X1_401/CTRL2 0.11fF
C39612 POR2X1_220/A POR2X1_532/A 0.01fF
C39613 POR2X1_287/B PAND2X1_122/CTRL 0.01fF
C39614 POR2X1_407/A POR2X1_407/CTRL 0.01fF
C39615 PAND2X1_195/O POR2X1_39/B 0.15fF
C39616 POR2X1_495/CTRL2 POR2X1_39/B 0.02fF
C39617 POR2X1_355/B POR2X1_564/B 0.05fF
C39618 POR2X1_108/CTRL POR2X1_387/Y 0.13fF
C39619 POR2X1_186/Y POR2X1_169/A 0.03fF
C39620 POR2X1_731/CTRL POR2X1_738/A 0.01fF
C39621 PAND2X1_63/B PAND2X1_32/B 0.03fF
C39622 PAND2X1_831/Y POR2X1_91/Y 0.03fF
C39623 PAND2X1_143/CTRL2 PAND2X1_8/Y 0.00fF
C39624 PAND2X1_215/B POR2X1_394/A 0.07fF
C39625 PAND2X1_865/Y PAND2X1_473/B 0.07fF
C39626 POR2X1_72/B PAND2X1_207/A 0.01fF
C39627 POR2X1_865/CTRL2 POR2X1_101/Y 0.03fF
C39628 POR2X1_684/Y VDD 0.12fF
C39629 POR2X1_275/O POR2X1_129/Y 0.01fF
C39630 POR2X1_341/Y POR2X1_351/CTRL 0.01fF
C39631 POR2X1_20/B PAND2X1_206/B 0.07fF
C39632 POR2X1_814/B PAND2X1_102/CTRL 0.08fF
C39633 POR2X1_130/CTRL2 PAND2X1_6/Y 0.02fF
C39634 VDD POR2X1_552/A 0.00fF
C39635 POR2X1_532/A POR2X1_569/A 0.07fF
C39636 POR2X1_327/Y PAND2X1_23/Y 0.06fF
C39637 POR2X1_177/CTRL PAND2X1_552/B 0.01fF
C39638 PAND2X1_427/O PAND2X1_72/A 0.01fF
C39639 POR2X1_456/B POR2X1_112/Y 0.03fF
C39640 POR2X1_86/CTRL2 VDD 0.00fF
C39641 POR2X1_124/B POR2X1_768/CTRL2 0.01fF
C39642 PAND2X1_270/O POR2X1_283/A 0.05fF
C39643 PAND2X1_620/CTRL PAND2X1_651/Y 0.00fF
C39644 POR2X1_614/A POR2X1_210/B 0.01fF
C39645 PAND2X1_698/CTRL POR2X1_532/A 0.01fF
C39646 POR2X1_68/B POR2X1_773/B 0.20fF
C39647 POR2X1_809/A POR2X1_803/A 0.25fF
C39648 PAND2X1_6/A POR2X1_394/A 0.17fF
C39649 POR2X1_407/Y POR2X1_596/O 0.01fF
C39650 PAND2X1_612/B POR2X1_814/A 0.00fF
C39651 PAND2X1_704/CTRL POR2X1_90/Y 0.01fF
C39652 PAND2X1_482/CTRL2 POR2X1_786/Y 0.02fF
C39653 POR2X1_54/Y POR2X1_624/B 0.00fF
C39654 POR2X1_780/B POR2X1_796/A 0.04fF
C39655 POR2X1_507/B D_GATE_741 0.04fF
C39656 POR2X1_813/Y PAND2X1_63/B 0.01fF
C39657 PAND2X1_341/B PAND2X1_341/O 0.01fF
C39658 POR2X1_45/Y PAND2X1_199/B 0.00fF
C39659 PAND2X1_82/Y PAND2X1_397/O 0.01fF
C39660 POR2X1_849/A PAND2X1_202/a_16_344# 0.07fF
C39661 POR2X1_477/A POR2X1_188/Y 0.03fF
C39662 POR2X1_57/A PAND2X1_722/CTRL2 0.03fF
C39663 POR2X1_514/O PAND2X1_48/A 0.09fF
C39664 PAND2X1_457/Y PAND2X1_464/B 0.02fF
C39665 POR2X1_527/CTRL PAND2X1_549/B 0.01fF
C39666 VDD POR2X1_342/A -0.00fF
C39667 POR2X1_116/A PAND2X1_39/B 0.02fF
C39668 POR2X1_199/a_56_344# POR2X1_199/B 0.00fF
C39669 POR2X1_54/Y POR2X1_859/CTRL2 0.03fF
C39670 PAND2X1_6/Y POR2X1_552/O 0.02fF
C39671 POR2X1_54/Y POR2X1_88/A 0.04fF
C39672 PAND2X1_657/B POR2X1_816/A 0.04fF
C39673 POR2X1_218/CTRL POR2X1_362/A 0.01fF
C39674 POR2X1_218/O POR2X1_276/Y 0.01fF
C39675 POR2X1_673/Y PAND2X1_63/B 0.03fF
C39676 POR2X1_101/Y POR2X1_249/Y 0.05fF
C39677 D_INPUT_5 PAND2X1_425/Y 0.04fF
C39678 POR2X1_609/Y POR2X1_399/Y 0.00fF
C39679 PAND2X1_87/O D_INPUT_0 0.15fF
C39680 POR2X1_239/a_16_28# POR2X1_153/Y 0.06fF
C39681 POR2X1_346/a_16_28# POR2X1_507/A 0.06fF
C39682 POR2X1_110/Y POR2X1_417/CTRL 0.01fF
C39683 POR2X1_411/B PAND2X1_340/B 0.03fF
C39684 POR2X1_385/Y PAND2X1_389/O 0.04fF
C39685 POR2X1_110/O POR2X1_73/Y 0.02fF
C39686 POR2X1_305/CTRL2 POR2X1_55/Y 0.01fF
C39687 POR2X1_41/B POR2X1_416/B 0.31fF
C39688 POR2X1_702/O POR2X1_186/B 0.01fF
C39689 PAND2X1_651/Y PAND2X1_500/CTRL2 0.06fF
C39690 POR2X1_740/Y POR2X1_568/B 0.05fF
C39691 PAND2X1_453/CTRL2 POR2X1_77/Y 0.10fF
C39692 POR2X1_510/Y POR2X1_553/O 0.02fF
C39693 POR2X1_48/A PAND2X1_447/a_16_344# 0.02fF
C39694 PAND2X1_96/B PAND2X1_759/CTRL2 0.01fF
C39695 POR2X1_567/A POR2X1_341/Y 0.22fF
C39696 POR2X1_441/a_16_28# POR2X1_669/B 0.02fF
C39697 PAND2X1_521/m4_208_n4# PAND2X1_522/m4_208_n4# 0.13fF
C39698 POR2X1_280/Y POR2X1_394/A 1.50fF
C39699 POR2X1_860/CTRL POR2X1_244/Y 0.01fF
C39700 POR2X1_445/A POR2X1_446/B 0.03fF
C39701 POR2X1_528/Y PAND2X1_156/A 0.46fF
C39702 POR2X1_453/Y POR2X1_436/B 0.01fF
C39703 POR2X1_802/B PAND2X1_72/A 0.98fF
C39704 POR2X1_520/a_16_28# POR2X1_559/A 0.01fF
C39705 POR2X1_57/A PAND2X1_352/O 0.01fF
C39706 POR2X1_119/Y PAND2X1_469/Y 0.15fF
C39707 PAND2X1_718/CTRL POR2X1_77/Y 0.01fF
C39708 POR2X1_212/CTRL POR2X1_191/Y 0.21fF
C39709 PAND2X1_682/CTRL2 POR2X1_728/A 0.00fF
C39710 PAND2X1_476/A POR2X1_235/CTRL2 0.00fF
C39711 POR2X1_760/A PAND2X1_361/CTRL2 0.03fF
C39712 PAND2X1_94/A PAND2X1_527/CTRL 0.01fF
C39713 POR2X1_84/B POR2X1_84/A 0.08fF
C39714 POR2X1_294/Y POR2X1_294/CTRL2 0.00fF
C39715 POR2X1_695/O POR2X1_23/Y 0.01fF
C39716 POR2X1_309/CTRL2 POR2X1_411/B 0.01fF
C39717 POR2X1_383/A POR2X1_383/a_16_28# 0.02fF
C39718 POR2X1_222/Y PAND2X1_72/A 0.03fF
C39719 D_GATE_222 PAND2X1_52/B 0.07fF
C39720 POR2X1_23/Y PAND2X1_477/CTRL2 0.15fF
C39721 POR2X1_25/Y POR2X1_26/CTRL 0.01fF
C39722 POR2X1_65/CTRL POR2X1_40/Y 0.01fF
C39723 POR2X1_416/B POR2X1_256/Y 0.06fF
C39724 POR2X1_68/A POR2X1_717/B 0.03fF
C39725 POR2X1_119/Y PAND2X1_123/a_16_344# 0.04fF
C39726 PAND2X1_483/CTRL POR2X1_252/Y 0.01fF
C39727 PAND2X1_483/CTRL2 PAND2X1_631/A 0.00fF
C39728 POR2X1_102/Y POR2X1_411/B 6.68fF
C39729 POR2X1_837/A VDD 0.00fF
C39730 PAND2X1_411/a_76_28# PAND2X1_52/B 0.02fF
C39731 POR2X1_848/O PAND2X1_90/Y 0.01fF
C39732 POR2X1_67/Y PAND2X1_381/CTRL 0.01fF
C39733 POR2X1_598/a_16_28# POR2X1_294/A 0.03fF
C39734 POR2X1_327/Y POR2X1_809/A 0.02fF
C39735 PAND2X1_213/Y POR2X1_77/Y 0.00fF
C39736 POR2X1_23/Y PAND2X1_214/CTRL 0.01fF
C39737 PAND2X1_72/a_16_344# PAND2X1_72/A 0.02fF
C39738 POR2X1_9/Y POR2X1_625/Y 0.04fF
C39739 POR2X1_728/CTRL2 POR2X1_814/A 0.02fF
C39740 POR2X1_343/Y PAND2X1_60/B 0.05fF
C39741 PAND2X1_635/Y INPUT_5 0.03fF
C39742 POR2X1_509/O POR2X1_532/A 0.02fF
C39743 PAND2X1_586/O PAND2X1_48/A 0.04fF
C39744 POR2X1_20/B POR2X1_750/B 0.03fF
C39745 POR2X1_99/B POR2X1_259/B 0.22fF
C39746 POR2X1_119/Y POR2X1_394/A 0.97fF
C39747 POR2X1_532/A PAND2X1_72/A 7.82fF
C39748 POR2X1_137/B POR2X1_734/A 0.03fF
C39749 POR2X1_284/B POR2X1_284/a_16_28# 0.08fF
C39750 POR2X1_153/Y PAND2X1_199/CTRL 0.08fF
C39751 POR2X1_477/B POR2X1_477/a_16_28# 0.02fF
C39752 POR2X1_116/A POR2X1_814/B 0.49fF
C39753 POR2X1_257/A POR2X1_40/Y 0.08fF
C39754 PAND2X1_220/Y POR2X1_20/B 0.03fF
C39755 PAND2X1_431/CTRL POR2X1_590/A 0.00fF
C39756 PAND2X1_39/B POR2X1_94/A 0.09fF
C39757 POR2X1_809/CTRL POR2X1_121/B 0.04fF
C39758 POR2X1_110/Y PAND2X1_716/B 0.03fF
C39759 POR2X1_260/B POR2X1_811/B 0.03fF
C39760 POR2X1_814/A POR2X1_220/Y 0.11fF
C39761 POR2X1_686/a_16_28# PAND2X1_72/A 0.02fF
C39762 PAND2X1_116/O POR2X1_150/Y 0.09fF
C39763 PAND2X1_472/CTRL POR2X1_39/B 0.09fF
C39764 PAND2X1_170/CTRL2 PAND2X1_326/B 0.01fF
C39765 POR2X1_263/Y POR2X1_669/B 0.02fF
C39766 POR2X1_49/a_16_28# POR2X1_38/B 0.03fF
C39767 POR2X1_411/A VDD 0.03fF
C39768 PAND2X1_677/CTRL2 POR2X1_260/B 0.01fF
C39769 POR2X1_399/CTRL2 POR2X1_20/B 0.01fF
C39770 POR2X1_834/Y PAND2X1_56/A 0.05fF
C39771 PAND2X1_65/B POR2X1_818/CTRL2 0.09fF
C39772 POR2X1_826/Y POR2X1_826/O 0.01fF
C39773 POR2X1_116/A POR2X1_325/A 0.03fF
C39774 PAND2X1_858/CTRL2 PAND2X1_850/Y 0.05fF
C39775 POR2X1_48/A POR2X1_764/m4_208_n4# 0.08fF
C39776 POR2X1_150/Y PAND2X1_140/Y 0.03fF
C39777 POR2X1_383/A POR2X1_343/B 0.03fF
C39778 POR2X1_96/A POR2X1_760/A 0.50fF
C39779 PAND2X1_444/m4_208_n4# PAND2X1_727/m4_208_n4# 0.05fF
C39780 PAND2X1_193/Y POR2X1_591/Y 0.01fF
C39781 POR2X1_685/CTRL2 POR2X1_452/Y 0.01fF
C39782 POR2X1_323/a_16_28# POR2X1_20/B 0.02fF
C39783 POR2X1_416/B PAND2X1_308/Y 0.03fF
C39784 POR2X1_150/Y PAND2X1_795/B 0.03fF
C39785 PAND2X1_273/CTRL POR2X1_814/A 0.01fF
C39786 POR2X1_376/B PAND2X1_340/B 0.02fF
C39787 PAND2X1_48/A PAND2X1_136/O 0.04fF
C39788 POR2X1_49/Y PAND2X1_477/O 0.16fF
C39789 POR2X1_327/Y POR2X1_711/Y 0.10fF
C39790 PAND2X1_405/CTRL2 POR2X1_38/Y 0.00fF
C39791 PAND2X1_847/CTRL POR2X1_394/A 0.01fF
C39792 POR2X1_655/A PAND2X1_90/Y 0.00fF
C39793 POR2X1_273/Y PAND2X1_717/A 0.03fF
C39794 POR2X1_8/Y POR2X1_8/CTRL2 0.01fF
C39795 INPUT_1 POR2X1_49/O 0.02fF
C39796 PAND2X1_6/Y PAND2X1_32/CTRL2 0.01fF
C39797 POR2X1_176/CTRL POR2X1_77/Y 0.01fF
C39798 POR2X1_9/Y POR2X1_245/CTRL 0.07fF
C39799 POR2X1_78/A POR2X1_264/CTRL2 0.02fF
C39800 PAND2X1_231/CTRL POR2X1_263/Y 0.01fF
C39801 POR2X1_76/Y POR2X1_341/A 0.19fF
C39802 POR2X1_97/A PAND2X1_41/B 0.03fF
C39803 PAND2X1_217/O PAND2X1_364/B 0.05fF
C39804 POR2X1_681/Y INPUT_0 0.05fF
C39805 PAND2X1_839/CTRL2 POR2X1_20/B 0.01fF
C39806 POR2X1_271/Y POR2X1_102/Y 0.03fF
C39807 PAND2X1_217/B POR2X1_32/A 0.10fF
C39808 PAND2X1_20/A POR2X1_638/A 0.02fF
C39809 POR2X1_423/CTRL2 POR2X1_423/Y 0.01fF
C39810 PAND2X1_644/CTRL2 POR2X1_597/Y 0.03fF
C39811 POR2X1_296/B POR2X1_355/A 0.00fF
C39812 POR2X1_263/Y POR2X1_230/O 0.00fF
C39813 POR2X1_33/A PAND2X1_14/CTRL 0.00fF
C39814 POR2X1_481/Y POR2X1_20/B 0.17fF
C39815 POR2X1_78/A POR2X1_734/A 0.07fF
C39816 PAND2X1_392/O POR2X1_5/Y 0.36fF
C39817 POR2X1_564/Y POR2X1_319/A 0.03fF
C39818 PAND2X1_20/A POR2X1_94/A 0.22fF
C39819 POR2X1_341/A POR2X1_740/Y 0.10fF
C39820 POR2X1_834/Y POR2X1_661/A 0.10fF
C39821 POR2X1_567/B VDD 6.63fF
C39822 PAND2X1_408/O PAND2X1_408/Y 0.00fF
C39823 POR2X1_41/B POR2X1_265/CTRL 0.00fF
C39824 POR2X1_356/A POR2X1_446/CTRL 0.31fF
C39825 POR2X1_356/A POR2X1_148/O 0.06fF
C39826 POR2X1_661/O POR2X1_78/A 0.01fF
C39827 POR2X1_83/B POR2X1_677/O 0.15fF
C39828 POR2X1_136/Y PAND2X1_717/A 0.03fF
C39829 POR2X1_458/Y PAND2X1_368/CTRL2 0.05fF
C39830 PAND2X1_631/CTRL POR2X1_20/B 0.01fF
C39831 POR2X1_385/Y POR2X1_331/O 0.04fF
C39832 POR2X1_864/A PAND2X1_69/A 0.03fF
C39833 POR2X1_267/B POR2X1_267/A 0.02fF
C39834 POR2X1_54/Y PAND2X1_283/CTRL2 0.03fF
C39835 POR2X1_376/B POR2X1_102/Y 0.52fF
C39836 POR2X1_260/B POR2X1_783/B 0.02fF
C39837 POR2X1_244/B POR2X1_66/A 0.03fF
C39838 PAND2X1_124/Y PAND2X1_364/B 0.03fF
C39839 PAND2X1_492/CTRL2 POR2X1_78/A 0.01fF
C39840 PAND2X1_479/A D_INPUT_0 0.03fF
C39841 POR2X1_542/B POR2X1_556/A 0.03fF
C39842 POR2X1_49/Y POR2X1_40/Y 0.49fF
C39843 POR2X1_32/A VDD 5.03fF
C39844 POR2X1_485/Y POR2X1_526/Y 0.06fF
C39845 PAND2X1_93/B PAND2X1_144/CTRL2 0.03fF
C39846 POR2X1_760/A POR2X1_7/A 0.03fF
C39847 PAND2X1_497/O POR2X1_294/B 0.22fF
C39848 POR2X1_83/B POR2X1_701/Y 0.01fF
C39849 POR2X1_814/B POR2X1_94/A 0.12fF
C39850 POR2X1_376/B PAND2X1_436/A 0.10fF
C39851 PAND2X1_416/O POR2X1_816/A 0.01fF
C39852 POR2X1_43/B POR2X1_827/Y 0.01fF
C39853 POR2X1_356/A POR2X1_220/B 0.07fF
C39854 PAND2X1_6/Y POR2X1_808/CTRL 0.01fF
C39855 POR2X1_805/O POR2X1_805/A 0.07fF
C39856 POR2X1_348/A POR2X1_814/B 0.02fF
C39857 POR2X1_287/B POR2X1_389/Y 0.03fF
C39858 POR2X1_416/B POR2X1_77/Y 0.15fF
C39859 POR2X1_824/Y POR2X1_20/B 0.00fF
C39860 POR2X1_266/m4_208_n4# POR2X1_294/B 0.06fF
C39861 POR2X1_650/A PAND2X1_41/B 0.05fF
C39862 D_INPUT_3 POR2X1_263/a_76_344# 0.04fF
C39863 POR2X1_49/Y PAND2X1_849/O 0.17fF
C39864 POR2X1_48/A PAND2X1_552/B 0.03fF
C39865 POR2X1_846/A POR2X1_129/Y 0.00fF
C39866 PAND2X1_76/Y POR2X1_423/Y 0.03fF
C39867 PAND2X1_487/CTRL PAND2X1_69/A 0.01fF
C39868 PAND2X1_65/B POR2X1_461/CTRL2 0.03fF
C39869 POR2X1_308/O POR2X1_794/B 0.01fF
C39870 PAND2X1_423/O POR2X1_807/A 0.02fF
C39871 PAND2X1_706/O PAND2X1_713/B 0.01fF
C39872 POR2X1_78/B POR2X1_200/O 0.02fF
C39873 POR2X1_389/A PAND2X1_39/B 0.03fF
C39874 PAND2X1_286/O PAND2X1_805/A 0.06fF
C39875 POR2X1_102/Y PAND2X1_598/O 0.05fF
C39876 POR2X1_614/A POR2X1_796/Y 0.03fF
C39877 POR2X1_311/Y POR2X1_96/A 0.09fF
C39878 POR2X1_417/Y VDD 0.43fF
C39879 POR2X1_419/Y VDD 0.18fF
C39880 POR2X1_244/CTRL2 POR2X1_243/Y 0.04fF
C39881 POR2X1_20/B POR2X1_751/a_16_28# 0.03fF
C39882 D_INPUT_3 POR2X1_54/Y 0.03fF
C39883 POR2X1_13/A PAND2X1_244/O 0.06fF
C39884 POR2X1_590/A PAND2X1_152/O 0.08fF
C39885 PAND2X1_93/B POR2X1_786/Y 0.07fF
C39886 PAND2X1_781/Y VDD 0.13fF
C39887 POR2X1_48/A PAND2X1_705/O 0.04fF
C39888 POR2X1_3/A PAND2X1_12/CTRL 0.18fF
C39889 POR2X1_83/B PAND2X1_364/B 0.19fF
C39890 POR2X1_52/A POR2X1_102/Y 5.51fF
C39891 PAND2X1_866/A GATE_741 0.03fF
C39892 PAND2X1_48/B POR2X1_590/A 0.35fF
C39893 POR2X1_645/CTRL2 POR2X1_718/A 0.01fF
C39894 PAND2X1_9/Y PAND2X1_63/B 0.01fF
C39895 POR2X1_432/CTRL2 PAND2X1_658/B 0.20fF
C39896 POR2X1_624/Y PAND2X1_60/B 0.31fF
C39897 POR2X1_391/A VDD 0.22fF
C39898 POR2X1_829/A PAND2X1_200/O 0.00fF
C39899 PAND2X1_212/CTRL POR2X1_142/Y 0.00fF
C39900 POR2X1_567/B PAND2X1_32/B 0.05fF
C39901 POR2X1_102/Y PAND2X1_398/CTRL2 0.01fF
C39902 PAND2X1_93/B POR2X1_788/B 0.23fF
C39903 POR2X1_250/Y PAND2X1_360/Y 0.02fF
C39904 POR2X1_556/A POR2X1_218/a_16_28# 0.02fF
C39905 PAND2X1_640/B POR2X1_73/Y 0.07fF
C39906 POR2X1_13/CTRL POR2X1_595/Y 0.00fF
C39907 POR2X1_60/A PAND2X1_254/O 0.17fF
C39908 POR2X1_541/B POR2X1_456/B 0.00fF
C39909 POR2X1_284/CTRL POR2X1_330/Y 0.00fF
C39910 POR2X1_260/B POR2X1_140/a_16_28# 0.02fF
C39911 POR2X1_852/B POR2X1_220/Y 0.07fF
C39912 POR2X1_23/a_16_28# POR2X1_42/Y 0.02fF
C39913 POR2X1_413/A POR2X1_413/a_16_28# 0.03fF
C39914 POR2X1_383/A POR2X1_643/Y 0.14fF
C39915 POR2X1_669/B PAND2X1_6/A 0.31fF
C39916 PAND2X1_553/B POR2X1_40/Y 0.58fF
C39917 POR2X1_298/Y PAND2X1_302/a_76_28# 0.02fF
C39918 POR2X1_330/Y PAND2X1_369/CTRL2 0.15fF
C39919 POR2X1_262/O POR2X1_40/Y 0.01fF
C39920 POR2X1_315/Y PAND2X1_469/CTRL 0.06fF
C39921 POR2X1_43/B POR2X1_516/Y 0.03fF
C39922 POR2X1_121/A PAND2X1_58/A 0.02fF
C39923 PAND2X1_94/A POR2X1_473/CTRL 0.01fF
C39924 PAND2X1_793/Y PAND2X1_474/A 0.00fF
C39925 PAND2X1_41/B POR2X1_208/CTRL 0.01fF
C39926 POR2X1_734/A PAND2X1_132/CTRL 0.27fF
C39927 POR2X1_708/O PAND2X1_65/B 0.01fF
C39928 PAND2X1_741/B VDD 0.26fF
C39929 PAND2X1_73/Y POR2X1_804/A 0.05fF
C39930 POR2X1_78/B VDD 5.35fF
C39931 PAND2X1_859/B POR2X1_60/Y 0.01fF
C39932 POR2X1_96/A POR2X1_485/CTRL2 0.00fF
C39933 POR2X1_205/CTRL2 POR2X1_330/Y 0.01fF
C39934 POR2X1_330/Y POR2X1_363/CTRL 0.00fF
C39935 POR2X1_220/B POR2X1_220/A 0.03fF
C39936 POR2X1_468/a_56_344# PAND2X1_41/B 0.00fF
C39937 POR2X1_366/Y PAND2X1_41/B 0.07fF
C39938 PAND2X1_41/B POR2X1_294/B 0.22fF
C39939 PAND2X1_417/a_76_28# POR2X1_186/B 0.02fF
C39940 POR2X1_48/A POR2X1_416/CTRL2 0.03fF
C39941 PAND2X1_431/a_76_28# PAND2X1_60/B 0.01fF
C39942 POR2X1_360/A PAND2X1_85/Y 1.28fF
C39943 POR2X1_13/A POR2X1_481/A 0.02fF
C39944 POR2X1_251/Y PAND2X1_347/Y 0.00fF
C39945 PAND2X1_565/CTRL POR2X1_40/Y 0.01fF
C39946 POR2X1_624/B POR2X1_4/Y 0.10fF
C39947 POR2X1_811/B POR2X1_407/Y 0.03fF
C39948 PAND2X1_217/B POR2X1_184/Y 0.05fF
C39949 PAND2X1_35/Y VDD 0.00fF
C39950 POR2X1_333/A POR2X1_775/a_76_344# 0.02fF
C39951 POR2X1_334/Y PAND2X1_39/B 0.03fF
C39952 POR2X1_389/A POR2X1_805/Y 0.01fF
C39953 PAND2X1_390/Y POR2X1_56/Y 0.03fF
C39954 POR2X1_130/a_16_28# POR2X1_318/A 0.07fF
C39955 POR2X1_236/Y POR2X1_531/O 0.18fF
C39956 POR2X1_186/Y POR2X1_782/A 0.05fF
C39957 POR2X1_49/Y PAND2X1_848/B 0.03fF
C39958 PAND2X1_115/O PAND2X1_787/Y 0.10fF
C39959 POR2X1_740/CTRL2 POR2X1_740/Y 0.00fF
C39960 POR2X1_865/B POR2X1_474/CTRL 0.00fF
C39961 POR2X1_483/A POR2X1_833/CTRL2 0.01fF
C39962 POR2X1_57/CTRL VDD 0.00fF
C39963 POR2X1_389/A PAND2X1_20/A 0.20fF
C39964 POR2X1_41/B PAND2X1_738/Y 0.10fF
C39965 POR2X1_355/B POR2X1_192/Y 0.37fF
C39966 POR2X1_16/A PAND2X1_644/Y 0.03fF
C39967 PAND2X1_642/CTRL2 POR2X1_48/A 0.03fF
C39968 POR2X1_141/CTRL POR2X1_514/Y 0.01fF
C39969 PAND2X1_592/Y PAND2X1_362/B 0.05fF
C39970 POR2X1_378/Y PAND2X1_459/Y 0.01fF
C39971 POR2X1_304/a_16_28# POR2X1_56/B 0.01fF
C39972 PAND2X1_17/a_76_28# INPUT_7 0.01fF
C39973 POR2X1_813/Y POR2X1_32/A 0.01fF
C39974 PAND2X1_459/Y POR2X1_7/B 0.00fF
C39975 POR2X1_529/CTRL VDD 0.00fF
C39976 PAND2X1_249/a_16_344# POR2X1_38/Y 0.04fF
C39977 POR2X1_391/A PAND2X1_32/B 0.02fF
C39978 PAND2X1_414/CTRL POR2X1_39/B 0.01fF
C39979 PAND2X1_859/A PAND2X1_509/CTRL2 0.01fF
C39980 PAND2X1_96/B POR2X1_186/Y 0.08fF
C39981 POR2X1_777/B POR2X1_458/B 0.03fF
C39982 POR2X1_78/B POR2X1_741/Y 0.08fF
C39983 POR2X1_97/A POR2X1_502/CTRL 0.06fF
C39984 POR2X1_566/A POR2X1_555/m4_208_n4# 0.06fF
C39985 POR2X1_189/Y VDD 0.00fF
C39986 INPUT_4 POR2X1_7/B 0.10fF
C39987 PAND2X1_859/A POR2X1_38/Y 0.01fF
C39988 POR2X1_51/A POR2X1_64/a_16_28# 0.07fF
C39989 POR2X1_65/A PAND2X1_341/A 0.03fF
C39990 POR2X1_403/a_56_344# PAND2X1_69/A 0.00fF
C39991 POR2X1_78/B PAND2X1_81/B 0.02fF
C39992 POR2X1_518/Y POR2X1_236/Y 0.09fF
C39993 POR2X1_72/B POR2X1_511/O 0.01fF
C39994 PAND2X1_620/Y POR2X1_93/A 5.53fF
C39995 POR2X1_362/B PAND2X1_69/A 0.03fF
C39996 PAND2X1_472/A POR2X1_236/Y 0.03fF
C39997 POR2X1_86/Y PAND2X1_206/B 0.07fF
C39998 POR2X1_669/B POR2X1_523/CTRL2 0.04fF
C39999 POR2X1_724/O POR2X1_732/B 0.01fF
C40000 PAND2X1_351/O POR2X1_293/Y 0.01fF
C40001 POR2X1_184/Y VDD 1.12fF
C40002 POR2X1_244/B POR2X1_222/Y 0.03fF
C40003 POR2X1_375/Y POR2X1_584/Y 0.09fF
C40004 POR2X1_48/A PAND2X1_713/O 0.03fF
C40005 POR2X1_65/A POR2X1_93/A 0.02fF
C40006 PAND2X1_849/B POR2X1_83/B 0.01fF
C40007 PAND2X1_115/B POR2X1_7/B 0.01fF
C40008 POR2X1_389/A POR2X1_814/B 0.06fF
C40009 POR2X1_828/Y POR2X1_686/CTRL 0.01fF
C40010 POR2X1_59/O POR2X1_32/A 0.01fF
C40011 POR2X1_72/B PAND2X1_656/A 0.06fF
C40012 PAND2X1_41/B PAND2X1_111/B 0.03fF
C40013 POR2X1_800/A POR2X1_783/A 0.00fF
C40014 POR2X1_400/A POR2X1_208/Y 0.07fF
C40015 POR2X1_78/B PAND2X1_125/a_76_28# 0.03fF
C40016 POR2X1_344/A POR2X1_68/A 0.03fF
C40017 POR2X1_121/B POR2X1_260/A 0.03fF
C40018 PAND2X1_65/B PAND2X1_518/a_16_344# 0.02fF
C40019 PAND2X1_651/Y VDD 6.24fF
C40020 POR2X1_632/A POR2X1_532/A 0.00fF
C40021 POR2X1_78/B PAND2X1_32/B 0.28fF
C40022 POR2X1_537/Y POR2X1_851/A 0.20fF
C40023 PAND2X1_695/O POR2X1_407/Y 0.02fF
C40024 PAND2X1_94/A POR2X1_634/A 0.10fF
C40025 PAND2X1_658/A POR2X1_7/B 0.01fF
C40026 POR2X1_102/Y PAND2X1_508/a_16_344# 0.00fF
C40027 POR2X1_614/A POR2X1_728/B 0.01fF
C40028 POR2X1_66/B POR2X1_456/B 0.06fF
C40029 D_GATE_741 POR2X1_776/B 0.07fF
C40030 POR2X1_507/CTRL POR2X1_355/A 0.01fF
C40031 POR2X1_66/A POR2X1_722/CTRL 0.01fF
C40032 POR2X1_789/A POR2X1_790/O 0.09fF
C40033 POR2X1_807/A POR2X1_590/CTRL2 0.01fF
C40034 POR2X1_83/A PAND2X1_243/B 1.24fF
C40035 POR2X1_65/A PAND2X1_559/CTRL2 0.01fF
C40036 PAND2X1_57/B POR2X1_112/Y 14.52fF
C40037 POR2X1_537/Y POR2X1_66/A 0.12fF
C40038 PAND2X1_844/B VDD 0.03fF
C40039 D_INPUT_3 PAND2X1_14/O 0.01fF
C40040 POR2X1_335/A PAND2X1_23/Y 0.03fF
C40041 PAND2X1_65/B POR2X1_222/A 0.03fF
C40042 POR2X1_566/A POR2X1_447/CTRL 0.14fF
C40043 POR2X1_250/A PAND2X1_537/CTRL2 0.01fF
C40044 POR2X1_188/A POR2X1_456/B 0.00fF
C40045 POR2X1_13/A PAND2X1_645/B 0.01fF
C40046 PAND2X1_347/Y PAND2X1_568/B 0.45fF
C40047 POR2X1_447/B POR2X1_836/O 0.16fF
C40048 POR2X1_508/B POR2X1_836/CTRL 0.00fF
C40049 PAND2X1_58/A POR2X1_720/CTRL 0.00fF
C40050 POR2X1_41/O POR2X1_40/Y 0.06fF
C40051 INPUT_1 PAND2X1_859/A 0.03fF
C40052 POR2X1_334/Y PAND2X1_20/A 0.02fF
C40053 POR2X1_96/A POR2X1_38/Y 1.82fF
C40054 POR2X1_693/a_16_28# PAND2X1_565/A 0.04fF
C40055 PAND2X1_652/A PAND2X1_798/B 0.44fF
C40056 POR2X1_251/A PAND2X1_348/A 0.03fF
C40057 POR2X1_65/A PAND2X1_545/Y 0.04fF
C40058 POR2X1_13/A INPUT_6 0.10fF
C40059 POR2X1_7/B POR2X1_73/Y 0.06fF
C40060 PAND2X1_535/CTRL VDD 0.00fF
C40061 POR2X1_273/O POR2X1_39/B 0.01fF
C40062 PAND2X1_845/O POR2X1_55/Y 0.13fF
C40063 POR2X1_861/a_16_28# POR2X1_572/B 0.03fF
C40064 PAND2X1_119/CTRL2 POR2X1_294/B 0.16fF
C40065 POR2X1_391/CTRL VDD 0.00fF
C40066 POR2X1_407/Y POR2X1_783/B 0.02fF
C40067 POR2X1_119/Y POR2X1_669/B 0.17fF
C40068 PAND2X1_563/O PAND2X1_566/Y 0.15fF
C40069 PAND2X1_139/B POR2X1_283/A 0.03fF
C40070 PAND2X1_350/O POR2X1_88/Y 0.17fF
C40071 POR2X1_38/Y POR2X1_406/CTRL 0.01fF
C40072 PAND2X1_307/O POR2X1_153/Y 0.07fF
C40073 VDD POR2X1_503/Y 0.03fF
C40074 PAND2X1_65/B PAND2X1_103/O 0.01fF
C40075 POR2X1_140/B POR2X1_574/O 0.00fF
C40076 POR2X1_36/B INPUT_5 0.19fF
C40077 POR2X1_54/Y PAND2X1_52/B 0.03fF
C40078 POR2X1_447/B PAND2X1_39/O 0.09fF
C40079 POR2X1_563/CTRL POR2X1_456/B 0.07fF
C40080 POR2X1_109/CTRL POR2X1_77/Y 0.01fF
C40081 VDD POR2X1_141/A 0.00fF
C40082 POR2X1_515/m4_208_n4# PAND2X1_60/B 0.07fF
C40083 PAND2X1_453/CTRL2 PAND2X1_241/Y 0.01fF
C40084 POR2X1_668/a_76_344# POR2X1_260/A 0.01fF
C40085 PAND2X1_219/A PAND2X1_737/CTRL2 0.03fF
C40086 PAND2X1_530/a_16_344# PAND2X1_32/B 0.02fF
C40087 POR2X1_460/O PAND2X1_32/B 0.18fF
C40088 POR2X1_808/CTRL PAND2X1_52/B 0.01fF
C40089 PAND2X1_94/A POR2X1_130/A 0.07fF
C40090 POR2X1_165/Y POR2X1_376/B 0.02fF
C40091 POR2X1_13/A POR2X1_521/Y 0.02fF
C40092 POR2X1_334/Y POR2X1_814/B 1.70fF
C40093 POR2X1_57/A POR2X1_399/A 0.01fF
C40094 POR2X1_813/Y PAND2X1_35/Y 0.02fF
C40095 POR2X1_16/A PAND2X1_556/B 0.03fF
C40096 POR2X1_366/Y POR2X1_228/Y 0.03fF
C40097 POR2X1_294/B POR2X1_228/Y 0.10fF
C40098 POR2X1_22/A POR2X1_3/a_56_344# 0.00fF
C40099 POR2X1_192/Y PAND2X1_315/a_76_28# 0.03fF
C40100 PAND2X1_725/B POR2X1_394/A 0.15fF
C40101 PAND2X1_536/CTRL2 PAND2X1_60/B 0.00fF
C40102 POR2X1_99/B POR2X1_244/CTRL 0.00fF
C40103 POR2X1_68/A POR2X1_844/CTRL 0.01fF
C40104 POR2X1_516/a_76_344# PAND2X1_651/Y 0.10fF
C40105 POR2X1_317/CTRL2 POR2X1_854/B 0.17fF
C40106 PAND2X1_477/B POR2X1_73/Y 0.03fF
C40107 POR2X1_550/A POR2X1_294/B 0.00fF
C40108 POR2X1_52/A POR2X1_92/m4_208_n4# 0.12fF
C40109 PAND2X1_152/a_76_28# PAND2X1_60/B 0.01fF
C40110 POR2X1_366/Y POR2X1_704/O 0.04fF
C40111 PAND2X1_216/B POR2X1_13/A 0.03fF
C40112 POR2X1_96/A INPUT_1 0.09fF
C40113 POR2X1_5/Y POR2X1_6/a_16_28# 0.02fF
C40114 POR2X1_573/A POR2X1_576/Y 0.02fF
C40115 PAND2X1_631/A POR2X1_72/B 0.03fF
C40116 POR2X1_52/A PAND2X1_160/O 0.01fF
C40117 POR2X1_163/A PAND2X1_160/CTRL 0.04fF
C40118 POR2X1_163/a_16_28# POR2X1_394/A 0.03fF
C40119 POR2X1_96/A PAND2X1_802/B 0.03fF
C40120 POR2X1_677/Y POR2X1_411/B 0.02fF
C40121 POR2X1_567/A PAND2X1_41/B 0.05fF
C40122 PAND2X1_643/Y PAND2X1_645/B 0.07fF
C40123 POR2X1_196/Y PAND2X1_88/Y 0.02fF
C40124 PAND2X1_798/B POR2X1_437/CTRL2 0.03fF
C40125 POR2X1_68/A POR2X1_845/CTRL 0.00fF
C40126 POR2X1_57/O PAND2X1_737/B 0.01fF
C40127 PAND2X1_72/CTRL PAND2X1_111/B 0.04fF
C40128 PAND2X1_809/A PAND2X1_539/Y 0.23fF
C40129 PAND2X1_23/Y POR2X1_249/Y 0.00fF
C40130 POR2X1_9/Y POR2X1_411/B 0.13fF
C40131 PAND2X1_137/Y POR2X1_103/CTRL2 0.01fF
C40132 POR2X1_332/B POR2X1_715/A 0.02fF
C40133 POR2X1_5/Y POR2X1_7/Y 0.02fF
C40134 POR2X1_180/O VDD 0.00fF
C40135 POR2X1_276/A POR2X1_515/Y 0.12fF
C40136 POR2X1_96/A POR2X1_153/Y 0.18fF
C40137 POR2X1_40/Y PAND2X1_169/CTRL 0.01fF
C40138 POR2X1_16/A POR2X1_488/Y 0.05fF
C40139 POR2X1_863/CTRL POR2X1_260/A 0.01fF
C40140 POR2X1_356/CTRL POR2X1_356/B 0.00fF
C40141 POR2X1_572/m4_208_n4# POR2X1_260/A 0.08fF
C40142 POR2X1_123/A PAND2X1_518/CTRL2 0.01fF
C40143 PAND2X1_835/Y PAND2X1_656/A 0.03fF
C40144 VDD POR2X1_294/A 5.67fF
C40145 POR2X1_748/A POR2X1_39/B 0.09fF
C40146 POR2X1_567/A POR2X1_456/m4_208_n4# 0.03fF
C40147 PAND2X1_205/B PAND2X1_853/B 0.03fF
C40148 POR2X1_153/O POR2X1_7/B 0.01fF
C40149 POR2X1_508/A PAND2X1_627/O 0.03fF
C40150 POR2X1_383/A PAND2X1_63/Y 0.32fF
C40151 POR2X1_391/CTRL PAND2X1_32/B 0.01fF
C40152 INPUT_0 PAND2X1_716/B 0.07fF
C40153 POR2X1_65/A PAND2X1_169/CTRL2 0.03fF
C40154 POR2X1_16/A POR2X1_599/A 0.01fF
C40155 PAND2X1_56/Y POR2X1_260/A 0.06fF
C40156 POR2X1_790/A POR2X1_750/Y 0.01fF
C40157 POR2X1_388/CTRL2 POR2X1_703/A 0.01fF
C40158 POR2X1_38/Y POR2X1_7/A 0.10fF
C40159 PAND2X1_94/A POR2X1_844/B 0.03fF
C40160 POR2X1_540/CTRL2 POR2X1_181/B 0.00fF
C40161 PAND2X1_58/A POR2X1_717/B 0.45fF
C40162 POR2X1_327/Y POR2X1_733/A 0.13fF
C40163 PAND2X1_596/CTRL2 POR2X1_761/A 0.01fF
C40164 PAND2X1_860/A D_INPUT_0 0.03fF
C40165 POR2X1_130/A PAND2X1_136/CTRL2 0.02fF
C40166 POR2X1_390/B POR2X1_840/B 0.05fF
C40167 POR2X1_57/a_16_28# POR2X1_394/A 0.02fF
C40168 POR2X1_190/Y POR2X1_188/Y 0.13fF
C40169 POR2X1_45/Y POR2X1_129/Y 0.03fF
C40170 PAND2X1_187/CTRL2 POR2X1_568/Y 0.34fF
C40171 PAND2X1_56/Y PAND2X1_142/O 0.02fF
C40172 INPUT_6 POR2X1_1/a_76_344# 0.01fF
C40173 POR2X1_462/O POR2X1_472/B 0.01fF
C40174 POR2X1_680/CTRL2 POR2X1_79/Y 0.01fF
C40175 PAND2X1_865/Y PAND2X1_793/Y 2.19fF
C40176 POR2X1_610/CTRL POR2X1_814/A 0.04fF
C40177 POR2X1_68/A POR2X1_370/O 0.02fF
C40178 PAND2X1_534/a_76_28# PAND2X1_60/B 0.01fF
C40179 PAND2X1_726/B POR2X1_526/Y 0.07fF
C40180 POR2X1_741/Y POR2X1_294/A 0.03fF
C40181 PAND2X1_342/O POR2X1_153/Y 0.17fF
C40182 PAND2X1_659/Y POR2X1_45/Y 0.03fF
C40183 PAND2X1_639/Y POR2X1_42/Y 0.02fF
C40184 POR2X1_530/O POR2X1_530/Y 0.02fF
C40185 POR2X1_841/B POR2X1_814/A 0.01fF
C40186 PAND2X1_725/A PAND2X1_725/a_56_28# 0.00fF
C40187 D_GATE_741 POR2X1_192/B 0.10fF
C40188 VDD POR2X1_387/CTRL 0.00fF
C40189 VDD PAND2X1_858/B 0.02fF
C40190 INPUT_1 POR2X1_7/A 19.54fF
C40191 PAND2X1_63/Y PAND2X1_71/Y 0.03fF
C40192 POR2X1_760/Y POR2X1_42/Y 0.04fF
C40193 PAND2X1_854/O PAND2X1_854/Y 0.00fF
C40194 POR2X1_537/O PAND2X1_60/B 0.01fF
C40195 PAND2X1_738/Y POR2X1_77/Y 0.05fF
C40196 POR2X1_383/A POR2X1_260/A 0.22fF
C40197 POR2X1_294/B PAND2X1_122/O 0.09fF
C40198 POR2X1_802/B POR2X1_532/O 0.03fF
C40199 POR2X1_294/A PAND2X1_32/B 0.21fF
C40200 POR2X1_457/B POR2X1_717/B 0.02fF
C40201 PAND2X1_6/Y POR2X1_4/Y 0.24fF
C40202 PAND2X1_193/Y POR2X1_72/B 0.00fF
C40203 PAND2X1_60/B POR2X1_186/B 0.15fF
C40204 POR2X1_677/Y POR2X1_271/Y 2.05fF
C40205 POR2X1_7/A POR2X1_153/Y 0.14fF
C40206 PAND2X1_5/CTRL2 POR2X1_4/Y 0.01fF
C40207 POR2X1_554/Y POR2X1_736/A 0.01fF
C40208 POR2X1_456/B PAND2X1_313/CTRL 0.01fF
C40209 PAND2X1_148/Y PAND2X1_797/Y 0.12fF
C40210 PAND2X1_798/B POR2X1_184/CTRL 0.01fF
C40211 POR2X1_245/Y PAND2X1_156/A 0.10fF
C40212 PAND2X1_82/O POR2X1_294/A 0.17fF
C40213 PAND2X1_309/CTRL2 POR2X1_717/B 0.01fF
C40214 POR2X1_737/CTRL POR2X1_186/B 0.09fF
C40215 POR2X1_81/CTRL PAND2X1_510/B 0.01fF
C40216 PAND2X1_222/B POR2X1_7/Y 0.05fF
C40217 PAND2X1_286/B POR2X1_282/Y 0.01fF
C40218 D_INPUT_3 POR2X1_4/Y 0.33fF
C40219 POR2X1_716/CTRL2 POR2X1_723/B 0.01fF
C40220 PAND2X1_497/CTRL2 POR2X1_624/Y 0.01fF
C40221 POR2X1_270/Y POR2X1_663/B 0.03fF
C40222 POR2X1_416/B POR2X1_426/CTRL2 0.00fF
C40223 POR2X1_158/CTRL2 POR2X1_425/Y 0.01fF
C40224 PAND2X1_618/O POR2X1_29/A 0.01fF
C40225 POR2X1_311/Y POR2X1_760/A 0.03fF
C40226 POR2X1_16/A POR2X1_599/O 0.04fF
C40227 PAND2X1_23/Y POR2X1_715/CTRL 0.00fF
C40228 POR2X1_54/Y POR2X1_126/a_16_28# 0.01fF
C40229 PAND2X1_69/A D_INPUT_4 0.03fF
C40230 POR2X1_376/B POR2X1_9/Y 0.19fF
C40231 POR2X1_730/Y POR2X1_326/A 0.03fF
C40232 POR2X1_532/A POR2X1_532/O 0.01fF
C40233 PAND2X1_824/B POR2X1_334/A 0.01fF
C40234 PAND2X1_674/CTRL PAND2X1_72/A 0.01fF
C40235 POR2X1_332/O POR2X1_186/B 0.06fF
C40236 PAND2X1_71/Y POR2X1_260/A 0.03fF
C40237 POR2X1_461/CTRL2 POR2X1_814/A 0.01fF
C40238 PAND2X1_93/B POR2X1_602/CTRL 0.01fF
C40239 PAND2X1_9/Y POR2X1_32/A 0.03fF
C40240 PAND2X1_672/O POR2X1_260/A 0.02fF
C40241 PAND2X1_29/CTRL PAND2X1_52/B 0.10fF
C40242 POR2X1_291/Y POR2X1_39/B 0.01fF
C40243 PAND2X1_813/O POR2X1_62/Y 0.05fF
C40244 POR2X1_532/A POR2X1_555/CTRL 0.01fF
C40245 PAND2X1_23/Y POR2X1_354/CTRL2 0.01fF
C40246 POR2X1_416/B POR2X1_258/a_56_344# 0.00fF
C40247 POR2X1_567/B PAND2X1_237/CTRL2 0.06fF
C40248 POR2X1_542/B POR2X1_325/B 0.06fF
C40249 PAND2X1_826/CTRL2 POR2X1_838/B 0.00fF
C40250 POR2X1_441/Y PAND2X1_169/Y 0.03fF
C40251 POR2X1_356/A PAND2X1_437/O 0.26fF
C40252 POR2X1_823/Y POR2X1_77/Y 0.01fF
C40253 POR2X1_68/B POR2X1_8/CTRL2 0.04fF
C40254 PAND2X1_864/B GATE_222 0.03fF
C40255 POR2X1_52/A POR2X1_9/Y 0.10fF
C40256 POR2X1_260/B POR2X1_296/B 0.12fF
C40257 POR2X1_519/CTRL POR2X1_39/B 0.01fF
C40258 POR2X1_88/CTRL2 POR2X1_14/Y 0.04fF
C40259 POR2X1_191/CTRL POR2X1_353/A 0.01fF
C40260 POR2X1_673/A POR2X1_624/B 0.03fF
C40261 POR2X1_533/Y POR2X1_534/Y 0.15fF
C40262 POR2X1_260/B POR2X1_605/O 0.01fF
C40263 POR2X1_442/a_16_28# POR2X1_40/Y 0.00fF
C40264 POR2X1_23/CTRL POR2X1_37/Y 0.01fF
C40265 POR2X1_16/CTRL POR2X1_73/Y 0.04fF
C40266 POR2X1_49/Y POR2X1_442/m4_208_n4# 0.15fF
C40267 POR2X1_116/A VDD 0.05fF
C40268 POR2X1_257/A POR2X1_5/Y 0.29fF
C40269 PAND2X1_487/CTRL2 POR2X1_287/B 0.01fF
C40270 POR2X1_78/B PAND2X1_9/Y 0.03fF
C40271 POR2X1_614/A PAND2X1_257/O 0.01fF
C40272 POR2X1_634/A POR2X1_637/CTRL2 0.08fF
C40273 POR2X1_48/A POR2X1_748/A 0.05fF
C40274 POR2X1_41/B POR2X1_263/CTRL2 0.00fF
C40275 POR2X1_632/B POR2X1_590/A 0.01fF
C40276 PAND2X1_6/Y POR2X1_458/Y 0.90fF
C40277 POR2X1_292/Y POR2X1_295/Y 0.03fF
C40278 POR2X1_286/B VDD 0.22fF
C40279 POR2X1_278/Y POR2X1_411/B 0.07fF
C40280 PAND2X1_93/B POR2X1_788/O 0.01fF
C40281 POR2X1_114/B POR2X1_814/A 0.06fF
C40282 POR2X1_98/a_16_28# PAND2X1_20/A 0.03fF
C40283 POR2X1_260/B PAND2X1_380/CTRL2 0.03fF
C40284 PAND2X1_9/Y PAND2X1_35/Y 0.00fF
C40285 POR2X1_445/CTRL2 POR2X1_341/A 0.04fF
C40286 PAND2X1_620/Y POR2X1_422/a_16_28# 0.03fF
C40287 POR2X1_447/B POR2X1_568/B 0.03fF
C40288 POR2X1_275/O POR2X1_275/A 0.02fF
C40289 POR2X1_850/B POR2X1_806/CTRL 0.01fF
C40290 POR2X1_631/O POR2X1_590/A 0.18fF
C40291 POR2X1_634/A PAND2X1_11/Y 0.23fF
C40292 POR2X1_329/A POR2X1_90/Y 0.24fF
C40293 POR2X1_41/B PAND2X1_838/B 0.03fF
C40294 POR2X1_760/A PAND2X1_218/A 0.03fF
C40295 PAND2X1_457/CTRL PAND2X1_464/B 0.02fF
C40296 PAND2X1_480/B PAND2X1_469/CTRL 0.17fF
C40297 POR2X1_49/Y PAND2X1_68/a_76_28# 0.01fF
C40298 POR2X1_814/A POR2X1_458/B 0.01fF
C40299 POR2X1_490/Y INPUT_0 0.02fF
C40300 POR2X1_63/Y POR2X1_55/Y 0.03fF
C40301 PAND2X1_206/B POR2X1_73/Y 0.03fF
C40302 PAND2X1_465/O POR2X1_83/B 0.07fF
C40303 POR2X1_78/A POR2X1_788/O 0.01fF
C40304 POR2X1_707/B POR2X1_707/A 0.00fF
C40305 PAND2X1_9/Y POR2X1_247/m4_208_n4# 0.15fF
C40306 POR2X1_66/CTRL PAND2X1_69/A 0.01fF
C40307 POR2X1_150/Y PAND2X1_357/Y 0.12fF
C40308 POR2X1_856/B PAND2X1_627/a_16_344# 0.02fF
C40309 PAND2X1_626/CTRL POR2X1_852/B 0.03fF
C40310 POR2X1_760/A POR2X1_38/Y 0.12fF
C40311 POR2X1_462/B POR2X1_859/CTRL2 0.01fF
C40312 POR2X1_20/Y POR2X1_20/B 0.00fF
C40313 POR2X1_83/B POR2X1_427/Y 0.24fF
C40314 POR2X1_218/Y POR2X1_217/O 0.03fF
C40315 POR2X1_4/Y PAND2X1_52/B 0.10fF
C40316 POR2X1_109/O POR2X1_46/Y 0.03fF
C40317 PAND2X1_600/a_16_344# POR2X1_130/A 0.06fF
C40318 POR2X1_814/A POR2X1_222/A 0.03fF
C40319 POR2X1_43/B POR2X1_628/Y 0.05fF
C40320 PAND2X1_206/A PAND2X1_101/O 0.02fF
C40321 POR2X1_23/Y PAND2X1_468/CTRL 0.01fF
C40322 PAND2X1_39/B POR2X1_218/A 0.02fF
C40323 PAND2X1_667/CTRL POR2X1_590/A 0.12fF
C40324 POR2X1_454/A POR2X1_294/B 0.01fF
C40325 POR2X1_466/A POR2X1_724/O 0.25fF
C40326 POR2X1_409/B PAND2X1_734/B 0.02fF
C40327 PAND2X1_651/Y PAND2X1_9/Y 0.08fF
C40328 INPUT_2 POR2X1_411/B 0.00fF
C40329 PAND2X1_139/O POR2X1_40/Y 0.04fF
C40330 PAND2X1_477/CTRL2 POR2X1_238/Y 0.01fF
C40331 POR2X1_186/Y POR2X1_355/A 0.04fF
C40332 PAND2X1_696/a_76_28# POR2X1_811/B 0.02fF
C40333 POR2X1_490/Y PAND2X1_218/CTRL 0.01fF
C40334 PAND2X1_244/B PAND2X1_206/B 2.27fF
C40335 POR2X1_558/O POR2X1_260/B 0.01fF
C40336 POR2X1_554/B POR2X1_510/Y 0.22fF
C40337 PAND2X1_841/CTRL POR2X1_23/Y 0.00fF
C40338 POR2X1_461/A PAND2X1_90/Y 0.01fF
C40339 POR2X1_814/A PAND2X1_103/O 0.04fF
C40340 INPUT_7 POR2X1_750/B 0.01fF
C40341 POR2X1_119/Y POR2X1_234/A 0.05fF
C40342 POR2X1_122/A POR2X1_40/Y 0.01fF
C40343 PAND2X1_65/B PAND2X1_46/CTRL 0.01fF
C40344 POR2X1_304/Y POR2X1_102/Y 0.09fF
C40345 D_INPUT_5 PAND2X1_752/Y 0.01fF
C40346 POR2X1_66/B PAND2X1_131/CTRL2 0.01fF
C40347 PAND2X1_265/O VDD 0.00fF
C40348 POR2X1_647/B POR2X1_865/CTRL 0.01fF
C40349 PAND2X1_48/B POR2X1_66/A 0.25fF
C40350 POR2X1_29/Y PAND2X1_35/A 0.02fF
C40351 POR2X1_260/B POR2X1_267/Y 0.01fF
C40352 POR2X1_220/Y PAND2X1_39/O 0.01fF
C40353 PAND2X1_862/B POR2X1_102/Y 0.03fF
C40354 POR2X1_638/A VDD 0.00fF
C40355 POR2X1_693/Y POR2X1_23/Y 0.03fF
C40356 POR2X1_49/Y POR2X1_5/Y 5.84fF
C40357 POR2X1_814/B POR2X1_475/A 7.42fF
C40358 POR2X1_753/Y POR2X1_7/B 3.03fF
C40359 POR2X1_822/O POR2X1_40/Y 0.02fF
C40360 POR2X1_78/B POR2X1_808/A 0.02fF
C40361 POR2X1_72/Y PAND2X1_657/CTRL2 0.01fF
C40362 POR2X1_862/Y PAND2X1_32/B 0.10fF
C40363 POR2X1_554/B POR2X1_276/Y 0.02fF
C40364 POR2X1_250/Y PAND2X1_343/a_16_344# 0.02fF
C40365 POR2X1_66/B PAND2X1_57/B 0.55fF
C40366 POR2X1_97/A POR2X1_350/CTRL2 0.10fF
C40367 POR2X1_94/A VDD 1.94fF
C40368 POR2X1_760/A PAND2X1_802/B 0.01fF
C40369 PAND2X1_731/B VDD 0.55fF
C40370 POR2X1_590/A POR2X1_717/Y 0.09fF
C40371 POR2X1_65/A PAND2X1_539/B 0.02fF
C40372 PAND2X1_55/Y POR2X1_296/B 1.62fF
C40373 POR2X1_362/B POR2X1_405/a_16_28# 0.03fF
C40374 PAND2X1_579/CTRL VDD 0.00fF
C40375 PAND2X1_810/B PAND2X1_539/Y 0.01fF
C40376 POR2X1_348/A VDD 0.00fF
C40377 PAND2X1_208/CTRL2 PAND2X1_35/Y 0.01fF
C40378 POR2X1_776/A POR2X1_566/B 0.12fF
C40379 POR2X1_415/A POR2X1_283/A 0.03fF
C40380 POR2X1_188/A PAND2X1_57/B 0.06fF
C40381 POR2X1_858/a_16_28# POR2X1_733/A 0.20fF
C40382 PAND2X1_803/A POR2X1_236/Y 0.06fF
C40383 PAND2X1_786/CTRL POR2X1_293/Y 0.05fF
C40384 POR2X1_32/A PAND2X1_717/O 0.01fF
C40385 PAND2X1_480/B POR2X1_423/Y 0.05fF
C40386 PAND2X1_205/Y INPUT_0 0.02fF
C40387 POR2X1_121/A POR2X1_608/Y 0.35fF
C40388 POR2X1_485/Y PAND2X1_726/B 0.07fF
C40389 POR2X1_16/A POR2X1_441/Y 0.05fF
C40390 POR2X1_750/B INPUT_4 0.10fF
C40391 POR2X1_788/Y POR2X1_296/B 0.04fF
C40392 POR2X1_263/Y PAND2X1_734/O 0.02fF
C40393 POR2X1_31/CTRL2 POR2X1_12/A 0.11fF
C40394 POR2X1_402/A POR2X1_296/B 0.09fF
C40395 POR2X1_579/Y POR2X1_330/Y 0.03fF
C40396 POR2X1_254/A POR2X1_785/A 0.03fF
C40397 PAND2X1_41/B PAND2X1_386/Y 0.03fF
C40398 PAND2X1_73/CTRL POR2X1_294/B 0.11fF
C40399 PAND2X1_70/CTRL VDD 0.00fF
C40400 POR2X1_110/Y POR2X1_329/A 0.10fF
C40401 POR2X1_687/A POR2X1_676/O 0.01fF
C40402 POR2X1_502/A POR2X1_830/A 0.01fF
C40403 PAND2X1_849/B PAND2X1_206/A 0.03fF
C40404 PAND2X1_115/CTRL2 PAND2X1_562/B 0.02fF
C40405 POR2X1_78/B POR2X1_403/A 0.01fF
C40406 POR2X1_122/CTRL2 POR2X1_411/B 0.01fF
C40407 POR2X1_814/A POR2X1_362/O 0.08fF
C40408 POR2X1_272/O POR2X1_42/Y 0.09fF
C40409 PAND2X1_390/Y POR2X1_42/Y 0.02fF
C40410 POR2X1_630/O POR2X1_510/Y 0.01fF
C40411 POR2X1_863/A POR2X1_181/Y 0.01fF
C40412 POR2X1_271/B POR2X1_129/Y 0.02fF
C40413 PAND2X1_73/Y POR2X1_570/B 0.03fF
C40414 POR2X1_267/A PAND2X1_767/CTRL 0.01fF
C40415 POR2X1_68/A PAND2X1_279/O -0.01fF
C40416 POR2X1_188/A POR2X1_285/A 0.01fF
C40417 POR2X1_68/A POR2X1_866/O 0.04fF
C40418 POR2X1_516/O POR2X1_60/A 0.18fF
C40419 POR2X1_52/A PAND2X1_736/CTRL2 0.00fF
C40420 POR2X1_43/B PAND2X1_556/a_76_28# 0.01fF
C40421 POR2X1_114/B POR2X1_405/CTRL2 0.01fF
C40422 PAND2X1_378/CTRL VDD 0.00fF
C40423 POR2X1_458/CTRL POR2X1_101/Y 0.07fF
C40424 POR2X1_130/A PAND2X1_56/CTRL2 0.01fF
C40425 PAND2X1_213/Y PAND2X1_220/A 0.00fF
C40426 POR2X1_383/A PAND2X1_65/O 0.04fF
C40427 PAND2X1_863/B PAND2X1_687/Y 0.01fF
C40428 POR2X1_294/CTRL POR2X1_507/A 0.04fF
C40429 POR2X1_264/a_16_28# POR2X1_294/B 0.03fF
C40430 POR2X1_435/Y POR2X1_794/O 0.05fF
C40431 PAND2X1_63/CTRL PAND2X1_63/B 0.01fF
C40432 POR2X1_569/CTRL POR2X1_853/A 0.01fF
C40433 PAND2X1_69/A POR2X1_720/a_16_28# 0.03fF
C40434 POR2X1_8/Y POR2X1_126/CTRL 0.01fF
C40435 PAND2X1_265/O PAND2X1_32/B 0.03fF
C40436 POR2X1_51/A VDD 0.13fF
C40437 POR2X1_23/Y PAND2X1_574/CTRL 0.03fF
C40438 POR2X1_251/A POR2X1_183/Y 0.04fF
C40439 POR2X1_60/A POR2X1_700/Y 0.03fF
C40440 POR2X1_13/A PAND2X1_768/CTRL2 0.00fF
C40441 POR2X1_614/A PAND2X1_677/O 0.04fF
C40442 POR2X1_614/A POR2X1_330/Y 0.06fF
C40443 PAND2X1_74/O POR2X1_702/A -0.00fF
C40444 POR2X1_14/Y POR2X1_750/CTRL2 0.10fF
C40445 POR2X1_476/Y POR2X1_294/B 0.03fF
C40446 POR2X1_12/A POR2X1_394/A 0.02fF
C40447 PAND2X1_92/CTRL INPUT_0 0.01fF
C40448 POR2X1_859/A PAND2X1_57/B 0.06fF
C40449 POR2X1_812/A POR2X1_532/A 0.01fF
C40450 POR2X1_175/A POR2X1_614/A 0.05fF
C40451 POR2X1_407/A PAND2X1_41/B 0.03fF
C40452 POR2X1_65/A PAND2X1_551/A 0.01fF
C40453 POR2X1_392/B POR2X1_391/Y 0.24fF
C40454 PAND2X1_437/O PAND2X1_72/A 0.02fF
C40455 PAND2X1_65/B POR2X1_732/B 0.03fF
C40456 POR2X1_558/B POR2X1_362/A 0.25fF
C40457 PAND2X1_653/Y POR2X1_40/Y 0.06fF
C40458 POR2X1_814/B POR2X1_218/A 0.12fF
C40459 PAND2X1_9/Y POR2X1_294/A 0.03fF
C40460 PAND2X1_652/Y VDD 0.12fF
C40461 POR2X1_464/CTRL PAND2X1_55/Y 0.00fF
C40462 POR2X1_94/A PAND2X1_32/B 0.03fF
C40463 PAND2X1_252/O POR2X1_750/B 0.02fF
C40464 POR2X1_19/a_76_344# POR2X1_4/Y 0.01fF
C40465 POR2X1_52/A POR2X1_278/Y 0.12fF
C40466 PAND2X1_798/B PAND2X1_76/Y 0.03fF
C40467 PAND2X1_6/Y PAND2X1_52/Y 0.04fF
C40468 POR2X1_848/A POR2X1_753/CTRL 0.04fF
C40469 POR2X1_51/A POR2X1_408/CTRL2 0.01fF
C40470 PAND2X1_852/A POR2X1_394/A 0.03fF
C40471 PAND2X1_828/O POR2X1_599/A 0.13fF
C40472 PAND2X1_785/Y POR2X1_7/B 0.00fF
C40473 PAND2X1_475/a_16_344# POR2X1_38/Y 0.02fF
C40474 POR2X1_654/B POR2X1_649/CTRL 0.03fF
C40475 PAND2X1_249/a_16_344# POR2X1_591/Y 0.01fF
C40476 PAND2X1_23/Y PAND2X1_293/CTRL 0.00fF
C40477 POR2X1_20/B PAND2X1_352/B 0.00fF
C40478 POR2X1_362/B POR2X1_723/B 0.06fF
C40479 POR2X1_508/B POR2X1_776/A 0.03fF
C40480 POR2X1_458/Y PAND2X1_52/B 0.03fF
C40481 POR2X1_121/B POR2X1_725/Y 0.64fF
C40482 POR2X1_566/A PAND2X1_441/CTRL 0.05fF
C40483 POR2X1_393/Y PAND2X1_656/A 0.01fF
C40484 PAND2X1_15/CTRL2 POR2X1_260/A 0.03fF
C40485 POR2X1_840/B POR2X1_274/Y 0.09fF
C40486 POR2X1_52/A POR2X1_829/A 0.04fF
C40487 PAND2X1_685/O INPUT_0 0.05fF
C40488 PAND2X1_218/a_16_344# PAND2X1_741/B 0.02fF
C40489 POR2X1_555/A PAND2X1_69/A 0.06fF
C40490 PAND2X1_844/CTRL2 D_INPUT_0 0.15fF
C40491 PAND2X1_860/A POR2X1_173/Y 0.01fF
C40492 POR2X1_65/A POR2X1_165/CTRL2 0.03fF
C40493 POR2X1_68/A PAND2X1_293/CTRL2 0.11fF
C40494 POR2X1_166/CTRL PAND2X1_714/A 0.01fF
C40495 PAND2X1_659/Y PAND2X1_205/CTRL2 0.01fF
C40496 PAND2X1_48/B PAND2X1_751/O 0.01fF
C40497 POR2X1_416/B PAND2X1_780/CTRL 0.03fF
C40498 POR2X1_78/A PAND2X1_528/a_16_344# 0.02fF
C40499 PAND2X1_813/CTRL2 POR2X1_78/A 0.03fF
C40500 POR2X1_272/CTRL PAND2X1_349/A 0.01fF
C40501 PAND2X1_48/B POR2X1_792/B 0.02fF
C40502 POR2X1_804/B VDD 0.03fF
C40503 PAND2X1_56/a_76_28# PAND2X1_55/Y 0.01fF
C40504 POR2X1_759/A POR2X1_236/Y 0.02fF
C40505 POR2X1_72/B PAND2X1_374/CTRL2 0.01fF
C40506 POR2X1_43/B PAND2X1_636/a_16_344# 0.02fF
C40507 POR2X1_65/A PAND2X1_338/B 0.03fF
C40508 PAND2X1_520/O POR2X1_518/Y 0.03fF
C40509 PAND2X1_520/CTRL PAND2X1_642/B 0.01fF
C40510 POR2X1_818/Y POR2X1_294/A 0.01fF
C40511 POR2X1_416/Y POR2X1_411/CTRL 0.01fF
C40512 POR2X1_303/O POR2X1_274/A 0.02fF
C40513 PAND2X1_594/CTRL POR2X1_151/Y 0.15fF
C40514 POR2X1_258/Y POR2X1_312/Y 0.10fF
C40515 PAND2X1_63/Y INPUT_0 0.13fF
C40516 POR2X1_537/Y POR2X1_858/CTRL2 0.01fF
C40517 POR2X1_323/a_16_28# POR2X1_73/Y 0.03fF
C40518 POR2X1_446/A POR2X1_568/B 0.02fF
C40519 POR2X1_68/A POR2X1_307/Y 0.05fF
C40520 PAND2X1_734/B POR2X1_229/CTRL2 0.01fF
C40521 PAND2X1_490/CTRL PAND2X1_57/B 0.01fF
C40522 POR2X1_833/O POR2X1_294/B 0.01fF
C40523 POR2X1_144/Y POR2X1_142/Y 0.01fF
C40524 POR2X1_41/B POR2X1_248/CTRL2 0.01fF
C40525 PAND2X1_48/B POR2X1_222/Y 0.03fF
C40526 POR2X1_234/CTRL POR2X1_293/Y 0.01fF
C40527 POR2X1_126/a_16_28# POR2X1_4/Y 0.02fF
C40528 PAND2X1_107/O POR2X1_640/Y 0.06fF
C40529 POR2X1_178/a_76_344# PAND2X1_738/Y 0.04fF
C40530 POR2X1_335/A POR2X1_733/A 0.03fF
C40531 POR2X1_198/CTRL2 POR2X1_68/A 0.01fF
C40532 POR2X1_389/A VDD 0.11fF
C40533 PAND2X1_20/A PAND2X1_586/CTRL2 0.00fF
C40534 POR2X1_16/A POR2X1_491/O 0.17fF
C40535 PAND2X1_6/Y POR2X1_84/CTRL2 0.00fF
C40536 PAND2X1_631/CTRL2 POR2X1_55/Y 0.03fF
C40537 PAND2X1_838/B POR2X1_77/Y 0.42fF
C40538 POR2X1_673/Y POR2X1_94/A 0.03fF
C40539 POR2X1_66/B POR2X1_259/B 0.03fF
C40540 PAND2X1_494/CTRL2 POR2X1_264/Y 0.01fF
C40541 POR2X1_72/CTRL2 POR2X1_23/Y 0.01fF
C40542 POR2X1_13/A POR2X1_597/CTRL2 0.01fF
C40543 PAND2X1_676/O PAND2X1_735/Y 0.09fF
C40544 POR2X1_220/Y PAND2X1_88/Y 0.03fF
C40545 PAND2X1_807/B PAND2X1_354/Y 0.01fF
C40546 PAND2X1_319/B PAND2X1_480/B 0.05fF
C40547 PAND2X1_562/B PAND2X1_348/O 0.10fF
C40548 POR2X1_707/O PAND2X1_41/B 0.01fF
C40549 POR2X1_302/A POR2X1_114/B 0.01fF
C40550 PAND2X1_523/O POR2X1_522/Y 0.01fF
C40551 PAND2X1_523/CTRL2 PAND2X1_844/B 0.01fF
C40552 POR2X1_140/B POR2X1_130/Y 0.04fF
C40553 POR2X1_43/B POR2X1_519/Y 0.01fF
C40554 INPUT_1 PAND2X1_42/O 0.02fF
C40555 POR2X1_130/A POR2X1_361/a_76_344# 0.02fF
C40556 PAND2X1_6/Y D_GATE_662 0.07fF
C40557 POR2X1_188/A PAND2X1_701/O 0.01fF
C40558 POR2X1_102/Y PAND2X1_716/B 0.06fF
C40559 PAND2X1_56/Y PAND2X1_111/a_16_344# 0.02fF
C40560 POR2X1_7/B PAND2X1_347/a_16_344# 0.02fF
C40561 POR2X1_404/Y PAND2X1_88/Y 0.03fF
C40562 POR2X1_750/B POR2X1_186/B 0.11fF
C40563 POR2X1_124/a_16_28# PAND2X1_32/B 0.02fF
C40564 PAND2X1_564/O POR2X1_765/Y 0.02fF
C40565 PAND2X1_48/B POR2X1_532/A 0.29fF
C40566 PAND2X1_684/CTRL2 PAND2X1_90/Y 0.05fF
C40567 PAND2X1_569/B PAND2X1_544/O 0.01fF
C40568 POR2X1_809/A POR2X1_866/a_56_344# 0.00fF
C40569 POR2X1_49/Y POR2X1_599/CTRL 0.01fF
C40570 PAND2X1_69/A PAND2X1_145/O 0.02fF
C40571 PAND2X1_7/m4_208_n4# POR2X1_222/Y 0.08fF
C40572 PAND2X1_445/O POR2X1_90/Y 0.02fF
C40573 POR2X1_730/Y POR2X1_480/A 0.07fF
C40574 POR2X1_66/A PAND2X1_529/CTRL2 0.03fF
C40575 POR2X1_555/A PAND2X1_824/B 0.07fF
C40576 POR2X1_188/A POR2X1_851/a_56_344# 0.00fF
C40577 POR2X1_68/A PAND2X1_72/O 0.02fF
C40578 POR2X1_78/B POR2X1_339/CTRL2 0.36fF
C40579 PAND2X1_832/O POR2X1_153/Y 0.17fF
C40580 POR2X1_65/A POR2X1_103/O 0.01fF
C40581 PAND2X1_360/CTRL POR2X1_385/Y 0.44fF
C40582 POR2X1_278/Y POR2X1_679/B 0.02fF
C40583 POR2X1_451/A POR2X1_635/CTRL 0.01fF
C40584 POR2X1_635/B POR2X1_635/O 0.01fF
C40585 POR2X1_62/Y PAND2X1_459/a_16_344# 0.02fF
C40586 POR2X1_263/Y POR2X1_39/B 0.05fF
C40587 PAND2X1_13/O POR2X1_186/B 0.02fF
C40588 POR2X1_750/B POR2X1_802/A 0.06fF
C40589 POR2X1_808/A POR2X1_294/A 0.06fF
C40590 POR2X1_213/O POR2X1_532/A 0.01fF
C40591 POR2X1_409/Y VDD 0.08fF
C40592 POR2X1_68/A POR2X1_68/B 10.11fF
C40593 POR2X1_853/A POR2X1_578/O 0.01fF
C40594 PAND2X1_169/Y PAND2X1_714/B 0.12fF
C40595 PAND2X1_613/a_16_344# PAND2X1_52/B 0.05fF
C40596 POR2X1_57/A POR2X1_83/A 0.02fF
C40597 PAND2X1_93/O PAND2X1_88/Y 0.02fF
C40598 POR2X1_517/CTRL POR2X1_83/B 0.01fF
C40599 POR2X1_311/CTRL POR2X1_7/B 0.01fF
C40600 POR2X1_394/A PAND2X1_738/a_16_344# 0.02fF
C40601 PAND2X1_691/Y PAND2X1_863/B 0.00fF
C40602 INPUT_0 POR2X1_260/A 0.16fF
C40603 POR2X1_550/A POR2X1_565/B 0.33fF
C40604 POR2X1_550/A POR2X1_546/B 0.01fF
C40605 PAND2X1_69/A POR2X1_705/O 0.01fF
C40606 D_INPUT_0 PAND2X1_339/O 0.08fF
C40607 POR2X1_7/B POR2X1_375/CTRL2 0.01fF
C40608 PAND2X1_251/O PAND2X1_52/B 0.01fF
C40609 POR2X1_193/Y POR2X1_228/O 0.08fF
C40610 POR2X1_72/B PAND2X1_199/CTRL 0.01fF
C40611 POR2X1_389/a_16_28# POR2X1_389/A 0.03fF
C40612 POR2X1_383/A PAND2X1_110/O 0.01fF
C40613 POR2X1_178/Y PAND2X1_553/B 0.18fF
C40614 POR2X1_857/B PAND2X1_503/CTRL2 0.03fF
C40615 PAND2X1_469/B POR2X1_387/Y 0.10fF
C40616 POR2X1_140/B POR2X1_228/Y 0.03fF
C40617 POR2X1_710/CTRL2 POR2X1_713/B 0.00fF
C40618 POR2X1_57/A POR2X1_90/Y 0.13fF
C40619 POR2X1_820/Y POR2X1_394/A 0.05fF
C40620 PAND2X1_90/A POR2X1_116/Y 0.05fF
C40621 POR2X1_334/Y VDD 0.00fF
C40622 POR2X1_796/a_16_28# POR2X1_783/Y -0.00fF
C40623 POR2X1_406/O PAND2X1_737/B 0.01fF
C40624 PAND2X1_56/Y POR2X1_725/Y 0.10fF
C40625 D_INPUT_3 D_INPUT_1 0.25fF
C40626 POR2X1_249/Y POR2X1_733/A 0.05fF
C40627 PAND2X1_830/Y PAND2X1_348/A 0.02fF
C40628 PAND2X1_484/O PAND2X1_57/B 0.09fF
C40629 POR2X1_614/A PAND2X1_158/CTRL 0.01fF
C40630 POR2X1_510/Y POR2X1_702/A 0.03fF
C40631 POR2X1_7/B PAND2X1_348/A 0.07fF
C40632 PAND2X1_723/Y POR2X1_7/Y 0.05fF
C40633 PAND2X1_810/a_76_28# POR2X1_7/B 0.01fF
C40634 PAND2X1_382/O POR2X1_816/A 0.01fF
C40635 POR2X1_516/O POR2X1_516/A 0.03fF
C40636 PAND2X1_547/O POR2X1_527/Y 0.02fF
C40637 POR2X1_403/A POR2X1_294/A 0.01fF
C40638 PAND2X1_79/Y PAND2X1_60/B 0.05fF
C40639 POR2X1_130/A POR2X1_561/Y 0.04fF
C40640 POR2X1_546/A POR2X1_550/B 0.00fF
C40641 POR2X1_411/B PAND2X1_269/CTRL 0.01fF
C40642 PAND2X1_390/Y POR2X1_589/a_76_344# 0.00fF
C40643 PAND2X1_55/Y POR2X1_590/Y 0.10fF
C40644 POR2X1_579/Y POR2X1_715/A 0.02fF
C40645 PAND2X1_6/Y PAND2X1_300/O 0.07fF
C40646 POR2X1_532/A PAND2X1_534/O 0.07fF
C40647 PAND2X1_649/A PAND2X1_688/CTRL 0.01fF
C40648 PAND2X1_139/CTRL PAND2X1_140/Y 0.01fF
C40649 PAND2X1_615/O PAND2X1_63/B 0.04fF
C40650 POR2X1_252/m4_208_n4# POR2X1_153/Y 0.03fF
C40651 INPUT_0 PAND2X1_517/CTRL2 0.06fF
C40652 POR2X1_832/A POR2X1_513/CTRL 0.05fF
C40653 PAND2X1_575/A POR2X1_394/A 0.15fF
C40654 PAND2X1_52/Y POR2X1_632/Y 0.03fF
C40655 POR2X1_54/Y POR2X1_848/O 0.01fF
C40656 POR2X1_580/a_16_28# POR2X1_191/Y 0.03fF
C40657 POR2X1_110/CTRL POR2X1_293/Y 0.01fF
C40658 POR2X1_450/B PAND2X1_72/A 0.00fF
C40659 POR2X1_54/Y PAND2X1_87/O 0.05fF
C40660 POR2X1_327/Y POR2X1_327/a_16_28# 0.02fF
C40661 POR2X1_215/A PAND2X1_88/Y 0.00fF
C40662 POR2X1_616/Y PAND2X1_621/Y 0.01fF
C40663 POR2X1_73/Y PAND2X1_840/m4_208_n4# 0.09fF
C40664 POR2X1_334/Y POR2X1_741/Y 0.07fF
C40665 POR2X1_609/Y PAND2X1_403/CTRL2 0.00fF
C40666 POR2X1_671/a_16_28# POR2X1_4/Y 0.03fF
C40667 PAND2X1_385/O PAND2X1_48/A 0.04fF
C40668 VDD POR2X1_343/CTRL -0.00fF
C40669 INPUT_1 POR2X1_38/Y 0.08fF
C40670 POR2X1_383/A POR2X1_725/Y 0.14fF
C40671 POR2X1_416/B POR2X1_106/Y 0.15fF
C40672 POR2X1_614/A POR2X1_715/A 0.02fF
C40673 PAND2X1_631/A POR2X1_7/B 0.03fF
C40674 PAND2X1_312/CTRL POR2X1_703/A 0.01fF
C40675 PAND2X1_671/a_76_28# INPUT_2 0.01fF
C40676 POR2X1_54/Y POR2X1_623/Y 0.08fF
C40677 POR2X1_57/A PAND2X1_732/A 1.48fF
C40678 POR2X1_780/A POR2X1_260/A 0.01fF
C40679 POR2X1_99/B POR2X1_294/B 0.03fF
C40680 PAND2X1_483/CTRL2 POR2X1_7/A 0.01fF
C40681 POR2X1_111/O POR2X1_111/Y 0.02fF
C40682 PAND2X1_484/CTRL PAND2X1_69/A 0.01fF
C40683 POR2X1_119/Y PAND2X1_466/O 0.16fF
C40684 PAND2X1_560/B POR2X1_73/Y 0.15fF
C40685 POR2X1_544/B POR2X1_540/A 0.42fF
C40686 POR2X1_548/CTRL PAND2X1_52/B 0.01fF
C40687 PAND2X1_501/CTRL2 PAND2X1_735/Y 0.05fF
C40688 POR2X1_38/Y POR2X1_153/Y 0.10fF
C40689 POR2X1_319/a_76_344# POR2X1_191/Y 0.01fF
C40690 POR2X1_416/B PAND2X1_580/B 0.03fF
C40691 POR2X1_570/Y POR2X1_854/B 0.05fF
C40692 POR2X1_561/Y POR2X1_844/B 0.00fF
C40693 POR2X1_108/a_16_28# PAND2X1_348/A 0.07fF
C40694 POR2X1_539/A POR2X1_675/Y 0.03fF
C40695 POR2X1_48/A POR2X1_600/CTRL 0.01fF
C40696 POR2X1_730/Y POR2X1_727/O 0.01fF
C40697 POR2X1_739/a_16_28# POR2X1_444/Y 0.03fF
C40698 PAND2X1_39/B PAND2X1_43/CTRL 0.01fF
C40699 POR2X1_290/CTRL2 POR2X1_234/A 0.01fF
C40700 POR2X1_57/A PAND2X1_360/Y 0.91fF
C40701 POR2X1_614/A POR2X1_337/Y 0.07fF
C40702 POR2X1_16/A PAND2X1_489/CTRL 0.06fF
C40703 POR2X1_147/CTRL2 POR2X1_435/Y 0.03fF
C40704 D_INPUT_6 PAND2X1_18/B 0.26fF
C40705 POR2X1_57/A PAND2X1_138/CTRL 0.01fF
C40706 PAND2X1_69/A PAND2X1_396/CTRL 0.08fF
C40707 POR2X1_539/A POR2X1_544/B 0.05fF
C40708 POR2X1_628/O POR2X1_39/B 0.02fF
C40709 POR2X1_57/A POR2X1_110/Y 0.08fF
C40710 POR2X1_324/O POR2X1_568/Y 0.09fF
C40711 POR2X1_662/Y POR2X1_736/A 0.07fF
C40712 PAND2X1_119/a_76_28# POR2X1_294/A 0.04fF
C40713 POR2X1_68/B PAND2X1_517/O 0.04fF
C40714 PAND2X1_6/A POR2X1_39/B 8.03fF
C40715 INPUT_1 POR2X1_153/Y 0.10fF
C40716 POR2X1_188/O POR2X1_188/Y 0.02fF
C40717 PAND2X1_731/CTRL2 POR2X1_39/B 0.01fF
C40718 POR2X1_416/B POR2X1_745/O 0.16fF
C40719 POR2X1_556/A POR2X1_269/CTRL2 0.01fF
C40720 POR2X1_863/A POR2X1_570/CTRL 0.00fF
C40721 POR2X1_130/O POR2X1_244/Y 0.02fF
C40722 PAND2X1_801/O POR2X1_761/Y 0.01fF
C40723 POR2X1_823/O POR2X1_77/Y 0.16fF
C40724 POR2X1_9/Y POR2X1_625/CTRL 0.09fF
C40725 PAND2X1_276/a_16_344# POR2X1_677/Y 0.01fF
C40726 POR2X1_248/CTRL2 POR2X1_77/Y 0.01fF
C40727 POR2X1_383/A PAND2X1_281/a_56_28# 0.00fF
C40728 PAND2X1_632/A PAND2X1_506/Y 0.12fF
C40729 D_GATE_662 PAND2X1_52/B 0.07fF
C40730 POR2X1_305/O PAND2X1_651/Y 0.00fF
C40731 POR2X1_566/B POR2X1_191/Y 0.07fF
C40732 PAND2X1_266/a_16_344# POR2X1_40/Y 0.01fF
C40733 D_INPUT_5 POR2X1_66/A 1.08fF
C40734 PAND2X1_621/O POR2X1_617/Y 0.03fF
C40735 PAND2X1_621/CTRL POR2X1_616/Y 0.01fF
C40736 PAND2X1_578/Y PAND2X1_771/Y 0.03fF
C40737 POR2X1_772/CTRL POR2X1_294/A 0.03fF
C40738 PAND2X1_601/CTRL2 POR2X1_66/A 0.01fF
C40739 POR2X1_688/Y D_INPUT_0 0.01fF
C40740 POR2X1_65/A PAND2X1_717/A 0.03fF
C40741 POR2X1_634/A POR2X1_705/B 0.03fF
C40742 POR2X1_220/CTRL POR2X1_220/B 0.01fF
C40743 PAND2X1_493/CTRL POR2X1_394/A 0.07fF
C40744 POR2X1_16/A PAND2X1_714/B 0.00fF
C40745 POR2X1_146/CTRL PAND2X1_797/Y 0.01fF
C40746 POR2X1_669/B PAND2X1_750/O 0.15fF
C40747 POR2X1_462/B PAND2X1_52/B 0.03fF
C40748 POR2X1_814/B POR2X1_621/a_56_344# 0.00fF
C40749 POR2X1_169/CTRL POR2X1_191/Y 0.10fF
C40750 POR2X1_169/O POR2X1_192/B 0.07fF
C40751 D_INPUT_1 PAND2X1_52/B 0.10fF
C40752 PAND2X1_193/Y POR2X1_7/B 0.01fF
C40753 POR2X1_343/Y POR2X1_318/A 0.10fF
C40754 POR2X1_411/B POR2X1_69/A 0.10fF
C40755 POR2X1_415/A POR2X1_14/Y 0.07fF
C40756 POR2X1_633/O POR2X1_734/A 0.04fF
C40757 POR2X1_20/B POR2X1_40/Y 0.58fF
C40758 POR2X1_812/A POR2X1_452/Y 1.95fF
C40759 POR2X1_383/A POR2X1_343/a_56_344# 0.00fF
C40760 POR2X1_811/CTRL D_INPUT_0 0.01fF
C40761 PAND2X1_9/Y POR2X1_94/A 0.04fF
C40762 POR2X1_329/A INPUT_0 0.13fF
C40763 POR2X1_416/B PAND2X1_349/A 0.03fF
C40764 POR2X1_422/CTRL POR2X1_422/Y 0.01fF
C40765 POR2X1_864/A POR2X1_828/Y 0.00fF
C40766 POR2X1_475/CTRL POR2X1_288/A 0.00fF
C40767 PAND2X1_48/A PAND2X1_692/O 0.07fF
C40768 POR2X1_490/Y POR2X1_102/Y 0.03fF
C40769 POR2X1_609/Y POR2X1_37/Y 0.05fF
C40770 POR2X1_416/B PAND2X1_114/B 0.03fF
C40771 POR2X1_801/CTRL2 POR2X1_452/Y 0.01fF
C40772 PAND2X1_849/O POR2X1_20/B 0.03fF
C40773 POR2X1_814/A POR2X1_405/Y 0.05fF
C40774 POR2X1_509/O POR2X1_854/B 0.33fF
C40775 POR2X1_13/A POR2X1_667/a_16_28# 0.02fF
C40776 POR2X1_814/A POR2X1_784/A 0.01fF
C40777 POR2X1_502/A PAND2X1_53/O 0.37fF
C40778 POR2X1_612/Y POR2X1_607/CTRL 0.08fF
C40779 POR2X1_502/A POR2X1_459/Y 0.01fF
C40780 POR2X1_508/B POR2X1_191/Y 0.05fF
C40781 PAND2X1_269/O POR2X1_55/Y 0.09fF
C40782 POR2X1_567/A POR2X1_99/B 0.05fF
C40783 POR2X1_260/B POR2X1_186/Y 0.03fF
C40784 POR2X1_666/O POR2X1_32/A 0.12fF
C40785 PAND2X1_20/A POR2X1_637/CTRL 0.00fF
C40786 PAND2X1_96/B POR2X1_643/CTRL 0.00fF
C40787 POR2X1_852/B POR2X1_629/CTRL 0.07fF
C40788 PAND2X1_717/A PAND2X1_303/a_56_28# 0.00fF
C40789 POR2X1_23/Y PAND2X1_658/CTRL 0.01fF
C40790 PAND2X1_796/B PAND2X1_778/O 0.00fF
C40791 PAND2X1_659/B POR2X1_20/B 0.02fF
C40792 PAND2X1_446/Y VDD -0.00fF
C40793 PAND2X1_808/Y POR2X1_250/Y 0.03fF
C40794 POR2X1_76/B POR2X1_366/A 0.05fF
C40795 POR2X1_133/O POR2X1_411/B 0.01fF
C40796 PAND2X1_48/B PAND2X1_417/CTRL2 0.01fF
C40797 POR2X1_854/CTRL VDD 0.00fF
C40798 PAND2X1_3/B D_INPUT_4 0.03fF
C40799 POR2X1_23/Y PAND2X1_61/Y 0.03fF
C40800 POR2X1_341/A POR2X1_220/Y 0.07fF
C40801 POR2X1_271/B POR2X1_293/Y 0.03fF
C40802 POR2X1_123/CTRL POR2X1_556/A 0.01fF
C40803 PAND2X1_851/O PAND2X1_841/Y 0.00fF
C40804 POR2X1_78/B POR2X1_648/m4_208_n4# 0.17fF
C40805 POR2X1_119/Y POR2X1_39/B 0.14fF
C40806 POR2X1_272/CTRL POR2X1_32/A 0.01fF
C40807 PAND2X1_404/Y PAND2X1_474/Y 0.04fF
C40808 POR2X1_590/A POR2X1_330/Y 0.08fF
C40809 PAND2X1_279/O PAND2X1_58/A 0.03fF
C40810 POR2X1_67/A PAND2X1_390/Y 0.03fF
C40811 POR2X1_753/Y POR2X1_750/B 0.07fF
C40812 POR2X1_60/A PAND2X1_786/CTRL 0.01fF
C40813 POR2X1_341/A POR2X1_404/Y 0.09fF
C40814 POR2X1_56/O POR2X1_423/Y 0.02fF
C40815 POR2X1_441/Y PAND2X1_324/Y 0.00fF
C40816 PAND2X1_65/B POR2X1_466/A 0.05fF
C40817 POR2X1_774/Y POR2X1_801/B 0.00fF
C40818 PAND2X1_404/Y POR2X1_13/A 0.05fF
C40819 POR2X1_45/Y POR2X1_275/A 0.12fF
C40820 POR2X1_620/B PAND2X1_52/B 0.05fF
C40821 POR2X1_261/A PAND2X1_771/Y 0.03fF
C40822 POR2X1_119/a_16_28# POR2X1_411/B 0.02fF
C40823 PAND2X1_287/Y PAND2X1_568/O 0.06fF
C40824 POR2X1_15/O PAND2X1_206/B 0.01fF
C40825 PAND2X1_68/a_56_28# POR2X1_5/Y 0.00fF
C40826 POR2X1_106/O POR2X1_106/Y 0.03fF
C40827 PAND2X1_39/B POR2X1_740/Y 0.06fF
C40828 POR2X1_681/Y POR2X1_829/A 0.53fF
C40829 PAND2X1_219/A PAND2X1_733/O 0.01fF
C40830 POR2X1_130/A PAND2X1_591/CTRL 0.01fF
C40831 POR2X1_102/Y PAND2X1_205/Y 0.02fF
C40832 POR2X1_846/CTRL2 POR2X1_129/Y 0.01fF
C40833 POR2X1_156/O POR2X1_728/A 0.00fF
C40834 PAND2X1_23/Y PAND2X1_826/O 0.03fF
C40835 POR2X1_814/A POR2X1_729/Y 0.33fF
C40836 PAND2X1_464/B POR2X1_91/Y 0.03fF
C40837 POR2X1_709/A PAND2X1_411/O 0.01fF
C40838 POR2X1_68/A PAND2X1_761/O 0.03fF
C40839 PAND2X1_404/Y PAND2X1_197/O 0.03fF
C40840 POR2X1_556/A POR2X1_501/B 0.03fF
C40841 PAND2X1_203/CTRL POR2X1_816/A 0.01fF
C40842 POR2X1_82/CTRL2 POR2X1_14/Y 0.03fF
C40843 POR2X1_288/a_16_28# POR2X1_286/Y -0.00fF
C40844 POR2X1_134/Y POR2X1_20/B 0.05fF
C40845 POR2X1_699/O POR2X1_7/B 0.01fF
C40846 POR2X1_621/A PAND2X1_6/A 0.08fF
C40847 POR2X1_502/A D_INPUT_0 0.08fF
C40848 POR2X1_68/A PAND2X1_826/CTRL 0.03fF
C40849 PAND2X1_5/CTRL2 INPUT_3 0.03fF
C40850 D_INPUT_0 POR2X1_783/A 0.01fF
C40851 PAND2X1_246/CTRL2 PAND2X1_63/B 0.01fF
C40852 PAND2X1_469/B POR2X1_273/CTRL 0.16fF
C40853 POR2X1_811/A POR2X1_783/A 0.27fF
C40854 PAND2X1_623/Y POR2X1_848/A 0.12fF
C40855 PAND2X1_23/Y POR2X1_458/CTRL 0.04fF
C40856 POR2X1_497/CTRL2 PAND2X1_501/B 0.01fF
C40857 D_INPUT_2 POR2X1_612/B 0.04fF
C40858 PAND2X1_677/CTRL PAND2X1_90/Y 0.03fF
C40859 PAND2X1_293/CTRL2 PAND2X1_58/A 0.00fF
C40860 POR2X1_243/A INPUT_0 0.02fF
C40861 POR2X1_476/Y POR2X1_643/A 0.04fF
C40862 POR2X1_121/A POR2X1_260/B 0.03fF
C40863 POR2X1_558/B POR2X1_572/B 0.02fF
C40864 POR2X1_20/B PAND2X1_840/CTRL2 0.02fF
C40865 POR2X1_654/B POR2X1_287/B 0.03fF
C40866 POR2X1_609/Y POR2X1_293/Y 0.06fF
C40867 PAND2X1_229/a_16_344# POR2X1_186/Y 0.02fF
C40868 POR2X1_448/a_16_28# POR2X1_448/A 0.05fF
C40869 PAND2X1_23/Y POR2X1_294/Y 0.27fF
C40870 D_INPUT_3 INPUT_3 0.50fF
C40871 POR2X1_677/Y PAND2X1_716/B 0.03fF
C40872 PAND2X1_236/CTRL POR2X1_94/A 0.01fF
C40873 PAND2X1_82/CTRL2 PAND2X1_39/B 0.05fF
C40874 POR2X1_487/Y PAND2X1_580/B 0.00fF
C40875 POR2X1_423/Y PAND2X1_473/B 0.12fF
C40876 POR2X1_356/A PAND2X1_73/Y 0.09fF
C40877 POR2X1_309/CTRL POR2X1_293/Y 0.01fF
C40878 POR2X1_287/B POR2X1_850/A 0.71fF
C40879 PAND2X1_6/Y PAND2X1_93/B 6.29fF
C40880 POR2X1_39/CTRL POR2X1_236/Y 0.03fF
C40881 POR2X1_307/Y PAND2X1_58/A 0.03fF
C40882 POR2X1_624/Y POR2X1_318/A 0.08fF
C40883 POR2X1_376/B POR2X1_743/CTRL 0.01fF
C40884 POR2X1_48/A PAND2X1_6/A 0.37fF
C40885 POR2X1_23/Y POR2X1_255/Y 0.10fF
C40886 POR2X1_623/O PAND2X1_6/A 0.07fF
C40887 POR2X1_48/A PAND2X1_731/CTRL2 0.03fF
C40888 PAND2X1_243/B POR2X1_102/Y 0.01fF
C40889 POR2X1_775/A POR2X1_97/A 0.07fF
C40890 POR2X1_56/B POR2X1_14/Y 0.03fF
C40891 POR2X1_660/O PAND2X1_55/Y 0.17fF
C40892 POR2X1_102/Y PAND2X1_219/CTRL2 0.01fF
C40893 POR2X1_502/A PAND2X1_278/CTRL2 0.01fF
C40894 POR2X1_405/CTRL2 POR2X1_405/Y 0.00fF
C40895 POR2X1_56/B PAND2X1_453/A 1.59fF
C40896 PAND2X1_65/B POR2X1_448/A 0.00fF
C40897 POR2X1_96/A POR2X1_72/B 0.14fF
C40898 PAND2X1_845/O POR2X1_37/Y 0.03fF
C40899 PAND2X1_394/m4_208_n4# POR2X1_207/m4_208_n4# 0.13fF
C40900 PAND2X1_217/B POR2X1_498/O 0.02fF
C40901 POR2X1_192/Y POR2X1_509/B 0.11fF
C40902 POR2X1_475/A VDD 0.51fF
C40903 PAND2X1_53/CTRL2 PAND2X1_48/A 0.14fF
C40904 POR2X1_511/Y PAND2X1_513/m4_208_n4# 0.08fF
C40905 PAND2X1_20/A POR2X1_740/Y 0.03fF
C40906 PAND2X1_859/O INPUT_0 0.14fF
C40907 POR2X1_16/A POR2X1_411/B 3.65fF
C40908 PAND2X1_638/B POR2X1_790/B 0.03fF
C40909 PAND2X1_35/a_76_28# POR2X1_394/A 0.02fF
C40910 POR2X1_5/Y PAND2X1_8/Y 0.07fF
C40911 POR2X1_97/B POR2X1_814/A 0.16fF
C40912 POR2X1_833/A POR2X1_541/B 0.46fF
C40913 POR2X1_687/A POR2X1_803/a_56_344# 0.00fF
C40914 POR2X1_45/Y POR2X1_60/A 0.03fF
C40915 PAND2X1_738/Y POR2X1_106/Y 0.05fF
C40916 POR2X1_409/Y PAND2X1_9/Y 0.01fF
C40917 POR2X1_78/CTRL2 POR2X1_78/A 0.00fF
C40918 PAND2X1_667/CTRL2 INPUT_0 0.03fF
C40919 POR2X1_327/Y POR2X1_554/B 0.02fF
C40920 POR2X1_41/B PAND2X1_620/Y 0.09fF
C40921 PAND2X1_714/O PAND2X1_731/B 0.02fF
C40922 POR2X1_355/a_56_344# POR2X1_192/Y 0.03fF
C40923 POR2X1_389/A PAND2X1_666/CTRL 0.00fF
C40924 PAND2X1_6/Y POR2X1_78/A 2.22fF
C40925 POR2X1_41/B POR2X1_65/A 4.14fF
C40926 PAND2X1_464/B POR2X1_109/Y 0.03fF
C40927 D_INPUT_3 POR2X1_14/CTRL 0.06fF
C40928 POR2X1_341/A POR2X1_332/CTRL 0.03fF
C40929 POR2X1_502/A PAND2X1_90/Y 0.27fF
C40930 PAND2X1_3/a_16_344# D_INPUT_5 0.01fF
C40931 POR2X1_856/B PAND2X1_60/B 0.03fF
C40932 PAND2X1_272/O POR2X1_573/A 0.04fF
C40933 POR2X1_66/B PAND2X1_612/CTRL2 0.00fF
C40934 PAND2X1_853/CTRL2 POR2X1_40/Y 0.02fF
C40935 PAND2X1_55/Y POR2X1_186/Y 0.76fF
C40936 POR2X1_750/B POR2X1_459/A 0.02fF
C40937 PAND2X1_118/CTRL2 PAND2X1_41/B 0.01fF
C40938 PAND2X1_738/Y PAND2X1_580/B 0.03fF
C40939 PAND2X1_808/Y POR2X1_488/CTRL2 0.01fF
C40940 PAND2X1_55/Y POR2X1_202/a_16_28# 0.03fF
C40941 POR2X1_272/CTRL POR2X1_184/Y 0.00fF
C40942 POR2X1_423/Y PAND2X1_390/O 0.02fF
C40943 POR2X1_632/B POR2X1_532/A 0.15fF
C40944 POR2X1_697/Y POR2X1_427/Y 0.04fF
C40945 PAND2X1_90/Y PAND2X1_176/O 0.01fF
C40946 POR2X1_46/Y PAND2X1_332/a_56_28# 0.00fF
C40947 POR2X1_814/B POR2X1_740/Y 0.03fF
C40948 POR2X1_687/O POR2X1_729/Y 0.01fF
C40949 PAND2X1_58/A POR2X1_68/B 0.76fF
C40950 POR2X1_686/B POR2X1_220/Y 0.03fF
C40951 POR2X1_464/Y PAND2X1_90/Y 0.08fF
C40952 POR2X1_624/Y POR2X1_574/Y 0.07fF
C40953 INPUT_1 POR2X1_248/A 0.01fF
C40954 POR2X1_48/A POR2X1_280/Y 0.43fF
C40955 PAND2X1_90/Y POR2X1_532/Y 0.05fF
C40956 POR2X1_82/CTRL2 POR2X1_55/Y 0.00fF
C40957 PAND2X1_39/B POR2X1_774/A 0.03fF
C40958 POR2X1_278/Y PAND2X1_862/B 0.12fF
C40959 POR2X1_327/CTRL VDD 0.00fF
C40960 POR2X1_863/B VDD 0.02fF
C40961 POR2X1_423/O POR2X1_387/Y 0.05fF
C40962 PAND2X1_531/O PAND2X1_111/B 0.01fF
C40963 PAND2X1_626/a_76_28# PAND2X1_96/B 0.01fF
C40964 PAND2X1_250/CTRL2 PAND2X1_32/B 0.02fF
C40965 POR2X1_809/A PAND2X1_761/a_16_344# 0.01fF
C40966 POR2X1_542/B POR2X1_750/B 0.03fF
C40967 PAND2X1_65/B POR2X1_341/CTRL 0.01fF
C40968 POR2X1_629/A VDD 0.00fF
C40969 POR2X1_740/Y POR2X1_325/A 0.05fF
C40970 PAND2X1_240/O POR2X1_232/Y 0.00fF
C40971 POR2X1_623/B PAND2X1_63/B 0.01fF
C40972 POR2X1_614/A POR2X1_543/A 0.08fF
C40973 POR2X1_66/B POR2X1_137/Y 0.03fF
C40974 PAND2X1_299/CTRL PAND2X1_32/B 0.01fF
C40975 PAND2X1_73/Y POR2X1_569/A 0.10fF
C40976 POR2X1_149/B PAND2X1_65/B 0.03fF
C40977 POR2X1_65/A PAND2X1_640/O 0.03fF
C40978 POR2X1_106/O PAND2X1_114/B 0.01fF
C40979 GATE_479 POR2X1_694/O 0.02fF
C40980 POR2X1_329/A POR2X1_522/CTRL2 0.01fF
C40981 POR2X1_614/A PAND2X1_679/O 0.16fF
C40982 POR2X1_332/B POR2X1_193/A 0.03fF
C40983 POR2X1_856/B POR2X1_353/A 0.03fF
C40984 POR2X1_194/A POR2X1_194/CTRL2 0.02fF
C40985 POR2X1_332/B POR2X1_579/Y 0.00fF
C40986 POR2X1_123/Y PAND2X1_41/B 0.01fF
C40987 POR2X1_49/Y PAND2X1_470/O 0.15fF
C40988 PAND2X1_471/B POR2X1_7/B 0.01fF
C40989 POR2X1_383/A POR2X1_811/B 0.14fF
C40990 POR2X1_68/A POR2X1_480/A 1.22fF
C40991 PAND2X1_213/Y POR2X1_417/Y 4.64fF
C40992 POR2X1_177/Y PAND2X1_566/Y 0.01fF
C40993 POR2X1_96/Y POR2X1_63/Y 0.03fF
C40994 POR2X1_29/A POR2X1_750/Y 0.03fF
C40995 POR2X1_333/Y PAND2X1_237/O 0.00fF
C40996 POR2X1_475/A PAND2X1_32/B 0.23fF
C40997 PAND2X1_775/CTRL POR2X1_7/B 0.01fF
C40998 POR2X1_119/Y PAND2X1_469/CTRL2 0.00fF
C40999 POR2X1_670/Y POR2X1_13/A 0.12fF
C41000 PAND2X1_41/B POR2X1_216/CTRL 0.00fF
C41001 PAND2X1_65/B POR2X1_644/A 0.05fF
C41002 PAND2X1_711/O POR2X1_763/A 0.08fF
C41003 PAND2X1_435/CTRL2 POR2X1_433/Y 0.02fF
C41004 PAND2X1_655/Y POR2X1_413/A 0.04fF
C41005 PAND2X1_480/B PAND2X1_798/B 0.05fF
C41006 POR2X1_72/B POR2X1_7/A 0.17fF
C41007 POR2X1_68/A POR2X1_243/Y 0.07fF
C41008 POR2X1_207/B POR2X1_207/A 0.36fF
C41009 POR2X1_10/CTRL2 POR2X1_83/B 0.00fF
C41010 PAND2X1_652/A POR2X1_79/Y 0.03fF
C41011 POR2X1_416/B POR2X1_411/A 0.03fF
C41012 POR2X1_435/CTRL VDD 0.00fF
C41013 POR2X1_57/A PAND2X1_756/CTRL2 0.03fF
C41014 POR2X1_471/A PAND2X1_179/O 0.08fF
C41015 PAND2X1_592/Y POR2X1_42/Y 0.93fF
C41016 PAND2X1_215/B PAND2X1_197/Y 0.07fF
C41017 POR2X1_383/A POR2X1_254/O 0.05fF
C41018 PAND2X1_654/A POR2X1_32/A 0.09fF
C41019 POR2X1_614/A POR2X1_332/B 0.04fF
C41020 PAND2X1_716/CTRL2 PAND2X1_364/B 0.05fF
C41021 POR2X1_144/CTRL2 POR2X1_669/B 0.03fF
C41022 POR2X1_348/O POR2X1_814/B 0.01fF
C41023 POR2X1_3/A POR2X1_2/CTRL 0.00fF
C41024 POR2X1_786/CTRL2 PAND2X1_60/B 0.06fF
C41025 POR2X1_52/A POR2X1_437/Y 0.01fF
C41026 PAND2X1_830/Y POR2X1_183/Y 0.02fF
C41027 POR2X1_41/Y PAND2X1_852/A 0.01fF
C41028 VDD POR2X1_140/CTRL 0.00fF
C41029 POR2X1_515/CTRL2 PAND2X1_60/B 0.10fF
C41030 POR2X1_119/Y POR2X1_48/A 0.19fF
C41031 POR2X1_350/Y POR2X1_776/B 0.07fF
C41032 POR2X1_549/O POR2X1_383/A 0.02fF
C41033 PAND2X1_766/CTRL2 POR2X1_260/A 0.01fF
C41034 POR2X1_83/B POR2X1_394/A 0.31fF
C41035 POR2X1_750/B PAND2X1_376/CTRL 0.01fF
C41036 POR2X1_57/A INPUT_0 0.06fF
C41037 POR2X1_225/a_76_344# POR2X1_129/Y 0.00fF
C41038 POR2X1_805/Y POR2X1_774/A 0.00fF
C41039 POR2X1_68/A PAND2X1_90/A 0.03fF
C41040 POR2X1_121/A PAND2X1_55/Y 0.07fF
C41041 PAND2X1_340/a_76_28# POR2X1_408/Y 0.05fF
C41042 PAND2X1_715/B POR2X1_40/Y 0.01fF
C41043 POR2X1_172/Y VDD 0.28fF
C41044 D_INPUT_0 POR2X1_188/Y 10.80fF
C41045 POR2X1_137/B PAND2X1_52/B 0.72fF
C41046 POR2X1_750/B POR2X1_754/O 0.05fF
C41047 PAND2X1_20/A POR2X1_774/A 0.06fF
C41048 PAND2X1_41/B PAND2X1_503/O 0.08fF
C41049 POR2X1_212/CTRL2 VDD -0.00fF
C41050 PAND2X1_183/CTRL POR2X1_540/A 0.01fF
C41051 PAND2X1_787/A PAND2X1_151/O 0.05fF
C41052 POR2X1_634/O POR2X1_559/A 0.02fF
C41053 PAND2X1_840/A PAND2X1_840/B 0.20fF
C41054 POR2X1_65/A POR2X1_291/O 0.01fF
C41055 PAND2X1_207/CTRL2 PAND2X1_207/A 0.01fF
C41056 PAND2X1_214/A POR2X1_153/Y 0.03fF
C41057 PAND2X1_107/CTRL PAND2X1_65/B 0.01fF
C41058 PAND2X1_568/B PAND2X1_568/CTRL 0.01fF
C41059 POR2X1_43/B PAND2X1_339/Y 0.14fF
C41060 PAND2X1_137/O POR2X1_132/Y 0.01fF
C41061 POR2X1_16/A POR2X1_376/B 0.05fF
C41062 POR2X1_85/O POR2X1_23/Y 0.01fF
C41063 POR2X1_32/A POR2X1_701/a_56_344# 0.01fF
C41064 PAND2X1_20/A POR2X1_550/B 0.01fF
C41065 POR2X1_832/A PAND2X1_57/B 0.15fF
C41066 PAND2X1_738/Y PAND2X1_349/A 0.05fF
C41067 POR2X1_73/CTRL VDD 0.00fF
C41068 PAND2X1_736/A PAND2X1_186/CTRL2 0.02fF
C41069 POR2X1_722/Y PAND2X1_60/B 0.01fF
C41070 POR2X1_65/A PAND2X1_308/Y 0.03fF
C41071 POR2X1_356/A PAND2X1_173/CTRL2 0.15fF
C41072 PAND2X1_57/B POR2X1_780/B 0.01fF
C41073 PAND2X1_220/Y PAND2X1_348/A 0.12fF
C41074 POR2X1_244/B POR2X1_854/B 0.05fF
C41075 POR2X1_219/a_76_344# POR2X1_294/B 0.00fF
C41076 PAND2X1_93/B POR2X1_632/Y 0.04fF
C41077 PAND2X1_370/CTRL POR2X1_309/Y 0.01fF
C41078 PAND2X1_599/a_16_344# PAND2X1_69/A 0.01fF
C41079 POR2X1_750/A POR2X1_749/a_16_28# 0.03fF
C41080 PAND2X1_23/Y POR2X1_544/CTRL 0.01fF
C41081 PAND2X1_82/Y PAND2X1_57/B 0.03fF
C41082 PAND2X1_23/Y POR2X1_249/a_16_28# 0.02fF
C41083 POR2X1_389/CTRL2 POR2X1_537/B 0.06fF
C41084 PAND2X1_242/Y POR2X1_271/B 0.05fF
C41085 POR2X1_390/B POR2X1_335/O 0.00fF
C41086 POR2X1_87/B PAND2X1_39/B 0.02fF
C41087 POR2X1_814/B POR2X1_774/A 0.03fF
C41088 POR2X1_138/O POR2X1_318/A 0.02fF
C41089 POR2X1_365/Y POR2X1_319/Y 0.03fF
C41090 D_INPUT_3 POR2X1_119/a_76_344# 0.01fF
C41091 POR2X1_468/a_16_28# POR2X1_478/B 0.00fF
C41092 POR2X1_538/A POR2X1_193/A 0.01fF
C41093 PAND2X1_847/CTRL POR2X1_48/A 0.03fF
C41094 PAND2X1_94/A POR2X1_124/CTRL 0.14fF
C41095 POR2X1_445/A POR2X1_863/A 0.01fF
C41096 PAND2X1_724/CTRL POR2X1_73/Y 0.01fF
C41097 VDD POR2X1_724/B 0.05fF
C41098 POR2X1_121/A POR2X1_121/a_56_344# 0.00fF
C41099 POR2X1_722/Y POR2X1_353/A 0.06fF
C41100 INPUT_0 POR2X1_559/A 0.17fF
C41101 PAND2X1_96/B POR2X1_68/B 0.03fF
C41102 POR2X1_78/B PAND2X1_399/O 0.04fF
C41103 PAND2X1_139/B POR2X1_129/Y 0.05fF
C41104 POR2X1_52/A POR2X1_16/A 0.28fF
C41105 PAND2X1_330/a_56_28# POR2X1_385/Y 0.00fF
C41106 POR2X1_416/B POR2X1_32/A 0.28fF
C41107 POR2X1_557/B VDD 0.33fF
C41108 PAND2X1_795/B POR2X1_394/A 0.09fF
C41109 POR2X1_442/Y POR2X1_39/B 0.05fF
C41110 PAND2X1_659/Y PAND2X1_736/CTRL 0.00fF
C41111 PAND2X1_194/CTRL2 POR2X1_73/Y 0.03fF
C41112 POR2X1_865/B POR2X1_458/B 0.03fF
C41113 PAND2X1_318/a_76_28# POR2X1_315/Y 0.02fF
C41114 POR2X1_38/Y POR2X1_591/Y 0.03fF
C41115 PAND2X1_498/O POR2X1_260/A 0.16fF
C41116 PAND2X1_343/CTRL2 POR2X1_42/Y 0.01fF
C41117 POR2X1_186/Y POR2X1_741/O 0.02fF
C41118 PAND2X1_90/Y POR2X1_188/Y 0.05fF
C41119 POR2X1_572/B POR2X1_362/A 0.01fF
C41120 POR2X1_224/a_16_28# POR2X1_394/A 0.09fF
C41121 POR2X1_16/A POR2X1_152/A 0.03fF
C41122 PAND2X1_440/CTRL POR2X1_60/A 0.01fF
C41123 PAND2X1_341/B PAND2X1_206/CTRL2 0.01fF
C41124 POR2X1_326/A POR2X1_435/Y 0.08fF
C41125 POR2X1_219/B POR2X1_215/Y 0.02fF
C41126 PAND2X1_592/a_16_344# PAND2X1_853/B 0.01fF
C41127 PAND2X1_65/B PAND2X1_179/CTRL2 0.01fF
C41128 POR2X1_254/Y PAND2X1_48/A 0.00fF
C41129 PAND2X1_73/Y PAND2X1_72/A 0.23fF
C41130 POR2X1_78/A PAND2X1_52/B 0.15fF
C41131 POR2X1_438/a_16_28# POR2X1_142/Y 0.01fF
C41132 POR2X1_102/Y PAND2X1_862/CTRL 0.01fF
C41133 POR2X1_278/Y PAND2X1_716/B 0.07fF
C41134 POR2X1_346/B POR2X1_68/A 0.08fF
C41135 POR2X1_614/A POR2X1_520/a_56_344# 0.00fF
C41136 PAND2X1_772/a_76_28# POR2X1_77/Y 0.01fF
C41137 POR2X1_416/B POR2X1_417/Y 0.03fF
C41138 POR2X1_222/A PAND2X1_88/Y 0.04fF
C41139 PAND2X1_390/Y PAND2X1_840/Y 0.00fF
C41140 PAND2X1_511/a_76_28# PAND2X1_48/A 0.01fF
C41141 POR2X1_840/B POR2X1_141/A 0.03fF
C41142 PAND2X1_69/A PAND2X1_528/O 0.00fF
C41143 POR2X1_833/CTRL2 POR2X1_186/B 0.01fF
C41144 POR2X1_831/CTRL POR2X1_814/A 0.01fF
C41145 POR2X1_93/A POR2X1_283/A 0.14fF
C41146 POR2X1_123/B POR2X1_123/A 0.30fF
C41147 POR2X1_717/CTRL2 POR2X1_101/Y 0.13fF
C41148 POR2X1_283/A POR2X1_91/Y 0.07fF
C41149 POR2X1_564/Y POR2X1_337/Y 0.06fF
C41150 POR2X1_86/Y POR2X1_40/Y 0.01fF
C41151 PAND2X1_491/O PAND2X1_94/A 0.04fF
C41152 POR2X1_503/A POR2X1_77/Y 0.05fF
C41153 POR2X1_559/O POR2X1_673/Y 0.02fF
C41154 PAND2X1_800/a_16_344# POR2X1_42/Y 0.02fF
C41155 POR2X1_65/A POR2X1_77/Y 3.07fF
C41156 POR2X1_706/B POR2X1_711/Y 0.01fF
C41157 PAND2X1_69/A POR2X1_675/Y 0.03fF
C41158 PAND2X1_341/A PAND2X1_100/O 0.02fF
C41159 POR2X1_575/B PAND2X1_48/A 0.76fF
C41160 POR2X1_65/A POR2X1_85/Y 0.02fF
C41161 POR2X1_422/Y POR2X1_386/Y 0.03fF
C41162 PAND2X1_38/a_76_28# POR2X1_4/Y 0.03fF
C41163 POR2X1_740/Y POR2X1_726/CTRL 0.00fF
C41164 PAND2X1_654/A PAND2X1_651/Y 0.00fF
C41165 POR2X1_119/Y PAND2X1_197/Y 0.05fF
C41166 PAND2X1_661/CTRL2 POR2X1_761/A 0.01fF
C41167 POR2X1_96/A POR2X1_304/CTRL 0.01fF
C41168 PAND2X1_652/A PAND2X1_730/A 0.03fF
C41169 POR2X1_592/Y POR2X1_220/Y 0.00fF
C41170 POR2X1_78/B PAND2X1_56/A 0.03fF
C41171 POR2X1_416/B PAND2X1_741/B 0.03fF
C41172 PAND2X1_551/O PAND2X1_545/Y 0.00fF
C41173 POR2X1_62/Y PAND2X1_6/A 0.26fF
C41174 POR2X1_557/B PAND2X1_32/B 0.06fF
C41175 POR2X1_43/B PAND2X1_338/CTRL2 0.01fF
C41176 POR2X1_567/A POR2X1_775/A 0.03fF
C41177 POR2X1_350/Y POR2X1_192/B 0.18fF
C41178 POR2X1_465/O POR2X1_454/A 0.09fF
C41179 POR2X1_326/A PAND2X1_96/B 0.12fF
C41180 POR2X1_244/Y PAND2X1_60/B 0.03fF
C41181 POR2X1_843/CTRL POR2X1_458/Y 0.01fF
C41182 POR2X1_96/A POR2X1_305/CTRL 0.02fF
C41183 PAND2X1_715/m4_208_n4# POR2X1_39/B 0.15fF
C41184 POR2X1_359/B POR2X1_532/A 0.14fF
C41185 PAND2X1_285/CTRL POR2X1_282/Y 0.01fF
C41186 POR2X1_40/Y POR2X1_321/CTRL 0.01fF
C41187 POR2X1_394/A POR2X1_380/A 0.02fF
C41188 PAND2X1_492/CTRL PAND2X1_72/A 0.04fF
C41189 POR2X1_318/A POR2X1_186/B 0.07fF
C41190 POR2X1_796/A POR2X1_260/A 0.03fF
C41191 PAND2X1_59/O PAND2X1_18/B 0.04fF
C41192 PAND2X1_683/O PAND2X1_69/A 0.03fF
C41193 PAND2X1_659/Y POR2X1_498/A 0.00fF
C41194 INPUT_1 PAND2X1_483/CTRL2 0.01fF
C41195 POR2X1_416/B PAND2X1_35/Y 0.05fF
C41196 PAND2X1_631/CTRL PAND2X1_631/A 0.02fF
C41197 PAND2X1_560/B PAND2X1_656/A 0.03fF
C41198 POR2X1_353/A POR2X1_151/CTRL2 0.01fF
C41199 POR2X1_347/O POR2X1_402/A 0.01fF
C41200 POR2X1_416/B POR2X1_57/CTRL 0.08fF
C41201 POR2X1_325/O POR2X1_544/B 0.01fF
C41202 POR2X1_614/A POR2X1_560/a_16_28# 0.03fF
C41203 POR2X1_188/a_16_28# POR2X1_733/Y 0.02fF
C41204 POR2X1_840/Y POR2X1_513/Y 0.01fF
C41205 PAND2X1_334/CTRL POR2X1_39/B 0.01fF
C41206 POR2X1_102/Y POR2X1_329/A 1.89fF
C41207 PAND2X1_350/CTRL2 POR2X1_4/Y 0.03fF
C41208 POR2X1_648/Y POR2X1_811/B 0.03fF
C41209 POR2X1_150/Y D_INPUT_0 0.03fF
C41210 POR2X1_110/O POR2X1_7/A 0.04fF
C41211 POR2X1_609/Y POR2X1_412/O 0.01fF
C41212 POR2X1_384/A POR2X1_384/a_16_28# 0.03fF
C41213 POR2X1_68/A POR2X1_716/CTRL 0.14fF
C41214 POR2X1_78/a_16_28# D_INPUT_0 0.03fF
C41215 POR2X1_796/Y POR2X1_808/CTRL2 0.01fF
C41216 POR2X1_63/Y POR2X1_37/Y 0.03fF
C41217 POR2X1_78/B POR2X1_661/A 0.07fF
C41218 POR2X1_416/B POR2X1_184/Y 0.05fF
C41219 POR2X1_451/A POR2X1_635/Y 0.01fF
C41220 PAND2X1_569/B POR2X1_373/CTRL 0.03fF
C41221 POR2X1_75/CTRL POR2X1_416/B 0.01fF
C41222 POR2X1_54/Y PAND2X1_669/CTRL 0.28fF
C41223 PAND2X1_651/Y POR2X1_416/B 0.03fF
C41224 POR2X1_509/O POR2X1_509/A 0.06fF
C41225 POR2X1_510/A PAND2X1_52/B 0.03fF
C41226 PAND2X1_55/Y POR2X1_556/CTRL 0.01fF
C41227 POR2X1_77/Y PAND2X1_359/B 0.03fF
C41228 PAND2X1_32/a_76_28# POR2X1_94/A 0.01fF
C41229 POR2X1_60/A POR2X1_271/B 0.03fF
C41230 POR2X1_760/A POR2X1_72/B 0.23fF
C41231 PAND2X1_606/CTRL POR2X1_37/Y 0.03fF
C41232 POR2X1_27/CTRL POR2X1_5/Y 0.01fF
C41233 PAND2X1_857/A POR2X1_761/A 0.03fF
C41234 POR2X1_52/O POR2X1_7/A 0.01fF
C41235 POR2X1_191/Y POR2X1_353/A 0.01fF
C41236 POR2X1_65/A PAND2X1_449/O 0.04fF
C41237 PAND2X1_399/O POR2X1_294/A 0.15fF
C41238 PAND2X1_173/CTRL2 PAND2X1_72/A 0.00fF
C41239 PAND2X1_106/O POR2X1_343/Y 0.00fF
C41240 POR2X1_357/CTRL POR2X1_191/Y 0.12fF
C41241 POR2X1_357/O POR2X1_192/B 0.07fF
C41242 POR2X1_669/B PAND2X1_124/Y 0.63fF
C41243 POR2X1_127/Y POR2X1_411/B 0.03fF
C41244 PAND2X1_58/A POR2X1_606/O 0.01fF
C41245 POR2X1_630/CTRL POR2X1_590/A 0.01fF
C41246 PAND2X1_39/B POR2X1_780/O 0.12fF
C41247 POR2X1_278/Y POR2X1_250/Y 0.10fF
C41248 POR2X1_558/B POR2X1_590/A 0.17fF
C41249 POR2X1_475/A POR2X1_475/CTRL2 0.01fF
C41250 POR2X1_327/Y POR2X1_741/CTRL 0.06fF
C41251 POR2X1_848/A PAND2X1_58/A 0.10fF
C41252 PAND2X1_108/a_76_28# POR2X1_814/A 0.04fF
C41253 PAND2X1_65/B POR2X1_633/a_16_28# 0.03fF
C41254 POR2X1_20/B POR2X1_5/Y 0.15fF
C41255 PAND2X1_163/O PAND2X1_72/A 0.01fF
C41256 POR2X1_149/CTRL2 PAND2X1_90/Y 0.01fF
C41257 PAND2X1_257/O POR2X1_222/Y 0.10fF
C41258 POR2X1_191/O POR2X1_191/B 0.04fF
C41259 POR2X1_648/Y POR2X1_783/B 0.01fF
C41260 POR2X1_445/A POR2X1_456/CTRL 0.10fF
C41261 POR2X1_760/A PAND2X1_216/CTRL 0.03fF
C41262 POR2X1_43/CTRL PAND2X1_560/B 0.03fF
C41263 POR2X1_66/B POR2X1_286/CTRL 0.01fF
C41264 POR2X1_456/B POR2X1_181/Y 0.03fF
C41265 POR2X1_65/CTRL2 POR2X1_55/Y 0.21fF
C41266 POR2X1_63/Y POR2X1_406/Y 0.63fF
C41267 PAND2X1_23/Y PAND2X1_45/CTRL2 0.01fF
C41268 POR2X1_83/B POR2X1_669/B 15.12fF
C41269 POR2X1_121/B POR2X1_296/B 0.03fF
C41270 POR2X1_48/A PAND2X1_456/CTRL2 0.14fF
C41271 PAND2X1_677/O POR2X1_66/A 0.05fF
C41272 POR2X1_66/A POR2X1_330/Y 0.11fF
C41273 POR2X1_856/B POR2X1_750/B 0.13fF
C41274 POR2X1_559/Y POR2X1_814/A 0.01fF
C41275 POR2X1_313/Y POR2X1_167/Y 0.08fF
C41276 PAND2X1_2/O D_INPUT_4 0.10fF
C41277 POR2X1_820/B PAND2X1_340/B 0.00fF
C41278 POR2X1_174/B POR2X1_836/A 0.03fF
C41279 POR2X1_462/B POR2X1_848/O 0.01fF
C41280 PAND2X1_639/m4_208_n4# POR2X1_583/m4_208_n4# 0.13fF
C41281 POR2X1_20/CTRL POR2X1_20/B 0.01fF
C41282 POR2X1_624/Y PAND2X1_131/O 0.01fF
C41283 POR2X1_728/B POR2X1_452/Y 0.07fF
C41284 POR2X1_669/B POR2X1_626/Y -0.02fF
C41285 POR2X1_467/Y POR2X1_78/A 0.03fF
C41286 POR2X1_294/A PAND2X1_56/A 0.03fF
C41287 POR2X1_63/Y POR2X1_293/Y 0.03fF
C41288 POR2X1_863/A POR2X1_260/A 0.45fF
C41289 POR2X1_541/B POR2X1_294/B 0.17fF
C41290 POR2X1_729/m4_208_n4# POR2X1_814/A 0.06fF
C41291 POR2X1_54/Y POR2X1_790/CTRL 0.01fF
C41292 POR2X1_48/A PAND2X1_725/B 0.01fF
C41293 POR2X1_257/A INPUT_5 1.43fF
C41294 PAND2X1_654/CTRL2 PAND2X1_9/Y 0.01fF
C41295 POR2X1_311/Y POR2X1_251/A 0.01fF
C41296 POR2X1_186/Y PAND2X1_331/CTRL 0.01fF
C41297 POR2X1_792/O PAND2X1_41/B 0.05fF
C41298 PAND2X1_695/a_16_344# PAND2X1_59/B 0.03fF
C41299 POR2X1_480/a_16_28# POR2X1_480/A -0.00fF
C41300 POR2X1_186/Y POR2X1_174/A 0.04fF
C41301 POR2X1_814/B PAND2X1_15/CTRL 0.02fF
C41302 PAND2X1_688/CTRL POR2X1_48/A 0.01fF
C41303 D_GATE_662 POR2X1_444/O 0.05fF
C41304 POR2X1_278/Y POR2X1_490/Y 0.05fF
C41305 POR2X1_866/A PAND2X1_511/a_16_344# 0.02fF
C41306 PAND2X1_326/B POR2X1_39/B 0.03fF
C41307 POR2X1_477/A POR2X1_477/a_16_28# 0.03fF
C41308 D_INPUT_7 POR2X1_1/O 0.08fF
C41309 POR2X1_265/CTRL PAND2X1_35/Y 0.01fF
C41310 PAND2X1_307/a_56_28# POR2X1_102/Y 0.00fF
C41311 POR2X1_49/Y POR2X1_421/Y 0.12fF
C41312 D_INPUT_5 PAND2X1_17/O 0.17fF
C41313 POR2X1_614/A PAND2X1_425/Y 1.04fF
C41314 PAND2X1_205/A POR2X1_79/Y 0.17fF
C41315 POR2X1_637/CTRL VDD 0.00fF
C41316 POR2X1_23/Y POR2X1_46/Y 0.12fF
C41317 POR2X1_257/A POR2X1_426/O 0.01fF
C41318 PAND2X1_475/a_16_344# POR2X1_72/B 0.02fF
C41319 POR2X1_9/Y POR2X1_260/A 0.07fF
C41320 POR2X1_116/A POR2X1_840/B 0.05fF
C41321 PAND2X1_73/Y POR2X1_285/O 0.02fF
C41322 POR2X1_67/Y POR2X1_391/a_56_344# 0.00fF
C41323 POR2X1_102/Y PAND2X1_795/m4_208_n4# 0.09fF
C41324 POR2X1_77/Y PAND2X1_169/O 0.01fF
C41325 POR2X1_66/B POR2X1_650/A 0.01fF
C41326 POR2X1_568/A POR2X1_551/A 0.03fF
C41327 POR2X1_760/A PAND2X1_799/O 0.02fF
C41328 PAND2X1_58/A POR2X1_480/A 0.07fF
C41329 PAND2X1_48/B PAND2X1_251/CTRL 0.00fF
C41330 POR2X1_159/CTRL POR2X1_376/B 0.01fF
C41331 POR2X1_20/B POR2X1_299/O 0.01fF
C41332 PAND2X1_24/CTRL2 D_INPUT_1 0.01fF
C41333 POR2X1_547/a_76_344# POR2X1_624/Y 0.01fF
C41334 PAND2X1_809/O PAND2X1_539/Y 0.02fF
C41335 D_INPUT_0 PAND2X1_364/B 0.23fF
C41336 POR2X1_287/B POR2X1_777/B 0.05fF
C41337 PAND2X1_78/m4_208_n4# PAND2X1_772/m4_208_n4# 0.13fF
C41338 POR2X1_590/A POR2X1_214/CTRL 0.01fF
C41339 PAND2X1_557/A PAND2X1_740/a_76_28# 0.01fF
C41340 POR2X1_541/B PAND2X1_111/B 0.03fF
C41341 POR2X1_76/A POR2X1_513/Y 0.03fF
C41342 PAND2X1_826/CTRL PAND2X1_96/B 0.01fF
C41343 POR2X1_411/B PAND2X1_388/Y 0.03fF
C41344 PAND2X1_793/Y POR2X1_487/a_16_28# 0.02fF
C41345 PAND2X1_6/Y POR2X1_84/A 0.18fF
C41346 PAND2X1_406/CTRL PAND2X1_32/B 0.00fF
C41347 PAND2X1_79/CTRL D_INPUT_0 0.01fF
C41348 POR2X1_411/B PAND2X1_549/B 0.03fF
C41349 POR2X1_607/A POR2X1_411/CTRL2 0.00fF
C41350 POR2X1_287/B PAND2X1_65/B 0.00fF
C41351 POR2X1_202/O POR2X1_206/A 0.01fF
C41352 POR2X1_502/A POR2X1_634/CTRL 0.12fF
C41353 POR2X1_341/A POR2X1_222/A 0.07fF
C41354 POR2X1_188/A POR2X1_285/a_76_344# 0.00fF
C41355 PAND2X1_623/a_56_28# POR2X1_615/Y 0.00fF
C41356 POR2X1_72/B POR2X1_372/m4_208_n4# 0.15fF
C41357 POR2X1_50/a_76_344# INPUT_7 0.01fF
C41358 POR2X1_366/O POR2X1_116/A 0.00fF
C41359 POR2X1_315/Y POR2X1_442/CTRL 0.05fF
C41360 POR2X1_194/B PAND2X1_41/B 0.05fF
C41361 PAND2X1_90/A PAND2X1_58/A 0.05fF
C41362 POR2X1_48/A POR2X1_258/CTRL2 0.01fF
C41363 POR2X1_483/A PAND2X1_65/B 0.02fF
C41364 POR2X1_70/O POR2X1_40/Y 0.02fF
C41365 POR2X1_222/Y POR2X1_555/B 0.03fF
C41366 POR2X1_74/CTRL POR2X1_20/B 0.01fF
C41367 PAND2X1_56/Y POR2X1_296/B 0.05fF
C41368 POR2X1_106/CTRL POR2X1_183/Y 0.00fF
C41369 POR2X1_60/A POR2X1_700/O 0.00fF
C41370 POR2X1_278/Y PAND2X1_205/Y 0.03fF
C41371 POR2X1_449/Y VDD 0.00fF
C41372 POR2X1_76/A POR2X1_366/A 0.04fF
C41373 POR2X1_866/A PAND2X1_60/B 0.04fF
C41374 PAND2X1_291/CTRL PAND2X1_93/B 0.01fF
C41375 POR2X1_66/B POR2X1_294/B 0.31fF
C41376 POR2X1_355/B POR2X1_798/CTRL 0.10fF
C41377 PAND2X1_445/O POR2X1_102/Y 0.02fF
C41378 POR2X1_763/Y POR2X1_40/Y 0.03fF
C41379 POR2X1_811/O POR2X1_532/A 0.01fF
C41380 POR2X1_319/A POR2X1_854/B 0.05fF
C41381 POR2X1_155/a_16_28# POR2X1_750/B 0.02fF
C41382 POR2X1_558/B POR2X1_361/CTRL 0.00fF
C41383 POR2X1_523/Y POR2X1_14/Y 0.03fF
C41384 POR2X1_102/Y PAND2X1_723/CTRL2 0.01fF
C41385 POR2X1_188/A POR2X1_294/B 0.03fF
C41386 POR2X1_48/A PAND2X1_350/CTRL 0.09fF
C41387 POR2X1_616/CTRL POR2X1_7/A 0.03fF
C41388 POR2X1_41/B POR2X1_278/O 0.00fF
C41389 POR2X1_329/Y PAND2X1_355/O 0.01fF
C41390 PAND2X1_73/Y PAND2X1_743/a_16_344# 0.02fF
C41391 POR2X1_495/a_56_344# POR2X1_55/Y 0.00fF
C41392 POR2X1_840/O POR2X1_660/Y 0.02fF
C41393 POR2X1_49/Y PAND2X1_724/B 0.07fF
C41394 PAND2X1_280/CTRL PAND2X1_90/Y 0.11fF
C41395 PAND2X1_84/Y INPUT_0 0.03fF
C41396 POR2X1_83/B PAND2X1_370/O 0.02fF
C41397 PAND2X1_659/B PAND2X1_735/CTRL 0.00fF
C41398 PAND2X1_658/CTRL PAND2X1_658/B 0.05fF
C41399 PAND2X1_845/O POR2X1_60/A 0.04fF
C41400 POR2X1_532/A POR2X1_555/B 0.04fF
C41401 POR2X1_130/A PAND2X1_511/CTRL 0.01fF
C41402 POR2X1_41/B POR2X1_122/Y 0.03fF
C41403 POR2X1_43/B POR2X1_39/CTRL2 0.01fF
C41404 POR2X1_614/A POR2X1_864/O 0.06fF
C41405 POR2X1_52/A PAND2X1_828/O 0.11fF
C41406 PAND2X1_23/Y POR2X1_402/CTRL 0.00fF
C41407 POR2X1_849/A POR2X1_550/Y 0.82fF
C41408 POR2X1_76/Y VDD 0.27fF
C41409 PAND2X1_860/A POR2X1_173/CTRL 0.01fF
C41410 POR2X1_56/B POR2X1_511/Y 0.07fF
C41411 POR2X1_274/A POR2X1_260/A 0.03fF
C41412 D_INPUT_0 PAND2X1_28/CTRL2 0.01fF
C41413 POR2X1_532/A PAND2X1_394/CTRL 0.01fF
C41414 POR2X1_57/A POR2X1_102/Y 0.25fF
C41415 PAND2X1_39/B POR2X1_398/CTRL 0.08fF
C41416 POR2X1_329/A POR2X1_761/A 0.00fF
C41417 POR2X1_566/A POR2X1_192/Y 0.83fF
C41418 POR2X1_356/A POR2X1_552/Y 0.03fF
C41419 POR2X1_290/Y PAND2X1_404/A 0.09fF
C41420 POR2X1_68/A POR2X1_402/CTRL2 0.01fF
C41421 POR2X1_523/Y POR2X1_849/CTRL2 0.01fF
C41422 PAND2X1_758/O POR2X1_236/Y 0.03fF
C41423 POR2X1_251/Y POR2X1_13/A 0.02fF
C41424 INPUT_7 POR2X1_587/Y 0.01fF
C41425 PAND2X1_796/B POR2X1_371/CTRL 0.00fF
C41426 POR2X1_383/A POR2X1_296/B 0.27fF
C41427 POR2X1_40/Y POR2X1_73/Y 7.86fF
C41428 D_INPUT_0 POR2X1_276/Y 0.03fF
C41429 PAND2X1_849/B D_INPUT_0 0.03fF
C41430 PAND2X1_90/A PAND2X1_667/O 0.01fF
C41431 PAND2X1_84/Y PAND2X1_717/CTRL2 0.01fF
C41432 POR2X1_818/O POR2X1_294/A 0.03fF
C41433 POR2X1_532/A POR2X1_330/Y 0.11fF
C41434 POR2X1_99/A POR2X1_68/B 0.04fF
C41435 PAND2X1_739/O POR2X1_42/Y 0.07fF
C41436 POR2X1_258/CTRL POR2X1_312/Y 0.06fF
C41437 POR2X1_38/Y POR2X1_72/B 0.77fF
C41438 PAND2X1_265/a_16_344# PAND2X1_60/B 0.02fF
C41439 POR2X1_646/Y POR2X1_101/Y 0.01fF
C41440 PAND2X1_6/Y PAND2X1_65/Y 0.03fF
C41441 PAND2X1_798/B PAND2X1_473/B 0.15fF
C41442 PAND2X1_11/CTRL2 INPUT_5 0.03fF
C41443 POR2X1_96/A POR2X1_7/B 0.19fF
C41444 POR2X1_740/Y VDD 6.44fF
C41445 PAND2X1_615/O POR2X1_94/A 0.15fF
C41446 POR2X1_67/A POR2X1_172/CTRL 0.02fF
C41447 POR2X1_748/A POR2X1_245/O 0.01fF
C41448 POR2X1_447/B PAND2X1_39/B 0.09fF
C41449 POR2X1_15/a_16_28# POR2X1_69/A 0.02fF
C41450 POR2X1_344/CTRL POR2X1_205/A 0.04fF
C41451 PAND2X1_810/A PAND2X1_811/Y 0.14fF
C41452 POR2X1_614/A PAND2X1_263/O 0.16fF
C41453 POR2X1_590/a_16_28# POR2X1_296/B 0.04fF
C41454 POR2X1_214/CTRL POR2X1_214/B 0.01fF
C41455 POR2X1_78/A PAND2X1_373/a_16_344# 0.02fF
C41456 PAND2X1_365/CTRL VDD -0.00fF
C41457 PAND2X1_65/B PAND2X1_59/CTRL2 0.01fF
C41458 POR2X1_614/A D_GATE_865 0.03fF
C41459 POR2X1_215/CTRL POR2X1_741/Y 0.24fF
C41460 PAND2X1_73/CTRL2 PAND2X1_63/B 0.01fF
C41461 POR2X1_590/A POR2X1_362/A 0.00fF
C41462 POR2X1_7/B PAND2X1_335/O 0.15fF
C41463 POR2X1_863/B POR2X1_149/Y 0.00fF
C41464 PAND2X1_830/O POR2X1_60/A 0.15fF
C41465 PAND2X1_48/B POR2X1_651/CTRL 0.01fF
C41466 POR2X1_16/A PAND2X1_404/CTRL2 0.01fF
C41467 PAND2X1_48/B PAND2X1_131/a_76_28# 0.02fF
C41468 POR2X1_193/A POR2X1_579/Y 0.03fF
C41469 PAND2X1_93/B POR2X1_722/CTRL2 0.02fF
C41470 PAND2X1_653/Y PAND2X1_723/Y 0.03fF
C41471 POR2X1_509/A POR2X1_244/B 0.03fF
C41472 POR2X1_90/Y POR2X1_236/Y 0.31fF
C41473 POR2X1_76/Y POR2X1_741/Y 1.85fF
C41474 POR2X1_65/A PAND2X1_241/Y 0.03fF
C41475 POR2X1_502/A D_GATE_222 0.12fF
C41476 PAND2X1_441/a_16_344# PAND2X1_52/B 0.01fF
C41477 POR2X1_614/A POR2X1_471/CTRL 0.01fF
C41478 PAND2X1_76/Y PAND2X1_785/A 0.03fF
C41479 POR2X1_346/B PAND2X1_58/A 0.01fF
C41480 PAND2X1_96/B POR2X1_480/A 0.08fF
C41481 PAND2X1_65/B POR2X1_209/A 0.03fF
C41482 POR2X1_97/a_16_28# POR2X1_97/A 0.01fF
C41483 POR2X1_22/A POR2X1_22/O 0.10fF
C41484 PAND2X1_651/Y PAND2X1_512/Y 0.02fF
C41485 POR2X1_7/B PAND2X1_506/CTRL 0.01fF
C41486 POR2X1_730/Y POR2X1_333/A 0.05fF
C41487 PAND2X1_685/O POR2X1_829/A 0.00fF
C41488 POR2X1_445/CTRL POR2X1_455/A 0.01fF
C41489 POR2X1_59/a_16_28# POR2X1_394/A 0.02fF
C41490 INPUT_4 POR2X1_587/Y 0.07fF
C41491 PAND2X1_244/B POR2X1_40/Y 0.03fF
C41492 POR2X1_78/B PAND2X1_314/CTRL2 0.05fF
C41493 POR2X1_78/A POR2X1_216/Y 0.01fF
C41494 POR2X1_861/O POR2X1_404/Y 0.01fF
C41495 PAND2X1_614/a_76_28# POR2X1_245/Y 0.01fF
C41496 PAND2X1_23/Y POR2X1_662/Y 0.05fF
C41497 POR2X1_244/B POR2X1_631/B 0.03fF
C41498 POR2X1_43/CTRL2 PAND2X1_838/B 0.01fF
C41499 POR2X1_776/A POR2X1_567/CTRL2 0.01fF
C41500 POR2X1_66/A POR2X1_703/O 0.01fF
C41501 POR2X1_502/A PAND2X1_411/a_76_28# 0.01fF
C41502 PAND2X1_645/B VDD 0.19fF
C41503 POR2X1_855/B POR2X1_774/Y 0.02fF
C41504 POR2X1_356/A POR2X1_35/Y 0.05fF
C41505 PAND2X1_659/B POR2X1_73/Y 0.19fF
C41506 PAND2X1_7/CTRL2 POR2X1_222/Y 0.09fF
C41507 PAND2X1_631/CTRL2 POR2X1_293/Y 0.03fF
C41508 POR2X1_376/B PAND2X1_549/B 0.10fF
C41509 POR2X1_41/Y PAND2X1_124/Y 0.06fF
C41510 PAND2X1_783/a_16_344# PAND2X1_779/Y 0.01fF
C41511 POR2X1_76/Y PAND2X1_32/B 0.04fF
C41512 POR2X1_66/A POR2X1_337/Y 0.38fF
C41513 POR2X1_355/B PAND2X1_69/A 0.01fF
C41514 POR2X1_394/A PAND2X1_545/CTRL2 0.05fF
C41515 POR2X1_785/A POR2X1_341/O 0.01fF
C41516 INPUT_0 POR2X1_9/CTRL2 0.03fF
C41517 INPUT_1 PAND2X1_614/CTRL 0.01fF
C41518 INPUT_1 POR2X1_72/B 0.07fF
C41519 INPUT_6 VDD 0.72fF
C41520 POR2X1_278/Y PAND2X1_676/CTRL 0.01fF
C41521 POR2X1_296/B PAND2X1_71/Y 0.03fF
C41522 POR2X1_503/CTRL2 POR2X1_65/A 0.00fF
C41523 POR2X1_614/A POR2X1_193/A 8.50fF
C41524 POR2X1_614/A POR2X1_579/Y 0.03fF
C41525 POR2X1_267/A POR2X1_557/B 0.32fF
C41526 PAND2X1_20/A POR2X1_398/CTRL 0.02fF
C41527 PAND2X1_671/a_16_344# POR2X1_35/B 0.02fF
C41528 PAND2X1_391/a_76_28# POR2X1_384/Y 0.04fF
C41529 PAND2X1_48/B POR2X1_778/B 0.15fF
C41530 PAND2X1_490/CTRL POR2X1_294/B 0.01fF
C41531 PAND2X1_90/Y POR2X1_520/O 0.02fF
C41532 POR2X1_537/Y PAND2X1_73/Y 0.01fF
C41533 POR2X1_383/A POR2X1_547/B 0.03fF
C41534 POR2X1_348/O VDD 0.00fF
C41535 PAND2X1_409/a_16_344# PAND2X1_408/Y 0.02fF
C41536 PAND2X1_409/O POR2X1_407/Y 0.01fF
C41537 PAND2X1_20/A PAND2X1_692/CTRL2 0.01fF
C41538 POR2X1_404/Y POR2X1_500/Y 0.03fF
C41539 POR2X1_7/B POR2X1_386/O 0.02fF
C41540 POR2X1_376/B POR2X1_428/O 0.03fF
C41541 PAND2X1_69/A POR2X1_55/Y 0.03fF
C41542 POR2X1_46/O POR2X1_153/Y 0.04fF
C41543 PAND2X1_150/CTRL POR2X1_404/Y 0.00fF
C41544 POR2X1_390/B POR2X1_362/B 0.03fF
C41545 PAND2X1_90/A PAND2X1_96/B 0.03fF
C41546 POR2X1_72/B POR2X1_153/Y 0.16fF
C41547 POR2X1_677/Y POR2X1_329/A 0.03fF
C41548 POR2X1_247/O POR2X1_532/A 0.01fF
C41549 PAND2X1_48/Y POR2X1_260/A 0.01fF
C41550 PAND2X1_795/O POR2X1_394/A 0.12fF
C41551 POR2X1_806/O POR2X1_737/A 0.01fF
C41552 PAND2X1_341/A POR2X1_55/Y 0.03fF
C41553 POR2X1_740/Y PAND2X1_32/B 0.36fF
C41554 POR2X1_285/B POR2X1_862/A 0.03fF
C41555 POR2X1_296/B POR2X1_788/CTRL 0.06fF
C41556 POR2X1_433/Y POR2X1_56/Y 0.00fF
C41557 PAND2X1_284/Y PAND2X1_555/A 1.72fF
C41558 POR2X1_8/Y POR2X1_381/CTRL2 0.10fF
C41559 POR2X1_538/CTRL PAND2X1_69/A 0.01fF
C41560 PAND2X1_853/CTRL PAND2X1_653/Y 0.03fF
C41561 POR2X1_590/A POR2X1_557/a_16_28# 0.01fF
C41562 PAND2X1_90/Y POR2X1_543/O 0.03fF
C41563 PAND2X1_659/B PAND2X1_244/B 0.01fF
C41564 POR2X1_93/A POR2X1_55/Y 0.24fF
C41565 POR2X1_123/CTRL PAND2X1_60/B 0.01fF
C41566 POR2X1_140/B POR2X1_112/Y 0.04fF
C41567 PAND2X1_698/a_76_28# PAND2X1_65/B 0.01fF
C41568 POR2X1_55/Y POR2X1_91/Y 0.03fF
C41569 POR2X1_566/A POR2X1_568/Y 0.10fF
C41570 PAND2X1_137/Y POR2X1_103/Y 0.01fF
C41571 PAND2X1_737/B VDD 0.05fF
C41572 PAND2X1_857/A POR2X1_829/A 0.03fF
C41573 POR2X1_559/CTRL2 POR2X1_38/B 0.02fF
C41574 POR2X1_52/A PAND2X1_549/B 0.03fF
C41575 POR2X1_7/B POR2X1_7/A 7.43fF
C41576 PAND2X1_810/A PAND2X1_812/A 0.01fF
C41577 POR2X1_150/Y POR2X1_173/Y 0.04fF
C41578 PAND2X1_194/CTRL POR2X1_42/Y 0.01fF
C41579 POR2X1_66/B POR2X1_567/A 0.02fF
C41580 PAND2X1_216/B VDD 0.73fF
C41581 PAND2X1_491/CTRL2 PAND2X1_32/B 0.01fF
C41582 PAND2X1_41/B PAND2X1_48/A 0.12fF
C41583 POR2X1_327/Y POR2X1_830/A 0.09fF
C41584 POR2X1_68/A POR2X1_219/a_16_28# 0.03fF
C41585 POR2X1_81/A POR2X1_83/B 0.62fF
C41586 PAND2X1_787/Y PAND2X1_853/B 1.82fF
C41587 PAND2X1_99/B PAND2X1_333/Y 0.03fF
C41588 PAND2X1_58/A PAND2X1_304/O 0.02fF
C41589 POR2X1_517/CTRL POR2X1_667/A 0.01fF
C41590 POR2X1_268/O POR2X1_39/B 0.02fF
C41591 PAND2X1_48/B POR2X1_854/B 8.49fF
C41592 POR2X1_614/A POR2X1_38/B 8.58fF
C41593 POR2X1_832/B POR2X1_592/O 0.01fF
C41594 PAND2X1_41/B POR2X1_192/B 0.14fF
C41595 POR2X1_57/A POR2X1_531/Y 0.00fF
C41596 POR2X1_188/A POR2X1_567/A 0.01fF
C41597 POR2X1_45/Y PAND2X1_175/B 0.03fF
C41598 POR2X1_71/O PAND2X1_84/Y 0.01fF
C41599 POR2X1_677/Y POR2X1_275/Y 0.00fF
C41600 PAND2X1_709/CTRL2 POR2X1_158/B 0.04fF
C41601 PAND2X1_551/O PAND2X1_551/A 0.02fF
C41602 POR2X1_558/A PAND2X1_494/O 0.00fF
C41603 POR2X1_802/a_16_28# POR2X1_802/B 0.01fF
C41604 POR2X1_285/B PAND2X1_73/Y 0.11fF
C41605 POR2X1_486/B POR2X1_634/A 1.29fF
C41606 POR2X1_774/A VDD 0.56fF
C41607 POR2X1_56/Y PAND2X1_840/CTRL 0.01fF
C41608 PAND2X1_308/CTRL2 POR2X1_56/B 0.02fF
C41609 POR2X1_327/Y POR2X1_532/m4_208_n4# 0.03fF
C41610 PAND2X1_50/O PAND2X1_18/B 0.09fF
C41611 INPUT_6 PAND2X1_32/B 0.01fF
C41612 POR2X1_199/a_56_344# POR2X1_260/A 0.00fF
C41613 POR2X1_102/Y PAND2X1_339/CTRL 0.01fF
C41614 POR2X1_78/B POR2X1_737/A 0.03fF
C41615 PAND2X1_71/Y POR2X1_547/B 0.01fF
C41616 POR2X1_366/Y PAND2X1_313/CTRL 0.02fF
C41617 POR2X1_383/A POR2X1_267/Y 0.00fF
C41618 PAND2X1_359/Y VDD 0.15fF
C41619 POR2X1_502/A POR2X1_544/Y 0.01fF
C41620 POR2X1_532/A POR2X1_148/A 0.01fF
C41621 POR2X1_283/A POR2X1_310/CTRL 0.06fF
C41622 POR2X1_110/Y POR2X1_236/Y 7.84fF
C41623 INPUT_3 PAND2X1_19/Y 0.02fF
C41624 POR2X1_332/B POR2X1_332/a_16_28# 0.05fF
C41625 PAND2X1_150/CTRL2 PAND2X1_60/B 0.02fF
C41626 PAND2X1_79/Y POR2X1_318/A 0.03fF
C41627 PAND2X1_778/CTRL PAND2X1_506/Y 0.00fF
C41628 POR2X1_671/CTRL2 POR2X1_4/Y 0.15fF
C41629 VDD POR2X1_550/B 0.04fF
C41630 POR2X1_68/B POR2X1_380/Y 0.02fF
C41631 POR2X1_83/B PAND2X1_327/O 0.00fF
C41632 POR2X1_336/CTRL2 POR2X1_538/A 0.00fF
C41633 PAND2X1_469/B PAND2X1_353/a_56_28# 0.00fF
C41634 POR2X1_40/Y PAND2X1_207/A 0.03fF
C41635 POR2X1_41/B PAND2X1_508/Y 0.07fF
C41636 POR2X1_285/Y PAND2X1_52/B 1.39fF
C41637 PAND2X1_367/O PAND2X1_366/Y 0.00fF
C41638 PAND2X1_744/CTRL POR2X1_260/A 0.01fF
C41639 POR2X1_391/m4_208_n4# POR2X1_816/A 0.15fF
C41640 POR2X1_643/CTRL POR2X1_260/B 0.01fF
C41641 POR2X1_697/Y POR2X1_394/A 0.00fF
C41642 INPUT_3 PAND2X1_87/O 0.12fF
C41643 POR2X1_739/CTRL POR2X1_568/Y 0.35fF
C41644 PAND2X1_559/O POR2X1_73/Y 0.09fF
C41645 PAND2X1_73/Y POR2X1_579/CTRL 0.01fF
C41646 PAND2X1_484/O POR2X1_294/B 0.07fF
C41647 PAND2X1_373/CTRL POR2X1_540/A 0.00fF
C41648 POR2X1_119/Y PAND2X1_549/O 0.02fF
C41649 POR2X1_376/A PAND2X1_63/B 0.00fF
C41650 POR2X1_844/B POR2X1_546/CTRL2 0.01fF
C41651 PAND2X1_452/A POR2X1_425/Y 0.07fF
C41652 POR2X1_750/B PAND2X1_681/CTRL2 0.01fF
C41653 POR2X1_68/A POR2X1_507/A 0.01fF
C41654 POR2X1_5/Y POR2X1_372/CTRL2 0.01fF
C41655 POR2X1_571/CTRL2 POR2X1_844/B 0.01fF
C41656 POR2X1_346/B PAND2X1_96/B 0.07fF
C41657 PAND2X1_191/O PAND2X1_730/A 0.00fF
C41658 PAND2X1_569/A PAND2X1_569/O 0.00fF
C41659 PAND2X1_715/B POR2X1_310/O 0.00fF
C41660 POR2X1_798/CTRL2 PAND2X1_52/B 0.01fF
C41661 POR2X1_802/a_16_28# POR2X1_532/A 0.03fF
C41662 POR2X1_730/Y POR2X1_788/B 0.03fF
C41663 PAND2X1_863/B PAND2X1_729/O 0.02fF
C41664 POR2X1_574/Y POR2X1_515/Y 0.01fF
C41665 POR2X1_52/A PAND2X1_330/CTRL -0.00fF
C41666 PAND2X1_643/A PAND2X1_364/B 0.03fF
C41667 PAND2X1_857/A PAND2X1_857/B 0.14fF
C41668 PAND2X1_171/CTRL D_GATE_741 0.01fF
C41669 POR2X1_83/B POR2X1_234/A 0.18fF
C41670 INPUT_0 PAND2X1_136/a_16_344# 0.02fF
C41671 POR2X1_119/Y POR2X1_119/O 0.02fF
C41672 PAND2X1_346/O POR2X1_295/Y 0.15fF
C41673 POR2X1_122/Y POR2X1_77/Y 0.03fF
C41674 POR2X1_68/A POR2X1_266/A 0.03fF
C41675 PAND2X1_127/CTRL POR2X1_318/A 0.08fF
C41676 POR2X1_796/A POR2X1_725/Y 0.02fF
C41677 POR2X1_16/A PAND2X1_216/m4_208_n4# 0.06fF
C41678 POR2X1_343/Y POR2X1_778/O 0.04fF
C41679 PAND2X1_803/O POR2X1_90/Y 0.17fF
C41680 POR2X1_702/A POR2X1_332/a_76_344# 0.03fF
C41681 POR2X1_730/Y PAND2X1_163/CTRL 0.01fF
C41682 PAND2X1_108/CTRL VDD -0.00fF
C41683 POR2X1_774/A PAND2X1_32/B 0.03fF
C41684 PAND2X1_61/a_16_344# POR2X1_9/Y 0.02fF
C41685 POR2X1_57/A POR2X1_165/Y 0.01fF
C41686 PAND2X1_72/CTRL PAND2X1_48/A 0.01fF
C41687 POR2X1_327/Y POR2X1_596/A 0.23fF
C41688 POR2X1_294/B POR2X1_199/B 0.01fF
C41689 D_INPUT_1 PAND2X1_527/O 0.04fF
C41690 POR2X1_51/A POR2X1_416/B 0.01fF
C41691 PAND2X1_140/A POR2X1_394/A 0.03fF
C41692 POR2X1_383/A POR2X1_590/Y 0.07fF
C41693 POR2X1_776/B POR2X1_567/O 0.02fF
C41694 POR2X1_657/Y POR2X1_222/O 0.02fF
C41695 POR2X1_528/Y POR2X1_394/A 0.01fF
C41696 PAND2X1_514/CTRL2 PAND2X1_348/A 0.01fF
C41697 PAND2X1_755/O PAND2X1_72/A 0.03fF
C41698 POR2X1_67/Y POR2X1_29/A 0.06fF
C41699 PAND2X1_563/A PAND2X1_346/Y 0.03fF
C41700 POR2X1_83/B POR2X1_667/CTRL2 0.00fF
C41701 POR2X1_62/Y PAND2X1_350/CTRL 0.01fF
C41702 POR2X1_102/CTRL2 INPUT_2 0.01fF
C41703 POR2X1_87/B VDD 0.38fF
C41704 POR2X1_102/CTRL D_INPUT_1 0.01fF
C41705 PAND2X1_20/A PAND2X1_607/a_76_28# 0.01fF
C41706 POR2X1_736/A PAND2X1_178/O 0.04fF
C41707 POR2X1_16/A PAND2X1_704/CTRL 0.01fF
C41708 PAND2X1_773/m4_208_n4# POR2X1_767/m4_208_n4# 0.13fF
C41709 PAND2X1_773/CTRL POR2X1_767/Y 0.01fF
C41710 POR2X1_652/Y PAND2X1_72/A 0.01fF
C41711 POR2X1_144/Y PAND2X1_147/O 0.00fF
C41712 PAND2X1_57/B PAND2X1_135/O 0.01fF
C41713 POR2X1_110/Y POR2X1_111/a_16_28# 0.03fF
C41714 PAND2X1_643/CTRL POR2X1_416/B 0.01fF
C41715 POR2X1_48/A POR2X1_253/O 0.02fF
C41716 POR2X1_48/A PAND2X1_750/O 0.01fF
C41717 PAND2X1_348/O PAND2X1_345/Y -0.00fF
C41718 POR2X1_593/CTRL2 POR2X1_449/A 0.01fF
C41719 POR2X1_49/Y POR2X1_441/CTRL2 0.01fF
C41720 POR2X1_688/O POR2X1_121/B 0.02fF
C41721 PAND2X1_661/Y PAND2X1_120/m4_208_n4# 0.09fF
C41722 POR2X1_57/A POR2X1_761/A 0.03fF
C41723 PAND2X1_94/A POR2X1_113/B 0.05fF
C41724 POR2X1_673/Y POR2X1_550/B 0.03fF
C41725 POR2X1_509/O POR2X1_35/Y 0.01fF
C41726 POR2X1_212/A POR2X1_220/B 0.01fF
C41727 POR2X1_35/Y PAND2X1_72/A 0.03fF
C41728 PAND2X1_631/A PAND2X1_514/CTRL2 0.02fF
C41729 POR2X1_257/A POR2X1_496/Y 0.03fF
C41730 POR2X1_287/B POR2X1_814/A 0.10fF
C41731 POR2X1_73/a_76_344# PAND2X1_341/B 0.00fF
C41732 POR2X1_545/CTRL2 POR2X1_551/A 0.01fF
C41733 PAND2X1_67/CTRL2 POR2X1_296/B 0.00fF
C41734 POR2X1_322/Y POR2X1_39/B 0.07fF
C41735 POR2X1_389/A PAND2X1_56/A 0.03fF
C41736 PAND2X1_856/B PAND2X1_854/Y 0.70fF
C41737 POR2X1_63/Y POR2X1_60/A 0.06fF
C41738 POR2X1_825/CTRL2 POR2X1_20/B 0.01fF
C41739 POR2X1_715/CTRL POR2X1_702/A 0.00fF
C41740 PAND2X1_129/CTRL POR2X1_814/A 0.01fF
C41741 POR2X1_814/A POR2X1_778/CTRL 0.01fF
C41742 POR2X1_243/A POR2X1_243/B 0.35fF
C41743 POR2X1_568/Y POR2X1_568/CTRL2 0.02fF
C41744 POR2X1_77/O POR2X1_83/B 0.18fF
C41745 POR2X1_87/B PAND2X1_32/B 0.21fF
C41746 POR2X1_643/CTRL PAND2X1_55/Y 0.03fF
C41747 PAND2X1_612/B PAND2X1_20/A 0.03fF
C41748 POR2X1_754/CTRL2 POR2X1_39/B 0.03fF
C41749 POR2X1_452/Y POR2X1_330/Y 0.01fF
C41750 POR2X1_461/Y PAND2X1_41/B 0.03fF
C41751 POR2X1_423/Y POR2X1_253/CTRL 0.01fF
C41752 POR2X1_651/Y POR2X1_712/Y 0.03fF
C41753 POR2X1_278/Y POR2X1_329/A 0.05fF
C41754 POR2X1_67/Y POR2X1_546/A 0.01fF
C41755 POR2X1_634/A POR2X1_610/CTRL2 0.01fF
C41756 POR2X1_130/A POR2X1_646/B 0.04fF
C41757 POR2X1_482/CTRL2 POR2X1_669/B 0.03fF
C41758 POR2X1_814/A PAND2X1_89/CTRL 0.07fF
C41759 POR2X1_123/A PAND2X1_72/A 0.01fF
C41760 POR2X1_304/CTRL POR2X1_153/Y 0.03fF
C41761 POR2X1_67/Y PAND2X1_754/O 0.03fF
C41762 PAND2X1_834/CTRL2 POR2X1_153/Y 0.05fF
C41763 POR2X1_446/B POR2X1_186/Y 0.03fF
C41764 PAND2X1_272/CTRL POR2X1_296/B 0.01fF
C41765 POR2X1_707/B PAND2X1_59/B 0.01fF
C41766 POR2X1_98/O POR2X1_590/A 0.16fF
C41767 POR2X1_41/B PAND2X1_464/B 0.02fF
C41768 POR2X1_65/A POR2X1_253/a_16_28# 0.01fF
C41769 POR2X1_20/B PAND2X1_347/Y 0.03fF
C41770 PAND2X1_147/CTRL2 POR2X1_142/Y 0.01fF
C41771 PAND2X1_475/CTRL2 D_INPUT_0 0.06fF
C41772 POR2X1_433/O POR2X1_37/Y 0.02fF
C41773 POR2X1_736/A POR2X1_741/B 0.03fF
C41774 POR2X1_48/A PAND2X1_820/B 0.00fF
C41775 POR2X1_624/Y POR2X1_5/Y 0.03fF
C41776 POR2X1_263/CTRL2 PAND2X1_35/Y 0.01fF
C41777 POR2X1_760/A POR2X1_7/B 0.05fF
C41778 POR2X1_168/O POR2X1_191/Y 0.01fF
C41779 PAND2X1_255/O POR2X1_786/Y 0.24fF
C41780 POR2X1_150/Y PAND2X1_735/Y 0.00fF
C41781 POR2X1_389/A POR2X1_661/A 1.24fF
C41782 POR2X1_46/CTRL2 POR2X1_409/B 0.01fF
C41783 PAND2X1_609/CTRL2 PAND2X1_90/Y 0.09fF
C41784 POR2X1_351/m4_208_n4# PAND2X1_72/A 0.17fF
C41785 PAND2X1_435/O POR2X1_20/B 0.03fF
C41786 POR2X1_102/Y PAND2X1_215/CTRL2 0.01fF
C41787 POR2X1_812/A PAND2X1_73/Y 0.01fF
C41788 PAND2X1_508/Y POR2X1_77/Y 0.03fF
C41789 POR2X1_769/CTRL2 PAND2X1_52/B 0.03fF
C41790 POR2X1_541/B PAND2X1_48/a_76_28# 0.01fF
C41791 PAND2X1_21/O PAND2X1_26/A 0.02fF
C41792 POR2X1_525/O POR2X1_23/Y 0.09fF
C41793 POR2X1_660/Y POR2X1_330/Y 0.05fF
C41794 PAND2X1_458/O POR2X1_91/Y 0.08fF
C41795 PAND2X1_39/B POR2X1_220/Y 0.10fF
C41796 POR2X1_257/A PAND2X1_804/B 0.03fF
C41797 PAND2X1_381/Y POR2X1_750/B 0.03fF
C41798 POR2X1_502/A POR2X1_54/Y 0.03fF
C41799 POR2X1_227/CTRL PAND2X1_52/B 0.01fF
C41800 POR2X1_150/Y PAND2X1_493/Y 0.88fF
C41801 PAND2X1_318/O POR2X1_20/B 0.22fF
C41802 POR2X1_23/Y PAND2X1_787/Y 0.00fF
C41803 POR2X1_49/Y POR2X1_496/Y 0.07fF
C41804 POR2X1_415/A POR2X1_415/a_16_28# 0.01fF
C41805 PAND2X1_769/Y VDD 0.00fF
C41806 POR2X1_18/CTRL2 D_INPUT_6 0.01fF
C41807 POR2X1_306/CTRL POR2X1_329/A 0.04fF
C41808 PAND2X1_39/B POR2X1_404/Y 0.03fF
C41809 POR2X1_636/CTRL POR2X1_750/B 0.01fF
C41810 POR2X1_38/a_16_28# POR2X1_5/Y 0.01fF
C41811 POR2X1_376/B PAND2X1_68/O 0.05fF
C41812 PAND2X1_841/O POR2X1_411/B 0.02fF
C41813 POR2X1_841/O POR2X1_733/A 0.04fF
C41814 POR2X1_13/A PAND2X1_410/O 0.04fF
C41815 POR2X1_66/B POR2X1_643/A 0.06fF
C41816 PAND2X1_20/A POR2X1_141/Y 0.03fF
C41817 POR2X1_479/B POR2X1_476/Y 0.02fF
C41818 POR2X1_423/Y POR2X1_516/Y 0.01fF
C41819 POR2X1_260/B PAND2X1_751/CTRL2 0.03fF
C41820 PAND2X1_622/O POR2X1_29/A 0.03fF
C41821 POR2X1_16/A PAND2X1_403/CTRL 0.01fF
C41822 POR2X1_476/Y PAND2X1_595/O 0.17fF
C41823 POR2X1_804/CTRL2 POR2X1_435/Y 0.05fF
C41824 POR2X1_820/Y POR2X1_48/A 0.03fF
C41825 POR2X1_257/A PAND2X1_514/Y 0.10fF
C41826 PAND2X1_58/A POR2X1_402/CTRL2 0.00fF
C41827 POR2X1_411/B PAND2X1_570/O 0.05fF
C41828 POR2X1_188/A POR2X1_643/A 0.00fF
C41829 PAND2X1_214/A POR2X1_72/B 0.01fF
C41830 PAND2X1_105/a_16_344# POR2X1_411/B 0.02fF
C41831 POR2X1_602/CTRL2 POR2X1_294/B 0.03fF
C41832 POR2X1_487/CTRL PAND2X1_580/B 0.00fF
C41833 POR2X1_274/A PAND2X1_516/a_76_28# 0.01fF
C41834 POR2X1_831/CTRL2 POR2X1_513/Y 0.03fF
C41835 PAND2X1_717/A POR2X1_283/A 0.08fF
C41836 PAND2X1_48/B POR2X1_862/A 0.07fF
C41837 PAND2X1_206/B POR2X1_7/A 0.11fF
C41838 POR2X1_843/m4_208_n4# POR2X1_343/A 0.01fF
C41839 POR2X1_843/a_16_28# POR2X1_287/B 0.00fF
C41840 PAND2X1_750/CTRL POR2X1_816/A 0.01fF
C41841 POR2X1_49/Y PAND2X1_733/A 0.03fF
C41842 POR2X1_832/Y PAND2X1_55/Y 0.06fF
C41843 POR2X1_624/Y PAND2X1_316/CTRL 0.01fF
C41844 PAND2X1_3/A INPUT_4 0.06fF
C41845 PAND2X1_849/CTRL2 POR2X1_60/Y 0.01fF
C41846 POR2X1_23/Y POR2X1_256/a_76_344# 0.03fF
C41847 POR2X1_20/B POR2X1_245/CTRL2 0.03fF
C41848 INPUT_0 POR2X1_296/B 0.08fF
C41849 POR2X1_257/A PAND2X1_324/CTRL 0.01fF
C41850 POR2X1_149/CTRL POR2X1_532/A 0.00fF
C41851 POR2X1_102/Y PAND2X1_84/Y 0.03fF
C41852 POR2X1_188/A POR2X1_807/A 0.02fF
C41853 POR2X1_313/Y PAND2X1_439/CTRL 0.01fF
C41854 PAND2X1_58/A POR2X1_459/CTRL2 0.00fF
C41855 POR2X1_639/a_16_28# POR2X1_750/B 0.03fF
C41856 POR2X1_241/B POR2X1_192/Y 0.05fF
C41857 PAND2X1_411/O POR2X1_260/B 0.04fF
C41858 POR2X1_630/CTRL POR2X1_222/Y 0.00fF
C41859 PAND2X1_272/O POR2X1_465/B 0.10fF
C41860 PAND2X1_23/Y POR2X1_444/A 0.09fF
C41861 POR2X1_16/A POR2X1_250/Y 0.07fF
C41862 POR2X1_193/Y PAND2X1_41/B 0.03fF
C41863 POR2X1_141/Y POR2X1_325/A 0.03fF
C41864 PAND2X1_804/A POR2X1_40/Y 0.09fF
C41865 POR2X1_65/A POR2X1_106/Y 0.03fF
C41866 PAND2X1_20/A POR2X1_220/Y 0.03fF
C41867 POR2X1_78/B POR2X1_302/B 0.03fF
C41868 POR2X1_45/Y POR2X1_409/B 0.00fF
C41869 POR2X1_590/A POR2X1_579/Y 0.03fF
C41870 PAND2X1_487/O PAND2X1_96/B 0.04fF
C41871 POR2X1_207/O POR2X1_330/Y 0.01fF
C41872 PAND2X1_48/B PAND2X1_73/Y 0.17fF
C41873 POR2X1_697/Y POR2X1_669/B 0.04fF
C41874 POR2X1_632/A POR2X1_61/Y 0.01fF
C41875 POR2X1_260/B POR2X1_68/B 0.03fF
C41876 POR2X1_415/A POR2X1_408/Y 0.10fF
C41877 POR2X1_48/A PAND2X1_506/a_76_28# 0.01fF
C41878 POR2X1_311/Y POR2X1_7/B 0.32fF
C41879 POR2X1_99/A POR2X1_243/Y 0.25fF
C41880 PAND2X1_20/A POR2X1_404/Y 0.03fF
C41881 POR2X1_20/B PAND2X1_346/Y 0.13fF
C41882 PAND2X1_59/B PAND2X1_26/CTRL2 0.03fF
C41883 POR2X1_20/B PAND2X1_100/CTRL 0.00fF
C41884 POR2X1_65/A PAND2X1_580/B 0.03fF
C41885 POR2X1_603/Y POR2X1_42/Y 0.12fF
C41886 PAND2X1_669/CTRL POR2X1_816/A 0.01fF
C41887 POR2X1_677/CTRL INPUT_0 0.05fF
C41888 POR2X1_476/A PAND2X1_69/A 0.07fF
C41889 POR2X1_596/A POR2X1_644/Y 0.04fF
C41890 PAND2X1_473/Y PAND2X1_576/O 0.01fF
C41891 PAND2X1_736/A POR2X1_674/Y 0.03fF
C41892 PAND2X1_648/O PAND2X1_645/Y 0.02fF
C41893 PAND2X1_669/CTRL D_INPUT_1 0.02fF
C41894 POR2X1_305/Y POR2X1_32/A 0.02fF
C41895 PAND2X1_36/CTRL2 PAND2X1_32/B 0.01fF
C41896 POR2X1_66/B POR2X1_138/CTRL2 0.01fF
C41897 POR2X1_804/a_16_28# POR2X1_804/B 0.01fF
C41898 POR2X1_43/B PAND2X1_244/CTRL2 0.03fF
C41899 INPUT_1 PAND2X1_247/CTRL 0.01fF
C41900 POR2X1_48/A POR2X1_280/CTRL 0.03fF
C41901 POR2X1_244/B POR2X1_61/Y 0.03fF
C41902 POR2X1_789/A POR2X1_590/A 0.03fF
C41903 POR2X1_88/O POR2X1_7/A 0.01fF
C41904 PAND2X1_456/CTRL PAND2X1_254/Y 0.01fF
C41905 POR2X1_121/A POR2X1_121/B 3.12fF
C41906 POR2X1_814/B POR2X1_220/Y 0.03fF
C41907 POR2X1_96/A PAND2X1_220/Y 0.13fF
C41908 POR2X1_614/A POR2X1_590/A 0.13fF
C41909 PAND2X1_459/Y POR2X1_5/Y 0.00fF
C41910 POR2X1_407/A POR2X1_390/O 0.00fF
C41911 INPUT_1 PAND2X1_407/CTRL2 0.01fF
C41912 INPUT_0 POR2X1_236/Y 0.57fF
C41913 POR2X1_477/A POR2X1_675/a_16_28# 0.01fF
C41914 POR2X1_814/B POR2X1_404/Y 0.05fF
C41915 POR2X1_66/B POR2X1_140/B 0.02fF
C41916 POR2X1_49/Y PAND2X1_454/O 0.24fF
C41917 POR2X1_445/A POR2X1_456/B 0.75fF
C41918 POR2X1_383/A PAND2X1_237/O 0.04fF
C41919 POR2X1_590/A POR2X1_38/B 0.21fF
C41920 POR2X1_102/Y POR2X1_239/CTRL 0.01fF
C41921 POR2X1_66/B POR2X1_407/A 0.03fF
C41922 POR2X1_262/m4_208_n4# POR2X1_7/Y 0.07fF
C41923 POR2X1_251/O PAND2X1_190/Y 0.01fF
C41924 POR2X1_220/Y POR2X1_325/A 0.03fF
C41925 PAND2X1_6/Y POR2X1_244/CTRL2 0.01fF
C41926 PAND2X1_220/a_16_344# POR2X1_417/Y 0.02fF
C41927 PAND2X1_296/m4_208_n4# PAND2X1_349/m4_208_n4# 0.13fF
C41928 POR2X1_186/Y POR2X1_795/B 0.07fF
C41929 POR2X1_66/B PAND2X1_252/CTRL2 0.03fF
C41930 POR2X1_538/A POR2X1_66/A 0.06fF
C41931 PAND2X1_39/B PAND2X1_399/CTRL 0.01fF
C41932 PAND2X1_407/CTRL2 POR2X1_153/Y 0.05fF
C41933 POR2X1_270/Y PAND2X1_368/CTRL 0.01fF
C41934 POR2X1_16/A POR2X1_490/Y 0.05fF
C41935 POR2X1_188/A POR2X1_407/A 0.03fF
C41936 PAND2X1_229/CTRL D_GATE_222 0.04fF
C41937 PAND2X1_449/Y POR2X1_72/B 0.10fF
C41938 GATE_479 PAND2X1_546/Y 0.05fF
C41939 PAND2X1_214/a_76_28# PAND2X1_656/A 0.01fF
C41940 POR2X1_96/A PAND2X1_739/Y 0.01fF
C41941 POR2X1_43/B PAND2X1_474/A 8.39fF
C41942 POR2X1_32/Y POR2X1_27/Y 0.08fF
C41943 POR2X1_13/A POR2X1_13/a_76_344# 0.02fF
C41944 POR2X1_264/Y PAND2X1_65/B 0.11fF
C41945 PAND2X1_658/A POR2X1_5/Y 0.05fF
C41946 PAND2X1_552/A PAND2X1_552/B 0.06fF
C41947 POR2X1_14/Y PAND2X1_338/B 0.05fF
C41948 PAND2X1_74/a_16_344# POR2X1_532/A 0.01fF
C41949 POR2X1_847/B PAND2X1_6/A 0.12fF
C41950 PAND2X1_827/CTRL2 POR2X1_507/A 0.03fF
C41951 PAND2X1_293/CTRL2 PAND2X1_55/Y 0.01fF
C41952 PAND2X1_573/CTRL2 POR2X1_494/Y 0.00fF
C41953 POR2X1_66/Y POR2X1_294/A 0.21fF
C41954 POR2X1_440/Y POR2X1_590/A 0.03fF
C41955 POR2X1_45/Y POR2X1_272/Y 0.06fF
C41956 POR2X1_72/B POR2X1_591/Y 0.03fF
C41957 POR2X1_632/A POR2X1_35/Y 0.00fF
C41958 POR2X1_423/Y PAND2X1_702/O 0.02fF
C41959 POR2X1_69/CTRL2 POR2X1_7/A 0.01fF
C41960 PAND2X1_96/B POR2X1_402/CTRL2 0.03fF
C41961 POR2X1_817/O POR2X1_394/A 0.08fF
C41962 POR2X1_16/A PAND2X1_561/O 0.14fF
C41963 POR2X1_712/A PAND2X1_90/Y 0.06fF
C41964 POR2X1_40/Y POR2X1_511/O 0.02fF
C41965 PAND2X1_218/O VDD 0.00fF
C41966 POR2X1_558/O INPUT_0 0.09fF
C41967 POR2X1_606/CTRL POR2X1_294/A 0.01fF
C41968 POR2X1_280/O POR2X1_312/Y 0.01fF
C41969 POR2X1_41/B POR2X1_525/Y 0.01fF
C41970 PAND2X1_640/B POR2X1_153/Y 0.01fF
C41971 PAND2X1_464/B POR2X1_77/Y 0.03fF
C41972 D_INPUT_3 POR2X1_293/CTRL 0.01fF
C41973 PAND2X1_190/Y PAND2X1_580/B 0.03fF
C41974 POR2X1_859/A POR2X1_415/Y 0.17fF
C41975 POR2X1_56/B POR2X1_293/Y 0.10fF
C41976 POR2X1_167/a_16_28# POR2X1_669/B 0.05fF
C41977 POR2X1_332/B POR2X1_222/Y 0.03fF
C41978 POR2X1_40/Y PAND2X1_656/A 0.03fF
C41979 POR2X1_5/Y POR2X1_73/Y 0.11fF
C41980 POR2X1_857/B POR2X1_579/Y 0.05fF
C41981 POR2X1_307/Y PAND2X1_55/Y 0.03fF
C41982 POR2X1_459/B VDD 0.10fF
C41983 POR2X1_23/Y PAND2X1_708/O 0.05fF
C41984 POR2X1_750/B POR2X1_7/A 0.03fF
C41985 PAND2X1_218/CTRL2 PAND2X1_364/B 0.02fF
C41986 POR2X1_244/B POR2X1_35/Y 0.07fF
C41987 PAND2X1_41/B PAND2X1_670/O 0.01fF
C41988 POR2X1_327/Y D_INPUT_0 0.06fF
C41989 INPUT_0 POR2X1_267/Y 0.02fF
C41990 POR2X1_557/A PAND2X1_20/A 0.03fF
C41991 PAND2X1_440/CTRL2 POR2X1_150/Y 0.01fF
C41992 POR2X1_564/Y POR2X1_545/A 0.34fF
C41993 POR2X1_383/A POR2X1_186/Y 0.17fF
C41994 PAND2X1_793/Y PAND2X1_798/B 0.25fF
C41995 POR2X1_43/B POR2X1_275/CTRL2 0.00fF
C41996 POR2X1_638/Y VDD 0.37fF
C41997 PAND2X1_65/B POR2X1_712/CTRL 0.01fF
C41998 POR2X1_196/Y VDD 0.25fF
C41999 POR2X1_193/Y POR2X1_228/Y 0.35fF
C42000 PAND2X1_20/A POR2X1_546/CTRL 0.01fF
C42001 POR2X1_96/A PAND2X1_631/CTRL 0.01fF
C42002 POR2X1_65/A PAND2X1_349/A 0.03fF
C42003 POR2X1_290/Y PAND2X1_334/O 0.02fF
C42004 PAND2X1_57/B PAND2X1_743/CTRL -0.00fF
C42005 INPUT_0 PAND2X1_858/Y 0.01fF
C42006 PAND2X1_254/Y POR2X1_56/Y 0.01fF
C42007 POR2X1_539/CTRL POR2X1_750/B 0.00fF
C42008 POR2X1_66/B POR2X1_537/CTRL 0.00fF
C42009 PAND2X1_58/A POR2X1_507/A 0.01fF
C42010 PAND2X1_20/A POR2X1_571/CTRL 0.01fF
C42011 POR2X1_633/O PAND2X1_52/B 0.01fF
C42012 POR2X1_462/B POR2X1_790/CTRL 0.01fF
C42013 POR2X1_750/B POR2X1_703/A 5.71fF
C42014 PAND2X1_857/CTRL POR2X1_23/Y 0.01fF
C42015 PAND2X1_738/Y PAND2X1_113/O 0.29fF
C42016 PAND2X1_748/CTRL POR2X1_752/Y 0.00fF
C42017 PAND2X1_778/O POR2X1_387/Y 0.07fF
C42018 POR2X1_853/A POR2X1_563/Y 0.59fF
C42019 POR2X1_57/A POR2X1_278/Y 0.10fF
C42020 POR2X1_537/CTRL POR2X1_188/A 0.01fF
C42021 PAND2X1_48/B PAND2X1_145/a_56_28# 0.00fF
C42022 POR2X1_750/Y PAND2X1_526/CTRL 0.25fF
C42023 PAND2X1_244/B POR2X1_5/Y 0.03fF
C42024 PAND2X1_354/A PAND2X1_563/A 0.03fF
C42025 POR2X1_40/Y PAND2X1_348/A 0.14fF
C42026 PAND2X1_48/B POR2X1_631/B 0.03fF
C42027 PAND2X1_773/a_56_28# POR2X1_7/B 0.00fF
C42028 POR2X1_502/A POR2X1_544/O 0.02fF
C42029 PAND2X1_115/B POR2X1_310/O 0.02fF
C42030 PAND2X1_650/CTRL2 POR2X1_46/Y 0.01fF
C42031 PAND2X1_90/Y POR2X1_407/O 0.04fF
C42032 POR2X1_49/Y PAND2X1_480/CTRL 0.01fF
C42033 PAND2X1_23/Y POR2X1_804/A 1.32fF
C42034 POR2X1_575/B POR2X1_576/Y 0.03fF
C42035 POR2X1_57/A POR2X1_829/A 0.03fF
C42036 POR2X1_38/Y POR2X1_7/B 0.08fF
C42037 VDD POR2X1_169/Y -0.00fF
C42038 POR2X1_853/A POR2X1_211/O 0.02fF
C42039 PAND2X1_124/Y POR2X1_39/B 0.04fF
C42040 POR2X1_469/CTRL2 POR2X1_478/B 0.00fF
C42041 PAND2X1_126/m4_208_n4# POR2X1_5/Y 0.09fF
C42042 PAND2X1_55/Y POR2X1_68/B 0.17fF
C42043 POR2X1_301/a_16_28# PAND2X1_23/Y 0.03fF
C42044 POR2X1_68/A POR2X1_786/Y 0.10fF
C42045 POR2X1_383/A POR2X1_483/O 0.07fF
C42046 POR2X1_335/CTRL2 POR2X1_260/A 0.00fF
C42047 POR2X1_196/Y POR2X1_741/Y 0.05fF
C42048 POR2X1_305/Y PAND2X1_651/Y 0.02fF
C42049 POR2X1_635/A PAND2X1_72/A 0.16fF
C42050 VDD POR2X1_352/CTRL 0.00fF
C42051 POR2X1_750/Y VDD 0.49fF
C42052 POR2X1_41/B POR2X1_283/A 2.26fF
C42053 POR2X1_618/CTRL POR2X1_7/A 0.02fF
C42054 POR2X1_722/B POR2X1_832/A 0.01fF
C42055 POR2X1_663/CTRL2 POR2X1_544/B 0.01fF
C42056 POR2X1_572/B POR2X1_361/CTRL 0.01fF
C42057 POR2X1_68/A POR2X1_788/B 0.03fF
C42058 PAND2X1_784/O POR2X1_387/Y 0.08fF
C42059 PAND2X1_90/Y POR2X1_317/B 0.88fF
C42060 PAND2X1_69/A POR2X1_513/Y 0.03fF
C42061 POR2X1_515/CTRL2 POR2X1_574/Y 0.01fF
C42062 POR2X1_394/A PAND2X1_712/B 0.01fF
C42063 POR2X1_402/A POR2X1_68/B 0.04fF
C42064 D_INPUT_3 PAND2X1_341/a_16_344# 0.04fF
C42065 POR2X1_327/Y PAND2X1_90/Y 0.13fF
C42066 PAND2X1_20/A POR2X1_554/CTRL 0.01fF
C42067 PAND2X1_496/CTRL POR2X1_569/A 0.05fF
C42068 POR2X1_687/A PAND2X1_760/a_76_28# 0.05fF
C42069 POR2X1_796/A POR2X1_783/B 0.00fF
C42070 PAND2X1_831/Y POR2X1_184/Y 0.02fF
C42071 POR2X1_135/CTRL POR2X1_423/Y 0.01fF
C42072 PAND2X1_631/A POR2X1_40/Y 0.07fF
C42073 PAND2X1_678/O POR2X1_677/Y 0.02fF
C42074 POR2X1_651/Y PAND2X1_39/B 0.03fF
C42075 D_GATE_222 POR2X1_510/Y 0.03fF
C42076 POR2X1_646/Y POR2X1_711/Y 0.07fF
C42077 POR2X1_219/CTRL PAND2X1_88/Y 0.01fF
C42078 POR2X1_333/A POR2X1_169/A 0.03fF
C42079 INPUT_1 POR2X1_7/B 0.19fF
C42080 POR2X1_83/B POR2X1_39/B 0.33fF
C42081 POR2X1_205/A PAND2X1_69/A 0.07fF
C42082 PAND2X1_190/Y PAND2X1_349/A 0.05fF
C42083 PAND2X1_65/B POR2X1_502/Y 0.05fF
C42084 POR2X1_16/A PAND2X1_243/B 0.01fF
C42085 PAND2X1_216/B PAND2X1_216/O 0.00fF
C42086 POR2X1_86/CTRL POR2X1_40/Y 0.01fF
C42087 POR2X1_41/B POR2X1_385/a_16_28# 0.01fF
C42088 PAND2X1_825/CTRL2 POR2X1_402/A 0.01fF
C42089 POR2X1_371/CTRL POR2X1_372/A 0.01fF
C42090 POR2X1_244/B POR2X1_227/CTRL2 0.01fF
C42091 POR2X1_165/CTRL POR2X1_73/Y 0.01fF
C42092 POR2X1_119/Y PAND2X1_76/Y 0.15fF
C42093 POR2X1_96/A PAND2X1_560/B 0.03fF
C42094 PAND2X1_389/O POR2X1_387/Y 0.12fF
C42095 POR2X1_565/B POR2X1_6/CTRL 0.00fF
C42096 PAND2X1_442/O POR2X1_191/Y 0.09fF
C42097 PAND2X1_442/a_16_344# POR2X1_192/B 0.02fF
C42098 PAND2X1_25/O PAND2X1_52/B 0.01fF
C42099 POR2X1_65/A POR2X1_86/CTRL2 -0.00fF
C42100 POR2X1_186/CTRL PAND2X1_55/Y -0.00fF
C42101 PAND2X1_691/Y POR2X1_665/Y 0.05fF
C42102 POR2X1_855/B POR2X1_796/a_76_344# 0.00fF
C42103 POR2X1_78/O POR2X1_569/A 0.01fF
C42104 POR2X1_280/Y PAND2X1_566/Y 0.01fF
C42105 POR2X1_7/B POR2X1_153/Y 0.69fF
C42106 PAND2X1_60/B POR2X1_140/O 0.13fF
C42107 POR2X1_677/Y POR2X1_271/CTRL2 0.00fF
C42108 POR2X1_463/a_16_28# POR2X1_460/Y 0.02fF
C42109 POR2X1_719/CTRL2 PAND2X1_60/B 0.01fF
C42110 POR2X1_166/a_16_28# POR2X1_73/Y 0.02fF
C42111 POR2X1_23/Y POR2X1_825/Y 0.00fF
C42112 POR2X1_447/B VDD 0.19fF
C42113 POR2X1_96/A PAND2X1_538/a_16_344# 0.01fF
C42114 POR2X1_92/CTRL POR2X1_408/Y 0.00fF
C42115 POR2X1_38/B POR2X1_384/O 0.01fF
C42116 PAND2X1_658/A PAND2X1_789/CTRL 0.01fF
C42117 POR2X1_43/B POR2X1_39/Y 0.01fF
C42118 POR2X1_57/A PAND2X1_857/B 0.01fF
C42119 POR2X1_750/Y PAND2X1_32/B 0.05fF
C42120 D_INPUT_6 PAND2X1_1/O 0.03fF
C42121 PAND2X1_63/Y POR2X1_456/B 0.11fF
C42122 POR2X1_326/A PAND2X1_55/Y 0.90fF
C42123 POR2X1_43/B PAND2X1_566/O 0.05fF
C42124 PAND2X1_476/A PAND2X1_734/B 0.00fF
C42125 POR2X1_136/CTRL2 PAND2X1_348/A 0.02fF
C42126 POR2X1_38/Y PAND2X1_194/m4_208_n4# 0.01fF
C42127 POR2X1_96/A PAND2X1_802/a_56_28# 0.00fF
C42128 PAND2X1_322/O POR2X1_188/Y 0.03fF
C42129 POR2X1_731/m4_208_n4# POR2X1_854/B 0.07fF
C42130 POR2X1_575/CTRL POR2X1_569/A 0.04fF
C42131 PAND2X1_39/B POR2X1_646/A 0.01fF
C42132 PAND2X1_65/B POR2X1_779/O 0.01fF
C42133 POR2X1_523/A POR2X1_7/B 0.01fF
C42134 POR2X1_16/A PAND2X1_655/B 0.01fF
C42135 POR2X1_394/A POR2X1_321/O 0.03fF
C42136 POR2X1_343/Y PAND2X1_65/B 0.05fF
C42137 PAND2X1_824/B POR2X1_219/B 0.04fF
C42138 POR2X1_651/Y POR2X1_805/Y 0.01fF
C42139 PAND2X1_530/CTRL2 POR2X1_4/Y 0.02fF
C42140 PAND2X1_96/B POR2X1_507/A 0.01fF
C42141 POR2X1_832/CTRL POR2X1_711/Y 0.04fF
C42142 POR2X1_8/Y POR2X1_619/A 0.01fF
C42143 POR2X1_713/O PAND2X1_48/A 0.02fF
C42144 INPUT_1 PAND2X1_60/B 0.95fF
C42145 PAND2X1_20/A POR2X1_651/Y 0.05fF
C42146 POR2X1_447/B POR2X1_741/Y 0.10fF
C42147 POR2X1_57/A POR2X1_122/CTRL2 0.03fF
C42148 PAND2X1_793/Y POR2X1_184/O 0.01fF
C42149 POR2X1_244/Y POR2X1_318/A 0.07fF
C42150 VDD POR2X1_747/CTRL 0.00fF
C42151 POR2X1_334/B PAND2X1_134/CTRL 0.05fF
C42152 POR2X1_420/CTRL2 POR2X1_329/A 0.03fF
C42153 PAND2X1_857/A POR2X1_16/A 0.07fF
C42154 PAND2X1_730/a_76_28# PAND2X1_730/A 0.01fF
C42155 POR2X1_527/CTRL PAND2X1_550/B 0.01fF
C42156 POR2X1_93/A POR2X1_129/Y 0.10fF
C42157 POR2X1_648/Y POR2X1_807/CTRL 0.03fF
C42158 PAND2X1_700/CTRL PAND2X1_52/B 0.14fF
C42159 POR2X1_129/Y POR2X1_91/Y 0.03fF
C42160 POR2X1_327/Y POR2X1_361/O 0.01fF
C42161 PAND2X1_639/Y POR2X1_584/O 0.14fF
C42162 PAND2X1_357/Y PAND2X1_353/Y 0.09fF
C42163 PAND2X1_182/A POR2X1_77/Y 0.01fF
C42164 PAND2X1_586/CTRL PAND2X1_60/B 0.01fF
C42165 PAND2X1_631/A POR2X1_136/CTRL2 0.03fF
C42166 PAND2X1_687/a_16_344# PAND2X1_643/Y 0.02fF
C42167 PAND2X1_90/CTRL POR2X1_68/B 0.01fF
C42168 POR2X1_7/A PAND2X1_560/B 0.03fF
C42169 POR2X1_48/A PAND2X1_35/a_76_28# 0.01fF
C42170 POR2X1_532/A POR2X1_342/O 0.01fF
C42171 POR2X1_814/B POR2X1_651/Y 0.03fF
C42172 POR2X1_333/CTRL POR2X1_333/Y 0.00fF
C42173 POR2X1_456/B POR2X1_260/A 0.03fF
C42174 POR2X1_153/Y PAND2X1_123/CTRL 0.08fF
C42175 PAND2X1_70/CTRL2 POR2X1_451/A 0.01fF
C42176 POR2X1_96/Y PAND2X1_341/A 0.03fF
C42177 POR2X1_555/A PAND2X1_628/CTRL 0.02fF
C42178 PAND2X1_20/A POR2X1_67/Y 0.03fF
C42179 POR2X1_785/m4_208_n4# POR2X1_191/Y 0.04fF
C42180 POR2X1_841/B PAND2X1_39/B 0.03fF
C42181 POR2X1_416/B PAND2X1_35/CTRL 0.01fF
C42182 POR2X1_646/A POR2X1_805/Y 0.07fF
C42183 POR2X1_333/Y POR2X1_502/O 0.00fF
C42184 POR2X1_35/Y POR2X1_555/CTRL 0.01fF
C42185 POR2X1_304/a_56_344# POR2X1_90/Y 0.00fF
C42186 PAND2X1_458/CTRL2 POR2X1_5/Y 0.01fF
C42187 POR2X1_553/A POR2X1_553/a_16_28# 0.03fF
C42188 POR2X1_773/A POR2X1_773/CTRL2 0.01fF
C42189 POR2X1_119/Y POR2X1_315/Y 0.17fF
C42190 POR2X1_804/A POR2X1_711/Y 0.10fF
C42191 POR2X1_97/a_76_344# POR2X1_186/B 0.00fF
C42192 POR2X1_835/CTRL VDD 0.00fF
C42193 POR2X1_740/Y POR2X1_568/A 0.03fF
C42194 POR2X1_848/A POR2X1_260/B 0.07fF
C42195 POR2X1_332/Y POR2X1_332/CTRL 0.00fF
C42196 PAND2X1_593/Y POR2X1_385/Y 1.43fF
C42197 PAND2X1_56/Y POR2X1_717/B 0.03fF
C42198 POR2X1_376/B POR2X1_27/CTRL2 0.03fF
C42199 POR2X1_56/B PAND2X1_242/Y 0.30fF
C42200 PAND2X1_635/Y VDD 0.49fF
C42201 PAND2X1_20/A POR2X1_296/a_16_28# 0.02fF
C42202 POR2X1_421/Y POR2X1_20/B 0.96fF
C42203 POR2X1_356/A POR2X1_535/a_56_344# 0.03fF
C42204 PAND2X1_731/m4_208_n4# POR2X1_77/Y 0.12fF
C42205 POR2X1_241/CTRL POR2X1_776/A 0.01fF
C42206 POR2X1_474/O POR2X1_556/A 0.01fF
C42207 POR2X1_711/Y PAND2X1_306/CTRL2 0.03fF
C42208 POR2X1_39/B PAND2X1_509/m4_208_n4# 0.03fF
C42209 POR2X1_814/B POR2X1_646/A 0.01fF
C42210 POR2X1_647/B POR2X1_78/A 0.03fF
C42211 PAND2X1_649/A POR2X1_394/CTRL2 0.01fF
C42212 POR2X1_118/Y POR2X1_37/Y 0.03fF
C42213 POR2X1_537/Y POR2X1_851/O 0.01fF
C42214 POR2X1_463/O VDD 0.00fF
C42215 POR2X1_3/B PAND2X1_18/B 0.04fF
C42216 POR2X1_46/CTRL PAND2X1_9/Y 0.01fF
C42217 POR2X1_20/B PAND2X1_354/A 27.34fF
C42218 POR2X1_283/A POR2X1_77/Y 1.36fF
C42219 PAND2X1_85/O INPUT_0 0.15fF
C42220 PAND2X1_31/a_56_28# PAND2X1_3/A 0.00fF
C42221 POR2X1_285/Y POR2X1_655/A 0.01fF
C42222 PAND2X1_469/B PAND2X1_860/A 0.03fF
C42223 POR2X1_814/A PAND2X1_372/CTRL2 0.01fF
C42224 PAND2X1_600/CTRL POR2X1_121/B 0.07fF
C42225 POR2X1_777/B POR2X1_624/Y 0.03fF
C42226 POR2X1_129/CTRL POR2X1_67/A 0.05fF
C42227 POR2X1_569/A POR2X1_500/O 0.03fF
C42228 POR2X1_383/A POR2X1_717/B 0.03fF
C42229 POR2X1_48/A POR2X1_83/B 0.13fF
C42230 POR2X1_37/O POR2X1_612/Y 0.03fF
C42231 POR2X1_86/Y PAND2X1_100/CTRL 0.01fF
C42232 PAND2X1_48/A PAND2X1_304/CTRL 0.04fF
C42233 POR2X1_499/A POR2X1_130/A 0.07fF
C42234 PAND2X1_201/O POR2X1_88/Y 0.17fF
C42235 PAND2X1_489/O POR2X1_487/Y -0.00fF
C42236 PAND2X1_717/A POR2X1_55/Y 8.14fF
C42237 PAND2X1_65/B POR2X1_624/Y 0.03fF
C42238 POR2X1_129/O POR2X1_83/B 0.17fF
C42239 PAND2X1_829/CTRL PAND2X1_73/Y 0.01fF
C42240 PAND2X1_435/CTRL2 POR2X1_411/B 0.01fF
C42241 POR2X1_48/A POR2X1_626/Y 0.00fF
C42242 POR2X1_264/Y POR2X1_814/A 0.03fF
C42243 POR2X1_604/Y POR2X1_32/A 0.32fF
C42244 POR2X1_640/Y POR2X1_476/A 0.03fF
C42245 POR2X1_669/B POR2X1_667/A 0.04fF
C42246 POR2X1_163/CTRL2 POR2X1_23/Y 0.01fF
C42247 PAND2X1_340/B POR2X1_236/Y 0.05fF
C42248 PAND2X1_837/O POR2X1_42/Y 0.02fF
C42249 POR2X1_66/A POR2X1_404/CTRL 0.01fF
C42250 POR2X1_49/Y PAND2X1_448/CTRL2 0.05fF
C42251 POR2X1_20/B INPUT_5 0.03fF
C42252 POR2X1_708/O PAND2X1_39/B 0.02fF
C42253 PAND2X1_414/CTRL2 PAND2X1_6/A 0.01fF
C42254 POR2X1_13/A POR2X1_257/A 0.19fF
C42255 PAND2X1_776/Y PAND2X1_803/A 0.02fF
C42256 PAND2X1_124/Y PAND2X1_199/A 1.83fF
C42257 POR2X1_260/B POR2X1_480/A 0.03fF
C42258 POR2X1_98/B POR2X1_98/A 0.02fF
C42259 PAND2X1_205/A PAND2X1_204/CTRL2 0.00fF
C42260 POR2X1_644/Y PAND2X1_90/Y 0.02fF
C42261 POR2X1_54/Y POR2X1_668/Y 0.03fF
C42262 PAND2X1_612/B VDD 0.01fF
C42263 POR2X1_68/A PAND2X1_617/a_16_344# 0.02fF
C42264 POR2X1_105/Y PAND2X1_251/a_16_344# 0.02fF
C42265 PAND2X1_404/Y VDD 0.58fF
C42266 PAND2X1_116/O POR2X1_48/A 0.04fF
C42267 POR2X1_20/B PAND2X1_724/B 0.02fF
C42268 PAND2X1_58/A POR2X1_720/m4_208_n4# 0.08fF
C42269 POR2X1_841/B POR2X1_325/A 0.03fF
C42270 POR2X1_102/Y PAND2X1_795/CTRL2 0.11fF
C42271 PAND2X1_792/a_16_344# POR2X1_533/A 0.03fF
C42272 PAND2X1_629/CTRL POR2X1_496/Y 0.06fF
C42273 POR2X1_66/B POR2X1_641/O 0.01fF
C42274 PAND2X1_32/a_16_344# PAND2X1_32/B 0.02fF
C42275 PAND2X1_206/B POR2X1_38/Y 0.07fF
C42276 POR2X1_65/A POR2X1_32/A 0.23fF
C42277 POR2X1_492/Y POR2X1_491/Y 0.00fF
C42278 PAND2X1_94/A POR2X1_643/CTRL2 0.01fF
C42279 PAND2X1_217/O PAND2X1_197/Y 0.00fF
C42280 PAND2X1_644/a_16_344# PAND2X1_643/Y 0.01fF
C42281 PAND2X1_266/a_56_28# POR2X1_73/Y 0.00fF
C42282 PAND2X1_826/CTRL PAND2X1_55/Y 0.01fF
C42283 POR2X1_32/A PAND2X1_558/CTRL 0.01fF
C42284 POR2X1_753/Y POR2X1_5/Y 0.07fF
C42285 POR2X1_471/CTRL POR2X1_66/A 0.03fF
C42286 POR2X1_311/Y PAND2X1_220/Y 0.03fF
C42287 POR2X1_650/CTRL PAND2X1_65/B 0.01fF
C42288 POR2X1_669/B PAND2X1_712/B 0.02fF
C42289 POR2X1_260/B PAND2X1_753/O 0.01fF
C42290 POR2X1_858/O VDD 0.00fF
C42291 POR2X1_114/B PAND2X1_39/B 0.07fF
C42292 POR2X1_39/B PAND2X1_841/Y 0.01fF
C42293 PAND2X1_90/A POR2X1_260/B 6.93fF
C42294 POR2X1_175/O POR2X1_78/A 0.02fF
C42295 PAND2X1_436/A POR2X1_677/CTRL 0.04fF
C42296 POR2X1_440/Y POR2X1_440/B 0.16fF
C42297 POR2X1_402/A POR2X1_68/Y 0.01fF
C42298 POR2X1_102/Y POR2X1_236/Y 2.00fF
C42299 PAND2X1_271/CTRL2 POR2X1_804/A 0.14fF
C42300 PAND2X1_20/A POR2X1_402/m4_208_n4# 0.15fF
C42301 PAND2X1_124/Y PAND2X1_197/Y 0.02fF
C42302 PAND2X1_42/CTRL PAND2X1_41/B 0.01fF
C42303 PAND2X1_787/A POR2X1_150/Y 0.07fF
C42304 POR2X1_409/B POR2X1_277/CTRL 0.01fF
C42305 PAND2X1_16/O PAND2X1_41/B 0.01fF
C42306 POR2X1_814/B POR2X1_461/CTRL2 0.03fF
C42307 PAND2X1_644/Y POR2X1_42/Y 0.00fF
C42308 POR2X1_49/Y PAND2X1_576/O 0.19fF
C42309 POR2X1_193/A POR2X1_66/A 0.00fF
C42310 POR2X1_66/A POR2X1_579/Y 0.03fF
C42311 INPUT_1 PAND2X1_608/CTRL2 0.03fF
C42312 PAND2X1_658/O POR2X1_376/B 0.08fF
C42313 POR2X1_692/a_16_28# POR2X1_46/Y 0.03fF
C42314 POR2X1_311/Y PAND2X1_739/Y 0.01fF
C42315 POR2X1_16/A POR2X1_329/A 0.05fF
C42316 POR2X1_394/Y VDD 0.15fF
C42317 PAND2X1_697/CTRL POR2X1_260/B 0.00fF
C42318 PAND2X1_494/O POR2X1_260/B 0.05fF
C42319 INPUT_1 PAND2X1_206/B 0.07fF
C42320 PAND2X1_6/Y PAND2X1_248/CTRL2 0.00fF
C42321 POR2X1_283/Y VDD 0.00fF
C42322 POR2X1_669/B POR2X1_252/O 0.06fF
C42323 PAND2X1_254/CTRL2 POR2X1_669/B 0.03fF
C42324 POR2X1_155/CTRL2 POR2X1_750/B 0.01fF
C42325 POR2X1_355/B POR2X1_836/A 0.05fF
C42326 POR2X1_857/B POR2X1_590/A 0.03fF
C42327 PAND2X1_88/O POR2X1_87/Y 0.00fF
C42328 POR2X1_76/A POR2X1_573/A 0.02fF
C42329 POR2X1_141/Y VDD 0.22fF
C42330 POR2X1_445/A POR2X1_540/O 0.04fF
C42331 POR2X1_335/A D_INPUT_0 0.03fF
C42332 POR2X1_66/A PAND2X1_385/a_56_28# 0.00fF
C42333 PAND2X1_472/A POR2X1_23/Y 0.07fF
C42334 PAND2X1_433/CTRL2 POR2X1_78/A 0.01fF
C42335 POR2X1_411/B PAND2X1_717/Y 0.08fF
C42336 PAND2X1_573/B POR2X1_293/Y 0.03fF
C42337 POR2X1_660/m4_208_n4# POR2X1_307/Y 0.01fF
C42338 PAND2X1_257/CTRL2 POR2X1_750/B 0.14fF
C42339 POR2X1_590/A POR2X1_214/B 0.61fF
C42340 POR2X1_56/B POR2X1_60/A 0.07fF
C42341 POR2X1_451/O POR2X1_635/Y 0.01fF
C42342 POR2X1_341/A POR2X1_274/B 0.01fF
C42343 POR2X1_614/A POR2X1_66/A 0.43fF
C42344 POR2X1_404/B POR2X1_404/O 0.01fF
C42345 POR2X1_49/Y POR2X1_13/A 0.08fF
C42346 POR2X1_56/a_16_28# POR2X1_55/Y 0.03fF
C42347 POR2X1_330/Y PAND2X1_131/a_76_28# 0.02fF
C42348 POR2X1_675/A VDD 0.00fF
C42349 POR2X1_458/Y POR2X1_188/Y 0.03fF
C42350 POR2X1_634/A PAND2X1_132/O 0.02fF
C42351 POR2X1_248/A POR2X1_248/a_16_28# 0.05fF
C42352 POR2X1_257/A POR2X1_321/Y 0.02fF
C42353 POR2X1_846/Y POR2X1_753/a_56_344# 0.00fF
C42354 POR2X1_748/A PAND2X1_784/CTRL 0.14fF
C42355 POR2X1_856/CTRL POR2X1_855/Y 0.01fF
C42356 PAND2X1_341/A POR2X1_37/Y 0.03fF
C42357 POR2X1_814/A POR2X1_502/Y 0.05fF
C42358 POR2X1_66/A POR2X1_38/B 0.26fF
C42359 POR2X1_66/B POR2X1_42/Y 0.19fF
C42360 PAND2X1_798/B POR2X1_516/Y 0.03fF
C42361 POR2X1_669/B POR2X1_321/O 0.05fF
C42362 POR2X1_682/CTRL2 POR2X1_829/A 0.00fF
C42363 POR2X1_283/a_16_28# PAND2X1_365/B 0.05fF
C42364 POR2X1_290/Y PAND2X1_402/O 0.05fF
C42365 PAND2X1_793/Y PAND2X1_185/O 0.01fF
C42366 POR2X1_423/Y POR2X1_372/Y 0.09fF
C42367 POR2X1_65/A PAND2X1_35/Y 0.04fF
C42368 POR2X1_275/O PAND2X1_390/Y 0.01fF
C42369 PAND2X1_23/Y POR2X1_794/B 0.01fF
C42370 PAND2X1_307/m4_208_n4# POR2X1_304/m4_208_n4# 0.05fF
C42371 PAND2X1_137/a_16_344# PAND2X1_354/A 0.02fF
C42372 POR2X1_93/A POR2X1_37/Y 0.08fF
C42373 PAND2X1_785/Y POR2X1_5/Y 0.02fF
C42374 POR2X1_333/A POR2X1_782/A 0.34fF
C42375 POR2X1_43/B PAND2X1_478/B 0.16fF
C42376 POR2X1_102/Y POR2X1_232/Y 0.34fF
C42377 POR2X1_455/CTRL POR2X1_76/Y 0.01fF
C42378 POR2X1_411/B PAND2X1_502/CTRL2 0.01fF
C42379 POR2X1_680/Y PAND2X1_205/Y 0.01fF
C42380 PAND2X1_615/a_76_28# D_INPUT_0 0.02fF
C42381 POR2X1_647/O POR2X1_101/Y 0.07fF
C42382 POR2X1_614/A POR2X1_634/CTRL2 0.03fF
C42383 POR2X1_79/Y PAND2X1_473/B 0.03fF
C42384 POR2X1_278/Y PAND2X1_84/Y 0.03fF
C42385 POR2X1_96/A PAND2X1_739/CTRL2 0.01fF
C42386 PAND2X1_511/O VDD 0.00fF
C42387 POR2X1_307/B POR2X1_513/B 0.12fF
C42388 PAND2X1_721/a_16_344# POR2X1_7/B 0.03fF
C42389 PAND2X1_48/B POR2X1_61/Y 0.09fF
C42390 POR2X1_102/Y PAND2X1_858/Y 0.03fF
C42391 POR2X1_455/A POR2X1_750/B 0.05fF
C42392 POR2X1_614/A PAND2X1_427/O 0.04fF
C42393 POR2X1_41/B POR2X1_48/O 0.01fF
C42394 POR2X1_614/A PAND2X1_230/a_56_28# 0.00fF
C42395 PAND2X1_403/Y POR2X1_293/Y 0.01fF
C42396 POR2X1_646/O POR2X1_480/A 0.03fF
C42397 D_INPUT_3 POR2X1_414/CTRL 0.01fF
C42398 POR2X1_220/Y VDD 1.57fF
C42399 POR2X1_183/Y POR2X1_40/Y 0.04fF
C42400 POR2X1_864/A POR2X1_294/A 0.00fF
C42401 PAND2X1_65/B POR2X1_785/A 0.06fF
C42402 POR2X1_631/O POR2X1_631/B 0.02fF
C42403 POR2X1_818/Y POR2X1_750/Y 0.00fF
C42404 POR2X1_156/B POR2X1_467/Y 0.03fF
C42405 POR2X1_83/CTRL POR2X1_23/Y 0.01fF
C42406 POR2X1_66/B POR2X1_123/Y 0.01fF
C42407 POR2X1_253/Y POR2X1_423/Y 0.01fF
C42408 POR2X1_37/Y POR2X1_416/O 0.01fF
C42409 POR2X1_669/B POR2X1_245/Y 0.07fF
C42410 POR2X1_368/CTRL POR2X1_372/Y 0.06fF
C42411 POR2X1_502/A POR2X1_459/O 0.01fF
C42412 POR2X1_114/B PAND2X1_299/a_16_344# 0.01fF
C42413 PAND2X1_55/Y POR2X1_480/A 0.14fF
C42414 POR2X1_404/Y VDD 0.57fF
C42415 POR2X1_66/A PAND2X1_393/a_76_28# 0.04fF
C42416 PAND2X1_96/B POR2X1_479/a_16_28# 0.03fF
C42417 PAND2X1_659/CTRL POR2X1_494/Y 0.00fF
C42418 D_INPUT_0 POR2X1_249/Y 0.03fF
C42419 POR2X1_119/Y POR2X1_442/CTRL2 0.00fF
C42420 PAND2X1_651/Y PAND2X1_620/Y 0.02fF
C42421 PAND2X1_778/a_16_344# POR2X1_55/Y 0.02fF
C42422 POR2X1_814/A POR2X1_779/O 0.31fF
C42423 POR2X1_13/A PAND2X1_553/B 0.01fF
C42424 POR2X1_290/Y POR2X1_233/CTRL2 0.02fF
C42425 POR2X1_750/CTRL2 POR2X1_750/A 0.01fF
C42426 POR2X1_78/A POR2X1_218/CTRL2 0.01fF
C42427 POR2X1_710/A POR2X1_710/O 0.02fF
C42428 PAND2X1_724/O PAND2X1_731/B 0.02fF
C42429 POR2X1_57/A PAND2X1_169/Y 0.03fF
C42430 POR2X1_65/A PAND2X1_651/Y 0.03fF
C42431 POR2X1_49/Y PAND2X1_661/B 1.40fF
C42432 PAND2X1_96/B POR2X1_734/A 0.07fF
C42433 POR2X1_796/A POR2X1_296/B 2.02fF
C42434 POR2X1_343/Y POR2X1_814/A 0.27fF
C42435 POR2X1_590/A POR2X1_590/a_56_344# 0.00fF
C42436 PAND2X1_20/A POR2X1_222/A 0.03fF
C42437 POR2X1_287/CTRL2 POR2X1_249/Y 0.01fF
C42438 PAND2X1_339/Y POR2X1_497/Y 0.03fF
C42439 POR2X1_289/CTRL2 VDD 0.00fF
C42440 PAND2X1_641/Y POR2X1_409/B 0.00fF
C42441 POR2X1_814/B PAND2X1_177/CTRL2 0.01fF
C42442 POR2X1_227/a_16_28# POR2X1_854/B 0.05fF
C42443 POR2X1_315/Y POR2X1_442/Y 0.11fF
C42444 POR2X1_236/Y POR2X1_531/Y 0.01fF
C42445 POR2X1_41/B POR2X1_55/Y 0.25fF
C42446 POR2X1_865/B POR2X1_287/B 0.03fF
C42447 PAND2X1_69/A POR2X1_786/CTRL 0.01fF
C42448 POR2X1_300/CTRL POR2X1_46/Y 0.24fF
C42449 POR2X1_502/A D_GATE_662 0.09fF
C42450 D_INPUT_0 POR2X1_394/A 0.10fF
C42451 POR2X1_355/B POR2X1_853/A 0.03fF
C42452 PAND2X1_684/CTRL2 POR2X1_78/A 0.03fF
C42453 PAND2X1_374/CTRL2 POR2X1_40/Y 0.01fF
C42454 PAND2X1_464/Y VDD 0.00fF
C42455 POR2X1_220/Y POR2X1_741/Y 0.03fF
C42456 PAND2X1_55/Y POR2X1_553/Y 0.01fF
C42457 POR2X1_192/Y D_GATE_741 0.10fF
C42458 PAND2X1_96/B POR2X1_563/O 0.01fF
C42459 POR2X1_14/Y POR2X1_419/O 0.18fF
C42460 POR2X1_102/Y POR2X1_757/Y 0.04fF
C42461 POR2X1_231/O POR2X1_785/A 0.15fF
C42462 POR2X1_260/B POR2X1_572/Y 0.12fF
C42463 POR2X1_66/B PAND2X1_376/CTRL2 0.11fF
C42464 POR2X1_802/O POR2X1_750/B 0.03fF
C42465 PAND2X1_467/Y POR2X1_418/Y 0.05fF
C42466 POR2X1_197/a_16_28# POR2X1_741/Y 0.03fF
C42467 PAND2X1_453/A POR2X1_419/O 0.01fF
C42468 PAND2X1_857/A PAND2X1_200/a_76_28# 0.01fF
C42469 POR2X1_66/B PAND2X1_127/CTRL2 0.01fF
C42470 POR2X1_821/Y POR2X1_236/Y 0.04fF
C42471 POR2X1_775/A POR2X1_776/B 0.00fF
C42472 PAND2X1_90/A PAND2X1_55/Y 0.06fF
C42473 PAND2X1_581/a_76_28# PAND2X1_3/B 0.02fF
C42474 POR2X1_617/Y POR2X1_48/A 0.03fF
C42475 POR2X1_96/A PAND2X1_734/CTRL2 0.03fF
C42476 POR2X1_832/A POR2X1_807/A 0.04fF
C42477 POR2X1_78/B POR2X1_194/O 0.02fF
C42478 POR2X1_488/Y POR2X1_42/Y 0.04fF
C42479 PAND2X1_738/Y PAND2X1_182/O 0.25fF
C42480 POR2X1_222/Y POR2X1_579/Y 0.03fF
C42481 D_GATE_222 POR2X1_578/Y 0.07fF
C42482 POR2X1_502/A POR2X1_462/B 0.03fF
C42483 PAND2X1_139/a_16_344# PAND2X1_349/A 0.01fF
C42484 POR2X1_14/Y PAND2X1_308/Y 0.04fF
C42485 POR2X1_754/A PAND2X1_6/A 0.03fF
C42486 POR2X1_65/A POR2X1_503/Y 0.01fF
C42487 POR2X1_278/Y POR2X1_594/A 0.12fF
C42488 POR2X1_502/A D_INPUT_1 0.10fF
C42489 PAND2X1_453/A PAND2X1_308/Y 0.01fF
C42490 PAND2X1_564/O POR2X1_73/Y 0.07fF
C42491 POR2X1_43/B POR2X1_494/Y 0.03fF
C42492 POR2X1_5/Y PAND2X1_656/A 0.05fF
C42493 PAND2X1_6/A PAND2X1_375/CTRL 0.01fF
C42494 POR2X1_220/Y PAND2X1_32/B 0.06fF
C42495 VDD POR2X1_395/Y 0.03fF
C42496 POR2X1_435/Y POR2X1_788/B 0.03fF
C42497 PAND2X1_31/m4_208_n4# PAND2X1_18/B 0.15fF
C42498 INPUT_1 POR2X1_750/B 0.03fF
C42499 PAND2X1_48/B POR2X1_35/Y 0.04fF
C42500 PAND2X1_94/A PAND2X1_41/B 0.18fF
C42501 POR2X1_36/B VDD 0.43fF
C42502 POR2X1_673/A PAND2X1_4/a_16_344# 0.02fF
C42503 PAND2X1_206/A POR2X1_39/B 0.17fF
C42504 POR2X1_814/A POR2X1_579/m4_208_n4# 0.06fF
C42505 PAND2X1_23/Y POR2X1_638/B 0.06fF
C42506 POR2X1_41/B PAND2X1_186/CTRL 0.02fF
C42507 POR2X1_13/A PAND2X1_778/Y 0.01fF
C42508 POR2X1_227/B PAND2X1_52/B 0.03fF
C42509 POR2X1_150/Y POR2X1_173/CTRL 0.01fF
C42510 POR2X1_498/a_16_28# POR2X1_498/A 0.08fF
C42511 POR2X1_404/Y PAND2X1_32/B 0.03fF
C42512 INPUT_0 POR2X1_597/O 0.36fF
C42513 PAND2X1_652/A PAND2X1_794/B 0.04fF
C42514 POR2X1_62/Y POR2X1_83/B 0.15fF
C42515 PAND2X1_341/A POR2X1_293/Y 0.03fF
C42516 POR2X1_256/Y POR2X1_55/Y 0.02fF
C42517 POR2X1_804/A POR2X1_733/A 0.10fF
C42518 POR2X1_355/A POR2X1_507/A 0.34fF
C42519 POR2X1_7/B POR2X1_591/Y 0.03fF
C42520 POR2X1_832/B PAND2X1_69/A 0.10fF
C42521 POR2X1_55/Y PAND2X1_548/O 0.03fF
C42522 POR2X1_193/A POR2X1_532/A 0.03fF
C42523 POR2X1_327/Y PAND2X1_279/a_56_28# 0.00fF
C42524 POR2X1_614/A POR2X1_222/Y 0.06fF
C42525 POR2X1_130/A POR2X1_537/A 0.02fF
C42526 POR2X1_532/A POR2X1_579/Y 0.06fF
C42527 PAND2X1_572/a_16_344# POR2X1_46/Y 0.02fF
C42528 PAND2X1_561/A PAND2X1_853/B 0.12fF
C42529 PAND2X1_799/a_76_28# INPUT_0 0.01fF
C42530 POR2X1_93/A POR2X1_293/Y 5.34fF
C42531 POR2X1_482/Y PAND2X1_508/Y 0.00fF
C42532 POR2X1_46/Y POR2X1_387/Y 0.10fF
C42533 PAND2X1_490/O POR2X1_334/B 0.44fF
C42534 PAND2X1_687/O POR2X1_60/A 0.03fF
C42535 PAND2X1_434/CTRL2 INPUT_0 0.03fF
C42536 POR2X1_777/B POR2X1_186/B 0.05fF
C42537 POR2X1_344/A POR2X1_383/A 0.04fF
C42538 POR2X1_293/Y POR2X1_91/Y 1.74fF
C42539 VDD POR2X1_577/Y 0.00fF
C42540 PAND2X1_793/Y POR2X1_530/Y 0.02fF
C42541 POR2X1_539/A POR2X1_566/A 0.04fF
C42542 POR2X1_333/m4_208_n4# PAND2X1_32/B 0.17fF
C42543 POR2X1_13/A PAND2X1_720/O 0.02fF
C42544 POR2X1_130/Y POR2X1_140/CTRL2 0.04fF
C42545 POR2X1_773/CTRL VDD 0.00fF
C42546 POR2X1_700/a_16_28# POR2X1_700/Y 0.02fF
C42547 PAND2X1_44/O PAND2X1_18/B 0.15fF
C42548 PAND2X1_104/CTRL2 POR2X1_4/Y 0.05fF
C42549 POR2X1_557/A VDD 0.42fF
C42550 POR2X1_258/CTRL2 PAND2X1_566/Y 0.01fF
C42551 POR2X1_237/CTRL PAND2X1_308/Y 0.01fF
C42552 PAND2X1_718/CTRL2 POR2X1_591/Y 0.01fF
C42553 POR2X1_527/CTRL2 POR2X1_96/A 0.00fF
C42554 PAND2X1_79/Y PAND2X1_316/CTRL 0.03fF
C42555 POR2X1_619/A POR2X1_619/O 0.11fF
C42556 PAND2X1_480/B PAND2X1_112/O 0.00fF
C42557 POR2X1_559/CTRL POR2X1_68/B 0.07fF
C42558 POR2X1_52/A PAND2X1_717/Y 0.03fF
C42559 PAND2X1_65/B POR2X1_186/B 0.10fF
C42560 POR2X1_294/B POR2X1_550/Y 0.17fF
C42561 POR2X1_614/A POR2X1_532/A 0.21fF
C42562 POR2X1_416/O POR2X1_293/Y 0.01fF
C42563 PAND2X1_57/B POR2X1_260/A 2.64fF
C42564 POR2X1_48/CTRL2 PAND2X1_123/Y 0.01fF
C42565 INPUT_0 POR2X1_171/a_16_28# 0.11fF
C42566 POR2X1_750/B PAND2X1_680/CTRL 0.01fF
C42567 POR2X1_523/Y PAND2X1_521/O 0.02fF
C42568 PAND2X1_742/B POR2X1_283/A 0.06fF
C42569 POR2X1_286/CTRL2 PAND2X1_52/B 0.01fF
C42570 PAND2X1_572/CTRL POR2X1_52/Y 0.01fF
C42571 POR2X1_638/Y POR2X1_639/Y 0.00fF
C42572 PAND2X1_23/Y PAND2X1_823/CTRL2 0.03fF
C42573 POR2X1_83/Y PAND2X1_61/Y 0.02fF
C42574 POR2X1_259/O POR2X1_785/A 0.01fF
C42575 PAND2X1_850/Y POR2X1_40/Y 0.05fF
C42576 POR2X1_407/A POR2X1_832/A 0.03fF
C42577 PAND2X1_215/B POR2X1_7/O 0.05fF
C42578 POR2X1_38/B POR2X1_532/A 0.10fF
C42579 POR2X1_316/CTRL POR2X1_13/A 0.01fF
C42580 POR2X1_437/CTRL2 PAND2X1_794/B 0.01fF
C42581 POR2X1_307/CTRL POR2X1_711/Y 0.08fF
C42582 POR2X1_709/B VDD 0.01fF
C42583 POR2X1_501/B POR2X1_318/A 0.07fF
C42584 POR2X1_99/B POR2X1_193/Y 0.02fF
C42585 POR2X1_346/B PAND2X1_55/Y 0.03fF
C42586 PAND2X1_57/B POR2X1_363/A 0.48fF
C42587 PAND2X1_6/Y POR2X1_850/a_16_28# 0.01fF
C42588 PAND2X1_30/O POR2X1_635/A 0.00fF
C42589 POR2X1_14/Y POR2X1_77/Y 0.09fF
C42590 PAND2X1_659/Y POR2X1_822/CTRL 0.00fF
C42591 PAND2X1_57/B PAND2X1_142/O 0.02fF
C42592 POR2X1_315/Y POR2X1_237/Y 0.03fF
C42593 PAND2X1_631/A POR2X1_5/Y 0.03fF
C42594 POR2X1_52/A PAND2X1_502/CTRL2 0.01fF
C42595 PAND2X1_94/A PAND2X1_411/CTRL 0.01fF
C42596 PAND2X1_126/CTRL PAND2X1_69/A 0.01fF
C42597 POR2X1_685/A POR2X1_828/A 0.00fF
C42598 INPUT_0 PAND2X1_851/CTRL 0.03fF
C42599 PAND2X1_724/B PAND2X1_303/Y 0.25fF
C42600 POR2X1_794/B POR2X1_711/Y 0.07fF
C42601 POR2X1_740/Y POR2X1_444/Y 0.03fF
C42602 PAND2X1_831/CTRL POR2X1_39/B 0.01fF
C42603 POR2X1_93/A POR2X1_408/Y 0.10fF
C42604 POR2X1_796/A POR2X1_796/a_16_28# -0.00fF
C42605 POR2X1_502/A POR2X1_620/B 0.07fF
C42606 POR2X1_784/O POR2X1_725/Y 0.03fF
C42607 D_INPUT_6 POR2X1_1/O 0.01fF
C42608 POR2X1_41/B PAND2X1_199/B 0.03fF
C42609 POR2X1_119/Y PAND2X1_480/B 0.00fF
C42610 PAND2X1_641/O PAND2X1_651/Y 0.02fF
C42611 POR2X1_828/A POR2X1_260/A 0.01fF
C42612 POR2X1_294/B POR2X1_195/CTRL 0.01fF
C42613 POR2X1_814/A POR2X1_624/Y 0.07fF
C42614 PAND2X1_605/CTRL POR2X1_73/Y 0.04fF
C42615 POR2X1_145/Y POR2X1_146/O 0.00fF
C42616 POR2X1_383/A POR2X1_338/CTRL 0.00fF
C42617 POR2X1_236/Y POR2X1_761/A 0.08fF
C42618 PAND2X1_530/CTRL2 POR2X1_620/B 0.01fF
C42619 PAND2X1_75/CTRL POR2X1_624/Y 0.05fF
C42620 POR2X1_502/A POR2X1_374/CTRL 0.01fF
C42621 POR2X1_383/A PAND2X1_824/O 0.05fF
C42622 PAND2X1_90/A PAND2X1_90/CTRL 0.03fF
C42623 POR2X1_57/A POR2X1_16/A 0.35fF
C42624 PAND2X1_651/a_76_28# POR2X1_43/B 0.01fF
C42625 PAND2X1_493/O POR2X1_599/A 0.06fF
C42626 PAND2X1_44/a_56_28# PAND2X1_72/A 0.00fF
C42627 POR2X1_234/A POR2X1_667/A 0.02fF
C42628 POR2X1_503/CTRL2 POR2X1_283/A 0.03fF
C42629 POR2X1_119/Y PAND2X1_398/CTRL 0.01fF
C42630 POR2X1_101/Y POR2X1_569/A 0.10fF
C42631 POR2X1_343/A POR2X1_343/B 0.01fF
C42632 POR2X1_38/Y PAND2X1_560/B 0.03fF
C42633 PAND2X1_467/Y PAND2X1_550/B 0.03fF
C42634 POR2X1_863/A POR2X1_436/O 0.00fF
C42635 POR2X1_714/O POR2X1_703/Y 0.02fF
C42636 POR2X1_66/B POR2X1_814/CTRL2 0.00fF
C42637 POR2X1_416/B POR2X1_481/A 0.06fF
C42638 POR2X1_176/O POR2X1_90/Y 0.02fF
C42639 POR2X1_513/B POR2X1_513/A 0.00fF
C42640 PAND2X1_55/Y PAND2X1_304/O 0.01fF
C42641 POR2X1_169/CTRL POR2X1_566/B 0.07fF
C42642 POR2X1_43/B PAND2X1_352/Y 0.01fF
C42643 POR2X1_687/CTRL POR2X1_814/A 0.06fF
C42644 POR2X1_816/A POR2X1_171/Y 0.03fF
C42645 PAND2X1_472/B POR2X1_77/Y 0.11fF
C42646 D_INPUT_7 PAND2X1_11/Y 0.07fF
C42647 PAND2X1_358/A PAND2X1_99/Y 0.01fF
C42648 POR2X1_257/A PAND2X1_562/Y 0.09fF
C42649 POR2X1_707/Y POR2X1_260/A 0.02fF
C42650 PAND2X1_575/A POR2X1_184/CTRL 0.01fF
C42651 POR2X1_862/A POR2X1_649/O 0.00fF
C42652 PAND2X1_661/Y PAND2X1_120/CTRL2 0.06fF
C42653 POR2X1_614/A PAND2X1_143/a_16_344# 0.01fF
C42654 POR2X1_697/Y POR2X1_39/B 0.02fF
C42655 PAND2X1_404/Y PAND2X1_9/Y 0.03fF
C42656 POR2X1_440/B POR2X1_590/A 0.01fF
C42657 PAND2X1_6/Y POR2X1_542/CTRL 0.01fF
C42658 POR2X1_505/Y PAND2X1_630/B 0.05fF
C42659 POR2X1_371/CTRL POR2X1_387/Y 0.07fF
C42660 PAND2X1_238/CTRL2 PAND2X1_52/B 0.03fF
C42661 POR2X1_55/Y POR2X1_77/Y 0.30fF
C42662 POR2X1_673/Y POR2X1_546/CTRL 0.02fF
C42663 POR2X1_458/Y POR2X1_457/CTRL 0.04fF
C42664 POR2X1_103/a_76_344# PAND2X1_349/A 0.00fF
C42665 POR2X1_178/Y PAND2X1_348/A 0.02fF
C42666 PAND2X1_508/Y PAND2X1_349/A 0.03fF
C42667 POR2X1_259/B POR2X1_260/A 0.07fF
C42668 POR2X1_136/Y POR2X1_183/a_16_28# 0.03fF
C42669 PAND2X1_357/Y POR2X1_39/B 0.03fF
C42670 PAND2X1_109/CTRL2 PAND2X1_32/B 0.01fF
C42671 POR2X1_65/CTRL2 POR2X1_60/A 0.06fF
C42672 POR2X1_10/O POR2X1_394/A 0.17fF
C42673 POR2X1_651/Y VDD 0.13fF
C42674 POR2X1_677/Y POR2X1_236/Y 0.02fF
C42675 POR2X1_496/Y POR2X1_20/B 0.08fF
C42676 POR2X1_846/A POR2X1_793/CTRL2 0.00fF
C42677 POR2X1_508/B POR2X1_566/B 0.05fF
C42678 PAND2X1_687/A PAND2X1_687/B 0.00fF
C42679 PAND2X1_560/B POR2X1_153/Y 0.07fF
C42680 POR2X1_9/Y POR2X1_236/Y 0.10fF
C42681 POR2X1_394/A PAND2X1_162/A 0.01fF
C42682 POR2X1_250/Y PAND2X1_742/a_76_28# 0.03fF
C42683 POR2X1_90/Y PAND2X1_326/CTRL2 0.03fF
C42684 POR2X1_67/Y PAND2X1_526/CTRL 0.01fF
C42685 POR2X1_290/Y POR2X1_825/Y 0.03fF
C42686 POR2X1_257/A POR2X1_163/Y 0.96fF
C42687 POR2X1_257/A POR2X1_29/A 1.11fF
C42688 POR2X1_294/B POR2X1_535/CTRL 0.01fF
C42689 POR2X1_54/Y POR2X1_104/CTRL2 0.01fF
C42690 POR2X1_274/A POR2X1_274/O 0.02fF
C42691 PAND2X1_94/A PAND2X1_122/O 0.27fF
C42692 POR2X1_20/B PAND2X1_733/A 0.00fF
C42693 POR2X1_571/a_16_28# POR2X1_560/Y -0.00fF
C42694 POR2X1_571/a_76_344# POR2X1_561/Y 0.02fF
C42695 POR2X1_647/B POR2X1_285/Y 0.00fF
C42696 POR2X1_48/A POR2X1_482/CTRL2 0.01fF
C42697 POR2X1_23/Y POR2X1_482/CTRL 0.02fF
C42698 POR2X1_528/Y POR2X1_39/B 0.07fF
C42699 POR2X1_282/Y PAND2X1_805/A 0.05fF
C42700 POR2X1_41/B PAND2X1_458/O 0.03fF
C42701 POR2X1_376/B PAND2X1_449/CTRL 0.10fF
C42702 POR2X1_274/A POR2X1_296/B 0.03fF
C42703 POR2X1_661/A POR2X1_740/Y 0.00fF
C42704 PAND2X1_338/B PAND2X1_333/Y 0.02fF
C42705 POR2X1_736/A POR2X1_736/a_16_28# 0.09fF
C42706 POR2X1_203/CTRL PAND2X1_72/A 0.01fF
C42707 POR2X1_67/Y VDD 0.80fF
C42708 POR2X1_834/a_16_28# POR2X1_260/B 0.03fF
C42709 PAND2X1_294/CTRL2 POR2X1_40/Y 0.00fF
C42710 POR2X1_851/A POR2X1_590/A 0.00fF
C42711 POR2X1_646/A VDD -0.00fF
C42712 POR2X1_323/O POR2X1_485/Y 0.01fF
C42713 POR2X1_411/B POR2X1_226/Y 0.01fF
C42714 POR2X1_90/Y POR2X1_91/CTRL2 0.00fF
C42715 POR2X1_41/B POR2X1_441/CTRL 0.02fF
C42716 POR2X1_351/CTRL2 PAND2X1_72/A 0.10fF
C42717 POR2X1_116/A POR2X1_362/B 0.00fF
C42718 POR2X1_174/B POR2X1_567/B 0.10fF
C42719 POR2X1_669/B D_INPUT_0 0.12fF
C42720 POR2X1_811/O PAND2X1_73/Y 0.01fF
C42721 POR2X1_614/A POR2X1_452/A 0.00fF
C42722 POR2X1_66/A POR2X1_590/A 0.37fF
C42723 POR2X1_68/CTRL POR2X1_296/B 0.01fF
C42724 POR2X1_416/B PAND2X1_737/B 0.12fF
C42725 POR2X1_411/B PAND2X1_793/O 0.02fF
C42726 POR2X1_101/Y PAND2X1_72/A 0.05fF
C42727 POR2X1_477/CTRL2 VDD 0.00fF
C42728 POR2X1_814/A POR2X1_785/A 0.07fF
C42729 PAND2X1_454/B PAND2X1_803/A 0.00fF
C42730 D_GATE_865 POR2X1_452/Y 0.05fF
C42731 POR2X1_730/Y PAND2X1_52/B 0.05fF
C42732 PAND2X1_56/Y POR2X1_260/CTRL2 0.04fF
C42733 PAND2X1_207/A PAND2X1_123/Y 0.61fF
C42734 POR2X1_602/A POR2X1_296/B -0.00fF
C42735 POR2X1_502/A POR2X1_137/B 0.10fF
C42736 POR2X1_866/CTRL POR2X1_801/B 0.01fF
C42737 POR2X1_174/O PAND2X1_72/A 0.01fF
C42738 POR2X1_443/A VDD 0.04fF
C42739 POR2X1_302/Y POR2X1_831/O 0.03fF
C42740 POR2X1_709/A POR2X1_410/O 0.01fF
C42741 PAND2X1_93/B PAND2X1_387/CTRL 0.03fF
C42742 POR2X1_774/A PAND2X1_56/A 0.03fF
C42743 PAND2X1_9/O POR2X1_29/A 0.03fF
C42744 POR2X1_431/m4_208_n4# POR2X1_55/Y 0.08fF
C42745 POR2X1_257/A POR2X1_256/CTRL 0.01fF
C42746 PAND2X1_427/CTRL POR2X1_121/B 0.08fF
C42747 PAND2X1_231/CTRL D_INPUT_0 0.00fF
C42748 POR2X1_504/a_16_28# POR2X1_416/B 0.04fF
C42749 POR2X1_477/Y PAND2X1_41/B 0.01fF
C42750 POR2X1_698/CTRL2 POR2X1_32/A 0.03fF
C42751 POR2X1_23/Y PAND2X1_803/A 0.05fF
C42752 POR2X1_629/a_16_28# POR2X1_186/Y 0.03fF
C42753 POR2X1_601/Y POR2X1_601/O 0.00fF
C42754 POR2X1_68/A POR2X1_624/B 0.07fF
C42755 PAND2X1_39/B POR2X1_405/Y 0.02fF
C42756 PAND2X1_73/Y POR2X1_330/Y 0.08fF
C42757 PAND2X1_292/O POR2X1_186/B 0.03fF
C42758 POR2X1_843/CTRL2 POR2X1_343/A 0.01fF
C42759 POR2X1_67/Y PAND2X1_32/B 0.00fF
C42760 POR2X1_284/a_16_28# PAND2X1_69/A 0.01fF
C42761 POR2X1_175/A PAND2X1_73/Y 0.01fF
C42762 POR2X1_260/B POR2X1_459/CTRL2 0.09fF
C42763 POR2X1_49/Y POR2X1_29/A 0.04fF
C42764 PAND2X1_79/CTRL POR2X1_78/Y 0.01fF
C42765 POR2X1_841/B VDD 0.12fF
C42766 POR2X1_20/B PAND2X1_514/Y 0.03fF
C42767 POR2X1_630/B PAND2X1_88/Y 0.01fF
C42768 POR2X1_674/Y POR2X1_331/Y 0.01fF
C42769 POR2X1_114/CTRL2 POR2X1_499/A 0.01fF
C42770 POR2X1_809/B POR2X1_809/O 0.00fF
C42771 PAND2X1_11/Y PAND2X1_41/B 0.01fF
C42772 POR2X1_514/O POR2X1_499/A 0.01fF
C42773 POR2X1_569/O POR2X1_174/A 0.03fF
C42774 POR2X1_639/CTRL2 POR2X1_750/B 0.01fF
C42775 POR2X1_656/a_16_28# POR2X1_647/Y 0.03fF
C42776 PAND2X1_65/B PAND2X1_245/CTRL2 0.01fF
C42777 POR2X1_428/Y PAND2X1_709/CTRL2 0.01fF
C42778 POR2X1_23/Y PAND2X1_673/Y 0.10fF
C42779 POR2X1_632/B POR2X1_61/Y 0.01fF
C42780 POR2X1_644/O POR2X1_513/B 0.07fF
C42781 POR2X1_502/A PAND2X1_93/B 3.30fF
C42782 PAND2X1_545/O POR2X1_40/Y 0.03fF
C42783 POR2X1_19/a_16_28# PAND2X1_6/A 0.07fF
C42784 POR2X1_150/Y POR2X1_816/A 5.39fF
C42785 PAND2X1_550/CTRL2 POR2X1_32/A 0.03fF
C42786 POR2X1_341/A PAND2X1_316/CTRL2 0.05fF
C42787 POR2X1_411/B POR2X1_56/Y 0.03fF
C42788 POR2X1_383/A POR2X1_260/CTRL2 0.06fF
C42789 PAND2X1_307/O POR2X1_40/Y 0.03fF
C42790 PAND2X1_213/a_56_28# PAND2X1_213/A 0.00fF
C42791 POR2X1_329/A PAND2X1_549/B 0.07fF
C42792 PAND2X1_10/CTRL PAND2X1_8/Y 0.02fF
C42793 POR2X1_447/B POR2X1_568/A 0.03fF
C42794 POR2X1_480/A POR2X1_174/A 0.01fF
C42795 PAND2X1_474/a_76_28# POR2X1_43/B 0.02fF
C42796 PAND2X1_859/A POR2X1_40/Y 0.03fF
C42797 PAND2X1_56/Y POR2X1_76/O 0.26fF
C42798 POR2X1_66/B PAND2X1_815/CTRL2 0.03fF
C42799 PAND2X1_250/CTRL POR2X1_389/Y 0.00fF
C42800 POR2X1_614/A POR2X1_452/Y 0.04fF
C42801 POR2X1_271/A POR2X1_677/Y 0.00fF
C42802 POR2X1_847/B PAND2X1_820/B 0.04fF
C42803 INPUT_3 POR2X1_409/O 0.02fF
C42804 POR2X1_436/B POR2X1_435/Y 0.00fF
C42805 PAND2X1_39/B POR2X1_249/O 0.01fF
C42806 POR2X1_504/CTRL POR2X1_846/A 0.01fF
C42807 POR2X1_60/Y PAND2X1_61/Y 0.02fF
C42808 POR2X1_65/A PAND2X1_731/B 0.02fF
C42809 POR2X1_49/Y POR2X1_820/A 0.11fF
C42810 PAND2X1_77/O PAND2X1_8/Y 0.05fF
C42811 PAND2X1_626/CTRL VDD 0.00fF
C42812 POR2X1_556/A PAND2X1_60/B 2.29fF
C42813 POR2X1_114/B PAND2X1_406/a_16_344# 0.01fF
C42814 PAND2X1_803/Y POR2X1_411/B 0.02fF
C42815 POR2X1_502/A POR2X1_78/A 0.31fF
C42816 POR2X1_52/A POR2X1_89/Y 0.01fF
C42817 PAND2X1_751/O POR2X1_590/A 0.04fF
C42818 POR2X1_66/B PAND2X1_377/CTRL 0.00fF
C42819 PAND2X1_467/B PAND2X1_707/O 0.02fF
C42820 PAND2X1_576/B POR2X1_599/A 0.05fF
C42821 POR2X1_276/O POR2X1_218/Y 0.03fF
C42822 POR2X1_376/B POR2X1_226/Y 0.02fF
C42823 POR2X1_66/B POR2X1_194/B 0.05fF
C42824 POR2X1_66/B POR2X1_415/O 0.03fF
C42825 POR2X1_590/A POR2X1_802/B 0.01fF
C42826 POR2X1_447/O POR2X1_447/A 0.01fF
C42827 POR2X1_48/A PAND2X1_357/Y 0.03fF
C42828 POR2X1_821/CTRL POR2X1_40/Y 0.00fF
C42829 POR2X1_760/A PAND2X1_537/O 0.01fF
C42830 POR2X1_476/A POR2X1_391/Y 0.01fF
C42831 POR2X1_220/B POR2X1_545/A 0.03fF
C42832 POR2X1_186/Y POR2X1_742/O 0.01fF
C42833 PAND2X1_594/O POR2X1_740/Y 0.00fF
C42834 POR2X1_448/CTRL2 POR2X1_294/B 0.05fF
C42835 POR2X1_841/B PAND2X1_32/B 0.03fF
C42836 POR2X1_814/A POR2X1_186/B 0.21fF
C42837 POR2X1_388/O PAND2X1_93/B 0.01fF
C42838 PAND2X1_717/A POR2X1_129/Y 0.03fF
C42839 PAND2X1_465/CTRL2 POR2X1_7/B 0.00fF
C42840 POR2X1_781/CTRL2 POR2X1_781/A 0.01fF
C42841 POR2X1_96/A POR2X1_40/Y 0.14fF
C42842 PAND2X1_65/CTRL PAND2X1_69/A 0.03fF
C42843 POR2X1_52/A POR2X1_497/O 0.18fF
C42844 POR2X1_480/m4_208_n4# POR2X1_469/m4_208_n4# 0.13fF
C42845 PAND2X1_6/Y POR2X1_218/Y 0.10fF
C42846 POR2X1_502/A POR2X1_830/a_16_28# 0.01fF
C42847 POR2X1_78/B POR2X1_555/A 0.13fF
C42848 POR2X1_590/A POR2X1_222/Y 0.03fF
C42849 PAND2X1_139/O POR2X1_13/A 0.04fF
C42850 PAND2X1_279/CTRL POR2X1_740/Y 0.03fF
C42851 POR2X1_23/Y POR2X1_229/a_16_28# 0.04fF
C42852 POR2X1_557/A PAND2X1_9/Y 0.02fF
C42853 PAND2X1_602/Y POR2X1_102/Y 0.03fF
C42854 POR2X1_83/B PAND2X1_652/A 0.00fF
C42855 POR2X1_13/A POR2X1_278/CTRL 0.01fF
C42856 POR2X1_40/Y PAND2X1_335/O 0.05fF
C42857 POR2X1_65/A POR2X1_51/A 0.04fF
C42858 POR2X1_72/B POR2X1_7/B 0.06fF
C42859 POR2X1_614/A POR2X1_660/Y 0.03fF
C42860 POR2X1_632/B POR2X1_35/Y 0.00fF
C42861 POR2X1_517/O POR2X1_13/A 0.01fF
C42862 POR2X1_307/B VDD 0.11fF
C42863 PAND2X1_57/B POR2X1_718/A 3.02fF
C42864 POR2X1_526/CTRL POR2X1_32/A 0.01fF
C42865 PAND2X1_659/Y PAND2X1_717/A 0.03fF
C42866 POR2X1_611/CTRL2 POR2X1_293/Y 0.01fF
C42867 POR2X1_306/Y POR2X1_56/B 0.12fF
C42868 POR2X1_483/A PAND2X1_48/CTRL 0.01fF
C42869 PAND2X1_230/O POR2X1_795/B 0.08fF
C42870 POR2X1_794/B POR2X1_733/A 0.26fF
C42871 POR2X1_825/O POR2X1_42/Y 0.01fF
C42872 PAND2X1_93/B POR2X1_140/m4_208_n4# 0.12fF
C42873 POR2X1_556/A POR2X1_787/a_16_28# -0.00fF
C42874 POR2X1_48/A POR2X1_278/A 0.01fF
C42875 POR2X1_52/A POR2X1_290/CTRL 0.01fF
C42876 POR2X1_719/O PAND2X1_93/B 0.02fF
C42877 POR2X1_555/B POR2X1_631/B 0.03fF
C42878 PAND2X1_56/Y PAND2X1_279/O 0.02fF
C42879 POR2X1_40/Y PAND2X1_506/CTRL 0.01fF
C42880 POR2X1_278/O PAND2X1_35/Y 0.01fF
C42881 POR2X1_52/A POR2X1_226/Y 0.01fF
C42882 INPUT_7 INPUT_5 0.05fF
C42883 POR2X1_672/O POR2X1_102/Y 0.01fF
C42884 POR2X1_294/O POR2X1_260/A 0.01fF
C42885 PAND2X1_474/CTRL POR2X1_153/Y 0.11fF
C42886 PAND2X1_347/Y PAND2X1_568/CTRL2 0.01fF
C42887 PAND2X1_140/A POR2X1_48/A 0.05fF
C42888 POR2X1_852/B POR2X1_785/A 0.07fF
C42889 PAND2X1_73/Y PAND2X1_519/a_76_28# 0.03fF
C42890 PAND2X1_474/A POR2X1_494/Y 0.03fF
C42891 PAND2X1_469/B PAND2X1_556/a_56_28# 0.00fF
C42892 POR2X1_150/Y PAND2X1_357/CTRL 0.07fF
C42893 PAND2X1_90/A POR2X1_860/A 0.03fF
C42894 POR2X1_45/Y PAND2X1_390/Y 0.03fF
C42895 POR2X1_590/A POR2X1_532/A 3.69fF
C42896 POR2X1_481/A PAND2X1_738/Y 0.05fF
C42897 POR2X1_41/B POR2X1_511/Y 0.07fF
C42898 POR2X1_528/Y POR2X1_48/A 0.10fF
C42899 PAND2X1_55/Y POR2X1_402/CTRL2 0.01fF
C42900 POR2X1_500/A PAND2X1_316/CTRL2 0.00fF
C42901 POR2X1_407/A POR2X1_843/m4_208_n4# 0.12fF
C42902 PAND2X1_284/O POR2X1_279/Y 0.01fF
C42903 POR2X1_338/O POR2X1_66/A 0.01fF
C42904 POR2X1_88/Y INPUT_0 0.05fF
C42905 POR2X1_52/A POR2X1_238/O 0.02fF
C42906 POR2X1_20/B POR2X1_75/Y 0.02fF
C42907 POR2X1_814/B POR2X1_732/B 0.10fF
C42908 POR2X1_634/A PAND2X1_69/A 0.08fF
C42909 PAND2X1_824/a_16_344# POR2X1_66/A 0.02fF
C42910 POR2X1_251/Y VDD 0.18fF
C42911 PAND2X1_674/O POR2X1_186/Y 0.08fF
C42912 POR2X1_60/A PAND2X1_341/A 0.03fF
C42913 POR2X1_541/B PAND2X1_48/A 1.32fF
C42914 PAND2X1_412/CTRL2 POR2X1_391/Y 0.01fF
C42915 POR2X1_859/A POR2X1_415/O 0.01fF
C42916 PAND2X1_272/a_16_344# PAND2X1_60/B 0.01fF
C42917 PAND2X1_848/B PAND2X1_859/A 0.01fF
C42918 POR2X1_78/B PAND2X1_89/O 0.03fF
C42919 PAND2X1_460/Y PAND2X1_472/B 0.04fF
C42920 POR2X1_60/a_56_344# POR2X1_60/A 0.00fF
C42921 POR2X1_308/CTRL2 PAND2X1_55/Y 0.00fF
C42922 POR2X1_440/Y POR2X1_220/B 0.03fF
C42923 POR2X1_66/B POR2X1_21/CTRL2 0.03fF
C42924 PAND2X1_793/Y POR2X1_79/A 0.04fF
C42925 PAND2X1_241/Y POR2X1_14/Y 0.13fF
C42926 POR2X1_60/A POR2X1_91/Y 0.07fF
C42927 POR2X1_255/Y PAND2X1_541/O -0.00fF
C42928 PAND2X1_207/CTRL2 POR2X1_153/Y 0.01fF
C42929 POR2X1_48/A POR2X1_394/CTRL2 0.03fF
C42930 POR2X1_68/A POR2X1_849/O 0.16fF
C42931 POR2X1_593/B POR2X1_804/A 0.05fF
C42932 PAND2X1_241/Y PAND2X1_453/A 0.00fF
C42933 POR2X1_40/CTRL2 POR2X1_32/A 0.03fF
C42934 PAND2X1_793/Y PAND2X1_468/CTRL2 0.01fF
C42935 PAND2X1_329/CTRL POR2X1_149/A 0.00fF
C42936 POR2X1_201/a_56_344# PAND2X1_88/Y 0.00fF
C42937 POR2X1_146/O POR2X1_669/B 0.00fF
C42938 POR2X1_651/m4_208_n4# PAND2X1_90/Y 0.09fF
C42939 POR2X1_72/O POR2X1_816/A 0.01fF
C42940 POR2X1_62/Y PAND2X1_206/A 0.01fF
C42941 POR2X1_78/B POR2X1_659/CTRL 0.02fF
C42942 POR2X1_119/Y PAND2X1_203/O 0.22fF
C42943 INPUT_4 INPUT_5 0.92fF
C42944 POR2X1_251/CTRL POR2X1_387/Y 0.01fF
C42945 PAND2X1_632/CTRL POR2X1_496/Y 0.03fF
C42946 POR2X1_66/B POR2X1_537/B 0.02fF
C42947 POR2X1_43/B POR2X1_497/Y 0.01fF
C42948 PAND2X1_90/A POR2X1_327/CTRL2 0.03fF
C42949 POR2X1_750/B PAND2X1_312/CTRL 0.00fF
C42950 POR2X1_98/B PAND2X1_41/B 0.02fF
C42951 POR2X1_128/A POR2X1_318/A 0.04fF
C42952 POR2X1_556/A POR2X1_554/O 0.08fF
C42953 POR2X1_383/A PAND2X1_279/O -0.01fF
C42954 POR2X1_499/A PAND2X1_136/O 0.06fF
C42955 POR2X1_853/A POR2X1_570/CTRL2 0.01fF
C42956 POR2X1_65/A PAND2X1_113/O 0.01fF
C42957 POR2X1_625/Y POR2X1_42/Y 1.75fF
C42958 POR2X1_49/Y POR2X1_583/O 0.11fF
C42959 POR2X1_114/B VDD 0.78fF
C42960 POR2X1_482/Y POR2X1_283/A 0.00fF
C42961 PAND2X1_465/B POR2X1_372/Y 0.02fF
C42962 POR2X1_188/A POR2X1_537/B 0.03fF
C42963 POR2X1_608/O POR2X1_712/Y 0.03fF
C42964 POR2X1_40/O POR2X1_83/B 0.16fF
C42965 POR2X1_10/O POR2X1_669/B 0.01fF
C42966 POR2X1_40/Y POR2X1_7/A 0.10fF
C42967 POR2X1_330/Y PAND2X1_163/O 0.02fF
C42968 POR2X1_52/A PAND2X1_736/Y 0.01fF
C42969 POR2X1_557/A POR2X1_267/A 0.07fF
C42970 POR2X1_654/CTRL POR2X1_725/Y 0.01fF
C42971 POR2X1_356/A PAND2X1_23/Y 0.05fF
C42972 PAND2X1_95/B POR2X1_638/CTRL 0.01fF
C42973 PAND2X1_691/Y POR2X1_829/CTRL 0.01fF
C42974 POR2X1_40/Y PAND2X1_130/O 0.01fF
C42975 PAND2X1_115/B PAND2X1_724/B 0.03fF
C42976 POR2X1_573/a_16_28# POR2X1_576/Y 0.01fF
C42977 POR2X1_306/CTRL POR2X1_236/Y 0.01fF
C42978 PAND2X1_863/B PAND2X1_794/B 0.03fF
C42979 PAND2X1_52/Y POR2X1_510/Y 0.03fF
C42980 POR2X1_48/A POR2X1_117/Y 0.01fF
C42981 POR2X1_72/B PAND2X1_123/CTRL 0.01fF
C42982 POR2X1_130/A PAND2X1_69/A 0.13fF
C42983 POR2X1_262/Y PAND2X1_339/O 0.01fF
C42984 POR2X1_668/Y POR2X1_816/A 0.01fF
C42985 PAND2X1_623/O POR2X1_129/Y 0.02fF
C42986 POR2X1_730/Y POR2X1_467/Y 0.07fF
C42987 PAND2X1_93/B POR2X1_188/Y 0.03fF
C42988 POR2X1_649/B VDD 0.41fF
C42989 PAND2X1_620/a_16_344# POR2X1_422/Y 0.02fF
C42990 POR2X1_668/Y D_INPUT_1 0.03fF
C42991 POR2X1_259/A POR2X1_259/CTRL 0.01fF
C42992 POR2X1_536/a_16_28# POR2X1_102/Y 0.03fF
C42993 PAND2X1_73/Y POR2X1_715/A 0.02fF
C42994 POR2X1_458/B VDD 0.00fF
C42995 PAND2X1_787/Y POR2X1_387/Y 0.10fF
C42996 PAND2X1_653/Y POR2X1_13/A 0.12fF
C42997 POR2X1_708/O PAND2X1_32/B 0.01fF
C42998 POR2X1_566/A PAND2X1_69/A 2.90fF
C42999 POR2X1_131/CTRL PAND2X1_137/Y 0.06fF
C43000 PAND2X1_645/a_16_344# PAND2X1_645/B 0.02fF
C43001 POR2X1_52/A POR2X1_56/Y 0.03fF
C43002 POR2X1_283/A POR2X1_106/Y 0.03fF
C43003 PAND2X1_786/CTRL2 POR2X1_394/A 0.05fF
C43004 POR2X1_134/Y POR2X1_96/A 0.60fF
C43005 PAND2X1_649/A PAND2X1_590/CTRL 0.01fF
C43006 PAND2X1_94/A PAND2X1_46/a_56_28# 0.00fF
C43007 POR2X1_186/Y POR2X1_727/m4_208_n4# 0.04fF
C43008 POR2X1_614/A POR2X1_786/A 0.36fF
C43009 POR2X1_293/Y POR2X1_310/CTRL 0.02fF
C43010 POR2X1_559/CTRL PAND2X1_90/A 0.01fF
C43011 POR2X1_785/A PAND2X1_504/a_16_344# 0.02fF
C43012 PAND2X1_568/B VDD 0.73fF
C43013 POR2X1_539/A POR2X1_733/O 0.00fF
C43014 POR2X1_346/B POR2X1_404/a_56_344# 0.00fF
C43015 POR2X1_43/B PAND2X1_466/a_16_344# 0.01fF
C43016 POR2X1_816/Y POR2X1_39/B 0.15fF
C43017 POR2X1_254/Y POR2X1_702/CTRL 0.03fF
C43018 PAND2X1_329/CTRL VDD 0.00fF
C43019 POR2X1_288/A POR2X1_734/O 0.00fF
C43020 POR2X1_693/a_16_28# POR2X1_73/Y 0.03fF
C43021 POR2X1_786/A POR2X1_38/B 0.23fF
C43022 PAND2X1_563/B PAND2X1_346/Y 0.03fF
C43023 POR2X1_222/A VDD 0.64fF
C43024 POR2X1_502/A PAND2X1_306/O 0.08fF
C43025 POR2X1_283/A PAND2X1_580/B 0.03fF
C43026 PAND2X1_209/A PAND2X1_213/A 0.06fF
C43027 PAND2X1_461/CTRL2 D_INPUT_0 0.00fF
C43028 POR2X1_857/B POR2X1_532/A 0.03fF
C43029 POR2X1_43/B POR2X1_118/CTRL2 0.01fF
C43030 PAND2X1_94/A POR2X1_476/Y 0.01fF
C43031 PAND2X1_659/Y PAND2X1_200/CTRL2 0.00fF
C43032 PAND2X1_724/B POR2X1_73/Y 0.00fF
C43033 POR2X1_78/A POR2X1_188/Y 0.03fF
C43034 PAND2X1_65/B POR2X1_218/a_16_28# 0.03fF
C43035 POR2X1_97/B PAND2X1_20/A 0.02fF
C43036 POR2X1_104/CTRL2 POR2X1_4/Y 0.03fF
C43037 POR2X1_618/O POR2X1_382/Y 0.01fF
C43038 PAND2X1_317/Y POR2X1_258/O 0.03fF
C43039 POR2X1_66/B PAND2X1_48/A 0.10fF
C43040 POR2X1_57/A POR2X1_680/Y 0.03fF
C43041 POR2X1_119/Y PAND2X1_404/CTRL 0.01fF
C43042 PAND2X1_6/Y POR2X1_68/A 1.16fF
C43043 POR2X1_52/A PAND2X1_803/Y 0.03fF
C43044 POR2X1_364/A D_GATE_222 0.07fF
C43045 POR2X1_523/Y POR2X1_844/B 0.07fF
C43046 PAND2X1_85/Y POR2X1_260/A 0.07fF
C43047 POR2X1_280/CTRL2 PAND2X1_552/B 0.00fF
C43048 PAND2X1_550/B PAND2X1_549/CTRL 0.01fF
C43049 PAND2X1_57/B POR2X1_725/Y 0.07fF
C43050 POR2X1_82/CTRL INPUT_1 0.01fF
C43051 POR2X1_164/Y VDD 0.10fF
C43052 PAND2X1_139/CTRL2 POR2X1_102/Y 0.01fF
C43053 PAND2X1_26/A PAND2X1_52/B 0.05fF
C43054 PAND2X1_90/Y POR2X1_721/O 0.16fF
C43055 POR2X1_114/B PAND2X1_32/B 0.03fF
C43056 POR2X1_220/O PAND2X1_52/B 0.01fF
C43057 PAND2X1_707/Y POR2X1_526/Y 0.00fF
C43058 POR2X1_188/A PAND2X1_48/A 0.03fF
C43059 POR2X1_551/O VDD 0.00fF
C43060 POR2X1_511/Y PAND2X1_308/Y 0.03fF
C43061 POR2X1_590/A POR2X1_510/CTRL2 0.00fF
C43062 PAND2X1_793/Y PAND2X1_574/CTRL2 0.01fF
C43063 POR2X1_687/A POR2X1_220/Y 0.01fF
C43064 POR2X1_49/Y POR2X1_146/Y 0.06fF
C43065 POR2X1_785/a_76_344# POR2X1_566/B 0.03fF
C43066 POR2X1_565/B POR2X1_550/Y 0.00fF
C43067 POR2X1_546/B POR2X1_550/Y 0.01fF
C43068 POR2X1_300/CTRL2 PAND2X1_349/A 0.01fF
C43069 PAND2X1_553/a_76_28# POR2X1_55/Y 0.01fF
C43070 PAND2X1_809/B PAND2X1_223/B 0.05fF
C43071 POR2X1_38/Y PAND2X1_734/CTRL2 0.00fF
C43072 PAND2X1_41/B PAND2X1_328/CTRL2 0.01fF
C43073 POR2X1_82/CTRL POR2X1_153/Y 0.03fF
C43074 POR2X1_743/a_56_344# POR2X1_153/Y 0.00fF
C43075 POR2X1_8/Y INPUT_0 0.07fF
C43076 POR2X1_213/a_16_28# POR2X1_210/Y 0.03fF
C43077 PAND2X1_653/Y PAND2X1_661/B 0.14fF
C43078 PAND2X1_433/O POR2X1_832/A 0.02fF
C43079 PAND2X1_57/B POR2X1_596/O 0.16fF
C43080 POR2X1_771/O PAND2X1_32/B 0.01fF
C43081 PAND2X1_96/B POR2X1_556/Y 0.03fF
C43082 POR2X1_360/A PAND2X1_94/A 0.04fF
C43083 PAND2X1_23/Y POR2X1_569/A 0.07fF
C43084 PAND2X1_752/Y POR2X1_532/A 0.02fF
C43085 POR2X1_13/A PAND2X1_563/A 0.03fF
C43086 POR2X1_458/B PAND2X1_32/B 0.03fF
C43087 POR2X1_349/CTRL PAND2X1_65/Y 0.00fF
C43088 PAND2X1_69/A PAND2X1_150/O 0.15fF
C43089 POR2X1_119/Y PAND2X1_541/a_16_344# 0.02fF
C43090 POR2X1_566/A PAND2X1_824/B 0.10fF
C43091 POR2X1_122/CTRL VDD -0.00fF
C43092 PAND2X1_848/B POR2X1_7/A 0.11fF
C43093 PAND2X1_663/CTRL POR2X1_413/A 0.01fF
C43094 POR2X1_667/A POR2X1_39/B 0.03fF
C43095 PAND2X1_735/Y POR2X1_394/A 0.10fF
C43096 PAND2X1_57/B POR2X1_559/A 0.12fF
C43097 POR2X1_355/B POR2X1_209/CTRL2 0.01fF
C43098 D_INPUT_3 POR2X1_63/a_16_28# 0.09fF
C43099 PAND2X1_48/B POR2X1_463/Y 0.05fF
C43100 POR2X1_367/m4_208_n4# POR2X1_568/Y 0.08fF
C43101 POR2X1_41/B POR2X1_129/Y 0.07fF
C43102 PAND2X1_605/O POR2X1_42/Y 0.02fF
C43103 POR2X1_318/A POR2X1_140/O 0.03fF
C43104 POR2X1_92/O POR2X1_38/Y 0.01fF
C43105 POR2X1_16/A PAND2X1_649/CTRL 0.01fF
C43106 POR2X1_43/B POR2X1_310/Y 0.05fF
C43107 POR2X1_222/A PAND2X1_32/B 0.03fF
C43108 POR2X1_57/A PAND2X1_388/Y 0.06fF
C43109 POR2X1_486/O POR2X1_556/A 0.01fF
C43110 POR2X1_178/Y POR2X1_183/Y 0.01fF
C43111 POR2X1_96/A POR2X1_533/O 0.01fF
C43112 PAND2X1_55/Y POR2X1_507/A 0.47fF
C43113 PAND2X1_141/a_16_344# POR2X1_39/B 0.02fF
C43114 PAND2X1_572/CTRL2 PAND2X1_656/A 0.01fF
C43115 POR2X1_383/A POR2X1_68/B 0.09fF
C43116 INPUT_0 POR2X1_385/Y 0.04fF
C43117 POR2X1_510/Y POR2X1_724/A 0.04fF
C43118 POR2X1_301/CTRL POR2X1_260/A 0.01fF
C43119 PAND2X1_859/B POR2X1_394/A 0.10fF
C43120 POR2X1_394/A PAND2X1_493/Y 0.18fF
C43121 PAND2X1_72/m4_208_n4# PAND2X1_60/B 0.17fF
C43122 POR2X1_57/A PAND2X1_549/B 1.18fF
C43123 INPUT_1 POR2X1_20/Y 0.03fF
C43124 POR2X1_307/A PAND2X1_305/CTRL 0.00fF
C43125 PAND2X1_481/CTRL2 D_GATE_741 0.01fF
C43126 D_INPUT_1 POR2X1_276/Y 0.03fF
C43127 POR2X1_345/CTRL2 PAND2X1_6/Y 0.00fF
C43128 POR2X1_41/B PAND2X1_659/Y 0.03fF
C43129 POR2X1_52/A POR2X1_824/CTRL2 0.01fF
C43130 POR2X1_276/A PAND2X1_60/B 0.02fF
C43131 PAND2X1_96/B POR2X1_259/a_16_28# 0.02fF
C43132 POR2X1_852/A POR2X1_191/Y 0.33fF
C43133 POR2X1_740/Y POR2X1_737/A 0.03fF
C43134 POR2X1_283/A PAND2X1_349/A 0.03fF
C43135 POR2X1_41/B POR2X1_96/Y 0.03fF
C43136 POR2X1_407/A PAND2X1_310/CTRL 0.00fF
C43137 PAND2X1_180/CTRL POR2X1_77/Y 0.01fF
C43138 PAND2X1_531/CTRL2 D_INPUT_1 0.05fF
C43139 PAND2X1_226/a_76_28# POR2X1_192/B 0.05fF
C43140 PAND2X1_61/Y PAND2X1_351/A 0.79fF
C43141 POR2X1_511/Y POR2X1_77/Y 21.11fF
C43142 POR2X1_137/Y POR2X1_260/A 0.03fF
C43143 POR2X1_366/Y POR2X1_540/Y 0.10fF
C43144 PAND2X1_543/CTRL POR2X1_77/Y 0.00fF
C43145 PAND2X1_301/CTRL POR2X1_91/Y 0.03fF
C43146 POR2X1_41/B PAND2X1_857/a_56_28# 0.00fF
C43147 PAND2X1_8/Y PAND2X1_102/a_16_344# 0.02fF
C43148 PAND2X1_101/B PAND2X1_101/O 0.00fF
C43149 POR2X1_577/a_16_28# POR2X1_569/Y -0.00fF
C43150 POR2X1_579/B POR2X1_576/Y 0.27fF
C43151 POR2X1_383/A POR2X1_561/O 0.03fF
C43152 INPUT_1 POR2X1_713/B 0.05fF
C43153 POR2X1_158/Y PAND2X1_210/a_76_28# 0.02fF
C43154 POR2X1_667/CTRL2 D_INPUT_0 0.09fF
C43155 PAND2X1_94/A PAND2X1_748/CTRL2 0.00fF
C43156 POR2X1_863/A POR2X1_186/Y 0.07fF
C43157 POR2X1_775/CTRL2 POR2X1_191/Y 0.18fF
C43158 POR2X1_68/B PAND2X1_71/Y 0.01fF
C43159 POR2X1_66/Y PAND2X1_43/CTRL 0.01fF
C43160 POR2X1_305/CTRL POR2X1_7/B 0.01fF
C43161 POR2X1_169/O POR2X1_568/Y 0.03fF
C43162 POR2X1_816/A POR2X1_749/Y 0.00fF
C43163 POR2X1_461/Y POR2X1_848/Y 0.01fF
C43164 PAND2X1_575/a_76_28# POR2X1_394/A 0.05fF
C43165 POR2X1_228/m4_208_n4# POR2X1_193/m4_208_n4# 0.13fF
C43166 POR2X1_633/A POR2X1_9/Y 0.01fF
C43167 D_INPUT_1 POR2X1_749/Y 0.03fF
C43168 PAND2X1_808/Y POR2X1_767/Y 0.61fF
C43169 PAND2X1_115/CTRL2 POR2X1_416/B 0.01fF
C43170 POR2X1_356/A POR2X1_711/Y 0.28fF
C43171 PAND2X1_353/CTRL PAND2X1_303/Y 0.01fF
C43172 PAND2X1_353/O PAND2X1_308/Y 0.04fF
C43173 PAND2X1_443/a_16_344# POR2X1_441/Y 0.02fF
C43174 POR2X1_369/CTRL2 POR2X1_315/Y 0.05fF
C43175 PAND2X1_656/A PAND2X1_123/Y 0.03fF
C43176 PAND2X1_48/B POR2X1_736/A 0.12fF
C43177 POR2X1_57/A POR2X1_397/CTRL 0.01fF
C43178 POR2X1_566/CTRL POR2X1_854/B 0.01fF
C43179 PAND2X1_569/B POR2X1_394/A 0.07fF
C43180 POR2X1_852/a_16_28# POR2X1_568/A 0.03fF
C43181 POR2X1_326/A POR2X1_383/A 0.02fF
C43182 POR2X1_394/A POR2X1_158/B 0.02fF
C43183 POR2X1_833/A POR2X1_260/A 0.01fF
C43184 PAND2X1_319/B PAND2X1_352/CTRL 0.03fF
C43185 POR2X1_411/B PAND2X1_771/Y 0.05fF
C43186 POR2X1_68/A POR2X1_632/Y 0.57fF
C43187 POR2X1_447/B PAND2X1_824/CTRL 0.00fF
C43188 PAND2X1_124/CTRL2 PAND2X1_123/Y 0.02fF
C43189 POR2X1_753/Y POR2X1_846/Y 0.08fF
C43190 PAND2X1_779/CTRL PAND2X1_550/B 0.01fF
C43191 PAND2X1_821/CTRL2 PAND2X1_52/B 0.00fF
C43192 POR2X1_725/Y POR2X1_512/CTRL2 0.05fF
C43193 PAND2X1_23/Y POR2X1_509/O 0.01fF
C43194 PAND2X1_360/Y PAND2X1_343/CTRL 0.01fF
C43195 PAND2X1_405/CTRL2 POR2X1_5/Y 0.01fF
C43196 PAND2X1_23/Y PAND2X1_72/A 0.13fF
C43197 POR2X1_542/B POR2X1_542/a_16_28# -0.00fF
C43198 PAND2X1_273/CTRL2 POR2X1_717/B 0.01fF
C43199 POR2X1_318/A PAND2X1_136/CTRL 0.04fF
C43200 POR2X1_456/B POR2X1_703/CTRL 0.01fF
C43201 POR2X1_20/B POR2X1_279/CTRL2 0.00fF
C43202 POR2X1_1/a_16_28# PAND2X1_18/B 0.06fF
C43203 POR2X1_186/a_16_28# POR2X1_353/A 0.03fF
C43204 POR2X1_71/CTRL POR2X1_394/A 0.04fF
C43205 PAND2X1_94/A POR2X1_571/Y 0.03fF
C43206 POR2X1_276/Y POR2X1_362/CTRL2 0.01fF
C43207 POR2X1_435/a_16_28# POR2X1_296/B 0.10fF
C43208 PAND2X1_18/B POR2X1_260/A 0.11fF
C43209 POR2X1_417/Y PAND2X1_464/B 0.02fF
C43210 PAND2X1_761/a_16_344# D_INPUT_0 0.02fF
C43211 POR2X1_68/A PAND2X1_52/B 11.27fF
C43212 POR2X1_149/CTRL2 POR2X1_78/A 0.03fF
C43213 POR2X1_638/Y PAND2X1_56/A 0.01fF
C43214 PAND2X1_849/B PAND2X1_101/B 0.00fF
C43215 POR2X1_760/A POR2X1_40/Y 0.08fF
C43216 POR2X1_597/O POR2X1_761/A 0.01fF
C43217 POR2X1_186/B POR2X1_151/Y 0.01fF
C43218 POR2X1_411/B PAND2X1_719/Y 0.57fF
C43219 POR2X1_48/A POR2X1_817/O 0.07fF
C43220 PAND2X1_269/CTRL POR2X1_236/Y 0.01fF
C43221 POR2X1_245/Y POR2X1_39/B 0.02fF
C43222 POR2X1_66/B POR2X1_461/Y 0.01fF
C43223 POR2X1_383/A POR2X1_862/CTRL2 0.01fF
C43224 PAND2X1_127/a_16_344# POR2X1_567/A -0.03fF
C43225 POR2X1_705/B PAND2X1_41/B 0.03fF
C43226 PAND2X1_88/Y POR2X1_555/a_76_344# 0.00fF
C43227 POR2X1_147/O POR2X1_532/A 0.01fF
C43228 POR2X1_90/Y POR2X1_167/Y 0.07fF
C43229 POR2X1_257/A PAND2X1_161/CTRL 0.01fF
C43230 POR2X1_567/B POR2X1_434/A 0.03fF
C43231 POR2X1_250/Y PAND2X1_362/B 0.17fF
C43232 POR2X1_816/m4_208_n4# POR2X1_750/B 0.08fF
C43233 POR2X1_77/Y PAND2X1_112/CTRL2 0.01fF
C43234 POR2X1_604/CTRL POR2X1_72/B 0.01fF
C43235 POR2X1_606/O POR2X1_121/B 0.03fF
C43236 POR2X1_406/Y PAND2X1_266/O 0.08fF
C43237 POR2X1_590/A POR2X1_458/O 0.01fF
C43238 POR2X1_670/CTRL POR2X1_20/B 0.01fF
C43239 POR2X1_472/CTRL PAND2X1_52/B 0.01fF
C43240 POR2X1_20/B PAND2X1_562/B 0.07fF
C43241 PAND2X1_449/O POR2X1_511/Y 0.01fF
C43242 PAND2X1_64/CTRL PAND2X1_11/Y 0.09fF
C43243 POR2X1_493/A POR2X1_78/A 0.01fF
C43244 POR2X1_858/CTRL2 POR2X1_590/A 0.03fF
C43245 POR2X1_65/A PAND2X1_446/Y 0.03fF
C43246 POR2X1_567/B POR2X1_857/CTRL 0.28fF
C43247 POR2X1_564/B POR2X1_564/a_16_28# -0.00fF
C43248 PAND2X1_246/O INPUT_0 0.05fF
C43249 POR2X1_815/A POR2X1_750/A 0.07fF
C43250 PAND2X1_227/O POR2X1_236/Y 0.04fF
C43251 PAND2X1_39/B POR2X1_403/CTRL 0.04fF
C43252 PAND2X1_569/B PAND2X1_326/CTRL 0.02fF
C43253 PAND2X1_139/m4_208_n4# POR2X1_150/Y 0.15fF
C43254 PAND2X1_124/Y PAND2X1_195/CTRL 0.01fF
C43255 PAND2X1_65/B POR2X1_776/A 0.12fF
C43256 POR2X1_48/A POR2X1_667/A 5.62fF
C43257 PAND2X1_507/CTRL POR2X1_39/B 0.03fF
C43258 PAND2X1_717/A POR2X1_293/Y 0.28fF
C43259 POR2X1_9/Y POR2X1_617/a_16_28# 0.06fF
C43260 POR2X1_48/A POR2X1_607/A 0.01fF
C43261 PAND2X1_704/CTRL2 POR2X1_77/Y 0.01fF
C43262 PAND2X1_476/CTRL2 PAND2X1_571/A 0.01fF
C43263 PAND2X1_474/Y POR2X1_20/B 0.16fF
C43264 PAND2X1_73/Y PAND2X1_413/O 0.11fF
C43265 POR2X1_52/A PAND2X1_97/Y 0.01fF
C43266 POR2X1_49/Y PAND2X1_444/CTRL -0.05fF
C43267 POR2X1_260/B POR2X1_734/A 0.03fF
C43268 PAND2X1_630/B POR2X1_90/Y 0.03fF
C43269 POR2X1_119/Y POR2X1_518/CTRL 0.11fF
C43270 PAND2X1_841/O POR2X1_329/A 0.06fF
C43271 D_INPUT_5 PAND2X1_18/CTRL 0.01fF
C43272 POR2X1_228/Y POR2X1_303/B 0.01fF
C43273 POR2X1_826/Y VDD 0.15fF
C43274 PAND2X1_170/O POR2X1_39/B 0.01fF
C43275 PAND2X1_833/O POR2X1_257/A 0.03fF
C43276 PAND2X1_159/CTRL2 POR2X1_29/A 0.01fF
C43277 POR2X1_13/A POR2X1_20/B 0.25fF
C43278 POR2X1_129/Y POR2X1_77/Y 0.08fF
C43279 POR2X1_479/B POR2X1_288/m4_208_n4# 0.01fF
C43280 POR2X1_461/Y POR2X1_859/A 0.20fF
C43281 POR2X1_428/Y POR2X1_701/Y 0.00fF
C43282 PAND2X1_410/CTRL POR2X1_236/Y 0.01fF
C43283 POR2X1_106/CTRL POR2X1_251/A 0.01fF
C43284 POR2X1_117/O POR2X1_48/A 0.01fF
C43285 PAND2X1_94/Y PAND2X1_60/B 0.03fF
C43286 POR2X1_814/B POR2X1_466/A 0.10fF
C43287 POR2X1_485/Y PAND2X1_707/Y 0.00fF
C43288 PAND2X1_108/a_76_28# PAND2X1_39/B 0.01fF
C43289 PAND2X1_659/Y POR2X1_77/Y 0.03fF
C43290 PAND2X1_340/B POR2X1_88/Y 0.07fF
C43291 POR2X1_629/CTRL VDD 0.00fF
C43292 POR2X1_856/B PAND2X1_65/B 0.10fF
C43293 POR2X1_112/O POR2X1_632/Y 0.02fF
C43294 POR2X1_48/A PAND2X1_712/B 0.28fF
C43295 PAND2X1_459/CTRL PAND2X1_58/A 0.11fF
C43296 POR2X1_411/B POR2X1_42/Y 13.18fF
C43297 POR2X1_82/CTRL2 POR2X1_409/B 0.01fF
C43298 POR2X1_311/Y POR2X1_40/Y 0.03fF
C43299 PAND2X1_675/A POR2X1_150/Y 0.79fF
C43300 POR2X1_852/B PAND2X1_39/CTRL 0.07fF
C43301 POR2X1_88/a_76_344# INPUT_0 0.02fF
C43302 PAND2X1_469/B POR2X1_150/Y 0.21fF
C43303 POR2X1_96/Y POR2X1_77/Y 0.01fF
C43304 POR2X1_411/B PAND2X1_562/CTRL 0.01fF
C43305 POR2X1_554/B POR2X1_804/A 0.01fF
C43306 POR2X1_61/Y POR2X1_555/B 0.03fF
C43307 PAND2X1_205/A PAND2X1_795/B 0.01fF
C43308 POR2X1_474/CTRL2 PAND2X1_41/B 0.00fF
C43309 POR2X1_240/A PAND2X1_88/Y 0.01fF
C43310 POR2X1_640/Y POR2X1_634/A 0.12fF
C43311 POR2X1_114/B POR2X1_475/CTRL2 0.04fF
C43312 POR2X1_66/Y POR2X1_740/Y 0.25fF
C43313 POR2X1_411/B POR2X1_309/Y 0.44fF
C43314 POR2X1_366/Y POR2X1_445/A 0.10fF
C43315 POR2X1_112/CTRL PAND2X1_72/A 0.01fF
C43316 POR2X1_61/Y PAND2X1_394/CTRL 0.07fF
C43317 PAND2X1_392/O VDD 0.00fF
C43318 POR2X1_662/O PAND2X1_55/Y 0.15fF
C43319 PAND2X1_95/B PAND2X1_26/A 0.05fF
C43320 POR2X1_593/B POR2X1_794/B 0.03fF
C43321 PAND2X1_435/Y PAND2X1_499/Y 0.91fF
C43322 PAND2X1_761/CTRL2 PAND2X1_32/B 0.01fF
C43323 POR2X1_86/a_56_344# POR2X1_85/Y 0.01fF
C43324 PAND2X1_675/O POR2X1_416/B 0.05fF
C43325 POR2X1_480/A POR2X1_121/B 0.15fF
C43326 POR2X1_262/Y PAND2X1_716/a_76_28# 0.02fF
C43327 POR2X1_490/Y PAND2X1_228/CTRL 0.01fF
C43328 POR2X1_251/A PAND2X1_220/Y 0.03fF
C43329 POR2X1_432/O VDD 0.00fF
C43330 POR2X1_43/B PAND2X1_469/CTRL 0.01fF
C43331 POR2X1_29/A PAND2X1_8/Y 0.73fF
C43332 POR2X1_48/A POR2X1_252/O 0.02fF
C43333 POR2X1_41/B POR2X1_37/Y 0.04fF
C43334 POR2X1_61/Y POR2X1_330/Y 0.07fF
C43335 POR2X1_590/A POR2X1_207/O 0.16fF
C43336 POR2X1_48/A PAND2X1_254/CTRL2 0.01fF
C43337 POR2X1_23/Y PAND2X1_254/CTRL 0.03fF
C43338 POR2X1_341/A POR2X1_541/CTRL2 0.03fF
C43339 POR2X1_465/CTRL2 POR2X1_569/A 0.02fF
C43340 PAND2X1_48/B POR2X1_270/Y 0.03fF
C43341 POR2X1_169/A PAND2X1_52/B 0.03fF
C43342 PAND2X1_39/B POR2X1_644/A 0.07fF
C43343 POR2X1_834/CTRL POR2X1_513/B 0.01fF
C43344 POR2X1_52/A POR2X1_754/Y 0.07fF
C43345 POR2X1_416/B POR2X1_747/CTRL 0.00fF
C43346 PAND2X1_354/A PAND2X1_563/B 0.00fF
C43347 POR2X1_355/B POR2X1_470/a_16_28# 0.02fF
C43348 PAND2X1_564/B PAND2X1_564/O 0.01fF
C43349 PAND2X1_859/A POR2X1_5/Y 0.03fF
C43350 POR2X1_77/Y PAND2X1_333/Y 0.06fF
C43351 POR2X1_725/O POR2X1_711/Y 0.01fF
C43352 POR2X1_327/Y POR2X1_458/Y 0.07fF
C43353 POR2X1_260/B POR2X1_786/Y 0.15fF
C43354 PAND2X1_57/B POR2X1_811/B 0.03fF
C43355 PAND2X1_863/B POR2X1_83/B 0.01fF
C43356 POR2X1_423/CTRL POR2X1_372/Y 0.04fF
C43357 POR2X1_669/B POR2X1_617/CTRL 0.32fF
C43358 POR2X1_786/A POR2X1_590/A 0.03fF
C43359 POR2X1_66/A POR2X1_222/Y 0.03fF
C43360 PAND2X1_72/A POR2X1_711/Y 0.07fF
C43361 POR2X1_124/O POR2X1_78/A 0.02fF
C43362 PAND2X1_220/A POR2X1_55/Y 0.01fF
C43363 POR2X1_300/CTRL2 POR2X1_32/A 0.02fF
C43364 PAND2X1_65/B PAND2X1_386/O 0.03fF
C43365 POR2X1_83/B POR2X1_669/CTRL 0.01fF
C43366 POR2X1_67/Y POR2X1_751/Y 0.02fF
C43367 PAND2X1_443/CTRL2 POR2X1_91/Y 0.01fF
C43368 POR2X1_68/A POR2X1_632/a_16_28# 0.03fF
C43369 PAND2X1_93/B POR2X1_243/CTRL2 0.01fF
C43370 POR2X1_848/A POR2X1_90/Y 0.01fF
C43371 POR2X1_78/A POR2X1_725/a_16_28# 0.01fF
C43372 POR2X1_20/B PAND2X1_510/B 2.23fF
C43373 PAND2X1_776/Y POR2X1_90/Y 0.02fF
C43374 INPUT_3 PAND2X1_28/CTRL2 0.05fF
C43375 POR2X1_260/B POR2X1_788/B 0.03fF
C43376 PAND2X1_217/B PAND2X1_473/Y 0.05fF
C43377 POR2X1_846/Y POR2X1_754/O 0.01fF
C43378 POR2X1_60/A PAND2X1_468/a_16_344# 0.01fF
C43379 PAND2X1_104/a_56_28# PAND2X1_8/Y 0.00fF
C43380 PAND2X1_72/A POR2X1_728/A 0.03fF
C43381 POR2X1_308/CTRL POR2X1_830/A 0.00fF
C43382 PAND2X1_674/CTRL POR2X1_590/A 0.01fF
C43383 POR2X1_814/B POR2X1_608/O 0.02fF
C43384 POR2X1_445/CTRL POR2X1_750/B 0.12fF
C43385 PAND2X1_73/Y PAND2X1_79/O 0.20fF
C43386 POR2X1_594/Y POR2X1_594/O 0.01fF
C43387 POR2X1_296/B PAND2X1_144/O 0.07fF
C43388 POR2X1_43/B POR2X1_586/Y 0.14fF
C43389 POR2X1_555/B POR2X1_35/Y 0.02fF
C43390 POR2X1_413/A POR2X1_607/A 0.52fF
C43391 POR2X1_482/Y POR2X1_55/Y 0.08fF
C43392 POR2X1_54/Y POR2X1_249/Y 0.02fF
C43393 PAND2X1_48/B POR2X1_477/B 0.06fF
C43394 POR2X1_66/A POR2X1_532/A 0.20fF
C43395 PAND2X1_572/a_76_28# PAND2X1_267/Y 0.03fF
C43396 PAND2X1_572/O PAND2X1_576/B 0.02fF
C43397 PAND2X1_84/O POR2X1_497/Y 0.09fF
C43398 PAND2X1_713/B VDD 0.18fF
C43399 POR2X1_814/A POR2X1_383/O 0.02fF
C43400 PAND2X1_394/CTRL POR2X1_35/Y 0.01fF
C43401 PAND2X1_93/B POR2X1_510/Y 0.03fF
C43402 POR2X1_83/B PAND2X1_566/Y 0.02fF
C43403 POR2X1_104/CTRL2 D_INPUT_1 0.01fF
C43404 POR2X1_376/B POR2X1_817/A 0.86fF
C43405 POR2X1_559/Y PAND2X1_20/A 0.04fF
C43406 POR2X1_259/A POR2X1_785/A 0.03fF
C43407 POR2X1_490/Y PAND2X1_717/Y 0.03fF
C43408 POR2X1_96/A POR2X1_826/O 0.01fF
C43409 POR2X1_96/A POR2X1_5/Y 0.86fF
C43410 PAND2X1_6/Y PAND2X1_58/A 0.71fF
C43411 POR2X1_302/B POR2X1_740/Y 0.08fF
C43412 POR2X1_278/Y PAND2X1_659/CTRL2 0.02fF
C43413 PAND2X1_93/B PAND2X1_312/a_76_28# 0.01fF
C43414 PAND2X1_192/CTRL PAND2X1_191/Y 0.01fF
C43415 POR2X1_164/O POR2X1_83/B 0.01fF
C43416 POR2X1_68/A POR2X1_467/Y 0.03fF
C43417 POR2X1_48/A POR2X1_245/Y 0.03fF
C43418 POR2X1_133/O POR2X1_236/Y 0.11fF
C43419 PAND2X1_695/O PAND2X1_57/B 0.17fF
C43420 PAND2X1_473/Y VDD 0.17fF
C43421 POR2X1_784/O POR2X1_296/B 0.04fF
C43422 PAND2X1_592/O PAND2X1_473/B 0.05fF
C43423 POR2X1_523/Y POR2X1_750/A 0.02fF
C43424 POR2X1_330/Y POR2X1_35/Y 0.03fF
C43425 PAND2X1_208/m4_208_n4# PAND2X1_198/m4_208_n4# 0.05fF
C43426 POR2X1_29/Y POR2X1_159/CTRL2 0.01fF
C43427 POR2X1_406/CTRL POR2X1_5/Y 0.01fF
C43428 POR2X1_614/A POR2X1_450/B 0.82fF
C43429 POR2X1_141/O POR2X1_139/Y 0.00fF
C43430 POR2X1_124/B POR2X1_650/a_16_28# 0.01fF
C43431 POR2X1_96/A PAND2X1_549/CTRL2 0.00fF
C43432 POR2X1_8/Y PAND2X1_340/B 0.03fF
C43433 PAND2X1_272/O POR2X1_228/Y 0.14fF
C43434 POR2X1_43/B POR2X1_423/Y 0.03fF
C43435 POR2X1_54/Y POR2X1_394/A 0.34fF
C43436 PAND2X1_493/O POR2X1_411/B 0.02fF
C43437 POR2X1_387/a_16_28# POR2X1_386/Y 0.02fF
C43438 PAND2X1_93/B POR2X1_276/Y 0.03fF
C43439 POR2X1_106/Y POR2X1_55/Y 0.03fF
C43440 POR2X1_65/A POR2X1_591/O 0.01fF
C43441 POR2X1_376/B POR2X1_42/Y 0.04fF
C43442 POR2X1_478/CTRL POR2X1_444/Y 0.03fF
C43443 PAND2X1_357/Y PAND2X1_349/B 0.03fF
C43444 POR2X1_405/Y VDD 0.06fF
C43445 POR2X1_15/CTRL POR2X1_14/Y 0.01fF
C43446 PAND2X1_632/B POR2X1_23/Y 0.00fF
C43447 PAND2X1_623/O POR2X1_408/Y 0.04fF
C43448 POR2X1_41/B PAND2X1_715/O 0.07fF
C43449 PAND2X1_58/A POR2X1_791/A 0.60fF
C43450 POR2X1_12/CTRL POR2X1_587/Y 0.00fF
C43451 POR2X1_784/A VDD 0.43fF
C43452 PAND2X1_803/A POR2X1_238/Y 0.06fF
C43453 PAND2X1_57/CTRL POR2X1_404/Y 0.03fF
C43454 POR2X1_83/B POR2X1_245/O 0.04fF
C43455 POR2X1_102/Y POR2X1_757/CTRL 0.01fF
C43456 POR2X1_257/A PAND2X1_345/Y 0.03fF
C43457 PAND2X1_733/A POR2X1_73/Y 0.07fF
C43458 PAND2X1_478/CTRL2 POR2X1_236/Y 0.01fF
C43459 PAND2X1_654/A PAND2X1_404/Y 0.00fF
C43460 POR2X1_840/B POR2X1_141/Y 0.05fF
C43461 PAND2X1_57/B POR2X1_247/CTRL2 0.02fF
C43462 PAND2X1_435/CTRL POR2X1_293/Y 0.00fF
C43463 POR2X1_121/B PAND2X1_305/O 0.01fF
C43464 POR2X1_38/Y POR2X1_40/Y 0.96fF
C43465 POR2X1_78/B POR2X1_563/Y 0.01fF
C43466 PAND2X1_56/Y POR2X1_480/A 0.07fF
C43467 D_INPUT_0 PAND2X1_514/O 0.02fF
C43468 POR2X1_669/B PAND2X1_569/B 0.07fF
C43469 PAND2X1_57/B POR2X1_783/B 0.02fF
C43470 PAND2X1_736/A VDD 0.11fF
C43471 PAND2X1_281/CTRL2 POR2X1_862/A 0.06fF
C43472 POR2X1_453/CTRL PAND2X1_60/B 0.03fF
C43473 PAND2X1_687/A POR2X1_60/A 0.04fF
C43474 POR2X1_335/CTRL POR2X1_741/Y 0.00fF
C43475 POR2X1_335/O POR2X1_740/Y 0.05fF
C43476 VDD POR2X1_732/B 2.36fF
C43477 PAND2X1_48/O POR2X1_294/B 0.03fF
C43478 POR2X1_14/Y PAND2X1_63/B 0.03fF
C43479 PAND2X1_23/Y POR2X1_244/B 0.01fF
C43480 POR2X1_539/A POR2X1_457/CTRL2 0.08fF
C43481 PAND2X1_411/CTRL POR2X1_461/B 0.00fF
C43482 PAND2X1_63/Y POR2X1_650/A 0.07fF
C43483 POR2X1_315/Y POR2X1_83/B 0.07fF
C43484 POR2X1_41/B POR2X1_293/Y 1.67fF
C43485 POR2X1_496/Y PAND2X1_508/CTRL 0.05fF
C43486 POR2X1_567/B POR2X1_544/B 0.03fF
C43487 POR2X1_347/a_16_28# POR2X1_402/A 0.01fF
C43488 PAND2X1_263/CTRL D_INPUT_1 0.06fF
C43489 POR2X1_697/CTRL2 PAND2X1_565/A 0.00fF
C43490 POR2X1_52/A POR2X1_71/Y 0.57fF
C43491 PAND2X1_207/a_16_344# POR2X1_394/A 0.02fF
C43492 PAND2X1_835/O VDD 0.00fF
C43493 PAND2X1_31/CTRL2 PAND2X1_18/B 0.04fF
C43494 POR2X1_26/CTRL POR2X1_32/A 0.01fF
C43495 POR2X1_78/A POR2X1_276/Y 0.11fF
C43496 POR2X1_823/CTRL2 VDD 0.00fF
C43497 PAND2X1_6/Y POR2X1_457/B 0.01fF
C43498 POR2X1_307/a_16_28# POR2X1_307/A 0.03fF
C43499 POR2X1_296/B POR2X1_456/B 0.03fF
C43500 PAND2X1_342/O POR2X1_5/Y 0.04fF
C43501 PAND2X1_94/A PAND2X1_531/O 0.03fF
C43502 PAND2X1_622/CTRL POR2X1_619/Y 0.01fF
C43503 POR2X1_853/O POR2X1_785/A 0.16fF
C43504 PAND2X1_65/B POR2X1_577/CTRL 0.03fF
C43505 POR2X1_257/A POR2X1_524/CTRL2 0.00fF
C43506 POR2X1_567/A POR2X1_445/A 6.17fF
C43507 POR2X1_417/Y POR2X1_283/A -0.01fF
C43508 POR2X1_291/a_16_28# POR2X1_32/A 0.01fF
C43509 PAND2X1_393/CTRL PAND2X1_41/B 0.01fF
C43510 POR2X1_231/B POR2X1_785/A 0.02fF
C43511 PAND2X1_90/Y POR2X1_758/CTRL 0.03fF
C43512 POR2X1_52/A POR2X1_42/Y 0.54fF
C43513 PAND2X1_6/Y POR2X1_435/Y 0.07fF
C43514 POR2X1_113/Y POR2X1_650/A 0.00fF
C43515 POR2X1_48/A POR2X1_183/O 0.02fF
C43516 PAND2X1_862/B POR2X1_56/Y 0.03fF
C43517 D_INPUT_0 POR2X1_5/CTRL2 -0.00fF
C43518 POR2X1_376/B PAND2X1_99/Y 0.05fF
C43519 PAND2X1_106/CTRL POR2X1_105/Y 0.01fF
C43520 POR2X1_806/O POR2X1_675/Y 0.02fF
C43521 PAND2X1_74/CTRL POR2X1_456/B 0.01fF
C43522 POR2X1_139/A POR2X1_130/A 0.02fF
C43523 POR2X1_346/B POR2X1_630/A 0.02fF
C43524 POR2X1_335/A PAND2X1_498/CTRL 0.01fF
C43525 PAND2X1_241/Y POR2X1_511/Y 0.03fF
C43526 PAND2X1_472/A POR2X1_669/CTRL2 0.01fF
C43527 POR2X1_68/B INPUT_0 0.44fF
C43528 POR2X1_65/A POR2X1_73/CTRL 0.01fF
C43529 POR2X1_538/a_16_28# POR2X1_566/A 0.02fF
C43530 POR2X1_20/B POR2X1_387/O 0.01fF
C43531 INPUT_1 POR2X1_40/Y 0.18fF
C43532 POR2X1_7/A POR2X1_5/Y 1.23fF
C43533 PAND2X1_298/CTRL POR2X1_750/B 0.03fF
C43534 POR2X1_300/CTRL2 POR2X1_184/Y 0.00fF
C43535 POR2X1_333/A POR2X1_333/Y 0.00fF
C43536 PAND2X1_716/CTRL2 PAND2X1_197/Y 0.00fF
C43537 PAND2X1_90/Y PAND2X1_305/a_16_344# 0.02fF
C43538 POR2X1_343/Y POR2X1_341/A 0.10fF
C43539 POR2X1_192/Y POR2X1_341/Y 0.05fF
C43540 POR2X1_405/Y PAND2X1_32/B 0.03fF
C43541 INPUT_1 POR2X1_35/B 0.03fF
C43542 PAND2X1_730/a_16_344# POR2X1_42/Y 0.01fF
C43543 PAND2X1_563/A PAND2X1_554/O 0.02fF
C43544 PAND2X1_640/O POR2X1_293/Y 0.08fF
C43545 POR2X1_383/A POR2X1_480/A 0.09fF
C43546 PAND2X1_575/a_16_344# INPUT_0 0.02fF
C43547 POR2X1_644/A POR2X1_513/B 0.42fF
C43548 POR2X1_763/Y PAND2X1_324/CTRL 0.01fF
C43549 POR2X1_784/A PAND2X1_32/B 0.03fF
C43550 POR2X1_96/A PAND2X1_739/B 0.03fF
C43551 POR2X1_804/A PAND2X1_369/CTRL 0.01fF
C43552 PAND2X1_462/B POR2X1_232/Y 0.03fF
C43553 PAND2X1_55/Y POR2X1_786/Y 0.05fF
C43554 PAND2X1_862/Y POR2X1_102/Y 0.01fF
C43555 PAND2X1_753/a_16_344# PAND2X1_752/Y 0.05fF
C43556 POR2X1_49/Y PAND2X1_620/CTRL 0.00fF
C43557 PAND2X1_63/Y POR2X1_294/B 0.10fF
C43558 POR2X1_40/Y POR2X1_153/Y 0.28fF
C43559 POR2X1_765/Y VDD 0.00fF
C43560 POR2X1_532/A POR2X1_802/B 0.41fF
C43561 POR2X1_709/A PAND2X1_52/B 0.03fF
C43562 POR2X1_650/A POR2X1_260/A 0.03fF
C43563 POR2X1_732/a_56_344# POR2X1_732/B 0.03fF
C43564 POR2X1_384/A POR2X1_40/Y 0.07fF
C43565 POR2X1_325/CTRL POR2X1_502/A 0.01fF
C43566 POR2X1_785/A PAND2X1_88/Y 0.03fF
C43567 PAND2X1_95/B POR2X1_460/A 0.01fF
C43568 POR2X1_41/B POR2X1_408/Y 0.10fF
C43569 POR2X1_186/a_16_28# POR2X1_750/B 0.02fF
C43570 POR2X1_115/O POR2X1_366/A 0.02fF
C43571 POR2X1_16/A POR2X1_236/Y 1.84fF
C43572 POR2X1_198/CTRL POR2X1_532/A 0.01fF
C43573 PAND2X1_283/CTRL2 PAND2X1_96/B 0.09fF
C43574 POR2X1_443/A POR2X1_568/A 0.01fF
C43575 POR2X1_351/Y POR2X1_350/a_16_28# 0.01fF
C43576 PAND2X1_41/B POR2X1_564/B 0.01fF
C43577 PAND2X1_65/B POR2X1_244/Y 0.03fF
C43578 PAND2X1_220/Y PAND2X1_343/a_76_28# 0.03fF
C43579 POR2X1_78/B POR2X1_675/Y 0.03fF
C43580 POR2X1_402/A PAND2X1_69/CTRL 0.01fF
C43581 POR2X1_853/A POR2X1_577/O 0.01fF
C43582 POR2X1_222/Y POR2X1_532/A 0.06fF
C43583 POR2X1_89/a_16_28# POR2X1_77/Y 0.05fF
C43584 POR2X1_423/Y POR2X1_183/CTRL 0.01fF
C43585 POR2X1_113/Y POR2X1_294/B 0.03fF
C43586 D_INPUT_0 POR2X1_39/B 0.09fF
C43587 POR2X1_78/CTRL2 PAND2X1_96/B 0.01fF
C43588 PAND2X1_534/CTRL POR2X1_294/B 0.06fF
C43589 POR2X1_570/B POR2X1_562/B 0.00fF
C43590 POR2X1_388/CTRL PAND2X1_69/A 0.01fF
C43591 PAND2X1_848/B POR2X1_38/Y 0.03fF
C43592 PAND2X1_6/Y PAND2X1_96/B 0.14fF
C43593 PAND2X1_319/B POR2X1_43/B 0.07fF
C43594 POR2X1_579/Y POR2X1_854/B 0.03fF
C43595 POR2X1_804/A POR2X1_702/A 0.15fF
C43596 POR2X1_37/Y POR2X1_77/Y 0.20fF
C43597 POR2X1_274/A POR2X1_717/B 0.01fF
C43598 PAND2X1_319/B POR2X1_312/O 0.05fF
C43599 PAND2X1_90/A POR2X1_383/A 0.16fF
C43600 PAND2X1_349/A POR2X1_55/Y 0.02fF
C43601 POR2X1_754/A POR2X1_754/CTRL2 0.01fF
C43602 POR2X1_84/a_16_28# POR2X1_532/A 0.02fF
C43603 PAND2X1_537/CTRL2 PAND2X1_364/B 0.03fF
C43604 PAND2X1_63/B POR2X1_55/Y 0.03fF
C43605 PAND2X1_705/O POR2X1_526/Y 0.00fF
C43606 POR2X1_85/Y POR2X1_37/Y 0.05fF
C43607 POR2X1_652/Y POR2X1_799/O 0.02fF
C43608 INPUT_1 POR2X1_586/CTRL 0.01fF
C43609 POR2X1_617/Y POR2X1_847/B 0.02fF
C43610 POR2X1_179/O POR2X1_387/Y 0.02fF
C43611 PAND2X1_48/B POR2X1_101/Y 0.13fF
C43612 POR2X1_334/B POR2X1_569/A 0.10fF
C43613 PAND2X1_148/CTRL2 PAND2X1_148/Y 0.02fF
C43614 POR2X1_559/B POR2X1_264/Y 0.01fF
C43615 POR2X1_192/Y POR2X1_731/A 0.03fF
C43616 PAND2X1_72/a_16_344# POR2X1_532/A 0.01fF
C43617 PAND2X1_80/CTRL2 PAND2X1_71/Y 0.01fF
C43618 PAND2X1_659/B POR2X1_153/Y 0.03fF
C43619 POR2X1_545/A POR2X1_854/B 0.05fF
C43620 POR2X1_191/B VDD 0.02fF
C43621 POR2X1_687/Y POR2X1_614/A 0.69fF
C43622 POR2X1_283/A POR2X1_184/Y 0.03fF
C43623 POR2X1_252/Y POR2X1_376/B 0.03fF
C43624 POR2X1_383/A PAND2X1_494/O 0.01fF
C43625 PAND2X1_63/Y PAND2X1_111/B 0.03fF
C43626 POR2X1_619/A POR2X1_751/CTRL 0.04fF
C43627 PAND2X1_65/B POR2X1_191/Y 0.05fF
C43628 POR2X1_294/B POR2X1_260/A 2.22fF
C43629 PAND2X1_493/CTRL PAND2X1_480/B 0.02fF
C43630 PAND2X1_56/Y POR2X1_787/CTRL 0.00fF
C43631 POR2X1_156/a_16_28# POR2X1_750/B 0.02fF
C43632 PAND2X1_651/Y POR2X1_283/A 0.03fF
C43633 POR2X1_208/A PAND2X1_69/A 0.03fF
C43634 PAND2X1_683/O POR2X1_78/B 0.01fF
C43635 POR2X1_96/A PAND2X1_779/CTRL2 0.00fF
C43636 POR2X1_97/B VDD 0.15fF
C43637 POR2X1_220/Y POR2X1_210/A 0.00fF
C43638 POR2X1_207/A PAND2X1_41/Y 0.00fF
C43639 VDD POR2X1_7/Y 0.60fF
C43640 POR2X1_711/CTRL POR2X1_713/B 0.01fF
C43641 PAND2X1_477/A POR2X1_43/B 0.01fF
C43642 POR2X1_231/B POR2X1_186/B 0.01fF
C43643 POR2X1_334/Y PAND2X1_89/O 0.08fF
C43644 PAND2X1_58/A PAND2X1_52/B 0.08fF
C43645 POR2X1_404/Y PAND2X1_399/O 0.01fF
C43646 POR2X1_390/B POR2X1_513/Y 0.03fF
C43647 PAND2X1_738/B POR2X1_39/B 0.04fF
C43648 PAND2X1_175/B POR2X1_91/Y 0.03fF
C43649 POR2X1_287/B POR2X1_343/O 0.01fF
C43650 PAND2X1_177/CTRL POR2X1_180/A 0.01fF
C43651 POR2X1_13/A PAND2X1_141/O 0.04fF
C43652 POR2X1_16/A POR2X1_232/Y 0.00fF
C43653 PAND2X1_371/CTRL POR2X1_773/A 0.03fF
C43654 PAND2X1_60/B POR2X1_758/a_16_28# 0.02fF
C43655 PAND2X1_90/A PAND2X1_71/Y 0.03fF
C43656 POR2X1_119/Y PAND2X1_793/Y 0.05fF
C43657 PAND2X1_473/CTRL2 PAND2X1_216/B 0.00fF
C43658 POR2X1_101/a_16_28# PAND2X1_69/A 0.00fF
C43659 POR2X1_670/O POR2X1_77/Y 0.09fF
C43660 POR2X1_90/Y POR2X1_766/a_16_28# 0.01fF
C43661 PAND2X1_48/B POR2X1_722/O 0.01fF
C43662 POR2X1_227/B POR2X1_227/A 0.03fF
C43663 POR2X1_548/B PAND2X1_143/CTRL2 0.03fF
C43664 POR2X1_283/A POR2X1_503/Y 0.32fF
C43665 POR2X1_440/Y POR2X1_854/B 0.03fF
C43666 POR2X1_327/Y D_INPUT_1 0.03fF
C43667 POR2X1_590/CTRL POR2X1_796/A 0.02fF
C43668 POR2X1_809/A POR2X1_810/a_56_344# 0.00fF
C43669 PAND2X1_42/a_76_28# POR2X1_267/A 0.04fF
C43670 PAND2X1_437/O POR2X1_590/A 0.01fF
C43671 POR2X1_822/Y POR2X1_394/A 0.06fF
C43672 PAND2X1_48/B PAND2X1_696/CTRL2 0.03fF
C43673 PAND2X1_111/B POR2X1_260/A 0.03fF
C43674 POR2X1_13/A POR2X1_372/CTRL2 0.00fF
C43675 PAND2X1_48/B POR2X1_542/CTRL2 0.10fF
C43676 POR2X1_178/a_16_28# PAND2X1_348/A 0.08fF
C43677 PAND2X1_60/B POR2X1_353/A 0.03fF
C43678 D_INPUT_3 POR2X1_4/O 0.01fF
C43679 PAND2X1_88/Y POR2X1_186/B 0.03fF
C43680 POR2X1_614/A POR2X1_845/A 0.01fF
C43681 PAND2X1_60/B POR2X1_332/O 0.00fF
C43682 POR2X1_856/B POR2X1_814/A 0.10fF
C43683 POR2X1_303/CTRL2 POR2X1_513/Y 0.03fF
C43684 PAND2X1_511/O PAND2X1_56/A 0.02fF
C43685 PAND2X1_787/A POR2X1_394/A 0.03fF
C43686 POR2X1_773/A PAND2X1_69/A 0.07fF
C43687 POR2X1_140/B POR2X1_540/Y 0.32fF
C43688 POR2X1_568/Y POR2X1_545/CTRL 0.01fF
C43689 PAND2X1_211/O POR2X1_20/B 0.15fF
C43690 POR2X1_228/a_16_28# POR2X1_631/B 0.01fF
C43691 POR2X1_208/A PAND2X1_824/B 0.03fF
C43692 POR2X1_85/a_16_28# PAND2X1_35/Y 0.02fF
C43693 PAND2X1_194/O POR2X1_16/Y -0.00fF
C43694 PAND2X1_501/O PAND2X1_862/B 0.02fF
C43695 POR2X1_785/A POR2X1_568/B 0.03fF
C43696 POR2X1_624/Y POR2X1_341/A 0.03fF
C43697 PAND2X1_290/CTRL POR2X1_334/B 0.02fF
C43698 POR2X1_322/Y POR2X1_373/Y 0.71fF
C43699 POR2X1_609/Y PAND2X1_608/O 0.00fF
C43700 POR2X1_119/Y PAND2X1_711/A 0.06fF
C43701 POR2X1_762/a_56_344# D_INPUT_6 0.00fF
C43702 POR2X1_669/B POR2X1_667/O 0.10fF
C43703 PAND2X1_189/CTRL2 POR2X1_854/B 0.08fF
C43704 POR2X1_293/Y POR2X1_77/Y 0.10fF
C43705 PAND2X1_858/O POR2X1_91/Y 0.06fF
C43706 POR2X1_85/Y POR2X1_293/Y 0.03fF
C43707 POR2X1_66/Y PAND2X1_67/O 0.07fF
C43708 POR2X1_832/A PAND2X1_48/A 0.07fF
C43709 POR2X1_224/Y POR2X1_77/Y 0.11fF
C43710 PAND2X1_160/CTRL POR2X1_394/A 0.01fF
C43711 POR2X1_553/O POR2X1_569/A 0.05fF
C43712 POR2X1_281/Y PAND2X1_805/A 0.03fF
C43713 POR2X1_329/A PAND2X1_561/Y 0.01fF
C43714 POR2X1_670/Y POR2X1_416/B 0.00fF
C43715 POR2X1_357/O POR2X1_568/Y 0.04fF
C43716 POR2X1_68/A POR2X1_555/CTRL2 0.01fF
C43717 POR2X1_203/a_16_28# PAND2X1_48/A 0.02fF
C43718 POR2X1_270/a_16_28# POR2X1_567/A -0.00fF
C43719 PAND2X1_680/CTRL2 POR2X1_162/Y 0.01fF
C43720 PAND2X1_6/Y POR2X1_342/B 0.02fF
C43721 POR2X1_86/O POR2X1_73/Y 0.01fF
C43722 POR2X1_16/A PAND2X1_803/O 0.03fF
C43723 PAND2X1_433/CTRL PAND2X1_72/A 0.01fF
C43724 POR2X1_733/A PAND2X1_72/A 1.43fF
C43725 POR2X1_20/B PAND2X1_722/O 0.04fF
C43726 POR2X1_647/B POR2X1_286/CTRL2 0.01fF
C43727 POR2X1_334/B PAND2X1_72/A 0.03fF
C43728 PAND2X1_65/B PAND2X1_224/CTRL 0.01fF
C43729 POR2X1_20/B POR2X1_29/A 0.06fF
C43730 POR2X1_411/B POR2X1_67/A 0.07fF
C43731 POR2X1_41/B PAND2X1_242/Y 0.10fF
C43732 POR2X1_74/a_16_28# POR2X1_271/A 0.02fF
C43733 POR2X1_416/B PAND2X1_565/A 0.03fF
C43734 POR2X1_537/CTRL2 POR2X1_537/Y 0.01fF
C43735 PAND2X1_47/O PAND2X1_11/Y 0.04fF
C43736 POR2X1_782/A PAND2X1_52/B 0.03fF
C43737 POR2X1_168/O POR2X1_566/B 0.35fF
C43738 POR2X1_383/A PAND2X1_304/O 0.18fF
C43739 POR2X1_104/CTRL2 INPUT_3 0.05fF
C43740 PAND2X1_634/O POR2X1_607/A 0.00fF
C43741 POR2X1_411/B POR2X1_226/O 0.01fF
C43742 POR2X1_54/Y POR2X1_669/B 0.16fF
C43743 POR2X1_329/A PAND2X1_733/m4_208_n4# 0.08fF
C43744 POR2X1_84/A POR2X1_240/m4_208_n4# 0.09fF
C43745 POR2X1_394/A POR2X1_701/CTRL2 0.01fF
C43746 POR2X1_567/A POR2X1_260/A 0.05fF
C43747 POR2X1_48/A PAND2X1_590/CTRL 0.01fF
C43748 POR2X1_9/Y POR2X1_88/Y 0.10fF
C43749 POR2X1_76/B POR2X1_575/B 0.00fF
C43750 POR2X1_846/Y POR2X1_615/CTRL 0.00fF
C43751 PAND2X1_96/B PAND2X1_52/B 0.06fF
C43752 POR2X1_36/B POR2X1_416/B 0.54fF
C43753 PAND2X1_358/O PAND2X1_656/A 0.02fF
C43754 PAND2X1_35/A PAND2X1_34/O 0.03fF
C43755 PAND2X1_651/CTRL PAND2X1_639/Y 0.12fF
C43756 POR2X1_648/Y POR2X1_480/A 0.07fF
C43757 POR2X1_78/A PAND2X1_609/CTRL2 0.01fF
C43758 POR2X1_566/B POR2X1_567/CTRL2 0.02fF
C43759 PAND2X1_644/O POR2X1_236/Y 0.01fF
C43760 POR2X1_760/A POR2X1_5/Y 0.12fF
C43761 POR2X1_48/A D_INPUT_0 0.10fF
C43762 POR2X1_329/A PAND2X1_362/B 0.01fF
C43763 POR2X1_394/A POR2X1_4/Y 0.08fF
C43764 POR2X1_748/A POR2X1_628/Y 0.18fF
C43765 PAND2X1_86/CTRL2 POR2X1_243/Y -0.02fF
C43766 POR2X1_373/Y POR2X1_373/O 0.03fF
C43767 PAND2X1_199/CTRL PAND2X1_123/Y 0.01fF
C43768 POR2X1_257/A PAND2X1_217/B 0.07fF
C43769 POR2X1_852/B POR2X1_776/A 0.46fF
C43770 POR2X1_624/Y POR2X1_500/A 0.01fF
C43771 POR2X1_78/A POR2X1_807/O 0.02fF
C43772 POR2X1_287/B PAND2X1_39/B 0.02fF
C43773 POR2X1_257/A PAND2X1_392/B 0.02fF
C43774 PAND2X1_207/CTRL2 POR2X1_72/B 0.02fF
C43775 PAND2X1_206/B POR2X1_7/B 0.07fF
C43776 PAND2X1_246/CTRL2 POR2X1_404/Y 0.10fF
C43777 POR2X1_650/A POR2X1_473/O 0.01fF
C43778 PAND2X1_267/a_16_344# POR2X1_72/B 0.01fF
C43779 PAND2X1_628/O PAND2X1_88/Y 0.02fF
C43780 POR2X1_553/a_56_344# POR2X1_632/Y 0.00fF
C43781 POR2X1_14/Y POR2X1_32/A 0.03fF
C43782 PAND2X1_96/B PAND2X1_628/m4_208_n4# 0.15fF
C43783 POR2X1_257/A VDD 3.84fF
C43784 PAND2X1_406/CTRL POR2X1_362/B 0.01fF
C43785 PAND2X1_39/B PAND2X1_8/Y 0.18fF
C43786 POR2X1_376/B POR2X1_699/CTRL 0.01fF
C43787 POR2X1_54/Y PAND2X1_293/CTRL 0.03fF
C43788 POR2X1_262/Y PAND2X1_364/B 0.07fF
C43789 POR2X1_866/A PAND2X1_65/B 0.03fF
C43790 POR2X1_48/A PAND2X1_738/B 0.05fF
C43791 POR2X1_856/B POR2X1_852/B 0.07fF
C43792 POR2X1_60/A PAND2X1_200/CTRL2 0.01fF
C43793 PAND2X1_439/CTRL POR2X1_90/Y 0.01fF
C43794 PAND2X1_66/a_56_28# POR2X1_5/Y 0.00fF
C43795 POR2X1_290/O POR2X1_37/Y 0.02fF
C43796 POR2X1_566/A POR2X1_454/CTRL 0.01fF
C43797 POR2X1_102/Y POR2X1_609/CTRL2 0.01fF
C43798 POR2X1_68/A POR2X1_623/Y 0.03fF
C43799 POR2X1_612/B VDD 0.05fF
C43800 PAND2X1_621/Y POR2X1_415/A 0.02fF
C43801 POR2X1_260/B POR2X1_410/O 0.02fF
C43802 POR2X1_202/A POR2X1_404/B 0.02fF
C43803 POR2X1_417/Y POR2X1_14/Y 0.18fF
C43804 PAND2X1_222/a_76_28# INPUT_0 0.01fF
C43805 POR2X1_14/Y POR2X1_419/Y 0.03fF
C43806 POR2X1_436/B POR2X1_436/a_76_344# 0.01fF
C43807 D_INPUT_5 POR2X1_638/CTRL2 0.00fF
C43808 POR2X1_754/Y POR2X1_625/CTRL 0.00fF
C43809 PAND2X1_453/A POR2X1_419/Y 0.06fF
C43810 POR2X1_49/Y PAND2X1_848/O 0.02fF
C43811 POR2X1_485/Y PAND2X1_705/O 0.04fF
C43812 PAND2X1_286/B PAND2X1_286/a_16_344# 0.03fF
C43813 PAND2X1_203/O PAND2X1_575/A 0.01fF
C43814 POR2X1_462/a_76_344# PAND2X1_69/A 0.01fF
C43815 PAND2X1_658/a_16_344# POR2X1_60/A 0.02fF
C43816 POR2X1_23/Y POR2X1_697/m4_208_n4# 0.12fF
C43817 POR2X1_492/O POR2X1_60/A 0.02fF
C43818 POR2X1_812/A POR2X1_801/CTRL 0.01fF
C43819 PAND2X1_214/A POR2X1_40/Y 0.12fF
C43820 POR2X1_52/A POR2X1_89/CTRL 0.01fF
C43821 POR2X1_466/A VDD 3.58fF
C43822 PAND2X1_78/O PAND2X1_354/A 0.02fF
C43823 POR2X1_119/Y PAND2X1_862/O 0.03fF
C43824 PAND2X1_263/CTRL POR2X1_78/A 0.01fF
C43825 POR2X1_411/B PAND2X1_642/B 0.02fF
C43826 POR2X1_620/O PAND2X1_9/Y 0.01fF
C43827 PAND2X1_20/A POR2X1_287/B 0.03fF
C43828 POR2X1_253/CTRL PAND2X1_6/A 0.05fF
C43829 POR2X1_48/O POR2X1_32/A 0.02fF
C43830 POR2X1_66/B PAND2X1_16/O 0.03fF
C43831 POR2X1_49/Y POR2X1_820/O 0.18fF
C43832 POR2X1_834/CTRL VDD 0.00fF
C43833 POR2X1_329/A PAND2X1_717/Y 0.03fF
C43834 POR2X1_260/B POR2X1_715/a_76_344# 0.01fF
C43835 POR2X1_322/CTRL2 POR2X1_23/Y 0.01fF
C43836 POR2X1_8/Y POR2X1_9/Y 0.27fF
C43837 POR2X1_473/CTRL POR2X1_391/Y 0.06fF
C43838 POR2X1_49/Y PAND2X1_217/B 0.05fF
C43839 PAND2X1_796/B POR2X1_90/Y 0.02fF
C43840 POR2X1_641/a_16_28# POR2X1_267/B 0.03fF
C43841 PAND2X1_454/B POR2X1_90/Y 0.03fF
C43842 POR2X1_556/A POR2X1_318/A 0.07fF
C43843 PAND2X1_57/B POR2X1_296/B 3.77fF
C43844 POR2X1_439/Y PAND2X1_41/B 0.01fF
C43845 POR2X1_694/a_16_28# POR2X1_257/A 0.01fF
C43846 PAND2X1_250/O POR2X1_287/B 0.01fF
C43847 POR2X1_814/B POR2X1_287/B 0.03fF
C43848 POR2X1_141/Y POR2X1_217/CTRL 0.00fF
C43849 POR2X1_673/A POR2X1_673/O 0.18fF
C43850 POR2X1_199/O POR2X1_590/A 0.18fF
C43851 POR2X1_413/A D_INPUT_0 0.01fF
C43852 PAND2X1_195/a_56_28# POR2X1_236/Y 0.00fF
C43853 POR2X1_814/A POR2X1_244/Y 0.12fF
C43854 POR2X1_516/CTRL POR2X1_48/A 0.01fF
C43855 PAND2X1_73/Y POR2X1_193/A 0.03fF
C43856 PAND2X1_73/Y POR2X1_579/Y 0.01fF
C43857 POR2X1_674/Y POR2X1_331/A 0.02fF
C43858 PAND2X1_862/B PAND2X1_575/B 0.03fF
C43859 PAND2X1_275/O D_INPUT_0 0.03fF
C43860 POR2X1_148/O POR2X1_532/A 0.01fF
C43861 PAND2X1_20/A PAND2X1_89/CTRL 0.01fF
C43862 POR2X1_41/B POR2X1_60/A 0.67fF
C43863 POR2X1_32/A POR2X1_55/Y 0.71fF
C43864 POR2X1_413/A PAND2X1_656/O 0.02fF
C43865 POR2X1_52/A POR2X1_226/O 0.02fF
C43866 POR2X1_250/CTRL2 POR2X1_250/A 0.00fF
C43867 INPUT_7 POR2X1_2/CTRL2 0.03fF
C43868 POR2X1_49/Y VDD 1.69fF
C43869 POR2X1_23/Y POR2X1_90/Y 0.05fF
C43870 POR2X1_39/B POR2X1_90/O 0.01fF
C43871 PAND2X1_20/A PAND2X1_226/O 0.04fF
C43872 PAND2X1_630/O POR2X1_496/Y 0.09fF
C43873 PAND2X1_807/B POR2X1_42/Y 0.30fF
C43874 POR2X1_407/A POR2X1_843/CTRL2 0.10fF
C43875 POR2X1_528/a_16_28# POR2X1_48/A 0.00fF
C43876 PAND2X1_80/a_16_344# PAND2X1_41/B 0.01fF
C43877 POR2X1_65/A POR2X1_481/A 0.03fF
C43878 POR2X1_814/B PAND2X1_8/Y 0.21fF
C43879 POR2X1_614/a_16_28# PAND2X1_69/A 0.03fF
C43880 POR2X1_192/Y PAND2X1_41/B 0.24fF
C43881 POR2X1_254/Y PAND2X1_13/CTRL 0.03fF
C43882 POR2X1_378/Y POR2X1_750/B 0.03fF
C43883 PAND2X1_340/CTRL2 INPUT_0 0.05fF
C43884 POR2X1_353/Y VDD 0.10fF
C43885 PAND2X1_581/Y VDD 0.13fF
C43886 POR2X1_753/Y POR2X1_790/A 0.08fF
C43887 PAND2X1_848/B PAND2X1_848/CTRL 0.01fF
C43888 POR2X1_257/A PAND2X1_467/O 0.17fF
C43889 PAND2X1_242/Y POR2X1_77/Y 0.01fF
C43890 PAND2X1_434/O POR2X1_172/Y 0.04fF
C43891 PAND2X1_621/CTRL POR2X1_415/A 0.06fF
C43892 POR2X1_614/A PAND2X1_73/Y 0.24fF
C43893 POR2X1_417/Y POR2X1_55/Y 0.18fF
C43894 POR2X1_419/Y POR2X1_55/Y 0.00fF
C43895 POR2X1_220/B POR2X1_532/A 0.03fF
C43896 POR2X1_590/A POR2X1_778/B 0.59fF
C43897 POR2X1_651/Y PAND2X1_56/A 0.03fF
C43898 PAND2X1_96/B POR2X1_288/CTRL 0.01fF
C43899 PAND2X1_6/A POR2X1_516/Y 0.04fF
C43900 PAND2X1_220/Y POR2X1_7/B 0.03fF
C43901 POR2X1_32/A PAND2X1_186/CTRL 0.01fF
C43902 PAND2X1_735/Y PAND2X1_499/Y 0.10fF
C43903 POR2X1_510/B POR2X1_567/B 0.91fF
C43904 PAND2X1_217/B PAND2X1_188/O 0.20fF
C43905 POR2X1_651/CTRL2 PAND2X1_90/Y 0.10fF
C43906 POR2X1_634/A POR2X1_391/Y 0.07fF
C43907 PAND2X1_651/Y POR2X1_14/Y 0.02fF
C43908 PAND2X1_73/Y POR2X1_38/B 0.16fF
C43909 POR2X1_62/Y PAND2X1_201/CTRL 0.01fF
C43910 PAND2X1_319/B POR2X1_298/Y 0.07fF
C43911 POR2X1_730/O POR2X1_330/Y 0.01fF
C43912 POR2X1_502/A PAND2X1_700/CTRL 0.07fF
C43913 POR2X1_322/O POR2X1_49/Y 0.01fF
C43914 POR2X1_814/A POR2X1_330/CTRL 0.06fF
C43915 POR2X1_66/B PAND2X1_385/m4_208_n4# 0.15fF
C43916 POR2X1_66/A PAND2X1_397/CTRL 0.01fF
C43917 POR2X1_60/A POR2X1_256/Y 0.01fF
C43918 POR2X1_355/B POR2X1_78/B 0.07fF
C43919 POR2X1_96/A PAND2X1_347/Y 0.03fF
C43920 PAND2X1_804/A PAND2X1_804/B 0.02fF
C43921 POR2X1_718/A POR2X1_294/B 0.07fF
C43922 POR2X1_243/Y INPUT_0 0.18fF
C43923 POR2X1_516/CTRL2 POR2X1_423/Y 0.01fF
C43924 POR2X1_341/A POR2X1_186/B 0.10fF
C43925 PAND2X1_11/Y D_INPUT_6 0.03fF
C43926 POR2X1_48/A POR2X1_108/Y 0.00fF
C43927 PAND2X1_454/CTRL POR2X1_511/Y 0.03fF
C43928 PAND2X1_219/B PAND2X1_219/O 0.00fF
C43929 POR2X1_66/B POR2X1_140/CTRL2 0.01fF
C43930 PAND2X1_553/B VDD 0.00fF
C43931 PAND2X1_371/O VDD 0.00fF
C43932 PAND2X1_833/CTRL2 PAND2X1_658/B 0.02fF
C43933 PAND2X1_29/O PAND2X1_41/B 0.03fF
C43934 POR2X1_13/A INPUT_4 0.03fF
C43935 POR2X1_65/A POR2X1_93/CTRL2 0.00fF
C43936 PAND2X1_715/CTRL PAND2X1_115/B 0.01fF
C43937 POR2X1_23/Y PAND2X1_732/A 0.03fF
C43938 PAND2X1_650/A D_INPUT_0 0.05fF
C43939 POR2X1_311/Y PAND2X1_222/B 0.10fF
C43940 POR2X1_52/A PAND2X1_455/Y 0.01fF
C43941 POR2X1_312/Y POR2X1_90/Y 0.33fF
C43942 POR2X1_590/A POR2X1_854/B 0.05fF
C43943 POR2X1_105/Y POR2X1_723/B 0.19fF
C43944 VDD PAND2X1_303/O 0.00fF
C43945 PAND2X1_824/B POR2X1_240/a_16_28# 0.02fF
C43946 PAND2X1_56/Y POR2X1_308/CTRL2 0.16fF
C43947 POR2X1_10/O POR2X1_48/A 0.01fF
C43948 POR2X1_777/B PAND2X1_150/CTRL2 0.11fF
C43949 PAND2X1_245/O PAND2X1_63/B 0.05fF
C43950 POR2X1_71/Y PAND2X1_862/B 0.03fF
C43951 PAND2X1_23/Y PAND2X1_58/O 0.00fF
C43952 PAND2X1_438/O PAND2X1_72/A 0.15fF
C43953 POR2X1_40/Y POR2X1_591/Y 0.03fF
C43954 PAND2X1_90/A INPUT_0 1.79fF
C43955 POR2X1_668/CTRL POR2X1_816/A 0.04fF
C43956 VDD PAND2X1_188/O -0.00fF
C43957 POR2X1_392/B PAND2X1_153/CTRL2 0.05fF
C43958 POR2X1_78/B POR2X1_538/CTRL 0.03fF
C43959 PAND2X1_852/a_16_344# POR2X1_122/Y 0.02fF
C43960 POR2X1_254/A PAND2X1_60/B 0.02fF
C43961 PAND2X1_794/B PAND2X1_473/B 0.08fF
C43962 PAND2X1_318/O POR2X1_96/A 0.02fF
C43963 POR2X1_327/Y PAND2X1_93/B 0.13fF
C43964 PAND2X1_57/B POR2X1_363/CTRL2 0.03fF
C43965 PAND2X1_264/CTRL2 POR2X1_83/B 0.01fF
C43966 POR2X1_447/B POR2X1_66/Y 0.06fF
C43967 POR2X1_273/a_16_28# POR2X1_153/Y 0.01fF
C43968 PAND2X1_206/CTRL2 PAND2X1_6/A 0.02fF
C43969 PAND2X1_35/Y POR2X1_55/Y 0.03fF
C43970 POR2X1_750/B PAND2X1_60/B 0.08fF
C43971 POR2X1_335/B POR2X1_543/A 0.13fF
C43972 POR2X1_706/CTRL INPUT_1 0.01fF
C43973 POR2X1_706/O PAND2X1_94/A 0.01fF
C43974 POR2X1_44/CTRL2 INPUT_6 0.03fF
C43975 POR2X1_276/a_16_28# POR2X1_325/A 0.00fF
C43976 PAND2X1_785/Y PAND2X1_514/Y 0.03fF
C43977 POR2X1_149/B VDD 0.38fF
C43978 POR2X1_13/A PAND2X1_658/A 0.03fF
C43979 POR2X1_853/A POR2X1_566/A 0.05fF
C43980 POR2X1_362/Y POR2X1_276/Y 0.40fF
C43981 POR2X1_302/O PAND2X1_6/Y 0.02fF
C43982 PAND2X1_565/CTRL VDD -0.00fF
C43983 POR2X1_559/Y VDD 0.20fF
C43984 POR2X1_102/Y POR2X1_172/O 0.03fF
C43985 POR2X1_840/B POR2X1_217/CTRL2 0.12fF
C43986 POR2X1_664/a_56_344# PAND2X1_73/Y 0.00fF
C43987 POR2X1_664/O POR2X1_78/A 0.08fF
C43988 POR2X1_45/Y PAND2X1_479/B 0.01fF
C43989 PAND2X1_494/O INPUT_0 0.16fF
C43990 POR2X1_315/Y PAND2X1_444/Y 0.08fF
C43991 POR2X1_38/Y POR2X1_5/Y 1.30fF
C43992 POR2X1_816/O POR2X1_39/B 0.06fF
C43993 POR2X1_406/Y POR2X1_52/Y 0.03fF
C43994 POR2X1_356/A POR2X1_477/A 0.03fF
C43995 POR2X1_32/A PAND2X1_727/a_16_344# 0.05fF
C43996 PAND2X1_673/O POR2X1_38/B 0.10fF
C43997 POR2X1_25/CTRL D_INPUT_6 0.01fF
C43998 POR2X1_66/B PAND2X1_94/A 0.10fF
C43999 POR2X1_355/B POR2X1_508/a_56_344# 0.00fF
C44000 PAND2X1_262/a_76_28# POR2X1_38/B 0.02fF
C44001 PAND2X1_209/A PAND2X1_209/O -0.00fF
C44002 PAND2X1_48/B PAND2X1_23/Y 1.77fF
C44003 PAND2X1_474/Y POR2X1_73/Y 0.03fF
C44004 POR2X1_110/Y POR2X1_23/Y 0.21fF
C44005 POR2X1_407/A POR2X1_114/Y 0.16fF
C44006 POR2X1_447/B POR2X1_629/O 0.06fF
C44007 PAND2X1_55/Y PAND2X1_178/CTRL 0.00fF
C44008 POR2X1_644/A VDD 0.19fF
C44009 POR2X1_376/B PAND2X1_168/O 0.15fF
C44010 POR2X1_294/B PAND2X1_110/O 0.31fF
C44011 POR2X1_661/A POR2X1_655/CTRL 0.06fF
C44012 POR2X1_62/Y D_INPUT_0 0.25fF
C44013 POR2X1_411/B PAND2X1_840/Y 0.03fF
C44014 POR2X1_156/B POR2X1_155/O 0.02fF
C44015 POR2X1_60/A PAND2X1_308/Y 0.03fF
C44016 PAND2X1_223/B PAND2X1_538/CTRL 0.01fF
C44017 POR2X1_188/A PAND2X1_94/A 0.17fF
C44018 POR2X1_327/Y POR2X1_78/A 0.10fF
C44019 POR2X1_272/Y POR2X1_91/Y 0.03fF
C44020 PAND2X1_778/Y VDD 0.17fF
C44021 POR2X1_13/A POR2X1_73/Y 0.54fF
C44022 POR2X1_52/A PAND2X1_642/B 0.04fF
C44023 PAND2X1_388/Y POR2X1_236/Y 0.01fF
C44024 PAND2X1_4/CTRL PAND2X1_8/Y 0.04fF
C44025 PAND2X1_219/A POR2X1_394/A 0.03fF
C44026 POR2X1_184/Y POR2X1_55/Y 0.09fF
C44027 POR2X1_478/B VDD 0.00fF
C44028 POR2X1_495/Y PAND2X1_840/A 0.01fF
C44029 PAND2X1_593/Y POR2X1_250/A 0.04fF
C44030 POR2X1_186/Y POR2X1_456/B 0.06fF
C44031 PAND2X1_90/Y POR2X1_181/B 0.03fF
C44032 POR2X1_376/B PAND2X1_550/B 0.05fF
C44033 PAND2X1_723/Y POR2X1_7/A 0.10fF
C44034 POR2X1_511/Y PAND2X1_349/A 0.00fF
C44035 POR2X1_83/B POR2X1_373/Y 0.05fF
C44036 POR2X1_750/B POR2X1_353/A 0.03fF
C44037 PAND2X1_215/B PAND2X1_723/CTRL 0.03fF
C44038 POR2X1_316/Y PAND2X1_436/O 0.01fF
C44039 POR2X1_781/A POR2X1_568/Y 0.04fF
C44040 POR2X1_193/A POR2X1_631/B 0.03fF
C44041 POR2X1_32/A PAND2X1_199/B 0.00fF
C44042 PAND2X1_549/B POR2X1_236/Y 0.10fF
C44043 POR2X1_294/B POR2X1_713/Y 0.00fF
C44044 PAND2X1_371/O PAND2X1_32/B 0.01fF
C44045 POR2X1_805/A POR2X1_710/CTRL2 0.00fF
C44046 PAND2X1_6/Y PAND2X1_7/CTRL 0.01fF
C44047 POR2X1_43/B PAND2X1_798/B 0.01fF
C44048 PAND2X1_651/Y POR2X1_55/Y 0.09fF
C44049 POR2X1_41/B POR2X1_152/m4_208_n4# 0.01fF
C44050 PAND2X1_662/O POR2X1_413/A 0.02fF
C44051 POR2X1_809/A POR2X1_812/A 0.08fF
C44052 PAND2X1_55/Y POR2X1_556/Y 0.59fF
C44053 POR2X1_198/B PAND2X1_69/A 0.03fF
C44054 PAND2X1_437/O POR2X1_440/B 0.01fF
C44055 PAND2X1_65/B POR2X1_703/A 0.05fF
C44056 POR2X1_356/A PAND2X1_747/CTRL 0.04fF
C44057 POR2X1_669/B POR2X1_4/Y 0.03fF
C44058 PAND2X1_631/A POR2X1_496/Y 0.03fF
C44059 POR2X1_274/B VDD 0.00fF
C44060 POR2X1_791/CTRL2 POR2X1_791/A 0.01fF
C44061 PAND2X1_844/O POR2X1_60/Y 0.02fF
C44062 PAND2X1_844/CTRL2 PAND2X1_61/Y 0.01fF
C44063 INPUT_1 POR2X1_5/Y 0.42fF
C44064 PAND2X1_341/A PAND2X1_101/CTRL 0.01fF
C44065 POR2X1_78/B PAND2X1_232/CTRL -0.04fF
C44066 POR2X1_579/Y PAND2X1_173/CTRL2 0.00fF
C44067 POR2X1_192/Y POR2X1_704/O 0.02fF
C44068 PAND2X1_575/B PAND2X1_716/B 0.03fF
C44069 POR2X1_428/O POR2X1_236/Y 0.01fF
C44070 POR2X1_337/a_16_28# POR2X1_335/Y -0.00fF
C44071 POR2X1_121/B POR2X1_691/A 0.03fF
C44072 PAND2X1_835/O PAND2X1_852/B 0.05fF
C44073 PAND2X1_551/Y POR2X1_90/Y 0.01fF
C44074 POR2X1_60/CTRL PAND2X1_339/Y 0.01fF
C44075 POR2X1_13/A PAND2X1_244/B 0.06fF
C44076 POR2X1_654/B POR2X1_768/Y 0.02fF
C44077 POR2X1_114/B POR2X1_840/B 0.05fF
C44078 POR2X1_76/Y POR2X1_553/A 0.02fF
C44079 POR2X1_834/Y POR2X1_130/A 0.05fF
C44080 POR2X1_46/Y PAND2X1_723/A 0.07fF
C44081 POR2X1_751/a_16_28# POR2X1_7/B 0.02fF
C44082 PAND2X1_488/CTRL POR2X1_294/A 0.03fF
C44083 POR2X1_5/Y POR2X1_153/Y 0.37fF
C44084 POR2X1_96/A PAND2X1_346/Y 0.03fF
C44085 PAND2X1_243/B POR2X1_235/Y 0.00fF
C44086 POR2X1_16/A PAND2X1_520/O 0.15fF
C44087 PAND2X1_72/Y VDD 0.14fF
C44088 POR2X1_384/A POR2X1_5/Y 0.05fF
C44089 PAND2X1_23/Y PAND2X1_757/a_16_344# 0.01fF
C44090 POR2X1_52/A PAND2X1_550/B 0.03fF
C44091 PAND2X1_642/O VDD 0.00fF
C44092 POR2X1_66/B PAND2X1_136/CTRL2 0.01fF
C44093 POR2X1_435/Y PAND2X1_533/CTRL2 0.05fF
C44094 POR2X1_763/Y POR2X1_321/Y 0.03fF
C44095 PAND2X1_209/A PAND2X1_161/Y 0.00fF
C44096 PAND2X1_661/B POR2X1_73/Y 0.03fF
C44097 POR2X1_347/A POR2X1_404/B 0.05fF
C44098 PAND2X1_643/Y POR2X1_73/Y 3.87fF
C44099 POR2X1_212/a_16_28# POR2X1_568/A 0.03fF
C44100 POR2X1_407/A POR2X1_113/Y 0.01fF
C44101 PAND2X1_386/Y POR2X1_260/A 0.01fF
C44102 POR2X1_101/Y POR2X1_717/Y 0.03fF
C44103 PAND2X1_72/CTRL2 PAND2X1_60/B 0.10fF
C44104 INPUT_1 POR2X1_20/CTRL 0.01fF
C44105 POR2X1_844/O D_INPUT_1 0.02fF
C44106 PAND2X1_672/O PAND2X1_671/Y 0.00fF
C44107 PAND2X1_48/CTRL POR2X1_186/B 0.01fF
C44108 POR2X1_78/B POR2X1_195/CTRL2 0.01fF
C44109 POR2X1_741/Y POR2X1_274/B 0.10fF
C44110 POR2X1_740/Y POR2X1_553/A 0.05fF
C44111 PAND2X1_140/A PAND2X1_566/Y 0.03fF
C44112 INPUT_0 PAND2X1_853/B 0.03fF
C44113 PAND2X1_79/Y POR2X1_84/Y 0.10fF
C44114 POR2X1_51/B POR2X1_587/Y 0.01fF
C44115 PAND2X1_126/O POR2X1_68/A 0.08fF
C44116 PAND2X1_449/CTRL POR2X1_329/A 0.02fF
C44117 PAND2X1_65/B PAND2X1_167/CTRL2 0.01fF
C44118 POR2X1_110/Y POR2X1_368/CTRL2 0.01fF
C44119 POR2X1_685/A POR2X1_407/A 0.02fF
C44120 POR2X1_839/O POR2X1_191/Y 0.33fF
C44121 POR2X1_60/A POR2X1_77/Y 13.94fF
C44122 POR2X1_845/O D_INPUT_1 0.04fF
C44123 POR2X1_415/Y POR2X1_260/A 0.02fF
C44124 POR2X1_719/B PAND2X1_48/B 0.04fF
C44125 POR2X1_16/A PAND2X1_602/Y 0.03fF
C44126 PAND2X1_824/B POR2X1_198/B 0.71fF
C44127 POR2X1_505/CTRL2 PAND2X1_6/A 0.04fF
C44128 POR2X1_407/Y PAND2X1_765/CTRL2 0.01fF
C44129 POR2X1_220/Y POR2X1_737/A 0.03fF
C44130 PAND2X1_57/B POR2X1_342/CTRL 0.01fF
C44131 POR2X1_591/A POR2X1_77/Y 0.00fF
C44132 POR2X1_274/B PAND2X1_32/B 0.05fF
C44133 POR2X1_327/Y PAND2X1_604/CTRL2 0.00fF
C44134 PAND2X1_794/B POR2X1_534/Y 0.35fF
C44135 INPUT_0 POR2X1_572/Y 0.04fF
C44136 PAND2X1_467/Y POR2X1_694/O 0.01fF
C44137 POR2X1_277/O PAND2X1_560/B 0.01fF
C44138 POR2X1_294/B POR2X1_559/A 0.06fF
C44139 POR2X1_52/A PAND2X1_620/a_76_28# 0.01fF
C44140 POR2X1_278/Y POR2X1_385/Y 0.10fF
C44141 PAND2X1_723/a_76_28# PAND2X1_656/A 0.01fF
C44142 PAND2X1_348/A PAND2X1_514/Y 0.11fF
C44143 POR2X1_407/A POR2X1_260/A 0.08fF
C44144 POR2X1_73/Y PAND2X1_510/B 0.00fF
C44145 PAND2X1_330/O VDD 0.00fF
C44146 PAND2X1_651/Y PAND2X1_510/CTRL2 0.04fF
C44147 POR2X1_205/A PAND2X1_63/B 0.01fF
C44148 POR2X1_280/CTRL2 POR2X1_280/Y 0.01fF
C44149 POR2X1_276/A POR2X1_318/A 0.02fF
C44150 POR2X1_316/Y PAND2X1_499/Y 5.61fF
C44151 PAND2X1_563/a_16_344# POR2X1_394/A 0.02fF
C44152 PAND2X1_784/O PAND2X1_156/A 0.02fF
C44153 POR2X1_143/O PAND2X1_341/B 0.02fF
C44154 POR2X1_65/Y PAND2X1_206/B 0.00fF
C44155 PAND2X1_61/Y PAND2X1_339/O 0.02fF
C44156 POR2X1_132/a_16_28# POR2X1_96/A 0.06fF
C44157 PAND2X1_859/CTRL POR2X1_77/Y 0.01fF
C44158 POR2X1_293/Y POR2X1_371/O 0.15fF
C44159 POR2X1_52/A POR2X1_616/Y 0.06fF
C44160 POR2X1_832/B POR2X1_652/A 0.05fF
C44161 POR2X1_57/A POR2X1_291/CTRL 0.01fF
C44162 POR2X1_8/Y INPUT_2 0.02fF
C44163 POR2X1_394/A POR2X1_816/A 0.22fF
C44164 POR2X1_537/Y POR2X1_733/A 0.25fF
C44165 POR2X1_188/CTRL2 POR2X1_456/B 0.00fF
C44166 POR2X1_68/A PAND2X1_142/a_16_344# 0.01fF
C44167 D_INPUT_1 POR2X1_394/A 0.01fF
C44168 POR2X1_307/B PAND2X1_56/A 0.01fF
C44169 D_INPUT_1 POR2X1_749/CTRL 0.01fF
C44170 POR2X1_88/O PAND2X1_206/B 0.00fF
C44171 POR2X1_687/A POR2X1_729/Y 0.04fF
C44172 POR2X1_862/O POR2X1_480/A 0.20fF
C44173 POR2X1_318/CTRL POR2X1_471/A 0.16fF
C44174 POR2X1_101/Y POR2X1_218/CTRL 0.05fF
C44175 PAND2X1_244/B PAND2X1_510/B 0.03fF
C44176 POR2X1_78/B POR2X1_500/CTRL2 0.08fF
C44177 POR2X1_130/O POR2X1_318/A 0.03fF
C44178 PAND2X1_631/A PAND2X1_514/Y 0.01fF
C44179 PAND2X1_69/A POR2X1_342/CTRL2 0.03fF
C44180 POR2X1_192/Y POR2X1_567/O 0.00fF
C44181 PAND2X1_847/CTRL2 POR2X1_820/Y 0.01fF
C44182 POR2X1_304/O POR2X1_56/B 0.00fF
C44183 POR2X1_730/Y POR2X1_738/A 0.03fF
C44184 POR2X1_293/Y PAND2X1_358/CTRL2 0.03fF
C44185 PAND2X1_193/Y PAND2X1_733/A 0.01fF
C44186 PAND2X1_734/m4_208_n4# PAND2X1_560/B 0.07fF
C44187 POR2X1_537/a_76_344# POR2X1_537/B 0.01fF
C44188 POR2X1_251/Y POR2X1_416/B 2.80fF
C44189 POR2X1_566/A PAND2X1_292/CTRL 0.11fF
C44190 POR2X1_276/A POR2X1_574/Y 0.02fF
C44191 PAND2X1_152/O POR2X1_711/Y 0.08fF
C44192 PAND2X1_349/A POR2X1_129/Y 0.03fF
C44193 POR2X1_51/A POR2X1_64/CTRL 0.01fF
C44194 PAND2X1_474/O PAND2X1_404/Y 0.01fF
C44195 PAND2X1_48/B POR2X1_711/Y 0.20fF
C44196 PAND2X1_785/Y PAND2X1_332/Y 0.03fF
C44197 POR2X1_54/Y POR2X1_77/O 0.03fF
C44198 PAND2X1_849/B PAND2X1_100/a_76_28# 0.01fF
C44199 POR2X1_383/A POR2X1_266/A 0.03fF
C44200 PAND2X1_47/a_16_344# PAND2X1_59/B 0.03fF
C44201 POR2X1_78/B PAND2X1_125/O 0.09fF
C44202 POR2X1_151/CTRL POR2X1_186/B 0.01fF
C44203 PAND2X1_787/A PAND2X1_353/Y 0.12fF
C44204 POR2X1_69/CTRL2 PAND2X1_206/B 0.00fF
C44205 PAND2X1_62/CTRL2 POR2X1_9/Y 0.03fF
C44206 POR2X1_69/CTRL POR2X1_67/Y 0.01fF
C44207 POR2X1_307/B POR2X1_661/A 0.01fF
C44208 PAND2X1_813/a_76_28# POR2X1_673/Y 0.02fF
C44209 POR2X1_504/Y POR2X1_846/A 0.01fF
C44210 POR2X1_477/A PAND2X1_72/A 0.06fF
C44211 PAND2X1_530/O PAND2X1_52/B 0.04fF
C44212 PAND2X1_94/A POR2X1_54/O 0.18fF
C44213 POR2X1_130/O POR2X1_574/Y 0.01fF
C44214 PAND2X1_287/Y PAND2X1_578/Y 0.01fF
C44215 POR2X1_840/B POR2X1_513/A 0.00fF
C44216 PAND2X1_665/CTRL PAND2X1_60/B 0.01fF
C44217 POR2X1_567/A POR2X1_725/Y 0.07fF
C44218 POR2X1_597/Y POR2X1_669/B 0.00fF
C44219 PAND2X1_206/B POR2X1_750/B 0.03fF
C44220 POR2X1_60/A PAND2X1_449/O 0.01fF
C44221 POR2X1_96/Y PAND2X1_63/B 0.03fF
C44222 POR2X1_78/B PAND2X1_628/a_56_28# 0.00fF
C44223 POR2X1_567/B POR2X1_434/CTRL2 0.17fF
C44224 PAND2X1_22/CTRL PAND2X1_3/A 0.01fF
C44225 PAND2X1_860/A POR2X1_46/Y 0.05fF
C44226 POR2X1_66/B POR2X1_460/Y 0.03fF
C44227 INPUT_6 D_INPUT_4 0.93fF
C44228 POR2X1_407/A PAND2X1_681/O 0.05fF
C44229 POR2X1_294/Y POR2X1_202/A 0.00fF
C44230 POR2X1_13/A PAND2X1_458/CTRL2 0.00fF
C44231 POR2X1_624/Y POR2X1_29/A 0.03fF
C44232 POR2X1_815/a_76_344# POR2X1_750/A 0.00fF
C44233 POR2X1_66/B PAND2X1_43/CTRL2 0.03fF
C44234 PAND2X1_9/O PAND2X1_9/Y 0.02fF
C44235 POR2X1_9/Y PAND2X1_751/CTRL2 0.03fF
C44236 POR2X1_864/A POR2X1_780/O 0.00fF
C44237 POR2X1_300/Y POR2X1_75/Y 0.00fF
C44238 POR2X1_726/Y POR2X1_568/B 0.02fF
C44239 POR2X1_294/A POR2X1_195/CTRL2 0.04fF
C44240 POR2X1_862/A POR2X1_590/A 0.08fF
C44241 PAND2X1_96/B POR2X1_579/CTRL2 0.00fF
C44242 POR2X1_63/Y PAND2X1_231/CTRL2 0.01fF
C44243 PAND2X1_109/a_16_344# POR2X1_854/B 0.07fF
C44244 PAND2X1_569/B POR2X1_39/B 0.07fF
C44245 POR2X1_302/Y POR2X1_814/A 0.02fF
C44246 POR2X1_158/B POR2X1_39/B 0.02fF
C44247 PAND2X1_405/O POR2X1_46/Y 0.06fF
C44248 POR2X1_16/A POR2X1_767/Y 0.08fF
C44249 POR2X1_703/A POR2X1_542/a_16_28# 0.03fF
C44250 POR2X1_741/CTRL POR2X1_741/B 0.04fF
C44251 PAND2X1_831/O POR2X1_411/B 0.03fF
C44252 POR2X1_49/Y PAND2X1_9/Y 0.10fF
C44253 POR2X1_54/Y PAND2X1_35/B 0.02fF
C44254 POR2X1_63/Y POR2X1_230/CTRL2 0.01fF
C44255 POR2X1_39/B POR2X1_172/a_16_28# 0.01fF
C44256 POR2X1_835/B POR2X1_835/Y 0.01fF
C44257 POR2X1_610/CTRL2 PAND2X1_41/B 0.03fF
C44258 POR2X1_260/B POR2X1_405/O 0.02fF
C44259 POR2X1_621/B POR2X1_621/A 0.12fF
C44260 PAND2X1_499/m4_208_n4# POR2X1_20/B 0.09fF
C44261 POR2X1_250/Y POR2X1_42/Y 0.03fF
C44262 PAND2X1_73/Y POR2X1_590/A 0.30fF
C44263 POR2X1_67/Y POR2X1_619/CTRL2 0.01fF
C44264 POR2X1_728/A POR2X1_210/B 0.02fF
C44265 POR2X1_195/A POR2X1_852/B 0.03fF
C44266 POR2X1_566/A POR2X1_443/O 0.05fF
C44267 POR2X1_56/O POR2X1_83/B 0.02fF
C44268 POR2X1_354/O POR2X1_319/Y 0.01fF
C44269 POR2X1_144/m4_208_n4# PAND2X1_797/Y 0.09fF
C44270 PAND2X1_20/A POR2X1_33/CTRL 0.01fF
C44271 POR2X1_703/A PAND2X1_178/CTRL2 0.01fF
C44272 POR2X1_9/Y POR2X1_68/B 0.00fF
C44273 POR2X1_191/O POR2X1_191/Y 0.06fF
C44274 PAND2X1_234/CTRL PAND2X1_88/Y 0.01fF
C44275 PAND2X1_317/CTRL POR2X1_167/Y 0.01fF
C44276 POR2X1_707/B PAND2X1_25/O 0.01fF
C44277 POR2X1_248/A POR2X1_5/Y 0.01fF
C44278 PAND2X1_844/O PAND2X1_351/A 0.00fF
C44279 POR2X1_373/CTRL2 POR2X1_77/Y 0.01fF
C44280 POR2X1_66/B PAND2X1_11/Y 0.01fF
C44281 POR2X1_499/A POR2X1_575/B 0.05fF
C44282 POR2X1_736/A POR2X1_337/Y 0.10fF
C44283 POR2X1_180/CTRL POR2X1_181/Y 0.01fF
C44284 POR2X1_814/A POR2X1_501/B 0.03fF
C44285 POR2X1_66/B POR2X1_606/Y 0.03fF
C44286 POR2X1_548/CTRL2 POR2X1_66/A 0.03fF
C44287 POR2X1_260/B POR2X1_596/Y 0.01fF
C44288 POR2X1_27/O POR2X1_38/Y 0.05fF
C44289 POR2X1_343/A POR2X1_296/B 0.01fF
C44290 POR2X1_464/Y POR2X1_471/A 0.10fF
C44291 POR2X1_300/Y PAND2X1_332/Y 0.00fF
C44292 POR2X1_450/B PAND2X1_427/O 0.08fF
C44293 POR2X1_557/A PAND2X1_42/m4_208_n4# 0.01fF
C44294 POR2X1_14/Y POR2X1_94/A 1.20fF
C44295 PAND2X1_48/B PAND2X1_271/CTRL2 0.02fF
C44296 PAND2X1_211/CTRL POR2X1_55/Y 0.01fF
C44297 POR2X1_669/B PAND2X1_714/A 0.02fF
C44298 POR2X1_809/A PAND2X1_681/a_16_344# 0.01fF
C44299 PAND2X1_626/O POR2X1_750/B 0.05fF
C44300 POR2X1_624/Y PAND2X1_110/CTRL 0.01fF
C44301 POR2X1_23/Y INPUT_0 0.49fF
C44302 POR2X1_680/Y POR2X1_679/Y 0.02fF
C44303 POR2X1_679/O POR2X1_816/A 0.01fF
C44304 POR2X1_316/Y POR2X1_39/B 0.03fF
C44305 PAND2X1_23/Y D_INPUT_5 0.03fF
C44306 POR2X1_41/B PAND2X1_444/O 0.05fF
C44307 POR2X1_254/A POR2X1_750/B 0.03fF
C44308 PAND2X1_48/B POR2X1_632/CTRL2 0.01fF
C44309 PAND2X1_225/a_16_344# POR2X1_750/B 0.01fF
C44310 PAND2X1_717/A PAND2X1_175/B 0.03fF
C44311 POR2X1_326/A POR2X1_863/A 0.04fF
C44312 PAND2X1_85/Y POR2X1_296/B 0.00fF
C44313 POR2X1_260/B POR2X1_795/CTRL2 0.00fF
C44314 PAND2X1_793/Y POR2X1_67/a_16_28# 0.02fF
C44315 POR2X1_72/B POR2X1_40/Y 0.21fF
C44316 POR2X1_861/O POR2X1_624/Y 0.02fF
C44317 POR2X1_13/A POR2X1_299/Y 0.02fF
C44318 POR2X1_614/A POR2X1_452/O 0.01fF
C44319 PAND2X1_215/B PAND2X1_267/Y 0.01fF
C44320 PAND2X1_212/O POR2X1_55/Y 0.04fF
C44321 POR2X1_628/Y PAND2X1_6/A 0.03fF
C44322 POR2X1_67/CTRL2 PAND2X1_658/A 0.01fF
C44323 POR2X1_706/CTRL2 VDD -0.00fF
C44324 PAND2X1_58/A PAND2X1_589/O 0.02fF
C44325 PAND2X1_6/Y POR2X1_803/CTRL 0.01fF
C44326 PAND2X1_531/O POR2X1_549/B 0.00fF
C44327 POR2X1_675/O POR2X1_675/A 0.01fF
C44328 POR2X1_655/Y POR2X1_660/A 0.28fF
C44329 POR2X1_83/B POR2X1_397/Y 0.03fF
C44330 POR2X1_651/CTRL POR2X1_66/A 0.01fF
C44331 POR2X1_849/CTRL2 POR2X1_94/A 0.00fF
C44332 POR2X1_311/Y PAND2X1_347/Y 0.03fF
C44333 POR2X1_794/B POR2X1_830/A 0.01fF
C44334 PAND2X1_73/Y PAND2X1_760/CTRL 0.01fF
C44335 PAND2X1_13/O POR2X1_750/B 0.02fF
C44336 POR2X1_413/Y D_INPUT_0 0.01fF
C44337 PAND2X1_630/a_76_28# POR2X1_628/Y 0.02fF
C44338 POR2X1_814/A POR2X1_703/A 0.07fF
C44339 POR2X1_341/A PAND2X1_79/Y 2.56fF
C44340 POR2X1_260/B PAND2X1_536/O 0.09fF
C44341 PAND2X1_11/Y PAND2X1_18/a_76_28# 0.07fF
C44342 POR2X1_12/A PAND2X1_711/A 0.28fF
C44343 PAND2X1_6/Y POR2X1_260/B 3.89fF
C44344 PAND2X1_448/O POR2X1_42/Y 0.06fF
C44345 PAND2X1_106/O POR2X1_556/A 0.02fF
C44346 PAND2X1_137/Y POR2X1_102/Y 0.55fF
C44347 PAND2X1_560/a_76_28# POR2X1_73/Y 0.01fF
C44348 PAND2X1_777/a_76_28# POR2X1_7/B 0.01fF
C44349 POR2X1_706/B POR2X1_706/A 0.04fF
C44350 POR2X1_69/A POR2X1_88/Y 0.49fF
C44351 PAND2X1_661/Y POR2X1_411/B 0.03fF
C44352 POR2X1_376/B POR2X1_381/CTRL 0.01fF
C44353 POR2X1_331/Y VDD 0.27fF
C44354 POR2X1_760/A POR2X1_385/a_76_344# 0.00fF
C44355 PAND2X1_659/B POR2X1_72/B 0.15fF
C44356 POR2X1_814/A POR2X1_768/m4_208_n4# 0.09fF
C44357 POR2X1_502/A POR2X1_640/O 0.04fF
C44358 POR2X1_351/B POR2X1_814/A 0.04fF
C44359 PAND2X1_658/A POR2X1_29/A 0.04fF
C44360 PAND2X1_787/A POR2X1_298/CTRL2 0.03fF
C44361 POR2X1_477/m4_208_n4# POR2X1_854/B 0.07fF
C44362 POR2X1_626/Y POR2X1_627/Y 0.01fF
C44363 POR2X1_302/B POR2X1_220/Y 0.01fF
C44364 POR2X1_96/A PAND2X1_354/A 0.03fF
C44365 POR2X1_811/B POR2X1_294/B 0.01fF
C44366 PAND2X1_472/B POR2X1_94/A 1.08fF
C44367 POR2X1_66/A PAND2X1_518/CTRL 0.01fF
C44368 POR2X1_287/B VDD 0.71fF
C44369 D_INPUT_0 POR2X1_804/A 0.05fF
C44370 POR2X1_8/Y PAND2X1_227/O 0.04fF
C44371 PAND2X1_801/B VDD 0.03fF
C44372 POR2X1_804/CTRL POR2X1_532/A 0.01fF
C44373 PAND2X1_714/CTRL POR2X1_40/Y 0.01fF
C44374 POR2X1_62/O PAND2X1_58/A 0.01fF
C44375 POR2X1_122/A VDD -0.00fF
C44376 POR2X1_830/CTRL2 POR2X1_740/Y 0.01fF
C44377 POR2X1_49/Y PAND2X1_523/CTRL2 0.00fF
C44378 PAND2X1_20/A POR2X1_264/Y 0.03fF
C44379 POR2X1_525/CTRL2 POR2X1_46/Y 0.01fF
C44380 POR2X1_856/B PAND2X1_88/Y 0.36fF
C44381 POR2X1_626/CTRL2 POR2X1_93/A 0.01fF
C44382 POR2X1_669/B POR2X1_816/A 0.05fF
C44383 POR2X1_661/A POR2X1_513/A 0.08fF
C44384 PAND2X1_295/a_76_28# PAND2X1_60/B 0.01fF
C44385 PAND2X1_272/O POR2X1_112/Y 0.01fF
C44386 POR2X1_333/A POR2X1_795/B 0.03fF
C44387 POR2X1_483/A VDD 0.45fF
C44388 POR2X1_669/B D_INPUT_1 0.16fF
C44389 POR2X1_41/B GATE_479 0.03fF
C44390 POR2X1_62/a_16_28# POR2X1_29/A 0.03fF
C44391 POR2X1_475/A PAND2X1_372/CTRL 0.02fF
C44392 POR2X1_114/B PAND2X1_279/CTRL 0.01fF
C44393 POR2X1_590/A POR2X1_631/B 0.12fF
C44394 INPUT_0 PAND2X1_558/O 0.04fF
C44395 POR2X1_65/A PAND2X1_714/CTRL2 0.03fF
C44396 POR2X1_94/A POR2X1_55/Y 0.04fF
C44397 POR2X1_822/O VDD 0.00fF
C44398 POR2X1_763/Y PAND2X1_738/CTRL2 0.05fF
C44399 PAND2X1_61/Y POR2X1_58/Y 0.01fF
C44400 PAND2X1_56/Y POR2X1_830/O 0.02fF
C44401 PAND2X1_593/CTRL INPUT_0 0.01fF
C44402 PAND2X1_211/A PAND2X1_724/B 0.25fF
C44403 POR2X1_43/B PAND2X1_195/O 0.04fF
C44404 PAND2X1_8/Y VDD 0.85fF
C44405 POR2X1_409/B PAND2X1_338/B 0.03fF
C44406 POR2X1_60/A POR2X1_52/Y 0.03fF
C44407 POR2X1_121/A POR2X1_654/CTRL 0.00fF
C44408 POR2X1_850/B PAND2X1_69/A 0.03fF
C44409 PAND2X1_67/CTRL2 POR2X1_507/A 0.02fF
C44410 POR2X1_661/CTRL2 POR2X1_740/Y 0.00fF
C44411 PAND2X1_63/Y POR2X1_641/O 0.11fF
C44412 POR2X1_514/CTRL POR2X1_777/B 0.00fF
C44413 POR2X1_37/Y PAND2X1_349/A 0.01fF
C44414 POR2X1_294/B PAND2X1_525/O -0.00fF
C44415 PAND2X1_675/A PAND2X1_540/O 0.04fF
C44416 POR2X1_57/A PAND2X1_721/B 0.03fF
C44417 POR2X1_20/B PAND2X1_345/Y 0.01fF
C44418 POR2X1_404/CTRL POR2X1_35/Y 0.01fF
C44419 POR2X1_37/Y PAND2X1_63/B 0.03fF
C44420 PAND2X1_382/CTRL2 POR2X1_29/A 0.01fF
C44421 INPUT_2 POR2X1_609/CTRL2 0.01fF
C44422 POR2X1_48/A PAND2X1_569/B 0.07fF
C44423 POR2X1_170/B VDD 0.14fF
C44424 POR2X1_267/CTRL POR2X1_318/A 0.04fF
C44425 POR2X1_14/Y POR2X1_583/CTRL 0.01fF
C44426 PAND2X1_225/CTRL2 POR2X1_68/B 0.01fF
C44427 POR2X1_174/CTRL2 POR2X1_567/B 0.05fF
C44428 POR2X1_428/Y POR2X1_394/A 0.01fF
C44429 POR2X1_345/A PAND2X1_6/Y 0.00fF
C44430 POR2X1_13/A PAND2X1_785/Y 0.16fF
C44431 POR2X1_493/A POR2X1_773/B 0.08fF
C44432 POR2X1_251/Y PAND2X1_738/Y 0.30fF
C44433 POR2X1_296/B POR2X1_575/O 0.02fF
C44434 POR2X1_66/B POR2X1_98/B 0.02fF
C44435 PAND2X1_241/Y POR2X1_60/A 0.08fF
C44436 PAND2X1_58/A PAND2X1_757/O 0.17fF
C44437 POR2X1_808/A POR2X1_644/A 0.01fF
C44438 PAND2X1_206/a_56_28# POR2X1_293/Y 0.00fF
C44439 PAND2X1_790/Y VDD 0.12fF
C44440 POR2X1_52/A PAND2X1_445/Y 0.23fF
C44441 PAND2X1_420/CTRL2 POR2X1_510/Y 0.01fF
C44442 POR2X1_483/A POR2X1_741/Y 0.03fF
C44443 POR2X1_500/A PAND2X1_79/Y 0.64fF
C44444 POR2X1_388/CTRL2 PAND2X1_65/B 0.01fF
C44445 POR2X1_502/A POR2X1_638/CTRL 0.02fF
C44446 POR2X1_93/Y POR2X1_394/A 0.07fF
C44447 POR2X1_138/CTRL POR2X1_130/A 0.04fF
C44448 POR2X1_78/A POR2X1_590/O 0.02fF
C44449 PAND2X1_476/A POR2X1_63/Y 0.04fF
C44450 POR2X1_365/Y POR2X1_502/A 0.03fF
C44451 POR2X1_287/B PAND2X1_32/B 0.07fF
C44452 POR2X1_660/Y POR2X1_308/B 0.01fF
C44453 POR2X1_754/Y POR2X1_260/A 0.07fF
C44454 POR2X1_376/B POR2X1_386/CTRL2 0.00fF
C44455 POR2X1_208/A POR2X1_201/O 0.00fF
C44456 POR2X1_809/A POR2X1_796/Y 0.14fF
C44457 PAND2X1_673/a_76_28# POR2X1_670/Y 0.02fF
C44458 POR2X1_61/B VDD 0.22fF
C44459 POR2X1_65/A POR2X1_597/CTRL2 0.03fF
C44460 PAND2X1_651/Y POR2X1_511/Y 0.03fF
C44461 PAND2X1_553/CTRL POR2X1_106/Y 0.01fF
C44462 POR2X1_56/B PAND2X1_453/CTRL 0.06fF
C44463 POR2X1_78/B PAND2X1_743/CTRL2 0.03fF
C44464 POR2X1_52/A PAND2X1_506/CTRL2 0.03fF
C44465 POR2X1_841/B POR2X1_737/A 0.03fF
C44466 POR2X1_247/CTRL2 POR2X1_294/B 0.01fF
C44467 INPUT_1 PAND2X1_623/a_16_344# 0.01fF
C44468 POR2X1_389/Y PAND2X1_60/B 0.03fF
C44469 POR2X1_68/A POR2X1_676/Y 0.03fF
C44470 POR2X1_833/A POR2X1_296/B 0.06fF
C44471 PAND2X1_793/Y PAND2X1_575/A 0.00fF
C44472 PAND2X1_462/B POR2X1_232/O 0.32fF
C44473 POR2X1_84/Y POR2X1_786/CTRL2 0.01fF
C44474 POR2X1_119/Y POR2X1_271/CTRL 0.06fF
C44475 PAND2X1_243/B POR2X1_42/Y 0.03fF
C44476 D_INPUT_3 POR2X1_381/CTRL2 0.13fF
C44477 PAND2X1_6/Y POR2X1_464/a_16_28# 0.03fF
C44478 POR2X1_244/B POR2X1_562/B 0.02fF
C44479 POR2X1_193/A POR2X1_193/CTRL 0.02fF
C44480 POR2X1_409/Y POR2X1_14/Y 0.03fF
C44481 PAND2X1_653/Y VDD 0.29fF
C44482 POR2X1_38/Y PAND2X1_723/Y 0.00fF
C44483 PAND2X1_362/B POR2X1_594/A 0.02fF
C44484 POR2X1_776/A POR2X1_568/B 0.01fF
C44485 PAND2X1_40/a_16_344# PAND2X1_587/Y 0.02fF
C44486 PAND2X1_8/Y PAND2X1_32/B 0.14fF
C44487 POR2X1_476/A POR2X1_294/A 0.07fF
C44488 PAND2X1_48/B POR2X1_334/B 0.07fF
C44489 PAND2X1_793/Y PAND2X1_794/B 0.00fF
C44490 POR2X1_32/A POR2X1_129/Y 0.03fF
C44491 POR2X1_261/A PAND2X1_284/Y 0.00fF
C44492 POR2X1_509/A POR2X1_857/B 0.12fF
C44493 PAND2X1_140/A POR2X1_107/CTRL2 0.01fF
C44494 PAND2X1_439/a_76_28# POR2X1_167/Y 0.01fF
C44495 POR2X1_407/Y POR2X1_596/Y 0.01fF
C44496 POR2X1_508/A POR2X1_856/B 2.44fF
C44497 POR2X1_134/Y PAND2X1_768/CTRL 0.01fF
C44498 POR2X1_807/A POR2X1_725/Y 0.02fF
C44499 POR2X1_209/A VDD 0.42fF
C44500 POR2X1_554/B PAND2X1_72/A 0.56fF
C44501 POR2X1_579/Y POR2X1_35/Y 0.03fF
C44502 POR2X1_20/Y POR2X1_7/B 0.02fF
C44503 PAND2X1_182/A PAND2X1_182/O 0.03fF
C44504 POR2X1_54/Y POR2X1_39/B 0.07fF
C44505 POR2X1_102/Y PAND2X1_853/B 0.06fF
C44506 POR2X1_620/A POR2X1_620/B 0.01fF
C44507 PAND2X1_200/CTRL POR2X1_153/Y 0.08fF
C44508 PAND2X1_55/Y PAND2X1_536/O 0.07fF
C44509 PAND2X1_661/Y PAND2X1_596/CTRL2 0.00fF
C44510 PAND2X1_833/CTRL POR2X1_283/A 0.01fF
C44511 POR2X1_709/CTRL PAND2X1_90/Y 0.01fF
C44512 POR2X1_343/Y PAND2X1_39/B 0.02fF
C44513 POR2X1_836/a_76_344# POR2X1_192/B 0.02fF
C44514 POR2X1_836/O POR2X1_191/Y -0.01fF
C44515 PAND2X1_6/Y POR2X1_205/Y 0.03fF
C44516 POR2X1_174/O POR2X1_175/A 0.01fF
C44517 PAND2X1_6/Y PAND2X1_369/O 0.02fF
C44518 POR2X1_562/CTRL POR2X1_562/B 0.01fF
C44519 PAND2X1_814/CTRL POR2X1_7/B 0.01fF
C44520 PAND2X1_58/A PAND2X1_142/a_16_344# 0.01fF
C44521 PAND2X1_6/Y PAND2X1_55/Y 5.57fF
C44522 PAND2X1_659/Y POR2X1_32/A 0.06fF
C44523 PAND2X1_48/B POR2X1_124/B 0.01fF
C44524 POR2X1_57/A POR2X1_693/O 0.02fF
C44525 PAND2X1_226/O PAND2X1_32/B 0.07fF
C44526 PAND2X1_727/a_76_28# PAND2X1_444/Y 0.04fF
C44527 POR2X1_297/Y PAND2X1_854/A 0.02fF
C44528 POR2X1_480/A POR2X1_796/A 0.07fF
C44529 PAND2X1_81/B PAND2X1_316/CTRL2 0.02fF
C44530 POR2X1_250/CTRL POR2X1_283/A 0.01fF
C44531 POR2X1_260/B POR2X1_632/Y 0.03fF
C44532 POR2X1_188/A POR2X1_733/Y 0.58fF
C44533 POR2X1_547/CTRL POR2X1_614/A 0.04fF
C44534 PAND2X1_84/Y PAND2X1_717/Y 0.01fF
C44535 POR2X1_316/Y POR2X1_48/A 0.03fF
C44536 POR2X1_41/B POR2X1_142/Y 0.12fF
C44537 PAND2X1_56/Y POR2X1_786/Y 0.10fF
C44538 POR2X1_13/A PAND2X1_656/A 0.05fF
C44539 INPUT_1 PAND2X1_65/B 0.03fF
C44540 POR2X1_786/Y POR2X1_795/B 0.05fF
C44541 PAND2X1_20/A POR2X1_502/Y 0.00fF
C44542 POR2X1_238/Y POR2X1_90/Y 0.06fF
C44543 POR2X1_96/Y POR2X1_32/A 0.03fF
C44544 PAND2X1_562/B PAND2X1_348/A 2.57fF
C44545 POR2X1_92/O POR2X1_7/B 0.01fF
C44546 PAND2X1_90/Y PAND2X1_313/O 0.01fF
C44547 POR2X1_192/Y POR2X1_727/CTRL 0.05fF
C44548 PAND2X1_625/CTRL2 PAND2X1_96/B 0.00fF
C44549 POR2X1_253/Y PAND2X1_6/A 0.02fF
C44550 POR2X1_119/Y PAND2X1_446/m4_208_n4# 0.08fF
C44551 POR2X1_145/O PAND2X1_213/Y 0.01fF
C44552 PAND2X1_214/B PAND2X1_656/A 0.02fF
C44553 POR2X1_29/Y PAND2X1_6/A 0.05fF
C44554 POR2X1_390/B POR2X1_130/A 0.03fF
C44555 POR2X1_89/O PAND2X1_333/Y 0.02fF
C44556 POR2X1_833/CTRL2 PAND2X1_60/B 0.03fF
C44557 POR2X1_536/Y POR2X1_385/Y 0.09fF
C44558 PAND2X1_275/a_16_344# POR2X1_532/A 0.01fF
C44559 POR2X1_260/B PAND2X1_52/B 0.18fF
C44560 PAND2X1_349/A POR2X1_293/Y 0.03fF
C44561 POR2X1_673/Y PAND2X1_8/Y 0.04fF
C44562 PAND2X1_127/O POR2X1_78/B 0.16fF
C44563 POR2X1_156/CTRL2 POR2X1_750/B 0.01fF
C44564 POR2X1_319/O POR2X1_319/Y 0.01fF
C44565 POR2X1_390/B POR2X1_566/A 0.03fF
C44566 POR2X1_730/Y POR2X1_155/O 0.01fF
C44567 PAND2X1_197/O PAND2X1_656/A 0.02fF
C44568 PAND2X1_220/O PAND2X1_213/Y 0.09fF
C44569 POR2X1_16/A POR2X1_88/Y 0.00fF
C44570 PAND2X1_35/B POR2X1_4/Y 0.00fF
C44571 PAND2X1_857/A POR2X1_42/Y 0.10fF
C44572 POR2X1_614/A POR2X1_335/B 0.07fF
C44573 PAND2X1_6/Y POR2X1_783/Y 0.01fF
C44574 INPUT_2 POR2X1_68/B 0.03fF
C44575 POR2X1_368/Y POR2X1_91/Y 0.02fF
C44576 POR2X1_137/Y POR2X1_267/Y 0.02fF
C44577 POR2X1_157/a_16_28# POR2X1_36/B 0.03fF
C44578 POR2X1_409/Y PAND2X1_472/B 0.02fF
C44579 POR2X1_334/CTRL POR2X1_360/A 0.01fF
C44580 POR2X1_124/O POR2X1_773/B -0.02fF
C44581 PAND2X1_808/Y PAND2X1_363/CTRL 0.01fF
C44582 POR2X1_68/B PAND2X1_518/O 0.07fF
C44583 PAND2X1_732/O POR2X1_39/B 0.03fF
C44584 POR2X1_13/A PAND2X1_348/A 0.08fF
C44585 POR2X1_691/O POR2X1_855/B 0.01fF
C44586 POR2X1_567/A POR2X1_776/CTRL 0.02fF
C44587 POR2X1_832/A POR2X1_435/CTRL2 0.00fF
C44588 POR2X1_299/a_76_344# POR2X1_90/Y 0.00fF
C44589 PAND2X1_552/O PAND2X1_552/B 0.04fF
C44590 POR2X1_131/A PAND2X1_140/Y 0.00fF
C44591 POR2X1_777/B PAND2X1_136/CTRL 0.00fF
C44592 POR2X1_595/Y PAND2X1_643/A 0.04fF
C44593 PAND2X1_435/O POR2X1_153/Y 0.15fF
C44594 POR2X1_730/Y POR2X1_532/Y 0.73fF
C44595 POR2X1_407/A POR2X1_725/Y 0.07fF
C44596 POR2X1_614/A POR2X1_123/A 0.03fF
C44597 PAND2X1_784/A POR2X1_39/B 0.03fF
C44598 POR2X1_409/Y POR2X1_55/Y 0.01fF
C44599 PAND2X1_693/O PAND2X1_94/A 0.01fF
C44600 POR2X1_42/Y POR2X1_260/A 0.07fF
C44601 POR2X1_383/A POR2X1_786/Y 0.07fF
C44602 POR2X1_101/CTRL2 PAND2X1_69/A 0.04fF
C44603 POR2X1_343/Y PAND2X1_20/A 0.05fF
C44604 POR2X1_816/A POR2X1_171/CTRL2 0.01fF
C44605 POR2X1_13/A POR2X1_300/Y 0.83fF
C44606 POR2X1_145/CTRL2 POR2X1_394/A 0.01fF
C44607 POR2X1_147/CTRL POR2X1_78/A 0.03fF
C44608 POR2X1_57/A PAND2X1_803/Y 0.05fF
C44609 PAND2X1_661/B PAND2X1_656/A 0.03fF
C44610 PAND2X1_691/Y POR2X1_683/Y 1.25fF
C44611 INPUT_1 D_INPUT_2 0.02fF
C44612 POR2X1_809/A POR2X1_728/B 0.01fF
C44613 POR2X1_537/Y POR2X1_733/a_16_28# 0.02fF
C44614 POR2X1_75/a_76_344# PAND2X1_349/A 0.00fF
C44615 POR2X1_305/CTRL POR2X1_40/Y 0.01fF
C44616 POR2X1_110/Y PAND2X1_471/CTRL 0.00fF
C44617 POR2X1_569/A POR2X1_702/A 0.03fF
C44618 PAND2X1_659/Y PAND2X1_741/O 0.10fF
C44619 POR2X1_278/Y POR2X1_265/Y 0.05fF
C44620 PAND2X1_850/Y PAND2X1_276/CTRL 0.01fF
C44621 PAND2X1_297/CTRL2 PAND2X1_69/A 0.03fF
C44622 PAND2X1_60/B POR2X1_318/A 0.08fF
C44623 POR2X1_532/A POR2X1_854/B 0.05fF
C44624 POR2X1_532/A POR2X1_710/B 0.01fF
C44625 PAND2X1_841/O POR2X1_271/A 0.03fF
C44626 POR2X1_596/A PAND2X1_765/CTRL 0.01fF
C44627 POR2X1_242/CTRL2 PAND2X1_52/B 0.02fF
C44628 PAND2X1_651/Y PAND2X1_861/CTRL 0.00fF
C44629 POR2X1_245/O POR2X1_245/Y 0.03fF
C44630 POR2X1_178/CTRL2 PAND2X1_348/A 0.03fF
C44631 PAND2X1_568/B PAND2X1_578/CTRL2 0.02fF
C44632 PAND2X1_23/Y POR2X1_359/B 0.03fF
C44633 POR2X1_543/A POR2X1_736/A 0.05fF
C44634 POR2X1_366/Y POR2X1_703/CTRL 0.06fF
C44635 POR2X1_614/A PAND2X1_813/O 0.17fF
C44636 PAND2X1_631/A POR2X1_13/A 0.07fF
C44637 POR2X1_343/Y POR2X1_814/B 0.05fF
C44638 POR2X1_128/O POR2X1_540/Y 0.30fF
C44639 POR2X1_848/A POR2X1_9/Y 0.78fF
C44640 POR2X1_95/O POR2X1_51/A 0.01fF
C44641 POR2X1_408/Y PAND2X1_63/B 0.05fF
C44642 POR2X1_119/Y POR2X1_372/Y 0.03fF
C44643 PAND2X1_696/CTRL POR2X1_502/A 0.06fF
C44644 POR2X1_96/Y PAND2X1_35/Y 0.03fF
C44645 POR2X1_184/Y POR2X1_129/Y 0.05fF
C44646 POR2X1_347/O PAND2X1_57/B 0.01fF
C44647 PAND2X1_716/B PAND2X1_302/CTRL2 0.01fF
C44648 PAND2X1_350/a_56_28# POR2X1_7/A 0.00fF
C44649 PAND2X1_48/B POR2X1_349/O 0.01fF
C44650 POR2X1_322/a_16_28# POR2X1_373/Y 0.02fF
C44651 POR2X1_7/B PAND2X1_352/B 0.01fF
C44652 PAND2X1_651/Y POR2X1_129/Y 0.05fF
C44653 PAND2X1_107/a_56_28# POR2X1_532/A 0.00fF
C44654 POR2X1_496/CTRL2 POR2X1_20/B 0.03fF
C44655 POR2X1_114/B POR2X1_737/A 0.04fF
C44656 PAND2X1_229/O PAND2X1_72/A 0.17fF
C44657 PAND2X1_793/Y PAND2X1_860/O 0.02fF
C44658 POR2X1_368/Y POR2X1_109/Y 0.02fF
C44659 POR2X1_119/Y POR2X1_519/Y 0.44fF
C44660 PAND2X1_658/B PAND2X1_185/CTRL2 0.09fF
C44661 PAND2X1_150/CTRL POR2X1_186/B 0.01fF
C44662 POR2X1_119/Y POR2X1_416/Y 0.00fF
C44663 PAND2X1_425/Y POR2X1_635/A 0.01fF
C44664 POR2X1_293/Y PAND2X1_860/a_76_28# 0.01fF
C44665 PAND2X1_865/Y PAND2X1_798/B 0.00fF
C44666 POR2X1_257/A PAND2X1_247/O 0.02fF
C44667 PAND2X1_290/CTRL2 PAND2X1_55/Y 0.03fF
C44668 POR2X1_574/Y PAND2X1_60/B 0.03fF
C44669 POR2X1_779/O POR2X1_513/B 0.02fF
C44670 POR2X1_773/B POR2X1_276/Y 0.30fF
C44671 PAND2X1_47/B D_INPUT_7 1.19fF
C44672 POR2X1_845/A POR2X1_532/A 0.33fF
C44673 POR2X1_728/B POR2X1_728/A 0.02fF
C44674 PAND2X1_39/B POR2X1_624/Y 0.07fF
C44675 INPUT_1 PAND2X1_632/O 0.01fF
C44676 POR2X1_431/CTRL2 POR2X1_67/A 0.12fF
C44677 PAND2X1_55/Y POR2X1_632/Y 0.03fF
C44678 POR2X1_649/a_16_28# POR2X1_643/Y 0.03fF
C44679 POR2X1_186/B POR2X1_128/B 0.00fF
C44680 POR2X1_205/A POR2X1_294/A 0.72fF
C44681 POR2X1_66/B POR2X1_846/A 0.03fF
C44682 POR2X1_96/A POR2X1_759/CTRL2 0.03fF
C44683 POR2X1_9/Y POR2X1_27/Y 0.01fF
C44684 POR2X1_411/A POR2X1_37/Y 0.08fF
C44685 POR2X1_863/A POR2X1_480/A 0.07fF
C44686 POR2X1_81/A POR2X1_816/A 0.03fF
C44687 POR2X1_190/Y PAND2X1_72/A 0.01fF
C44688 PAND2X1_57/B POR2X1_717/B 0.03fF
C44689 POR2X1_8/Y POR2X1_16/A 0.02fF
C44690 PAND2X1_860/A PAND2X1_787/Y 0.05fF
C44691 POR2X1_44/CTRL2 PAND2X1_635/Y 0.01fF
C44692 PAND2X1_736/A POR2X1_416/B 0.19fF
C44693 POR2X1_599/A PAND2X1_198/O 0.02fF
C44694 PAND2X1_865/CTRL2 PAND2X1_862/Y 0.03fF
C44695 POR2X1_66/a_16_28# POR2X1_66/A 0.10fF
C44696 POR2X1_83/B POR2X1_431/O 0.18fF
C44697 PAND2X1_319/B PAND2X1_352/Y 0.06fF
C44698 POR2X1_416/B POR2X1_395/a_16_28# 0.01fF
C44699 POR2X1_9/Y PAND2X1_340/CTRL2 0.04fF
C44700 PAND2X1_55/Y PAND2X1_52/B 0.12fF
C44701 POR2X1_158/Y PAND2X1_725/A 1.43fF
C44702 POR2X1_655/Y POR2X1_814/A 0.24fF
C44703 POR2X1_54/Y POR2X1_48/A 0.14fF
C44704 POR2X1_191/B POR2X1_444/Y 0.01fF
C44705 POR2X1_329/A PAND2X1_361/a_76_28# 0.03fF
C44706 POR2X1_13/A PAND2X1_193/Y 0.78fF
C44707 INPUT_3 POR2X1_669/B 0.05fF
C44708 POR2X1_452/CTRL2 POR2X1_121/B 0.05fF
C44709 POR2X1_633/A POR2X1_633/a_56_344# 0.00fF
C44710 POR2X1_16/A POR2X1_385/Y 0.10fF
C44711 POR2X1_312/m4_208_n4# POR2X1_77/Y 0.12fF
C44712 POR2X1_153/Y PAND2X1_123/Y 0.09fF
C44713 POR2X1_490/Y PAND2X1_576/B 0.04fF
C44714 PAND2X1_787/A POR2X1_39/B 0.03fF
C44715 PAND2X1_159/CTRL2 PAND2X1_9/Y 0.03fF
C44716 POR2X1_862/A POR2X1_66/A 0.04fF
C44717 POR2X1_65/A POR2X1_667/a_16_28# 0.02fF
C44718 POR2X1_71/CTRL POR2X1_62/Y 0.01fF
C44719 POR2X1_814/B POR2X1_240/A 0.03fF
C44720 POR2X1_428/Y POR2X1_669/B 0.06fF
C44721 PAND2X1_72/A POR2X1_702/A 0.06fF
C44722 POR2X1_102/Y PAND2X1_796/B 0.05fF
C44723 POR2X1_77/Y POR2X1_142/Y 14.50fF
C44724 POR2X1_113/A POR2X1_113/B 0.00fF
C44725 POR2X1_359/CTRL2 POR2X1_363/A 0.01fF
C44726 POR2X1_804/A POR2X1_715/O 0.00fF
C44727 POR2X1_143/CTRL POR2X1_9/Y 0.06fF
C44728 POR2X1_116/A POR2X1_269/Y 0.00fF
C44729 PAND2X1_454/B POR2X1_102/Y 0.06fF
C44730 INPUT_1 POR2X1_585/CTRL2 0.01fF
C44731 PAND2X1_205/A D_INPUT_0 0.03fF
C44732 PAND2X1_717/A POR2X1_272/Y 0.03fF
C44733 PAND2X1_20/A POR2X1_624/Y 0.06fF
C44734 POR2X1_632/B POR2X1_632/CTRL2 0.01fF
C44735 POR2X1_523/A POR2X1_523/a_16_28# 0.03fF
C44736 POR2X1_783/Y PAND2X1_52/B 0.04fF
C44737 POR2X1_499/A PAND2X1_41/B 0.03fF
C44738 PAND2X1_26/O PAND2X1_72/A 0.01fF
C44739 POR2X1_630/B VDD 0.02fF
C44740 POR2X1_814/A PAND2X1_257/CTRL2 0.06fF
C44741 PAND2X1_832/CTRL POR2X1_411/B 0.01fF
C44742 PAND2X1_23/Y PAND2X1_438/CTRL 0.01fF
C44743 PAND2X1_41/CTRL PAND2X1_41/B 0.01fF
C44744 POR2X1_567/A POR2X1_703/CTRL 0.11fF
C44745 POR2X1_502/A POR2X1_848/a_16_28# 0.00fF
C44746 POR2X1_37/Y POR2X1_32/A 0.27fF
C44747 POR2X1_467/Y POR2X1_260/B 0.03fF
C44748 POR2X1_23/Y POR2X1_102/Y 0.19fF
C44749 PAND2X1_73/Y POR2X1_66/A 0.45fF
C44750 POR2X1_48/A PAND2X1_732/O 0.01fF
C44751 POR2X1_20/B PAND2X1_721/a_56_28# 0.00fF
C44752 POR2X1_71/Y POR2X1_329/A 0.16fF
C44753 POR2X1_119/Y PAND2X1_858/a_76_28# 0.03fF
C44754 POR2X1_814/B POR2X1_624/Y 0.03fF
C44755 POR2X1_13/A POR2X1_669/Y 0.74fF
C44756 POR2X1_411/B PAND2X1_719/CTRL2 0.01fF
C44757 POR2X1_257/A POR2X1_697/CTRL2 0.01fF
C44758 POR2X1_841/B POR2X1_302/B 0.03fF
C44759 POR2X1_20/B VDD 5.87fF
C44760 POR2X1_456/B POR2X1_715/CTRL2 0.02fF
C44761 POR2X1_316/a_16_28# POR2X1_81/A 0.01fF
C44762 POR2X1_65/A PAND2X1_404/Y 0.02fF
C44763 POR2X1_202/A POR2X1_402/CTRL 0.04fF
C44764 POR2X1_864/A POR2X1_220/Y 0.03fF
C44765 PAND2X1_9/Y PAND2X1_8/Y 5.13fF
C44766 POR2X1_83/B POR2X1_667/Y 0.15fF
C44767 POR2X1_838/B POR2X1_296/B 0.01fF
C44768 POR2X1_411/A POR2X1_293/Y 0.12fF
C44769 PAND2X1_242/Y PAND2X1_349/A 0.05fF
C44770 POR2X1_129/Y PAND2X1_858/B 0.01fF
C44771 POR2X1_624/Y POR2X1_325/A 0.07fF
C44772 POR2X1_696/CTRL2 POR2X1_32/A 0.03fF
C44773 POR2X1_805/CTRL POR2X1_805/B 0.01fF
C44774 POR2X1_567/B POR2X1_509/B 0.05fF
C44775 POR2X1_528/Y POR2X1_386/Y 0.19fF
C44776 POR2X1_270/Y POR2X1_543/A 0.03fF
C44777 POR2X1_333/Y PAND2X1_52/B 0.03fF
C44778 PAND2X1_230/a_16_344# POR2X1_78/A 0.00fF
C44779 PAND2X1_797/Y PAND2X1_326/B 0.03fF
C44780 POR2X1_99/Y POR2X1_243/Y 0.02fF
C44781 PAND2X1_865/Y POR2X1_184/O 0.00fF
C44782 POR2X1_113/A POR2X1_768/A 0.01fF
C44783 POR2X1_4/Y POR2X1_39/B 0.03fF
C44784 POR2X1_16/A POR2X1_91/CTRL2 0.01fF
C44785 PAND2X1_288/CTRL POR2X1_7/B 0.09fF
C44786 PAND2X1_281/CTRL PAND2X1_52/B 0.01fF
C44787 POR2X1_78/B POR2X1_222/a_16_28# 0.09fF
C44788 POR2X1_49/Y PAND2X1_796/O 0.12fF
C44789 POR2X1_416/B POR2X1_7/Y 0.02fF
C44790 POR2X1_482/Y POR2X1_60/A 0.14fF
C44791 POR2X1_60/A PAND2X1_360/O 0.02fF
C44792 POR2X1_60/A POR2X1_251/O 0.01fF
C44793 POR2X1_591/A PAND2X1_718/Y 0.02fF
C44794 PAND2X1_447/CTRL POR2X1_90/Y 0.01fF
C44795 POR2X1_433/Y POR2X1_271/B 0.01fF
C44796 POR2X1_590/A POR2X1_61/Y 0.02fF
C44797 PAND2X1_222/A PAND2X1_592/Y 0.00fF
C44798 PAND2X1_48/A POR2X1_343/B 0.01fF
C44799 POR2X1_16/A POR2X1_16/a_76_344# 0.01fF
C44800 PAND2X1_90/A POR2X1_243/B 0.30fF
C44801 PAND2X1_485/CTRL PAND2X1_57/B 0.02fF
C44802 POR2X1_43/B POR2X1_442/CTRL 0.01fF
C44803 POR2X1_116/A POR2X1_513/Y 0.03fF
C44804 POR2X1_43/B POR2X1_424/Y 0.12fF
C44805 PAND2X1_249/a_16_344# PAND2X1_733/A 0.02fF
C44806 POR2X1_308/O POR2X1_660/Y 0.02fF
C44807 POR2X1_807/A POR2X1_811/B 0.01fF
C44808 PAND2X1_97/CTRL POR2X1_293/Y 0.04fF
C44809 POR2X1_48/A POR2X1_277/CTRL2 0.01fF
C44810 POR2X1_63/Y PAND2X1_734/CTRL 0.01fF
C44811 POR2X1_65/A POR2X1_283/Y 0.01fF
C44812 POR2X1_334/B POR2X1_473/a_76_344# 0.10fF
C44813 POR2X1_60/A POR2X1_106/Y 0.03fF
C44814 PAND2X1_215/a_76_28# PAND2X1_205/Y 0.05fF
C44815 POR2X1_857/CTRL2 VDD -0.00fF
C44816 POR2X1_33/CTRL VDD 0.00fF
C44817 POR2X1_32/A PAND2X1_151/CTRL2 0.01fF
C44818 POR2X1_37/Y PAND2X1_35/Y 0.04fF
C44819 POR2X1_76/A POR2X1_130/Y 0.01fF
C44820 POR2X1_102/Y PAND2X1_558/O 0.05fF
C44821 POR2X1_20/B PAND2X1_344/CTRL2 0.03fF
C44822 POR2X1_41/B POR2X1_409/B 0.03fF
C44823 PAND2X1_850/Y PAND2X1_332/Y 0.07fF
C44824 POR2X1_750/B POR2X1_720/A 0.03fF
C44825 POR2X1_43/B POR2X1_273/O 0.01fF
C44826 POR2X1_96/A POR2X1_496/Y 0.07fF
C44827 POR2X1_614/A POR2X1_635/A 0.01fF
C44828 POR2X1_356/A PAND2X1_237/a_76_28# 0.03fF
C44829 POR2X1_860/CTRL POR2X1_814/A 0.00fF
C44830 PAND2X1_806/O POR2X1_42/Y 0.03fF
C44831 POR2X1_65/A POR2X1_295/a_76_344# 0.01fF
C44832 POR2X1_663/B POR2X1_724/A 0.03fF
C44833 POR2X1_60/A PAND2X1_580/B 0.03fF
C44834 POR2X1_66/B POR2X1_461/B 0.00fF
C44835 PAND2X1_614/CTRL POR2X1_5/Y 0.01fF
C44836 POR2X1_72/B POR2X1_5/Y 1.34fF
C44837 PAND2X1_289/O POR2X1_210/Y 0.02fF
C44838 PAND2X1_289/CTRL POR2X1_220/A 0.00fF
C44839 POR2X1_647/B PAND2X1_96/B 0.68fF
C44840 POR2X1_674/O PAND2X1_742/B 0.01fF
C44841 POR2X1_264/CTRL2 INPUT_0 0.06fF
C44842 POR2X1_717/a_16_28# POR2X1_499/A 0.03fF
C44843 POR2X1_52/A POR2X1_626/m4_208_n4# 0.12fF
C44844 POR2X1_116/A POR2X1_366/A 0.02fF
C44845 POR2X1_66/A PAND2X1_144/CTRL 0.01fF
C44846 POR2X1_270/CTRL2 POR2X1_445/A 0.03fF
C44847 POR2X1_639/A POR2X1_639/a_16_28# 0.01fF
C44848 PAND2X1_463/CTRL2 PAND2X1_460/Y 0.01fF
C44849 POR2X1_32/A POR2X1_293/Y 0.05fF
C44850 POR2X1_257/A PAND2X1_213/Y 0.01fF
C44851 POR2X1_300/O D_INPUT_0 0.01fF
C44852 POR2X1_656/CTRL POR2X1_733/A 0.15fF
C44853 POR2X1_417/Y PAND2X1_151/CTRL2 0.01fF
C44854 POR2X1_260/B PAND2X1_743/O 0.02fF
C44855 PAND2X1_793/Y POR2X1_83/B 0.03fF
C44856 POR2X1_722/B POR2X1_296/B 0.03fF
C44857 PAND2X1_477/B PAND2X1_477/O 0.00fF
C44858 POR2X1_687/Y POR2X1_452/Y 0.01fF
C44859 PAND2X1_845/CTRL POR2X1_23/Y 0.01fF
C44860 POR2X1_296/B POR2X1_294/B 3.19fF
C44861 PAND2X1_848/A POR2X1_669/B 0.12fF
C44862 PAND2X1_485/CTRL2 PAND2X1_69/A 0.03fF
C44863 POR2X1_862/A POR2X1_532/A 0.22fF
C44864 POR2X1_16/A POR2X1_679/CTRL 0.25fF
C44865 INPUT_0 POR2X1_734/A 0.10fF
C44866 PAND2X1_512/CTRL2 POR2X1_7/B 0.00fF
C44867 PAND2X1_319/B POR2X1_298/CTRL 0.01fF
C44868 POR2X1_718/a_16_28# POR2X1_718/A 0.02fF
C44869 POR2X1_814/A POR2X1_768/Y 0.01fF
C44870 POR2X1_66/B PAND2X1_385/CTRL2 0.04fF
C44871 PAND2X1_73/Y POR2X1_222/Y 0.03fF
C44872 PAND2X1_20/A POR2X1_785/A 0.10fF
C44873 POR2X1_76/A POR2X1_228/Y 0.03fF
C44874 INPUT_0 POR2X1_250/A 0.03fF
C44875 PAND2X1_651/Y POR2X1_37/Y 0.12fF
C44876 POR2X1_685/A POR2X1_676/CTRL 0.01fF
C44877 POR2X1_130/A POR2X1_267/B 0.07fF
C44878 POR2X1_790/A PAND2X1_381/Y 0.01fF
C44879 POR2X1_590/A POR2X1_35/Y 0.12fF
C44880 POR2X1_68/A POR2X1_202/B 0.00fF
C44881 POR2X1_224/O POR2X1_226/Y 0.00fF
C44882 POR2X1_40/Y POR2X1_7/B 0.16fF
C44883 POR2X1_78/B POR2X1_786/CTRL 0.03fF
C44884 POR2X1_417/Y POR2X1_293/Y 0.08fF
C44885 POR2X1_814/B PAND2X1_183/CTRL2 0.01fF
C44886 POR2X1_857/O POR2X1_795/B 0.01fF
C44887 PAND2X1_204/O PAND2X1_84/Y 0.00fF
C44888 POR2X1_198/B POR2X1_201/O 0.01fF
C44889 PAND2X1_661/Y POR2X1_681/Y 0.03fF
C44890 PAND2X1_755/CTRL PAND2X1_90/Y 0.00fF
C44891 PAND2X1_23/Y POR2X1_330/Y 0.18fF
C44892 POR2X1_12/O INPUT_4 0.03fF
C44893 PAND2X1_236/CTRL PAND2X1_8/Y 0.01fF
C44894 PAND2X1_484/O POR2X1_705/B 0.00fF
C44895 POR2X1_262/Y POR2X1_394/A 0.01fF
C44896 POR2X1_407/A POR2X1_811/B 0.03fF
C44897 INPUT_0 POR2X1_372/A 0.06fF
C44898 POR2X1_60/A POR2X1_406/A 0.01fF
C44899 PAND2X1_20/A POR2X1_139/CTRL 0.01fF
C44900 POR2X1_60/A PAND2X1_337/A 0.23fF
C44901 POR2X1_341/A POR2X1_244/Y 0.07fF
C44902 PAND2X1_836/O POR2X1_102/Y 0.02fF
C44903 PAND2X1_119/O PAND2X1_73/Y 0.01fF
C44904 POR2X1_43/B POR2X1_748/A 0.03fF
C44905 PAND2X1_73/Y POR2X1_532/A 1.09fF
C44906 POR2X1_502/A PAND2X1_589/a_76_28# 0.01fF
C44907 PAND2X1_48/B PAND2X1_387/O 0.01fF
C44908 POR2X1_447/B POR2X1_66/CTRL 0.08fF
C44909 POR2X1_538/CTRL2 POR2X1_814/B 0.03fF
C44910 POR2X1_114/B POR2X1_302/B 0.00fF
C44911 POR2X1_302/A PAND2X1_299/O 0.14fF
C44912 POR2X1_57/A PAND2X1_296/CTRL 0.01fF
C44913 POR2X1_548/B POR2X1_5/Y 0.10fF
C44914 POR2X1_118/Y PAND2X1_123/O 0.00fF
C44915 POR2X1_317/CTRL2 PAND2X1_90/Y 0.03fF
C44916 PAND2X1_752/a_76_28# PAND2X1_32/B 0.02fF
C44917 PAND2X1_39/B POR2X1_186/B 0.03fF
C44918 PAND2X1_640/B PAND2X1_559/O 0.03fF
C44919 POR2X1_558/B POR2X1_101/Y 0.12fF
C44920 POR2X1_220/B POR2X1_854/B 0.03fF
C44921 POR2X1_49/Y POR2X1_528/O 0.03fF
C44922 POR2X1_296/B PAND2X1_111/B 0.04fF
C44923 PAND2X1_140/A POR2X1_127/a_56_344# 0.00fF
C44924 POR2X1_23/Y PAND2X1_160/O 0.03fF
C44925 POR2X1_32/A POR2X1_408/Y 0.08fF
C44926 POR2X1_496/Y POR2X1_7/A 0.23fF
C44927 POR2X1_686/a_16_28# PAND2X1_73/Y 0.03fF
C44928 POR2X1_57/A PAND2X1_719/Y 0.62fF
C44929 PAND2X1_793/Y PAND2X1_795/B 0.03fF
C44930 POR2X1_78/B POR2X1_832/B 0.03fF
C44931 POR2X1_294/B POR2X1_547/B 0.05fF
C44932 POR2X1_62/Y POR2X1_54/Y 0.05fF
C44933 POR2X1_68/A POR2X1_866/B 0.12fF
C44934 POR2X1_672/CTRL2 POR2X1_5/Y 0.02fF
C44935 POR2X1_65/A PAND2X1_565/A 0.01fF
C44936 PAND2X1_865/m4_208_n4# POR2X1_23/Y 0.07fF
C44937 POR2X1_93/A PAND2X1_390/Y 0.02fF
C44938 PAND2X1_35/Y POR2X1_293/Y 0.03fF
C44939 PAND2X1_41/B POR2X1_206/CTRL 0.09fF
C44940 POR2X1_264/Y VDD 0.81fF
C44941 POR2X1_60/A PAND2X1_349/A 0.07fF
C44942 PAND2X1_853/CTRL2 VDD -0.00fF
C44943 POR2X1_60/A PAND2X1_63/B 0.03fF
C44944 PAND2X1_390/Y POR2X1_91/Y 0.03fF
C44945 POR2X1_750/B POR2X1_318/A 0.10fF
C44946 PAND2X1_658/B INPUT_0 0.10fF
C44947 POR2X1_274/Y POR2X1_573/A 0.01fF
C44948 PAND2X1_499/Y POR2X1_816/A 0.05fF
C44949 POR2X1_476/A POR2X1_768/a_16_28# 0.03fF
C44950 POR2X1_49/Y PAND2X1_213/Y 0.03fF
C44951 POR2X1_60/A PAND2X1_114/B 0.03fF
C44952 POR2X1_775/A POR2X1_192/Y 0.03fF
C44953 POR2X1_46/a_76_344# PAND2X1_338/B 0.01fF
C44954 PAND2X1_228/CTRL2 PAND2X1_364/B 0.03fF
C44955 POR2X1_96/A PAND2X1_514/Y 0.03fF
C44956 POR2X1_102/Y POR2X1_530/CTRL 0.01fF
C44957 POR2X1_485/CTRL POR2X1_73/Y 0.01fF
C44958 PAND2X1_61/Y PAND2X1_560/CTRL 0.01fF
C44959 PAND2X1_80/CTRL D_INPUT_1 0.06fF
C44960 POR2X1_750/O POR2X1_720/A 0.01fF
C44961 POR2X1_193/A POR2X1_795/O 0.02fF
C44962 PAND2X1_424/CTRL2 POR2X1_480/A 0.02fF
C44963 POR2X1_68/A POR2X1_502/A 0.14fF
C44964 POR2X1_786/Y INPUT_0 0.46fF
C44965 PAND2X1_613/O POR2X1_4/Y 0.00fF
C44966 POR2X1_403/O PAND2X1_60/B 0.01fF
C44967 PAND2X1_48/B POR2X1_477/A 0.04fF
C44968 PAND2X1_213/B PAND2X1_162/O 0.02fF
C44969 POR2X1_178/Y POR2X1_251/A 0.00fF
C44970 POR2X1_7/B POR2X1_587/Y 0.00fF
C44971 PAND2X1_93/m4_208_n4# PAND2X1_57/B 0.15fF
C44972 POR2X1_130/CTRL POR2X1_66/B 0.01fF
C44973 POR2X1_558/O POR2X1_294/B 0.05fF
C44974 POR2X1_851/O POR2X1_590/A 0.01fF
C44975 POR2X1_857/B POR2X1_35/Y 0.03fF
C44976 POR2X1_41/B POR2X1_229/CTRL2 0.00fF
C44977 POR2X1_74/Y POR2X1_23/Y 0.01fF
C44978 POR2X1_68/A POR2X1_464/Y 0.00fF
C44979 POR2X1_407/A POR2X1_783/B 0.01fF
C44980 POR2X1_48/A POR2X1_4/Y 0.03fF
C44981 PAND2X1_36/O PAND2X1_18/B 0.05fF
C44982 POR2X1_365/Y POR2X1_357/Y 0.21fF
C44983 POR2X1_547/B PAND2X1_111/B 0.01fF
C44984 PAND2X1_20/A POR2X1_186/B 0.10fF
C44985 POR2X1_220/Y POR2X1_194/O 0.06fF
C44986 PAND2X1_849/B PAND2X1_61/Y 0.00fF
C44987 PAND2X1_651/Y POR2X1_293/Y 0.19fF
C44988 POR2X1_76/Y POR2X1_541/O 0.01fF
C44989 POR2X1_502/A POR2X1_565/m4_208_n4# 0.06fF
C44990 POR2X1_52/A PAND2X1_209/A 0.00fF
C44991 POR2X1_416/B POR2X1_257/A 27.69fF
C44992 POR2X1_369/a_56_344# POR2X1_60/A 0.03fF
C44993 POR2X1_45/Y POR2X1_599/A 0.01fF
C44994 POR2X1_214/a_16_28# POR2X1_208/Y 0.05fF
C44995 PAND2X1_811/Y VDD 0.00fF
C44996 PAND2X1_386/CTRL2 POR2X1_260/A 0.01fF
C44997 PAND2X1_200/O PAND2X1_200/B 0.00fF
C44998 POR2X1_852/O POR2X1_854/B 0.04fF
C44999 POR2X1_614/A POR2X1_795/O 0.01fF
C45000 POR2X1_134/Y POR2X1_7/B 0.10fF
C45001 POR2X1_390/B POR2X1_105/Y 0.03fF
C45002 PAND2X1_131/O PAND2X1_60/B 0.16fF
C45003 PAND2X1_94/A PAND2X1_55/O 0.04fF
C45004 PAND2X1_486/CTRL2 POR2X1_526/Y 0.03fF
C45005 PAND2X1_182/O POR2X1_55/Y 0.04fF
C45006 PAND2X1_214/A PAND2X1_123/Y 0.03fF
C45007 PAND2X1_631/A POR2X1_482/a_16_28# 0.03fF
C45008 PAND2X1_702/CTRL POR2X1_42/Y 0.02fF
C45009 POR2X1_347/A POR2X1_402/CTRL 0.01fF
C45010 POR2X1_149/Y POR2X1_209/A 0.04fF
C45011 POR2X1_174/B POR2X1_447/B 0.03fF
C45012 PAND2X1_95/B POR2X1_407/Y 0.00fF
C45013 POR2X1_156/B POR2X1_803/A 0.01fF
C45014 POR2X1_407/A POR2X1_114/CTRL 0.00fF
C45015 POR2X1_264/Y PAND2X1_32/B 0.05fF
C45016 POR2X1_721/a_16_28# POR2X1_720/Y 0.03fF
C45017 POR2X1_809/A POR2X1_330/Y 0.05fF
C45018 POR2X1_308/O POR2X1_308/B 0.01fF
C45019 POR2X1_57/A POR2X1_42/Y 1.10fF
C45020 POR2X1_685/a_16_28# POR2X1_687/A 0.02fF
C45021 PAND2X1_632/CTRL VDD -0.00fF
C45022 POR2X1_55/Y POR2X1_172/Y 0.13fF
C45023 POR2X1_814/B POR2X1_186/B 0.03fF
C45024 D_GATE_662 POR2X1_544/CTRL 0.03fF
C45025 PAND2X1_275/CTRL2 PAND2X1_60/B 0.03fF
C45026 POR2X1_68/A PAND2X1_747/CTRL2 0.02fF
C45027 POR2X1_220/Y POR2X1_553/A 0.03fF
C45028 POR2X1_640/Y POR2X1_113/B 0.02fF
C45029 POR2X1_509/A POR2X1_532/A 0.03fF
C45030 POR2X1_523/Y POR2X1_844/CTRL2 0.01fF
C45031 PAND2X1_715/B VDD 0.23fF
C45032 PAND2X1_864/O GATE_741 0.01fF
C45033 POR2X1_390/B POR2X1_337/CTRL2 0.00fF
C45034 POR2X1_409/B POR2X1_77/Y 0.07fF
C45035 POR2X1_48/CTRL POR2X1_153/Y 0.06fF
C45036 POR2X1_57/A POR2X1_309/Y 6.61fF
C45037 PAND2X1_716/a_16_344# POR2X1_73/Y 0.01fF
C45038 PAND2X1_90/Y PAND2X1_384/O 0.02fF
C45039 PAND2X1_303/Y VDD 0.13fF
C45040 POR2X1_407/Y PAND2X1_743/O 0.02fF
C45041 PAND2X1_662/Y PAND2X1_660/B 0.01fF
C45042 PAND2X1_364/B POR2X1_385/O 0.04fF
C45043 POR2X1_541/CTRL2 PAND2X1_32/B 0.01fF
C45044 POR2X1_532/A POR2X1_631/B 0.03fF
C45045 POR2X1_60/Y PAND2X1_338/CTRL 0.01fF
C45046 POR2X1_68/A POR2X1_140/m4_208_n4# 0.06fF
C45047 PAND2X1_749/a_16_344# PAND2X1_8/Y 0.02fF
C45048 POR2X1_584/Y POR2X1_42/Y 0.03fF
C45049 PAND2X1_386/a_76_28# PAND2X1_48/A 0.03fF
C45050 PAND2X1_636/m4_208_n4# POR2X1_260/A 0.09fF
C45051 POR2X1_110/O POR2X1_5/Y 0.02fF
C45052 POR2X1_407/Y POR2X1_770/a_56_344# 0.00fF
C45053 POR2X1_204/CTRL PAND2X1_63/B 0.01fF
C45054 POR2X1_356/A POR2X1_782/CTRL2 0.04fF
C45055 POR2X1_555/A POR2X1_447/B 0.07fF
C45056 POR2X1_278/Y PAND2X1_853/B 0.07fF
C45057 POR2X1_93/CTRL2 POR2X1_283/A 0.01fF
C45058 PAND2X1_651/Y POR2X1_408/Y 0.05fF
C45059 POR2X1_356/A POR2X1_703/Y 0.05fF
C45060 POR2X1_90/Y POR2X1_387/Y 0.07fF
C45061 PAND2X1_675/A PAND2X1_181/a_16_344# 0.01fF
C45062 POR2X1_519/CTRL POR2X1_43/B 0.01fF
C45063 POR2X1_68/A POR2X1_799/CTRL 0.06fF
C45064 POR2X1_3/A D_INPUT_6 0.72fF
C45065 POR2X1_740/Y POR2X1_675/Y 0.03fF
C45066 POR2X1_247/a_16_28# POR2X1_260/A 0.02fF
C45067 POR2X1_174/A PAND2X1_52/B 0.03fF
C45068 POR2X1_264/Y POR2X1_673/Y 0.03fF
C45069 POR2X1_502/Y VDD 0.15fF
C45070 PAND2X1_659/Y POR2X1_821/CTRL2 0.11fF
C45071 PAND2X1_48/O PAND2X1_48/A 0.01fF
C45072 POR2X1_111/O POR2X1_387/Y 0.06fF
C45073 POR2X1_461/Y POR2X1_848/CTRL 0.01fF
C45074 POR2X1_790/B POR2X1_789/B 0.03fF
C45075 POR2X1_334/A POR2X1_404/Y 0.05fF
C45076 POR2X1_857/B POR2X1_227/CTRL2 0.03fF
C45077 PAND2X1_812/A VDD 0.18fF
C45078 POR2X1_96/A POR2X1_75/Y 0.07fF
C45079 PAND2X1_94/A PAND2X1_49/O 0.03fF
C45080 POR2X1_330/Y POR2X1_711/Y 0.10fF
C45081 POR2X1_114/Y PAND2X1_48/A 0.01fF
C45082 POR2X1_405/Y POR2X1_737/A 0.02fF
C45083 PAND2X1_150/O PAND2X1_63/B 0.01fF
C45084 PAND2X1_23/Y POR2X1_715/A 0.15fF
C45085 POR2X1_23/Y POR2X1_677/Y 0.03fF
C45086 POR2X1_330/Y POR2X1_728/A 0.02fF
C45087 POR2X1_332/Y POR2X1_785/A 0.06fF
C45088 PAND2X1_649/A POR2X1_393/O 0.01fF
C45089 POR2X1_49/Y POR2X1_416/B 0.48fF
C45090 PAND2X1_843/Y PAND2X1_842/Y 0.20fF
C45091 PAND2X1_55/Y POR2X1_722/CTRL2 0.00fF
C45092 POR2X1_16/A PAND2X1_401/m4_208_n4# 0.15fF
C45093 POR2X1_730/Y POR2X1_732/a_16_28# 0.02fF
C45094 POR2X1_294/B POR2X1_342/CTRL 0.01fF
C45095 POR2X1_492/Y VDD 0.14fF
C45096 POR2X1_21/CTRL2 POR2X1_260/A 0.01fF
C45097 PAND2X1_850/Y POR2X1_13/A 0.07fF
C45098 PAND2X1_611/O POR2X1_54/Y 0.01fF
C45099 POR2X1_640/Y POR2X1_768/A 0.03fF
C45100 POR2X1_568/Y POR2X1_162/Y 0.03fF
C45101 PAND2X1_191/a_76_28# POR2X1_385/Y 0.06fF
C45102 POR2X1_189/O VDD 0.00fF
C45103 POR2X1_343/A POR2X1_717/B 0.03fF
C45104 PAND2X1_569/B POR2X1_766/CTRL2 0.01fF
C45105 POR2X1_763/Y POR2X1_524/CTRL2 0.01fF
C45106 POR2X1_20/B PAND2X1_9/Y 0.03fF
C45107 POR2X1_560/a_56_344# POR2X1_294/B 0.00fF
C45108 POR2X1_478/B POR2X1_444/Y 0.03fF
C45109 POR2X1_608/O PAND2X1_56/A 0.01fF
C45110 POR2X1_343/Y VDD 3.45fF
C45111 POR2X1_830/A PAND2X1_72/A 0.01fF
C45112 POR2X1_68/A POR2X1_188/Y 0.05fF
C45113 PAND2X1_127/m4_208_n4# PAND2X1_125/m4_208_n4# 0.13fF
C45114 PAND2X1_349/A PAND2X1_301/CTRL 0.01fF
C45115 POR2X1_86/Y VDD -0.00fF
C45116 PAND2X1_63/Y PAND2X1_48/A 0.04fF
C45117 POR2X1_1/O POR2X1_260/A 0.01fF
C45118 POR2X1_447/a_76_344# POR2X1_186/B 0.00fF
C45119 POR2X1_333/Y POR2X1_350/B 0.95fF
C45120 POR2X1_42/Y POR2X1_589/CTRL 0.01fF
C45121 POR2X1_101/Y POR2X1_362/A 0.10fF
C45122 POR2X1_116/Y POR2X1_276/Y 0.44fF
C45123 POR2X1_711/B PAND2X1_69/A 0.01fF
C45124 PAND2X1_841/B PAND2X1_841/Y 0.04fF
C45125 POR2X1_153/CTRL POR2X1_96/B 0.01fF
C45126 POR2X1_835/B PAND2X1_239/O 0.01fF
C45127 PAND2X1_738/A POR2X1_394/A 0.05fF
C45128 POR2X1_471/O PAND2X1_72/A 0.08fF
C45129 POR2X1_25/Y D_INPUT_6 0.01fF
C45130 POR2X1_52/CTRL POR2X1_599/A 0.01fF
C45131 POR2X1_711/B POR2X1_710/a_16_28# 0.03fF
C45132 POR2X1_43/Y VDD 0.01fF
C45133 POR2X1_293/Y POR2X1_387/CTRL -0.02fF
C45134 POR2X1_416/B PAND2X1_553/B 0.07fF
C45135 PAND2X1_644/CTRL POR2X1_669/B 0.01fF
C45136 POR2X1_113/Y PAND2X1_48/A 0.07fF
C45137 VDD POR2X1_589/Y 0.01fF
C45138 POR2X1_132/CTRL PAND2X1_140/A 0.01fF
C45139 POR2X1_96/A PAND2X1_332/Y 0.96fF
C45140 POR2X1_257/A POR2X1_109/CTRL 0.05fF
C45141 POR2X1_121/O POR2X1_537/Y 0.01fF
C45142 POR2X1_119/Y PAND2X1_344/O 0.02fF
C45143 POR2X1_110/Y POR2X1_387/Y 0.06fF
C45144 POR2X1_119/Y PAND2X1_560/O 0.23fF
C45145 POR2X1_428/CTRL POR2X1_394/A 0.01fF
C45146 POR2X1_55/O POR2X1_624/B 0.14fF
C45147 POR2X1_799/CTRL2 POR2X1_652/A 0.00fF
C45148 PAND2X1_288/a_16_344# PAND2X1_287/Y 0.02fF
C45149 POR2X1_159/a_76_344# POR2X1_9/Y 0.01fF
C45150 PAND2X1_326/CTRL2 PAND2X1_324/Y 0.00fF
C45151 PAND2X1_466/A POR2X1_669/B 0.00fF
C45152 POR2X1_816/A POR2X1_39/B 0.08fF
C45153 POR2X1_533/Y POR2X1_759/Y 0.01fF
C45154 POR2X1_260/B POR2X1_655/A 0.06fF
C45155 D_INPUT_1 POR2X1_39/B 0.03fF
C45156 POR2X1_614/A POR2X1_736/A 0.05fF
C45157 POR2X1_326/A POR2X1_456/B 0.17fF
C45158 PAND2X1_206/B POR2X1_40/Y 0.14fF
C45159 PAND2X1_634/CTRL POR2X1_102/Y 0.01fF
C45160 POR2X1_93/O POR2X1_77/Y 0.01fF
C45161 PAND2X1_48/A POR2X1_260/A 2.81fF
C45162 POR2X1_343/Y PAND2X1_32/B 0.07fF
C45163 POR2X1_16/A POR2X1_767/CTRL 0.01fF
C45164 POR2X1_86/O POR2X1_7/A 0.02fF
C45165 PAND2X1_295/O POR2X1_294/Y 0.00fF
C45166 POR2X1_78/A POR2X1_663/B 0.00fF
C45167 POR2X1_286/B PAND2X1_595/m4_208_n4# 0.01fF
C45168 POR2X1_739/m4_208_n4# POR2X1_738/m4_208_n4# 0.05fF
C45169 POR2X1_332/Y POR2X1_186/B 0.13fF
C45170 POR2X1_698/Y PAND2X1_709/CTRL2 0.03fF
C45171 POR2X1_344/Y POR2X1_359/CTRL 0.00fF
C45172 PAND2X1_275/CTRL POR2X1_76/B 0.01fF
C45173 POR2X1_520/CTRL2 POR2X1_383/Y 0.01fF
C45174 POR2X1_513/A POR2X1_513/a_16_28# 0.06fF
C45175 POR2X1_408/Y POR2X1_387/CTRL 0.01fF
C45176 POR2X1_13/A PAND2X1_99/O 0.02fF
C45177 POR2X1_777/B POR2X1_556/A 0.03fF
C45178 POR2X1_596/A PAND2X1_72/A 0.06fF
C45179 POR2X1_48/A POR2X1_695/Y 0.01fF
C45180 PAND2X1_12/O PAND2X1_11/Y 0.02fF
C45181 POR2X1_702/A POR2X1_579/CTRL 0.01fF
C45182 POR2X1_567/A POR2X1_566/CTRL2 0.03fF
C45183 POR2X1_604/CTRL POR2X1_40/Y 0.01fF
C45184 POR2X1_359/B POR2X1_349/O 0.00fF
C45185 POR2X1_614/A PAND2X1_135/a_76_28# 0.01fF
C45186 POR2X1_65/Y POR2X1_40/Y 0.01fF
C45187 PAND2X1_271/CTRL2 POR2X1_330/Y 0.31fF
C45188 POR2X1_431/a_16_28# POR2X1_236/Y 0.06fF
C45189 PAND2X1_651/Y PAND2X1_242/Y 0.02fF
C45190 PAND2X1_449/CTRL POR2X1_236/Y 0.01fF
C45191 POR2X1_728/A PAND2X1_158/CTRL 0.00fF
C45192 PAND2X1_43/O POR2X1_852/B 0.08fF
C45193 POR2X1_96/CTRL2 POR2X1_77/Y 0.00fF
C45194 POR2X1_89/O POR2X1_60/A 0.02fF
C45195 PAND2X1_65/B POR2X1_556/A 0.08fF
C45196 POR2X1_60/A PAND2X1_97/CTRL 0.01fF
C45197 POR2X1_62/Y POR2X1_4/Y 0.08fF
C45198 POR2X1_530/a_76_344# POR2X1_39/B 0.00fF
C45199 POR2X1_486/a_16_28# PAND2X1_57/B 0.02fF
C45200 PAND2X1_247/CTRL POR2X1_5/Y 0.01fF
C45201 POR2X1_115/CTRL2 POR2X1_554/B 0.03fF
C45202 POR2X1_265/CTRL2 POR2X1_40/Y 0.03fF
C45203 PAND2X1_241/O POR2X1_329/A 0.06fF
C45204 PAND2X1_446/Y POR2X1_511/Y 0.03fF
C45205 PAND2X1_358/O POR2X1_153/Y 0.26fF
C45206 POR2X1_627/O POR2X1_628/Y 0.00fF
C45207 POR2X1_669/B POR2X1_423/O 0.01fF
C45208 POR2X1_471/CTRL2 POR2X1_471/A 0.00fF
C45209 PAND2X1_797/Y POR2X1_373/O 0.08fF
C45210 POR2X1_12/A POR2X1_12/a_16_28# 0.07fF
C45211 POR2X1_150/Y POR2X1_46/Y 0.05fF
C45212 POR2X1_60/A POR2X1_32/A 1.50fF
C45213 POR2X1_703/Y PAND2X1_72/A 0.03fF
C45214 PAND2X1_717/A PAND2X1_717/a_16_344# 0.01fF
C45215 POR2X1_16/A POR2X1_167/Y 0.27fF
C45216 POR2X1_94/A POR2X1_37/Y 0.06fF
C45217 PAND2X1_48/B POR2X1_554/B 0.03fF
C45218 POR2X1_624/Y VDD 2.17fF
C45219 PAND2X1_645/CTRL POR2X1_600/Y 0.01fF
C45220 POR2X1_449/A PAND2X1_72/A 0.04fF
C45221 D_INPUT_0 PAND2X1_558/Y 0.00fF
C45222 POR2X1_257/A PAND2X1_738/Y 0.01fF
C45223 POR2X1_603/O POR2X1_597/A 0.00fF
C45224 POR2X1_502/A POR2X1_709/A 0.03fF
C45225 POR2X1_257/A POR2X1_425/CTRL 0.01fF
C45226 POR2X1_66/A POR2X1_61/Y 0.07fF
C45227 PAND2X1_645/CTRL2 POR2X1_48/A 0.00fF
C45228 POR2X1_687/B POR2X1_452/Y 0.01fF
C45229 PAND2X1_463/CTRL PAND2X1_58/A 0.02fF
C45230 POR2X1_502/A PAND2X1_601/O 0.03fF
C45231 POR2X1_60/A POR2X1_417/Y 0.03fF
C45232 POR2X1_135/Y POR2X1_48/A 0.28fF
C45233 POR2X1_121/B POR2X1_405/O 0.16fF
C45234 PAND2X1_810/O PAND2X1_221/Y 0.01fF
C45235 PAND2X1_200/CTRL POR2X1_72/B 0.01fF
C45236 POR2X1_807/A POR2X1_296/B 0.03fF
C45237 POR2X1_102/Y POR2X1_250/A 0.03fF
C45238 PAND2X1_205/A PAND2X1_735/Y 0.02fF
C45239 POR2X1_474/O POR2X1_777/B 0.02fF
C45240 POR2X1_278/Y POR2X1_23/Y 0.01fF
C45241 POR2X1_624/Y POR2X1_501/CTRL2 0.03fF
C45242 POR2X1_12/A PAND2X1_709/CTRL 0.02fF
C45243 PAND2X1_443/Y PAND2X1_803/A 0.02fF
C45244 POR2X1_491/CTRL POR2X1_72/B 0.01fF
C45245 POR2X1_458/Y PAND2X1_300/CTRL2 0.01fF
C45246 PAND2X1_338/O PAND2X1_333/Y 0.02fF
C45247 POR2X1_566/A POR2X1_567/B 0.46fF
C45248 POR2X1_446/B POR2X1_276/O 0.01fF
C45249 POR2X1_257/A POR2X1_273/Y 0.03fF
C45250 POR2X1_624/Y POR2X1_741/Y 0.07fF
C45251 POR2X1_686/A POR2X1_467/Y 0.09fF
C45252 PAND2X1_55/Y POR2X1_655/A 0.07fF
C45253 PAND2X1_277/O PAND2X1_57/B 0.12fF
C45254 POR2X1_689/A PAND2X1_590/CTRL2 0.01fF
C45255 POR2X1_69/A PAND2X1_340/CTRL2 0.03fF
C45256 PAND2X1_68/m4_208_n4# PAND2X1_340/m4_208_n4# 0.04fF
C45257 PAND2X1_852/B POR2X1_20/B 0.01fF
C45258 PAND2X1_81/B POR2X1_624/Y 0.02fF
C45259 POR2X1_22/A POR2X1_12/A 0.00fF
C45260 POR2X1_270/Y POR2X1_193/A 4.09fF
C45261 PAND2X1_220/Y POR2X1_40/Y 0.03fF
C45262 PAND2X1_39/B POR2X1_208/Y 0.21fF
C45263 PAND2X1_20/A POR2X1_489/a_16_28# 0.03fF
C45264 POR2X1_102/Y POR2X1_372/A 0.05fF
C45265 POR2X1_411/B POR2X1_382/Y 0.02fF
C45266 PAND2X1_6/Y POR2X1_446/B 0.03fF
C45267 POR2X1_41/B PAND2X1_804/a_16_344# 0.01fF
C45268 PAND2X1_7/Y PAND2X1_52/Y 0.29fF
C45269 POR2X1_174/B POR2X1_852/a_16_28# 0.01fF
C45270 POR2X1_807/CTRL POR2X1_294/B 0.01fF
C45271 POR2X1_624/Y PAND2X1_32/B 7.02fF
C45272 POR2X1_343/CTRL2 POR2X1_343/B 0.01fF
C45273 POR2X1_3/A PAND2X1_635/m4_208_n4# 0.01fF
C45274 PAND2X1_814/a_16_344# INPUT_3 0.04fF
C45275 POR2X1_306/CTRL PAND2X1_454/B 0.01fF
C45276 POR2X1_78/A PAND2X1_322/CTRL2 0.04fF
C45277 POR2X1_106/O PAND2X1_553/B 0.03fF
C45278 PAND2X1_116/CTRL2 POR2X1_106/Y 0.01fF
C45279 POR2X1_502/A PAND2X1_58/A 16.81fF
C45280 POR2X1_142/O PAND2X1_738/Y 0.04fF
C45281 POR2X1_96/A POR2X1_674/Y 0.03fF
C45282 POR2X1_786/A PAND2X1_73/Y 0.14fF
C45283 POR2X1_62/CTRL2 POR2X1_29/A 0.08fF
C45284 POR2X1_278/Y PAND2X1_221/O 0.07fF
C45285 POR2X1_60/A PAND2X1_35/Y 0.06fF
C45286 PAND2X1_279/O PAND2X1_57/B 0.17fF
C45287 POR2X1_138/CTRL2 POR2X1_296/B 0.01fF
C45288 POR2X1_43/B POR2X1_263/Y 0.05fF
C45289 POR2X1_290/CTRL POR2X1_236/Y 0.01fF
C45290 PAND2X1_116/CTRL PAND2X1_787/Y 0.29fF
C45291 PAND2X1_699/O POR2X1_260/A 0.02fF
C45292 POR2X1_290/Y POR2X1_102/Y 0.12fF
C45293 POR2X1_614/A POR2X1_270/Y 0.03fF
C45294 POR2X1_66/A POR2X1_35/Y 1.97fF
C45295 INPUT_1 POR2X1_19/CTRL 0.01fF
C45296 POR2X1_48/A POR2X1_816/A 0.03fF
C45297 POR2X1_48/A PAND2X1_569/A 0.03fF
C45298 POR2X1_119/CTRL POR2X1_102/Y 0.01fF
C45299 POR2X1_48/A D_INPUT_1 0.06fF
C45300 PAND2X1_700/CTRL2 PAND2X1_90/Y 0.07fF
C45301 D_INPUT_5 POR2X1_1/CTRL 0.05fF
C45302 PAND2X1_685/CTRL2 POR2X1_60/A 0.01fF
C45303 POR2X1_78/CTRL D_INPUT_0 0.01fF
C45304 POR2X1_602/B POR2X1_722/Y 0.01fF
C45305 POR2X1_49/Y PAND2X1_738/Y 0.03fF
C45306 PAND2X1_456/O VDD 0.00fF
C45307 POR2X1_750/B POR2X1_586/CTRL 0.00fF
C45308 PAND2X1_235/CTRL PAND2X1_55/Y 0.01fF
C45309 POR2X1_76/CTRL2 POR2X1_274/B 0.01fF
C45310 PAND2X1_810/A POR2X1_7/B 0.09fF
C45311 PAND2X1_833/CTRL POR2X1_511/Y 0.02fF
C45312 POR2X1_37/Y PAND2X1_342/CTRL 0.01fF
C45313 INPUT_7 VDD 0.68fF
C45314 POR2X1_271/Y POR2X1_275/O 0.00fF
C45315 POR2X1_102/Y POR2X1_238/Y 1.46fF
C45316 POR2X1_189/Y POR2X1_60/A 0.03fF
C45317 POR2X1_407/A POR2X1_296/B 0.10fF
C45318 POR2X1_102/Y PAND2X1_658/B 0.05fF
C45319 POR2X1_461/Y POR2X1_260/A 0.03fF
C45320 PAND2X1_755/a_76_28# PAND2X1_41/B 0.01fF
C45321 POR2X1_707/A PAND2X1_48/B 0.02fF
C45322 POR2X1_94/A POR2X1_293/Y 0.03fF
C45323 POR2X1_278/Y PAND2X1_740/O 0.12fF
C45324 PAND2X1_843/a_56_28# PAND2X1_738/Y 0.00fF
C45325 POR2X1_121/B PAND2X1_536/O 0.01fF
C45326 POR2X1_675/O POR2X1_732/B 0.28fF
C45327 PAND2X1_863/B PAND2X1_805/A 0.07fF
C45328 POR2X1_330/Y POR2X1_733/A 0.10fF
C45329 POR2X1_60/A POR2X1_184/Y 0.04fF
C45330 PAND2X1_242/a_16_344# POR2X1_60/A 0.01fF
C45331 PAND2X1_6/Y POR2X1_121/B 0.11fF
C45332 POR2X1_808/A PAND2X1_599/CTRL 0.06fF
C45333 POR2X1_78/B POR2X1_130/A 0.07fF
C45334 POR2X1_62/CTRL POR2X1_94/A 0.01fF
C45335 PAND2X1_20/A POR2X1_515/Y 0.01fF
C45336 POR2X1_832/A PAND2X1_591/CTRL 0.03fF
C45337 POR2X1_366/Y POR2X1_186/Y 0.07fF
C45338 POR2X1_186/Y POR2X1_294/B 0.03fF
C45339 PAND2X1_61/Y PAND2X1_523/O 0.01fF
C45340 PAND2X1_96/B POR2X1_202/B 0.04fF
C45341 PAND2X1_436/A PAND2X1_658/B 0.10fF
C45342 POR2X1_254/A POR2X1_341/O 0.01fF
C45343 PAND2X1_579/B VDD 0.37fF
C45344 POR2X1_75/CTRL POR2X1_60/A 0.01fF
C45345 POR2X1_502/A PAND2X1_588/a_76_28# 0.01fF
C45346 POR2X1_48/A PAND2X1_854/A 0.02fF
C45347 POR2X1_346/B POR2X1_629/CTRL2 0.01fF
C45348 POR2X1_78/B POR2X1_566/A 0.13fF
C45349 PAND2X1_651/Y POR2X1_60/A 0.09fF
C45350 POR2X1_509/B POR2X1_340/O 0.03fF
C45351 PAND2X1_63/Y PAND2X1_265/CTRL 0.28fF
C45352 PAND2X1_857/B POR2X1_23/Y 0.03fF
C45353 POR2X1_7/B POR2X1_5/Y 8.12fF
C45354 POR2X1_356/A PAND2X1_90/Y 0.07fF
C45355 PAND2X1_459/Y VDD 0.00fF
C45356 PAND2X1_6/Y POR2X1_630/A 0.03fF
C45357 PAND2X1_804/CTRL POR2X1_283/A 0.01fF
C45358 POR2X1_96/A PAND2X1_474/Y 0.02fF
C45359 POR2X1_123/A POR2X1_66/A 0.03fF
C45360 POR2X1_738/Y VDD 0.10fF
C45361 POR2X1_631/A POR2X1_590/A 0.12fF
C45362 POR2X1_13/Y POR2X1_595/Y 0.01fF
C45363 POR2X1_198/CTRL POR2X1_61/Y 0.01fF
C45364 PAND2X1_805/A PAND2X1_567/O 0.02fF
C45365 POR2X1_69/O PAND2X1_69/A 0.01fF
C45366 PAND2X1_732/CTRL2 PAND2X1_731/A 0.01fF
C45367 PAND2X1_732/O POR2X1_152/Y 0.02fF
C45368 INPUT_4 VDD 0.67fF
C45369 PAND2X1_20/A PAND2X1_79/Y 0.02fF
C45370 POR2X1_502/A POR2X1_435/Y 0.07fF
C45371 PAND2X1_126/CTRL2 POR2X1_29/A 0.12fF
C45372 D_INPUT_0 POR2X1_569/A 0.29fF
C45373 POR2X1_61/Y POR2X1_222/Y 0.07fF
C45374 POR2X1_331/A VDD 0.00fF
C45375 POR2X1_504/Y PAND2X1_631/CTRL2 0.01fF
C45376 POR2X1_71/Y PAND2X1_84/Y 0.10fF
C45377 POR2X1_16/A PAND2X1_776/Y 0.01fF
C45378 POR2X1_96/A POR2X1_13/A 0.15fF
C45379 POR2X1_407/A PAND2X1_679/CTRL2 0.02fF
C45380 POR2X1_68/A PAND2X1_679/CTRL 0.03fF
C45381 PAND2X1_57/B PAND2X1_751/CTRL2 0.18fF
C45382 PAND2X1_254/a_16_344# POR2X1_511/Y 0.02fF
C45383 POR2X1_565/B POR2X1_547/B 0.02fF
C45384 PAND2X1_115/B VDD 0.35fF
C45385 PAND2X1_738/Y PAND2X1_553/B 0.10fF
C45386 POR2X1_218/Y POR2X1_276/Y 0.03fF
C45387 POR2X1_38/Y PAND2X1_733/A 0.23fF
C45388 POR2X1_785/A VDD 0.30fF
C45389 PAND2X1_217/B POR2X1_73/Y 0.03fF
C45390 PAND2X1_41/B PAND2X1_69/A 8.17fF
C45391 POR2X1_481/A POR2X1_55/Y 0.03fF
C45392 PAND2X1_48/B POR2X1_723/CTRL 0.00fF
C45393 POR2X1_329/A PAND2X1_840/Y 0.03fF
C45394 POR2X1_114/B POR2X1_362/B 0.08fF
C45395 PAND2X1_243/B PAND2X1_734/B 0.06fF
C45396 POR2X1_13/CTRL2 POR2X1_13/Y 0.01fF
C45397 POR2X1_46/Y PAND2X1_364/B 0.07fF
C45398 PAND2X1_476/A PAND2X1_267/B 0.00fF
C45399 POR2X1_435/Y POR2X1_532/Y 0.15fF
C45400 PAND2X1_258/CTRL2 POR2X1_186/B 0.03fF
C45401 PAND2X1_658/A VDD 0.09fF
C45402 POR2X1_669/B POR2X1_428/CTRL 0.04fF
C45403 PAND2X1_23/Y POR2X1_332/B 0.04fF
C45404 POR2X1_483/O POR2X1_294/B 0.08fF
C45405 POR2X1_413/A POR2X1_607/Y 0.01fF
C45406 INPUT_1 POR2X1_496/Y 0.14fF
C45407 POR2X1_94/A PAND2X1_521/O 0.05fF
C45408 POR2X1_287/B POR2X1_840/B 0.13fF
C45409 PAND2X1_20/O POR2X1_68/B 0.04fF
C45410 POR2X1_325/A POR2X1_515/Y 0.01fF
C45411 POR2X1_481/O POR2X1_481/Y 0.01fF
C45412 PAND2X1_613/O POR2X1_620/B 0.05fF
C45413 PAND2X1_172/O POR2X1_174/A 0.02fF
C45414 POR2X1_61/Y POR2X1_532/A 1.30fF
C45415 POR2X1_355/B POR2X1_740/Y 0.03fF
C45416 POR2X1_174/CTRL POR2X1_174/A 0.01fF
C45417 PAND2X1_504/O VDD 0.00fF
C45418 POR2X1_32/A PAND2X1_301/CTRL 0.01fF
C45419 POR2X1_463/Y POR2X1_590/A 0.03fF
C45420 POR2X1_78/B POR2X1_844/B 0.04fF
C45421 PAND2X1_65/B PAND2X1_153/CTRL 0.01fF
C45422 PAND2X1_23/Y POR2X1_284/CTRL 0.01fF
C45423 PAND2X1_614/CTRL2 POR2X1_283/A 0.01fF
C45424 POR2X1_476/A POR2X1_557/B 3.53fF
C45425 POR2X1_410/Y PAND2X1_65/B 0.01fF
C45426 PAND2X1_274/O POR2X1_273/Y 0.02fF
C45427 POR2X1_483/A POR2X1_840/B 0.01fF
C45428 POR2X1_237/O POR2X1_90/Y 0.01fF
C45429 POR2X1_130/A PAND2X1_767/CTRL 0.03fF
C45430 POR2X1_383/A POR2X1_405/O 0.04fF
C45431 POR2X1_57/A PAND2X1_319/CTRL 0.01fF
C45432 PAND2X1_436/a_76_28# PAND2X1_508/Y 0.02fF
C45433 POR2X1_542/B POR2X1_325/A 0.00fF
C45434 POR2X1_477/B POR2X1_440/Y 0.00fF
C45435 PAND2X1_349/A PAND2X1_140/O 0.02fF
C45436 POR2X1_496/Y POR2X1_153/Y 0.10fF
C45437 POR2X1_57/A PAND2X1_733/Y 0.19fF
C45438 POR2X1_850/A PAND2X1_60/B 0.01fF
C45439 POR2X1_73/Y VDD 1.47fF
C45440 PAND2X1_203/m4_208_n4# PAND2X1_575/A 0.17fF
C45441 POR2X1_278/Y PAND2X1_359/CTRL 0.01fF
C45442 PAND2X1_793/Y PAND2X1_357/Y 0.03fF
C45443 INPUT_3 POR2X1_39/B 0.75fF
C45444 PAND2X1_859/A PAND2X1_510/B 0.65fF
C45445 PAND2X1_807/CTRL VDD 0.00fF
C45446 POR2X1_41/B POR2X1_368/Y 0.02fF
C45447 PAND2X1_23/Y POR2X1_363/CTRL 0.01fF
C45448 PAND2X1_48/B POR2X1_205/CTRL 0.10fF
C45449 POR2X1_252/CTRL PAND2X1_6/A 0.03fF
C45450 PAND2X1_556/CTRL PAND2X1_348/A 0.04fF
C45451 POR2X1_43/B PAND2X1_215/B 0.05fF
C45452 PAND2X1_366/A PAND2X1_363/Y 0.13fF
C45453 PAND2X1_803/Y POR2X1_236/Y 0.02fF
C45454 POR2X1_592/A POR2X1_794/B 0.00fF
C45455 POR2X1_121/A POR2X1_294/B 0.01fF
C45456 POR2X1_502/A PAND2X1_96/B 0.06fF
C45457 PAND2X1_65/B POR2X1_407/CTRL2 0.01fF
C45458 PAND2X1_57/B POR2X1_68/B 0.22fF
C45459 POR2X1_493/CTRL VDD 0.00fF
C45460 INPUT_4 PAND2X1_32/B 0.03fF
C45461 POR2X1_65/A POR2X1_164/Y 0.03fF
C45462 POR2X1_42/Y POR2X1_396/CTRL 0.01fF
C45463 POR2X1_326/CTRL PAND2X1_41/B 0.03fF
C45464 PAND2X1_11/Y POR2X1_3/B 0.01fF
C45465 PAND2X1_821/a_76_28# POR2X1_857/B 0.02fF
C45466 PAND2X1_65/B POR2X1_566/B 0.05fF
C45467 POR2X1_198/CTRL POR2X1_35/Y 0.01fF
C45468 PAND2X1_823/O PAND2X1_41/B 0.08fF
C45469 POR2X1_93/CTRL2 POR2X1_55/Y 0.32fF
C45470 PAND2X1_572/a_16_344# INPUT_0 0.01fF
C45471 POR2X1_96/A PAND2X1_243/a_16_344# 0.02fF
C45472 POR2X1_301/CTRL2 POR2X1_335/A 0.01fF
C45473 INPUT_0 POR2X1_387/Y 0.09fF
C45474 POR2X1_388/a_16_28# POR2X1_566/A 0.02fF
C45475 PAND2X1_48/B POR2X1_731/CTRL 0.01fF
C45476 POR2X1_222/Y POR2X1_35/Y 0.03fF
C45477 PAND2X1_776/a_76_28# POR2X1_238/Y 0.02fF
C45478 POR2X1_16/A PAND2X1_340/CTRL2 0.00fF
C45479 PAND2X1_96/B PAND2X1_176/O 0.01fF
C45480 PAND2X1_48/B POR2X1_702/A 0.03fF
C45481 POR2X1_220/Y PAND2X1_163/CTRL2 0.00fF
C45482 POR2X1_785/A PAND2X1_32/B 1.28fF
C45483 POR2X1_464/Y PAND2X1_96/B 0.01fF
C45484 POR2X1_52/A POR2X1_382/Y 0.02fF
C45485 POR2X1_40/Y PAND2X1_560/B 0.03fF
C45486 PAND2X1_824/B PAND2X1_41/B 0.22fF
C45487 POR2X1_193/Y POR2X1_260/A 0.03fF
C45488 PAND2X1_96/B POR2X1_532/Y 0.10fF
C45489 POR2X1_43/B PAND2X1_6/A 0.10fF
C45490 PAND2X1_56/Y PAND2X1_6/Y 0.32fF
C45491 PAND2X1_6/Y POR2X1_795/B 0.15fF
C45492 POR2X1_51/A POR2X1_408/Y 0.01fF
C45493 POR2X1_138/O PAND2X1_32/B 0.01fF
C45494 POR2X1_860/A POR2X1_216/Y 0.03fF
C45495 POR2X1_157/CTRL2 POR2X1_36/B 0.01fF
C45496 PAND2X1_825/CTRL2 PAND2X1_57/B 0.01fF
C45497 POR2X1_13/A POR2X1_7/A 0.26fF
C45498 PAND2X1_857/CTRL2 POR2X1_83/B 0.01fF
C45499 PAND2X1_244/B VDD 0.48fF
C45500 POR2X1_391/O POR2X1_546/A 0.01fF
C45501 POR2X1_324/CTRL POR2X1_324/A 0.01fF
C45502 POR2X1_93/A POR2X1_618/O 0.01fF
C45503 POR2X1_7/B POR2X1_665/A 0.00fF
C45504 POR2X1_203/CTRL POR2X1_579/Y 0.00fF
C45505 POR2X1_634/A POR2X1_294/A 0.07fF
C45506 POR2X1_72/B PAND2X1_123/Y 0.10fF
C45507 POR2X1_807/A POR2X1_590/Y 0.01fF
C45508 PAND2X1_58/A POR2X1_188/Y 0.03fF
C45509 POR2X1_60/A PAND2X1_199/CTRL2 0.01fF
C45510 POR2X1_78/B POR2X1_596/CTRL 0.01fF
C45511 POR2X1_136/Y PAND2X1_553/B 0.07fF
C45512 POR2X1_65/A PAND2X1_800/O 0.05fF
C45513 PAND2X1_866/A PAND2X1_866/a_76_28# 0.04fF
C45514 D_GATE_222 POR2X1_570/B 0.07fF
C45515 PAND2X1_115/CTRL2 POR2X1_283/A 0.03fF
C45516 PAND2X1_422/CTRL2 POR2X1_294/B 0.05fF
C45517 PAND2X1_631/A PAND2X1_556/CTRL 0.00fF
C45518 POR2X1_25/Y POR2X1_698/CTRL 0.01fF
C45519 PAND2X1_784/CTRL POR2X1_245/Y 0.00fF
C45520 POR2X1_518/CTRL POR2X1_667/A 0.01fF
C45521 POR2X1_489/CTRL2 POR2X1_294/A 0.02fF
C45522 POR2X1_782/A PAND2X1_747/CTRL2 0.01fF
C45523 PAND2X1_797/Y POR2X1_83/B 0.03fF
C45524 POR2X1_532/A POR2X1_35/Y 5.49fF
C45525 PAND2X1_727/O VDD 0.00fF
C45526 POR2X1_38/B PAND2X1_6/A 0.11fF
C45527 POR2X1_96/A PAND2X1_728/O 0.04fF
C45528 POR2X1_68/A PAND2X1_670/CTRL2 0.00fF
C45529 PAND2X1_808/Y PAND2X1_774/O 0.02fF
C45530 POR2X1_755/a_16_28# PAND2X1_645/B 0.01fF
C45531 POR2X1_809/A PAND2X1_679/O 0.01fF
C45532 PAND2X1_632/a_16_344# INPUT_0 0.02fF
C45533 PAND2X1_119/m4_208_n4# POR2X1_294/B 0.03fF
C45534 PAND2X1_744/a_76_28# POR2X1_644/A 0.02fF
C45535 PAND2X1_605/a_16_344# INPUT_0 0.01fF
C45536 PAND2X1_219/a_76_28# POR2X1_591/Y 0.01fF
C45537 POR2X1_326/CTRL2 POR2X1_468/B 0.03fF
C45538 POR2X1_718/A PAND2X1_48/A 0.03fF
C45539 POR2X1_57/A PAND2X1_642/B 0.06fF
C45540 POR2X1_119/Y PAND2X1_240/CTRL 0.04fF
C45541 PAND2X1_486/CTRL2 PAND2X1_726/B 0.05fF
C45542 POR2X1_567/A POR2X1_186/Y 0.05fF
C45543 POR2X1_614/A POR2X1_203/CTRL 0.01fF
C45544 POR2X1_119/Y PAND2X1_786/a_76_28# 0.04fF
C45545 POR2X1_209/CTRL VDD 0.00fF
C45546 PAND2X1_631/O POR2X1_93/A 0.07fF
C45547 POR2X1_68/A POR2X1_510/Y 0.03fF
C45548 POR2X1_168/A POR2X1_97/A 0.05fF
C45549 VDD POR2X1_186/B 1.58fF
C45550 POR2X1_63/O POR2X1_7/A 0.01fF
C45551 POR2X1_516/Y PAND2X1_841/Y 0.05fF
C45552 POR2X1_537/Y POR2X1_830/A 0.00fF
C45553 POR2X1_101/Y POR2X1_572/B 0.03fF
C45554 POR2X1_367/CTRL2 POR2X1_191/Y 0.12fF
C45555 PAND2X1_23/Y POR2X1_507/O 0.01fF
C45556 POR2X1_334/Y PAND2X1_261/CTRL 0.04fF
C45557 PAND2X1_362/B POR2X1_594/CTRL2 0.01fF
C45558 D_INPUT_0 PAND2X1_72/A 0.11fF
C45559 POR2X1_43/B POR2X1_588/Y 0.06fF
C45560 PAND2X1_90/A POR2X1_456/B 0.03fF
C45561 POR2X1_824/CTRL2 POR2X1_236/Y 0.01fF
C45562 POR2X1_516/A POR2X1_184/Y 0.03fF
C45563 PAND2X1_6/Y POR2X1_383/A 0.24fF
C45564 POR2X1_186/Y POR2X1_542/O 0.01fF
C45565 POR2X1_730/Y POR2X1_803/A 0.03fF
C45566 POR2X1_362/B POR2X1_362/O 0.02fF
C45567 POR2X1_491/Y POR2X1_72/B 0.01fF
C45568 POR2X1_802/A VDD 0.10fF
C45569 POR2X1_110/Y POR2X1_237/O 0.06fF
C45570 PAND2X1_94/A POR2X1_790/B 0.03fF
C45571 POR2X1_130/A POR2X1_294/A 0.24fF
C45572 POR2X1_68/A POR2X1_276/Y 0.05fF
C45573 POR2X1_197/Y PAND2X1_88/Y 0.02fF
C45574 POR2X1_516/A PAND2X1_651/Y 0.10fF
C45575 POR2X1_72/B POR2X1_372/CTRL 0.13fF
C45576 POR2X1_824/CTRL VDD -0.00fF
C45577 POR2X1_614/A POR2X1_101/Y 0.10fF
C45578 POR2X1_121/B PAND2X1_52/B 0.09fF
C45579 POR2X1_814/A POR2X1_556/A 0.10fF
C45580 PAND2X1_465/CTRL POR2X1_77/Y 0.01fF
C45581 POR2X1_7/B PAND2X1_337/O 0.17fF
C45582 POR2X1_49/O POR2X1_29/A 0.01fF
C45583 POR2X1_164/Y PAND2X1_565/O 0.02fF
C45584 POR2X1_94/A PAND2X1_102/a_56_28# 0.00fF
C45585 POR2X1_123/A POR2X1_532/A 0.07fF
C45586 PAND2X1_649/A POR2X1_689/O 0.01fF
C45587 PAND2X1_315/a_16_344# PAND2X1_32/B 0.02fF
C45588 POR2X1_184/Y PAND2X1_301/CTRL 0.00fF
C45589 POR2X1_131/a_76_344# PAND2X1_349/A 0.00fF
C45590 POR2X1_68/A POR2X1_543/O 0.02fF
C45591 PAND2X1_659/Y POR2X1_498/O 0.18fF
C45592 POR2X1_416/B POR2X1_331/Y 0.03fF
C45593 POR2X1_43/B POR2X1_583/Y 0.06fF
C45594 POR2X1_112/CTRL POR2X1_332/B 0.01fF
C45595 POR2X1_307/Y POR2X1_512/CTRL2 0.01fF
C45596 PAND2X1_432/CTRL2 PAND2X1_72/A 0.01fF
C45597 POR2X1_264/Y POR2X1_558/Y 0.01fF
C45598 PAND2X1_865/Y POR2X1_79/A 0.00fF
C45599 POR2X1_57/A PAND2X1_550/B 0.06fF
C45600 POR2X1_664/a_16_28# POR2X1_651/Y 0.03fF
C45601 POR2X1_693/Y POR2X1_394/A 0.02fF
C45602 POR2X1_407/A POR2X1_590/Y 0.55fF
C45603 PAND2X1_359/Y POR2X1_55/Y 0.03fF
C45604 POR2X1_741/Y POR2X1_186/B 0.06fF
C45605 PAND2X1_162/A PAND2X1_162/CTRL 0.01fF
C45606 POR2X1_537/B POR2X1_725/Y 0.07fF
C45607 PAND2X1_865/Y PAND2X1_468/CTRL2 0.00fF
C45608 PAND2X1_55/Y PAND2X1_527/O 0.02fF
C45609 PAND2X1_857/A PAND2X1_661/Y 0.14fF
C45610 VDD PAND2X1_358/CTRL -0.00fF
C45611 PAND2X1_679/O POR2X1_728/A 0.00fF
C45612 POR2X1_222/A POR2X1_553/A 0.03fF
C45613 VDD PAND2X1_207/A 0.00fF
C45614 POR2X1_186/B PAND2X1_32/B 0.06fF
C45615 POR2X1_260/A PAND2X1_670/O 0.01fF
C45616 PAND2X1_716/CTRL PAND2X1_716/B 0.01fF
C45617 PAND2X1_48/A POR2X1_713/Y 0.01fF
C45618 POR2X1_119/Y POR2X1_43/B 6.05fF
C45619 PAND2X1_90/Y PAND2X1_72/A 0.27fF
C45620 POR2X1_62/Y D_INPUT_1 0.10fF
C45621 PAND2X1_675/a_76_28# POR2X1_416/B 0.02fF
C45622 POR2X1_574/Y POR2X1_318/A 0.07fF
C45623 PAND2X1_319/B PAND2X1_357/CTRL2 0.01fF
C45624 POR2X1_129/Y POR2X1_172/Y 0.00fF
C45625 PAND2X1_9/Y POR2X1_624/Y 0.02fF
C45626 POR2X1_680/CTRL PAND2X1_652/A 0.02fF
C45627 PAND2X1_20/A PAND2X1_234/CTRL 0.03fF
C45628 PAND2X1_96/B POR2X1_188/Y 0.03fF
C45629 PAND2X1_493/m4_208_n4# PAND2X1_717/m4_208_n4# 0.05fF
C45630 POR2X1_258/Y POR2X1_394/A 0.03fF
C45631 PAND2X1_490/O POR2X1_4/Y 0.04fF
C45632 POR2X1_110/CTRL2 POR2X1_387/Y 0.04fF
C45633 PAND2X1_838/O POR2X1_827/Y -0.00fF
C45634 PAND2X1_187/a_76_28# POR2X1_444/Y 0.01fF
C45635 POR2X1_736/CTRL2 POR2X1_188/Y 0.01fF
C45636 POR2X1_383/A PAND2X1_310/O 0.07fF
C45637 POR2X1_803/CTRL2 POR2X1_796/Y 0.01fF
C45638 POR2X1_795/B POR2X1_632/Y 0.07fF
C45639 POR2X1_20/B POR2X1_616/O 0.01fF
C45640 PAND2X1_217/CTRL PAND2X1_124/Y 0.00fF
C45641 PAND2X1_217/O PAND2X1_267/Y 0.02fF
C45642 PAND2X1_798/Y PAND2X1_354/O 0.02fF
C45643 PAND2X1_69/A PAND2X1_122/O 0.12fF
C45644 PAND2X1_94/A POR2X1_673/B 0.01fF
C45645 POR2X1_9/Y POR2X1_734/A 0.10fF
C45646 PAND2X1_469/B POR2X1_39/B 0.03fF
C45647 PAND2X1_356/O PAND2X1_354/Y 0.04fF
C45648 POR2X1_505/a_16_28# PAND2X1_632/B 0.02fF
C45649 POR2X1_647/B POR2X1_260/B 0.03fF
C45650 POR2X1_725/Y PAND2X1_48/A 0.07fF
C45651 POR2X1_859/O POR2X1_66/A 0.02fF
C45652 PAND2X1_253/O POR2X1_186/B 0.04fF
C45653 POR2X1_730/Y POR2X1_327/Y 0.06fF
C45654 POR2X1_16/A PAND2X1_853/B 0.07fF
C45655 POR2X1_48/A INPUT_3 0.05fF
C45656 POR2X1_814/B PAND2X1_234/CTRL 0.04fF
C45657 PAND2X1_175/a_76_28# PAND2X1_853/B 0.02fF
C45658 POR2X1_112/O POR2X1_510/Y 0.02fF
C45659 PAND2X1_447/CTRL POR2X1_102/Y 0.01fF
C45660 POR2X1_368/Y POR2X1_77/Y 0.02fF
C45661 POR2X1_754/A POR2X1_90/O 0.00fF
C45662 POR2X1_528/Y POR2X1_613/Y 0.01fF
C45663 PAND2X1_717/A PAND2X1_390/Y 0.03fF
C45664 POR2X1_795/B PAND2X1_52/B 0.03fF
C45665 PAND2X1_646/CTRL POR2X1_612/Y 0.01fF
C45666 PAND2X1_628/O VDD 0.00fF
C45667 POR2X1_41/B POR2X1_310/CTRL2 0.05fF
C45668 POR2X1_416/B POR2X1_765/a_16_28# 0.01fF
C45669 PAND2X1_653/Y POR2X1_416/B 0.07fF
C45670 PAND2X1_267/Y PAND2X1_124/Y 0.02fF
C45671 PAND2X1_47/B PAND2X1_47/O 0.00fF
C45672 POR2X1_837/a_16_28# POR2X1_837/A 0.10fF
C45673 PAND2X1_641/CTRL2 PAND2X1_476/A 0.00fF
C45674 POR2X1_812/A POR2X1_688/a_16_28# 0.05fF
C45675 PAND2X1_348/A PAND2X1_345/Y 0.02fF
C45676 POR2X1_41/B PAND2X1_147/O 0.05fF
C45677 POR2X1_27/m4_208_n4# POR2X1_27/Y 0.12fF
C45678 POR2X1_391/Y POR2X1_768/A 0.07fF
C45679 POR2X1_287/B POR2X1_486/a_56_344# 0.00fF
C45680 PAND2X1_731/A POR2X1_39/B 0.07fF
C45681 POR2X1_643/CTRL2 POR2X1_121/Y 0.00fF
C45682 POR2X1_864/A POR2X1_783/O 0.02fF
C45683 PAND2X1_675/O POR2X1_283/A 0.05fF
C45684 POR2X1_416/B POR2X1_426/Y 0.15fF
C45685 POR2X1_158/Y POR2X1_425/Y 2.05fF
C45686 PAND2X1_403/B POR2X1_20/B 0.16fF
C45687 PAND2X1_206/B POR2X1_5/Y 0.07fF
C45688 POR2X1_567/A POR2X1_339/O -0.01fF
C45689 POR2X1_315/Y POR2X1_316/Y 0.00fF
C45690 POR2X1_383/A POR2X1_632/Y 0.07fF
C45691 PAND2X1_26/A PAND2X1_36/a_16_344# 0.05fF
C45692 POR2X1_624/Y POR2X1_267/A 0.03fF
C45693 POR2X1_78/A POR2X1_266/CTRL 0.01fF
C45694 POR2X1_6/O POR2X1_4/Y 0.00fF
C45695 POR2X1_102/Y PAND2X1_791/a_56_28# 0.00fF
C45696 POR2X1_648/A PAND2X1_57/B 0.07fF
C45697 POR2X1_38/Y PAND2X1_332/Y 0.05fF
C45698 POR2X1_626/Y POR2X1_628/Y 0.06fF
C45699 POR2X1_62/Y POR2X1_620/B 0.53fF
C45700 POR2X1_825/Y POR2X1_396/O 0.00fF
C45701 POR2X1_361/O PAND2X1_72/A 0.02fF
C45702 PAND2X1_445/Y POR2X1_329/A 0.09fF
C45703 PAND2X1_827/CTRL POR2X1_296/B 0.01fF
C45704 POR2X1_66/B POR2X1_610/CTRL2 0.00fF
C45705 POR2X1_83/B PAND2X1_267/Y 0.23fF
C45706 POR2X1_62/Y PAND2X1_101/B 0.01fF
C45707 POR2X1_677/Y PAND2X1_658/B 0.04fF
C45708 POR2X1_65/A POR2X1_826/Y 0.03fF
C45709 PAND2X1_780/O VDD 0.00fF
C45710 POR2X1_150/Y PAND2X1_787/Y 0.05fF
C45711 POR2X1_863/A POR2X1_788/B 0.01fF
C45712 POR2X1_630/O POR2X1_632/B 0.02fF
C45713 POR2X1_383/A PAND2X1_52/B 0.19fF
C45714 POR2X1_624/B INPUT_0 0.03fF
C45715 POR2X1_567/B POR2X1_241/B 0.05fF
C45716 POR2X1_479/CTRL POR2X1_66/A 0.00fF
C45717 PAND2X1_207/CTRL2 POR2X1_40/Y 0.09fF
C45718 POR2X1_673/Y PAND2X1_529/a_16_344# 0.01fF
C45719 POR2X1_602/B POR2X1_866/A 0.03fF
C45720 PAND2X1_20/A POR2X1_856/B 0.03fF
C45721 POR2X1_99/CTRL POR2X1_243/Y 0.02fF
C45722 PAND2X1_381/Y POR2X1_29/A 1.61fF
C45723 POR2X1_113/a_76_344# POR2X1_768/A 0.01fF
C45724 POR2X1_116/A POR2X1_130/A 0.03fF
C45725 PAND2X1_20/A POR2X1_35/CTRL2 0.01fF
C45726 POR2X1_88/A INPUT_0 0.02fF
C45727 POR2X1_614/A PAND2X1_255/CTRL 0.08fF
C45728 POR2X1_431/Y INPUT_0 0.21fF
C45729 POR2X1_121/B POR2X1_288/CTRL 0.06fF
C45730 POR2X1_675/O POR2X1_466/A 0.31fF
C45731 POR2X1_458/Y POR2X1_804/A 0.10fF
C45732 PAND2X1_3/A POR2X1_750/B 0.03fF
C45733 POR2X1_399/a_16_28# POR2X1_411/B 0.01fF
C45734 PAND2X1_459/Y PAND2X1_9/Y 0.01fF
C45735 PAND2X1_95/B PAND2X1_53/a_16_344# 0.02fF
C45736 PAND2X1_222/A PAND2X1_593/CTRL2 0.00fF
C45737 POR2X1_461/Y POR2X1_790/CTRL2 0.02fF
C45738 POR2X1_23/O POR2X1_14/Y 0.03fF
C45739 PAND2X1_73/Y PAND2X1_531/a_56_28# 0.00fF
C45740 POR2X1_814/B POR2X1_856/B 0.10fF
C45741 POR2X1_83/B PAND2X1_215/O 0.02fF
C45742 POR2X1_568/B PAND2X1_680/CTRL 0.31fF
C45743 POR2X1_807/A POR2X1_807/CTRL 0.01fF
C45744 PAND2X1_466/A PAND2X1_466/O -0.00fF
C45745 PAND2X1_57/B POR2X1_68/Y 0.01fF
C45746 POR2X1_153/Y PAND2X1_332/Y 0.03fF
C45747 POR2X1_65/A POR2X1_283/CTRL 0.01fF
C45748 PAND2X1_415/CTRL POR2X1_293/Y 0.01fF
C45749 PAND2X1_52/CTRL2 POR2X1_532/A 0.01fF
C45750 GATE_479 POR2X1_32/A 0.03fF
C45751 PAND2X1_394/O POR2X1_330/Y 0.03fF
C45752 POR2X1_45/Y POR2X1_411/B 0.03fF
C45753 POR2X1_60/A PAND2X1_731/B 0.08fF
C45754 POR2X1_360/A PAND2X1_82/a_76_28# 0.02fF
C45755 PAND2X1_790/CTRL2 POR2X1_42/Y 0.08fF
C45756 POR2X1_48/A POR2X1_393/O 0.16fF
C45757 POR2X1_299/Y VDD 0.08fF
C45758 POR2X1_567/B PAND2X1_438/CTRL2 0.15fF
C45759 POR2X1_411/B POR2X1_234/CTRL 0.01fF
C45760 POR2X1_311/Y PAND2X1_562/B 0.07fF
C45761 POR2X1_455/A POR2X1_341/A 0.05fF
C45762 PAND2X1_223/CTRL2 POR2X1_283/Y 0.01fF
C45763 PAND2X1_651/Y POR2X1_490/CTRL2 0.05fF
C45764 POR2X1_636/B POR2X1_636/A 0.27fF
C45765 POR2X1_66/B PAND2X1_13/CTRL 0.03fF
C45766 POR2X1_639/A POR2X1_639/CTRL2 0.01fF
C45767 PAND2X1_117/CTRL2 POR2X1_493/A 0.01fF
C45768 POR2X1_448/CTRL PAND2X1_90/Y 0.27fF
C45769 POR2X1_555/A PAND2X1_626/CTRL 0.22fF
C45770 POR2X1_593/B POR2X1_330/Y 0.05fF
C45771 PAND2X1_661/Y POR2X1_329/A 0.00fF
C45772 PAND2X1_658/CTRL2 PAND2X1_474/A -0.00fF
C45773 POR2X1_257/A POR2X1_248/CTRL2 0.07fF
C45774 POR2X1_78/B POR2X1_241/B 0.01fF
C45775 POR2X1_16/A POR2X1_827/CTRL 0.01fF
C45776 POR2X1_515/CTRL2 PAND2X1_20/A 0.01fF
C45777 POR2X1_753/Y VDD 0.92fF
C45778 PAND2X1_93/B POR2X1_662/Y 0.03fF
C45779 PAND2X1_794/CTRL PAND2X1_580/B 0.00fF
C45780 POR2X1_411/Y POR2X1_48/A 0.01fF
C45781 POR2X1_796/Y POR2X1_800/A 0.02fF
C45782 POR2X1_800/CTRL2 D_GATE_865 0.20fF
C45783 POR2X1_16/A PAND2X1_439/CTRL 0.01fF
C45784 POR2X1_814/A POR2X1_772/CTRL2 0.01fF
C45785 POR2X1_78/B POR2X1_719/A 0.03fF
C45786 POR2X1_60/A POR2X1_256/CTRL2 0.00fF
C45787 POR2X1_457/CTRL2 POR2X1_370/Y 0.02fF
C45788 POR2X1_334/B POR2X1_558/B 0.05fF
C45789 PAND2X1_848/A POR2X1_48/A 0.01fF
C45790 POR2X1_490/Y PAND2X1_716/CTRL 0.01fF
C45791 PAND2X1_93/B PAND2X1_275/O 0.03fF
C45792 PAND2X1_557/A POR2X1_250/CTRL2 0.01fF
C45793 POR2X1_76/A POR2X1_112/Y 0.03fF
C45794 POR2X1_311/Y POR2X1_13/A 0.03fF
C45795 POR2X1_48/CTRL POR2X1_72/B 0.01fF
C45796 PAND2X1_675/A POR2X1_48/A 5.13fF
C45797 POR2X1_437/Y POR2X1_23/Y 0.01fF
C45798 D_GATE_662 POR2X1_444/A 0.08fF
C45799 PAND2X1_247/CTRL2 POR2X1_283/A 0.01fF
C45800 POR2X1_48/A PAND2X1_469/B 0.05fF
C45801 PAND2X1_412/O PAND2X1_90/Y 0.04fF
C45802 POR2X1_813/CTRL POR2X1_7/A 0.01fF
C45803 PAND2X1_475/a_16_344# PAND2X1_474/Y 0.03fF
C45804 POR2X1_83/B POR2X1_372/Y 0.07fF
C45805 PAND2X1_283/O POR2X1_66/A 0.03fF
C45806 POR2X1_57/A PAND2X1_212/CTRL 0.01fF
C45807 D_INPUT_7 PAND2X1_3/B 0.09fF
C45808 POR2X1_411/B PAND2X1_383/a_56_28# 0.00fF
C45809 PAND2X1_20/A POR2X1_128/a_56_344# 0.00fF
C45810 POR2X1_630/CTRL2 PAND2X1_96/B 0.03fF
C45811 PAND2X1_649/CTRL2 POR2X1_32/A 0.03fF
C45812 POR2X1_43/B PAND2X1_97/a_76_28# 0.02fF
C45813 POR2X1_47/CTRL2 POR2X1_83/B 0.00fF
C45814 POR2X1_662/Y POR2X1_78/A 0.00fF
C45815 POR2X1_13/A PAND2X1_140/CTRL2 0.00fF
C45816 POR2X1_493/A PAND2X1_96/B 0.03fF
C45817 PAND2X1_90/A PAND2X1_9/CTRL 0.01fF
C45818 PAND2X1_808/Y PAND2X1_772/CTRL2 0.01fF
C45819 POR2X1_476/CTRL2 POR2X1_121/Y 0.11fF
C45820 POR2X1_55/CTRL2 PAND2X1_6/A 0.03fF
C45821 POR2X1_300/CTRL POR2X1_102/Y 0.01fF
C45822 POR2X1_433/Y POR2X1_432/CTRL 0.01fF
C45823 POR2X1_351/Y POR2X1_97/A 0.03fF
C45824 PAND2X1_563/B VDD 0.03fF
C45825 POR2X1_83/B POR2X1_519/Y 0.04fF
C45826 POR2X1_407/A POR2X1_660/O 0.01fF
C45827 PAND2X1_581/a_76_28# INPUT_6 0.01fF
C45828 POR2X1_43/B POR2X1_442/Y 0.06fF
C45829 POR2X1_43/B POR2X1_497/CTRL 0.01fF
C45830 PAND2X1_639/B PAND2X1_639/CTRL2 0.01fF
C45831 POR2X1_427/Y POR2X1_46/Y 0.08fF
C45832 POR2X1_72/Y PAND2X1_659/A 0.01fF
C45833 POR2X1_48/A PAND2X1_731/A 0.01fF
C45834 POR2X1_631/A POR2X1_66/A 0.06fF
C45835 PAND2X1_73/Y PAND2X1_518/CTRL 0.03fF
C45836 PAND2X1_790/a_76_28# POR2X1_7/A 0.02fF
C45837 POR2X1_45/Y POR2X1_271/Y 0.03fF
C45838 PAND2X1_558/Y PAND2X1_493/Y 0.27fF
C45839 PAND2X1_65/B POR2X1_572/O 0.01fF
C45840 POR2X1_37/Y POR2X1_172/Y 0.03fF
C45841 POR2X1_68/A POR2X1_864/CTRL 0.05fF
C45842 POR2X1_77/Y PAND2X1_147/O 0.09fF
C45843 PAND2X1_94/A POR2X1_643/Y 0.00fF
C45844 POR2X1_744/Y POR2X1_394/A 0.01fF
C45845 PAND2X1_57/B POR2X1_480/A 0.10fF
C45846 POR2X1_362/B POR2X1_405/Y 0.36fF
C45847 POR2X1_461/Y POR2X1_559/A 0.00fF
C45848 POR2X1_121/B PAND2X1_743/O 0.15fF
C45849 PAND2X1_39/B POR2X1_244/Y 0.12fF
C45850 PAND2X1_482/CTRL POR2X1_541/B 0.07fF
C45851 POR2X1_233/CTRL POR2X1_236/Y 0.01fF
C45852 POR2X1_618/CTRL POR2X1_5/Y 0.00fF
C45853 PAND2X1_865/CTRL2 POR2X1_23/Y 0.09fF
C45854 POR2X1_814/B POR2X1_791/O 0.02fF
C45855 POR2X1_362/B POR2X1_784/A 0.03fF
C45856 POR2X1_614/A POR2X1_800/CTRL2 0.03fF
C45857 PAND2X1_431/O POR2X1_440/Y 0.04fF
C45858 PAND2X1_785/Y VDD 0.42fF
C45859 POR2X1_65/A PAND2X1_736/A 0.01fF
C45860 POR2X1_338/CTRL POR2X1_97/A 0.01fF
C45861 PAND2X1_684/CTRL2 POR2X1_260/B 0.01fF
C45862 PAND2X1_3/CTRL2 PAND2X1_3/A 0.01fF
C45863 PAND2X1_723/Y POR2X1_7/B 0.22fF
C45864 POR2X1_309/CTRL2 POR2X1_387/Y 0.06fF
C45865 PAND2X1_57/B POR2X1_243/Y 0.07fF
C45866 POR2X1_853/CTRL VDD 0.00fF
C45867 PAND2X1_73/CTRL PAND2X1_69/A 0.00fF
C45868 POR2X1_319/A POR2X1_703/Y 0.02fF
C45869 PAND2X1_44/CTRL2 PAND2X1_32/B 0.00fF
C45870 PAND2X1_833/CTRL2 POR2X1_495/Y 0.00fF
C45871 PAND2X1_480/B PAND2X1_735/Y 0.09fF
C45872 PAND2X1_347/Y POR2X1_7/B 0.03fF
C45873 PAND2X1_272/CTRL2 POR2X1_569/A 0.02fF
C45874 PAND2X1_598/a_16_344# INPUT_0 0.02fF
C45875 POR2X1_493/B POR2X1_493/A 0.00fF
C45876 PAND2X1_48/B POR2X1_542/m4_208_n4# 0.08fF
C45877 POR2X1_32/A PAND2X1_175/B 0.03fF
C45878 PAND2X1_824/B POR2X1_454/A 0.04fF
C45879 PAND2X1_96/B PAND2X1_74/O 0.17fF
C45880 POR2X1_62/Y INPUT_3 0.12fF
C45881 POR2X1_29/A POR2X1_7/A 0.06fF
C45882 POR2X1_16/A POR2X1_23/Y 0.53fF
C45883 PAND2X1_428/O PAND2X1_32/B 0.03fF
C45884 PAND2X1_496/CTRL2 INPUT_0 0.03fF
C45885 POR2X1_306/Y PAND2X1_651/Y 0.00fF
C45886 POR2X1_42/Y POR2X1_236/Y 0.13fF
C45887 POR2X1_614/A POR2X1_801/CTRL 0.01fF
C45888 POR2X1_72/B PAND2X1_186/CTRL2 0.04fF
C45889 POR2X1_102/Y POR2X1_387/Y 2.31fF
C45890 POR2X1_255/a_16_28# POR2X1_184/Y 0.03fF
C45891 PAND2X1_281/CTRL POR2X1_647/B 0.01fF
C45892 POR2X1_502/A POR2X1_708/B 0.03fF
C45893 PAND2X1_733/A POR2X1_591/Y 12.84fF
C45894 POR2X1_137/B PAND2X1_134/CTRL 0.01fF
C45895 PAND2X1_48/B POR2X1_471/O 0.01fF
C45896 POR2X1_722/Y POR2X1_513/B 0.02fF
C45897 POR2X1_78/A POR2X1_181/B 0.03fF
C45898 PAND2X1_341/CTRL INPUT_0 0.07fF
C45899 POR2X1_734/A PAND2X1_518/O 0.12fF
C45900 PAND2X1_656/a_76_28# PAND2X1_656/A 0.01fF
C45901 POR2X1_793/A PAND2X1_90/Y 0.02fF
C45902 PAND2X1_48/Y POR2X1_786/Y 0.03fF
C45903 POR2X1_49/Y PAND2X1_724/O 0.04fF
C45904 POR2X1_590/A POR2X1_101/Y 0.08fF
C45905 PAND2X1_654/CTRL POR2X1_13/A 0.16fF
C45906 POR2X1_96/A POR2X1_406/O 0.01fF
C45907 POR2X1_356/A PAND2X1_524/O 0.19fF
C45908 POR2X1_417/Y POR2X1_142/Y 0.03fF
C45909 PAND2X1_97/O POR2X1_153/Y 0.16fF
C45910 POR2X1_459/A VDD -0.00fF
C45911 PAND2X1_794/B PAND2X1_366/Y 0.03fF
C45912 PAND2X1_90/A PAND2X1_57/B 0.86fF
C45913 POR2X1_74/a_16_28# POR2X1_23/Y 0.10fF
C45914 PAND2X1_6/Y PAND2X1_627/CTRL2 0.01fF
C45915 POR2X1_68/A POR2X1_471/CTRL2 0.01fF
C45916 POR2X1_102/Y PAND2X1_121/O 0.02fF
C45917 POR2X1_625/O POR2X1_90/Y 0.01fF
C45918 POR2X1_596/A PAND2X1_597/CTRL2 0.01fF
C45919 POR2X1_814/B PAND2X1_757/CTRL2 0.01fF
C45920 POR2X1_777/B PAND2X1_60/B 0.08fF
C45921 POR2X1_270/O POR2X1_814/B 0.05fF
C45922 POR2X1_634/A POR2X1_710/Y 0.30fF
C45923 POR2X1_515/Y VDD 0.12fF
C45924 POR2X1_719/a_16_28# POR2X1_719/A 0.05fF
C45925 POR2X1_14/Y POR2X1_750/Y 0.03fF
C45926 POR2X1_158/CTRL2 POR2X1_257/A 0.03fF
C45927 PAND2X1_115/O PAND2X1_115/Y 0.02fF
C45928 POR2X1_406/Y PAND2X1_716/O 0.07fF
C45929 PAND2X1_217/B PAND2X1_656/A 0.00fF
C45930 POR2X1_327/Y POR2X1_218/Y 0.03fF
C45931 INPUT_1 PAND2X1_77/O 0.03fF
C45932 POR2X1_390/B POR2X1_105/CTRL 0.00fF
C45933 PAND2X1_6/Y INPUT_0 0.06fF
C45934 POR2X1_32/A PAND2X1_777/CTRL 0.01fF
C45935 PAND2X1_23/Y POR2X1_193/A 0.03fF
C45936 POR2X1_466/A PAND2X1_313/m4_208_n4# 0.06fF
C45937 PAND2X1_23/Y POR2X1_579/Y 0.43fF
C45938 POR2X1_230/CTRL2 PAND2X1_338/B 0.03fF
C45939 POR2X1_770/O POR2X1_770/A 0.01fF
C45940 POR2X1_52/A POR2X1_45/Y 0.03fF
C45941 PAND2X1_557/A PAND2X1_593/Y 0.00fF
C45942 POR2X1_542/B VDD 0.31fF
C45943 PAND2X1_483/CTRL POR2X1_482/Y 0.01fF
C45944 POR2X1_65/A POR2X1_765/Y 0.03fF
C45945 POR2X1_356/A D_GATE_222 0.10fF
C45946 POR2X1_219/B POR2X1_215/CTRL 0.05fF
C45947 PAND2X1_65/B PAND2X1_60/B 0.13fF
C45948 POR2X1_154/a_16_28# POR2X1_803/A 0.02fF
C45949 PAND2X1_474/Y POR2X1_38/Y 0.05fF
C45950 PAND2X1_79/Y VDD 0.26fF
C45951 PAND2X1_20/A POR2X1_244/Y 0.03fF
C45952 POR2X1_416/B POR2X1_20/B 2.22fF
C45953 POR2X1_537/Y D_INPUT_0 0.03fF
C45954 POR2X1_15/O VDD 0.00fF
C45955 PAND2X1_48/B PAND2X1_146/O 0.05fF
C45956 POR2X1_389/A POR2X1_130/A 0.07fF
C45957 POR2X1_215/O PAND2X1_88/Y 0.01fF
C45958 POR2X1_13/A POR2X1_38/Y 0.07fF
C45959 PAND2X1_660/Y PAND2X1_660/B 0.01fF
C45960 POR2X1_16/A POR2X1_312/Y 0.03fF
C45961 POR2X1_360/A PAND2X1_69/A 0.07fF
C45962 D_INPUT_3 INPUT_0 0.49fF
C45963 POR2X1_178/Y PAND2X1_220/Y 0.43fF
C45964 PAND2X1_131/O POR2X1_318/A 0.05fF
C45965 POR2X1_859/A POR2X1_750/CTRL2 0.03fF
C45966 POR2X1_42/Y PAND2X1_850/O 0.03fF
C45967 POR2X1_68/A POR2X1_803/A 0.04fF
C45968 PAND2X1_682/CTRL2 POR2X1_68/A 0.13fF
C45969 POR2X1_839/O POR2X1_566/B 0.04fF
C45970 PAND2X1_20/A PAND2X1_527/CTRL2 0.02fF
C45971 POR2X1_62/Y POR2X1_78/A 0.05fF
C45972 POR2X1_124/O PAND2X1_96/B 0.02fF
C45973 POR2X1_272/Y PAND2X1_349/A 0.04fF
C45974 VDD PAND2X1_656/A 0.45fF
C45975 POR2X1_614/A PAND2X1_23/Y 0.77fF
C45976 PAND2X1_117/O PAND2X1_32/B 0.01fF
C45977 INPUT_2 POR2X1_119/CTRL 0.01fF
C45978 PAND2X1_367/A PAND2X1_366/Y 0.01fF
C45979 PAND2X1_714/O POR2X1_73/Y 0.02fF
C45980 POR2X1_556/A PAND2X1_135/CTRL2 0.01fF
C45981 POR2X1_525/CTRL PAND2X1_726/B 0.03fF
C45982 POR2X1_811/B PAND2X1_48/A 0.03fF
C45983 POR2X1_492/CTRL2 POR2X1_394/A 0.05fF
C45984 POR2X1_516/CTRL2 PAND2X1_6/A 0.10fF
C45985 POR2X1_256/CTRL POR2X1_7/A 0.02fF
C45986 PAND2X1_137/Y PAND2X1_388/Y 0.07fF
C45987 POR2X1_57/O POR2X1_38/Y 0.15fF
C45988 POR2X1_219/B POR2X1_740/Y 0.10fF
C45989 POR2X1_809/A POR2X1_864/O 0.01fF
C45990 POR2X1_133/a_16_28# POR2X1_93/A 0.03fF
C45991 POR2X1_814/B POR2X1_244/Y 0.05fF
C45992 PAND2X1_734/B POR2X1_229/Y 0.01fF
C45993 POR2X1_348/A POR2X1_344/Y 0.03fF
C45994 POR2X1_726/Y VDD 0.10fF
C45995 POR2X1_76/Y POR2X1_366/A 0.03fF
C45996 POR2X1_861/O POR2X1_501/B 0.03fF
C45997 POR2X1_542/B POR2X1_741/Y 0.03fF
C45998 PAND2X1_467/Y PAND2X1_707/CTRL2 0.01fF
C45999 POR2X1_164/CTRL2 PAND2X1_565/A 0.00fF
C46000 PAND2X1_20/A POR2X1_191/Y 0.05fF
C46001 POR2X1_205/O POR2X1_203/Y 0.00fF
C46002 PAND2X1_217/B POR2X1_300/Y 0.06fF
C46003 PAND2X1_376/CTRL VDD 0.00fF
C46004 PAND2X1_776/O POR2X1_91/Y 0.01fF
C46005 POR2X1_562/a_16_28# POR2X1_341/Y 0.03fF
C46006 POR2X1_775/A POR2X1_775/a_16_28# 0.03fF
C46007 POR2X1_63/O POR2X1_38/Y 0.03fF
C46008 POR2X1_13/A POR2X1_597/m4_208_n4# 0.07fF
C46009 PAND2X1_560/B POR2X1_5/Y 0.02fF
C46010 PAND2X1_81/B PAND2X1_79/Y 0.03fF
C46011 POR2X1_128/A POR2X1_735/O 0.00fF
C46012 POR2X1_51/A POR2X1_744/CTRL 0.01fF
C46013 POR2X1_66/A POR2X1_736/A 0.03fF
C46014 POR2X1_228/Y POR2X1_556/O 0.06fF
C46015 POR2X1_78/A PAND2X1_179/a_16_344# 0.01fF
C46016 INPUT_1 POR2X1_13/A 0.97fF
C46017 POR2X1_793/A POR2X1_789/O 0.01fF
C46018 POR2X1_383/A PAND2X1_95/B 0.03fF
C46019 POR2X1_369/O POR2X1_236/Y 0.01fF
C46020 PAND2X1_59/B PAND2X1_72/A 0.06fF
C46021 POR2X1_220/Y POR2X1_675/Y 0.03fF
C46022 INPUT_1 PAND2X1_38/O 0.03fF
C46023 POR2X1_7/B PAND2X1_346/Y 0.03fF
C46024 PAND2X1_787/A PAND2X1_566/Y 0.29fF
C46025 PAND2X1_852/B POR2X1_73/Y 0.01fF
C46026 POR2X1_501/B POR2X1_500/Y 0.08fF
C46027 POR2X1_855/Y POR2X1_260/A 0.03fF
C46028 PAND2X1_605/CTRL POR2X1_7/B 0.01fF
C46029 POR2X1_228/Y POR2X1_723/B 0.01fF
C46030 POR2X1_809/A D_GATE_865 0.01fF
C46031 PAND2X1_397/CTRL POR2X1_35/Y 0.01fF
C46032 POR2X1_184/Y PAND2X1_175/B 0.02fF
C46033 PAND2X1_793/Y PAND2X1_579/A 0.01fF
C46034 POR2X1_188/A POR2X1_840/Y 0.02fF
C46035 POR2X1_13/A POR2X1_153/Y 0.19fF
C46036 POR2X1_292/CTRL POR2X1_411/B 0.03fF
C46037 POR2X1_300/Y VDD 0.21fF
C46038 POR2X1_220/Y POR2X1_544/B 0.03fF
C46039 POR2X1_327/Y POR2X1_115/CTRL 0.01fF
C46040 POR2X1_360/A PAND2X1_824/B 0.03fF
C46041 POR2X1_13/A POR2X1_384/A 0.01fF
C46042 POR2X1_123/A PAND2X1_132/m4_208_n4# 0.08fF
C46043 PAND2X1_6/A POR2X1_384/O 0.01fF
C46044 PAND2X1_651/Y PAND2X1_175/B 0.05fF
C46045 POR2X1_7/B PAND2X1_112/a_76_28# 0.07fF
C46046 POR2X1_566/A POR2X1_334/Y 0.10fF
C46047 PAND2X1_467/Y PAND2X1_725/A 0.36fF
C46048 PAND2X1_662/Y VDD 0.13fF
C46049 POR2X1_623/A PAND2X1_6/A 0.03fF
C46050 PAND2X1_96/B POR2X1_510/Y 1.18fF
C46051 POR2X1_445/O POR2X1_186/B 0.01fF
C46052 PAND2X1_858/CTRL2 POR2X1_13/A 0.03fF
C46053 POR2X1_614/A POR2X1_520/A 0.04fF
C46054 POR2X1_302/O POR2X1_188/Y 0.01fF
C46055 POR2X1_495/CTRL POR2X1_39/B 0.01fF
C46056 POR2X1_448/Y POR2X1_532/CTRL 0.02fF
C46057 PAND2X1_362/B POR2X1_385/Y 0.03fF
C46058 POR2X1_108/O POR2X1_387/Y 0.28fF
C46059 PAND2X1_455/CTRL2 POR2X1_77/Y 0.01fF
C46060 POR2X1_680/Y PAND2X1_853/B 0.08fF
C46061 POR2X1_375/CTRL2 PAND2X1_32/B 0.00fF
C46062 POR2X1_57/A PAND2X1_130/CTRL 0.01fF
C46063 PAND2X1_390/Y POR2X1_77/Y 0.03fF
C46064 POR2X1_327/Y PAND2X1_152/a_16_344# 0.04fF
C46065 POR2X1_814/B PAND2X1_102/O 0.09fF
C46066 PAND2X1_658/A POR2X1_751/Y 0.00fF
C46067 POR2X1_57/A PAND2X1_661/Y 0.10fF
C46068 PAND2X1_94/A PAND2X1_63/Y 0.16fF
C46069 POR2X1_469/a_16_28# POR2X1_444/Y -0.00fF
C46070 POR2X1_863/A POR2X1_436/B 3.48fF
C46071 POR2X1_355/B POR2X1_447/B 0.03fF
C46072 POR2X1_529/O POR2X1_384/A 0.01fF
C46073 POR2X1_175/B POR2X1_570/B 0.02fF
C46074 POR2X1_177/O PAND2X1_552/B 0.18fF
C46075 POR2X1_61/O PAND2X1_69/A 0.01fF
C46076 POR2X1_66/A PAND2X1_125/a_56_28# 0.00fF
C46077 POR2X1_315/Y PAND2X1_787/A 0.00fF
C46078 POR2X1_86/CTRL VDD 0.00fF
C46079 POR2X1_124/B POR2X1_768/CTRL 0.00fF
C46080 PAND2X1_620/O PAND2X1_651/Y 0.00fF
C46081 POR2X1_327/Y POR2X1_68/A 0.32fF
C46082 POR2X1_216/CTRL2 POR2X1_276/Y 0.01fF
C46083 PAND2X1_698/O POR2X1_532/A 0.13fF
C46084 PAND2X1_699/CTRL2 POR2X1_628/Y 0.00fF
C46085 POR2X1_463/Y POR2X1_532/A 0.10fF
C46086 D_INPUT_1 POR2X1_6/O 0.03fF
C46087 POR2X1_62/Y POR2X1_620/CTRL2 0.00fF
C46088 PAND2X1_704/O POR2X1_90/Y 0.17fF
C46089 POR2X1_833/A POR2X1_68/B 0.03fF
C46090 POR2X1_112/CTRL POR2X1_579/Y 0.00fF
C46091 PAND2X1_94/A POR2X1_113/Y 0.05fF
C46092 POR2X1_411/B POR2X1_271/B 0.03fF
C46093 PAND2X1_274/CTRL2 POR2X1_39/B 0.03fF
C46094 PAND2X1_649/A POR2X1_689/A 0.93fF
C46095 PAND2X1_853/a_76_28# PAND2X1_853/B 0.02fF
C46096 POR2X1_614/A POR2X1_809/A 0.04fF
C46097 PAND2X1_555/Y POR2X1_394/A 2.03fF
C46098 POR2X1_837/B POR2X1_296/B 2.24fF
C46099 POR2X1_54/Y POR2X1_859/CTRL 0.01fF
C46100 PAND2X1_655/Y POR2X1_690/CTRL 0.01fF
C46101 POR2X1_218/O POR2X1_362/A 0.00fF
C46102 POR2X1_218/m4_208_n4# POR2X1_361/m4_208_n4# 0.15fF
C46103 POR2X1_52/A POR2X1_305/CTRL2 0.03fF
C46104 POR2X1_732/B PAND2X1_179/CTRL 0.03fF
C46105 POR2X1_675/Y POR2X1_737/CTRL2 0.01fF
C46106 INPUT_0 PAND2X1_52/B 0.12fF
C46107 PAND2X1_425/Y PAND2X1_581/CTRL 0.01fF
C46108 POR2X1_110/Y POR2X1_417/O 0.01fF
C46109 PAND2X1_94/A POR2X1_260/A 0.46fF
C46110 PAND2X1_651/Y PAND2X1_500/CTRL 0.01fF
C46111 POR2X1_257/A POR2X1_694/Y 0.01fF
C46112 PAND2X1_453/CTRL POR2X1_77/Y 0.00fF
C46113 PAND2X1_39/B PAND2X1_27/O 0.06fF
C46114 POR2X1_153/Y PAND2X1_510/B 0.03fF
C46115 PAND2X1_631/A PAND2X1_344/CTRL2 0.05fF
C46116 POR2X1_384/A PAND2X1_510/B 0.00fF
C46117 POR2X1_452/a_16_28# POR2X1_450/Y -0.00fF
C46118 POR2X1_866/A PAND2X1_39/B 0.12fF
C46119 PAND2X1_569/B POR2X1_373/Y 0.02fF
C46120 POR2X1_119/Y PAND2X1_711/a_76_28# 0.01fF
C46121 PAND2X1_39/B POR2X1_195/A 0.01fF
C46122 POR2X1_447/B POR2X1_510/B 0.12fF
C46123 PAND2X1_476/A PAND2X1_338/B 0.03fF
C46124 PAND2X1_718/O POR2X1_77/Y 0.17fF
C46125 PAND2X1_216/B POR2X1_129/Y 0.11fF
C46126 PAND2X1_475/O POR2X1_329/A 0.03fF
C46127 PAND2X1_221/Y PAND2X1_366/Y 0.03fF
C46128 POR2X1_609/Y POR2X1_411/B 4.58fF
C46129 POR2X1_212/O POR2X1_191/Y 0.01fF
C46130 PAND2X1_193/Y VDD 0.28fF
C46131 POR2X1_760/A PAND2X1_361/CTRL 0.01fF
C46132 PAND2X1_476/A POR2X1_235/CTRL 0.00fF
C46133 POR2X1_614/A POR2X1_711/Y 0.07fF
C46134 POR2X1_785/A POR2X1_568/A 0.03fF
C46135 PAND2X1_50/CTRL2 D_INPUT_7 0.01fF
C46136 POR2X1_294/Y POR2X1_294/CTRL 0.00fF
C46137 POR2X1_438/CTRL POR2X1_77/Y 0.00fF
C46138 POR2X1_695/O POR2X1_48/A 0.14fF
C46139 POR2X1_309/CTRL POR2X1_411/B 0.01fF
C46140 POR2X1_485/Y POR2X1_83/B 0.03fF
C46141 D_GATE_222 PAND2X1_72/A 0.08fF
C46142 PAND2X1_659/Y PAND2X1_737/B 0.24fF
C46143 POR2X1_25/Y POR2X1_26/O 0.01fF
C46144 POR2X1_65/O POR2X1_40/Y 0.01fF
C46145 POR2X1_614/A POR2X1_728/A 0.01fF
C46146 POR2X1_532/A POR2X1_736/A 0.01fF
C46147 PAND2X1_659/Y PAND2X1_216/B 0.06fF
C46148 POR2X1_119/Y PAND2X1_123/a_56_28# 0.00fF
C46149 POR2X1_407/A POR2X1_717/B 0.07fF
C46150 POR2X1_554/B POR2X1_330/Y 0.03fF
C46151 POR2X1_66/B POR2X1_499/A 0.03fF
C46152 POR2X1_510/B POR2X1_510/O 0.07fF
C46153 PAND2X1_446/Y POR2X1_60/A 0.06fF
C46154 PAND2X1_738/A POR2X1_39/B 0.18fF
C46155 POR2X1_23/Y PAND2X1_214/O 0.03fF
C46156 PAND2X1_138/O POR2X1_129/Y 0.01fF
C46157 POR2X1_270/Y POR2X1_66/A 0.03fF
C46158 POR2X1_192/a_16_28# POR2X1_191/Y 0.03fF
C46159 POR2X1_66/B POR2X1_415/A 0.17fF
C46160 POR2X1_655/A POR2X1_121/B 0.04fF
C46161 POR2X1_327/Y POR2X1_861/A 0.01fF
C46162 POR2X1_153/Y PAND2X1_199/O 0.09fF
C46163 POR2X1_440/Y POR2X1_711/Y 0.35fF
C46164 POR2X1_773/A POR2X1_294/A 0.03fF
C46165 POR2X1_116/A POR2X1_105/Y 0.00fF
C46166 POR2X1_333/A POR2X1_212/a_56_344# 0.00fF
C46167 POR2X1_376/B POR2X1_271/B 0.03fF
C46168 POR2X1_66/B POR2X1_76/A 0.00fF
C46169 PAND2X1_431/O POR2X1_590/A 0.12fF
C46170 POR2X1_809/O POR2X1_121/B 0.03fF
C46171 POR2X1_815/CTRL INPUT_0 0.09fF
C46172 PAND2X1_20/A POR2X1_866/A 0.12fF
C46173 POR2X1_409/B POR2X1_32/A 0.03fF
C46174 POR2X1_180/A POR2X1_180/Y 0.09fF
C46175 POR2X1_669/Y VDD 0.01fF
C46176 PAND2X1_170/CTRL PAND2X1_326/B 0.01fF
C46177 POR2X1_65/A POR2X1_257/A 0.10fF
C46178 PAND2X1_677/m4_208_n4# POR2X1_678/m4_208_n4# 0.05fF
C46179 PAND2X1_677/CTRL POR2X1_260/B 0.01fF
C46180 POR2X1_399/CTRL POR2X1_20/B 0.01fF
C46181 POR2X1_149/A POR2X1_856/B 0.02fF
C46182 PAND2X1_65/B POR2X1_818/CTRL 0.00fF
C46183 POR2X1_169/A POR2X1_317/B 0.04fF
C46184 POR2X1_20/B PAND2X1_773/B 0.01fF
C46185 POR2X1_846/A POR2X1_790/B 0.03fF
C46186 PAND2X1_858/CTRL PAND2X1_850/Y 0.06fF
C46187 POR2X1_416/B PAND2X1_715/B 0.02fF
C46188 POR2X1_119/Y PAND2X1_865/Y 0.05fF
C46189 POR2X1_835/B POR2X1_776/B 0.01fF
C46190 PAND2X1_245/m4_208_n4# POR2X1_66/A 0.15fF
C46191 POR2X1_685/CTRL POR2X1_452/Y 0.01fF
C46192 POR2X1_78/A POR2X1_646/Y 0.00fF
C46193 POR2X1_812/A D_INPUT_0 0.01fF
C46194 PAND2X1_443/CTRL PAND2X1_803/A 0.00fF
C46195 POR2X1_20/B PAND2X1_738/Y 0.05fF
C46196 POR2X1_486/a_16_28# POR2X1_294/B 0.07fF
C46197 PAND2X1_48/B PAND2X1_53/O 0.01fF
C46198 POR2X1_776/A VDD 0.22fF
C46199 PAND2X1_467/B POR2X1_163/Y 0.10fF
C46200 POR2X1_594/Y POR2X1_760/A -0.00fF
C46201 POR2X1_319/A PAND2X1_90/Y 0.03fF
C46202 POR2X1_679/A PAND2X1_580/B 0.17fF
C46203 POR2X1_8/Y POR2X1_8/CTRL 0.01fF
C46204 POR2X1_39/B POR2X1_397/CTRL2 0.00fF
C46205 PAND2X1_6/Y PAND2X1_32/CTRL 0.01fF
C46206 POR2X1_83/B PAND2X1_249/CTRL2 0.01fF
C46207 PAND2X1_309/O POR2X1_556/A 0.01fF
C46208 POR2X1_415/A POR2X1_859/A 0.07fF
C46209 POR2X1_566/A POR2X1_854/CTRL 0.03fF
C46210 POR2X1_355/B POR2X1_446/A 0.11fF
C46211 POR2X1_496/Y POR2X1_72/B 0.25fF
C46212 PAND2X1_634/a_16_344# POR2X1_290/Y 0.01fF
C46213 PAND2X1_476/CTRL2 POR2X1_102/Y 0.01fF
C46214 POR2X1_262/Y PAND2X1_197/Y 0.23fF
C46215 PAND2X1_128/CTRL POR2X1_411/B 0.01fF
C46216 POR2X1_84/B PAND2X1_57/B 0.03fF
C46217 PAND2X1_839/CTRL POR2X1_20/B 0.01fF
C46218 POR2X1_54/Y POR2X1_754/A 1.16fF
C46219 POR2X1_659/A POR2X1_220/Y 0.03fF
C46220 POR2X1_423/CTRL POR2X1_423/Y 0.03fF
C46221 POR2X1_376/B PAND2X1_796/CTRL2 0.00fF
C46222 POR2X1_263/Y POR2X1_230/a_56_344# 0.00fF
C46223 PAND2X1_51/CTRL POR2X1_451/A 0.01fF
C46224 POR2X1_48/A POR2X1_689/O 0.18fF
C46225 PAND2X1_487/O PAND2X1_57/B 0.02fF
C46226 POR2X1_738/O POR2X1_731/Y 0.00fF
C46227 POR2X1_33/A PAND2X1_14/O 0.00fF
C46228 POR2X1_502/A POR2X1_260/B 0.18fF
C46229 POR2X1_179/O POR2X1_150/Y 0.01fF
C46230 POR2X1_416/A VDD 0.00fF
C46231 PAND2X1_410/CTRL POR2X1_290/Y 0.06fF
C46232 PAND2X1_463/CTRL2 POR2X1_94/A 0.01fF
C46233 POR2X1_836/A PAND2X1_41/B 0.04fF
C46234 POR2X1_856/B VDD 10.80fF
C46235 PAND2X1_73/Y POR2X1_573/CTRL2 0.01fF
C46236 POR2X1_814/A PAND2X1_60/B 0.22fF
C46237 POR2X1_196/O POR2X1_702/B 0.02fF
C46238 POR2X1_24/Y POR2X1_42/Y 0.03fF
C46239 POR2X1_41/B POR2X1_265/O 0.00fF
C46240 PAND2X1_75/CTRL PAND2X1_60/B 0.01fF
C46241 POR2X1_356/A POR2X1_446/O 0.04fF
C46242 POR2X1_866/A POR2X1_513/B 0.20fF
C46243 POR2X1_72/B PAND2X1_733/A 0.03fF
C46244 POR2X1_94/A POR2X1_750/A 0.03fF
C46245 POR2X1_458/Y PAND2X1_368/CTRL 0.06fF
C46246 POR2X1_65/A POR2X1_423/a_16_28# 0.06fF
C46247 POR2X1_452/Y POR2X1_730/O 0.01fF
C46248 POR2X1_251/A POR2X1_251/a_56_344# 0.00fF
C46249 POR2X1_142/O POR2X1_65/A 0.02fF
C46250 POR2X1_67/A POR2X1_236/Y 0.07fF
C46251 POR2X1_864/A POR2X1_644/A 0.03fF
C46252 POR2X1_54/Y PAND2X1_283/CTRL 0.01fF
C46253 POR2X1_67/Y POR2X1_283/A 0.03fF
C46254 POR2X1_272/Y POR2X1_32/A 0.07fF
C46255 PAND2X1_492/CTRL PAND2X1_73/Y 0.05fF
C46256 POR2X1_770/B VDD 0.02fF
C46257 PAND2X1_695/CTRL2 POR2X1_634/A 0.15fF
C46258 POR2X1_848/A POR2X1_615/Y 0.02fF
C46259 POR2X1_194/A POR2X1_750/B 0.36fF
C46260 POR2X1_865/B POR2X1_556/A 0.03fF
C46261 POR2X1_776/A PAND2X1_32/B 0.03fF
C46262 PAND2X1_793/Y D_INPUT_0 0.03fF
C46263 POR2X1_102/Y POR2X1_237/O 0.01fF
C46264 POR2X1_638/CTRL2 POR2X1_66/A 0.01fF
C46265 PAND2X1_65/B POR2X1_254/A 0.01fF
C46266 POR2X1_813/CTRL POR2X1_38/Y 0.03fF
C46267 POR2X1_274/m4_208_n4# POR2X1_325/A 0.01fF
C46268 POR2X1_298/a_16_28# POR2X1_55/Y 0.03fF
C46269 PAND2X1_39/B POR2X1_501/B 0.06fF
C46270 PAND2X1_9/Y PAND2X1_79/Y 0.00fF
C46271 PAND2X1_564/B VDD 0.18fF
C46272 POR2X1_49/Y POR2X1_65/A 0.44fF
C46273 POR2X1_266/CTRL2 PAND2X1_69/A 0.01fF
C46274 PAND2X1_206/B PAND2X1_100/CTRL 0.01fF
C46275 POR2X1_43/B PAND2X1_211/a_76_28# 0.02fF
C46276 PAND2X1_65/B POR2X1_750/B 0.14fF
C46277 PAND2X1_6/Y POR2X1_808/O 0.18fF
C46278 POR2X1_840/B POR2X1_624/Y 0.10fF
C46279 POR2X1_823/Y POR2X1_20/B 0.00fF
C46280 PAND2X1_48/B D_INPUT_0 0.08fF
C46281 POR2X1_270/Y POR2X1_222/Y 0.01fF
C46282 D_INPUT_3 POR2X1_263/a_16_28# 0.09fF
C46283 POR2X1_640/CTRL2 INPUT_0 0.06fF
C46284 PAND2X1_73/CTRL2 PAND2X1_8/Y 0.01fF
C46285 PAND2X1_65/B POR2X1_461/CTRL 0.03fF
C46286 PAND2X1_706/a_56_28# POR2X1_692/Y 0.00fF
C46287 POR2X1_567/B D_GATE_741 0.07fF
C46288 POR2X1_102/Y PAND2X1_598/a_16_344# 0.02fF
C46289 POR2X1_862/O PAND2X1_52/B 0.01fF
C46290 POR2X1_244/CTRL POR2X1_243/Y 0.07fF
C46291 PAND2X1_205/A POR2X1_816/A 0.01fF
C46292 POR2X1_13/A PAND2X1_244/a_16_344# 0.01fF
C46293 PAND2X1_556/B PAND2X1_168/Y 0.03fF
C46294 POR2X1_632/m4_208_n4# POR2X1_222/Y 0.15fF
C46295 PAND2X1_93/B POR2X1_804/A 0.05fF
C46296 PAND2X1_20/A PAND2X1_516/a_16_344# 0.01fF
C46297 POR2X1_3/A PAND2X1_12/O 0.01fF
C46298 POR2X1_13/A PAND2X1_214/A 0.02fF
C46299 PAND2X1_23/Y POR2X1_590/A 0.21fF
C46300 PAND2X1_55/Y POR2X1_202/B 0.84fF
C46301 D_INPUT_3 PAND2X1_340/B 0.00fF
C46302 POR2X1_645/CTRL POR2X1_718/A 0.01fF
C46303 POR2X1_416/B POR2X1_43/Y 0.01fF
C46304 PAND2X1_859/A POR2X1_224/CTRL2 0.01fF
C46305 POR2X1_181/a_16_28# POR2X1_181/A 0.03fF
C46306 PAND2X1_220/Y PAND2X1_347/Y 0.03fF
C46307 POR2X1_615/CTRL VDD -0.00fF
C46308 PAND2X1_454/B PAND2X1_549/B 0.01fF
C46309 PAND2X1_96/B POR2X1_499/CTRL2 -0.00fF
C46310 PAND2X1_804/B POR2X1_72/B 0.01fF
C46311 PAND2X1_244/O POR2X1_293/Y 0.07fF
C46312 PAND2X1_651/Y POR2X1_409/B 0.00fF
C46313 PAND2X1_212/O POR2X1_142/Y 0.03fF
C46314 POR2X1_856/B PAND2X1_32/B 0.03fF
C46315 PAND2X1_214/A PAND2X1_214/B 0.01fF
C46316 POR2X1_669/A POR2X1_669/B 0.02fF
C46317 POR2X1_302/Y POR2X1_814/B 0.00fF
C46318 POR2X1_763/A VDD 0.00fF
C46319 POR2X1_670/Y POR2X1_14/Y 0.00fF
C46320 POR2X1_13/O POR2X1_595/Y 0.00fF
C46321 POR2X1_624/CTRL2 POR2X1_94/A 0.01fF
C46322 POR2X1_528/CTRL POR2X1_14/Y 0.01fF
C46323 PAND2X1_354/A POR2X1_7/B 0.03fF
C46324 POR2X1_330/Y PAND2X1_369/CTRL 0.10fF
C46325 POR2X1_383/A POR2X1_655/A 0.01fF
C46326 POR2X1_528/CTRL PAND2X1_453/A 0.01fF
C46327 POR2X1_379/CTRL POR2X1_260/B 0.01fF
C46328 POR2X1_315/Y PAND2X1_469/O 0.06fF
C46329 POR2X1_105/Y POR2X1_723/a_76_344# 0.01fF
C46330 POR2X1_105/a_16_28# POR2X1_717/Y 0.03fF
C46331 POR2X1_96/A PAND2X1_363/Y 0.02fF
C46332 POR2X1_141/Y POR2X1_276/CTRL 0.01fF
C46333 PAND2X1_83/a_76_28# POR2X1_66/A 0.05fF
C46334 PAND2X1_94/A POR2X1_473/O 0.02fF
C46335 PAND2X1_41/B POR2X1_208/O 0.01fF
C46336 PAND2X1_85/Y POR2X1_243/Y 0.03fF
C46337 POR2X1_78/A POR2X1_804/A 0.05fF
C46338 POR2X1_218/Y POR2X1_361/CTRL2 0.06fF
C46339 POR2X1_185/a_16_28# PAND2X1_73/Y 0.03fF
C46340 PAND2X1_844/Y PAND2X1_61/Y 0.99fF
C46341 POR2X1_302/Y POR2X1_325/A 0.03fF
C46342 PAND2X1_464/Y POR2X1_14/Y 0.01fF
C46343 POR2X1_96/A POR2X1_485/CTRL 0.00fF
C46344 PAND2X1_473/B PAND2X1_735/Y 0.07fF
C46345 POR2X1_205/CTRL POR2X1_330/Y 0.00fF
C46346 PAND2X1_443/Y POR2X1_90/Y 0.01fF
C46347 POR2X1_835/B POR2X1_192/B 0.03fF
C46348 POR2X1_800/A POR2X1_330/Y 0.05fF
C46349 POR2X1_23/Y PAND2X1_549/B 0.07fF
C46350 POR2X1_48/A PAND2X1_738/A 0.01fF
C46351 POR2X1_38/Y POR2X1_29/A 0.05fF
C46352 POR2X1_14/Y PAND2X1_565/A 0.03fF
C46353 POR2X1_242/m4_208_n4# POR2X1_578/Y 0.07fF
C46354 POR2X1_401/CTRL POR2X1_401/B -0.00fF
C46355 POR2X1_122/O POR2X1_20/B 0.02fF
C46356 POR2X1_853/A PAND2X1_41/B 0.03fF
C46357 PAND2X1_20/A POR2X1_501/B 0.03fF
C46358 POR2X1_413/A POR2X1_607/a_16_28# 0.01fF
C46359 POR2X1_136/CTRL2 POR2X1_40/Y 0.03fF
C46360 PAND2X1_471/B VDD 0.11fF
C46361 POR2X1_722/Y VDD 0.49fF
C46362 POR2X1_267/A PAND2X1_79/Y 0.00fF
C46363 POR2X1_853/m4_208_n4# PAND2X1_41/B 0.12fF
C46364 POR2X1_234/Y VDD 0.13fF
C46365 PAND2X1_48/B PAND2X1_90/Y 0.24fF
C46366 POR2X1_78/B POR2X1_465/B 0.03fF
C46367 POR2X1_355/CTRL D_GATE_741 0.06fF
C46368 POR2X1_836/O POR2X1_566/B 0.34fF
C46369 POR2X1_841/B POR2X1_675/Y 0.03fF
C46370 PAND2X1_41/B POR2X1_391/Y 0.07fF
C46371 POR2X1_330/Y POR2X1_702/A 0.03fF
C46372 POR2X1_66/A POR2X1_101/Y 0.10fF
C46373 D_INPUT_3 POR2X1_102/Y 0.03fF
C46374 POR2X1_14/Y POR2X1_395/Y 0.06fF
C46375 PAND2X1_115/a_16_344# PAND2X1_787/Y 0.03fF
C46376 POR2X1_740/CTRL POR2X1_740/Y 0.00fF
C46377 PAND2X1_661/B PAND2X1_214/A 0.02fF
C46378 PAND2X1_859/A PAND2X1_227/CTRL2 0.01fF
C46379 POR2X1_865/B POR2X1_474/O 0.01fF
C46380 POR2X1_483/A POR2X1_833/CTRL 0.01fF
C46381 POR2X1_141/O POR2X1_514/Y 0.16fF
C46382 POR2X1_12/A POR2X1_762/CTRL 0.01fF
C46383 PAND2X1_472/O POR2X1_23/Y 0.01fF
C46384 POR2X1_63/CTRL2 POR2X1_236/Y 0.15fF
C46385 PAND2X1_62/CTRL PAND2X1_6/A 0.09fF
C46386 POR2X1_72/CTRL PAND2X1_651/Y 0.01fF
C46387 POR2X1_791/O VDD 0.00fF
C46388 PAND2X1_659/CTRL PAND2X1_575/A 0.03fF
C46389 POR2X1_174/A POR2X1_738/A 0.02fF
C46390 POR2X1_20/Y POR2X1_5/Y 0.01fF
C46391 PAND2X1_414/O POR2X1_39/B 0.17fF
C46392 POR2X1_283/A POR2X1_225/a_16_28# 0.02fF
C46393 POR2X1_566/A POR2X1_629/A 0.22fF
C46394 PAND2X1_859/A PAND2X1_509/CTRL 0.01fF
C46395 POR2X1_463/CTRL2 PAND2X1_52/B 0.26fF
C46396 POR2X1_814/B POR2X1_501/B 0.03fF
C46397 POR2X1_820/A POR2X1_38/Y 0.01fF
C46398 POR2X1_97/A POR2X1_502/O 0.01fF
C46399 PAND2X1_216/B PAND2X1_561/CTRL 0.01fF
C46400 POR2X1_41/B PAND2X1_592/Y 0.03fF
C46401 PAND2X1_76/Y POR2X1_816/A 0.18fF
C46402 POR2X1_663/a_16_28# POR2X1_662/Y 0.08fF
C46403 INPUT_5 POR2X1_7/B 0.02fF
C46404 POR2X1_272/Y POR2X1_184/Y 0.03fF
C46405 POR2X1_690/a_16_28# POR2X1_413/A 0.03fF
C46406 POR2X1_502/A PAND2X1_55/Y 0.10fF
C46407 POR2X1_403/a_76_344# PAND2X1_69/A 0.00fF
C46408 POR2X1_537/CTRL2 POR2X1_590/A 0.01fF
C46409 POR2X1_504/Y POR2X1_93/A 0.03fF
C46410 INPUT_1 POR2X1_29/A 0.42fF
C46411 PAND2X1_642/B POR2X1_236/Y 1.68fF
C46412 POR2X1_130/A POR2X1_218/A 0.10fF
C46413 POR2X1_413/Y POR2X1_411/Y 0.01fF
C46414 POR2X1_102/Y POR2X1_7/CTRL 0.01fF
C46415 POR2X1_669/B POR2X1_523/CTRL 0.01fF
C46416 PAND2X1_417/CTRL2 POR2X1_736/A 0.15fF
C46417 POR2X1_244/B D_GATE_222 0.03fF
C46418 POR2X1_183/Y VDD 0.55fF
C46419 POR2X1_740/Y PAND2X1_152/CTRL2 0.00fF
C46420 POR2X1_697/Y POR2X1_531/CTRL 0.01fF
C46421 PAND2X1_724/B POR2X1_7/B 0.02fF
C46422 POR2X1_741/Y POR2X1_722/Y 0.00fF
C46423 PAND2X1_787/A PAND2X1_787/O 0.04fF
C46424 POR2X1_828/Y POR2X1_686/O 0.18fF
C46425 PAND2X1_65/B POR2X1_686/CTRL2 0.01fF
C46426 PAND2X1_11/Y POR2X1_260/A 0.20fF
C46427 PAND2X1_23/Y POR2X1_857/B 0.11fF
C46428 PAND2X1_55/CTRL2 PAND2X1_60/B 0.01fF
C46429 POR2X1_128/A POR2X1_128/B 0.12fF
C46430 POR2X1_188/A POR2X1_539/A 0.02fF
C46431 POR2X1_188/A POR2X1_537/A 0.01fF
C46432 POR2X1_260/B POR2X1_188/Y 0.45fF
C46433 PAND2X1_631/CTRL2 POR2X1_625/Y 0.02fF
C46434 POR2X1_832/O POR2X1_804/A 0.35fF
C46435 POR2X1_671/CTRL POR2X1_38/B 0.01fF
C46436 PAND2X1_695/a_16_344# POR2X1_407/Y 0.00fF
C46437 POR2X1_29/A POR2X1_153/Y 0.09fF
C46438 POR2X1_57/A PAND2X1_719/CTRL2 0.03fF
C46439 POR2X1_860/A POR2X1_218/CTRL2 0.01fF
C46440 POR2X1_29/A POR2X1_384/A 0.64fF
C46441 POR2X1_96/A PAND2X1_779/Y 0.01fF
C46442 PAND2X1_35/Y POR2X1_229/CTRL2 0.01fF
C46443 POR2X1_119/Y POR2X1_265/a_76_344# 0.04fF
C46444 POR2X1_400/A PAND2X1_88/Y 0.01fF
C46445 POR2X1_66/A POR2X1_722/O 0.01fF
C46446 POR2X1_807/A POR2X1_590/CTRL 0.01fF
C46447 POR2X1_65/A PAND2X1_559/CTRL 0.01fF
C46448 POR2X1_141/m4_208_n4# POR2X1_574/Y 0.17fF
C46449 POR2X1_192/Y POR2X1_190/CTRL 0.31fF
C46450 PAND2X1_341/B POR2X1_263/Y 0.03fF
C46451 POR2X1_327/Y PAND2X1_58/A 0.10fF
C46452 POR2X1_376/A PAND2X1_8/Y 0.13fF
C46453 PAND2X1_535/CTRL2 POR2X1_236/Y 0.04fF
C46454 POR2X1_566/A POR2X1_447/O 0.25fF
C46455 POR2X1_526/a_16_28# PAND2X1_556/B 0.02fF
C46456 PAND2X1_484/a_16_344# PAND2X1_73/Y 0.01fF
C46457 POR2X1_383/A PAND2X1_386/m4_208_n4# 0.12fF
C46458 POR2X1_13/A POR2X1_591/Y 0.03fF
C46459 POR2X1_296/B PAND2X1_48/A 1.26fF
C46460 PAND2X1_372/a_16_344# D_INPUT_1 0.02fF
C46461 POR2X1_508/B POR2X1_836/O 0.00fF
C46462 POR2X1_32/A POR2X1_150/CTRL 0.01fF
C46463 PAND2X1_6/Y PAND2X1_273/CTRL2 0.08fF
C46464 PAND2X1_803/a_16_344# POR2X1_83/B 0.01fF
C46465 POR2X1_814/B POR2X1_703/A 0.03fF
C46466 POR2X1_351/B PAND2X1_20/A 0.01fF
C46467 PAND2X1_696/CTRL2 POR2X1_66/A 0.01fF
C46468 PAND2X1_551/Y PAND2X1_324/Y 0.01fF
C46469 PAND2X1_480/B PAND2X1_787/A 0.10fF
C46470 POR2X1_335/A POR2X1_68/A 0.03fF
C46471 POR2X1_614/A POR2X1_733/A 0.07fF
C46472 PAND2X1_65/B POR2X1_502/CTRL2 0.00fF
C46473 POR2X1_368/O POR2X1_387/Y 0.04fF
C46474 PAND2X1_119/CTRL POR2X1_294/B 0.04fF
C46475 POR2X1_614/A POR2X1_334/B 0.39fF
C46476 POR2X1_833/A PAND2X1_46/a_76_28# 0.02fF
C46477 PAND2X1_550/B POR2X1_236/Y 0.06fF
C46478 POR2X1_57/A PAND2X1_520/a_76_28# 0.02fF
C46479 PAND2X1_807/O POR2X1_7/B 0.04fF
C46480 PAND2X1_614/CTRL2 POR2X1_129/Y 0.01fF
C46481 PAND2X1_563/a_16_344# PAND2X1_566/Y 0.04fF
C46482 POR2X1_65/A POR2X1_41/O 0.01fF
C46483 POR2X1_38/Y POR2X1_406/O 0.17fF
C46484 PAND2X1_691/Y PAND2X1_687/Y 0.06fF
C46485 POR2X1_68/B POR2X1_294/B 0.18fF
C46486 INPUT_0 POR2X1_385/CTRL2 0.01fF
C46487 POR2X1_563/O POR2X1_456/B 0.01fF
C46488 PAND2X1_469/Y POR2X1_46/Y 0.05fF
C46489 POR2X1_596/Y POR2X1_796/A 0.01fF
C46490 PAND2X1_213/Y POR2X1_763/Y 0.07fF
C46491 POR2X1_334/B POR2X1_38/B 0.27fF
C46492 PAND2X1_863/B PAND2X1_854/A 0.02fF
C46493 POR2X1_516/Y PAND2X1_851/a_16_344# 0.01fF
C46494 PAND2X1_453/CTRL PAND2X1_241/Y 0.01fF
C46495 POR2X1_668/a_16_28# POR2X1_260/A 0.01fF
C46496 POR2X1_814/A POR2X1_655/O 0.35fF
C46497 POR2X1_518/O POR2X1_669/B 0.33fF
C46498 PAND2X1_219/A PAND2X1_737/CTRL 0.01fF
C46499 PAND2X1_90/A POR2X1_137/Y 0.03fF
C46500 PAND2X1_339/Y POR2X1_522/Y 0.01fF
C46501 PAND2X1_216/O PAND2X1_656/A 0.01fF
C46502 POR2X1_119/Y PAND2X1_478/B 0.04fF
C46503 POR2X1_808/O PAND2X1_52/B 0.05fF
C46504 POR2X1_853/A POR2X1_170/m4_208_n4# 0.01fF
C46505 POR2X1_406/Y PAND2X1_737/B 0.14fF
C46506 POR2X1_507/B POR2X1_186/Y 0.10fF
C46507 POR2X1_119/Y POR2X1_609/CTRL 0.04fF
C46508 POR2X1_647/Y POR2X1_737/A 0.01fF
C46509 POR2X1_22/A POR2X1_3/a_76_344# 0.00fF
C46510 POR2X1_68/A POR2X1_844/O 0.16fF
C46511 POR2X1_198/a_76_344# PAND2X1_88/Y 0.00fF
C46512 POR2X1_317/CTRL POR2X1_854/B 0.29fF
C46513 POR2X1_3/A PAND2X1_635/CTRL2 0.00fF
C46514 POR2X1_244/Y VDD 0.40fF
C46515 POR2X1_703/A PAND2X1_176/CTRL2 0.00fF
C46516 POR2X1_196/Y POR2X1_219/B 0.12fF
C46517 PAND2X1_316/CTRL POR2X1_318/A 0.02fF
C46518 POR2X1_57/A PAND2X1_182/CTRL 0.01fF
C46519 POR2X1_581/a_16_28# D_INPUT_6 0.04fF
C46520 POR2X1_344/Y POR2X1_349/Y 0.00fF
C46521 POR2X1_376/B POR2X1_701/CTRL 0.07fF
C46522 POR2X1_163/A PAND2X1_160/O 0.04fF
C46523 D_INPUT_6 PAND2X1_69/A 0.01fF
C46524 POR2X1_199/CTRL2 PAND2X1_824/B 0.06fF
C46525 POR2X1_9/Y POR2X1_88/A 0.00fF
C46526 POR2X1_590/A POR2X1_711/Y 0.14fF
C46527 POR2X1_16/A POR2X1_290/Y 0.03fF
C46528 PAND2X1_675/A POR2X1_437/CTRL2 0.00fF
C46529 PAND2X1_800/CTRL2 PAND2X1_863/B 0.01fF
C46530 PAND2X1_192/O PAND2X1_730/A 0.00fF
C46531 PAND2X1_850/Y PAND2X1_217/B 0.10fF
C46532 POR2X1_68/A POR2X1_845/O 0.01fF
C46533 POR2X1_130/A POR2X1_557/B 0.15fF
C46534 POR2X1_327/Y POR2X1_435/Y 0.10fF
C46535 POR2X1_35/Y POR2X1_854/B 0.05fF
C46536 POR2X1_502/A POR2X1_333/Y 0.00fF
C46537 PAND2X1_566/Y PAND2X1_854/A 0.03fF
C46538 PAND2X1_72/O PAND2X1_111/B 0.02fF
C46539 PAND2X1_474/Y POR2X1_150/CTRL2 0.00fF
C46540 PAND2X1_94/A PAND2X1_110/O 0.05fF
C46541 PAND2X1_137/Y POR2X1_103/CTRL 0.01fF
C46542 PAND2X1_213/Y POR2X1_73/Y 0.03fF
C46543 PAND2X1_354/O PAND2X1_854/A -0.00fF
C46544 POR2X1_394/A POR2X1_46/Y 0.24fF
C46545 PAND2X1_533/CTRL POR2X1_802/B 0.04fF
C46546 POR2X1_334/Y PAND2X1_257/CTRL 0.08fF
C46547 POR2X1_366/CTRL2 PAND2X1_6/Y 0.07fF
C46548 POR2X1_863/O POR2X1_260/A 0.02fF
C46549 POR2X1_356/O POR2X1_356/B 0.09fF
C46550 PAND2X1_90/A POR2X1_833/A 0.27fF
C46551 POR2X1_730/a_16_28# POR2X1_729/Y 0.05fF
C46552 POR2X1_383/A POR2X1_548/m4_208_n4# 0.07fF
C46553 PAND2X1_252/a_16_344# PAND2X1_60/B 0.03fF
C46554 POR2X1_68/B PAND2X1_111/B 0.01fF
C46555 PAND2X1_115/CTRL PAND2X1_348/A 0.04fF
C46556 PAND2X1_863/A PAND2X1_805/A 4.97fF
C46557 POR2X1_776/B POR2X1_566/CTRL2 0.03fF
C46558 POR2X1_123/A PAND2X1_518/CTRL 0.01fF
C46559 PAND2X1_317/Y PAND2X1_317/O 0.00fF
C46560 POR2X1_366/a_16_28# PAND2X1_48/B 0.01fF
C46561 POR2X1_16/A POR2X1_238/Y 0.10fF
C46562 PAND2X1_6/Y POR2X1_796/A 0.92fF
C46563 POR2X1_508/A PAND2X1_627/a_16_344# 0.02fF
C46564 PAND2X1_41/B POR2X1_383/Y 0.03fF
C46565 POR2X1_152/Y PAND2X1_731/A 0.01fF
C46566 POR2X1_391/O PAND2X1_32/B 0.16fF
C46567 INPUT_1 POR2X1_805/A 0.03fF
C46568 POR2X1_546/B POR2X1_546/a_16_28# 0.06fF
C46569 POR2X1_65/A PAND2X1_169/CTRL 0.01fF
C46570 VDD POR2X1_191/Y 2.61fF
C46571 POR2X1_114/B POR2X1_675/Y 0.02fF
C46572 VDD PAND2X1_199/CTRL 0.00fF
C46573 POR2X1_510/B PAND2X1_824/CTRL2 0.12fF
C46574 POR2X1_81/CTRL POR2X1_293/Y 0.03fF
C46575 POR2X1_540/CTRL POR2X1_181/B 0.01fF
C46576 POR2X1_584/O POR2X1_260/A 0.01fF
C46577 POR2X1_532/A POR2X1_101/Y 0.08fF
C46578 POR2X1_83/A POR2X1_83/a_16_28# 0.01fF
C46579 PAND2X1_596/CTRL POR2X1_761/A 0.01fF
C46580 PAND2X1_850/Y VDD -0.00fF
C46581 POR2X1_725/Y POR2X1_307/A 0.05fF
C46582 POR2X1_556/A POR2X1_658/CTRL2 0.04fF
C46583 POR2X1_532/A PAND2X1_690/CTRL2 0.03fF
C46584 POR2X1_41/B PAND2X1_476/A 0.02fF
C46585 PAND2X1_292/CTRL PAND2X1_41/B 0.01fF
C46586 POR2X1_85/Y POR2X1_230/CTRL2 0.01fF
C46587 PAND2X1_341/B PAND2X1_215/B 0.01fF
C46588 POR2X1_75/CTRL2 POR2X1_271/A 0.03fF
C46589 PAND2X1_187/CTRL POR2X1_568/Y 0.30fF
C46590 POR2X1_462/a_16_28# POR2X1_461/Y 0.05fF
C46591 POR2X1_119/Y POR2X1_494/Y 0.03fF
C46592 POR2X1_72/B PAND2X1_332/Y 0.03fF
C46593 POR2X1_244/Y PAND2X1_32/B 0.03fF
C46594 POR2X1_158/Y PAND2X1_712/CTRL2 0.00fF
C46595 POR2X1_98/B POR2X1_260/A 0.07fF
C46596 POR2X1_547/O POR2X1_266/A 0.01fF
C46597 POR2X1_648/Y POR2X1_655/A 0.05fF
C46598 POR2X1_416/B POR2X1_48/CTRL2 0.31fF
C46599 PAND2X1_55/Y POR2X1_188/Y 0.02fF
C46600 POR2X1_112/a_16_28# POR2X1_220/Y 0.01fF
C46601 POR2X1_532/A PAND2X1_533/CTRL 0.01fF
C46602 POR2X1_715/A POR2X1_702/A 0.38fF
C46603 POR2X1_505/CTRL2 POR2X1_245/Y 0.03fF
C46604 POR2X1_326/CTRL2 POR2X1_319/Y 0.03fF
C46605 D_GATE_741 POR2X1_294/A 0.02fF
C46606 PAND2X1_659/Y PAND2X1_218/O 0.01fF
C46607 POR2X1_274/B POR2X1_553/A 0.50fF
C46608 POR2X1_327/Y PAND2X1_96/B 0.07fF
C46609 POR2X1_556/A POR2X1_341/A 0.07fF
C46610 POR2X1_840/B POR2X1_186/B 0.06fF
C46611 POR2X1_267/Y PAND2X1_48/A 0.20fF
C46612 POR2X1_136/Y PAND2X1_715/B 0.73fF
C46613 POR2X1_809/A PAND2X1_583/O 0.02fF
C46614 POR2X1_306/a_16_28# PAND2X1_308/Y 0.07fF
C46615 PAND2X1_341/B PAND2X1_6/A 0.07fF
C46616 PAND2X1_350/O POR2X1_394/A 0.02fF
C46617 POR2X1_3/A POR2X1_3/B 0.10fF
C46618 POR2X1_369/Y PAND2X1_370/O -0.00fF
C46619 POR2X1_41/B PAND2X1_327/CTRL2 0.00fF
C46620 POR2X1_191/Y PAND2X1_32/B 0.05fF
C46621 PAND2X1_857/A PAND2X1_200/B 0.01fF
C46622 POR2X1_43/B PAND2X1_860/O 0.06fF
C46623 PAND2X1_841/CTRL POR2X1_39/B 0.01fF
C46624 POR2X1_192/Y POR2X1_181/Y 0.05fF
C46625 PAND2X1_60/O PAND2X1_39/B -0.00fF
C46626 PAND2X1_174/CTRL2 POR2X1_77/Y 0.04fF
C46627 POR2X1_49/O VDD 0.00fF
C46628 POR2X1_416/B POR2X1_763/Y 0.26fF
C46629 D_INPUT_3 POR2X1_5/O 0.01fF
C46630 PAND2X1_798/B POR2X1_184/O 0.01fF
C46631 POR2X1_575/a_76_344# POR2X1_574/Y 0.01fF
C46632 POR2X1_416/B PAND2X1_115/B 0.00fF
C46633 POR2X1_14/Y POR2X1_67/Y 0.03fF
C46634 POR2X1_737/O POR2X1_186/B 0.01fF
C46635 PAND2X1_404/A POR2X1_234/A 0.02fF
C46636 PAND2X1_497/CTRL POR2X1_624/Y 0.01fF
C46637 POR2X1_257/A PAND2X1_434/O 0.03fF
C46638 PAND2X1_632/B PAND2X1_156/A 0.05fF
C46639 POR2X1_416/B POR2X1_426/CTRL 0.01fF
C46640 POR2X1_158/Y POR2X1_426/CTRL2 0.00fF
C46641 POR2X1_158/CTRL POR2X1_425/Y 0.01fF
C46642 POR2X1_814/A POR2X1_750/B 0.17fF
C46643 POR2X1_353/A POR2X1_151/Y 0.01fF
C46644 POR2X1_461/CTRL POR2X1_814/A 0.01fF
C46645 PAND2X1_93/B POR2X1_602/O 0.01fF
C46646 PAND2X1_612/B POR2X1_476/A 0.03fF
C46647 POR2X1_67/Y POR2X1_849/CTRL2 0.03fF
C46648 POR2X1_416/B POR2X1_73/Y 0.21fF
C46649 POR2X1_326/A PAND2X1_533/O 0.17fF
C46650 PAND2X1_224/CTRL VDD -0.00fF
C46651 PAND2X1_681/CTRL2 PAND2X1_32/B 0.01fF
C46652 POR2X1_590/Y PAND2X1_48/A 0.11fF
C46653 POR2X1_846/Y POR2X1_750/B 0.03fF
C46654 PAND2X1_23/Y POR2X1_354/CTRL 0.00fF
C46655 POR2X1_567/B PAND2X1_237/CTRL 0.01fF
C46656 PAND2X1_834/CTRL PAND2X1_349/A 0.01fF
C46657 PAND2X1_826/CTRL POR2X1_838/B 0.00fF
C46658 POR2X1_796/Y POR2X1_811/A 0.01fF
C46659 POR2X1_647/B POR2X1_121/B 0.03fF
C46660 POR2X1_566/B POR2X1_568/B 0.02fF
C46661 POR2X1_180/A POR2X1_568/B 0.03fF
C46662 POR2X1_77/Y PAND2X1_348/Y 1.85fF
C46663 POR2X1_149/A POR2X1_149/a_16_28# 0.02fF
C46664 PAND2X1_714/Y PAND2X1_326/B 0.01fF
C46665 POR2X1_814/B PAND2X1_85/m4_208_n4# 0.15fF
C46666 POR2X1_68/B POR2X1_8/CTRL 0.03fF
C46667 POR2X1_635/a_16_28# POR2X1_750/B 0.02fF
C46668 PAND2X1_71/Y PAND2X1_527/O 0.02fF
C46669 POR2X1_88/CTRL POR2X1_14/Y 0.00fF
C46670 POR2X1_655/Y PAND2X1_39/B 0.10fF
C46671 POR2X1_191/O POR2X1_353/A 0.01fF
C46672 POR2X1_721/CTRL POR2X1_383/Y 0.01fF
C46673 POR2X1_424/Y POR2X1_423/Y 0.22fF
C46674 POR2X1_567/A POR2X1_326/A 0.03fF
C46675 POR2X1_281/CTRL2 POR2X1_416/B 0.01fF
C46676 POR2X1_261/A POR2X1_261/a_16_28# 0.03fF
C46677 POR2X1_760/A POR2X1_250/O 0.07fF
C46678 POR2X1_329/O POR2X1_250/Y 0.01fF
C46679 PAND2X1_20/A PAND2X1_609/a_76_28# 0.01fF
C46680 POR2X1_796/A PAND2X1_52/B -0.00fF
C46681 POR2X1_23/O POR2X1_37/Y 0.01fF
C46682 POR2X1_508/B POR2X1_508/A 0.18fF
C46683 POR2X1_609/Y PAND2X1_404/CTRL2 0.00fF
C46684 POR2X1_16/O POR2X1_73/Y 0.03fF
C46685 D_INPUT_5 POR2X1_25/CTRL2 0.03fF
C46686 PAND2X1_798/Y PAND2X1_366/O 0.10fF
C46687 PAND2X1_487/CTRL POR2X1_287/B 0.01fF
C46688 PAND2X1_235/O POR2X1_66/A 0.03fF
C46689 POR2X1_175/B PAND2X1_72/A 0.01fF
C46690 INPUT_3 PAND2X1_381/a_16_344# 0.01fF
C46691 POR2X1_862/B POR2X1_260/B 0.03fF
C46692 POR2X1_634/A POR2X1_637/CTRL 0.01fF
C46693 POR2X1_41/B POR2X1_263/CTRL 0.00fF
C46694 PAND2X1_208/O PAND2X1_124/Y 0.05fF
C46695 POR2X1_153/O POR2X1_416/B 0.04fF
C46696 PAND2X1_39/B POR2X1_206/A 0.12fF
C46697 POR2X1_472/B VDD 0.11fF
C46698 POR2X1_45/a_16_28# POR2X1_411/B 0.01fF
C46699 PAND2X1_402/CTRL2 D_INPUT_0 0.05fF
C46700 POR2X1_24/a_16_28# POR2X1_23/Y 0.05fF
C46701 POR2X1_508/B POR2X1_568/B 0.05fF
C46702 POR2X1_445/CTRL POR2X1_341/A 0.05fF
C46703 D_INPUT_3 POR2X1_9/Y 0.10fF
C46704 POR2X1_241/B POR2X1_254/CTRL2 0.01fF
C46705 POR2X1_850/B POR2X1_806/O 0.01fF
C46706 POR2X1_78/A POR2X1_794/B 0.03fF
C46707 POR2X1_157/CTRL2 POR2X1_257/A 0.03fF
C46708 POR2X1_866/A VDD 2.89fF
C46709 PAND2X1_457/O PAND2X1_464/B 0.06fF
C46710 PAND2X1_480/B PAND2X1_469/O 0.16fF
C46711 POR2X1_303/B POR2X1_260/A 0.01fF
C46712 POR2X1_288/A POR2X1_296/B 0.03fF
C46713 PAND2X1_476/A POR2X1_77/Y 0.01fF
C46714 PAND2X1_416/a_76_28# POR2X1_859/A 0.04fF
C46715 POR2X1_128/A PAND2X1_20/A 0.00fF
C46716 POR2X1_48/A PAND2X1_456/m4_208_n4# 0.09fF
C46717 D_INPUT_0 PAND2X1_206/CTRL2 0.05fF
C46718 POR2X1_83/B PAND2X1_208/O 0.04fF
C46719 PAND2X1_476/A POR2X1_85/Y 0.02fF
C46720 POR2X1_52/A PAND2X1_457/Y 0.06fF
C46721 POR2X1_66/O PAND2X1_69/A 0.01fF
C46722 POR2X1_78/CTRL POR2X1_78/Y 0.02fF
C46723 PAND2X1_43/m4_208_n4# PAND2X1_55/Y 0.12fF
C46724 PAND2X1_626/O POR2X1_852/B 0.17fF
C46725 POR2X1_462/B POR2X1_859/CTRL 0.01fF
C46726 POR2X1_42/CTRL2 POR2X1_20/B 0.01fF
C46727 POR2X1_189/Y POR2X1_679/A 0.00fF
C46728 PAND2X1_286/CTRL POR2X1_283/Y 0.01fF
C46729 PAND2X1_405/CTRL PAND2X1_737/B 0.01fF
C46730 POR2X1_23/Y PAND2X1_468/O 0.01fF
C46731 POR2X1_66/B POR2X1_286/Y 0.01fF
C46732 POR2X1_777/B PAND2X1_46/O 0.01fF
C46733 PAND2X1_381/Y VDD 0.01fF
C46734 POR2X1_54/Y POR2X1_793/A 0.01fF
C46735 POR2X1_439/O PAND2X1_41/B 0.15fF
C46736 POR2X1_852/B POR2X1_750/B 0.07fF
C46737 POR2X1_251/A PAND2X1_562/B 0.03fF
C46738 PAND2X1_48/B PAND2X1_59/B 0.12fF
C46739 POR2X1_78/B POR2X1_850/B 0.12fF
C46740 POR2X1_636/CTRL VDD 0.00fF
C46741 POR2X1_65/A POR2X1_331/Y 0.03fF
C46742 PAND2X1_284/Y POR2X1_411/B 0.03fF
C46743 POR2X1_490/Y POR2X1_45/Y 0.03fF
C46744 POR2X1_689/A POR2X1_48/A 0.01fF
C46745 POR2X1_856/B POR2X1_149/Y 0.01fF
C46746 PAND2X1_678/CTRL2 PAND2X1_175/B 0.01fF
C46747 PAND2X1_831/a_16_344# PAND2X1_217/B 0.12fF
C46748 PAND2X1_841/O POR2X1_23/Y 0.07fF
C46749 PAND2X1_540/CTRL2 POR2X1_106/Y 0.01fF
C46750 POR2X1_40/Y POR2X1_5/Y 0.08fF
C46751 PAND2X1_48/B POR2X1_610/a_16_28# 0.03fF
C46752 POR2X1_502/A POR2X1_174/A 0.03fF
C46753 POR2X1_669/B POR2X1_46/Y 0.29fF
C46754 PAND2X1_65/B PAND2X1_46/O 0.03fF
C46755 POR2X1_60/A POR2X1_481/A 0.04fF
C46756 POR2X1_43/B PAND2X1_124/Y 0.04fF
C46757 PAND2X1_23/Y POR2X1_66/A 0.19fF
C46758 POR2X1_496/Y POR2X1_7/B 0.07fF
C46759 POR2X1_65/A POR2X1_517/O 0.02fF
C46760 POR2X1_344/O PAND2X1_65/B 0.16fF
C46761 PAND2X1_109/m4_208_n4# POR2X1_78/A 0.09fF
C46762 POR2X1_76/A PAND2X1_311/CTRL2 0.01fF
C46763 POR2X1_811/B POR2X1_779/m4_208_n4# 0.09fF
C46764 PAND2X1_738/B PAND2X1_738/O 0.00fF
C46765 POR2X1_672/Y POR2X1_38/B 0.01fF
C46766 POR2X1_260/a_56_344# POR2X1_260/A 0.00fF
C46767 POR2X1_78/Y POR2X1_569/A 0.02fF
C46768 POR2X1_502/A POR2X1_375/Y 0.00fF
C46769 PAND2X1_474/Y POR2X1_72/B 0.01fF
C46770 POR2X1_72/Y PAND2X1_657/CTRL 0.02fF
C46771 POR2X1_71/Y PAND2X1_657/O 0.04fF
C46772 POR2X1_23/Y PAND2X1_726/m4_208_n4# 0.08fF
C46773 POR2X1_287/B POR2X1_362/B 0.03fF
C46774 POR2X1_866/A PAND2X1_32/B 0.07fF
C46775 POR2X1_269/CTRL2 POR2X1_741/Y 0.09fF
C46776 POR2X1_269/O POR2X1_740/Y 0.02fF
C46777 PAND2X1_223/B POR2X1_42/Y 0.03fF
C46778 POR2X1_97/A POR2X1_350/CTRL 0.00fF
C46779 POR2X1_628/Y POR2X1_245/Y 0.03fF
C46780 POR2X1_590/A POR2X1_733/A 0.03fF
C46781 POR2X1_462/CTRL2 POR2X1_559/A 0.00fF
C46782 PAND2X1_211/A VDD 0.30fF
C46783 PAND2X1_230/CTRL2 POR2X1_785/A 0.00fF
C46784 POR2X1_33/A D_INPUT_1 0.01fF
C46785 POR2X1_13/A POR2X1_72/B 5.06fF
C46786 POR2X1_547/CTRL2 POR2X1_78/A 0.03fF
C46787 POR2X1_705/B POR2X1_260/A 0.06fF
C46788 POR2X1_383/A POR2X1_647/B 3.45fF
C46789 PAND2X1_48/B PAND2X1_594/a_76_28# 0.01fF
C46790 PAND2X1_648/Y PAND2X1_655/B 0.01fF
C46791 POR2X1_121/CTRL POR2X1_260/B 0.01fF
C46792 POR2X1_96/A PAND2X1_217/B 0.06fF
C46793 PAND2X1_57/B POR2X1_734/A 0.08fF
C46794 POR2X1_659/A POR2X1_222/A 3.88fF
C46795 POR2X1_750/B INPUT_5 0.07fF
C46796 PAND2X1_733/A POR2X1_7/B 0.00fF
C46797 PAND2X1_866/A PAND2X1_288/A 0.10fF
C46798 POR2X1_263/Y PAND2X1_734/a_16_344# 0.01fF
C46799 POR2X1_260/B POR2X1_510/Y 0.03fF
C46800 POR2X1_245/m4_208_n4# POR2X1_245/Y 0.07fF
C46801 POR2X1_496/CTRL POR2X1_789/B 0.00fF
C46802 POR2X1_14/Y POR2X1_586/m4_208_n4# 0.01fF
C46803 POR2X1_207/A VDD 0.23fF
C46804 POR2X1_31/CTRL POR2X1_12/A 0.00fF
C46805 POR2X1_43/B POR2X1_83/B 0.53fF
C46806 PAND2X1_73/O POR2X1_294/B 0.14fF
C46807 POR2X1_860/CTRL PAND2X1_39/B 0.12fF
C46808 POR2X1_840/O D_INPUT_0 0.01fF
C46809 POR2X1_667/A POR2X1_519/Y 0.87fF
C46810 POR2X1_514/CTRL PAND2X1_20/A 0.01fF
C46811 POR2X1_814/B POR2X1_471/a_16_28# 0.03fF
C46812 INPUT_1 PAND2X1_39/B 0.01fF
C46813 POR2X1_307/Y POR2X1_807/A 0.02fF
C46814 POR2X1_499/m4_208_n4# POR2X1_576/Y 0.01fF
C46815 PAND2X1_20/A PAND2X1_519/O 0.04fF
C46816 PAND2X1_793/Y PAND2X1_805/A 0.02fF
C46817 POR2X1_63/a_16_28# POR2X1_669/B 0.02fF
C46818 POR2X1_416/Y POR2X1_607/A 0.01fF
C46819 POR2X1_642/CTRL2 POR2X1_734/A 0.03fF
C46820 POR2X1_54/Y POR2X1_753/CTRL2 0.04fF
C46821 POR2X1_272/a_56_344# POR2X1_42/Y 0.00fF
C46822 POR2X1_481/Y PAND2X1_354/A 0.03fF
C46823 POR2X1_78/A POR2X1_570/B 0.03fF
C46824 POR2X1_135/Y PAND2X1_480/B 0.05fF
C46825 POR2X1_302/Y VDD 0.29fF
C46826 PAND2X1_821/CTRL PAND2X1_41/B 0.03fF
C46827 POR2X1_52/A PAND2X1_736/CTRL 0.01fF
C46828 POR2X1_628/Y PAND2X1_507/CTRL 0.00fF
C46829 POR2X1_114/B POR2X1_405/CTRL 0.01fF
C46830 POR2X1_287/B PAND2X1_371/a_16_344# 0.01fF
C46831 POR2X1_458/O POR2X1_101/Y 0.02fF
C46832 PAND2X1_777/O POR2X1_387/Y 0.05fF
C46833 POR2X1_130/A PAND2X1_56/CTRL 0.01fF
C46834 POR2X1_83/B POR2X1_38/B 0.03fF
C46835 POR2X1_294/O POR2X1_507/A 0.03fF
C46836 PAND2X1_843/CTRL PAND2X1_675/A 0.02fF
C46837 PAND2X1_63/O PAND2X1_63/B 0.04fF
C46838 POR2X1_123/B POR2X1_78/A 0.00fF
C46839 POR2X1_368/Y POR2X1_417/Y 0.05fF
C46840 POR2X1_96/A VDD 3.70fF
C46841 POR2X1_66/B POR2X1_649/CTRL2 0.00fF
C46842 PAND2X1_90/A PAND2X1_412/a_16_344# 0.02fF
C46843 PAND2X1_651/Y PAND2X1_465/CTRL 0.00fF
C46844 POR2X1_66/B PAND2X1_69/A 2.31fF
C46845 POR2X1_60/A PAND2X1_645/B 0.02fF
C46846 POR2X1_13/A PAND2X1_768/CTRL 0.01fF
C46847 POR2X1_707/B POR2X1_407/Y 0.02fF
C46848 PAND2X1_209/A PAND2X1_161/O 0.03fF
C46849 POR2X1_141/Y POR2X1_513/Y 0.03fF
C46850 POR2X1_14/Y POR2X1_750/CTRL 0.00fF
C46851 POR2X1_40/Y POR2X1_310/O 0.04fF
C46852 POR2X1_480/A POR2X1_294/B 0.10fF
C46853 PAND2X1_92/O INPUT_0 0.17fF
C46854 POR2X1_257/A PAND2X1_508/Y 0.06fF
C46855 PAND2X1_738/Y PAND2X1_544/m4_208_n4# 0.04fF
C46856 POR2X1_614/A POR2X1_593/B 0.03fF
C46857 POR2X1_388/CTRL2 POR2X1_814/B 0.03fF
C46858 POR2X1_188/A PAND2X1_69/A 0.10fF
C46859 PAND2X1_661/B POR2X1_72/B 0.05fF
C46860 POR2X1_123/A PAND2X1_73/Y 0.19fF
C46861 POR2X1_207/A POR2X1_741/Y 0.05fF
C46862 POR2X1_9/Y PAND2X1_52/B 0.15fF
C46863 POR2X1_464/O PAND2X1_55/Y 0.01fF
C46864 PAND2X1_61/Y POR2X1_521/O 0.01fF
C46865 POR2X1_596/A POR2X1_330/Y 0.05fF
C46866 PAND2X1_206/B PAND2X1_358/O 0.00fF
C46867 PAND2X1_738/Y POR2X1_763/Y 0.04fF
C46868 POR2X1_257/A POR2X1_320/CTRL 0.01fF
C46869 PAND2X1_848/B POR2X1_5/Y 0.03fF
C46870 POR2X1_81/Y PAND2X1_573/a_16_344# 0.05fF
C46871 PAND2X1_207/CTRL2 PAND2X1_123/Y 0.01fF
C46872 POR2X1_549/A POR2X1_549/a_16_28# 0.02fF
C46873 POR2X1_188/A POR2X1_710/a_16_28# 0.01fF
C46874 POR2X1_61/Y POR2X1_631/B 0.07fF
C46875 PAND2X1_23/Y PAND2X1_293/O 0.00fF
C46876 POR2X1_566/A PAND2X1_441/O 0.03fF
C46877 POR2X1_88/Y POR2X1_42/Y 0.05fF
C46878 POR2X1_719/B POR2X1_66/A 0.00fF
C46879 POR2X1_777/B POR2X1_318/A 0.10fF
C46880 POR2X1_566/A POR2X1_740/Y 0.03fF
C46881 PAND2X1_434/CTRL POR2X1_83/B 0.01fF
C46882 PAND2X1_842/CTRL2 PAND2X1_389/Y 0.03fF
C46883 PAND2X1_280/CTRL PAND2X1_55/Y 0.01fF
C46884 POR2X1_186/Y PAND2X1_747/O 0.04fF
C46885 POR2X1_131/CTRL2 PAND2X1_140/Y 0.03fF
C46886 POR2X1_68/A PAND2X1_293/CTRL 0.03fF
C46887 POR2X1_448/B POR2X1_788/B 0.04fF
C46888 PAND2X1_659/Y PAND2X1_205/CTRL 0.03fF
C46889 POR2X1_416/B PAND2X1_780/O 0.05fF
C46890 POR2X1_166/a_16_28# POR2X1_40/Y 0.09fF
C46891 POR2X1_141/Y POR2X1_366/A 0.03fF
C46892 PAND2X1_813/CTRL POR2X1_78/A 0.01fF
C46893 POR2X1_272/O PAND2X1_349/A 0.01fF
C46894 POR2X1_333/A POR2X1_326/CTRL2 0.08fF
C46895 POR2X1_68/A POR2X1_404/B 0.01fF
C46896 POR2X1_523/Y POR2X1_859/A 0.01fF
C46897 POR2X1_68/A PAND2X1_524/CTRL2 0.01fF
C46898 POR2X1_60/A PAND2X1_737/B 0.03fF
C46899 POR2X1_516/B POR2X1_56/Y 0.03fF
C46900 POR2X1_102/Y PAND2X1_861/O 0.01fF
C46901 POR2X1_489/B POR2X1_260/A 0.02fF
C46902 PAND2X1_742/B PAND2X1_592/Y 0.03fF
C46903 POR2X1_599/A PAND2X1_198/m4_208_n4# 0.06fF
C46904 INPUT_1 PAND2X1_20/A 0.06fF
C46905 PAND2X1_520/O PAND2X1_642/B 0.02fF
C46906 POR2X1_66/B PAND2X1_765/a_76_28# 0.02fF
C46907 PAND2X1_90/A POR2X1_294/B 0.19fF
C46908 POR2X1_744/Y POR2X1_39/B 0.01fF
C46909 POR2X1_356/A D_GATE_662 0.10fF
C46910 PAND2X1_216/B POR2X1_60/A 0.03fF
C46911 POR2X1_72/B PAND2X1_510/B 0.01fF
C46912 PAND2X1_65/B POR2X1_318/A 0.07fF
C46913 POR2X1_16/A PAND2X1_195/CTRL2 -0.03fF
C46914 POR2X1_508/CTRL POR2X1_579/Y 0.00fF
C46915 PAND2X1_540/CTRL2 PAND2X1_114/B 0.04fF
C46916 VDD POR2X1_501/B 0.28fF
C46917 PAND2X1_771/Y POR2X1_766/Y 0.16fF
C46918 PAND2X1_57/B POR2X1_786/Y 0.07fF
C46919 PAND2X1_480/B POR2X1_816/A 0.05fF
C46920 POR2X1_302/Y PAND2X1_32/B 0.01fF
C46921 POR2X1_178/Y POR2X1_40/Y 0.02fF
C46922 POR2X1_582/a_16_28# INPUT_7 0.03fF
C46923 PAND2X1_734/B POR2X1_229/CTRL 0.01fF
C46924 PAND2X1_57/B PAND2X1_69/CTRL 0.01fF
C46925 POR2X1_332/B POR2X1_702/A 0.29fF
C46926 POR2X1_143/O PAND2X1_6/A 0.04fF
C46927 POR2X1_330/Y POR2X1_598/O 0.02fF
C46928 PAND2X1_738/Y POR2X1_73/Y 0.05fF
C46929 POR2X1_100/CTRL2 POR2X1_243/Y 0.03fF
C46930 PAND2X1_80/CTRL2 PAND2X1_111/B 0.01fF
C46931 PAND2X1_23/Y POR2X1_222/Y 0.06fF
C46932 PAND2X1_48/B D_GATE_222 0.03fF
C46933 PAND2X1_865/Y PAND2X1_773/Y 0.23fF
C46934 POR2X1_327/a_16_28# POR2X1_572/B 0.03fF
C46935 VDD POR2X1_689/Y 0.00fF
C46936 POR2X1_66/B PAND2X1_824/B 0.07fF
C46937 PAND2X1_230/CTRL2 POR2X1_186/B 0.09fF
C46938 POR2X1_780/CTRL POR2X1_260/A 0.01fF
C46939 POR2X1_234/O POR2X1_293/Y 0.16fF
C46940 PAND2X1_350/CTRL2 INPUT_0 0.06fF
C46941 POR2X1_435/O POR2X1_513/B 0.01fF
C46942 POR2X1_390/B PAND2X1_41/B 0.03fF
C46943 PAND2X1_254/CTRL2 POR2X1_253/Y 0.10fF
C46944 PAND2X1_556/B POR2X1_91/Y 0.03fF
C46945 POR2X1_136/m4_208_n4# PAND2X1_480/B 0.04fF
C46946 PAND2X1_20/A PAND2X1_586/CTRL 0.00fF
C46947 PAND2X1_494/O POR2X1_294/B 0.05fF
C46948 POR2X1_76/Y POR2X1_573/A 0.01fF
C46949 PAND2X1_494/CTRL POR2X1_264/Y 0.01fF
C46950 PAND2X1_220/CTRL2 PAND2X1_566/Y 0.00fF
C46951 POR2X1_740/Y PAND2X1_111/O 0.15fF
C46952 PAND2X1_707/Y PAND2X1_705/O 0.01fF
C46953 PAND2X1_492/CTRL POR2X1_123/A 0.01fF
C46954 PAND2X1_661/Y POR2X1_236/Y 0.07fF
C46955 POR2X1_634/A POR2X1_774/A 0.19fF
C46956 INPUT_1 POR2X1_814/B 0.16fF
C46957 POR2X1_7/A VDD 3.19fF
C46958 POR2X1_614/A POR2X1_477/A 0.01fF
C46959 POR2X1_509/A POR2X1_35/Y 0.03fF
C46960 POR2X1_193/CTRL POR2X1_631/B 0.03fF
C46961 POR2X1_130/A POR2X1_361/a_16_28# 0.03fF
C46962 PAND2X1_675/A PAND2X1_566/Y 0.07fF
C46963 POR2X1_174/A POR2X1_188/Y 0.03fF
C46964 POR2X1_16/A POR2X1_689/CTRL2 0.01fF
C46965 POR2X1_78/B POR2X1_317/A 0.25fF
C46966 PAND2X1_278/CTRL POR2X1_559/A 0.00fF
C46967 POR2X1_49/O PAND2X1_9/Y 0.01fF
C46968 POR2X1_205/A POR2X1_404/Y 0.07fF
C46969 PAND2X1_660/Y VDD -0.00fF
C46970 POR2X1_43/Y PAND2X1_838/B 1.65fF
C46971 POR2X1_776/A POR2X1_568/A 0.06fF
C46972 PAND2X1_23/Y POR2X1_532/A 9.00fF
C46973 PAND2X1_684/CTRL PAND2X1_90/Y 0.16fF
C46974 POR2X1_809/A POR2X1_866/a_76_344# 0.00fF
C46975 POR2X1_740/Y POR2X1_573/A 0.03fF
C46976 POR2X1_35/Y POR2X1_631/B 0.03fF
C46977 POR2X1_703/A VDD 0.35fF
C46978 POR2X1_78/B POR2X1_339/CTRL 0.00fF
C46979 POR2X1_121/CTRL PAND2X1_55/Y 0.03fF
C46980 PAND2X1_90/A PAND2X1_111/B 0.07fF
C46981 POR2X1_74/Y PAND2X1_76/CTRL 0.01fF
C46982 POR2X1_451/A POR2X1_635/O 0.01fF
C46983 POR2X1_566/A PAND2X1_253/CTRL 0.01fF
C46984 POR2X1_413/A PAND2X1_647/CTRL2 0.01fF
C46985 PAND2X1_499/Y PAND2X1_861/a_56_28# 0.00fF
C46986 POR2X1_407/A POR2X1_68/B 0.00fF
C46987 POR2X1_66/A POR2X1_711/Y 0.23fF
C46988 PAND2X1_6/Y PAND2X1_424/CTRL2 0.00fF
C46989 PAND2X1_55/Y POR2X1_510/Y 0.03fF
C46990 POR2X1_356/A POR2X1_356/B 0.06fF
C46991 PAND2X1_93/a_16_344# PAND2X1_88/Y 0.00fF
C46992 POR2X1_311/O POR2X1_7/B 0.18fF
C46993 PAND2X1_691/a_76_28# POR2X1_689/Y 0.02fF
C46994 D_INPUT_0 PAND2X1_339/a_16_344# 0.05fF
C46995 POR2X1_7/B POR2X1_375/CTRL 0.01fF
C46996 POR2X1_501/B PAND2X1_32/B 0.03fF
C46997 PAND2X1_736/A POR2X1_283/A 0.07fF
C46998 POR2X1_68/A PAND2X1_177/a_76_28# 0.02fF
C46999 POR2X1_72/B PAND2X1_199/O 0.01fF
C47000 POR2X1_327/Y POR2X1_302/O 0.01fF
C47001 POR2X1_440/Y POR2X1_477/A 0.03fF
C47002 PAND2X1_658/B PAND2X1_549/B 0.03fF
C47003 POR2X1_449/A POR2X1_449/a_16_28# 0.03fF
C47004 POR2X1_22/a_76_344# POR2X1_260/A 0.00fF
C47005 POR2X1_130/A POR2X1_774/A 0.07fF
C47006 POR2X1_351/B VDD 0.19fF
C47007 D_INPUT_3 INPUT_2 0.14fF
C47008 VDD POR2X1_384/Y 0.00fF
C47009 POR2X1_346/B POR2X1_294/B 0.05fF
C47010 PAND2X1_797/Y PAND2X1_738/B 0.09fF
C47011 POR2X1_539/CTRL POR2X1_741/Y 0.00fF
C47012 POR2X1_614/A PAND2X1_158/O 0.17fF
C47013 POR2X1_255/CTRL2 PAND2X1_840/Y 0.03fF
C47014 POR2X1_741/Y POR2X1_703/A 0.47fF
C47015 POR2X1_732/B POR2X1_675/Y 0.33fF
C47016 POR2X1_8/Y POR2X1_42/Y 0.08fF
C47017 PAND2X1_88/Y PAND2X1_60/B 0.03fF
C47018 D_INPUT_1 POR2X1_569/A 0.07fF
C47019 POR2X1_84/Y PAND2X1_60/B 0.51fF
C47020 POR2X1_268/Y POR2X1_39/B 0.01fF
C47021 POR2X1_383/A POR2X1_203/Y 0.05fF
C47022 INPUT_1 POR2X1_32/a_16_28# 0.01fF
C47023 POR2X1_411/B PAND2X1_269/O 0.03fF
C47024 PAND2X1_804/CTRL2 PAND2X1_860/A 0.01fF
C47025 POR2X1_110/O POR2X1_13/A 0.18fF
C47026 POR2X1_860/O POR2X1_218/A 0.02fF
C47027 POR2X1_278/Y POR2X1_187/Y 0.03fF
C47028 PAND2X1_649/A PAND2X1_688/O 0.01fF
C47029 PAND2X1_61/Y POR2X1_39/B 0.03fF
C47030 POR2X1_544/B POR2X1_732/B 0.10fF
C47031 POR2X1_219/B POR2X1_215/A 0.12fF
C47032 POR2X1_72/B POR2X1_387/O 0.01fF
C47033 POR2X1_832/A POR2X1_513/O 0.02fF
C47034 POR2X1_569/A POR2X1_724/A 0.14fF
C47035 PAND2X1_414/CTRL2 INPUT_3 0.01fF
C47036 PAND2X1_96/B POR2X1_249/Y 0.02fF
C47037 PAND2X1_467/Y POR2X1_425/Y 0.05fF
C47038 PAND2X1_21/CTRL2 D_INPUT_4 0.00fF
C47039 POR2X1_141/CTRL2 POR2X1_343/Y 0.02fF
C47040 POR2X1_257/A PAND2X1_464/B 0.14fF
C47041 POR2X1_609/Y PAND2X1_403/CTRL 0.00fF
C47042 POR2X1_813/Y POR2X1_7/A 0.01fF
C47043 POR2X1_385/Y POR2X1_42/Y 0.05fF
C47044 POR2X1_336/a_16_28# POR2X1_703/A 0.03fF
C47045 POR2X1_121/A PAND2X1_48/A 0.03fF
C47046 PAND2X1_312/O POR2X1_703/A 0.02fF
C47047 POR2X1_467/Y POR2X1_863/A 0.03fF
C47048 POR2X1_702/CTRL POR2X1_260/A 0.13fF
C47049 PAND2X1_484/O PAND2X1_69/A 0.01fF
C47050 POR2X1_779/A POR2X1_294/A 0.03fF
C47051 PAND2X1_341/A PAND2X1_358/A 0.33fF
C47052 POR2X1_90/Y PAND2X1_156/A 0.07fF
C47053 POR2X1_673/Y POR2X1_7/A 0.03fF
C47054 POR2X1_844/B POR2X1_550/B 0.67fF
C47055 POR2X1_319/a_16_28# POR2X1_191/Y 0.04fF
C47056 POR2X1_652/O POR2X1_652/A 0.00fF
C47057 PAND2X1_865/Y PAND2X1_575/A 0.00fF
C47058 POR2X1_616/Y POR2X1_617/a_16_28# 0.03fF
C47059 POR2X1_834/Y POR2X1_513/m4_208_n4# 0.04fF
C47060 POR2X1_48/A POR2X1_600/O 0.16fF
C47061 PAND2X1_440/CTRL2 PAND2X1_793/Y 0.01fF
C47062 POR2X1_416/B PAND2X1_785/Y 0.03fF
C47063 PAND2X1_39/B PAND2X1_43/O 0.04fF
C47064 PAND2X1_352/CTRL PAND2X1_357/Y 0.01fF
C47065 POR2X1_809/A POR2X1_532/A 0.00fF
C47066 POR2X1_411/B PAND2X1_222/A 0.01fF
C47067 PAND2X1_865/Y PAND2X1_794/B 0.00fF
C47068 POR2X1_703/A POR2X1_543/CTRL2 0.04fF
C47069 POR2X1_147/CTRL POR2X1_435/Y 0.06fF
C47070 PAND2X1_476/A POR2X1_52/Y 0.03fF
C47071 D_INPUT_6 PAND2X1_3/B 0.03fF
C47072 PAND2X1_501/CTRL POR2X1_494/Y 0.00fF
C47073 POR2X1_46/Y PAND2X1_327/O 0.05fF
C47074 POR2X1_628/a_56_344# POR2X1_39/B 0.00fF
C47075 POR2X1_168/A POR2X1_776/B 0.00fF
C47076 POR2X1_20/B POR2X1_612/Y 0.07fF
C47077 POR2X1_303/CTRL2 POR2X1_228/Y 0.01fF
C47078 POR2X1_60/Y POR2X1_9/Y 0.04fF
C47079 POR2X1_43/B PAND2X1_841/Y 0.02fF
C47080 POR2X1_824/O POR2X1_824/Y 0.01fF
C47081 PAND2X1_804/B POR2X1_173/a_16_28# 0.08fF
C47082 POR2X1_186/CTRL2 POR2X1_186/B 0.03fF
C47083 POR2X1_68/B PAND2X1_517/a_16_344# 0.02fF
C47084 PAND2X1_731/CTRL POR2X1_39/B 0.01fF
C47085 POR2X1_556/A POR2X1_269/CTRL 0.01fF
C47086 PAND2X1_59/CTRL2 D_INPUT_4 0.00fF
C47087 POR2X1_863/A POR2X1_570/O 0.11fF
C47088 PAND2X1_860/A INPUT_0 0.03fF
C47089 POR2X1_83/B PAND2X1_201/CTRL2 0.03fF
C47090 POR2X1_394/A POR2X1_744/a_16_28# 0.01fF
C47091 POR2X1_9/Y POR2X1_625/O 0.17fF
C47092 POR2X1_411/B POR2X1_432/CTRL 0.01fF
C47093 D_GATE_662 PAND2X1_72/A 0.12fF
C47094 POR2X1_99/B POR2X1_259/CTRL2 0.00fF
C47095 POR2X1_814/A POR2X1_389/Y 0.02fF
C47096 PAND2X1_64/O PAND2X1_26/A 0.02fF
C47097 PAND2X1_367/A PAND2X1_367/O 0.01fF
C47098 POR2X1_327/Y POR2X1_860/a_16_28# 0.01fF
C47099 POR2X1_772/O POR2X1_294/A 0.05fF
C47100 PAND2X1_601/CTRL POR2X1_66/A 0.01fF
C47101 POR2X1_78/B POR2X1_98/A 1.05fF
C47102 POR2X1_532/A POR2X1_711/Y 0.02fF
C47103 POR2X1_67/Y PAND2X1_793/A 0.01fF
C47104 POR2X1_394/A PAND2X1_708/O 0.02fF
C47105 POR2X1_760/A PAND2X1_217/B 0.08fF
C47106 POR2X1_146/O PAND2X1_797/Y 0.01fF
C47107 POR2X1_346/B POR2X1_567/A 0.03fF
C47108 PAND2X1_404/Y POR2X1_37/Y 0.07fF
C47109 POR2X1_88/A POR2X1_69/A 0.02fF
C47110 D_INPUT_1 PAND2X1_72/A 0.03fF
C47111 PAND2X1_518/O PAND2X1_52/B 0.06fF
C47112 POR2X1_114/a_16_28# POR2X1_717/B 0.01fF
C47113 POR2X1_633/a_56_344# POR2X1_734/A 0.03fF
C47114 POR2X1_688/Y POR2X1_121/B 0.13fF
C47115 POR2X1_800/CTRL2 POR2X1_452/Y 0.01fF
C47116 POR2X1_383/A POR2X1_343/a_76_344# 0.00fF
C47117 POR2X1_416/B PAND2X1_656/A 0.07fF
C47118 POR2X1_41/B POR2X1_827/CTRL2 0.01fF
C47119 POR2X1_577/CTRL POR2X1_568/A 0.03fF
C47120 INPUT_3 POR2X1_293/CTRL2 0.01fF
C47121 PAND2X1_189/O POR2X1_188/Y 0.00fF
C47122 POR2X1_811/O D_INPUT_0 0.16fF
C47123 PAND2X1_620/Y POR2X1_20/B 0.03fF
C47124 POR2X1_291/CTRL2 POR2X1_39/B 0.00fF
C47125 PAND2X1_824/B POR2X1_199/B 0.02fF
C47126 POR2X1_422/O POR2X1_422/Y 0.01fF
C47127 POR2X1_466/A POR2X1_434/A 0.25fF
C47128 POR2X1_582/Y POR2X1_748/A 0.22fF
C47129 POR2X1_65/A POR2X1_20/B 1.25fF
C47130 POR2X1_294/A POR2X1_113/B 0.03fF
C47131 POR2X1_475/O POR2X1_288/A 0.00fF
C47132 POR2X1_568/B POR2X1_353/A 0.05fF
C47133 POR2X1_760/A VDD 1.65fF
C47134 POR2X1_801/CTRL POR2X1_452/Y 0.01fF
C47135 POR2X1_176/Y POR2X1_77/Y 0.01fF
C47136 POR2X1_455/CTRL2 POR2X1_341/A 0.06fF
C47137 PAND2X1_47/B PAND2X1_25/CTRL2 0.01fF
C47138 PAND2X1_120/CTRL2 POR2X1_77/Y 0.00fF
C47139 POR2X1_416/B PAND2X1_348/A 0.89fF
C47140 PAND2X1_20/A POR2X1_637/O 0.00fF
C47141 PAND2X1_96/B POR2X1_643/O 0.10fF
C47142 POR2X1_23/Y PAND2X1_658/O 0.04fF
C47143 PAND2X1_717/A PAND2X1_303/a_76_28# 0.01fF
C47144 POR2X1_45/Y POR2X1_329/A 0.03fF
C47145 PAND2X1_466/B VDD 0.00fF
C47146 D_INPUT_0 POR2X1_330/Y 0.05fF
C47147 PAND2X1_415/O VDD 0.00fF
C47148 POR2X1_811/A POR2X1_330/Y 0.05fF
C47149 PAND2X1_48/B PAND2X1_417/CTRL 0.01fF
C47150 POR2X1_96/A PAND2X1_9/Y 0.03fF
C47151 PAND2X1_699/CTRL2 POR2X1_43/B 0.09fF
C47152 POR2X1_554/B POR2X1_572/B 0.06fF
C47153 POR2X1_376/B PAND2X1_99/B 0.01fF
C47154 POR2X1_496/Y POR2X1_750/B 0.07fF
C47155 PAND2X1_58/O POR2X1_202/A 0.12fF
C47156 PAND2X1_578/Y PAND2X1_580/B 0.03fF
C47157 POR2X1_272/O POR2X1_32/A 0.01fF
C47158 PAND2X1_635/Y POR2X1_408/Y 0.12fF
C47159 POR2X1_855/CTRL2 POR2X1_855/A 0.00fF
C47160 PAND2X1_390/Y POR2X1_32/A 0.03fF
C47161 POR2X1_49/Y POR2X1_751/A 0.01fF
C47162 POR2X1_52/A POR2X1_415/A 0.61fF
C47163 POR2X1_168/A POR2X1_192/B 0.05fF
C47164 POR2X1_525/Y POR2X1_257/A 0.03fF
C47165 POR2X1_117/a_16_28# POR2X1_409/B 0.02fF
C47166 POR2X1_792/CTRL2 PAND2X1_90/Y 0.10fF
C47167 POR2X1_376/B POR2X1_432/CTRL 0.06fF
C47168 POR2X1_814/A POR2X1_318/A 0.07fF
C47169 PAND2X1_48/B POR2X1_54/Y 0.20fF
C47170 PAND2X1_631/A POR2X1_416/B 0.68fF
C47171 PAND2X1_75/CTRL POR2X1_318/A 0.04fF
C47172 PAND2X1_68/a_76_28# POR2X1_5/Y 0.01fF
C47173 POR2X1_66/B POR2X1_640/Y 0.06fF
C47174 POR2X1_294/A POR2X1_768/A 0.08fF
C47175 PAND2X1_836/CTRL2 POR2X1_20/B 0.01fF
C47176 POR2X1_814/A POR2X1_713/B 0.05fF
C47177 POR2X1_68/A POR2X1_663/B 0.03fF
C47178 POR2X1_84/B POR2X1_294/B 0.02fF
C47179 PAND2X1_404/Y POR2X1_293/Y 0.11fF
C47180 PAND2X1_640/B POR2X1_13/A 0.07fF
C47181 POR2X1_846/CTRL POR2X1_129/Y 0.01fF
C47182 POR2X1_579/B POR2X1_579/a_16_28# 0.07fF
C47183 PAND2X1_487/O POR2X1_294/B 0.05fF
C47184 PAND2X1_832/a_76_28# PAND2X1_435/Y 0.01fF
C47185 POR2X1_709/A PAND2X1_411/a_16_344# 0.03fF
C47186 POR2X1_407/A PAND2X1_761/O 0.04fF
C47187 PAND2X1_203/O POR2X1_816/A 0.01fF
C47188 PAND2X1_695/O PAND2X1_11/Y 0.01fF
C47189 POR2X1_632/CTRL2 POR2X1_222/Y 0.10fF
C47190 POR2X1_132/Y POR2X1_20/B 0.11fF
C47191 POR2X1_68/A PAND2X1_826/O 0.00fF
C47192 PAND2X1_246/CTRL PAND2X1_63/B 0.01fF
C47193 POR2X1_639/A POR2X1_750/B 0.54fF
C47194 POR2X1_416/B POR2X1_43/CTRL 0.00fF
C47195 POR2X1_851/A POR2X1_733/A 0.04fF
C47196 POR2X1_658/CTRL2 PAND2X1_60/B 0.06fF
C47197 PAND2X1_23/Y POR2X1_458/O 0.00fF
C47198 POR2X1_441/Y POR2X1_91/Y 0.01fF
C47199 PAND2X1_635/O POR2X1_582/Y 0.06fF
C47200 PAND2X1_838/B POR2X1_73/Y 0.11fF
C47201 POR2X1_311/Y VDD 0.80fF
C47202 POR2X1_376/B PAND2X1_168/Y 0.01fF
C47203 POR2X1_48/A PAND2X1_784/O 0.06fF
C47204 PAND2X1_677/O PAND2X1_90/Y 0.07fF
C47205 PAND2X1_90/Y POR2X1_330/Y 0.10fF
C47206 PAND2X1_467/B VDD 0.01fF
C47207 PAND2X1_654/CTRL2 POR2X1_409/B 0.01fF
C47208 PAND2X1_293/CTRL PAND2X1_58/A 0.01fF
C47209 PAND2X1_6/Y POR2X1_629/CTRL2 0.01fF
C47210 POR2X1_428/Y POR2X1_426/m4_208_n4# 0.09fF
C47211 POR2X1_609/Y PAND2X1_243/B 0.02fF
C47212 PAND2X1_443/CTRL POR2X1_90/Y 0.01fF
C47213 PAND2X1_326/B POR2X1_166/Y 0.01fF
C47214 PAND2X1_723/Y POR2X1_40/Y 0.03fF
C47215 POR2X1_502/A POR2X1_121/B 0.10fF
C47216 PAND2X1_58/A POR2X1_404/B 0.01fF
C47217 POR2X1_712/A POR2X1_260/B 0.03fF
C47218 PAND2X1_392/O POR2X1_55/Y 0.25fF
C47219 PAND2X1_23/Y POR2X1_220/B 0.03fF
C47220 POR2X1_334/B POR2X1_66/A 0.69fF
C47221 POR2X1_647/Y POR2X1_362/B 0.01fF
C47222 POR2X1_341/A PAND2X1_60/B 0.14fF
C47223 POR2X1_41/B POR2X1_603/Y 0.03fF
C47224 POR2X1_655/Y VDD 0.00fF
C47225 PAND2X1_236/O POR2X1_94/A 0.03fF
C47226 PAND2X1_82/CTRL PAND2X1_39/B 0.08fF
C47227 POR2X1_356/A POR2X1_78/A 0.07fF
C47228 POR2X1_632/CTRL2 POR2X1_532/A 0.01fF
C47229 POR2X1_309/O POR2X1_293/Y 0.02fF
C47230 POR2X1_376/B POR2X1_743/O 0.17fF
C47231 POR2X1_68/A POR2X1_294/Y 0.00fF
C47232 POR2X1_13/A POR2X1_272/CTRL2 0.01fF
C47233 POR2X1_98/A POR2X1_294/A 0.02fF
C47234 POR2X1_66/B POR2X1_121/Y 6.63fF
C47235 POR2X1_666/Y PAND2X1_719/CTRL 0.01fF
C47236 PAND2X1_42/CTRL POR2X1_547/B 0.02fF
C47237 POR2X1_48/A POR2X1_255/Y 0.02fF
C47238 PAND2X1_562/Y PAND2X1_570/B 0.01fF
C47239 POR2X1_416/Y D_INPUT_0 0.03fF
C47240 POR2X1_807/A POR2X1_480/A 0.04fF
C47241 POR2X1_477/A POR2X1_590/A 0.03fF
C47242 POR2X1_48/A PAND2X1_731/CTRL 0.01fF
C47243 POR2X1_54/Y PAND2X1_521/a_76_28# 0.05fF
C47244 POR2X1_257/A POR2X1_283/A 0.14fF
C47245 PAND2X1_299/O VDD 0.00fF
C47246 POR2X1_590/A POR2X1_565/CTRL2 0.01fF
C47247 POR2X1_441/Y PAND2X1_545/Y 0.02fF
C47248 POR2X1_242/CTRL2 POR2X1_578/Y 0.09fF
C47249 POR2X1_180/B POR2X1_663/B 0.03fF
C47250 POR2X1_16/A POR2X1_88/A 0.02fF
C47251 PAND2X1_42/O VDD 0.00fF
C47252 POR2X1_405/CTRL POR2X1_405/Y 0.00fF
C47253 POR2X1_569/CTRL2 POR2X1_355/B 0.04fF
C47254 POR2X1_188/A POR2X1_121/Y 0.01fF
C47255 PAND2X1_452/A POR2X1_257/A 0.01fF
C47256 POR2X1_32/A PAND2X1_718/O 0.07fF
C47257 POR2X1_29/Y D_INPUT_0 0.02fF
C47258 POR2X1_567/B POR2X1_341/Y 0.05fF
C47259 POR2X1_118/O POR2X1_37/Y 0.01fF
C47260 POR2X1_649/B POR2X1_476/A 0.50fF
C47261 PAND2X1_422/CTRL POR2X1_260/B 0.00fF
C47262 POR2X1_52/A PAND2X1_168/Y 0.12fF
C47263 PAND2X1_671/CTRL2 POR2X1_54/Y 0.01fF
C47264 POR2X1_41/B POR2X1_504/Y 0.00fF
C47265 POR2X1_705/B POR2X1_559/A 0.05fF
C47266 POR2X1_78/CTRL POR2X1_78/A 0.01fF
C47267 PAND2X1_714/a_16_344# PAND2X1_731/B 0.01fF
C47268 POR2X1_389/A PAND2X1_666/O 0.06fF
C47269 PAND2X1_808/Y PAND2X1_557/A 0.02fF
C47270 PAND2X1_830/Y PAND2X1_562/B 0.02fF
C47271 PAND2X1_249/m4_208_n4# PAND2X1_193/m4_208_n4# 0.05fF
C47272 PAND2X1_23/Y PAND2X1_23/CTRL2 0.00fF
C47273 PAND2X1_168/Y POR2X1_152/A 0.03fF
C47274 POR2X1_206/A VDD 0.24fF
C47275 POR2X1_416/B PAND2X1_193/Y 0.04fF
C47276 PAND2X1_562/B POR2X1_7/B 0.07fF
C47277 POR2X1_341/A POR2X1_332/O 0.01fF
C47278 D_INPUT_2 POR2X1_40/Y 0.03fF
C47279 POR2X1_254/Y PAND2X1_48/CTRL2 0.07fF
C47280 POR2X1_43/B PAND2X1_444/Y 0.01fF
C47281 PAND2X1_3/a_56_28# D_INPUT_5 0.00fF
C47282 PAND2X1_616/CTRL2 PAND2X1_6/A 0.01fF
C47283 PAND2X1_229/O POR2X1_579/Y 0.00fF
C47284 POR2X1_66/B PAND2X1_612/CTRL 0.01fF
C47285 PAND2X1_93/B POR2X1_569/A 0.07fF
C47286 POR2X1_56/B POR2X1_376/B 0.09fF
C47287 PAND2X1_853/CTRL POR2X1_40/Y 0.01fF
C47288 PAND2X1_6/Y POR2X1_783/CTRL2 0.00fF
C47289 POR2X1_566/A PAND2X1_627/O 0.30fF
C47290 POR2X1_777/B PAND2X1_372/m4_208_n4# 0.05fF
C47291 POR2X1_304/CTRL2 POR2X1_329/A 0.03fF
C47292 PAND2X1_118/CTRL PAND2X1_41/B 0.01fF
C47293 POR2X1_272/O POR2X1_184/Y 0.00fF
C47294 PAND2X1_390/Y POR2X1_184/Y 0.02fF
C47295 PAND2X1_467/B POR2X1_694/a_16_28# 0.02fF
C47296 POR2X1_463/Y POR2X1_862/A 0.02fF
C47297 POR2X1_296/B POR2X1_307/A 0.03fF
C47298 PAND2X1_36/m4_208_n4# PAND2X1_32/B 0.01fF
C47299 POR2X1_66/B POR2X1_139/A 0.01fF
C47300 POR2X1_423/Y PAND2X1_6/A 0.07fF
C47301 POR2X1_407/A POR2X1_783/m4_208_n4# 0.12fF
C47302 POR2X1_30/CTRL2 INPUT_7 0.00fF
C47303 POR2X1_83/CTRL2 D_INPUT_0 0.03fF
C47304 PAND2X1_651/Y PAND2X1_390/Y 0.05fF
C47305 POR2X1_809/A POR2X1_452/Y 0.02fF
C47306 POR2X1_741/Y POR2X1_733/CTRL2 0.00fF
C47307 PAND2X1_469/B PAND2X1_787/O 0.06fF
C47308 POR2X1_177/Y PAND2X1_552/B 0.04fF
C47309 PAND2X1_592/Y PAND2X1_580/B 0.03fF
C47310 POR2X1_61/Y POR2X1_35/Y 1.01fF
C47311 POR2X1_89/CTRL2 POR2X1_394/A 0.05fF
C47312 POR2X1_377/O POR2X1_5/Y 0.01fF
C47313 PAND2X1_531/a_16_344# PAND2X1_111/B 0.03fF
C47314 PAND2X1_97/CTRL2 POR2X1_394/A 0.04fF
C47315 POR2X1_83/B PAND2X1_154/CTRL2 0.00fF
C47316 PAND2X1_830/Y POR2X1_13/A 0.03fF
C47317 PAND2X1_250/CTRL PAND2X1_32/B 0.01fF
C47318 POR2X1_719/O POR2X1_121/B 0.02fF
C47319 POR2X1_447/A POR2X1_186/B 0.03fF
C47320 PAND2X1_65/B POR2X1_341/O 0.17fF
C47321 POR2X1_13/A POR2X1_7/B 10.35fF
C47322 POR2X1_186/Y POR2X1_731/O 0.25fF
C47323 POR2X1_327/Y POR2X1_260/B 0.01fF
C47324 PAND2X1_299/O PAND2X1_32/B 0.03fF
C47325 POR2X1_750/B PAND2X1_88/Y 0.05fF
C47326 POR2X1_78/A POR2X1_569/A 0.18fF
C47327 PAND2X1_217/B POR2X1_38/Y 0.02fF
C47328 POR2X1_32/A PAND2X1_123/O 0.04fF
C47329 POR2X1_194/A POR2X1_194/CTRL 0.03fF
C47330 PAND2X1_244/O PAND2X1_175/B 0.05fF
C47331 POR2X1_407/A POR2X1_480/A 0.07fF
C47332 PAND2X1_751/m4_208_n4# POR2X1_546/A 0.03fF
C47333 POR2X1_52/A PAND2X1_776/CTRL2 0.01fF
C47334 PAND2X1_253/CTRL POR2X1_241/B 0.01fF
C47335 PAND2X1_94/A POR2X1_296/B 0.24fF
C47336 POR2X1_102/Y PAND2X1_723/A 0.11fF
C47337 PAND2X1_260/a_16_344# PAND2X1_555/Y 0.01fF
C47338 POR2X1_514/CTRL VDD 0.00fF
C47339 POR2X1_220/Y POR2X1_832/B 0.03fF
C47340 POR2X1_52/A POR2X1_56/B 0.03fF
C47341 POR2X1_97/CTRL POR2X1_78/A 0.01fF
C47342 POR2X1_505/CTRL POR2X1_669/B 0.02fF
C47343 POR2X1_500/A PAND2X1_60/B 0.03fF
C47344 POR2X1_455/A VDD -0.00fF
C47345 PAND2X1_775/O POR2X1_7/B 0.17fF
C47346 PAND2X1_473/B POR2X1_816/A 0.03fF
C47347 POR2X1_119/Y PAND2X1_469/CTRL 0.01fF
C47348 POR2X1_466/A POR2X1_544/B 0.01fF
C47349 PAND2X1_73/Y POR2X1_463/Y 0.07fF
C47350 PAND2X1_218/A VDD 0.00fF
C47351 PAND2X1_41/B POR2X1_216/O 0.15fF
C47352 POR2X1_502/A POR2X1_795/B 0.03fF
C47353 PAND2X1_56/Y POR2X1_502/A 0.04fF
C47354 PAND2X1_467/B PAND2X1_467/O 0.08fF
C47355 PAND2X1_183/CTRL POR2X1_732/B 0.30fF
C47356 POR2X1_131/Y POR2X1_102/Y 0.71fF
C47357 POR2X1_477/B POR2X1_854/B 0.10fF
C47358 PAND2X1_435/CTRL POR2X1_433/Y 0.01fF
C47359 POR2X1_83/B PAND2X1_714/Y 0.67fF
C47360 POR2X1_303/O POR2X1_76/A 0.07fF
C47361 PAND2X1_468/CTRL2 PAND2X1_798/B 0.01fF
C47362 POR2X1_65/A PAND2X1_551/CTRL2 0.03fF
C47363 POR2X1_10/CTRL POR2X1_83/B 0.01fF
C47364 POR2X1_805/Y POR2X1_758/Y 0.01fF
C47365 POR2X1_20/B D_INPUT_4 0.03fF
C47366 POR2X1_663/B POR2X1_169/A 0.02fF
C47367 POR2X1_57/A PAND2X1_756/CTRL 0.01fF
C47368 POR2X1_49/Y POR2X1_283/A 0.01fF
C47369 PAND2X1_41/B PAND2X1_63/B 0.03fF
C47370 PAND2X1_228/CTRL2 PAND2X1_197/Y 0.00fF
C47371 POR2X1_838/B POR2X1_507/A 0.03fF
C47372 PAND2X1_575/A POR2X1_494/Y 1.34fF
C47373 POR2X1_144/CTRL POR2X1_669/B 0.03fF
C47374 POR2X1_3/A POR2X1_2/O 0.01fF
C47375 POR2X1_106/Y PAND2X1_348/Y 0.11fF
C47376 POR2X1_467/O PAND2X1_52/B 0.01fF
C47377 POR2X1_38/Y VDD 2.80fF
C47378 PAND2X1_478/a_56_28# POR2X1_46/Y 0.00fF
C47379 POR2X1_78/B PAND2X1_697/m4_208_n4# 0.15fF
C47380 PAND2X1_96/B POR2X1_404/B 0.01fF
C47381 POR2X1_669/B PAND2X1_708/O 0.04fF
C47382 POR2X1_351/Y POR2X1_776/B 0.03fF
C47383 PAND2X1_766/CTRL POR2X1_260/A 0.01fF
C47384 POR2X1_129/a_16_28# POR2X1_129/Y 0.06fF
C47385 POR2X1_66/B PAND2X1_413/CTRL2 -0.00fF
C47386 POR2X1_750/B PAND2X1_376/O 0.02fF
C47387 POR2X1_52/A PAND2X1_814/CTRL2 0.01fF
C47388 POR2X1_302/CTRL2 POR2X1_383/A 0.06fF
C47389 POR2X1_853/A POR2X1_775/A 0.06fF
C47390 POR2X1_860/A POR2X1_276/Y 0.03fF
C47391 POR2X1_407/A PAND2X1_90/A 0.06fF
C47392 POR2X1_481/A POR2X1_142/Y 0.03fF
C47393 POR2X1_197/Y VDD 0.25fF
C47394 PAND2X1_795/m4_208_n4# PAND2X1_575/m4_208_n4# 0.13fF
C47395 POR2X1_193/A POR2X1_702/A 0.03fF
C47396 POR2X1_625/Y POR2X1_93/A 0.08fF
C47397 POR2X1_579/Y POR2X1_702/A 4.80fF
C47398 PAND2X1_643/Y POR2X1_7/B 0.04fF
C47399 POR2X1_212/CTRL VDD 0.00fF
C47400 POR2X1_862/O POR2X1_647/B 0.01fF
C47401 POR2X1_700/CTRL2 PAND2X1_711/A 0.01fF
C47402 POR2X1_68/A PAND2X1_29/CTRL2 0.00fF
C47403 PAND2X1_568/B PAND2X1_568/O 0.01fF
C47404 POR2X1_452/Y POR2X1_728/A 0.02fF
C47405 PAND2X1_661/B POR2X1_277/O 0.01fF
C47406 PAND2X1_137/Y PAND2X1_803/Y 0.07fF
C47407 POR2X1_52/A POR2X1_92/CTRL 0.00fF
C47408 POR2X1_43/B PAND2X1_357/Y 0.03fF
C47409 PAND2X1_217/B POR2X1_153/Y 0.05fF
C47410 POR2X1_614/A POR2X1_800/A 0.03fF
C47411 POR2X1_5/Y POR2X1_6/CTRL2 0.01fF
C47412 POR2X1_289/Y POR2X1_77/Y 0.02fF
C47413 POR2X1_52/A POR2X1_526/a_16_28# 0.02fF
C47414 POR2X1_40/Y PAND2X1_123/Y 0.03fF
C47415 PAND2X1_736/A PAND2X1_186/CTRL 0.06fF
C47416 POR2X1_356/A PAND2X1_173/CTRL 0.18fF
C47417 POR2X1_121/B POR2X1_188/Y 0.03fF
C47418 POR2X1_163/CTRL2 POR2X1_394/A 0.01fF
C47419 PAND2X1_57/B PAND2X1_765/CTRL2 0.00fF
C47420 POR2X1_219/a_16_28# POR2X1_294/B 0.00fF
C47421 POR2X1_502/A POR2X1_383/A 0.27fF
C47422 PAND2X1_726/B PAND2X1_712/B 0.02fF
C47423 POR2X1_16/A POR2X1_290/a_16_28# 0.08fF
C47424 POR2X1_114/B POR2X1_513/Y 0.03fF
C47425 PAND2X1_94/A POR2X1_547/B 0.01fF
C47426 PAND2X1_20/A POR2X1_560/CTRL2 0.01fF
C47427 POR2X1_296/B PAND2X1_136/CTRL2 0.01fF
C47428 POR2X1_334/B POR2X1_532/A 0.14fF
C47429 POR2X1_514/CTRL PAND2X1_32/B 0.01fF
C47430 POR2X1_462/B POR2X1_793/A 0.01fF
C47431 POR2X1_720/B PAND2X1_69/A 0.03fF
C47432 PAND2X1_484/CTRL POR2X1_287/B 0.12fF
C47433 POR2X1_389/A PAND2X1_385/O 0.02fF
C47434 POR2X1_416/B POR2X1_699/O 0.01fF
C47435 POR2X1_283/A PAND2X1_553/B 0.07fF
C47436 INPUT_1 VDD 2.89fF
C47437 PAND2X1_392/B POR2X1_384/A 0.01fF
C47438 POR2X1_416/B POR2X1_416/A 0.01fF
C47439 POR2X1_614/A POR2X1_702/A 0.01fF
C47440 PAND2X1_462/O POR2X1_48/A 0.01fF
C47441 PAND2X1_802/B VDD 0.11fF
C47442 POR2X1_383/A PAND2X1_530/CTRL2 0.01fF
C47443 D_INPUT_3 POR2X1_119/a_16_28# 0.03fF
C47444 POR2X1_68/B PAND2X1_110/a_76_28# 0.02fF
C47445 POR2X1_572/CTRL POR2X1_260/A 0.00fF
C47446 POR2X1_62/Y PAND2X1_61/Y 0.07fF
C47447 POR2X1_43/B POR2X1_278/A 0.03fF
C47448 POR2X1_119/Y POR2X1_423/Y 0.03fF
C47449 PAND2X1_93/B PAND2X1_72/A 0.06fF
C47450 PAND2X1_593/Y PAND2X1_364/B 0.07fF
C47451 POR2X1_46/Y PAND2X1_514/O 0.05fF
C47452 PAND2X1_738/Y PAND2X1_348/A 0.10fF
C47453 VDD POR2X1_153/Y 5.65fF
C47454 PAND2X1_724/O POR2X1_73/Y 0.02fF
C47455 POR2X1_631/A POR2X1_631/B 0.71fF
C47456 PAND2X1_90/Y POR2X1_703/O 0.05fF
C47457 POR2X1_835/a_16_28# POR2X1_835/A 0.08fF
C47458 POR2X1_719/CTRL2 PAND2X1_32/B 0.03fF
C47459 POR2X1_528/Y POR2X1_43/B 0.03fF
C47460 PAND2X1_55/Y POR2X1_407/O 0.03fF
C47461 PAND2X1_798/B PAND2X1_574/CTRL2 0.01fF
C47462 PAND2X1_659/Y PAND2X1_736/O 0.02fF
C47463 PAND2X1_90/Y POR2X1_337/Y 0.02fF
C47464 PAND2X1_41/B PAND2X1_166/CTRL2 0.02fF
C47465 PAND2X1_23/Y POR2X1_787/O 0.01fF
C47466 POR2X1_16/A PAND2X1_341/CTRL 0.00fF
C47467 POR2X1_190/Y PAND2X1_189/CTRL2 0.00fF
C47468 POR2X1_38/B PAND2X1_670/CTRL 0.01fF
C47469 PAND2X1_343/CTRL POR2X1_42/Y 0.01fF
C47470 PAND2X1_495/CTRL PAND2X1_60/B 0.00fF
C47471 POR2X1_447/CTRL2 POR2X1_510/Y 0.01fF
C47472 PAND2X1_580/B POR2X1_767/CTRL2 0.00fF
C47473 POR2X1_750/B POR2X1_568/B 0.05fF
C47474 PAND2X1_341/B PAND2X1_206/CTRL 0.01fF
C47475 POR2X1_333/Y POR2X1_578/Y 0.03fF
C47476 POR2X1_57/A POR2X1_396/Y 0.01fF
C47477 PAND2X1_297/CTRL POR2X1_402/A 0.01fF
C47478 POR2X1_379/O PAND2X1_752/Y 0.03fF
C47479 POR2X1_329/A POR2X1_271/B 0.03fF
C47480 POR2X1_294/B POR2X1_507/A 0.01fF
C47481 POR2X1_78/A PAND2X1_72/A 0.46fF
C47482 POR2X1_778/B POR2X1_101/Y 0.03fF
C47483 POR2X1_502/A POR2X1_560/Y 0.59fF
C47484 PAND2X1_824/B POR2X1_208/m4_208_n4# 0.09fF
C47485 POR2X1_702/a_16_28# POR2X1_702/A 0.10fF
C47486 PAND2X1_726/B PAND2X1_546/CTRL2 0.02fF
C47487 PAND2X1_736/Y PAND2X1_853/B 0.07fF
C47488 PAND2X1_388/Y POR2X1_387/Y 0.07fF
C47489 PAND2X1_6/Y POR2X1_456/B 0.03fF
C47490 POR2X1_327/Y PAND2X1_55/Y 0.02fF
C47491 PAND2X1_390/Y PAND2X1_858/B 0.01fF
C47492 POR2X1_783/CTRL2 PAND2X1_52/B 0.03fF
C47493 POR2X1_813/Y POR2X1_38/Y 0.03fF
C47494 POR2X1_134/Y PAND2X1_346/Y 0.01fF
C47495 POR2X1_447/B POR2X1_566/A 0.10fF
C47496 POR2X1_833/CTRL POR2X1_186/B 0.01fF
C47497 POR2X1_831/O POR2X1_814/A 0.17fF
C47498 PAND2X1_29/O POR2X1_260/A 0.01fF
C47499 PAND2X1_513/CTRL2 POR2X1_77/Y 0.03fF
C47500 PAND2X1_865/Y PAND2X1_795/B 0.12fF
C47501 POR2X1_559/a_56_344# POR2X1_673/Y 0.00fF
C47502 PAND2X1_549/B POR2X1_387/Y 0.07fF
C47503 POR2X1_833/A POR2X1_786/Y 1.15fF
C47504 VDD PAND2X1_136/CTRL 0.00fF
C47505 INPUT_1 PAND2X1_32/B 0.03fF
C47506 POR2X1_62/Y PAND2X1_228/CTRL2 0.01fF
C47507 POR2X1_825/Y POR2X1_669/B 0.03fF
C47508 POR2X1_416/B POR2X1_763/A 0.07fF
C47509 POR2X1_163/CTRL POR2X1_158/Y 0.00fF
C47510 POR2X1_65/A POR2X1_86/Y 0.01fF
C47511 POR2X1_96/O POR2X1_38/B 0.10fF
C47512 POR2X1_343/Y POR2X1_362/B 0.07fF
C47513 POR2X1_242/O POR2X1_568/A 0.06fF
C47514 POR2X1_273/Y POR2X1_300/Y 0.02fF
C47515 POR2X1_3/A POR2X1_260/A 1.16fF
C47516 POR2X1_220/Y POR2X1_330/O 0.00fF
C47517 POR2X1_16/A D_INPUT_3 0.01fF
C47518 PAND2X1_860/A POR2X1_102/Y 0.04fF
C47519 PAND2X1_551/a_16_344# PAND2X1_545/Y 0.03fF
C47520 PAND2X1_56/Y POR2X1_188/Y 0.03fF
C47521 PAND2X1_39/B POR2X1_556/A 0.02fF
C47522 POR2X1_38/B PAND2X1_531/CTRL 0.04fF
C47523 PAND2X1_216/B PAND2X1_175/B 0.01fF
C47524 POR2X1_351/Y POR2X1_192/B 0.15fF
C47525 POR2X1_46/Y POR2X1_39/B 0.05fF
C47526 POR2X1_391/Y PAND2X1_134/CTRL2 0.02fF
C47527 POR2X1_136/Y PAND2X1_348/A 0.02fF
C47528 POR2X1_96/A POR2X1_305/O 0.01fF
C47529 PAND2X1_285/O POR2X1_282/Y 0.04fF
C47530 PAND2X1_607/CTRL2 PAND2X1_58/A 0.01fF
C47531 POR2X1_722/Y PAND2X1_56/A 0.02fF
C47532 PAND2X1_492/O PAND2X1_72/A 0.05fF
C47533 PAND2X1_358/A PAND2X1_338/B 0.07fF
C47534 POR2X1_751/Y POR2X1_7/A 0.03fF
C47535 INPUT_1 PAND2X1_637/CTRL2 0.01fF
C47536 PAND2X1_476/A POR2X1_406/A 0.00fF
C47537 PAND2X1_90/CTRL2 POR2X1_38/B 0.00fF
C47538 PAND2X1_187/CTRL2 POR2X1_191/B 0.00fF
C47539 POR2X1_101/CTRL2 POR2X1_334/Y 0.01fF
C47540 PAND2X1_623/Y POR2X1_39/B 0.03fF
C47541 POR2X1_54/Y POR2X1_126/CTRL2 0.01fF
C47542 POR2X1_353/A POR2X1_151/CTRL 0.01fF
C47543 POR2X1_394/A POR2X1_527/Y 0.65fF
C47544 INPUT_1 POR2X1_673/Y 0.03fF
C47545 POR2X1_349/O POR2X1_532/A 0.01fF
C47546 POR2X1_327/Y POR2X1_337/A 0.46fF
C47547 POR2X1_732/B POR2X1_181/a_16_28# 0.05fF
C47548 PAND2X1_334/O POR2X1_39/B 0.17fF
C47549 PAND2X1_840/A POR2X1_39/B 0.01fF
C47550 POR2X1_420/Y POR2X1_329/A 0.02fF
C47551 POR2X1_68/A POR2X1_39/B 0.03fF
C47552 POR2X1_566/A POR2X1_181/A 0.05fF
C47553 PAND2X1_641/Y POR2X1_83/a_76_344# 0.01fF
C47554 POR2X1_513/Y POR2X1_513/A 0.38fF
C47555 POR2X1_433/Y POR2X1_77/Y 0.03fF
C47556 POR2X1_383/A POR2X1_188/Y 0.10fF
C47557 PAND2X1_631/A POR2X1_136/Y 0.04fF
C47558 POR2X1_796/Y POR2X1_808/CTRL 0.01fF
C47559 PAND2X1_63/B PAND2X1_143/CTRL 0.01fF
C47560 POR2X1_713/a_16_28# POR2X1_711/Y 0.02fF
C47561 PAND2X1_341/Y PAND2X1_358/A 0.10fF
C47562 POR2X1_36/CTRL2 POR2X1_39/B 0.00fF
C47563 POR2X1_7/CTRL2 POR2X1_7/Y 0.01fF
C47564 PAND2X1_476/A PAND2X1_63/B 0.02fF
C47565 POR2X1_75/O POR2X1_416/B 0.01fF
C47566 PAND2X1_863/A PAND2X1_854/A 0.03fF
C47567 POR2X1_187/O POR2X1_385/Y 0.04fF
C47568 POR2X1_260/B POR2X1_644/Y 0.01fF
C47569 POR2X1_54/Y PAND2X1_669/O 0.03fF
C47570 POR2X1_510/A PAND2X1_72/A 0.07fF
C47571 POR2X1_751/Y POR2X1_384/Y 0.00fF
C47572 POR2X1_191/Y POR2X1_545/CTRL2 0.03fF
C47573 PAND2X1_20/A POR2X1_556/A 0.05fF
C47574 PAND2X1_485/O POR2X1_260/B 0.05fF
C47575 POR2X1_661/A POR2X1_722/Y 0.03fF
C47576 PAND2X1_477/A POR2X1_119/Y 0.01fF
C47577 PAND2X1_407/CTRL2 POR2X1_29/A 0.01fF
C47578 POR2X1_555/A POR2X1_630/B 0.01fF
C47579 PAND2X1_165/m4_208_n4# POR2X1_854/B 0.04fF
C47580 PAND2X1_797/Y PAND2X1_569/B 0.07fF
C47581 POR2X1_27/O POR2X1_5/Y 0.00fF
C47582 PAND2X1_827/CTRL2 POR2X1_294/Y 0.00fF
C47583 PAND2X1_678/CTRL POR2X1_72/B 0.00fF
C47584 POR2X1_345/CTRL POR2X1_99/B 0.00fF
C47585 POR2X1_567/A POR2X1_507/A 0.10fF
C47586 POR2X1_122/CTRL PAND2X1_659/Y 0.00fF
C47587 POR2X1_254/A POR2X1_341/A 0.00fF
C47588 POR2X1_848/A POR2X1_754/Y 1.77fF
C47589 POR2X1_65/A PAND2X1_449/a_16_344# 0.01fF
C47590 PAND2X1_399/a_16_344# POR2X1_294/A 0.02fF
C47591 PAND2X1_717/A PAND2X1_556/B 0.11fF
C47592 PAND2X1_173/CTRL PAND2X1_72/A 0.01fF
C47593 POR2X1_341/A POR2X1_750/B 0.10fF
C47594 POR2X1_357/a_56_344# POR2X1_192/B 0.00fF
C47595 POR2X1_814/B POR2X1_556/A 0.06fF
C47596 PAND2X1_630/B POR2X1_42/Y 0.03fF
C47597 POR2X1_486/B POR2X1_260/A 0.11fF
C47598 PAND2X1_404/Y POR2X1_60/A 0.03fF
C47599 PAND2X1_629/O POR2X1_20/B 0.09fF
C47600 POR2X1_502/A POR2X1_648/Y 0.07fF
C47601 POR2X1_630/O POR2X1_590/A 0.18fF
C47602 POR2X1_456/B POR2X1_632/Y 0.03fF
C47603 POR2X1_475/A POR2X1_475/CTRL 0.01fF
C47604 POR2X1_327/Y POR2X1_741/O 0.26fF
C47605 POR2X1_711/Y POR2X1_308/B 0.03fF
C47606 POR2X1_210/A POR2X1_330/CTRL 0.01fF
C47607 PAND2X1_403/Y POR2X1_411/B 0.01fF
C47608 POR2X1_149/CTRL PAND2X1_90/Y 0.01fF
C47609 POR2X1_122/Y POR2X1_20/B 0.01fF
C47610 PAND2X1_666/CTRL2 PAND2X1_20/A 0.00fF
C47611 POR2X1_556/A POR2X1_325/A 0.03fF
C47612 POR2X1_129/a_16_28# POR2X1_37/Y 0.05fF
C47613 POR2X1_294/Y PAND2X1_58/A 0.00fF
C47614 POR2X1_161/a_16_28# POR2X1_162/Y 0.02fF
C47615 POR2X1_445/A POR2X1_456/O 0.01fF
C47616 POR2X1_43/O PAND2X1_560/B 0.01fF
C47617 POR2X1_760/A PAND2X1_216/O 0.05fF
C47618 POR2X1_66/B POR2X1_286/O 0.18fF
C47619 POR2X1_333/A POR2X1_97/A 2.81fF
C47620 POR2X1_240/B POR2X1_590/A 0.01fF
C47621 PAND2X1_274/CTRL POR2X1_411/B 0.01fF
C47622 POR2X1_65/CTRL POR2X1_55/Y 0.15fF
C47623 PAND2X1_23/Y PAND2X1_45/CTRL 0.01fF
C47624 PAND2X1_39/B POR2X1_400/A 0.04fF
C47625 PAND2X1_717/A POR2X1_599/A 2.07fF
C47626 POR2X1_856/B POR2X1_856/CTRL2 0.12fF
C47627 PAND2X1_52/CTRL2 POR2X1_35/Y 0.01fF
C47628 PAND2X1_677/a_16_344# POR2X1_66/A 0.01fF
C47629 POR2X1_567/B PAND2X1_41/B 0.06fF
C47630 PAND2X1_313/a_16_344# PAND2X1_72/A 0.02fF
C47631 POR2X1_188/A PAND2X1_282/CTRL2 0.01fF
C47632 PAND2X1_10/CTRL2 PAND2X1_41/B 0.01fF
C47633 POR2X1_20/O POR2X1_20/B 0.02fF
C47634 POR2X1_20/A PAND2X1_8/Y 0.10fF
C47635 POR2X1_189/Y POR2X1_679/CTRL2 0.01fF
C47636 PAND2X1_231/CTRL2 POR2X1_32/A 0.01fF
C47637 PAND2X1_93/B POR2X1_632/A 0.00fF
C47638 POR2X1_760/A PAND2X1_218/a_16_344# 0.02fF
C47639 POR2X1_768/a_16_28# POR2X1_768/A -0.00fF
C47640 POR2X1_66/A PAND2X1_387/O 0.03fF
C47641 POR2X1_715/A POR2X1_715/O 0.05fF
C47642 POR2X1_846/CTRL2 POR2X1_260/A 0.04fF
C47643 POR2X1_23/Y POR2X1_238/O 0.02fF
C47644 POR2X1_54/Y POR2X1_790/O 0.01fF
C47645 PAND2X1_654/CTRL PAND2X1_9/Y 0.01fF
C47646 POR2X1_23/Y PAND2X1_735/CTRL2 0.01fF
C47647 POR2X1_248/A VDD 0.00fF
C47648 POR2X1_13/A POR2X1_265/CTRL2 0.01fF
C47649 PAND2X1_47/B PAND2X1_44/O 0.00fF
C47650 POR2X1_186/Y PAND2X1_331/O 0.02fF
C47651 POR2X1_441/Y PAND2X1_551/A 0.01fF
C47652 PAND2X1_213/B PAND2X1_213/O 0.00fF
C47653 POR2X1_230/CTRL2 POR2X1_32/A 0.01fF
C47654 PAND2X1_688/O POR2X1_48/A 0.17fF
C47655 POR2X1_257/A POR2X1_55/Y 0.29fF
C47656 POR2X1_52/A POR2X1_815/A 0.01fF
C47657 POR2X1_448/Y POR2X1_296/B 0.04fF
C47658 POR2X1_862/B POR2X1_121/B 0.03fF
C47659 POR2X1_682/a_56_344# POR2X1_669/B 0.00fF
C47660 POR2X1_49/Y POR2X1_14/Y 0.32fF
C47661 POR2X1_265/O PAND2X1_35/Y 0.01fF
C47662 PAND2X1_822/O POR2X1_835/A 0.01fF
C47663 POR2X1_49/Y PAND2X1_453/A 0.11fF
C47664 PAND2X1_267/CTRL2 PAND2X1_215/B 0.02fF
C47665 PAND2X1_42/O POR2X1_267/A 0.15fF
C47666 POR2X1_67/Y POR2X1_408/Y 0.03fF
C47667 POR2X1_35/B POR2X1_34/Y 0.01fF
C47668 PAND2X1_557/A PAND2X1_221/m4_208_n4# 0.07fF
C47669 PAND2X1_219/A PAND2X1_219/B 0.01fF
C47670 PAND2X1_205/A PAND2X1_205/B 0.20fF
C47671 PAND2X1_790/a_76_28# POR2X1_7/B 0.01fF
C47672 POR2X1_48/A POR2X1_46/Y 3.06fF
C47673 PAND2X1_218/CTRL2 PAND2X1_267/Y 0.01fF
C47674 POR2X1_67/Y POR2X1_391/a_76_344# 0.00fF
C47675 POR2X1_130/A POR2X1_267/CTRL2 0.02fF
C47676 PAND2X1_48/B PAND2X1_251/O 0.06fF
C47677 PAND2X1_96/B POR2X1_663/B 10.51fF
C47678 POR2X1_159/O POR2X1_376/B 0.01fF
C47679 POR2X1_454/B VDD 0.00fF
C47680 PAND2X1_24/CTRL D_INPUT_1 0.01fF
C47681 PAND2X1_9/Y POR2X1_38/Y 0.03fF
C47682 POR2X1_411/B POR2X1_93/A 0.44fF
C47683 POR2X1_16/A POR2X1_600/CTRL2 0.01fF
C47684 POR2X1_78/A POR2X1_244/B 0.03fF
C47685 POR2X1_411/B POR2X1_91/Y 0.03fF
C47686 POR2X1_590/A POR2X1_214/O 0.18fF
C47687 PAND2X1_786/CTRL PAND2X1_84/Y 0.02fF
C47688 POR2X1_66/A PAND2X1_176/a_16_344# 0.02fF
C47689 PAND2X1_40/CTRL2 PAND2X1_59/B 0.01fF
C47690 POR2X1_44/CTRL2 INPUT_7 0.00fF
C47691 PAND2X1_220/Y PAND2X1_562/B 0.07fF
C47692 PAND2X1_826/O PAND2X1_96/B 0.01fF
C47693 POR2X1_643/CTRL2 POR2X1_294/A 0.03fF
C47694 D_INPUT_0 POR2X1_500/a_16_28# 0.02fF
C47695 PAND2X1_22/CTRL PAND2X1_32/B 0.11fF
C47696 POR2X1_654/B PAND2X1_65/B 0.01fF
C47697 POR2X1_29/A POR2X1_7/B 0.06fF
C47698 PAND2X1_391/CTRL POR2X1_42/Y 0.12fF
C47699 POR2X1_850/A POR2X1_660/A 0.01fF
C47700 POR2X1_865/CTRL2 POR2X1_260/B 0.02fF
C47701 PAND2X1_592/Y POR2X1_32/A 10.50fF
C47702 PAND2X1_214/A VDD 0.12fF
C47703 POR2X1_816/Y POR2X1_38/B 0.03fF
C47704 PAND2X1_406/O PAND2X1_32/B 0.03fF
C47705 POR2X1_23/Y POR2X1_56/Y 0.03fF
C47706 PAND2X1_79/O D_INPUT_0 0.02fF
C47707 POR2X1_607/A POR2X1_411/CTRL 0.00fF
C47708 PAND2X1_247/O POR2X1_7/A 0.05fF
C47709 POR2X1_56/a_16_28# PAND2X1_254/Y 0.02fF
C47710 POR2X1_278/Y PAND2X1_557/A 5.94fF
C47711 POR2X1_686/B POR2X1_750/B 0.03fF
C47712 POR2X1_814/B PAND2X1_236/CTRL2 0.03fF
C47713 POR2X1_78/B PAND2X1_41/B 5.12fF
C47714 D_INPUT_0 PAND2X1_339/Y 0.05fF
C47715 POR2X1_502/A POR2X1_634/O 0.30fF
C47716 PAND2X1_39/B PAND2X1_393/O 0.04fF
C47717 POR2X1_78/A POR2X1_562/CTRL 0.08fF
C47718 POR2X1_644/Y POR2X1_407/Y 0.01fF
C47719 PAND2X1_736/A PAND2X1_362/A 0.00fF
C47720 POR2X1_446/B POR2X1_510/Y 0.22fF
C47721 POR2X1_333/A POR2X1_468/a_56_344# 0.00fF
C47722 POR2X1_315/Y POR2X1_442/O 0.05fF
C47723 POR2X1_154/O POR2X1_750/B 0.01fF
C47724 POR2X1_48/A POR2X1_258/CTRL 0.00fF
C47725 POR2X1_333/A POR2X1_366/Y 0.10fF
C47726 D_GATE_222 POR2X1_555/B 0.03fF
C47727 PAND2X1_475/a_76_28# INPUT_0 0.01fF
C47728 POR2X1_264/CTRL2 POR2X1_294/B 0.12fF
C47729 PAND2X1_554/O POR2X1_7/B 0.05fF
C47730 POR2X1_106/O POR2X1_183/Y 0.00fF
C47731 POR2X1_669/B POR2X1_518/Y 0.03fF
C47732 POR2X1_97/A POR2X1_775/O 0.02fF
C47733 POR2X1_13/A PAND2X1_220/Y 0.03fF
C47734 POR2X1_609/a_16_28# POR2X1_609/A 0.03fF
C47735 POR2X1_294/Y PAND2X1_96/B 0.00fF
C47736 POR2X1_709/A PAND2X1_748/CTRL 0.01fF
C47737 PAND2X1_472/A POR2X1_669/B 0.14fF
C47738 INPUT_1 PAND2X1_9/Y 4.88fF
C47739 POR2X1_60/A POR2X1_289/CTRL2 0.01fF
C47740 POR2X1_720/B POR2X1_720/O 0.01fF
C47741 POR2X1_52/A PAND2X1_195/a_76_28# 0.02fF
C47742 POR2X1_567/B POR2X1_714/CTRL 0.28fF
C47743 POR2X1_457/m4_208_n4# POR2X1_220/Y 0.08fF
C47744 POR2X1_27/Y POR2X1_42/Y 0.13fF
C47745 POR2X1_43/B POR2X1_667/A 0.03fF
C47746 POR2X1_558/B POR2X1_361/O 0.00fF
C47747 POR2X1_434/A POR2X1_209/A 0.03fF
C47748 POR2X1_446/B POR2X1_276/Y 0.01fF
C47749 POR2X1_471/A PAND2X1_313/O 0.07fF
C47750 POR2X1_781/CTRL VDD -0.00fF
C47751 POR2X1_57/A POR2X1_609/Y 0.06fF
C47752 POR2X1_48/A PAND2X1_350/O 0.01fF
C47753 POR2X1_222/a_16_28# POR2X1_222/A -0.00fF
C47754 POR2X1_616/O POR2X1_7/A 0.02fF
C47755 POR2X1_294/B POR2X1_734/A 0.10fF
C47756 POR2X1_49/Y POR2X1_55/Y 0.09fF
C47757 POR2X1_383/A POR2X1_493/A 0.04fF
C47758 POR2X1_66/B POR2X1_391/Y 0.07fF
C47759 PAND2X1_280/O PAND2X1_90/Y 0.23fF
C47760 POR2X1_23/Y POR2X1_235/Y 0.12fF
C47761 PAND2X1_9/Y POR2X1_153/Y 0.05fF
C47762 POR2X1_604/Y POR2X1_73/Y 0.10fF
C47763 POR2X1_567/B POR2X1_704/O 0.57fF
C47764 POR2X1_814/B PAND2X1_385/CTRL 0.00fF
C47765 PAND2X1_658/O PAND2X1_658/B 0.05fF
C47766 POR2X1_610/CTRL2 POR2X1_260/A 0.03fF
C47767 POR2X1_130/A PAND2X1_511/O 0.06fF
C47768 POR2X1_20/B PAND2X1_508/Y 0.03fF
C47769 D_INPUT_2 POR2X1_611/CTRL 0.03fF
C47770 PAND2X1_57/B POR2X1_596/Y 0.01fF
C47771 POR2X1_416/B PAND2X1_405/CTRL2 0.01fF
C47772 PAND2X1_23/Y POR2X1_402/O 0.01fF
C47773 POR2X1_502/A INPUT_0 0.14fF
C47774 PAND2X1_423/a_16_344# PAND2X1_55/Y 0.01fF
C47775 PAND2X1_860/A POR2X1_173/O 0.02fF
C47776 D_INPUT_0 PAND2X1_28/CTRL 0.01fF
C47777 POR2X1_301/A POR2X1_260/A 0.02fF
C47778 POR2X1_848/A POR2X1_754/CTRL 0.03fF
C47779 POR2X1_532/A PAND2X1_394/O 0.04fF
C47780 POR2X1_41/B PAND2X1_556/B 0.04fF
C47781 POR2X1_57/A POR2X1_420/Y 0.00fF
C47782 PAND2X1_39/B POR2X1_398/O 0.06fF
C47783 PAND2X1_859/A POR2X1_382/a_16_28# 0.02fF
C47784 POR2X1_121/O POR2X1_590/A 0.01fF
C47785 POR2X1_566/A POR2X1_220/Y 0.03fF
C47786 D_INPUT_2 POR2X1_5/Y 0.17fF
C47787 POR2X1_68/A POR2X1_402/CTRL 0.01fF
C47788 POR2X1_523/Y POR2X1_849/CTRL 0.01fF
C47789 POR2X1_304/Y POR2X1_56/B 0.02fF
C47790 POR2X1_130/A POR2X1_404/Y 0.07fF
C47791 POR2X1_58/Y INPUT_0 0.03fF
C47792 PAND2X1_460/CTRL2 POR2X1_94/A 0.01fF
C47793 PAND2X1_84/a_76_28# POR2X1_81/Y 0.03fF
C47794 POR2X1_134/Y PAND2X1_354/A 0.06fF
C47795 POR2X1_376/B PAND2X1_565/CTRL2 0.00fF
C47796 PAND2X1_433/O POR2X1_480/A 0.01fF
C47797 PAND2X1_42/CTRL2 POR2X1_38/B 0.02fF
C47798 POR2X1_41/B PAND2X1_254/Y 0.05fF
C47799 PAND2X1_425/CTRL2 INPUT_6 0.01fF
C47800 POR2X1_76/Y POR2X1_465/B 0.01fF
C47801 POR2X1_271/Y POR2X1_91/Y 0.14fF
C47802 POR2X1_777/B PAND2X1_536/m4_208_n4# 0.07fF
C47803 PAND2X1_795/B POR2X1_494/Y 0.10fF
C47804 POR2X1_234/A POR2X1_825/Y 0.02fF
C47805 POR2X1_258/O POR2X1_312/Y 0.31fF
C47806 POR2X1_323/CTRL2 POR2X1_73/Y 0.01fF
C47807 PAND2X1_73/Y POR2X1_101/Y 0.05fF
C47808 PAND2X1_469/B PAND2X1_473/B 0.08fF
C47809 PAND2X1_20/A POR2X1_276/A 0.03fF
C47810 POR2X1_45/Y PAND2X1_84/Y 0.03fF
C47811 POR2X1_614/A POR2X1_640/A 0.02fF
C47812 POR2X1_67/A POR2X1_172/O 0.01fF
C47813 POR2X1_65/A POR2X1_73/Y 6.03fF
C47814 POR2X1_630/A POR2X1_510/Y 0.00fF
C47815 POR2X1_602/B PAND2X1_60/B 0.02fF
C47816 PAND2X1_20/A POR2X1_566/B 0.03fF
C47817 POR2X1_814/B POR2X1_410/Y 0.00fF
C47818 POR2X1_126/CTRL2 POR2X1_4/Y 0.03fF
C47819 POR2X1_214/O POR2X1_214/B 0.01fF
C47820 D_INPUT_3 POR2X1_414/Y 0.02fF
C47821 POR2X1_376/B PAND2X1_341/A 0.02fF
C47822 POR2X1_215/O POR2X1_741/Y 0.02fF
C47823 PAND2X1_73/CTRL PAND2X1_63/B 0.01fF
C47824 POR2X1_46/Y PAND2X1_197/Y 0.03fF
C47825 POR2X1_128/CTRL2 POR2X1_222/Y 0.03fF
C47826 PAND2X1_449/Y VDD 0.05fF
C47827 POR2X1_174/O PAND2X1_73/Y 0.02fF
C47828 PAND2X1_553/B POR2X1_55/Y 0.09fF
C47829 PAND2X1_860/A POR2X1_677/Y 0.11fF
C47830 PAND2X1_93/B POR2X1_722/CTRL 0.06fF
C47831 POR2X1_809/A POR2X1_636/B 0.07fF
C47832 POR2X1_283/A POR2X1_331/Y 0.03fF
C47833 INPUT_1 POR2X1_267/A 0.20fF
C47834 POR2X1_614/A POR2X1_471/O 0.01fF
C47835 POR2X1_334/B POR2X1_786/A 0.10fF
C47836 POR2X1_401/a_16_28# POR2X1_401/A 0.03fF
C47837 POR2X1_537/Y PAND2X1_93/B 0.01fF
C47838 POR2X1_7/B PAND2X1_506/O 0.17fF
C47839 PAND2X1_151/m4_208_n4# PAND2X1_303/m4_208_n4# 0.15fF
C47840 POR2X1_294/B PAND2X1_144/CTRL2 0.02fF
C47841 INPUT_5 POR2X1_587/Y 0.03fF
C47842 POR2X1_445/O POR2X1_455/A 0.01fF
C47843 PAND2X1_139/O POR2X1_283/A 0.02fF
C47844 PAND2X1_6/Y PAND2X1_57/B 5.16fF
C47845 POR2X1_383/A POR2X1_862/B 0.03fF
C47846 POR2X1_333/a_16_28# PAND2X1_20/A 0.01fF
C47847 POR2X1_38/B POR2X1_236/a_16_28# 0.03fF
C47848 POR2X1_78/B PAND2X1_314/CTRL 0.06fF
C47849 POR2X1_750/Y POR2X1_750/A 0.01fF
C47850 PAND2X1_865/a_76_28# POR2X1_516/Y 0.02fF
C47851 POR2X1_174/A POR2X1_317/B 0.03fF
C47852 POR2X1_87/Y POR2X1_38/B 0.01fF
C47853 POR2X1_432/O POR2X1_129/Y 0.00fF
C47854 PAND2X1_469/Y PAND2X1_803/A 0.00fF
C47855 PAND2X1_643/O POR2X1_7/B 0.03fF
C47856 POR2X1_43/CTRL PAND2X1_838/B 0.01fF
C47857 POR2X1_776/A POR2X1_567/CTRL 0.01fF
C47858 POR2X1_686/B POR2X1_686/CTRL2 0.03fF
C47859 POR2X1_591/Y VDD 0.36fF
C47860 PAND2X1_793/Y POR2X1_816/A 0.01fF
C47861 POR2X1_65/A PAND2X1_244/B 0.03fF
C47862 POR2X1_115/O POR2X1_112/Y 0.02fF
C47863 POR2X1_814/B POR2X1_180/A 0.04fF
C47864 PAND2X1_254/Y POR2X1_256/Y 0.16fF
C47865 INPUT_0 POR2X1_9/CTRL 0.03fF
C47866 POR2X1_393/Y POR2X1_394/a_16_28# 0.03fF
C47867 INPUT_1 PAND2X1_614/O 0.04fF
C47868 POR2X1_278/Y PAND2X1_676/O 0.12fF
C47869 POR2X1_505/Y PAND2X1_507/CTRL2 0.00fF
C47870 POR2X1_220/Y POR2X1_573/A 0.03fF
C47871 POR2X1_857/A PAND2X1_52/B 0.00fF
C47872 POR2X1_101/Y POR2X1_573/CTRL2 0.23fF
C47873 POR2X1_367/CTRL POR2X1_568/Y 0.01fF
C47874 POR2X1_72/B PAND2X1_777/CTRL2 0.03fF
C47875 PAND2X1_48/B POR2X1_816/A 0.03fF
C47876 POR2X1_102/Y PAND2X1_156/A 0.03fF
C47877 PAND2X1_290/CTRL POR2X1_84/A 0.08fF
C47878 PAND2X1_20/A POR2X1_398/O 0.01fF
C47879 POR2X1_786/Y POR2X1_294/B 0.75fF
C47880 POR2X1_276/A POR2X1_325/A 0.01fF
C47881 PAND2X1_48/B POR2X1_462/B 0.04fF
C47882 PAND2X1_96/B POR2X1_554/Y 0.01fF
C47883 POR2X1_783/A POR2X1_780/A 0.06fF
C47884 POR2X1_68/A PAND2X1_275/O 0.15fF
C47885 PAND2X1_48/B D_INPUT_1 0.08fF
C47886 PAND2X1_23/Y POR2X1_778/B 0.03fF
C47887 POR2X1_537/Y POR2X1_78/A 0.10fF
C47888 POR2X1_558/CTRL2 PAND2X1_32/B 0.01fF
C47889 POR2X1_394/A PAND2X1_561/A 0.03fF
C47890 POR2X1_174/B POR2X1_502/Y 0.02fF
C47891 POR2X1_404/Y POR2X1_573/A 0.09fF
C47892 PAND2X1_150/O POR2X1_404/Y 0.08fF
C47893 POR2X1_52/A POR2X1_93/A 0.09fF
C47894 PAND2X1_73/Y PAND2X1_323/CTRL2 0.01fF
C47895 PAND2X1_675/a_76_28# POR2X1_283/A 0.02fF
C47896 PAND2X1_476/A POR2X1_32/A 0.02fF
C47897 PAND2X1_682/CTRL POR2X1_614/A 0.00fF
C47898 POR2X1_294/B POR2X1_788/B 0.12fF
C47899 POR2X1_52/A POR2X1_91/Y 0.15fF
C47900 POR2X1_51/B VDD 0.24fF
C47901 PAND2X1_65/B POR2X1_576/O 0.01fF
C47902 PAND2X1_341/B POR2X1_83/B 0.03fF
C47903 POR2X1_164/O POR2X1_693/Y 0.01fF
C47904 POR2X1_866/A PAND2X1_56/A 0.03fF
C47905 POR2X1_532/A PAND2X1_530/CTRL 0.01fF
C47906 POR2X1_8/Y POR2X1_381/CTRL 0.00fF
C47907 POR2X1_383/A PAND2X1_280/CTRL 0.03fF
C47908 POR2X1_327/Y POR2X1_686/A 0.02fF
C47909 POR2X1_327/Y POR2X1_860/A 0.11fF
C47910 PAND2X1_793/Y PAND2X1_854/A 0.02fF
C47911 POR2X1_590/A POR2X1_741/CTRL 0.01fF
C47912 POR2X1_83/B PAND2X1_352/Y 0.02fF
C47913 POR2X1_407/CTRL2 POR2X1_513/B 0.01fF
C47914 PAND2X1_6/Y POR2X1_828/A 0.26fF
C47915 PAND2X1_803/A POR2X1_394/A 0.03fF
C47916 POR2X1_152/A POR2X1_91/Y 0.03fF
C47917 POR2X1_557/A POR2X1_130/A 0.04fF
C47918 POR2X1_750/B POR2X1_735/O 0.04fF
C47919 POR2X1_38/B POR2X1_380/CTRL2 0.11fF
C47920 POR2X1_537/Y POR2X1_830/a_16_28# 0.02fF
C47921 PAND2X1_194/O POR2X1_42/Y 0.02fF
C47922 POR2X1_336/a_76_344# POR2X1_741/Y 0.01fF
C47923 PAND2X1_491/CTRL PAND2X1_32/B 0.01fF
C47924 VDD POR2X1_758/Y 0.01fF
C47925 POR2X1_855/B POR2X1_783/B 0.19fF
C47926 PAND2X1_41/B POR2X1_294/A 2.21fF
C47927 PAND2X1_632/B POR2X1_252/CTRL2 0.01fF
C47928 PAND2X1_231/a_76_28# POR2X1_153/Y 0.05fF
C47929 PAND2X1_650/A POR2X1_46/Y 0.02fF
C47930 POR2X1_532/A POR2X1_562/B 0.01fF
C47931 PAND2X1_655/Y PAND2X1_691/Y 0.04fF
C47932 PAND2X1_556/B PAND2X1_308/Y 0.03fF
C47933 PAND2X1_200/B POR2X1_236/Y 0.02fF
C47934 PAND2X1_23/Y POR2X1_854/B 0.09fF
C47935 POR2X1_614/A POR2X1_596/A 0.03fF
C47936 POR2X1_805/A PAND2X1_60/B 0.23fF
C47937 POR2X1_95/CTRL POR2X1_40/Y 0.01fF
C47938 POR2X1_795/B POR2X1_510/Y 0.07fF
C47939 PAND2X1_56/Y POR2X1_510/Y 0.05fF
C47940 PAND2X1_60/B POR2X1_712/Y 0.06fF
C47941 POR2X1_114/a_16_28# POR2X1_68/B 0.03fF
C47942 PAND2X1_96/B POR2X1_758/CTRL 0.01fF
C47943 POR2X1_776/B POR2X1_502/O 0.07fF
C47944 VDD POR2X1_741/A -0.00fF
C47945 PAND2X1_709/CTRL POR2X1_158/B 0.02fF
C47946 PAND2X1_61/a_76_28# POR2X1_39/B 0.03fF
C47947 PAND2X1_58/A POR2X1_39/B 0.03fF
C47948 POR2X1_502/A POR2X1_502/a_76_344# 0.03fF
C47949 PAND2X1_840/A PAND2X1_840/O -0.00fF
C47950 POR2X1_859/A POR2X1_753/O 0.33fF
C47951 POR2X1_51/A POR2X1_752/a_16_28# -0.00fF
C47952 POR2X1_13/A PAND2X1_560/B 0.03fF
C47953 POR2X1_130/Y POR2X1_141/A 0.09fF
C47954 GATE_741 PAND2X1_366/CTRL 0.01fF
C47955 PAND2X1_308/CTRL POR2X1_56/B 0.03fF
C47956 POR2X1_102/Y PAND2X1_339/O 0.02fF
C47957 POR2X1_327/Y POR2X1_327/CTRL2 0.01fF
C47958 POR2X1_846/A POR2X1_496/CTRL 0.01fF
C47959 POR2X1_548/A PAND2X1_69/A 0.01fF
C47960 PAND2X1_150/CTRL PAND2X1_60/B 0.01fF
C47961 PAND2X1_778/O PAND2X1_506/Y 0.07fF
C47962 POR2X1_695/CTRL2 POR2X1_425/Y 0.01fF
C47963 POR2X1_315/Y POR2X1_299/CTRL2 0.03fF
C47964 POR2X1_336/CTRL POR2X1_538/A 0.00fF
C47965 PAND2X1_469/B PAND2X1_353/a_76_28# 0.04fF
C47966 POR2X1_866/A POR2X1_661/A 0.07fF
C47967 PAND2X1_90/Y PAND2X1_759/CTRL 0.02fF
C47968 POR2X1_122/CTRL POR2X1_293/Y 0.01fF
C47969 POR2X1_362/Y PAND2X1_72/A 0.19fF
C47970 POR2X1_416/B PAND2X1_545/O 0.02fF
C47971 PAND2X1_108/CTRL2 POR2X1_862/B 0.00fF
C47972 PAND2X1_744/O POR2X1_260/A 0.04fF
C47973 POR2X1_557/A POR2X1_844/B 0.03fF
C47974 PAND2X1_771/B PAND2X1_771/a_16_344# 0.03fF
C47975 POR2X1_643/O POR2X1_260/B 0.02fF
C47976 POR2X1_379/O POR2X1_532/A 0.02fF
C47977 POR2X1_42/Y PAND2X1_853/B 0.03fF
C47978 INPUT_3 PAND2X1_87/a_16_344# 0.03fF
C47979 PAND2X1_504/CTRL POR2X1_507/A 0.04fF
C47980 PAND2X1_73/Y POR2X1_579/O 0.02fF
C47981 PAND2X1_464/B POR2X1_20/B 3.89fF
C47982 PAND2X1_373/O POR2X1_540/A 0.08fF
C47983 POR2X1_565/B POR2X1_266/A 0.00fF
C47984 POR2X1_119/Y PAND2X1_549/a_16_344# 0.02fF
C47985 INPUT_7 D_INPUT_4 0.03fF
C47986 POR2X1_844/B POR2X1_546/CTRL 0.01fF
C47987 PAND2X1_832/a_76_28# POR2X1_316/Y 0.02fF
C47988 POR2X1_614/A POR2X1_703/Y 0.03fF
C47989 POR2X1_750/B PAND2X1_681/CTRL 0.01fF
C47990 PAND2X1_333/CTRL2 POR2X1_77/Y 0.03fF
C47991 POR2X1_741/Y POR2X1_741/A 0.02fF
C47992 POR2X1_5/Y POR2X1_372/CTRL 0.01fF
C47993 POR2X1_383/A POR2X1_510/Y 0.07fF
C47994 POR2X1_571/CTRL POR2X1_844/B 0.01fF
C47995 PAND2X1_787/Y POR2X1_39/B 0.03fF
C47996 PAND2X1_476/A PAND2X1_35/Y 0.02fF
C47997 PAND2X1_6/Y POR2X1_259/B 0.06fF
C47998 POR2X1_477/A POR2X1_552/CTRL 0.15fF
C47999 POR2X1_612/A POR2X1_612/B 0.02fF
C48000 PAND2X1_691/Y PAND2X1_664/m4_208_n4# 0.12fF
C48001 PAND2X1_480/a_76_28# POR2X1_238/Y 0.02fF
C48002 PAND2X1_457/Y POR2X1_329/A 0.01fF
C48003 POR2X1_364/A POR2X1_333/Y 0.21fF
C48004 PAND2X1_171/O D_GATE_741 0.13fF
C48005 PAND2X1_555/O POR2X1_394/A 0.08fF
C48006 POR2X1_68/A POR2X1_62/Y 0.03fF
C48007 PAND2X1_661/B PAND2X1_560/B 0.03fF
C48008 POR2X1_180/B POR2X1_181/B 0.02fF
C48009 POR2X1_383/A POR2X1_276/Y 0.07fF
C48010 PAND2X1_23/Y POR2X1_374/CTRL2 0.01fF
C48011 POR2X1_702/A POR2X1_332/a_16_28# 0.01fF
C48012 POR2X1_324/A POR2X1_568/A 0.05fF
C48013 POR2X1_119/Y PAND2X1_798/B 0.05fF
C48014 PAND2X1_556/B POR2X1_77/Y 0.02fF
C48015 POR2X1_215/Y POR2X1_260/A 0.11fF
C48016 POR2X1_316/Y POR2X1_372/Y 0.07fF
C48017 PAND2X1_72/O PAND2X1_48/A 0.02fF
C48018 POR2X1_325/A POR2X1_325/B 0.04fF
C48019 INPUT_4 D_INPUT_4 0.33fF
C48020 POR2X1_63/Y POR2X1_813/O 0.03fF
C48021 POR2X1_442/a_76_344# POR2X1_411/B 0.01fF
C48022 PAND2X1_641/Y POR2X1_229/Y 0.02fF
C48023 POR2X1_63/a_16_28# POR2X1_62/Y 0.02fF
C48024 POR2X1_98/a_16_28# POR2X1_98/A 0.03fF
C48025 POR2X1_20/B POR2X1_20/A 0.01fF
C48026 POR2X1_68/B PAND2X1_48/A 0.04fF
C48027 POR2X1_96/A POR2X1_416/B 12.14fF
C48028 PAND2X1_865/Y PAND2X1_357/Y 0.07fF
C48029 PAND2X1_35/Y PAND2X1_327/CTRL2 0.01fF
C48030 POR2X1_338/CTRL2 POR2X1_334/Y 0.05fF
C48031 PAND2X1_476/A PAND2X1_651/Y 0.05fF
C48032 PAND2X1_57/B PAND2X1_52/B 0.06fF
C48033 PAND2X1_206/B POR2X1_29/A 0.03fF
C48034 POR2X1_610/Y POR2X1_610/CTRL2 0.01fF
C48035 POR2X1_83/B POR2X1_667/CTRL 0.00fF
C48036 POR2X1_62/Y PAND2X1_350/O 0.02fF
C48037 POR2X1_318/a_16_28# POR2X1_454/A 0.03fF
C48038 POR2X1_102/CTRL INPUT_2 0.01fF
C48039 POR2X1_102/O D_INPUT_1 0.02fF
C48040 PAND2X1_358/A PAND2X1_100/CTRL2 0.02fF
C48041 PAND2X1_481/CTRL2 POR2X1_260/A 0.03fF
C48042 INPUT_1 POR2X1_751/Y 0.03fF
C48043 POR2X1_16/A PAND2X1_704/O 0.04fF
C48044 POR2X1_66/B PAND2X1_75/CTRL2 0.01fF
C48045 PAND2X1_474/CTRL2 POR2X1_37/Y 0.03fF
C48046 PAND2X1_773/O POR2X1_767/Y 0.02fF
C48047 D_INPUT_1 PAND2X1_529/CTRL2 0.01fF
C48048 POR2X1_441/CTRL2 POR2X1_40/Y 0.03fF
C48049 POR2X1_490/Y PAND2X1_222/A 0.01fF
C48050 PAND2X1_182/B PAND2X1_336/a_76_28# 0.04fF
C48051 POR2X1_711/B POR2X1_710/Y 0.01fF
C48052 PAND2X1_482/CTRL POR2X1_260/A 0.01fF
C48053 POR2X1_130/A POR2X1_651/Y 0.07fF
C48054 PAND2X1_722/CTRL2 POR2X1_394/A 0.09fF
C48055 PAND2X1_126/a_56_28# POR2X1_62/Y 0.00fF
C48056 POR2X1_48/A PAND2X1_750/a_16_344# 0.02fF
C48057 POR2X1_704/Y POR2X1_317/B 0.01fF
C48058 POR2X1_73/Y PAND2X1_169/O 0.02fF
C48059 POR2X1_20/B POR2X1_751/A 0.06fF
C48060 POR2X1_593/CTRL POR2X1_449/A 0.01fF
C48061 POR2X1_49/Y POR2X1_441/CTRL 0.01fF
C48062 POR2X1_654/B POR2X1_814/A 0.02fF
C48063 PAND2X1_123/a_56_28# POR2X1_117/Y 0.00fF
C48064 PAND2X1_432/a_56_28# POR2X1_648/Y 0.00fF
C48065 PAND2X1_810/B POR2X1_283/Y 0.03fF
C48066 POR2X1_828/A PAND2X1_52/B 0.05fF
C48067 POR2X1_545/CTRL POR2X1_551/A 0.01fF
C48068 PAND2X1_67/CTRL POR2X1_296/B 0.07fF
C48069 PAND2X1_277/a_16_344# POR2X1_260/B 0.02fF
C48070 PAND2X1_856/B PAND2X1_863/A 0.18fF
C48071 POR2X1_825/CTRL POR2X1_20/B 0.01fF
C48072 POR2X1_38/Y POR2X1_522/O 0.10fF
C48073 POR2X1_814/A POR2X1_778/O 0.02fF
C48074 POR2X1_182/m4_208_n4# POR2X1_854/B 0.04fF
C48075 POR2X1_669/B POR2X1_260/B 0.05fF
C48076 POR2X1_557/B POR2X1_113/B 0.09fF
C48077 POR2X1_319/A POR2X1_78/A 0.10fF
C48078 POR2X1_116/A PAND2X1_41/B 0.03fF
C48079 PAND2X1_207/CTRL POR2X1_32/A 0.01fF
C48080 POR2X1_502/A POR2X1_463/CTRL2 0.01fF
C48081 POR2X1_568/Y POR2X1_568/CTRL 0.01fF
C48082 POR2X1_416/B POR2X1_7/A 0.06fF
C48083 PAND2X1_652/a_16_344# PAND2X1_593/Y 0.02fF
C48084 POR2X1_234/A POR2X1_518/Y 0.03fF
C48085 POR2X1_643/O PAND2X1_55/Y 0.03fF
C48086 POR2X1_423/Y POR2X1_253/O 0.01fF
C48087 POR2X1_257/A PAND2X1_541/CTRL 0.01fF
C48088 POR2X1_130/A POR2X1_646/A 0.02fF
C48089 POR2X1_634/A POR2X1_610/CTRL 0.01fF
C48090 POR2X1_482/CTRL POR2X1_669/B 0.02fF
C48091 PAND2X1_659/Y POR2X1_7/Y 0.03fF
C48092 D_INPUT_0 PAND2X1_591/a_76_28# 0.02fF
C48093 POR2X1_240/B POR2X1_66/A 0.27fF
C48094 POR2X1_356/A PAND2X1_52/CTRL 0.31fF
C48095 POR2X1_259/B POR2X1_632/Y 0.15fF
C48096 PAND2X1_205/Y PAND2X1_222/A 0.16fF
C48097 PAND2X1_272/O POR2X1_296/B 0.01fF
C48098 POR2X1_23/Y PAND2X1_575/B 0.04fF
C48099 POR2X1_556/A VDD 0.70fF
C48100 PAND2X1_639/a_56_28# POR2X1_408/Y 0.00fF
C48101 POR2X1_150/Y INPUT_0 0.03fF
C48102 POR2X1_257/A PAND2X1_276/O 0.01fF
C48103 POR2X1_257/A POR2X1_511/Y 0.03fF
C48104 POR2X1_294/A PAND2X1_122/O 0.02fF
C48105 POR2X1_848/A POR2X1_615/CTRL2 0.02fF
C48106 POR2X1_341/A POR2X1_573/a_76_344# 0.02fF
C48107 POR2X1_263/CTRL PAND2X1_35/Y 0.01fF
C48108 POR2X1_257/A POR2X1_524/Y 0.01fF
C48109 POR2X1_864/CTRL2 POR2X1_801/B 0.01fF
C48110 POR2X1_678/Y POR2X1_750/B 0.00fF
C48111 PAND2X1_358/A POR2X1_77/Y 0.03fF
C48112 POR2X1_46/CTRL POR2X1_409/B 0.01fF
C48113 POR2X1_863/A POR2X1_738/A 0.03fF
C48114 POR2X1_41/B POR2X1_441/Y 0.02fF
C48115 POR2X1_62/Y PAND2X1_529/CTRL 0.03fF
C48116 PAND2X1_609/CTRL PAND2X1_90/Y 0.01fF
C48117 POR2X1_69/CTRL2 POR2X1_29/A 0.11fF
C48118 PAND2X1_771/Y POR2X1_312/Y 0.23fF
C48119 POR2X1_456/B POR2X1_579/CTRL2 0.01fF
C48120 POR2X1_20/B PAND2X1_182/A 0.14fF
C48121 POR2X1_294/Y POR2X1_355/A 0.03fF
C48122 POR2X1_102/Y PAND2X1_215/CTRL 0.01fF
C48123 PAND2X1_474/CTRL2 POR2X1_293/Y 0.03fF
C48124 POR2X1_566/A POR2X1_443/A 0.04fF
C48125 POR2X1_78/B POR2X1_454/A 0.07fF
C48126 POR2X1_150/Y PAND2X1_717/CTRL2 0.01fF
C48127 POR2X1_525/Y POR2X1_20/B 0.03fF
C48128 POR2X1_202/CTRL2 POR2X1_296/B 0.02fF
C48129 POR2X1_814/B POR2X1_606/m4_208_n4# 0.15fF
C48130 POR2X1_826/Y POR2X1_293/Y 0.03fF
C48131 POR2X1_29/A POR2X1_750/B 0.10fF
C48132 POR2X1_227/O PAND2X1_52/B 0.09fF
C48133 POR2X1_13/A PAND2X1_436/CTRL2 0.03fF
C48134 PAND2X1_318/a_16_344# POR2X1_20/B 0.01fF
C48135 POR2X1_48/A PAND2X1_787/Y 0.05fF
C48136 PAND2X1_137/a_56_28# POR2X1_20/B 0.00fF
C48137 POR2X1_557/B POR2X1_768/A 0.16fF
C48138 POR2X1_18/CTRL D_INPUT_6 0.03fF
C48139 POR2X1_306/O POR2X1_329/A 0.03fF
C48140 POR2X1_556/A POR2X1_741/Y 4.54fF
C48141 POR2X1_376/B PAND2X1_68/a_16_344# 0.02fF
C48142 POR2X1_636/O POR2X1_750/B 0.01fF
C48143 POR2X1_89/m4_208_n4# PAND2X1_333/m4_208_n4# 0.13fF
C48144 POR2X1_68/A POR2X1_66/a_76_344# 0.01fF
C48145 D_INPUT_2 POR2X1_612/CTRL2 0.01fF
C48146 POR2X1_13/A PAND2X1_410/a_16_344# 0.01fF
C48147 POR2X1_479/B POR2X1_480/A 0.01fF
C48148 POR2X1_814/B POR2X1_267/CTRL 0.32fF
C48149 POR2X1_110/a_16_28# POR2X1_14/Y 0.02fF
C48150 POR2X1_669/B PAND2X1_803/A 0.03fF
C48151 POR2X1_260/B PAND2X1_751/CTRL 0.03fF
C48152 POR2X1_16/A PAND2X1_403/O 0.02fF
C48153 PAND2X1_742/CTRL POR2X1_331/Y 0.01fF
C48154 POR2X1_590/A POR2X1_830/A 0.03fF
C48155 PAND2X1_733/A POR2X1_40/Y 0.03fF
C48156 PAND2X1_58/A POR2X1_402/CTRL 0.01fF
C48157 POR2X1_788/A POR2X1_718/A 0.00fF
C48158 POR2X1_814/B POR2X1_673/CTRL2 0.07fF
C48159 POR2X1_411/B POR2X1_310/CTRL 0.01fF
C48160 POR2X1_602/CTRL POR2X1_294/B 0.04fF
C48161 POR2X1_556/A PAND2X1_32/B 0.11fF
C48162 PAND2X1_217/B POR2X1_72/B 0.60fF
C48163 POR2X1_487/O PAND2X1_580/B 0.00fF
C48164 POR2X1_831/CTRL POR2X1_513/Y 0.02fF
C48165 PAND2X1_23/Y POR2X1_862/A 1.40fF
C48166 POR2X1_613/CTRL POR2X1_55/Y 0.02fF
C48167 POR2X1_71/Y POR2X1_23/Y 0.67fF
C48168 POR2X1_12/A POR2X1_587/O 0.01fF
C48169 POR2X1_94/A PAND2X1_41/B 0.04fF
C48170 POR2X1_678/A POR2X1_718/A 0.03fF
C48171 POR2X1_87/Y POR2X1_590/A 0.01fF
C48172 POR2X1_624/Y PAND2X1_316/O 0.01fF
C48173 POR2X1_658/CTRL2 POR2X1_318/A 0.02fF
C48174 POR2X1_260/B POR2X1_459/m4_208_n4# 0.08fF
C48175 PAND2X1_3/A INPUT_5 0.06fF
C48176 POR2X1_467/Y POR2X1_448/B 0.00fF
C48177 PAND2X1_48/B PAND2X1_93/B 3.27fF
C48178 POR2X1_669/B PAND2X1_673/Y 0.19fF
C48179 POR2X1_314/O POR2X1_48/A 0.02fF
C48180 POR2X1_29/Y POR2X1_54/Y 0.04fF
C48181 POR2X1_257/A PAND2X1_324/O 0.16fF
C48182 POR2X1_126/CTRL2 D_INPUT_1 0.01fF
C48183 POR2X1_149/O POR2X1_532/A 0.01fF
C48184 POR2X1_113/Y POR2X1_499/A 0.15fF
C48185 POR2X1_23/Y POR2X1_42/Y 0.04fF
C48186 PAND2X1_20/A POR2X1_401/CTRL 0.01fF
C48187 POR2X1_313/Y PAND2X1_439/O 0.02fF
C48188 PAND2X1_630/CTRL2 POR2X1_48/A 0.01fF
C48189 PAND2X1_58/A POR2X1_459/CTRL 0.00fF
C48190 PAND2X1_104/CTRL2 INPUT_0 0.01fF
C48191 PAND2X1_95/CTRL2 POR2X1_66/A 0.01fF
C48192 POR2X1_428/Y PAND2X1_711/A 0.01fF
C48193 PAND2X1_65/B POR2X1_777/B 0.04fF
C48194 POR2X1_630/O POR2X1_222/Y 0.01fF
C48195 PAND2X1_651/Y PAND2X1_436/CTRL 0.01fF
C48196 PAND2X1_862/B PAND2X1_573/B 0.01fF
C48197 POR2X1_9/Y PAND2X1_156/A 0.10fF
C48198 PAND2X1_70/O POR2X1_750/B 0.02fF
C48199 D_INPUT_0 POR2X1_572/B 0.06fF
C48200 POR2X1_863/A PAND2X1_167/O 0.01fF
C48201 POR2X1_445/A POR2X1_540/A 0.02fF
C48202 POR2X1_49/Y POR2X1_511/Y 0.07fF
C48203 POR2X1_251/A VDD 0.24fF
C48204 POR2X1_20/B POR2X1_283/A 18.47fF
C48205 PAND2X1_557/A GATE_741 0.07fF
C48206 POR2X1_20/B PAND2X1_121/CTRL 0.01fF
C48207 PAND2X1_39/B PAND2X1_60/B 5.85fF
C48208 POR2X1_63/Y POR2X1_229/Y 0.71fF
C48209 POR2X1_72/B VDD 3.40fF
C48210 POR2X1_202/O VDD 0.00fF
C48211 POR2X1_43/B D_INPUT_0 0.15fF
C48212 PAND2X1_48/B POR2X1_78/A 0.13fF
C48213 PAND2X1_23/Y PAND2X1_73/Y 0.13fF
C48214 POR2X1_174/B POR2X1_785/A 0.05fF
C48215 POR2X1_517/Y POR2X1_83/B 0.01fF
C48216 POR2X1_648/A PAND2X1_48/A 0.00fF
C48217 PAND2X1_805/A PAND2X1_366/Y 0.01fF
C48218 PAND2X1_159/CTRL2 POR2X1_55/Y 0.00fF
C48219 PAND2X1_804/B POR2X1_40/Y 0.07fF
C48220 POR2X1_257/A PAND2X1_112/CTRL2 0.06fF
C48221 POR2X1_614/A D_INPUT_0 0.27fF
C48222 POR2X1_499/A POR2X1_260/A 0.03fF
C48223 PAND2X1_59/B PAND2X1_26/CTRL 0.01fF
C48224 POR2X1_614/A POR2X1_811/A 0.03fF
C48225 POR2X1_20/B PAND2X1_100/O 0.01fF
C48226 PAND2X1_669/O POR2X1_816/A 0.02fF
C48227 POR2X1_677/O INPUT_0 0.04fF
C48228 POR2X1_850/B POR2X1_740/Y 0.03fF
C48229 POR2X1_218/Y POR2X1_804/A 0.10fF
C48230 POR2X1_472/CTRL2 POR2X1_862/A 0.02fF
C48231 POR2X1_825/Y POR2X1_39/B 0.09fF
C48232 PAND2X1_669/O D_INPUT_1 0.01fF
C48233 POR2X1_43/B PAND2X1_435/Y 0.02fF
C48234 POR2X1_192/Y POR2X1_776/CTRL 0.01fF
C48235 POR2X1_66/B POR2X1_138/CTRL 0.01fF
C48236 POR2X1_814/B POR2X1_572/O 0.34fF
C48237 INPUT_1 PAND2X1_247/O 0.04fF
C48238 POR2X1_48/A POR2X1_280/O 0.03fF
C48239 D_INPUT_0 POR2X1_38/B 0.06fF
C48240 POR2X1_549/B POR2X1_547/B 0.27fF
C48241 INPUT_3 POR2X1_376/CTRL 0.06fF
C48242 POR2X1_852/B POR2X1_852/A 0.02fF
C48243 PAND2X1_20/A POR2X1_574/CTRL 0.01fF
C48244 PAND2X1_845/CTRL2 POR2X1_83/B 0.03fF
C48245 POR2X1_123/CTRL2 PAND2X1_41/B 0.00fF
C48246 POR2X1_96/A PAND2X1_192/Y 0.05fF
C48247 POR2X1_307/B POR2X1_130/A 0.01fF
C48248 POR2X1_46/Y PAND2X1_706/m4_208_n4# 0.09fF
C48249 PAND2X1_798/B PAND2X1_798/a_76_28# 0.02fF
C48250 POR2X1_290/CTRL POR2X1_290/Y 0.08fF
C48251 POR2X1_781/a_16_28# POR2X1_781/B 0.06fF
C48252 PAND2X1_51/CTRL2 POR2X1_635/A 0.01fF
C48253 INPUT_1 PAND2X1_407/CTRL 0.01fF
C48254 POR2X1_400/A VDD 0.06fF
C48255 POR2X1_322/O POR2X1_72/B 0.01fF
C48256 POR2X1_294/B POR2X1_788/O 0.04fF
C48257 POR2X1_839/a_16_28# POR2X1_835/Y 0.02fF
C48258 POR2X1_852/CTRL2 POR2X1_776/B 0.04fF
C48259 POR2X1_76/A POR2X1_260/A 0.03fF
C48260 PAND2X1_810/B PAND2X1_365/A 0.01fF
C48261 PAND2X1_6/Y POR2X1_244/CTRL 0.00fF
C48262 POR2X1_555/A POR2X1_785/A 0.07fF
C48263 PAND2X1_275/CTRL POR2X1_274/Y 0.02fF
C48264 PAND2X1_573/CTRL2 PAND2X1_735/Y 0.03fF
C48265 POR2X1_66/B PAND2X1_252/CTRL 0.03fF
C48266 POR2X1_257/A POR2X1_129/Y 0.21fF
C48267 POR2X1_634/A POR2X1_771/O 0.10fF
C48268 POR2X1_78/B POR2X1_360/A 0.20fF
C48269 PAND2X1_472/B PAND2X1_8/Y 0.05fF
C48270 PAND2X1_407/CTRL POR2X1_153/Y 0.03fF
C48271 POR2X1_270/Y PAND2X1_368/O 0.18fF
C48272 PAND2X1_635/O POR2X1_748/A 0.01fF
C48273 POR2X1_96/A PAND2X1_738/Y 0.05fF
C48274 POR2X1_83/A POR2X1_46/a_16_28# 0.03fF
C48275 PAND2X1_216/CTRL VDD 0.00fF
C48276 POR2X1_446/B POR2X1_317/B 0.00fF
C48277 POR2X1_302/A POR2X1_850/A 0.43fF
C48278 POR2X1_470/O POR2X1_854/B 0.08fF
C48279 POR2X1_805/Y PAND2X1_60/B 0.02fF
C48280 INPUT_0 PAND2X1_364/B 0.42fF
C48281 POR2X1_48/A PAND2X1_114/O 0.04fF
C48282 PAND2X1_58/A POR2X1_550/a_16_28# 0.03fF
C48283 POR2X1_505/CTRL POR2X1_48/A 0.01fF
C48284 POR2X1_13/A POR2X1_13/a_16_28# 0.10fF
C48285 POR2X1_45/O POR2X1_42/Y 0.08fF
C48286 POR2X1_548/B VDD 0.23fF
C48287 POR2X1_41/B POR2X1_625/Y 0.07fF
C48288 PAND2X1_20/A PAND2X1_60/B 4.16fF
C48289 POR2X1_52/A POR2X1_418/a_16_28# 0.03fF
C48290 POR2X1_323/Y VDD 0.05fF
C48291 PAND2X1_74/a_56_28# POR2X1_532/A 0.00fF
C48292 GATE_479 PAND2X1_565/A 0.03fF
C48293 POR2X1_55/Y PAND2X1_8/Y 0.03fF
C48294 PAND2X1_827/CTRL POR2X1_507/A 0.04fF
C48295 PAND2X1_293/CTRL PAND2X1_55/Y 0.02fF
C48296 POR2X1_60/O POR2X1_60/Y 0.01fF
C48297 PAND2X1_573/CTRL POR2X1_494/Y 0.00fF
C48298 PAND2X1_659/Y POR2X1_257/A 0.09fF
C48299 PAND2X1_76/Y POR2X1_255/Y 0.00fF
C48300 POR2X1_262/CTRL2 PAND2X1_215/B 0.00fF
C48301 PAND2X1_612/B POR2X1_773/A 0.00fF
C48302 POR2X1_500/A POR2X1_318/A 0.17fF
C48303 PAND2X1_55/Y POR2X1_404/B 0.01fF
C48304 POR2X1_69/CTRL POR2X1_7/A 0.01fF
C48305 POR2X1_614/A PAND2X1_90/Y 0.29fF
C48306 PAND2X1_6/Y PAND2X1_85/Y 0.00fF
C48307 PAND2X1_96/B POR2X1_402/CTRL 0.01fF
C48308 POR2X1_317/Y PAND2X1_90/Y 0.04fF
C48309 PAND2X1_390/Y POR2X1_172/Y 0.03fF
C48310 PAND2X1_865/a_16_344# POR2X1_32/A 0.01fF
C48311 PAND2X1_95/B PAND2X1_57/B 0.88fF
C48312 PAND2X1_223/B PAND2X1_539/Y 0.03fF
C48313 PAND2X1_341/B PAND2X1_206/A 0.00fF
C48314 POR2X1_606/O PAND2X1_48/A 0.01fF
C48315 PAND2X1_96/CTRL PAND2X1_60/B 0.01fF
C48316 POR2X1_672/CTRL2 VDD 0.00fF
C48317 PAND2X1_652/Y PAND2X1_592/Y 0.01fF
C48318 POR2X1_416/B POR2X1_760/A 4.98fF
C48319 POR2X1_332/B D_GATE_222 0.12fF
C48320 POR2X1_16/A PAND2X1_443/Y 0.01fF
C48321 PAND2X1_89/O POR2X1_785/A 0.01fF
C48322 POR2X1_38/B PAND2X1_90/Y 0.03fF
C48323 POR2X1_122/Y POR2X1_73/Y 0.07fF
C48324 POR2X1_57/A PAND2X1_768/Y 0.02fF
C48325 PAND2X1_52/O PAND2X1_52/B 0.00fF
C48326 PAND2X1_218/CTRL PAND2X1_364/B 0.03fF
C48327 POR2X1_814/B PAND2X1_60/B 0.29fF
C48328 POR2X1_719/B PAND2X1_73/Y 0.01fF
C48329 POR2X1_294/B POR2X1_193/CTRL2 0.04fF
C48330 PAND2X1_835/Y VDD 0.00fF
C48331 PAND2X1_675/A PAND2X1_793/Y 0.03fF
C48332 POR2X1_243/CTRL2 INPUT_0 0.00fF
C48333 POR2X1_135/Y PAND2X1_702/O 0.01fF
C48334 POR2X1_65/A PAND2X1_656/A 0.03fF
C48335 PAND2X1_793/Y PAND2X1_469/B 0.03fF
C48336 POR2X1_441/Y POR2X1_77/Y 0.03fF
C48337 PAND2X1_380/O POR2X1_532/A 0.01fF
C48338 PAND2X1_65/B POR2X1_712/O 0.01fF
C48339 POR2X1_85/a_16_28# POR2X1_20/B 0.02fF
C48340 POR2X1_207/B VDD 0.03fF
C48341 POR2X1_115/CTRL POR2X1_804/A 0.14fF
C48342 PAND2X1_20/A POR2X1_546/O 0.01fF
C48343 POR2X1_40/Y PAND2X1_124/CTRL 0.09fF
C48344 POR2X1_8/Y POR2X1_104/O 0.01fF
C48345 POR2X1_16/A PAND2X1_557/A 0.10fF
C48346 POR2X1_252/Y POR2X1_23/Y 0.09fF
C48347 POR2X1_410/Y VDD 0.11fF
C48348 PAND2X1_57/B PAND2X1_743/O 0.15fF
C48349 POR2X1_57/A PAND2X1_139/B 0.05fF
C48350 PAND2X1_20/A POR2X1_571/O 0.01fF
C48351 POR2X1_396/Y POR2X1_236/Y 0.00fF
C48352 POR2X1_175/A POR2X1_175/B 0.01fF
C48353 PAND2X1_568/a_76_28# PAND2X1_566/Y 0.02fF
C48354 POR2X1_462/B POR2X1_790/O 0.01fF
C48355 POR2X1_327/Y POR2X1_121/B 0.04fF
C48356 POR2X1_480/A POR2X1_537/B 0.01fF
C48357 POR2X1_325/A PAND2X1_60/B 0.03fF
C48358 POR2X1_239/CTRL2 POR2X1_7/B 0.00fF
C48359 POR2X1_809/A PAND2X1_73/Y 0.02fF
C48360 PAND2X1_23/Y POR2X1_249/CTRL2 0.03fF
C48361 POR2X1_135/O POR2X1_48/A 0.02fF
C48362 PAND2X1_471/CTRL2 PAND2X1_241/Y 0.01fF
C48363 POR2X1_220/B POR2X1_357/B 0.09fF
C48364 POR2X1_57/A POR2X1_45/a_16_28# 0.05fF
C48365 PAND2X1_48/B PAND2X1_145/a_76_28# 0.01fF
C48366 POR2X1_355/B POR2X1_209/A 0.03fF
C48367 POR2X1_570/a_16_28# POR2X1_570/B 0.03fF
C48368 POR2X1_750/Y PAND2X1_526/O -0.01fF
C48369 PAND2X1_862/B POR2X1_91/Y 0.01fF
C48370 PAND2X1_570/B VDD 0.04fF
C48371 PAND2X1_393/O VDD 0.00fF
C48372 POR2X1_137/O PAND2X1_32/B 0.18fF
C48373 POR2X1_16/A POR2X1_238/CTRL2 0.01fF
C48374 PAND2X1_773/a_76_28# POR2X1_7/B 0.01fF
C48375 POR2X1_62/Y PAND2X1_58/A 0.07fF
C48376 PAND2X1_691/Y POR2X1_829/Y 0.01fF
C48377 POR2X1_276/A VDD 0.21fF
C48378 POR2X1_43/B POR2X1_277/a_16_28# 0.02fF
C48379 PAND2X1_650/CTRL POR2X1_46/Y 0.01fF
C48380 POR2X1_334/O POR2X1_814/B 0.01fF
C48381 PAND2X1_783/m4_208_n4# POR2X1_90/Y 0.15fF
C48382 VDD POR2X1_566/B 2.77fF
C48383 POR2X1_662/Y PAND2X1_96/B 6.95fF
C48384 POR2X1_271/O POR2X1_39/B 0.01fF
C48385 POR2X1_301/CTRL PAND2X1_6/Y 0.15fF
C48386 POR2X1_102/Y POR2X1_171/Y 0.16fF
C48387 VDD POR2X1_180/A 0.19fF
C48388 POR2X1_178/O PAND2X1_675/A 0.01fF
C48389 POR2X1_222/Y POR2X1_702/A 0.03fF
C48390 POR2X1_65/A PAND2X1_348/A 0.07fF
C48391 POR2X1_717/CTRL POR2X1_717/Y 0.01fF
C48392 POR2X1_513/B PAND2X1_60/B 0.03fF
C48393 POR2X1_469/CTRL POR2X1_478/B 0.00fF
C48394 POR2X1_49/Y POR2X1_129/Y 0.03fF
C48395 POR2X1_835/CTRL2 POR2X1_835/B 0.03fF
C48396 POR2X1_790/B PAND2X1_69/A 0.03fF
C48397 POR2X1_68/A POR2X1_804/A 0.05fF
C48398 PAND2X1_651/Y POR2X1_521/CTRL 0.01fF
C48399 POR2X1_722/Y POR2X1_513/a_16_28# 0.02fF
C48400 POR2X1_502/A POR2X1_796/A 0.03fF
C48401 PAND2X1_444/a_76_28# POR2X1_39/B 0.02fF
C48402 POR2X1_166/m4_208_n4# PAND2X1_544/m4_208_n4# 0.05fF
C48403 POR2X1_783/A POR2X1_796/A 0.04fF
C48404 PAND2X1_532/CTRL VDD 0.00fF
C48405 POR2X1_663/CTRL POR2X1_544/B 0.02fF
C48406 POR2X1_188/a_16_28# POR2X1_220/Y 0.01fF
C48407 POR2X1_110/Y PAND2X1_465/O 0.01fF
C48408 POR2X1_572/B POR2X1_361/O 0.02fF
C48409 PAND2X1_844/B POR2X1_521/CTRL 0.01fF
C48410 POR2X1_787/a_16_28# POR2X1_325/A 0.02fF
C48411 PAND2X1_555/Y PAND2X1_566/Y 0.34fF
C48412 POR2X1_49/Y PAND2X1_659/Y 0.03fF
C48413 PAND2X1_20/A POR2X1_554/O 0.01fF
C48414 POR2X1_691/B POR2X1_800/A 0.00fF
C48415 PAND2X1_496/O POR2X1_569/A 0.10fF
C48416 POR2X1_741/Y POR2X1_702/O 0.01fF
C48417 POR2X1_532/A POR2X1_702/A 0.03fF
C48418 PAND2X1_291/O POR2X1_35/Y 0.02fF
C48419 PAND2X1_678/a_16_344# POR2X1_677/Y 0.02fF
C48420 POR2X1_219/O PAND2X1_88/Y 0.01fF
C48421 PAND2X1_73/Y POR2X1_711/Y 0.03fF
C48422 PAND2X1_291/CTRL2 PAND2X1_69/A 0.03fF
C48423 POR2X1_564/Y POR2X1_703/Y 0.07fF
C48424 PAND2X1_95/B POR2X1_707/Y 0.01fF
C48425 PAND2X1_139/Y PAND2X1_853/B 0.00fF
C48426 POR2X1_49/Y POR2X1_96/Y 0.03fF
C48427 POR2X1_476/Y POR2X1_294/A 0.02fF
C48428 POR2X1_480/A PAND2X1_48/A 2.89fF
C48429 PAND2X1_602/Y POR2X1_755/m4_208_n4# 0.12fF
C48430 POR2X1_280/Y PAND2X1_552/B 0.03fF
C48431 PAND2X1_216/B PAND2X1_216/a_16_344# 0.05fF
C48432 POR2X1_433/Y PAND2X1_349/A 0.03fF
C48433 POR2X1_65/A PAND2X1_631/A 0.03fF
C48434 POR2X1_86/O POR2X1_40/Y 0.01fF
C48435 PAND2X1_825/CTRL POR2X1_402/A 0.01fF
C48436 PAND2X1_96/B POR2X1_194/a_16_28# 0.01fF
C48437 POR2X1_139/a_16_28# POR2X1_137/Y -0.00fF
C48438 POR2X1_244/B POR2X1_227/CTRL 0.01fF
C48439 POR2X1_119/Y POR2X1_666/A 0.20fF
C48440 POR2X1_416/B PAND2X1_556/CTRL2 0.01fF
C48441 POR2X1_712/A POR2X1_383/A 0.00fF
C48442 POR2X1_327/Y PAND2X1_760/a_16_344# 0.02fF
C48443 POR2X1_311/Y POR2X1_416/B 0.03fF
C48444 POR2X1_78/B POR2X1_571/Y 0.53fF
C48445 PAND2X1_389/a_16_344# POR2X1_387/Y 0.01fF
C48446 POR2X1_702/O PAND2X1_32/B 0.06fF
C48447 PAND2X1_797/Y PAND2X1_714/A 0.01fF
C48448 PAND2X1_25/O PAND2X1_72/A 0.01fF
C48449 POR2X1_65/A POR2X1_86/CTRL 0.01fF
C48450 POR2X1_399/Y POR2X1_20/B 0.02fF
C48451 POR2X1_68/A PAND2X1_6/CTRL2 0.10fF
C48452 PAND2X1_283/CTRL POR2X1_773/B 0.08fF
C48453 POR2X1_78/B POR2X1_99/B 0.05fF
C48454 POR2X1_406/Y POR2X1_7/Y 0.03fF
C48455 PAND2X1_213/B PAND2X1_162/A 0.02fF
C48456 POR2X1_422/Y POR2X1_387/a_16_28# 0.01fF
C48457 PAND2X1_96/B POR2X1_181/B 0.01fF
C48458 POR2X1_566/B PAND2X1_32/B 4.88fF
C48459 POR2X1_148/B POR2X1_148/A 0.05fF
C48460 POR2X1_222/A POR2X1_573/A 0.03fF
C48461 POR2X1_265/Y PAND2X1_734/B 0.00fF
C48462 POR2X1_508/B VDD 0.01fF
C48463 PAND2X1_653/Y POR2X1_7/CTRL2 0.04fF
C48464 PAND2X1_717/A POR2X1_411/B 0.03fF
C48465 PAND2X1_285/O POR2X1_281/Y 0.00fF
C48466 POR2X1_554/Y POR2X1_735/CTRL2 0.01fF
C48467 POR2X1_798/O POR2X1_568/B 0.33fF
C48468 POR2X1_79/Y PAND2X1_730/A 0.12fF
C48469 PAND2X1_290/CTRL2 PAND2X1_85/Y 0.03fF
C48470 POR2X1_360/A POR2X1_294/A 0.10fF
C48471 POR2X1_814/A PAND2X1_268/CTRL 0.01fF
C48472 POR2X1_772/CTRL2 PAND2X1_32/B 0.08fF
C48473 PAND2X1_298/CTRL PAND2X1_32/B 0.01fF
C48474 POR2X1_600/a_56_344# POR2X1_411/B 0.00fF
C48475 POR2X1_136/Y POR2X1_7/A 0.00fF
C48476 POR2X1_327/Y PAND2X1_56/Y 0.10fF
C48477 PAND2X1_349/A PAND2X1_840/CTRL 0.01fF
C48478 PAND2X1_90/A PAND2X1_48/A 0.08fF
C48479 POR2X1_763/Y POR2X1_320/CTRL 0.06fF
C48480 POR2X1_49/Y PAND2X1_333/Y 0.09fF
C48481 POR2X1_136/CTRL PAND2X1_348/A 0.04fF
C48482 POR2X1_329/A PAND2X1_222/A 0.03fF
C48483 POR2X1_96/A PAND2X1_802/a_76_28# 0.01fF
C48484 POR2X1_274/B POR2X1_366/A 0.03fF
C48485 PAND2X1_476/A POR2X1_406/CTRL2 0.00fF
C48486 POR2X1_343/A PAND2X1_52/B 0.00fF
C48487 POR2X1_16/A PAND2X1_350/CTRL2 0.00fF
C48488 PAND2X1_844/Y PAND2X1_338/CTRL 0.01fF
C48489 PAND2X1_498/O POR2X1_188/Y 0.00fF
C48490 POR2X1_208/A POR2X1_215/A 0.17fF
C48491 POR2X1_713/O POR2X1_294/A 0.02fF
C48492 POR2X1_567/A POR2X1_231/a_76_344# 0.01fF
C48493 PAND2X1_291/CTRL2 PAND2X1_824/B 0.01fF
C48494 POR2X1_834/Y POR2X1_832/A 0.07fF
C48495 POR2X1_270/m4_208_n4# POR2X1_456/B 0.08fF
C48496 POR2X1_569/A POR2X1_576/CTRL2 0.03fF
C48497 POR2X1_327/Y POR2X1_336/O 0.02fF
C48498 PAND2X1_7/O POR2X1_99/B 0.00fF
C48499 PAND2X1_18/O PAND2X1_52/B 0.24fF
C48500 PAND2X1_480/O POR2X1_91/Y 0.04fF
C48501 POR2X1_420/CTRL POR2X1_329/A 0.04fF
C48502 PAND2X1_508/Y POR2X1_73/Y 0.10fF
C48503 POR2X1_539/A POR2X1_260/A 0.06fF
C48504 POR2X1_283/A PAND2X1_715/B 0.01fF
C48505 POR2X1_416/B POR2X1_609/A 0.03fF
C48506 PAND2X1_788/a_76_28# POR2X1_533/Y 0.05fF
C48507 POR2X1_648/Y POR2X1_807/O 0.02fF
C48508 POR2X1_369/Y PAND2X1_566/Y 0.00fF
C48509 VDD POR2X1_325/B 0.11fF
C48510 POR2X1_248/m4_208_n4# POR2X1_153/Y 0.03fF
C48511 POR2X1_655/Y POR2X1_661/A 0.02fF
C48512 PAND2X1_341/A PAND2X1_716/B 0.00fF
C48513 PAND2X1_357/Y PAND2X1_352/Y 0.01fF
C48514 PAND2X1_838/B PAND2X1_838/a_76_28# 0.02fF
C48515 POR2X1_334/Y POR2X1_228/Y 0.03fF
C48516 PAND2X1_631/A POR2X1_136/CTRL 0.08fF
C48517 POR2X1_567/A POR2X1_556/Y 0.05fF
C48518 PAND2X1_69/A POR2X1_540/Y 0.03fF
C48519 PAND2X1_90/O POR2X1_68/B 0.03fF
C48520 POR2X1_327/Y POR2X1_383/A 0.61fF
C48521 POR2X1_639/Y PAND2X1_328/O 0.04fF
C48522 POR2X1_38/Y PAND2X1_120/a_76_28# 0.02fF
C48523 POR2X1_332/Y PAND2X1_60/B 0.03fF
C48524 PAND2X1_716/B POR2X1_91/Y 0.03fF
C48525 POR2X1_283/A PAND2X1_502/CTRL 0.04fF
C48526 POR2X1_245/a_16_28# POR2X1_129/Y 0.02fF
C48527 POR2X1_12/A POR2X1_582/Y 0.00fF
C48528 POR2X1_735/O POR2X1_318/A 0.04fF
C48529 PAND2X1_96/B PAND2X1_134/CTRL 0.01fF
C48530 POR2X1_461/Y POR2X1_848/A 0.25fF
C48531 POR2X1_540/A POR2X1_181/CTRL2 0.03fF
C48532 POR2X1_458/Y POR2X1_330/Y 0.10fF
C48533 POR2X1_567/A POR2X1_854/CTRL2 -0.00fF
C48534 POR2X1_555/A PAND2X1_628/O 0.06fF
C48535 PAND2X1_165/CTRL2 POR2X1_854/B 0.18fF
C48536 POR2X1_680/O POR2X1_594/A 0.10fF
C48537 PAND2X1_394/CTRL2 POR2X1_215/A 0.05fF
C48538 POR2X1_842/CTRL2 PAND2X1_39/B 0.03fF
C48539 PAND2X1_472/A POR2X1_39/B 0.10fF
C48540 POR2X1_66/Y POR2X1_195/A 0.01fF
C48541 PAND2X1_717/A POR2X1_271/Y 0.03fF
C48542 PAND2X1_20/O PAND2X1_19/Y 0.00fF
C48543 POR2X1_840/CTRL2 POR2X1_513/A 0.00fF
C48544 POR2X1_502/A POR2X1_863/A 0.03fF
C48545 POR2X1_309/CTRL2 POR2X1_150/Y 0.03fF
C48546 PAND2X1_458/CTRL POR2X1_5/Y 0.01fF
C48547 PAND2X1_601/CTRL2 PAND2X1_93/B 0.03fF
C48548 POR2X1_396/a_16_28# POR2X1_39/B 0.01fF
C48549 POR2X1_773/A POR2X1_773/CTRL 0.00fF
C48550 POR2X1_257/A POR2X1_37/Y 0.87fF
C48551 POR2X1_814/A POR2X1_777/B 0.03fF
C48552 POR2X1_514/Y PAND2X1_72/A 0.03fF
C48553 POR2X1_369/Y POR2X1_315/Y 0.01fF
C48554 POR2X1_316/CTRL POR2X1_129/Y 0.01fF
C48555 POR2X1_150/Y POR2X1_102/Y 1.93fF
C48556 POR2X1_332/Y POR2X1_332/O 0.00fF
C48557 PAND2X1_94/Y VDD 0.11fF
C48558 PAND2X1_189/m4_208_n4# POR2X1_353/A 0.12fF
C48559 POR2X1_840/Y POR2X1_725/Y 0.01fF
C48560 POR2X1_14/Y POR2X1_20/B 0.15fF
C48561 POR2X1_507/B POR2X1_507/A 0.05fF
C48562 POR2X1_416/B POR2X1_38/Y 0.06fF
C48563 PAND2X1_404/Y POR2X1_409/B 0.03fF
C48564 POR2X1_376/B PAND2X1_717/A 0.01fF
C48565 POR2X1_325/B PAND2X1_32/B 0.01fF
C48566 PAND2X1_65/B POR2X1_814/A 0.22fF
C48567 POR2X1_241/O POR2X1_776/A 0.03fF
C48568 POR2X1_711/Y PAND2X1_306/CTRL 0.04fF
C48569 POR2X1_502/A POR2X1_9/Y 0.41fF
C48570 POR2X1_478/a_16_28# POR2X1_477/Y 0.03fF
C48571 PAND2X1_649/A POR2X1_394/CTRL 0.01fF
C48572 POR2X1_551/a_16_28# POR2X1_551/A 0.06fF
C48573 PAND2X1_865/Y PAND2X1_579/A 0.00fF
C48574 PAND2X1_69/A POR2X1_343/B 0.03fF
C48575 PAND2X1_65/B PAND2X1_256/CTRL2 0.00fF
C48576 POR2X1_20/B POR2X1_279/Y 0.01fF
C48577 POR2X1_527/Y POR2X1_39/B 0.00fF
C48578 POR2X1_46/O PAND2X1_9/Y 0.01fF
C48579 PAND2X1_65/B POR2X1_846/Y 0.03fF
C48580 POR2X1_58/Y POR2X1_9/Y 0.05fF
C48581 POR2X1_19/CTRL POR2X1_5/Y 0.01fF
C48582 PAND2X1_31/a_76_28# PAND2X1_3/A 0.01fF
C48583 PAND2X1_47/B PAND2X1_31/CTRL2 0.00fF
C48584 PAND2X1_716/B POR2X1_109/Y 0.03fF
C48585 PAND2X1_93/B POR2X1_632/B 0.18fF
C48586 PAND2X1_313/O POR2X1_169/A 0.02fF
C48587 D_GATE_662 PAND2X1_438/CTRL 0.03fF
C48588 POR2X1_52/A PAND2X1_717/A 0.08fF
C48589 D_INPUT_0 POR2X1_590/A 1.07fF
C48590 POR2X1_271/B POR2X1_236/Y 0.87fF
C48591 POR2X1_56/B POR2X1_329/A 0.09fF
C48592 POR2X1_707/B PAND2X1_762/a_16_344# 0.01fF
C48593 INPUT_1 POR2X1_416/B 0.14fF
C48594 POR2X1_19/O PAND2X1_8/Y 0.06fF
C48595 POR2X1_83/B POR2X1_427/CTRL2 0.03fF
C48596 POR2X1_86/Y PAND2X1_100/O 0.18fF
C48597 PAND2X1_611/a_76_28# POR2X1_130/A 0.04fF
C48598 POR2X1_669/B POR2X1_626/a_16_28# 0.09fF
C48599 POR2X1_286/B POR2X1_476/Y 0.06fF
C48600 PAND2X1_48/A PAND2X1_304/O 0.03fF
C48601 PAND2X1_717/A POR2X1_152/A 0.01fF
C48602 POR2X1_773/B PAND2X1_72/A 0.03fF
C48603 PAND2X1_435/CTRL POR2X1_411/B 0.01fF
C48604 PAND2X1_698/a_16_344# PAND2X1_52/B 0.05fF
C48605 POR2X1_603/Y POR2X1_32/A 0.09fF
C48606 POR2X1_804/O POR2X1_330/Y 0.09fF
C48607 POR2X1_416/B POR2X1_153/Y 0.10fF
C48608 POR2X1_60/A POR2X1_432/O 0.03fF
C48609 POR2X1_66/A PAND2X1_16/CTRL2 0.01fF
C48610 POR2X1_41/B POR2X1_411/B 1.30fF
C48611 POR2X1_66/B PAND2X1_39/CTRL2 0.03fF
C48612 POR2X1_66/A POR2X1_404/O 0.00fF
C48613 PAND2X1_865/CTRL2 PAND2X1_860/A 0.01fF
C48614 POR2X1_49/Y PAND2X1_448/CTRL 0.08fF
C48615 POR2X1_49/Y POR2X1_37/Y 0.12fF
C48616 PAND2X1_414/CTRL PAND2X1_6/A 0.01fF
C48617 POR2X1_614/A PAND2X1_426/CTRL2 0.00fF
C48618 POR2X1_287/B POR2X1_476/A 0.03fF
C48619 PAND2X1_205/A PAND2X1_204/CTRL 0.00fF
C48620 POR2X1_505/Y POR2X1_669/B 0.03fF
C48621 POR2X1_20/B POR2X1_55/Y 1.73fF
C48622 POR2X1_311/Y POR2X1_487/Y 0.00fF
C48623 POR2X1_39/CTRL POR2X1_669/B 0.01fF
C48624 POR2X1_629/B POR2X1_630/A 0.05fF
C48625 PAND2X1_20/A POR2X1_254/A 0.03fF
C48626 POR2X1_586/Y POR2X1_752/Y 0.03fF
C48627 PAND2X1_52/B PAND2X1_18/B 0.05fF
C48628 POR2X1_257/A POR2X1_293/Y 0.10fF
C48629 POR2X1_257/A PAND2X1_555/A 0.05fF
C48630 PAND2X1_20/A POR2X1_750/B 0.08fF
C48631 POR2X1_83/B POR2X1_423/Y 5.19fF
C48632 POR2X1_459/Y PAND2X1_752/Y 0.02fF
C48633 POR2X1_555/B PAND2X1_52/Y 2.43fF
C48634 PAND2X1_71/a_16_344# PAND2X1_39/B 0.01fF
C48635 PAND2X1_94/A POR2X1_643/CTRL 0.00fF
C48636 PAND2X1_640/B VDD 0.92fF
C48637 POR2X1_496/Y POR2X1_5/Y 0.07fF
C48638 PAND2X1_266/a_76_28# POR2X1_73/Y 0.01fF
C48639 POR2X1_254/A POR2X1_254/CTRL 0.01fF
C48640 POR2X1_800/A POR2X1_452/Y 0.12fF
C48641 POR2X1_65/A PAND2X1_564/B 0.03fF
C48642 PAND2X1_826/O PAND2X1_55/Y 0.02fF
C48643 POR2X1_23/Y PAND2X1_198/Y 0.06fF
C48644 POR2X1_590/A PAND2X1_90/Y 0.08fF
C48645 POR2X1_471/O POR2X1_66/A 0.02fF
C48646 POR2X1_311/Y PAND2X1_192/Y 0.03fF
C48647 POR2X1_341/A POR2X1_341/O 0.14fF
C48648 POR2X1_370/a_16_28# POR2X1_717/B 0.02fF
C48649 PAND2X1_416/O POR2X1_415/Y -0.00fF
C48650 PAND2X1_217/B POR2X1_272/CTRL2 -0.00fF
C48651 POR2X1_157/O POR2X1_12/A 0.06fF
C48652 PAND2X1_205/A POR2X1_46/Y 0.03fF
C48653 POR2X1_612/B POR2X1_293/Y 0.01fF
C48654 POR2X1_650/O PAND2X1_65/B 0.01fF
C48655 POR2X1_23/Y PAND2X1_775/CTRL2 0.15fF
C48656 POR2X1_254/CTRL POR2X1_750/B 0.01fF
C48657 POR2X1_492/CTRL2 PAND2X1_558/Y 0.03fF
C48658 PAND2X1_796/CTRL VDD 0.00fF
C48659 POR2X1_800/A POR2X1_808/CTRL2 0.00fF
C48660 PAND2X1_647/B VDD 0.03fF
C48661 POR2X1_66/B POR2X1_267/B 0.05fF
C48662 POR2X1_94/O POR2X1_24/Y 0.01fF
C48663 POR2X1_220/B POR2X1_190/Y 0.03fF
C48664 PAND2X1_436/A POR2X1_677/O -0.02fF
C48665 POR2X1_670/CTRL POR2X1_40/Y -0.00fF
C48666 POR2X1_837/B POR2X1_507/A 0.01fF
C48667 PAND2X1_562/B POR2X1_40/Y 0.07fF
C48668 PAND2X1_811/a_76_28# PAND2X1_811/A 0.04fF
C48669 POR2X1_814/B POR2X1_750/B 1.39fF
C48670 POR2X1_648/Y POR2X1_407/O 0.01fF
C48671 POR2X1_863/A POR2X1_188/Y 0.03fF
C48672 PAND2X1_271/CTRL POR2X1_804/A 0.05fF
C48673 POR2X1_852/B POR2X1_194/A 0.04fF
C48674 POR2X1_814/B POR2X1_461/CTRL 0.01fF
C48675 POR2X1_49/Y PAND2X1_576/a_16_344# 0.01fF
C48676 PAND2X1_272/CTRL2 POR2X1_193/A 0.03fF
C48677 INPUT_1 PAND2X1_608/CTRL 0.03fF
C48678 POR2X1_475/A PAND2X1_41/B 0.01fF
C48679 PAND2X1_695/CTRL2 PAND2X1_41/B 0.01fF
C48680 POR2X1_311/Y PAND2X1_738/Y 0.05fF
C48681 POR2X1_445/A PAND2X1_69/A 0.67fF
C48682 PAND2X1_279/O POR2X1_284/B 0.01fF
C48683 POR2X1_502/A POR2X1_602/A 0.01fF
C48684 POR2X1_294/Y PAND2X1_55/Y 0.01fF
C48685 POR2X1_393/Y VDD 0.00fF
C48686 POR2X1_52/A PAND2X1_623/O 0.02fF
C48687 POR2X1_775/A POR2X1_567/B 0.03fF
C48688 PAND2X1_6/Y PAND2X1_248/CTRL 0.01fF
C48689 POR2X1_174/B POR2X1_853/CTRL 0.28fF
C48690 POR2X1_272/CTRL2 VDD -0.00fF
C48691 PAND2X1_354/A PAND2X1_347/Y 0.03fF
C48692 PAND2X1_254/CTRL POR2X1_669/B 0.08fF
C48693 POR2X1_57/A PAND2X1_222/A 0.01fF
C48694 PAND2X1_409/O PAND2X1_11/Y 0.02fF
C48695 POR2X1_423/Y PAND2X1_140/Y 0.03fF
C48696 PAND2X1_90/A POR2X1_614/Y 0.02fF
C48697 POR2X1_102/Y PAND2X1_364/B 0.07fF
C48698 PAND2X1_472/A POR2X1_48/A 0.01fF
C48699 POR2X1_857/CTRL POR2X1_785/A 0.01fF
C48700 POR2X1_490/Y PAND2X1_341/A 0.03fF
C48701 POR2X1_302/Y POR2X1_302/B 0.39fF
C48702 PAND2X1_68/CTRL2 PAND2X1_6/A 0.02fF
C48703 POR2X1_49/Y POR2X1_406/Y 0.06fF
C48704 POR2X1_13/A POR2X1_40/Y 1.15fF
C48705 POR2X1_389/CTRL POR2X1_121/B 0.01fF
C48706 POR2X1_334/B PAND2X1_73/Y 0.10fF
C48707 POR2X1_362/Y PAND2X1_48/B 0.35fF
C48708 POR2X1_23/Y PAND2X1_243/CTRL2 0.01fF
C48709 PAND2X1_771/Y PAND2X1_577/O 0.33fF
C48710 POR2X1_471/A POR2X1_569/A 0.02fF
C48711 POR2X1_465/A POR2X1_186/Y 0.11fF
C48712 POR2X1_590/A POR2X1_732/CTRL2 0.01fF
C48713 POR2X1_750/B PAND2X1_176/CTRL2 0.01fF
C48714 PAND2X1_6/Y POR2X1_97/A 0.03fF
C48715 POR2X1_616/a_16_28# POR2X1_90/Y 0.01fF
C48716 POR2X1_609/Y POR2X1_232/Y 0.00fF
C48717 PAND2X1_214/B POR2X1_40/Y 0.05fF
C48718 POR2X1_81/a_16_28# POR2X1_293/Y 0.02fF
C48719 POR2X1_606/m4_208_n4# PAND2X1_32/B 0.15fF
C48720 POR2X1_801/B PAND2X1_583/CTRL 0.00fF
C48721 POR2X1_682/CTRL POR2X1_829/A 0.00fF
C48722 POR2X1_49/Y POR2X1_293/Y 0.10fF
C48723 POR2X1_403/B POR2X1_403/Y 0.03fF
C48724 PAND2X1_774/O PAND2X1_771/Y 0.03fF
C48725 POR2X1_271/A POR2X1_271/B 0.16fF
C48726 POR2X1_41/B POR2X1_376/B 0.21fF
C48727 POR2X1_529/O POR2X1_40/Y 0.01fF
C48728 POR2X1_564/Y PAND2X1_90/Y 0.03fF
C48729 PAND2X1_573/O PAND2X1_499/Y 0.05fF
C48730 PAND2X1_60/CTRL2 POR2X1_66/A 0.01fF
C48731 POR2X1_495/Y POR2X1_495/O 0.00fF
C48732 POR2X1_41/B PAND2X1_596/CTRL2 0.01fF
C48733 PAND2X1_822/O POR2X1_590/A -0.00fF
C48734 POR2X1_455/O POR2X1_76/Y -0.00fF
C48735 PAND2X1_58/A POR2X1_804/A 0.06fF
C48736 POR2X1_68/A POR2X1_794/B 0.07fF
C48737 PAND2X1_7/CTRL2 PAND2X1_52/Y 0.01fF
C48738 PAND2X1_790/Y PAND2X1_793/A 0.01fF
C48739 POR2X1_72/B PAND2X1_717/O 0.03fF
C48740 PAND2X1_659/CTRL PAND2X1_735/Y 0.08fF
C48741 PAND2X1_50/CTRL INPUT_5 0.11fF
C48742 POR2X1_614/A POR2X1_634/CTRL 0.05fF
C48743 PAND2X1_512/Y POR2X1_372/m4_208_n4# 0.01fF
C48744 POR2X1_748/A PAND2X1_6/A 0.10fF
C48745 PAND2X1_623/Y POR2X1_847/B 0.03fF
C48746 POR2X1_96/A PAND2X1_739/CTRL 0.01fF
C48747 POR2X1_23/Y PAND2X1_550/B 0.03fF
C48748 PAND2X1_23/Y POR2X1_61/Y 0.03fF
C48749 PAND2X1_48/B PAND2X1_65/Y 0.40fF
C48750 POR2X1_614/A PAND2X1_230/a_76_28# 0.01fF
C48751 POR2X1_13/A PAND2X1_659/B 0.03fF
C48752 PAND2X1_651/Y PAND2X1_512/CTRL 0.00fF
C48753 POR2X1_378/Y VDD 0.00fF
C48754 D_INPUT_3 POR2X1_414/O 0.01fF
C48755 POR2X1_260/Y PAND2X1_65/B 0.01fF
C48756 PAND2X1_696/a_16_344# POR2X1_814/A 0.04fF
C48757 PAND2X1_319/B POR2X1_83/B 0.07fF
C48758 POR2X1_37/Y PAND2X1_559/CTRL 0.28fF
C48759 PAND2X1_41/B POR2X1_218/A 0.00fF
C48760 POR2X1_829/CTRL2 POR2X1_761/Y 0.01fF
C48761 PAND2X1_830/Y VDD 0.23fF
C48762 PAND2X1_466/O PAND2X1_803/A 0.00fF
C48763 POR2X1_83/O POR2X1_23/Y 0.01fF
C48764 PAND2X1_630/a_76_28# POR2X1_748/A 0.03fF
C48765 POR2X1_7/B VDD 4.00fF
C48766 POR2X1_806/m4_208_n4# PAND2X1_69/A 0.09fF
C48767 PAND2X1_95/B PAND2X1_18/O 0.05fF
C48768 POR2X1_580/O POR2X1_578/Y 0.01fF
C48769 PAND2X1_661/B POR2X1_40/Y 0.03fF
C48770 PAND2X1_643/Y POR2X1_40/Y 0.03fF
C48771 POR2X1_66/B PAND2X1_638/m4_208_n4# 0.08fF
C48772 PAND2X1_652/A PAND2X1_787/Y 0.00fF
C48773 POR2X1_277/O VDD 0.00fF
C48774 POR2X1_334/B PAND2X1_262/a_76_28# 0.03fF
C48775 POR2X1_549/A POR2X1_549/B 0.29fF
C48776 POR2X1_197/O POR2X1_205/Y 0.01fF
C48777 POR2X1_488/Y PAND2X1_580/B 0.03fF
C48778 POR2X1_119/Y POR2X1_442/CTRL 0.01fF
C48779 POR2X1_465/B POR2X1_220/Y 0.03fF
C48780 POR2X1_334/Y POR2X1_454/A 0.03fF
C48781 POR2X1_596/Y POR2X1_294/B 0.00fF
C48782 POR2X1_290/Y POR2X1_233/CTRL 0.06fF
C48783 POR2X1_293/Y POR2X1_586/CTRL2 0.02fF
C48784 PAND2X1_467/Y POR2X1_32/A 0.03fF
C48785 POR2X1_750/CTRL POR2X1_750/A 0.01fF
C48786 POR2X1_78/A POR2X1_218/CTRL 0.01fF
C48787 POR2X1_502/A POR2X1_651/O 0.31fF
C48788 POR2X1_57/A PAND2X1_168/Y 0.00fF
C48789 POR2X1_78/B POR2X1_775/A 0.01fF
C48790 POR2X1_681/O POR2X1_39/B 0.05fF
C48791 PAND2X1_42/CTRL POR2X1_68/B 0.01fF
C48792 POR2X1_41/B POR2X1_52/A 0.16fF
C48793 PAND2X1_632/B POR2X1_669/B 0.03fF
C48794 POR2X1_254/CTRL2 POR2X1_228/Y 0.10fF
C48795 POR2X1_254/Y POR2X1_740/Y 0.10fF
C48796 POR2X1_287/CTRL POR2X1_249/Y 0.01fF
C48797 POR2X1_113/CTRL POR2X1_640/Y 0.01fF
C48798 PAND2X1_48/B PAND2X1_371/CTRL2 0.00fF
C48799 POR2X1_814/B PAND2X1_177/CTRL 0.01fF
C48800 POR2X1_359/B PAND2X1_93/B 0.03fF
C48801 POR2X1_566/A POR2X1_732/B 0.10fF
C48802 POR2X1_742/a_16_28# POR2X1_740/Y 0.08fF
C48803 POR2X1_121/B POR2X1_249/Y 0.06fF
C48804 POR2X1_96/Y PAND2X1_98/a_76_28# 0.04fF
C48805 POR2X1_525/Y POR2X1_763/Y 0.12fF
C48806 PAND2X1_69/A POR2X1_786/O 0.18fF
C48807 POR2X1_300/O POR2X1_46/Y 0.04fF
C48808 PAND2X1_58/CTRL PAND2X1_69/A 0.06fF
C48809 POR2X1_49/Y POR2X1_408/Y 0.15fF
C48810 POR2X1_290/Y POR2X1_42/Y 0.12fF
C48811 POR2X1_795/CTRL2 POR2X1_294/B 0.00fF
C48812 PAND2X1_684/CTRL POR2X1_78/A 0.01fF
C48813 POR2X1_220/Y D_GATE_741 0.07fF
C48814 PAND2X1_55/Y POR2X1_554/Y 0.03fF
C48815 PAND2X1_477/B VDD 0.17fF
C48816 PAND2X1_391/CTRL2 POR2X1_384/Y 0.03fF
C48817 POR2X1_780/a_16_28# POR2X1_780/A 0.02fF
C48818 POR2X1_96/A POR2X1_305/Y 0.03fF
C48819 POR2X1_40/Y POR2X1_321/Y 0.01fF
C48820 POR2X1_435/Y POR2X1_804/A 0.22fF
C48821 PAND2X1_456/O POR2X1_283/A 0.10fF
C48822 PAND2X1_354/A PAND2X1_346/Y 0.05fF
C48823 D_GATE_222 POR2X1_579/Y 0.07fF
C48824 POR2X1_411/B POR2X1_77/Y 1.47fF
C48825 POR2X1_650/A POR2X1_493/a_76_344# 0.02fF
C48826 POR2X1_353/Y POR2X1_353/O 0.02fF
C48827 POR2X1_134/Y POR2X1_13/A 0.00fF
C48828 PAND2X1_365/O POR2X1_7/B 0.04fF
C48829 POR2X1_572/O PAND2X1_32/B 0.01fF
C48830 PAND2X1_55/Y PAND2X1_29/CTRL2 0.09fF
C48831 POR2X1_43/B PAND2X1_859/B 0.01fF
C48832 POR2X1_376/Y PAND2X1_63/B 0.01fF
C48833 PAND2X1_200/Y POR2X1_394/A 0.01fF
C48834 PAND2X1_23/Y POR2X1_35/Y 0.08fF
C48835 PAND2X1_216/B PAND2X1_390/Y 0.20fF
C48836 PAND2X1_623/Y POR2X1_90/m4_208_n4# 0.01fF
C48837 PAND2X1_40/a_76_28# PAND2X1_57/B 0.03fF
C48838 POR2X1_483/A POR2X1_366/A 0.02fF
C48839 PAND2X1_798/B PAND2X1_575/A 0.51fF
C48840 PAND2X1_693/a_56_28# PAND2X1_48/B 0.00fF
C48841 VDD PAND2X1_60/B 2.59fF
C48842 POR2X1_305/Y PAND2X1_506/CTRL 0.01fF
C48843 PAND2X1_6/Y POR2X1_294/B 0.38fF
C48844 POR2X1_41/B PAND2X1_186/O 0.05fF
C48845 POR2X1_740/Y POR2X1_574/O 0.03fF
C48846 POR2X1_741/Y POR2X1_574/CTRL 0.00fF
C48847 POR2X1_7/B PAND2X1_32/B 0.02fF
C48848 POR2X1_150/Y POR2X1_173/O 0.01fF
C48849 PAND2X1_865/Y D_INPUT_0 0.03fF
C48850 PAND2X1_831/Y POR2X1_96/A 0.03fF
C48851 POR2X1_260/B POR2X1_39/B 0.03fF
C48852 PAND2X1_798/B PAND2X1_794/B 0.03fF
C48853 PAND2X1_787/Y PAND2X1_175/O 0.15fF
C48854 PAND2X1_57/B PAND2X1_757/O 0.02fF
C48855 PAND2X1_701/CTRL2 POR2X1_710/A 0.01fF
C48856 POR2X1_57/A POR2X1_56/B 0.02fF
C48857 POR2X1_471/A PAND2X1_72/A 0.06fF
C48858 PAND2X1_778/Y POR2X1_293/Y 0.03fF
C48859 POR2X1_614/A D_GATE_222 0.10fF
C48860 POR2X1_332/Y POR2X1_254/A 0.02fF
C48861 POR2X1_174/B PAND2X1_165/O 0.16fF
C48862 POR2X1_278/Y POR2X1_187/CTRL2 0.05fF
C48863 POR2X1_376/B PAND2X1_308/Y 0.19fF
C48864 VDD POR2X1_737/CTRL 0.00fF
C48865 POR2X1_60/A POR2X1_7/Y 0.03fF
C48866 PAND2X1_659/B PAND2X1_510/B 0.02fF
C48867 PAND2X1_94/A PAND2X1_293/CTRL2 0.01fF
C48868 PAND2X1_41/B POR2X1_557/B 0.03fF
C48869 POR2X1_335/a_16_28# POR2X1_538/A 0.03fF
C48870 POR2X1_788/Y PAND2X1_144/m4_208_n4# 0.02fF
C48871 POR2X1_270/Y POR2X1_736/A 0.08fF
C48872 POR2X1_130/Y POR2X1_140/CTRL -0.00fF
C48873 PAND2X1_810/CTRL GATE_741 0.01fF
C48874 PAND2X1_643/Y POR2X1_761/a_16_28# 0.01fF
C48875 PAND2X1_44/O PAND2X1_3/B 0.01fF
C48876 POR2X1_315/Y POR2X1_46/Y 0.03fF
C48877 POR2X1_258/CTRL PAND2X1_566/Y 0.03fF
C48878 PAND2X1_718/CTRL POR2X1_591/Y 0.01fF
C48879 POR2X1_532/A PAND2X1_146/O 0.01fF
C48880 POR2X1_334/O VDD 0.00fF
C48881 PAND2X1_23/Y POR2X1_325/CTRL2 0.01fF
C48882 PAND2X1_252/CTRL2 POR2X1_556/Y 0.00fF
C48883 VDD POR2X1_353/A 0.38fF
C48884 PAND2X1_79/Y PAND2X1_316/O 0.02fF
C48885 POR2X1_283/A PAND2X1_115/B 0.02fF
C48886 PAND2X1_713/O PAND2X1_725/B 0.00fF
C48887 PAND2X1_63/Y PAND2X1_69/A 0.03fF
C48888 PAND2X1_96/B POR2X1_804/A 0.03fF
C48889 POR2X1_257/A PAND2X1_242/Y 0.03fF
C48890 POR2X1_741/Y PAND2X1_60/B 0.03fF
C48891 POR2X1_495/Y PAND2X1_549/B 0.01fF
C48892 POR2X1_48/CTRL PAND2X1_123/Y 0.01fF
C48893 POR2X1_314/CTRL2 POR2X1_16/A 0.03fF
C48894 POR2X1_750/B PAND2X1_680/O 0.02fF
C48895 PAND2X1_81/B PAND2X1_60/B 0.68fF
C48896 PAND2X1_675/A PAND2X1_843/Y 0.07fF
C48897 POR2X1_286/CTRL PAND2X1_52/B 0.01fF
C48898 POR2X1_57/A PAND2X1_724/CTRL2 0.01fF
C48899 POR2X1_805/A POR2X1_713/B 0.03fF
C48900 PAND2X1_575/B POR2X1_184/CTRL2 0.01fF
C48901 PAND2X1_572/O POR2X1_52/Y 0.17fF
C48902 POR2X1_348/A POR2X1_99/B 0.27fF
C48903 PAND2X1_495/O PAND2X1_69/A 0.16fF
C48904 POR2X1_730/Y POR2X1_356/A 0.05fF
C48905 PAND2X1_6/Y PAND2X1_111/B 1.52fF
C48906 POR2X1_198/B POR2X1_215/A 0.48fF
C48907 POR2X1_305/Y POR2X1_7/A 0.46fF
C48908 POR2X1_192/Y POR2X1_566/CTRL2 0.01fF
C48909 POR2X1_596/A POR2X1_532/A 0.04fF
C48910 POR2X1_549/a_16_28# POR2X1_266/A 0.03fF
C48911 POR2X1_97/A PAND2X1_52/B 0.09fF
C48912 POR2X1_566/A PAND2X1_313/a_76_28# 0.05fF
C48913 POR2X1_52/A PAND2X1_308/Y 0.02fF
C48914 POR2X1_270/a_16_28# PAND2X1_69/A 0.03fF
C48915 POR2X1_276/a_16_28# POR2X1_366/A 0.02fF
C48916 POR2X1_701/CTRL POR2X1_236/Y 0.00fF
C48917 PAND2X1_60/B PAND2X1_32/B 0.24fF
C48918 PAND2X1_95/B PAND2X1_51/CTRL 0.01fF
C48919 POR2X1_383/A POR2X1_865/CTRL2 0.01fF
C48920 PAND2X1_659/Y POR2X1_822/O 0.01fF
C48921 POR2X1_802/CTRL2 POR2X1_532/A 0.01fF
C48922 PAND2X1_691/Y PAND2X1_664/CTRL 0.10fF
C48923 POR2X1_316/CTRL POR2X1_293/Y 0.03fF
C48924 PAND2X1_23/Y PAND2X1_701/CTRL 0.13fF
C48925 PAND2X1_94/A PAND2X1_411/O 0.15fF
C48926 POR2X1_360/A POR2X1_334/Y 0.20fF
C48927 POR2X1_283/A POR2X1_73/Y 0.06fF
C48928 PAND2X1_308/Y POR2X1_152/A 4.64fF
C48929 POR2X1_87/m4_208_n4# POR2X1_590/A 0.12fF
C48930 INPUT_0 PAND2X1_851/O 0.03fF
C48931 POR2X1_685/A PAND2X1_69/A 0.01fF
C48932 POR2X1_519/a_16_28# POR2X1_42/Y 0.01fF
C48933 POR2X1_667/A PAND2X1_327/a_16_344# 0.02fF
C48934 POR2X1_740/Y POR2X1_731/A 0.02fF
C48935 POR2X1_40/Y POR2X1_524/m4_208_n4# 0.09fF
C48936 POR2X1_566/A POR2X1_97/B 0.03fF
C48937 PAND2X1_803/Y POR2X1_387/Y 0.03fF
C48938 PAND2X1_23/Y POR2X1_227/CTRL2 0.06fF
C48939 POR2X1_383/A POR2X1_361/CTRL2 0.01fF
C48940 PAND2X1_386/O D_INPUT_4 0.01fF
C48941 POR2X1_76/B POR2X1_274/O 0.16fF
C48942 POR2X1_71/Y PAND2X1_657/B 0.01fF
C48943 POR2X1_390/B PAND2X1_311/CTRL2 0.00fF
C48944 PAND2X1_787/CTRL2 POR2X1_77/Y 0.01fF
C48945 INPUT_1 PAND2X1_401/a_76_28# 0.02fF
C48946 PAND2X1_803/A POR2X1_39/B 0.03fF
C48947 PAND2X1_94/A POR2X1_68/B 0.97fF
C48948 PAND2X1_69/A POR2X1_260/A 10.78fF
C48949 POR2X1_273/Y POR2X1_153/Y 0.03fF
C48950 POR2X1_294/B POR2X1_195/O 0.01fF
C48951 PAND2X1_661/Y PAND2X1_194/O 0.04fF
C48952 POR2X1_76/B POR2X1_296/B 1.94fF
C48953 PAND2X1_95/B PAND2X1_18/B 0.32fF
C48954 POR2X1_376/B POR2X1_77/Y 5.64fF
C48955 PAND2X1_90/A PAND2X1_90/O 0.03fF
C48956 POR2X1_394/A POR2X1_90/Y 0.17fF
C48957 POR2X1_8/Y POR2X1_382/Y 0.02fF
C48958 POR2X1_145/CTRL2 PAND2X1_797/Y 0.01fF
C48959 POR2X1_383/A POR2X1_249/Y 0.10fF
C48960 PAND2X1_673/Y POR2X1_39/B 0.09fF
C48961 POR2X1_252/Y PAND2X1_658/B 0.05fF
C48962 POR2X1_137/Y POR2X1_216/Y 0.00fF
C48963 POR2X1_66/B POR2X1_814/CTRL 0.01fF
C48964 PAND2X1_9/Y PAND2X1_407/CTRL2 0.01fF
C48965 POR2X1_168/m4_208_n4# POR2X1_578/Y 0.07fF
C48966 POR2X1_317/CTRL2 POR2X1_169/A 0.01fF
C48967 PAND2X1_653/Y PAND2X1_659/Y 6.64fF
C48968 POR2X1_687/O POR2X1_814/A 0.35fF
C48969 PAND2X1_6/Y POR2X1_567/A 0.32fF
C48970 PAND2X1_65/B POR2X1_535/CTRL2 0.01fF
C48971 PAND2X1_6/Y PAND2X1_323/O 0.07fF
C48972 PAND2X1_53/O POR2X1_66/A 0.03fF
C48973 POR2X1_52/A POR2X1_77/Y 0.13fF
C48974 PAND2X1_575/A POR2X1_184/O 0.08fF
C48975 POR2X1_294/B POR2X1_632/Y 0.03fF
C48976 POR2X1_119/Y PAND2X1_785/A 0.01fF
C48977 POR2X1_316/Y POR2X1_43/B 0.01fF
C48978 PAND2X1_6/Y POR2X1_542/O 0.01fF
C48979 POR2X1_54/Y PAND2X1_35/A 0.03fF
C48980 POR2X1_673/Y POR2X1_546/O 0.02fF
C48981 POR2X1_458/Y POR2X1_457/O 0.05fF
C48982 POR2X1_329/A PAND2X1_573/B 0.10fF
C48983 PAND2X1_824/B POR2X1_260/A 0.10fF
C48984 POR2X1_677/O POR2X1_677/Y 0.02fF
C48985 POR2X1_51/CTRL2 INPUT_6 0.03fF
C48986 PAND2X1_63/CTRL2 PAND2X1_9/Y 0.00fF
C48987 PAND2X1_508/Y PAND2X1_861/CTRL2 0.01fF
C48988 POR2X1_113/A POR2X1_260/A 0.00fF
C48989 POR2X1_366/Y PAND2X1_52/B 0.07fF
C48990 POR2X1_294/B PAND2X1_52/B 0.34fF
C48991 PAND2X1_856/B PAND2X1_856/a_76_28# 0.03fF
C48992 POR2X1_65/CTRL POR2X1_60/A 0.06fF
C48993 POR2X1_675/Y POR2X1_186/B 0.06fF
C48994 PAND2X1_308/Y PAND2X1_727/a_56_28# 0.00fF
C48995 POR2X1_817/CTRL2 PAND2X1_340/B 0.01fF
C48996 POR2X1_357/B POR2X1_854/B 0.32fF
C48997 PAND2X1_289/CTRL POR2X1_220/B 0.01fF
C48998 PAND2X1_488/CTRL2 POR2X1_814/A 0.01fF
C48999 PAND2X1_797/Y PAND2X1_731/A 0.03fF
C49000 POR2X1_458/Y POR2X1_543/A 0.01fF
C49001 POR2X1_518/a_16_28# POR2X1_73/Y 0.12fF
C49002 POR2X1_510/Y POR2X1_554/CTRL2 0.00fF
C49003 PAND2X1_56/Y POR2X1_715/CTRL 0.01fF
C49004 POR2X1_78/A POR2X1_649/O 0.01fF
C49005 POR2X1_544/B POR2X1_186/B 0.03fF
C49006 POR2X1_8/Y POR2X1_749/a_16_28# -0.00fF
C49007 POR2X1_55/Y PAND2X1_349/O 0.02fF
C49008 POR2X1_48/A POR2X1_260/B 0.03fF
C49009 POR2X1_90/Y PAND2X1_326/CTRL 0.03fF
C49010 POR2X1_67/Y PAND2X1_526/O 0.02fF
C49011 POR2X1_174/B POR2X1_776/A 10.87fF
C49012 POR2X1_416/B POR2X1_591/Y 0.07fF
C49013 POR2X1_110/Y POR2X1_394/A 0.03fF
C49014 PAND2X1_484/a_76_28# POR2X1_559/A 0.10fF
C49015 POR2X1_257/A POR2X1_60/A 14.58fF
C49016 POR2X1_456/B PAND2X1_167/O 0.01fF
C49017 POR2X1_571/a_16_28# POR2X1_561/Y -0.00fF
C49018 POR2X1_48/A POR2X1_482/CTRL 0.01fF
C49019 POR2X1_23/Y POR2X1_482/O 0.03fF
C49020 POR2X1_20/B PAND2X1_541/CTRL 0.02fF
C49021 POR2X1_376/B PAND2X1_449/O 0.06fF
C49022 PAND2X1_206/B VDD 0.06fF
C49023 D_INPUT_0 POR2X1_66/A 0.06fF
C49024 POR2X1_334/Y POR2X1_99/B 0.04fF
C49025 PAND2X1_294/CTRL POR2X1_40/Y 0.01fF
C49026 PAND2X1_798/B PAND2X1_221/Y 0.03fF
C49027 POR2X1_150/Y PAND2X1_736/CTRL2 0.01fF
C49028 POR2X1_458/Y PAND2X1_369/CTRL2 0.02fF
C49029 POR2X1_210/Y POR2X1_161/a_16_28# 0.02fF
C49030 PAND2X1_211/O POR2X1_40/Y 0.05fF
C49031 PAND2X1_809/CTRL POR2X1_7/B 0.09fF
C49032 POR2X1_41/B POR2X1_441/O 0.02fF
C49033 PAND2X1_251/a_16_344# POR2X1_296/B 0.06fF
C49034 POR2X1_90/Y POR2X1_91/CTRL 0.00fF
C49035 PAND2X1_631/A PAND2X1_508/Y 0.02fF
C49036 PAND2X1_93/B PAND2X1_394/CTRL 0.01fF
C49037 POR2X1_610/a_16_28# POR2X1_590/A 0.02fF
C49038 POR2X1_681/CTRL2 POR2X1_829/A 0.00fF
C49039 POR2X1_68/O POR2X1_296/B 0.18fF
C49040 POR2X1_503/O POR2X1_77/Y 0.01fF
C49041 POR2X1_477/CTRL VDD 0.00fF
C49042 POR2X1_260/Y POR2X1_814/A 0.05fF
C49043 POR2X1_566/B POR2X1_568/A 0.03fF
C49044 PAND2X1_93/B POR2X1_330/Y 0.12fF
C49045 PAND2X1_206/B PAND2X1_101/CTRL2 0.01fF
C49046 POR2X1_808/A POR2X1_808/a_16_28# 0.04fF
C49047 POR2X1_411/B PAND2X1_571/Y 0.03fF
C49048 POR2X1_16/O POR2X1_591/Y 0.02fF
C49049 POR2X1_632/CTRL2 POR2X1_61/Y 0.02fF
C49050 POR2X1_278/Y POR2X1_150/Y 0.07fF
C49051 POR2X1_730/Y PAND2X1_72/A 0.40fF
C49052 PAND2X1_55/Y PAND2X1_45/CTRL2 0.01fF
C49053 POR2X1_227/B POR2X1_244/B 0.08fF
C49054 PAND2X1_56/Y POR2X1_260/CTRL 0.01fF
C49055 POR2X1_38/CTRL2 POR2X1_5/Y 0.03fF
C49056 POR2X1_23/Y PAND2X1_579/CTRL2 0.03fF
C49057 POR2X1_788/A POR2X1_296/B 0.02fF
C49058 POR2X1_65/Y VDD 0.01fF
C49059 POR2X1_866/O POR2X1_801/B 0.01fF
C49060 PAND2X1_571/a_76_28# PAND2X1_561/Y 0.04fF
C49061 POR2X1_479/B POR2X1_479/a_16_28# 0.02fF
C49062 POR2X1_846/A POR2X1_789/CTRL2 0.00fF
C49063 PAND2X1_673/O POR2X1_672/Y 0.13fF
C49064 POR2X1_302/Y POR2X1_831/a_56_344# 0.01fF
C49065 POR2X1_466/O POR2X1_453/Y 0.00fF
C49066 PAND2X1_475/CTRL2 POR2X1_102/Y 0.01fF
C49067 POR2X1_20/B POR2X1_628/CTRL2 0.03fF
C49068 POR2X1_378/Y PAND2X1_9/Y 0.04fF
C49069 POR2X1_479/B POR2X1_734/A 0.02fF
C49070 PAND2X1_258/O PAND2X1_52/Y 0.01fF
C49071 PAND2X1_97/O POR2X1_5/Y 0.15fF
C49072 POR2X1_29/A POR2X1_40/Y 0.05fF
C49073 POR2X1_638/Y PAND2X1_53/CTRL2 0.06fF
C49074 POR2X1_698/CTRL POR2X1_32/A 0.01fF
C49075 D_INPUT_7 INPUT_6 0.25fF
C49076 PAND2X1_9/Y POR2X1_7/B 0.03fF
C49077 POR2X1_88/O VDD 0.00fF
C49078 POR2X1_49/Y PAND2X1_61/O 0.17fF
C49079 PAND2X1_292/a_16_344# POR2X1_186/B 0.02fF
C49080 PAND2X1_657/CTRL2 POR2X1_72/B 0.00fF
C49081 POR2X1_78/A POR2X1_330/Y 0.05fF
C49082 PAND2X1_458/CTRL2 POR2X1_283/A 0.02fF
C49083 PAND2X1_62/CTRL D_INPUT_0 0.01fF
C49084 POR2X1_843/CTRL POR2X1_343/A 0.01fF
C49085 PAND2X1_58/A POR2X1_794/B 3.01fF
C49086 PAND2X1_45/m4_208_n4# POR2X1_741/Y 0.12fF
C49087 POR2X1_175/A POR2X1_78/A 0.07fF
C49088 POR2X1_260/B POR2X1_459/CTRL 0.00fF
C49089 POR2X1_66/A PAND2X1_90/Y 0.21fF
C49090 POR2X1_643/Y POR2X1_121/Y 0.11fF
C49091 PAND2X1_79/O POR2X1_78/Y 0.01fF
C49092 PAND2X1_240/CTRL2 POR2X1_102/Y 0.01fF
C49093 PAND2X1_23/Y POR2X1_294/CTRL2 0.01fF
C49094 POR2X1_329/A POR2X1_91/Y 0.07fF
C49095 POR2X1_114/CTRL POR2X1_499/A 0.00fF
C49096 POR2X1_660/Y POR2X1_830/A 0.03fF
C49097 POR2X1_188/A PAND2X1_701/m4_208_n4# 0.07fF
C49098 POR2X1_49/Y POR2X1_60/A 0.13fF
C49099 POR2X1_376/Y POR2X1_32/A 0.02fF
C49100 POR2X1_383/A POR2X1_655/m4_208_n4# 0.09fF
C49101 POR2X1_428/Y PAND2X1_709/CTRL 0.01fF
C49102 PAND2X1_237/O POR2X1_192/Y 0.03fF
C49103 PAND2X1_65/B PAND2X1_245/CTRL 0.01fF
C49104 POR2X1_427/O POR2X1_236/Y 0.18fF
C49105 PAND2X1_849/B POR2X1_9/Y 0.07fF
C49106 POR2X1_23/Y PAND2X1_734/B 0.02fF
C49107 POR2X1_76/CTRL POR2X1_740/Y 0.19fF
C49108 POR2X1_200/CTRL2 PAND2X1_41/B 0.03fF
C49109 POR2X1_341/A PAND2X1_316/CTRL 0.01fF
C49110 PAND2X1_550/CTRL POR2X1_32/A 0.01fF
C49111 POR2X1_383/A POR2X1_260/CTRL 0.07fF
C49112 POR2X1_116/A POR2X1_112/Y 0.01fF
C49113 PAND2X1_307/a_16_344# POR2X1_40/Y 0.00fF
C49114 POR2X1_833/A PAND2X1_255/CTRL2 0.05fF
C49115 POR2X1_54/Y POR2X1_43/B 0.40fF
C49116 POR2X1_566/A POR2X1_466/A 0.10fF
C49117 POR2X1_840/B POR2X1_556/A 0.05fF
C49118 POR2X1_508/B POR2X1_568/A 0.03fF
C49119 POR2X1_54/Y POR2X1_789/A 0.03fF
C49120 POR2X1_66/B PAND2X1_815/CTRL 0.02fF
C49121 PAND2X1_556/B POR2X1_32/A 1.20fF
C49122 PAND2X1_235/CTRL PAND2X1_85/Y 0.01fF
C49123 POR2X1_29/Y INPUT_3 1.27fF
C49124 PAND2X1_673/O POR2X1_83/B 0.17fF
C49125 POR2X1_41/B POR2X1_484/CTRL2 0.01fF
C49126 POR2X1_812/A POR2X1_801/A 0.05fF
C49127 PAND2X1_250/O POR2X1_389/Y 0.01fF
C49128 POR2X1_632/CTRL2 POR2X1_35/Y 0.01fF
C49129 POR2X1_750/B PAND2X1_526/CTRL 0.00fF
C49130 PAND2X1_278/O PAND2X1_41/B 0.02fF
C49131 POR2X1_435/O POR2X1_435/B 0.00fF
C49132 PAND2X1_630/B PAND2X1_507/O 0.02fF
C49133 POR2X1_610/Y PAND2X1_69/A 0.03fF
C49134 PAND2X1_30/CTRL2 PAND2X1_3/B 0.01fF
C49135 POR2X1_814/B POR2X1_389/Y 0.13fF
C49136 POR2X1_65/A PAND2X1_859/A 0.03fF
C49137 POR2X1_439/Y POR2X1_186/Y 0.07fF
C49138 POR2X1_263/Y PAND2X1_215/B 0.00fF
C49139 POR2X1_65/A PAND2X1_211/A 0.03fF
C49140 PAND2X1_77/a_16_344# PAND2X1_8/Y 0.02fF
C49141 POR2X1_66/B POR2X1_78/B 0.47fF
C49142 POR2X1_666/a_16_28# INPUT_0 0.01fF
C49143 POR2X1_697/Y POR2X1_427/CTRL2 0.01fF
C49144 POR2X1_697/CTRL2 POR2X1_72/B 0.01fF
C49145 POR2X1_54/Y POR2X1_38/B 0.10fF
C49146 PAND2X1_733/A PAND2X1_723/Y 0.00fF
C49147 PAND2X1_471/O POR2X1_83/B 0.02fF
C49148 POR2X1_812/A POR2X1_809/B 0.01fF
C49149 POR2X1_102/Y POR2X1_411/CTRL2 0.00fF
C49150 PAND2X1_9/Y PAND2X1_60/B 0.12fF
C49151 PAND2X1_39/B POR2X1_318/A 0.07fF
C49152 POR2X1_78/B PAND2X1_420/m4_208_n4# 0.03fF
C49153 POR2X1_188/A POR2X1_78/B 0.03fF
C49154 POR2X1_96/A PAND2X1_221/CTRL2 0.01fF
C49155 PAND2X1_71/O POR2X1_296/B 0.06fF
C49156 POR2X1_832/O POR2X1_330/Y 0.04fF
C49157 POR2X1_417/Y PAND2X1_556/B 0.03fF
C49158 PAND2X1_56/Y POR2X1_842/a_56_344# 0.03fF
C49159 POR2X1_783/A POR2X1_783/CTRL2 0.01fF
C49160 POR2X1_750/B VDD 5.12fF
C49161 POR2X1_435/Y POR2X1_794/B 0.01fF
C49162 POR2X1_821/O POR2X1_40/Y 0.05fF
C49163 POR2X1_333/A POR2X1_776/B 0.05fF
C49164 POR2X1_60/A PAND2X1_553/B 0.08fF
C49165 POR2X1_220/O POR2X1_220/A 0.03fF
C49166 POR2X1_558/B D_INPUT_1 0.03fF
C49167 POR2X1_446/B POR2X1_714/O 0.01fF
C49168 POR2X1_502/A POR2X1_264/O 0.06fF
C49169 POR2X1_503/CTRL2 POR2X1_411/B 0.01fF
C49170 POR2X1_366/O POR2X1_556/A 0.01fF
C49171 POR2X1_517/Y POR2X1_667/A 0.07fF
C49172 POR2X1_96/A PAND2X1_772/a_76_28# 0.02fF
C49173 PAND2X1_220/Y VDD 2.14fF
C49174 POR2X1_516/A POR2X1_257/A 0.63fF
C49175 PAND2X1_254/Y POR2X1_417/Y 0.09fF
C49176 POR2X1_32/A POR2X1_599/A 0.03fF
C49177 PAND2X1_502/a_16_344# POR2X1_42/Y 0.06fF
C49178 POR2X1_192/Y POR2X1_186/Y 1.71fF
C49179 PAND2X1_65/O PAND2X1_69/A 0.02fF
C49180 POR2X1_590/A D_GATE_222 0.03fF
C49181 PAND2X1_37/CTRL2 PAND2X1_6/A 0.01fF
C49182 PAND2X1_785/a_16_344# PAND2X1_776/Y 0.03fF
C49183 PAND2X1_558/Y POR2X1_46/Y 0.02fF
C49184 POR2X1_467/Y POR2X1_294/B 0.07fF
C49185 PAND2X1_717/A PAND2X1_716/B 0.06fF
C49186 PAND2X1_20/A POR2X1_713/CTRL2 0.01fF
C49187 POR2X1_65/A POR2X1_96/A 5.44fF
C49188 PAND2X1_65/B PAND2X1_587/Y 0.03fF
C49189 POR2X1_353/Y POR2X1_566/A 0.03fF
C49190 D_INPUT_0 POR2X1_532/A 3.20fF
C49191 POR2X1_669/B POR2X1_90/Y 0.21fF
C49192 POR2X1_811/A POR2X1_532/A 0.00fF
C49193 PAND2X1_496/m4_208_n4# PAND2X1_48/A 0.08fF
C49194 POR2X1_13/A POR2X1_5/Y 0.76fF
C49195 POR2X1_66/B PAND2X1_7/O 0.04fF
C49196 POR2X1_52/A POR2X1_290/O 0.02fF
C49197 POR2X1_66/B POR2X1_460/O 0.02fF
C49198 PAND2X1_204/CTRL2 POR2X1_79/Y 0.01fF
C49199 POR2X1_509/A POR2X1_227/m4_208_n4# 0.17fF
C49200 PAND2X1_90/A PAND2X1_42/CTRL 0.03fF
C49201 POR2X1_40/Y PAND2X1_506/O 0.03fF
C49202 PAND2X1_645/O VDD 0.00fF
C49203 POR2X1_362/B POR2X1_723/a_16_28# 0.02fF
C49204 POR2X1_814/B POR2X1_756/CTRL2 0.01fF
C49205 POR2X1_20/B POR2X1_129/Y 0.14fF
C49206 PAND2X1_474/O POR2X1_153/Y 0.20fF
C49207 POR2X1_806/CTRL2 POR2X1_804/A 0.13fF
C49208 PAND2X1_739/Y VDD 0.04fF
C49209 PAND2X1_347/Y PAND2X1_568/CTRL 0.03fF
C49210 POR2X1_16/A PAND2X1_443/CTRL 0.01fF
C49211 PAND2X1_41/B POR2X1_740/Y 0.06fF
C49212 POR2X1_750/B POR2X1_741/Y 0.03fF
C49213 PAND2X1_279/CTRL2 PAND2X1_32/B 0.01fF
C49214 PAND2X1_469/B PAND2X1_556/a_76_28# 0.04fF
C49215 POR2X1_797/A POR2X1_149/Y 0.02fF
C49216 POR2X1_333/A POR2X1_577/CTRL2 0.05fF
C49217 POR2X1_150/Y PAND2X1_357/O 0.13fF
C49218 POR2X1_97/A POR2X1_350/B 0.02fF
C49219 PAND2X1_456/O POR2X1_55/Y 0.15fF
C49220 POR2X1_122/A POR2X1_293/Y 0.03fF
C49221 POR2X1_66/B PAND2X1_767/CTRL 0.01fF
C49222 PAND2X1_90/Y POR2X1_792/B 0.07fF
C49223 PAND2X1_90/Y POR2X1_802/B 0.10fF
C49224 POR2X1_41/CTRL2 PAND2X1_852/A 0.01fF
C49225 PAND2X1_55/Y POR2X1_402/CTRL 0.01fF
C49226 POR2X1_500/A PAND2X1_316/CTRL 0.00fF
C49227 POR2X1_615/a_16_28# POR2X1_754/A 0.05fF
C49228 POR2X1_14/Y POR2X1_73/Y 0.06fF
C49229 POR2X1_57/O POR2X1_5/Y 0.02fF
C49230 PAND2X1_576/CTRL2 POR2X1_599/A 0.29fF
C49231 PAND2X1_412/CTRL POR2X1_391/Y 0.01fF
C49232 POR2X1_48/a_16_28# POR2X1_46/Y 0.05fF
C49233 POR2X1_52/A PAND2X1_571/Y 0.02fF
C49234 PAND2X1_659/Y POR2X1_20/B 0.03fF
C49235 POR2X1_529/O POR2X1_5/Y 0.22fF
C49236 POR2X1_308/CTRL PAND2X1_55/Y 0.01fF
C49237 PAND2X1_480/B POR2X1_46/Y 0.07fF
C49238 PAND2X1_20/A POR2X1_318/A 0.17fF
C49239 POR2X1_753/Y POR2X1_283/A 0.07fF
C49240 POR2X1_750/B PAND2X1_32/B 3.30fF
C49241 POR2X1_267/A PAND2X1_60/B 0.03fF
C49242 POR2X1_278/Y PAND2X1_364/B 0.10fF
C49243 POR2X1_48/A POR2X1_394/CTRL 0.01fF
C49244 PAND2X1_839/CTRL2 VDD -0.00fF
C49245 PAND2X1_118/O PAND2X1_65/B 0.03fF
C49246 PAND2X1_6/Y POR2X1_807/A 0.03fF
C49247 PAND2X1_793/Y PAND2X1_468/CTRL 0.01fF
C49248 PAND2X1_329/O POR2X1_149/A 0.00fF
C49249 POR2X1_441/Y POR2X1_373/a_76_344# 0.00fF
C49250 POR2X1_235/a_16_28# POR2X1_32/A 0.03fF
C49251 POR2X1_201/a_76_344# PAND2X1_88/Y 0.00fF
C49252 PAND2X1_20/A POR2X1_713/B 0.75fF
C49253 PAND2X1_278/CTRL POR2X1_68/B 0.01fF
C49254 PAND2X1_217/B PAND2X1_575/CTRL 0.01fF
C49255 PAND2X1_41/B POR2X1_711/CTRL2 0.10fF
C49256 POR2X1_865/B POR2X1_777/B 3.71fF
C49257 POR2X1_78/B POR2X1_659/O 0.06fF
C49258 POR2X1_119/Y PAND2X1_203/a_16_344# 0.04fF
C49259 POR2X1_481/Y VDD 0.03fF
C49260 PAND2X1_459/Y POR2X1_55/Y 0.01fF
C49261 POR2X1_718/A PAND2X1_69/A 0.06fF
C49262 PAND2X1_632/O POR2X1_496/Y 0.09fF
C49263 PAND2X1_13/O PAND2X1_32/B 0.01fF
C49264 PAND2X1_213/Y POR2X1_72/B 0.03fF
C49265 POR2X1_43/B PAND2X1_501/B 0.85fF
C49266 POR2X1_355/B POR2X1_785/A 0.03fF
C49267 POR2X1_750/B PAND2X1_312/O 0.09fF
C49268 POR2X1_113/Y POR2X1_640/Y 0.01fF
C49269 POR2X1_808/A PAND2X1_60/B 0.02fF
C49270 PAND2X1_3/O PAND2X1_11/Y 0.02fF
C49271 PAND2X1_623/Y POR2X1_754/A 0.02fF
C49272 POR2X1_853/A POR2X1_570/CTRL 0.01fF
C49273 POR2X1_362/B POR2X1_501/B 0.05fF
C49274 POR2X1_669/B PAND2X1_732/A 0.07fF
C49275 PAND2X1_798/B PAND2X1_795/B 0.03fF
C49276 POR2X1_66/B POR2X1_141/A 0.01fF
C49277 POR2X1_502/A PAND2X1_144/O 0.06fF
C49278 POR2X1_814/B POR2X1_318/A 0.10fF
C49279 PAND2X1_841/CTRL PAND2X1_841/B 0.02fF
C49280 POR2X1_532/A PAND2X1_90/Y 0.63fF
C49281 PAND2X1_35/A POR2X1_4/Y 0.03fF
C49282 POR2X1_102/a_16_28# POR2X1_411/B 0.01fF
C49283 POR2X1_542/B POR2X1_663/O 0.05fF
C49284 PAND2X1_35/Y POR2X1_599/A 0.05fF
C49285 POR2X1_848/m4_208_n4# PAND2X1_52/B 0.12fF
C49286 POR2X1_358/a_76_344# POR2X1_578/Y 0.01fF
C49287 POR2X1_96/A PAND2X1_190/Y 0.54fF
C49288 POR2X1_113/CTRL2 PAND2X1_65/B 0.01fF
C49289 PAND2X1_95/B POR2X1_638/O 0.02fF
C49290 POR2X1_376/B PAND2X1_241/Y 0.03fF
C49291 POR2X1_763/Y PAND2X1_726/CTRL2 0.01fF
C49292 PAND2X1_691/Y POR2X1_829/O 0.04fF
C49293 PAND2X1_620/Y POR2X1_7/A 0.03fF
C49294 POR2X1_814/B POR2X1_713/B 0.06fF
C49295 PAND2X1_93/B POR2X1_337/Y 0.07fF
C49296 PAND2X1_202/CTRL2 D_INPUT_1 0.05fF
C49297 PAND2X1_824/B POR2X1_243/A 0.04fF
C49298 PAND2X1_254/Y POR2X1_184/Y 0.17fF
C49299 POR2X1_306/O POR2X1_236/Y 0.01fF
C49300 POR2X1_65/A POR2X1_7/A 1.31fF
C49301 POR2X1_662/Y PAND2X1_55/Y 0.04fF
C49302 POR2X1_143/a_56_344# POR2X1_43/B 0.00fF
C49303 POR2X1_356/A POR2X1_68/A 0.09fF
C49304 PAND2X1_658/A POR2X1_55/Y 1.21fF
C49305 POR2X1_259/A POR2X1_259/O 0.01fF
C49306 POR2X1_325/A POR2X1_318/A 0.07fF
C49307 PAND2X1_651/Y PAND2X1_254/Y 0.03fF
C49308 PAND2X1_824/B POR2X1_631/CTRL2 0.06fF
C49309 PAND2X1_474/A POR2X1_171/CTRL 0.01fF
C49310 POR2X1_411/Y POR2X1_416/Y 0.01fF
C49311 POR2X1_846/a_16_28# POR2X1_846/A 0.02fF
C49312 POR2X1_290/Y PAND2X1_642/B 0.23fF
C49313 PAND2X1_215/B PAND2X1_6/A 0.03fF
C49314 POR2X1_61/A POR2X1_66/A 0.01fF
C49315 PAND2X1_341/B D_INPUT_0 0.07fF
C49316 POR2X1_20/B PAND2X1_333/Y 0.00fF
C49317 PAND2X1_20/A POR2X1_574/Y 0.01fF
C49318 POR2X1_640/Y POR2X1_260/A 0.03fF
C49319 POR2X1_775/O POR2X1_776/B 0.00fF
C49320 POR2X1_132/Y POR2X1_96/A 0.00fF
C49321 POR2X1_13/A POR2X1_299/O 0.01fF
C49322 POR2X1_824/Y VDD 0.00fF
C49323 PAND2X1_649/A PAND2X1_590/O 0.02fF
C49324 PAND2X1_94/A PAND2X1_46/a_76_28# 0.01fF
C49325 POR2X1_780/a_16_28# POR2X1_796/A 0.00fF
C49326 PAND2X1_710/O POR2X1_763/A 0.04fF
C49327 PAND2X1_553/B PAND2X1_702/CTRL2 0.01fF
C49328 PAND2X1_854/A PAND2X1_366/Y 0.02fF
C49329 POR2X1_628/O PAND2X1_6/A 0.04fF
C49330 POR2X1_178/Y PAND2X1_562/B 0.01fF
C49331 POR2X1_346/B PAND2X1_16/O 0.03fF
C49332 POR2X1_5/Y PAND2X1_510/B 0.03fF
C49333 POR2X1_110/Y POR2X1_669/B 0.14fF
C49334 POR2X1_170/B POR2X1_577/O 0.01fF
C49335 POR2X1_433/a_16_28# POR2X1_153/Y -0.00fF
C49336 PAND2X1_804/A POR2X1_283/A 0.00fF
C49337 POR2X1_364/A POR2X1_319/O 0.02fF
C49338 PAND2X1_329/O VDD 0.00fF
C49339 POR2X1_830/A POR2X1_308/B 0.04fF
C49340 POR2X1_78/A POR2X1_337/Y 0.07fF
C49341 POR2X1_76/Y POR2X1_228/Y 0.03fF
C49342 POR2X1_502/A PAND2X1_306/a_16_344# 0.02fF
C49343 POR2X1_55/Y POR2X1_73/Y 0.12fF
C49344 POR2X1_408/m4_208_n4# POR2X1_587/Y 0.01fF
C49345 PAND2X1_713/A VDD 0.00fF
C49346 PAND2X1_94/A PAND2X1_80/CTRL2 0.01fF
C49347 POR2X1_66/B POR2X1_735/CTRL 0.01fF
C49348 POR2X1_52/A PAND2X1_241/Y 0.04fF
C49349 POR2X1_46/Y PAND2X1_303/B 0.00fF
C49350 POR2X1_333/A POR2X1_192/B 0.16fF
C49351 PAND2X1_852/CTRL2 POR2X1_821/Y 0.01fF
C49352 PAND2X1_488/a_76_28# POR2X1_260/A 0.02fF
C49353 POR2X1_765/CTRL2 POR2X1_73/Y 0.05fF
C49354 PAND2X1_785/Y POR2X1_283/A 0.02fF
C49355 POR2X1_38/B POR2X1_382/CTRL2 0.03fF
C49356 PAND2X1_6/Y POR2X1_407/A 0.03fF
C49357 POR2X1_66/B POR2X1_294/A 1.04fF
C49358 POR2X1_559/Y POR2X1_844/B 0.00fF
C49359 POR2X1_529/Y PAND2X1_793/Y 0.00fF
C49360 PAND2X1_489/CTRL PAND2X1_580/B 0.00fF
C49361 POR2X1_389/A POR2X1_664/Y 0.22fF
C49362 POR2X1_190/Y POR2X1_854/B 0.05fF
C49363 POR2X1_280/CTRL PAND2X1_552/B 0.01fF
C49364 PAND2X1_139/CTRL POR2X1_102/Y 0.01fF
C49365 POR2X1_465/B POR2X1_222/A 0.03fF
C49366 POR2X1_188/A POR2X1_294/A 0.03fF
C49367 PAND2X1_756/CTRL2 POR2X1_394/A 0.10fF
C49368 POR2X1_192/Y POR2X1_192/CTRL2 0.01fF
C49369 PAND2X1_62/O POR2X1_394/A 0.20fF
C49370 POR2X1_42/Y POR2X1_387/Y 0.10fF
C49371 POR2X1_734/A PAND2X1_48/A 0.07fF
C49372 PAND2X1_793/Y PAND2X1_574/CTRL 0.01fF
C49373 POR2X1_38/B PAND2X1_29/CTRL 0.01fF
C49374 POR2X1_740/Y POR2X1_228/Y 0.03fF
C49375 POR2X1_326/A POR2X1_448/Y 0.03fF
C49376 PAND2X1_591/O PAND2X1_56/A 0.01fF
C49377 POR2X1_177/a_16_28# POR2X1_72/B 0.00fF
C49378 POR2X1_785/a_16_28# POR2X1_566/B 0.02fF
C49379 PAND2X1_220/O POR2X1_142/Y 0.01fF
C49380 PAND2X1_403/CTRL2 POR2X1_20/B 0.06fF
C49381 POR2X1_502/A POR2X1_456/B 0.03fF
C49382 POR2X1_43/B PAND2X1_787/A 0.03fF
C49383 POR2X1_687/Y POR2X1_800/A 0.00fF
C49384 PAND2X1_41/B PAND2X1_328/CTRL 0.01fF
C49385 POR2X1_503/CTRL2 POR2X1_52/A 0.01fF
C49386 POR2X1_356/A POR2X1_180/B 0.70fF
C49387 PAND2X1_319/B PAND2X1_357/Y 0.01fF
C49388 POR2X1_325/A POR2X1_574/Y 0.03fF
C49389 POR2X1_96/A PAND2X1_641/O 0.01fF
C49390 PAND2X1_284/CTRL2 POR2X1_258/Y 0.01fF
C49391 POR2X1_7/B PAND2X1_155/CTRL2 0.03fF
C49392 POR2X1_166/CTRL2 POR2X1_73/Y 0.01fF
C49393 POR2X1_228/a_16_28# PAND2X1_52/Y -0.00fF
C49394 PAND2X1_239/O PAND2X1_52/B -0.00fF
C49395 PAND2X1_560/B VDD 0.41fF
C49396 POR2X1_387/Y POR2X1_309/Y 0.02fF
C49397 POR2X1_394/A INPUT_0 0.48fF
C49398 POR2X1_579/Y POR2X1_175/B 0.02fF
C49399 POR2X1_383/A PAND2X1_71/a_76_28# 0.02fF
C49400 PAND2X1_90/A PAND2X1_94/A 3.11fF
C49401 POR2X1_48/Y PAND2X1_196/O 0.04fF
C49402 POR2X1_218/Y PAND2X1_72/A 0.07fF
C49403 PAND2X1_48/B POR2X1_773/B 0.03fF
C49404 POR2X1_13/A POR2X1_599/CTRL 0.01fF
C49405 POR2X1_98/B POR2X1_68/B 0.02fF
C49406 PAND2X1_663/O POR2X1_413/A 0.02fF
C49407 POR2X1_68/A POR2X1_569/A 0.10fF
C49408 POR2X1_153/O PAND2X1_472/B 0.02fF
C49409 POR2X1_55/Y PAND2X1_508/CTRL 0.03fF
C49410 POR2X1_355/B POR2X1_209/CTRL 0.01fF
C49411 POR2X1_100/O PAND2X1_88/Y 0.08fF
C49412 PAND2X1_805/A PAND2X1_367/O 0.01fF
C49413 PAND2X1_865/Y PAND2X1_805/A 0.03fF
C49414 PAND2X1_23/Y POR2X1_463/Y 0.03fF
C49415 PAND2X1_476/A PAND2X1_721/O 0.03fF
C49416 POR2X1_751/Y POR2X1_7/B 0.04fF
C49417 PAND2X1_460/a_16_344# POR2X1_68/B 0.02fF
C49418 PAND2X1_23/Y POR2X1_756/Y 0.06fF
C49419 POR2X1_505/Y POR2X1_39/B 0.03fF
C49420 PAND2X1_81/O PAND2X1_63/B 0.04fF
C49421 PAND2X1_69/A POR2X1_725/Y 0.07fF
C49422 POR2X1_16/A PAND2X1_649/O 0.03fF
C49423 PAND2X1_832/CTRL2 POR2X1_39/B 0.06fF
C49424 POR2X1_486/a_16_28# POR2X1_705/B 0.03fF
C49425 POR2X1_349/CTRL PAND2X1_57/B 0.01fF
C49426 POR2X1_416/B POR2X1_251/A 0.03fF
C49427 PAND2X1_572/CTRL PAND2X1_656/A 0.01fF
C49428 POR2X1_574/A POR2X1_724/A 0.03fF
C49429 VDD PAND2X1_539/CTRL 0.00fF
C49430 POR2X1_614/A POR2X1_175/B 0.05fF
C49431 POR2X1_274/B POR2X1_573/A 0.01fF
C49432 INPUT_1 POR2X1_248/CTRL2 0.01fF
C49433 POR2X1_41/B PAND2X1_716/B 0.07fF
C49434 POR2X1_416/B POR2X1_72/B 0.14fF
C49435 POR2X1_845/a_76_344# POR2X1_532/A 0.00fF
C49436 POR2X1_851/O POR2X1_733/A 0.04fF
C49437 POR2X1_307/A PAND2X1_305/O 0.02fF
C49438 D_INPUT_1 POR2X1_362/A 0.03fF
C49439 PAND2X1_481/CTRL D_GATE_741 0.01fF
C49440 POR2X1_300/CTRL2 POR2X1_300/Y 0.01fF
C49441 POR2X1_78/B POR2X1_199/B 0.01fF
C49442 PAND2X1_65/B POR2X1_568/B 0.11fF
C49443 POR2X1_643/A PAND2X1_52/B 0.03fF
C49444 POR2X1_532/A PAND2X1_133/CTRL 0.01fF
C49445 POR2X1_722/B POR2X1_722/CTRL2 0.01fF
C49446 PAND2X1_833/CTRL2 POR2X1_39/B 0.03fF
C49447 POR2X1_294/B POR2X1_722/CTRL2 0.03fF
C49448 PAND2X1_510/CTRL2 POR2X1_73/Y 0.00fF
C49449 POR2X1_566/A PAND2X1_179/CTRL2 0.04fF
C49450 POR2X1_327/Y PAND2X1_674/O 0.01fF
C49451 POR2X1_62/Y PAND2X1_55/Y 1.16fF
C49452 D_GATE_222 POR2X1_332/a_16_28# 0.04fF
C49453 POR2X1_248/CTRL2 POR2X1_153/Y 0.15fF
C49454 POR2X1_119/Y PAND2X1_215/B 0.05fF
C49455 PAND2X1_357/Y PAND2X1_357/CTRL2 0.01fF
C49456 POR2X1_407/A PAND2X1_310/O 0.00fF
C49457 PAND2X1_180/O POR2X1_77/Y 0.17fF
C49458 INPUT_1 POR2X1_376/A 0.00fF
C49459 PAND2X1_865/CTRL PAND2X1_175/B 0.01fF
C49460 PAND2X1_96/B POR2X1_741/B 0.01fF
C49461 PAND2X1_69/A POR2X1_559/A 0.08fF
C49462 POR2X1_736/O POR2X1_675/Y 0.01fF
C49463 POR2X1_334/Y POR2X1_193/a_16_28# 0.06fF
C49464 POR2X1_542/B POR2X1_544/B 0.02fF
C49465 PAND2X1_661/B POR2X1_599/CTRL 0.01fF
C49466 POR2X1_540/m4_208_n4# POR2X1_703/A 0.15fF
C49467 PAND2X1_543/O POR2X1_77/Y 0.01fF
C49468 PAND2X1_301/O POR2X1_91/Y 0.07fF
C49469 POR2X1_577/a_16_28# POR2X1_570/Y 0.03fF
C49470 POR2X1_87/B PAND2X1_41/B 0.01fF
C49471 POR2X1_786/Y PAND2X1_48/A 0.02fF
C49472 POR2X1_3/A POR2X1_762/CTRL2 0.00fF
C49473 POR2X1_667/CTRL D_INPUT_0 0.00fF
C49474 POR2X1_356/A POR2X1_169/A 0.05fF
C49475 PAND2X1_831/Y POR2X1_153/Y 0.05fF
C49476 PAND2X1_862/B POR2X1_77/Y 0.04fF
C49477 POR2X1_64/O POR2X1_39/B 0.16fF
C49478 POR2X1_83/Y POR2X1_56/Y 0.19fF
C49479 POR2X1_775/CTRL POR2X1_191/Y 0.19fF
C49480 POR2X1_775/O POR2X1_192/B 0.24fF
C49481 POR2X1_66/Y PAND2X1_43/O 0.02fF
C49482 POR2X1_283/A PAND2X1_348/A 0.07fF
C49483 POR2X1_614/A POR2X1_4/Y 0.07fF
C49484 POR2X1_68/B POR2X1_561/Y 0.00fF
C49485 POR2X1_588/Y POR2X1_583/Y 0.18fF
C49486 POR2X1_446/B POR2X1_663/B 0.01fF
C49487 POR2X1_305/O POR2X1_7/B 0.18fF
C49488 POR2X1_126/O POR2X1_411/B 0.01fF
C49489 POR2X1_576/CTRL POR2X1_260/A 0.11fF
C49490 POR2X1_673/Y POR2X1_721/CTRL2 0.04fF
C49491 PAND2X1_353/a_16_344# PAND2X1_308/Y 0.01fF
C49492 PAND2X1_353/O PAND2X1_303/Y 0.03fF
C49493 POR2X1_369/CTRL POR2X1_315/Y 0.08fF
C49494 POR2X1_38/B POR2X1_4/Y 0.39fF
C49495 POR2X1_245/a_76_344# PAND2X1_156/A 0.03fF
C49496 PAND2X1_23/Y POR2X1_736/A 0.05fF
C49497 POR2X1_57/A POR2X1_397/O 0.01fF
C49498 POR2X1_566/O POR2X1_854/B 0.02fF
C49499 POR2X1_329/A POR2X1_594/CTRL 0.01fF
C49500 POR2X1_550/A POR2X1_550/B 0.05fF
C49501 PAND2X1_816/CTRL2 PAND2X1_52/B 0.01fF
C49502 POR2X1_565/B PAND2X1_52/B 0.01fF
C49503 POR2X1_20/B POR2X1_37/Y 4.40fF
C49504 PAND2X1_124/CTRL PAND2X1_123/Y 0.02fF
C49505 PAND2X1_779/O POR2X1_527/Y 0.02fF
C49506 POR2X1_416/B PAND2X1_547/CTRL2 0.03fF
C49507 POR2X1_62/Y PAND2X1_28/O 0.05fF
C49508 POR2X1_725/Y POR2X1_512/CTRL 0.08fF
C49509 PAND2X1_152/a_16_344# PAND2X1_72/A 0.02fF
C49510 POR2X1_83/B POR2X1_27/a_16_28# 0.03fF
C49511 POR2X1_166/O PAND2X1_326/B 0.01fF
C49512 POR2X1_499/A POR2X1_296/B 0.05fF
C49513 PAND2X1_631/A POR2X1_283/A 0.15fF
C49514 POR2X1_20/B POR2X1_279/CTRL 0.01fF
C49515 POR2X1_71/O POR2X1_394/A 0.03fF
C49516 PAND2X1_3/B POR2X1_260/A 0.01fF
C49517 POR2X1_407/A PAND2X1_52/B 0.05fF
C49518 POR2X1_68/A PAND2X1_72/A 20.46fF
C49519 POR2X1_149/CTRL POR2X1_78/A 0.01fF
C49520 POR2X1_54/Y POR2X1_55/CTRL2 0.01fF
C49521 POR2X1_619/A POR2X1_39/B 0.10fF
C49522 POR2X1_285/Y POR2X1_649/O 0.01fF
C49523 POR2X1_111/Y POR2X1_109/Y 0.02fF
C49524 POR2X1_456/B POR2X1_188/Y 0.44fF
C49525 PAND2X1_308/Y PAND2X1_716/B 0.00fF
C49526 POR2X1_54/Y POR2X1_590/A 0.03fF
C49527 PAND2X1_404/m4_208_n4# POR2X1_411/A 0.01fF
C49528 POR2X1_343/Y POR2X1_205/A 0.10fF
C49529 POR2X1_411/B PAND2X1_718/Y 0.05fF
C49530 POR2X1_313/CTRL2 POR2X1_167/Y 0.01fF
C49531 POR2X1_65/A POR2X1_760/A 2.31fF
C49532 PAND2X1_269/O POR2X1_236/Y 0.04fF
C49533 POR2X1_76/A POR2X1_296/B 0.02fF
C49534 POR2X1_661/A PAND2X1_385/CTRL -0.03fF
C49535 PAND2X1_59/B POR2X1_66/A 0.01fF
C49536 POR2X1_66/B POR2X1_286/B 0.31fF
C49537 PAND2X1_467/B POR2X1_694/Y 0.07fF
C49538 PAND2X1_9/Y POR2X1_750/B 0.03fF
C49539 POR2X1_856/B POR2X1_434/A 0.01fF
C49540 POR2X1_461/Y POR2X1_734/A 0.05fF
C49541 PAND2X1_632/B POR2X1_39/B 0.03fF
C49542 POR2X1_777/B POR2X1_341/A 0.07fF
C49543 POR2X1_604/O POR2X1_72/B 0.01fF
C49544 PAND2X1_497/CTRL2 POR2X1_267/A 0.03fF
C49545 POR2X1_670/O POR2X1_20/B 0.02fF
C49546 POR2X1_12/A POR2X1_748/A 0.03fF
C49547 POR2X1_394/A PAND2X1_379/CTRL2 0.12fF
C49548 POR2X1_472/O PAND2X1_52/B 0.01fF
C49549 POR2X1_841/B POR2X1_850/B 0.03fF
C49550 POR2X1_558/B POR2X1_78/A 0.05fF
C49551 POR2X1_660/Y D_INPUT_0 1.31fF
C49552 PAND2X1_72/A PAND2X1_315/CTRL2 0.01fF
C49553 POR2X1_49/Y PAND2X1_443/CTRL2 0.11fF
C49554 POR2X1_83/B PAND2X1_214/CTRL2 0.01fF
C49555 PAND2X1_246/a_16_344# INPUT_0 0.01fF
C49556 GATE_479 POR2X1_257/A 0.03fF
C49557 PAND2X1_207/O PAND2X1_200/Y 0.00fF
C49558 PAND2X1_39/B POR2X1_403/O 0.01fF
C49559 PAND2X1_569/B PAND2X1_326/O 0.01fF
C49560 POR2X1_816/CTRL2 INPUT_0 -0.00fF
C49561 PAND2X1_309/O POR2X1_814/A 0.17fF
C49562 PAND2X1_65/B POR2X1_341/A 0.09fF
C49563 PAND2X1_124/Y PAND2X1_195/O 0.06fF
C49564 POR2X1_180/B PAND2X1_72/A 0.03fF
C49565 POR2X1_648/CTRL2 PAND2X1_90/Y 0.06fF
C49566 PAND2X1_652/CTRL2 POR2X1_385/Y 0.01fF
C49567 POR2X1_20/B PAND2X1_151/CTRL2 0.00fF
C49568 PAND2X1_704/CTRL POR2X1_77/Y 0.00fF
C49569 POR2X1_411/B PAND2X1_580/B 0.03fF
C49570 POR2X1_49/Y PAND2X1_444/O 0.11fF
C49571 POR2X1_818/Y POR2X1_750/B 0.03fF
C49572 POR2X1_66/B POR2X1_630/a_16_28# 0.01fF
C49573 POR2X1_505/Y POR2X1_48/A 0.01fF
C49574 POR2X1_614/A POR2X1_458/Y 0.07fF
C49575 PAND2X1_226/CTRL2 POR2X1_227/A 0.00fF
C49576 POR2X1_14/Y POR2X1_753/Y 0.07fF
C49577 POR2X1_416/B PAND2X1_343/a_76_28# 0.02fF
C49578 PAND2X1_93/B POR2X1_543/A 0.03fF
C49579 POR2X1_814/A POR2X1_790/A 0.02fF
C49580 POR2X1_63/Y POR2X1_230/Y 0.03fF
C49581 PAND2X1_200/O POR2X1_32/A 0.04fF
C49582 POR2X1_666/a_16_28# POR2X1_102/Y 0.03fF
C49583 POR2X1_78/B POR2X1_602/CTRL2 0.02fF
C49584 POR2X1_568/A POR2X1_353/A 0.03fF
C49585 POR2X1_838/B POR2X1_838/a_16_28# 0.02fF
C49586 POR2X1_106/O POR2X1_251/A 0.08fF
C49587 POR2X1_20/B POR2X1_293/Y 0.34fF
C49588 PAND2X1_46/CTRL2 POR2X1_296/B 0.00fF
C49589 PAND2X1_716/B POR2X1_77/Y 0.03fF
C49590 POR2X1_383/a_16_28# POR2X1_383/Y 0.01fF
C49591 PAND2X1_207/CTRL2 VDD 0.00fF
C49592 POR2X1_491/O POR2X1_32/A 0.01fF
C49593 POR2X1_20/B PAND2X1_555/A 0.16fF
C49594 POR2X1_664/CTRL2 POR2X1_651/Y 0.01fF
C49595 POR2X1_846/Y POR2X1_790/A 0.03fF
C49596 PAND2X1_73/a_76_28# POR2X1_590/A 0.02fF
C49597 PAND2X1_459/O PAND2X1_58/A 0.01fF
C49598 PAND2X1_865/Y PAND2X1_440/CTRL2 0.00fF
C49599 POR2X1_518/CTRL2 POR2X1_77/Y 0.01fF
C49600 POR2X1_865/B POR2X1_814/A 0.03fF
C49601 POR2X1_220/B PAND2X1_90/Y 0.03fF
C49602 PAND2X1_6/Y POR2X1_287/A 0.01fF
C49603 PAND2X1_48/B POR2X1_471/A 0.34fF
C49604 POR2X1_586/Y POR2X1_585/CTRL 0.01fF
C49605 POR2X1_48/A PAND2X1_818/CTRL2 0.03fF
C49606 POR2X1_437/Y POR2X1_150/Y 0.04fF
C49607 POR2X1_852/B PAND2X1_39/O 0.16fF
C49608 POR2X1_477/Y POR2X1_480/A 0.08fF
C49609 POR2X1_863/A POR2X1_317/B 0.01fF
C49610 PAND2X1_20/A POR2X1_35/B 0.04fF
C49611 D_INPUT_0 POR2X1_497/Y 0.07fF
C49612 POR2X1_411/B PAND2X1_562/O 0.04fF
C49613 POR2X1_692/CTRL2 POR2X1_46/Y 0.01fF
C49614 POR2X1_29/A POR2X1_5/Y 0.21fF
C49615 POR2X1_474/CTRL PAND2X1_41/B 0.01fF
C49616 POR2X1_114/B POR2X1_475/CTRL 0.03fF
C49617 POR2X1_311/Y POR2X1_65/A 0.06fF
C49618 PAND2X1_400/CTRL2 VDD 0.00fF
C49619 POR2X1_349/a_16_28# POR2X1_343/Y 0.04fF
C49620 D_INPUT_0 PAND2X1_332/a_76_28# 0.02fF
C49621 POR2X1_411/B PAND2X1_337/A 0.08fF
C49622 POR2X1_861/A PAND2X1_72/A 0.01fF
C49623 POR2X1_432/CTRL POR2X1_236/Y 0.01fF
C49624 POR2X1_112/O PAND2X1_72/A 0.18fF
C49625 POR2X1_61/Y PAND2X1_394/O 0.13fF
C49626 PAND2X1_621/O POR2X1_9/Y 0.05fF
C49627 PAND2X1_48/B PAND2X1_248/CTRL2 0.01fF
C49628 POR2X1_287/B POR2X1_634/A 0.03fF
C49629 POR2X1_177/Y POR2X1_83/B 0.05fF
C49630 POR2X1_48/A POR2X1_411/O 0.01fF
C49631 POR2X1_669/B INPUT_0 0.29fF
C49632 POR2X1_490/Y PAND2X1_228/O 0.01fF
C49633 POR2X1_79/O PAND2X1_798/B 0.11fF
C49634 POR2X1_376/B POR2X1_482/Y 0.20fF
C49635 POR2X1_43/B PAND2X1_469/O 0.01fF
C49636 POR2X1_143/O D_INPUT_0 0.02fF
C49637 POR2X1_288/A POR2X1_734/A 0.00fF
C49638 POR2X1_23/Y PAND2X1_254/O 0.02fF
C49639 POR2X1_48/A PAND2X1_254/CTRL 0.01fF
C49640 POR2X1_35/B POR2X1_814/B 0.90fF
C49641 POR2X1_181/O PAND2X1_72/A 0.02fF
C49642 POR2X1_341/A POR2X1_541/CTRL 0.03fF
C49643 POR2X1_465/CTRL POR2X1_569/A 0.04fF
C49644 POR2X1_456/O POR2X1_186/Y 0.06fF
C49645 POR2X1_49/Y GATE_479 0.02fF
C49646 POR2X1_12/A PAND2X1_635/O 0.02fF
C49647 PAND2X1_65/B POR2X1_500/A 0.03fF
C49648 POR2X1_169/A PAND2X1_72/A 1.39fF
C49649 POR2X1_295/CTRL2 POR2X1_481/A 0.01fF
C49650 POR2X1_834/O POR2X1_513/B 0.01fF
C49651 POR2X1_675/CTRL VDD 0.00fF
C49652 POR2X1_78/A POR2X1_646/CTRL2 0.01fF
C49653 POR2X1_606/CTRL2 PAND2X1_32/B 0.05fF
C49654 POR2X1_399/A POR2X1_48/A 0.01fF
C49655 POR2X1_614/A POR2X1_266/O 0.05fF
C49656 POR2X1_20/B POR2X1_408/Y 0.01fF
C49657 POR2X1_330/a_16_28# PAND2X1_72/A 0.03fF
C49658 PAND2X1_259/CTRL2 POR2X1_258/Y 0.01fF
C49659 PAND2X1_557/A PAND2X1_362/B 0.03fF
C49660 POR2X1_260/B POR2X1_804/A 0.17fF
C49661 POR2X1_65/A POR2X1_485/CTRL2 0.03fF
C49662 POR2X1_260/B PAND2X1_316/a_76_28# 0.02fF
C49663 POR2X1_411/B PAND2X1_349/A 0.03fF
C49664 PAND2X1_498/CTRL POR2X1_590/A 0.01fF
C49665 POR2X1_49/Y PAND2X1_208/m4_208_n4# 0.08fF
C49666 POR2X1_669/B POR2X1_617/O 0.04fF
C49667 POR2X1_423/O POR2X1_372/Y 0.04fF
C49668 POR2X1_411/B PAND2X1_63/B 0.03fF
C49669 POR2X1_66/A D_GATE_222 0.10fF
C49670 PAND2X1_55/Y POR2X1_646/Y 0.07fF
C49671 POR2X1_72/B PAND2X1_512/Y 3.08fF
C49672 POR2X1_251/A PAND2X1_738/Y 0.05fF
C49673 POR2X1_83/B POR2X1_669/O 0.16fF
C49674 PAND2X1_6/Y POR2X1_808/B 0.01fF
C49675 POR2X1_257/A PAND2X1_175/B 0.03fF
C49676 POR2X1_389/Y VDD 0.46fF
C49677 PAND2X1_738/Y POR2X1_72/B 0.05fF
C49678 PAND2X1_93/B POR2X1_243/CTRL 0.01fF
C49679 INPUT_3 PAND2X1_28/CTRL 0.06fF
C49680 POR2X1_83/B PAND2X1_435/a_76_28# 0.01fF
C49681 POR2X1_846/Y POR2X1_754/a_56_344# 0.00fF
C49682 POR2X1_51/CTRL2 PAND2X1_635/Y 0.01fF
C49683 POR2X1_859/A POR2X1_94/A 0.02fF
C49684 POR2X1_624/Y POR2X1_366/A 0.07fF
C49685 PAND2X1_841/CTRL POR2X1_516/Y 0.09fF
C49686 POR2X1_720/A VDD 0.00fF
C49687 POR2X1_16/A POR2X1_150/Y 0.12fF
C49688 PAND2X1_73/Y POR2X1_800/A 0.00fF
C49689 POR2X1_308/O POR2X1_830/A 0.01fF
C49690 POR2X1_536/Y PAND2X1_364/B 0.02fF
C49691 POR2X1_130/A POR2X1_287/B 0.05fF
C49692 POR2X1_346/B PAND2X1_43/CTRL2 0.00fF
C49693 POR2X1_445/O POR2X1_750/B 0.09fF
C49694 PAND2X1_73/Y PAND2X1_79/a_16_344# 0.04fF
C49695 POR2X1_241/B POR2X1_341/CTRL 0.01fF
C49696 POR2X1_620/CTRL POR2X1_296/B 0.01fF
C49697 POR2X1_96/A PAND2X1_356/B 0.02fF
C49698 POR2X1_610/a_16_28# POR2X1_532/A 0.04fF
C49699 POR2X1_41/B PAND2X1_205/Y 7.19fF
C49700 PAND2X1_56/Y POR2X1_657/a_76_344# 0.03fF
C49701 POR2X1_66/B POR2X1_124/a_16_28# 0.01fF
C49702 POR2X1_114/B POR2X1_850/B 0.02fF
C49703 POR2X1_81/Y PAND2X1_500/a_16_344# 0.04fF
C49704 PAND2X1_116/CTRL2 PAND2X1_553/B 0.01fF
C49705 PAND2X1_394/O POR2X1_35/Y 0.02fF
C49706 POR2X1_66/B PAND2X1_638/CTRL2 0.10fF
C49707 PAND2X1_73/Y POR2X1_702/A 0.03fF
C49708 PAND2X1_96/B POR2X1_479/CTRL2 0.01fF
C49709 INPUT_2 POR2X1_104/CTRL2 0.01fF
C49710 D_INPUT_2 POR2X1_37/a_76_344# 0.02fF
C49711 PAND2X1_834/O POR2X1_677/Y 0.05fF
C49712 PAND2X1_622/O PAND2X1_621/Y 0.00fF
C49713 POR2X1_428/Y PAND2X1_726/B 0.07fF
C49714 POR2X1_407/A POR2X1_467/Y 0.16fF
C49715 PAND2X1_430/O PAND2X1_429/Y 0.00fF
C49716 PAND2X1_787/A POR2X1_298/Y 0.01fF
C49717 POR2X1_378/A D_INPUT_0 0.01fF
C49718 POR2X1_406/O POR2X1_5/Y 0.02fF
C49719 PAND2X1_643/CTRL2 POR2X1_595/Y 0.01fF
C49720 POR2X1_489/B POR2X1_68/B 0.04fF
C49721 POR2X1_748/A PAND2X1_506/a_76_28# 0.03fF
C49722 POR2X1_614/A POR2X1_450/A 0.01fF
C49723 POR2X1_347/B VDD 0.71fF
C49724 POR2X1_295/CTRL POR2X1_90/Y 0.10fF
C49725 POR2X1_566/A POR2X1_724/CTRL 0.28fF
C49726 POR2X1_56/B POR2X1_236/Y 0.33fF
C49727 PAND2X1_493/a_16_344# POR2X1_411/B 0.02fF
C49728 PAND2X1_658/A PAND2X1_793/A 0.01fF
C49729 POR2X1_60/Y POR2X1_56/Y 0.03fF
C49730 POR2X1_478/O POR2X1_444/Y 0.11fF
C49731 POR2X1_254/Y POR2X1_220/Y 0.07fF
C49732 INPUT_1 POR2X1_612/Y 0.07fF
C49733 POR2X1_15/O POR2X1_14/Y 0.05fF
C49734 PAND2X1_632/B POR2X1_48/A 0.04fF
C49735 POR2X1_525/a_16_28# POR2X1_763/Y 0.09fF
C49736 POR2X1_763/Y POR2X1_524/Y 0.01fF
C49737 PAND2X1_730/B PAND2X1_364/B 0.10fF
C49738 POR2X1_814/A POR2X1_568/B 0.18fF
C49739 PAND2X1_659/B PAND2X1_659/a_56_28# 0.00fF
C49740 POR2X1_52/A PAND2X1_580/B 0.03fF
C49741 PAND2X1_340/B POR2X1_394/A 0.09fF
C49742 POR2X1_502/A PAND2X1_57/B 1.12fF
C49743 POR2X1_12/O POR2X1_587/Y 0.10fF
C49744 POR2X1_416/B POR2X1_292/O 0.01fF
C49745 POR2X1_8/Y POR2X1_77/a_16_28# 0.00fF
C49746 PAND2X1_57/O POR2X1_404/Y 0.09fF
C49747 POR2X1_780/CTRL2 POR2X1_532/A 0.03fF
C49748 POR2X1_102/Y POR2X1_757/O 0.01fF
C49749 POR2X1_66/B POR2X1_389/A 0.03fF
C49750 POR2X1_590/A POR2X1_201/Y 0.18fF
C49751 POR2X1_96/A POR2X1_305/a_16_28# 0.02fF
C49752 POR2X1_528/Y POR2X1_422/Y 0.01fF
C49753 POR2X1_197/CTRL POR2X1_740/Y 0.01fF
C49754 D_INPUT_0 POR2X1_308/B 0.00fF
C49755 POR2X1_389/Y PAND2X1_32/B 0.08fF
C49756 POR2X1_327/Y POR2X1_274/A 0.03fF
C49757 POR2X1_639/Y POR2X1_750/B 0.01fF
C49758 PAND2X1_57/B POR2X1_247/CTRL 0.01fF
C49759 POR2X1_68/A POR2X1_632/A 0.02fF
C49760 PAND2X1_645/CTRL PAND2X1_602/Y 0.02fF
C49761 PAND2X1_735/Y POR2X1_494/Y 0.06fF
C49762 POR2X1_312/a_16_28# POR2X1_65/A 0.07fF
C49763 POR2X1_135/Y POR2X1_43/B 0.03fF
C49764 POR2X1_453/O PAND2X1_60/B 0.02fF
C49765 PAND2X1_58/A PAND2X1_382/a_16_344# 0.02fF
C49766 PAND2X1_697/O PAND2X1_90/Y 0.15fF
C49767 PAND2X1_785/Y POR2X1_55/Y 0.06fF
C49768 POR2X1_41/B PAND2X1_243/B 0.00fF
C49769 PAND2X1_58/A POR2X1_569/A 0.01fF
C49770 PAND2X1_478/O VDD -0.00fF
C49771 PAND2X1_411/O POR2X1_461/B 0.00fF
C49772 POR2X1_197/O PAND2X1_56/Y 0.06fF
C49773 POR2X1_856/B POR2X1_544/B 0.02fF
C49774 POR2X1_65/A POR2X1_38/Y 0.13fF
C49775 PAND2X1_263/O D_INPUT_1 0.01fF
C49776 PAND2X1_71/CTRL POR2X1_579/Y 0.00fF
C49777 POR2X1_697/CTRL PAND2X1_565/A 0.00fF
C49778 POR2X1_26/O POR2X1_32/A 0.01fF
C49779 POR2X1_83/B POR2X1_428/CTRL2 0.00fF
C49780 POR2X1_823/CTRL VDD -0.00fF
C49781 PAND2X1_605/O POR2X1_32/A 0.04fF
C49782 POR2X1_49/Y POR2X1_142/Y 0.82fF
C49783 PAND2X1_342/a_16_344# POR2X1_5/Y 0.00fF
C49784 POR2X1_20/Y VDD 0.11fF
C49785 POR2X1_257/A POR2X1_524/CTRL 0.01fF
C49786 POR2X1_79/A PAND2X1_794/B 0.01fF
C49787 POR2X1_38/Y PAND2X1_558/CTRL 0.00fF
C49788 POR2X1_471/A POR2X1_181/CTRL 0.00fF
C49789 PAND2X1_803/Y PAND2X1_360/a_76_28# 0.01fF
C49790 POR2X1_547/O POR2X1_502/A 0.03fF
C49791 POR2X1_708/O POR2X1_779/A 0.01fF
C49792 POR2X1_78/B PAND2X1_81/O 0.04fF
C49793 VDD POR2X1_747/Y 0.00fF
C49794 POR2X1_404/Y POR2X1_575/B 0.07fF
C49795 PAND2X1_90/Y POR2X1_758/O 0.03fF
C49796 POR2X1_188/A POR2X1_121/a_76_344# -0.00fF
C49797 POR2X1_68/B POR2X1_549/B 0.26fF
C49798 POR2X1_494/Y PAND2X1_493/Y 0.00fF
C49799 POR2X1_16/A PAND2X1_794/O 0.08fF
C49800 POR2X1_14/Y POR2X1_754/O 0.09fF
C49801 POR2X1_188/A POR2X1_710/Y 0.01fF
C49802 POR2X1_546/A POR2X1_705/CTRL 0.02fF
C49803 POR2X1_673/A POR2X1_38/B 0.03fF
C49804 POR2X1_73/O POR2X1_40/Y 0.01fF
C49805 POR2X1_72/B POR2X1_172/CTRL2 0.09fF
C49806 D_INPUT_0 POR2X1_5/CTRL 0.01fF
C49807 PAND2X1_629/O POR2X1_7/A 0.01fF
C49808 POR2X1_687/A POR2X1_750/B 0.03fF
C49809 PAND2X1_74/O POR2X1_456/B 0.02fF
C49810 POR2X1_706/B POR2X1_383/A 0.00fF
C49811 POR2X1_52/A POR2X1_315/CTRL 0.01fF
C49812 POR2X1_455/CTRL PAND2X1_60/B 0.09fF
C49813 POR2X1_335/A PAND2X1_498/O 0.02fF
C49814 POR2X1_95/a_76_344# POR2X1_12/A 0.00fF
C49815 POR2X1_376/B PAND2X1_349/A 0.03fF
C49816 PAND2X1_472/A POR2X1_669/CTRL 0.00fF
C49817 POR2X1_356/A POR2X1_782/A 0.11fF
C49818 POR2X1_278/A POR2X1_278/a_76_344# 0.01fF
C49819 POR2X1_102/Y POR2X1_394/A 0.27fF
C49820 POR2X1_376/B PAND2X1_63/B 0.03fF
C49821 VDD POR2X1_578/CTRL 0.00fF
C49822 PAND2X1_793/Y PAND2X1_548/CTRL2 0.01fF
C49823 POR2X1_614/A PAND2X1_71/CTRL 0.02fF
C49824 PAND2X1_84/Y POR2X1_91/Y 0.05fF
C49825 PAND2X1_93/a_76_28# POR2X1_404/Y 0.02fF
C49826 VDD POR2X1_318/A 0.05fF
C49827 POR2X1_559/B PAND2X1_65/B 0.01fF
C49828 PAND2X1_803/Y PAND2X1_543/a_16_344# 0.04fF
C49829 PAND2X1_562/B PAND2X1_346/Y 0.68fF
C49830 PAND2X1_69/A PAND2X1_176/CTRL 0.01fF
C49831 PAND2X1_730/a_56_28# POR2X1_42/Y 0.00fF
C49832 PAND2X1_23/Y PAND2X1_6/A 0.00fF
C49833 POR2X1_78/B POR2X1_780/B 0.01fF
C49834 POR2X1_284/O POR2X1_804/A 0.54fF
C49835 INPUT_1 PAND2X1_620/Y 0.06fF
C49836 POR2X1_96/A POR2X1_299/a_56_344# 0.00fF
C49837 PAND2X1_287/Y POR2X1_767/Y 0.03fF
C49838 POR2X1_763/Y PAND2X1_324/O 0.06fF
C49839 POR2X1_356/A PAND2X1_96/B 0.05fF
C49840 VDD POR2X1_713/B 1.55fF
C49841 POR2X1_66/B POR2X1_334/Y 0.07fF
C49842 POR2X1_804/A PAND2X1_369/O 0.16fF
C49843 POR2X1_283/A PAND2X1_715/CTRL2 0.03fF
C49844 PAND2X1_55/Y POR2X1_804/A 0.05fF
C49845 POR2X1_632/CTRL POR2X1_632/Y 0.01fF
C49846 POR2X1_49/Y PAND2X1_620/O 0.04fF
C49847 POR2X1_358/a_16_28# POR2X1_351/Y 0.02fF
C49848 POR2X1_828/Y POR2X1_260/A 0.01fF
C49849 PAND2X1_798/B PAND2X1_357/Y 0.07fF
C49850 POR2X1_440/CTRL2 POR2X1_440/B 0.02fF
C49851 D_INPUT_1 POR2X1_572/B 0.03fF
C49852 POR2X1_193/A POR2X1_724/A 0.07fF
C49853 POR2X1_590/A POR2X1_4/Y 0.07fF
C49854 POR2X1_854/CTRL2 POR2X1_776/B 0.02fF
C49855 POR2X1_35/Y POR2X1_562/B 0.01fF
C49856 PAND2X1_17/CTRL2 INPUT_6 0.01fF
C49857 PAND2X1_624/a_76_28# POR2X1_283/A 0.02fF
C49858 POR2X1_43/B POR2X1_816/A 0.03fF
C49859 PAND2X1_498/a_16_344# POR2X1_840/B 0.07fF
C49860 POR2X1_66/B PAND2X1_281/O 0.03fF
C49861 POR2X1_651/a_76_344# POR2X1_639/Y 0.01fF
C49862 PAND2X1_494/CTRL2 PAND2X1_32/B 0.01fF
C49863 PAND2X1_260/CTRL2 PAND2X1_345/Y 0.01fF
C49864 POR2X1_119/Y POR2X1_442/Y 0.01fF
C49865 POR2X1_383/A PAND2X1_322/CTRL2 0.10fF
C49866 POR2X1_65/A POR2X1_153/Y 0.12fF
C49867 POR2X1_462/B POR2X1_789/A 0.03fF
C49868 POR2X1_41/B PAND2X1_857/A 0.06fF
C49869 PAND2X1_864/B PAND2X1_568/B 6.83fF
C49870 PAND2X1_283/CTRL PAND2X1_96/B 0.00fF
C49871 POR2X1_38/Y PAND2X1_188/a_56_28# 0.00fF
C49872 PAND2X1_63/Y PAND2X1_81/CTRL2 0.01fF
C49873 POR2X1_306/CTRL2 POR2X1_43/B 0.02fF
C49874 POR2X1_407/A PAND2X1_743/O 0.08fF
C49875 D_INPUT_3 POR2X1_42/Y 0.03fF
C49876 PAND2X1_242/Y POR2X1_20/B 0.05fF
C49877 POR2X1_52/A PAND2X1_349/A 0.03fF
C49878 PAND2X1_450/CTRL2 POR2X1_425/Y 0.01fF
C49879 POR2X1_402/A PAND2X1_69/O 0.02fF
C49880 POR2X1_276/CTRL2 POR2X1_366/A 0.01fF
C49881 D_GATE_222 POR2X1_532/A 0.03fF
C49882 POR2X1_355/B POR2X1_726/Y 0.01fF
C49883 POR2X1_423/Y POR2X1_183/O 0.01fF
C49884 POR2X1_13/A PAND2X1_346/Y 0.01fF
C49885 POR2X1_614/A D_INPUT_1 0.15fF
C49886 POR2X1_57/A PAND2X1_837/CTRL2 0.03fF
C49887 POR2X1_416/B PAND2X1_640/B 0.01fF
C49888 POR2X1_41/B PAND2X1_374/O 0.05fF
C49889 POR2X1_78/CTRL PAND2X1_96/B 0.00fF
C49890 PAND2X1_715/B PAND2X1_715/O 0.00fF
C49891 POR2X1_741/Y POR2X1_318/A 0.07fF
C49892 PAND2X1_866/CTRL VDD -0.00fF
C49893 POR2X1_345/CTRL2 POR2X1_244/B 0.01fF
C49894 POR2X1_532/A POR2X1_140/A 0.01fF
C49895 POR2X1_301/A POR2X1_717/B 0.02fF
C49896 PAND2X1_319/B PAND2X1_182/CTRL2 0.05fF
C49897 PAND2X1_273/O PAND2X1_60/B 0.08fF
C49898 POR2X1_476/Y POR2X1_774/A 0.03fF
C49899 POR2X1_254/Y POR2X1_332/CTRL 0.02fF
C49900 POR2X1_38/B D_INPUT_1 1.98fF
C49901 POR2X1_508/A POR2X1_852/B 0.09fF
C49902 PAND2X1_705/a_16_344# POR2X1_526/Y 0.03fF
C49903 POR2X1_447/B PAND2X1_41/B 1.37fF
C49904 POR2X1_86/Y POR2X1_37/Y 0.06fF
C49905 POR2X1_669/B POR2X1_747/CTRL2 0.01fF
C49906 POR2X1_614/A POR2X1_724/A 0.01fF
C49907 POR2X1_41/B POR2X1_260/A 0.07fF
C49908 POR2X1_574/Y VDD 0.04fF
C49909 PAND2X1_341/B PAND2X1_231/O 0.00fF
C49910 POR2X1_489/A POR2X1_260/A 0.08fF
C49911 POR2X1_16/A PAND2X1_364/B 0.10fF
C49912 PAND2X1_23/Y POR2X1_101/Y 0.10fF
C49913 POR2X1_740/Y POR2X1_787/CTRL2 0.01fF
C49914 PAND2X1_96/B POR2X1_190/O 0.01fF
C49915 PAND2X1_90/A PAND2X1_133/O 0.04fF
C49916 PAND2X1_80/CTRL PAND2X1_71/Y 0.01fF
C49917 POR2X1_730/Y PAND2X1_48/B 0.03fF
C49918 POR2X1_318/A PAND2X1_32/B 0.07fF
C49919 PAND2X1_715/B POR2X1_293/Y 0.02fF
C49920 POR2X1_57/A POR2X1_165/CTRL2 0.01fF
C49921 POR2X1_283/A POR2X1_183/Y 0.03fF
C49922 POR2X1_383/A POR2X1_713/a_76_344# 0.01fF
C49923 POR2X1_618/m4_208_n4# POR2X1_751/m4_208_n4# 0.04fF
C49924 POR2X1_707/O PAND2X1_95/B 0.01fF
C49925 POR2X1_840/B PAND2X1_60/B 0.06fF
C49926 POR2X1_729/Y POR2X1_685/B 0.12fF
C49927 POR2X1_57/A PAND2X1_338/B -0.00fF
C49928 POR2X1_55/Y PAND2X1_348/A 0.50fF
C49929 PAND2X1_659/Y PAND2X1_579/B 0.03fF
C49930 POR2X1_852/B POR2X1_568/B 0.03fF
C49931 POR2X1_711/O POR2X1_713/B 0.18fF
C49932 POR2X1_383/A POR2X1_758/CTRL 0.01fF
C49933 PAND2X1_717/A POR2X1_275/Y 0.03fF
C49934 PAND2X1_96/B POR2X1_569/A 0.21fF
C49935 PAND2X1_58/A PAND2X1_72/A 0.06fF
C49936 PAND2X1_472/CTRL2 PAND2X1_472/A 0.02fF
C49937 POR2X1_391/Y POR2X1_260/A 0.07fF
C49938 PAND2X1_372/O PAND2X1_48/A 0.05fF
C49939 VDD PAND2X1_352/B 0.19fF
C49940 POR2X1_814/A POR2X1_341/A 0.10fF
C49941 POR2X1_52/A PAND2X1_708/a_16_344# 0.01fF
C49942 PAND2X1_57/B POR2X1_188/Y 0.04fF
C49943 PAND2X1_805/A POR2X1_533/Y 0.06fF
C49944 POR2X1_137/Y POR2X1_218/CTRL2 0.00fF
C49945 PAND2X1_177/O POR2X1_180/A 0.01fF
C49946 PAND2X1_649/A INPUT_0 0.03fF
C49947 PAND2X1_371/O POR2X1_773/A 0.04fF
C49948 POR2X1_411/B POR2X1_411/A 0.06fF
C49949 POR2X1_81/A INPUT_0 0.11fF
C49950 POR2X1_548/A PAND2X1_63/B 0.00fF
C49951 PAND2X1_90/A POR2X1_561/Y -0.00fF
C49952 POR2X1_576/O POR2X1_500/Y 0.18fF
C49953 PAND2X1_641/O POR2X1_38/Y 0.13fF
C49954 POR2X1_837/B PAND2X1_419/CTRL 0.01fF
C49955 POR2X1_172/Y POR2X1_530/CTRL2 0.01fF
C49956 POR2X1_712/CTRL2 POR2X1_260/A 0.01fF
C49957 POR2X1_750/B POR2X1_568/A 0.03fF
C49958 POR2X1_366/O PAND2X1_60/B 0.07fF
C49959 POR2X1_653/CTRL2 POR2X1_711/Y 0.02fF
C49960 PAND2X1_348/Y PAND2X1_348/O 0.01fF
C49961 POR2X1_177/CTRL POR2X1_90/Y 0.08fF
C49962 PAND2X1_717/Y PAND2X1_723/A 1.54fF
C49963 POR2X1_590/O POR2X1_796/A 0.12fF
C49964 POR2X1_99/B POR2X1_740/Y 0.05fF
C49965 PAND2X1_631/A POR2X1_55/Y 2.66fF
C49966 POR2X1_510/Y POR2X1_456/B 0.03fF
C49967 POR2X1_129/Y POR2X1_73/Y 0.03fF
C49968 POR2X1_537/Y POR2X1_68/A 0.05fF
C49969 POR2X1_821/Y POR2X1_394/A 4.07fF
C49970 PAND2X1_48/B PAND2X1_696/CTRL 0.01fF
C49971 POR2X1_13/A POR2X1_372/CTRL 0.01fF
C49972 PAND2X1_6/Y POR2X1_359/CTRL2 0.03fF
C49973 PAND2X1_48/B POR2X1_542/CTRL 0.00fF
C49974 PAND2X1_610/CTRL2 D_INPUT_2 0.03fF
C49975 PAND2X1_716/B POR2X1_52/Y 0.00fF
C49976 PAND2X1_23/Y POR2X1_359/a_16_28# 0.02fF
C49977 PAND2X1_511/a_16_344# PAND2X1_56/A 0.01fF
C49978 POR2X1_259/CTRL2 POR2X1_260/A 0.03fF
C49979 POR2X1_293/Y POR2X1_372/CTRL2 0.01fF
C49980 POR2X1_568/Y POR2X1_545/O 0.04fF
C49981 POR2X1_16/A PAND2X1_849/B 0.03fF
C49982 PAND2X1_659/Y POR2X1_73/Y 0.07fF
C49983 POR2X1_7/B POR2X1_588/CTRL 0.01fF
C49984 PAND2X1_830/Y POR2X1_416/B 0.01fF
C49985 PAND2X1_691/Y PAND2X1_686/O 0.05fF
C49986 POR2X1_366/A POR2X1_186/B 0.03fF
C49987 PAND2X1_243/B POR2X1_77/Y 0.03fF
C49988 POR2X1_435/Y PAND2X1_72/A 0.17fF
C49989 POR2X1_416/B POR2X1_7/B 3.07fF
C49990 PAND2X1_189/CTRL POR2X1_854/B 0.01fF
C49991 POR2X1_730/Y POR2X1_151/a_16_28# 0.02fF
C49992 PAND2X1_508/Y POR2X1_7/A 0.03fF
C49993 PAND2X1_527/O PAND2X1_111/B 0.02fF
C49994 PAND2X1_690/O POR2X1_260/A 0.00fF
C49995 PAND2X1_687/B POR2X1_73/Y 0.02fF
C49996 POR2X1_83/A POR2X1_39/B 0.61fF
C49997 PAND2X1_160/O POR2X1_394/A 0.02fF
C49998 POR2X1_780/B POR2X1_294/A 0.01fF
C49999 POR2X1_353/A POR2X1_444/Y 0.16fF
C50000 POR2X1_677/Y POR2X1_432/Y 0.02fF
C50001 PAND2X1_742/B POR2X1_331/CTRL2 0.01fF
C50002 POR2X1_68/A POR2X1_555/CTRL 0.01fF
C50003 PAND2X1_82/Y POR2X1_294/A 0.01fF
C50004 PAND2X1_549/B POR2X1_171/Y 0.19fF
C50005 PAND2X1_175/B PAND2X1_865/A 0.01fF
C50006 POR2X1_90/Y POR2X1_39/B 0.25fF
C50007 POR2X1_67/Y PAND2X1_390/Y 0.02fF
C50008 POR2X1_78/Y POR2X1_590/A 0.03fF
C50009 POR2X1_647/B POR2X1_286/CTRL 0.01fF
C50010 PAND2X1_73/Y POR2X1_688/a_16_28# 0.02fF
C50011 POR2X1_294/Y PAND2X1_67/CTRL2 0.00fF
C50012 POR2X1_411/B POR2X1_32/A 0.29fF
C50013 POR2X1_54/Y POR2X1_66/A 0.03fF
C50014 PAND2X1_169/CTRL POR2X1_142/Y 0.03fF
C50015 POR2X1_813/a_76_344# POR2X1_263/Y 0.01fF
C50016 PAND2X1_850/Y POR2X1_283/A 0.03fF
C50017 POR2X1_334/Y POR2X1_97/a_16_28# 0.05fF
C50018 POR2X1_316/O POR2X1_153/Y 0.01fF
C50019 PAND2X1_221/Y POR2X1_79/Y 0.02fF
C50020 POR2X1_60/A POR2X1_20/B 0.16fF
C50021 PAND2X1_79/Y POR2X1_500/CTRL2 0.00fF
C50022 INPUT_1 POR2X1_397/a_16_28# 0.01fF
C50023 POR2X1_48/A PAND2X1_590/O 0.17fF
C50024 POR2X1_20/B POR2X1_591/A 0.02fF
C50025 PAND2X1_96/B PAND2X1_72/A 0.16fF
C50026 PAND2X1_60/B PAND2X1_56/A 0.05fF
C50027 PAND2X1_35/A PAND2X1_34/a_16_344# 0.03fF
C50028 POR2X1_417/Y POR2X1_411/B 0.03fF
C50029 POR2X1_441/Y PAND2X1_731/B 0.05fF
C50030 POR2X1_416/B POR2X1_108/a_16_28# 0.03fF
C50031 POR2X1_590/A POR2X1_266/O 0.07fF
C50032 PAND2X1_417/m4_208_n4# POR2X1_750/B 0.03fF
C50033 POR2X1_78/A PAND2X1_609/CTRL 0.01fF
C50034 PAND2X1_261/CTRL2 POR2X1_814/A 0.04fF
C50035 POR2X1_566/B POR2X1_567/CTRL 0.06fF
C50036 POR2X1_66/B PAND2X1_60/CTRL 0.01fF
C50037 POR2X1_38/a_16_28# POR2X1_37/Y 0.03fF
C50038 POR2X1_356/A PAND2X1_438/a_16_344# 0.05fF
C50039 PAND2X1_86/CTRL POR2X1_243/Y 0.02fF
C50040 POR2X1_491/a_16_28# POR2X1_150/Y 0.03fF
C50041 PAND2X1_800/O POR2X1_760/Y 0.00fF
C50042 PAND2X1_199/O PAND2X1_123/Y 0.02fF
C50043 POR2X1_602/a_16_28# POR2X1_296/B 0.04fF
C50044 POR2X1_41/B POR2X1_329/A 0.11fF
C50045 PAND2X1_732/A POR2X1_39/B 0.23fF
C50046 POR2X1_96/A PAND2X1_464/B 0.07fF
C50047 POR2X1_460/Y POR2X1_459/CTRL2 0.01fF
C50048 POR2X1_850/A PAND2X1_39/B 0.02fF
C50049 POR2X1_411/B PAND2X1_741/B 0.03fF
C50050 POR2X1_82/CTRL PAND2X1_9/Y 0.01fF
C50051 POR2X1_335/O POR2X1_556/A 0.02fF
C50052 PAND2X1_246/CTRL POR2X1_404/Y 0.00fF
C50053 POR2X1_493/B PAND2X1_72/A 0.06fF
C50054 PAND2X1_503/O PAND2X1_52/B 0.07fF
C50055 POR2X1_257/A POR2X1_272/Y 0.03fF
C50056 POR2X1_669/B POR2X1_102/Y 0.12fF
C50057 PAND2X1_628/a_16_344# PAND2X1_88/Y 0.01fF
C50058 PAND2X1_138/CTRL POR2X1_39/B 0.11fF
C50059 POR2X1_89/O POR2X1_376/B 0.07fF
C50060 PAND2X1_406/O POR2X1_362/B 0.02fF
C50061 POR2X1_106/a_76_344# POR2X1_102/Y 0.01fF
C50062 PAND2X1_56/Y PAND2X1_45/CTRL2 0.40fF
C50063 POR2X1_423/Y D_INPUT_0 0.03fF
C50064 POR2X1_54/Y PAND2X1_293/O -0.00fF
C50065 PAND2X1_807/a_76_28# PAND2X1_221/Y 0.02fF
C50066 POR2X1_110/Y POR2X1_39/B 0.20fF
C50067 POR2X1_49/Y POR2X1_409/B 0.02fF
C50068 POR2X1_470/a_16_28# POR2X1_466/Y -0.00fF
C50069 POR2X1_680/Y POR2X1_150/Y 1.72fF
C50070 POR2X1_66/B POR2X1_98/a_16_28# 0.02fF
C50071 PAND2X1_439/O POR2X1_90/Y 0.17fF
C50072 PAND2X1_65/B PAND2X1_65/CTRL2 0.00fF
C50073 PAND2X1_66/a_76_28# POR2X1_5/Y 0.01fF
C50074 PAND2X1_65/B POR2X1_678/Y 0.03fF
C50075 POR2X1_566/A POR2X1_454/O 0.04fF
C50076 PAND2X1_73/Y PAND2X1_42/CTRL2 0.03fF
C50077 POR2X1_83/B POR2X1_748/A 0.15fF
C50078 PAND2X1_436/O INPUT_0 0.02fF
C50079 POR2X1_812/A POR2X1_800/CTRL 0.05fF
C50080 POR2X1_189/Y POR2X1_411/B 0.02fF
C50081 POR2X1_57/A PAND2X1_717/A 0.03fF
C50082 D_INPUT_5 POR2X1_638/CTRL 0.01fF
C50083 POR2X1_754/Y POR2X1_625/O 0.06fF
C50084 POR2X1_753/Y POR2X1_625/CTRL2 0.04fF
C50085 POR2X1_168/CTRL POR2X1_168/A 0.01fF
C50086 POR2X1_485/Y PAND2X1_705/a_16_344# 0.01fF
C50087 POR2X1_376/B POR2X1_32/A 0.13fF
C50088 POR2X1_647/B POR2X1_294/B 0.03fF
C50089 POR2X1_411/B POR2X1_184/Y 0.05fF
C50090 POR2X1_597/Y POR2X1_683/Y 0.00fF
C50091 POR2X1_462/a_16_28# PAND2X1_69/A 0.03fF
C50092 PAND2X1_23/Y PAND2X1_24/O 0.00fF
C50093 PAND2X1_73/Y POR2X1_640/A 0.02fF
C50094 POR2X1_399/O POR2X1_609/Y 0.09fF
C50095 POR2X1_614/A POR2X1_137/B 0.01fF
C50096 POR2X1_847/A POR2X1_49/Y 0.11fF
C50097 POR2X1_109/CTRL POR2X1_7/B 0.00fF
C50098 POR2X1_296/B POR2X1_788/a_16_28# 0.09fF
C50099 POR2X1_812/A POR2X1_801/O 0.01fF
C50100 POR2X1_52/A POR2X1_89/O 0.01fF
C50101 POR2X1_52/A PAND2X1_97/CTRL 0.01fF
C50102 POR2X1_115/CTRL2 POR2X1_218/Y 0.07fF
C50103 POR2X1_10/CTRL2 POR2X1_9/Y 0.01fF
C50104 PAND2X1_263/O POR2X1_78/A 0.01fF
C50105 PAND2X1_651/Y POR2X1_411/B 0.05fF
C50106 POR2X1_559/B POR2X1_814/A 0.02fF
C50107 POR2X1_355/B POR2X1_856/B 0.03fF
C50108 POR2X1_253/O PAND2X1_6/A 0.02fF
C50109 POR2X1_834/O VDD 0.00fF
C50110 PAND2X1_93/B POR2X1_193/A 0.03fF
C50111 PAND2X1_93/B POR2X1_579/Y 0.03fF
C50112 PAND2X1_766/O PAND2X1_41/B 0.01fF
C50113 POR2X1_677/Y POR2X1_394/A 0.05fF
C50114 POR2X1_335/a_16_28# POR2X1_66/A 0.03fF
C50115 POR2X1_473/O POR2X1_391/Y 0.04fF
C50116 POR2X1_568/B POR2X1_180/Y 0.02fF
C50117 POR2X1_335/A POR2X1_274/A 0.03fF
C50118 PAND2X1_354/A PAND2X1_562/B 0.07fF
C50119 POR2X1_241/CTRL VDD -0.00fF
C50120 POR2X1_399/CTRL2 PAND2X1_403/B 0.07fF
C50121 PAND2X1_93/B POR2X1_572/B 0.06fF
C50122 POR2X1_517/a_16_28# POR2X1_667/A 0.05fF
C50123 INPUT_3 POR2X1_38/B 0.18fF
C50124 POR2X1_83/B POR2X1_418/O 0.02fF
C50125 POR2X1_9/Y POR2X1_394/A 0.33fF
C50126 POR2X1_150/Y PAND2X1_388/Y 0.07fF
C50127 POR2X1_262/Y PAND2X1_560/O 0.05fF
C50128 POR2X1_602/B PAND2X1_65/B 0.03fF
C50129 PAND2X1_250/a_16_344# POR2X1_287/B 0.01fF
C50130 POR2X1_130/A POR2X1_288/a_76_344# 0.04fF
C50131 PAND2X1_48/B POR2X1_218/Y 0.07fF
C50132 POR2X1_360/A PAND2X1_15/CTRL 0.06fF
C50133 POR2X1_54/Y POR2X1_532/A 0.03fF
C50134 PAND2X1_221/Y PAND2X1_730/A 0.14fF
C50135 POR2X1_14/Y PAND2X1_377/O 0.00fF
C50136 POR2X1_52/A POR2X1_32/A 5.64fF
C50137 PAND2X1_790/CTRL2 POR2X1_93/A 0.00fF
C50138 POR2X1_490/Y POR2X1_52/Y 2.58fF
C50139 POR2X1_329/A PAND2X1_308/Y 0.02fF
C50140 POR2X1_111/Y PAND2X1_717/A 0.05fF
C50141 PAND2X1_471/B POR2X1_14/Y 0.00fF
C50142 PAND2X1_658/A POR2X1_37/Y 0.03fF
C50143 PAND2X1_195/a_76_28# POR2X1_236/Y 0.01fF
C50144 POR2X1_600/Y PAND2X1_645/B 0.00fF
C50145 PAND2X1_402/O POR2X1_397/Y 0.06fF
C50146 POR2X1_40/Y VDD 4.89fF
C50147 POR2X1_707/B PAND2X1_57/B 0.00fF
C50148 POR2X1_614/A PAND2X1_93/B 0.10fF
C50149 POR2X1_516/O POR2X1_23/Y 0.01fF
C50150 POR2X1_78/A POR2X1_579/Y 0.06fF
C50151 POR2X1_569/m4_208_n4# PAND2X1_41/B 0.07fF
C50152 POR2X1_81/Y PAND2X1_573/B 0.01fF
C50153 POR2X1_35/B VDD 0.50fF
C50154 PAND2X1_275/a_16_344# D_INPUT_0 0.02fF
C50155 PAND2X1_863/B PAND2X1_249/CTRL 0.01fF
C50156 PAND2X1_23/Y POR2X1_843/O 0.03fF
C50157 POR2X1_196/O POR2X1_205/Y 0.02fF
C50158 POR2X1_41/B PAND2X1_361/O 0.02fF
C50159 PAND2X1_217/B PAND2X1_659/B 0.00fF
C50160 INPUT_7 POR2X1_2/CTRL 0.00fF
C50161 POR2X1_13/A PAND2X1_354/A 0.03fF
C50162 POR2X1_78/A POR2X1_572/B 0.01fF
C50163 POR2X1_120/CTRL2 PAND2X1_90/Y 0.09fF
C50164 POR2X1_48/A POR2X1_90/Y 0.10fF
C50165 PAND2X1_93/B POR2X1_38/B 0.13fF
C50166 POR2X1_102/Y PAND2X1_174/CTRL 0.01fF
C50167 PAND2X1_20/A PAND2X1_226/a_16_344# 0.02fF
C50168 PAND2X1_787/Y PAND2X1_473/B 0.49fF
C50169 POR2X1_407/A POR2X1_843/CTRL 0.00fF
C50170 POR2X1_567/B POR2X1_190/CTRL 0.14fF
C50171 POR2X1_632/a_56_344# PAND2X1_88/Y 0.00fF
C50172 PAND2X1_46/m4_208_n4# INPUT_0 0.15fF
C50173 PAND2X1_80/a_56_28# PAND2X1_41/B 0.00fF
C50174 POR2X1_147/A POR2X1_296/B 0.04fF
C50175 POR2X1_52/A POR2X1_417/Y 0.02fF
C50176 POR2X1_52/A POR2X1_419/Y 0.04fF
C50177 POR2X1_708/CTRL2 PAND2X1_90/Y 0.06fF
C50178 POR2X1_220/Y PAND2X1_41/B 0.03fF
C50179 PAND2X1_340/CTRL INPUT_0 0.07fF
C50180 POR2X1_49/Y PAND2X1_351/Y 0.02fF
C50181 PAND2X1_222/A PAND2X1_799/a_76_28# 0.01fF
C50182 POR2X1_37/Y POR2X1_73/Y 0.15fF
C50183 POR2X1_716/CTRL POR2X1_303/B 0.01fF
C50184 POR2X1_129/O POR2X1_90/Y 0.10fF
C50185 POR2X1_47/CTRL POR2X1_748/A 0.09fF
C50186 POR2X1_356/A POR2X1_355/A 0.01fF
C50187 PAND2X1_848/B PAND2X1_848/O 0.04fF
C50188 PAND2X1_55/Y POR2X1_794/B 0.03fF
C50189 PAND2X1_463/a_76_28# PAND2X1_459/Y 0.02fF
C50190 PAND2X1_65/B POR2X1_546/A 0.55fF
C50191 POR2X1_462/B POR2X1_590/A 0.06fF
C50192 PAND2X1_422/O PAND2X1_93/B -0.00fF
C50193 POR2X1_748/A PAND2X1_709/O 0.00fF
C50194 PAND2X1_499/Y INPUT_0 0.07fF
C50195 POR2X1_614/A POR2X1_78/A 20.78fF
C50196 PAND2X1_818/O POR2X1_5/Y 0.02fF
C50197 PAND2X1_41/B POR2X1_404/Y 0.03fF
C50198 POR2X1_417/Y POR2X1_152/A 0.01fF
C50199 PAND2X1_20/A POR2X1_775/CTRL2 0.02fF
C50200 POR2X1_590/A D_INPUT_1 0.26fF
C50201 POR2X1_68/A POR2X1_812/A 0.19fF
C50202 PAND2X1_69/A POR2X1_296/B 2.19fF
C50203 POR2X1_322/O POR2X1_40/Y 0.00fF
C50204 POR2X1_255/Y POR2X1_516/Y 0.03fF
C50205 POR2X1_32/A PAND2X1_186/O 0.01fF
C50206 POR2X1_821/Y POR2X1_669/B 0.01fF
C50207 POR2X1_271/Y POR2X1_184/Y 0.02fF
C50208 POR2X1_594/CTRL POR2X1_594/A 0.01fF
C50209 PAND2X1_274/O POR2X1_272/Y 0.05fF
C50210 PAND2X1_659/B VDD 0.00fF
C50211 POR2X1_78/A POR2X1_38/B 0.07fF
C50212 POR2X1_596/A PAND2X1_73/Y 0.03fF
C50213 POR2X1_62/Y PAND2X1_201/O 0.02fF
C50214 POR2X1_327/Y POR2X1_276/B 0.02fF
C50215 POR2X1_481/O VDD 0.00fF
C50216 PAND2X1_205/Y PAND2X1_742/B 0.03fF
C50217 POR2X1_305/Y POR2X1_72/B 0.04fF
C50218 PAND2X1_583/CTRL2 POR2X1_750/B 0.01fF
C50219 POR2X1_516/CTRL POR2X1_423/Y 0.01fF
C50220 POR2X1_791/O POR2X1_637/B 0.04fF
C50221 POR2X1_113/Y POR2X1_650/CTRL2 0.00fF
C50222 PAND2X1_244/B POR2X1_37/Y 0.07fF
C50223 PAND2X1_319/O PAND2X1_317/Y 0.01fF
C50224 POR2X1_499/CTRL2 POR2X1_456/B 0.01fF
C50225 POR2X1_66/B POR2X1_140/CTRL 0.01fF
C50226 POR2X1_267/A POR2X1_318/A 0.03fF
C50227 PAND2X1_707/Y PAND2X1_712/B 0.00fF
C50228 PAND2X1_735/CTRL POR2X1_293/Y 0.03fF
C50229 PAND2X1_512/Y POR2X1_7/B 0.01fF
C50230 PAND2X1_501/B POR2X1_494/Y 0.00fF
C50231 PAND2X1_738/Y POR2X1_7/B 0.05fF
C50232 POR2X1_13/A INPUT_5 0.03fF
C50233 PAND2X1_787/Y PAND2X1_390/O 0.04fF
C50234 POR2X1_376/B PAND2X1_242/a_16_344# 0.02fF
C50235 PAND2X1_275/CTRL2 VDD -0.00fF
C50236 POR2X1_41/B PAND2X1_515/CTRL 0.31fF
C50237 PAND2X1_474/A POR2X1_816/A 0.35fF
C50238 PAND2X1_715/O PAND2X1_115/B 0.02fF
C50239 POR2X1_186/Y PAND2X1_146/m4_208_n4# 0.08fF
C50240 POR2X1_48/A PAND2X1_732/A -0.00fF
C50241 PAND2X1_23/Y POR2X1_740/a_16_28# 0.03fF
C50242 PAND2X1_793/Y POR2X1_46/Y 0.03fF
C50243 POR2X1_777/B POR2X1_500/Y 0.05fF
C50244 PAND2X1_108/O PAND2X1_55/Y 0.14fF
C50245 PAND2X1_56/Y POR2X1_308/CTRL 0.14fF
C50246 PAND2X1_679/CTRL2 PAND2X1_69/A 0.01fF
C50247 POR2X1_824/Y PAND2X1_403/B 0.07fF
C50248 POR2X1_777/B PAND2X1_150/CTRL 0.12fF
C50249 PAND2X1_65/B POR2X1_712/Y 0.01fF
C50250 POR2X1_329/A POR2X1_77/Y 0.10fF
C50251 POR2X1_52/A PAND2X1_35/Y 0.02fF
C50252 POR2X1_186/Y POR2X1_540/A 0.03fF
C50253 PAND2X1_48/B POR2X1_115/CTRL 0.00fF
C50254 POR2X1_668/O POR2X1_816/A 0.02fF
C50255 POR2X1_443/a_16_28# POR2X1_192/B 0.04fF
C50256 PAND2X1_651/Y POR2X1_376/B 0.03fF
C50257 POR2X1_392/B PAND2X1_153/CTRL 0.08fF
C50258 POR2X1_49/Y PAND2X1_560/CTRL2 0.00fF
C50259 POR2X1_536/CTRL2 POR2X1_102/Y 0.01fF
C50260 POR2X1_121/B PAND2X1_300/CTRL2 0.03fF
C50261 POR2X1_463/Y POR2X1_792/CTRL 0.09fF
C50262 PAND2X1_318/a_16_344# POR2X1_96/A 0.01fF
C50263 PAND2X1_264/CTRL POR2X1_83/B 0.00fF
C50264 VDD POR2X1_587/Y 0.09fF
C50265 POR2X1_199/CTRL2 POR2X1_740/Y 0.51fF
C50266 POR2X1_290/a_16_28# PAND2X1_642/B 0.01fF
C50267 PAND2X1_73/Y POR2X1_598/O 0.01fF
C50268 PAND2X1_824/CTRL2 PAND2X1_41/B 0.03fF
C50269 PAND2X1_206/CTRL PAND2X1_6/A 0.04fF
C50270 POR2X1_68/A PAND2X1_58/O 0.04fF
C50271 POR2X1_60/Y PAND2X1_99/Y 0.02fF
C50272 POR2X1_65/A POR2X1_591/Y 0.01fF
C50273 POR2X1_300/a_16_28# POR2X1_272/Y 0.02fF
C50274 POR2X1_153/O POR2X1_37/Y 0.01fF
C50275 PAND2X1_848/B VDD 0.26fF
C50276 POR2X1_44/CTRL INPUT_6 0.01fF
C50277 POR2X1_197/Y POR2X1_244/a_56_344# 0.01fF
C50278 PAND2X1_65/B POR2X1_500/Y 0.03fF
C50279 PAND2X1_115/B POR2X1_293/Y 0.82fF
C50280 POR2X1_102/Y POR2X1_172/a_56_344# 0.00fF
C50281 PAND2X1_213/Y PAND2X1_220/Y 0.00fF
C50282 POR2X1_718/CTRL2 POR2X1_832/A 0.02fF
C50283 POR2X1_664/a_76_344# PAND2X1_73/Y 0.00fF
C50284 PAND2X1_6/Y POR2X1_194/B 0.02fF
C50285 POR2X1_401/CTRL2 POR2X1_68/B 0.01fF
C50286 PAND2X1_341/A POR2X1_236/Y 0.03fF
C50287 PAND2X1_859/A POR2X1_283/A 0.02fF
C50288 PAND2X1_476/A PAND2X1_404/Y 0.03fF
C50289 PAND2X1_20/A POR2X1_576/O 0.05fF
C50290 PAND2X1_97/Y PAND2X1_351/A 0.00fF
C50291 POR2X1_614/A PAND2X1_129/a_76_28# 0.01fF
C50292 POR2X1_134/Y VDD 0.12fF
C50293 PAND2X1_658/A POR2X1_293/Y 0.03fF
C50294 PAND2X1_13/a_16_344# PAND2X1_60/B 0.03fF
C50295 POR2X1_78/A POR2X1_772/a_16_28# 0.01fF
C50296 POR2X1_406/Y POR2X1_73/Y 0.05fF
C50297 POR2X1_93/A POR2X1_236/Y 0.06fF
C50298 POR2X1_550/CTRL VDD 0.00fF
C50299 PAND2X1_55/Y PAND2X1_178/O 0.04fF
C50300 INPUT_1 POR2X1_49/CTRL2 0.01fF
C50301 PAND2X1_23/Y PAND2X1_504/CTRL2 0.01fF
C50302 POR2X1_236/Y POR2X1_91/Y 0.03fF
C50303 POR2X1_661/A POR2X1_655/O 0.05fF
C50304 PAND2X1_96/B POR2X1_244/B 0.03fF
C50305 POR2X1_65/A POR2X1_167/O 0.01fF
C50306 POR2X1_76/Y POR2X1_112/Y 0.06fF
C50307 PAND2X1_254/O PAND2X1_658/B 0.01fF
C50308 POR2X1_510/A POR2X1_579/Y 0.03fF
C50309 POR2X1_790/a_16_28# POR2X1_790/B 0.03fF
C50310 PAND2X1_94/A POR2X1_734/A 0.15fF
C50311 PAND2X1_48/B POR2X1_68/A 3.16fF
C50312 POR2X1_16/A PAND2X1_240/CTRL2 0.11fF
C50313 PAND2X1_90/Y POR2X1_854/B 0.05fF
C50314 PAND2X1_4/O PAND2X1_8/Y 0.04fF
C50315 POR2X1_52/A PAND2X1_651/Y 0.05fF
C50316 POR2X1_315/Y PAND2X1_803/A 0.14fF
C50317 POR2X1_557/A PAND2X1_41/B 0.03fF
C50318 PAND2X1_281/CTRL2 POR2X1_285/Y 0.09fF
C50319 PAND2X1_90/Y POR2X1_710/B 0.12fF
C50320 POR2X1_455/O POR2X1_222/A 0.02fF
C50321 POR2X1_319/A POR2X1_169/A 0.03fF
C50322 POR2X1_66/A POR2X1_4/Y 0.19fF
C50323 POR2X1_499/A POR2X1_717/B 0.79fF
C50324 POR2X1_590/A POR2X1_620/B 0.01fF
C50325 PAND2X1_215/B PAND2X1_723/O 0.06fF
C50326 POR2X1_41/B POR2X1_57/A 0.19fF
C50327 PAND2X1_41/B PAND2X1_184/O 0.01fF
C50328 POR2X1_590/A POR2X1_362/CTRL2 0.01fF
C50329 POR2X1_293/Y POR2X1_73/Y 0.28fF
C50330 POR2X1_66/B POR2X1_557/B 0.03fF
C50331 PAND2X1_106/O VDD 0.00fF
C50332 PAND2X1_170/CTRL2 PAND2X1_169/Y 0.00fF
C50333 POR2X1_43/B PAND2X1_469/B 1.37fF
C50334 PAND2X1_57/B POR2X1_711/a_16_28# 0.02fF
C50335 POR2X1_718/O POR2X1_834/Y 0.13fF
C50336 POR2X1_220/Y POR2X1_228/Y 0.07fF
C50337 POR2X1_203/Y POR2X1_294/B 0.02fF
C50338 PAND2X1_57/B POR2X1_510/Y 0.03fF
C50339 POR2X1_740/Y POR2X1_112/Y 0.01fF
C50340 POR2X1_21/O INPUT_4 0.04fF
C50341 POR2X1_537/Y PAND2X1_58/A 0.03fF
C50342 POR2X1_254/Y POR2X1_222/A 0.07fF
C50343 POR2X1_81/Y POR2X1_91/Y 0.01fF
C50344 POR2X1_791/O POR2X1_791/B 0.00fF
C50345 POR2X1_791/CTRL POR2X1_791/A 0.01fF
C50346 PAND2X1_848/A POR2X1_38/B 0.01fF
C50347 PAND2X1_20/A PAND2X1_396/CTRL2 0.01fF
C50348 POR2X1_416/B PAND2X1_606/O 0.04fF
C50349 POR2X1_96/A POR2X1_283/A 0.20fF
C50350 POR2X1_78/B PAND2X1_232/O 0.12fF
C50351 POR2X1_579/Y PAND2X1_173/CTRL 0.00fF
C50352 POR2X1_297/CTRL2 PAND2X1_359/Y 0.01fF
C50353 POR2X1_96/A POR2X1_134/CTRL 0.01fF
C50354 POR2X1_531/a_16_28# POR2X1_73/Y 0.03fF
C50355 POR2X1_41/B POR2X1_229/Y 0.11fF
C50356 POR2X1_515/Y POR2X1_513/Y 0.00fF
C50357 POR2X1_136/Y POR2X1_7/B 0.04fF
C50358 PAND2X1_65/B POR2X1_520/B 0.01fF
C50359 POR2X1_368/Y PAND2X1_457/O -0.00fF
C50360 PAND2X1_835/a_16_344# PAND2X1_852/B 0.02fF
C50361 INPUT_6 POR2X1_587/CTRL2 0.03fF
C50362 PAND2X1_649/A POR2X1_102/Y 0.00fF
C50363 PAND2X1_555/O PAND2X1_566/Y 0.17fF
C50364 POR2X1_52/A POR2X1_503/Y 0.01fF
C50365 PAND2X1_866/a_16_344# PAND2X1_805/A 0.02fF
C50366 POR2X1_187/CTRL POR2X1_79/Y 0.01fF
C50367 PAND2X1_472/CTRL2 PAND2X1_673/Y 0.04fF
C50368 PAND2X1_276/CTRL2 POR2X1_129/Y 0.01fF
C50369 POR2X1_504/a_16_28# POR2X1_504/Y 0.02fF
C50370 POR2X1_669/B POR2X1_761/A 0.00fF
C50371 PAND2X1_832/O PAND2X1_508/Y 0.03fF
C50372 POR2X1_81/A POR2X1_102/Y 0.03fF
C50373 POR2X1_807/A PAND2X1_142/a_16_344# 0.03fF
C50374 PAND2X1_714/B PAND2X1_731/B 0.35fF
C50375 POR2X1_390/B POR2X1_114/Y 0.31fF
C50376 POR2X1_730/Y POR2X1_728/B 0.44fF
C50377 PAND2X1_29/O POR2X1_68/B 0.13fF
C50378 POR2X1_383/A POR2X1_662/Y 0.07fF
C50379 POR2X1_287/B POR2X1_773/A 0.03fF
C50380 PAND2X1_824/B POR2X1_214/CTRL2 0.05fF
C50381 POR2X1_567/B POR2X1_181/Y 0.05fF
C50382 POR2X1_492/Y POR2X1_60/A 0.17fF
C50383 POR2X1_712/O POR2X1_712/Y 0.00fF
C50384 POR2X1_180/B PAND2X1_48/B 0.14fF
C50385 POR2X1_304/a_16_28# POR2X1_153/Y 0.02fF
C50386 POR2X1_8/Y POR2X1_618/CTRL2 0.00fF
C50387 POR2X1_81/A PAND2X1_436/A 0.02fF
C50388 PAND2X1_63/Y POR2X1_493/CTRL2 0.02fF
C50389 INPUT_1 POR2X1_20/O 0.18fF
C50390 POR2X1_278/Y POR2X1_394/A 0.19fF
C50391 POR2X1_41/B POR2X1_111/Y 0.03fF
C50392 POR2X1_78/B POR2X1_195/CTRL 0.01fF
C50393 POR2X1_189/Y POR2X1_679/B 0.09fF
C50394 PAND2X1_858/Y POR2X1_91/Y 1.97fF
C50395 PAND2X1_785/Y POR2X1_129/Y 0.03fF
C50396 VDD POR2X1_533/O 0.00fF
C50397 POR2X1_203/O POR2X1_203/Y 0.00fF
C50398 PAND2X1_449/O POR2X1_329/A 0.06fF
C50399 POR2X1_203/Y PAND2X1_111/B 0.01fF
C50400 PAND2X1_652/A PAND2X1_593/Y 0.01fF
C50401 INPUT_6 D_INPUT_6 0.44fF
C50402 POR2X1_829/A POR2X1_394/A 0.03fF
C50403 PAND2X1_109/CTRL2 PAND2X1_41/B 0.01fF
C50404 POR2X1_113/O PAND2X1_96/B 0.01fF
C50405 POR2X1_567/B POR2X1_535/CTRL 0.00fF
C50406 PAND2X1_675/A PAND2X1_336/O 0.07fF
C50407 PAND2X1_631/A POR2X1_511/Y 0.32fF
C50408 POR2X1_532/A POR2X1_148/B 0.05fF
C50409 PAND2X1_71/CTRL2 PAND2X1_71/Y 0.01fF
C50410 POR2X1_9/Y POR2X1_818/a_16_28# 0.09fF
C50411 POR2X1_21/a_76_344# POR2X1_460/A 0.03fF
C50412 POR2X1_407/Y PAND2X1_765/CTRL 0.01fF
C50413 POR2X1_327/Y PAND2X1_604/CTRL 0.01fF
C50414 PAND2X1_94/A POR2X1_786/Y 0.03fF
C50415 PAND2X1_798/B PAND2X1_579/A 0.04fF
C50416 PAND2X1_445/O PAND2X1_308/Y 0.04fF
C50417 POR2X1_664/Y POR2X1_774/A 0.03fF
C50418 POR2X1_416/B POR2X1_750/B 0.06fF
C50419 PAND2X1_633/CTRL2 POR2X1_77/Y 0.00fF
C50420 PAND2X1_496/CTRL2 PAND2X1_48/A 0.08fF
C50421 INPUT_1 PAND2X1_341/m4_208_n4# 0.12fF
C50422 POR2X1_539/A POR2X1_188/CTRL2 0.09fF
C50423 POR2X1_68/B POR2X1_773/CTRL2 0.00fF
C50424 POR2X1_49/O POR2X1_14/Y 0.01fF
C50425 POR2X1_622/A POR2X1_622/a_16_28# 0.03fF
C50426 PAND2X1_651/Y PAND2X1_510/CTRL 0.01fF
C50427 POR2X1_280/CTRL POR2X1_280/Y 0.01fF
C50428 POR2X1_840/CTRL POR2X1_834/Y 0.01fF
C50429 POR2X1_302/B POR2X1_325/B 0.12fF
C50430 POR2X1_416/B PAND2X1_220/Y 6.80fF
C50431 PAND2X1_859/O POR2X1_77/Y 0.03fF
C50432 POR2X1_335/Y POR2X1_260/A 0.01fF
C50433 POR2X1_391/Y POR2X1_559/A 0.10fF
C50434 POR2X1_832/B POR2X1_802/A 0.28fF
C50435 POR2X1_283/A POR2X1_7/A 0.27fF
C50436 POR2X1_57/A POR2X1_291/O 0.01fF
C50437 POR2X1_25/O D_INPUT_4 0.01fF
C50438 POR2X1_68/B POR2X1_571/CTRL2 0.09fF
C50439 POR2X1_283/A PAND2X1_130/O 0.05fF
C50440 POR2X1_493/CTRL2 POR2X1_260/A 0.03fF
C50441 PAND2X1_106/CTRL2 POR2X1_276/Y 0.01fF
C50442 POR2X1_390/B POR2X1_113/Y 0.04fF
C50443 POR2X1_131/Y PAND2X1_803/Y 0.03fF
C50444 POR2X1_461/Y POR2X1_859/CTRL2 0.01fF
C50445 POR2X1_435/Y POR2X1_532/O 0.05fF
C50446 POR2X1_188/CTRL POR2X1_456/B 0.01fF
C50447 INPUT_2 POR2X1_394/A 0.01fF
C50448 PAND2X1_94/A PAND2X1_27/CTRL2 0.11fF
C50449 PAND2X1_23/Y POR2X1_112/CTRL 0.01fF
C50450 D_INPUT_1 POR2X1_749/O 0.02fF
C50451 POR2X1_119/Y PAND2X1_575/A 0.03fF
C50452 INPUT_0 POR2X1_39/B 0.28fF
C50453 PAND2X1_661/Y PAND2X1_121/O 0.02fF
C50454 PAND2X1_6/Y PAND2X1_48/A 0.03fF
C50455 POR2X1_318/O POR2X1_471/A 0.06fF
C50456 POR2X1_281/Y POR2X1_102/Y 0.01fF
C50457 POR2X1_101/Y POR2X1_218/O 0.05fF
C50458 POR2X1_669/B POR2X1_9/Y 0.15fF
C50459 POR2X1_834/Y POR2X1_725/Y 0.22fF
C50460 PAND2X1_69/A POR2X1_342/CTRL 0.02fF
C50461 POR2X1_503/O POR2X1_503/Y 0.01fF
C50462 PAND2X1_847/CTRL POR2X1_820/Y 0.01fF
C50463 PAND2X1_525/a_76_28# PAND2X1_52/B 0.02fF
C50464 POR2X1_259/B POR2X1_510/Y 0.03fF
C50465 POR2X1_416/B POR2X1_425/CTRL2 0.00fF
C50466 POR2X1_293/Y PAND2X1_358/CTRL 0.03fF
C50467 POR2X1_856/O POR2X1_863/A 0.00fF
C50468 PAND2X1_48/B POR2X1_169/A 0.03fF
C50469 POR2X1_791/A PAND2X1_48/A 0.05fF
C50470 POR2X1_390/B POR2X1_260/A 0.02fF
C50471 POR2X1_669/B POR2X1_827/a_16_28# 0.02fF
C50472 POR2X1_814/A POR2X1_29/A 0.01fF
C50473 POR2X1_196/Y POR2X1_99/B 0.02fF
C50474 POR2X1_737/A PAND2X1_60/B 1.68fF
C50475 POR2X1_186/CTRL2 POR2X1_353/A 0.01fF
C50476 PAND2X1_854/A POR2X1_314/Y 0.02fF
C50477 POR2X1_532/A POR2X1_4/Y 0.08fF
C50478 POR2X1_776/B PAND2X1_52/B 0.06fF
C50479 POR2X1_713/B PAND2X1_692/CTRL 0.01fF
C50480 POR2X1_383/A POR2X1_62/Y 0.03fF
C50481 POR2X1_43/a_16_28# POR2X1_42/Y 0.05fF
C50482 POR2X1_397/Y POR2X1_825/Y 0.29fF
C50483 PAND2X1_286/O GATE_222 0.02fF
C50484 PAND2X1_349/A PAND2X1_716/B 0.04fF
C50485 POR2X1_456/B POR2X1_317/B 0.01fF
C50486 POR2X1_305/CTRL POR2X1_305/Y 0.01fF
C50487 POR2X1_151/O POR2X1_186/B 0.09fF
C50488 PAND2X1_404/CTRL2 POR2X1_411/A 0.08fF
C50489 POR2X1_69/CTRL PAND2X1_206/B 0.00fF
C50490 POR2X1_69/O POR2X1_67/Y 0.01fF
C50491 PAND2X1_787/A PAND2X1_352/Y 0.00fF
C50492 PAND2X1_838/B PAND2X1_640/B 0.01fF
C50493 POR2X1_602/B POR2X1_814/A 0.05fF
C50494 POR2X1_835/B POR2X1_506/B 0.01fF
C50495 INPUT_1 PAND2X1_508/Y 0.03fF
C50496 POR2X1_270/Y POR2X1_222/CTRL2 0.01fF
C50497 PAND2X1_631/CTRL POR2X1_416/B 0.01fF
C50498 PAND2X1_865/Y PAND2X1_854/A 0.02fF
C50499 POR2X1_49/O POR2X1_55/Y 0.16fF
C50500 POR2X1_122/CTRL2 POR2X1_394/A 0.09fF
C50501 POR2X1_532/A POR2X1_160/a_16_28# -0.00fF
C50502 POR2X1_565/CTRL PAND2X1_52/B 0.03fF
C50503 POR2X1_747/O POR2X1_747/Y 0.01fF
C50504 POR2X1_78/B PAND2X1_628/a_76_28# 0.04fF
C50505 POR2X1_567/B POR2X1_434/CTRL 0.14fF
C50506 POR2X1_462/CTRL2 POR2X1_734/A 0.03fF
C50507 PAND2X1_22/O PAND2X1_3/A 0.04fF
C50508 POR2X1_343/Y POR2X1_573/A 0.05fF
C50509 POR2X1_61/O POR2X1_447/B 0.06fF
C50510 POR2X1_57/A POR2X1_77/Y 0.24fF
C50511 PAND2X1_508/Y POR2X1_153/Y 0.36fF
C50512 POR2X1_13/A PAND2X1_458/CTRL 0.01fF
C50513 POR2X1_180/B POR2X1_181/CTRL 0.00fF
C50514 POR2X1_539/a_56_344# POR2X1_567/A 0.00fF
C50515 POR2X1_66/B PAND2X1_43/CTRL 0.01fF
C50516 POR2X1_681/Y POR2X1_32/A 0.08fF
C50517 POR2X1_9/Y PAND2X1_751/CTRL 0.04fF
C50518 POR2X1_826/a_16_28# POR2X1_55/Y 0.07fF
C50519 PAND2X1_458/CTRL2 POR2X1_293/Y 0.01fF
C50520 POR2X1_411/B POR2X1_94/A 0.06fF
C50521 PAND2X1_717/A PAND2X1_84/Y 0.12fF
C50522 POR2X1_9/Y POR2X1_617/CTRL2 0.03fF
C50523 PAND2X1_9/Y POR2X1_40/Y 0.03fF
C50524 PAND2X1_747/O PAND2X1_52/B 0.01fF
C50525 POR2X1_294/A POR2X1_195/CTRL 0.00fF
C50526 PAND2X1_96/B POR2X1_579/CTRL 0.01fF
C50527 POR2X1_250/Y PAND2X1_580/B 0.03fF
C50528 POR2X1_629/CTRL2 POR2X1_629/B 0.02fF
C50529 PAND2X1_643/A PAND2X1_538/CTRL2 0.01fF
C50530 POR2X1_647/B POR2X1_643/A 0.20fF
C50531 POR2X1_814/A POR2X1_546/A 0.03fF
C50532 PAND2X1_405/a_16_344# POR2X1_46/Y 0.02fF
C50533 POR2X1_741/O POR2X1_741/B 0.25fF
C50534 PAND2X1_93/B POR2X1_590/A 0.03fF
C50535 POR2X1_430/O POR2X1_669/B 0.02fF
C50536 PAND2X1_860/A POR2X1_56/Y 0.00fF
C50537 PAND2X1_662/Y PAND2X1_659/Y 0.01fF
C50538 POR2X1_54/Y PAND2X1_23/CTRL2 0.09fF
C50539 POR2X1_556/A POR2X1_362/B 0.00fF
C50540 POR2X1_479/B POR2X1_288/CTRL 0.02fF
C50541 POR2X1_63/Y POR2X1_230/CTRL 0.01fF
C50542 POR2X1_753/Y POR2X1_37/Y 0.05fF
C50543 PAND2X1_73/Y D_INPUT_0 0.11fF
C50544 POR2X1_12/A POR2X1_429/a_16_28# 0.05fF
C50545 POR2X1_559/A POR2X1_383/Y 0.16fF
C50546 PAND2X1_73/Y POR2X1_811/A 0.02fF
C50547 POR2X1_83/B POR2X1_263/Y 0.05fF
C50548 POR2X1_111/Y POR2X1_77/Y 0.02fF
C50549 POR2X1_610/CTRL PAND2X1_41/B 0.01fF
C50550 PAND2X1_65/B PAND2X1_39/B 0.17fF
C50551 POR2X1_333/A POR2X1_477/Y 0.02fF
C50552 POR2X1_79/a_16_28# PAND2X1_354/A 0.01fF
C50553 PAND2X1_803/Y PAND2X1_860/A 2.49fF
C50554 PAND2X1_400/O POR2X1_394/Y -0.00fF
C50555 POR2X1_78/A POR2X1_590/A 0.22fF
C50556 POR2X1_14/Y PAND2X1_381/Y 0.03fF
C50557 POR2X1_838/B POR2X1_202/B 0.31fF
C50558 POR2X1_67/Y POR2X1_619/CTRL 0.01fF
C50559 POR2X1_129/Y POR2X1_589/a_16_28# 0.04fF
C50560 POR2X1_541/B POR2X1_76/Y 0.12fF
C50561 POR2X1_657/Y POR2X1_220/Y 0.03fF
C50562 POR2X1_478/CTRL2 POR2X1_480/A 0.04fF
C50563 POR2X1_681/Y POR2X1_682/a_16_28# 0.03fF
C50564 PAND2X1_20/A POR2X1_33/O 0.01fF
C50565 POR2X1_49/Y POR2X1_626/CTRL2 0.00fF
C50566 POR2X1_508/A POR2X1_568/B 0.06fF
C50567 POR2X1_130/A POR2X1_624/Y 0.07fF
C50568 PAND2X1_244/B PAND2X1_242/Y 0.28fF
C50569 PAND2X1_234/O PAND2X1_88/Y 0.02fF
C50570 PAND2X1_317/O POR2X1_167/Y 0.06fF
C50571 POR2X1_707/B PAND2X1_25/a_16_344# 0.01fF
C50572 POR2X1_456/CTRL2 POR2X1_66/A 0.10fF
C50573 POR2X1_834/O POR2X1_808/A 0.02fF
C50574 POR2X1_66/A PAND2X1_52/Y 0.11fF
C50575 POR2X1_20/B PAND2X1_269/CTRL2 0.03fF
C50576 PAND2X1_73/Y PAND2X1_278/CTRL2 0.01fF
C50577 PAND2X1_48/A POR2X1_725/CTRL 0.01fF
C50578 POR2X1_48/A PAND2X1_62/O 0.06fF
C50579 POR2X1_180/O POR2X1_181/Y 0.01fF
C50580 POR2X1_43/B PAND2X1_466/A 0.04fF
C50581 POR2X1_604/Y POR2X1_72/B 0.01fF
C50582 POR2X1_548/CTRL POR2X1_66/A 0.03fF
C50583 POR2X1_693/Y POR2X1_485/Y 0.00fF
C50584 PAND2X1_262/CTRL POR2X1_296/B 0.12fF
C50585 PAND2X1_48/A PAND2X1_52/B 0.03fF
C50586 PAND2X1_622/CTRL POR2X1_669/B 0.00fF
C50587 PAND2X1_307/O POR2X1_14/Y 0.16fF
C50588 POR2X1_866/CTRL2 POR2X1_750/B 0.01fF
C50589 POR2X1_75/Y PAND2X1_332/Y 0.03fF
C50590 POR2X1_753/Y POR2X1_615/O 0.02fF
C50591 POR2X1_192/B PAND2X1_52/B 0.18fF
C50592 PAND2X1_307/O PAND2X1_453/A 0.03fF
C50593 PAND2X1_20/A POR2X1_777/B 0.05fF
C50594 POR2X1_365/Y POR2X1_212/A 0.03fF
C50595 POR2X1_20/B POR2X1_396/CTRL2 0.01fF
C50596 PAND2X1_48/B PAND2X1_271/CTRL 0.01fF
C50597 PAND2X1_241/Y POR2X1_329/A 0.01fF
C50598 POR2X1_816/CTRL POR2X1_816/A 0.01fF
C50599 POR2X1_498/CTRL2 PAND2X1_205/A 0.00fF
C50600 POR2X1_48/A INPUT_0 0.15fF
C50601 POR2X1_405/a_16_28# POR2X1_296/B 0.11fF
C50602 PAND2X1_3/A VDD 0.20fF
C50603 PAND2X1_208/CTRL2 POR2X1_40/Y 0.03fF
C50604 PAND2X1_73/Y PAND2X1_90/Y 0.14fF
C50605 POR2X1_856/B POR2X1_570/CTRL2 0.03fF
C50606 POR2X1_330/CTRL2 PAND2X1_52/B 0.01fF
C50607 POR2X1_496/a_16_28# POR2X1_55/Y -0.00fF
C50608 POR2X1_260/B POR2X1_795/CTRL 0.01fF
C50609 PAND2X1_558/Y PAND2X1_561/A 0.03fF
C50610 PAND2X1_20/A PAND2X1_65/B 5.46fF
C50611 PAND2X1_215/B PAND2X1_124/Y 0.07fF
C50612 POR2X1_368/Y POR2X1_257/A 0.04fF
C50613 POR2X1_102/Y PAND2X1_499/Y 0.03fF
C50614 POR2X1_67/CTRL PAND2X1_658/A 0.01fF
C50615 POR2X1_706/CTRL VDD 0.00fF
C50616 POR2X1_20/B PAND2X1_546/m4_208_n4# 0.07fF
C50617 PAND2X1_6/Y POR2X1_803/O 0.17fF
C50618 POR2X1_48/CTRL2 POR2X1_60/A 0.01fF
C50619 PAND2X1_659/CTRL POR2X1_498/Y 0.01fF
C50620 PAND2X1_620/Y POR2X1_72/B 0.03fF
C50621 POR2X1_502/A POR2X1_97/A 0.08fF
C50622 POR2X1_43/B PAND2X1_477/CTRL2 0.03fF
C50623 POR2X1_65/A POR2X1_72/B 2.59fF
C50624 POR2X1_624/Y POR2X1_844/B 0.01fF
C50625 POR2X1_13/A POR2X1_496/Y 0.00fF
C50626 POR2X1_186/Y POR2X1_798/CTRL 0.13fF
C50627 POR2X1_760/A POR2X1_283/A 0.06fF
C50628 POR2X1_814/B POR2X1_777/B 0.03fF
C50629 POR2X1_849/CTRL POR2X1_94/A 0.04fF
C50630 PAND2X1_862/B POR2X1_32/A 0.03fF
C50631 PAND2X1_58/A PAND2X1_58/O 0.05fF
C50632 PAND2X1_55/O POR2X1_94/A 0.01fF
C50633 PAND2X1_73/Y PAND2X1_760/O 0.02fF
C50634 POR2X1_633/Y POR2X1_633/A 0.01fF
C50635 PAND2X1_65/B POR2X1_254/CTRL 0.01fF
C50636 POR2X1_20/B POR2X1_142/Y 0.03fF
C50637 POR2X1_446/B POR2X1_804/A 0.03fF
C50638 POR2X1_72/B PAND2X1_558/CTRL 0.01fF
C50639 PAND2X1_436/A PAND2X1_499/Y 0.50fF
C50640 POR2X1_60/A PAND2X1_579/B 0.02fF
C50641 POR2X1_45/Y POR2X1_23/Y 0.07fF
C50642 PAND2X1_635/m4_208_n4# INPUT_6 0.12fF
C50643 PAND2X1_61/CTRL POR2X1_55/Y 0.14fF
C50644 PAND2X1_220/Y PAND2X1_192/Y 0.01fF
C50645 POR2X1_829/A POR2X1_669/B 0.00fF
C50646 POR2X1_20/B PAND2X1_785/a_76_28# 0.01fF
C50647 PAND2X1_250/O PAND2X1_65/B 0.00fF
C50648 D_INPUT_5 POR2X1_460/A 0.02fF
C50649 POR2X1_624/Y POR2X1_573/A 0.03fF
C50650 POR2X1_49/Y POR2X1_58/CTRL2 0.00fF
C50651 POR2X1_20/B PAND2X1_175/B 0.02fF
C50652 PAND2X1_810/A VDD 0.07fF
C50653 POR2X1_94/O POR2X1_23/Y 0.01fF
C50654 POR2X1_753/Y POR2X1_293/Y 0.00fF
C50655 D_GATE_662 POR2X1_66/A 0.08fF
C50656 POR2X1_96/A POR2X1_14/Y 0.25fF
C50657 POR2X1_814/B PAND2X1_65/B 0.10fF
C50658 POR2X1_96/A PAND2X1_453/A 0.03fF
C50659 POR2X1_857/B POR2X1_78/A 0.03fF
C50660 POR2X1_71/Y POR2X1_497/CTRL2 0.01fF
C50661 POR2X1_863/CTRL2 PAND2X1_73/Y 0.01fF
C50662 PAND2X1_798/B D_INPUT_0 0.03fF
C50663 PAND2X1_512/O INPUT_0 0.01fF
C50664 POR2X1_556/A POR2X1_553/A 0.03fF
C50665 POR2X1_376/B POR2X1_381/O 0.02fF
C50666 POR2X1_843/O POR2X1_733/A 0.02fF
C50667 POR2X1_13/A PAND2X1_733/A 0.03fF
C50668 POR2X1_83/B PAND2X1_215/B 0.72fF
C50669 POR2X1_654/B VDD 0.37fF
C50670 POR2X1_378/A POR2X1_54/Y 0.01fF
C50671 POR2X1_428/Y PAND2X1_711/a_76_28# 0.01fF
C50672 POR2X1_344/CTRL POR2X1_344/A 0.01fF
C50673 POR2X1_155/a_76_344# POR2X1_467/Y 0.01fF
C50674 PAND2X1_48/B PAND2X1_58/A 0.06fF
C50675 PAND2X1_578/Y PAND2X1_568/B 0.03fF
C50676 POR2X1_334/A PAND2X1_86/O 0.00fF
C50677 POR2X1_462/B POR2X1_66/A 0.03fF
C50678 PAND2X1_787/A POR2X1_298/CTRL 0.04fF
C50679 PAND2X1_3/A PAND2X1_32/B 0.10fF
C50680 PAND2X1_49/CTRL2 POR2X1_29/A 0.03fF
C50681 POR2X1_66/A D_INPUT_1 0.07fF
C50682 POR2X1_148/O POR2X1_148/B 0.00fF
C50683 PAND2X1_192/Y PAND2X1_739/Y 0.01fF
C50684 POR2X1_614/A POR2X1_450/CTRL2 0.03fF
C50685 POR2X1_850/A VDD 0.19fF
C50686 POR2X1_692/CTRL POR2X1_526/Y 0.01fF
C50687 POR2X1_510/A POR2X1_590/A 0.00fF
C50688 POR2X1_5/Y VDD 4.08fF
C50689 POR2X1_296/B POR2X1_723/B 0.17fF
C50690 PAND2X1_816/O POR2X1_634/A 0.17fF
C50691 POR2X1_68/A POR2X1_632/B 0.03fF
C50692 POR2X1_804/O POR2X1_532/A 0.01fF
C50693 PAND2X1_714/O POR2X1_40/Y 0.03fF
C50694 PAND2X1_658/A POR2X1_60/A 0.08fF
C50695 POR2X1_830/CTRL POR2X1_740/Y 0.00fF
C50696 POR2X1_66/B POR2X1_740/Y 0.07fF
C50697 PAND2X1_116/m4_208_n4# POR2X1_106/Y 0.15fF
C50698 PAND2X1_557/A POR2X1_42/Y 0.03fF
C50699 PAND2X1_227/O POR2X1_394/A 0.07fF
C50700 PAND2X1_36/CTRL2 D_INPUT_6 0.01fF
C50701 POR2X1_497/Y PAND2X1_501/B 0.02fF
C50702 POR2X1_626/CTRL POR2X1_93/A 0.02fF
C50703 PAND2X1_480/B PAND2X1_803/A 0.00fF
C50704 POR2X1_66/A POR2X1_724/A 0.07fF
C50705 POR2X1_83/B PAND2X1_6/A 0.14fF
C50706 POR2X1_81/a_56_344# POR2X1_43/B 0.00fF
C50707 POR2X1_477/B POR2X1_477/A 0.18fF
C50708 POR2X1_260/B POR2X1_569/A 0.14fF
C50709 INPUT_0 PAND2X1_558/a_16_344# 0.02fF
C50710 PAND2X1_287/Y PAND2X1_578/CTRL 0.01fF
C50711 POR2X1_65/A PAND2X1_714/CTRL 0.01fF
C50712 POR2X1_139/A POR2X1_296/B 0.01fF
C50713 POR2X1_188/A POR2X1_740/Y 0.03fF
C50714 PAND2X1_65/B PAND2X1_176/CTRL2 0.01fF
C50715 POR2X1_751/A POR2X1_38/Y 0.06fF
C50716 PAND2X1_859/A POR2X1_55/Y 0.05fF
C50717 POR2X1_652/Y POR2X1_653/B 0.10fF
C50718 PAND2X1_211/A POR2X1_55/Y 0.00fF
C50719 INPUT_1 POR2X1_20/A 0.01fF
C50720 PAND2X1_593/O INPUT_0 0.02fF
C50721 PAND2X1_65/B POR2X1_513/B 0.10fF
C50722 PAND2X1_793/Y PAND2X1_787/Y 0.17fF
C50723 PAND2X1_433/CTRL2 POR2X1_807/A 0.01fF
C50724 POR2X1_237/a_16_28# POR2X1_236/Y 0.05fF
C50725 POR2X1_251/A PAND2X1_190/Y 0.00fF
C50726 PAND2X1_13/CTRL2 POR2X1_222/Y 0.09fF
C50727 POR2X1_66/B PAND2X1_491/CTRL2 0.01fF
C50728 PAND2X1_90/Y PAND2X1_132/CTRL2 0.01fF
C50729 POR2X1_323/Y POR2X1_65/A 0.05fF
C50730 POR2X1_278/Y POR2X1_297/Y 0.00fF
C50731 PAND2X1_739/Y PAND2X1_738/Y 0.05fF
C50732 POR2X1_626/Y PAND2X1_6/A -0.05fF
C50733 PAND2X1_58/A POR2X1_565/a_16_28# 0.03fF
C50734 POR2X1_661/CTRL POR2X1_740/Y 0.00fF
C50735 PAND2X1_67/CTRL POR2X1_507/A 0.04fF
C50736 POR2X1_43/B PAND2X1_849/CTRL2 0.03fF
C50737 POR2X1_60/A POR2X1_73/Y 0.18fF
C50738 POR2X1_16/A PAND2X1_590/CTRL2 0.05fF
C50739 POR2X1_49/Y POR2X1_617/a_76_344# 0.01fF
C50740 POR2X1_48/A PAND2X1_348/CTRL 0.00fF
C50741 POR2X1_404/O POR2X1_35/Y 0.00fF
C50742 POR2X1_222/Y PAND2X1_52/Y 0.03fF
C50743 PAND2X1_382/CTRL PAND2X1_381/Y 0.01fF
C50744 POR2X1_23/Y POR2X1_171/O 0.02fF
C50745 POR2X1_852/A VDD -0.00fF
C50746 POR2X1_72/B PAND2X1_565/O 0.03fF
C50747 POR2X1_753/Y POR2X1_408/Y 0.10fF
C50748 PAND2X1_225/CTRL POR2X1_68/B 0.01fF
C50749 POR2X1_65/A PAND2X1_547/CTRL2 0.03fF
C50750 POR2X1_13/A PAND2X1_804/B 0.09fF
C50751 POR2X1_308/a_16_28# POR2X1_307/Y 0.04fF
C50752 POR2X1_558/B POR2X1_773/B 0.05fF
C50753 POR2X1_265/Y POR2X1_63/Y 0.04fF
C50754 POR2X1_814/A POR2X1_343/O 0.03fF
C50755 POR2X1_383/A POR2X1_646/Y 0.01fF
C50756 PAND2X1_852/B POR2X1_40/Y 0.00fF
C50757 PAND2X1_827/O POR2X1_260/A 0.05fF
C50758 POR2X1_573/a_16_28# POR2X1_404/Y 0.01fF
C50759 POR2X1_96/A PAND2X1_472/B 0.19fF
C50760 POR2X1_186/Y PAND2X1_69/A 5.70fF
C50761 POR2X1_52/A POR2X1_51/A 0.04fF
C50762 PAND2X1_206/a_76_28# POR2X1_293/Y 0.01fF
C50763 POR2X1_436/CTRL POR2X1_209/A 0.00fF
C50764 PAND2X1_771/Y PAND2X1_569/O 0.02fF
C50765 PAND2X1_785/Y POR2X1_293/Y 0.02fF
C50766 PAND2X1_6/Y POR2X1_193/Y 0.06fF
C50767 POR2X1_471/A POR2X1_337/Y 0.07fF
C50768 PAND2X1_420/CTRL POR2X1_510/Y 0.01fF
C50769 POR2X1_829/Y PAND2X1_794/B 0.03fF
C50770 PAND2X1_41/B PAND2X1_177/CTRL2 0.00fF
C50771 POR2X1_14/Y POR2X1_7/A 1.24fF
C50772 VDD PAND2X1_145/CTRL 0.00fF
C50773 POR2X1_311/Y POR2X1_283/A 0.03fF
C50774 POR2X1_413/A INPUT_0 0.12fF
C50775 POR2X1_502/A POR2X1_638/O 0.14fF
C50776 POR2X1_138/O POR2X1_130/A 0.02fF
C50777 POR2X1_722/B POR2X1_502/A 0.00fF
C50778 POR2X1_566/A POR2X1_785/A 0.05fF
C50779 PAND2X1_453/A POR2X1_7/A 0.00fF
C50780 PAND2X1_592/CTRL2 POR2X1_42/Y 0.01fF
C50781 POR2X1_502/A POR2X1_294/B 0.24fF
C50782 PAND2X1_222/CTRL2 PAND2X1_643/A 0.03fF
C50783 POR2X1_603/CTRL2 POR2X1_761/A 0.01fF
C50784 PAND2X1_7/CTRL POR2X1_244/B 0.02fF
C50785 POR2X1_850/A PAND2X1_32/B 0.03fF
C50786 POR2X1_360/A POR2X1_404/Y 0.12fF
C50787 POR2X1_96/A POR2X1_55/Y 1.11fF
C50788 POR2X1_538/CTRL2 POR2X1_566/A 0.01fF
C50789 POR2X1_532/A PAND2X1_52/Y 0.01fF
C50790 PAND2X1_222/A POR2X1_385/Y 0.00fF
C50791 POR2X1_448/Y POR2X1_788/B 0.01fF
C50792 POR2X1_376/B POR2X1_386/CTRL 0.01fF
C50793 POR2X1_13/A PAND2X1_514/Y 0.01fF
C50794 POR2X1_60/A PAND2X1_244/B 0.06fF
C50795 POR2X1_853/a_56_344# POR2X1_776/B 0.00fF
C50796 POR2X1_528/Y POR2X1_748/A 0.46fF
C50797 D_INPUT_0 POR2X1_576/a_16_28# 0.03fF
C50798 POR2X1_56/B PAND2X1_453/O 0.07fF
C50799 POR2X1_78/B PAND2X1_743/CTRL 0.00fF
C50800 POR2X1_247/CTRL POR2X1_294/B 0.01fF
C50801 POR2X1_94/A POR2X1_550/Y 0.35fF
C50802 POR2X1_445/A POR2X1_552/A -0.02fF
C50803 POR2X1_842/CTRL2 POR2X1_737/A 0.01fF
C50804 PAND2X1_287/Y POR2X1_767/CTRL 0.02fF
C50805 POR2X1_304/CTRL2 PAND2X1_454/B 0.01fF
C50806 POR2X1_68/A POR2X1_728/B 0.02fF
C50807 POR2X1_407/A POR2X1_676/Y 0.06fF
C50808 POR2X1_548/O POR2X1_68/B 0.07fF
C50809 PAND2X1_388/CTRL POR2X1_236/Y 0.01fF
C50810 POR2X1_356/A POR2X1_466/a_76_344# 0.09fF
C50811 D_INPUT_3 POR2X1_381/CTRL 0.01fF
C50812 PAND2X1_652/A PAND2X1_191/Y 0.03fF
C50813 POR2X1_79/Y PAND2X1_357/Y 0.03fF
C50814 PAND2X1_96/B PAND2X1_58/O 0.01fF
C50815 POR2X1_588/Y POR2X1_752/Y 0.08fF
C50816 PAND2X1_93/B POR2X1_788/CTRL2 0.03fF
C50817 PAND2X1_23/Y POR2X1_733/A 0.10fF
C50818 POR2X1_55/Y PAND2X1_506/CTRL 0.01fF
C50819 PAND2X1_651/Y PAND2X1_862/B 0.05fF
C50820 POR2X1_66/A POR2X1_620/B 0.07fF
C50821 POR2X1_722/Y POR2X1_513/Y 0.01fF
C50822 POR2X1_305/Y POR2X1_7/B 0.79fF
C50823 POR2X1_510/A POR2X1_857/B 0.03fF
C50824 PAND2X1_739/B VDD 0.00fF
C50825 PAND2X1_140/A POR2X1_107/CTRL 0.01fF
C50826 POR2X1_730/Y POR2X1_330/Y 0.31fF
C50827 POR2X1_288/CTRL PAND2X1_48/A 0.04fF
C50828 POR2X1_665/A VDD -0.00fF
C50829 PAND2X1_48/B POR2X1_782/A 0.06fF
C50830 PAND2X1_661/Y PAND2X1_596/CTRL 0.00fF
C50831 PAND2X1_222/B VDD 0.02fF
C50832 POR2X1_32/A PAND2X1_716/B 0.07fF
C50833 PAND2X1_710/CTRL2 POR2X1_701/Y 0.03fF
C50834 POR2X1_836/a_16_28# POR2X1_192/B 0.05fF
C50835 POR2X1_202/CTRL2 POR2X1_507/A 0.03fF
C50836 POR2X1_461/Y PAND2X1_52/B 0.03fF
C50837 POR2X1_562/O POR2X1_562/B 0.02fF
C50838 PAND2X1_814/O POR2X1_7/B 0.01fF
C50839 POR2X1_406/Y PAND2X1_656/A 0.03fF
C50840 POR2X1_66/B POR2X1_774/A 0.03fF
C50841 POR2X1_480/A POR2X1_568/Y 0.10fF
C50842 POR2X1_730/B POR2X1_730/CTRL 0.01fF
C50843 POR2X1_606/CTRL2 PAND2X1_56/A 0.01fF
C50844 POR2X1_241/B POR2X1_502/Y 0.01fF
C50845 PAND2X1_23/Y POR2X1_124/B 0.02fF
C50846 PAND2X1_824/B POR2X1_186/Y 0.07fF
C50847 PAND2X1_391/O POR2X1_4/Y 0.02fF
C50848 POR2X1_831/CTRL2 POR2X1_717/B 0.01fF
C50849 POR2X1_52/A POR2X1_583/CTRL 0.01fF
C50850 POR2X1_51/A POR2X1_36/a_16_28# 0.02fF
C50851 PAND2X1_81/B PAND2X1_316/CTRL 0.00fF
C50852 PAND2X1_48/B PAND2X1_96/B 1.05fF
C50853 POR2X1_84/CTRL2 POR2X1_532/A 0.01fF
C50854 POR2X1_57/A PAND2X1_114/Y 0.01fF
C50855 PAND2X1_48/B POR2X1_736/CTRL2 0.09fF
C50856 PAND2X1_674/a_76_28# POR2X1_732/B 0.05fF
C50857 POR2X1_673/Y POR2X1_5/Y 0.03fF
C50858 POR2X1_124/O POR2X1_137/Y 0.00fF
C50859 POR2X1_417/a_16_28# POR2X1_372/Y 0.06fF
C50860 POR2X1_41/B PAND2X1_149/A 0.04fF
C50861 PAND2X1_56/Y POR2X1_804/A 0.10fF
C50862 POR2X1_188/A POR2X1_774/A 0.03fF
C50863 POR2X1_119/Y POR2X1_83/B 0.12fF
C50864 PAND2X1_360/Y PAND2X1_349/B 0.01fF
C50865 POR2X1_345/a_16_28# POR2X1_345/A 0.02fF
C50866 POR2X1_192/Y POR2X1_727/O 0.04fF
C50867 POR2X1_57/A PAND2X1_742/B 0.01fF
C50868 PAND2X1_625/CTRL PAND2X1_96/B 0.01fF
C50869 POR2X1_178/Y VDD 0.11fF
C50870 PAND2X1_308/a_76_28# POR2X1_306/Y 0.01fF
C50871 PAND2X1_425/CTRL PAND2X1_18/B 0.01fF
C50872 PAND2X1_94/A POR2X1_410/O 0.29fF
C50873 POR2X1_417/Y PAND2X1_716/B 0.03fF
C50874 PAND2X1_440/CTRL POR2X1_23/Y 0.01fF
C50875 PAND2X1_442/O POR2X1_444/Y 0.04fF
C50876 POR2X1_750/B POR2X1_737/A 0.06fF
C50877 POR2X1_775/CTRL2 PAND2X1_32/B 0.01fF
C50878 PAND2X1_744/CTRL2 POR2X1_532/A 0.03fF
C50879 POR2X1_293/Y PAND2X1_656/A 0.06fF
C50880 PAND2X1_297/CTRL PAND2X1_57/B 0.01fF
C50881 POR2X1_222/Y POR2X1_724/A 0.03fF
C50882 INPUT_0 POR2X1_530/O 0.05fF
C50883 POR2X1_833/CTRL PAND2X1_60/B 0.01fF
C50884 POR2X1_327/Y POR2X1_448/B 0.01fF
C50885 POR2X1_135/a_16_28# POR2X1_32/A 0.00fF
C50886 POR2X1_260/B PAND2X1_72/A 0.20fF
C50887 PAND2X1_127/a_16_344# POR2X1_78/B 0.02fF
C50888 POR2X1_30/CTRL POR2X1_3/A 0.30fF
C50889 POR2X1_55/Y POR2X1_7/A 0.20fF
C50890 PAND2X1_108/CTRL2 POR2X1_646/Y 0.07fF
C50891 PAND2X1_696/O POR2X1_811/B 0.02fF
C50892 POR2X1_532/A POR2X1_771/CTRL2 0.03fF
C50893 POR2X1_85/CTRL POR2X1_83/B 0.01fF
C50894 POR2X1_309/CTRL2 POR2X1_39/B 0.03fF
C50895 POR2X1_462/B POR2X1_532/A 0.11fF
C50896 POR2X1_332/Y PAND2X1_65/B 0.02fF
C50897 POR2X1_207/A POR2X1_195/CTRL2 0.01fF
C50898 POR2X1_65/A POR2X1_110/O 0.03fF
C50899 PAND2X1_55/Y POR2X1_569/A 0.14fF
C50900 POR2X1_532/A D_INPUT_1 0.09fF
C50901 POR2X1_266/A POR2X1_549/B 0.02fF
C50902 PAND2X1_785/CTRL2 POR2X1_91/Y 0.01fF
C50903 POR2X1_635/B PAND2X1_47/m4_208_n4# 0.07fF
C50904 POR2X1_102/Y POR2X1_39/B 8.55fF
C50905 D_GATE_222 POR2X1_854/B 0.10fF
C50906 PAND2X1_117/CTRL POR2X1_260/A 0.01fF
C50907 POR2X1_811/B POR2X1_779/CTRL 0.08fF
C50908 POR2X1_60/A PAND2X1_207/A 0.63fF
C50909 POR2X1_555/B POR2X1_555/O 0.04fF
C50910 POR2X1_832/A POR2X1_435/CTRL 0.01fF
C50911 POR2X1_840/B POR2X1_318/A 0.10fF
C50912 POR2X1_532/A POR2X1_724/A 0.03fF
C50913 PAND2X1_383/O POR2X1_816/A 0.02fF
C50914 POR2X1_327/Y PAND2X1_57/B 0.12fF
C50915 POR2X1_566/A POR2X1_186/B 0.08fF
C50916 POR2X1_317/a_16_28# POR2X1_317/A 0.10fF
C50917 POR2X1_316/Y POR2X1_423/Y 0.04fF
C50918 POR2X1_383/A POR2X1_804/A 0.12fF
C50919 POR2X1_538/CTRL POR2X1_703/A 0.03fF
C50920 PAND2X1_693/CTRL INPUT_1 0.01fF
C50921 POR2X1_72/B PAND2X1_169/O 0.02fF
C50922 PAND2X1_737/B POR2X1_599/A 0.05fF
C50923 POR2X1_13/A POR2X1_75/Y 0.05fF
C50924 PAND2X1_63/Y PAND2X1_63/B 0.04fF
C50925 POR2X1_147/O POR2X1_78/A 0.04fF
C50926 POR2X1_78/B POR2X1_540/Y 0.10fF
C50927 POR2X1_712/A POR2X1_707/Y 0.06fF
C50928 PAND2X1_73/Y POR2X1_715/O 0.02fF
C50929 POR2X1_305/O POR2X1_40/Y 0.02fF
C50930 PAND2X1_533/O POR2X1_532/Y 0.02fF
C50931 POR2X1_49/Y POR2X1_52/a_56_344# 0.00fF
C50932 PAND2X1_850/Y PAND2X1_276/O 0.09fF
C50933 POR2X1_188/A PAND2X1_108/CTRL 0.01fF
C50934 POR2X1_38/Y POR2X1_283/A 0.03fF
C50935 POR2X1_824/Y POR2X1_823/Y 0.14fF
C50936 POR2X1_110/Y PAND2X1_549/O 0.15fF
C50937 POR2X1_38/Y PAND2X1_121/CTRL 0.02fF
C50938 VDD PAND2X1_41/Y 0.10fF
C50939 POR2X1_596/A PAND2X1_765/O 0.02fF
C50940 POR2X1_83/Y PAND2X1_734/B 0.01fF
C50941 POR2X1_814/A PAND2X1_39/B 0.23fF
C50942 POR2X1_567/A POR2X1_502/A 0.05fF
C50943 POR2X1_99/B POR2X1_220/Y 0.03fF
C50944 POR2X1_222/A POR2X1_228/Y 3.11fF
C50945 PAND2X1_95/B PAND2X1_48/A 0.01fF
C50946 POR2X1_343/Y POR2X1_105/Y 0.05fF
C50947 POR2X1_78/B PAND2X1_166/O 0.06fF
C50948 PAND2X1_74/a_76_28# PAND2X1_72/A 0.02fF
C50949 POR2X1_288/A PAND2X1_52/B 0.03fF
C50950 PAND2X1_716/B PAND2X1_302/CTRL 0.01fF
C50951 POR2X1_68/A POR2X1_359/B 0.07fF
C50952 PAND2X1_350/a_76_28# POR2X1_7/A 0.01fF
C50953 POR2X1_567/A POR2X1_464/Y 0.05fF
C50954 PAND2X1_631/A POR2X1_293/Y 0.04fF
C50955 PAND2X1_732/A POR2X1_152/Y 0.00fF
C50956 POR2X1_92/CTRL POR2X1_8/Y 0.01fF
C50957 POR2X1_840/Y POR2X1_307/Y 0.01fF
C50958 PAND2X1_310/CTRL2 POR2X1_501/B 0.01fF
C50959 POR2X1_840/B POR2X1_574/Y 0.05fF
C50960 POR2X1_158/Y PAND2X1_713/B 0.00fF
C50961 POR2X1_184/Y PAND2X1_716/B 0.12fF
C50962 POR2X1_617/Y PAND2X1_6/A 0.03fF
C50963 POR2X1_205/A POR2X1_244/Y 0.07fF
C50964 PAND2X1_63/B POR2X1_376/CTRL2 0.01fF
C50965 PAND2X1_833/a_16_344# POR2X1_77/Y 0.02fF
C50966 PAND2X1_357/Y PAND2X1_730/A 0.03fF
C50967 PAND2X1_785/CTRL2 POR2X1_109/Y 0.03fF
C50968 PAND2X1_150/O POR2X1_186/B 0.01fF
C50969 INPUT_1 POR2X1_283/A 0.10fF
C50970 PAND2X1_408/O PAND2X1_26/A 0.00fF
C50971 PAND2X1_63/B POR2X1_260/A 0.12fF
C50972 POR2X1_727/CTRL2 POR2X1_353/A 0.00fF
C50973 PAND2X1_779/O POR2X1_90/Y 0.04fF
C50974 PAND2X1_865/Y PAND2X1_675/A 0.07fF
C50975 PAND2X1_714/A POR2X1_166/Y 0.12fF
C50976 PAND2X1_26/CTRL2 PAND2X1_18/B 0.01fF
C50977 PAND2X1_79/Y PAND2X1_527/CTRL 0.08fF
C50978 POR2X1_363/A POR2X1_359/Y 0.02fF
C50979 POR2X1_861/A POR2X1_861/a_16_28# 0.01fF
C50980 PAND2X1_290/CTRL PAND2X1_55/Y 0.01fF
C50981 INPUT_1 PAND2X1_528/O 0.01fF
C50982 POR2X1_518/O POR2X1_519/Y 0.09fF
C50983 POR2X1_518/CTRL POR2X1_518/Y 0.02fF
C50984 PAND2X1_630/CTRL PAND2X1_508/B 0.01fF
C50985 PAND2X1_474/Y PAND2X1_332/Y 0.97fF
C50986 POR2X1_532/A POR2X1_620/B 0.68fF
C50987 PAND2X1_48/B POR2X1_342/B 0.02fF
C50988 POR2X1_283/A POR2X1_153/Y 0.05fF
C50989 POR2X1_49/Y PAND2X1_147/O 0.02fF
C50990 POR2X1_648/Y POR2X1_646/Y 0.06fF
C50991 POR2X1_692/CTRL POR2X1_485/Y 0.01fF
C50992 POR2X1_42/a_56_344# POR2X1_4/Y 0.00fF
C50993 POR2X1_13/A PAND2X1_332/Y 0.06fF
C50994 POR2X1_23/Y POR2X1_271/B 0.03fF
C50995 POR2X1_74/CTRL2 POR2X1_271/A 0.04fF
C50996 PAND2X1_501/CTRL PAND2X1_575/A 0.01fF
C50997 POR2X1_334/Y POR2X1_97/CTRL2 0.05fF
C50998 POR2X1_539/A POR2X1_370/O 0.08fF
C50999 PAND2X1_20/A POR2X1_814/A 0.18fF
C51000 POR2X1_508/a_76_344# POR2X1_568/B 0.03fF
C51001 POR2X1_44/CTRL PAND2X1_635/Y 0.01fF
C51002 POR2X1_137/B POR2X1_66/A 0.07fF
C51003 POR2X1_16/A POR2X1_394/A 0.33fF
C51004 POR2X1_532/A PAND2X1_134/O 0.16fF
C51005 POR2X1_531/Y POR2X1_39/B 0.00fF
C51006 POR2X1_20/B POR2X1_409/B 0.03fF
C51007 PAND2X1_483/CTRL2 PAND2X1_508/Y 0.00fF
C51008 PAND2X1_845/CTRL POR2X1_39/B 0.00fF
C51009 POR2X1_484/Y POR2X1_484/O 0.01fF
C51010 POR2X1_789/Y PAND2X1_52/B 0.04fF
C51011 PAND2X1_55/Y PAND2X1_72/A 0.13fF
C51012 PAND2X1_346/Y PAND2X1_345/Y 0.06fF
C51013 PAND2X1_462/O POR2X1_416/Y 0.02fF
C51014 POR2X1_9/Y PAND2X1_340/CTRL 0.07fF
C51015 INPUT_3 POR2X1_66/A 0.02fF
C51016 POR2X1_677/Y PAND2X1_499/Y 0.03fF
C51017 POR2X1_65/A POR2X1_292/O 0.02fF
C51018 POR2X1_96/A PAND2X1_862/m4_208_n4# 0.01fF
C51019 POR2X1_416/B POR2X1_747/Y 0.01fF
C51020 PAND2X1_857/A PAND2X1_857/O -0.00fF
C51021 POR2X1_709/a_16_28# POR2X1_709/B 0.08fF
C51022 POR2X1_48/A PAND2X1_340/B 0.03fF
C51023 POR2X1_821/Y POR2X1_39/B 0.01fF
C51024 POR2X1_557/A POR2X1_571/Y 0.03fF
C51025 POR2X1_814/B POR2X1_814/A 0.11fF
C51026 POR2X1_452/CTRL POR2X1_121/B 0.08fF
C51027 POR2X1_633/A POR2X1_633/a_76_344# 0.01fF
C51028 POR2X1_137/B POR2X1_634/CTRL2 0.00fF
C51029 POR2X1_77/a_76_344# POR2X1_48/A 0.01fF
C51030 PAND2X1_418/CTRL PAND2X1_41/B 0.10fF
C51031 PAND2X1_60/B POR2X1_716/CTRL2 0.09fF
C51032 POR2X1_847/A POR2X1_20/B 0.01fF
C51033 POR2X1_731/O PAND2X1_52/B 0.02fF
C51034 PAND2X1_69/A POR2X1_717/B 0.08fF
C51035 PAND2X1_93/B POR2X1_66/A 0.49fF
C51036 PAND2X1_860/A POR2X1_42/Y 0.06fF
C51037 POR2X1_407/Y PAND2X1_72/A 0.03fF
C51038 POR2X1_814/A POR2X1_325/A 0.03fF
C51039 POR2X1_705/B POR2X1_734/A 0.05fF
C51040 PAND2X1_717/A POR2X1_236/Y 0.03fF
C51041 POR2X1_359/CTRL POR2X1_363/A 0.04fF
C51042 POR2X1_825/Y PAND2X1_334/CTRL2 0.00fF
C51043 D_INPUT_5 PAND2X1_58/A 0.02fF
C51044 POR2X1_646/B POR2X1_480/A 0.00fF
C51045 POR2X1_600/Y POR2X1_601/a_16_28# 0.02fF
C51046 POR2X1_96/B POR2X1_77/Y 0.03fF
C51047 PAND2X1_647/B POR2X1_612/Y 0.14fF
C51048 PAND2X1_761/CTRL POR2X1_750/B 0.01fF
C51049 PAND2X1_617/CTRL2 VDD 0.00fF
C51050 POR2X1_500/A POR2X1_341/A 0.07fF
C51051 POR2X1_84/A POR2X1_590/A 0.03fF
C51052 PAND2X1_3/A PAND2X1_36/CTRL 0.01fF
C51053 POR2X1_257/A PAND2X1_390/Y 0.07fF
C51054 POR2X1_416/B PAND2X1_514/CTRL2 0.01fF
C51055 PAND2X1_69/A PAND2X1_146/CTRL 0.01fF
C51056 POR2X1_567/m4_208_n4# POR2X1_854/B 0.06fF
C51057 PAND2X1_23/Y PAND2X1_438/O 0.02fF
C51058 POR2X1_60/A POR2X1_813/m4_208_n4# 0.09fF
C51059 PAND2X1_41/O PAND2X1_41/B 0.01fF
C51060 PAND2X1_691/O POR2X1_689/Y 0.02fF
C51061 PAND2X1_850/Y POR2X1_129/Y 0.19fF
C51062 PAND2X1_357/O PAND2X1_353/Y 0.08fF
C51063 PAND2X1_39/B POR2X1_852/B 0.20fF
C51064 POR2X1_814/A POR2X1_513/B 0.06fF
C51065 PAND2X1_497/a_76_28# POR2X1_78/A 0.02fF
C51066 PAND2X1_446/Y POR2X1_376/B 0.08fF
C51067 POR2X1_48/A POR2X1_102/Y 3.44fF
C51068 PAND2X1_9/Y POR2X1_5/Y 0.06fF
C51069 PAND2X1_807/B PAND2X1_805/Y 0.00fF
C51070 POR2X1_78/A POR2X1_66/A 11.30fF
C51071 POR2X1_20/B PAND2X1_721/a_76_28# 0.01fF
C51072 POR2X1_72/Y POR2X1_329/A 0.03fF
C51073 POR2X1_416/B PAND2X1_537/O 0.05fF
C51074 POR2X1_20/B POR2X1_272/Y 0.03fF
C51075 POR2X1_567/A POR2X1_188/Y 0.03fF
C51076 POR2X1_88/a_16_28# POR2X1_69/A 0.02fF
C51077 POR2X1_257/A POR2X1_697/CTRL 0.01fF
C51078 POR2X1_456/B POR2X1_715/CTRL 0.01fF
C51079 POR2X1_520/m4_208_n4# PAND2X1_52/B 0.09fF
C51080 PAND2X1_434/O POR2X1_72/B 0.02fF
C51081 POR2X1_202/A POR2X1_402/O 0.03fF
C51082 PAND2X1_412/O POR2X1_260/B 0.02fF
C51083 PAND2X1_416/CTRL2 VDD -0.00fF
C51084 POR2X1_362/Y POR2X1_590/A 0.01fF
C51085 POR2X1_285/Y POR2X1_590/A 0.01fF
C51086 POR2X1_20/B PAND2X1_351/Y 0.02fF
C51087 POR2X1_218/Y POR2X1_330/Y 0.10fF
C51088 PAND2X1_791/CTRL VDD -0.00fF
C51089 POR2X1_814/A POR2X1_467/CTRL2 0.02fF
C51090 POR2X1_696/CTRL POR2X1_32/A 0.01fF
C51091 POR2X1_805/O POR2X1_805/B 0.03fF
C51092 POR2X1_78/B POR2X1_445/A 0.23fF
C51093 PAND2X1_644/CTRL POR2X1_683/Y 0.00fF
C51094 POR2X1_326/O POR2X1_568/A 0.01fF
C51095 POR2X1_669/B POR2X1_69/A 0.30fF
C51096 POR2X1_650/A POR2X1_493/A 0.03fF
C51097 POR2X1_65/A PAND2X1_640/B 0.42fF
C51098 POR2X1_333/Y PAND2X1_72/A 0.05fF
C51099 PAND2X1_73/Y POR2X1_780/CTRL2 0.01fF
C51100 POR2X1_322/CTRL POR2X1_441/Y 0.01fF
C51101 POR2X1_490/Y PAND2X1_741/B 0.03fF
C51102 POR2X1_260/B POR2X1_285/O 0.02fF
C51103 PAND2X1_699/CTRL2 PAND2X1_6/A 0.01fF
C51104 PAND2X1_20/A POR2X1_34/Y 0.96fF
C51105 POR2X1_16/A POR2X1_91/CTRL 0.01fF
C51106 PAND2X1_288/O POR2X1_7/B 0.01fF
C51107 PAND2X1_205/Y POR2X1_32/A 0.03fF
C51108 POR2X1_302/B PAND2X1_279/CTRL2 0.01fF
C51109 PAND2X1_808/Y PAND2X1_580/a_76_28# 0.01fF
C51110 POR2X1_60/A PAND2X1_541/CTRL2 0.00fF
C51111 POR2X1_556/A POR2X1_556/a_16_28# 0.04fF
C51112 POR2X1_634/A PAND2X1_428/O 0.17fF
C51113 PAND2X1_447/O POR2X1_90/Y 0.02fF
C51114 PAND2X1_57/B POR2X1_644/Y 0.06fF
C51115 PAND2X1_267/Y POR2X1_46/Y 0.13fF
C51116 POR2X1_302/A PAND2X1_39/B 0.02fF
C51117 POR2X1_16/A POR2X1_16/a_16_28# 0.01fF
C51118 POR2X1_786/A POR2X1_266/O 0.02fF
C51119 PAND2X1_485/O PAND2X1_57/B 0.08fF
C51120 POR2X1_43/B POR2X1_442/O 0.01fF
C51121 PAND2X1_234/CTRL2 POR2X1_260/A 0.03fF
C51122 POR2X1_329/A PAND2X1_349/A 0.03fF
C51123 POR2X1_499/A POR2X1_68/B 0.03fF
C51124 POR2X1_490/CTRL2 POR2X1_73/Y 0.01fF
C51125 POR2X1_137/B POR2X1_532/A 0.10fF
C51126 POR2X1_32/A PAND2X1_151/CTRL 0.03fF
C51127 POR2X1_416/A POR2X1_293/Y 0.05fF
C51128 PAND2X1_206/A PAND2X1_6/A 0.00fF
C51129 PAND2X1_90/A POR2X1_28/O 0.02fF
C51130 PAND2X1_657/CTRL2 PAND2X1_659/B 0.00fF
C51131 POR2X1_493/A POR2X1_294/B 0.05fF
C51132 POR2X1_829/O POR2X1_829/Y 0.02fF
C51133 POR2X1_198/CTRL PAND2X1_93/B 0.01fF
C51134 POR2X1_60/A PAND2X1_804/A 0.01fF
C51135 POR2X1_697/CTRL2 POR2X1_40/Y 0.01fF
C51136 PAND2X1_93/B POR2X1_222/Y 0.03fF
C51137 PAND2X1_200/CTRL VDD -0.00fF
C51138 POR2X1_65/A POR2X1_295/a_16_28# 0.02fF
C51139 PAND2X1_614/O POR2X1_5/Y 0.17fF
C51140 PAND2X1_631/A PAND2X1_242/Y 0.05fF
C51141 PAND2X1_20/A POR2X1_401/B 0.02fF
C51142 PAND2X1_94/A POR2X1_624/B 0.26fF
C51143 POR2X1_60/A PAND2X1_785/Y 0.06fF
C51144 POR2X1_355/a_16_28# POR2X1_355/A 0.05fF
C51145 POR2X1_270/CTRL POR2X1_445/A 0.02fF
C51146 POR2X1_657/Y POR2X1_222/A 0.03fF
C51147 POR2X1_150/Y PAND2X1_717/Y 0.21fF
C51148 D_GATE_662 POR2X1_220/B 0.07fF
C51149 POR2X1_656/O POR2X1_733/A 0.24fF
C51150 POR2X1_604/Y POR2X1_7/B 0.10fF
C51151 PAND2X1_793/Y PAND2X1_78/CTRL2 0.01fF
C51152 POR2X1_417/Y PAND2X1_151/CTRL 0.01fF
C51153 POR2X1_66/B POR2X1_445/CTRL2 0.11fF
C51154 PAND2X1_477/B PAND2X1_477/a_16_344# 0.03fF
C51155 POR2X1_777/B VDD 3.36fF
C51156 POR2X1_482/CTRL2 PAND2X1_6/A 0.13fF
C51157 PAND2X1_845/O POR2X1_23/Y 0.02fF
C51158 POR2X1_236/CTRL2 POR2X1_5/Y 0.03fF
C51159 POR2X1_241/B POR2X1_785/A 0.03fF
C51160 PAND2X1_485/CTRL PAND2X1_69/A 0.01fF
C51161 POR2X1_194/A VDD -0.00fF
C51162 POR2X1_813/O PAND2X1_63/B 0.02fF
C51163 PAND2X1_192/Y PAND2X1_739/CTRL2 0.01fF
C51164 PAND2X1_685/O POR2X1_32/A 0.02fF
C51165 POR2X1_345/A POR2X1_244/B 0.02fF
C51166 POR2X1_16/A POR2X1_679/O 0.01fF
C51167 POR2X1_660/A VDD 0.13fF
C51168 PAND2X1_319/B POR2X1_298/O 0.01fF
C51169 POR2X1_311/Y POR2X1_55/Y 14.12fF
C51170 POR2X1_102/Y PAND2X1_197/Y 0.06fF
C51171 PAND2X1_93/B POR2X1_532/A 1.58fF
C51172 POR2X1_413/A POR2X1_102/Y 0.03fF
C51173 PAND2X1_811/O PAND2X1_805/A 0.02fF
C51174 POR2X1_655/A POR2X1_537/B 0.01fF
C51175 INPUT_0 POR2X1_595/Y 0.03fF
C51176 PAND2X1_48/B PAND2X1_394/a_16_344# 0.01fF
C51177 POR2X1_763/A POR2X1_763/a_16_28# 0.05fF
C51178 POR2X1_196/O PAND2X1_56/Y 0.04fF
C51179 POR2X1_685/A POR2X1_676/O 0.01fF
C51180 POR2X1_790/A POR2X1_29/A 7.65fF
C51181 POR2X1_60/CTRL D_INPUT_0 0.07fF
C51182 PAND2X1_540/CTRL2 PAND2X1_553/B 0.05fF
C51183 PAND2X1_65/B VDD 3.06fF
C51184 PAND2X1_391/O POR2X1_816/A 0.02fF
C51185 POR2X1_13/A PAND2X1_562/B 0.07fF
C51186 POR2X1_78/B POR2X1_786/O 0.03fF
C51187 PAND2X1_50/CTRL VDD 0.00fF
C51188 POR2X1_417/Y PAND2X1_775/a_16_344# 0.03fF
C51189 PAND2X1_204/a_16_344# PAND2X1_84/Y 0.05fF
C51190 POR2X1_68/A PAND2X1_394/CTRL 0.01fF
C51191 PAND2X1_723/Y VDD 0.07fF
C51192 POR2X1_14/O POR2X1_68/B 0.01fF
C51193 PAND2X1_755/O PAND2X1_90/Y 0.09fF
C51194 POR2X1_248/A POR2X1_283/A 0.01fF
C51195 POR2X1_237/Y POR2X1_83/B 0.01fF
C51196 PAND2X1_347/Y VDD 0.31fF
C51197 PAND2X1_236/O PAND2X1_8/Y 0.03fF
C51198 POR2X1_65/A POR2X1_7/B 0.15fF
C51199 PAND2X1_137/Y PAND2X1_768/Y 0.04fF
C51200 PAND2X1_362/A PAND2X1_362/O 0.01fF
C51201 GATE_479 POR2X1_763/Y 0.07fF
C51202 POR2X1_57/A PAND2X1_220/A 0.01fF
C51203 PAND2X1_656/B PAND2X1_656/A 0.02fF
C51204 PAND2X1_20/A POR2X1_139/O 0.01fF
C51205 POR2X1_96/A POR2X1_511/Y 0.12fF
C51206 PAND2X1_857/O POR2X1_329/A 0.03fF
C51207 PAND2X1_655/B POR2X1_32/A 0.01fF
C51208 PAND2X1_119/O POR2X1_78/A 0.01fF
C51209 POR2X1_9/Y POR2X1_39/B 0.42fF
C51210 POR2X1_68/A POR2X1_330/Y 0.17fF
C51211 POR2X1_260/Y POR2X1_814/B 0.01fF
C51212 POR2X1_78/A POR2X1_532/A 0.36fF
C51213 POR2X1_174/A POR2X1_190/O 0.07fF
C51214 POR2X1_41/B POR2X1_236/Y 0.22fF
C51215 PAND2X1_805/O PAND2X1_793/Y 0.05fF
C51216 PAND2X1_838/B PAND2X1_560/B 0.02fF
C51217 PAND2X1_576/B PAND2X1_723/A 0.15fF
C51218 POR2X1_447/B POR2X1_66/O 0.06fF
C51219 POR2X1_273/CTRL2 POR2X1_153/Y 0.00fF
C51220 POR2X1_296/B PAND2X1_505/O 0.15fF
C51221 POR2X1_116/a_16_28# POR2X1_114/Y 0.07fF
C51222 PAND2X1_139/B PAND2X1_137/Y 0.06fF
C51223 POR2X1_14/Y POR2X1_38/Y 0.03fF
C51224 POR2X1_57/A PAND2X1_296/O 0.01fF
C51225 POR2X1_376/B PAND2X1_254/a_16_344# 0.02fF
C51226 POR2X1_317/CTRL PAND2X1_90/Y 0.01fF
C51227 POR2X1_614/A PAND2X1_262/CTRL2 0.05fF
C51228 POR2X1_548/O PAND2X1_90/A 0.01fF
C51229 POR2X1_178/CTRL2 PAND2X1_562/B 0.05fF
C51230 PAND2X1_715/CTRL2 POR2X1_293/Y 0.01fF
C51231 POR2X1_444/CTRL2 POR2X1_191/Y 0.01fF
C51232 POR2X1_444/O POR2X1_192/B 0.06fF
C51233 POR2X1_23/Y PAND2X1_160/a_16_344# 0.02fF
C51234 POR2X1_692/CTRL PAND2X1_726/B 0.04fF
C51235 POR2X1_141/Y POR2X1_112/Y 0.70fF
C51236 PAND2X1_857/A POR2X1_32/A 0.03fF
C51237 PAND2X1_46/CTRL2 POR2X1_68/B 0.00fF
C51238 PAND2X1_65/B POR2X1_741/Y 0.03fF
C51239 POR2X1_597/A INPUT_0 0.05fF
C51240 POR2X1_57/A PAND2X1_718/Y 0.00fF
C51241 PAND2X1_55/Y POR2X1_285/O 0.03fF
C51242 POR2X1_502/A PAND2X1_386/Y 0.01fF
C51243 POR2X1_777/B PAND2X1_32/B 0.09fF
C51244 POR2X1_451/a_16_28# POR2X1_451/A 0.02fF
C51245 POR2X1_78/A PAND2X1_424/a_76_28# 0.02fF
C51246 POR2X1_56/B POR2X1_516/B 0.00fF
C51247 PAND2X1_641/Y POR2X1_23/Y 0.55fF
C51248 PAND2X1_99/O PAND2X1_333/Y 0.02fF
C51249 POR2X1_57/A PAND2X1_360/O 0.01fF
C51250 PAND2X1_653/CTRL POR2X1_760/A 0.02fF
C51251 POR2X1_68/A PAND2X1_525/a_16_344# 0.02fF
C51252 POR2X1_174/A POR2X1_569/A 0.45fF
C51253 POR2X1_46/Y POR2X1_531/CTRL 0.08fF
C51254 PAND2X1_805/A POR2X1_759/Y 0.02fF
C51255 POR2X1_244/B POR2X1_340/CTRL 0.01fF
C51256 POR2X1_244/B POR2X1_205/Y 0.03fF
C51257 POR2X1_60/A PAND2X1_656/A 0.06fF
C51258 POR2X1_652/CTRL2 POR2X1_480/A 0.03fF
C51259 PAND2X1_159/a_76_28# POR2X1_68/B 0.07fF
C51260 POR2X1_62/Y PAND2X1_340/B 0.06fF
C51261 POR2X1_565/B POR2X1_502/A 0.05fF
C51262 PAND2X1_243/B PAND2X1_35/Y 0.00fF
C51263 PAND2X1_360/CTRL PAND2X1_843/Y 0.01fF
C51264 PAND2X1_213/Y POR2X1_40/Y 0.03fF
C51265 D_INPUT_2 VDD 0.78fF
C51266 POR2X1_234/Y POR2X1_293/Y 0.09fF
C51267 GATE_479 POR2X1_73/Y 0.03fF
C51268 PAND2X1_55/Y POR2X1_244/B 0.03fF
C51269 POR2X1_655/A PAND2X1_48/A 0.03fF
C51270 POR2X1_614/A POR2X1_801/A 0.01fF
C51271 PAND2X1_41/B POR2X1_206/O 0.02fF
C51272 POR2X1_643/Y POR2X1_294/A 0.02fF
C51273 PAND2X1_853/CTRL VDD 0.00fF
C51274 PAND2X1_226/CTRL2 POR2X1_578/Y 0.03fF
C51275 POR2X1_16/A POR2X1_669/B 0.51fF
C51276 POR2X1_748/A POR2X1_245/Y 0.07fF
C51277 POR2X1_834/Y POR2X1_296/B 0.10fF
C51278 PAND2X1_65/B PAND2X1_32/B 0.23fF
C51279 POR2X1_174/A POR2X1_570/Y 0.07fF
C51280 POR2X1_383/A POR2X1_794/B 0.02fF
C51281 PAND2X1_48/B POR2X1_708/B 0.01fF
C51282 PAND2X1_14/CTRL D_INPUT_1 0.01fF
C51283 POR2X1_537/Y POR2X1_260/B 0.05fF
C51284 POR2X1_775/A POR2X1_220/Y 0.07fF
C51285 PAND2X1_228/CTRL PAND2X1_364/B 0.03fF
C51286 POR2X1_211/CTRL VDD -0.00fF
C51287 PAND2X1_90/Y POR2X1_540/CTRL2 0.01fF
C51288 PAND2X1_61/Y PAND2X1_560/O 0.03fF
C51289 POR2X1_102/Y POR2X1_530/O 0.01fF
C51290 POR2X1_485/O POR2X1_73/Y 0.01fF
C51291 POR2X1_684/CTRL POR2X1_42/Y 0.01fF
C51292 POR2X1_346/B PAND2X1_626/CTRL2 0.00fF
C51293 PAND2X1_541/CTRL POR2X1_7/A 0.01fF
C51294 POR2X1_57/A POR2X1_106/Y 0.03fF
C51295 POR2X1_78/B PAND2X1_63/Y 0.03fF
C51296 POR2X1_790/A POR2X1_546/A 0.03fF
C51297 POR2X1_326/a_16_28# POR2X1_220/B 0.00fF
C51298 INPUT_1 POR2X1_14/Y 15.27fF
C51299 POR2X1_294/B POR2X1_725/a_16_28# 0.01fF
C51300 PAND2X1_736/A PAND2X1_592/Y 0.07fF
C51301 POR2X1_614/A POR2X1_809/B 0.04fF
C51302 POR2X1_333/a_16_28# POR2X1_174/B -0.00fF
C51303 POR2X1_66/B POR2X1_750/Y 0.01fF
C51304 POR2X1_302/Y POR2X1_513/Y 0.03fF
C51305 POR2X1_407/A POR2X1_502/A 0.03fF
C51306 POR2X1_407/A POR2X1_783/A 0.09fF
C51307 POR2X1_41/B POR2X1_152/CTRL 0.03fF
C51308 POR2X1_28/CTRL2 POR2X1_4/Y 0.06fF
C51309 POR2X1_41/B PAND2X1_850/O 0.01fF
C51310 POR2X1_43/B PAND2X1_735/a_76_28# 0.01fF
C51311 PAND2X1_65/B PAND2X1_312/O 0.00fF
C51312 PAND2X1_23/Y POR2X1_477/A 0.03fF
C51313 PAND2X1_492/O POR2X1_532/A 0.10fF
C51314 PAND2X1_84/CTRL2 POR2X1_91/Y 0.01fF
C51315 POR2X1_362/B PAND2X1_60/B 0.06fF
C51316 PAND2X1_95/B PAND2X1_95/O 0.01fF
C51317 PAND2X1_50/O INPUT_6 0.15fF
C51318 POR2X1_278/Y PAND2X1_734/O 0.23fF
C51319 PAND2X1_241/CTRL2 POR2X1_237/Y 0.01fF
C51320 POR2X1_60/A PAND2X1_348/A 0.07fF
C51321 POR2X1_241/B POR2X1_186/B 0.06fF
C51322 POR2X1_57/A PAND2X1_580/B 0.03fF
C51323 POR2X1_220/Y POR2X1_112/Y 0.03fF
C51324 PAND2X1_661/B POR2X1_13/A 2.75fF
C51325 POR2X1_391/A POR2X1_391/a_16_28# -0.00fF
C51326 POR2X1_142/CTRL2 POR2X1_394/A 0.05fF
C51327 POR2X1_13/A PAND2X1_643/Y 0.03fF
C51328 PAND2X1_341/A POR2X1_88/Y 0.01fF
C51329 POR2X1_558/CTRL POR2X1_264/Y 0.01fF
C51330 POR2X1_41/B POR2X1_229/CTRL 0.00fF
C51331 POR2X1_345/CTRL2 POR2X1_330/Y 0.03fF
C51332 PAND2X1_402/B POR2X1_5/Y 0.01fF
C51333 POR2X1_14/Y POR2X1_153/Y 0.32fF
C51334 PAND2X1_516/a_16_344# POR2X1_513/Y 0.02fF
C51335 POR2X1_123/A PAND2X1_90/Y 0.03fF
C51336 POR2X1_722/A POR2X1_811/B 0.72fF
C51337 POR2X1_511/Y POR2X1_7/A 0.07fF
C51338 PAND2X1_453/A POR2X1_153/Y 0.03fF
C51339 POR2X1_846/B POR2X1_43/B 0.02fF
C51340 PAND2X1_472/B POR2X1_38/Y 0.07fF
C51341 POR2X1_536/O POR2X1_250/A 0.01fF
C51342 POR2X1_52/A POR2X1_131/O 0.01fF
C51343 POR2X1_391/A POR2X1_260/A 0.03fF
C51344 POR2X1_76/Y POR2X1_541/a_56_344# 0.00fF
C51345 POR2X1_650/A POR2X1_276/Y 0.03fF
C51346 POR2X1_158/Y POR2X1_257/A 0.04fF
C51347 POR2X1_369/a_76_344# POR2X1_60/A 0.03fF
C51348 PAND2X1_386/CTRL POR2X1_260/A 0.01fF
C51349 POR2X1_231/O PAND2X1_32/B 0.01fF
C51350 POR2X1_96/Y PAND2X1_61/CTRL 0.09fF
C51351 POR2X1_60/A POR2X1_300/Y 0.09fF
C51352 POR2X1_132/Y POR2X1_7/B 0.01fF
C51353 POR2X1_62/Y POR2X1_102/Y 0.06fF
C51354 POR2X1_379/Y PAND2X1_20/A 0.00fF
C51355 POR2X1_46/Y POR2X1_526/Y 0.00fF
C51356 PAND2X1_108/O POR2X1_383/A 0.05fF
C51357 POR2X1_316/CTRL PAND2X1_390/Y 0.01fF
C51358 POR2X1_334/B POR2X1_124/B 0.07fF
C51359 PAND2X1_65/B PAND2X1_253/O 0.17fF
C51360 PAND2X1_289/O PAND2X1_52/B 0.02fF
C51361 PAND2X1_742/B POR2X1_594/A 0.02fF
C51362 POR2X1_296/B POR2X1_722/a_16_28# 0.21fF
C51363 POR2X1_55/Y PAND2X1_509/CTRL2 0.15fF
C51364 POR2X1_68/B PAND2X1_132/O 0.01fF
C51365 POR2X1_457/Y POR2X1_458/Y 0.03fF
C51366 PAND2X1_212/B PAND2X1_352/CTRL 0.01fF
C51367 PAND2X1_65/B POR2X1_673/Y 0.03fF
C51368 POR2X1_285/B POR2X1_260/B 0.00fF
C51369 PAND2X1_209/A PAND2X1_162/CTRL2 0.09fF
C51370 POR2X1_220/Y POR2X1_162/Y 0.02fF
C51371 POR2X1_38/Y POR2X1_55/Y 0.13fF
C51372 POR2X1_347/A POR2X1_402/O 0.01fF
C51373 PAND2X1_491/O POR2X1_264/Y 0.02fF
C51374 POR2X1_174/B POR2X1_508/B 0.03fF
C51375 POR2X1_407/A POR2X1_114/O 0.00fF
C51376 POR2X1_544/A POR2X1_180/A 0.19fF
C51377 POR2X1_72/B PAND2X1_508/Y 0.03fF
C51378 VDD PAND2X1_346/Y 0.30fF
C51379 POR2X1_795/B POR2X1_570/B 0.19fF
C51380 POR2X1_22/A POR2X1_36/CTRL2 0.01fF
C51381 POR2X1_13/A PAND2X1_510/B 0.03fF
C51382 PAND2X1_354/A PAND2X1_345/Y 0.01fF
C51383 PAND2X1_48/CTRL2 POR2X1_260/A 0.01fF
C51384 POR2X1_78/B POR2X1_260/A 0.15fF
C51385 PAND2X1_632/O VDD 0.00fF
C51386 POR2X1_751/Y POR2X1_5/Y 0.05fF
C51387 POR2X1_66/B POR2X1_447/B 0.10fF
C51388 PAND2X1_566/Y POR2X1_90/Y 0.04fF
C51389 POR2X1_861/O POR2X1_865/B 0.03fF
C51390 POR2X1_12/CTRL2 POR2X1_3/B 0.00fF
C51391 POR2X1_119/Y PAND2X1_444/Y 0.01fF
C51392 PAND2X1_631/A POR2X1_60/A 2.10fF
C51393 POR2X1_859/A POR2X1_750/Y 0.03fF
C51394 PAND2X1_308/Y POR2X1_236/Y 0.09fF
C51395 POR2X1_48/A POR2X1_320/Y 0.01fF
C51396 PAND2X1_17/m4_208_n4# POR2X1_581/m4_208_n4# 0.13fF
C51397 PAND2X1_717/Y PAND2X1_364/B 0.07fF
C51398 POR2X1_294/B POR2X1_510/Y 1.24fF
C51399 POR2X1_523/Y POR2X1_844/CTRL 0.01fF
C51400 PAND2X1_736/CTRL PAND2X1_853/B 0.11fF
C51401 POR2X1_614/A POR2X1_156/B 0.00fF
C51402 POR2X1_510/A POR2X1_532/A 0.01fF
C51403 PAND2X1_6/Y POR2X1_140/CTRL2 0.08fF
C51404 D_GATE_222 PAND2X1_173/CTRL2 0.03fF
C51405 POR2X1_407/m4_208_n4# PAND2X1_597/m4_208_n4# 0.13fF
C51406 POR2X1_83/B PAND2X1_326/B 0.03fF
C51407 POR2X1_357/O POR2X1_353/Y 0.03fF
C51408 PAND2X1_524/CTRL2 POR2X1_456/B 0.01fF
C51409 POR2X1_57/A PAND2X1_337/A 0.01fF
C51410 POR2X1_48/O POR2X1_153/Y 0.04fF
C51411 PAND2X1_79/Y POR2X1_844/B 0.91fF
C51412 PAND2X1_55/Y POR2X1_736/a_16_28# 0.02fF
C51413 INPUT_1 PAND2X1_472/B 0.09fF
C51414 PAND2X1_658/A PAND2X1_175/B 0.03fF
C51415 POR2X1_205/A POR2X1_205/a_16_28# 0.03fF
C51416 PAND2X1_90/Y PAND2X1_384/a_16_344# 0.02fF
C51417 POR2X1_541/CTRL PAND2X1_32/B 0.01fF
C51418 POR2X1_407/Y PAND2X1_743/a_16_344# 0.01fF
C51419 POR2X1_65/a_16_28# POR2X1_9/Y 0.02fF
C51420 PAND2X1_61/Y PAND2X1_338/CTRL2 0.01fF
C51421 POR2X1_303/CTRL POR2X1_814/B 0.01fF
C51422 PAND2X1_139/B PAND2X1_853/B 0.01fF
C51423 POR2X1_170/B POR2X1_169/O 0.02fF
C51424 POR2X1_786/Y POR2X1_702/CTRL 0.06fF
C51425 PAND2X1_735/O POR2X1_153/Y 0.11fF
C51426 POR2X1_529/O PAND2X1_510/B 0.02fF
C51427 POR2X1_157/O POR2X1_158/B 0.01fF
C51428 POR2X1_110/Y PAND2X1_76/Y 0.03fF
C51429 POR2X1_294/B POR2X1_276/Y 0.05fF
C51430 PAND2X1_410/CTRL POR2X1_234/A 0.01fF
C51431 INPUT_1 PAND2X1_341/CTRL2 0.10fF
C51432 VDD PAND2X1_123/Y 0.04fF
C51433 POR2X1_245/O POR2X1_90/Y 0.01fF
C51434 PAND2X1_6/Y POR2X1_802/CTRL 0.00fF
C51435 POR2X1_204/O PAND2X1_63/B 0.02fF
C51436 INPUT_1 POR2X1_55/Y 0.21fF
C51437 POR2X1_73/Y POR2X1_142/Y 0.03fF
C51438 PAND2X1_472/B POR2X1_153/Y 0.02fF
C51439 POR2X1_96/A POR2X1_129/Y 0.03fF
C51440 POR2X1_41/B POR2X1_271/A 0.12fF
C51441 PAND2X1_94/A PAND2X1_283/CTRL2 0.17fF
C51442 POR2X1_68/A POR2X1_799/O 0.05fF
C51443 POR2X1_36/B D_INPUT_6 0.44fF
C51444 POR2X1_417/CTRL2 POR2X1_7/A 0.03fF
C51445 PAND2X1_319/B PAND2X1_787/A 0.03fF
C51446 PAND2X1_175/B POR2X1_73/Y 0.03fF
C51447 POR2X1_66/B PAND2X1_665/m4_208_n4# 0.15fF
C51448 POR2X1_330/Y POR2X1_330/a_16_28# 0.06fF
C51449 POR2X1_383/A POR2X1_570/B 0.02fF
C51450 POR2X1_174/A PAND2X1_72/A 0.12fF
C51451 PAND2X1_7/O POR2X1_260/A 0.01fF
C51452 PAND2X1_659/Y POR2X1_821/CTRL 0.00fF
C51453 POR2X1_174/m4_208_n4# PAND2X1_72/A 0.12fF
C51454 POR2X1_315/Y POR2X1_90/Y 0.01fF
C51455 POR2X1_461/Y POR2X1_848/O 0.01fF
C51456 PAND2X1_467/Y PAND2X1_565/A 0.01fF
C51457 PAND2X1_6/Y PAND2X1_94/A 0.35fF
C51458 POR2X1_857/B POR2X1_227/CTRL 0.03fF
C51459 POR2X1_775/A POR2X1_332/CTRL 0.01fF
C51460 POR2X1_55/Y POR2X1_153/Y 0.46fF
C51461 POR2X1_93/A POR2X1_384/CTRL 0.01fF
C51462 POR2X1_114/Y POR2X1_294/A 0.05fF
C51463 POR2X1_57/A PAND2X1_349/A 0.03fF
C51464 POR2X1_123/B POR2X1_383/A 0.01fF
C51465 POR2X1_416/B POR2X1_40/Y 0.99fF
C51466 POR2X1_502/A PAND2X1_142/a_76_28# 0.02fF
C51467 POR2X1_384/A POR2X1_55/Y 0.03fF
C51468 POR2X1_96/A PAND2X1_659/Y 0.06fF
C51469 PAND2X1_150/a_16_344# PAND2X1_63/B 0.02fF
C51470 PAND2X1_476/A PAND2X1_473/Y 0.01fF
C51471 POR2X1_394/A PAND2X1_324/Y 0.03fF
C51472 POR2X1_544/O POR2X1_854/B 0.04fF
C51473 POR2X1_213/B POR2X1_568/B 0.05fF
C51474 PAND2X1_495/CTRL2 POR2X1_260/A 0.02fF
C51475 POR2X1_278/Y POR2X1_680/CTRL2 0.05fF
C51476 PAND2X1_631/A PAND2X1_515/CTRL2 0.04fF
C51477 POR2X1_762/a_16_28# INPUT_4 0.02fF
C51478 POR2X1_96/A POR2X1_96/Y 0.01fF
C51479 PAND2X1_55/Y POR2X1_722/CTRL 0.00fF
C51480 POR2X1_228/a_76_344# POR2X1_294/B 0.00fF
C51481 POR2X1_48/A POR2X1_9/Y 0.18fF
C51482 POR2X1_553/A PAND2X1_60/B 0.03fF
C51483 POR2X1_537/Y PAND2X1_55/Y 0.02fF
C51484 POR2X1_568/Y POR2X1_319/Y 0.05fF
C51485 POR2X1_8/Y PAND2X1_341/A 0.01fF
C51486 PAND2X1_6/O POR2X1_68/B 0.09fF
C51487 PAND2X1_20/A PAND2X1_125/CTRL 0.01fF
C51488 PAND2X1_244/B PAND2X1_175/B 0.01fF
C51489 POR2X1_119/Y POR2X1_697/Y 0.03fF
C51490 POR2X1_686/A PAND2X1_72/A 0.00fF
C51491 POR2X1_860/A PAND2X1_72/A 0.00fF
C51492 PAND2X1_47/B POR2X1_451/A 0.04fF
C51493 POR2X1_236/Y POR2X1_77/Y 0.24fF
C51494 POR2X1_8/Y POR2X1_93/A 0.01fF
C51495 PAND2X1_569/B POR2X1_766/CTRL 0.03fF
C51496 POR2X1_763/Y POR2X1_524/CTRL 0.01fF
C51497 POR2X1_60/A PAND2X1_193/Y 0.23fF
C51498 POR2X1_815/O POR2X1_816/Y 0.00fF
C51499 POR2X1_608/a_56_344# PAND2X1_56/A 0.00fF
C51500 POR2X1_391/CTRL POR2X1_260/A 0.11fF
C51501 POR2X1_556/A PAND2X1_268/O 0.01fF
C51502 POR2X1_383/A POR2X1_351/a_16_28# 0.03fF
C51503 POR2X1_240/A POR2X1_240/a_16_28# 0.05fF
C51504 PAND2X1_866/O PAND2X1_568/B 0.02fF
C51505 POR2X1_316/Y PAND2X1_465/B 0.04fF
C51506 POR2X1_778/CTRL2 POR2X1_717/B 0.01fF
C51507 POR2X1_407/A POR2X1_188/Y 0.03fF
C51508 PAND2X1_531/CTRL2 PAND2X1_111/B 0.00fF
C51509 PAND2X1_349/A PAND2X1_301/O 0.02fF
C51510 POR2X1_383/A PAND2X1_701/CTRL2 0.01fF
C51511 PAND2X1_63/Y POR2X1_294/A 0.03fF
C51512 POR2X1_327/Y POR2X1_137/Y 0.03fF
C51513 PAND2X1_824/B PAND2X1_824/O 0.04fF
C51514 POR2X1_829/A POR2X1_39/B 0.06fF
C51515 POR2X1_447/a_16_28# POR2X1_186/B 0.00fF
C51516 POR2X1_13/A POR2X1_387/O 0.16fF
C51517 PAND2X1_787/A PAND2X1_357/CTRL2 0.00fF
C51518 POR2X1_334/A PAND2X1_60/B 0.17fF
C51519 PAND2X1_323/CTRL2 POR2X1_702/A 0.00fF
C51520 PAND2X1_109/CTRL2 POR2X1_775/A 0.01fF
C51521 POR2X1_7/A POR2X1_129/Y 0.75fF
C51522 POR2X1_329/A POR2X1_32/A 21.02fF
C51523 POR2X1_327/CTRL2 PAND2X1_72/A 0.01fF
C51524 PAND2X1_644/O POR2X1_669/B 0.02fF
C51525 PAND2X1_130/O POR2X1_129/Y -0.00fF
C51526 POR2X1_113/Y POR2X1_294/A 0.07fF
C51527 POR2X1_191/Y POR2X1_577/O 0.29fF
C51528 POR2X1_285/B PAND2X1_55/Y 0.01fF
C51529 POR2X1_477/A POR2X1_711/Y 0.07fF
C51530 POR2X1_132/O PAND2X1_140/A 0.01fF
C51531 PAND2X1_440/CTRL2 PAND2X1_798/B 0.02fF
C51532 POR2X1_54/Y POR2X1_862/A 0.01fF
C51533 POR2X1_20/B POR2X1_626/CTRL2 0.03fF
C51534 POR2X1_119/Y PAND2X1_344/a_16_344# 0.02fF
C51535 POR2X1_63/Y POR2X1_23/Y 0.23fF
C51536 POR2X1_428/O POR2X1_394/A 0.01fF
C51537 POR2X1_831/a_16_28# POR2X1_301/A 0.11fF
C51538 POR2X1_852/A POR2X1_568/A 0.01fF
C51539 POR2X1_567/A POR2X1_510/Y 0.05fF
C51540 PAND2X1_222/a_76_28# PAND2X1_222/A 0.01fF
C51541 POR2X1_675/Y POR2X1_741/A 0.01fF
C51542 PAND2X1_326/CTRL PAND2X1_324/Y 0.01fF
C51543 POR2X1_417/Y POR2X1_329/A 0.25fF
C51544 POR2X1_329/A POR2X1_419/Y 0.04fF
C51545 POR2X1_99/B POR2X1_222/A 0.02fF
C51546 POR2X1_681/a_16_28# POR2X1_32/A 0.01fF
C51547 POR2X1_416/B POR2X1_136/CTRL2 0.01fF
C51548 POR2X1_96/Y POR2X1_7/A 0.03fF
C51549 POR2X1_180/B POR2X1_337/Y 0.01fF
C51550 PAND2X1_301/CTRL2 POR2X1_75/Y 0.01fF
C51551 POR2X1_30/a_16_28# D_INPUT_4 0.05fF
C51552 POR2X1_48/A PAND2X1_606/CTRL2 0.03fF
C51553 POR2X1_57/A POR2X1_43/CTRL2 0.03fF
C51554 POR2X1_516/A PAND2X1_631/A 0.01fF
C51555 PAND2X1_634/O POR2X1_102/Y 0.17fF
C51556 POR2X1_294/A POR2X1_260/A 0.25fF
C51557 POR2X1_813/O POR2X1_32/A 0.01fF
C51558 POR2X1_16/A POR2X1_767/O 0.01fF
C51559 POR2X1_65/A PAND2X1_206/B 0.11fF
C51560 PAND2X1_60/B D_INPUT_4 0.01fF
C51561 POR2X1_54/Y PAND2X1_73/Y 0.03fF
C51562 PAND2X1_39/B PAND2X1_39/O 0.01fF
C51563 POR2X1_16/A POR2X1_41/Y 0.00fF
C51564 POR2X1_14/m4_208_n4# INPUT_3 0.01fF
C51565 POR2X1_567/A POR2X1_543/O 0.14fF
C51566 POR2X1_651/Y POR2X1_664/Y 0.13fF
C51567 POR2X1_84/A POR2X1_66/A 0.06fF
C51568 PAND2X1_199/B POR2X1_153/Y 0.05fF
C51569 POR2X1_864/A POR2X1_750/B 0.03fF
C51570 POR2X1_16/A PAND2X1_649/A 0.00fF
C51571 POR2X1_698/Y PAND2X1_709/CTRL 0.00fF
C51572 POR2X1_520/CTRL POR2X1_383/Y 0.01fF
C51573 POR2X1_539/A POR2X1_374/a_16_28# 0.02fF
C51574 POR2X1_329/A PAND2X1_741/B 0.03fF
C51575 PAND2X1_290/CTRL2 PAND2X1_94/A 0.00fF
C51576 PAND2X1_798/Y PAND2X1_356/a_16_344# 0.03fF
C51577 POR2X1_12/A POR2X1_83/B 0.05fF
C51578 POR2X1_558/B POR2X1_218/Y 0.06fF
C51579 D_INPUT_7 PAND2X1_11/CTRL2 0.00fF
C51580 POR2X1_814/A VDD 11.18fF
C51581 POR2X1_702/A POR2X1_579/O 0.01fF
C51582 PAND2X1_68/CTRL2 D_INPUT_0 0.01fF
C51583 POR2X1_777/B PAND2X1_9/Y 0.09fF
C51584 POR2X1_604/O POR2X1_40/Y 0.01fF
C51585 PAND2X1_271/CTRL POR2X1_330/Y 0.01fF
C51586 POR2X1_66/B PAND2X1_612/B 0.15fF
C51587 POR2X1_369/m4_208_n4# PAND2X1_803/m4_208_n4# 0.13fF
C51588 PAND2X1_449/O POR2X1_236/Y 0.02fF
C51589 POR2X1_728/A PAND2X1_158/O 0.00fF
C51590 PAND2X1_221/Y PAND2X1_794/B 0.03fF
C51591 POR2X1_119/Y POR2X1_117/Y 0.64fF
C51592 POR2X1_144/CTRL PAND2X1_797/Y 0.09fF
C51593 POR2X1_846/Y VDD 0.30fF
C51594 POR2X1_863/m4_208_n4# POR2X1_797/m4_208_n4# 0.13fF
C51595 PAND2X1_247/O POR2X1_5/Y 0.15fF
C51596 POR2X1_265/CTRL POR2X1_40/Y 0.01fF
C51597 POR2X1_91/CTRL2 POR2X1_91/Y 0.01fF
C51598 PAND2X1_476/A POR2X1_7/Y 0.03fF
C51599 PAND2X1_94/A PAND2X1_52/B 0.30fF
C51600 POR2X1_660/Y POR2X1_78/A 0.03fF
C51601 POR2X1_411/B POR2X1_481/A 0.01fF
C51602 POR2X1_567/A POR2X1_741/CTRL2 0.01fF
C51603 POR2X1_586/Y POR2X1_585/Y 0.01fF
C51604 PAND2X1_678/CTRL PAND2X1_804/B 0.01fF
C51605 POR2X1_260/B PAND2X1_597/CTRL2 0.01fF
C51606 POR2X1_814/A POR2X1_741/Y 0.10fF
C51607 POR2X1_261/A POR2X1_257/A 0.03fF
C51608 POR2X1_142/CTRL2 POR2X1_669/B 0.03fF
C51609 POR2X1_485/Y POR2X1_46/Y 0.51fF
C51610 PAND2X1_75/O POR2X1_740/Y 0.02fF
C51611 PAND2X1_75/CTRL POR2X1_741/Y 0.00fF
C51612 POR2X1_703/O POR2X1_169/A 0.01fF
C51613 POR2X1_116/A POR2X1_114/Y 0.17fF
C51614 POR2X1_471/CTRL POR2X1_471/A 0.01fF
C51615 PAND2X1_301/CTRL2 PAND2X1_332/Y 0.03fF
C51616 PAND2X1_357/O POR2X1_39/B 0.04fF
C51617 POR2X1_227/A POR2X1_776/B 0.03fF
C51618 PAND2X1_420/CTRL2 POR2X1_590/A 0.00fF
C51619 POR2X1_329/A POR2X1_184/Y 0.03fF
C51620 POR2X1_311/Y PAND2X1_362/A 1.68fF
C51621 POR2X1_517/a_56_344# PAND2X1_404/Y 0.00fF
C51622 POR2X1_169/A POR2X1_337/Y 0.04fF
C51623 POR2X1_566/A POR2X1_776/A 0.73fF
C51624 PAND2X1_23/Y POR2X1_554/B 0.03fF
C51625 POR2X1_159/CTRL POR2X1_669/B 0.01fF
C51626 POR2X1_66/B POR2X1_267/CTRL2 0.01fF
C51627 POR2X1_842/m4_208_n4# POR2X1_794/B 0.08fF
C51628 PAND2X1_65/B PAND2X1_237/CTRL2 -0.00fF
C51629 PAND2X1_859/A POR2X1_37/Y 0.11fF
C51630 POR2X1_466/A PAND2X1_41/B 0.35fF
C51631 POR2X1_188/A POR2X1_858/O 0.01fF
C51632 POR2X1_444/B VDD 0.05fF
C51633 POR2X1_834/a_16_28# POR2X1_678/A 0.05fF
C51634 POR2X1_150/Y PAND2X1_736/Y 0.01fF
C51635 POR2X1_257/A POR2X1_425/O 0.01fF
C51636 POR2X1_814/A PAND2X1_32/B 0.22fF
C51637 PAND2X1_34/a_76_28# POR2X1_27/Y 0.02fF
C51638 POR2X1_593/O PAND2X1_72/A 0.01fF
C51639 PAND2X1_633/CTRL2 POR2X1_32/A 0.01fF
C51640 POR2X1_16/A POR2X1_234/A 0.04fF
C51641 PAND2X1_58/A POR2X1_330/Y 0.07fF
C51642 POR2X1_312/CTRL2 POR2X1_20/B 0.00fF
C51643 POR2X1_660/CTRL2 POR2X1_660/A 0.01fF
C51644 POR2X1_271/B PAND2X1_658/B 0.05fF
C51645 PAND2X1_65/B PAND2X1_591/a_16_344# 0.01fF
C51646 PAND2X1_205/A INPUT_0 0.03fF
C51647 POR2X1_356/A POR2X1_446/B 0.05fF
C51648 POR2X1_450/B POR2X1_450/A 0.01fF
C51649 PAND2X1_52/B PAND2X1_680/CTRL2 0.02fF
C51650 PAND2X1_771/Y PAND2X1_345/O 0.23fF
C51651 POR2X1_102/Y POR2X1_595/Y 0.02fF
C51652 POR2X1_84/CTRL POR2X1_84/B 0.00fF
C51653 PAND2X1_609/CTRL2 POR2X1_294/B 0.03fF
C51654 POR2X1_624/Y POR2X1_501/CTRL 0.03fF
C51655 POR2X1_12/A PAND2X1_709/O 0.02fF
C51656 POR2X1_687/O VDD 0.00fF
C51657 PAND2X1_223/B PAND2X1_539/B 0.01fF
C51658 POR2X1_458/Y PAND2X1_300/CTRL 0.01fF
C51659 POR2X1_566/A POR2X1_856/B 0.11fF
C51660 POR2X1_60/A POR2X1_763/A 0.02fF
C51661 PAND2X1_81/CTRL PAND2X1_9/Y 0.01fF
C51662 POR2X1_487/CTRL2 PAND2X1_738/Y 0.17fF
C51663 PAND2X1_48/B POR2X1_260/B 5.24fF
C51664 POR2X1_20/B POR2X1_234/a_16_28# 0.01fF
C51665 POR2X1_864/A POR2X1_686/CTRL2 0.00fF
C51666 PAND2X1_277/a_16_344# PAND2X1_57/B 0.03fF
C51667 POR2X1_96/A POR2X1_37/Y 0.03fF
C51668 POR2X1_706/a_16_28# POR2X1_706/B 0.02fF
C51669 POR2X1_69/A PAND2X1_340/CTRL 0.00fF
C51670 POR2X1_614/A POR2X1_471/A 0.34fF
C51671 POR2X1_96/A POR2X1_271/a_16_28# 0.02fF
C51672 PAND2X1_80/O PAND2X1_73/Y 0.04fF
C51673 POR2X1_423/CTRL2 INPUT_0 0.13fF
C51674 POR2X1_377/a_16_28# POR2X1_54/Y 0.03fF
C51675 POR2X1_13/CTRL2 POR2X1_102/Y 0.00fF
C51676 POR2X1_13/A POR2X1_29/A 0.00fF
C51677 POR2X1_341/A POR2X1_500/Y 0.01fF
C51678 PAND2X1_803/Y POR2X1_150/Y 0.02fF
C51679 POR2X1_609/Y POR2X1_290/Y 0.03fF
C51680 PAND2X1_58/A POR2X1_585/m4_208_n4# 0.05fF
C51681 PAND2X1_65/B POR2X1_808/A 0.03fF
C51682 POR2X1_673/Y POR2X1_814/A 0.03fF
C51683 PAND2X1_496/CTRL D_INPUT_0 0.01fF
C51684 POR2X1_807/O POR2X1_294/B 0.01fF
C51685 PAND2X1_39/B PAND2X1_88/Y 0.03fF
C51686 POR2X1_343/CTRL POR2X1_343/B 0.01fF
C51687 POR2X1_306/O PAND2X1_454/B 0.01fF
C51688 POR2X1_673/CTRL PAND2X1_8/Y 0.09fF
C51689 POR2X1_34/Y VDD -0.00fF
C51690 POR2X1_78/A PAND2X1_322/CTRL 0.02fF
C51691 POR2X1_307/a_16_28# POR2X1_307/B -0.00fF
C51692 POR2X1_333/A POR2X1_192/Y 0.17fF
C51693 PAND2X1_668/CTRL2 POR2X1_83/B 0.00fF
C51694 POR2X1_84/a_16_28# POR2X1_84/A 0.03fF
C51695 PAND2X1_833/a_16_344# POR2X1_482/Y 0.02fF
C51696 PAND2X1_489/a_76_28# POR2X1_42/Y 0.01fF
C51697 POR2X1_28/CTRL2 D_INPUT_1 0.03fF
C51698 POR2X1_817/O PAND2X1_6/A 0.07fF
C51699 POR2X1_62/Y POR2X1_9/Y 1.68fF
C51700 POR2X1_135/Y POR2X1_423/Y 0.01fF
C51701 POR2X1_832/Y PAND2X1_69/A 3.56fF
C51702 POR2X1_786/A POR2X1_78/A 0.67fF
C51703 PAND2X1_354/A VDD 0.68fF
C51704 POR2X1_66/B POR2X1_220/Y 0.06fF
C51705 POR2X1_498/Y POR2X1_494/Y 0.02fF
C51706 POR2X1_435/Y POR2X1_330/Y 0.10fF
C51707 PAND2X1_738/Y POR2X1_40/Y 0.09fF
C51708 POR2X1_138/CTRL POR2X1_296/B 0.01fF
C51709 POR2X1_290/O POR2X1_236/Y 0.01fF
C51710 POR2X1_653/CTRL2 POR2X1_653/B 0.01fF
C51711 PAND2X1_20/A POR2X1_231/B 0.03fF
C51712 POR2X1_92/a_16_28# INPUT_3 0.03fF
C51713 POR2X1_529/O POR2X1_29/A 0.04fF
C51714 POR2X1_669/B PAND2X1_324/Y 0.03fF
C51715 INPUT_1 POR2X1_19/O 0.18fF
C51716 POR2X1_852/B VDD 2.24fF
C51717 PAND2X1_217/B PAND2X1_598/CTRL2 0.32fF
C51718 POR2X1_78/B POR2X1_718/A 0.07fF
C51719 POR2X1_84/A POR2X1_532/A 0.00fF
C51720 POR2X1_96/A PAND2X1_78/a_16_344# 0.01fF
C51721 POR2X1_23/Y PAND2X1_575/CTRL2 0.03fF
C51722 INPUT_2 POR2X1_48/A 0.05fF
C51723 POR2X1_119/O POR2X1_102/Y 0.01fF
C51724 POR2X1_188/A POR2X1_220/Y 0.13fF
C51725 POR2X1_66/B POR2X1_404/Y 0.40fF
C51726 POR2X1_78/O D_INPUT_0 0.01fF
C51727 PAND2X1_96/B POR2X1_734/B 0.01fF
C51728 POR2X1_65/A PAND2X1_739/Y 0.03fF
C51729 POR2X1_301/CTRL2 POR2X1_590/A 0.03fF
C51730 POR2X1_76/CTRL POR2X1_274/B 0.01fF
C51731 PAND2X1_224/O POR2X1_191/Y 0.01fF
C51732 POR2X1_49/Y PAND2X1_149/CTRL 0.01fF
C51733 POR2X1_37/Y PAND2X1_342/O 0.00fF
C51734 POR2X1_17/CTRL2 INPUT_5 0.01fF
C51735 POR2X1_305/Y PAND2X1_777/a_76_28# 0.04fF
C51736 POR2X1_409/B POR2X1_73/Y 0.03fF
C51737 PAND2X1_90/A PAND2X1_46/CTRL2 0.03fF
C51738 PAND2X1_76/Y INPUT_0 0.07fF
C51739 POR2X1_798/CTRL POR2X1_468/B 0.01fF
C51740 PAND2X1_65/B POR2X1_483/CTRL2 0.00fF
C51741 PAND2X1_96/B POR2X1_792/CTRL2 0.01fF
C51742 PAND2X1_843/a_76_28# PAND2X1_738/Y 0.04fF
C51743 POR2X1_383/A POR2X1_647/O 0.03fF
C51744 D_INPUT_0 POR2X1_291/Y 0.02fF
C51745 PAND2X1_129/m4_208_n4# POR2X1_264/m4_208_n4# 0.13fF
C51746 POR2X1_41/B PAND2X1_499/CTRL 0.07fF
C51747 PAND2X1_474/A PAND2X1_735/a_76_28# 0.01fF
C51748 PAND2X1_449/Y POR2X1_14/Y 0.02fF
C51749 PAND2X1_20/A POR2X1_790/A 0.02fF
C51750 POR2X1_254/Y POR2X1_483/A 0.06fF
C51751 PAND2X1_25/CTRL2 INPUT_6 0.00fF
C51752 POR2X1_60/A POR2X1_183/Y 0.03fF
C51753 POR2X1_808/A PAND2X1_599/O 0.09fF
C51754 PAND2X1_96/B POR2X1_555/B 0.03fF
C51755 PAND2X1_449/Y PAND2X1_453/A 0.02fF
C51756 PAND2X1_659/Y POR2X1_760/A 0.07fF
C51757 POR2X1_232/CTRL2 POR2X1_5/Y 0.03fF
C51758 PAND2X1_682/O POR2X1_467/Y 0.02fF
C51759 PAND2X1_859/A POR2X1_224/Y 0.01fF
C51760 POR2X1_419/Y PAND2X1_506/a_16_344# 0.03fF
C51761 D_INPUT_0 POR2X1_575/CTRL 0.01fF
C51762 POR2X1_690/a_76_344# INPUT_0 0.02fF
C51763 POR2X1_662/CTRL POR2X1_353/A 0.01fF
C51764 POR2X1_57/A POR2X1_32/A 1.20fF
C51765 PAND2X1_20/A PAND2X1_83/O 0.03fF
C51766 POR2X1_75/O POR2X1_60/A 0.20fF
C51767 POR2X1_401/B VDD 0.02fF
C51768 PAND2X1_63/Y PAND2X1_265/O 0.04fF
C51769 POR2X1_37/Y POR2X1_7/A 0.10fF
C51770 PAND2X1_425/Y PAND2X1_2/CTRL 0.01fF
C51771 POR2X1_322/CTRL POR2X1_376/B 0.01fF
C51772 POR2X1_227/A POR2X1_192/B 0.05fF
C51773 POR2X1_164/CTRL2 POR2X1_72/B 0.01fF
C51774 POR2X1_852/B POR2X1_741/Y 0.10fF
C51775 PAND2X1_804/O POR2X1_283/A 0.02fF
C51776 POR2X1_287/A POR2X1_188/Y 0.00fF
C51777 PAND2X1_452/A PAND2X1_452/a_76_28# 0.02fF
C51778 POR2X1_96/A POR2X1_406/Y 0.03fF
C51779 PAND2X1_473/Y PAND2X1_479/B -0.00fF
C51780 POR2X1_130/A POR2X1_722/Y 0.02fF
C51781 PAND2X1_863/B INPUT_0 0.03fF
C51782 PAND2X1_805/A PAND2X1_567/a_16_344# 0.02fF
C51783 PAND2X1_20/A PAND2X1_88/Y 0.03fF
C51784 PAND2X1_732/CTRL PAND2X1_731/A 0.01fF
C51785 PAND2X1_732/a_16_344# POR2X1_152/Y 0.01fF
C51786 PAND2X1_20/A POR2X1_84/Y 0.00fF
C51787 POR2X1_43/B PAND2X1_61/Y 0.09fF
C51788 POR2X1_405/CTRL2 PAND2X1_32/B 0.01fF
C51789 POR2X1_528/a_16_28# POR2X1_748/A 0.06fF
C51790 INPUT_5 VDD 0.91fF
C51791 POR2X1_16/A PAND2X1_207/O -0.00fF
C51792 POR2X1_68/A POR2X1_543/A 0.29fF
C51793 POR2X1_61/Y D_GATE_222 0.07fF
C51794 POR2X1_265/Y PAND2X1_267/B 0.02fF
C51795 POR2X1_32/A POR2X1_229/Y 0.65fF
C51796 POR2X1_669/B PAND2X1_720/CTRL2 -0.02fF
C51797 PAND2X1_269/CTRL POR2X1_39/B 0.08fF
C51798 POR2X1_634/A PAND2X1_757/CTRL2 0.17fF
C51799 POR2X1_669/B PAND2X1_549/B 0.10fF
C51800 PAND2X1_96/B POR2X1_330/Y 0.12fF
C51801 PAND2X1_57/B PAND2X1_751/CTRL 0.00fF
C51802 POR2X1_322/Y POR2X1_83/B 0.01fF
C51803 POR2X1_407/A PAND2X1_679/CTRL 0.03fF
C51804 POR2X1_68/A PAND2X1_679/O 0.03fF
C51805 PAND2X1_9/a_76_28# D_INPUT_1 0.02fF
C51806 POR2X1_33/B POR2X1_68/B 0.04fF
C51807 PAND2X1_724/B VDD 0.49fF
C51808 POR2X1_647/B PAND2X1_48/A 0.03fF
C51809 POR2X1_57/A POR2X1_417/Y 0.03fF
C51810 POR2X1_260/Y VDD 0.08fF
C51811 POR2X1_218/Y POR2X1_362/A 0.01fF
C51812 POR2X1_57/A POR2X1_419/Y 0.03fF
C51813 PAND2X1_470/A POR2X1_14/Y 0.05fF
C51814 PAND2X1_55/Y PAND2X1_58/O 0.02fF
C51815 PAND2X1_652/A PAND2X1_192/a_16_344# 0.01fF
C51816 PAND2X1_41/B POR2X1_194/CTRL2 0.03fF
C51817 POR2X1_750/B POR2X1_194/O 0.06fF
C51818 POR2X1_38/Y PAND2X1_733/CTRL2 0.00fF
C51819 POR2X1_29/A PAND2X1_510/B 0.00fF
C51820 PAND2X1_659/A POR2X1_73/Y 0.96fF
C51821 POR2X1_5/Y POR2X1_382/a_16_28# 0.01fF
C51822 PAND2X1_48/B POR2X1_723/O 0.11fF
C51823 POR2X1_733/a_16_28# POR2X1_733/A 0.04fF
C51824 POR2X1_96/A POR2X1_293/Y 0.21fF
C51825 POR2X1_13/CTRL POR2X1_13/Y 0.01fF
C51826 PAND2X1_55/Y POR2X1_483/B 0.01fF
C51827 POR2X1_60/A PAND2X1_535/O 0.03fF
C51828 PAND2X1_850/Y POR2X1_275/A 0.16fF
C51829 PAND2X1_48/B PAND2X1_516/CTRL 0.09fF
C51830 POR2X1_302/A VDD 0.04fF
C51831 POR2X1_407/Y PAND2X1_597/CTRL2 0.01fF
C51832 POR2X1_408/CTRL2 INPUT_5 0.00fF
C51833 POR2X1_278/Y PAND2X1_197/Y 0.05fF
C51834 PAND2X1_131/CTRL POR2X1_130/Y 0.01fF
C51835 POR2X1_390/B POR2X1_296/B 0.03fF
C51836 POR2X1_16/A POR2X1_601/O 0.00fF
C51837 POR2X1_107/CTRL2 POR2X1_90/Y 0.02fF
C51838 PAND2X1_387/a_76_28# POR2X1_712/Y 0.00fF
C51839 POR2X1_669/B POR2X1_428/O 0.03fF
C51840 PAND2X1_795/B PAND2X1_575/A 0.03fF
C51841 PAND2X1_855/CTRL2 POR2X1_236/Y 0.04fF
C51842 PAND2X1_73/Y POR2X1_175/B 0.02fF
C51843 POR2X1_136/Y POR2X1_40/Y 0.43fF
C51844 PAND2X1_118/CTRL2 POR2X1_502/A 0.43fF
C51845 POR2X1_850/A POR2X1_840/B 1.27fF
C51846 POR2X1_865/B POR2X1_814/B 0.03fF
C51847 POR2X1_814/B PAND2X1_88/Y 0.10fF
C51848 POR2X1_478/B PAND2X1_41/B 1.50fF
C51849 POR2X1_97/B POR2X1_454/A 0.03fF
C51850 PAND2X1_65/Y POR2X1_532/A 0.38fF
C51851 POR2X1_32/A PAND2X1_301/O 0.01fF
C51852 PAND2X1_181/CTRL2 POR2X1_40/Y 0.00fF
C51853 POR2X1_639/Y PAND2X1_65/B 0.03fF
C51854 POR2X1_109/O POR2X1_109/Y 0.02fF
C51855 PAND2X1_48/B PAND2X1_280/a_16_344# 0.01fF
C51856 PAND2X1_471/CTRL2 PAND2X1_464/Y 0.01fF
C51857 POR2X1_72/B POR2X1_283/A 0.03fF
C51858 PAND2X1_859/A POR2X1_408/Y 0.58fF
C51859 PAND2X1_614/CTRL POR2X1_283/A 0.01fF
C51860 POR2X1_68/A POR2X1_214/CTRL 0.03fF
C51861 POR2X1_139/O VDD 0.00fF
C51862 PAND2X1_855/CTRL VDD -0.00fF
C51863 POR2X1_237/a_56_344# POR2X1_90/Y 0.00fF
C51864 POR2X1_529/Y PAND2X1_474/A 0.06fF
C51865 POR2X1_57/A PAND2X1_319/O 0.01fF
C51866 PAND2X1_48/B PAND2X1_55/Y 8.98fF
C51867 PAND2X1_549/O POR2X1_531/Y -0.00fF
C51868 PAND2X1_349/A PAND2X1_140/a_16_344# 0.01fF
C51869 POR2X1_356/A POR2X1_795/B 0.05fF
C51870 POR2X1_57/A PAND2X1_741/B 0.01fF
C51871 POR2X1_278/Y PAND2X1_359/O 0.17fF
C51872 PAND2X1_480/B POR2X1_90/Y 0.07fF
C51873 PAND2X1_241/Y POR2X1_236/Y 0.02fF
C51874 PAND2X1_48/B POR2X1_205/O 0.01fF
C51875 POR2X1_52/A POR2X1_93/CTRL2 0.01fF
C51876 POR2X1_773/CTRL2 POR2X1_734/A 0.05fF
C51877 POR2X1_252/O PAND2X1_6/A 0.03fF
C51878 PAND2X1_48/B POR2X1_363/O 0.02fF
C51879 POR2X1_56/Y PAND2X1_364/B 0.08fF
C51880 D_GATE_741 POR2X1_785/A 0.07fF
C51881 PAND2X1_556/O PAND2X1_348/A 0.05fF
C51882 POR2X1_66/B PAND2X1_748/a_56_28# 0.00fF
C51883 POR2X1_67/A PAND2X1_156/A 0.04fF
C51884 PAND2X1_254/CTRL2 PAND2X1_6/A 0.10fF
C51885 PAND2X1_96/B POR2X1_449/a_16_28# 0.02fF
C51886 POR2X1_614/A POR2X1_570/a_16_28# 0.03fF
C51887 POR2X1_754/A POR2X1_90/Y 0.03fF
C51888 POR2X1_94/A POR2X1_260/A 0.03fF
C51889 INPUT_4 POR2X1_3/CTRL2 0.05fF
C51890 POR2X1_307/Y PAND2X1_69/A 0.03fF
C51891 INPUT_5 PAND2X1_32/B 0.05fF
C51892 POR2X1_480/A POR2X1_537/A 0.01fF
C51893 POR2X1_42/Y POR2X1_396/O 0.01fF
C51894 POR2X1_13/A POR2X1_583/O 0.01fF
C51895 POR2X1_301/CTRL POR2X1_335/A 0.01fF
C51896 POR2X1_537/CTRL POR2X1_862/B 0.00fF
C51897 PAND2X1_65/B POR2X1_687/A 0.01fF
C51898 POR2X1_78/B POR2X1_725/Y 0.07fF
C51899 POR2X1_406/Y POR2X1_7/A 0.03fF
C51900 D_GATE_222 POR2X1_35/Y 0.03fF
C51901 PAND2X1_421/O PAND2X1_69/A 0.03fF
C51902 POR2X1_16/A PAND2X1_340/CTRL 0.00fF
C51903 PAND2X1_23/Y POR2X1_702/A 0.12fF
C51904 D_GATE_741 PAND2X1_504/O 0.31fF
C51905 PAND2X1_48/B POR2X1_407/Y 0.02fF
C51906 PAND2X1_65/B POR2X1_352/O 0.01fF
C51907 PAND2X1_698/O PAND2X1_90/Y 0.21fF
C51908 PAND2X1_785/Y PAND2X1_175/B 0.00fF
C51909 POR2X1_52/A INPUT_6 0.01fF
C51910 POR2X1_96/A POR2X1_408/Y 0.01fF
C51911 PAND2X1_229/CTRL2 POR2X1_186/B 0.03fF
C51912 POR2X1_594/CTRL POR2X1_385/Y 0.00fF
C51913 PAND2X1_6/Y POR2X1_796/CTRL2 0.00fF
C51914 POR2X1_463/Y PAND2X1_90/Y 0.07fF
C51915 PAND2X1_825/CTRL PAND2X1_57/B 0.01fF
C51916 POR2X1_302/A PAND2X1_32/B 0.30fF
C51917 POR2X1_324/O POR2X1_324/A 0.01fF
C51918 POR2X1_83/B POR2X1_373/O -0.01fF
C51919 POR2X1_119/Y POR2X1_667/A 0.09fF
C51920 PAND2X1_35/Y POR2X1_229/Y 0.03fF
C51921 POR2X1_188/A POR2X1_709/B 0.01fF
C51922 PAND2X1_89/O PAND2X1_60/B 0.04fF
C51923 POR2X1_446/B PAND2X1_72/A 0.13fF
C51924 POR2X1_65/A PAND2X1_560/B 0.01fF
C51925 POR2X1_141/CTRL2 POR2X1_574/Y 0.02fF
C51926 POR2X1_57/A POR2X1_189/Y 0.03fF
C51927 POR2X1_60/A PAND2X1_199/CTRL 0.01fF
C51928 PAND2X1_392/CTRL POR2X1_39/B 0.31fF
C51929 POR2X1_78/B POR2X1_596/O 0.01fF
C51930 POR2X1_111/m4_208_n4# POR2X1_46/Y 0.06fF
C51931 POR2X1_326/A POR2X1_798/CTRL 0.01fF
C51932 PAND2X1_422/CTRL POR2X1_294/B 0.04fF
C51933 PAND2X1_244/B PAND2X1_351/Y 1.42fF
C51934 POR2X1_356/A POR2X1_383/A 0.32fF
C51935 PAND2X1_631/A PAND2X1_556/O 0.02fF
C51936 POR2X1_7/A POR2X1_293/Y 0.29fF
C51937 POR2X1_502/A PAND2X1_376/CTRL2 0.01fF
C51938 POR2X1_25/Y POR2X1_698/O 0.01fF
C51939 POR2X1_778/B D_INPUT_1 0.15fF
C51940 POR2X1_489/CTRL POR2X1_294/A 0.03fF
C51941 PAND2X1_777/O POR2X1_39/B 0.01fF
C51942 POR2X1_57/A POR2X1_184/Y 0.03fF
C51943 POR2X1_511/Y POR2X1_153/Y 0.18fF
C51944 POR2X1_51/A POR2X1_260/A 0.12fF
C51945 VDD PAND2X1_157/O 0.00fF
C51946 PAND2X1_635/CTRL2 INPUT_6 0.10fF
C51947 POR2X1_130/A POR2X1_244/Y 0.39fF
C51948 POR2X1_68/B PAND2X1_69/A 3.27fF
C51949 PAND2X1_341/Y POR2X1_88/Y 0.60fF
C51950 POR2X1_52/A PAND2X1_737/B 0.02fF
C51951 D_GATE_662 POR2X1_854/B 0.10fF
C51952 PAND2X1_726/B POR2X1_46/Y 0.39fF
C51953 POR2X1_751/O POR2X1_816/A 0.01fF
C51954 PAND2X1_20/A POR2X1_568/B 0.03fF
C51955 POR2X1_140/B POR2X1_510/Y 0.01fF
C51956 POR2X1_49/Y PAND2X1_476/A 0.03fF
C51957 PAND2X1_483/CTRL2 POR2X1_55/Y 0.02fF
C51958 POR2X1_136/CTRL2 POR2X1_136/Y 0.03fF
C51959 POR2X1_52/A PAND2X1_216/B 1.87fF
C51960 POR2X1_750/B PAND2X1_179/CTRL 0.01fF
C51961 VDD POR2X1_151/Y 0.12fF
C51962 D_INPUT_0 POR2X1_500/O 0.01fF
C51963 PAND2X1_56/Y POR2X1_569/A 0.10fF
C51964 PAND2X1_6/A POR2X1_245/Y 0.07fF
C51965 PAND2X1_6/Y POR2X1_348/CTRL 0.03fF
C51966 PAND2X1_388/Y PAND2X1_370/O 0.02fF
C51967 POR2X1_334/Y PAND2X1_261/O 0.09fF
C51968 POR2X1_43/B PAND2X1_651/A 0.05fF
C51969 POR2X1_379/Y VDD 0.04fF
C51970 POR2X1_69/A POR2X1_39/B 0.00fF
C51971 POR2X1_222/A POR2X1_112/Y 0.03fF
C51972 PAND2X1_169/Y POR2X1_39/B 0.03fF
C51973 POR2X1_582/O POR2X1_582/A -0.00fF
C51974 POR2X1_137/Y POR2X1_361/CTRL2 0.11fF
C51975 POR2X1_211/O POR2X1_566/B 0.00fF
C51976 PAND2X1_190/O POR2X1_131/A 0.06fF
C51977 PAND2X1_469/B POR2X1_310/Y 0.05fF
C51978 POR2X1_750/B D_INPUT_4 0.03fF
C51979 POR2X1_278/Y POR2X1_62/Y 0.03fF
C51980 POR2X1_465/B POR2X1_186/B 0.03fF
C51981 PAND2X1_11/Y PAND2X1_52/B 0.08fF
C51982 POR2X1_346/O PAND2X1_60/B 0.01fF
C51983 PAND2X1_578/O PAND2X1_578/A 0.00fF
C51984 POR2X1_824/O VDD 0.00fF
C51985 POR2X1_322/Y PAND2X1_168/CTRL2 0.00fF
C51986 POR2X1_121/B PAND2X1_72/A 0.12fF
C51987 POR2X1_219/a_16_28# POR2X1_215/Y 0.05fF
C51988 POR2X1_322/CTRL2 POR2X1_373/Y 0.01fF
C51989 PAND2X1_801/CTRL2 POR2X1_236/Y 0.04fF
C51990 POR2X1_366/Y POR2X1_317/B 0.02fF
C51991 POR2X1_814/B POR2X1_568/B 0.10fF
C51992 POR2X1_23/Y POR2X1_485/a_76_344# 0.01fF
C51993 POR2X1_327/Y POR2X1_366/Y 0.03fF
C51994 POR2X1_327/Y POR2X1_294/B 0.07fF
C51995 POR2X1_94/A PAND2X1_102/a_76_28# 0.01fF
C51996 POR2X1_730/Y POR2X1_614/A 0.03fF
C51997 POR2X1_184/Y PAND2X1_301/O 0.00fF
C51998 POR2X1_566/A POR2X1_191/Y 0.10fF
C51999 POR2X1_707/CTRL2 POR2X1_407/Y 0.01fF
C52000 POR2X1_112/O POR2X1_332/B 0.01fF
C52001 POR2X1_307/Y POR2X1_512/CTRL 0.01fF
C52002 PAND2X1_801/CTRL VDD 0.00fF
C52003 POR2X1_311/CTRL POR2X1_142/Y 0.00fF
C52004 POR2X1_408/Y POR2X1_7/A 0.09fF
C52005 POR2X1_740/Y POR2X1_195/CTRL 0.26fF
C52006 POR2X1_274/B POR2X1_228/Y 0.22fF
C52007 PAND2X1_865/Y PAND2X1_468/CTRL 0.01fF
C52008 PAND2X1_93/B POR2X1_457/Y 0.01fF
C52009 POR2X1_809/A POR2X1_800/A 0.03fF
C52010 PAND2X1_90/Y POR2X1_736/A 0.10fF
C52011 POR2X1_383/A POR2X1_569/A 0.14fF
C52012 POR2X1_416/B POR2X1_5/Y 0.16fF
C52013 PAND2X1_175/B PAND2X1_861/CTRL2 0.01fF
C52014 PAND2X1_306/O POR2X1_308/B 0.01fF
C52015 VDD PAND2X1_358/O 0.00fF
C52016 POR2X1_771/A POR2X1_771/a_16_28# 0.03fF
C52017 POR2X1_244/Y POR2X1_573/A 0.03fF
C52018 POR2X1_29/a_16_28# POR2X1_29/A 0.05fF
C52019 POR2X1_119/Y PAND2X1_716/CTRL2 0.13fF
C52020 POR2X1_11/O POR2X1_12/A 0.03fF
C52021 PAND2X1_716/O PAND2X1_716/B 0.04fF
C52022 PAND2X1_348/A POR2X1_142/Y 0.01fF
C52023 PAND2X1_48/B POR2X1_741/O 0.01fF
C52024 POR2X1_834/m4_208_n4# POR2X1_645/m4_208_n4# 0.15fF
C52025 POR2X1_475/A POR2X1_343/B 0.02fF
C52026 POR2X1_597/A POR2X1_761/A 0.31fF
C52027 POR2X1_845/A D_INPUT_1 0.06fF
C52028 VDD POR2X1_180/Y 0.10fF
C52029 POR2X1_730/Y POR2X1_440/Y 0.03fF
C52030 PAND2X1_65/B POR2X1_568/A 24.27fF
C52031 POR2X1_203/Y PAND2X1_48/A 0.34fF
C52032 PAND2X1_39/B POR2X1_341/A 0.07fF
C52033 PAND2X1_319/B PAND2X1_357/CTRL 0.01fF
C52034 VDD POR2X1_759/CTRL2 0.00fF
C52035 INPUT_6 POR2X1_3/B 1.01fF
C52036 PAND2X1_96/B POR2X1_337/Y 0.07fF
C52037 PAND2X1_20/A PAND2X1_234/O 0.08fF
C52038 PAND2X1_659/Y POR2X1_38/Y 0.06fF
C52039 POR2X1_691/a_16_28# POR2X1_691/A 0.05fF
C52040 POR2X1_544/B POR2X1_180/A 0.03fF
C52041 POR2X1_110/CTRL POR2X1_387/Y 0.05fF
C52042 POR2X1_736/CTRL POR2X1_188/Y 0.01fF
C52043 PAND2X1_270/a_16_344# PAND2X1_508/Y 0.02fF
C52044 POR2X1_803/CTRL POR2X1_796/Y 0.01fF
C52045 POR2X1_96/Y POR2X1_38/Y 0.07fF
C52046 PAND2X1_217/O PAND2X1_124/Y 0.05fF
C52047 POR2X1_550/Y POR2X1_550/B 0.02fF
C52048 PAND2X1_481/CTRL2 POR2X1_507/A 0.03fF
C52049 INPUT_1 POR2X1_129/Y 0.10fF
C52050 POR2X1_814/B PAND2X1_234/O 0.07fF
C52051 POR2X1_334/Y POR2X1_260/A 0.07fF
C52052 PAND2X1_551/A PAND2X1_326/CTRL2 0.01fF
C52053 POR2X1_40/CTRL POR2X1_25/Y 0.01fF
C52054 PAND2X1_409/a_76_28# PAND2X1_52/B 0.04fF
C52055 PAND2X1_732/A POR2X1_373/Y 0.03fF
C52056 PAND2X1_447/O POR2X1_102/Y 0.03fF
C52057 PAND2X1_73/Y POR2X1_78/Y 0.15fF
C52058 PAND2X1_785/CTRL2 POR2X1_77/Y 0.01fF
C52059 POR2X1_795/B PAND2X1_72/A 0.03fF
C52060 PAND2X1_56/Y PAND2X1_72/A 0.06fF
C52061 POR2X1_796/CTRL2 PAND2X1_52/B 0.03fF
C52062 PAND2X1_646/O POR2X1_612/Y 0.04fF
C52063 POR2X1_468/a_16_28# POR2X1_568/A 0.01fF
C52064 POR2X1_129/Y POR2X1_153/Y 0.06fF
C52065 POR2X1_334/Y POR2X1_363/A 0.01fF
C52066 PAND2X1_641/CTRL PAND2X1_476/A 0.00fF
C52067 POR2X1_287/B POR2X1_486/a_76_344# 0.00fF
C52068 PAND2X1_858/CTRL2 POR2X1_129/Y 0.01fF
C52069 POR2X1_643/CTRL POR2X1_121/Y 0.00fF
C52070 PAND2X1_20/A POR2X1_341/A 0.10fF
C52071 POR2X1_559/A POR2X1_294/A 0.10fF
C52072 INPUT_1 POR2X1_96/Y 0.03fF
C52073 POR2X1_158/Y POR2X1_426/Y 0.00fF
C52074 POR2X1_496/O PAND2X1_58/A 0.02fF
C52075 POR2X1_865/O PAND2X1_52/B 0.01fF
C52076 PAND2X1_659/Y POR2X1_153/Y 0.07fF
C52077 POR2X1_416/B PAND2X1_222/B 0.03fF
C52078 POR2X1_634/A PAND2X1_59/a_16_344# 0.06fF
C52079 POR2X1_20/B PAND2X1_390/Y 0.02fF
C52080 POR2X1_319/A POR2X1_174/A 0.03fF
C52081 POR2X1_672/Y POR2X1_83/B 0.00fF
C52082 POR2X1_102/Y PAND2X1_791/a_76_28# 0.01fF
C52083 POR2X1_327/Y POR2X1_567/A 0.09fF
C52084 POR2X1_263/Y D_INPUT_0 0.03fF
C52085 PAND2X1_6/Y POR2X1_303/B 0.03fF
C52086 POR2X1_96/Y POR2X1_153/Y 0.28fF
C52087 POR2X1_616/Y PAND2X1_156/A 0.03fF
C52088 POR2X1_60/A POR2X1_437/CTRL 0.02fF
C52089 POR2X1_67/Y POR2X1_859/A 0.03fF
C52090 POR2X1_51/A POR2X1_329/A 0.00fF
C52091 PAND2X1_827/O POR2X1_296/B 0.17fF
C52092 POR2X1_16/A POR2X1_39/B 0.44fF
C52093 POR2X1_66/B POR2X1_610/CTRL 0.01fF
C52094 POR2X1_83/B PAND2X1_124/Y 0.03fF
C52095 POR2X1_102/Y PAND2X1_205/A 0.03fF
C52096 POR2X1_814/B POR2X1_341/A 0.07fF
C52097 POR2X1_178/Y POR2X1_416/B 1.23fF
C52098 POR2X1_383/A PAND2X1_72/A 7.86fF
C52099 POR2X1_863/A POR2X1_535/A 0.01fF
C52100 POR2X1_78/B POR2X1_318/CTRL2 0.03fF
C52101 POR2X1_856/B POR2X1_241/B 0.03fF
C52102 POR2X1_97/B POR2X1_99/B 0.03fF
C52103 POR2X1_338/a_56_344# PAND2X1_72/A 0.00fF
C52104 POR2X1_99/O POR2X1_243/Y 0.01fF
C52105 PAND2X1_464/B POR2X1_7/B 0.03fF
C52106 POR2X1_188/A POR2X1_841/B 0.00fF
C52107 PAND2X1_20/A POR2X1_35/CTRL 0.01fF
C52108 POR2X1_341/A POR2X1_325/A 0.04fF
C52109 POR2X1_614/A PAND2X1_255/O 0.08fF
C52110 PAND2X1_242/Y POR2X1_7/A 0.07fF
C52111 POR2X1_411/B PAND2X1_216/CTRL2 0.01fF
C52112 PAND2X1_222/A PAND2X1_593/CTRL 0.00fF
C52113 POR2X1_544/B POR2X1_325/B 0.08fF
C52114 POR2X1_461/Y POR2X1_790/CTRL 0.03fF
C52115 POR2X1_23/Y PAND2X1_332/CTRL 0.01fF
C52116 POR2X1_23/a_56_344# POR2X1_14/Y 0.01fF
C52117 PAND2X1_850/Y POR2X1_589/CTRL2 0.03fF
C52118 POR2X1_424/Y POR2X1_424/CTRL 0.00fF
C52119 POR2X1_43/B PAND2X1_449/CTRL2 0.01fF
C52120 POR2X1_83/B PAND2X1_215/a_16_344# 0.02fF
C52121 POR2X1_568/B PAND2X1_680/O 0.02fF
C52122 POR2X1_807/A POR2X1_807/O 0.09fF
C52123 POR2X1_150/Y POR2X1_42/Y 0.03fF
C52124 PAND2X1_838/CTRL2 POR2X1_42/Y 0.01fF
C52125 POR2X1_682/CTRL2 POR2X1_32/A 0.01fF
C52126 POR2X1_65/A POR2X1_283/O 0.01fF
C52127 POR2X1_56/B PAND2X1_796/B 0.02fF
C52128 POR2X1_130/A POR2X1_866/A 0.03fF
C52129 PAND2X1_71/Y PAND2X1_72/A 0.02fF
C52130 PAND2X1_415/O POR2X1_293/Y 0.03fF
C52131 PAND2X1_73/Y POR2X1_456/CTRL2 0.01fF
C52132 POR2X1_56/B PAND2X1_454/B 0.03fF
C52133 PAND2X1_52/CTRL POR2X1_532/A 0.01fF
C52134 POR2X1_14/Y POR2X1_72/B 0.03fF
C52135 PAND2X1_20/A POR2X1_500/A 0.06fF
C52136 POR2X1_257/A PAND2X1_213/A 0.00fF
C52137 POR2X1_274/Y POR2X1_296/B 0.03fF
C52138 POR2X1_411/B PAND2X1_218/O 0.03fF
C52139 POR2X1_150/Y POR2X1_309/Y 0.06fF
C52140 PAND2X1_453/A POR2X1_72/B 0.03fF
C52141 PAND2X1_790/CTRL POR2X1_42/Y 0.05fF
C52142 PAND2X1_58/A POR2X1_543/A 0.46fF
C52143 POR2X1_66/B POR2X1_461/CTRL2 0.00fF
C52144 POR2X1_411/B POR2X1_234/O 0.01fF
C52145 POR2X1_814/B PAND2X1_585/CTRL2 0.01fF
C52146 POR2X1_451/CTRL POR2X1_750/B 0.01fF
C52147 POR2X1_37/Y POR2X1_609/A 0.00fF
C52148 PAND2X1_223/CTRL POR2X1_283/Y 0.01fF
C52149 PAND2X1_651/Y POR2X1_490/CTRL 0.01fF
C52150 POR2X1_120/CTRL2 POR2X1_78/A 0.01fF
C52151 PAND2X1_76/Y POR2X1_102/Y 0.03fF
C52152 PAND2X1_117/CTRL2 POR2X1_558/B 0.00fF
C52153 POR2X1_496/Y VDD 3.22fF
C52154 PAND2X1_84/Y POR2X1_32/A 0.03fF
C52155 POR2X1_448/O PAND2X1_90/Y 0.02fF
C52156 POR2X1_555/A PAND2X1_626/O 0.05fF
C52157 POR2X1_467/Y POR2X1_448/Y 0.03fF
C52158 POR2X1_631/CTRL POR2X1_193/Y 0.02fF
C52159 PAND2X1_658/CTRL PAND2X1_474/A 0.01fF
C52160 POR2X1_16/A POR2X1_827/O 0.05fF
C52161 PAND2X1_239/O POR2X1_578/Y 0.05fF
C52162 POR2X1_687/A POR2X1_814/A 0.02fF
C52163 POR2X1_841/a_76_344# POR2X1_804/A 0.03fF
C52164 POR2X1_29/A POR2X1_546/A 0.03fF
C52165 POR2X1_224/O POR2X1_32/A 0.01fF
C52166 POR2X1_78/B POR2X1_811/B 0.03fF
C52167 PAND2X1_462/B POR2X1_48/A 0.12fF
C52168 POR2X1_800/CTRL D_GATE_865 0.01fF
C52169 POR2X1_68/Y PAND2X1_69/A 0.04fF
C52170 POR2X1_16/A PAND2X1_439/O 0.04fF
C52171 POR2X1_193/A POR2X1_218/Y 0.17fF
C52172 POR2X1_814/A POR2X1_772/CTRL 0.01fF
C52173 POR2X1_148/CTRL PAND2X1_69/A 0.01fF
C52174 POR2X1_457/O POR2X1_457/B 0.04fF
C52175 PAND2X1_660/CTRL PAND2X1_660/B 0.01fF
C52176 POR2X1_857/O POR2X1_192/Y 0.09fF
C52177 POR2X1_490/Y PAND2X1_716/O 0.01fF
C52178 PAND2X1_754/O POR2X1_29/A 0.02fF
C52179 POR2X1_751/A POR2X1_7/B 0.03fF
C52180 POR2X1_23/Y PAND2X1_725/A 0.01fF
C52181 POR2X1_695/Y PAND2X1_707/Y 0.35fF
C52182 POR2X1_590/A POR2X1_208/CTRL2 0.00fF
C52183 POR2X1_302/O POR2X1_330/Y 0.31fF
C52184 POR2X1_582/O POR2X1_582/Y 0.01fF
C52185 POR2X1_462/B POR2X1_862/A 0.01fF
C52186 PAND2X1_863/B POR2X1_102/Y 0.03fF
C52187 POR2X1_48/O POR2X1_72/B 0.01fF
C52188 POR2X1_218/Y POR2X1_572/B 0.06fF
C52189 PAND2X1_65/B PAND2X1_423/CTRL 0.01fF
C52190 PAND2X1_44/CTRL VDD 0.00fF
C52191 PAND2X1_827/m4_208_n4# POR2X1_740/Y 0.06fF
C52192 POR2X1_669/B POR2X1_615/Y 0.03fF
C52193 POR2X1_96/A POR2X1_60/A 0.51fF
C52194 PAND2X1_733/A VDD 0.29fF
C52195 POR2X1_458/CTRL2 PAND2X1_69/A 0.01fF
C52196 PAND2X1_247/CTRL POR2X1_283/A 0.01fF
C52197 POR2X1_859/A PAND2X1_225/O 0.02fF
C52198 POR2X1_23/Y PAND2X1_457/CTRL 0.01fF
C52199 PAND2X1_241/CTRL2 POR2X1_83/B 0.06fF
C52200 POR2X1_67/Y PAND2X1_789/O 0.02fF
C52201 PAND2X1_48/B POR2X1_174/A 0.02fF
C52202 POR2X1_143/CTRL2 POR2X1_40/Y 0.03fF
C52203 POR2X1_480/A POR2X1_286/Y 0.01fF
C52204 PAND2X1_640/CTRL2 D_INPUT_0 0.09fF
C52205 PAND2X1_58/A PAND2X1_369/CTRL2 0.01fF
C52206 POR2X1_57/A PAND2X1_212/O 0.01fF
C52207 PAND2X1_41/B PAND2X1_8/Y 6.35fF
C52208 PAND2X1_20/A POR2X1_128/a_76_344# 0.00fF
C52209 D_INPUT_0 PAND2X1_6/A 0.61fF
C52210 PAND2X1_7/CTRL POR2X1_555/B 0.01fF
C52211 POR2X1_630/CTRL PAND2X1_96/B 0.01fF
C52212 PAND2X1_649/CTRL POR2X1_32/A 0.01fF
C52213 POR2X1_788/A PAND2X1_144/CTRL2 0.01fF
C52214 POR2X1_47/CTRL POR2X1_83/B 0.01fF
C52215 POR2X1_278/Y PAND2X1_349/B 0.34fF
C52216 PAND2X1_95/B PAND2X1_11/Y 0.13fF
C52217 POR2X1_240/a_76_344# PAND2X1_88/Y 0.00fF
C52218 POR2X1_13/A PAND2X1_140/CTRL 0.01fF
C52219 POR2X1_655/A POR2X1_307/A 0.01fF
C52220 POR2X1_639/A VDD 0.00fF
C52221 POR2X1_558/B PAND2X1_96/B 0.03fF
C52222 POR2X1_629/B POR2X1_294/B 0.05fF
C52223 POR2X1_411/B PAND2X1_348/O 0.04fF
C52224 PAND2X1_73/Y PAND2X1_744/CTRL2 0.01fF
C52225 POR2X1_848/A POR2X1_93/A 0.08fF
C52226 POR2X1_55/CTRL PAND2X1_6/A 0.03fF
C52227 POR2X1_300/O POR2X1_102/Y 0.01fF
C52228 POR2X1_37/Y POR2X1_380/a_76_344# 0.01fF
C52229 POR2X1_49/Y PAND2X1_479/B 0.00fF
C52230 POR2X1_433/Y POR2X1_432/O 0.01fF
C52231 PAND2X1_512/Y POR2X1_5/Y 0.03fF
C52232 PAND2X1_276/CTRL VDD 0.00fF
C52233 PAND2X1_776/Y POR2X1_91/Y 0.00fF
C52234 PAND2X1_48/B PAND2X1_15/a_76_28# 0.02fF
C52235 PAND2X1_94/A PAND2X1_24/CTRL2 0.00fF
C52236 PAND2X1_309/CTRL2 POR2X1_543/A 0.01fF
C52237 POR2X1_12/O POR2X1_13/A 0.01fF
C52238 POR2X1_38/Y POR2X1_37/Y 0.11fF
C52239 POR2X1_504/CTRL POR2X1_20/B 0.01fF
C52240 POR2X1_117/CTRL POR2X1_46/Y 0.00fF
C52241 POR2X1_251/A POR2X1_55/Y 0.05fF
C52242 POR2X1_462/B PAND2X1_73/Y 0.03fF
C52243 POR2X1_128/A POR2X1_128/a_16_28# 0.03fF
C52244 POR2X1_32/A POR2X1_594/A 0.02fF
C52245 POR2X1_72/B POR2X1_55/Y 0.13fF
C52246 PAND2X1_73/Y D_INPUT_1 0.16fF
C52247 PAND2X1_558/Y PAND2X1_717/CTRL2 0.00fF
C52248 POR2X1_558/A POR2X1_558/B 0.02fF
C52249 POR2X1_49/Y PAND2X1_466/CTRL 0.02fF
C52250 PAND2X1_849/B POR2X1_813/a_16_28# 0.07fF
C52251 POR2X1_72/O POR2X1_71/Y 0.03fF
C52252 POR2X1_68/A POR2X1_864/O 0.04fF
C52253 POR2X1_272/Y PAND2X1_785/Y 0.03fF
C52254 PAND2X1_792/a_76_28# POR2X1_759/Y 0.03fF
C52255 PAND2X1_587/Y VDD 0.16fF
C52256 POR2X1_231/A POR2X1_785/A 0.01fF
C52257 PAND2X1_482/O POR2X1_541/B 0.09fF
C52258 PAND2X1_568/CTRL VDD 0.00fF
C52259 POR2X1_233/O POR2X1_236/Y 0.01fF
C52260 PAND2X1_73/Y POR2X1_724/A 0.01fF
C52261 POR2X1_305/Y POR2X1_40/Y 0.04fF
C52262 POR2X1_614/A POR2X1_800/CTRL 0.01fF
C52263 PAND2X1_6/Y POR2X1_605/B 0.10fF
C52264 POR2X1_188/A POR2X1_114/B 0.01fF
C52265 PAND2X1_804/B VDD 0.02fF
C52266 POR2X1_866/A POR2X1_596/CTRL 0.12fF
C52267 PAND2X1_469/B POR2X1_423/Y 0.05fF
C52268 POR2X1_48/A POR2X1_766/O 0.01fF
C52269 PAND2X1_684/CTRL POR2X1_260/B 0.01fF
C52270 PAND2X1_3/CTRL PAND2X1_3/A 0.01fF
C52271 POR2X1_309/CTRL POR2X1_387/Y 0.07fF
C52272 POR2X1_49/Y POR2X1_521/CTRL 0.01fF
C52273 POR2X1_319/A POR2X1_704/Y 0.00fF
C52274 POR2X1_332/Y POR2X1_341/A 1.07fF
C52275 PAND2X1_73/O PAND2X1_69/A 0.01fF
C52276 POR2X1_66/B POR2X1_649/B 0.12fF
C52277 PAND2X1_44/CTRL PAND2X1_32/B 0.01fF
C52278 POR2X1_78/B POR2X1_783/B 0.02fF
C52279 POR2X1_83/B PAND2X1_168/CTRL2 0.03fF
C52280 PAND2X1_272/CTRL POR2X1_569/A 0.02fF
C52281 POR2X1_493/B POR2X1_558/B 0.00fF
C52282 PAND2X1_116/CTRL2 POR2X1_183/Y 0.00fF
C52283 D_INPUT_0 POR2X1_101/Y 0.05fF
C52284 POR2X1_231/B VDD 0.04fF
C52285 POR2X1_79/Y PAND2X1_735/Y 0.17fF
C52286 PAND2X1_499/a_76_28# POR2X1_293/Y 0.01fF
C52287 PAND2X1_731/CTRL2 PAND2X1_738/B 0.00fF
C52288 POR2X1_16/A POR2X1_48/A 0.13fF
C52289 POR2X1_449/O POR2X1_832/B 0.00fF
C52290 POR2X1_614/A POR2X1_801/O 0.01fF
C52291 POR2X1_296/B PAND2X1_63/B 0.10fF
C52292 POR2X1_378/O D_INPUT_1 0.01fF
C52293 POR2X1_72/B PAND2X1_186/CTRL 0.02fF
C52294 PAND2X1_840/A PAND2X1_499/O 0.04fF
C52295 PAND2X1_724/O POR2X1_40/Y 0.05fF
C52296 POR2X1_66/A POR2X1_773/B 0.00fF
C52297 D_INPUT_0 PAND2X1_690/CTRL2 0.00fF
C52298 POR2X1_502/A POR2X1_776/B 0.02fF
C52299 POR2X1_78/A POR2X1_854/B 0.03fF
C52300 POR2X1_846/A PAND2X1_52/B 1.01fF
C52301 INPUT_1 POR2X1_37/Y 0.57fF
C52302 PAND2X1_52/Y POR2X1_631/B 0.10fF
C52303 POR2X1_858/B POR2X1_858/O 0.00fF
C52304 POR2X1_57/A PAND2X1_731/B 0.03fF
C52305 POR2X1_68/A D_GATE_865 0.04fF
C52306 POR2X1_83/A POR2X1_397/Y 0.01fF
C52307 PAND2X1_341/O INPUT_0 0.09fF
C52308 POR2X1_60/A POR2X1_7/A 1.97fF
C52309 PAND2X1_514/Y VDD 0.18fF
C52310 PAND2X1_96/B POR2X1_543/A 0.03fF
C52311 POR2X1_840/B POR2X1_660/A 0.16fF
C52312 PAND2X1_58/A PAND2X1_28/CTRL 0.06fF
C52313 PAND2X1_264/O POR2X1_669/B 0.28fF
C52314 POR2X1_65/A PAND2X1_724/CTRL 0.01fF
C52315 PAND2X1_232/m4_208_n4# POR2X1_66/A 0.08fF
C52316 PAND2X1_654/O POR2X1_13/A 0.06fF
C52317 PAND2X1_495/CTRL POR2X1_814/B 0.00fF
C52318 POR2X1_356/A PAND2X1_524/a_16_344# 0.04fF
C52319 POR2X1_460/B VDD 0.02fF
C52320 POR2X1_829/A POR2X1_597/A 0.86fF
C52321 PAND2X1_97/a_16_344# POR2X1_153/Y 0.05fF
C52322 POR2X1_66/B POR2X1_222/A 0.03fF
C52323 POR2X1_174/B POR2X1_502/CTRL2 0.15fF
C52324 PAND2X1_6/Y PAND2X1_627/CTRL 0.01fF
C52325 POR2X1_68/A POR2X1_471/CTRL 0.01fF
C52326 POR2X1_730/Y POR2X1_590/A 0.03fF
C52327 POR2X1_596/A PAND2X1_597/CTRL 0.01fF
C52328 POR2X1_278/Y PAND2X1_652/A 0.07fF
C52329 PAND2X1_56/Y POR2X1_244/B 0.11fF
C52330 POR2X1_612/a_16_28# POR2X1_4/Y 0.02fF
C52331 PAND2X1_192/Y PAND2X1_739/B 0.12fF
C52332 POR2X1_327/Y PAND2X1_431/a_16_344# 0.04fF
C52333 POR2X1_37/Y POR2X1_153/Y 0.61fF
C52334 POR2X1_790/A VDD 0.64fF
C52335 POR2X1_480/A PAND2X1_69/A 0.07fF
C52336 PAND2X1_94/A PAND2X1_235/CTRL 0.01fF
C52337 POR2X1_37/Y POR2X1_384/A 0.03fF
C52338 POR2X1_648/Y PAND2X1_72/A 0.03fF
C52339 POR2X1_158/CTRL POR2X1_257/A 0.01fF
C52340 PAND2X1_776/Y POR2X1_109/Y 0.03fF
C52341 POR2X1_52/A PAND2X1_717/CTRL 0.01fF
C52342 POR2X1_390/B POR2X1_105/O 0.00fF
C52343 PAND2X1_624/A PAND2X1_623/Y 0.01fF
C52344 POR2X1_814/A POR2X1_568/A 0.41fF
C52345 POR2X1_113/Y POR2X1_475/A 0.07fF
C52346 POR2X1_43/B POR2X1_46/Y 0.16fF
C52347 POR2X1_811/CTRL2 POR2X1_294/A 0.05fF
C52348 POR2X1_230/CTRL PAND2X1_338/B 0.03fF
C52349 PAND2X1_864/CTRL PAND2X1_810/A 0.01fF
C52350 POR2X1_130/A POR2X1_501/B 0.07fF
C52351 PAND2X1_309/O POR2X1_741/Y 0.03fF
C52352 PAND2X1_587/Y PAND2X1_32/B 0.03fF
C52353 POR2X1_243/Y PAND2X1_69/A 0.07fF
C52354 PAND2X1_96/B PAND2X1_516/CTRL2 0.01fF
C52355 POR2X1_219/B POR2X1_215/O 0.02fF
C52356 POR2X1_567/B POR2X1_726/O 0.02fF
C52357 VDD PAND2X1_88/Y 1.00fF
C52358 POR2X1_406/Y POR2X1_38/Y 0.02fF
C52359 POR2X1_865/B VDD 0.42fF
C52360 POR2X1_127/a_16_28# POR2X1_394/A 0.01fF
C52361 POR2X1_68/A POR2X1_579/Y 0.03fF
C52362 POR2X1_332/B PAND2X1_96/B 0.07fF
C52363 POR2X1_84/Y VDD 0.14fF
C52364 POR2X1_705/B PAND2X1_52/B 0.03fF
C52365 POR2X1_483/A POR2X1_228/Y 0.06fF
C52366 POR2X1_66/A POR2X1_195/a_16_28# 0.02fF
C52367 POR2X1_65/A POR2X1_527/CTRL2 0.09fF
C52368 POR2X1_119/Y D_INPUT_0 0.17fF
C52369 POR2X1_327/CTRL PAND2X1_63/Y 0.03fF
C52370 PAND2X1_738/Y PAND2X1_388/O 0.10fF
C52371 PAND2X1_48/B PAND2X1_146/a_16_344# 0.01fF
C52372 POR2X1_215/a_56_344# PAND2X1_88/Y 0.00fF
C52373 POR2X1_57/A POR2X1_51/A 0.02fF
C52374 PAND2X1_349/A POR2X1_236/Y 0.03fF
C52375 POR2X1_859/A POR2X1_750/CTRL 0.03fF
C52376 POR2X1_124/a_56_344# POR2X1_124/B 0.00fF
C52377 PAND2X1_63/B POR2X1_236/Y 0.05fF
C52378 POR2X1_231/B PAND2X1_32/B 0.04fF
C52379 PAND2X1_682/CTRL2 POR2X1_407/A 0.02fF
C52380 POR2X1_854/CTRL2 POR2X1_192/Y 0.01fF
C52381 POR2X1_392/O PAND2X1_32/B 0.01fF
C52382 POR2X1_845/A POR2X1_78/A 0.01fF
C52383 PAND2X1_64/CTRL2 D_INPUT_4 0.00fF
C52384 PAND2X1_90/A PAND2X1_69/A 8.54fF
C52385 POR2X1_68/A POR2X1_545/A 0.04fF
C52386 INPUT_2 POR2X1_119/O 0.01fF
C52387 POR2X1_475/A POR2X1_260/A 0.03fF
C52388 POR2X1_38/Y POR2X1_293/Y 2.71fF
C52389 POR2X1_556/A PAND2X1_135/CTRL 0.00fF
C52390 POR2X1_537/Y POR2X1_121/B 0.03fF
C52391 POR2X1_525/O PAND2X1_726/B 0.02fF
C52392 PAND2X1_484/CTRL2 PAND2X1_41/B 0.09fF
C52393 PAND2X1_654/a_16_344# PAND2X1_651/Y 0.09fF
C52394 POR2X1_492/CTRL POR2X1_394/A 0.06fF
C52395 POR2X1_516/CTRL PAND2X1_6/A 0.05fF
C52396 POR2X1_16/A PAND2X1_199/A 0.01fF
C52397 PAND2X1_353/CTRL VDD -0.00fF
C52398 POR2X1_49/Y POR2X1_177/CTRL2 0.03fF
C52399 POR2X1_241/B POR2X1_191/Y 0.05fF
C52400 PAND2X1_794/B PAND2X1_357/Y 0.03fF
C52401 POR2X1_383/A POR2X1_244/B 0.03fF
C52402 INPUT_0 POR2X1_569/A 0.07fF
C52403 POR2X1_7/A PAND2X1_515/CTRL2 0.01fF
C52404 POR2X1_62/Y POR2X1_69/A 0.03fF
C52405 POR2X1_416/Y PAND2X1_472/A 0.01fF
C52406 POR2X1_840/O PAND2X1_55/Y 0.18fF
C52407 POR2X1_809/A POR2X1_864/a_56_344# 0.00fF
C52408 POR2X1_614/A POR2X1_68/A 6.86fF
C52409 PAND2X1_351/Y PAND2X1_656/A 0.00fF
C52410 PAND2X1_344/CTRL2 PAND2X1_514/Y 0.03fF
C52411 POR2X1_78/A POR2X1_374/CTRL2 0.00fF
C52412 POR2X1_460/B PAND2X1_32/B 0.03fF
C52413 POR2X1_712/A POR2X1_407/A 0.05fF
C52414 POR2X1_567/A POR2X1_629/B 0.05fF
C52415 PAND2X1_467/Y PAND2X1_707/CTRL 0.01fF
C52416 PAND2X1_290/O POR2X1_66/A 0.04fF
C52417 PAND2X1_480/CTRL2 POR2X1_236/Y 0.01fF
C52418 POR2X1_164/CTRL PAND2X1_565/A 0.00fF
C52419 POR2X1_63/a_16_28# POR2X1_43/B 0.02fF
C52420 POR2X1_327/Y POR2X1_807/A 0.03fF
C52421 POR2X1_355/B POR2X1_180/A 0.03fF
C52422 POR2X1_790/A PAND2X1_32/B 0.03fF
C52423 POR2X1_741/Y PAND2X1_88/Y 0.03fF
C52424 PAND2X1_602/Y PAND2X1_648/O 0.04fF
C52425 PAND2X1_376/O VDD 0.00fF
C52426 POR2X1_278/O PAND2X1_560/B 0.02fF
C52427 POR2X1_72/B PAND2X1_199/B 0.04fF
C52428 POR2X1_68/A POR2X1_38/B 0.07fF
C52429 POR2X1_283/A POR2X1_7/B 5.51fF
C52430 PAND2X1_319/B PAND2X1_675/A 0.07fF
C52431 PAND2X1_651/Y POR2X1_239/CTRL 0.00fF
C52432 PAND2X1_824/B POR2X1_207/CTRL2 0.06fF
C52433 PAND2X1_81/B POR2X1_84/Y 0.07fF
C52434 POR2X1_276/A POR2X1_276/CTRL 0.04fF
C52435 POR2X1_566/A POR2X1_703/A 0.07fF
C52436 POR2X1_51/A POR2X1_744/O 0.01fF
C52437 PAND2X1_319/B PAND2X1_469/B 0.05fF
C52438 PAND2X1_101/O PAND2X1_99/Y 0.04fF
C52439 POR2X1_66/B PAND2X1_665/CTRL2 0.00fF
C52440 PAND2X1_94/A PAND2X1_92/O 0.05fF
C52441 POR2X1_590/A POR2X1_532/a_56_344# 0.03fF
C52442 POR2X1_850/A POR2X1_737/A 0.00fF
C52443 POR2X1_29/Y POR2X1_409/a_16_28# 0.02fF
C52444 POR2X1_13/A PAND2X1_777/CTRL2 0.00fF
C52445 POR2X1_327/CTRL POR2X1_260/A 0.01fF
C52446 POR2X1_68/A PAND2X1_422/O 0.01fF
C52447 POR2X1_865/B PAND2X1_32/B 0.03fF
C52448 POR2X1_501/B POR2X1_573/A 0.12fF
C52449 POR2X1_349/Y POR2X1_363/A 0.01fF
C52450 POR2X1_272/Y POR2X1_300/Y 0.01fF
C52451 POR2X1_863/B POR2X1_260/A 0.01fF
C52452 POR2X1_41/B POR2X1_8/Y 0.07fF
C52453 INPUT_1 POR2X1_293/Y 0.27fF
C52454 POR2X1_201/Y POR2X1_35/Y 0.01fF
C52455 POR2X1_510/A POR2X1_854/B 0.37fF
C52456 PAND2X1_357/Y POR2X1_107/Y 0.00fF
C52457 POR2X1_814/B POR2X1_703/m4_208_n4# 0.01fF
C52458 POR2X1_42/Y PAND2X1_154/a_76_28# 0.02fF
C52459 POR2X1_75/Y VDD 0.03fF
C52460 POR2X1_662/Y POR2X1_456/B 0.03fF
C52461 PAND2X1_686/CTRL POR2X1_42/Y 0.01fF
C52462 POR2X1_614/A PAND2X1_315/CTRL2 0.01fF
C52463 POR2X1_74/Y PAND2X1_76/Y 0.26fF
C52464 PAND2X1_6/Y POR2X1_855/B 0.01fF
C52465 POR2X1_96/A POR2X1_96/a_16_28# 0.01fF
C52466 POR2X1_81/CTRL PAND2X1_862/B 0.01fF
C52467 POR2X1_16/A PAND2X1_401/CTRL 0.00fF
C52468 PAND2X1_702/CTRL2 POR2X1_7/A 0.03fF
C52469 PAND2X1_54/CTRL2 POR2X1_4/Y 0.02fF
C52470 PAND2X1_564/m4_208_n4# POR2X1_766/m4_208_n4# 0.13fF
C52471 PAND2X1_96/B POR2X1_574/A 0.52fF
C52472 PAND2X1_858/CTRL POR2X1_13/A 0.01fF
C52473 POR2X1_287/B PAND2X1_122/O 0.02fF
C52474 POR2X1_13/A PAND2X1_345/Y 0.00fF
C52475 POR2X1_293/Y POR2X1_153/Y 5.62fF
C52476 POR2X1_508/A VDD 0.11fF
C52477 PAND2X1_797/Y PAND2X1_803/A -0.00fF
C52478 POR2X1_407/A POR2X1_407/O 0.17fF
C52479 POR2X1_38/Y POR2X1_408/Y 0.12fF
C52480 POR2X1_180/B POR2X1_614/A 0.03fF
C52481 PAND2X1_90/Y POR2X1_542/CTRL2 0.17fF
C52482 POR2X1_502/A PAND2X1_48/A 0.13fF
C52483 POR2X1_495/O POR2X1_39/B 0.01fF
C52484 PAND2X1_474/Y PAND2X1_500/CTRL2 0.00fF
C52485 POR2X1_731/O POR2X1_738/A 0.16fF
C52486 PAND2X1_143/CTRL PAND2X1_8/Y 0.01fF
C52487 POR2X1_218/A POR2X1_260/A 0.07fF
C52488 POR2X1_502/A POR2X1_192/B 0.14fF
C52489 POR2X1_865/CTRL POR2X1_101/Y 0.03fF
C52490 POR2X1_375/CTRL PAND2X1_32/B 0.01fF
C52491 POR2X1_341/Y POR2X1_351/O 0.01fF
C52492 POR2X1_130/CTRL PAND2X1_6/Y 0.01fF
C52493 POR2X1_389/A POR2X1_725/Y 0.18fF
C52494 POR2X1_283/A POR2X1_248/a_16_28# 0.02fF
C52495 POR2X1_346/B PAND2X1_69/A 0.03fF
C52496 POR2X1_355/B POR2X1_508/B 0.11fF
C52497 POR2X1_783/B POR2X1_294/A 0.03fF
C52498 POR2X1_653/B POR2X1_711/Y 0.02fF
C52499 PAND2X1_140/A POR2X1_107/Y 0.01fF
C52500 PAND2X1_837/O POR2X1_826/Y 0.00fF
C52501 POR2X1_124/B POR2X1_768/O 0.01fF
C52502 POR2X1_830/A POR2X1_711/Y 0.07fF
C52503 PAND2X1_4/CTRL2 POR2X1_260/A 0.03fF
C52504 PAND2X1_90/A PAND2X1_384/m4_208_n4# 0.20fF
C52505 POR2X1_327/Y POR2X1_407/A 0.03fF
C52506 POR2X1_216/CTRL POR2X1_276/Y 0.01fF
C52507 PAND2X1_699/CTRL POR2X1_628/Y 0.00fF
C52508 PAND2X1_452/B VDD 0.02fF
C52509 PAND2X1_65/B PAND2X1_56/A 0.15fF
C52510 VDD POR2X1_568/B 9.28fF
C52511 POR2X1_407/Y POR2X1_596/a_56_344# 0.00fF
C52512 PAND2X1_217/B PAND2X1_332/Y 0.03fF
C52513 POR2X1_112/O POR2X1_579/Y 0.00fF
C52514 PAND2X1_482/CTRL POR2X1_786/Y 0.05fF
C52515 PAND2X1_56/Y POR2X1_537/Y 0.05fF
C52516 POR2X1_416/B PAND2X1_723/Y 0.02fF
C52517 PAND2X1_691/Y PAND2X1_854/A 0.14fF
C52518 PAND2X1_354/O PAND2X1_354/Y 0.00fF
C52519 PAND2X1_390/Y POR2X1_589/Y 0.04fF
C52520 POR2X1_711/B POR2X1_710/CTRL2 0.03fF
C52521 POR2X1_43/O VDD 0.00fF
C52522 PAND2X1_847/m4_208_n4# POR2X1_4/Y 0.07fF
C52523 POR2X1_861/A POR2X1_572/B 0.10fF
C52524 POR2X1_852/B POR2X1_568/A 0.54fF
C52525 PAND2X1_798/Y POR2X1_79/Y 0.01fF
C52526 POR2X1_416/B PAND2X1_347/Y 0.03fF
C52527 INPUT_1 POR2X1_408/Y 0.04fF
C52528 POR2X1_527/O PAND2X1_549/B 0.01fF
C52529 POR2X1_356/A POR2X1_510/CTRL 0.16fF
C52530 POR2X1_837/A POR2X1_296/B 0.03fF
C52531 POR2X1_54/Y POR2X1_859/O 0.01fF
C52532 PAND2X1_563/A PAND2X1_348/Y 0.03fF
C52533 POR2X1_88/Y POR2X1_77/Y 0.03fF
C52534 POR2X1_461/B PAND2X1_52/B 0.02fF
C52535 POR2X1_809/A POR2X1_596/A 0.02fF
C52536 POR2X1_27/CTRL2 POR2X1_669/B 0.01fF
C52537 POR2X1_466/A POR2X1_466/a_16_28# 0.01fF
C52538 POR2X1_675/Y POR2X1_737/CTRL 0.01fF
C52539 POR2X1_113/Y POR2X1_557/B 0.01fF
C52540 POR2X1_271/A PAND2X1_349/A 0.03fF
C52541 INPUT_0 PAND2X1_72/A 0.05fF
C52542 PAND2X1_425/Y PAND2X1_581/O 0.02fF
C52543 VDD PAND2X1_332/Y 0.57fF
C52544 POR2X1_360/a_76_344# POR2X1_244/Y 0.01fF
C52545 PAND2X1_404/Y POR2X1_411/B 0.03fF
C52546 POR2X1_385/Y PAND2X1_389/a_56_28# 0.00fF
C52547 PAND2X1_800/CTRL2 PAND2X1_691/Y 0.00fF
C52548 POR2X1_305/CTRL POR2X1_55/Y 0.01fF
C52549 PAND2X1_717/Y POR2X1_394/A 0.07fF
C52550 PAND2X1_453/O POR2X1_77/Y 0.01fF
C52551 POR2X1_582/Y POR2X1_428/Y 0.08fF
C52552 POR2X1_510/Y POR2X1_553/a_76_344# 0.01fF
C52553 POR2X1_343/Y POR2X1_575/B 0.02fF
C52554 PAND2X1_96/B PAND2X1_759/CTRL 0.01fF
C52555 POR2X1_614/A POR2X1_181/O 0.09fF
C52556 PAND2X1_351/O PAND2X1_351/A 0.02fF
C52557 POR2X1_860/O POR2X1_244/Y 0.18fF
C52558 POR2X1_319/A POR2X1_446/B 0.05fF
C52559 POR2X1_614/A POR2X1_169/A 0.03fF
C52560 POR2X1_317/Y POR2X1_169/A 0.02fF
C52561 POR2X1_537/Y POR2X1_383/A 0.03fF
C52562 POR2X1_677/Y PAND2X1_76/Y 0.03fF
C52563 POR2X1_376/B PAND2X1_635/Y 0.03fF
C52564 POR2X1_14/CTRL2 INPUT_3 0.01fF
C52565 PAND2X1_39/B POR2X1_678/Y 0.07fF
C52566 POR2X1_568/B PAND2X1_32/B 0.03fF
C52567 POR2X1_416/B POR2X1_628/a_16_28# 0.03fF
C52568 POR2X1_557/B POR2X1_260/A 0.03fF
C52569 POR2X1_471/A POR2X1_66/A 0.03fF
C52570 PAND2X1_3/O PAND2X1_3/B -0.00fF
C52571 PAND2X1_682/CTRL POR2X1_728/A 0.00fF
C52572 POR2X1_666/CTRL2 POR2X1_411/B 0.01fF
C52573 PAND2X1_476/A POR2X1_235/O 0.00fF
C52574 POR2X1_54/Y PAND2X1_68/CTRL2 0.09fF
C52575 PAND2X1_762/Y PAND2X1_52/B 0.04fF
C52576 POR2X1_137/B PAND2X1_73/Y 0.07fF
C52577 PAND2X1_94/A PAND2X1_527/O 0.04fF
C52578 POR2X1_16/A POR2X1_62/Y 0.04fF
C52579 POR2X1_294/Y POR2X1_294/O 0.00fF
C52580 POR2X1_438/O POR2X1_77/Y 0.02fF
C52581 PAND2X1_611/CTRL2 POR2X1_389/Y 0.00fF
C52582 POR2X1_309/O POR2X1_411/B 0.01fF
C52583 POR2X1_23/Y PAND2X1_477/CTRL 0.10fF
C52584 POR2X1_260/B POR2X1_734/B 0.04fF
C52585 PAND2X1_388/Y POR2X1_39/B 0.03fF
C52586 PAND2X1_483/CTRL PAND2X1_631/A 0.01fF
C52587 PAND2X1_483/O POR2X1_252/Y 0.02fF
C52588 POR2X1_65/A POR2X1_65/O 0.00fF
C52589 POR2X1_67/Y PAND2X1_381/O 0.02fF
C52590 PAND2X1_466/A POR2X1_423/Y 0.10fF
C52591 POR2X1_556/A POR2X1_269/Y 0.01fF
C52592 PAND2X1_549/B POR2X1_39/B 0.03fF
C52593 POR2X1_14/Y PAND2X1_407/CTRL2 0.03fF
C52594 PAND2X1_618/Y POR2X1_29/A 0.04fF
C52595 POR2X1_52/A PAND2X1_635/Y 0.01fF
C52596 POR2X1_728/CTRL POR2X1_814/A 0.06fF
C52597 POR2X1_78/A POR2X1_862/A 0.03fF
C52598 POR2X1_602/B PAND2X1_39/B 0.10fF
C52599 PAND2X1_93/B PAND2X1_73/Y 0.10fF
C52600 PAND2X1_260/O POR2X1_257/A 0.08fF
C52601 POR2X1_411/A POR2X1_236/Y 0.01fF
C52602 POR2X1_863/A POR2X1_570/B 6.09fF
C52603 PAND2X1_221/Y PAND2X1_357/Y 0.00fF
C52604 PAND2X1_57/B PAND2X1_45/CTRL2 0.03fF
C52605 POR2X1_416/B PAND2X1_346/Y 0.01fF
C52606 POR2X1_855/B PAND2X1_52/B 0.03fF
C52607 PAND2X1_10/CTRL2 POR2X1_296/B 0.01fF
C52608 PAND2X1_472/O POR2X1_39/B 0.01fF
C52609 POR2X1_23/Y PAND2X1_573/B 0.03fF
C52610 PAND2X1_170/O PAND2X1_326/B 0.02fF
C52611 PAND2X1_677/O POR2X1_260/B 0.02fF
C52612 POR2X1_260/B POR2X1_330/Y 0.08fF
C52613 POR2X1_352/CTRL2 PAND2X1_52/B 0.03fF
C52614 PAND2X1_224/m4_208_n4# POR2X1_578/Y 0.05fF
C52615 PAND2X1_65/B POR2X1_818/O 0.01fF
C52616 POR2X1_416/B POR2X1_419/a_56_344# 0.00fF
C52617 PAND2X1_222/A POR2X1_250/A 0.03fF
C52618 POR2X1_8/Y POR2X1_77/Y 0.12fF
C52619 POR2X1_411/B PAND2X1_340/m4_208_n4# 0.07fF
C52620 POR2X1_383/A POR2X1_579/CTRL 0.08fF
C52621 POR2X1_352/CTRL2 POR2X1_212/B 0.03fF
C52622 POR2X1_499/A POR2X1_778/a_16_28# 0.03fF
C52623 PAND2X1_858/O PAND2X1_850/Y 0.12fF
C52624 POR2X1_801/A POR2X1_452/Y 0.17fF
C52625 PAND2X1_221/Y PAND2X1_365/a_76_28# 0.02fF
C52626 POR2X1_96/A POR2X1_329/Y 0.01fF
C52627 POR2X1_685/O POR2X1_452/Y 0.01fF
C52628 POR2X1_390/B POR2X1_717/B 0.03fF
C52629 PAND2X1_73/Y POR2X1_78/A 4.52fF
C52630 POR2X1_567/B POR2X1_436/O 0.01fF
C52631 POR2X1_341/A VDD 2.94fF
C52632 PAND2X1_273/O POR2X1_814/A 0.15fF
C52633 POR2X1_774/Y POR2X1_866/A 0.08fF
C52634 POR2X1_640/O POR2X1_66/A 0.02fF
C52635 PAND2X1_20/A POR2X1_29/A 0.03fF
C52636 POR2X1_502/A POR2X1_461/Y 0.03fF
C52637 POR2X1_48/A POR2X1_414/Y 0.45fF
C52638 POR2X1_809/B POR2X1_452/Y 0.01fF
C52639 POR2X1_416/B PAND2X1_123/Y 0.05fF
C52640 POR2X1_137/B PAND2X1_132/CTRL2 0.02fF
C52641 PAND2X1_405/CTRL POR2X1_38/Y 0.01fF
C52642 PAND2X1_847/O POR2X1_394/A 0.02fF
C52643 POR2X1_537/Y PAND2X1_108/CTRL2 0.01fF
C52644 POR2X1_8/Y POR2X1_8/O 0.01fF
C52645 POR2X1_115/CTRL2 POR2X1_446/B 0.01fF
C52646 POR2X1_176/O POR2X1_77/Y 0.18fF
C52647 POR2X1_39/B POR2X1_397/CTRL 0.01fF
C52648 PAND2X1_6/Y PAND2X1_32/O 0.02fF
C52649 POR2X1_311/Y POR2X1_60/A 0.03fF
C52650 POR2X1_9/Y POR2X1_245/O 0.07fF
C52651 POR2X1_78/A POR2X1_264/CTRL 0.02fF
C52652 POR2X1_566/A POR2X1_854/O 0.01fF
C52653 PAND2X1_231/O POR2X1_263/Y 0.02fF
C52654 POR2X1_564/B PAND2X1_52/B 0.11fF
C52655 POR2X1_840/B POR2X1_814/A 0.05fF
C52656 POR2X1_604/Y POR2X1_40/Y 0.01fF
C52657 POR2X1_345/A POR2X1_555/B 0.03fF
C52658 PAND2X1_839/O POR2X1_20/B 0.04fF
C52659 POR2X1_423/O POR2X1_423/Y 0.05fF
C52660 POR2X1_102/Y PAND2X1_558/Y 0.01fF
C52661 POR2X1_20/B POR2X1_619/CTRL 0.09fF
C52662 POR2X1_602/B PAND2X1_20/A 0.01fF
C52663 POR2X1_801/CTRL2 POR2X1_121/B -0.00fF
C52664 POR2X1_814/B POR2X1_29/A 0.12fF
C52665 POR2X1_263/Y POR2X1_230/a_76_344# 0.00fF
C52666 PAND2X1_51/O POR2X1_451/A 0.03fF
C52667 POR2X1_60/A PAND2X1_140/CTRL2 0.01fF
C52668 PAND2X1_407/CTRL2 POR2X1_55/Y 0.00fF
C52669 PAND2X1_624/CTRL2 POR2X1_29/A 0.01fF
C52670 POR2X1_788/A POR2X1_788/O 0.09fF
C52671 POR2X1_278/Y PAND2X1_205/A 0.13fF
C52672 POR2X1_394/A POR2X1_321/CTRL2 0.05fF
C52673 POR2X1_52/A PAND2X1_404/Y 0.03fF
C52674 POR2X1_341/A POR2X1_741/Y 0.07fF
C52675 PAND2X1_242/Y POR2X1_153/Y 0.10fF
C52676 POR2X1_624/Y POR2X1_575/B 0.08fF
C52677 POR2X1_817/CTRL2 POR2X1_817/A 0.01fF
C52678 PAND2X1_48/B POR2X1_446/B 0.04fF
C52679 PAND2X1_73/Y POR2X1_573/CTRL 0.01fF
C52680 POR2X1_776/A D_GATE_741 0.07fF
C52681 POR2X1_196/a_56_344# POR2X1_702/B 0.00fF
C52682 POR2X1_556/A POR2X1_513/Y 0.03fF
C52683 PAND2X1_81/B POR2X1_341/A 0.05fF
C52684 PAND2X1_99/B PAND2X1_99/CTRL2 0.01fF
C52685 POR2X1_32/A POR2X1_236/Y 0.21fF
C52686 POR2X1_458/Y PAND2X1_368/O 0.11fF
C52687 PAND2X1_631/O POR2X1_20/B 0.01fF
C52688 POR2X1_142/a_56_344# POR2X1_65/A 0.00fF
C52689 PAND2X1_39/B POR2X1_712/Y 0.03fF
C52690 POR2X1_257/A POR2X1_433/Y 0.03fF
C52691 POR2X1_40/Y POR2X1_503/A 0.01fF
C52692 POR2X1_54/Y PAND2X1_283/O 0.01fF
C52693 POR2X1_78/B POR2X1_296/B 0.11fF
C52694 PAND2X1_576/B PAND2X1_364/B 0.11fF
C52695 PAND2X1_492/CTRL POR2X1_78/A 0.01fF
C52696 PAND2X1_492/O PAND2X1_73/Y 0.05fF
C52697 POR2X1_65/A POR2X1_40/Y 3.68fF
C52698 POR2X1_227/B POR2X1_532/A 0.01fF
C52699 PAND2X1_61/CTRL2 POR2X1_58/Y 0.01fF
C52700 POR2X1_341/A PAND2X1_32/B 0.10fF
C52701 POR2X1_210/CTRL2 POR2X1_220/Y 0.00fF
C52702 POR2X1_865/B POR2X1_475/CTRL2 0.02fF
C52703 POR2X1_504/Y POR2X1_49/Y 0.03fF
C52704 POR2X1_638/CTRL POR2X1_66/A 0.01fF
C52705 POR2X1_451/A PAND2X1_3/B 0.04fF
C52706 POR2X1_484/Y POR2X1_526/Y 0.03fF
C52707 POR2X1_674/Y VDD 0.00fF
C52708 POR2X1_78/B POR2X1_605/O 0.08fF
C52709 PAND2X1_93/B PAND2X1_144/CTRL 0.01fF
C52710 POR2X1_22/A POR2X1_260/B 0.04fF
C52711 PAND2X1_9/Y POR2X1_84/Y 0.27fF
C52712 POR2X1_730/Y POR2X1_440/B 0.00fF
C52713 PAND2X1_206/B PAND2X1_100/O 0.00fF
C52714 PAND2X1_48/B PAND2X1_485/a_76_28# 0.02fF
C52715 PAND2X1_480/B POR2X1_102/Y 0.06fF
C52716 POR2X1_417/Y POR2X1_236/Y 0.03fF
C52717 POR2X1_429/CTRL2 VDD 0.00fF
C52718 POR2X1_48/A PAND2X1_324/Y 0.01fF
C52719 PAND2X1_20/A POR2X1_546/A 0.54fF
C52720 POR2X1_61/Y PAND2X1_52/Y 0.03fF
C52721 PAND2X1_839/B POR2X1_20/B 0.01fF
C52722 POR2X1_60/A POR2X1_609/A 0.17fF
C52723 PAND2X1_23/Y D_INPUT_0 0.03fF
C52724 POR2X1_72/B POR2X1_511/Y 0.20fF
C52725 POR2X1_556/A POR2X1_216/a_16_28# 0.02fF
C52726 POR2X1_490/CTRL2 POR2X1_7/A 0.01fF
C52727 POR2X1_556/A POR2X1_366/A 0.02fF
C52728 PAND2X1_73/CTRL PAND2X1_8/Y 0.01fF
C52729 PAND2X1_487/O PAND2X1_69/A 0.16fF
C52730 PAND2X1_65/B POR2X1_461/O 0.03fF
C52731 PAND2X1_706/a_76_28# POR2X1_692/Y 0.01fF
C52732 POR2X1_818/Y POR2X1_790/A 0.03fF
C52733 PAND2X1_423/a_16_344# POR2X1_807/A 0.01fF
C52734 POR2X1_856/B D_GATE_741 0.03fF
C52735 PAND2X1_251/CTRL2 PAND2X1_69/A 0.01fF
C52736 POR2X1_500/A VDD 0.00fF
C52737 POR2X1_205/Y POR2X1_555/B 0.03fF
C52738 PAND2X1_821/CTRL2 POR2X1_590/A -0.00fF
C52739 PAND2X1_93/B POR2X1_631/B 0.03fF
C52740 POR2X1_14/Y POR2X1_7/B 1.73fF
C52741 PAND2X1_55/Y POR2X1_555/B 0.03fF
C52742 PAND2X1_248/CTRL2 POR2X1_532/A 0.01fF
C52743 POR2X1_330/Y PAND2X1_516/CTRL 0.01fF
C52744 POR2X1_297/A POR2X1_297/a_16_28# 0.03fF
C52745 PAND2X1_48/B POR2X1_121/B 0.03fF
C52746 POR2X1_645/O POR2X1_718/A 0.13fF
C52747 PAND2X1_453/A POR2X1_7/B 0.03fF
C52748 PAND2X1_859/A POR2X1_224/CTRL 0.01fF
C52749 PAND2X1_795/O PAND2X1_795/B 0.00fF
C52750 POR2X1_432/CTRL PAND2X1_658/B -0.01fF
C52751 POR2X1_416/B POR2X1_32/CTRL2 0.01fF
C52752 POR2X1_653/m4_208_n4# POR2X1_750/B 0.15fF
C52753 POR2X1_814/A POR2X1_210/A 0.08fF
C52754 POR2X1_13/A PAND2X1_217/B 0.10fF
C52755 POR2X1_83/B POR2X1_697/Y 0.03fF
C52756 POR2X1_595/Y PAND2X1_730/B 0.02fF
C52757 POR2X1_23/Y PAND2X1_341/A 0.03fF
C52758 PAND2X1_96/B POR2X1_499/CTRL 0.01fF
C52759 PAND2X1_562/B VDD 0.02fF
C52760 POR2X1_602/B POR2X1_513/B 0.03fF
C52761 POR2X1_261/Y PAND2X1_569/Y 0.02fF
C52762 POR2X1_102/Y PAND2X1_398/CTRL 0.09fF
C52763 PAND2X1_467/Y POR2X1_257/A 0.07fF
C52764 POR2X1_68/A POR2X1_590/A 0.20fF
C52765 POR2X1_188/A POR2X1_784/A 0.02fF
C52766 POR2X1_284/O POR2X1_330/Y 0.04fF
C52767 PAND2X1_58/CTRL2 VDD -0.00fF
C52768 POR2X1_23/Y POR2X1_91/Y 0.16fF
C52769 PAND2X1_262/CTRL2 POR2X1_786/A 0.05fF
C52770 POR2X1_192/Y POR2X1_439/a_16_28# 0.10fF
C52771 GATE_479 POR2X1_96/A 5.15fF
C52772 PAND2X1_220/Y PAND2X1_182/A 0.05fF
C52773 POR2X1_805/Y POR2X1_712/Y 0.01fF
C52774 PAND2X1_47/B PAND2X1_587/CTRL2 0.01fF
C52775 POR2X1_330/Y PAND2X1_369/O 0.22fF
C52776 POR2X1_368/O PAND2X1_76/Y 0.07fF
C52777 PAND2X1_94/A POR2X1_647/B 0.03fF
C52778 PAND2X1_55/Y POR2X1_330/Y 0.08fF
C52779 POR2X1_78/B POR2X1_547/B 0.03fF
C52780 POR2X1_83/B PAND2X1_357/Y 0.03fF
C52781 POR2X1_105/Y POR2X1_723/a_16_28# 0.03fF
C52782 POR2X1_48/A PAND2X1_388/Y 0.03fF
C52783 PAND2X1_20/A POR2X1_712/Y 0.03fF
C52784 POR2X1_275/A POR2X1_153/Y 0.01fF
C52785 POR2X1_33/CTRL2 POR2X1_68/B 0.01fF
C52786 PAND2X1_474/Y VDD 0.18fF
C52787 POR2X1_614/A PAND2X1_58/A 7.73fF
C52788 POR2X1_734/A PAND2X1_132/O 0.02fF
C52789 POR2X1_218/Y POR2X1_361/CTRL 0.00fF
C52790 POR2X1_686/B VDD 0.19fF
C52791 PAND2X1_738/Y PAND2X1_347/Y 0.05fF
C52792 PAND2X1_477/B POR2X1_14/Y 0.04fF
C52793 POR2X1_96/A POR2X1_485/O 0.00fF
C52794 POR2X1_205/O POR2X1_330/Y 0.01fF
C52795 PAND2X1_658/A PAND2X1_390/Y 0.02fF
C52796 POR2X1_330/Y POR2X1_363/O 0.01fF
C52797 POR2X1_329/CTRL2 PAND2X1_362/B 0.01fF
C52798 POR2X1_48/A PAND2X1_549/B 0.03fF
C52799 PAND2X1_35/Y POR2X1_236/Y 0.05fF
C52800 POR2X1_264/Y PAND2X1_41/B 0.07fF
C52801 POR2X1_13/A VDD 3.41fF
C52802 PAND2X1_81/B POR2X1_500/A 0.00fF
C52803 POR2X1_485/Y PAND2X1_325/O 0.01fF
C52804 POR2X1_33/m4_208_n4# D_INPUT_1 0.08fF
C52805 POR2X1_48/A POR2X1_416/CTRL 0.01fF
C52806 PAND2X1_58/A POR2X1_38/B 0.13fF
C52807 PAND2X1_94/A PAND2X1_27/m4_208_n4# 0.12fF
C52808 POR2X1_60/A PAND2X1_509/CTRL2 0.02fF
C52809 POR2X1_78/A PAND2X1_173/CTRL2 0.01fF
C52810 PAND2X1_20/A POR2X1_500/Y 1.02fF
C52811 PAND2X1_115/O POR2X1_106/Y 0.02fF
C52812 PAND2X1_552/B PAND2X1_714/A 0.01fF
C52813 POR2X1_136/CTRL POR2X1_40/Y 0.03fF
C52814 PAND2X1_216/B POR2X1_490/Y 0.04fF
C52815 PAND2X1_565/O POR2X1_40/Y 0.04fF
C52816 POR2X1_814/B POR2X1_204/CTRL2 0.11fF
C52817 POR2X1_60/A POR2X1_38/Y 0.41fF
C52818 POR2X1_424/a_16_28# POR2X1_511/Y 0.01fF
C52819 PAND2X1_23/Y PAND2X1_90/Y 0.12fF
C52820 PAND2X1_214/B VDD 0.04fF
C52821 POR2X1_355/O D_GATE_741 0.31fF
C52822 POR2X1_333/A POR2X1_775/a_16_28# 0.10fF
C52823 POR2X1_751/A POR2X1_751/a_16_28# 0.09fF
C52824 POR2X1_842/CTRL2 POR2X1_675/Y 0.01fF
C52825 PAND2X1_52/Y POR2X1_35/Y 0.01fF
C52826 POR2X1_814/B POR2X1_712/Y 0.03fF
C52827 PAND2X1_859/A PAND2X1_227/CTRL 0.01fF
C52828 POR2X1_740/O POR2X1_740/Y 0.01fF
C52829 POR2X1_407/Y POR2X1_330/Y 0.05fF
C52830 POR2X1_57/O VDD 0.00fF
C52831 POR2X1_483/A POR2X1_833/O 0.01fF
C52832 PAND2X1_390/Y POR2X1_73/Y 0.03fF
C52833 PAND2X1_642/CTRL POR2X1_48/A 0.01fF
C52834 PAND2X1_643/Y POR2X1_666/Y 0.03fF
C52835 POR2X1_43/B PAND2X1_787/Y 0.03fF
C52836 POR2X1_63/CTRL POR2X1_236/Y 0.14fF
C52837 PAND2X1_476/A POR2X1_20/B 0.03fF
C52838 POR2X1_260/B POR2X1_715/A 0.06fF
C52839 POR2X1_814/A PAND2X1_56/A 0.05fF
C52840 POR2X1_809/Y POR2X1_750/B 0.66fF
C52841 POR2X1_254/Y POR2X1_785/A 0.39fF
C52842 POR2X1_248/CTRL2 POR2X1_5/Y 0.08fF
C52843 PAND2X1_472/B POR2X1_7/B 0.19fF
C52844 POR2X1_621/B PAND2X1_6/A 0.11fF
C52845 PAND2X1_20/A POR2X1_128/B 0.01fF
C52846 POR2X1_376/B PAND2X1_565/A 0.00fF
C52847 PAND2X1_205/m4_208_n4# PAND2X1_728/m4_208_n4# 0.13fF
C52848 PAND2X1_859/A PAND2X1_509/O 0.02fF
C52849 POR2X1_255/CTRL2 PAND2X1_349/A 0.01fF
C52850 POR2X1_463/CTRL PAND2X1_52/B 0.27fF
C52851 POR2X1_814/B POR2X1_500/Y 0.05fF
C52852 POR2X1_105/Y POR2X1_501/B 0.01fF
C52853 POR2X1_567/B POR2X1_566/CTRL2 0.03fF
C52854 POR2X1_639/Y POR2X1_639/A 0.01fF
C52855 PAND2X1_216/B PAND2X1_561/O 0.16fF
C52856 PAND2X1_56/O POR2X1_832/B 0.03fF
C52857 POR2X1_502/A POR2X1_789/Y 0.00fF
C52858 PAND2X1_473/Y POR2X1_599/A 0.05fF
C52859 POR2X1_63/O VDD 0.00fF
C52860 POR2X1_855/B POR2X1_467/Y 0.06fF
C52861 POR2X1_378/Y POR2X1_55/Y 0.78fF
C52862 POR2X1_502/A PAND2X1_95/O 0.05fF
C52863 PAND2X1_671/Y PAND2X1_69/A 0.01fF
C52864 POR2X1_750/A POR2X1_7/A 0.02fF
C52865 POR2X1_403/a_16_28# PAND2X1_69/A 0.01fF
C52866 PAND2X1_651/Y PAND2X1_455/m4_208_n4# 0.09fF
C52867 PAND2X1_651/Y POR2X1_236/Y 0.02fF
C52868 POR2X1_102/Y POR2X1_7/O 0.01fF
C52869 POR2X1_669/B POR2X1_523/O 0.64fF
C52870 PAND2X1_417/CTRL POR2X1_736/A 0.09fF
C52871 POR2X1_55/Y POR2X1_7/B 0.22fF
C52872 POR2X1_740/Y PAND2X1_152/CTRL 0.00fF
C52873 PAND2X1_127/a_76_28# POR2X1_66/A 0.02fF
C52874 POR2X1_493/A PAND2X1_48/A 0.01fF
C52875 POR2X1_862/B POR2X1_537/B 0.00fF
C52876 PAND2X1_787/A PAND2X1_787/a_16_344# 0.01fF
C52877 PAND2X1_64/O PAND2X1_18/B 0.07fF
C52878 PAND2X1_65/B POR2X1_686/CTRL 0.01fF
C52879 POR2X1_23/Y POR2X1_109/Y 0.05fF
C52880 POR2X1_278/Y PAND2X1_566/Y 0.05fF
C52881 POR2X1_36/B POR2X1_376/B 0.00fF
C52882 POR2X1_66/B POR2X1_61/CTRL2 0.00fF
C52883 POR2X1_388/CTRL2 POR2X1_566/A 0.01fF
C52884 PAND2X1_55/CTRL PAND2X1_60/B 0.01fF
C52885 POR2X1_52/A POR2X1_289/CTRL2 0.02fF
C52886 POR2X1_89/Y POR2X1_394/A 0.06fF
C52887 INPUT_1 POR2X1_60/A 0.06fF
C52888 POR2X1_564/Y POR2X1_68/A 0.02fF
C52889 POR2X1_400/A POR2X1_219/B 0.04fF
C52890 POR2X1_504/CTRL2 POR2X1_14/Y 0.00fF
C52891 POR2X1_791/Y PAND2X1_60/B 0.28fF
C52892 POR2X1_614/A POR2X1_435/Y 0.07fF
C52893 PAND2X1_661/B VDD 0.21fF
C52894 POR2X1_271/A POR2X1_32/A 0.04fF
C52895 POR2X1_809/A D_INPUT_0 0.03fF
C52896 INPUT_1 POR2X1_634/A 0.05fF
C52897 POR2X1_637/B PAND2X1_60/B 0.02fF
C52898 PAND2X1_852/CTRL2 POR2X1_42/Y 0.01fF
C52899 PAND2X1_643/Y VDD 0.26fF
C52900 POR2X1_347/B PAND2X1_69/CTRL2 0.13fF
C52901 PAND2X1_495/CTRL VDD -0.00fF
C52902 PAND2X1_220/Y POR2X1_283/A 0.05fF
C52903 POR2X1_614/A PAND2X1_309/CTRL2 0.03fF
C52904 POR2X1_860/A POR2X1_218/CTRL 0.01fF
C52905 PAND2X1_56/Y PAND2X1_48/B 0.05fF
C52906 POR2X1_507/O POR2X1_355/A 0.01fF
C52907 POR2X1_49/Y PAND2X1_467/Y 0.02fF
C52908 PAND2X1_35/Y POR2X1_229/CTRL 0.01fF
C52909 POR2X1_807/A POR2X1_590/O 0.01fF
C52910 POR2X1_65/A PAND2X1_559/O 0.04fF
C52911 PAND2X1_793/Y POR2X1_90/Y 0.11fF
C52912 POR2X1_52/A PAND2X1_565/A 0.03fF
C52913 POR2X1_750/B POR2X1_675/Y 0.03fF
C52914 POR2X1_60/A POR2X1_153/Y 2.40fF
C52915 PAND2X1_535/CTRL POR2X1_236/Y 0.03fF
C52916 D_INPUT_3 PAND2X1_14/a_16_344# 0.02fF
C52917 POR2X1_68/A POR2X1_214/B 0.03fF
C52918 POR2X1_267/m4_208_n4# POR2X1_260/A 0.15fF
C52919 POR2X1_220/Y POR2X1_210/Y 0.61fF
C52920 PAND2X1_863/B POR2X1_761/Y 0.00fF
C52921 POR2X1_250/A PAND2X1_537/CTRL 0.04fF
C52922 POR2X1_296/B POR2X1_294/A 0.03fF
C52923 INPUT_0 POR2X1_239/Y 0.12fF
C52924 POR2X1_72/B PAND2X1_704/CTRL2 0.03fF
C52925 PAND2X1_90/Y POR2X1_520/A 0.00fF
C52926 POR2X1_489/A POR2X1_68/B 0.01fF
C52927 PAND2X1_675/A PAND2X1_798/B 0.07fF
C52928 PAND2X1_803/a_56_28# POR2X1_83/B 0.00fF
C52929 PAND2X1_696/CTRL POR2X1_66/A 0.01fF
C52930 POR2X1_271/A POR2X1_417/Y 0.04fF
C52931 PAND2X1_96/B POR2X1_193/A 0.03fF
C52932 POR2X1_661/A POR2X1_814/A 0.10fF
C52933 PAND2X1_96/B POR2X1_579/Y 0.04fF
C52934 PAND2X1_798/B PAND2X1_469/B 0.01fF
C52935 POR2X1_335/A POR2X1_407/A 0.03fF
C52936 POR2X1_750/B POR2X1_544/B 0.03fF
C52937 POR2X1_559/B VDD 0.02fF
C52938 POR2X1_259/B PAND2X1_7/Y 0.03fF
C52939 POR2X1_696/a_16_28# POR2X1_394/A 0.03fF
C52940 POR2X1_383/A POR2X1_483/B 0.08fF
C52941 POR2X1_72/B POR2X1_129/Y 0.14fF
C52942 PAND2X1_614/CTRL POR2X1_129/Y 0.01fF
C52943 POR2X1_96/A PAND2X1_785/a_76_28# 0.01fF
C52944 POR2X1_52/A POR2X1_36/B 0.09fF
C52945 VDD PAND2X1_510/B 0.58fF
C52946 POR2X1_96/A PAND2X1_175/B 0.02fF
C52947 PAND2X1_726/B POR2X1_763/CTRL2 0.03fF
C52948 VDD POR2X1_321/Y 0.10fF
C52949 POR2X1_128/O POR2X1_510/Y 0.04fF
C52950 PAND2X1_212/B PAND2X1_352/Y 0.17fF
C52951 POR2X1_302/A POR2X1_840/B 0.50fF
C52952 PAND2X1_728/O VDD 0.00fF
C52953 POR2X1_109/O POR2X1_77/Y 0.02fF
C52954 POR2X1_226/Y POR2X1_394/A 0.06fF
C52955 PAND2X1_453/O PAND2X1_241/Y 0.03fF
C52956 PAND2X1_40/CTRL2 POR2X1_407/Y 0.01fF
C52957 INPUT_1 POR2X1_381/a_16_28# 0.03fF
C52958 PAND2X1_569/CTRL2 VDD 0.00fF
C52959 POR2X1_770/A POR2X1_260/A 0.01fF
C52960 PAND2X1_219/A PAND2X1_737/O 0.01fF
C52961 POR2X1_417/Y PAND2X1_352/CTRL2 0.01fF
C52962 PAND2X1_651/Y POR2X1_229/CTRL 0.27fF
C52963 POR2X1_68/B POR2X1_391/Y 0.07fF
C52964 POR2X1_383/A PAND2X1_38/m4_208_n4# 0.07fF
C52965 POR2X1_446/a_56_344# PAND2X1_72/A 0.00fF
C52966 PAND2X1_659/Y POR2X1_72/B 0.92fF
C52967 POR2X1_862/B PAND2X1_48/A 0.03fF
C52968 D_INPUT_0 POR2X1_711/Y 0.07fF
C52969 POR2X1_119/Y POR2X1_609/O 0.03fF
C52970 POR2X1_614/A PAND2X1_96/B 0.22fF
C52971 PAND2X1_48/B POR2X1_383/A 0.76fF
C52972 POR2X1_660/A POR2X1_737/A 0.03fF
C52973 PAND2X1_536/CTRL PAND2X1_60/B 0.01fF
C52974 POR2X1_90/Y PAND2X1_711/A 0.06fF
C52975 POR2X1_99/B POR2X1_244/O 0.00fF
C52976 PAND2X1_292/CTRL2 POR2X1_66/A 0.01fF
C52977 POR2X1_516/a_16_28# PAND2X1_651/Y 0.10fF
C52978 PAND2X1_552/B PAND2X1_854/A 0.02fF
C52979 POR2X1_317/O POR2X1_854/B 0.04fF
C52980 POR2X1_3/A PAND2X1_635/CTRL 0.01fF
C52981 PAND2X1_316/O POR2X1_318/A 0.00fF
C52982 POR2X1_809/A PAND2X1_90/Y 0.02fF
C52983 POR2X1_134/Y POR2X1_132/Y 0.06fF
C52984 POR2X1_834/Y POR2X1_307/Y 0.17fF
C52985 POR2X1_549/A PAND2X1_63/B 0.01fF
C52986 POR2X1_57/A PAND2X1_182/O 0.01fF
C52987 POR2X1_355/B POR2X1_353/A 0.03fF
C52988 POR2X1_186/Y POR2X1_552/A 0.03fF
C52989 PAND2X1_254/m4_208_n4# POR2X1_7/A 0.08fF
C52990 POR2X1_730/Y POR2X1_802/B 0.07fF
C52991 POR2X1_376/B POR2X1_701/O 0.05fF
C52992 PAND2X1_800/CTRL PAND2X1_863/B 0.01fF
C52993 POR2X1_254/Y POR2X1_186/B 0.03fF
C52994 POR2X1_51/CTRL2 INPUT_7 0.00fF
C52995 PAND2X1_137/Y POR2X1_103/O 0.01fF
C52996 POR2X1_68/A POR2X1_623/A 0.01fF
C52997 POR2X1_49/O POR2X1_409/B 0.03fF
C52998 POR2X1_504/CTRL2 POR2X1_55/Y 0.01fF
C52999 POR2X1_740/Y POR2X1_260/A 0.07fF
C53000 POR2X1_40/Y PAND2X1_169/O 0.03fF
C53001 POR2X1_791/B PAND2X1_60/B 0.01fF
C53002 POR2X1_42/Y PAND2X1_507/CTRL2 0.04fF
C53003 POR2X1_16/A PAND2X1_652/A 0.27fF
C53004 POR2X1_407/A POR2X1_249/Y 0.03fF
C53005 POR2X1_354/a_16_28# POR2X1_854/B 0.03fF
C53006 POR2X1_858/A POR2X1_660/A 0.02fF
C53007 POR2X1_51/A POR2X1_328/CTRL2 0.01fF
C53008 POR2X1_96/A PAND2X1_858/O 0.04fF
C53009 POR2X1_411/B POR2X1_67/Y 0.03fF
C53010 POR2X1_468/Y POR2X1_319/Y 0.02fF
C53011 POR2X1_388/CTRL POR2X1_703/A 0.03fF
C53012 POR2X1_416/B PAND2X1_354/A 0.03fF
C53013 POR2X1_41/B POR2X1_265/Y 0.02fF
C53014 POR2X1_119/Y PAND2X1_735/Y 0.10fF
C53015 POR2X1_540/O POR2X1_181/B 0.17fF
C53016 POR2X1_73/Y PAND2X1_123/O 0.02fF
C53017 POR2X1_584/a_56_344# POR2X1_260/A 0.00fF
C53018 POR2X1_804/A POR2X1_456/B 0.05fF
C53019 PAND2X1_65/B PAND2X1_134/a_76_28# 0.02fF
C53020 POR2X1_669/B POR2X1_321/CTRL2 0.05fF
C53021 PAND2X1_596/O POR2X1_761/A 0.02fF
C53022 PAND2X1_844/O POR2X1_43/B 0.04fF
C53023 PAND2X1_793/Y PAND2X1_185/CTRL2 0.01fF
C53024 POR2X1_271/A POR2X1_184/Y 0.03fF
C53025 POR2X1_130/A PAND2X1_136/CTRL 0.03fF
C53026 POR2X1_730/Y POR2X1_532/A 0.03fF
C53027 PAND2X1_865/Y POR2X1_46/Y 0.03fF
C53028 POR2X1_276/A POR2X1_366/A 0.25fF
C53029 POR2X1_394/A POR2X1_56/Y 0.07fF
C53030 POR2X1_556/A POR2X1_658/CTRL 0.03fF
C53031 POR2X1_532/A PAND2X1_690/CTRL 0.01fF
C53032 PAND2X1_580/B POR2X1_767/Y 0.02fF
C53033 POR2X1_283/A POR2X1_751/a_16_28# 0.01fF
C53034 PAND2X1_90/Y POR2X1_711/Y 0.10fF
C53035 POR2X1_416/B POR2X1_290/a_56_344# 0.00fF
C53036 POR2X1_485/Y POR2X1_484/Y 0.01fF
C53037 POR2X1_85/Y POR2X1_230/CTRL 0.08fF
C53038 POR2X1_75/CTRL POR2X1_271/A 0.03fF
C53039 PAND2X1_69/A POR2X1_507/A 0.07fF
C53040 PAND2X1_55/Y POR2X1_337/Y 0.07fF
C53041 POR2X1_680/CTRL POR2X1_79/Y 0.01fF
C53042 PAND2X1_742/B POR2X1_385/Y 0.05fF
C53043 INPUT_6 POR2X1_260/A 0.01fF
C53044 POR2X1_610/O POR2X1_814/A 0.00fF
C53045 POR2X1_416/B POR2X1_48/CTRL 0.01fF
C53046 POR2X1_326/CTRL POR2X1_319/Y 0.00fF
C53047 PAND2X1_823/CTRL POR2X1_854/B 0.15fF
C53048 POR2X1_52/CTRL2 PAND2X1_215/B 0.03fF
C53049 POR2X1_599/A POR2X1_7/Y 0.05fF
C53050 POR2X1_564/Y POR2X1_169/A 0.03fF
C53051 POR2X1_267/Y POR2X1_294/A 0.09fF
C53052 POR2X1_341/Y POR2X1_186/B 0.03fF
C53053 PAND2X1_725/A PAND2X1_725/a_76_28# 0.02fF
C53054 POR2X1_16/A POR2X1_437/CTRL2 0.01fF
C53055 D_GATE_741 POR2X1_191/Y 0.10fF
C53056 POR2X1_809/A PAND2X1_583/a_16_344# 0.01fF
C53057 POR2X1_505/CTRL2 PAND2X1_632/B 0.01fF
C53058 POR2X1_615/Y POR2X1_39/B 0.01fF
C53059 POR2X1_760/A POR2X1_674/O 0.06fF
C53060 POR2X1_370/Y POR2X1_717/B 0.02fF
C53061 POR2X1_416/B INPUT_5 0.06fF
C53062 POR2X1_41/B PAND2X1_327/CTRL 0.00fF
C53063 POR2X1_192/Y PAND2X1_52/B 0.10fF
C53064 POR2X1_503/CTRL2 POR2X1_8/Y 0.03fF
C53065 POR2X1_43/B PAND2X1_860/a_16_344# 0.01fF
C53066 PAND2X1_5/CTRL POR2X1_4/Y 0.01fF
C53067 PAND2X1_841/O POR2X1_39/B 0.01fF
C53068 POR2X1_456/B PAND2X1_313/O 0.04fF
C53069 POR2X1_316/Y PAND2X1_6/A 0.07fF
C53070 PAND2X1_309/CTRL POR2X1_717/B 0.01fF
C53071 POR2X1_305/a_56_344# POR2X1_42/Y 0.00fF
C53072 POR2X1_14/Y PAND2X1_206/B 0.07fF
C53073 PAND2X1_498/O PAND2X1_72/A 0.01fF
C53074 POR2X1_837/A POR2X1_202/a_16_28# 0.10fF
C53075 POR2X1_716/CTRL POR2X1_723/B 0.01fF
C53076 PAND2X1_497/O POR2X1_624/Y 0.02fF
C53077 POR2X1_416/B POR2X1_426/O 0.18fF
C53078 POR2X1_158/Y POR2X1_426/CTRL 0.00fF
C53079 POR2X1_158/O POR2X1_425/Y 0.01fF
C53080 POR2X1_774/A POR2X1_260/A 0.03fF
C53081 POR2X1_68/B POR2X1_383/Y 0.04fF
C53082 POR2X1_276/Y PAND2X1_48/A 0.08fF
C53083 PAND2X1_139/CTRL2 PAND2X1_349/A 0.01fF
C53084 POR2X1_116/A POR2X1_296/B 0.05fF
C53085 PAND2X1_23/Y POR2X1_715/O 0.01fF
C53086 POR2X1_311/Y POR2X1_329/Y 0.03fF
C53087 POR2X1_356/A POR2X1_863/A 0.29fF
C53088 POR2X1_502/Y POR2X1_502/CTRL 0.00fF
C53089 PAND2X1_674/O PAND2X1_72/A 0.03fF
C53090 POR2X1_38/Y PAND2X1_339/CTRL2 0.06fF
C53091 POR2X1_461/O POR2X1_814/A 0.00fF
C53092 POR2X1_68/A POR2X1_87/a_16_28# 0.03fF
C53093 POR2X1_46/Y POR2X1_91/O 0.01fF
C53094 POR2X1_96/a_16_28# POR2X1_153/Y 0.02fF
C53095 POR2X1_67/Y POR2X1_849/CTRL 0.03fF
C53096 PAND2X1_29/O PAND2X1_52/B 0.12fF
C53097 PAND2X1_813/a_16_344# POR2X1_62/Y 0.01fF
C53098 PAND2X1_681/CTRL PAND2X1_32/B 0.01fF
C53099 POR2X1_532/A POR2X1_555/O 0.02fF
C53100 PAND2X1_39/B POR2X1_805/Y 0.01fF
C53101 POR2X1_341/A POR2X1_267/A 0.09fF
C53102 POR2X1_178/a_16_28# POR2X1_416/B 0.03fF
C53103 PAND2X1_641/Y POR2X1_83/Y 0.01fF
C53104 POR2X1_567/B PAND2X1_237/O 0.48fF
C53105 POR2X1_416/B POR2X1_258/a_16_28# 0.03fF
C53106 POR2X1_159/CTRL2 INPUT_3 0.15fF
C53107 PAND2X1_20/A PAND2X1_39/B 0.17fF
C53108 PAND2X1_826/O POR2X1_838/B 0.01fF
C53109 PAND2X1_841/CTRL2 POR2X1_677/Y 0.00fF
C53110 PAND2X1_60/B POR2X1_500/CTRL2 0.03fF
C53111 D_INPUT_7 INPUT_4 0.03fF
C53112 POR2X1_54/Y PAND2X1_817/O 0.21fF
C53113 POR2X1_68/B POR2X1_8/O 0.03fF
C53114 PAND2X1_71/Y PAND2X1_527/a_16_344# 0.01fF
C53115 PAND2X1_6/Y POR2X1_76/B 0.03fF
C53116 POR2X1_519/O POR2X1_39/B 0.16fF
C53117 POR2X1_88/O POR2X1_14/Y 0.00fF
C53118 POR2X1_862/A POR2X1_285/Y -0.00fF
C53119 POR2X1_505/Y POR2X1_628/Y 0.02fF
C53120 POR2X1_656/O D_INPUT_0 0.01fF
C53121 POR2X1_624/Y PAND2X1_41/B 0.03fF
C53122 POR2X1_281/CTRL POR2X1_416/B 0.01fF
C53123 POR2X1_659/A POR2X1_750/B 0.26fF
C53124 POR2X1_814/B PAND2X1_39/B 0.12fF
C53125 POR2X1_52/A POR2X1_67/Y 0.06fF
C53126 POR2X1_838/B POR2X1_294/Y 0.21fF
C53127 POR2X1_796/A PAND2X1_72/A 0.03fF
C53128 PAND2X1_206/B PAND2X1_341/CTRL2 0.00fF
C53129 PAND2X1_48/B POR2X1_648/Y 0.03fF
C53130 PAND2X1_206/B POR2X1_55/Y 0.10fF
C53131 PAND2X1_432/a_16_344# POR2X1_866/A 0.04fF
C53132 POR2X1_669/B PAND2X1_721/B 0.02fF
C53133 PAND2X1_72/A POR2X1_332/CTRL2 0.00fF
C53134 POR2X1_634/A POR2X1_637/O 0.04fF
C53135 POR2X1_542/Y POR2X1_552/A 0.01fF
C53136 POR2X1_863/A POR2X1_569/A 0.07fF
C53137 POR2X1_41/B POR2X1_263/O 0.00fF
C53138 PAND2X1_73/Y POR2X1_285/Y 0.03fF
C53139 PAND2X1_58/A POR2X1_590/A 0.15fF
C53140 PAND2X1_562/Y VDD 0.00fF
C53141 POR2X1_567/B POR2X1_186/Y 0.10fF
C53142 POR2X1_60/A PAND2X1_794/CTRL2 0.01fF
C53143 POR2X1_499/A PAND2X1_372/O 0.01fF
C53144 POR2X1_150/Y PAND2X1_335/CTRL2 0.15fF
C53145 POR2X1_13/A PAND2X1_9/Y 0.04fF
C53146 POR2X1_119/Y POR2X1_316/Y 0.05fF
C53147 POR2X1_23/Y POR2X1_278/CTRL2 0.01fF
C53148 POR2X1_37/Y POR2X1_72/B 0.65fF
C53149 PAND2X1_93/B POR2X1_61/Y 0.05fF
C53150 PAND2X1_402/CTRL D_INPUT_0 0.02fF
C53151 PAND2X1_20/A POR2X1_805/Y 0.01fF
C53152 POR2X1_87/B POR2X1_260/A 0.04fF
C53153 POR2X1_83/B POR2X1_667/A 1.09fF
C53154 POR2X1_612/Y POR2X1_5/Y 0.02fF
C53155 PAND2X1_613/CTRL2 PAND2X1_8/Y 0.04fF
C53156 POR2X1_260/B PAND2X1_380/CTRL 0.01fF
C53157 POR2X1_445/O POR2X1_341/A 0.06fF
C53158 POR2X1_257/A PAND2X1_254/Y 0.01fF
C53159 POR2X1_696/a_16_28# POR2X1_669/B 0.09fF
C53160 POR2X1_94/A POR2X1_296/B 0.05fF
C53161 POR2X1_445/A POR2X1_445/CTRL2 0.01fF
C53162 POR2X1_20/B PAND2X1_776/O 0.01fF
C53163 POR2X1_175/A POR2X1_174/A 0.47fF
C53164 PAND2X1_608/O POR2X1_73/Y 0.04fF
C53165 POR2X1_366/Y POR2X1_663/B 0.03fF
C53166 POR2X1_60/A PAND2X1_214/A 0.01fF
C53167 PAND2X1_404/Y PAND2X1_862/B 0.03fF
C53168 POR2X1_332/B POR2X1_260/B 0.22fF
C53169 PAND2X1_218/B INPUT_0 0.01fF
C53170 POR2X1_14/Y POR2X1_750/B 0.04fF
C53171 PAND2X1_392/B POR2X1_29/A 0.03fF
C53172 POR2X1_466/a_16_28# POR2X1_209/A 0.03fF
C53173 POR2X1_678/Y VDD 0.20fF
C53174 POR2X1_814/B POR2X1_805/Y 0.01fF
C53175 D_INPUT_0 PAND2X1_206/CTRL 0.06fF
C53176 POR2X1_490/Y PAND2X1_216/CTRL2 0.03fF
C53177 POR2X1_78/A POR2X1_61/Y 0.03fF
C53178 PAND2X1_846/a_76_28# POR2X1_815/Y 0.05fF
C53179 POR2X1_655/A PAND2X1_385/CTRL2 0.00fF
C53180 POR2X1_78/O POR2X1_78/Y 0.00fF
C53181 GATE_479 PAND2X1_467/B 0.03fF
C53182 POR2X1_856/B PAND2X1_627/a_76_28# 0.02fF
C53183 PAND2X1_20/A POR2X1_814/B 0.26fF
C53184 PAND2X1_811/A VDD 0.00fF
C53185 POR2X1_36/B POR2X1_18/a_16_28# 0.03fF
C53186 POR2X1_462/B POR2X1_859/O 0.01fF
C53187 POR2X1_42/CTRL POR2X1_20/B 0.01fF
C53188 POR2X1_624/Y POR2X1_130/Y 0.51fF
C53189 POR2X1_189/Y POR2X1_679/Y 0.16fF
C53190 POR2X1_102/Y POR2X1_760/CTRL2 0.03fF
C53191 PAND2X1_661/Y POR2X1_681/CTRL2 0.03fF
C53192 PAND2X1_93/B POR2X1_652/Y 0.09fF
C53193 POR2X1_96/A POR2X1_409/B 0.09fF
C53194 POR2X1_29/A VDD 2.49fF
C53195 POR2X1_54/Y PAND2X1_6/A 1.34fF
C53196 PAND2X1_667/O POR2X1_590/A 0.01fF
C53197 POR2X1_163/Y VDD 0.01fF
C53198 POR2X1_614/A POR2X1_676/CTRL2 0.00fF
C53199 PAND2X1_661/B PAND2X1_9/Y 0.01fF
C53200 POR2X1_834/Y POR2X1_648/A 0.00fF
C53201 PAND2X1_139/a_16_344# POR2X1_40/Y 0.01fF
C53202 PAND2X1_477/CTRL POR2X1_238/Y 0.01fF
C53203 PAND2X1_20/A POR2X1_325/A 0.03fF
C53204 PAND2X1_691/Y PAND2X1_644/CTRL 0.09fF
C53205 PAND2X1_23/Y PAND2X1_59/B 2.57fF
C53206 POR2X1_490/Y PAND2X1_218/O 0.01fF
C53207 POR2X1_590/A POR2X1_435/Y 0.01fF
C53208 POR2X1_473/CTRL2 PAND2X1_32/B 0.02fF
C53209 POR2X1_257/A PAND2X1_161/Y 0.92fF
C53210 POR2X1_230/Y POR2X1_32/A 0.29fF
C53211 PAND2X1_276/CTRL2 PAND2X1_390/Y 0.01fF
C53212 POR2X1_645/CTRL2 POR2X1_330/Y 0.15fF
C53213 PAND2X1_540/CTRL POR2X1_106/Y 0.01fF
C53214 POR2X1_365/Y POR2X1_220/B 0.02fF
C53215 POR2X1_566/A POR2X1_454/B 0.05fF
C53216 POR2X1_294/Y POR2X1_294/B 0.01fF
C53217 PAND2X1_216/B POR2X1_329/A 1.41fF
C53218 POR2X1_122/Y POR2X1_40/Y 0.03fF
C53219 POR2X1_593/B POR2X1_830/A 0.02fF
C53220 POR2X1_66/B PAND2X1_131/CTRL 0.01fF
C53221 POR2X1_647/B POR2X1_865/O 0.01fF
C53222 D_INPUT_0 POR2X1_733/A 0.07fF
C53223 PAND2X1_93/B POR2X1_35/Y 0.07fF
C53224 PAND2X1_6/Y POR2X1_301/A 0.01fF
C53225 POR2X1_568/B POR2X1_568/A 0.00fF
C53226 PAND2X1_65/B POR2X1_392/B 0.04fF
C53227 PAND2X1_773/B PAND2X1_354/A 0.13fF
C53228 POR2X1_123/A POR2X1_137/B 0.03fF
C53229 POR2X1_32/Y PAND2X1_35/A 0.03fF
C53230 POR2X1_334/B D_INPUT_0 0.03fF
C53231 POR2X1_76/A PAND2X1_311/CTRL 0.00fF
C53232 POR2X1_65/A POR2X1_5/Y 0.03fF
C53233 POR2X1_287/A POR2X1_249/Y 0.09fF
C53234 POR2X1_602/B VDD 0.30fF
C53235 POR2X1_541/B POR2X1_274/B 0.00fF
C53236 POR2X1_78/B POR2X1_186/Y 0.07fF
C53237 POR2X1_822/a_76_344# POR2X1_40/Y 0.01fF
C53238 POR2X1_558/a_76_344# POR2X1_558/B 0.01fF
C53239 POR2X1_406/Y POR2X1_72/B 0.03fF
C53240 POR2X1_68/A POR2X1_66/A 0.28fF
C53241 POR2X1_72/Y PAND2X1_657/O 0.02fF
C53242 POR2X1_71/Y PAND2X1_657/a_16_344# 0.02fF
C53243 POR2X1_287/CTRL2 POR2X1_733/A 0.15fF
C53244 POR2X1_850/A POR2X1_362/B 0.95fF
C53245 POR2X1_624/Y POR2X1_228/Y 0.10fF
C53246 PAND2X1_61/Y POR2X1_497/Y 0.62fF
C53247 POR2X1_269/CTRL POR2X1_741/Y 0.00fF
C53248 PAND2X1_478/B POR2X1_46/Y 1.49fF
C53249 POR2X1_814/B POR2X1_325/A 0.03fF
C53250 POR2X1_49/Y PAND2X1_556/B 0.07fF
C53251 POR2X1_97/A POR2X1_350/O 0.01fF
C53252 PAND2X1_220/Y POR2X1_488/a_16_28# 0.06fF
C53253 PAND2X1_785/Y PAND2X1_390/Y 0.03fF
C53254 POR2X1_329/O PAND2X1_557/A 0.01fF
C53255 POR2X1_462/CTRL POR2X1_559/A 0.01fF
C53256 POR2X1_718/CTRL VDD 0.00fF
C53257 POR2X1_65/A PAND2X1_549/CTRL2 0.03fF
C53258 PAND2X1_230/CTRL POR2X1_785/A 0.01fF
C53259 PAND2X1_31/CTRL2 INPUT_6 0.00fF
C53260 POR2X1_547/CTRL POR2X1_78/A 0.01fF
C53261 PAND2X1_97/Y POR2X1_394/A 0.04fF
C53262 PAND2X1_208/CTRL PAND2X1_35/Y 0.01fF
C53263 POR2X1_568/A POR2X1_161/CTRL2 0.03fF
C53264 PAND2X1_660/B VDD 0.01fF
C53265 POR2X1_381/O POR2X1_236/Y 0.08fF
C53266 PAND2X1_786/O POR2X1_293/Y 0.05fF
C53267 POR2X1_303/a_16_28# POR2X1_302/Y 0.02fF
C53268 POR2X1_23/Y POR2X1_425/Y 0.00fF
C53269 POR2X1_484/Y PAND2X1_726/B 0.12fF
C53270 POR2X1_213/B VDD 0.07fF
C53271 POR2X1_541/B PAND2X1_72/Y 0.03fF
C53272 PAND2X1_733/CTRL2 POR2X1_7/B 0.01fF
C53273 POR2X1_274/CTRL2 POR2X1_573/A 0.01fF
C53274 PAND2X1_658/B PAND2X1_573/B 0.00fF
C53275 POR2X1_72/B POR2X1_293/Y 0.30fF
C53276 POR2X1_814/B PAND2X1_176/CTRL2 0.03fF
C53277 POR2X1_31/O POR2X1_12/A 0.01fF
C53278 PAND2X1_204/CTRL2 PAND2X1_735/Y 0.03fF
C53279 POR2X1_730/Y POR2X1_452/Y 0.60fF
C53280 POR2X1_23/Y PAND2X1_338/B 0.03fF
C53281 POR2X1_821/CTRL2 POR2X1_236/Y 0.11fF
C53282 PAND2X1_73/a_16_344# POR2X1_294/B 0.03fF
C53283 POR2X1_750/B POR2X1_55/Y 0.06fF
C53284 POR2X1_274/A POR2X1_569/A 0.18fF
C53285 POR2X1_29/A PAND2X1_32/B 0.03fF
C53286 PAND2X1_6/Y PAND2X1_626/CTRL2 0.11fF
C53287 PAND2X1_449/Y POR2X1_60/A 0.06fF
C53288 PAND2X1_20/A PAND2X1_519/a_16_344# 0.01fF
C53289 POR2X1_255/CTRL2 POR2X1_184/Y 0.00fF
C53290 POR2X1_614/A POR2X1_806/CTRL2 0.01fF
C53291 PAND2X1_41/B POR2X1_785/A 0.06fF
C53292 POR2X1_863/A PAND2X1_72/A 0.13fF
C53293 PAND2X1_96/B POR2X1_590/A 0.68fF
C53294 POR2X1_642/CTRL POR2X1_734/A 0.04fF
C53295 PAND2X1_115/CTRL PAND2X1_562/B 0.06fF
C53296 POR2X1_122/CTRL POR2X1_411/B 0.01fF
C53297 POR2X1_72/B POR2X1_531/a_16_28# 0.02fF
C53298 PAND2X1_58/A PAND2X1_752/Y 0.02fF
C53299 POR2X1_267/A PAND2X1_767/O 0.17fF
C53300 POR2X1_68/A PAND2X1_279/a_16_344# -0.01fF
C53301 PAND2X1_220/Y POR2X1_55/Y 0.03fF
C53302 POR2X1_96/A POR2X1_272/Y 0.03fF
C53303 POR2X1_546/A VDD 0.26fF
C53304 PAND2X1_55/Y POR2X1_543/A 0.40fF
C53305 POR2X1_333/A PAND2X1_69/A 0.03fF
C53306 POR2X1_682/Y INPUT_0 0.05fF
C53307 POR2X1_52/A PAND2X1_736/O 0.16fF
C53308 POR2X1_502/A POR2X1_284/B 0.01fF
C53309 POR2X1_49/Y POR2X1_599/A 0.08fF
C53310 POR2X1_511/Y POR2X1_7/B 0.03fF
C53311 POR2X1_41/B PAND2X1_842/a_76_28# 0.01fF
C53312 POR2X1_74/CTRL2 POR2X1_23/Y 0.03fF
C53313 POR2X1_130/A PAND2X1_56/O 0.04fF
C53314 PAND2X1_863/B PAND2X1_730/B 0.01fF
C53315 PAND2X1_843/O PAND2X1_675/A 0.01fF
C53316 POR2X1_569/O POR2X1_853/A 0.01fF
C53317 POR2X1_8/Y POR2X1_126/O 0.01fF
C53318 POR2X1_66/B POR2X1_194/CTRL2 0.02fF
C53319 POR2X1_23/Y PAND2X1_574/O 0.04fF
C53320 POR2X1_66/B POR2X1_649/CTRL 0.01fF
C53321 POR2X1_278/Y PAND2X1_480/B 0.07fF
C53322 POR2X1_558/A POR2X1_590/A 0.01fF
C53323 POR2X1_60/A POR2X1_591/Y 0.03fF
C53324 POR2X1_16/A PAND2X1_205/A 0.05fF
C53325 PAND2X1_793/Y INPUT_0 0.08fF
C53326 POR2X1_48/A PAND2X1_264/O 0.02fF
C53327 POR2X1_180/B POR2X1_66/A 0.04fF
C53328 PAND2X1_675/O POR2X1_250/Y 0.11fF
C53329 POR2X1_325/CTRL2 POR2X1_78/A 0.00fF
C53330 PAND2X1_92/a_16_344# INPUT_0 0.02fF
C53331 POR2X1_14/Y POR2X1_750/O 0.01fF
C53332 POR2X1_40/Y POR2X1_310/a_56_344# 0.00fF
C53333 POR2X1_102/Y POR2X1_239/Y 0.38fF
C53334 PAND2X1_776/Y PAND2X1_308/Y 0.03fF
C53335 POR2X1_591/A POR2X1_591/Y 0.05fF
C53336 POR2X1_466/A PAND2X1_313/CTRL 0.01fF
C53337 POR2X1_41/B PAND2X1_137/Y 0.07fF
C53338 PAND2X1_69/A POR2X1_734/A 0.12fF
C53339 POR2X1_123/A POR2X1_78/A 1.71fF
C53340 POR2X1_83/Y POR2X1_63/Y 0.02fF
C53341 POR2X1_594/Y VDD -0.00fF
C53342 POR2X1_83/B POR2X1_245/Y 0.01fF
C53343 PAND2X1_48/B INPUT_0 0.09fF
C53344 PAND2X1_568/O POR2X1_7/B 0.03fF
C53345 POR2X1_730/Y POR2X1_220/B 0.03fF
C53346 POR2X1_848/A POR2X1_753/O 0.02fF
C53347 POR2X1_257/A POR2X1_320/O 0.16fF
C53348 POR2X1_51/A POR2X1_408/CTRL 0.01fF
C53349 PAND2X1_828/a_16_344# POR2X1_599/A 0.06fF
C53350 POR2X1_121/A POR2X1_78/B 0.02fF
C53351 POR2X1_154/CTRL2 POR2X1_803/A 0.01fF
C53352 POR2X1_332/B PAND2X1_55/Y 0.19fF
C53353 PAND2X1_249/a_56_28# POR2X1_591/Y 0.00fF
C53354 POR2X1_578/Y POR2X1_776/B 0.03fF
C53355 POR2X1_805/A VDD 0.15fF
C53356 PAND2X1_129/a_16_344# POR2X1_559/Y 0.05fF
C53357 POR2X1_532/A POR2X1_710/A 0.01fF
C53358 PAND2X1_15/CTRL POR2X1_260/A 0.03fF
C53359 POR2X1_673/Y POR2X1_29/A 0.07fF
C53360 PAND2X1_479/A POR2X1_45/Y 0.01fF
C53361 PAND2X1_685/a_16_344# INPUT_0 0.01fF
C53362 PAND2X1_844/CTRL D_INPUT_0 0.10fF
C53363 PAND2X1_280/O PAND2X1_55/Y 0.04fF
C53364 VDD POR2X1_712/Y 0.21fF
C53365 POR2X1_72/B POR2X1_408/Y 0.05fF
C53366 PAND2X1_483/CTRL2 POR2X1_60/A 0.01fF
C53367 POR2X1_65/A POR2X1_165/CTRL 0.01fF
C53368 POR2X1_68/A PAND2X1_293/O 0.02fF
C53369 POR2X1_166/O PAND2X1_714/A 0.15fF
C53370 PAND2X1_659/Y PAND2X1_205/O 0.10fF
C53371 PAND2X1_813/O POR2X1_78/A 0.01fF
C53372 POR2X1_272/a_56_344# PAND2X1_349/A 0.00fF
C53373 POR2X1_333/A POR2X1_326/CTRL 0.08fF
C53374 POR2X1_68/A PAND2X1_524/CTRL 0.01fF
C53375 POR2X1_72/B PAND2X1_374/CTRL 0.01fF
C53376 POR2X1_43/B PAND2X1_636/a_76_28# 0.02fF
C53377 PAND2X1_520/a_16_344# POR2X1_518/Y 0.01fF
C53378 POR2X1_807/O PAND2X1_48/A 0.01fF
C53379 POR2X1_16/A PAND2X1_195/CTRL 0.01fF
C53380 PAND2X1_540/CTRL PAND2X1_114/B 0.04fF
C53381 POR2X1_65/A POR2X1_166/a_16_28# 0.00fF
C53382 POR2X1_508/O POR2X1_579/Y 0.11fF
C53383 POR2X1_725/a_56_344# POR2X1_712/Y 0.00fF
C53384 POR2X1_416/Y POR2X1_411/O 0.01fF
C53385 PAND2X1_57/B POR2X1_804/A 0.08fF
C53386 PAND2X1_594/O POR2X1_151/Y 0.14fF
C53387 POR2X1_79/Y POR2X1_816/A 0.03fF
C53388 POR2X1_133/CTRL2 POR2X1_93/A 0.01fF
C53389 POR2X1_546/A PAND2X1_32/B 0.04fF
C53390 POR2X1_68/A POR2X1_802/B 0.07fF
C53391 POR2X1_794/B POR2X1_456/B 0.03fF
C53392 POR2X1_537/Y POR2X1_858/CTRL 0.01fF
C53393 PAND2X1_734/B POR2X1_229/O 0.01fF
C53394 PAND2X1_57/B PAND2X1_69/O 0.02fF
C53395 POR2X1_584/CTRL2 POR2X1_42/Y 0.05fF
C53396 PAND2X1_490/O PAND2X1_57/B 0.01fF
C53397 PAND2X1_593/m4_208_n4# PAND2X1_219/m4_208_n4# 0.13fF
C53398 PAND2X1_803/CTRL2 POR2X1_60/A 0.13fF
C53399 POR2X1_100/CTRL POR2X1_243/Y 0.04fF
C53400 POR2X1_41/B POR2X1_248/CTRL 0.03fF
C53401 PAND2X1_80/CTRL PAND2X1_111/B 0.01fF
C53402 PAND2X1_23/Y D_GATE_222 0.03fF
C53403 PAND2X1_57/B POR2X1_705/a_16_28# 0.01fF
C53404 PAND2X1_675/A PAND2X1_552/B 0.03fF
C53405 PAND2X1_230/CTRL POR2X1_186/B 0.00fF
C53406 PAND2X1_90/A POR2X1_391/Y 0.06fF
C53407 POR2X1_780/O POR2X1_260/A 0.02fF
C53408 PAND2X1_254/CTRL POR2X1_253/Y 0.03fF
C53409 POR2X1_178/a_16_28# PAND2X1_738/Y 0.08fF
C53410 POR2X1_198/CTRL POR2X1_68/A 0.00fF
C53411 PAND2X1_719/Y POR2X1_394/A 0.22fF
C53412 PAND2X1_575/B POR2X1_394/A 0.22fF
C53413 PAND2X1_6/Y POR2X1_84/CTRL 0.01fF
C53414 POR2X1_272/Y POR2X1_7/A 0.03fF
C53415 PAND2X1_835/Y POR2X1_293/Y 0.00fF
C53416 PAND2X1_220/CTRL PAND2X1_566/Y 0.01fF
C53417 POR2X1_164/Y POR2X1_376/B 0.01fF
C53418 POR2X1_740/Y PAND2X1_111/a_16_344# 0.06fF
C53419 PAND2X1_23/Y POR2X1_140/A 0.02fF
C53420 POR2X1_102/Y POR2X1_131/A 0.04fF
C53421 POR2X1_774/CTRL VDD 0.00fF
C53422 POR2X1_13/A POR2X1_597/CTRL 0.01fF
C53423 POR2X1_68/A POR2X1_222/Y 0.03fF
C53424 PAND2X1_492/O POR2X1_123/A 0.04fF
C53425 POR2X1_192/Y POR2X1_350/B 0.81fF
C53426 POR2X1_32/O POR2X1_29/Y 0.03fF
C53427 VDD POR2X1_128/B 0.02fF
C53428 POR2X1_174/A POR2X1_337/Y 0.07fF
C53429 PAND2X1_552/A PAND2X1_569/Y 0.15fF
C53430 PAND2X1_523/CTRL PAND2X1_844/B 0.01fF
C53431 POR2X1_414/CTRL2 POR2X1_4/Y 0.01fF
C53432 POR2X1_66/A PAND2X1_517/O 0.08fF
C53433 POR2X1_79/A PAND2X1_854/A 0.02fF
C53434 POR2X1_510/A POR2X1_35/Y 0.01fF
C53435 POR2X1_7/B PAND2X1_347/a_56_28# 0.00fF
C53436 POR2X1_16/A POR2X1_689/CTRL 0.01fF
C53437 PAND2X1_278/O POR2X1_559/A 0.04fF
C53438 POR2X1_633/A POR2X1_294/A 0.14fF
C53439 PAND2X1_834/CTRL2 POR2X1_37/Y 0.01fF
C53440 POR2X1_49/Y PAND2X1_358/A 0.07fF
C53441 POR2X1_834/Y POR2X1_480/A 0.10fF
C53442 PAND2X1_41/B POR2X1_186/B 0.14fF
C53443 POR2X1_66/A POR2X1_169/A 0.03fF
C53444 POR2X1_686/B POR2X1_687/A 0.01fF
C53445 POR2X1_56/B POR2X1_387/Y 0.10fF
C53446 POR2X1_49/Y POR2X1_599/O 0.01fF
C53447 PAND2X1_3/A D_INPUT_4 0.12fF
C53448 POR2X1_66/A PAND2X1_529/CTRL 0.03fF
C53449 POR2X1_188/A POR2X1_851/a_76_344# 0.00fF
C53450 POR2X1_65/A PAND2X1_779/CTRL2 0.03fF
C53451 POR2X1_78/B POR2X1_339/O 0.02fF
C53452 PAND2X1_217/CTRL2 POR2X1_599/A 0.32fF
C53453 PAND2X1_360/O POR2X1_385/Y 0.04fF
C53454 PAND2X1_863/A POR2X1_102/Y 0.05fF
C53455 POR2X1_123/A PAND2X1_132/CTRL 0.02fF
C53456 POR2X1_74/Y PAND2X1_76/O 0.04fF
C53457 POR2X1_154/a_56_344# POR2X1_855/B 0.00fF
C53458 POR2X1_68/A POR2X1_532/A 0.08fF
C53459 POR2X1_413/A PAND2X1_647/CTRL 0.01fF
C53460 POR2X1_786/Y PAND2X1_69/A 1.10fF
C53461 POR2X1_502/A PAND2X1_94/A 0.07fF
C53462 POR2X1_96/A POR2X1_96/CTRL2 0.01fF
C53463 POR2X1_7/B PAND2X1_112/CTRL2 0.00fF
C53464 POR2X1_238/Y POR2X1_91/Y 1.49fF
C53465 POR2X1_523/A POR2X1_750/A 0.02fF
C53466 POR2X1_383/A POR2X1_717/Y 0.03fF
C53467 PAND2X1_613/a_76_28# PAND2X1_52/B 0.05fF
C53468 PAND2X1_652/CTRL2 PAND2X1_557/A 0.01fF
C53469 POR2X1_520/B VDD 0.02fF
C53470 PAND2X1_299/CTRL2 POR2X1_188/Y 0.01fF
C53471 POR2X1_617/a_56_344# POR2X1_408/Y 0.03fF
C53472 POR2X1_52/A POR2X1_164/Y 0.12fF
C53473 PAND2X1_408/Y POR2X1_407/Y 0.78fF
C53474 PAND2X1_55/Y PAND2X1_312/m4_208_n4# 0.15fF
C53475 POR2X1_484/a_16_28# POR2X1_39/B 0.03fF
C53476 POR2X1_271/A POR2X1_256/CTRL2 0.08fF
C53477 POR2X1_7/B POR2X1_375/O 0.02fF
C53478 POR2X1_740/Y POR2X1_725/Y 0.07fF
C53479 PAND2X1_94/A POR2X1_247/CTRL 0.10fF
C53480 INPUT_1 POR2X1_624/CTRL2 0.01fF
C53481 POR2X1_416/B POR2X1_496/Y 0.07fF
C53482 POR2X1_857/B PAND2X1_503/CTRL 0.03fF
C53483 POR2X1_62/Y PAND2X1_85/Y 0.29fF
C53484 PAND2X1_140/A PAND2X1_357/Y 0.03fF
C53485 POR2X1_710/CTRL POR2X1_713/B 0.01fF
C53486 PAND2X1_691/Y POR2X1_761/CTRL 0.10fF
C53487 POR2X1_45/Y PAND2X1_723/A 0.07fF
C53488 POR2X1_57/A PAND2X1_645/B 0.08fF
C53489 POR2X1_22/a_16_28# POR2X1_260/A 0.03fF
C53490 POR2X1_113/Y PAND2X1_153/CTRL2 0.00fF
C53491 PAND2X1_173/O POR2X1_570/B 0.05fF
C53492 POR2X1_394/A POR2X1_817/A 0.03fF
C53493 POR2X1_146/Y VDD 0.06fF
C53494 POR2X1_102/Y PAND2X1_861/B 0.02fF
C53495 POR2X1_57/A INPUT_6 0.01fF
C53496 POR2X1_41/B PAND2X1_853/B 0.03fF
C53497 POR2X1_38/B POR2X1_380/Y 0.02fF
C53498 POR2X1_71/Y POR2X1_394/A 0.02fF
C53499 POR2X1_709/CTRL2 PAND2X1_69/A 0.00fF
C53500 PAND2X1_865/Y PAND2X1_787/Y 0.12fF
C53501 POR2X1_130/A POR2X1_557/CTRL2 0.01fF
C53502 PAND2X1_474/A PAND2X1_860/a_16_344# 0.02fF
C53503 POR2X1_13/A PAND2X1_851/CTRL2 0.03fF
C53504 POR2X1_7/B POR2X1_129/Y 0.03fF
C53505 PAND2X1_580/B POR2X1_385/Y 0.03fF
C53506 POR2X1_13/A POR2X1_595/O 0.12fF
C53507 POR2X1_754/Y POR2X1_90/CTRL2 0.01fF
C53508 POR2X1_284/B POR2X1_188/Y 0.01fF
C53509 POR2X1_205/A PAND2X1_60/B 0.07fF
C53510 PAND2X1_6/A PAND2X1_748/O 0.00fF
C53511 POR2X1_394/A POR2X1_42/Y 0.06fF
C53512 POR2X1_416/B PAND2X1_733/A 0.09fF
C53513 PAND2X1_23/Y POR2X1_544/Y 0.01fF
C53514 POR2X1_860/a_16_28# POR2X1_572/B 0.02fF
C53515 INPUT_1 POR2X1_409/CTRL2 0.01fF
C53516 INPUT_0 PAND2X1_517/CTRL 0.07fF
C53517 POR2X1_814/A POR2X1_435/B 0.35fF
C53518 PAND2X1_60/B POR2X1_366/A 0.06fF
C53519 POR2X1_216/a_16_28# PAND2X1_60/B 0.01fF
C53520 PAND2X1_414/CTRL INPUT_3 0.01fF
C53521 POR2X1_220/Y POR2X1_540/Y 1.40fF
C53522 POR2X1_390/B POR2X1_68/B 0.02fF
C53523 PAND2X1_659/Y POR2X1_7/B 0.03fF
C53524 POR2X1_578/Y POR2X1_192/B 3.24fF
C53525 POR2X1_110/O POR2X1_293/Y 0.15fF
C53526 PAND2X1_467/Y POR2X1_426/Y 0.01fF
C53527 PAND2X1_233/O POR2X1_66/A 0.06fF
C53528 POR2X1_196/Y POR2X1_260/A 2.48fF
C53529 POR2X1_509/A POR2X1_227/CTRL 0.09fF
C53530 POR2X1_57/A PAND2X1_737/B 0.79fF
C53531 POR2X1_609/Y PAND2X1_403/O 0.00fF
C53532 VDD POR2X1_561/B 0.04fF
C53533 POR2X1_57/A PAND2X1_216/B 0.03fF
C53534 VDD POR2X1_343/O 0.00fF
C53535 POR2X1_270/Y POR2X1_458/Y 0.07fF
C53536 POR2X1_96/Y POR2X1_7/B 0.01fF
C53537 POR2X1_346/CTRL2 POR2X1_507/A 0.03fF
C53538 PAND2X1_6/Y PAND2X1_482/CTRL 0.02fF
C53539 POR2X1_538/A POR2X1_337/A 0.10fF
C53540 PAND2X1_687/B POR2X1_7/B 0.01fF
C53541 POR2X1_121/A POR2X1_294/A 0.02fF
C53542 PAND2X1_483/CTRL POR2X1_7/A 0.01fF
C53543 POR2X1_23/Y PAND2X1_717/A 0.06fF
C53544 PAND2X1_228/a_76_28# POR2X1_7/Y 0.01fF
C53545 POR2X1_548/O PAND2X1_52/B 0.02fF
C53546 PAND2X1_501/CTRL PAND2X1_735/Y 0.06fF
C53547 PAND2X1_730/A POR2X1_816/A 0.06fF
C53548 PAND2X1_242/Y POR2X1_72/B 0.05fF
C53549 POR2X1_804/A POR2X1_512/CTRL2 0.46fF
C53550 POR2X1_16/A POR2X1_315/Y 0.01fF
C53551 POR2X1_222/Y POR2X1_735/m4_208_n4# 0.15fF
C53552 PAND2X1_139/CTRL2 POR2X1_184/Y 0.00fF
C53553 POR2X1_560/CTRL2 POR2X1_844/B 0.01fF
C53554 POR2X1_8/Y PAND2X1_63/B 0.60fF
C53555 PAND2X1_794/B PAND2X1_643/A 0.03fF
C53556 PAND2X1_6/A POR2X1_4/Y 0.21fF
C53557 POR2X1_16/O PAND2X1_733/A 0.01fF
C53558 PAND2X1_137/Y POR2X1_77/Y 0.01fF
C53559 POR2X1_57/A PAND2X1_359/Y 0.02fF
C53560 POR2X1_78/B POR2X1_717/B 0.06fF
C53561 POR2X1_290/CTRL POR2X1_234/A 0.01fF
C53562 POR2X1_508/B POR2X1_508/a_16_28# 0.02fF
C53563 POR2X1_228/Y POR2X1_186/B 0.03fF
C53564 PAND2X1_175/B POR2X1_153/Y 0.03fF
C53565 POR2X1_750/Y POR2X1_260/A 0.05fF
C53566 POR2X1_147/O POR2X1_435/Y 0.05fF
C53567 PAND2X1_360/Y PAND2X1_843/Y 0.01fF
C53568 POR2X1_57/A PAND2X1_138/O 0.02fF
C53569 POR2X1_726/Y POR2X1_731/A 0.03fF
C53570 PAND2X1_69/A PAND2X1_396/O 0.02fF
C53571 POR2X1_46/Y PAND2X1_327/a_16_344# 0.02fF
C53572 PAND2X1_6/Y POR2X1_840/Y 0.14fF
C53573 PAND2X1_476/A POR2X1_73/Y 0.03fF
C53574 POR2X1_774/A POR2X1_725/Y 0.03fF
C53575 PAND2X1_797/Y POR2X1_90/Y 0.53fF
C53576 POR2X1_324/a_56_344# POR2X1_568/Y 0.03fF
C53577 POR2X1_119/Y PAND2X1_787/A 0.03fF
C53578 POR2X1_456/B POR2X1_741/B 0.01fF
C53579 POR2X1_343/Y POR2X1_833/O 0.04fF
C53580 PAND2X1_779/O PAND2X1_549/B 0.02fF
C53581 POR2X1_416/B PAND2X1_514/Y 0.04fF
C53582 POR2X1_145/a_76_344# POR2X1_77/Y 0.01fF
C53583 POR2X1_561/B PAND2X1_32/B 0.00fF
C53584 POR2X1_180/a_16_28# POR2X1_180/A 0.03fF
C53585 POR2X1_343/O PAND2X1_32/B 0.03fF
C53586 POR2X1_556/A POR2X1_269/O 0.02fF
C53587 PAND2X1_731/O POR2X1_39/B 0.03fF
C53588 POR2X1_313/Y POR2X1_314/Y 0.00fF
C53589 POR2X1_83/B PAND2X1_201/CTRL 0.02fF
C53590 POR2X1_532/CTRL2 PAND2X1_60/B 0.09fF
C53591 POR2X1_248/CTRL POR2X1_77/Y 0.01fF
C53592 PAND2X1_276/a_76_28# POR2X1_677/Y 0.07fF
C53593 POR2X1_383/A PAND2X1_281/a_76_28# 0.01fF
C53594 POR2X1_411/B POR2X1_432/O 0.01fF
C53595 POR2X1_99/B POR2X1_259/CTRL 0.00fF
C53596 PAND2X1_9/Y POR2X1_29/A 0.22fF
C53597 PAND2X1_476/A PAND2X1_244/B 0.03fF
C53598 POR2X1_101/Y POR2X1_4/Y 0.05fF
C53599 PAND2X1_621/O POR2X1_616/Y 0.02fF
C53600 POR2X1_866/A POR2X1_807/CTRL2 0.06fF
C53601 PAND2X1_601/O POR2X1_66/A 0.01fF
C53602 POR2X1_736/A POR2X1_724/A 0.07fF
C53603 POR2X1_447/B POR2X1_260/A 0.07fF
C53604 PAND2X1_493/O POR2X1_394/A 0.08fF
C53605 POR2X1_220/O POR2X1_220/B 0.02fF
C53606 POR2X1_52/A POR2X1_485/a_16_28# 0.00fF
C53607 POR2X1_814/B POR2X1_621/a_76_344# 0.00fF
C53608 PAND2X1_569/B PAND2X1_326/B 0.05fF
C53609 POR2X1_169/O POR2X1_191/Y 0.26fF
C53610 POR2X1_169/a_56_344# POR2X1_192/B 0.00fF
C53611 POR2X1_327/Y PAND2X1_48/A 0.04fF
C53612 PAND2X1_366/O PAND2X1_354/Y 0.05fF
C53613 POR2X1_813/a_16_28# POR2X1_669/B 0.01fF
C53614 PAND2X1_424/CTRL2 PAND2X1_72/A 0.01fF
C53615 POR2X1_326/A POR2X1_652/A 0.03fF
C53616 POR2X1_633/a_76_344# POR2X1_734/A 0.03fF
C53617 PAND2X1_640/B POR2X1_37/Y 0.03fF
C53618 POR2X1_49/Y POR2X1_441/Y 0.04fF
C53619 POR2X1_45/Y PAND2X1_860/A 0.03fF
C53620 POR2X1_800/CTRL POR2X1_452/Y 0.01fF
C53621 POR2X1_335/O POR2X1_814/A 0.01fF
C53622 POR2X1_41/B POR2X1_827/CTRL 0.00fF
C53623 POR2X1_612/Y POR2X1_413/CTRL2 0.05fF
C53624 POR2X1_16/a_16_28# POR2X1_42/Y 0.03fF
C53625 POR2X1_504/Y POR2X1_20/B 0.04fF
C53626 POR2X1_647/a_16_28# POR2X1_646/Y 0.02fF
C53627 POR2X1_291/CTRL POR2X1_39/B 0.01fF
C53628 PAND2X1_639/B PAND2X1_635/Y 0.11fF
C53629 POR2X1_428/Y POR2X1_748/A 0.17fF
C53630 POR2X1_864/A PAND2X1_65/B 0.00fF
C53631 POR2X1_446/B POR2X1_330/Y 0.05fF
C53632 PAND2X1_48/A PAND2X1_692/a_16_344# 0.01fF
C53633 POR2X1_24/Y POR2X1_94/A 0.03fF
C53634 POR2X1_801/O POR2X1_452/Y 0.01fF
C53635 POR2X1_66/Y POR2X1_852/B 0.05fF
C53636 POR2X1_734/B POR2X1_121/B 0.01fF
C53637 POR2X1_483/A POR2X1_541/B 0.11fF
C53638 POR2X1_669/B POR2X1_754/Y 0.10fF
C53639 POR2X1_612/Y POR2X1_607/O 0.04fF
C53640 PAND2X1_58/A POR2X1_66/A 0.10fF
C53641 POR2X1_455/CTRL POR2X1_341/A 0.06fF
C53642 POR2X1_83/B D_INPUT_0 0.06fF
C53643 PAND2X1_446/Y POR2X1_236/Y 0.03fF
C53644 POR2X1_130/A POR2X1_556/A 0.03fF
C53645 POR2X1_502/A POR2X1_460/Y 0.04fF
C53646 PAND2X1_473/Y POR2X1_411/B 0.03fF
C53647 POR2X1_666/a_76_344# POR2X1_32/A 0.02fF
C53648 POR2X1_808/A POR2X1_678/Y 0.50fF
C53649 POR2X1_566/A POR2X1_556/A 0.03fF
C53650 PAND2X1_853/B POR2X1_77/Y 0.03fF
C53651 POR2X1_852/B POR2X1_629/O 0.09fF
C53652 PAND2X1_39/B VDD 2.16fF
C53653 PAND2X1_444/CTRL2 POR2X1_236/Y 0.01fF
C53654 POR2X1_558/B POR2X1_860/A 0.02fF
C53655 PAND2X1_48/B PAND2X1_417/O 0.02fF
C53656 PAND2X1_699/CTRL POR2X1_43/B 0.00fF
C53657 POR2X1_220/CTRL2 POR2X1_220/Y 0.00fF
C53658 POR2X1_123/O POR2X1_556/A 0.01fF
C53659 PAND2X1_618/Y VDD 0.12fF
C53660 POR2X1_96/A POR2X1_679/A 0.03fF
C53661 POR2X1_99/A POR2X1_590/A 0.01fF
C53662 PAND2X1_444/CTRL VDD 0.00fF
C53663 POR2X1_855/CTRL POR2X1_855/A 0.00fF
C53664 POR2X1_60/A PAND2X1_786/O 0.04fF
C53665 POR2X1_251/A POR2X1_60/A 0.06fF
C53666 PAND2X1_432/O POR2X1_811/B 0.13fF
C53667 POR2X1_866/B POR2X1_801/B 0.01fF
C53668 POR2X1_60/A POR2X1_72/B 23.07fF
C53669 POR2X1_411/B POR2X1_395/a_16_28# 0.04fF
C53670 POR2X1_274/CTRL POR2X1_325/A 0.09fF
C53671 POR2X1_792/CTRL PAND2X1_90/Y 0.04fF
C53672 PAND2X1_9/Y POR2X1_204/CTRL2 0.00fF
C53673 POR2X1_376/B POR2X1_432/O 0.16fF
C53674 PAND2X1_666/CTRL2 POR2X1_130/A 0.09fF
C53675 POR2X1_818/Y POR2X1_546/A 0.08fF
C53676 POR2X1_416/B POR2X1_746/a_16_28# -0.00fF
C53677 PAND2X1_23/Y POR2X1_54/Y 0.09fF
C53678 POR2X1_634/A POR2X1_634/a_16_28# 0.09fF
C53679 POR2X1_433/Y POR2X1_20/B 1.53fF
C53680 PAND2X1_224/O POR2X1_566/B 0.12fF
C53681 PAND2X1_39/B POR2X1_741/Y 0.06fF
C53682 POR2X1_14/Y POR2X1_720/A 0.03fF
C53683 POR2X1_130/A PAND2X1_591/O 0.03fF
C53684 PAND2X1_836/CTRL POR2X1_20/B 0.01fF
C53685 POR2X1_102/Y PAND2X1_219/B 0.01fF
C53686 POR2X1_327/CTRL2 POR2X1_558/B 0.00fF
C53687 POR2X1_602/B POR2X1_808/A 0.02fF
C53688 POR2X1_260/B POR2X1_193/A 0.04fF
C53689 POR2X1_260/B POR2X1_579/Y 0.03fF
C53690 POR2X1_846/O POR2X1_129/Y 0.01fF
C53691 POR2X1_454/A POR2X1_785/A 0.03fF
C53692 POR2X1_41/B POR2X1_23/Y 0.42fF
C53693 PAND2X1_23/Y POR2X1_202/A 0.06fF
C53694 POR2X1_96/A POR2X1_626/CTRL2 0.00fF
C53695 POR2X1_496/Y PAND2X1_512/Y 0.08fF
C53696 POR2X1_66/B POR2X1_287/B 0.03fF
C53697 POR2X1_595/a_16_28# POR2X1_250/A 0.05fF
C53698 POR2X1_556/A POR2X1_573/A 0.03fF
C53699 POR2X1_82/CTRL POR2X1_14/Y 0.01fF
C53700 PAND2X1_640/B POR2X1_293/Y 0.06fF
C53701 PAND2X1_5/CTRL INPUT_3 0.01fF
C53702 POR2X1_20/B D_INPUT_6 0.01fF
C53703 POR2X1_628/Y POR2X1_90/Y 0.03fF
C53704 POR2X1_32/A POR2X1_88/Y 0.03fF
C53705 POR2X1_805/Y VDD 0.96fF
C53706 POR2X1_840/B POR2X1_341/A 0.10fF
C53707 PAND2X1_246/O PAND2X1_63/B 0.06fF
C53708 PAND2X1_469/B POR2X1_273/O 0.02fF
C53709 POR2X1_37/Y POR2X1_7/B 0.05fF
C53710 POR2X1_416/B POR2X1_43/O 0.00fF
C53711 PAND2X1_39/B PAND2X1_32/B 0.36fF
C53712 POR2X1_658/CTRL PAND2X1_60/B 0.00fF
C53713 POR2X1_181/CTRL2 POR2X1_181/A 0.01fF
C53714 POR2X1_497/CTRL PAND2X1_501/B 0.01fF
C53715 POR2X1_43/B POR2X1_260/B 0.03fF
C53716 D_INPUT_2 POR2X1_612/Y 0.01fF
C53717 PAND2X1_556/CTRL VDD -0.00fF
C53718 PAND2X1_582/O PAND2X1_581/Y -0.00fF
C53719 PAND2X1_416/O PAND2X1_69/A 0.01fF
C53720 PAND2X1_635/O POR2X1_428/Y 0.03fF
C53721 POR2X1_516/Y INPUT_0 0.07fF
C53722 PAND2X1_20/A VDD 2.64fF
C53723 PAND2X1_654/CTRL POR2X1_409/B 0.01fF
C53724 PAND2X1_293/O PAND2X1_58/A 0.25fF
C53725 POR2X1_779/A POR2X1_866/A 0.02fF
C53726 PAND2X1_621/Y PAND2X1_381/Y 0.03fF
C53727 PAND2X1_268/a_16_344# PAND2X1_69/A 0.02fF
C53728 POR2X1_84/A POR2X1_35/Y 0.15fF
C53729 POR2X1_502/A PAND2X1_11/Y 0.05fF
C53730 POR2X1_493/A PAND2X1_519/CTRL 0.01fF
C53731 POR2X1_20/B PAND2X1_840/CTRL 0.00fF
C53732 POR2X1_461/B POR2X1_461/A 0.00fF
C53733 POR2X1_614/A POR2X1_260/B 0.33fF
C53734 PAND2X1_23/Y POR2X1_346/A 0.02fF
C53735 D_INPUT_0 POR2X1_565/CTRL2 0.01fF
C53736 POR2X1_383/A POR2X1_649/O 0.01fF
C53737 POR2X1_174/B POR2X1_852/A 0.08fF
C53738 PAND2X1_793/Y POR2X1_102/Y 0.03fF
C53739 POR2X1_227/B POR2X1_854/B 0.26fF
C53740 POR2X1_660/A POR2X1_362/B 0.01fF
C53741 POR2X1_257/A POR2X1_695/CTRL2 0.03fF
C53742 PAND2X1_82/O PAND2X1_39/B 0.09fF
C53743 POR2X1_83/B PAND2X1_364/CTRL2 0.01fF
C53744 PAND2X1_601/O POR2X1_532/A 0.07fF
C53745 POR2X1_669/B POR2X1_42/Y 0.30fF
C53746 POR2X1_444/O POR2X1_568/Y 0.08fF
C53747 PAND2X1_57/B POR2X1_794/B 2.23fF
C53748 POR2X1_810/a_16_28# POR2X1_636/B 0.01fF
C53749 POR2X1_39/O POR2X1_236/Y 0.03fF
C53750 POR2X1_293/a_76_344# POR2X1_5/Y 0.01fF
C53751 POR2X1_659/A POR2X1_318/A 0.03fF
C53752 POR2X1_13/A POR2X1_272/CTRL 0.01fF
C53753 POR2X1_60/A PAND2X1_714/CTRL 0.05fF
C53754 POR2X1_174/B PAND2X1_226/a_16_344# 0.03fF
C53755 POR2X1_65/A PAND2X1_347/Y 0.03fF
C53756 PAND2X1_473/B PAND2X1_736/CTRL2 0.11fF
C53757 POR2X1_590/A PAND2X1_530/O 0.04fF
C53758 POR2X1_48/A PAND2X1_731/O 0.01fF
C53759 POR2X1_814/B VDD 3.02fF
C53760 POR2X1_102/Y PAND2X1_219/CTRL 0.01fF
C53761 PAND2X1_94/A POR2X1_78/a_16_28# 0.01fF
C53762 POR2X1_502/A PAND2X1_278/CTRL 0.01fF
C53763 POR2X1_68/A POR2X1_660/Y 0.05fF
C53764 PAND2X1_56/Y POR2X1_555/B 0.00fF
C53765 PAND2X1_363/Y VDD 0.32fF
C53766 POR2X1_218/A POR2X1_296/B 0.05fF
C53767 POR2X1_413/A POR2X1_607/CTRL2 0.01fF
C53768 POR2X1_65/A PAND2X1_564/O 0.03fF
C53769 POR2X1_734/A POR2X1_121/Y 0.07fF
C53770 D_INPUT_0 POR2X1_522/Y 0.02fF
C53771 PAND2X1_96/B POR2X1_66/A 0.81fF
C53772 POR2X1_856/B POR2X1_341/Y 0.03fF
C53773 POR2X1_270/Y POR2X1_724/A 0.03fF
C53774 PAND2X1_422/O POR2X1_260/B 0.07fF
C53775 POR2X1_376/Y PAND2X1_8/Y 0.03fF
C53776 POR2X1_853/CTRL PAND2X1_41/B 0.09fF
C53777 PAND2X1_283/O POR2X1_78/A 0.08fF
C53778 PAND2X1_738/Y PAND2X1_180/CTRL2 0.14fF
C53779 PAND2X1_53/CTRL PAND2X1_48/A 0.13fF
C53780 PAND2X1_20/A POR2X1_741/Y 0.03fF
C53781 PAND2X1_859/a_16_344# INPUT_0 0.04fF
C53782 POR2X1_409/B POR2X1_38/Y 0.07fF
C53783 POR2X1_102/Y POR2X1_665/Y 0.03fF
C53784 POR2X1_12/A POR2X1_158/B 0.06fF
C53785 POR2X1_687/A POR2X1_803/a_16_28# 0.03fF
C53786 POR2X1_325/A VDD 0.46fF
C53787 POR2X1_78/O POR2X1_78/A 0.18fF
C53788 PAND2X1_667/CTRL INPUT_0 0.05fF
C53789 POR2X1_20/Y POR2X1_14/Y 0.16fF
C53790 POR2X1_278/Y PAND2X1_473/B 0.07fF
C53791 POR2X1_114/a_76_344# POR2X1_590/A 0.01fF
C53792 PAND2X1_23/Y PAND2X1_23/CTRL 0.00fF
C53793 POR2X1_66/B POR2X1_61/B 0.37fF
C53794 PAND2X1_7/Y POR2X1_294/B 0.03fF
C53795 PAND2X1_824/O POR2X1_567/B 0.02fF
C53796 POR2X1_805/Y PAND2X1_32/B 0.01fF
C53797 D_INPUT_3 POR2X1_14/O 0.18fF
C53798 POR2X1_302/A POR2X1_302/B 0.18fF
C53799 POR2X1_810/CTRL2 POR2X1_750/B 0.01fF
C53800 POR2X1_5/Y POR2X1_395/CTRL2 0.00fF
C53801 PAND2X1_454/B PAND2X1_308/Y 0.65fF
C53802 POR2X1_96/Y PAND2X1_206/B 0.07fF
C53803 PAND2X1_616/CTRL PAND2X1_6/A 0.01fF
C53804 PAND2X1_6/Y POR2X1_783/CTRL 0.01fF
C53805 POR2X1_448/Y POR2X1_532/Y 0.09fF
C53806 POR2X1_41/B POR2X1_368/CTRL2 0.02fF
C53807 PAND2X1_319/B PAND2X1_212/B 0.03fF
C53808 PAND2X1_20/A PAND2X1_32/B 0.59fF
C53809 POR2X1_164/CTRL2 POR2X1_40/Y 0.01fF
C53810 PAND2X1_817/O D_INPUT_1 0.01fF
C53811 PAND2X1_808/Y POR2X1_488/CTRL 0.01fF
C53812 PAND2X1_58/A POR2X1_532/A 0.13fF
C53813 POR2X1_79/Y PAND2X1_740/Y 0.00fF
C53814 PAND2X1_658/CTRL2 POR2X1_816/A 0.01fF
C53815 PAND2X1_96/B POR2X1_634/CTRL2 0.05fF
C53816 PAND2X1_479/B PAND2X1_579/B 0.02fF
C53817 PAND2X1_94/A POR2X1_493/A 0.05fF
C53818 PAND2X1_90/Y PAND2X1_176/a_16_344# 0.05fF
C53819 POR2X1_46/Y PAND2X1_332/a_76_28# 0.04fF
C53820 POR2X1_687/A POR2X1_678/Y 0.04fF
C53821 POR2X1_814/B POR2X1_741/Y 0.03fF
C53822 POR2X1_748/A POR2X1_748/CTRL2 0.00fF
C53823 VDD POR2X1_513/B 0.51fF
C53824 POR2X1_423/Y POR2X1_255/Y 0.54fF
C53825 PAND2X1_639/a_16_344# POR2X1_386/Y 0.04fF
C53826 POR2X1_82/CTRL POR2X1_55/Y 0.01fF
C53827 POR2X1_52/A PAND2X1_473/Y 0.02fF
C53828 PAND2X1_669/CTRL2 POR2X1_750/Y 0.14fF
C53829 POR2X1_763/A POR2X1_700/a_16_28# 0.06fF
C53830 PAND2X1_469/B PAND2X1_787/a_16_344# 0.07fF
C53831 POR2X1_208/Y PAND2X1_41/B 0.09fF
C53832 POR2X1_741/Y POR2X1_733/CTRL 0.00fF
C53833 POR2X1_479/B POR2X1_249/Y 0.03fF
C53834 PAND2X1_65/Y POR2X1_35/Y 0.03fF
C53835 POR2X1_89/CTRL POR2X1_394/A 0.07fF
C53836 POR2X1_435/Y POR2X1_802/B 0.98fF
C53837 PAND2X1_805/m4_208_n4# POR2X1_7/B 0.09fF
C53838 POR2X1_454/A POR2X1_186/B 0.03fF
C53839 PAND2X1_250/O PAND2X1_32/B 0.01fF
C53840 POR2X1_23/Y PAND2X1_308/Y 0.05fF
C53841 INPUT_1 POR2X1_409/B 0.13fF
C53842 POR2X1_741/Y POR2X1_325/A 0.03fF
C53843 PAND2X1_417/CTRL2 POR2X1_169/A 0.06fF
C53844 POR2X1_814/B PAND2X1_32/B 15.85fF
C53845 PAND2X1_79/Y PAND2X1_41/B 0.03fF
C53846 GATE_479 POR2X1_694/a_76_344# 0.01fF
C53847 POR2X1_329/A POR2X1_522/CTRL 0.01fF
C53848 POR2X1_194/A POR2X1_194/O 0.13fF
C53849 POR2X1_43/Y POR2X1_827/CTRL2 0.00fF
C53850 PAND2X1_478/CTRL2 PAND2X1_480/B 0.06fF
C53851 PAND2X1_499/Y POR2X1_56/Y 0.25fF
C53852 PAND2X1_347/Y PAND2X1_190/Y 0.05fF
C53853 POR2X1_673/A PAND2X1_6/A 0.03fF
C53854 POR2X1_96/Y POR2X1_65/Y 1.34fF
C53855 PAND2X1_575/A PAND2X1_735/Y 0.01fF
C53856 POR2X1_7/B POR2X1_293/Y 0.07fF
C53857 PAND2X1_651/Y PAND2X1_84/CTRL2 0.03fF
C53858 POR2X1_267/CTRL2 POR2X1_260/A 0.12fF
C53859 POR2X1_119/Y PAND2X1_469/O 0.16fF
C53860 POR2X1_409/B POR2X1_153/Y 0.14fF
C53861 POR2X1_383/A POR2X1_330/Y 0.21fF
C53862 PAND2X1_490/O PAND2X1_85/Y 0.00fF
C53863 POR2X1_283/A POR2X1_40/Y 0.13fF
C53864 POR2X1_8/Y POR2X1_32/A 0.03fF
C53865 PAND2X1_779/Y VDD 0.06fF
C53866 POR2X1_52/A PAND2X1_736/A 0.17fF
C53867 PAND2X1_675/A POR2X1_79/Y 0.03fF
C53868 POR2X1_325/A PAND2X1_32/B 0.01fF
C53869 PAND2X1_55/Y POR2X1_193/A 0.03fF
C53870 PAND2X1_655/Y POR2X1_690/Y 0.04fF
C53871 PAND2X1_55/Y POR2X1_579/Y 0.03fF
C53872 PAND2X1_418/CTRL2 PAND2X1_52/B 0.03fF
C53873 PAND2X1_468/CTRL PAND2X1_798/B 0.01fF
C53874 POR2X1_65/A PAND2X1_551/CTRL 0.01fF
C53875 PAND2X1_20/A POR2X1_673/Y 0.03fF
C53876 POR2X1_10/O POR2X1_83/B 0.17fF
C53877 PAND2X1_55/Y POR2X1_445/m4_208_n4# 0.15fF
C53878 POR2X1_20/Y PAND2X1_472/B 0.09fF
C53879 POR2X1_52/A POR2X1_823/CTRL2 0.01fF
C53880 PAND2X1_228/CTRL PAND2X1_197/Y 0.00fF
C53881 VDD PAND2X1_509/CTRL 0.00fF
C53882 POR2X1_407/A PAND2X1_498/CTRL2 0.01fF
C53883 POR2X1_459/a_16_28# POR2X1_459/A 0.09fF
C53884 PAND2X1_716/CTRL PAND2X1_364/B 0.07fF
C53885 POR2X1_140/B POR2X1_554/Y 0.11fF
C53886 POR2X1_157/a_16_28# INPUT_5 0.02fF
C53887 POR2X1_786/CTRL PAND2X1_60/B 0.01fF
C53888 PAND2X1_478/a_76_28# POR2X1_46/Y 0.01fF
C53889 PAND2X1_4/CTRL VDD 0.00fF
C53890 PAND2X1_805/A PAND2X1_367/A 0.05fF
C53891 POR2X1_515/CTRL PAND2X1_60/B 0.00fF
C53892 POR2X1_435/Y POR2X1_532/A 0.09fF
C53893 POR2X1_16/A PAND2X1_558/Y 0.05fF
C53894 PAND2X1_862/Y POR2X1_32/A 0.00fF
C53895 POR2X1_364/A POR2X1_776/B 0.19fF
C53896 PAND2X1_766/O POR2X1_260/A 0.02fF
C53897 POR2X1_302/CTRL POR2X1_383/A 0.03fF
C53898 POR2X1_860/A POR2X1_362/A 0.00fF
C53899 POR2X1_416/Y POR2X1_232/a_16_28# 0.02fF
C53900 PAND2X1_6/Y PAND2X1_604/O 0.01fF
C53901 PAND2X1_63/Y POR2X1_404/Y 0.03fF
C53902 PAND2X1_96/B POR2X1_792/B 0.01fF
C53903 POR2X1_614/A PAND2X1_55/Y 0.22fF
C53904 POR2X1_32/A POR2X1_385/Y 0.03fF
C53905 PAND2X1_96/B POR2X1_802/B 0.01fF
C53906 POR2X1_814/B POR2X1_673/Y 0.02fF
C53907 POR2X1_656/a_16_28# POR2X1_737/A 0.02fF
C53908 PAND2X1_183/O POR2X1_540/A 0.02fF
C53909 POR2X1_700/CTRL PAND2X1_711/A 0.01fF
C53910 POR2X1_252/Y POR2X1_669/B 0.21fF
C53911 PAND2X1_124/Y PAND2X1_198/CTRL 0.09fF
C53912 PAND2X1_207/CTRL PAND2X1_207/A 0.01fF
C53913 PAND2X1_71/CTRL2 PAND2X1_111/B 0.01fF
C53914 PAND2X1_107/O PAND2X1_65/B 0.04fF
C53915 POR2X1_439/m4_208_n4# POR2X1_456/B 0.09fF
C53916 POR2X1_795/a_16_28# POR2X1_786/Y -0.00fF
C53917 POR2X1_750/B POR2X1_129/Y 0.07fF
C53918 PAND2X1_724/O PAND2X1_724/B 0.00fF
C53919 INPUT_1 POR2X1_29/CTRL2 0.01fF
C53920 POR2X1_218/A POR2X1_267/Y 0.00fF
C53921 PAND2X1_182/CTRL2 PAND2X1_357/Y 0.02fF
C53922 PAND2X1_55/Y POR2X1_38/B 0.06fF
C53923 PAND2X1_736/A PAND2X1_186/O 0.06fF
C53924 POR2X1_334/Y POR2X1_186/Y 0.07fF
C53925 POR2X1_356/A PAND2X1_173/O 0.02fF
C53926 PAND2X1_57/B PAND2X1_765/CTRL 0.01fF
C53927 PAND2X1_844/Y PAND2X1_99/Y 0.02fF
C53928 PAND2X1_96/B POR2X1_222/Y 0.10fF
C53929 POR2X1_9/Y PAND2X1_87/a_16_344# 0.02fF
C53930 PAND2X1_6/A POR2X1_816/A 0.03fF
C53931 PAND2X1_370/O POR2X1_309/Y 0.02fF
C53932 PAND2X1_599/a_76_28# PAND2X1_69/A 0.02fF
C53933 POR2X1_566/A POR2X1_566/B 0.02fF
C53934 PAND2X1_20/A POR2X1_560/CTRL 0.01fF
C53935 POR2X1_408/Y POR2X1_7/B 0.08fF
C53936 POR2X1_566/A POR2X1_180/A 0.07fF
C53937 PAND2X1_23/Y POR2X1_544/O 0.01fF
C53938 POR2X1_23/Y POR2X1_77/Y 0.27fF
C53939 PAND2X1_6/A D_INPUT_1 0.18fF
C53940 POR2X1_66/A POR2X1_342/B 0.02fF
C53941 POR2X1_72/B POR2X1_373/CTRL2 0.01fF
C53942 PAND2X1_865/Y PAND2X1_78/CTRL2 0.00fF
C53943 PAND2X1_484/O POR2X1_287/B 0.01fF
C53944 POR2X1_662/CTRL2 PAND2X1_55/Y 0.00fF
C53945 POR2X1_389/CTRL POR2X1_537/B 0.02fF
C53946 POR2X1_197/Y POR2X1_198/B 0.33fF
C53947 POR2X1_416/B POR2X1_699/a_56_344# 0.00fF
C53948 POR2X1_85/Y POR2X1_23/Y 0.01fF
C53949 PAND2X1_6/Y POR2X1_540/A 0.03fF
C53950 POR2X1_614/A POR2X1_407/Y 0.03fF
C53951 POR2X1_366/CTRL2 PAND2X1_48/B 0.01fF
C53952 POR2X1_272/Y POR2X1_153/Y 0.03fF
C53953 POR2X1_220/Y POR2X1_260/A 0.13fF
C53954 PAND2X1_847/O POR2X1_48/A 0.08fF
C53955 PAND2X1_508/Y POR2X1_5/Y 0.03fF
C53956 PAND2X1_94/A POR2X1_124/O 0.02fF
C53957 PAND2X1_48/B POR2X1_796/A 0.03fF
C53958 PAND2X1_57/B PAND2X1_701/CTRL2 0.01fF
C53959 PAND2X1_41/B PAND2X1_165/O 0.05fF
C53960 PAND2X1_119/O PAND2X1_96/B 0.04fF
C53961 POR2X1_55/Y PAND2X1_514/CTRL2 0.00fF
C53962 POR2X1_46/Y PAND2X1_514/a_16_344# 0.09fF
C53963 PAND2X1_388/Y PAND2X1_566/Y 0.03fF
C53964 POR2X1_197/a_16_28# POR2X1_260/A 0.03fF
C53965 POR2X1_661/Y POR2X1_711/Y 0.02fF
C53966 PAND2X1_721/B POR2X1_39/B 0.03fF
C53967 POR2X1_319/A POR2X1_863/A 0.03fF
C53968 PAND2X1_96/B POR2X1_532/A 3.80fF
C53969 POR2X1_356/A POR2X1_456/B 0.09fF
C53970 POR2X1_757/A POR2X1_757/a_16_28# 0.03fF
C53971 POR2X1_480/A POR2X1_652/A 0.10fF
C53972 POR2X1_78/A POR2X1_736/A 0.05fF
C53973 POR2X1_404/Y POR2X1_260/A 0.03fF
C53974 PAND2X1_850/Y PAND2X1_390/Y 0.00fF
C53975 PAND2X1_330/a_76_28# POR2X1_385/Y 0.05fF
C53976 POR2X1_213/CTRL POR2X1_568/Y 0.33fF
C53977 POR2X1_332/Y VDD 0.14fF
C53978 PAND2X1_798/B PAND2X1_574/CTRL 0.01fF
C53979 VDD PAND2X1_345/Y 0.29fF
C53980 POR2X1_539/A PAND2X1_6/Y 0.03fF
C53981 PAND2X1_194/CTRL POR2X1_73/Y 0.04fF
C53982 POR2X1_16/A PAND2X1_341/O 0.00fF
C53983 POR2X1_190/Y PAND2X1_189/CTRL 0.01fF
C53984 PAND2X1_585/CTRL2 PAND2X1_56/A 0.01fF
C53985 PAND2X1_863/O PAND2X1_863/A 0.00fF
C53986 POR2X1_447/CTRL POR2X1_510/Y 0.01fF
C53987 VDD POR2X1_726/CTRL 0.00fF
C53988 PAND2X1_580/B POR2X1_767/CTRL 0.00fF
C53989 POR2X1_347/A PAND2X1_23/Y 1.88fF
C53990 PAND2X1_440/O POR2X1_60/A 0.04fF
C53991 PAND2X1_341/B PAND2X1_206/O 0.02fF
C53992 POR2X1_333/Y POR2X1_579/Y 0.03fF
C53993 POR2X1_68/A POR2X1_308/B 0.03fF
C53994 PAND2X1_592/a_76_28# PAND2X1_853/B 0.02fF
C53995 PAND2X1_651/Y PAND2X1_270/a_76_28# 0.07fF
C53996 POR2X1_575/B POR2X1_244/Y 0.01fF
C53997 PAND2X1_47/B PAND2X1_52/B 0.05fF
C53998 PAND2X1_65/B PAND2X1_179/CTRL 0.01fF
C53999 PAND2X1_297/O POR2X1_402/A 0.02fF
C54000 PAND2X1_640/O PAND2X1_633/Y -0.00fF
C54001 D_INPUT_1 POR2X1_101/Y 0.07fF
C54002 POR2X1_387/Y POR2X1_91/Y 0.07fF
C54003 POR2X1_68/B PAND2X1_63/B 0.09fF
C54004 POR2X1_276/A POR2X1_573/A 0.01fF
C54005 POR2X1_102/Y PAND2X1_862/O 0.02fF
C54006 PAND2X1_726/B PAND2X1_546/CTRL 0.03fF
C54007 POR2X1_614/A POR2X1_520/a_16_28# 0.00fF
C54008 POR2X1_312/Y POR2X1_77/Y 0.12fF
C54009 POR2X1_783/CTRL PAND2X1_52/B 0.01fF
C54010 POR2X1_833/O POR2X1_186/B 0.01fF
C54011 POR2X1_717/CTRL POR2X1_101/Y 0.11fF
C54012 PAND2X1_839/B PAND2X1_656/A 0.01fF
C54013 PAND2X1_513/CTRL POR2X1_77/Y 0.03fF
C54014 POR2X1_110/Y POR2X1_372/Y 1.06fF
C54015 PAND2X1_65/B D_INPUT_4 2.04fF
C54016 POR2X1_62/Y POR2X1_294/B 0.01fF
C54017 POR2X1_52/A POR2X1_7/Y 0.02fF
C54018 POR2X1_13/A PAND2X1_346/CTRL2 0.01fF
C54019 POR2X1_62/Y PAND2X1_228/CTRL 0.01fF
C54020 POR2X1_416/B PAND2X1_562/B 0.18fF
C54021 POR2X1_322/Y PAND2X1_569/B 0.29fF
C54022 POR2X1_190/O POR2X1_456/B 0.12fF
C54023 POR2X1_760/Y POR2X1_96/A 0.04fF
C54024 POR2X1_68/A PAND2X1_6/m4_208_n4# 0.07fF
C54025 POR2X1_99/B POR2X1_785/A 0.03fF
C54026 POR2X1_740/Y POR2X1_726/O 0.00fF
C54027 POR2X1_567/A POR2X1_662/Y 0.07fF
C54028 PAND2X1_675/A PAND2X1_730/A 0.03fF
C54029 POR2X1_847/a_16_28# POR2X1_20/B 0.01fF
C54030 PAND2X1_661/CTRL POR2X1_761/A 0.01fF
C54031 PAND2X1_319/a_16_344# POR2X1_416/B 0.02fF
C54032 POR2X1_55/Y PAND2X1_352/B 0.02fF
C54033 POR2X1_96/A POR2X1_304/O 0.01fF
C54034 POR2X1_41/Y POR2X1_42/Y 0.01fF
C54035 POR2X1_265/Y POR2X1_406/A 0.10fF
C54036 POR2X1_740/A POR2X1_319/Y 0.07fF
C54037 POR2X1_730/Y POR2X1_854/B 0.03fF
C54038 POR2X1_78/B POR2X1_147/CTRL2 0.04fF
C54039 POR2X1_332/Y PAND2X1_32/B 0.02fF
C54040 POR2X1_257/A POR2X1_411/B 0.10fF
C54041 POR2X1_43/B PAND2X1_338/CTRL 0.01fF
C54042 PAND2X1_651/CTRL2 POR2X1_588/Y 0.01fF
C54043 POR2X1_456/B POR2X1_569/A 0.15fF
C54044 POR2X1_213/B POR2X1_568/A 0.05fF
C54045 PAND2X1_348/A PAND2X1_348/Y 0.03fF
C54046 POR2X1_416/B POR2X1_13/A 0.34fF
C54047 POR2X1_843/O POR2X1_458/Y 0.01fF
C54048 POR2X1_119/Y POR2X1_816/A 0.05fF
C54049 PAND2X1_206/B POR2X1_37/Y 0.07fF
C54050 PAND2X1_607/CTRL PAND2X1_58/A 0.01fF
C54051 PAND2X1_90/CTRL POR2X1_38/B 0.03fF
C54052 PAND2X1_187/CTRL POR2X1_191/B 0.00fF
C54053 POR2X1_213/B PAND2X1_146/CTRL2 -0.00fF
C54054 POR2X1_361/CTRL2 PAND2X1_48/A 0.00fF
C54055 INPUT_1 PAND2X1_483/CTRL 0.00fF
C54056 PAND2X1_631/O PAND2X1_631/A 0.07fF
C54057 POR2X1_353/A POR2X1_151/O 0.01fF
C54058 POR2X1_407/A PAND2X1_304/a_16_344# 0.02fF
C54059 POR2X1_415/Y POR2X1_39/B 0.01fF
C54060 POR2X1_416/B POR2X1_57/O 0.06fF
C54061 POR2X1_394/A PAND2X1_550/B 0.01fF
C54062 PAND2X1_612/B POR2X1_610/Y 0.03fF
C54063 PAND2X1_20/A PAND2X1_85/CTRL2 0.01fF
C54064 POR2X1_554/B D_INPUT_0 0.03fF
C54065 POR2X1_327/Y POR2X1_539/CTRL2 0.01fF
C54066 PAND2X1_94/A PAND2X1_531/CTRL2 0.01fF
C54067 POR2X1_96/CTRL2 POR2X1_153/Y 0.01fF
C54068 PAND2X1_440/CTRL2 PAND2X1_794/B 0.01fF
C54069 POR2X1_66/B POR2X1_630/B 0.05fF
C54070 PAND2X1_350/CTRL POR2X1_4/Y 0.03fF
C54071 POR2X1_56/Y POR2X1_39/B 0.08fF
C54072 PAND2X1_132/O PAND2X1_52/B 0.03fF
C54073 POR2X1_502/A POR2X1_364/a_16_28# 0.01fF
C54074 POR2X1_178/CTRL2 POR2X1_416/B 0.01fF
C54075 POR2X1_97/CTRL2 POR2X1_97/B 0.01fF
C54076 POR2X1_68/A POR2X1_716/O 0.33fF
C54077 PAND2X1_639/Y POR2X1_7/A 0.04fF
C54078 POR2X1_249/Y PAND2X1_48/A 0.03fF
C54079 PAND2X1_476/A PAND2X1_656/A 0.03fF
C54080 POR2X1_796/Y POR2X1_808/O 0.02fF
C54081 POR2X1_567/A POR2X1_181/B 0.03fF
C54082 PAND2X1_63/B PAND2X1_143/O 0.03fF
C54083 POR2X1_36/CTRL POR2X1_39/B 0.01fF
C54084 POR2X1_814/B PAND2X1_85/CTRL2 0.12fF
C54085 POR2X1_452/A POR2X1_635/Y 0.01fF
C54086 POR2X1_532/A POR2X1_342/B 0.38fF
C54087 PAND2X1_569/B POR2X1_373/O 0.01fF
C54088 PAND2X1_206/A D_INPUT_0 0.00fF
C54089 PAND2X1_242/Y POR2X1_7/B 0.01fF
C54090 PAND2X1_661/B POR2X1_416/B 0.05fF
C54091 POR2X1_416/B PAND2X1_643/Y 0.01fF
C54092 POR2X1_862/A POR2X1_286/CTRL2 0.00fF
C54093 PAND2X1_48/B POR2X1_863/A 0.06fF
C54094 POR2X1_191/Y POR2X1_545/CTRL 0.02fF
C54095 PAND2X1_803/Y POR2X1_39/B 0.02fF
C54096 PAND2X1_485/a_16_344# POR2X1_260/B 0.01fF
C54097 POR2X1_114/B POR2X1_343/B 0.03fF
C54098 PAND2X1_407/CTRL POR2X1_29/A 0.01fF
C54099 POR2X1_270/Y PAND2X1_93/B 0.03fF
C54100 PAND2X1_20/A PAND2X1_9/Y 0.03fF
C54101 POR2X1_234/A POR2X1_42/Y 0.02fF
C54102 POR2X1_814/A POR2X1_362/B 0.11fF
C54103 PAND2X1_606/O POR2X1_37/Y 0.10fF
C54104 POR2X1_66/B POR2X1_20/B 0.03fF
C54105 POR2X1_830/Y PAND2X1_39/B 0.00fF
C54106 POR2X1_502/A POR2X1_846/A 0.03fF
C54107 PAND2X1_827/CTRL POR2X1_294/Y 0.00fF
C54108 PAND2X1_841/B POR2X1_677/Y 0.00fF
C54109 POR2X1_345/O POR2X1_99/B 0.00fF
C54110 PAND2X1_464/B POR2X1_5/Y 0.01fF
C54111 POR2X1_188/Y POR2X1_733/Y 0.00fF
C54112 POR2X1_257/A POR2X1_271/Y 0.08fF
C54113 POR2X1_260/B POR2X1_590/A 7.94fF
C54114 POR2X1_65/A PAND2X1_449/a_56_28# 0.00fF
C54115 POR2X1_109/O POR2X1_32/A 0.00fF
C54116 POR2X1_49/Y POR2X1_411/B 0.10fF
C54117 POR2X1_458/B POR2X1_343/B 0.11fF
C54118 PAND2X1_173/O PAND2X1_72/A 0.19fF
C54119 POR2X1_357/O POR2X1_191/Y 0.26fF
C54120 PAND2X1_48/B POR2X1_9/Y 0.07fF
C54121 PAND2X1_39/B POR2X1_808/A 0.07fF
C54122 PAND2X1_67/CTRL2 POR2X1_330/Y 0.03fF
C54123 POR2X1_105/Y POR2X1_556/A 0.00fF
C54124 PAND2X1_633/Y POR2X1_77/Y 0.01fF
C54125 POR2X1_416/B POR2X1_321/Y 0.02fF
C54126 POR2X1_814/B PAND2X1_9/Y 3.86fF
C54127 PAND2X1_374/a_76_28# POR2X1_39/B 0.02fF
C54128 POR2X1_251/Y POR2X1_250/Y 0.21fF
C54129 PAND2X1_23/Y POR2X1_458/Y 0.22fF
C54130 POR2X1_475/A POR2X1_475/O 0.01fF
C54131 POR2X1_149/O PAND2X1_90/Y 0.02fF
C54132 POR2X1_676/a_16_28# POR2X1_750/B 0.03fF
C54133 POR2X1_257/A POR2X1_376/B 3.31fF
C54134 PAND2X1_666/CTRL PAND2X1_20/A 0.01fF
C54135 POR2X1_558/Y POR2X1_561/B 0.12fF
C54136 POR2X1_20/B PAND2X1_556/B 0.03fF
C54137 POR2X1_648/a_76_344# POR2X1_718/A 0.01fF
C54138 POR2X1_502/A POR2X1_705/B 0.03fF
C54139 POR2X1_760/A PAND2X1_216/a_16_344# 0.02fF
C54140 POR2X1_456/B PAND2X1_72/A 0.10fF
C54141 POR2X1_691/CTRL POR2X1_814/A 0.30fF
C54142 POR2X1_660/Y PAND2X1_58/A 0.03fF
C54143 PAND2X1_217/CTRL INPUT_0 0.01fF
C54144 POR2X1_65/O POR2X1_55/Y 0.02fF
C54145 PAND2X1_274/O POR2X1_411/B 0.03fF
C54146 POR2X1_674/O POR2X1_72/B 0.00fF
C54147 PAND2X1_23/Y PAND2X1_45/O 0.03fF
C54148 PAND2X1_39/B POR2X1_403/A 0.13fF
C54149 POR2X1_99/A POR2X1_66/A 0.02fF
C54150 POR2X1_57/A PAND2X1_635/Y 0.01fF
C54151 POR2X1_856/B POR2X1_856/CTRL 0.05fF
C54152 PAND2X1_20/A PAND2X1_15/O 0.01fF
C54153 PAND2X1_52/CTRL POR2X1_35/Y 0.01fF
C54154 POR2X1_856/B PAND2X1_41/B 0.04fF
C54155 PAND2X1_410/CTRL2 PAND2X1_404/A 0.00fF
C54156 POR2X1_102/Y POR2X1_516/Y 0.03fF
C54157 POR2X1_849/B POR2X1_849/O 0.00fF
C54158 POR2X1_188/A PAND2X1_282/CTRL 0.01fF
C54159 PAND2X1_20/A POR2X1_267/A 0.03fF
C54160 POR2X1_411/B PAND2X1_553/B 0.46fF
C54161 POR2X1_23/Y PAND2X1_712/CTRL2 0.01fF
C54162 POR2X1_707/B PAND2X1_11/Y 0.00fF
C54163 POR2X1_189/Y POR2X1_679/CTRL 0.01fF
C54164 POR2X1_148/a_16_28# POR2X1_213/B 0.08fF
C54165 POR2X1_52/A POR2X1_257/A 0.18fF
C54166 POR2X1_846/CTRL POR2X1_260/A 0.03fF
C54167 POR2X1_669/B PAND2X1_161/a_76_28# 0.04fF
C54168 PAND2X1_654/O PAND2X1_9/Y 0.02fF
C54169 PAND2X1_267/Y INPUT_0 2.77fF
C54170 POR2X1_14/Y POR2X1_40/Y 0.10fF
C54171 PAND2X1_58/A PAND2X1_23/CTRL2 0.01fF
C54172 POR2X1_13/A POR2X1_265/CTRL 0.01fF
C54173 POR2X1_673/a_16_28# POR2X1_296/B 0.03fF
C54174 PAND2X1_453/A POR2X1_40/Y 0.03fF
C54175 POR2X1_814/B PAND2X1_15/O 0.05fF
C54176 POR2X1_230/CTRL POR2X1_32/A 0.01fF
C54177 POR2X1_257/A POR2X1_152/A 0.03fF
C54178 POR2X1_866/A PAND2X1_511/a_76_28# 0.02fF
C54179 D_INPUT_7 POR2X1_1/a_56_344# 0.00fF
C54180 POR2X1_274/CTRL VDD -0.00fF
C54181 POR2X1_105/CTRL2 POR2X1_814/B 0.03fF
C54182 PAND2X1_307/a_76_28# POR2X1_102/Y 0.01fF
C54183 PAND2X1_42/a_16_344# POR2X1_267/A 0.04fF
C54184 PAND2X1_206/B POR2X1_408/Y 0.10fF
C54185 POR2X1_174/B PAND2X1_65/B 0.15fF
C54186 INPUT_3 PAND2X1_6/A 0.24fF
C54187 PAND2X1_48/B POR2X1_274/A 0.03fF
C54188 POR2X1_287/A POR2X1_249/a_16_28# 0.02fF
C54189 PAND2X1_115/Y POR2X1_48/A 0.03fF
C54190 PAND2X1_218/CTRL PAND2X1_267/Y 0.01fF
C54191 GATE_479 POR2X1_72/B 0.03fF
C54192 POR2X1_708/B POR2X1_66/A 0.01fF
C54193 POR2X1_130/A POR2X1_267/CTRL 0.04fF
C54194 PAND2X1_557/A PAND2X1_768/Y 0.00fF
C54195 POR2X1_464/m4_208_n4# POR2X1_186/B 0.21fF
C54196 PAND2X1_209/A PAND2X1_213/CTRL2 0.01fF
C54197 PAND2X1_24/O D_INPUT_1 0.03fF
C54198 POR2X1_624/Y POR2X1_112/Y 0.23fF
C54199 POR2X1_486/CTRL POR2X1_260/A 0.06fF
C54200 POR2X1_76/Y POR2X1_296/B 0.01fF
C54201 POR2X1_123/A POR2X1_633/O 0.01fF
C54202 POR2X1_814/A POR2X1_734/CTRL 0.00fF
C54203 POR2X1_49/Y POR2X1_376/B 0.94fF
C54204 POR2X1_44/CTRL INPUT_7 0.01fF
C54205 POR2X1_49/Y PAND2X1_596/CTRL2 0.01fF
C54206 POR2X1_541/B POR2X1_203/a_56_344# 0.00fF
C54207 POR2X1_646/O POR2X1_590/A 0.03fF
C54208 POR2X1_646/CTRL2 POR2X1_121/B 0.10fF
C54209 POR2X1_643/CTRL POR2X1_294/A 0.01fF
C54210 PAND2X1_22/O PAND2X1_32/B 0.01fF
C54211 POR2X1_847/a_76_344# POR2X1_283/A 0.01fF
C54212 POR2X1_649/B POR2X1_643/Y 0.02fF
C54213 POR2X1_14/Y POR2X1_586/CTRL 0.00fF
C54214 POR2X1_260/B PAND2X1_752/Y 0.02fF
C54215 POR2X1_800/A D_INPUT_0 0.03fF
C54216 PAND2X1_48/B POR2X1_269/A 0.03fF
C54217 POR2X1_646/Y POR2X1_294/B 0.01fF
C54218 POR2X1_23/Y POR2X1_52/Y 0.03fF
C54219 POR2X1_48/A POR2X1_56/Y 0.02fF
C54220 PAND2X1_217/B VDD 3.08fF
C54221 POR2X1_666/Y VDD 0.01fF
C54222 PAND2X1_247/a_16_344# POR2X1_7/A 0.01fF
C54223 POR2X1_20/B POR2X1_235/a_16_28# 0.03fF
C54224 POR2X1_814/B PAND2X1_236/CTRL 0.08fF
C54225 POR2X1_499/CTRL2 POR2X1_576/Y 0.01fF
C54226 PAND2X1_55/Y POR2X1_590/A 2.68fF
C54227 POR2X1_57/A PAND2X1_404/Y 0.02fF
C54228 POR2X1_63/CTRL2 POR2X1_669/B 0.01fF
C54229 POR2X1_296/B POR2X1_740/Y 0.07fF
C54230 POR2X1_60/A POR2X1_7/B 0.16fF
C54231 POR2X1_438/Y POR2X1_73/Y 0.03fF
C54232 POR2X1_220/B POR2X1_782/A 0.05fF
C54233 D_INPUT_0 POR2X1_501/a_16_28# 0.03fF
C54234 POR2X1_422/CTRL2 POR2X1_93/A 0.03fF
C54235 POR2X1_78/A POR2X1_562/O 0.01fF
C54236 PAND2X1_472/B POR2X1_40/Y 0.07fF
C54237 PAND2X1_526/CTRL VDD 0.00fF
C54238 PAND2X1_95/B PAND2X1_47/B 0.04fF
C54239 POR2X1_96/A PAND2X1_390/Y 0.03fF
C54240 PAND2X1_623/a_76_28# POR2X1_615/Y 0.01fF
C54241 PAND2X1_392/B VDD 0.00fF
C54242 POR2X1_48/A POR2X1_258/O 0.11fF
C54243 D_INPUT_0 POR2X1_702/A 0.02fF
C54244 POR2X1_174/A POR2X1_545/A 0.03fF
C54245 PAND2X1_738/Y PAND2X1_562/B 0.10fF
C54246 POR2X1_808/A POR2X1_513/B 0.03fF
C54247 POR2X1_423/Y POR2X1_46/Y 0.05fF
C54248 POR2X1_74/O POR2X1_20/B 0.01fF
C54249 PAND2X1_554/a_16_344# POR2X1_7/B 0.01fF
C54250 POR2X1_687/A PAND2X1_39/B 0.02fF
C54251 POR2X1_333/A POR2X1_853/A 0.03fF
C54252 POR2X1_669/B PAND2X1_642/B 0.01fF
C54253 PAND2X1_222/A POR2X1_385/CTRL2 0.00fF
C54254 POR2X1_498/a_16_28# POR2X1_72/B 0.02fF
C54255 PAND2X1_404/Y POR2X1_229/Y 1.33fF
C54256 POR2X1_54/Y POR2X1_754/CTRL2 0.01fF
C54257 POR2X1_750/B POR2X1_293/Y 0.07fF
C54258 POR2X1_57/a_16_28# PAND2X1_219/A 0.07fF
C54259 PAND2X1_6/Y POR2X1_247/Y 0.03fF
C54260 POR2X1_41/B POR2X1_250/A 1.16fF
C54261 PAND2X1_291/O PAND2X1_93/B 0.15fF
C54262 POR2X1_52/A POR2X1_49/Y 19.11fF
C54263 PAND2X1_269/CTRL2 POR2X1_72/B 0.11fF
C54264 POR2X1_355/B POR2X1_798/O 0.01fF
C54265 POR2X1_66/B POR2X1_264/Y 0.03fF
C54266 POR2X1_40/Y POR2X1_55/Y 0.18fF
C54267 POR2X1_48/A PAND2X1_803/Y 0.03fF
C54268 POR2X1_832/B POR2X1_750/B 0.03fF
C54269 POR2X1_43/B POR2X1_375/Y 0.09fF
C54270 POR2X1_52/A PAND2X1_558/CTRL2 0.00fF
C54271 POR2X1_102/Y PAND2X1_723/CTRL 0.01fF
C54272 PAND2X1_118/a_76_28# POR2X1_78/A 0.01fF
C54273 POR2X1_20/B PAND2X1_358/A 0.07fF
C54274 POR2X1_57/A POR2X1_666/CTRL2 0.03fF
C54275 POR2X1_49/Y POR2X1_152/A 0.07fF
C54276 POR2X1_383/A POR2X1_558/B 0.04fF
C54277 POR2X1_502/A POR2X1_461/B 0.16fF
C54278 PAND2X1_11/Y PAND2X1_26/CTRL2 0.03fF
C54279 POR2X1_65/A PAND2X1_724/B 0.05fF
C54280 POR2X1_828/Y POR2X1_828/O 0.01fF
C54281 PAND2X1_65/B POR2X1_828/CTRL2 0.01fF
C54282 POR2X1_222/Y POR2X1_355/A 0.03fF
C54283 PAND2X1_90/A POR2X1_267/B 0.01fF
C54284 POR2X1_603/Y POR2X1_73/Y 0.07fF
C54285 POR2X1_188/A POR2X1_710/CTRL2 0.01fF
C54286 POR2X1_13/A PAND2X1_512/Y 0.06fF
C54287 POR2X1_860/A POR2X1_572/B 0.02fF
C54288 POR2X1_610/CTRL POR2X1_260/A 0.03fF
C54289 PAND2X1_659/B PAND2X1_735/O 0.00fF
C54290 POR2X1_57/A POR2X1_309/O 0.05fF
C54291 POR2X1_702/B PAND2X1_23/Y 0.01fF
C54292 POR2X1_399/CTRL2 POR2X1_293/Y 0.00fF
C54293 POR2X1_130/A PAND2X1_511/a_16_344# 0.01fF
C54294 PAND2X1_340/CTRL POR2X1_42/Y 0.27fF
C54295 POR2X1_110/Y POR2X1_485/Y 0.01fF
C54296 POR2X1_43/B POR2X1_39/CTRL 0.01fF
C54297 POR2X1_13/A PAND2X1_738/Y 0.05fF
C54298 INPUT_7 POR2X1_587/CTRL2 0.00fF
C54299 PAND2X1_795/B PAND2X1_735/Y 0.07fF
C54300 PAND2X1_56/Y POR2X1_543/A 0.03fF
C54301 POR2X1_734/A POR2X1_391/Y 0.10fF
C54302 PAND2X1_436/CTRL2 POR2X1_129/Y 0.01fF
C54303 PAND2X1_612/B POR2X1_559/A 0.00fF
C54304 POR2X1_166/CTRL2 POR2X1_40/Y 0.01fF
C54305 POR2X1_68/A POR2X1_797/CTRL2 0.03fF
C54306 POR2X1_278/Y PAND2X1_793/Y 0.03fF
C54307 INPUT_0 POR2X1_372/Y 0.06fF
C54308 POR2X1_32/A PAND2X1_550/Y 0.01fF
C54309 POR2X1_682/Y POR2X1_829/A 0.00fF
C54310 POR2X1_817/Y POR2X1_376/B 0.01fF
C54311 POR2X1_68/A POR2X1_402/O 0.02fF
C54312 POR2X1_523/Y POR2X1_849/O 0.01fF
C54313 POR2X1_108/a_16_28# POR2X1_60/A 0.03fF
C54314 POR2X1_376/B PAND2X1_565/CTRL 0.00fF
C54315 POR2X1_132/Y PAND2X1_354/A 0.17fF
C54316 POR2X1_651/CTRL2 PAND2X1_386/Y 0.01fF
C54317 POR2X1_669/B PAND2X1_550/B 0.04fF
C54318 PAND2X1_84/Y PAND2X1_717/CTRL 0.01fF
C54319 POR2X1_634/A PAND2X1_60/B 0.05fF
C54320 PAND2X1_575/A PAND2X1_501/B 0.00fF
C54321 POR2X1_322/O VDD 0.00fF
C54322 POR2X1_844/CTRL POR2X1_94/A 0.16fF
C54323 POR2X1_440/Y POR2X1_174/A 0.02fF
C54324 POR2X1_241/B POR2X1_566/B 0.03fF
C54325 POR2X1_334/B PAND2X1_80/O 0.08fF
C54326 POR2X1_684/CTRL2 POR2X1_7/B 0.03fF
C54327 POR2X1_260/B POR2X1_332/a_16_28# 0.03fF
C54328 PAND2X1_526/CTRL PAND2X1_32/B 0.01fF
C54329 POR2X1_641/a_16_28# POR2X1_318/A 0.06fF
C54330 PAND2X1_265/a_76_28# PAND2X1_60/B 0.02fF
C54331 PAND2X1_580/CTRL2 VDD 0.00fF
C54332 POR2X1_741/Y VDD 1.77fF
C54333 POR2X1_78/A POR2X1_101/Y 0.23fF
C54334 VDD PAND2X1_850/CTRL -0.00fF
C54335 PAND2X1_65/B POR2X1_705/O 0.02fF
C54336 POR2X1_72/B POR2X1_142/Y 1.58fF
C54337 POR2X1_119/Y POR2X1_428/Y 1.97fF
C54338 POR2X1_83/B PAND2X1_569/B 0.07fF
C54339 POR2X1_83/B POR2X1_158/B 0.03fF
C54340 POR2X1_344/O POR2X1_205/A 0.00fF
C54341 POR2X1_346/B PAND2X1_39/CTRL2 0.00fF
C54342 POR2X1_327/CTRL2 POR2X1_572/B 0.01fF
C54343 POR2X1_730/Y PAND2X1_73/Y 0.03fF
C54344 PAND2X1_81/B VDD 0.42fF
C54345 POR2X1_178/CTRL2 PAND2X1_738/Y 0.13fF
C54346 PAND2X1_56/Y POR2X1_332/B 0.03fF
C54347 POR2X1_27/Y PAND2X1_63/B 0.01fF
C54348 PAND2X1_365/O VDD 0.00fF
C54349 PAND2X1_73/O PAND2X1_63/B 0.04fF
C54350 PAND2X1_65/B PAND2X1_59/CTRL 0.01fF
C54351 POR2X1_72/B PAND2X1_175/B 0.08fF
C54352 INPUT_7 D_INPUT_6 0.01fF
C54353 POR2X1_128/CTRL POR2X1_222/Y 0.04fF
C54354 PAND2X1_58/A POR2X1_308/B 0.03fF
C54355 POR2X1_326/A POR2X1_567/B 0.03fF
C54356 PAND2X1_839/CTRL2 POR2X1_293/Y 0.00fF
C54357 PAND2X1_48/B POR2X1_651/O 0.01fF
C54358 POR2X1_855/Y POR2X1_803/A 0.12fF
C54359 POR2X1_16/A PAND2X1_404/CTRL 0.01fF
C54360 POR2X1_179/Y POR2X1_40/Y 0.02fF
C54361 POR2X1_41/B PAND2X1_658/B 0.10fF
C54362 PAND2X1_93/B POR2X1_722/O 0.28fF
C54363 POR2X1_700/Y POR2X1_701/Y 0.02fF
C54364 VDD PAND2X1_32/B 2.24fF
C54365 POR2X1_78/B POR2X1_68/B 0.12fF
C54366 POR2X1_22/A POR2X1_22/a_56_344# 0.00fF
C54367 POR2X1_481/Y PAND2X1_555/A 0.15fF
C54368 POR2X1_343/Y POR2X1_541/B 0.21fF
C54369 POR2X1_78/B PAND2X1_314/O 0.12fF
C54370 PAND2X1_23/Y D_GATE_662 0.01fF
C54371 POR2X1_43/O PAND2X1_838/B 0.01fF
C54372 POR2X1_776/A POR2X1_567/O 0.03fF
C54373 PAND2X1_696/CTRL2 PAND2X1_93/B 0.02fF
C54374 POR2X1_686/B POR2X1_686/CTRL 0.01fF
C54375 PAND2X1_38/CTRL2 POR2X1_68/B 0.03fF
C54376 POR2X1_288/A POR2X1_249/Y 1.72fF
C54377 POR2X1_855/B POR2X1_866/B 0.24fF
C54378 PAND2X1_7/CTRL POR2X1_222/Y 0.00fF
C54379 POR2X1_283/A POR2X1_5/Y 0.16fF
C54380 POR2X1_829/Y PAND2X1_854/A 0.06fF
C54381 PAND2X1_631/CTRL POR2X1_293/Y 0.03fF
C54382 POR2X1_52/CTRL2 PAND2X1_124/Y 0.07fF
C54383 POR2X1_394/A PAND2X1_545/CTRL 0.06fF
C54384 INPUT_0 POR2X1_9/O 0.05fF
C54385 POR2X1_8/Y POR2X1_94/A 0.03fF
C54386 POR2X1_593/B POR2X1_592/A 0.01fF
C54387 POR2X1_101/Y POR2X1_573/CTRL 0.22fF
C54388 POR2X1_503/CTRL POR2X1_65/A 0.01fF
C54389 POR2X1_130/A PAND2X1_60/B 0.20fF
C54390 POR2X1_208/A POR2X1_400/A 0.20fF
C54391 POR2X1_72/B PAND2X1_777/CTRL 0.01fF
C54392 D_INPUT_6 INPUT_4 0.03fF
C54393 POR2X1_420/Y PAND2X1_156/A 0.01fF
C54394 POR2X1_616/Y POR2X1_669/B 0.03fF
C54395 POR2X1_812/B POR2X1_812/O 0.00fF
C54396 POR2X1_808/A POR2X1_598/a_16_28# 0.00fF
C54397 PAND2X1_23/Y POR2X1_462/B 0.05fF
C54398 POR2X1_366/Y POR2X1_804/A 0.03fF
C54399 PAND2X1_319/B POR2X1_46/Y 0.05fF
C54400 POR2X1_804/A POR2X1_294/B 0.07fF
C54401 PAND2X1_23/Y D_INPUT_1 0.02fF
C54402 PAND2X1_787/Y POR2X1_310/Y 0.02fF
C54403 PAND2X1_490/O POR2X1_294/B 0.01fF
C54404 PAND2X1_409/a_16_344# POR2X1_407/Y 0.01fF
C54405 PAND2X1_401/CTRL2 POR2X1_73/Y 0.01fF
C54406 PAND2X1_20/A PAND2X1_692/CTRL 0.01fF
C54407 PAND2X1_552/B PAND2X1_388/CTRL2 0.00fF
C54408 POR2X1_813/Y VDD 0.03fF
C54409 POR2X1_575/B POR2X1_501/B 0.18fF
C54410 PAND2X1_73/Y PAND2X1_323/CTRL 0.01fF
C54411 POR2X1_501/CTRL2 PAND2X1_32/B 0.04fF
C54412 POR2X1_327/Y PAND2X1_299/CTRL2 0.01fF
C54413 PAND2X1_831/O POR2X1_394/A 0.02fF
C54414 POR2X1_294/B POR2X1_535/A 0.08fF
C54415 PAND2X1_795/a_16_344# POR2X1_394/A 0.04fF
C54416 POR2X1_16/A PAND2X1_473/B 0.07fF
C54417 POR2X1_741/Y PAND2X1_32/B 6.23fF
C54418 POR2X1_824/Y POR2X1_293/Y 0.11fF
C54419 PAND2X1_137/Y PAND2X1_349/A 0.00fF
C54420 POR2X1_855/B POR2X1_783/A 0.00fF
C54421 PAND2X1_23/Y POR2X1_724/A 0.07fF
C54422 POR2X1_220/Y POR2X1_725/Y 0.07fF
C54423 PAND2X1_57/B POR2X1_569/A 0.07fF
C54424 POR2X1_532/A PAND2X1_530/O 0.02fF
C54425 POR2X1_8/Y POR2X1_381/O 0.01fF
C54426 POR2X1_538/O PAND2X1_69/A 0.01fF
C54427 POR2X1_383/A PAND2X1_280/O 0.03fF
C54428 PAND2X1_853/O PAND2X1_653/Y 0.09fF
C54429 PAND2X1_55/Y PAND2X1_29/m4_208_n4# 0.07fF
C54430 D_INPUT_3 PAND2X1_8/O 0.02fF
C54431 POR2X1_590/A POR2X1_741/O 0.00fF
C54432 POR2X1_383/A POR2X1_340/CTRL2 0.01fF
C54433 POR2X1_123/O PAND2X1_60/B 0.01fF
C54434 POR2X1_433/Y POR2X1_73/Y 0.01fF
C54435 POR2X1_673/Y VDD 0.82fF
C54436 PAND2X1_6/Y PAND2X1_69/A 1.97fF
C54437 POR2X1_106/Y PAND2X1_853/B 1.54fF
C54438 PAND2X1_556/B PAND2X1_715/B 0.02fF
C54439 POR2X1_559/CTRL POR2X1_38/B 0.06fF
C54440 POR2X1_754/Y POR2X1_39/B 0.23fF
C54441 POR2X1_336/a_16_28# POR2X1_741/Y 0.01fF
C54442 PAND2X1_90/A PAND2X1_63/B 4.44fF
C54443 PAND2X1_632/B POR2X1_252/CTRL 0.01fF
C54444 PAND2X1_556/B PAND2X1_303/Y 0.01fF
C54445 POR2X1_383/A POR2X1_205/CTRL2 0.06fF
C54446 PAND2X1_798/Y POR2X1_83/B 0.10fF
C54447 POR2X1_122/Y PAND2X1_123/Y 0.00fF
C54448 POR2X1_57/A PAND2X1_565/A 0.01fF
C54449 PAND2X1_746/CTRL VDD 0.00fF
C54450 POR2X1_95/O POR2X1_40/Y 0.01fF
C54451 POR2X1_327/Y POR2X1_284/B 0.03fF
C54452 PAND2X1_56/Y POR2X1_574/A 0.16fF
C54453 PAND2X1_840/B PAND2X1_349/A 0.01fF
C54454 POR2X1_406/Y PAND2X1_560/B 0.03fF
C54455 POR2X1_267/B POR2X1_572/Y 0.02fF
C54456 PAND2X1_580/B PAND2X1_853/B 0.03fF
C54457 PAND2X1_56/Y POR2X1_538/A 0.20fF
C54458 POR2X1_416/B POR2X1_29/A 0.05fF
C54459 PAND2X1_96/B POR2X1_758/O 0.03fF
C54460 POR2X1_313/a_76_344# POR2X1_90/Y 0.01fF
C54461 POR2X1_208/Y POR2X1_206/a_16_28# 0.07fF
C54462 POR2X1_387/Y POR2X1_310/CTRL 0.07fF
C54463 PAND2X1_709/O POR2X1_158/B 0.03fF
C54464 POR2X1_198/a_16_28# POR2X1_197/Y 0.03fF
C54465 PAND2X1_23/Y PAND2X1_300/O 0.01fF
C54466 PAND2X1_373/O POR2X1_732/B 0.12fF
C54467 PAND2X1_764/CTRL2 PAND2X1_32/B 0.01fF
C54468 D_INPUT_3 PAND2X1_341/A 0.11fF
C54469 GATE_741 PAND2X1_366/O 0.02fF
C54470 POR2X1_56/Y PAND2X1_840/O 0.03fF
C54471 POR2X1_366/Y PAND2X1_313/O 0.06fF
C54472 POR2X1_73/Y PAND2X1_840/CTRL 0.08fF
C54473 POR2X1_283/A POR2X1_310/O 0.04fF
C54474 PAND2X1_60/B POR2X1_573/A 0.06fF
C54475 POR2X1_333/Y POR2X1_857/B 0.03fF
C54476 PAND2X1_382/O PAND2X1_69/A 0.05fF
C54477 POR2X1_66/B POR2X1_343/Y 0.05fF
C54478 PAND2X1_150/O PAND2X1_60/B 0.01fF
C54479 POR2X1_550/CTRL2 POR2X1_550/Y 0.00fF
C54480 POR2X1_574/a_16_28# POR2X1_574/A 0.06fF
C54481 POR2X1_734/A POR2X1_383/Y 0.07fF
C54482 POR2X1_528/a_16_28# POR2X1_528/Y 0.02fF
C54483 PAND2X1_714/A PAND2X1_326/B 0.00fF
C54484 POR2X1_671/CTRL POR2X1_4/Y 0.00fF
C54485 POR2X1_36/B POR2X1_386/a_16_28# 0.02fF
C54486 POR2X1_695/CTRL POR2X1_425/Y 0.01fF
C54487 PAND2X1_90/Y POR2X1_741/CTRL 0.29fF
C54488 PAND2X1_90/Y PAND2X1_759/O 0.03fF
C54489 POR2X1_114/B POR2X1_260/A 0.00fF
C54490 PAND2X1_751/CTRL2 POR2X1_294/A 0.01fF
C54491 POR2X1_238/Y PAND2X1_308/Y 0.09fF
C54492 POR2X1_265/Y PAND2X1_35/Y 0.03fF
C54493 POR2X1_542/B POR2X1_787/CTRL2 0.03fF
C54494 POR2X1_110/CTRL2 POR2X1_372/Y 0.05fF
C54495 POR2X1_820/Y POR2X1_4/Y 0.03fF
C54496 PAND2X1_467/Y POR2X1_73/Y 0.03fF
C54497 POR2X1_366/A POR2X1_318/A 0.07fF
C54498 POR2X1_739/O POR2X1_568/Y 0.04fF
C54499 INPUT_3 PAND2X1_87/a_56_28# 0.00fF
C54500 POR2X1_529/Y POR2X1_530/Y 0.17fF
C54501 PAND2X1_20/A POR2X1_568/A 0.06fF
C54502 POR2X1_775/A POR2X1_186/B 0.07fF
C54503 POR2X1_845/CTRL2 POR2X1_7/A 0.01fF
C54504 POR2X1_844/B POR2X1_546/O 0.01fF
C54505 POR2X1_616/Y POR2X1_617/CTRL2 0.01fF
C54506 PAND2X1_6/Y PAND2X1_824/B 0.03fF
C54507 PAND2X1_333/CTRL POR2X1_77/Y 0.02fF
C54508 PAND2X1_569/B PAND2X1_168/CTRL2 0.00fF
C54509 POR2X1_571/O POR2X1_844/B 0.01fF
C54510 POR2X1_333/A POR2X1_161/a_16_28# 0.01fF
C54511 POR2X1_477/A POR2X1_552/O 0.01fF
C54512 POR2X1_777/O PAND2X1_48/A 0.05fF
C54513 POR2X1_798/CTRL PAND2X1_52/B 0.00fF
C54514 POR2X1_294/Y POR2X1_837/B 0.04fF
C54515 POR2X1_574/Y POR2X1_513/Y 0.00fF
C54516 PAND2X1_182/B PAND2X1_182/O 0.03fF
C54517 POR2X1_52/A PAND2X1_330/O 0.15fF
C54518 POR2X1_286/Y PAND2X1_52/B 0.01fF
C54519 PAND2X1_850/Y PAND2X1_592/Y 0.02fF
C54520 POR2X1_334/B POR2X1_4/Y 0.10fF
C54521 POR2X1_62/Y POR2X1_56/Y 0.12fF
C54522 PAND2X1_127/O POR2X1_318/A 0.07fF
C54523 POR2X1_383/A POR2X1_362/A 0.01fF
C54524 PAND2X1_23/Y POR2X1_374/CTRL 0.01fF
C54525 POR2X1_814/B POR2X1_568/A 0.07fF
C54526 POR2X1_730/Y PAND2X1_163/O 0.01fF
C54527 PAND2X1_607/m4_208_n4# PAND2X1_609/m4_208_n4# 0.13fF
C54528 POR2X1_677/Y POR2X1_516/Y 0.03fF
C54529 POR2X1_119/Y PAND2X1_469/B 0.00fF
C54530 POR2X1_222/A POR2X1_260/A 0.02fF
C54531 POR2X1_532/A POR2X1_735/CTRL2 0.01fF
C54532 INPUT_5 D_INPUT_4 5.09fF
C54533 POR2X1_442/a_16_28# POR2X1_411/B -0.00fF
C54534 POR2X1_68/B POR2X1_294/A 0.55fF
C54535 PAND2X1_35/Y PAND2X1_327/CTRL 0.01fF
C54536 POR2X1_204/a_16_28# POR2X1_4/Y 0.03fF
C54537 POR2X1_574/Y POR2X1_366/A 0.01fF
C54538 POR2X1_338/CTRL POR2X1_334/Y 0.07fF
C54539 PAND2X1_79/Y POR2X1_571/Y 0.01fF
C54540 PAND2X1_349/A PAND2X1_853/B 0.03fF
C54541 PAND2X1_661/Y POR2X1_394/A 0.07fF
C54542 POR2X1_42/Y POR2X1_39/B 1.20fF
C54543 POR2X1_83/Y PAND2X1_341/A 0.02fF
C54544 PAND2X1_57/B PAND2X1_72/A 2.05fF
C54545 PAND2X1_514/CTRL PAND2X1_348/A 0.02fF
C54546 POR2X1_174/B POR2X1_814/A 0.20fF
C54547 POR2X1_410/a_16_28# PAND2X1_52/B 0.01fF
C54548 POR2X1_610/Y POR2X1_610/CTRL 0.01fF
C54549 POR2X1_83/B POR2X1_667/O 0.16fF
C54550 POR2X1_102/O INPUT_2 0.01fF
C54551 POR2X1_327/Y POR2X1_860/CTRL2 0.01fF
C54552 POR2X1_83/Y POR2X1_91/Y 0.00fF
C54553 PAND2X1_481/CTRL POR2X1_260/A 0.01fF
C54554 PAND2X1_580/a_76_28# PAND2X1_771/Y 0.02fF
C54555 POR2X1_263/Y POR2X1_262/Y 0.00fF
C54556 POR2X1_309/Y POR2X1_39/B 0.01fF
C54557 PAND2X1_658/B POR2X1_77/Y 0.79fF
C54558 POR2X1_60/A PAND2X1_206/B 0.07fF
C54559 PAND2X1_474/CTRL POR2X1_37/Y 0.03fF
C54560 POR2X1_441/CTRL POR2X1_40/Y 0.06fF
C54561 POR2X1_784/A POR2X1_343/B 0.03fF
C54562 POR2X1_394/A POR2X1_394/O 0.07fF
C54563 POR2X1_712/Y PAND2X1_56/A 0.03fF
C54564 PAND2X1_643/O POR2X1_416/B 0.03fF
C54565 POR2X1_707/B PAND2X1_426/O 0.04fF
C54566 PAND2X1_632/O PAND2X1_508/Y 0.03fF
C54567 POR2X1_333/CTRL2 POR2X1_191/Y 0.12fF
C54568 PAND2X1_482/O POR2X1_260/A 0.04fF
C54569 POR2X1_49/Y POR2X1_441/O 0.01fF
C54570 POR2X1_523/Y PAND2X1_52/B 0.03fF
C54571 POR2X1_127/O POR2X1_257/A 0.10fF
C54572 POR2X1_171/O POR2X1_171/Y 0.00fF
C54573 PAND2X1_425/Y POR2X1_121/B 0.00fF
C54574 PAND2X1_631/A PAND2X1_514/CTRL 0.04fF
C54575 PAND2X1_432/a_76_28# POR2X1_648/Y 0.01fF
C54576 POR2X1_339/Y POR2X1_186/B 0.03fF
C54577 POR2X1_649/CTRL2 PAND2X1_52/B 0.01fF
C54578 PAND2X1_69/A PAND2X1_52/B 0.37fF
C54579 POR2X1_260/B POR2X1_66/A 0.26fF
C54580 POR2X1_169/A POR2X1_854/B 0.05fF
C54581 POR2X1_545/O POR2X1_551/A 0.01fF
C54582 PAND2X1_67/O POR2X1_296/B 0.17fF
C54583 POR2X1_825/O POR2X1_20/B 0.02fF
C54584 POR2X1_54/Y POR2X1_83/B 0.14fF
C54585 POR2X1_715/O POR2X1_702/A 0.00fF
C54586 PAND2X1_129/O POR2X1_814/A 0.02fF
C54587 PAND2X1_699/m4_208_n4# POR2X1_750/B 0.08fF
C54588 POR2X1_364/a_16_28# POR2X1_357/Y 0.08fF
C54589 POR2X1_768/Y POR2X1_113/B 0.01fF
C54590 POR2X1_66/B POR2X1_624/Y 0.03fF
C54591 POR2X1_502/A POR2X1_463/CTRL 0.10fF
C54592 POR2X1_568/Y POR2X1_568/O 0.00fF
C54593 POR2X1_48/A POR2X1_754/Y 0.07fF
C54594 POR2X1_234/A PAND2X1_642/B 0.04fF
C54595 PAND2X1_831/Y PAND2X1_332/Y 0.05fF
C54596 POR2X1_102/Y PAND2X1_267/Y 0.01fF
C54597 POR2X1_754/CTRL POR2X1_39/B 0.01fF
C54598 POR2X1_634/CTRL2 POR2X1_260/B 0.03fF
C54599 POR2X1_122/A POR2X1_411/B 0.04fF
C54600 POR2X1_54/Y POR2X1_752/Y 0.07fF
C54601 POR2X1_482/O POR2X1_669/B 0.04fF
C54602 POR2X1_458/Y POR2X1_733/A 0.03fF
C54603 POR2X1_814/A PAND2X1_89/O 0.13fF
C54604 POR2X1_304/O POR2X1_153/Y 0.02fF
C54605 PAND2X1_834/CTRL POR2X1_153/Y 0.06fF
C54606 POR2X1_356/A PAND2X1_52/O 0.04fF
C54607 POR2X1_417/Y PAND2X1_776/Y 0.02fF
C54608 POR2X1_96/A POR2X1_679/CTRL2 0.01fF
C54609 POR2X1_23/Y POR2X1_482/Y 0.02fF
C54610 POR2X1_623/B POR2X1_29/A 0.03fF
C54611 POR2X1_257/A PAND2X1_276/a_16_344# 0.01fF
C54612 PAND2X1_147/CTRL POR2X1_142/Y 0.01fF
C54613 PAND2X1_475/CTRL D_INPUT_0 0.07fF
C54614 POR2X1_269/A POR2X1_269/a_16_28# 0.07fF
C54615 PAND2X1_318/O PAND2X1_464/B 0.06fF
C54616 PAND2X1_736/A POR2X1_250/Y 0.10fF
C54617 PAND2X1_9/Y VDD 1.57fF
C54618 POR2X1_590/A POR2X1_174/A 0.02fF
C54619 POR2X1_263/O PAND2X1_35/Y 0.01fF
C54620 POR2X1_195/A PAND2X1_41/B 0.00fF
C54621 POR2X1_586/Y PAND2X1_58/A 0.05fF
C54622 POR2X1_864/CTRL POR2X1_801/B 0.01fF
C54623 POR2X1_124/CTRL POR2X1_556/A 0.01fF
C54624 POR2X1_20/B POR2X1_625/Y 0.03fF
C54625 POR2X1_46/O POR2X1_409/B 0.01fF
C54626 POR2X1_409/B POR2X1_72/B 0.02fF
C54627 PAND2X1_609/O PAND2X1_90/Y 0.03fF
C54628 POR2X1_69/CTRL POR2X1_29/A 0.00fF
C54629 POR2X1_86/Y PAND2X1_358/A 0.08fF
C54630 POR2X1_456/B POR2X1_579/CTRL 0.01fF
C54631 POR2X1_556/A POR2X1_465/B 0.77fF
C54632 POR2X1_27/Y POR2X1_32/A 0.01fF
C54633 POR2X1_262/Y PAND2X1_215/B 0.01fF
C54634 POR2X1_102/Y PAND2X1_215/O 0.02fF
C54635 PAND2X1_474/CTRL POR2X1_293/Y 0.03fF
C54636 POR2X1_769/CTRL PAND2X1_52/B 0.01fF
C54637 POR2X1_260/m4_208_n4# POR2X1_740/Y 0.06fF
C54638 POR2X1_202/CTRL POR2X1_296/B 0.06fF
C54639 PAND2X1_620/Y POR2X1_496/Y 0.07fF
C54640 PAND2X1_48/B POR2X1_276/B 0.01fF
C54641 POR2X1_567/B POR2X1_480/A 0.10fF
C54642 POR2X1_45/Y POR2X1_150/Y 0.03fF
C54643 PAND2X1_237/CTRL2 VDD -0.00fF
C54644 POR2X1_854/a_16_28# POR2X1_192/Y 0.02fF
C54645 POR2X1_18/O D_INPUT_6 0.05fF
C54646 POR2X1_860/A POR2X1_590/A 0.65fF
C54647 PAND2X1_263/a_16_344# D_INPUT_0 0.02fF
C54648 POR2X1_68/A POR2X1_66/a_16_28# 0.01fF
C54649 POR2X1_23/Y PAND2X1_580/B 0.01fF
C54650 POR2X1_688/CTRL2 PAND2X1_32/B 0.11fF
C54651 POR2X1_814/A PAND2X1_163/CTRL2 0.02fF
C54652 POR2X1_174/B POR2X1_852/B 0.21fF
C54653 POR2X1_446/B POR2X1_193/A 0.03fF
C54654 D_INPUT_2 POR2X1_612/CTRL 0.01fF
C54655 POR2X1_227/B POR2X1_35/Y 0.02fF
C54656 POR2X1_558/B INPUT_0 0.15fF
C54657 POR2X1_260/B PAND2X1_751/O 0.09fF
C54658 PAND2X1_277/CTRL2 POR2X1_546/A 0.03fF
C54659 PAND2X1_717/A POR2X1_387/Y 0.08fF
C54660 PAND2X1_81/B PAND2X1_9/Y 0.09fF
C54661 POR2X1_804/CTRL POR2X1_435/Y 0.08fF
C54662 POR2X1_60/A PAND2X1_220/Y 0.03fF
C54663 PAND2X1_742/O POR2X1_331/Y 0.01fF
C54664 PAND2X1_58/A POR2X1_402/O 0.15fF
C54665 POR2X1_314/a_16_28# POR2X1_257/A 0.03fF
C54666 POR2X1_411/B PAND2X1_570/a_16_344# 0.01fF
C54667 POR2X1_48/A POR2X1_817/A 0.02fF
C54668 PAND2X1_202/O POR2X1_66/A 0.02fF
C54669 PAND2X1_653/Y POR2X1_411/B 0.03fF
C54670 POR2X1_14/Y POR2X1_5/Y 2.29fF
C54671 POR2X1_602/O POR2X1_294/B 0.03fF
C54672 PAND2X1_659/A POR2X1_72/B 0.03fF
C54673 POR2X1_831/O POR2X1_513/Y 0.01fF
C54674 PAND2X1_413/O INPUT_0 0.06fF
C54675 PAND2X1_478/B PAND2X1_803/A 1.31fF
C54676 PAND2X1_9/Y PAND2X1_32/B 0.03fF
C54677 POR2X1_65/A PAND2X1_733/A 0.02fF
C54678 POR2X1_72/Y POR2X1_23/Y 0.08fF
C54679 PAND2X1_750/O POR2X1_816/A 0.02fF
C54680 POR2X1_72/CTRL POR2X1_72/B 0.01fF
C54681 POR2X1_596/A POR2X1_678/CTRL2 0.01fF
C54682 POR2X1_658/CTRL POR2X1_318/A 0.03fF
C54683 PAND2X1_849/CTRL POR2X1_60/Y 0.01fF
C54684 POR2X1_23/Y POR2X1_256/a_16_28# 0.02fF
C54685 POR2X1_260/B POR2X1_222/Y 0.03fF
C54686 PAND2X1_23/Y PAND2X1_93/B 8.82fF
C54687 POR2X1_20/B POR2X1_245/CTRL 0.03fF
C54688 POR2X1_614/A POR2X1_446/B 0.03fF
C54689 POR2X1_105/CTRL2 VDD -0.00fF
C54690 POR2X1_840/B PAND2X1_39/B 0.05fF
C54691 INPUT_2 POR2X1_126/CTRL2 0.01fF
C54692 POR2X1_267/A VDD 0.27fF
C54693 POR2X1_441/Y PAND2X1_551/CTRL2 0.01fF
C54694 POR2X1_48/A POR2X1_42/Y 0.16fF
C54695 PAND2X1_20/A POR2X1_401/O 0.01fF
C54696 PAND2X1_55/Y POR2X1_66/A 1.18fF
C54697 POR2X1_564/Y POR2X1_174/A 11.83fF
C54698 POR2X1_511/Y POR2X1_40/Y 0.01fF
C54699 POR2X1_555/A POR2X1_852/B 0.03fF
C54700 POR2X1_811/B PAND2X1_511/O 0.03fF
C54701 PAND2X1_95/CTRL POR2X1_66/A 0.01fF
C54702 POR2X1_423/Y PAND2X1_787/Y 0.22fF
C54703 POR2X1_524/Y POR2X1_40/Y 0.00fF
C54704 POR2X1_207/A PAND2X1_41/B 0.01fF
C54705 POR2X1_863/A PAND2X1_167/a_16_344# 0.02fF
C54706 POR2X1_808/A VDD 0.23fF
C54707 PAND2X1_90/A PAND2X1_77/CTRL2 0.03fF
C54708 POR2X1_66/B INPUT_4 0.07fF
C54709 POR2X1_149/A POR2X1_149/Y 0.03fF
C54710 POR2X1_260/B POR2X1_532/A 0.58fF
C54711 PAND2X1_23/Y POR2X1_78/A 0.11fF
C54712 POR2X1_566/A POR2X1_750/B 0.08fF
C54713 PAND2X1_463/CTRL2 POR2X1_7/B 0.00fF
C54714 POR2X1_96/A PAND2X1_231/CTRL2 0.03fF
C54715 POR2X1_777/B PAND2X1_372/CTRL 0.14fF
C54716 PAND2X1_59/B PAND2X1_26/O 0.12fF
C54717 POR2X1_750/A POR2X1_7/B 0.04fF
C54718 POR2X1_66/B POR2X1_785/A 0.03fF
C54719 POR2X1_68/A PAND2X1_73/Y 0.06fF
C54720 PAND2X1_669/a_16_344# POR2X1_816/A 0.01fF
C54721 POR2X1_84/B PAND2X1_63/B 0.01fF
C54722 POR2X1_830/Y POR2X1_741/Y 0.08fF
C54723 PAND2X1_412/O PAND2X1_57/B 0.09fF
C54724 POR2X1_472/CTRL POR2X1_862/A 0.06fF
C54725 POR2X1_102/Y POR2X1_757/A 0.01fF
C54726 POR2X1_78/B POR2X1_480/A 0.07fF
C54727 POR2X1_673/Y PAND2X1_9/Y 0.03fF
C54728 PAND2X1_36/CTRL PAND2X1_32/B 0.08fF
C54729 POR2X1_66/B POR2X1_138/O 0.01fF
C54730 POR2X1_472/Y VDD 0.17fF
C54731 POR2X1_306/Y POR2X1_7/B 0.00fF
C54732 POR2X1_416/Y POR2X1_102/Y 0.00fF
C54733 POR2X1_96/A POR2X1_230/CTRL2 0.03fF
C54734 POR2X1_43/B PAND2X1_244/CTRL 0.03fF
C54735 POR2X1_596/A D_INPUT_0 0.03fF
C54736 PAND2X1_9/CTRL2 PAND2X1_6/A 0.00fF
C54737 POR2X1_127/a_16_28# PAND2X1_566/Y 0.08fF
C54738 PAND2X1_456/O PAND2X1_254/Y 0.02fF
C54739 POR2X1_707/B PAND2X1_762/Y 0.03fF
C54740 POR2X1_123/CTRL PAND2X1_41/B 0.01fF
C54741 POR2X1_475/a_16_28# POR2X1_249/Y 0.02fF
C54742 PAND2X1_319/B PAND2X1_352/A 0.10fF
C54743 POR2X1_614/A POR2X1_121/B 0.01fF
C54744 POR2X1_201/CTRL2 POR2X1_35/Y 0.01fF
C54745 POR2X1_290/O POR2X1_290/Y 0.35fF
C54746 POR2X1_188/A PAND2X1_816/O 0.01fF
C54747 POR2X1_590/A POR2X1_447/CTRL2 0.00fF
C54748 POR2X1_188/A PAND2X1_536/CTRL2 0.01fF
C54749 PAND2X1_472/B POR2X1_5/Y 0.41fF
C54750 POR2X1_541/B POR2X1_186/B 0.18fF
C54751 POR2X1_23/Y PAND2X1_349/A 0.03fF
C54752 INPUT_1 PAND2X1_407/O 0.03fF
C54753 PAND2X1_216/B POR2X1_679/Y 0.05fF
C54754 POR2X1_186/Y POR2X1_740/Y 0.13fF
C54755 POR2X1_65/A PAND2X1_454/O 0.01fF
C54756 PAND2X1_736/A PAND2X1_205/Y 0.07fF
C54757 POR2X1_839/a_16_28# POR2X1_836/Y 0.07fF
C54758 POR2X1_102/Y POR2X1_239/O 0.07fF
C54759 POR2X1_852/CTRL POR2X1_776/B 0.03fF
C54760 PAND2X1_20/A POR2X1_840/B 0.05fF
C54761 PAND2X1_573/CTRL PAND2X1_735/Y 0.04fF
C54762 POR2X1_467/Y PAND2X1_69/A 0.03fF
C54763 POR2X1_55/Y POR2X1_5/Y 0.41fF
C54764 POR2X1_66/B PAND2X1_252/O 0.09fF
C54765 POR2X1_653/CTRL2 POR2X1_661/B 0.01fF
C54766 POR2X1_51/A POR2X1_22/CTRL2 0.01fF
C54767 POR2X1_16/A PAND2X1_218/B 0.05fF
C54768 POR2X1_337/A POR2X1_66/A 0.38fF
C54769 POR2X1_680/Y PAND2X1_473/B 0.03fF
C54770 PAND2X1_39/B PAND2X1_399/O 0.02fF
C54771 POR2X1_502/A POR2X1_192/Y 0.05fF
C54772 PAND2X1_407/O POR2X1_153/Y 0.03fF
C54773 PAND2X1_229/O D_GATE_222 0.05fF
C54774 POR2X1_466/A PAND2X1_373/O 0.02fF
C54775 POR2X1_241/B PAND2X1_60/B 0.05fF
C54776 PAND2X1_216/O VDD 0.00fF
C54777 POR2X1_52/A POR2X1_52/a_16_28# 0.03fF
C54778 POR2X1_119/Y POR2X1_262/Y 0.10fF
C54779 POR2X1_78/B PAND2X1_90/A 0.06fF
C54780 PAND2X1_55/Y PAND2X1_13/a_76_28# 0.02fF
C54781 PAND2X1_556/B POR2X1_763/Y 0.03fF
C54782 POR2X1_149/Y VDD 0.18fF
C54783 PAND2X1_661/Y POR2X1_669/B 0.03fF
C54784 PAND2X1_556/B PAND2X1_115/B 0.02fF
C54785 PAND2X1_76/CTRL POR2X1_91/Y 0.10fF
C54786 POR2X1_257/A PAND2X1_716/B 0.10fF
C54787 POR2X1_79/Y PAND2X1_205/B 0.01fF
C54788 POR2X1_719/B PAND2X1_93/B 0.00fF
C54789 POR2X1_719/A PAND2X1_60/B 0.02fF
C54790 POR2X1_94/A POR2X1_68/B 0.30fF
C54791 POR2X1_832/a_16_28# POR2X1_722/Y 0.02fF
C54792 PAND2X1_41/B POR2X1_501/B 0.07fF
C54793 PAND2X1_74/a_76_28# POR2X1_532/A 0.01fF
C54794 POR2X1_43/B POR2X1_421/CTRL2 0.03fF
C54795 POR2X1_807/A POR2X1_804/A 0.05fF
C54796 POR2X1_96/A PAND2X1_592/Y 0.03fF
C54797 PAND2X1_90/A PAND2X1_38/CTRL2 0.03fF
C54798 PAND2X1_827/O POR2X1_507/A 0.05fF
C54799 PAND2X1_293/O PAND2X1_55/Y 0.03fF
C54800 PAND2X1_573/O POR2X1_494/Y 0.00fF
C54801 POR2X1_78/A POR2X1_520/A 0.03fF
C54802 POR2X1_508/CTRL2 POR2X1_192/Y 0.17fF
C54803 POR2X1_814/B POR2X1_840/B 0.05fF
C54804 POR2X1_157/CTRL2 INPUT_5 0.01fF
C54805 PAND2X1_211/CTRL2 PAND2X1_352/Y 0.01fF
C54806 POR2X1_355/B POR2X1_509/a_16_28# 0.02fF
C54807 PAND2X1_717/O VDD -0.00fF
C54808 POR2X1_52/A PAND2X1_440/a_76_28# 0.02fF
C54809 POR2X1_78/B PAND2X1_697/CTRL 0.11fF
C54810 D_INPUT_3 POR2X1_611/CTRL2 0.01fF
C54811 POR2X1_69/O POR2X1_7/A 0.01fF
C54812 POR2X1_754/A POR2X1_615/Y 0.12fF
C54813 PAND2X1_96/B POR2X1_402/O 0.01fF
C54814 POR2X1_817/a_76_344# POR2X1_394/A 0.01fF
C54815 PAND2X1_579/B POR2X1_599/A 0.21fF
C54816 POR2X1_129/CTRL2 POR2X1_129/Y 0.05fF
C54817 POR2X1_606/O POR2X1_294/A 0.03fF
C54818 PAND2X1_541/O POR2X1_91/Y 0.06fF
C54819 POR2X1_809/A PAND2X1_93/B 0.02fF
C54820 POR2X1_119/Y PAND2X1_477/CTRL2 0.00fF
C54821 POR2X1_406/Y PAND2X1_734/CTRL2 0.01fF
C54822 D_INPUT_3 POR2X1_293/O 0.02fF
C54823 POR2X1_474/CTRL2 POR2X1_276/Y 0.01fF
C54824 POR2X1_120/a_76_344# POR2X1_712/Y 0.00fF
C54825 POR2X1_596/A PAND2X1_90/Y 0.28fF
C54826 POR2X1_865/B POR2X1_362/B 0.02fF
C54827 POR2X1_490/Y POR2X1_7/Y 0.00fF
C54828 POR2X1_625/O POR2X1_93/A 0.02fF
C54829 POR2X1_305/Y POR2X1_13/A 0.02fF
C54830 POR2X1_23/Y PAND2X1_708/a_16_344# 0.01fF
C54831 PAND2X1_52/O PAND2X1_72/A 0.04fF
C54832 POR2X1_366/Y POR2X1_317/CTRL2 0.05fF
C54833 PAND2X1_798/B POR2X1_46/Y 0.03fF
C54834 POR2X1_45/Y PAND2X1_364/B 0.07fF
C54835 PAND2X1_137/Y POR2X1_184/Y 0.02fF
C54836 PAND2X1_440/CTRL POR2X1_150/Y 0.01fF
C54837 PAND2X1_852/B VDD 0.17fF
C54838 POR2X1_437/Y PAND2X1_793/Y 0.01fF
C54839 POR2X1_439/CTRL2 POR2X1_456/B 0.11fF
C54840 POR2X1_135/a_16_28# POR2X1_257/A 0.02fF
C54841 POR2X1_776/B POR2X1_350/O 0.08fF
C54842 POR2X1_243/CTRL INPUT_0 0.01fF
C54843 PAND2X1_556/B POR2X1_73/Y 0.03fF
C54844 POR2X1_32/A PAND2X1_853/B 0.03fF
C54845 POR2X1_193/A POR2X1_795/B 0.02fF
C54846 PAND2X1_56/Y POR2X1_579/Y 0.03fF
C54847 POR2X1_43/B POR2X1_275/CTRL 0.01fF
C54848 POR2X1_639/Y VDD 0.30fF
C54849 POR2X1_579/Y POR2X1_795/B 0.03fF
C54850 POR2X1_40/Y PAND2X1_124/O 0.01fF
C54851 POR2X1_96/A PAND2X1_631/O 0.16fF
C54852 PAND2X1_55/Y POR2X1_222/Y 2.23fF
C54853 POR2X1_252/Y POR2X1_48/A 0.01fF
C54854 POR2X1_638/O POR2X1_638/B 0.00fF
C54855 POR2X1_539/O POR2X1_750/B 0.01fF
C54856 POR2X1_66/B POR2X1_537/O 0.01fF
C54857 PAND2X1_857/O POR2X1_23/Y 0.01fF
C54858 PAND2X1_39/B PAND2X1_56/A 0.03fF
C54859 PAND2X1_23/Y POR2X1_510/A 0.03fF
C54860 POR2X1_809/A POR2X1_78/A 0.02fF
C54861 PAND2X1_254/Y POR2X1_73/Y 0.03fF
C54862 PAND2X1_748/O POR2X1_752/Y 0.09fF
C54863 PAND2X1_471/CTRL PAND2X1_241/Y 0.01fF
C54864 POR2X1_397/Y PAND2X1_720/CTRL2 0.11fF
C54865 POR2X1_57/A POR2X1_251/Y 0.01fF
C54866 POR2X1_537/O POR2X1_188/A 0.00fF
C54867 PAND2X1_831/Y POR2X1_13/A 0.00fF
C54868 POR2X1_66/B POR2X1_186/B 0.06fF
C54869 POR2X1_302/Y POR2X1_228/Y 0.00fF
C54870 POR2X1_548/A PAND2X1_8/Y 0.00fF
C54871 POR2X1_83/B POR2X1_701/CTRL2 0.00fF
C54872 PAND2X1_402/B VDD 0.10fF
C54873 PAND2X1_6/Y PAND2X1_183/a_76_28# 0.02fF
C54874 POR2X1_468/CTRL2 POR2X1_478/B 0.00fF
C54875 PAND2X1_575/A POR2X1_816/A 0.03fF
C54876 POR2X1_447/B POR2X1_296/B 0.09fF
C54877 POR2X1_119/Y POR2X1_498/Y 0.01fF
C54878 PAND2X1_390/Y POR2X1_153/Y 0.03fF
C54879 POR2X1_334/B D_INPUT_1 0.10fF
C54880 POR2X1_814/B POR2X1_444/Y 0.39fF
C54881 POR2X1_614/A POR2X1_795/B 0.07fF
C54882 PAND2X1_56/Y POR2X1_614/A 0.06fF
C54883 POR2X1_49/Y PAND2X1_480/O 0.14fF
C54884 POR2X1_532/A POR2X1_205/Y 0.12fF
C54885 POR2X1_96/A PAND2X1_348/Y 0.01fF
C54886 POR2X1_188/A POR2X1_186/B 0.00fF
C54887 POR2X1_41/B POR2X1_387/Y 0.19fF
C54888 POR2X1_769/Y VDD 0.00fF
C54889 PAND2X1_55/Y POR2X1_532/A 0.19fF
C54890 POR2X1_7/B POR2X1_142/Y 0.03fF
C54891 POR2X1_5/Y PAND2X1_508/O 0.08fF
C54892 PAND2X1_6/Y POR2X1_723/B 0.03fF
C54893 POR2X1_3/A PAND2X1_709/CTRL2 -0.00fF
C54894 D_GATE_222 POR2X1_702/A 0.01fF
C54895 POR2X1_717/O POR2X1_717/Y 0.00fF
C54896 POR2X1_687/A VDD 0.22fF
C54897 POR2X1_68/A POR2X1_631/B 0.03fF
C54898 POR2X1_140/B POR2X1_804/A 0.03fF
C54899 POR2X1_481/A PAND2X1_336/CTRL2 0.01fF
C54900 POR2X1_43/B POR2X1_90/Y 0.11fF
C54901 PAND2X1_93/B POR2X1_711/Y 0.07fF
C54902 POR2X1_83/B POR2X1_4/Y 0.06fF
C54903 POR2X1_562/a_16_28# POR2X1_556/Y 0.01fF
C54904 PAND2X1_90/Y POR2X1_703/Y 0.01fF
C54905 PAND2X1_392/B POR2X1_751/Y 0.01fF
C54906 POR2X1_312/O POR2X1_90/Y 0.01fF
C54907 POR2X1_835/CTRL POR2X1_835/B 0.01fF
C54908 PAND2X1_858/CTRL2 PAND2X1_390/Y 0.01fF
C54909 POR2X1_463/Y PAND2X1_700/CTRL 0.00fF
C54910 POR2X1_502/A POR2X1_568/Y 0.05fF
C54911 POR2X1_335/CTRL POR2X1_260/A 0.01fF
C54912 PAND2X1_569/Y PAND2X1_345/a_16_344# 0.02fF
C54913 POR2X1_532/A POR2X1_788/Y 0.02fF
C54914 PAND2X1_659/Y POR2X1_40/Y 0.06fF
C54915 POR2X1_502/A POR2X1_785/B 0.03fF
C54916 POR2X1_618/O POR2X1_7/A 0.02fF
C54917 PAND2X1_730/O PAND2X1_739/B 0.01fF
C54918 POR2X1_480/A PAND2X1_142/CTRL2 0.02fF
C54919 POR2X1_383/A POR2X1_193/A 0.07fF
C54920 POR2X1_383/A POR2X1_579/Y 0.03fF
C54921 PAND2X1_531/CTRL2 POR2X1_549/B 0.04fF
C54922 POR2X1_49/Y PAND2X1_716/B 0.03fF
C54923 PAND2X1_390/O PAND2X1_388/Y 0.00fF
C54924 POR2X1_394/A PAND2X1_719/CTRL2 0.10fF
C54925 D_INPUT_3 PAND2X1_341/a_56_28# 0.00fF
C54926 POR2X1_515/CTRL POR2X1_574/Y 0.01fF
C54927 POR2X1_706/B PAND2X1_48/A 0.01fF
C54928 POR2X1_67/A POR2X1_39/B 0.10fF
C54929 PAND2X1_96/B POR2X1_341/a_16_28# 0.01fF
C54930 PAND2X1_741/B PAND2X1_853/B 9.22fF
C54931 POR2X1_751/Y VDD 0.29fF
C54932 POR2X1_383/A POR2X1_572/B 3.03fF
C54933 POR2X1_8/Y POR2X1_58/m4_208_n4# 0.09fF
C54934 POR2X1_481/A PAND2X1_182/B 0.15fF
C54935 POR2X1_96/Y POR2X1_40/Y 0.03fF
C54936 POR2X1_426/a_16_28# POR2X1_425/Y 0.08fF
C54937 POR2X1_139/A POR2X1_139/a_16_28# 0.04fF
C54938 POR2X1_50/m4_208_n4# POR2X1_744/m4_208_n4# 0.13fF
C54939 PAND2X1_205/Y POR2X1_7/Y 0.00fF
C54940 POR2X1_16/A PAND2X1_793/Y 1.21fF
C54941 POR2X1_639/Y PAND2X1_32/B 0.03fF
C54942 PAND2X1_687/B POR2X1_40/Y 0.02fF
C54943 POR2X1_740/Y POR2X1_702/a_76_344# 0.04fF
C54944 POR2X1_755/a_16_28# POR2X1_665/A 0.05fF
C54945 POR2X1_135/O POR2X1_423/Y 0.01fF
C54946 POR2X1_244/B POR2X1_259/B 0.27fF
C54947 POR2X1_730/Y POR2X1_652/Y 0.05fF
C54948 POR2X1_407/Y POR2X1_532/A 0.06fF
C54949 POR2X1_439/Y POR2X1_188/Y 0.02fF
C54950 POR2X1_661/A PAND2X1_39/B 0.07fF
C54951 POR2X1_78/A POR2X1_711/Y 0.10fF
C54952 POR2X1_219/a_56_344# PAND2X1_88/Y 0.00fF
C54953 POR2X1_564/Y POR2X1_704/Y 0.05fF
C54954 PAND2X1_631/A PAND2X1_513/CTRL2 0.00fF
C54955 PAND2X1_291/CTRL PAND2X1_69/A 0.03fF
C54956 POR2X1_504/Y PAND2X1_631/A 0.00fF
C54957 PAND2X1_794/B PAND2X1_854/A 0.61fF
C54958 PAND2X1_209/A POR2X1_145/Y 0.04fF
C54959 PAND2X1_48/B POR2X1_456/B 0.06fF
C54960 D_GATE_741 POR2X1_566/B 0.10fF
C54961 POR2X1_539/A POR2X1_337/m4_208_n4# 0.01fF
C54962 POR2X1_360/A POR2X1_244/Y 0.04fF
C54963 PAND2X1_825/O POR2X1_402/A 0.02fF
C54964 POR2X1_244/B POR2X1_227/O 0.00fF
C54965 POR2X1_614/A POR2X1_383/A 0.52fF
C54966 POR2X1_371/O POR2X1_372/A 0.01fF
C54967 POR2X1_165/O POR2X1_73/Y 0.01fF
C54968 PAND2X1_35/Y PAND2X1_853/B 0.10fF
C54969 PAND2X1_20/A PAND2X1_56/A 0.05fF
C54970 POR2X1_416/B PAND2X1_556/CTRL 0.01fF
C54971 PAND2X1_41/B POR2X1_738/a_16_28# 0.08fF
C54972 POR2X1_614/A PAND2X1_253/CTRL2 0.03fF
C54973 POR2X1_322/Y PAND2X1_565/a_76_28# 0.01fF
C54974 PAND2X1_800/a_16_344# POR2X1_96/A 0.01fF
C54975 POR2X1_565/B POR2X1_6/O 0.03fF
C54976 PAND2X1_442/a_76_28# POR2X1_192/B 0.04fF
C54977 POR2X1_65/A POR2X1_86/O 0.16fF
C54978 POR2X1_186/O PAND2X1_55/Y 0.16fF
C54979 POR2X1_243/Y POR2X1_294/A 0.07fF
C54980 POR2X1_615/CTRL2 POR2X1_39/B 0.04fF
C54981 POR2X1_383/A POR2X1_38/B 0.07fF
C54982 POR2X1_7/B PAND2X1_156/B 0.01fF
C54983 POR2X1_677/Y POR2X1_271/CTRL 0.00fF
C54984 POR2X1_769/Y PAND2X1_32/B 0.02fF
C54985 POR2X1_537/Y PAND2X1_57/B 0.03fF
C54986 POR2X1_719/CTRL PAND2X1_60/B 0.01fF
C54987 POR2X1_506/B PAND2X1_52/B 0.05fF
C54988 POR2X1_579/Y PAND2X1_171/CTRL2 0.00fF
C54989 POR2X1_92/O POR2X1_408/Y 0.02fF
C54990 POR2X1_567/B PAND2X1_437/CTRL2 0.32fF
C54991 POR2X1_96/A PAND2X1_538/a_56_28# 0.00fF
C54992 POR2X1_192/Y POR2X1_188/Y 0.05fF
C54993 POR2X1_41/a_16_28# POR2X1_42/Y 0.02fF
C54994 PAND2X1_658/A PAND2X1_789/O 0.02fF
C54995 POR2X1_265/Y POR2X1_406/CTRL2 0.01fF
C54996 POR2X1_579/Y PAND2X1_71/Y 0.26fF
C54997 POR2X1_257/A POR2X1_431/CTRL2 0.01fF
C54998 POR2X1_189/Y PAND2X1_853/B 0.03fF
C54999 PAND2X1_290/CTRL PAND2X1_85/Y 0.05fF
C55000 PAND2X1_553/B PAND2X1_716/B 0.01fF
C55001 PAND2X1_549/B POR2X1_239/Y 0.03fF
C55002 POR2X1_814/A PAND2X1_268/O 0.01fF
C55003 POR2X1_772/CTRL PAND2X1_32/B 0.00fF
C55004 POR2X1_814/B PAND2X1_56/A 0.03fF
C55005 POR2X1_57/A POR2X1_164/Y 0.03fF
C55006 POR2X1_659/O POR2X1_186/B 0.01fF
C55007 POR2X1_96/A PAND2X1_476/A 0.03fF
C55008 POR2X1_62/Y POR2X1_42/Y 0.05fF
C55009 PAND2X1_90/A POR2X1_294/A 0.03fF
C55010 POR2X1_43/B PAND2X1_566/a_16_344# 0.02fF
C55011 POR2X1_763/Y POR2X1_320/O 0.04fF
C55012 POR2X1_550/A POR2X1_7/A 0.02fF
C55013 POR2X1_121/A POR2X1_774/A 0.00fF
C55014 POR2X1_184/Y PAND2X1_853/B 0.03fF
C55015 POR2X1_136/O PAND2X1_348/A 0.02fF
C55016 POR2X1_685/A POR2X1_729/Y 0.17fF
C55017 POR2X1_409/Y POR2X1_68/B 0.65fF
C55018 PAND2X1_219/CTRL2 POR2X1_7/Y 0.01fF
C55019 POR2X1_575/O POR2X1_569/A 0.03fF
C55020 PAND2X1_476/A POR2X1_406/CTRL 0.00fF
C55021 POR2X1_661/a_16_28# POR2X1_711/Y 0.08fF
C55022 POR2X1_467/CTRL2 POR2X1_210/A 0.03fF
C55023 PAND2X1_499/Y PAND2X1_840/Y 0.10fF
C55024 POR2X1_383/A POR2X1_440/Y 0.11fF
C55025 PAND2X1_209/A POR2X1_394/A 0.02fF
C55026 POR2X1_703/A POR2X1_228/Y 0.00fF
C55027 POR2X1_20/B POR2X1_411/B 0.22fF
C55028 POR2X1_528/Y POR2X1_158/B 0.02fF
C55029 PAND2X1_587/Y D_INPUT_4 0.03fF
C55030 POR2X1_558/Y PAND2X1_32/B 0.07fF
C55031 PAND2X1_139/Y POR2X1_39/B 0.04fF
C55032 PAND2X1_530/CTRL POR2X1_4/Y 0.03fF
C55033 POR2X1_110/Y POR2X1_43/B 0.15fF
C55034 POR2X1_614/A PAND2X1_71/Y 0.04fF
C55035 POR2X1_415/O POR2X1_39/B 0.01fF
C55036 POR2X1_832/O POR2X1_711/Y 0.03fF
C55037 PAND2X1_291/CTRL PAND2X1_824/B 0.01fF
C55038 POR2X1_178/Y POR2X1_179/Y 0.10fF
C55039 POR2X1_520/m4_208_n4# PAND2X1_518/m4_208_n4# 0.13fF
C55040 POR2X1_175/A POR2X1_863/A 0.03fF
C55041 POR2X1_334/A PAND2X1_88/Y 0.03fF
C55042 POR2X1_57/A POR2X1_122/CTRL 0.01fF
C55043 POR2X1_135/a_16_28# PAND2X1_553/B 0.06fF
C55044 POR2X1_334/B PAND2X1_134/O 0.05fF
C55045 PAND2X1_480/a_16_344# POR2X1_91/Y 0.02fF
C55046 POR2X1_420/O POR2X1_329/A 0.01fF
C55047 POR2X1_38/B PAND2X1_71/Y 0.00fF
C55048 POR2X1_566/A PAND2X1_179/m4_208_n4# 0.06fF
C55049 POR2X1_816/O POR2X1_816/Y 0.02fF
C55050 INPUT_3 PAND2X1_750/O 0.02fF
C55051 POR2X1_856/B POR2X1_466/a_16_28# 0.10fF
C55052 POR2X1_567/B POR2X1_466/m4_208_n4# 0.06fF
C55053 POR2X1_527/O PAND2X1_550/B 0.01fF
C55054 POR2X1_62/Y POR2X1_15/CTRL2 0.01fF
C55055 POR2X1_13/A POR2X1_80/CTRL2 0.00fF
C55056 PAND2X1_700/O PAND2X1_52/B 0.30fF
C55057 POR2X1_529/CTRL2 POR2X1_39/B 0.15fF
C55058 POR2X1_513/B PAND2X1_56/A 1.48fF
C55059 PAND2X1_586/O PAND2X1_60/B 0.02fF
C55060 PAND2X1_631/A POR2X1_136/O 0.03fF
C55061 PAND2X1_388/Y POR2X1_131/A 0.01fF
C55062 PAND2X1_687/a_76_28# PAND2X1_643/Y 0.02fF
C55063 VDD POR2X1_568/A 1.74fF
C55064 POR2X1_440/B POR2X1_174/A 0.04fF
C55065 POR2X1_639/Y PAND2X1_328/a_16_344# 0.02fF
C55066 POR2X1_121/Y PAND2X1_52/B 0.03fF
C55067 POR2X1_62/Y PAND2X1_99/Y 0.03fF
C55068 POR2X1_283/A PAND2X1_502/O 0.05fF
C55069 POR2X1_814/B POR2X1_661/A 0.07fF
C55070 POR2X1_333/O POR2X1_333/Y 0.00fF
C55071 POR2X1_12/A POR2X1_428/Y 0.03fF
C55072 PAND2X1_244/B PAND2X1_358/A 0.72fF
C55073 POR2X1_285/B POR2X1_285/A 0.05fF
C55074 POR2X1_153/Y PAND2X1_123/O 0.08fF
C55075 PAND2X1_70/CTRL POR2X1_451/A 0.01fF
C55076 PAND2X1_339/Y POR2X1_522/CTRL2 0.00fF
C55077 PAND2X1_271/CTRL2 PAND2X1_93/B 0.01fF
C55078 POR2X1_680/a_56_344# POR2X1_594/A 0.00fF
C55079 PAND2X1_52/B PAND2X1_145/CTRL2 0.01fF
C55080 POR2X1_416/B PAND2X1_35/O 0.26fF
C55081 POR2X1_842/CTRL PAND2X1_39/B 0.01fF
C55082 POR2X1_840/CTRL POR2X1_513/A 0.00fF
C55083 POR2X1_35/Y POR2X1_555/O 0.01fF
C55084 POR2X1_309/CTRL POR2X1_150/Y 0.12fF
C55085 PAND2X1_206/B POR2X1_750/A 0.02fF
C55086 PAND2X1_476/A POR2X1_7/A 0.08fF
C55087 PAND2X1_458/O POR2X1_5/Y 0.03fF
C55088 PAND2X1_601/CTRL PAND2X1_93/B 0.01fF
C55089 POR2X1_773/A POR2X1_773/O 0.10fF
C55090 POR2X1_740/Y POR2X1_717/B 0.03fF
C55091 PAND2X1_93/B POR2X1_632/CTRL2 0.00fF
C55092 PAND2X1_407/CTRL2 POR2X1_409/B 0.02fF
C55093 PAND2X1_251/a_76_28# PAND2X1_39/B 0.03fF
C55094 POR2X1_346/B POR2X1_294/A 0.03fF
C55095 POR2X1_327/Y POR2X1_733/Y 0.03fF
C55096 PAND2X1_661/Y PAND2X1_649/A 0.03fF
C55097 POR2X1_54/Y PAND2X1_819/a_76_28# 0.05fF
C55098 POR2X1_711/B INPUT_1 0.01fF
C55099 POR2X1_97/a_16_28# POR2X1_186/B 0.01fF
C55100 PAND2X1_9/Y PAND2X1_15/O 0.03fF
C55101 PAND2X1_796/B POR2X1_32/A 0.01fF
C55102 POR2X1_376/B POR2X1_27/CTRL 0.04fF
C55103 POR2X1_257/A POR2X1_279/O 0.02fF
C55104 PAND2X1_65/B PAND2X1_255/a_76_28# 0.02fF
C55105 POR2X1_711/Y POR2X1_513/CTRL2 0.03fF
C55106 POR2X1_661/A POR2X1_513/B 0.01fF
C55107 POR2X1_711/Y PAND2X1_306/O 0.04fF
C55108 POR2X1_387/Y POR2X1_77/Y 0.07fF
C55109 POR2X1_725/Y POR2X1_513/A 0.03fF
C55110 POR2X1_567/A POR2X1_741/B 0.05fF
C55111 POR2X1_99/B POR2X1_244/Y 0.02fF
C55112 PAND2X1_649/A POR2X1_394/O 0.01fF
C55113 POR2X1_568/A PAND2X1_32/B 0.03fF
C55114 POR2X1_129/CTRL2 POR2X1_37/Y 0.01fF
C55115 PAND2X1_65/B PAND2X1_256/CTRL 0.01fF
C55116 PAND2X1_550/B POR2X1_39/B 0.01fF
C55117 PAND2X1_473/Y POR2X1_329/A 0.01fF
C55118 POR2X1_137/Y PAND2X1_72/A 0.08fF
C55119 POR2X1_60/A PAND2X1_207/CTRL2 0.01fF
C55120 POR2X1_19/O POR2X1_5/Y 0.05fF
C55121 POR2X1_23/Y POR2X1_32/A 0.31fF
C55122 D_INPUT_0 POR2X1_811/A 0.03fF
C55123 POR2X1_333/A PAND2X1_91/O 0.06fF
C55124 POR2X1_814/A PAND2X1_372/CTRL 0.01fF
C55125 PAND2X1_510/B POR2X1_80/CTRL2 0.01fF
C55126 POR2X1_679/A POR2X1_72/B 0.01fF
C55127 POR2X1_376/B POR2X1_20/B 0.37fF
C55128 D_GATE_662 PAND2X1_438/O 0.02fF
C55129 PAND2X1_600/O POR2X1_121/B 0.16fF
C55130 POR2X1_274/A POR2X1_330/Y 0.01fF
C55131 POR2X1_129/O POR2X1_67/A 0.05fF
C55132 PAND2X1_86/a_76_28# INPUT_0 0.02fF
C55133 PAND2X1_175/B POR2X1_173/a_16_28# 0.02fF
C55134 POR2X1_83/B POR2X1_427/CTRL 0.01fF
C55135 POR2X1_686/B POR2X1_864/A 0.00fF
C55136 POR2X1_728/B POR2X1_467/O 0.03fF
C55137 PAND2X1_255/CTRL2 PAND2X1_69/A 0.01fF
C55138 POR2X1_23/Y POR2X1_417/Y 0.07fF
C55139 POR2X1_49/Y POR2X1_490/Y 0.03fF
C55140 POR2X1_29/Y POR2X1_9/Y 2.46fF
C55141 POR2X1_760/A PAND2X1_592/Y 0.03fF
C55142 POR2X1_729/CTRL POR2X1_814/A 0.01fF
C55143 POR2X1_483/CTRL POR2X1_556/A 0.09fF
C55144 PAND2X1_247/O VDD 0.00fF
C55145 PAND2X1_829/O PAND2X1_73/Y 0.02fF
C55146 POR2X1_48/A POR2X1_615/CTRL2 0.07fF
C55147 POR2X1_590/A POR2X1_121/B 0.06fF
C55148 PAND2X1_73/Y PAND2X1_58/A 0.06fF
C55149 POR2X1_37/Y POR2X1_40/Y 0.12fF
C55150 PAND2X1_417/CTRL2 PAND2X1_55/Y 0.03fF
C55151 POR2X1_78/B POR2X1_84/B 0.07fF
C55152 POR2X1_66/B POR2X1_753/Y 0.07fF
C55153 POR2X1_163/CTRL POR2X1_23/Y 0.01fF
C55154 PAND2X1_404/Y POR2X1_236/Y 0.02fF
C55155 POR2X1_83/B PAND2X1_219/A 0.04fF
C55156 POR2X1_66/A PAND2X1_16/CTRL 0.01fF
C55157 POR2X1_52/A POR2X1_20/B 0.13fF
C55158 POR2X1_66/B PAND2X1_39/CTRL 0.01fF
C55159 PAND2X1_221/Y PAND2X1_854/A 0.06fF
C55160 POR2X1_590/A POR2X1_630/A 0.64fF
C55161 POR2X1_49/Y PAND2X1_448/O 0.08fF
C55162 POR2X1_9/Y POR2X1_9/O 0.01fF
C55163 POR2X1_416/B PAND2X1_345/Y 0.07fF
C55164 POR2X1_438/Y PAND2X1_544/CTRL2 0.05fF
C55165 PAND2X1_414/O PAND2X1_6/A 0.04fF
C55166 POR2X1_614/A PAND2X1_426/CTRL 0.01fF
C55167 POR2X1_254/A POR2X1_241/B 0.01fF
C55168 PAND2X1_205/A PAND2X1_204/O 0.00fF
C55169 POR2X1_20/B PAND2X1_398/CTRL2 0.01fF
C55170 POR2X1_68/A PAND2X1_617/a_76_28# 0.02fF
C55171 PAND2X1_657/CTRL2 PAND2X1_217/B 0.01fF
C55172 PAND2X1_317/Y POR2X1_20/B 0.03fF
C55173 POR2X1_334/B POR2X1_137/B 0.76fF
C55174 POR2X1_241/B POR2X1_750/B 0.03fF
C55175 POR2X1_20/B POR2X1_152/A 0.01fF
C55176 PAND2X1_831/CTRL2 POR2X1_102/Y 0.00fF
C55177 POR2X1_102/Y PAND2X1_795/CTRL 0.00fF
C55178 D_INPUT_0 PAND2X1_90/Y 0.07fF
C55179 PAND2X1_52/B PAND2X1_3/B 0.04fF
C55180 PAND2X1_629/O POR2X1_496/Y 0.08fF
C55181 PAND2X1_72/A PAND2X1_18/B 0.06fF
C55182 PAND2X1_94/A POR2X1_643/O 0.01fF
C55183 PAND2X1_404/Y POR2X1_81/Y 0.08fF
C55184 POR2X1_144/Y POR2X1_669/B 0.03fF
C55185 POR2X1_32/A PAND2X1_558/O 0.01fF
C55186 POR2X1_23/Y PAND2X1_35/Y 5.10fF
C55187 PAND2X1_217/B POR2X1_272/CTRL 0.03fF
C55188 POR2X1_441/Y POR2X1_73/Y 0.03fF
C55189 POR2X1_492/CTRL PAND2X1_558/Y 0.04fF
C55190 POR2X1_650/a_16_28# POR2X1_650/A 0.10fF
C55191 POR2X1_800/A POR2X1_808/CTRL 0.00fF
C55192 POR2X1_39/B PAND2X1_840/Y 0.06fF
C55193 PAND2X1_651/Y PAND2X1_796/B 1.16fF
C55194 POR2X1_175/a_56_344# POR2X1_78/A 0.00fF
C55195 POR2X1_863/A POR2X1_337/Y 0.07fF
C55196 POR2X1_416/Y PAND2X1_606/CTRL2 0.01fF
C55197 D_INPUT_0 PAND2X1_351/CTRL2 0.14fF
C55198 POR2X1_670/O POR2X1_40/Y 0.01fF
C55199 POR2X1_78/B POR2X1_400/CTRL2 0.01fF
C55200 POR2X1_837/A POR2X1_507/A 0.03fF
C55201 POR2X1_96/A POR2X1_420/a_16_28# 0.01fF
C55202 POR2X1_753/Y POR2X1_859/A 0.54fF
C55203 POR2X1_453/a_16_28# POR2X1_448/Y -0.00fF
C55204 POR2X1_324/A PAND2X1_41/B 0.03fF
C55205 POR2X1_57/A POR2X1_826/Y 0.04fF
C55206 PAND2X1_271/O POR2X1_804/A 0.12fF
C55207 PAND2X1_576/B PAND2X1_197/Y 1.03fF
C55208 PAND2X1_736/A PAND2X1_806/O 0.00fF
C55209 POR2X1_220/Y POR2X1_296/B 0.07fF
C55210 PAND2X1_42/O PAND2X1_41/B 0.02fF
C55211 POR2X1_409/B POR2X1_277/O 0.01fF
C55212 POR2X1_356/A POR2X1_97/A 0.05fF
C55213 POR2X1_814/B POR2X1_461/O 0.02fF
C55214 PAND2X1_272/CTRL POR2X1_193/A 0.03fF
C55215 POR2X1_65/A PAND2X1_562/B 0.07fF
C55216 INPUT_1 PAND2X1_608/O 0.09fF
C55217 POR2X1_272/CTRL2 POR2X1_272/Y 0.04fF
C55218 POR2X1_241/Y POR2X1_506/B 0.00fF
C55219 POR2X1_368/CTRL2 POR2X1_417/Y 0.08fF
C55220 POR2X1_686/CTRL PAND2X1_39/B 0.04fF
C55221 POR2X1_502/A POR2X1_788/A 0.43fF
C55222 PAND2X1_697/O POR2X1_260/B 0.09fF
C55223 PAND2X1_403/B VDD 0.78fF
C55224 PAND2X1_494/a_16_344# POR2X1_260/B 0.01fF
C55225 POR2X1_453/O VDD 0.00fF
C55226 POR2X1_775/A POR2X1_856/B 0.03fF
C55227 POR2X1_296/B POR2X1_404/Y 0.06fF
C55228 PAND2X1_6/Y PAND2X1_248/O 0.16fF
C55229 POR2X1_411/B PAND2X1_121/CTRL2 0.01fF
C55230 POR2X1_23/Y POR2X1_184/Y 0.10fF
C55231 POR2X1_174/B POR2X1_853/O 0.02fF
C55232 POR2X1_272/CTRL VDD 0.00fF
C55233 POR2X1_222/CTRL2 POR2X1_724/A 0.03fF
C55234 POR2X1_406/Y POR2X1_40/Y 0.01fF
C55235 POR2X1_625/CTRL2 POR2X1_5/Y 0.07fF
C55236 PAND2X1_96/B POR2X1_862/A 0.03fF
C55237 PAND2X1_254/O POR2X1_669/B 0.05fF
C55238 POR2X1_660/Y PAND2X1_55/Y 0.01fF
C55239 POR2X1_155/CTRL POR2X1_750/B 0.01fF
C55240 POR2X1_206/A PAND2X1_41/B 0.21fF
C55241 POR2X1_48/A PAND2X1_642/B 0.08fF
C55242 PAND2X1_651/Y POR2X1_23/Y 0.19fF
C55243 POR2X1_445/A POR2X1_540/a_76_344# -0.01fF
C55244 POR2X1_66/A PAND2X1_385/a_76_28# 0.01fF
C55245 PAND2X1_68/CTRL PAND2X1_6/A 0.03fF
C55246 POR2X1_490/Y PAND2X1_217/CTRL2 0.03fF
C55247 POR2X1_130/A POR2X1_389/Y 0.05fF
C55248 PAND2X1_433/CTRL POR2X1_78/A 0.01fF
C55249 POR2X1_78/A POR2X1_733/A 0.06fF
C55250 POR2X1_511/Y POR2X1_5/Y 0.03fF
C55251 POR2X1_334/B POR2X1_78/A 0.12fF
C55252 PAND2X1_257/CTRL POR2X1_750/B 0.09fF
C55253 POR2X1_23/Y PAND2X1_243/CTRL 0.01fF
C55254 POR2X1_52/A POR2X1_491/CTRL2 0.00fF
C55255 POR2X1_49/Y PAND2X1_661/CTRL2 0.01fF
C55256 POR2X1_341/A POR2X1_553/A 0.03fF
C55257 PAND2X1_56/Y POR2X1_590/A 0.05fF
C55258 POR2X1_348/A POR2X1_243/Y 0.00fF
C55259 POR2X1_590/A POR2X1_732/CTRL 0.00fF
C55260 PAND2X1_620/Y POR2X1_13/A 0.65fF
C55261 POR2X1_23/Y PAND2X1_844/B 0.03fF
C55262 PAND2X1_90/Y POR2X1_793/O 0.05fF
C55263 PAND2X1_57/B PAND2X1_597/CTRL2 0.00fF
C55264 POR2X1_65/A POR2X1_13/A 1.91fF
C55265 POR2X1_40/Y POR2X1_293/Y 0.82fF
C55266 POR2X1_251/Y PAND2X1_140/a_16_344# 0.03fF
C55267 POR2X1_411/B PAND2X1_715/B 0.09fF
C55268 POR2X1_102/Y PAND2X1_339/Y 0.01fF
C55269 POR2X1_96/A PAND2X1_192/CTRL2 0.01fF
C55270 POR2X1_748/A PAND2X1_784/O 0.02fF
C55271 POR2X1_298/Y POR2X1_90/Y 0.00fF
C55272 POR2X1_329/A POR2X1_7/Y 0.03fF
C55273 POR2X1_856/O POR2X1_855/Y 0.02fF
C55274 PAND2X1_90/A POR2X1_94/A 0.37fF
C55275 PAND2X1_209/A POR2X1_669/B 0.03fF
C55276 POR2X1_682/O POR2X1_829/A 0.00fF
C55277 POR2X1_224/Y POR2X1_40/Y 0.01fF
C55278 PAND2X1_23/CTRL2 PAND2X1_55/Y 0.01fF
C55279 POR2X1_124/B POR2X1_78/A 0.02fF
C55280 POR2X1_275/a_56_344# PAND2X1_390/Y 0.00fF
C55281 POR2X1_355/B PAND2X1_65/B 0.10fF
C55282 POR2X1_830/a_16_28# POR2X1_733/A 0.07fF
C55283 POR2X1_83/B POR2X1_816/A 0.03fF
C55284 PAND2X1_349/B POR2X1_42/Y 0.01fF
C55285 POR2X1_37/Y PAND2X1_840/CTRL2 0.01fF
C55286 PAND2X1_96/B PAND2X1_73/Y 0.14fF
C55287 PAND2X1_573/a_16_344# PAND2X1_499/Y 0.09fF
C55288 POR2X1_121/B PAND2X1_583/O 0.05fF
C55289 POR2X1_41/B PAND2X1_596/CTRL 0.01fF
C55290 POR2X1_98/a_16_28# POR2X1_68/B 0.06fF
C55291 POR2X1_411/B PAND2X1_502/CTRL 0.01fF
C55292 POR2X1_777/B PAND2X1_536/CTRL 0.02fF
C55293 PAND2X1_242/O POR2X1_423/Y 0.06fF
C55294 POR2X1_29/A POR2X1_376/A 0.02fF
C55295 PAND2X1_652/A PAND2X1_361/a_76_28# 0.05fF
C55296 POR2X1_614/A POR2X1_634/O 0.09fF
C55297 POR2X1_16/A POR2X1_827/Y 0.02fF
C55298 PAND2X1_621/CTRL2 POR2X1_818/Y 0.01fF
C55299 POR2X1_96/A PAND2X1_739/O 0.04fF
C55300 POR2X1_625/m4_208_n4# POR2X1_754/A 0.01fF
C55301 POR2X1_814/B PAND2X1_411/CTRL2 0.00fF
C55302 PAND2X1_443/Y POR2X1_91/Y 0.04fF
C55303 POR2X1_558/A PAND2X1_73/Y 0.05fF
C55304 POR2X1_37/Y PAND2X1_559/O 0.02fF
C55305 POR2X1_829/CTRL POR2X1_761/Y 0.03fF
C55306 POR2X1_68/A POR2X1_61/Y 0.03fF
C55307 PAND2X1_39/B POR2X1_737/A 0.44fF
C55308 POR2X1_383/A POR2X1_590/A 0.25fF
C55309 PAND2X1_347/Y POR2X1_55/Y 0.00fF
C55310 PAND2X1_52/Y POR2X1_562/B 0.02fF
C55311 POR2X1_368/O POR2X1_372/Y 0.04fF
C55312 PAND2X1_659/B POR2X1_293/Y 0.03fF
C55313 INPUT_1 POR2X1_266/m4_208_n4# 0.12fF
C55314 PAND2X1_798/B PAND2X1_787/Y 0.14fF
C55315 PAND2X1_6/Y POR2X1_828/Y 0.03fF
C55316 PAND2X1_659/O POR2X1_494/Y 0.00fF
C55317 PAND2X1_231/CTRL2 POR2X1_38/Y 0.03fF
C55318 PAND2X1_578/O PAND2X1_577/Y 0.02fF
C55319 POR2X1_119/Y POR2X1_442/O 0.16fF
C55320 PAND2X1_633/Y POR2X1_32/A 0.01fF
C55321 POR2X1_293/Y POR2X1_586/CTRL 0.06fF
C55322 POR2X1_290/Y POR2X1_233/O 0.36fF
C55323 POR2X1_572/B INPUT_0 0.08fF
C55324 POR2X1_750/O POR2X1_750/A 0.02fF
C55325 POR2X1_78/A POR2X1_218/O 0.02fF
C55326 POR2X1_65/A PAND2X1_553/CTRL2 0.01fF
C55327 PAND2X1_724/a_16_344# PAND2X1_731/B 0.01fF
C55328 POR2X1_634/A POR2X1_713/B 0.03fF
C55329 PAND2X1_48/B PAND2X1_57/B 2.72fF
C55330 POR2X1_65/A PAND2X1_643/Y 0.03fF
C55331 PAND2X1_23/Y POR2X1_663/a_16_28# 0.02fF
C55332 POR2X1_241/B POR2X1_502/CTRL2 0.01fF
C55333 POR2X1_287/O POR2X1_249/Y 0.01fF
C55334 POR2X1_557/A POR2X1_296/B 0.00fF
C55335 PAND2X1_96/B POR2X1_573/CTRL2 0.00fF
C55336 POR2X1_289/CTRL VDD 0.00fF
C55337 POR2X1_417/CTRL2 POR2X1_5/Y 0.01fF
C55338 POR2X1_96/A PAND2X1_776/O 0.07fF
C55339 POR2X1_60/Y PAND2X1_338/B 0.16fF
C55340 POR2X1_814/B PAND2X1_177/O 0.12fF
C55341 POR2X1_475/A POR2X1_68/B 0.03fF
C55342 POR2X1_230/CTRL2 POR2X1_38/Y 0.02fF
C55343 PAND2X1_23/Y PAND2X1_371/CTRL2 0.02fF
C55344 POR2X1_43/B INPUT_0 0.26fF
C55345 POR2X1_236/Y PAND2X1_565/A 0.03fF
C55346 POR2X1_492/Y POR2X1_411/B 0.04fF
C55347 POR2X1_555/A PAND2X1_88/Y 0.00fF
C55348 POR2X1_593/B POR2X1_592/CTRL2 0.01fF
C55349 POR2X1_356/A POR2X1_294/B 0.13fF
C55350 POR2X1_356/A POR2X1_366/Y 0.10fF
C55351 PAND2X1_220/Y POR2X1_142/Y 0.03fF
C55352 POR2X1_13/A PAND2X1_190/Y 0.03fF
C55353 POR2X1_343/Y PAND2X1_256/O 0.16fF
C55354 POR2X1_856/B POR2X1_339/Y 0.03fF
C55355 POR2X1_850/CTRL2 POR2X1_850/A 0.01fF
C55356 POR2X1_750/B POR2X1_799/CTRL2 0.01fF
C55357 POR2X1_614/A INPUT_0 0.24fF
C55358 POR2X1_795/CTRL POR2X1_294/B 0.01fF
C55359 PAND2X1_374/CTRL POR2X1_40/Y 0.01fF
C55360 POR2X1_686/A POR2X1_686/a_16_28# 0.03fF
C55361 POR2X1_189/O POR2X1_411/B 0.08fF
C55362 PAND2X1_857/A POR2X1_49/Y 0.03fF
C55363 PAND2X1_558/Y PAND2X1_717/Y 0.23fF
C55364 POR2X1_550/A PAND2X1_525/CTRL2 0.01fF
C55365 POR2X1_66/B PAND2X1_376/CTRL 0.00fF
C55366 PAND2X1_795/B POR2X1_816/A 0.03fF
C55367 POR2X1_840/B VDD 4.81fF
C55368 POR2X1_236/Y POR2X1_395/Y 0.05fF
C55369 POR2X1_66/B PAND2X1_127/CTRL 0.01fF
C55370 POR2X1_616/Y POR2X1_48/A 0.03fF
C55371 POR2X1_96/A PAND2X1_734/CTRL 0.01fF
C55372 POR2X1_38/B INPUT_0 0.08fF
C55373 PAND2X1_615/O VDD 0.00fF
C55374 POR2X1_496/Y PAND2X1_508/Y 0.05fF
C55375 D_GATE_662 POR2X1_477/A 0.07fF
C55376 PAND2X1_734/B PAND2X1_734/O 0.00fF
C55377 POR2X1_650/A POR2X1_493/a_16_28# 0.02fF
C55378 PAND2X1_365/a_16_344# POR2X1_7/B 0.02fF
C55379 PAND2X1_213/Y VDD 0.32fF
C55380 PAND2X1_6/A PAND2X1_375/O 0.15fF
C55381 POR2X1_130/A POR2X1_318/A 1.68fF
C55382 POR2X1_194/B POR2X1_194/a_16_28# 0.02fF
C55383 PAND2X1_467/Y POR2X1_763/A 0.07fF
C55384 INPUT_1 PAND2X1_41/B 0.16fF
C55385 PAND2X1_6/Y PAND2X1_599/CTRL2 0.00fF
C55386 POR2X1_101/A POR2X1_99/A 0.01fF
C55387 PAND2X1_693/a_76_28# PAND2X1_48/B 0.01fF
C55388 POR2X1_305/Y PAND2X1_506/O 0.12fF
C55389 POR2X1_41/B PAND2X1_186/a_16_344# 0.01fF
C55390 PAND2X1_717/a_76_28# PAND2X1_493/Y 0.02fF
C55391 PAND2X1_808/Y PAND2X1_580/O 0.01fF
C55392 PAND2X1_723/Y POR2X1_7/CTRL2 0.00fF
C55393 PAND2X1_675/A PAND2X1_794/B 0.03fF
C55394 POR2X1_68/A POR2X1_35/Y 0.03fF
C55395 POR2X1_41/B D_INPUT_3 0.05fF
C55396 POR2X1_277/CTRL2 POR2X1_278/A 0.00fF
C55397 POR2X1_316/a_16_28# POR2X1_83/B 0.02fF
C55398 POR2X1_400/CTRL2 POR2X1_294/A 0.00fF
C55399 PAND2X1_787/Y PAND2X1_175/a_16_344# 0.06fF
C55400 POR2X1_124/CTRL PAND2X1_60/B 0.01fF
C55401 POR2X1_592/A POR2X1_830/A 0.02fF
C55402 PAND2X1_701/CTRL POR2X1_710/A 0.01fF
C55403 PAND2X1_625/CTRL2 PAND2X1_69/A 0.01fF
C55404 PAND2X1_56/Y POR2X1_574/a_76_344# 0.09fF
C55405 POR2X1_327/Y PAND2X1_279/a_76_28# 0.01fF
C55406 PAND2X1_572/a_76_28# POR2X1_46/Y 0.01fF
C55407 POR2X1_465/B PAND2X1_60/B 0.03fF
C55408 PAND2X1_837/a_76_28# POR2X1_825/Y 0.01fF
C55409 PAND2X1_480/B PAND2X1_717/Y 0.02fF
C55410 PAND2X1_434/CTRL INPUT_0 0.05fF
C55411 POR2X1_557/A POR2X1_547/B 0.09fF
C55412 POR2X1_57/A PAND2X1_736/A 0.07fF
C55413 INPUT_2 POR2X1_416/Y 0.02fF
C55414 PAND2X1_94/A PAND2X1_293/CTRL 0.01fF
C55415 PAND2X1_793/Y PAND2X1_549/B 0.07fF
C55416 PAND2X1_106/CTRL2 PAND2X1_48/B 0.00fF
C55417 POR2X1_130/Y POR2X1_140/O 0.01fF
C55418 PAND2X1_810/O GATE_741 0.02fF
C55419 POR2X1_707/CTRL2 PAND2X1_57/B 0.00fF
C55420 POR2X1_198/B PAND2X1_60/B 0.03fF
C55421 POR2X1_383/A POR2X1_857/B 0.05fF
C55422 POR2X1_725/Y POR2X1_784/A 0.09fF
C55423 PAND2X1_460/a_76_28# POR2X1_7/B 0.02fF
C55424 PAND2X1_104/CTRL POR2X1_4/Y 0.07fF
C55425 POR2X1_258/O PAND2X1_566/Y 0.01fF
C55426 POR2X1_237/O PAND2X1_308/Y 0.01fF
C55427 PAND2X1_718/a_16_344# PAND2X1_645/B 0.02fF
C55428 PAND2X1_718/O POR2X1_591/Y 0.03fF
C55429 POR2X1_335/B POR2X1_68/A 0.19fF
C55430 POR2X1_129/Y POR2X1_5/Y 0.08fF
C55431 POR2X1_527/CTRL POR2X1_96/A 0.00fF
C55432 POR2X1_215/a_16_28# POR2X1_215/A 0.05fF
C55433 PAND2X1_243/B PAND2X1_720/O 0.06fF
C55434 PAND2X1_23/Y POR2X1_325/CTRL 0.01fF
C55435 POR2X1_527/a_16_28# POR2X1_236/Y 0.03fF
C55436 PAND2X1_252/CTRL POR2X1_556/Y 0.01fF
C55437 POR2X1_332/B POR2X1_332/CTRL2 0.01fF
C55438 VDD POR2X1_444/Y 0.22fF
C55439 POR2X1_283/A PAND2X1_724/B 0.03fF
C55440 POR2X1_559/O POR2X1_68/B 0.03fF
C55441 POR2X1_614/Y POR2X1_39/B 0.02fF
C55442 POR2X1_447/B POR2X1_186/Y 0.07fF
C55443 PAND2X1_556/B PAND2X1_348/A 0.01fF
C55444 PAND2X1_108/CTRL2 POR2X1_590/A 0.03fF
C55445 POR2X1_174/B POR2X1_568/B 0.07fF
C55446 POR2X1_96/CTRL2 POR2X1_7/B 0.03fF
C55447 POR2X1_840/B PAND2X1_32/B 0.15fF
C55448 POR2X1_294/B POR2X1_569/A 0.01fF
C55449 PAND2X1_787/A PAND2X1_357/Y 0.05fF
C55450 PAND2X1_686/CTRL2 POR2X1_7/B 0.03fF
C55451 POR2X1_855/B POR2X1_803/A 0.00fF
C55452 PAND2X1_803/Y PAND2X1_566/Y 0.04fF
C55453 POR2X1_725/Y POR2X1_732/B 0.00fF
C55454 PAND2X1_797/Y PAND2X1_169/Y 0.03fF
C55455 POR2X1_599/A PAND2X1_656/A 0.08fF
C55456 POR2X1_48/O PAND2X1_123/Y 0.01fF
C55457 PAND2X1_496/O POR2X1_101/Y 0.25fF
C55458 PAND2X1_658/B PAND2X1_349/A 0.05fF
C55459 PAND2X1_8/Y POR2X1_673/B 0.04fF
C55460 POR2X1_286/O PAND2X1_52/B 0.01fF
C55461 PAND2X1_848/B POR2X1_408/Y 0.05fF
C55462 PAND2X1_575/B POR2X1_184/CTRL 0.01fF
C55463 POR2X1_333/a_76_344# POR2X1_578/Y 0.01fF
C55464 PAND2X1_399/O VDD -0.00fF
C55465 PAND2X1_23/Y PAND2X1_823/CTRL 0.02fF
C55466 POR2X1_210/A VDD 0.25fF
C55467 PAND2X1_55/Y POR2X1_308/B 0.66fF
C55468 POR2X1_97/A PAND2X1_72/A 0.03fF
C55469 POR2X1_316/O POR2X1_13/A 0.01fF
C55470 POR2X1_307/O POR2X1_711/Y 0.04fF
C55471 POR2X1_327/Y POR2X1_217/a_16_28# 0.02fF
C55472 POR2X1_701/O POR2X1_236/Y 0.02fF
C55473 POR2X1_853/A POR2X1_569/Y 0.02fF
C55474 POR2X1_786/Y PAND2X1_63/B 0.08fF
C55475 PAND2X1_95/B PAND2X1_51/O 0.01fF
C55476 PAND2X1_6/Y POR2X1_259/CTRL2 0.00fF
C55477 POR2X1_509/A PAND2X1_503/CTRL 0.00fF
C55478 PAND2X1_295/CTRL2 POR2X1_837/B 0.03fF
C55479 PAND2X1_480/CTRL2 POR2X1_238/Y 0.01fF
C55480 PAND2X1_126/O PAND2X1_69/A 0.03fF
C55481 POR2X1_52/A PAND2X1_502/CTRL 0.01fF
C55482 PAND2X1_303/Y POR2X1_152/A 0.11fF
C55483 PAND2X1_71/CTRL2 PAND2X1_48/A 0.01fF
C55484 POR2X1_836/A PAND2X1_52/B 0.09fF
C55485 PAND2X1_831/O POR2X1_39/B 0.01fF
C55486 POR2X1_56/B PAND2X1_156/A 1.12fF
C55487 POR2X1_68/A PAND2X1_813/O 0.07fF
C55488 PAND2X1_631/A PAND2X1_556/B 0.00fF
C55489 PAND2X1_23/Y POR2X1_227/CTRL 0.04fF
C55490 POR2X1_16/A PAND2X1_723/CTRL -0.01fF
C55491 POR2X1_180/B POR2X1_540/CTRL2 0.00fF
C55492 POR2X1_383/A POR2X1_361/CTRL 0.01fF
C55493 POR2X1_257/A POR2X1_329/A 0.03fF
C55494 POR2X1_72/Y PAND2X1_657/B 0.00fF
C55495 POR2X1_390/B PAND2X1_311/CTRL 0.00fF
C55496 PAND2X1_787/CTRL POR2X1_77/Y 0.01fF
C55497 PAND2X1_6/m4_208_n4# PAND2X1_55/Y 0.07fF
C55498 POR2X1_41/B POR2X1_83/Y 0.02fF
C55499 POR2X1_315/Y PAND2X1_803/Y 0.02fF
C55500 POR2X1_644/A POR2X1_260/A 0.03fF
C55501 PAND2X1_95/B PAND2X1_3/B 0.94fF
C55502 PAND2X1_605/O POR2X1_73/Y 0.05fF
C55503 PAND2X1_631/A PAND2X1_254/Y 1.37fF
C55504 POR2X1_383/A POR2X1_338/O 0.01fF
C55505 PAND2X1_75/O POR2X1_624/Y 0.05fF
C55506 PAND2X1_530/CTRL POR2X1_620/B 0.01fF
C55507 POR2X1_502/A POR2X1_374/O 0.02fF
C55508 POR2X1_544/A POR2X1_568/B 0.44fF
C55509 POR2X1_5/Y PAND2X1_333/Y 0.03fF
C55510 PAND2X1_242/Y POR2X1_423/m4_208_n4# 0.01fF
C55511 PAND2X1_44/a_76_28# PAND2X1_72/A 0.01fF
C55512 POR2X1_650/A PAND2X1_72/A 0.06fF
C55513 POR2X1_289/a_16_28# POR2X1_394/A 0.08fF
C55514 POR2X1_416/B PAND2X1_346/a_76_28# 0.01fF
C55515 PAND2X1_74/O POR2X1_76/B 0.01fF
C55516 POR2X1_574/Y POR2X1_573/A 0.03fF
C55517 POR2X1_503/CTRL POR2X1_283/A 0.03fF
C55518 VDD PAND2X1_56/A 0.51fF
C55519 POR2X1_52/A POR2X1_492/Y 0.02fF
C55520 POR2X1_119/Y PAND2X1_398/O 0.15fF
C55521 POR2X1_416/B VDD 5.83fF
C55522 POR2X1_257/A POR2X1_275/Y 0.04fF
C55523 POR2X1_287/B POR2X1_343/B 0.01fF
C55524 POR2X1_68/B POR2X1_557/B 0.94fF
C55525 PAND2X1_723/CTRL2 POR2X1_7/Y 0.01fF
C55526 POR2X1_41/B PAND2X1_653/O 0.05fF
C55527 POR2X1_863/A POR2X1_436/a_56_344# 0.00fF
C55528 POR2X1_66/B POR2X1_814/O 0.17fF
C55529 POR2X1_643/a_16_28# POR2X1_590/A 0.02fF
C55530 PAND2X1_9/Y PAND2X1_407/CTRL 0.01fF
C55531 POR2X1_169/O POR2X1_566/B 0.02fF
C55532 POR2X1_317/CTRL POR2X1_169/A 0.01fF
C55533 POR2X1_66/Y PAND2X1_39/B 0.56fF
C55534 PAND2X1_714/B POR2X1_73/Y 0.00fF
C55535 PAND2X1_358/A PAND2X1_656/A 0.12fF
C55536 PAND2X1_6/Y PAND2X1_323/a_16_344# 0.01fF
C55537 PAND2X1_831/CTRL2 POR2X1_677/Y 0.00fF
C55538 POR2X1_661/B POR2X1_711/Y 0.16fF
C55539 PAND2X1_745/O POR2X1_568/Y 0.38fF
C55540 POR2X1_76/Y POR2X1_715/CTRL2 0.19fF
C55541 PAND2X1_714/Y PAND2X1_732/A 0.02fF
C55542 POR2X1_648/Y POR2X1_590/A 0.03fF
C55543 POR2X1_57/A POR2X1_7/Y 0.03fF
C55544 PAND2X1_661/Y PAND2X1_120/CTRL 0.11fF
C55545 POR2X1_864/A POR2X1_678/Y 0.03fF
C55546 POR2X1_614/A PAND2X1_143/a_56_28# 0.00fF
C55547 POR2X1_54/Y POR2X1_816/Y 0.03fF
C55548 PAND2X1_476/A POR2X1_38/Y 0.05fF
C55549 POR2X1_371/O POR2X1_387/Y 0.06fF
C55550 PAND2X1_238/CTRL PAND2X1_52/B 0.01fF
C55551 POR2X1_59/CTRL2 POR2X1_394/A 0.01fF
C55552 POR2X1_51/CTRL INPUT_6 0.01fF
C55553 POR2X1_43/B POR2X1_522/CTRL2 0.13fF
C55554 POR2X1_52/A POR2X1_43/Y 0.08fF
C55555 POR2X1_722/B PAND2X1_72/A 0.08fF
C55556 PAND2X1_599/CTRL2 PAND2X1_52/B 0.03fF
C55557 PAND2X1_63/CTRL PAND2X1_9/Y 0.01fF
C55558 POR2X1_73/CTRL2 PAND2X1_341/B 0.01fF
C55559 POR2X1_294/B PAND2X1_72/A 0.17fF
C55560 POR2X1_366/Y PAND2X1_72/A 0.29fF
C55561 POR2X1_39/Y POR2X1_16/Y 0.02fF
C55562 PAND2X1_109/CTRL PAND2X1_32/B 0.01fF
C55563 PAND2X1_6/Y POR2X1_342/Y 0.01fF
C55564 POR2X1_65/O POR2X1_60/A 0.03fF
C55565 POR2X1_853/A PAND2X1_52/B 0.03fF
C55566 POR2X1_817/CTRL PAND2X1_340/B 0.01fF
C55567 POR2X1_14/Y POR2X1_846/Y 0.03fF
C55568 PAND2X1_488/CTRL POR2X1_814/A 0.01fF
C55569 POR2X1_567/A POR2X1_569/A 0.10fF
C55570 POR2X1_296/a_16_28# POR2X1_296/B 0.01fF
C55571 POR2X1_772/CTRL2 POR2X1_113/B 0.01fF
C55572 POR2X1_51/CTRL2 POR2X1_51/B 0.01fF
C55573 POR2X1_250/Y POR2X1_331/Y 0.03fF
C55574 POR2X1_49/Y POR2X1_329/A 0.07fF
C55575 PAND2X1_404/CTRL2 POR2X1_20/B 0.04fF
C55576 PAND2X1_56/A PAND2X1_32/B 0.03fF
C55577 POR2X1_446/B POR2X1_66/A 0.03fF
C55578 POR2X1_391/Y PAND2X1_52/B 0.07fF
C55579 POR2X1_846/A POR2X1_793/CTRL 0.01fF
C55580 POR2X1_847/m4_208_n4# POR2X1_67/A 0.01fF
C55581 POR2X1_55/Y PAND2X1_349/a_16_344# 0.02fF
C55582 POR2X1_416/B PAND2X1_344/CTRL2 0.01fF
C55583 POR2X1_467/O POR2X1_330/Y 0.03fF
C55584 POR2X1_67/Y PAND2X1_526/a_16_344# 0.01fF
C55585 POR2X1_90/Y PAND2X1_326/O 0.07fF
C55586 POR2X1_294/B POR2X1_535/O 0.01fF
C55587 D_INPUT_3 POR2X1_77/Y 0.06fF
C55588 INPUT_1 PAND2X1_476/A 0.02fF
C55589 POR2X1_54/Y PAND2X1_749/a_76_28# 0.05fF
C55590 POR2X1_464/a_16_28# POR2X1_457/Y -0.00fF
C55591 POR2X1_54/Y POR2X1_104/CTRL 0.01fF
C55592 PAND2X1_18/B PAND2X1_2/CTRL2 0.03fF
C55593 POR2X1_16/A PAND2X1_797/Y 0.56fF
C55594 PAND2X1_661/Y POR2X1_39/B 0.03fF
C55595 POR2X1_335/A POR2X1_303/B 0.01fF
C55596 POR2X1_428/Y POR2X1_83/B 0.01fF
C55597 PAND2X1_199/B PAND2X1_123/Y 0.02fF
C55598 POR2X1_586/Y POR2X1_260/B 0.16fF
C55599 POR2X1_48/A POR2X1_482/O 0.02fF
C55600 POR2X1_364/A POR2X1_364/a_16_28# -0.00fF
C55601 PAND2X1_476/A POR2X1_153/Y 0.05fF
C55602 PAND2X1_246/CTRL2 VDD -0.00fF
C55603 PAND2X1_675/a_76_28# POR2X1_250/Y 0.03fF
C55604 POR2X1_302/B PAND2X1_39/B 0.42fF
C55605 POR2X1_203/O PAND2X1_72/A 0.16fF
C55606 PAND2X1_111/B PAND2X1_72/A 0.04fF
C55607 PAND2X1_294/O POR2X1_40/Y 0.17fF
C55608 POR2X1_355/B POR2X1_814/A 0.07fF
C55609 POR2X1_150/Y PAND2X1_736/CTRL 0.01fF
C55610 PAND2X1_469/O PAND2X1_444/Y -0.00fF
C55611 POR2X1_458/Y PAND2X1_369/CTRL 0.02fF
C55612 PAND2X1_809/O POR2X1_7/B 0.01fF
C55613 POR2X1_90/Y POR2X1_91/O 0.17fF
C55614 POR2X1_351/CTRL PAND2X1_72/A 0.00fF
C55615 PAND2X1_93/B PAND2X1_394/O 0.16fF
C55616 POR2X1_257/A PAND2X1_738/CTRL 0.05fF
C55617 POR2X1_681/CTRL POR2X1_829/A 0.00fF
C55618 POR2X1_220/B POR2X1_174/A 0.05fF
C55619 PAND2X1_266/CTRL2 PAND2X1_215/B 0.00fF
C55620 POR2X1_66/A POR2X1_121/B 0.07fF
C55621 POR2X1_647/B POR2X1_286/Y 0.01fF
C55622 POR2X1_661/A PAND2X1_32/B 0.07fF
C55623 PAND2X1_139/B POR2X1_150/Y 0.03fF
C55624 D_INPUT_2 POR2X1_612/A 0.08fF
C55625 POR2X1_814/A POR2X1_730/CTRL2 0.02fF
C55626 POR2X1_604/CTRL2 POR2X1_236/Y 0.10fF
C55627 POR2X1_814/B POR2X1_606/CTRL 0.12fF
C55628 PAND2X1_860/A POR2X1_91/Y 0.03fF
C55629 PAND2X1_206/B PAND2X1_101/CTRL 0.03fF
C55630 POR2X1_552/a_16_28# POR2X1_542/Y -0.00fF
C55631 POR2X1_254/Y POR2X1_556/A 0.07fF
C55632 PAND2X1_535/Y POR2X1_281/Y 0.63fF
C55633 POR2X1_66/A POR2X1_630/A 0.06fF
C55634 POR2X1_290/Y POR2X1_411/A 0.03fF
C55635 POR2X1_23/Y PAND2X1_731/B 0.02fF
C55636 POR2X1_836/a_16_28# POR2X1_836/A 0.06fF
C55637 PAND2X1_93/B POR2X1_593/B 0.01fF
C55638 D_INPUT_0 POR2X1_780/CTRL2 0.00fF
C55639 PAND2X1_862/B POR2X1_20/B 0.02fF
C55640 PAND2X1_55/Y PAND2X1_45/CTRL 0.01fF
C55641 POR2X1_23/Y PAND2X1_579/CTRL 0.01fF
C55642 POR2X1_68/A PAND2X1_52/CTRL2 0.01fF
C55643 POR2X1_55/m4_208_n4# POR2X1_623/m4_208_n4# 0.05fF
C55644 PAND2X1_93/B PAND2X1_387/O 0.05fF
C55645 POR2X1_609/Y PAND2X1_240/CTRL2 0.00fF
C55646 POR2X1_257/A POR2X1_256/O 0.01fF
C55647 PAND2X1_20/A POR2X1_296/Y 0.01fF
C55648 POR2X1_14/Y POR2X1_421/Y 0.00fF
C55649 D_INPUT_5 PAND2X1_57/B 0.02fF
C55650 PAND2X1_427/O POR2X1_121/B 0.09fF
C55651 PAND2X1_231/O D_INPUT_0 0.07fF
C55652 POR2X1_411/B PAND2X1_115/B 0.70fF
C55653 POR2X1_698/O POR2X1_32/A 0.01fF
C55654 POR2X1_109/CTRL VDD -0.00fF
C55655 PAND2X1_65/B POR2X1_476/A 0.06fF
C55656 PAND2X1_657/CTRL POR2X1_72/B 0.01fF
C55657 POR2X1_610/O VDD 0.00fF
C55658 PAND2X1_458/CTRL POR2X1_283/A 0.04fF
C55659 POR2X1_843/CTRL2 POR2X1_287/B 0.01fF
C55660 PAND2X1_58/A PAND2X1_37/m4_208_n4# 0.15fF
C55661 POR2X1_37/Y POR2X1_5/Y 5.75fF
C55662 POR2X1_83/Y POR2X1_85/Y 0.02fF
C55663 POR2X1_78/A POR2X1_593/B 0.03fF
C55664 POR2X1_23/Y POR2X1_256/CTRL2 0.16fF
C55665 PAND2X1_658/A POR2X1_411/B 0.03fF
C55666 POR2X1_60/A POR2X1_40/Y 0.38fF
C55667 PAND2X1_240/CTRL POR2X1_102/Y 0.01fF
C55668 PAND2X1_23/Y POR2X1_294/CTRL 0.01fF
C55669 POR2X1_114/O POR2X1_499/A 0.12fF
C55670 POR2X1_54/Y POR2X1_8/a_16_28# 0.02fF
C55671 PAND2X1_450/CTRL2 POR2X1_257/A 0.03fF
C55672 POR2X1_43/B POR2X1_263/a_16_28# 0.02fF
C55673 POR2X1_639/CTRL POR2X1_750/B 0.01fF
C55674 POR2X1_251/A PAND2X1_540/CTRL2 0.01fF
C55675 PAND2X1_65/B PAND2X1_245/O 0.04fF
C55676 POR2X1_428/Y PAND2X1_709/O 0.04fF
C55677 PAND2X1_58/A POR2X1_61/Y 0.02fF
C55678 POR2X1_76/O POR2X1_740/Y 0.03fF
C55679 PAND2X1_438/CTRL POR2X1_456/B 0.02fF
C55680 POR2X1_567/A PAND2X1_72/A 0.05fF
C55681 POR2X1_307/B POR2X1_296/B 0.20fF
C55682 POR2X1_141/CTRL2 PAND2X1_20/A 0.01fF
C55683 POR2X1_200/CTRL PAND2X1_41/B 0.01fF
C55684 PAND2X1_9/a_56_28# POR2X1_94/A 0.00fF
C55685 POR2X1_341/A PAND2X1_316/O 0.11fF
C55686 POR2X1_32/A POR2X1_372/A 0.46fF
C55687 POR2X1_554/B POR2X1_724/A 0.03fF
C55688 POR2X1_72/B PAND2X1_390/Y 0.05fF
C55689 POR2X1_446/B POR2X1_222/Y 0.04fF
C55690 D_INPUT_0 PAND2X1_735/Y 0.07fF
C55691 PAND2X1_213/a_76_28# PAND2X1_213/A 0.01fF
C55692 POR2X1_467/Y POR2X1_828/Y 0.00fF
C55693 PAND2X1_10/O PAND2X1_8/Y -0.00fF
C55694 PAND2X1_594/a_76_28# PAND2X1_90/Y 0.06fF
C55695 POR2X1_411/B POR2X1_73/Y 0.07fF
C55696 POR2X1_720/A POR2X1_750/A 0.31fF
C55697 POR2X1_60/A PAND2X1_185/a_76_28# 0.02fF
C55698 POR2X1_623/B VDD 0.17fF
C55699 POR2X1_41/B POR2X1_484/CTRL 0.01fF
C55700 PAND2X1_76/Y PAND2X1_575/B 0.01fF
C55701 POR2X1_590/A INPUT_0 0.16fF
C55702 POR2X1_334/B POR2X1_84/A 0.07fF
C55703 POR2X1_78/A POR2X1_733/a_16_28# 0.01fF
C55704 POR2X1_750/B PAND2X1_526/O 0.05fF
C55705 POR2X1_383/Y PAND2X1_52/B 0.03fF
C55706 POR2X1_66/B POR2X1_254/m4_208_n4# 0.15fF
C55707 POR2X1_437/O PAND2X1_190/Y 0.06fF
C55708 POR2X1_647/B POR2X1_649/CTRL2 0.01fF
C55709 POR2X1_504/O POR2X1_846/A 0.18fF
C55710 PAND2X1_30/CTRL PAND2X1_3/B 0.01fF
C55711 PAND2X1_319/B PAND2X1_211/CTRL2 0.02fF
C55712 POR2X1_675/A POR2X1_186/Y 0.02fF
C55713 POR2X1_193/Y PAND2X1_7/Y 0.02fF
C55714 D_INPUT_0 PAND2X1_493/Y 0.03fF
C55715 POR2X1_57/A POR2X1_257/A 0.07fF
C55716 POR2X1_697/Y POR2X1_427/CTRL 0.01fF
C55717 POR2X1_697/CTRL POR2X1_72/B 0.01fF
C55718 PAND2X1_733/CTRL2 PAND2X1_723/Y 0.00fF
C55719 INPUT_3 POR2X1_380/A 0.14fF
C55720 POR2X1_102/Y POR2X1_411/CTRL 0.01fF
C55721 POR2X1_66/B PAND2X1_377/O 0.04fF
C55722 PAND2X1_39/B POR2X1_784/m4_208_n4# 0.12fF
C55723 POR2X1_796/Y POR2X1_828/A 0.03fF
C55724 PAND2X1_653/Y POR2X1_490/Y 0.47fF
C55725 POR2X1_66/A POR2X1_795/B 0.07fF
C55726 PAND2X1_56/Y POR2X1_66/A 0.01fF
C55727 POR2X1_96/A PAND2X1_221/CTRL 0.01fF
C55728 POR2X1_49/Y POR2X1_820/B 0.02fF
C55729 PAND2X1_319/B PAND2X1_212/CTRL2 0.02fF
C55730 PAND2X1_56/Y POR2X1_842/a_76_344# 0.03fF
C55731 POR2X1_783/A POR2X1_783/CTRL 0.01fF
C55732 POR2X1_125/a_16_28# POR2X1_411/B 0.02fF
C55733 POR2X1_448/CTRL POR2X1_294/B 0.08fF
C55734 PAND2X1_575/A POR2X1_498/Y 0.00fF
C55735 POR2X1_78/B POR2X1_661/O 0.08fF
C55736 PAND2X1_220/CTRL2 POR2X1_83/B 0.03fF
C55737 PAND2X1_474/A INPUT_0 0.05fF
C55738 POR2X1_188/A POR2X1_722/Y 0.02fF
C55739 PAND2X1_849/B POR2X1_63/Y 0.05fF
C55740 PAND2X1_465/CTRL POR2X1_7/B 0.00fF
C55741 POR2X1_781/CTRL POR2X1_781/A 0.01fF
C55742 POR2X1_220/Y POR2X1_186/Y 0.12fF
C55743 POR2X1_114/B POR2X1_296/B 0.03fF
C55744 PAND2X1_37/CTRL PAND2X1_6/A 0.01fF
C55745 POR2X1_783/O POR2X1_783/B 0.00fF
C55746 POR2X1_355/B POR2X1_852/B 0.07fF
C55747 POR2X1_474/a_16_28# POR2X1_404/Y 0.06fF
C55748 POR2X1_504/Y POR2X1_96/A 0.00fF
C55749 POR2X1_465/B POR2X1_750/B 0.05fF
C55750 POR2X1_406/Y POR2X1_5/Y 0.01fF
C55751 PAND2X1_675/A POR2X1_83/B 0.03fF
C55752 PAND2X1_279/O POR2X1_740/Y 0.01fF
C55753 PAND2X1_673/CTRL2 POR2X1_13/A 0.01fF
C55754 POR2X1_43/B POR2X1_102/Y 0.15fF
C55755 PAND2X1_798/B PAND2X1_78/CTRL2 0.02fF
C55756 POR2X1_661/CTRL POR2X1_722/Y 0.07fF
C55757 PAND2X1_20/A POR2X1_713/CTRL 0.01fF
C55758 POR2X1_596/A POR2X1_644/B 0.01fF
C55759 POR2X1_541/B POR2X1_244/Y 0.05fF
C55760 POR2X1_78/A POR2X1_562/B 0.03fF
C55761 POR2X1_13/A POR2X1_278/O 0.02fF
C55762 POR2X1_119/Y PAND2X1_266/CTRL2 0.15fF
C55763 PAND2X1_773/B VDD 0.03fF
C55764 POR2X1_131/CTRL2 POR2X1_102/Y 0.01fF
C55765 PAND2X1_180/CTRL2 PAND2X1_182/A 0.00fF
C55766 POR2X1_526/O POR2X1_32/A 0.01fF
C55767 POR2X1_611/CTRL POR2X1_293/Y 0.01fF
C55768 POR2X1_376/B INPUT_4 0.12fF
C55769 PAND2X1_480/O POR2X1_20/B 0.01fF
C55770 PAND2X1_782/a_76_28# POR2X1_747/Y 0.05fF
C55771 POR2X1_483/A PAND2X1_48/O 0.02fF
C55772 POR2X1_346/B PAND2X1_60/CTRL 0.00fF
C55773 POR2X1_66/B PAND2X1_7/a_16_344# 0.01fF
C55774 PAND2X1_204/CTRL POR2X1_79/Y 0.01fF
C55775 POR2X1_329/A PAND2X1_865/A 0.02fF
C55776 PAND2X1_512/Y VDD 0.15fF
C55777 POR2X1_111/Y POR2X1_257/A 0.02fF
C55778 PAND2X1_248/CTRL2 POR2X1_101/Y 0.06fF
C55779 POR2X1_832/CTRL2 POR2X1_722/Y 0.01fF
C55780 POR2X1_52/A INPUT_7 0.01fF
C55781 PAND2X1_654/A PAND2X1_9/Y 0.01fF
C55782 POR2X1_814/B POR2X1_756/CTRL 0.01fF
C55783 PAND2X1_230/CTRL2 PAND2X1_32/B 0.02fF
C55784 POR2X1_43/B PAND2X1_436/A 0.09fF
C55785 POR2X1_806/CTRL POR2X1_804/A 0.11fF
C55786 PAND2X1_738/Y VDD 4.15fF
C55787 PAND2X1_347/Y PAND2X1_568/O 0.05fF
C55788 POR2X1_71/Y PAND2X1_76/Y 0.05fF
C55789 PAND2X1_661/Y POR2X1_48/A 0.03fF
C55790 PAND2X1_279/CTRL PAND2X1_32/B 0.01fF
C55791 POR2X1_866/CTRL2 PAND2X1_32/B 0.01fF
C55792 POR2X1_293/Y POR2X1_5/Y 0.24fF
C55793 POR2X1_102/Y POR2X1_38/B 0.03fF
C55794 POR2X1_383/A POR2X1_66/A 0.21fF
C55795 PAND2X1_217/B POR2X1_273/Y 0.03fF
C55796 PAND2X1_545/a_76_28# PAND2X1_324/Y 0.03fF
C55797 POR2X1_121/B POR2X1_532/A 0.03fF
C55798 PAND2X1_478/B POR2X1_90/Y 0.03fF
C55799 PAND2X1_55/Y POR2X1_402/O 0.01fF
C55800 POR2X1_500/A PAND2X1_316/O 0.00fF
C55801 POR2X1_37/Y POR2X1_235/a_56_344# 0.00fF
C55802 PAND2X1_284/m4_208_n4# POR2X1_279/m4_208_n4# 0.05fF
C55803 POR2X1_16/A PAND2X1_267/Y 0.03fF
C55804 PAND2X1_576/CTRL POR2X1_599/A 0.27fF
C55805 PAND2X1_253/CTRL2 POR2X1_66/A 0.01fF
C55806 POR2X1_335/B PAND2X1_58/A 0.00fF
C55807 PAND2X1_350/A INPUT_0 0.05fF
C55808 POR2X1_20/B PAND2X1_716/B 0.03fF
C55809 PAND2X1_48/B PAND2X1_85/Y 0.07fF
C55810 PAND2X1_658/A POR2X1_376/B 0.03fF
C55811 PAND2X1_702/CTRL2 POR2X1_40/Y 0.03fF
C55812 POR2X1_496/Y POR2X1_283/A 0.00fF
C55813 PAND2X1_272/a_76_28# PAND2X1_60/B 0.01fF
C55814 POR2X1_52/A PAND2X1_579/B 0.03fF
C55815 POR2X1_78/B PAND2X1_144/CTRL2 0.01fF
C55816 PAND2X1_491/CTRL PAND2X1_41/B 0.06fF
C55817 POR2X1_308/O PAND2X1_55/Y 0.18fF
C55818 POR2X1_66/B POR2X1_21/CTRL 0.02fF
C55819 PAND2X1_480/B PAND2X1_151/m4_208_n4# 0.04fF
C55820 POR2X1_750/B POR2X1_685/B 0.01fF
C55821 PAND2X1_635/CTRL2 INPUT_7 0.01fF
C55822 PAND2X1_207/CTRL POR2X1_153/Y 0.04fF
C55823 POR2X1_48/A POR2X1_394/O 0.01fF
C55824 PAND2X1_839/CTRL VDD 0.00fF
C55825 POR2X1_422/m4_208_n4# POR2X1_260/A 0.08fF
C55826 POR2X1_410/CTRL2 POR2X1_790/B 0.03fF
C55827 PAND2X1_653/Y PAND2X1_205/Y 0.54fF
C55828 POR2X1_40/CTRL POR2X1_32/A 0.01fF
C55829 D_INPUT_0 PAND2X1_749/CTRL2 0.00fF
C55830 PAND2X1_793/Y PAND2X1_468/O 0.02fF
C55831 POR2X1_244/B POR2X1_294/B 0.03fF
C55832 POR2X1_578/Y POR2X1_785/O 0.01fF
C55833 PAND2X1_278/O POR2X1_68/B 0.01fF
C55834 PAND2X1_217/B PAND2X1_575/O 0.04fF
C55835 POR2X1_52/A POR2X1_331/A 0.01fF
C55836 PAND2X1_41/B POR2X1_711/CTRL 0.00fF
C55837 POR2X1_119/Y PAND2X1_203/a_56_28# 0.00fF
C55838 POR2X1_57/A POR2X1_49/Y 0.21fF
C55839 PAND2X1_96/B POR2X1_61/Y 7.46fF
C55840 POR2X1_251/O POR2X1_387/Y 0.03fF
C55841 POR2X1_245/Y PAND2X1_784/A 0.15fF
C55842 PAND2X1_206/A PAND2X1_101/B 0.01fF
C55843 POR2X1_52/A POR2X1_763/Y 0.10fF
C55844 POR2X1_376/B POR2X1_73/Y 0.03fF
C55845 PAND2X1_643/Y PAND2X1_729/m4_208_n4# 0.01fF
C55846 POR2X1_273/Y VDD 0.03fF
C55847 PAND2X1_863/B POR2X1_42/Y 0.03fF
C55848 PAND2X1_90/A POR2X1_327/CTRL 0.03fF
C55849 PAND2X1_48/CTRL2 POR2X1_786/Y 0.02fF
C55850 POR2X1_853/A POR2X1_570/O 0.01fF
C55851 D_INPUT_1 PAND2X1_526/m4_208_n4# 0.08fF
C55852 POR2X1_109/a_16_28# POR2X1_394/A 0.10fF
C55853 POR2X1_683/Y INPUT_0 0.06fF
C55854 POR2X1_409/B PAND2X1_560/B 0.03fF
C55855 POR2X1_65/A PAND2X1_113/a_56_28# 0.00fF
C55856 POR2X1_278/Y PAND2X1_339/Y 0.05fF
C55857 POR2X1_307/Y POR2X1_740/Y 0.00fF
C55858 PAND2X1_392/B PAND2X1_383/CTRL2 0.01fF
C55859 POR2X1_652/a_76_344# PAND2X1_90/Y 0.04fF
C55860 PAND2X1_841/O PAND2X1_841/B 0.07fF
C55861 POR2X1_510/B POR2X1_852/B 0.04fF
C55862 POR2X1_220/B PAND2X1_189/O 0.07fF
C55863 PAND2X1_65/B POR2X1_205/A 0.08fF
C55864 PAND2X1_724/B POR2X1_55/Y 0.02fF
C55865 POR2X1_358/a_16_28# POR2X1_578/Y 0.03fF
C55866 POR2X1_504/Y POR2X1_7/A 0.00fF
C55867 POR2X1_654/O POR2X1_725/Y 0.00fF
C55868 POR2X1_763/Y PAND2X1_726/CTRL 0.08fF
C55869 POR2X1_66/A PAND2X1_71/Y 0.00fF
C55870 POR2X1_669/B PAND2X1_200/B 0.02fF
C55871 PAND2X1_635/CTRL2 INPUT_4 0.01fF
C55872 PAND2X1_783/CTRL POR2X1_90/Y 0.12fF
C55873 POR2X1_106/Y POR2X1_387/Y 0.03fF
C55874 PAND2X1_202/CTRL D_INPUT_1 0.06fF
C55875 POR2X1_676/Y PAND2X1_69/A 0.04fF
C55876 POR2X1_72/B PAND2X1_123/O 0.01fF
C55877 PAND2X1_241/a_16_344# POR2X1_238/Y 0.02fF
C55878 POR2X1_408/Y POR2X1_5/Y 2.28fF
C55879 PAND2X1_623/a_16_344# POR2X1_129/Y 0.01fF
C55880 POR2X1_330/Y POR2X1_456/B 0.03fF
C55881 POR2X1_102/Y PAND2X1_532/a_56_28# 0.00fF
C55882 PAND2X1_65/B POR2X1_366/A 0.02fF
C55883 POR2X1_368/Y POR2X1_7/B 0.02fF
C55884 PAND2X1_126/CTRL POR2X1_5/Y 0.09fF
C55885 POR2X1_416/B PAND2X1_9/Y 0.05fF
C55886 POR2X1_66/B POR2X1_244/Y 0.03fF
C55887 PAND2X1_824/B POR2X1_631/CTRL 0.07fF
C55888 POR2X1_131/O PAND2X1_137/Y 0.06fF
C55889 POR2X1_646/Y PAND2X1_48/A 0.03fF
C55890 POR2X1_206/A POR2X1_206/a_16_28# 0.03fF
C55891 PAND2X1_462/B POR2X1_416/Y 0.05fF
C55892 POR2X1_502/A POR2X1_540/A 0.03fF
C55893 POR2X1_65/A POR2X1_744/CTRL2 0.03fF
C55894 POR2X1_32/A PAND2X1_657/B 0.10fF
C55895 POR2X1_62/Y POR2X1_614/Y 0.15fF
C55896 PAND2X1_786/CTRL POR2X1_394/A 0.07fF
C55897 POR2X1_222/Y POR2X1_795/B 0.07fF
C55898 POR2X1_823/Y VDD 0.00fF
C55899 POR2X1_392/a_16_28# POR2X1_391/Y 0.01fF
C55900 PAND2X1_309/CTRL2 POR2X1_335/B 0.01fF
C55901 POR2X1_865/B PAND2X1_372/CTRL 0.03fF
C55902 POR2X1_706/B PAND2X1_94/A 0.03fF
C55903 POR2X1_136/Y VDD 0.16fF
C55904 POR2X1_293/Y POR2X1_310/O 0.08fF
C55905 PAND2X1_553/B PAND2X1_702/CTRL 0.01fF
C55906 POR2X1_52/A POR2X1_73/Y 0.20fF
C55907 POR2X1_559/O PAND2X1_90/A 0.01fF
C55908 PAND2X1_96/B POR2X1_652/Y 0.11fF
C55909 PAND2X1_578/CTRL2 VDD 0.00fF
C55910 PAND2X1_41/B POR2X1_758/Y 0.03fF
C55911 POR2X1_346/B POR2X1_404/a_16_28# 0.00fF
C55912 POR2X1_463/Y POR2X1_710/A 0.10fF
C55913 POR2X1_287/B POR2X1_260/A 0.06fF
C55914 POR2X1_254/Y POR2X1_702/O 0.04fF
C55915 POR2X1_57/A PAND2X1_553/B 0.07fF
C55916 PAND2X1_83/CTRL2 POR2X1_35/Y 0.01fF
C55917 PAND2X1_477/A PAND2X1_803/A 0.00fF
C55918 PAND2X1_592/Y POR2X1_591/Y 0.01fF
C55919 PAND2X1_736/A POR2X1_594/A 0.03fF
C55920 POR2X1_685/A POR2X1_685/a_16_28# 0.05fF
C55921 PAND2X1_461/CTRL D_INPUT_0 0.01fF
C55922 PAND2X1_215/CTRL2 POR2X1_7/Y 0.01fF
C55923 POR2X1_370/Y PAND2X1_368/CTRL2 0.03fF
C55924 PAND2X1_21/CTRL2 POR2X1_260/A 0.01fF
C55925 POR2X1_152/A POR2X1_73/Y 0.03fF
C55926 POR2X1_43/B POR2X1_118/CTRL 0.00fF
C55927 PAND2X1_275/CTRL2 POR2X1_573/A 0.01fF
C55928 PAND2X1_566/Y POR2X1_309/Y 0.03fF
C55929 PAND2X1_94/A PAND2X1_80/CTRL 0.01fF
C55930 PAND2X1_659/Y PAND2X1_200/CTRL 0.00fF
C55931 POR2X1_313/Y POR2X1_177/Y 0.02fF
C55932 POR2X1_539/A POR2X1_502/A 0.03fF
C55933 PAND2X1_804/B POR2X1_283/A 0.00fF
C55934 PAND2X1_6/A POR2X1_255/Y 0.04fF
C55935 POR2X1_104/CTRL POR2X1_4/Y 0.01fF
C55936 POR2X1_483/A POR2X1_260/A 2.80fF
C55937 PAND2X1_63/Y PAND2X1_316/CTRL2 0.04fF
C55938 POR2X1_38/B POR2X1_382/CTRL 0.01fF
C55939 PAND2X1_317/Y POR2X1_258/a_76_344# 0.01fF
C55940 POR2X1_119/Y PAND2X1_404/O 0.15fF
C55941 POR2X1_280/O PAND2X1_552/B 0.16fF
C55942 POR2X1_82/O INPUT_1 0.04fF
C55943 POR2X1_539/A POR2X1_337/CTRL 0.01fF
C55944 PAND2X1_550/B PAND2X1_549/O 0.02fF
C55945 PAND2X1_96/B POR2X1_35/Y 0.03fF
C55946 POR2X1_513/B POR2X1_513/a_16_28# -0.00fF
C55947 PAND2X1_56/Y POR2X1_532/A 0.05fF
C55948 POR2X1_821/Y POR2X1_43/B 0.01fF
C55949 PAND2X1_467/Y POR2X1_96/A 0.03fF
C55950 PAND2X1_495/CTRL2 POR2X1_786/Y 0.01fF
C55951 PAND2X1_8/Y POR2X1_260/A 0.00fF
C55952 POR2X1_679/A POR2X1_173/a_16_28# 0.05fF
C55953 PAND2X1_334/O POR2X1_291/Y -0.00fF
C55954 PAND2X1_385/O PAND2X1_60/B 0.02fF
C55955 POR2X1_590/A POR2X1_510/CTRL 0.01fF
C55956 PAND2X1_756/CTRL POR2X1_394/A 0.03fF
C55957 POR2X1_192/Y POR2X1_192/CTRL 0.01fF
C55958 PAND2X1_41/B PAND2X1_171/a_16_344# 0.01fF
C55959 PAND2X1_62/a_16_344# POR2X1_394/A 0.04fF
C55960 POR2X1_734/A POR2X1_294/A 0.14fF
C55961 POR2X1_316/Y PAND2X1_435/Y 0.06fF
C55962 PAND2X1_390/CTRL2 POR2X1_283/A 0.01fF
C55963 POR2X1_52/A PAND2X1_244/B 0.03fF
C55964 INPUT_7 POR2X1_3/B 0.04fF
C55965 POR2X1_578/Y POR2X1_568/Y 0.00fF
C55966 PAND2X1_403/CTRL POR2X1_20/B 0.07fF
C55967 POR2X1_300/CTRL PAND2X1_349/A 0.01fF
C55968 PAND2X1_691/Y PAND2X1_719/a_76_28# 0.02fF
C55969 PAND2X1_41/B PAND2X1_328/O 0.03fF
C55970 POR2X1_38/Y PAND2X1_734/CTRL 0.01fF
C55971 POR2X1_7/B PAND2X1_155/CTRL 0.01fF
C55972 POR2X1_82/O POR2X1_153/Y -0.00fF
C55973 PAND2X1_661/Y POR2X1_413/A 0.03fF
C55974 POR2X1_119/Y PAND2X1_61/Y 0.05fF
C55975 POR2X1_539/CTRL2 POR2X1_662/Y 0.00fF
C55976 POR2X1_383/A POR2X1_222/Y 0.07fF
C55977 PAND2X1_431/a_16_344# PAND2X1_72/A 0.02fF
C55978 POR2X1_192/Y POR2X1_317/B 0.05fF
C55979 POR2X1_349/O PAND2X1_65/Y 0.02fF
C55980 POR2X1_579/Y POR2X1_332/CTRL2 0.00fF
C55981 POR2X1_458/a_16_28# POR2X1_717/B 0.09fF
C55982 POR2X1_111/Y PAND2X1_553/B 0.02fF
C55983 PAND2X1_23/Y POR2X1_773/B 0.10fF
C55984 PAND2X1_659/Y PAND2X1_723/Y 0.03fF
C55985 POR2X1_737/A VDD 0.21fF
C55986 POR2X1_809/A POR2X1_809/B 0.00fF
C55987 PAND2X1_383/O POR2X1_90/Y 0.07fF
C55988 POR2X1_41/B PAND2X1_114/m4_208_n4# 0.08fF
C55989 POR2X1_359/B PAND2X1_57/B 0.40fF
C55990 PAND2X1_710/CTRL2 PAND2X1_711/A 0.01fF
C55991 POR2X1_13/A PAND2X1_508/Y 0.03fF
C55992 POR2X1_38/Y PAND2X1_194/CTRL 0.01fF
C55993 PAND2X1_727/O POR2X1_152/A 0.01fF
C55994 POR2X1_203/CTRL2 PAND2X1_111/B 0.01fF
C55995 POR2X1_16/A POR2X1_519/Y 0.00fF
C55996 POR2X1_119/Y PAND2X1_404/A 0.01fF
C55997 POR2X1_3/B INPUT_4 0.05fF
C55998 POR2X1_541/CTRL POR2X1_366/A 0.09fF
C55999 POR2X1_133/a_16_28# POR2X1_384/A 0.02fF
C56000 POR2X1_383/A POR2X1_532/A 0.28fF
C56001 POR2X1_390/B PAND2X1_6/Y 0.03fF
C56002 POR2X1_81/CTRL2 POR2X1_494/Y 0.00fF
C56003 PAND2X1_832/CTRL POR2X1_39/B 0.01fF
C56004 PAND2X1_572/O PAND2X1_656/A 0.02fF
C56005 POR2X1_301/O POR2X1_260/A 0.16fF
C56006 POR2X1_814/B POR2X1_716/CTRL2 0.03fF
C56007 POR2X1_705/CTRL2 POR2X1_260/A 0.01fF
C56008 PAND2X1_389/Y PAND2X1_842/Y 0.04fF
C56009 PAND2X1_865/Y INPUT_0 0.03fF
C56010 POR2X1_567/A POR2X1_244/B 0.05fF
C56011 PAND2X1_857/m4_208_n4# PAND2X1_733/m4_208_n4# 0.05fF
C56012 POR2X1_834/Y PAND2X1_433/m4_208_n4# 0.04fF
C56013 POR2X1_45/Y POR2X1_394/A 0.07fF
C56014 POR2X1_845/a_16_28# POR2X1_532/A 0.02fF
C56015 PAND2X1_349/A POR2X1_387/Y 0.03fF
C56016 POR2X1_345/CTRL PAND2X1_6/Y 0.01fF
C56017 POR2X1_722/B POR2X1_722/CTRL 0.01fF
C56018 PAND2X1_59/CTRL2 POR2X1_260/A 0.01fF
C56019 PAND2X1_584/CTRL2 PAND2X1_52/B 0.03fF
C56020 PAND2X1_48/B PAND2X1_18/B 0.03fF
C56021 PAND2X1_140/A PAND2X1_854/A 0.02fF
C56022 POR2X1_326/A POR2X1_740/Y 0.03fF
C56023 POR2X1_52/A POR2X1_824/CTRL 0.01fF
C56024 PAND2X1_631/A POR2X1_625/Y 0.01fF
C56025 PAND2X1_510/CTRL POR2X1_73/Y 0.01fF
C56026 POR2X1_294/B POR2X1_722/CTRL 0.04fF
C56027 POR2X1_327/Y PAND2X1_674/a_16_344# 0.04fF
C56028 POR2X1_537/Y POR2X1_294/B 0.24fF
C56029 POR2X1_387/Y PAND2X1_114/B 0.03fF
C56030 POR2X1_741/Y POR2X1_737/A 0.03fF
C56031 POR2X1_513/B PAND2X1_304/CTRL2 0.00fF
C56032 POR2X1_41/B POR2X1_85/CTRL2 0.00fF
C56033 PAND2X1_357/Y PAND2X1_357/CTRL 0.01fF
C56034 PAND2X1_531/CTRL D_INPUT_1 0.04fF
C56035 POR2X1_193/A POR2X1_554/CTRL2 0.09fF
C56036 POR2X1_588/Y PAND2X1_651/A 0.01fF
C56037 POR2X1_760/Y POR2X1_7/B 0.01fF
C56038 POR2X1_807/A PAND2X1_72/A 0.00fF
C56039 PAND2X1_350/CTRL2 PAND2X1_341/Y 0.03fF
C56040 POR2X1_545/A POR2X1_564/O 0.00fF
C56041 POR2X1_327/Y POR2X1_605/A 0.01fF
C56042 POR2X1_864/A PAND2X1_39/B 0.05fF
C56043 POR2X1_452/A POR2X1_121/B 0.03fF
C56044 PAND2X1_6/Y POR2X1_652/A 0.07fF
C56045 POR2X1_41/B PAND2X1_857/a_76_28# 0.01fF
C56046 PAND2X1_678/O POR2X1_257/A 0.01fF
C56047 POR2X1_539/A POR2X1_733/m4_208_n4# 0.12fF
C56048 POR2X1_68/B POR2X1_774/A 0.01fF
C56049 POR2X1_786/Y POR2X1_294/A 0.03fF
C56050 POR2X1_383/A POR2X1_561/a_76_344# 0.01fF
C56051 POR2X1_476/A POR2X1_814/A 0.03fF
C56052 PAND2X1_200/O PAND2X1_193/Y 0.00fF
C56053 POR2X1_101/Y POR2X1_116/Y 0.06fF
C56054 PAND2X1_90/CTRL2 D_INPUT_1 0.00fF
C56055 POR2X1_737/A PAND2X1_32/B 0.02fF
C56056 POR2X1_648/Y POR2X1_66/A 0.03fF
C56057 POR2X1_667/O D_INPUT_0 0.01fF
C56058 POR2X1_119/Y POR2X1_255/Y 0.01fF
C56059 PAND2X1_94/A PAND2X1_748/CTRL 0.01fF
C56060 POR2X1_532/A PAND2X1_71/Y 0.02fF
C56061 PAND2X1_446/Y PAND2X1_454/B 0.01fF
C56062 POR2X1_52/A PAND2X1_207/A 0.01fF
C56063 PAND2X1_607/CTRL2 POR2X1_606/Y 0.01fF
C56064 POR2X1_93/A PAND2X1_156/A 0.11fF
C56065 POR2X1_66/Y PAND2X1_43/a_16_344# 0.01fF
C56066 POR2X1_554/B PAND2X1_93/B 0.03fF
C56067 POR2X1_333/Y POR2X1_854/B 0.05fF
C56068 POR2X1_355/B POR2X1_180/Y 0.01fF
C56069 PAND2X1_373/CTRL2 POR2X1_544/B 0.03fF
C56070 POR2X1_540/A POR2X1_188/Y 0.73fF
C56071 PAND2X1_242/Y POR2X1_5/Y 0.03fF
C56072 PAND2X1_115/CTRL POR2X1_416/B 0.01fF
C56073 POR2X1_369/O POR2X1_315/Y 0.03fF
C56074 PAND2X1_27/CTRL2 POR2X1_294/A 0.00fF
C56075 POR2X1_329/A POR2X1_594/O 0.01fF
C56076 PAND2X1_484/CTRL2 POR2X1_260/A 0.00fF
C56077 PAND2X1_508/Y PAND2X1_510/B 0.02fF
C56078 PAND2X1_223/a_76_28# PAND2X1_221/Y 0.02fF
C56079 PAND2X1_319/B PAND2X1_352/O 0.05fF
C56080 POR2X1_48/A PAND2X1_415/CTRL2 0.03fF
C56081 PAND2X1_816/CTRL PAND2X1_52/B 0.01fF
C56082 POR2X1_68/A POR2X1_736/A 0.05fF
C56083 POR2X1_447/B PAND2X1_824/O 0.15fF
C56084 POR2X1_456/B POR2X1_715/A 0.02fF
C56085 PAND2X1_448/O POR2X1_20/B 0.05fF
C56086 PAND2X1_124/O PAND2X1_123/Y 0.05fF
C56087 PAND2X1_779/O PAND2X1_550/B 0.02fF
C56088 PAND2X1_821/CTRL PAND2X1_52/B 0.01fF
C56089 POR2X1_551/A POR2X1_319/Y 0.15fF
C56090 POR2X1_539/A POR2X1_188/Y 0.94fF
C56091 POR2X1_725/Y POR2X1_512/O 0.04fF
C56092 PAND2X1_360/Y PAND2X1_343/O 0.17fF
C56093 PAND2X1_405/CTRL POR2X1_5/Y 0.01fF
C56094 PAND2X1_273/CTRL POR2X1_717/B 0.01fF
C56095 POR2X1_318/A PAND2X1_136/O 0.04fF
C56096 POR2X1_54/Y D_INPUT_0 0.53fF
C56097 POR2X1_265/Y PAND2X1_737/B 0.03fF
C56098 POR2X1_456/B POR2X1_703/O 0.04fF
C56099 POR2X1_20/B POR2X1_279/O 0.16fF
C56100 POR2X1_863/A POR2X1_579/Y 0.03fF
C56101 POR2X1_276/Y POR2X1_362/CTRL 0.01fF
C56102 POR2X1_623/B PAND2X1_9/Y 0.02fF
C56103 POR2X1_456/B POR2X1_337/Y 0.07fF
C56104 POR2X1_383/A POR2X1_510/CTRL2 0.10fF
C56105 POR2X1_407/A PAND2X1_72/A 0.22fF
C56106 POR2X1_149/O POR2X1_78/A 0.01fF
C56107 POR2X1_54/Y POR2X1_55/CTRL 0.01fF
C56108 POR2X1_156/B POR2X1_728/A 0.00fF
C56109 POR2X1_319/A POR2X1_97/A 0.03fF
C56110 POR2X1_452/Y POR2X1_121/B 0.29fF
C56111 POR2X1_351/B POR2X1_339/Y 0.00fF
C56112 PAND2X1_452/A PAND2X1_452/B 0.11fF
C56113 POR2X1_490/CTRL2 POR2X1_40/Y 0.03fF
C56114 POR2X1_66/B POR2X1_472/B 0.03fF
C56115 POR2X1_246/Y POR2X1_39/B 0.08fF
C56116 POR2X1_383/A POR2X1_862/CTRL 0.01fF
C56117 POR2X1_477/CTRL2 POR2X1_186/Y 0.16fF
C56118 POR2X1_270/Y POR2X1_218/Y 0.00fF
C56119 POR2X1_556/A PAND2X1_41/B 0.05fF
C56120 PAND2X1_73/Y POR2X1_260/B 0.26fF
C56121 POR2X1_257/A PAND2X1_161/O 0.19fF
C56122 POR2X1_614/A POR2X1_863/A 0.06fF
C56123 POR2X1_454/B POR2X1_454/A 0.14fF
C56124 POR2X1_121/A POR2X1_651/Y 0.02fF
C56125 POR2X1_87/B POR2X1_68/B 0.04fF
C56126 PAND2X1_717/A PAND2X1_151/O 0.02fF
C56127 POR2X1_180/B POR2X1_736/A 0.02fF
C56128 POR2X1_77/Y PAND2X1_112/CTRL 0.01fF
C56129 POR2X1_432/Y POR2X1_271/B 0.01fF
C56130 POR2X1_286/B POR2X1_734/A 0.02fF
C56131 PAND2X1_497/CTRL POR2X1_267/A 0.02fF
C56132 POR2X1_416/B PAND2X1_155/CTRL2 0.01fF
C56133 POR2X1_441/Y PAND2X1_544/CTRL2 0.01fF
C56134 POR2X1_43/B POR2X1_677/Y 0.03fF
C56135 POR2X1_394/A PAND2X1_379/CTRL 0.04fF
C56136 PAND2X1_64/O PAND2X1_11/Y 0.03fF
C56137 POR2X1_842/CTRL2 POR2X1_850/B 0.01fF
C56138 POR2X1_858/CTRL POR2X1_590/A 0.01fF
C56139 POR2X1_13/A PAND2X1_464/B 0.01fF
C56140 PAND2X1_72/A PAND2X1_315/CTRL 0.00fF
C56141 POR2X1_567/B POR2X1_857/O 0.02fF
C56142 POR2X1_537/Y POR2X1_567/A 0.03fF
C56143 POR2X1_83/B PAND2X1_214/CTRL 0.01fF
C56144 POR2X1_544/B POR2X1_568/B 0.01fF
C56145 POR2X1_43/B POR2X1_9/Y 0.10fF
C56146 POR2X1_66/B POR2X1_195/A 0.01fF
C56147 POR2X1_816/CTRL INPUT_0 0.03fF
C56148 POR2X1_18/a_16_28# INPUT_4 0.02fF
C56149 POR2X1_9/Y POR2X1_789/A 0.04fF
C56150 POR2X1_188/A POR2X1_866/A 0.03fF
C56151 PAND2X1_39/B POR2X1_362/B 0.96fF
C56152 POR2X1_648/CTRL PAND2X1_90/Y 0.06fF
C56153 PAND2X1_507/O POR2X1_39/B 0.02fF
C56154 POR2X1_54/Y PAND2X1_90/Y 0.03fF
C56155 PAND2X1_476/CTRL PAND2X1_571/A 0.01fF
C56156 PAND2X1_414/CTRL2 POR2X1_42/Y 0.16fF
C56157 POR2X1_20/B PAND2X1_151/CTRL 0.00fF
C56158 PAND2X1_704/O POR2X1_77/Y 0.11fF
C56159 POR2X1_119/Y POR2X1_518/O 0.08fF
C56160 POR2X1_14/Y POR2X1_496/Y 0.07fF
C56161 D_INPUT_5 PAND2X1_18/O 0.15fF
C56162 PAND2X1_838/B VDD 0.00fF
C56163 POR2X1_411/B PAND2X1_785/Y 0.03fF
C56164 POR2X1_440/Y POR2X1_863/A 3.01fF
C56165 PAND2X1_159/CTRL POR2X1_29/A 0.01fF
C56166 PAND2X1_226/CTRL POR2X1_227/A 0.00fF
C56167 POR2X1_9/Y POR2X1_38/B 0.23fF
C56168 PAND2X1_833/a_16_344# POR2X1_257/A 0.01fF
C56169 POR2X1_435/B VDD 0.10fF
C56170 PAND2X1_244/CTRL2 POR2X1_102/Y 0.01fF
C56171 POR2X1_83/B POR2X1_423/O 0.05fF
C56172 POR2X1_66/Y VDD 0.22fF
C56173 PAND2X1_223/B POR2X1_283/Y 0.06fF
C56174 POR2X1_49/CTRL2 POR2X1_29/A 0.01fF
C56175 POR2X1_568/A POR2X1_444/Y 0.03fF
C56176 POR2X1_814/A POR2X1_513/Y 0.03fF
C56177 POR2X1_78/B POR2X1_602/CTRL 0.06fF
C56178 PAND2X1_243/B POR2X1_20/B 0.03fF
C56179 PAND2X1_410/O POR2X1_236/Y 0.02fF
C56180 POR2X1_707/B PAND2X1_47/B 0.97fF
C56181 PAND2X1_46/CTRL POR2X1_296/B 0.00fF
C56182 POR2X1_647/B POR2X1_121/Y 0.03fF
C56183 POR2X1_98/A PAND2X1_60/B 0.01fF
C56184 PAND2X1_23/Y POR2X1_227/B 0.00fF
C56185 PAND2X1_362/A PAND2X1_354/A 0.09fF
C56186 POR2X1_427/O POR2X1_427/Y 0.02fF
C56187 POR2X1_664/CTRL POR2X1_651/Y 0.01fF
C56188 POR2X1_112/a_56_344# POR2X1_632/Y 0.00fF
C56189 POR2X1_695/Y PAND2X1_712/B 0.01fF
C56190 PAND2X1_222/A PAND2X1_364/B 0.03fF
C56191 POR2X1_814/A POR2X1_205/A 0.10fF
C56192 POR2X1_67/Y POR2X1_619/Y 0.00fF
C56193 POR2X1_82/CTRL POR2X1_409/B 0.01fF
C56194 PAND2X1_782/Y VDD 0.09fF
C56195 POR2X1_61/Y POR2X1_400/B 0.02fF
C56196 POR2X1_689/CTRL2 POR2X1_32/A 0.03fF
C56197 PAND2X1_392/O POR2X1_236/Y 0.02fF
C56198 POR2X1_260/B PAND2X1_132/CTRL2 0.03fF
C56199 POR2X1_474/O PAND2X1_41/B 0.16fF
C56200 POR2X1_66/A INPUT_0 0.22fF
C56201 POR2X1_114/B POR2X1_475/O 0.03fF
C56202 PAND2X1_256/CTRL2 POR2X1_205/A 0.05fF
C56203 POR2X1_96/A PAND2X1_644/Y 0.00fF
C56204 PAND2X1_400/CTRL VDD -0.00fF
C56205 POR2X1_432/O POR2X1_236/Y 0.01fF
C56206 POR2X1_736/A POR2X1_169/A 0.05fF
C56207 PAND2X1_48/B PAND2X1_248/CTRL 0.01fF
C56208 POR2X1_60/A POR2X1_5/Y 0.59fF
C56209 PAND2X1_116/CTRL2 POR2X1_40/Y 0.01fF
C56210 POR2X1_397/Y PAND2X1_721/B 0.10fF
C56211 POR2X1_614/A POR2X1_841/a_76_344# 0.01fF
C56212 GATE_479 POR2X1_40/Y 0.03fF
C56213 PAND2X1_761/CTRL PAND2X1_32/B 0.01fF
C56214 POR2X1_86/a_16_28# POR2X1_85/Y 0.04fF
C56215 POR2X1_859/A PAND2X1_381/Y 0.03fF
C56216 PAND2X1_257/O POR2X1_259/B 0.02fF
C56217 PAND2X1_570/a_76_28# PAND2X1_562/Y 0.02fF
C56218 POR2X1_484/CTRL2 POR2X1_763/Y 0.03fF
C56219 PAND2X1_795/B POR2X1_498/Y 0.03fF
C56220 POR2X1_754/Y POR2X1_754/A 0.01fF
C56221 POR2X1_48/A PAND2X1_254/O 0.03fF
C56222 POR2X1_296/Y VDD 0.30fF
C56223 POR2X1_341/A POR2X1_541/O 0.02fF
C56224 POR2X1_465/O POR2X1_569/A 0.02fF
C56225 POR2X1_181/a_56_344# PAND2X1_72/A 0.00fF
C56226 POR2X1_556/A POR2X1_228/Y 0.13fF
C56227 POR2X1_405/Y POR2X1_296/B 0.03fF
C56228 POR2X1_634/CTRL2 INPUT_0 0.30fF
C56229 POR2X1_816/Y D_INPUT_1 0.94fF
C56230 POR2X1_52/A POR2X1_753/Y 0.07fF
C56231 POR2X1_243/B POR2X1_38/B 0.01fF
C56232 POR2X1_330/Y PAND2X1_131/CTRL2 0.03fF
C56233 POR2X1_78/A POR2X1_646/CTRL 0.00fF
C56234 POR2X1_606/CTRL PAND2X1_32/B 0.01fF
C56235 POR2X1_416/B POR2X1_747/O 0.16fF
C56236 POR2X1_41/B PAND2X1_443/Y 0.05fF
C56237 POR2X1_68/A POR2X1_270/Y 0.03fF
C56238 POR2X1_411/B PAND2X1_656/A 0.37fF
C56239 D_INPUT_2 POR2X1_37/Y 0.12fF
C56240 PAND2X1_259/CTRL POR2X1_258/Y 0.01fF
C56241 POR2X1_57/A POR2X1_442/a_16_28# 0.03fF
C56242 POR2X1_102/Y POR2X1_275/CTRL2 0.01fF
C56243 POR2X1_814/B POR2X1_362/B 0.03fF
C56244 POR2X1_496/Y POR2X1_55/Y 0.24fF
C56245 POR2X1_65/A POR2X1_485/CTRL 0.01fF
C56246 POR2X1_257/A PAND2X1_149/A 0.03fF
C56247 POR2X1_302/B VDD 0.04fF
C56248 PAND2X1_498/O POR2X1_590/A 0.01fF
C56249 POR2X1_271/Y PAND2X1_785/Y 0.03fF
C56250 POR2X1_78/B POR2X1_788/O 0.08fF
C56251 POR2X1_300/CTRL POR2X1_32/A 0.01fF
C56252 PAND2X1_93/B POR2X1_702/A 0.03fF
C56253 PAND2X1_443/CTRL POR2X1_91/Y 0.01fF
C56254 POR2X1_400/A PAND2X1_41/B 0.03fF
C56255 PAND2X1_73/Y PAND2X1_55/Y 0.18fF
C56256 POR2X1_499/A POR2X1_276/Y 0.03fF
C56257 POR2X1_720/Y POR2X1_546/A 0.01fF
C56258 PAND2X1_57/B POR2X1_330/Y 0.08fF
C56259 POR2X1_343/Y POR2X1_343/B 0.01fF
C56260 POR2X1_392/B VDD 0.01fF
C56261 PAND2X1_93/B POR2X1_243/O 0.01fF
C56262 POR2X1_41/B PAND2X1_557/A 0.03fF
C56263 PAND2X1_56/Y POR2X1_660/Y 0.05fF
C56264 POR2X1_51/CTRL PAND2X1_635/Y 0.01fF
C56265 PAND2X1_84/Y PAND2X1_558/CTRL2 0.01fF
C56266 PAND2X1_104/a_76_28# PAND2X1_8/Y 0.03fF
C56267 POR2X1_141/CTRL2 VDD 0.00fF
C56268 PAND2X1_841/O POR2X1_516/Y 0.01fF
C56269 PAND2X1_674/O POR2X1_590/A 0.04fF
C56270 PAND2X1_455/CTRL2 POR2X1_7/B 0.00fF
C56271 POR2X1_150/Y PAND2X1_175/m4_208_n4# 0.08fF
C56272 POR2X1_20/B POR2X1_260/A 0.03fF
C56273 POR2X1_620/O POR2X1_296/B 0.02fF
C56274 POR2X1_346/B PAND2X1_43/CTRL 0.00fF
C56275 PAND2X1_73/Y PAND2X1_79/a_56_28# 0.00fF
C56276 POR2X1_241/B POR2X1_341/O 0.02fF
C56277 POR2X1_245/CTRL2 POR2X1_37/Y 0.00fF
C56278 POR2X1_846/Y POR2X1_129/Y 0.01fF
C56279 PAND2X1_592/Y POR2X1_72/B 0.03fF
C56280 PAND2X1_94/A POR2X1_621/A 0.02fF
C56281 POR2X1_72/B PAND2X1_174/CTRL2 0.03fF
C56282 POR2X1_854/CTRL2 POR2X1_567/B -0.00fF
C56283 PAND2X1_56/Y POR2X1_657/a_16_28# 0.08fF
C56284 POR2X1_411/B PAND2X1_348/A 0.09fF
C56285 GATE_741 PAND2X1_366/Y 0.01fF
C56286 POR2X1_814/A POR2X1_383/a_76_344# 0.01fF
C56287 POR2X1_66/B PAND2X1_638/CTRL 0.00fF
C56288 PAND2X1_76/Y PAND2X1_775/CTRL2 0.03fF
C56289 POR2X1_66/A PAND2X1_393/CTRL2 0.02fF
C56290 PAND2X1_96/B POR2X1_479/CTRL 0.01fF
C56291 PAND2X1_73/Y POR2X1_407/Y 0.03fF
C56292 PAND2X1_218/B PAND2X1_717/Y 0.05fF
C56293 POR2X1_104/CTRL D_INPUT_1 0.01fF
C56294 PAND2X1_469/B PAND2X1_444/Y 0.00fF
C56295 POR2X1_302/B POR2X1_741/Y 0.03fF
C56296 POR2X1_278/Y PAND2X1_659/CTRL 0.03fF
C56297 PAND2X1_192/O PAND2X1_191/Y 0.01fF
C56298 POR2X1_473/a_16_28# POR2X1_773/B 0.06fF
C56299 POR2X1_29/Y POR2X1_159/CTRL 0.00fF
C56300 POR2X1_396/Y POR2X1_669/B 0.09fF
C56301 PAND2X1_854/O PAND2X1_805/A 0.02fF
C56302 PAND2X1_225/CTRL2 POR2X1_38/B 0.01fF
C56303 POR2X1_32/A POR2X1_387/Y 0.12fF
C56304 PAND2X1_753/CTRL VDD -0.00fF
C56305 POR2X1_66/B POR2X1_501/B 0.03fF
C56306 POR2X1_295/O POR2X1_90/Y 0.01fF
C56307 PAND2X1_65/B POR2X1_832/B 0.01fF
C56308 POR2X1_96/A PAND2X1_549/CTRL 0.00fF
C56309 POR2X1_566/A POR2X1_724/O 0.04fF
C56310 PAND2X1_610/a_76_28# POR2X1_612/A 0.04fF
C56311 PAND2X1_736/Y PAND2X1_473/B 0.05fF
C56312 PAND2X1_42/CTRL2 D_INPUT_1 0.02fF
C56313 POR2X1_15/a_56_344# POR2X1_14/Y 0.00fF
C56314 POR2X1_218/Y POR2X1_101/Y 0.13fF
C56315 PAND2X1_451/O POR2X1_428/Y 0.01fF
C56316 PAND2X1_832/O POR2X1_433/Y 0.00fF
C56317 POR2X1_302/B PAND2X1_32/B 0.03fF
C56318 POR2X1_60/A POR2X1_665/A 0.00fF
C56319 POR2X1_312/Y PAND2X1_182/O 0.02fF
C56320 PAND2X1_6/Y POR2X1_274/Y 0.03fF
C56321 POR2X1_96/A PAND2X1_254/Y 0.06fF
C56322 POR2X1_174/A POR2X1_854/B 0.08fF
C56323 POR2X1_260/B POR2X1_576/a_16_28# 0.01fF
C56324 PAND2X1_478/CTRL POR2X1_236/Y 0.01fF
C56325 D_INPUT_5 PAND2X1_18/B 1.19fF
C56326 POR2X1_65/A PAND2X1_779/Y 0.01fF
C56327 POR2X1_557/A PAND2X1_63/a_16_344# 0.03fF
C56328 PAND2X1_631/A POR2X1_411/B 0.07fF
C56329 POR2X1_392/B PAND2X1_32/B 1.87fF
C56330 POR2X1_77/a_16_28# POR2X1_394/A 0.01fF
C56331 POR2X1_674/Y POR2X1_283/A 0.06fF
C56332 PAND2X1_435/O POR2X1_293/Y 0.07fF
C56333 POR2X1_590/A POR2X1_796/A 0.02fF
C56334 PAND2X1_57/B POR2X1_247/O 0.01fF
C56335 POR2X1_236/Y POR2X1_395/a_16_28# 0.02fF
C56336 POR2X1_300/CTRL2 POR2X1_13/A 0.01fF
C56337 POR2X1_823/CTRL2 POR2X1_236/Y 0.01fF
C56338 POR2X1_40/Y POR2X1_142/Y 0.06fF
C56339 PAND2X1_13/m4_208_n4# POR2X1_222/Y 0.08fF
C56340 PAND2X1_215/B POR2X1_46/Y 0.07fF
C56341 PAND2X1_281/CTRL POR2X1_862/A 0.07fF
C56342 PAND2X1_480/B POR2X1_42/Y 0.05fF
C56343 POR2X1_335/O POR2X1_741/Y 0.01fF
C56344 POR2X1_57/A PAND2X1_139/O 0.02fF
C56345 POR2X1_417/Y POR2X1_387/Y 0.08fF
C56346 POR2X1_65/A PAND2X1_509/CTRL 0.02fF
C56347 POR2X1_65/A POR2X1_321/a_16_28# 0.03fF
C56348 POR2X1_283/A POR2X1_226/a_16_28# 0.05fF
C56349 POR2X1_539/A POR2X1_457/CTRL 0.00fF
C56350 PAND2X1_467/Y PAND2X1_467/B 1.66fF
C56351 PAND2X1_23/Y PAND2X1_238/CTRL2 0.00fF
C56352 POR2X1_496/Y PAND2X1_508/O 0.07fF
C56353 POR2X1_305/Y VDD 0.15fF
C56354 POR2X1_697/O PAND2X1_565/A 0.00fF
C56355 POR2X1_754/A POR2X1_42/Y 0.19fF
C56356 PAND2X1_31/CTRL PAND2X1_18/B 0.03fF
C56357 POR2X1_83/B POR2X1_428/CTRL 0.01fF
C56358 POR2X1_823/O VDD 0.00fF
C56359 POR2X1_248/CTRL2 VDD 0.00fF
C56360 POR2X1_41/B POR2X1_495/Y 0.06fF
C56361 PAND2X1_40/CTRL2 PAND2X1_57/B 0.00fF
C56362 POR2X1_49/Y PAND2X1_149/A 0.09fF
C56363 PAND2X1_605/a_16_344# POR2X1_32/A 0.02fF
C56364 PAND2X1_6/Y POR2X1_370/Y 0.10fF
C56365 PAND2X1_622/O POR2X1_619/Y 0.02fF
C56366 POR2X1_178/Y POR2X1_60/A 0.01fF
C56367 POR2X1_78/B POR2X1_556/Y 0.05fF
C56368 POR2X1_57/A POR2X1_122/A 0.02fF
C56369 PAND2X1_65/B POR2X1_577/O 0.02fF
C56370 PAND2X1_810/A PAND2X1_810/CTRL2 0.01fF
C56371 POR2X1_722/B PAND2X1_48/B 0.04fF
C56372 POR2X1_463/Y PAND2X1_58/A 0.01fF
C56373 PAND2X1_393/O PAND2X1_41/B 0.01fF
C56374 POR2X1_78/B PAND2X1_81/a_16_344# 0.00fF
C56375 PAND2X1_48/B POR2X1_294/B 1.95fF
C56376 POR2X1_366/Y PAND2X1_48/B 2.21fF
C56377 POR2X1_259/B POR2X1_555/B 0.05fF
C56378 D_INPUT_2 POR2X1_293/Y 0.04fF
C56379 POR2X1_862/B POR2X1_537/A 0.00fF
C56380 PAND2X1_58/A POR2X1_756/Y 0.01fF
C56381 PAND2X1_814/O VDD -0.00fF
C56382 PAND2X1_65/B PAND2X1_534/CTRL2 0.01fF
C56383 POR2X1_72/B POR2X1_172/CTRL 0.01fF
C56384 POR2X1_283/A PAND2X1_562/B 0.07fF
C56385 POR2X1_55/Y PAND2X1_514/Y 0.93fF
C56386 PAND2X1_41/B POR2X1_180/A 0.06fF
C56387 PAND2X1_106/O POR2X1_105/Y 0.10fF
C56388 PAND2X1_23/Y POR2X1_469/a_56_344# 0.00fF
C56389 POR2X1_502/A PAND2X1_69/A 0.13fF
C56390 POR2X1_804/A PAND2X1_516/O 0.18fF
C56391 POR2X1_52/A POR2X1_315/O 0.01fF
C56392 PAND2X1_90/Y POR2X1_148/B 0.01fF
C56393 POR2X1_532/A INPUT_0 0.20fF
C56394 POR2X1_455/O PAND2X1_60/B 0.01fF
C56395 PAND2X1_862/B POR2X1_73/Y 0.03fF
C56396 PAND2X1_472/A POR2X1_669/O 0.01fF
C56397 POR2X1_376/A VDD -0.00fF
C56398 VDD POR2X1_578/O 0.00fF
C56399 PAND2X1_793/Y PAND2X1_548/CTRL 0.01fF
C56400 POR2X1_65/A POR2X1_73/O 0.16fF
C56401 PAND2X1_298/O POR2X1_750/B 0.09fF
C56402 POR2X1_43/B POR2X1_586/a_16_28# 0.01fF
C56403 POR2X1_788/Y PAND2X1_144/CTRL 0.00fF
C56404 POR2X1_300/CTRL POR2X1_184/Y 0.00fF
C56405 VDD PAND2X1_305/CTRL2 -0.00fF
C56406 POR2X1_155/CTRL2 POR2X1_162/Y 0.01fF
C56407 PAND2X1_716/CTRL PAND2X1_197/Y 0.00fF
C56408 POR2X1_60/A PAND2X1_337/O 0.19fF
C56409 D_INPUT_0 POR2X1_4/Y 0.10fF
C56410 POR2X1_504/Y INPUT_1 0.03fF
C56411 PAND2X1_460/CTRL2 POR2X1_7/B 0.00fF
C56412 PAND2X1_69/A PAND2X1_176/O 0.02fF
C56413 PAND2X1_717/A PAND2X1_860/A 0.03fF
C56414 PAND2X1_730/a_76_28# POR2X1_42/Y 0.01fF
C56415 POR2X1_830/Y POR2X1_737/A 0.02fF
C56416 PAND2X1_530/CTRL2 PAND2X1_69/A 0.01fF
C56417 PAND2X1_55/Y POR2X1_631/B 0.02fF
C56418 POR2X1_283/A PAND2X1_715/CTRL 0.02fF
C56419 PAND2X1_675/A PAND2X1_357/Y 0.03fF
C56420 POR2X1_632/O POR2X1_632/Y 0.01fF
C56421 PAND2X1_839/O PAND2X1_835/Y 0.00fF
C56422 POR2X1_440/CTRL POR2X1_440/B 0.01fF
C56423 PAND2X1_469/B PAND2X1_357/Y 0.36fF
C56424 POR2X1_832/A POR2X1_722/Y 0.60fF
C56425 PAND2X1_63/Y POR2X1_264/Y 0.31fF
C56426 POR2X1_13/A POR2X1_283/A 0.26fF
C56427 POR2X1_325/O POR2X1_502/A 0.02fF
C56428 PAND2X1_254/Y POR2X1_7/A 0.03fF
C56429 PAND2X1_494/CTRL PAND2X1_32/B 0.01fF
C56430 PAND2X1_260/CTRL PAND2X1_345/Y 0.01fF
C56431 POR2X1_260/Y POR2X1_205/A 0.00fF
C56432 POR2X1_383/A PAND2X1_322/CTRL 0.05fF
C56433 POR2X1_334/A POR2X1_814/B 0.02fF
C56434 POR2X1_52/A PAND2X1_656/A 0.02fF
C56435 POR2X1_537/Y POR2X1_643/A 0.04fF
C56436 PAND2X1_862/B PAND2X1_244/B 0.03fF
C56437 PAND2X1_865/Y POR2X1_102/Y 0.04fF
C56438 POR2X1_198/O POR2X1_532/A 0.01fF
C56439 POR2X1_333/A POR2X1_551/A 0.05fF
C56440 PAND2X1_48/B PAND2X1_111/B 0.03fF
C56441 PAND2X1_283/O PAND2X1_96/B 0.01fF
C56442 POR2X1_38/Y PAND2X1_188/a_76_28# 0.01fF
C56443 POR2X1_306/CTRL POR2X1_43/B 0.01fF
C56444 POR2X1_60/CTRL2 PAND2X1_651/Y 0.30fF
C56445 POR2X1_78/O PAND2X1_96/B 0.09fF
C56446 PAND2X1_534/O POR2X1_294/B 0.12fF
C56447 POR2X1_260/Y POR2X1_366/A 0.02fF
C56448 POR2X1_388/O PAND2X1_69/A 0.01fF
C56449 PAND2X1_715/B PAND2X1_715/a_16_344# 0.05fF
C56450 POR2X1_841/B POR2X1_717/B 0.03fF
C56451 POR2X1_754/A POR2X1_754/CTRL 0.01fF
C56452 PAND2X1_476/A POR2X1_72/B 0.03fF
C56453 PAND2X1_140/A PAND2X1_675/A 0.03fF
C56454 POR2X1_519/CTRL2 POR2X1_42/Y 0.03fF
C56455 POR2X1_254/Y POR2X1_332/O 0.09fF
C56456 PAND2X1_537/CTRL PAND2X1_364/B 0.03fF
C56457 POR2X1_315/Y PAND2X1_302/CTRL2 0.00fF
C56458 POR2X1_537/Y POR2X1_807/A 0.02fF
C56459 PAND2X1_264/CTRL2 POR2X1_42/Y 0.00fF
C56460 POR2X1_508/B PAND2X1_41/B 0.03fF
C56461 POR2X1_68/B PAND2X1_153/CTRL2 0.01fF
C56462 INPUT_1 POR2X1_586/O 0.01fF
C56463 POR2X1_57/A PAND2X1_653/Y 0.06fF
C56464 POR2X1_276/A POR2X1_130/Y 0.02fF
C56465 POR2X1_599/A POR2X1_7/A 0.03fF
C56466 POR2X1_566/A POR2X1_97/a_76_344# 0.03fF
C56467 POR2X1_40/Y POR2X1_524/CTRL 0.09fF
C56468 POR2X1_616/Y POR2X1_847/B 0.02fF
C56469 PAND2X1_148/CTRL PAND2X1_148/Y 0.01fF
C56470 POR2X1_740/Y POR2X1_787/CTRL 0.08fF
C56471 PAND2X1_651/Y POR2X1_387/Y 0.10fF
C56472 POR2X1_631/A PAND2X1_96/B -0.01fF
C56473 PAND2X1_72/a_56_28# POR2X1_532/A 0.00fF
C56474 PAND2X1_697/O POR2X1_383/A 0.00fF
C56475 POR2X1_346/B POR2X1_740/Y 0.05fF
C56476 POR2X1_532/A POR2X1_780/A 0.01fF
C56477 PAND2X1_631/A POR2X1_376/B 0.05fF
C56478 PAND2X1_839/B PAND2X1_835/Y 0.02fF
C56479 POR2X1_383/A POR2X1_713/a_16_28# 0.01fF
C56480 POR2X1_545/A POR2X1_551/CTRL2 0.01fF
C56481 POR2X1_619/A POR2X1_751/O 0.01fF
C56482 PAND2X1_56/Y POR2X1_308/B 0.03fF
C56483 PAND2X1_493/O PAND2X1_480/B 0.06fF
C56484 POR2X1_264/Y POR2X1_260/A 0.02fF
C56485 PAND2X1_56/Y POR2X1_787/O 0.03fF
C56486 POR2X1_60/a_16_28# POR2X1_38/Y 0.01fF
C56487 PAND2X1_7/CTRL2 POR2X1_259/B 0.01fF
C56488 POR2X1_96/A PAND2X1_779/CTRL 0.00fF
C56489 POR2X1_364/A POR2X1_568/Y 0.95fF
C56490 POR2X1_416/B PAND2X1_403/B 0.07fF
C56491 PAND2X1_557/A POR2X1_77/Y 0.05fF
C56492 POR2X1_20/B POR2X1_329/A 0.03fF
C56493 PAND2X1_341/B INPUT_0 0.02fF
C56494 POR2X1_364/A POR2X1_785/B 0.07fF
C56495 PAND2X1_105/CTRL2 PAND2X1_348/A 0.04fF
C56496 POR2X1_207/A POR2X1_199/B 0.04fF
C56497 PAND2X1_55/Y POR2X1_576/a_16_28# 0.03fF
C56498 POR2X1_383/A POR2X1_758/O 0.02fF
C56499 PAND2X1_472/CTRL PAND2X1_472/A 0.03fF
C56500 POR2X1_124/B POR2X1_773/B 0.05fF
C56501 POR2X1_355/B POR2X1_508/A 0.01fF
C56502 PAND2X1_372/a_16_344# PAND2X1_48/A 0.01fF
C56503 VDD PAND2X1_304/CTRL2 0.00fF
C56504 PAND2X1_546/Y POR2X1_394/A 0.12fF
C56505 D_INPUT_3 PAND2X1_63/B 0.03fF
C56506 PAND2X1_6/A POR2X1_376/O 0.07fF
C56507 POR2X1_287/B POR2X1_343/a_56_344# 0.00fF
C56508 POR2X1_119/Y POR2X1_46/Y 0.15fF
C56509 POR2X1_137/Y POR2X1_218/CTRL 0.00fF
C56510 POR2X1_669/B PAND2X1_147/CTRL2 0.03fF
C56511 POR2X1_863/A POR2X1_590/A 0.03fF
C56512 PAND2X1_96/B POR2X1_463/Y 0.05fF
C56513 POR2X1_433/Y POR2X1_153/Y 0.53fF
C56514 PAND2X1_473/CTRL PAND2X1_216/B 0.01fF
C56515 PAND2X1_96/B POR2X1_756/Y 0.02fF
C56516 POR2X1_172/Y POR2X1_530/CTRL 0.04fF
C56517 POR2X1_66/CTRL PAND2X1_39/B 0.01fF
C56518 POR2X1_548/B PAND2X1_143/CTRL 0.01fF
C56519 PAND2X1_481/a_76_28# POR2X1_222/Y 0.02fF
C56520 POR2X1_283/A PAND2X1_510/B 0.02fF
C56521 POR2X1_556/A POR2X1_657/Y 0.06fF
C56522 PAND2X1_48/B POR2X1_567/A 3.87fF
C56523 POR2X1_712/CTRL POR2X1_260/A 0.01fF
C56524 POR2X1_653/CTRL POR2X1_711/Y 0.04fF
C56525 POR2X1_703/Y POR2X1_724/A 0.04fF
C56526 POR2X1_177/O POR2X1_90/Y 0.02fF
C56527 POR2X1_458/Y D_INPUT_0 0.03fF
C56528 POR2X1_809/A POR2X1_810/a_16_28# 0.02fF
C56529 POR2X1_355/B POR2X1_568/B 26.70fF
C56530 POR2X1_13/Y PAND2X1_643/A 0.15fF
C56531 POR2X1_264/Y PAND2X1_517/CTRL2 0.01fF
C56532 POR2X1_537/Y POR2X1_407/A 0.03fF
C56533 POR2X1_658/O POR2X1_624/Y 0.01fF
C56534 POR2X1_3/A POR2X1_394/A 0.02fF
C56535 PAND2X1_808/Y PAND2X1_865/Y 0.23fF
C56536 PAND2X1_6/Y POR2X1_359/CTRL 0.00fF
C56537 POR2X1_9/Y POR2X1_590/A 0.07fF
C56538 PAND2X1_48/B POR2X1_542/O 0.01fF
C56539 POR2X1_249/Y POR2X1_773/CTRL2 0.01fF
C56540 POR2X1_704/CTRL2 POR2X1_317/B 0.00fF
C56541 POR2X1_303/CTRL POR2X1_513/Y 0.03fF
C56542 PAND2X1_716/B POR2X1_73/Y 0.03fF
C56543 POR2X1_293/Y POR2X1_372/CTRL 0.01fF
C56544 POR2X1_259/CTRL POR2X1_260/A 0.01fF
C56545 PAND2X1_6/Y POR2X1_552/A 0.33fF
C56546 POR2X1_123/B PAND2X1_48/A 0.01fF
C56547 PAND2X1_69/A POR2X1_188/Y 0.06fF
C56548 POR2X1_68/A POR2X1_359/a_16_28# 0.07fF
C56549 POR2X1_416/B POR2X1_232/CTRL2 0.01fF
C56550 POR2X1_7/B POR2X1_588/O 0.02fF
C56551 PAND2X1_290/O POR2X1_334/B 0.02fF
C56552 POR2X1_762/a_76_344# D_INPUT_6 0.00fF
C56553 POR2X1_518/CTRL2 POR2X1_73/Y 0.04fF
C56554 PAND2X1_330/O POR2X1_594/A 0.00fF
C56555 PAND2X1_189/O POR2X1_854/B 0.28fF
C56556 POR2X1_683/Y POR2X1_761/A 0.00fF
C56557 POR2X1_66/Y PAND2X1_67/a_16_344# 0.01fF
C56558 POR2X1_495/Y POR2X1_77/Y 0.18fF
C56559 PAND2X1_193/Y PAND2X1_596/CTRL2 0.03fF
C56560 POR2X1_78/Y D_INPUT_0 0.01fF
C56561 POR2X1_508/A POR2X1_510/B 0.01fF
C56562 PAND2X1_737/B PAND2X1_853/B 0.03fF
C56563 POR2X1_353/A POR2X1_731/A 0.01fF
C56564 POR2X1_71/Y PAND2X1_501/m4_208_n4# 0.12fF
C56565 PAND2X1_216/B PAND2X1_853/B 0.03fF
C56566 PAND2X1_680/CTRL POR2X1_162/Y 0.01fF
C56567 PAND2X1_6/Y POR2X1_342/A 0.01fF
C56568 PAND2X1_118/CTRL2 PAND2X1_72/A 0.01fF
C56569 POR2X1_362/Y POR2X1_554/B 0.02fF
C56570 PAND2X1_433/O PAND2X1_72/A 0.02fF
C56571 POR2X1_647/B POR2X1_286/O 0.01fF
C56572 POR2X1_463/a_16_28# POR2X1_750/B 0.03fF
C56573 PAND2X1_65/B PAND2X1_224/O 0.02fF
C56574 POR2X1_294/Y PAND2X1_67/CTRL 0.01fF
C56575 PAND2X1_96/B POR2X1_736/A 0.12fF
C56576 PAND2X1_472/a_76_28# POR2X1_153/Y 0.00fF
C56577 POR2X1_41/B PAND2X1_860/A 0.03fF
C56578 POR2X1_123/a_16_28# PAND2X1_72/A 0.09fF
C56579 PAND2X1_269/m4_208_n4# POR2X1_72/B 0.15fF
C56580 POR2X1_736/A POR2X1_736/CTRL2 0.02fF
C56581 POR2X1_67/Y POR2X1_668/CTRL2 0.10fF
C56582 POR2X1_74/m4_208_n4# POR2X1_271/A 0.07fF
C56583 POR2X1_537/CTRL POR2X1_537/Y 0.01fF
C56584 POR2X1_527/a_56_344# POR2X1_110/Y 0.01fF
C56585 POR2X1_114/B POR2X1_717/B 0.06fF
C56586 POR2X1_316/a_56_344# POR2X1_153/Y 0.03fF
C56587 POR2X1_42/Y PAND2X1_850/CTRL2 0.01fF
C56588 POR2X1_104/CTRL INPUT_3 0.00fF
C56589 POR2X1_441/Y PAND2X1_545/O 0.03fF
C56590 POR2X1_25/Y POR2X1_394/A 0.49fF
C56591 PAND2X1_815/O POR2X1_814/Y -0.00fF
C56592 POR2X1_394/A POR2X1_701/CTRL 0.01fF
C56593 POR2X1_42/Y POR2X1_386/Y 0.07fF
C56594 PAND2X1_73/CTRL2 PAND2X1_9/Y 0.01fF
C56595 POR2X1_123/Y PAND2X1_72/A 0.03fF
C56596 PAND2X1_458/a_16_344# PAND2X1_785/Y 0.03fF
C56597 POR2X1_9/Y PAND2X1_350/A 0.04fF
C56598 POR2X1_250/Y POR2X1_488/a_76_344# 0.01fF
C56599 POR2X1_846/Y POR2X1_615/O 0.03fF
C56600 PAND2X1_863/m4_208_n4# POR2X1_282/m4_208_n4# 0.13fF
C56601 PAND2X1_651/O PAND2X1_639/Y 0.05fF
C56602 POR2X1_458/B POR2X1_717/B 0.15fF
C56603 POR2X1_274/A POR2X1_590/A 0.03fF
C56604 POR2X1_78/A PAND2X1_609/O 0.02fF
C56605 PAND2X1_261/CTRL POR2X1_814/A 0.05fF
C56606 POR2X1_540/Y POR2X1_186/B 0.03fF
C56607 POR2X1_566/B POR2X1_567/O 0.28fF
C56608 POR2X1_66/B PAND2X1_60/O 0.15fF
C56609 POR2X1_99/B POR2X1_228/CTRL2 0.00fF
C56610 POR2X1_294/CTRL2 POR2X1_355/A 0.01fF
C56611 PAND2X1_629/CTRL2 POR2X1_628/Y 0.00fF
C56612 POR2X1_137/B POR2X1_640/A -0.01fF
C56613 PAND2X1_63/B PAND2X1_52/B 0.03fF
C56614 PAND2X1_60/B POR2X1_301/m4_208_n4# 0.15fF
C56615 POR2X1_479/B POR2X1_479/CTRL2 0.01fF
C56616 POR2X1_730/Y POR2X1_711/Y 0.07fF
C56617 POR2X1_343/Y POR2X1_260/A 0.09fF
C56618 POR2X1_14/Y PAND2X1_448/CTRL2 0.00fF
C56619 POR2X1_96/A PAND2X1_447/CTRL2 0.01fF
C56620 POR2X1_460/Y POR2X1_459/CTRL 0.01fF
C56621 POR2X1_864/A VDD 0.08fF
C56622 POR2X1_825/Y POR2X1_291/Y 0.00fF
C56623 PAND2X1_207/CTRL POR2X1_72/B 0.01fF
C56624 POR2X1_411/B PAND2X1_715/CTRL2 0.01fF
C56625 PAND2X1_200/B POR2X1_39/B 0.02fF
C56626 POR2X1_730/Y POR2X1_728/A 0.08fF
C56627 PAND2X1_246/O POR2X1_404/Y 0.01fF
C56628 PAND2X1_58/A PAND2X1_37/CTRL2 0.12fF
C56629 PAND2X1_73/Y POR2X1_174/A 0.00fF
C56630 POR2X1_257/A POR2X1_236/Y 0.25fF
C56631 POR2X1_101/Y POR2X1_138/A 0.05fF
C56632 POR2X1_175/m4_208_n4# POR2X1_465/m4_208_n4# 0.04fF
C56633 POR2X1_294/Y POR2X1_202/CTRL2 0.00fF
C56634 PAND2X1_267/a_56_28# POR2X1_72/B 0.00fF
C56635 POR2X1_409/B POR2X1_40/Y 0.07fF
C56636 POR2X1_234/Y POR2X1_411/B 0.01fF
C56637 POR2X1_553/a_16_28# POR2X1_632/Y 0.01fF
C56638 PAND2X1_93/B POR2X1_653/B 0.05fF
C56639 POR2X1_106/a_16_28# POR2X1_102/Y 0.03fF
C56640 POR2X1_174/B PAND2X1_20/A 0.03fF
C56641 PAND2X1_56/Y PAND2X1_45/CTRL 0.00fF
C56642 POR2X1_376/B POR2X1_699/O 0.18fF
C56643 POR2X1_470/a_16_28# POR2X1_467/Y 0.04fF
C56644 POR2X1_760/A POR2X1_599/A 0.10fF
C56645 POR2X1_463/CTRL2 POR2X1_532/A 0.03fF
C56646 POR2X1_60/A PAND2X1_200/CTRL 0.01fF
C56647 POR2X1_450/B POR2X1_121/B 0.01fF
C56648 PAND2X1_65/B PAND2X1_65/CTRL 0.01fF
C56649 POR2X1_815/Y VDD 0.00fF
C56650 PAND2X1_39/B POR2X1_828/CTRL2 0.02fF
C56651 POR2X1_102/Y POR2X1_609/CTRL 0.01fF
C56652 POR2X1_78/A PAND2X1_42/CTRL2 0.02fF
C56653 POR2X1_270/Y POR2X1_457/B 0.01fF
C56654 POR2X1_612/Y VDD 0.00fF
C56655 POR2X1_812/A POR2X1_800/O 0.00fF
C56656 INPUT_3 POR2X1_8/a_16_28# 0.03fF
C56657 PAND2X1_23/Y POR2X1_444/a_16_28# 0.03fF
C56658 D_INPUT_5 POR2X1_638/O 0.17fF
C56659 POR2X1_135/Y D_INPUT_0 1.94fF
C56660 POR2X1_838/a_16_28# POR2X1_837/Y 0.03fF
C56661 POR2X1_753/Y POR2X1_625/CTRL 0.05fF
C56662 PAND2X1_792/B VDD 0.10fF
C56663 POR2X1_673/A D_INPUT_0 1.79fF
C56664 POR2X1_416/B PAND2X1_346/CTRL2 0.03fF
C56665 POR2X1_696/Y POR2X1_32/A 0.01fF
C56666 POR2X1_66/B POR2X1_128/A 0.01fF
C56667 PAND2X1_601/CTRL2 POR2X1_294/B 0.02fF
C56668 POR2X1_496/Y POR2X1_511/Y 0.08fF
C56669 POR2X1_32/A PAND2X1_596/CTRL 0.08fF
C56670 PAND2X1_658/a_76_28# POR2X1_60/A 0.02fF
C56671 POR2X1_78/A POR2X1_830/A 0.01fF
C56672 POR2X1_448/A POR2X1_296/B 0.04fF
C56673 POR2X1_864/A PAND2X1_32/B 0.18fF
C56674 INPUT_3 POR2X1_380/CTRL2 0.04fF
C56675 POR2X1_10/CTRL POR2X1_9/Y 0.01fF
C56676 POR2X1_709/A PAND2X1_6/A 0.01fF
C56677 PAND2X1_815/O POR2X1_14/Y 0.06fF
C56678 PAND2X1_65/B POR2X1_634/A 0.08fF
C56679 PAND2X1_463/CTRL2 POR2X1_5/Y 0.03fF
C56680 POR2X1_260/B POR2X1_715/a_16_28# 0.03fF
C56681 POR2X1_322/CTRL POR2X1_23/Y 0.01fF
C56682 POR2X1_429/O INPUT_7 0.05fF
C56683 POR2X1_604/Y VDD 0.01fF
C56684 POR2X1_57/A POR2X1_20/B 13.47fF
C56685 PAND2X1_413/O PAND2X1_57/B 0.05fF
C56686 POR2X1_150/Y POR2X1_91/Y 0.14fF
C56687 POR2X1_471/O POR2X1_78/A 0.01fF
C56688 POR2X1_60/A PAND2X1_347/Y 0.03fF
C56689 POR2X1_241/O VDD 0.00fF
C56690 POR2X1_399/CTRL PAND2X1_403/B 0.03fF
C56691 PAND2X1_63/Y POR2X1_624/Y 0.03fF
C56692 POR2X1_856/m4_208_n4# POR2X1_782/m4_208_n4# 0.13fF
C56693 POR2X1_188/A POR2X1_733/CTRL2 0.01fF
C56694 POR2X1_830/a_16_28# POR2X1_830/A 0.02fF
C56695 POR2X1_475/A POR2X1_734/A 0.13fF
C56696 POR2X1_221/CTRL2 POR2X1_186/Y 0.01fF
C56697 PAND2X1_217/B PAND2X1_558/CTRL 0.27fF
C56698 POR2X1_66/B POR2X1_206/A 0.02fF
C56699 POR2X1_67/A POR2X1_754/A 0.00fF
C56700 PAND2X1_23/Y POR2X1_218/Y 0.07fF
C56701 POR2X1_13/A POR2X1_14/Y 0.05fF
C56702 PAND2X1_790/CTRL POR2X1_93/A 0.01fF
C56703 POR2X1_43/B POR2X1_420/CTRL2 0.03fF
C56704 PAND2X1_93/CTRL2 POR2X1_66/A 0.01fF
C56705 POR2X1_141/Y POR2X1_217/O 0.04fF
C56706 PAND2X1_612/B POR2X1_68/B 0.01fF
C56707 PAND2X1_260/CTRL VDD 0.00fF
C56708 POR2X1_49/Y POR2X1_236/Y 0.18fF
C56709 POR2X1_254/Y POR2X1_254/A 0.01fF
C56710 PAND2X1_402/a_16_344# POR2X1_397/Y 0.01fF
C56711 PAND2X1_57/CTRL2 PAND2X1_41/B 0.01fF
C56712 POR2X1_490/Y POR2X1_73/Y 0.06fF
C56713 POR2X1_516/O POR2X1_48/A 0.04fF
C56714 POR2X1_556/A POR2X1_787/CTRL2 0.03fF
C56715 POR2X1_130/A POR2X1_777/B 0.10fF
C56716 POR2X1_481/A POR2X1_312/Y 0.00fF
C56717 POR2X1_254/Y POR2X1_750/B 0.10fF
C56718 PAND2X1_20/A PAND2X1_89/O 0.17fF
C56719 PAND2X1_620/Y VDD 0.15fF
C56720 POR2X1_669/B PAND2X1_546/Y 0.08fF
C56721 POR2X1_250/CTRL POR2X1_250/A 0.06fF
C56722 PAND2X1_659/A PAND2X1_659/B 1.15fF
C56723 INPUT_7 POR2X1_2/O 0.01fF
C56724 POR2X1_270/Y PAND2X1_96/B 0.03fF
C56725 POR2X1_65/A VDD 4.59fF
C56726 POR2X1_311/Y POR2X1_488/Y 0.02fF
C56727 D_INPUT_0 POR2X1_816/A 0.03fF
C56728 POR2X1_72/CTRL PAND2X1_659/B 0.00fF
C56729 POR2X1_120/CTRL PAND2X1_90/Y 0.03fF
C56730 POR2X1_411/Y POR2X1_607/A 0.02fF
C56731 POR2X1_814/B POR2X1_544/A 0.01fF
C56732 D_INPUT_0 D_INPUT_1 8.37fF
C56733 POR2X1_615/CTRL2 POR2X1_754/A 0.01fF
C56734 POR2X1_149/B POR2X1_296/B 0.06fF
C56735 PAND2X1_57/B POR2X1_543/A 0.03fF
C56736 POR2X1_254/Y PAND2X1_13/O 0.05fF
C56737 PAND2X1_340/O INPUT_0 0.04fF
C56738 POR2X1_362/B VDD 0.38fF
C56739 POR2X1_525/CTRL2 POR2X1_41/B 0.01fF
C56740 POR2X1_693/Y POR2X1_83/B 0.02fF
C56741 POR2X1_130/A PAND2X1_65/B 0.10fF
C56742 POR2X1_631/O POR2X1_294/B 0.02fF
C56743 POR2X1_866/A POR2X1_780/B 0.10fF
C56744 POR2X1_47/O POR2X1_748/A 0.01fF
C56745 POR2X1_123/A POR2X1_260/B 0.06fF
C56746 PAND2X1_445/Y PAND2X1_76/Y 0.03fF
C56747 PAND2X1_621/O POR2X1_415/A 0.12fF
C56748 POR2X1_566/A PAND2X1_65/B 0.11fF
C56749 PAND2X1_58/A PAND2X1_6/A 0.07fF
C56750 POR2X1_523/Y POR2X1_819/a_16_28# 0.02fF
C56751 PAND2X1_434/a_16_344# POR2X1_172/Y 0.01fF
C56752 POR2X1_443/A POR2X1_545/O 0.00fF
C56753 POR2X1_327/Y POR2X1_499/A 0.03fF
C56754 POR2X1_372/A POR2X1_372/a_16_28# 0.03fF
C56755 POR2X1_260/B PAND2X1_765/O 0.02fF
C56756 POR2X1_78/B POR2X1_596/Y 0.04fF
C56757 POR2X1_66/B POR2X1_455/A 0.03fF
C56758 PAND2X1_20/A POR2X1_775/CTRL 0.01fF
C56759 POR2X1_54/Y PAND2X1_749/CTRL2 0.08fF
C56760 POR2X1_624/Y POR2X1_260/A 0.03fF
C56761 POR2X1_322/a_56_344# POR2X1_40/Y 0.00fF
C56762 PAND2X1_96/B POR2X1_288/O 0.01fF
C56763 POR2X1_146/m4_208_n4# POR2X1_257/A 0.07fF
C56764 PAND2X1_408/O PAND2X1_18/B 0.15fF
C56765 POR2X1_740/O POR2X1_738/Y 0.00fF
C56766 POR2X1_186/Y POR2X1_732/B 0.10fF
C56767 POR2X1_594/O POR2X1_594/A 0.02fF
C56768 PAND2X1_735/Y PAND2X1_501/B 0.02fF
C56769 POR2X1_61/Y POR2X1_205/Y 0.07fF
C56770 PAND2X1_562/B POR2X1_55/Y 0.08fF
C56771 PAND2X1_23/Y POR2X1_710/A 0.03fF
C56772 D_INPUT_3 POR2X1_32/A 0.03fF
C56773 POR2X1_271/A POR2X1_257/A 0.03fF
C56774 PAND2X1_55/Y POR2X1_61/Y 0.07fF
C56775 POR2X1_502/A PAND2X1_700/O 0.01fF
C56776 POR2X1_814/A POR2X1_330/O 0.33fF
C56777 POR2X1_646/Y POR2X1_307/A 0.04fF
C56778 POR2X1_23/Y POR2X1_521/Y 0.10fF
C56779 POR2X1_66/A PAND2X1_397/O 0.01fF
C56780 POR2X1_43/B PAND2X1_500/O 0.02fF
C56781 POR2X1_13/A PAND2X1_735/O 0.02fF
C56782 POR2X1_113/Y POR2X1_650/CTRL 0.01fF
C56783 POR2X1_481/a_16_28# POR2X1_481/A 0.03fF
C56784 POR2X1_66/A POR2X1_796/A 0.03fF
C56785 POR2X1_332/B PAND2X1_57/B 0.03fF
C56786 PAND2X1_137/Y PAND2X1_768/CTRL2 0.01fF
C56787 PAND2X1_454/O POR2X1_511/Y 0.09fF
C56788 POR2X1_445/A POR2X1_186/B 0.03fF
C56789 PAND2X1_473/B POR2X1_42/Y 0.05fF
C56790 POR2X1_623/A POR2X1_623/a_16_28# 0.06fF
C56791 POR2X1_283/A POR2X1_29/A 0.03fF
C56792 POR2X1_499/CTRL POR2X1_456/B 0.01fF
C56793 POR2X1_66/B POR2X1_140/O 0.01fF
C56794 POR2X1_96/A POR2X1_625/Y 0.00fF
C56795 POR2X1_327/Y POR2X1_76/A 0.03fF
C56796 PAND2X1_216/B POR2X1_23/Y 0.03fF
C56797 POR2X1_254/A POR2X1_341/Y 0.12fF
C56798 POR2X1_397/Y POR2X1_42/Y 0.26fF
C56799 POR2X1_423/Y POR2X1_90/Y 0.00fF
C56800 PAND2X1_824/B POR2X1_630/CTRL2 0.04fF
C56801 POR2X1_296/B POR2X1_274/B 0.04fF
C56802 PAND2X1_635/CTRL2 POR2X1_763/A 0.01fF
C56803 POR2X1_96/A PAND2X1_191/CTRL2 0.01fF
C56804 PAND2X1_833/CTRL PAND2X1_658/B -0.00fF
C56805 PAND2X1_93/B POR2X1_449/A 0.03fF
C56806 POR2X1_97/A PAND2X1_503/CTRL2 0.04fF
C56807 POR2X1_65/A POR2X1_93/CTRL 0.01fF
C56808 POR2X1_41/B PAND2X1_515/O 0.02fF
C56809 POR2X1_52/A PAND2X1_471/B 0.01fF
C56810 PAND2X1_56/Y POR2X1_308/O 0.29fF
C56811 PAND2X1_679/CTRL PAND2X1_69/A 0.01fF
C56812 POR2X1_777/B PAND2X1_150/O 0.01fF
C56813 POR2X1_13/A POR2X1_55/Y 0.17fF
C56814 POR2X1_78/B POR2X1_538/O 0.02fF
C56815 PAND2X1_850/Y POR2X1_411/B 0.07fF
C56816 POR2X1_462/B PAND2X1_90/Y 0.03fF
C56817 PAND2X1_391/CTRL2 POR2X1_751/Y 0.01fF
C56818 POR2X1_121/B PAND2X1_300/CTRL 0.01fF
C56819 POR2X1_192/Y POR2X1_221/Y 0.04fF
C56820 PAND2X1_190/Y VDD 1.36fF
C56821 PAND2X1_48/B PAND2X1_386/Y 0.90fF
C56822 PAND2X1_57/B POR2X1_363/CTRL 0.01fF
C56823 POR2X1_78/B PAND2X1_6/Y 0.16fF
C56824 POR2X1_362/B PAND2X1_32/B 0.06fF
C56825 PAND2X1_206/O PAND2X1_6/A 0.06fF
C56826 POR2X1_61/a_16_28# POR2X1_66/A 0.03fF
C56827 POR2X1_302/a_16_28# POR2X1_302/A 0.03fF
C56828 PAND2X1_41/B PAND2X1_60/B 6.80fF
C56829 POR2X1_706/O INPUT_1 0.01fF
C56830 POR2X1_44/O INPUT_6 0.01fF
C56831 PAND2X1_96/a_76_28# PAND2X1_94/Y 0.07fF
C56832 POR2X1_136/CTRL VDD 0.00fF
C56833 PAND2X1_724/B POR2X1_293/Y 0.01fF
C56834 PAND2X1_565/O VDD 0.00fF
C56835 POR2X1_840/B POR2X1_217/CTRL 0.13fF
C56836 POR2X1_102/Y POR2X1_172/a_76_344# 0.00fF
C56837 POR2X1_713/A POR2X1_532/A 0.02fF
C56838 PAND2X1_41/B POR2X1_758/a_16_28# 0.02fF
C56839 POR2X1_664/a_76_344# POR2X1_78/A 0.00fF
C56840 POR2X1_78/A POR2X1_703/Y 0.03fF
C56841 PAND2X1_821/CTRL2 PAND2X1_23/Y 0.04fF
C56842 POR2X1_496/Y POR2X1_129/Y 0.07fF
C56843 PAND2X1_859/CTRL2 POR2X1_283/A 0.00fF
C56844 POR2X1_471/CTRL2 POR2X1_540/A 0.01fF
C56845 POR2X1_830/A PAND2X1_306/O 0.02fF
C56846 POR2X1_25/O D_INPUT_6 0.01fF
C56847 POR2X1_66/B INPUT_1 0.03fF
C56848 POR2X1_132/Y VDD 0.00fF
C56849 PAND2X1_48/B POR2X1_415/Y 0.02fF
C56850 VDD PAND2X1_359/B 0.11fF
C56851 POR2X1_529/O POR2X1_55/Y 0.07fF
C56852 PAND2X1_793/Y POR2X1_56/Y 0.03fF
C56853 POR2X1_376/B PAND2X1_374/CTRL2 0.00fF
C56854 PAND2X1_63/Y POR2X1_786/m4_208_n4# 0.08fF
C56855 POR2X1_781/B POR2X1_568/Y 0.31fF
C56856 POR2X1_16/A POR2X1_39/CTRL2 0.01fF
C56857 PAND2X1_48/B POR2X1_140/B 0.03fF
C56858 POR2X1_205/Y POR2X1_35/Y 0.03fF
C56859 PAND2X1_254/a_16_344# PAND2X1_658/B -0.00fF
C56860 POR2X1_188/A INPUT_1 0.03fF
C56861 PAND2X1_223/B PAND2X1_538/O 0.02fF
C56862 POR2X1_43/B PAND2X1_478/CTRL2 0.03fF
C56863 PAND2X1_55/Y POR2X1_35/Y 0.03fF
C56864 PAND2X1_48/B POR2X1_407/A 0.06fF
C56865 PAND2X1_23/Y POR2X1_68/A 0.20fF
C56866 POR2X1_16/A PAND2X1_240/CTRL 0.02fF
C56867 POR2X1_383/A PAND2X1_759/a_76_28# 0.02fF
C56868 POR2X1_455/a_56_344# POR2X1_222/A 0.00fF
C56869 POR2X1_402/B PAND2X1_60/B 0.00fF
C56870 VDD POR2X1_161/Y -0.00fF
C56871 POR2X1_60/A PAND2X1_123/Y 0.08fF
C56872 PAND2X1_341/A PAND2X1_364/B 0.05fF
C56873 PAND2X1_41/B POR2X1_353/A 0.02fF
C56874 PAND2X1_243/B POR2X1_73/Y 0.07fF
C56875 POR2X1_68/B POR2X1_404/Y 0.03fF
C56876 D_INPUT_3 PAND2X1_35/Y 0.05fF
C56877 POR2X1_83/Y POR2X1_32/A 0.02fF
C56878 POR2X1_192/Y POR2X1_714/O 0.07fF
C56879 POR2X1_177/CTRL2 POR2X1_72/B 0.01fF
C56880 PAND2X1_631/A POR2X1_56/CTRL2 0.01fF
C56881 POR2X1_805/A POR2X1_710/CTRL 0.00fF
C56882 PAND2X1_170/CTRL PAND2X1_169/Y 0.01fF
C56883 INPUT_7 POR2X1_260/A 0.03fF
C56884 PAND2X1_6/Y PAND2X1_7/O 0.17fF
C56885 POR2X1_596/A PAND2X1_604/CTRL2 0.01fF
C56886 INPUT_1 POR2X1_376/Y 0.01fF
C56887 POR2X1_32/A POR2X1_371/a_16_28# 0.04fF
C56888 POR2X1_356/A PAND2X1_747/O 0.10fF
C56889 POR2X1_538/A PAND2X1_57/B 0.01fF
C56890 PAND2X1_844/CTRL PAND2X1_61/Y 0.01fF
C56891 PAND2X1_341/A PAND2X1_101/O 0.03fF
C56892 POR2X1_408/Y INPUT_5 0.01fF
C56893 POR2X1_404/B PAND2X1_397/a_16_344# 0.02fF
C56894 PAND2X1_20/A PAND2X1_396/CTRL 0.01fF
C56895 POR2X1_7/B PAND2X1_348/Y 1.30fF
C56896 POR2X1_579/Y PAND2X1_173/O 0.00fF
C56897 POR2X1_297/CTRL PAND2X1_359/Y 0.01fF
C56898 PAND2X1_722/CTRL2 POR2X1_666/A 0.00fF
C56899 POR2X1_38/Y POR2X1_599/A 0.05fF
C56900 POR2X1_344/Y PAND2X1_65/B 0.01fF
C56901 POR2X1_60/O PAND2X1_339/Y 0.16fF
C56902 INPUT_6 POR2X1_587/CTRL 0.01fF
C56903 POR2X1_239/m4_208_n4# POR2X1_55/Y 0.09fF
C56904 PAND2X1_472/CTRL PAND2X1_673/Y 0.04fF
C56905 PAND2X1_276/CTRL POR2X1_129/Y 0.01fF
C56906 POR2X1_97/B POR2X1_186/Y 0.05fF
C56907 PAND2X1_488/O POR2X1_294/A 0.03fF
C56908 POR2X1_740/Y POR2X1_319/Y 0.03fF
C56909 POR2X1_597/A POR2X1_597/a_16_28# 0.03fF
C56910 POR2X1_130/Y PAND2X1_60/B 1.19fF
C56911 PAND2X1_29/a_16_344# POR2X1_68/B 0.01fF
C56912 PAND2X1_741/B PAND2X1_557/O 0.02fF
C56913 POR2X1_55/Y POR2X1_9/m4_208_n4# 0.03fF
C56914 POR2X1_66/B PAND2X1_136/CTRL 0.01fF
C56915 PAND2X1_850/Y POR2X1_271/Y 0.15fF
C56916 POR2X1_435/Y PAND2X1_533/CTRL 0.06fF
C56917 INPUT_4 POR2X1_260/A 0.36fF
C56918 POR2X1_856/B POR2X1_181/Y 0.02fF
C56919 POR2X1_198/CTRL2 POR2X1_215/A 0.02fF
C56920 POR2X1_491/Y POR2X1_60/A 0.00fF
C56921 POR2X1_334/A VDD 0.11fF
C56922 POR2X1_51/B POR2X1_587/CTRL2 0.01fF
C56923 PAND2X1_319/B POR2X1_90/Y 0.12fF
C56924 POR2X1_219/B PAND2X1_88/Y 0.00fF
C56925 POR2X1_96/A POR2X1_419/a_76_344# 0.01fF
C56926 POR2X1_176/a_16_28# POR2X1_312/Y 0.02fF
C56927 POR2X1_795/B POR2X1_854/B 0.05fF
C56928 POR2X1_102/Y POR2X1_533/Y 0.14fF
C56929 PAND2X1_209/A POR2X1_152/Y 0.00fF
C56930 POR2X1_193/A POR2X1_456/B 0.03fF
C56931 PAND2X1_72/CTRL PAND2X1_60/B 0.00fF
C56932 POR2X1_579/Y POR2X1_456/B 0.01fF
C56933 PAND2X1_63/Y POR2X1_493/CTRL 0.01fF
C56934 POR2X1_844/a_76_344# D_INPUT_1 0.01fF
C56935 PAND2X1_48/O POR2X1_186/B 0.02fF
C56936 D_INPUT_1 POR2X1_361/O 0.02fF
C56937 POR2X1_78/B POR2X1_195/O 0.02fF
C56938 POR2X1_741/Y POR2X1_553/A 0.03fF
C56939 POR2X1_785/A POR2X1_260/A 0.08fF
C56940 PAND2X1_816/O POR2X1_260/A 0.02fF
C56941 PAND2X1_550/Y PAND2X1_565/A 0.00fF
C56942 PAND2X1_264/O POR2X1_519/Y 0.00fF
C56943 PAND2X1_65/B PAND2X1_167/CTRL 0.01fF
C56944 POR2X1_110/Y POR2X1_368/CTRL 0.01fF
C56945 D_GATE_222 POR2X1_175/B 0.02fF
C56946 PAND2X1_6/Y POR2X1_141/A 0.01fF
C56947 PAND2X1_723/A POR2X1_52/Y 0.01fF
C56948 PAND2X1_857/A POR2X1_73/Y 0.03fF
C56949 POR2X1_16/A POR2X1_43/B 0.34fF
C56950 POR2X1_41/B PAND2X1_156/A 0.10fF
C56951 POR2X1_13/A PAND2X1_199/B 0.01fF
C56952 POR2X1_740/Y POR2X1_507/A 0.10fF
C56953 PAND2X1_785/Y PAND2X1_716/B 0.10fF
C56954 POR2X1_57/A PAND2X1_121/CTRL2 0.03fF
C56955 POR2X1_505/CTRL PAND2X1_6/A 0.03fF
C56956 PAND2X1_57/B POR2X1_342/O 0.01fF
C56957 POR2X1_334/Y POR2X1_193/CTRL2 0.03fF
C56958 POR2X1_553/A PAND2X1_32/B 0.56fF
C56959 POR2X1_327/Y PAND2X1_604/O 0.17fF
C56960 POR2X1_407/Y PAND2X1_765/O 0.02fF
C56961 PAND2X1_60/B POR2X1_228/Y 0.29fF
C56962 PAND2X1_96/B POR2X1_101/Y 0.09fF
C56963 POR2X1_614/A POR2X1_456/B 0.03fF
C56964 POR2X1_264/Y POR2X1_559/A 0.03fF
C56965 POR2X1_532/A POR2X1_796/A 0.03fF
C56966 POR2X1_609/Y POR2X1_234/A 0.03fF
C56967 POR2X1_38/Y POR2X1_235/a_16_28# 0.06fF
C56968 POR2X1_87/CTRL2 PAND2X1_41/B 0.01fF
C56969 PAND2X1_625/m4_208_n4# POR2X1_260/A 0.09fF
C56970 POR2X1_539/A POR2X1_188/CTRL 0.00fF
C56971 PAND2X1_849/B PAND2X1_341/A 0.03fF
C56972 POR2X1_83/Y PAND2X1_35/Y 0.03fF
C56973 POR2X1_68/B POR2X1_773/CTRL 0.01fF
C56974 POR2X1_278/Y PAND2X1_865/Y 0.07fF
C56975 POR2X1_78/B PAND2X1_290/CTRL2 0.02fF
C56976 PAND2X1_651/Y PAND2X1_510/O 0.14fF
C56977 PAND2X1_218/O PAND2X1_853/B 0.04fF
C56978 POR2X1_216/CTRL2 POR2X1_101/Y 0.09fF
C56979 POR2X1_280/O POR2X1_280/Y 0.01fF
C56980 POR2X1_333/Y POR2X1_35/Y 0.03fF
C56981 POR2X1_557/A POR2X1_68/B 0.06fF
C56982 PAND2X1_42/a_56_28# POR2X1_590/A 0.00fF
C56983 PAND2X1_6/Y PAND2X1_142/CTRL2 0.00fF
C56984 POR2X1_416/B PAND2X1_192/Y 0.05fF
C56985 PAND2X1_476/A POR2X1_7/B 0.01fF
C56986 PAND2X1_467/Y PAND2X1_470/A 0.13fF
C56987 POR2X1_809/A POR2X1_68/A 0.00fF
C56988 PAND2X1_283/CTRL2 POR2X1_294/A 0.17fF
C56989 VDD D_INPUT_4 0.39fF
C56990 POR2X1_7/B PAND2X1_539/O 0.04fF
C56991 POR2X1_68/B POR2X1_571/CTRL 0.00fF
C56992 PAND2X1_417/a_16_344# POR2X1_663/B 0.03fF
C56993 POR2X1_283/A PAND2X1_130/a_16_344# 0.01fF
C56994 POR2X1_493/CTRL POR2X1_260/A 0.01fF
C56995 PAND2X1_106/CTRL POR2X1_276/Y 0.01fF
C56996 POR2X1_461/Y POR2X1_859/CTRL 0.01fF
C56997 PAND2X1_382/CTRL2 POR2X1_260/A 0.03fF
C56998 PAND2X1_94/A PAND2X1_27/CTRL 0.00fF
C56999 POR2X1_356/A POR2X1_726/a_16_28# 0.04fF
C57000 PAND2X1_23/Y POR2X1_112/O 0.02fF
C57001 PAND2X1_661/Y PAND2X1_121/a_16_344# 0.02fF
C57002 POR2X1_118/a_76_344# PAND2X1_560/B 0.01fF
C57003 PAND2X1_6/Y POR2X1_294/A 1.96fF
C57004 POR2X1_814/A PAND2X1_65/CTRL 0.30fF
C57005 POR2X1_78/B POR2X1_500/CTRL 0.00fF
C57006 PAND2X1_294/CTRL2 POR2X1_411/B 0.01fF
C57007 POR2X1_542/Y POR2X1_732/B 0.14fF
C57008 POR2X1_416/B PAND2X1_738/Y 0.03fF
C57009 PAND2X1_824/B POR2X1_510/Y 0.02fF
C57010 POR2X1_78/B PAND2X1_52/B 1.07fF
C57011 POR2X1_840/B POR2X1_737/A 0.05fF
C57012 PAND2X1_661/B PAND2X1_199/B 0.01fF
C57013 POR2X1_416/B POR2X1_425/CTRL 0.01fF
C57014 POR2X1_293/Y PAND2X1_358/O 0.03fF
C57015 POR2X1_559/Y POR2X1_560/a_56_344# 0.00fF
C57016 PAND2X1_38/CTRL2 PAND2X1_52/B 0.34fF
C57017 PAND2X1_96/B PAND2X1_323/CTRL2 0.05fF
C57018 POR2X1_327/Y POR2X1_539/A 0.01fF
C57019 POR2X1_566/A PAND2X1_292/O 0.20fF
C57020 PAND2X1_198/O PAND2X1_197/Y 0.02fF
C57021 POR2X1_209/A POR2X1_726/O 0.01fF
C57022 POR2X1_1/CTRL2 PAND2X1_18/B 0.04fF
C57023 POR2X1_83/Y PAND2X1_844/B 0.02fF
C57024 POR2X1_622/B POR2X1_29/A 0.02fF
C57025 PAND2X1_171/CTRL2 POR2X1_854/B 0.18fF
C57026 POR2X1_45/Y POR2X1_39/B 0.23fF
C57027 D_INPUT_7 POR2X1_750/B 0.01fF
C57028 POR2X1_54/Y POR2X1_77/a_56_344# 0.01fF
C57029 PAND2X1_716/B PAND2X1_656/A 0.00fF
C57030 POR2X1_713/B PAND2X1_692/O 0.17fF
C57031 POR2X1_326/A POR2X1_737/CTRL2 0.07fF
C57032 POR2X1_569/A PAND2X1_48/A 0.07fF
C57033 POR2X1_784/A POR2X1_717/B 0.03fF
C57034 POR2X1_634/A POR2X1_814/A 0.02fF
C57035 POR2X1_68/A POR2X1_711/Y 0.10fF
C57036 POR2X1_78/B PAND2X1_125/a_16_344# 0.03fF
C57037 POR2X1_305/O POR2X1_305/Y 0.01fF
C57038 INPUT_1 PAND2X1_358/A 0.03fF
C57039 PAND2X1_439/CTRL2 POR2X1_72/B 0.03fF
C57040 POR2X1_186/B POR2X1_260/A 0.04fF
C57041 POR2X1_858/A POR2X1_840/B 0.03fF
C57042 POR2X1_69/O PAND2X1_206/B 0.00fF
C57043 PAND2X1_62/CTRL POR2X1_9/Y 0.01fF
C57044 POR2X1_411/B PAND2X1_722/CTRL 0.01fF
C57045 PAND2X1_32/B D_INPUT_4 0.03fF
C57046 INPUT_3 D_INPUT_0 0.14fF
C57047 POR2X1_814/A POR2X1_489/CTRL2 0.01fF
C57048 PAND2X1_854/A PAND2X1_643/A 0.02fF
C57049 POR2X1_376/B PAND2X1_99/O 0.02fF
C57050 POR2X1_270/Y POR2X1_222/CTRL 0.01fF
C57051 POR2X1_68/A POR2X1_728/A 0.00fF
C57052 POR2X1_67/Y PAND2X1_225/m4_208_n4# 0.15fF
C57053 POR2X1_832/Y POR2X1_841/B 0.07fF
C57054 POR2X1_316/Y PAND2X1_787/A 0.35fF
C57055 PAND2X1_665/O PAND2X1_60/B 0.02fF
C57056 POR2X1_63/Y POR2X1_669/B 0.01fF
C57057 POR2X1_863/A POR2X1_802/B 0.03fF
C57058 POR2X1_243/B POR2X1_66/A 0.01fF
C57059 POR2X1_97/A POR2X1_212/A 0.03fF
C57060 PAND2X1_104/a_16_344# POR2X1_624/B 0.04fF
C57061 POR2X1_567/B POR2X1_434/O 0.02fF
C57062 POR2X1_624/B POR2X1_94/A 0.12fF
C57063 POR2X1_462/CTRL POR2X1_734/A 0.04fF
C57064 POR2X1_432/a_16_28# POR2X1_271/B 0.04fF
C57065 POR2X1_396/Y POR2X1_39/B 0.01fF
C57066 POR2X1_329/A POR2X1_237/CTRL2 0.03fF
C57067 PAND2X1_348/A PAND2X1_716/B 0.01fF
C57068 POR2X1_346/A POR2X1_202/A 0.04fF
C57069 POR2X1_13/A PAND2X1_458/O 0.21fF
C57070 POR2X1_864/A POR2X1_808/A 0.03fF
C57071 POR2X1_815/a_16_28# POR2X1_750/A 0.01fF
C57072 POR2X1_564/B POR2X1_564/CTRL2 0.03fF
C57073 PAND2X1_48/B PAND2X1_628/CTRL2 0.01fF
C57074 PAND2X1_93/B D_INPUT_0 11.61fF
C57075 POR2X1_66/B PAND2X1_43/O 0.01fF
C57076 POR2X1_360/A PAND2X1_94/Y 0.44fF
C57077 POR2X1_416/B POR2X1_136/Y 0.03fF
C57078 POR2X1_9/Y PAND2X1_751/O 0.07fF
C57079 PAND2X1_458/CTRL POR2X1_293/Y 0.01fF
C57080 PAND2X1_602/a_76_28# POR2X1_600/Y 0.02fF
C57081 POR2X1_130/A POR2X1_814/A 0.16fF
C57082 POR2X1_329/A PAND2X1_579/B 0.02fF
C57083 PAND2X1_859/A POR2X1_411/B 0.05fF
C57084 POR2X1_57/A POR2X1_43/Y 0.04fF
C57085 POR2X1_294/A POR2X1_195/O 0.09fF
C57086 POR2X1_63/Y PAND2X1_231/CTRL 0.01fF
C57087 PAND2X1_96/B POR2X1_579/O 0.17fF
C57088 POR2X1_411/B PAND2X1_579/O 0.08fF
C57089 POR2X1_566/A POR2X1_814/A 0.13fF
C57090 POR2X1_158/Y PAND2X1_713/A 0.00fF
C57091 POR2X1_65/A PAND2X1_9/Y 0.03fF
C57092 POR2X1_54/Y PAND2X1_23/CTRL 0.05fF
C57093 POR2X1_137/B PAND2X1_90/Y 0.01fF
C57094 POR2X1_863/A POR2X1_532/A 0.03fF
C57095 PAND2X1_436/CTRL2 PAND2X1_390/Y 0.01fF
C57096 POR2X1_271/B PAND2X1_499/Y 0.03fF
C57097 POR2X1_63/Y POR2X1_230/O 0.01fF
C57098 POR2X1_424/Y PAND2X1_803/A 0.25fF
C57099 PAND2X1_631/A PAND2X1_716/B 0.07fF
C57100 POR2X1_602/A POR2X1_66/A 0.03fF
C57101 POR2X1_78/A D_INPUT_0 0.10fF
C57102 POR2X1_379/a_76_344# PAND2X1_52/B 0.03fF
C57103 POR2X1_567/B POR2X1_467/Y 0.43fF
C57104 PAND2X1_70/CTRL2 POR2X1_635/A 0.01fF
C57105 PAND2X1_86/a_76_28# PAND2X1_57/B 0.02fF
C57106 POR2X1_438/Y POR2X1_72/B 0.03fF
C57107 PAND2X1_340/B PAND2X1_340/O 0.05fF
C57108 PAND2X1_73/Y POR2X1_121/B 0.03fF
C57109 POR2X1_83/B PAND2X1_212/B 0.03fF
C57110 POR2X1_14/Y POR2X1_29/A 0.08fF
C57111 POR2X1_67/Y POR2X1_619/O 0.01fF
C57112 POR2X1_442/a_16_28# POR2X1_236/Y 0.03fF
C57113 POR2X1_96/A POR2X1_411/B 0.06fF
C57114 POR2X1_56/a_56_344# POR2X1_83/B 0.00fF
C57115 POR2X1_478/CTRL POR2X1_480/A 0.08fF
C57116 PAND2X1_156/A POR2X1_77/Y 0.03fF
C57117 POR2X1_49/Y POR2X1_626/CTRL 0.00fF
C57118 POR2X1_466/A POR2X1_186/Y 0.10fF
C57119 PAND2X1_234/a_16_344# PAND2X1_88/Y 0.00fF
C57120 PAND2X1_317/a_16_344# POR2X1_167/Y 0.01fF
C57121 POR2X1_456/CTRL POR2X1_66/A 0.00fF
C57122 POR2X1_857/A POR2X1_579/Y 0.01fF
C57123 POR2X1_411/B PAND2X1_335/O 0.03fF
C57124 POR2X1_373/CTRL POR2X1_77/Y 0.01fF
C57125 POR2X1_649/O POR2X1_294/B 0.02fF
C57126 POR2X1_838/B POR2X1_330/Y 0.03fF
C57127 POR2X1_129/Y PAND2X1_332/Y 0.03fF
C57128 POR2X1_329/A POR2X1_73/Y 0.17fF
C57129 PAND2X1_48/A POR2X1_725/O 0.02fF
C57130 POR2X1_32/A PAND2X1_733/O 0.02fF
C57131 POR2X1_397/Y PAND2X1_720/m4_208_n4# 0.15fF
C57132 POR2X1_48/A PAND2X1_62/a_16_344# 0.02fF
C57133 POR2X1_67/Y POR2X1_68/B 0.03fF
C57134 POR2X1_813/CTRL POR2X1_55/Y 0.13fF
C57135 POR2X1_814/A POR2X1_573/A 0.05fF
C57136 POR2X1_603/Y POR2X1_72/B 0.03fF
C57137 POR2X1_294/A PAND2X1_52/B 0.10fF
C57138 PAND2X1_645/Y VDD 0.00fF
C57139 PAND2X1_48/A PAND2X1_72/A 0.19fF
C57140 POR2X1_262/Y PAND2X1_716/CTRL2 0.02fF
C57141 POR2X1_287/B POR2X1_296/B 0.03fF
C57142 POR2X1_866/CTRL POR2X1_750/B 0.01fF
C57143 POR2X1_20/B POR2X1_396/CTRL 0.01fF
C57144 PAND2X1_48/B PAND2X1_271/O 0.04fF
C57145 POR2X1_32/A PAND2X1_778/CTRL2 0.01fF
C57146 PAND2X1_211/O POR2X1_55/Y 0.03fF
C57147 PAND2X1_61/Y POR2X1_83/B 0.03fF
C57148 PAND2X1_6/Y POR2X1_116/A 0.03fF
C57149 POR2X1_816/O POR2X1_816/A 0.05fF
C57150 POR2X1_498/CTRL PAND2X1_205/A 0.00fF
C57151 PAND2X1_88/CTRL2 PAND2X1_41/B 0.01fF
C57152 POR2X1_624/Y PAND2X1_110/O 0.02fF
C57153 PAND2X1_659/Y PAND2X1_332/Y 0.14fF
C57154 POR2X1_67/CTRL2 POR2X1_55/Y 0.24fF
C57155 PAND2X1_65/B POR2X1_241/B 0.04fF
C57156 POR2X1_856/B POR2X1_570/CTRL 0.01fF
C57157 POR2X1_41/B PAND2X1_444/a_16_344# 0.01fF
C57158 POR2X1_78/A PAND2X1_90/Y 2.71fF
C57159 POR2X1_556/A POR2X1_112/Y 0.03fF
C57160 POR2X1_607/A POR2X1_607/a_16_28# 0.09fF
C57161 PAND2X1_48/B POR2X1_632/CTRL 0.01fF
C57162 POR2X1_260/B POR2X1_795/O 0.18fF
C57163 POR2X1_850/A POR2X1_287/a_16_28# 0.07fF
C57164 POR2X1_49/Y PAND2X1_208/CTRL 0.02fF
C57165 POR2X1_750/B PAND2X1_41/B 0.19fF
C57166 POR2X1_335/A POR2X1_76/A 0.03fF
C57167 POR2X1_296/B PAND2X1_8/Y 0.12fF
C57168 POR2X1_67/O PAND2X1_658/A 0.01fF
C57169 POR2X1_257/A PAND2X1_785/CTRL2 0.05fF
C57170 POR2X1_48/CTRL POR2X1_60/A 0.01fF
C57171 PAND2X1_23/Y PAND2X1_827/CTRL2 0.01fF
C57172 POR2X1_68/A POR2X1_632/CTRL2 0.01fF
C57173 POR2X1_174/B VDD 1.61fF
C57174 POR2X1_651/O POR2X1_66/A 0.01fF
C57175 POR2X1_849/O POR2X1_94/A 0.03fF
C57176 PAND2X1_23/Y POR2X1_480/a_16_28# 0.03fF
C57177 POR2X1_750/B POR2X1_781/A 0.54fF
C57178 PAND2X1_58/A PAND2X1_58/a_16_344# 0.01fF
C57179 PAND2X1_55/a_16_344# POR2X1_94/A 0.02fF
C57180 POR2X1_411/Y D_INPUT_0 0.00fF
C57181 PAND2X1_859/A POR2X1_376/B 0.02fF
C57182 POR2X1_14/Y POR2X1_546/A 0.01fF
C57183 POR2X1_60/A PAND2X1_598/CTRL2 0.01fF
C57184 POR2X1_45/Y POR2X1_48/A 0.03fF
C57185 PAND2X1_784/CTRL2 POR2X1_32/A 0.01fF
C57186 POR2X1_496/Y POR2X1_293/Y 2.79fF
C57187 PAND2X1_423/CTRL2 POR2X1_480/A 0.02fF
C57188 PAND2X1_557/A PAND2X1_580/B 0.99fF
C57189 POR2X1_49/Y POR2X1_58/CTRL 0.01fF
C57190 POR2X1_411/B POR2X1_7/A 0.10fF
C57191 POR2X1_96/B POR2X1_20/B 0.02fF
C57192 POR2X1_344/Y POR2X1_814/A 0.14fF
C57193 POR2X1_29/A POR2X1_55/Y 0.13fF
C57194 POR2X1_864/A POR2X1_687/A 0.02fF
C57195 POR2X1_863/CTRL PAND2X1_73/Y 0.01fF
C57196 POR2X1_341/A POR2X1_366/A 0.07fF
C57197 POR2X1_555/B POR2X1_294/B 0.03fF
C57198 POR2X1_274/A POR2X1_532/A 0.03fF
C57199 PAND2X1_341/B POR2X1_9/Y 0.07fF
C57200 PAND2X1_793/Y PAND2X1_575/B 0.88fF
C57201 POR2X1_423/Y INPUT_0 0.09fF
C57202 POR2X1_295/CTRL2 POR2X1_7/B 0.00fF
C57203 PAND2X1_356/B VDD 0.11fF
C57204 POR2X1_344/O POR2X1_254/Y 0.00fF
C57205 PAND2X1_23/Y PAND2X1_58/A 0.19fF
C57206 POR2X1_73/a_56_344# POR2X1_20/B 0.00fF
C57207 POR2X1_257/A PAND2X1_434/CTRL2 0.00fF
C57208 PAND2X1_56/Y PAND2X1_73/Y 0.03fF
C57209 PAND2X1_631/CTRL2 POR2X1_669/B 0.01fF
C57210 PAND2X1_787/A POR2X1_298/O 0.03fF
C57211 POR2X1_566/A POR2X1_852/B 0.10fF
C57212 PAND2X1_49/CTRL POR2X1_29/A 0.01fF
C57213 POR2X1_555/A VDD 0.16fF
C57214 POR2X1_333/A POR2X1_740/Y 0.05fF
C57215 PAND2X1_192/Y PAND2X1_738/Y 0.05fF
C57216 PAND2X1_20/A POR2X1_563/Y 0.05fF
C57217 POR2X1_614/A POR2X1_450/CTRL 0.01fF
C57218 POR2X1_66/A PAND2X1_518/O 0.01fF
C57219 PAND2X1_816/a_16_344# POR2X1_634/A 0.01fF
C57220 POR2X1_490/Y PAND2X1_656/A 0.02fF
C57221 POR2X1_387/CTRL2 POR2X1_386/Y 0.00fF
C57222 POR2X1_122/Y VDD 0.07fF
C57223 POR2X1_830/O POR2X1_740/Y 0.10fF
C57224 POR2X1_830/CTRL2 POR2X1_741/Y 0.00fF
C57225 POR2X1_137/Y POR2X1_558/B 2.11fF
C57226 POR2X1_669/A POR2X1_83/B 0.01fF
C57227 POR2X1_52/A PAND2X1_859/A 0.06fF
C57228 POR2X1_383/A POR2X1_862/A 0.03fF
C57229 PAND2X1_21/CTRL VDD 0.00fF
C57230 POR2X1_330/Y POR2X1_294/B 0.16fF
C57231 POR2X1_366/Y POR2X1_330/Y 0.05fF
C57232 POR2X1_49/Y PAND2X1_523/CTRL 0.01fF
C57233 POR2X1_495/Y POR2X1_482/Y 0.23fF
C57234 POR2X1_389/CTRL2 POR2X1_389/Y 0.01fF
C57235 POR2X1_525/CTRL POR2X1_46/Y 0.01fF
C57236 POR2X1_459/a_16_28# POR2X1_750/B 0.02fF
C57237 POR2X1_96/A POR2X1_376/B 0.06fF
C57238 POR2X1_502/A POR2X1_663/CTRL2 0.01fF
C57239 POR2X1_626/O POR2X1_93/A 0.14fF
C57240 PAND2X1_39/B POR2X1_675/Y 0.00fF
C57241 POR2X1_355/B POR2X1_213/B 0.01fF
C57242 POR2X1_475/A PAND2X1_372/O 0.04fF
C57243 PAND2X1_267/Y PAND2X1_717/Y 0.03fF
C57244 POR2X1_13/A POR2X1_511/Y 0.03fF
C57245 POR2X1_114/B PAND2X1_279/O 0.06fF
C57246 PAND2X1_787/Y PAND2X1_592/O 0.15fF
C57247 POR2X1_65/A PAND2X1_714/O 0.01fF
C57248 PAND2X1_214/A POR2X1_599/A 0.02fF
C57249 POR2X1_590/A POR2X1_206/CTRL2 0.00fF
C57250 POR2X1_480/A POR2X1_220/Y 0.07fF
C57251 POR2X1_763/Y PAND2X1_738/CTRL 0.08fF
C57252 PAND2X1_650/O D_INPUT_0 0.05fF
C57253 POR2X1_174/B PAND2X1_32/B 0.30fF
C57254 POR2X1_661/B POR2X1_653/B 0.59fF
C57255 POR2X1_544/A VDD -0.00fF
C57256 POR2X1_590/A POR2X1_784/O 0.02fF
C57257 POR2X1_221/a_16_28# POR2X1_192/Y 0.06fF
C57258 POR2X1_65/A POR2X1_424/m4_208_n4# 0.08fF
C57259 POR2X1_66/B PAND2X1_491/CTRL 0.00fF
C57260 PAND2X1_90/Y PAND2X1_132/CTRL 0.01fF
C57261 POR2X1_108/CTRL2 POR2X1_102/Y 0.01fF
C57262 POR2X1_814/A POR2X1_342/m4_208_n4# 0.06fF
C57263 POR2X1_602/A POR2X1_532/A 0.06fF
C57264 POR2X1_121/A POR2X1_654/O 0.13fF
C57265 POR2X1_114/CTRL2 POR2X1_777/B 0.15fF
C57266 POR2X1_433/Y POR2X1_72/B 0.07fF
C57267 POR2X1_463/Y POR2X1_260/B 0.03fF
C57268 PAND2X1_67/O POR2X1_507/A 0.04fF
C57269 POR2X1_661/O POR2X1_740/Y 0.00fF
C57270 POR2X1_347/A POR2X1_202/A 0.02fF
C57271 POR2X1_496/Y POR2X1_408/Y 0.10fF
C57272 POR2X1_514/O POR2X1_777/B 0.04fF
C57273 PAND2X1_6/Y POR2X1_94/A 0.03fF
C57274 POR2X1_49/Y POR2X1_617/a_16_28# 0.03fF
C57275 POR2X1_855/B POR2X1_855/a_16_28# -0.00fF
C57276 D_GATE_222 PAND2X1_52/Y 0.03fF
C57277 PAND2X1_382/CTRL POR2X1_29/A 0.01fF
C57278 INPUT_2 POR2X1_609/CTRL 0.01fF
C57279 POR2X1_267/O POR2X1_318/A 0.03fF
C57280 PAND2X1_225/O POR2X1_68/B 0.04fF
C57281 POR2X1_14/Y POR2X1_583/O 0.18fF
C57282 POR2X1_174/CTRL POR2X1_567/B 0.01fF
C57283 POR2X1_348/A PAND2X1_6/Y 0.01fF
C57284 POR2X1_383/A PAND2X1_73/Y 0.13fF
C57285 POR2X1_244/B POR2X1_776/B 0.05fF
C57286 PAND2X1_827/a_16_344# POR2X1_260/A 0.02fF
C57287 POR2X1_243/Y POR2X1_404/Y 0.07fF
C57288 POR2X1_366/a_16_28# PAND2X1_93/B 0.02fF
C57289 POR2X1_52/A POR2X1_96/A 0.18fF
C57290 PAND2X1_20/A PAND2X1_505/a_56_28# 0.00fF
C57291 POR2X1_436/O POR2X1_209/A 0.01fF
C57292 PAND2X1_57/B POR2X1_193/A 0.08fF
C57293 PAND2X1_57/B POR2X1_579/Y 0.03fF
C57294 PAND2X1_420/O POR2X1_510/Y 0.02fF
C57295 POR2X1_60/Y PAND2X1_844/B 0.02fF
C57296 PAND2X1_61/Y POR2X1_522/Y 0.03fF
C57297 PAND2X1_41/B PAND2X1_177/CTRL 0.01fF
C57298 POR2X1_65/A PAND2X1_852/B 0.04fF
C57299 POR2X1_659/CTRL VDD -0.00fF
C57300 POR2X1_388/CTRL PAND2X1_65/B 0.11fF
C57301 POR2X1_71/Y PAND2X1_793/Y 0.00fF
C57302 POR2X1_686/O POR2X1_750/B 0.02fF
C57303 POR2X1_254/A POR2X1_228/Y 0.01fF
C57304 POR2X1_330/Y PAND2X1_111/B 0.03fF
C57305 D_INPUT_3 POR2X1_94/A 0.03fF
C57306 POR2X1_713/A POR2X1_713/a_16_28# 0.11fF
C57307 POR2X1_49/Y POR2X1_619/Y 0.03fF
C57308 PAND2X1_592/CTRL POR2X1_42/Y 0.01fF
C57309 PAND2X1_222/CTRL PAND2X1_643/A 0.01fF
C57310 POR2X1_603/CTRL POR2X1_761/A 0.01fF
C57311 POR2X1_54/Y POR2X1_4/Y 0.23fF
C57312 POR2X1_750/B POR2X1_228/Y 0.10fF
C57313 POR2X1_515/O POR2X1_515/Y 0.00fF
C57314 POR2X1_753/Y POR2X1_260/A 0.07fF
C57315 POR2X1_853/A POR2X1_502/A 0.10fF
C57316 POR2X1_376/B POR2X1_386/O 0.18fF
C57317 PAND2X1_793/Y POR2X1_42/Y 0.03fF
C57318 POR2X1_775/CTRL VDD 0.00fF
C57319 POR2X1_57/A INPUT_7 0.01fF
C57320 PAND2X1_738/B PAND2X1_731/A 0.18fF
C57321 PAND2X1_90/A POR2X1_404/Y 0.03fF
C57322 POR2X1_65/A POR2X1_597/CTRL 0.01fF
C57323 PAND2X1_553/O POR2X1_106/Y 0.02fF
C57324 POR2X1_78/B PAND2X1_743/O 0.01fF
C57325 POR2X1_52/A PAND2X1_506/CTRL 0.01fF
C57326 POR2X1_526/CTRL VDD -0.00fF
C57327 POR2X1_247/O POR2X1_294/B 0.01fF
C57328 POR2X1_271/B POR2X1_39/B 0.04fF
C57329 POR2X1_842/CTRL POR2X1_737/A 0.01fF
C57330 PAND2X1_287/Y POR2X1_767/O 0.01fF
C57331 PAND2X1_57/B POR2X1_789/A 0.06fF
C57332 POR2X1_407/A POR2X1_728/B 0.02fF
C57333 POR2X1_502/A POR2X1_391/Y 0.10fF
C57334 POR2X1_84/Y POR2X1_786/CTRL 0.01fF
C57335 POR2X1_119/Y POR2X1_271/O 0.07fF
C57336 POR2X1_43/B POR2X1_262/CTRL 0.28fF
C57337 D_INPUT_3 POR2X1_381/O 0.07fF
C57338 PAND2X1_735/Y POR2X1_816/A 0.01fF
C57339 POR2X1_614/A PAND2X1_57/B 0.27fF
C57340 PAND2X1_467/Y POR2X1_72/B 0.03fF
C57341 POR2X1_193/A POR2X1_193/O 0.02fF
C57342 PAND2X1_41/B POR2X1_200/A -0.00fF
C57343 POR2X1_707/B PAND2X1_51/O 0.03fF
C57344 POR2X1_72/B POR2X1_530/CTRL2 0.03fF
C57345 POR2X1_55/Y PAND2X1_506/O 0.02fF
C57346 PAND2X1_805/A PAND2X1_854/A 0.03fF
C57347 PAND2X1_6/A POR2X1_224/m4_208_n4# 0.12fF
C57348 POR2X1_13/A POR2X1_417/CTRL2 0.00fF
C57349 POR2X1_376/B POR2X1_7/A 0.16fF
C57350 PAND2X1_714/Y PAND2X1_169/Y 0.23fF
C57351 PAND2X1_334/CTRL2 POR2X1_42/Y 0.01fF
C57352 PAND2X1_624/CTRL2 POR2X1_283/A 0.04fF
C57353 POR2X1_793/CTRL2 POR2X1_713/B 0.06fF
C57354 PAND2X1_41/B POR2X1_502/CTRL2 0.03fF
C57355 POR2X1_45/Y PAND2X1_197/Y 0.03fF
C57356 PAND2X1_774/CTRL2 VDD 0.00fF
C57357 POR2X1_693/Y POR2X1_697/Y 0.01fF
C57358 POR2X1_673/Y POR2X1_720/Y 0.02fF
C57359 POR2X1_134/Y PAND2X1_768/O 0.03fF
C57360 PAND2X1_57/B POR2X1_38/B 0.03fF
C57361 PAND2X1_73/Y PAND2X1_71/Y 0.03fF
C57362 PAND2X1_180/m4_208_n4# PAND2X1_182/m4_208_n4# 0.13fF
C57363 POR2X1_68/A POR2X1_733/A 0.10fF
C57364 POR2X1_416/B PAND2X1_838/B 0.04fF
C57365 POR2X1_755/Y VDD 0.00fF
C57366 PAND2X1_200/O POR2X1_153/Y 0.09fF
C57367 POR2X1_169/B POR2X1_97/A 0.01fF
C57368 PAND2X1_661/Y PAND2X1_596/O 0.06fF
C57369 PAND2X1_473/B PAND2X1_728/CTRL2 0.03fF
C57370 PAND2X1_833/O POR2X1_283/A 0.02fF
C57371 POR2X1_709/O PAND2X1_90/Y 0.02fF
C57372 PAND2X1_535/Y PAND2X1_863/B 0.02fF
C57373 POR2X1_202/CTRL POR2X1_507/A 0.03fF
C57374 POR2X1_786/Y POR2X1_740/Y 0.10fF
C57375 POR2X1_286/B PAND2X1_52/B 0.00fF
C57376 POR2X1_614/A POR2X1_341/CTRL2 0.03fF
C57377 POR2X1_562/a_56_344# POR2X1_562/B 0.00fF
C57378 PAND2X1_58/A PAND2X1_142/a_56_28# 0.00fF
C57379 POR2X1_606/CTRL PAND2X1_56/A 0.01fF
C57380 INPUT_4 POR2X1_386/a_16_28# 0.03fF
C57381 POR2X1_460/a_16_28# POR2X1_460/B 0.01fF
C57382 PAND2X1_391/a_16_344# POR2X1_4/Y 0.02fF
C57383 POR2X1_831/CTRL POR2X1_717/B 0.01fF
C57384 POR2X1_51/A POR2X1_36/m4_208_n4# 0.01fF
C57385 POR2X1_614/A POR2X1_193/O 0.04fF
C57386 POR2X1_479/a_16_28# POR2X1_774/A 0.03fF
C57387 PAND2X1_738/Y PAND2X1_181/CTRL2 0.17fF
C57388 POR2X1_322/Y POR2X1_46/Y 0.03fF
C57389 POR2X1_567/A POR2X1_555/B 0.40fF
C57390 PAND2X1_23/Y PAND2X1_96/B 0.38fF
C57391 PAND2X1_81/B PAND2X1_316/O 0.05fF
C57392 POR2X1_250/O POR2X1_283/A 0.01fF
C57393 PAND2X1_682/CTRL2 PAND2X1_69/A 0.01fF
C57394 POR2X1_547/O POR2X1_614/A 0.03fF
C57395 POR2X1_707/B PAND2X1_3/B 0.05fF
C57396 PAND2X1_48/B POR2X1_736/CTRL 0.00fF
C57397 POR2X1_152/a_16_28# POR2X1_152/A 0.00fF
C57398 POR2X1_360/A PAND2X1_60/B 0.09fF
C57399 POR2X1_369/Y POR2X1_83/B 0.04fF
C57400 POR2X1_814/B POR2X1_544/B 0.07fF
C57401 POR2X1_774/A POR2X1_734/A 0.03fF
C57402 PAND2X1_535/Y PAND2X1_567/O 0.00fF
C57403 PAND2X1_625/O PAND2X1_96/B 0.15fF
C57404 POR2X1_41/B PAND2X1_196/CTRL2 0.01fF
C57405 POR2X1_52/A POR2X1_7/A 0.15fF
C57406 PAND2X1_425/O PAND2X1_18/B 0.01fF
C57407 POR2X1_862/Y PAND2X1_52/B 0.04fF
C57408 POR2X1_614/A POR2X1_828/A 1.64fF
C57409 POR2X1_775/CTRL PAND2X1_32/B 0.01fF
C57410 POR2X1_96/A POR2X1_679/B 0.00fF
C57411 PAND2X1_744/CTRL POR2X1_532/A 0.01fF
C57412 PAND2X1_297/O PAND2X1_57/B 0.03fF
C57413 PAND2X1_808/CTRL2 POR2X1_283/A 0.01fF
C57414 POR2X1_833/O PAND2X1_60/B 0.01fF
C57415 PAND2X1_338/B PAND2X1_101/O 0.01fF
C57416 PAND2X1_56/Y PAND2X1_306/CTRL 0.05fF
C57417 POR2X1_156/CTRL POR2X1_750/B 0.01fF
C57418 POR2X1_346/B POR2X1_220/Y 0.03fF
C57419 POR2X1_502/A POR2X1_834/Y 0.05fF
C57420 INPUT_6 PAND2X1_587/CTRL2 0.00fF
C57421 POR2X1_544/B POR2X1_325/A 0.04fF
C57422 PAND2X1_220/a_16_344# PAND2X1_213/Y 0.01fF
C57423 INPUT_1 POR2X1_625/Y 0.03fF
C57424 PAND2X1_854/O PAND2X1_854/A 0.00fF
C57425 POR2X1_278/Y PAND2X1_343/O 0.07fF
C57426 POR2X1_309/CTRL POR2X1_39/B 0.01fF
C57427 POR2X1_532/A POR2X1_771/CTRL 0.01fF
C57428 POR2X1_85/O POR2X1_83/B 0.01fF
C57429 POR2X1_16/A PAND2X1_350/A 0.00fF
C57430 PAND2X1_542/CTRL2 VDD 0.00fF
C57431 POR2X1_207/A POR2X1_195/CTRL 0.01fF
C57432 PAND2X1_63/Y PAND2X1_79/Y 0.05fF
C57433 POR2X1_281/CTRL PAND2X1_809/A 0.03fF
C57434 POR2X1_43/B PAND2X1_549/B 0.03fF
C57435 POR2X1_334/O POR2X1_360/A 0.04fF
C57436 PAND2X1_808/Y PAND2X1_363/O 0.02fF
C57437 POR2X1_57/A POR2X1_73/Y 0.24fF
C57438 POR2X1_170/CTRL2 POR2X1_566/B 0.01fF
C57439 POR2X1_557/A PAND2X1_90/A 0.03fF
C57440 POR2X1_12/A POR2X1_698/Y 0.22fF
C57441 PAND2X1_117/O POR2X1_260/A 0.01fF
C57442 POR2X1_624/a_16_28# POR2X1_623/Y 0.03fF
C57443 PAND2X1_508/Y VDD 0.27fF
C57444 POR2X1_13/A POR2X1_129/Y 0.06fF
C57445 PAND2X1_58/A POR2X1_711/Y 0.08fF
C57446 POR2X1_811/B POR2X1_779/O 0.01fF
C57447 POR2X1_567/A POR2X1_776/O 0.08fF
C57448 POR2X1_832/A POR2X1_435/O 0.16fF
C57449 POR2X1_730/Y POR2X1_477/A 0.03fF
C57450 PAND2X1_539/Y PAND2X1_567/O 0.00fF
C57451 PAND2X1_383/a_16_344# POR2X1_816/A 0.01fF
C57452 POR2X1_304/O POR2X1_40/Y 0.08fF
C57453 POR2X1_463/Y PAND2X1_55/Y 0.07fF
C57454 POR2X1_777/B PAND2X1_136/O 0.04fF
C57455 POR2X1_383/A POR2X1_631/B 0.04fF
C57456 POR2X1_809/A POR2X1_435/Y -0.00fF
C57457 PAND2X1_329/CTRL2 POR2X1_532/A 0.03fF
C57458 POR2X1_101/CTRL PAND2X1_69/A 0.03fF
C57459 PAND2X1_693/a_16_344# PAND2X1_94/A 0.02fF
C57460 POR2X1_383/A POR2X1_784/CTRL2 0.01fF
C57461 PAND2X1_693/O INPUT_1 0.03fF
C57462 POR2X1_25/a_16_28# PAND2X1_18/B 0.09fF
C57463 PAND2X1_717/A POR2X1_150/Y 0.46fF
C57464 POR2X1_816/A POR2X1_171/CTRL 0.01fF
C57465 POR2X1_509/B POR2X1_568/B 0.01fF
C57466 POR2X1_145/CTRL POR2X1_394/A 0.01fF
C57467 PAND2X1_569/A PAND2X1_569/B 0.14fF
C57468 POR2X1_110/Y PAND2X1_471/O 0.07fF
C57469 PAND2X1_324/O POR2X1_321/Y 0.00fF
C57470 PAND2X1_659/Y POR2X1_13/A 0.03fF
C57471 POR2X1_294/B POR2X1_715/A 0.01fF
C57472 POR2X1_575/B POR2X1_574/Y 0.01fF
C57473 PAND2X1_297/CTRL PAND2X1_69/A 0.01fF
C57474 PAND2X1_57/B POR2X1_398/a_16_28# 0.01fF
C57475 PAND2X1_803/Y PAND2X1_843/Y 0.03fF
C57476 POR2X1_316/CTRL2 POR2X1_43/B 0.00fF
C57477 PAND2X1_841/a_16_344# POR2X1_271/A 0.01fF
C57478 POR2X1_242/CTRL PAND2X1_52/B 0.01fF
C57479 PAND2X1_651/Y PAND2X1_861/O 0.04fF
C57480 D_GATE_662 POR2X1_544/Y 0.04fF
C57481 PAND2X1_242/Y POR2X1_496/Y 0.09fF
C57482 POR2X1_760/A POR2X1_411/B 0.07fF
C57483 POR2X1_178/CTRL PAND2X1_348/A 0.03fF
C57484 POR2X1_96/Y POR2X1_13/A 0.02fF
C57485 PAND2X1_568/B PAND2X1_578/CTRL 0.01fF
C57486 PAND2X1_48/B POR2X1_359/CTRL2 0.01fF
C57487 POR2X1_110/Y PAND2X1_465/B 0.02fF
C57488 POR2X1_94/A PAND2X1_52/B 0.05fF
C57489 PAND2X1_687/B POR2X1_13/A 0.01fF
C57490 POR2X1_366/Y POR2X1_703/O 0.04fF
C57491 POR2X1_614/A POR2X1_259/B 0.01fF
C57492 POR2X1_578/a_16_28# POR2X1_568/Y -0.00fF
C57493 PAND2X1_696/O POR2X1_502/A 0.32fF
C57494 POR2X1_137/Y POR2X1_362/A 0.02fF
C57495 POR2X1_85/CTRL2 PAND2X1_35/Y 0.01fF
C57496 PAND2X1_716/B PAND2X1_302/O 0.03fF
C57497 PAND2X1_6/Y POR2X1_334/Y 0.14fF
C57498 PAND2X1_736/A POR2X1_385/Y 0.10fF
C57499 PAND2X1_569/B PAND2X1_854/A 0.14fF
C57500 POR2X1_327/Y PAND2X1_69/A 2.06fF
C57501 POR2X1_502/A POR2X1_383/Y 0.05fF
C57502 INPUT_3 PAND2X1_33/O 0.02fF
C57503 PAND2X1_864/O PAND2X1_568/B 0.05fF
C57504 POR2X1_164/Y PAND2X1_550/Y 0.00fF
C57505 PAND2X1_310/CTRL POR2X1_501/B 0.01fF
C57506 POR2X1_496/CTRL POR2X1_20/B 0.01fF
C57507 PAND2X1_107/a_76_28# POR2X1_532/A 0.06fF
C57508 PAND2X1_632/A PAND2X1_632/B 0.03fF
C57509 POR2X1_131/Y PAND2X1_349/A 0.01fF
C57510 PAND2X1_408/Y PAND2X1_18/B 0.01fF
C57511 POR2X1_614/A POR2X1_512/CTRL2 0.01fF
C57512 POR2X1_307/Y POR2X1_513/A 0.01fF
C57513 PAND2X1_860/A PAND2X1_360/O 0.03fF
C57514 PAND2X1_743/O POR2X1_294/A 0.01fF
C57515 POR2X1_119/Y PAND2X1_472/A 0.07fF
C57516 POR2X1_508/A POR2X1_508/a_16_28# 0.04fF
C57517 POR2X1_727/CTRL POR2X1_353/A 0.01fF
C57518 PAND2X1_865/Y POR2X1_437/Y 0.00fF
C57519 POR2X1_375/CTRL2 POR2X1_260/A 0.03fF
C57520 PAND2X1_26/CTRL PAND2X1_18/B 0.01fF
C57521 PAND2X1_653/O PAND2X1_652/Y 0.00fF
C57522 POR2X1_13/A PAND2X1_333/Y 0.03fF
C57523 POR2X1_203/CTRL2 PAND2X1_48/A 0.01fF
C57524 PAND2X1_630/O PAND2X1_508/B 0.03fF
C57525 POR2X1_406/Y PAND2X1_332/Y 0.01fF
C57526 POR2X1_725/Y POR2X1_186/B 0.09fF
C57527 POR2X1_431/O POR2X1_67/A 0.02fF
C57528 PAND2X1_55/Y POR2X1_736/A 1.61fF
C57529 PAND2X1_242/CTRL2 POR2X1_77/Y 0.08fF
C57530 POR2X1_96/A POR2X1_759/CTRL 0.01fF
C57531 POR2X1_42/a_76_344# POR2X1_4/Y 0.02fF
C57532 POR2X1_16/A POR2X1_39/Y 0.02fF
C57533 PAND2X1_687/B PAND2X1_643/Y 0.07fF
C57534 POR2X1_571/Y PAND2X1_60/B 0.03fF
C57535 POR2X1_537/Y POR2X1_537/B 0.00fF
C57536 POR2X1_711/B POR2X1_713/B 0.77fF
C57537 POR2X1_76/a_56_344# POR2X1_76/A 0.00fF
C57538 POR2X1_508/a_16_28# POR2X1_568/B 0.02fF
C57539 POR2X1_44/O PAND2X1_635/Y 0.01fF
C57540 POR2X1_262/Y D_INPUT_0 0.07fF
C57541 POR2X1_765/Y POR2X1_766/Y 0.02fF
C57542 POR2X1_532/A PAND2X1_134/a_16_344# 0.06fF
C57543 PAND2X1_865/CTRL PAND2X1_862/Y 0.01fF
C57544 POR2X1_293/Y PAND2X1_332/Y 0.19fF
C57545 POR2X1_83/B POR2X1_431/a_76_344# 0.00fF
C57546 PAND2X1_41/CTRL2 POR2X1_66/A 0.01fF
C57547 POR2X1_84/A POR2X1_240/CTRL 0.09fF
C57548 PAND2X1_845/O POR2X1_39/B 0.24fF
C57549 POR2X1_305/Y POR2X1_416/B 0.08fF
C57550 POR2X1_9/Y PAND2X1_340/O 0.09fF
C57551 PAND2X1_797/Y PAND2X1_803/Y 0.05fF
C57552 PAND2X1_111/CTRL2 PAND2X1_72/A 0.00fF
C57553 POR2X1_16/A POR2X1_314/Y 0.04fF
C57554 POR2X1_639/Y D_INPUT_4 0.12fF
C57555 POR2X1_445/A POR2X1_856/B 0.01fF
C57556 PAND2X1_404/Y POR2X1_23/Y 0.03fF
C57557 PAND2X1_96/B POR2X1_711/Y 0.19fF
C57558 POR2X1_506/CTRL2 POR2X1_508/B 0.00fF
C57559 POR2X1_774/Y POR2X1_814/A 0.05fF
C57560 POR2X1_38/CTRL2 POR2X1_37/Y 0.01fF
C57561 POR2X1_105/Y POR2X1_814/A 0.39fF
C57562 POR2X1_415/A POR2X1_669/B 0.10fF
C57563 POR2X1_311/Y POR2X1_411/B 0.03fF
C57564 POR2X1_796/Y POR2X1_808/B 0.01fF
C57565 POR2X1_156/a_16_28# POR2X1_162/Y 0.01fF
C57566 POR2X1_452/O POR2X1_121/B 0.06fF
C57567 POR2X1_633/A POR2X1_633/a_16_28# 0.00fF
C57568 POR2X1_137/B POR2X1_634/CTRL 0.02fF
C57569 POR2X1_77/a_16_28# POR2X1_48/A 0.02fF
C57570 POR2X1_66/B POR2X1_556/A 0.06fF
C57571 PAND2X1_270/O POR2X1_39/B 0.04fF
C57572 PAND2X1_159/CTRL PAND2X1_9/Y 0.01fF
C57573 PAND2X1_418/O PAND2X1_41/B 0.01fF
C57574 PAND2X1_865/Y POR2X1_16/A 0.51fF
C57575 POR2X1_649/O POR2X1_643/A 0.07fF
C57576 POR2X1_447/B POR2X1_507/A 0.02fF
C57577 POR2X1_394/A POR2X1_599/m4_208_n4# 0.15fF
C57578 POR2X1_49/CTRL2 PAND2X1_9/Y 0.01fF
C57579 PAND2X1_844/B PAND2X1_351/A 0.00fF
C57580 POR2X1_825/Y PAND2X1_334/CTRL 0.00fF
C57581 POR2X1_143/O POR2X1_9/Y 0.31fF
C57582 POR2X1_748/Y POR2X1_39/B 0.09fF
C57583 POR2X1_646/A POR2X1_480/A 0.07fF
C57584 PAND2X1_20/A POR2X1_659/A 0.03fF
C57585 POR2X1_632/B POR2X1_632/CTRL 0.00fF
C57586 POR2X1_609/Y POR2X1_48/A 0.03fF
C57587 POR2X1_600/Y POR2X1_601/m4_208_n4# 0.15fF
C57588 PAND2X1_476/A PAND2X1_560/B 0.03fF
C57589 PAND2X1_617/CTRL VDD 0.00fF
C57590 POR2X1_537/Y PAND2X1_48/A 0.03fF
C57591 POR2X1_257/A PAND2X1_725/Y 0.01fF
C57592 PAND2X1_806/CTRL2 PAND2X1_362/A 0.01fF
C57593 PAND2X1_464/B VDD 0.30fF
C57594 POR2X1_814/A PAND2X1_257/CTRL 0.06fF
C57595 PAND2X1_832/O POR2X1_411/B 0.02fF
C57596 POR2X1_477/CTRL2 POR2X1_480/A 0.03fF
C57597 POR2X1_254/A POR2X1_454/A 0.08fF
C57598 POR2X1_567/A POR2X1_703/O 0.01fF
C57599 POR2X1_849/A POR2X1_590/A 1.03fF
C57600 PAND2X1_448/a_16_344# POR2X1_32/A 0.03fF
C57601 POR2X1_48/A POR2X1_420/Y 0.01fF
C57602 POR2X1_567/A POR2X1_337/Y 0.07fF
C57603 POR2X1_20/B POR2X1_236/Y 0.13fF
C57604 PAND2X1_9/CTRL2 D_INPUT_0 0.01fF
C57605 POR2X1_362/Y D_INPUT_0 0.03fF
C57606 PAND2X1_477/a_76_28# POR2X1_102/Y 0.02fF
C57607 POR2X1_416/B PAND2X1_537/a_16_344# 0.02fF
C57608 PAND2X1_850/Y PAND2X1_716/B 0.07fF
C57609 POR2X1_52/A POR2X1_760/A 0.02fF
C57610 POR2X1_411/B PAND2X1_719/CTRL 0.01fF
C57611 PAND2X1_771/Y PAND2X1_542/a_76_28# 0.04fF
C57612 POR2X1_334/Y POR2X1_632/Y 0.07fF
C57613 POR2X1_257/A POR2X1_697/O 0.01fF
C57614 POR2X1_497/CTRL2 POR2X1_32/A 0.03fF
C57615 POR2X1_411/B POR2X1_609/A 0.55fF
C57616 PAND2X1_243/B POR2X1_669/Y 0.03fF
C57617 POR2X1_60/A POR2X1_496/Y 0.10fF
C57618 POR2X1_41/B POR2X1_150/Y 0.14fF
C57619 POR2X1_41/B PAND2X1_838/CTRL2 0.01fF
C57620 POR2X1_661/A PAND2X1_305/CTRL2 -0.02fF
C57621 POR2X1_96/A PAND2X1_203/CTRL2 0.01fF
C57622 POR2X1_814/A POR2X1_467/CTRL 0.06fF
C57623 PAND2X1_791/O VDD 0.00fF
C57624 POR2X1_696/O POR2X1_32/A 0.01fF
C57625 PAND2X1_857/A PAND2X1_193/Y 0.08fF
C57626 POR2X1_81/Y POR2X1_20/B 0.02fF
C57627 PAND2X1_644/O POR2X1_683/Y 0.00fF
C57628 PAND2X1_557/A POR2X1_32/A 0.03fF
C57629 POR2X1_857/B POR2X1_857/A 0.01fF
C57630 PAND2X1_73/Y POR2X1_634/O 0.01fF
C57631 POR2X1_830/CTRL2 POR2X1_830/Y 0.09fF
C57632 POR2X1_650/A POR2X1_558/B 0.03fF
C57633 PAND2X1_20/A POR2X1_14/Y 0.03fF
C57634 PAND2X1_207/m4_208_n4# POR2X1_40/Y 0.08fF
C57635 PAND2X1_230/a_76_28# POR2X1_78/A 0.00fF
C57636 PAND2X1_699/CTRL PAND2X1_6/A 0.01fF
C57637 POR2X1_77/Y POR2X1_171/Y 0.17fF
C57638 POR2X1_415/A POR2X1_617/CTRL2 0.05fF
C57639 POR2X1_16/A POR2X1_91/O 0.02fF
C57640 PAND2X1_281/O PAND2X1_52/B 0.03fF
C57641 POR2X1_60/A PAND2X1_733/A 0.03fF
C57642 POR2X1_335/CTRL2 POR2X1_66/A 0.04fF
C57643 POR2X1_302/B PAND2X1_279/CTRL 0.01fF
C57644 POR2X1_29/A PAND2X1_793/A 0.51fF
C57645 POR2X1_102/Y POR2X1_423/Y 0.18fF
C57646 PAND2X1_304/CTRL2 PAND2X1_56/A 0.01fF
C57647 POR2X1_69/a_16_28# POR2X1_69/A 0.04fF
C57648 PAND2X1_474/Y POR2X1_37/Y 0.03fF
C57649 PAND2X1_447/a_16_344# POR2X1_90/Y 0.01fF
C57650 POR2X1_158/CTRL2 POR2X1_416/B 0.00fF
C57651 POR2X1_805/Y POR2X1_791/Y 0.00fF
C57652 POR2X1_411/B PAND2X1_218/A 0.18fF
C57653 POR2X1_669/B POR2X1_692/Y 0.14fF
C57654 PAND2X1_124/Y POR2X1_46/Y 0.03fF
C57655 PAND2X1_20/A POR2X1_849/CTRL2 0.01fF
C57656 POR2X1_461/Y POR2X1_793/A 0.01fF
C57657 POR2X1_16/A POR2X1_16/m4_208_n4# 0.01fF
C57658 POR2X1_434/A VDD -0.00fF
C57659 POR2X1_850/B POR2X1_850/A 0.13fF
C57660 PAND2X1_234/CTRL POR2X1_260/A 0.01fF
C57661 POR2X1_705/B POR2X1_705/a_16_28# 0.08fF
C57662 POR2X1_13/A POR2X1_37/Y 0.10fF
C57663 PAND2X1_20/A POR2X1_637/B 0.00fF
C57664 POR2X1_827/Y POR2X1_42/Y 0.02fF
C57665 PAND2X1_97/O POR2X1_293/Y 0.08fF
C57666 POR2X1_490/CTRL POR2X1_73/Y 0.01fF
C57667 PAND2X1_859/B POR2X1_93/Y 0.03fF
C57668 POR2X1_48/A POR2X1_277/CTRL 0.01fF
C57669 POR2X1_63/Y PAND2X1_734/O 0.03fF
C57670 POR2X1_807/A POR2X1_330/Y 0.05fF
C57671 POR2X1_857/CTRL VDD 0.00fF
C57672 PAND2X1_73/Y INPUT_0 2.17fF
C57673 POR2X1_54/Y POR2X1_816/A 0.03fF
C57674 POR2X1_32/A PAND2X1_151/O 0.04fF
C57675 POR2X1_411/B POR2X1_38/Y 0.13fF
C57676 POR2X1_54/Y POR2X1_462/B 0.08fF
C57677 POR2X1_20/B PAND2X1_344/CTRL 0.02fF
C57678 PAND2X1_90/A PAND2X1_613/m4_208_n4# 0.12fF
C57679 POR2X1_54/Y D_INPUT_1 4.12fF
C57680 PAND2X1_657/CTRL PAND2X1_659/B 0.00fF
C57681 POR2X1_270/Y PAND2X1_55/Y 0.03fF
C57682 POR2X1_558/B POR2X1_294/B 0.09fF
C57683 PAND2X1_57/B POR2X1_590/A 0.68fF
C57684 POR2X1_431/Y POR2X1_172/Y 0.04fF
C57685 POR2X1_860/O POR2X1_814/A 0.01fF
C57686 PAND2X1_806/a_16_344# POR2X1_42/Y 0.02fF
C57687 POR2X1_697/CTRL POR2X1_40/Y 0.01fF
C57688 POR2X1_260/B PAND2X1_6/A 0.62fF
C57689 PAND2X1_793/Y POR2X1_67/A 0.02fF
C57690 PAND2X1_93/B D_GATE_222 0.03fF
C57691 POR2X1_814/B POR2X1_791/Y 0.01fF
C57692 PAND2X1_289/O POR2X1_220/A 0.01fF
C57693 POR2X1_56/B POR2X1_669/B 2.41fF
C57694 POR2X1_264/CTRL INPUT_0 0.07fF
C57695 POR2X1_814/B POR2X1_637/B 0.76fF
C57696 POR2X1_83/B POR2X1_46/Y 0.06fF
C57697 POR2X1_413/A POR2X1_609/Y 0.03fF
C57698 POR2X1_355/B PAND2X1_20/A 0.03fF
C57699 POR2X1_16/A PAND2X1_608/a_76_28# 0.02fF
C57700 POR2X1_66/A PAND2X1_144/O 0.03fF
C57701 POR2X1_270/O POR2X1_445/A 0.08fF
C57702 POR2X1_528/Y POR2X1_744/Y 0.03fF
C57703 PAND2X1_463/CTRL PAND2X1_460/Y 0.01fF
C57704 PAND2X1_307/O POR2X1_304/Y -0.00fF
C57705 POR2X1_72/B PAND2X1_556/B 0.05fF
C57706 POR2X1_603/Y POR2X1_7/B 0.00fF
C57707 POR2X1_417/Y PAND2X1_151/O 0.03fF
C57708 POR2X1_71/Y POR2X1_516/Y 0.05fF
C57709 PAND2X1_793/Y PAND2X1_78/CTRL 0.01fF
C57710 POR2X1_66/B POR2X1_445/CTRL 0.00fF
C57711 POR2X1_23/Y PAND2X1_565/A 0.03fF
C57712 POR2X1_458/CTRL2 POR2X1_458/B 0.01fF
C57713 POR2X1_482/CTRL PAND2X1_6/A 0.01fF
C57714 POR2X1_236/CTRL POR2X1_5/Y 0.01fF
C57715 POR2X1_146/CTRL2 POR2X1_257/A 0.10fF
C57716 POR2X1_285/A POR2X1_590/A 0.01fF
C57717 PAND2X1_412/CTRL2 POR2X1_546/A 0.03fF
C57718 PAND2X1_485/O PAND2X1_69/A 0.01fF
C57719 PAND2X1_192/Y PAND2X1_739/CTRL 0.01fF
C57720 POR2X1_49/Y POR2X1_88/Y 0.06fF
C57721 PAND2X1_58/A POR2X1_733/A 0.07fF
C57722 PAND2X1_454/O POR2X1_60/A 0.05fF
C57723 POR2X1_307/B POR2X1_480/A 0.07fF
C57724 PAND2X1_360/CTRL2 POR2X1_42/Y 0.01fF
C57725 PAND2X1_512/CTRL POR2X1_7/B 0.00fF
C57726 PAND2X1_864/B PAND2X1_810/A 0.00fF
C57727 PAND2X1_261/m4_208_n4# POR2X1_330/Y 0.12fF
C57728 POR2X1_814/A POR2X1_773/A 0.01fF
C57729 POR2X1_66/B PAND2X1_385/CTRL 0.01fF
C57730 INPUT_1 POR2X1_411/B 0.10fF
C57731 POR2X1_78/A D_GATE_222 0.15fF
C57732 PAND2X1_661/B POR2X1_37/Y 0.03fF
C57733 POR2X1_478/a_16_28# POR2X1_478/B 0.01fF
C57734 PAND2X1_478/B PAND2X1_478/CTRL2 0.01fF
C57735 PAND2X1_212/B PAND2X1_357/Y 0.01fF
C57736 PAND2X1_95/B POR2X1_638/A 0.00fF
C57737 D_INPUT_5 PAND2X1_1/O 0.04fF
C57738 PAND2X1_65/CTRL2 POR2X1_205/A 0.04fF
C57739 PAND2X1_540/CTRL PAND2X1_553/B 0.06fF
C57740 POR2X1_244/B POR2X1_193/Y 0.05fF
C57741 PAND2X1_840/A POR2X1_83/B 0.05fF
C57742 PAND2X1_391/a_16_344# POR2X1_816/A 0.01fF
C57743 POR2X1_355/B POR2X1_814/B 0.07fF
C57744 POR2X1_428/Y POR2X1_158/B 0.03fF
C57745 POR2X1_814/B PAND2X1_183/CTRL 0.06fF
C57746 POR2X1_32/a_16_28# POR2X1_14/Y 0.03fF
C57747 POR2X1_300/CTRL2 PAND2X1_217/B -0.01fF
C57748 POR2X1_68/A PAND2X1_394/O 0.02fF
C57749 POR2X1_271/A POR2X1_20/B 0.04fF
C57750 PAND2X1_23/Y POR2X1_355/A 4.33fF
C57751 POR2X1_355/CTRL2 PAND2X1_23/Y 0.01fF
C57752 PAND2X1_474/Y POR2X1_406/Y 0.01fF
C57753 POR2X1_529/a_16_28# POR2X1_83/B 0.06fF
C57754 PAND2X1_84/Y PAND2X1_579/B 0.03fF
C57755 PAND2X1_631/A POR2X1_329/A 0.07fF
C57756 POR2X1_411/B POR2X1_153/Y 4.41fF
C57757 PAND2X1_633/Y PAND2X1_404/Y 0.13fF
C57758 POR2X1_483/A POR2X1_483/O 0.08fF
C57759 POR2X1_49/Y POR2X1_743/Y 0.02fF
C57760 POR2X1_260/B POR2X1_101/Y 0.10fF
C57761 POR2X1_355/A PAND2X1_504/CTRL2 0.01fF
C57762 POR2X1_411/B POR2X1_384/A 0.03fF
C57763 PAND2X1_824/B POR2X1_240/CTRL2 0.01fF
C57764 PAND2X1_20/A POR2X1_139/a_56_344# 0.00fF
C57765 POR2X1_140/B POR2X1_330/Y 0.05fF
C57766 POR2X1_72/B POR2X1_599/A 0.03fF
C57767 POR2X1_629/B PAND2X1_69/A 0.60fF
C57768 POR2X1_32/A PAND2X1_350/CTRL2 0.01fF
C57769 POR2X1_337/A POR2X1_270/Y 0.06fF
C57770 POR2X1_407/A POR2X1_330/Y 0.05fF
C57771 POR2X1_463/Y POR2X1_805/CTRL2 0.00fF
C57772 POR2X1_526/a_16_28# POR2X1_669/B 0.09fF
C57773 PAND2X1_425/Y PAND2X1_18/B 0.03fF
C57774 PAND2X1_73/Y POR2X1_780/A 0.48fF
C57775 PAND2X1_372/CTRL VDD -0.00fF
C57776 POR2X1_192/Y POR2X1_223/CTRL2 0.01fF
C57777 POR2X1_304/Y POR2X1_96/A 0.01fF
C57778 POR2X1_538/CTRL POR2X1_814/B 0.01fF
C57779 PAND2X1_16/m4_208_n4# POR2X1_785/A 0.15fF
C57780 POR2X1_37/Y PAND2X1_510/B 0.03fF
C57781 POR2X1_317/O PAND2X1_90/Y 0.01fF
C57782 PAND2X1_57/B PAND2X1_57/a_76_28# 0.02fF
C57783 PAND2X1_94/A POR2X1_33/A 0.03fF
C57784 POR2X1_96/A PAND2X1_862/B 0.03fF
C57785 PAND2X1_474/Y POR2X1_293/Y 0.04fF
C57786 PAND2X1_715/CTRL POR2X1_293/Y 0.01fF
C57787 POR2X1_175/m4_208_n4# POR2X1_566/A 0.03fF
C57788 POR2X1_20/B PAND2X1_352/CTRL2 0.00fF
C57789 POR2X1_809/A POR2X1_676/CTRL2 0.01fF
C57790 POR2X1_444/CTRL POR2X1_191/Y 0.00fF
C57791 PAND2X1_140/A POR2X1_127/a_76_344# 0.00fF
C57792 POR2X1_251/Y PAND2X1_137/Y 0.04fF
C57793 PAND2X1_465/B INPUT_0 0.07fF
C57794 PAND2X1_46/CTRL POR2X1_68/B 0.01fF
C57795 POR2X1_856/B POR2X1_260/A 0.18fF
C57796 POR2X1_66/A POR2X1_456/B 0.03fF
C57797 POR2X1_257/A POR2X1_766/Y 0.03fF
C57798 POR2X1_13/A POR2X1_293/Y 0.85fF
C57799 POR2X1_566/A POR2X1_231/B 0.05fF
C57800 PAND2X1_787/Y PAND2X1_794/B 0.01fF
C57801 POR2X1_41/B PAND2X1_364/B 0.07fF
C57802 POR2X1_68/A PAND2X1_525/a_56_28# 0.00fF
C57803 PAND2X1_693/CTRL VDD 0.00fF
C57804 POR2X1_368/Y POR2X1_5/Y 0.01fF
C57805 POR2X1_672/CTRL POR2X1_5/Y 0.01fF
C57806 POR2X1_549/A PAND2X1_8/Y 0.01fF
C57807 POR2X1_356/A POR2X1_855/Y 0.05fF
C57808 POR2X1_646/CTRL2 POR2X1_294/B 0.03fF
C57809 POR2X1_814/B POR2X1_791/B 0.02fF
C57810 POR2X1_66/B POR2X1_276/A 0.02fF
C57811 PAND2X1_226/CTRL POR2X1_578/Y 0.03fF
C57812 PAND2X1_798/B INPUT_0 0.05fF
C57813 PAND2X1_808/B PAND2X1_803/Y 0.01fF
C57814 PAND2X1_20/A POR2X1_472/m4_208_n4# 0.12fF
C57815 POR2X1_177/Y POR2X1_90/Y 0.04fF
C57816 POR2X1_319/A POR2X1_192/B 0.03fF
C57817 POR2X1_425/Y POR2X1_427/Y 0.00fF
C57818 POR2X1_376/B POR2X1_38/Y 0.03fF
C57819 POR2X1_840/B POR2X1_362/B 0.05fF
C57820 POR2X1_65/A PAND2X1_213/Y 0.03fF
C57821 POR2X1_78/A POR2X1_592/A 0.00fF
C57822 PAND2X1_6/Y POR2X1_349/Y 0.02fF
C57823 PAND2X1_14/O D_INPUT_1 0.01fF
C57824 PAND2X1_477/A POR2X1_102/Y 0.05fF
C57825 PAND2X1_85/Y POR2X1_38/B 0.03fF
C57826 POR2X1_46/a_16_28# PAND2X1_338/B 0.03fF
C57827 PAND2X1_228/O PAND2X1_364/B 0.05fF
C57828 POR2X1_211/O VDD 0.00fF
C57829 PAND2X1_90/Y POR2X1_540/CTRL 0.00fF
C57830 PAND2X1_41/B POR2X1_713/B 0.03fF
C57831 POR2X1_684/O POR2X1_42/Y 0.03fF
C57832 POR2X1_346/B PAND2X1_626/CTRL 0.00fF
C57833 PAND2X1_80/O D_INPUT_1 0.06fF
C57834 PAND2X1_738/A PAND2X1_738/B 0.10fF
C57835 PAND2X1_525/CTRL2 POR2X1_550/Y 0.00fF
C57836 PAND2X1_424/CTRL POR2X1_480/A 0.03fF
C57837 PAND2X1_84/Y POR2X1_73/Y 0.03fF
C57838 POR2X1_614/A POR2X1_812/CTRL2 0.03fF
C57839 POR2X1_25/Y POR2X1_48/A 0.01fF
C57840 POR2X1_150/Y POR2X1_77/Y 0.05fF
C57841 PAND2X1_632/B POR2X1_748/A 0.03fF
C57842 POR2X1_63/Y POR2X1_39/B 0.05fF
C57843 POR2X1_28/CTRL POR2X1_4/Y 0.07fF
C57844 POR2X1_29/A POR2X1_129/Y 0.02fF
C57845 POR2X1_57/A PAND2X1_804/A 0.04fF
C57846 PAND2X1_65/B PAND2X1_312/a_16_344# 0.05fF
C57847 PAND2X1_84/CTRL POR2X1_91/Y 0.01fF
C57848 INPUT_1 POR2X1_24/CTRL2 0.01fF
C57849 POR2X1_45/Y POR2X1_48/Y 0.11fF
C57850 PAND2X1_241/CTRL POR2X1_237/Y 0.01fF
C57851 POR2X1_130/O POR2X1_66/B 0.01fF
C57852 POR2X1_142/CTRL POR2X1_394/A 0.08fF
C57853 POR2X1_558/O POR2X1_264/Y 0.01fF
C57854 POR2X1_41/B POR2X1_229/O 0.00fF
C57855 POR2X1_331/A POR2X1_594/A 0.07fF
C57856 PAND2X1_6/Y POR2X1_629/A 0.04fF
C57857 POR2X1_68/A POR2X1_477/A 0.01fF
C57858 POR2X1_566/A PAND2X1_88/Y 0.05fF
C57859 POR2X1_38/Y PAND2X1_598/O 0.05fF
C57860 PAND2X1_55/Y PAND2X1_6/A 0.00fF
C57861 POR2X1_793/A POR2X1_789/Y 0.01fF
C57862 POR2X1_106/Y PAND2X1_114/CTRL2 0.01fF
C57863 POR2X1_481/A POR2X1_387/Y 0.04fF
C57864 D_INPUT_3 POR2X1_58/m4_208_n4# 0.06fF
C57865 POR2X1_271/Y POR2X1_153/Y 0.01fF
C57866 PAND2X1_856/B PAND2X1_805/A 0.03fF
C57867 POR2X1_406/a_16_28# POR2X1_406/A 0.05fF
C57868 PAND2X1_193/Y POR2X1_329/A 0.03fF
C57869 POR2X1_504/CTRL2 POR2X1_504/Y 0.01fF
C57870 PAND2X1_551/O VDD 0.00fF
C57871 POR2X1_76/Y POR2X1_541/a_76_344# 0.00fF
C57872 POR2X1_8/Y POR2X1_49/Y 0.06fF
C57873 POR2X1_795/B POR2X1_35/Y 0.00fF
C57874 POR2X1_751/CTRL2 POR2X1_7/B 0.03fF
C57875 POR2X1_369/a_16_28# POR2X1_60/A 0.04fF
C57876 POR2X1_332/B PAND2X1_111/B 0.01fF
C57877 PAND2X1_386/O POR2X1_260/A 0.02fF
C57878 POR2X1_283/A VDD 1.24fF
C57879 POR2X1_52/A POR2X1_38/Y 3.37fF
C57880 POR2X1_60/A POR2X1_75/Y 0.71fF
C57881 POR2X1_66/B POR2X1_398/O 0.01fF
C57882 INPUT_1 POR2X1_376/B 0.84fF
C57883 POR2X1_13/A POR2X1_408/Y 0.03fF
C57884 PAND2X1_486/CTRL POR2X1_526/Y 0.02fF
C57885 PAND2X1_552/B POR2X1_90/Y 0.03fF
C57886 PAND2X1_182/a_16_344# POR2X1_55/Y 0.02fF
C57887 POR2X1_68/A POR2X1_562/B 0.01fF
C57888 POR2X1_55/Y PAND2X1_509/CTRL 0.14fF
C57889 POR2X1_96/Y POR2X1_29/A 0.03fF
C57890 POR2X1_334/B PAND2X1_96/B 0.11fF
C57891 PAND2X1_209/A PAND2X1_162/CTRL 0.00fF
C57892 POR2X1_335/A PAND2X1_69/A 0.03fF
C57893 PAND2X1_702/O POR2X1_42/Y 0.04fF
C57894 POR2X1_186/a_16_28# POR2X1_188/A 0.03fF
C57895 POR2X1_176/CTRL2 POR2X1_312/Y 0.01fF
C57896 PAND2X1_48/B PAND2X1_747/O 0.01fF
C57897 POR2X1_763/Y PAND2X1_149/A 0.03fF
C57898 POR2X1_22/A POR2X1_36/CTRL 0.10fF
C57899 PAND2X1_506/CTRL2 POR2X1_239/Y 0.01fF
C57900 POR2X1_664/Y PAND2X1_60/B 0.40fF
C57901 POR2X1_376/B POR2X1_153/Y 0.12fF
C57902 POR2X1_26/CTRL VDD 0.00fF
C57903 POR2X1_137/Y POR2X1_572/B 3.03fF
C57904 PAND2X1_56/Y POR2X1_335/B 0.03fF
C57905 POR2X1_327/Y POR2X1_405/a_16_28# 0.03fF
C57906 VDD POR2X1_675/Y 0.01fF
C57907 POR2X1_12/CTRL POR2X1_3/B 0.01fF
C57908 D_GATE_662 POR2X1_544/O 0.05fF
C57909 POR2X1_204/O PAND2X1_79/Y 0.00fF
C57910 PAND2X1_275/CTRL PAND2X1_60/B 0.03fF
C57911 POR2X1_42/Y PAND2X1_843/Y 0.99fF
C57912 POR2X1_130/Y POR2X1_318/A 0.03fF
C57913 POR2X1_68/A PAND2X1_747/CTRL 0.01fF
C57914 POR2X1_654/B POR2X1_113/B 0.02fF
C57915 POR2X1_523/Y POR2X1_844/O 0.01fF
C57916 PAND2X1_736/O PAND2X1_853/B 0.01fF
C57917 D_GATE_222 PAND2X1_173/CTRL 0.03fF
C57918 PAND2X1_6/Y POR2X1_140/CTRL 0.06fF
C57919 POR2X1_60/A POR2X1_373/a_16_28# 0.00fF
C57920 POR2X1_41/B PAND2X1_849/B 0.02fF
C57921 POR2X1_293/Y PAND2X1_510/B 0.03fF
C57922 POR2X1_124/B PAND2X1_96/B 0.93fF
C57923 POR2X1_357/a_56_344# POR2X1_353/Y 0.01fF
C57924 POR2X1_775/A PAND2X1_60/B 0.04fF
C57925 POR2X1_99/B POR2X1_750/B 0.05fF
C57926 POR2X1_390/B POR2X1_337/CTRL 0.00fF
C57927 PAND2X1_524/CTRL POR2X1_456/B 0.00fF
C57928 PAND2X1_716/a_56_28# POR2X1_73/Y 0.00fF
C57929 PAND2X1_484/m4_208_n4# PAND2X1_41/B 0.12fF
C57930 POR2X1_544/B VDD 0.22fF
C57931 PAND2X1_659/Y PAND2X1_660/B 0.12fF
C57932 POR2X1_541/O PAND2X1_32/B 0.01fF
C57933 POR2X1_60/Y PAND2X1_338/O 0.02fF
C57934 POR2X1_52/A INPUT_1 0.06fF
C57935 PAND2X1_836/m4_208_n4# POR2X1_823/m4_208_n4# 0.05fF
C57936 POR2X1_343/Y POR2X1_296/B 0.14fF
C57937 POR2X1_220/Y POR2X1_507/A 0.07fF
C57938 POR2X1_383/A POR2X1_35/Y 0.03fF
C57939 PAND2X1_735/a_16_344# POR2X1_153/Y 0.02fF
C57940 POR2X1_119/Y PAND2X1_803/A 0.03fF
C57941 POR2X1_36/B POR2X1_582/CTRL2 0.01fF
C57942 POR2X1_164/Y PAND2X1_776/a_16_344# 0.01fF
C57943 PAND2X1_480/O POR2X1_96/A 0.05fF
C57944 POR2X1_83/a_16_28# PAND2X1_35/Y 0.02fF
C57945 PAND2X1_392/CTRL2 POR2X1_55/Y 0.18fF
C57946 PAND2X1_854/O PAND2X1_856/B 0.03fF
C57947 PAND2X1_630/a_16_344# POR2X1_7/A 0.02fF
C57948 POR2X1_722/A POR2X1_502/A 0.08fF
C57949 POR2X1_621/m4_208_n4# POR2X1_622/m4_208_n4# 0.05fF
C57950 PAND2X1_60/B POR2X1_112/Y 0.04fF
C57951 POR2X1_407/Y POR2X1_770/a_76_344# 0.00fF
C57952 POR2X1_356/A POR2X1_782/CTRL 0.21fF
C57953 PAND2X1_56/Y PAND2X1_368/O 0.09fF
C57954 PAND2X1_20/A POR2X1_725/CTRL2 0.01fF
C57955 POR2X1_93/CTRL POR2X1_283/A 0.01fF
C57956 PAND2X1_675/A PAND2X1_181/a_76_28# 0.02fF
C57957 POR2X1_519/O POR2X1_43/B 0.02fF
C57958 PAND2X1_20/A POR2X1_500/CTRL2 0.01fF
C57959 PAND2X1_94/A PAND2X1_283/CTRL 0.06fF
C57960 POR2X1_52/A POR2X1_153/Y 0.14fF
C57961 POR2X1_222/Y POR2X1_456/B 0.03fF
C57962 POR2X1_417/CTRL POR2X1_7/A 0.03fF
C57963 POR2X1_569/A POR2X1_576/Y 0.02fF
C57964 POR2X1_741/Y POR2X1_675/Y 0.03fF
C57965 POR2X1_391/Y POR2X1_276/Y 0.09fF
C57966 PAND2X1_69/A PAND2X1_133/CTRL2 0.01fF
C57967 PAND2X1_659/Y POR2X1_821/O 0.01fF
C57968 POR2X1_57/A PAND2X1_656/A 0.03fF
C57969 POR2X1_228/Y POR2X1_318/A 0.10fF
C57970 POR2X1_96/A PAND2X1_716/B 0.27fF
C57971 POR2X1_857/B POR2X1_227/O 0.09fF
C57972 POR2X1_775/A POR2X1_332/O 0.01fF
C57973 POR2X1_307/B PAND2X1_304/O 0.01fF
C57974 INPUT_1 PAND2X1_49/O 0.02fF
C57975 POR2X1_328/CTRL2 INPUT_4 0.03fF
C57976 POR2X1_249/Y PAND2X1_69/A 0.01fF
C57977 POR2X1_687/A POR2X1_730/a_16_28# 0.02fF
C57978 POR2X1_174/B POR2X1_568/A 18.95fF
C57979 POR2X1_60/A PAND2X1_332/Y 0.54fF
C57980 POR2X1_122/m4_208_n4# POR2X1_822/m4_208_n4# 0.15fF
C57981 POR2X1_15/a_16_28# POR2X1_7/A 0.03fF
C57982 POR2X1_614/A POR2X1_833/A 1.01fF
C57983 POR2X1_416/B PAND2X1_620/Y 0.03fF
C57984 PAND2X1_48/B PAND2X1_48/A 0.12fF
C57985 POR2X1_677/O POR2X1_77/Y 0.02fF
C57986 POR2X1_65/A POR2X1_416/B 0.78fF
C57987 POR2X1_567/A PAND2X1_280/O 0.02fF
C57988 PAND2X1_631/A PAND2X1_515/CTRL 0.06fF
C57989 POR2X1_731/a_16_28# POR2X1_726/Y -0.00fF
C57990 PAND2X1_860/A POR2X1_32/A 0.03fF
C57991 POR2X1_532/A POR2X1_456/B 0.06fF
C57992 PAND2X1_55/Y POR2X1_722/O 0.09fF
C57993 POR2X1_228/a_16_28# POR2X1_294/B 0.00fF
C57994 POR2X1_294/B POR2X1_342/O 0.01fF
C57995 POR2X1_107/Y POR2X1_103/Y 0.00fF
C57996 PAND2X1_625/CTRL2 POR2X1_294/A 0.00fF
C57997 POR2X1_21/CTRL POR2X1_260/A 0.01fF
C57998 PAND2X1_610/CTRL2 POR2X1_293/Y 0.01fF
C57999 PAND2X1_20/A PAND2X1_125/O 0.02fF
C58000 POR2X1_156/a_16_28# POR2X1_155/Y 0.03fF
C58001 POR2X1_83/B POR2X1_698/Y 0.01fF
C58002 PAND2X1_86/Y PAND2X1_60/B 0.00fF
C58003 POR2X1_566/A POR2X1_568/B 0.10fF
C58004 PAND2X1_6/Y POR2X1_593/a_56_344# 0.00fF
C58005 POR2X1_57/A PAND2X1_348/A 0.07fF
C58006 POR2X1_287/B POR2X1_717/B 0.00fF
C58007 POR2X1_734/O PAND2X1_60/B 0.02fF
C58008 PAND2X1_94/A POR2X1_569/A 0.07fF
C58009 POR2X1_560/a_16_28# POR2X1_294/B 0.01fF
C58010 PAND2X1_461/O POR2X1_413/Y 0.00fF
C58011 PAND2X1_652/CTRL2 PAND2X1_652/A 0.03fF
C58012 POR2X1_608/a_76_344# PAND2X1_56/A 0.00fF
C58013 PAND2X1_849/B PAND2X1_100/CTRL2 0.01fF
C58014 POR2X1_391/O POR2X1_260/A 0.01fF
C58015 POR2X1_394/A POR2X1_91/Y 0.12fF
C58016 POR2X1_329/A PAND2X1_561/CTRL2 0.01fF
C58017 POR2X1_540/A POR2X1_552/CTRL2 0.03fF
C58018 POR2X1_778/CTRL POR2X1_717/B 0.01fF
C58019 PAND2X1_349/A PAND2X1_301/a_16_344# 0.00fF
C58020 POR2X1_383/A PAND2X1_701/CTRL 0.01fF
C58021 POR2X1_416/B POR2X1_481/a_56_344# 0.00fF
C58022 POR2X1_592/Y POR2X1_832/B 0.04fF
C58023 POR2X1_54/Y INPUT_3 0.11fF
C58024 POR2X1_456/B POR2X1_704/a_76_344# 0.01fF
C58025 POR2X1_64/CTRL VDD 0.00fF
C58026 PAND2X1_476/A PAND2X1_734/CTRL2 0.00fF
C58027 POR2X1_43/Y POR2X1_236/Y 1.55fF
C58028 POR2X1_42/Y POR2X1_589/O 0.01fF
C58029 PAND2X1_787/A PAND2X1_357/CTRL 0.00fF
C58030 POR2X1_4/Y POR2X1_816/A 0.03fF
C58031 POR2X1_719/O POR2X1_722/A 0.01fF
C58032 PAND2X1_841/B PAND2X1_840/Y 0.05fF
C58033 POR2X1_153/O POR2X1_96/B 0.02fF
C58034 D_INPUT_1 POR2X1_4/Y 1.38fF
C58035 PAND2X1_323/CTRL POR2X1_702/A 0.00fF
C58036 POR2X1_168/A POR2X1_170/B 0.01fF
C58037 PAND2X1_641/Y PAND2X1_650/A 0.00fF
C58038 POR2X1_286/B POR2X1_655/A 0.01fF
C58039 POR2X1_677/Y POR2X1_423/Y 0.00fF
C58040 POR2X1_52/O POR2X1_599/A 0.04fF
C58041 POR2X1_841/CTRL POR2X1_841/B 0.03fF
C58042 POR2X1_293/Y POR2X1_387/O 0.10fF
C58043 POR2X1_554/B POR2X1_218/Y 0.28fF
C58044 POR2X1_244/Y POR2X1_260/A 0.03fF
C58045 POR2X1_7/A PAND2X1_716/B 0.03fF
C58046 PAND2X1_545/Y POR2X1_394/A 0.03fF
C58047 POR2X1_814/A PAND2X1_310/m4_208_n4# 0.09fF
C58048 POR2X1_20/B POR2X1_626/CTRL 0.01fF
C58049 POR2X1_257/A POR2X1_109/O 0.10fF
C58050 POR2X1_588/O POR2X1_587/Y 0.01fF
C58051 POR2X1_119/Y PAND2X1_560/a_16_344# 0.06fF
C58052 POR2X1_799/CTRL POR2X1_652/A 0.00fF
C58053 POR2X1_111/Y PAND2X1_348/A 0.02fF
C58054 POR2X1_707/CTRL2 PAND2X1_48/A 0.08fF
C58055 PAND2X1_326/O PAND2X1_324/Y 0.17fF
C58056 POR2X1_13/A PAND2X1_242/Y 0.20fF
C58057 POR2X1_782/O POR2X1_782/B 0.00fF
C58058 POR2X1_416/B POR2X1_136/CTRL 0.01fF
C58059 POR2X1_244/Y POR2X1_363/A 0.01fF
C58060 PAND2X1_301/CTRL POR2X1_75/Y 0.01fF
C58061 PAND2X1_301/O POR2X1_300/Y 0.00fF
C58062 POR2X1_48/A PAND2X1_606/CTRL 0.01fF
C58063 POR2X1_750/CTRL2 POR2X1_39/B 0.03fF
C58064 POR2X1_57/A POR2X1_43/CTRL 0.01fF
C58065 POR2X1_390/B POR2X1_188/Y 0.00fF
C58066 PAND2X1_213/Y PAND2X1_169/O 0.05fF
C58067 PAND2X1_737/B PAND2X1_737/CTRL2 0.01fF
C58068 POR2X1_16/A PAND2X1_341/B 0.07fF
C58069 POR2X1_703/A POR2X1_540/Y 0.15fF
C58070 POR2X1_623/Y POR2X1_94/A 0.00fF
C58071 POR2X1_435/CTRL2 PAND2X1_72/A 0.01fF
C58072 POR2X1_624/Y POR2X1_296/B 0.12fF
C58073 POR2X1_604/Y POR2X1_604/O 0.01fF
C58074 POR2X1_394/A POR2X1_109/Y 0.05fF
C58075 POR2X1_54/Y POR2X1_78/A 0.03fF
C58076 PAND2X1_90/A PAND2X1_42/a_76_28# 0.02fF
C58077 POR2X1_257/A POR2X1_427/a_16_28# 0.03fF
C58078 PAND2X1_243/B POR2X1_826/a_16_28# 0.01fF
C58079 POR2X1_441/Y POR2X1_72/B 0.05fF
C58080 POR2X1_698/Y PAND2X1_709/O 0.05fF
C58081 PAND2X1_275/O POR2X1_76/B 0.15fF
C58082 POR2X1_520/O POR2X1_383/Y 0.01fF
C58083 POR2X1_111/Y PAND2X1_631/A 0.03fF
C58084 POR2X1_344/Y POR2X1_359/O 0.01fF
C58085 PAND2X1_290/CTRL PAND2X1_94/A 0.01fF
C58086 POR2X1_408/Y POR2X1_387/O 0.60fF
C58087 POR2X1_814/Y VDD 0.10fF
C58088 PAND2X1_267/CTRL2 POR2X1_102/Y 0.01fF
C58089 POR2X1_777/B POR2X1_475/CTRL 0.30fF
C58090 POR2X1_849/A POR2X1_66/A 0.03fF
C58091 PAND2X1_860/A POR2X1_184/Y 0.02fF
C58092 PAND2X1_68/CTRL D_INPUT_0 0.01fF
C58093 POR2X1_622/B VDD 0.14fF
C58094 POR2X1_567/A POR2X1_566/CTRL 0.04fF
C58095 POR2X1_633/O PAND2X1_90/Y 0.08fF
C58096 PAND2X1_499/CTRL POR2X1_20/B 0.03fF
C58097 PAND2X1_271/O POR2X1_330/Y 0.04fF
C58098 POR2X1_709/A POR2X1_752/Y 0.03fF
C58099 POR2X1_685/A PAND2X1_681/CTRL2 0.04fF
C58100 POR2X1_265/Y POR2X1_7/Y 0.03fF
C58101 PAND2X1_651/Y PAND2X1_860/A 0.05fF
C58102 POR2X1_96/A POR2X1_250/Y 0.10fF
C58103 PAND2X1_862/Y PAND2X1_865/A 0.00fF
C58104 POR2X1_37/Y POR2X1_29/A 0.06fF
C58105 POR2X1_96/CTRL POR2X1_77/Y 0.01fF
C58106 POR2X1_60/A PAND2X1_97/O 0.03fF
C58107 POR2X1_4/Y POR2X1_620/B 1.28fF
C58108 PAND2X1_612/B POR2X1_734/A 0.03fF
C58109 POR2X1_115/CTRL POR2X1_554/B 0.01fF
C58110 POR2X1_860/CTRL2 PAND2X1_72/A 0.01fF
C58111 POR2X1_257/A PAND2X1_210/CTRL2 0.00fF
C58112 POR2X1_265/O POR2X1_40/Y 0.01fF
C58113 POR2X1_119/Y POR2X1_150/a_76_344# 0.04fF
C58114 POR2X1_91/CTRL POR2X1_91/Y 0.01fF
C58115 POR2X1_57/A PAND2X1_193/Y 2.28fF
C58116 PAND2X1_330/O POR2X1_385/Y 0.17fF
C58117 PAND2X1_94/A PAND2X1_72/A 0.03fF
C58118 PAND2X1_678/m4_208_n4# PAND2X1_579/m4_208_n4# 0.15fF
C58119 POR2X1_661/Y POR2X1_78/A 0.03fF
C58120 POR2X1_586/Y PAND2X1_638/B 0.00fF
C58121 POR2X1_260/B PAND2X1_597/CTRL 0.01fF
C58122 POR2X1_142/CTRL POR2X1_669/B 0.04fF
C58123 POR2X1_471/O POR2X1_471/A 0.16fF
C58124 PAND2X1_301/CTRL PAND2X1_332/Y 0.02fF
C58125 PAND2X1_357/a_16_344# POR2X1_39/B 0.01fF
C58126 PAND2X1_486/CTRL2 POR2X1_484/Y 0.01fF
C58127 PAND2X1_689/a_16_344# POR2X1_121/B 0.03fF
C58128 PAND2X1_420/CTRL POR2X1_590/A 0.01fF
C58129 POR2X1_257/A POR2X1_516/B 0.02fF
C58130 POR2X1_159/O POR2X1_669/B 0.09fF
C58131 PAND2X1_645/O POR2X1_600/Y 0.02fF
C58132 POR2X1_66/B POR2X1_267/CTRL 0.01fF
C58133 POR2X1_659/A VDD 0.12fF
C58134 PAND2X1_65/B PAND2X1_237/CTRL 0.01fF
C58135 PAND2X1_859/CTRL2 POR2X1_37/Y 0.06fF
C58136 POR2X1_188/A POR2X1_858/a_56_344# 0.00fF
C58137 POR2X1_406/Y PAND2X1_560/a_76_28# 0.04fF
C58138 POR2X1_814/B POR2X1_288/CTRL2 0.03fF
C58139 POR2X1_496/CTRL2 POR2X1_55/Y 0.01fF
C58140 POR2X1_814/A POR2X1_685/B 0.08fF
C58141 POR2X1_68/A POR2X1_554/B 0.03fF
C58142 POR2X1_662/O POR2X1_220/Y 0.01fF
C58143 PAND2X1_645/CTRL POR2X1_48/A 0.01fF
C58144 PAND2X1_463/O PAND2X1_58/A 0.03fF
C58145 POR2X1_660/CTRL POR2X1_660/A 0.01fF
C58146 PAND2X1_251/a_76_28# POR2X1_362/B 0.01fF
C58147 POR2X1_96/A POR2X1_490/Y 0.02fF
C58148 POR2X1_628/Y POR2X1_42/Y 0.03fF
C58149 PAND2X1_58/A POR2X1_593/B 0.04fF
C58150 POR2X1_428/Y POR2X1_700/CTRL2 0.01fF
C58151 PAND2X1_810/a_16_344# PAND2X1_221/Y 0.02fF
C58152 PAND2X1_362/A PAND2X1_363/Y 0.02fF
C58153 PAND2X1_200/O POR2X1_72/B 0.01fF
C58154 PAND2X1_404/Y POR2X1_290/Y 0.03fF
C58155 POR2X1_568/B POR2X1_568/CTRL2 0.13fF
C58156 PAND2X1_221/CTRL2 PAND2X1_192/Y 0.01fF
C58157 POR2X1_60/A PAND2X1_562/B 0.08fF
C58158 POR2X1_383/A PAND2X1_52/CTRL2 0.10fF
C58159 PAND2X1_609/CTRL POR2X1_294/B 0.01fF
C58160 POR2X1_624/Y POR2X1_501/O 0.02fF
C58161 POR2X1_491/O POR2X1_72/B 0.01fF
C58162 POR2X1_458/Y PAND2X1_300/O 0.03fF
C58163 PAND2X1_57/B POR2X1_66/A 0.22fF
C58164 POR2X1_487/CTRL PAND2X1_738/Y 0.23fF
C58165 PAND2X1_23/Y POR2X1_260/B 5.73fF
C58166 POR2X1_65/A POR2X1_487/Y 0.06fF
C58167 PAND2X1_644/Y POR2X1_7/B 0.03fF
C58168 PAND2X1_277/a_56_28# PAND2X1_57/B 0.00fF
C58169 POR2X1_864/A POR2X1_686/CTRL 0.00fF
C58170 POR2X1_504/Y POR2X1_750/B 0.03fF
C58171 POR2X1_689/A PAND2X1_590/CTRL 0.01fF
C58172 PAND2X1_39/B POR2X1_513/Y 0.03fF
C58173 POR2X1_424/Y POR2X1_90/Y 0.03fF
C58174 D_INPUT_3 PAND2X1_618/O 0.00fF
C58175 POR2X1_69/A PAND2X1_340/O 0.09fF
C58176 POR2X1_423/CTRL INPUT_0 0.03fF
C58177 POR2X1_428/Y PAND2X1_711/CTRL2 0.06fF
C58178 POR2X1_13/CTRL POR2X1_102/Y 0.05fF
C58179 PAND2X1_474/Y POR2X1_60/A 0.02fF
C58180 POR2X1_42/a_76_344# INPUT_3 0.09fF
C58181 POR2X1_14/Y VDD 2.67fF
C58182 POR2X1_341/A POR2X1_573/A 0.02fF
C58183 PAND2X1_735/Y POR2X1_498/Y 0.05fF
C58184 POR2X1_642/CTRL2 POR2X1_66/A 0.01fF
C58185 PAND2X1_390/Y POR2X1_5/Y 0.05fF
C58186 POR2X1_45/Y PAND2X1_205/A 0.03fF
C58187 POR2X1_541/B PAND2X1_60/B 0.13fF
C58188 POR2X1_41/B PAND2X1_804/a_56_28# 0.00fF
C58189 PAND2X1_496/O D_INPUT_0 0.02fF
C58190 POR2X1_97/A POR2X1_579/Y 0.03fF
C58191 POR2X1_65/A PAND2X1_192/Y 0.03fF
C58192 POR2X1_21/CTRL2 D_INPUT_5 0.03fF
C58193 POR2X1_850/CTRL2 PAND2X1_39/B 0.16fF
C58194 PAND2X1_39/B POR2X1_205/A 0.07fF
C58195 POR2X1_355/B POR2X1_149/A 0.21fF
C58196 POR2X1_13/A POR2X1_60/A 1.11fF
C58197 PAND2X1_814/a_56_28# INPUT_3 0.00fF
C58198 POR2X1_78/A PAND2X1_322/O 0.04fF
C58199 PAND2X1_668/CTRL POR2X1_83/B 0.01fF
C58200 PAND2X1_631/CTRL2 POR2X1_48/A 0.01fF
C58201 PAND2X1_116/CTRL POR2X1_106/Y 0.03fF
C58202 POR2X1_514/Y D_INPUT_0 0.06fF
C58203 POR2X1_28/CTRL D_INPUT_1 0.01fF
C58204 PAND2X1_500/O POR2X1_497/Y 0.05fF
C58205 PAND2X1_500/a_16_344# PAND2X1_499/Y 0.10fF
C58206 POR2X1_681/Y POR2X1_38/Y 0.02fF
C58207 PAND2X1_26/A PAND2X1_26/O 0.02fF
C58208 POR2X1_62/CTRL POR2X1_29/A 0.03fF
C58209 POR2X1_355/B POR2X1_209/a_16_28# 0.03fF
C58210 POR2X1_389/A POR2X1_655/A 0.03fF
C58211 PAND2X1_48/B POR2X1_274/a_16_28# 0.02fF
C58212 POR2X1_138/O POR2X1_296/B 0.02fF
C58213 POR2X1_13/A PAND2X1_554/a_16_344# 0.02fF
C58214 PAND2X1_116/O PAND2X1_787/Y 0.04fF
C58215 POR2X1_653/CTRL POR2X1_653/B 0.01fF
C58216 PAND2X1_217/B PAND2X1_598/CTRL 0.01fF
C58217 POR2X1_454/A POR2X1_318/A 0.12fF
C58218 POR2X1_96/A PAND2X1_78/a_56_28# 0.00fF
C58219 POR2X1_791/Y VDD 0.00fF
C58220 POR2X1_460/A PAND2X1_22/a_76_28# 0.04fF
C58221 POR2X1_523/Y POR2X1_669/B 0.05fF
C58222 PAND2X1_700/CTRL PAND2X1_90/Y 0.04fF
C58223 D_INPUT_5 POR2X1_1/O 0.03fF
C58224 PAND2X1_685/CTRL POR2X1_60/A 0.01fF
C58225 PAND2X1_58/A POR2X1_565/CTRL2 0.01fF
C58226 POR2X1_301/CTRL POR2X1_590/A 0.01fF
C58227 POR2X1_65/A PAND2X1_738/Y 0.05fF
C58228 POR2X1_97/A POR2X1_317/Y 0.03fF
C58229 PAND2X1_652/Y PAND2X1_557/A 0.00fF
C58230 POR2X1_750/B POR2X1_586/O 0.01fF
C58231 POR2X1_637/B VDD 0.42fF
C58232 PAND2X1_787/Y PAND2X1_140/Y 0.05fF
C58233 POR2X1_76/O POR2X1_274/B 0.01fF
C58234 POR2X1_76/CTRL2 POR2X1_553/A 0.01fF
C58235 POR2X1_493/CTRL2 POR2X1_493/A 0.01fF
C58236 PAND2X1_793/Y PAND2X1_579/CTRL2 0.01fF
C58237 PAND2X1_96/B PAND2X1_595/CTRL2 0.01fF
C58238 PAND2X1_235/O PAND2X1_55/Y 0.01fF
C58239 PAND2X1_23/Y POR2X1_242/CTRL2 0.00fF
C58240 POR2X1_49/Y PAND2X1_149/O 0.03fF
C58241 PAND2X1_833/O POR2X1_511/Y 0.04fF
C58242 PAND2X1_592/Y POR2X1_40/Y 0.06fF
C58243 PAND2X1_798/B POR2X1_102/Y 0.05fF
C58244 POR2X1_490/Y POR2X1_7/A 0.01fF
C58245 INPUT_0 POR2X1_666/A 0.00fF
C58246 PAND2X1_90/A PAND2X1_46/CTRL 0.01fF
C58247 PAND2X1_54/CTRL2 INPUT_0 -0.00fF
C58248 POR2X1_178/CTRL2 POR2X1_60/A 0.03fF
C58249 PAND2X1_65/B POR2X1_483/CTRL 0.01fF
C58250 PAND2X1_96/B POR2X1_792/CTRL 0.01fF
C58251 PAND2X1_78/CTRL2 PAND2X1_794/B 0.01fF
C58252 POR2X1_20/B PAND2X1_182/B 0.00fF
C58253 POR2X1_260/B POR2X1_520/A 0.03fF
C58254 POR2X1_102/Y POR2X1_759/Y 0.03fF
C58255 POR2X1_471/A POR2X1_703/Y 0.03fF
C58256 POR2X1_445/A POR2X1_703/A 0.07fF
C58257 POR2X1_378/Y POR2X1_376/Y 0.32fF
C58258 PAND2X1_93/B POR2X1_201/Y 0.01fF
C58259 POR2X1_62/O POR2X1_94/A 0.01fF
C58260 PAND2X1_20/A POR2X1_513/Y 0.03fF
C58261 POR2X1_775/A POR2X1_750/B 0.05fF
C58262 POR2X1_832/A PAND2X1_591/O 0.08fF
C58263 POR2X1_232/CTRL POR2X1_5/Y 0.03fF
C58264 POR2X1_669/B POR2X1_93/A 0.17fF
C58265 POR2X1_376/Y POR2X1_7/B 0.03fF
C58266 POR2X1_14/Y PAND2X1_32/B 0.03fF
C58267 POR2X1_101/A POR2X1_99/Y 0.57fF
C58268 POR2X1_537/CTRL2 POR2X1_260/B 0.03fF
C58269 POR2X1_567/B POR2X1_738/A 0.05fF
C58270 PAND2X1_48/B POR2X1_193/Y 0.03fF
C58271 POR2X1_346/B POR2X1_629/CTRL 0.00fF
C58272 PAND2X1_661/B POR2X1_60/A 0.03fF
C58273 POR2X1_60/A PAND2X1_643/Y 0.03fF
C58274 POR2X1_505/Y PAND2X1_6/A 0.02fF
C58275 POR2X1_356/A POR2X1_781/CTRL2 -0.00fF
C58276 POR2X1_355/B VDD 1.44fF
C58277 POR2X1_650/A POR2X1_572/B 0.03fF
C58278 PAND2X1_472/B VDD 0.04fF
C58279 POR2X1_346/a_16_28# POR2X1_346/A 0.03fF
C58280 POR2X1_164/CTRL POR2X1_72/B 0.01fF
C58281 POR2X1_866/A POR2X1_260/A 0.03fF
C58282 POR2X1_861/A POR2X1_554/B 0.04fF
C58283 POR2X1_500/A POR2X1_844/B 0.27fF
C58284 POR2X1_444/A POR2X1_568/Y 0.05fF
C58285 POR2X1_748/A POR2X1_90/Y 0.06fF
C58286 POR2X1_29/A POR2X1_408/Y 0.12fF
C58287 PAND2X1_725/Y PAND2X1_162/m4_208_n4# 0.08fF
C58288 POR2X1_198/O POR2X1_61/Y 0.02fF
C58289 PAND2X1_732/O PAND2X1_731/A 0.06fF
C58290 POR2X1_405/CTRL PAND2X1_32/B 0.01fF
C58291 PAND2X1_126/CTRL POR2X1_29/A 0.04fF
C58292 D_INPUT_0 POR2X1_576/CTRL2 0.01fF
C58293 PAND2X1_556/B POR2X1_7/B 0.05fF
C58294 POR2X1_750/B POR2X1_112/Y 0.05fF
C58295 POR2X1_13/A POR2X1_684/CTRL2 0.00fF
C58296 POR2X1_504/Y PAND2X1_631/CTRL 0.02fF
C58297 POR2X1_78/A POR2X1_148/B 0.01fF
C58298 POR2X1_681/Y POR2X1_153/Y 0.17fF
C58299 PAND2X1_269/O POR2X1_39/B 0.05fF
C58300 POR2X1_669/B PAND2X1_720/CTRL 0.01fF
C58301 POR2X1_669/B PAND2X1_559/CTRL2 0.01fF
C58302 POR2X1_406/Y POR2X1_406/O 0.00fF
C58303 PAND2X1_57/B PAND2X1_751/O 0.03fF
C58304 POR2X1_407/A PAND2X1_679/O 0.02fF
C58305 POR2X1_110/Y POR2X1_424/Y 0.16fF
C58306 PAND2X1_254/a_76_28# POR2X1_511/Y 0.01fF
C58307 POR2X1_55/Y VDD 4.03fF
C58308 PAND2X1_449/Y POR2X1_376/B 0.01fF
C58309 PAND2X1_658/A POR2X1_236/Y 0.03fF
C58310 POR2X1_814/B POR2X1_513/Y 0.03fF
C58311 POR2X1_779/A PAND2X1_65/B 0.61fF
C58312 POR2X1_750/B D_INPUT_6 0.03fF
C58313 POR2X1_647/B POR2X1_294/A 0.03fF
C58314 PAND2X1_73/Y POR2X1_796/A 0.03fF
C58315 PAND2X1_41/B POR2X1_194/CTRL 0.01fF
C58316 POR2X1_66/B PAND2X1_60/B 2.84fF
C58317 PAND2X1_20/A POR2X1_366/A 0.03fF
C58318 POR2X1_38/Y PAND2X1_733/CTRL 0.01fF
C58319 PAND2X1_638/a_76_28# POR2X1_752/Y 0.02fF
C58320 PAND2X1_550/O PAND2X1_546/Y 0.01fF
C58321 POR2X1_96/A PAND2X1_243/B 0.03fF
C58322 POR2X1_62/Y POR2X1_88/CTRL2 0.01fF
C58323 INPUT_3 POR2X1_4/Y 0.55fF
C58324 PAND2X1_811/O PAND2X1_808/Y 0.00fF
C58325 POR2X1_13/O POR2X1_13/Y 0.01fF
C58326 PAND2X1_536/CTRL VDD -0.00fF
C58327 POR2X1_60/A PAND2X1_535/a_16_344# 0.02fF
C58328 PAND2X1_572/O POR2X1_72/B 0.01fF
C58329 PAND2X1_48/B PAND2X1_516/O 0.01fF
C58330 PAND2X1_850/Y POR2X1_275/Y 0.05fF
C58331 POR2X1_809/A POR2X1_260/B 0.02fF
C58332 POR2X1_407/Y PAND2X1_597/CTRL 0.01fF
C58333 PAND2X1_381/Y POR2X1_260/A 0.03fF
C58334 POR2X1_60/A POR2X1_9/m4_208_n4# 0.08fF
C58335 PAND2X1_131/O POR2X1_130/Y 0.01fF
C58336 POR2X1_693/Y POR2X1_697/a_16_28# 0.01fF
C58337 PAND2X1_258/CTRL POR2X1_186/B 0.02fF
C58338 PAND2X1_460/CTRL2 POR2X1_5/Y 0.01fF
C58339 POR2X1_60/A PAND2X1_510/B 0.04fF
C58340 POR2X1_188/A PAND2X1_60/B 0.03fF
C58341 PAND2X1_691/Y POR2X1_102/Y 0.03fF
C58342 POR2X1_78/A POR2X1_175/B 0.01fF
C58343 POR2X1_41/B PAND2X1_852/CTRL2 0.01fF
C58344 POR2X1_697/Y POR2X1_46/Y 0.03fF
C58345 PAND2X1_118/CTRL POR2X1_502/A 0.00fF
C58346 POR2X1_140/B PAND2X1_516/CTRL2 0.00fF
C58347 POR2X1_325/A POR2X1_513/Y 0.03fF
C58348 POR2X1_750/B POR2X1_162/Y 2.97fF
C58349 POR2X1_673/A D_INPUT_1 0.16fF
C58350 POR2X1_174/O POR2X1_174/A 0.03fF
C58351 POR2X1_169/m4_208_n4# PAND2X1_91/m4_208_n4# 0.13fF
C58352 PAND2X1_181/CTRL POR2X1_40/Y 0.01fF
C58353 POR2X1_366/Y POR2X1_193/A 0.03fF
C58354 POR2X1_193/A POR2X1_294/B 0.60fF
C58355 PAND2X1_471/CTRL PAND2X1_464/Y 0.01fF
C58356 POR2X1_579/Y POR2X1_294/B 0.03fF
C58357 POR2X1_830/Y POR2X1_675/Y 0.02fF
C58358 POR2X1_820/A POR2X1_408/Y 0.02fF
C58359 POR2X1_416/B PAND2X1_634/CTRL2 0.01fF
C58360 PAND2X1_65/B PAND2X1_153/O 0.02fF
C58361 POR2X1_832/Y POR2X1_512/O 0.02fF
C58362 POR2X1_236/Y POR2X1_73/Y 0.17fF
C58363 PAND2X1_23/Y POR2X1_284/O 0.01fF
C58364 PAND2X1_614/O POR2X1_283/A 0.01fF
C58365 POR2X1_68/A POR2X1_214/O 0.09fF
C58366 PAND2X1_855/O VDD 0.00fF
C58367 PAND2X1_23/Y POR2X1_205/Y 0.03fF
C58368 POR2X1_853/A POR2X1_578/Y 0.01fF
C58369 POR2X1_130/A PAND2X1_767/O 0.04fF
C58370 PAND2X1_499/CTRL2 POR2X1_283/A 0.01fF
C58371 POR2X1_532/A PAND2X1_131/CTRL2 0.01fF
C58372 POR2X1_139/Y POR2X1_514/Y 0.01fF
C58373 POR2X1_32/A PAND2X1_708/CTRL2 0.03fF
C58374 PAND2X1_23/Y PAND2X1_55/Y 5.05fF
C58375 POR2X1_572/B POR2X1_294/B 0.23fF
C58376 POR2X1_791/B VDD 0.25fF
C58377 PAND2X1_674/CTRL2 POR2X1_732/B 0.13fF
C58378 PAND2X1_543/CTRL2 POR2X1_142/Y 0.01fF
C58379 POR2X1_845/CTRL2 POR2X1_5/Y 0.01fF
C58380 POR2X1_795/O POR2X1_795/B 0.02fF
C58381 POR2X1_128/CTRL2 PAND2X1_96/B 0.01fF
C58382 POR2X1_415/A POR2X1_39/B 0.08fF
C58383 POR2X1_32/A PAND2X1_156/A 0.05fF
C58384 POR2X1_860/A POR2X1_101/Y 0.03fF
C58385 POR2X1_773/CTRL POR2X1_734/A 0.05fF
C58386 POR2X1_355/B PAND2X1_32/B 0.03fF
C58387 PAND2X1_23/Y POR2X1_363/O 0.01fF
C58388 POR2X1_52/Y PAND2X1_364/B 0.02fF
C58389 POR2X1_519/Y POR2X1_42/Y 0.01fF
C58390 PAND2X1_254/CTRL PAND2X1_6/A 0.03fF
C58391 POR2X1_786/Y POR2X1_404/Y 0.07fF
C58392 POR2X1_220/Y POR2X1_788/B 0.01fF
C58393 PAND2X1_57/B POR2X1_532/A 10.06fF
C58394 POR2X1_50/O POR2X1_158/B 0.00fF
C58395 INPUT_4 POR2X1_3/CTRL 0.06fF
C58396 PAND2X1_65/B POR2X1_598/CTRL2 0.01fF
C58397 PAND2X1_23/Y POR2X1_402/A 0.70fF
C58398 PAND2X1_65/B POR2X1_407/CTRL 0.01fF
C58399 POR2X1_325/A POR2X1_366/A 0.03fF
C58400 POR2X1_366/Y POR2X1_614/A 0.07fF
C58401 POR2X1_614/A POR2X1_294/B 8.25fF
C58402 POR2X1_567/B PAND2X1_167/O 0.02fF
C58403 POR2X1_326/O PAND2X1_41/B 0.10fF
C58404 POR2X1_446/B POR2X1_736/A 0.02fF
C58405 POR2X1_68/A POR2X1_800/A 0.07fF
C58406 POR2X1_510/B VDD 0.10fF
C58407 POR2X1_366/Y POR2X1_317/Y 0.03fF
C58408 PAND2X1_6/Y POR2X1_740/Y 0.07fF
C58409 POR2X1_198/O POR2X1_35/Y 0.01fF
C58410 POR2X1_93/CTRL POR2X1_55/Y 0.01fF
C58411 INPUT_0 POR2X1_530/Y 0.17fF
C58412 POR2X1_730/Y POR2X1_653/B 0.05fF
C58413 POR2X1_96/A PAND2X1_243/a_76_28# 0.02fF
C58414 POR2X1_29/Y POR2X1_42/Y 0.03fF
C58415 PAND2X1_371/O POR2X1_68/B 0.01fF
C58416 PAND2X1_48/B POR2X1_731/O 0.06fF
C58417 POR2X1_179/Y VDD 0.01fF
C58418 POR2X1_123/A INPUT_0 0.05fF
C58419 POR2X1_278/A POR2X1_46/Y 0.76fF
C58420 INPUT_1 POR2X1_625/CTRL 0.07fF
C58421 POR2X1_16/A PAND2X1_340/O 0.00fF
C58422 POR2X1_220/Y PAND2X1_163/CTRL 0.00fF
C58423 PAND2X1_339/Y POR2X1_56/Y 0.03fF
C58424 POR2X1_544/A POR2X1_544/a_16_28# 0.03fF
C58425 PAND2X1_632/A INPUT_0 0.05fF
C58426 POR2X1_55/Y PAND2X1_344/CTRL2 0.00fF
C58427 POR2X1_477/A PAND2X1_96/B 0.03fF
C58428 POR2X1_38/B POR2X1_294/B 0.23fF
C58429 POR2X1_260/B POR2X1_711/Y 0.07fF
C58430 PAND2X1_23/Y POR2X1_407/Y 0.00fF
C58431 VDD POR2X1_7/CTRL2 -0.00fF
C58432 PAND2X1_804/B PAND2X1_175/B 0.90fF
C58433 PAND2X1_470/CTRL2 POR2X1_43/B 0.03fF
C58434 POR2X1_207/A POR2X1_260/A 0.03fF
C58435 POR2X1_78/A POR2X1_4/Y 0.10fF
C58436 POR2X1_419/Y PAND2X1_156/A 0.01fF
C58437 POR2X1_594/O POR2X1_385/Y 0.10fF
C58438 PAND2X1_6/Y POR2X1_796/CTRL 0.01fF
C58439 POR2X1_502/A PAND2X1_63/B 0.01fF
C58440 POR2X1_157/CTRL POR2X1_36/B 0.01fF
C58441 PAND2X1_825/O PAND2X1_57/B 0.03fF
C58442 PAND2X1_857/CTRL POR2X1_83/B 0.01fF
C58443 PAND2X1_232/CTRL VDD 0.00fF
C58444 POR2X1_68/A POR2X1_702/A 0.03fF
C58445 POR2X1_203/O POR2X1_579/Y 0.00fF
C58446 POR2X1_725/Y POR2X1_722/Y 0.02fF
C58447 POR2X1_579/Y PAND2X1_111/B 0.03fF
C58448 PAND2X1_89/a_16_344# PAND2X1_60/B 0.01fF
C58449 POR2X1_281/O VDD 0.00fF
C58450 POR2X1_327/Y POR2X1_828/Y 0.09fF
C58451 POR2X1_60/A PAND2X1_199/O 0.03fF
C58452 D_INPUT_1 POR2X1_816/A 0.03fF
C58453 PAND2X1_422/O POR2X1_294/B 0.08fF
C58454 PAND2X1_115/CTRL POR2X1_283/A 0.02fF
C58455 POR2X1_559/Y POR2X1_68/B 0.01fF
C58456 POR2X1_302/Y POR2X1_260/A 0.02fF
C58457 POR2X1_865/B POR2X1_114/CTRL2 0.12fF
C58458 POR2X1_81/A PAND2X1_573/B 0.13fF
C58459 POR2X1_128/a_16_28# POR2X1_128/B 0.02fF
C58460 POR2X1_52/A POR2X1_51/B 0.01fF
C58461 PAND2X1_784/O POR2X1_245/Y 0.04fF
C58462 POR2X1_518/O POR2X1_667/A 0.01fF
C58463 POR2X1_782/A PAND2X1_747/CTRL 0.01fF
C58464 PAND2X1_777/a_16_344# POR2X1_39/B 0.02fF
C58465 POR2X1_57/A POR2X1_183/Y 0.03fF
C58466 POR2X1_619/A PAND2X1_6/A 0.03fF
C58467 PAND2X1_434/m4_208_n4# POR2X1_39/B 0.15fF
C58468 POR2X1_241/B POR2X1_568/B 0.03fF
C58469 POR2X1_68/A PAND2X1_670/CTRL 0.01fF
C58470 PAND2X1_469/B PAND2X1_787/A 0.12fF
C58471 PAND2X1_476/A POR2X1_40/Y 0.03fF
C58472 POR2X1_464/CTRL POR2X1_186/B 0.12fF
C58473 POR2X1_809/A PAND2X1_679/a_16_344# 0.01fF
C58474 POR2X1_93/CTRL2 D_INPUT_3 0.04fF
C58475 PAND2X1_632/a_56_28# INPUT_0 0.00fF
C58476 PAND2X1_635/CTRL INPUT_6 0.00fF
C58477 POR2X1_119/Y PAND2X1_240/O 0.04fF
C58478 POR2X1_362/B POR2X1_737/A 0.93fF
C58479 PAND2X1_486/CTRL PAND2X1_726/B 0.06fF
C58480 PAND2X1_473/Y PAND2X1_853/B 0.11fF
C58481 POR2X1_140/B POR2X1_574/A 0.00fF
C58482 POR2X1_637/CTRL2 PAND2X1_72/A 0.01fF
C58483 POR2X1_614/A POR2X1_203/O 0.01fF
C58484 POR2X1_614/A PAND2X1_111/B 0.03fF
C58485 POR2X1_136/CTRL POR2X1_136/Y 0.01fF
C58486 PAND2X1_862/B POR2X1_153/Y 0.03fF
C58487 POR2X1_73/CTRL2 PAND2X1_6/A -0.01fF
C58488 PAND2X1_6/Y POR2X1_348/O 0.02fF
C58489 POR2X1_516/Y PAND2X1_840/Y 0.05fF
C58490 POR2X1_537/CTRL2 PAND2X1_55/Y 0.02fF
C58491 POR2X1_760/A POR2X1_250/Y 0.36fF
C58492 POR2X1_367/CTRL POR2X1_191/Y 0.11fF
C58493 POR2X1_488/Y PAND2X1_363/a_76_28# 0.04fF
C58494 POR2X1_134/Y PAND2X1_348/Y 0.03fF
C58495 POR2X1_824/CTRL POR2X1_236/Y 0.01fF
C58496 POR2X1_38/B PAND2X1_111/B 0.00fF
C58497 PAND2X1_199/B VDD 0.03fF
C58498 POR2X1_197/CTRL2 POR2X1_99/B 0.00fF
C58499 POR2X1_596/A POR2X1_770/a_16_28# 0.02fF
C58500 POR2X1_137/Y POR2X1_361/CTRL 0.00fF
C58501 POR2X1_772/a_16_28# POR2X1_294/B 0.08fF
C58502 INPUT_1 POR2X1_790/B 0.03fF
C58503 PAND2X1_632/B PAND2X1_6/A 0.02fF
C58504 PAND2X1_11/Y PAND2X1_72/A 0.04fF
C58505 POR2X1_208/A PAND2X1_88/Y 0.01fF
C58506 POR2X1_778/B PAND2X1_103/CTRL2 0.09fF
C58507 POR2X1_119/Y PAND2X1_659/O 0.19fF
C58508 POR2X1_322/Y PAND2X1_168/CTRL 0.00fF
C58509 PAND2X1_465/O POR2X1_77/Y 0.03fF
C58510 PAND2X1_429/Y PAND2X1_3/B 0.02fF
C58511 POR2X1_40/Y PAND2X1_327/CTRL2 0.03fF
C58512 POR2X1_46/Y POR2X1_117/Y 0.07fF
C58513 POR2X1_502/A POR2X1_383/CTRL 0.30fF
C58514 POR2X1_52/A POR2X1_150/CTRL2 0.00fF
C58515 POR2X1_23/Y POR2X1_485/a_16_28# 0.02fF
C58516 POR2X1_222/Y POR2X1_259/B 0.03fF
C58517 POR2X1_8/Y PAND2X1_341/a_76_28# 0.05fF
C58518 PAND2X1_577/a_16_344# PAND2X1_569/Y 0.02fF
C58519 POR2X1_532/A POR2X1_707/Y 0.03fF
C58520 POR2X1_707/CTRL POR2X1_407/Y 0.01fF
C58521 PAND2X1_73/Y POR2X1_863/A 0.03fF
C58522 PAND2X1_191/Y PAND2X1_730/A 0.00fF
C58523 POR2X1_307/Y POR2X1_512/O 0.01fF
C58524 PAND2X1_432/CTRL PAND2X1_72/A 0.01fF
C58525 POR2X1_717/Y PAND2X1_48/A 0.15fF
C58526 POR2X1_311/O POR2X1_142/Y 0.09fF
C58527 POR2X1_501/B POR2X1_260/A 0.01fF
C58528 PAND2X1_150/CTRL2 POR2X1_260/A 0.01fF
C58529 POR2X1_730/Y POR2X1_596/A 0.03fF
C58530 PAND2X1_673/CTRL2 POR2X1_416/B 0.01fF
C58531 POR2X1_740/Y POR2X1_195/O 0.04fF
C58532 POR2X1_771/A POR2X1_532/A 0.02fF
C58533 PAND2X1_93/B POR2X1_458/Y 0.07fF
C58534 PAND2X1_865/Y PAND2X1_468/O 0.00fF
C58535 POR2X1_567/A POR2X1_579/Y 0.05fF
C58536 POR2X1_83/B POR2X1_825/Y 0.16fF
C58537 PAND2X1_6/Y POR2X1_774/A 0.31fF
C58538 POR2X1_464/Y POR2X1_552/A 0.01fF
C58539 D_INPUT_7 PAND2X1_3/A 0.00fF
C58540 POR2X1_49/Y POR2X1_167/Y 0.08fF
C58541 POR2X1_271/A POR2X1_73/Y 0.01fF
C58542 POR2X1_655/CTRL2 POR2X1_646/Y 0.01fF
C58543 POR2X1_399/A POR2X1_119/Y 0.02fF
C58544 POR2X1_551/CTRL2 POR2X1_854/B 0.16fF
C58545 POR2X1_725/Y POR2X1_151/CTRL2 0.02fF
C58546 PAND2X1_651/Y PAND2X1_156/A 0.05fF
C58547 POR2X1_71/CTRL2 POR2X1_91/Y 0.01fF
C58548 POR2X1_383/A POR2X1_463/Y 0.03fF
C58549 POR2X1_760/A POR2X1_490/Y 0.03fF
C58550 PAND2X1_358/O PAND2X1_351/Y 0.02fF
C58551 PAND2X1_65/B POR2X1_768/A 0.03fF
C58552 POR2X1_837/A POR2X1_202/B 0.22fF
C58553 POR2X1_520/a_16_28# POR2X1_520/A 0.05fF
C58554 PAND2X1_394/CTRL2 PAND2X1_88/Y 0.01fF
C58555 POR2X1_252/Y POR2X1_253/Y 0.01fF
C58556 POR2X1_610/Y POR2X1_472/B 0.01fF
C58557 POR2X1_614/A POR2X1_567/A 0.13fF
C58558 POR2X1_346/B POR2X1_61/CTRL2 0.00fF
C58559 POR2X1_647/B POR2X1_286/B 0.03fF
C58560 PAND2X1_319/B PAND2X1_357/O 0.02fF
C58561 PAND2X1_163/CTRL2 POR2X1_210/A 0.03fF
C58562 POR2X1_38/Y PAND2X1_716/B 0.07fF
C58563 POR2X1_305/a_16_28# POR2X1_416/B 0.00fF
C58564 POR2X1_680/O PAND2X1_652/A 0.01fF
C58565 POR2X1_793/a_76_344# PAND2X1_52/B 0.01fF
C58566 POR2X1_157/CTRL2 POR2X1_416/B 0.00fF
C58567 POR2X1_96/A PAND2X1_862/CTRL 0.10fF
C58568 POR2X1_661/CTRL2 POR2X1_661/A 0.05fF
C58569 POR2X1_322/Y PAND2X1_325/O 0.02fF
C58570 POR2X1_571/Y POR2X1_318/A 0.03fF
C58571 PAND2X1_55/Y POR2X1_711/Y 0.07fF
C58572 POR2X1_329/A PAND2X1_361/CTRL2 0.04fF
C58573 POR2X1_730/Y POR2X1_449/A 0.03fF
C58574 POR2X1_647/B POR2X1_862/Y 0.01fF
C58575 POR2X1_51/B POR2X1_3/B 0.12fF
C58576 POR2X1_803/O POR2X1_796/Y 0.02fF
C58577 POR2X1_156/CTRL2 POR2X1_162/Y 0.01fF
C58578 PAND2X1_217/CTRL PAND2X1_576/B 0.03fF
C58579 POR2X1_257/A PAND2X1_776/Y 0.03fF
C58580 POR2X1_312/CTRL POR2X1_77/Y 0.10fF
C58581 INPUT_1 POR2X1_673/B 0.01fF
C58582 PAND2X1_441/O PAND2X1_52/B 0.05fF
C58583 PAND2X1_535/Y PAND2X1_863/A 0.10fF
C58584 PAND2X1_356/a_16_344# PAND2X1_354/Y 0.01fF
C58585 POR2X1_57/A PAND2X1_850/Y 0.02fF
C58586 PAND2X1_388/Y PAND2X1_352/Y 0.01fF
C58587 POR2X1_740/Y PAND2X1_52/B 0.03fF
C58588 PAND2X1_481/CTRL POR2X1_507/A 0.04fF
C58589 PAND2X1_341/Y POR2X1_394/A 0.05fF
C58590 POR2X1_48/A POR2X1_415/A 0.07fF
C58591 POR2X1_814/B PAND2X1_234/a_16_344# 0.02fF
C58592 PAND2X1_551/A PAND2X1_326/CTRL 0.01fF
C58593 POR2X1_40/O POR2X1_25/Y 0.01fF
C58594 POR2X1_270/Y POR2X1_446/B 0.03fF
C58595 PAND2X1_447/O POR2X1_420/Y 0.00fF
C58596 POR2X1_78/A POR2X1_78/Y 0.04fF
C58597 POR2X1_600/Y POR2X1_601/CTRL2 0.01fF
C58598 POR2X1_796/CTRL PAND2X1_52/B 0.01fF
C58599 POR2X1_854/a_16_28# POR2X1_567/B 0.07fF
C58600 POR2X1_7/A PAND2X1_508/B 0.04fF
C58601 PAND2X1_267/Y PAND2X1_576/B 0.05fF
C58602 POR2X1_241/B POR2X1_341/A 0.11fF
C58603 POR2X1_14/Y PAND2X1_9/Y 0.04fF
C58604 POR2X1_60/A POR2X1_813/CTRL 0.07fF
C58605 POR2X1_760/A PAND2X1_205/Y 0.02fF
C58606 PAND2X1_858/CTRL POR2X1_129/Y 0.01fF
C58607 PAND2X1_716/B POR2X1_153/Y 0.03fF
C58608 POR2X1_612/A VDD 0.00fF
C58609 POR2X1_864/A POR2X1_783/a_76_344# 0.01fF
C58610 POR2X1_333/A POR2X1_443/A 0.03fF
C58611 PAND2X1_6/Y POR2X1_87/B 0.09fF
C58612 POR2X1_411/B POR2X1_72/B 0.10fF
C58613 PAND2X1_853/B POR2X1_7/Y 0.03fF
C58614 POR2X1_383/A POR2X1_736/A 0.10fF
C58615 INPUT_6 PAND2X1_52/B 1.51fF
C58616 POR2X1_78/A POR2X1_266/O 0.01fF
C58617 POR2X1_818/CTRL2 POR2X1_734/A 0.16fF
C58618 POR2X1_60/A POR2X1_437/O 0.10fF
C58619 POR2X1_150/Y POR2X1_106/Y 0.03fF
C58620 POR2X1_76/B POR2X1_804/A 0.05fF
C58621 POR2X1_77/CTRL2 POR2X1_40/Y 0.03fF
C58622 POR2X1_96/A POR2X1_329/A 0.09fF
C58623 PAND2X1_76/Y POR2X1_271/B 0.06fF
C58624 PAND2X1_175/B PAND2X1_332/Y 0.03fF
C58625 POR2X1_14/Y POR2X1_818/Y 0.03fF
C58626 POR2X1_65/A PAND2X1_838/B 0.06fF
C58627 POR2X1_78/B POR2X1_318/CTRL 0.03fF
C58628 POR2X1_863/A PAND2X1_173/CTRL2 0.00fF
C58629 POR2X1_479/O POR2X1_66/A 0.02fF
C58630 POR2X1_673/Y PAND2X1_529/a_56_28# 0.00fF
C58631 PAND2X1_207/CTRL POR2X1_40/Y 0.00fF
C58632 POR2X1_471/A PAND2X1_90/Y 0.03fF
C58633 POR2X1_411/B PAND2X1_756/O 0.03fF
C58634 POR2X1_150/Y PAND2X1_580/B 0.03fF
C58635 PAND2X1_245/CTRL2 POR2X1_296/B 0.00fF
C58636 POR2X1_769/O POR2X1_769/B 0.00fF
C58637 PAND2X1_489/O PAND2X1_557/A 0.02fF
C58638 POR2X1_859/O INPUT_0 0.03fF
C58639 POR2X1_113/a_16_28# POR2X1_768/A 0.02fF
C58640 PAND2X1_20/A POR2X1_35/O 0.01fF
C58641 POR2X1_49/Y POR2X1_848/A 0.07fF
C58642 POR2X1_121/B POR2X1_288/O 0.07fF
C58643 POR2X1_482/a_16_28# POR2X1_60/A 0.01fF
C58644 POR2X1_60/A POR2X1_29/A 0.07fF
C58645 PAND2X1_206/A PAND2X1_206/O -0.00fF
C58646 POR2X1_411/B PAND2X1_216/CTRL 0.01fF
C58647 PAND2X1_222/A PAND2X1_593/O 0.00fF
C58648 POR2X1_669/B PAND2X1_706/CTRL2 0.04fF
C58649 POR2X1_461/Y POR2X1_790/O 0.00fF
C58650 PAND2X1_97/Y PAND2X1_339/Y 0.00fF
C58651 PAND2X1_73/Y PAND2X1_531/a_76_28# 0.01fF
C58652 PAND2X1_850/Y POR2X1_589/CTRL 0.04fF
C58653 POR2X1_424/Y POR2X1_424/O 0.02fF
C58654 PAND2X1_61/Y D_INPUT_0 0.07fF
C58655 POR2X1_774/A PAND2X1_52/B 0.03fF
C58656 POR2X1_43/B PAND2X1_449/CTRL 0.01fF
C58657 POR2X1_111/CTRL2 PAND2X1_717/A -0.00fF
C58658 POR2X1_807/A POR2X1_807/a_56_344# 0.00fF
C58659 PAND2X1_838/CTRL POR2X1_42/Y 0.01fF
C58660 POR2X1_66/B PAND2X1_88/CTRL2 0.01fF
C58661 PAND2X1_446/a_76_28# POR2X1_417/Y 0.07fF
C58662 PAND2X1_859/B PAND2X1_98/O 0.02fF
C58663 PAND2X1_9/Y POR2X1_55/Y 1.45fF
C58664 POR2X1_682/CTRL POR2X1_32/A 0.01fF
C58665 PAND2X1_85/Y POR2X1_66/A 0.09fF
C58666 PAND2X1_73/Y POR2X1_456/CTRL 0.01fF
C58667 POR2X1_66/B POR2X1_254/A 0.03fF
C58668 POR2X1_466/A POR2X1_480/A 0.10fF
C58669 PAND2X1_52/O POR2X1_532/A 0.03fF
C58670 PAND2X1_645/O PAND2X1_644/Y 0.05fF
C58671 POR2X1_78/A PAND2X1_52/Y 0.00fF
C58672 POR2X1_441/Y POR2X1_438/CTRL2 0.01fF
C58673 POR2X1_476/A VDD 0.18fF
C58674 POR2X1_66/B POR2X1_750/B 0.12fF
C58675 POR2X1_96/A POR2X1_437/a_56_344# 0.00fF
C58676 PAND2X1_404/A D_INPUT_0 0.01fF
C58677 POR2X1_554/B PAND2X1_96/B 0.00fF
C58678 PAND2X1_412/a_16_344# POR2X1_590/A 0.02fF
C58679 PAND2X1_469/Y PAND2X1_717/A 0.09fF
C58680 POR2X1_502/A POR2X1_567/B 0.05fF
C58681 POR2X1_66/B POR2X1_461/CTRL 0.01fF
C58682 POR2X1_127/CTRL VDD -0.00fF
C58683 POR2X1_329/A POR2X1_7/A 0.07fF
C58684 POR2X1_814/B PAND2X1_585/CTRL 0.01fF
C58685 POR2X1_14/Y POR2X1_236/CTRL2 0.00fF
C58686 POR2X1_413/A PAND2X1_646/CTRL2 0.01fF
C58687 POR2X1_188/A POR2X1_750/B 0.06fF
C58688 PAND2X1_223/O POR2X1_283/Y 0.02fF
C58689 PAND2X1_65/B POR2X1_267/O 0.03fF
C58690 PAND2X1_835/Y POR2X1_411/B 0.05fF
C58691 PAND2X1_651/Y POR2X1_490/O 0.02fF
C58692 POR2X1_120/CTRL POR2X1_78/A 0.01fF
C58693 INPUT_3 POR2X1_816/A 0.03fF
C58694 POR2X1_66/B PAND2X1_13/O 0.08fF
C58695 POR2X1_102/Y POR2X1_666/A 0.06fF
C58696 POR2X1_639/A POR2X1_639/CTRL 0.01fF
C58697 PAND2X1_117/CTRL POR2X1_493/A 0.01fF
C58698 POR2X1_260/B POR2X1_733/A 0.05fF
C58699 PAND2X1_499/Y PAND2X1_573/B 0.25fF
C58700 PAND2X1_501/B POR2X1_498/Y 0.00fF
C58701 INPUT_3 D_INPUT_1 0.22fF
C58702 POR2X1_445/A POR2X1_455/A 0.48fF
C58703 POR2X1_663/B PAND2X1_69/A 0.03fF
C58704 POR2X1_334/B POR2X1_260/B 0.25fF
C58705 POR2X1_56/B POR2X1_48/A 0.03fF
C58706 POR2X1_631/O POR2X1_193/Y 0.01fF
C58707 PAND2X1_658/O PAND2X1_474/A 0.15fF
C58708 POR2X1_257/A POR2X1_248/CTRL 0.05fF
C58709 POR2X1_515/CTRL PAND2X1_20/A 0.01fF
C58710 POR2X1_660/Y PAND2X1_57/B 0.03fF
C58711 POR2X1_224/a_56_344# POR2X1_32/A 0.00fF
C58712 POR2X1_841/a_16_28# POR2X1_804/A 0.02fF
C58713 POR2X1_376/B POR2X1_72/B 3.72fF
C58714 PAND2X1_262/O PAND2X1_41/B 0.01fF
C58715 PAND2X1_794/O PAND2X1_580/B 0.00fF
C58716 POR2X1_376/Y POR2X1_750/B 0.00fF
C58717 PAND2X1_859/A PAND2X1_859/O 0.00fF
C58718 POR2X1_800/O D_GATE_865 0.01fF
C58719 POR2X1_857/B POR2X1_97/A 4.80fF
C58720 POR2X1_490/Y PAND2X1_218/A 0.01fF
C58721 POR2X1_814/A POR2X1_772/O 0.02fF
C58722 POR2X1_60/A POR2X1_256/CTRL 0.01fF
C58723 POR2X1_457/CTRL POR2X1_370/Y 0.04fF
C58724 PAND2X1_56/Y POR2X1_270/Y 0.07fF
C58725 POR2X1_150/Y PAND2X1_349/A 0.03fF
C58726 POR2X1_814/B PAND2X1_395/O 0.02fF
C58727 PAND2X1_557/A POR2X1_250/CTRL 0.03fF
C58728 POR2X1_411/B PAND2X1_570/B 0.03fF
C58729 POR2X1_48/A PAND2X1_725/A 0.01fF
C58730 POR2X1_590/A POR2X1_208/CTRL 0.01fF
C58731 PAND2X1_65/B PAND2X1_423/O 0.01fF
C58732 POR2X1_667/A POR2X1_46/Y 0.07fF
C58733 POR2X1_602/B POR2X1_130/A 0.02fF
C58734 POR2X1_458/CTRL PAND2X1_69/A 0.06fF
C58735 POR2X1_343/Y POR2X1_717/B 0.02fF
C58736 POR2X1_681/Y POR2X1_591/Y 0.03fF
C58737 PAND2X1_717/A POR2X1_394/A 0.03fF
C58738 PAND2X1_580/O PAND2X1_771/Y 0.04fF
C58739 PAND2X1_247/O POR2X1_283/A 0.02fF
C58740 POR2X1_590/A POR2X1_294/B 1.17fF
C58741 POR2X1_859/A PAND2X1_225/a_16_344# 0.02fF
C58742 POR2X1_23/Y PAND2X1_457/O 0.04fF
C58743 PAND2X1_241/CTRL POR2X1_83/B 0.01fF
C58744 POR2X1_813/O POR2X1_7/A 0.01fF
C58745 POR2X1_67/Y PAND2X1_789/a_16_344# 0.01fF
C58746 POR2X1_301/a_16_28# POR2X1_301/A 0.05fF
C58747 PAND2X1_23/Y POR2X1_174/A 0.03fF
C58748 PAND2X1_58/A PAND2X1_369/CTRL 0.01fF
C58749 POR2X1_52/A PAND2X1_465/CTRL2 0.03fF
C58750 PAND2X1_640/CTRL D_INPUT_0 0.00fF
C58751 POR2X1_859/A POR2X1_750/B 2.49fF
C58752 POR2X1_411/B PAND2X1_383/a_76_28# 0.01fF
C58753 PAND2X1_352/A PAND2X1_357/Y 0.02fF
C58754 POR2X1_155/Y POR2X1_750/B 0.01fF
C58755 POR2X1_43/B POR2X1_89/Y 0.01fF
C58756 PAND2X1_633/Y POR2X1_826/Y 0.01fF
C58757 POR2X1_630/O PAND2X1_96/B 0.07fF
C58758 PAND2X1_649/O POR2X1_32/A 0.01fF
C58759 POR2X1_602/CTRL2 PAND2X1_60/B 0.01fF
C58760 POR2X1_47/O POR2X1_83/B 0.16fF
C58761 POR2X1_669/B PAND2X1_551/A 0.03fF
C58762 POR2X1_476/A PAND2X1_32/B 0.01fF
C58763 D_GATE_662 POR2X1_78/A 0.21fF
C58764 POR2X1_13/A PAND2X1_140/O 0.17fF
C58765 POR2X1_294/Y PAND2X1_69/A 0.02fF
C58766 PAND2X1_90/A PAND2X1_9/O 0.03fF
C58767 PAND2X1_808/Y PAND2X1_772/CTRL 0.01fF
C58768 POR2X1_476/O POR2X1_121/Y 0.01fF
C58769 POR2X1_52/A POR2X1_251/A 0.21fF
C58770 PAND2X1_73/Y PAND2X1_744/CTRL 0.01fF
C58771 POR2X1_828/Y PAND2X1_760/CTRL2 0.00fF
C58772 PAND2X1_553/A POR2X1_106/Y 0.01fF
C58773 POR2X1_55/O PAND2X1_6/A 0.02fF
C58774 POR2X1_37/Y POR2X1_380/a_16_28# 0.03fF
C58775 POR2X1_52/A POR2X1_72/B 0.28fF
C58776 POR2X1_814/A POR2X1_113/B 1.95fF
C58777 POR2X1_288/CTRL2 PAND2X1_32/B 0.10fF
C58778 PAND2X1_139/B PAND2X1_139/a_76_28# 0.04fF
C58779 POR2X1_8/Y POR2X1_20/B 0.09fF
C58780 PAND2X1_229/CTRL2 POR2X1_231/B 0.00fF
C58781 POR2X1_78/B POR2X1_403/Y 0.01fF
C58782 PAND2X1_94/A PAND2X1_24/CTRL 0.01fF
C58783 POR2X1_511/Y VDD 0.23fF
C58784 POR2X1_254/Y PAND2X1_65/B 0.04fF
C58785 POR2X1_175/CTRL2 POR2X1_566/A 0.16fF
C58786 POR2X1_117/O POR2X1_46/Y 0.00fF
C58787 POR2X1_83/B POR2X1_518/Y 0.03fF
C58788 POR2X1_524/Y VDD 0.10fF
C58789 POR2X1_866/A POR2X1_725/Y 0.07fF
C58790 POR2X1_657/CTRL2 POR2X1_112/Y 0.01fF
C58791 PAND2X1_472/A POR2X1_83/B 0.09fF
C58792 POR2X1_72/B POR2X1_152/A 0.03fF
C58793 POR2X1_78/A D_INPUT_1 0.13fF
C58794 POR2X1_57/A PAND2X1_722/CTRL 0.01fF
C58795 POR2X1_186/Y POR2X1_785/A 0.04fF
C58796 POR2X1_43/B POR2X1_497/O 0.02fF
C58797 PAND2X1_639/B PAND2X1_639/CTRL 0.01fF
C58798 POR2X1_777/B POR2X1_575/B 0.15fF
C58799 PAND2X1_73/Y PAND2X1_518/O 0.05fF
C58800 POR2X1_383/A POR2X1_270/Y 0.55fF
C58801 POR2X1_114/B POR2X1_830/O 0.01fF
C58802 POR2X1_46/Y PAND2X1_712/B 0.02fF
C58803 PAND2X1_79/Y POR2X1_296/B 0.03fF
C58804 POR2X1_669/B POR2X1_425/Y 0.03fF
C58805 POR2X1_45/Y PAND2X1_558/Y 0.05fF
C58806 POR2X1_659/O POR2X1_750/B 0.10fF
C58807 POR2X1_78/B POR2X1_502/A 0.21fF
C58808 POR2X1_472/B POR2X1_559/A 0.00fF
C58809 POR2X1_618/O POR2X1_5/Y 0.01fF
C58810 PAND2X1_865/CTRL POR2X1_23/Y 0.00fF
C58811 POR2X1_78/A POR2X1_724/A 0.27fF
C58812 POR2X1_829/A PAND2X1_687/Y 0.02fF
C58813 POR2X1_65/Y PAND2X1_358/A 0.08fF
C58814 POR2X1_680/Y PAND2X1_192/O 0.02fF
C58815 POR2X1_614/A POR2X1_800/O 0.01fF
C58816 PAND2X1_687/CTRL2 POR2X1_597/Y 0.03fF
C58817 POR2X1_866/A POR2X1_596/O 0.11fF
C58818 POR2X1_114/B POR2X1_734/A 0.07fF
C58819 POR2X1_338/O POR2X1_97/A 0.01fF
C58820 POR2X1_186/Y PAND2X1_504/O 0.06fF
C58821 POR2X1_590/A PAND2X1_111/B 0.04fF
C58822 POR2X1_52/A PAND2X1_520/CTRL2 0.01fF
C58823 POR2X1_834/Y POR2X1_644/Y 0.30fF
C58824 POR2X1_309/O POR2X1_387/Y 0.05fF
C58825 POR2X1_83/B PAND2X1_168/CTRL 0.01fF
C58826 PAND2X1_272/O POR2X1_569/A 0.04fF
C58827 PAND2X1_833/CTRL POR2X1_495/Y 0.01fF
C58828 PAND2X1_205/B PAND2X1_735/Y 0.02fF
C58829 PAND2X1_119/CTRL2 POR2X1_654/B 0.06fF
C58830 PAND2X1_412/CTRL2 PAND2X1_32/B 0.00fF
C58831 POR2X1_102/Y POR2X1_530/Y 0.01fF
C58832 PAND2X1_731/CTRL PAND2X1_738/B 0.00fF
C58833 PAND2X1_496/CTRL INPUT_0 0.03fF
C58834 POR2X1_68/A POR2X1_830/A 0.03fF
C58835 POR2X1_760/a_16_28# POR2X1_7/B 0.01fF
C58836 POR2X1_72/B PAND2X1_186/O 0.05fF
C58837 POR2X1_614/A POR2X1_807/A 0.03fF
C58838 POR2X1_254/Y POR2X1_231/O 0.03fF
C58839 POR2X1_65/CTRL2 POR2X1_39/B 0.14fF
C58840 PAND2X1_281/O POR2X1_647/B 0.01fF
C58841 D_INPUT_0 PAND2X1_690/CTRL 0.01fF
C58842 POR2X1_625/Y POR2X1_7/B 0.07fF
C58843 POR2X1_350/Y PAND2X1_65/B 0.02fF
C58844 PAND2X1_402/B POR2X1_14/Y 0.01fF
C58845 POR2X1_649/B POR2X1_734/A 0.02fF
C58846 PAND2X1_632/A POR2X1_102/Y 0.03fF
C58847 POR2X1_43/B PAND2X1_735/CTRL2 0.03fF
C58848 POR2X1_212/A POR2X1_192/B 0.03fF
C58849 POR2X1_833/A POR2X1_66/A 0.07fF
C58850 POR2X1_137/B PAND2X1_134/O 0.16fF
C58851 POR2X1_355/B POR2X1_149/Y 0.29fF
C58852 POR2X1_135/Y PAND2X1_469/B 0.03fF
C58853 POR2X1_734/A PAND2X1_518/a_16_344# 0.04fF
C58854 PAND2X1_94/A POR2X1_35/a_76_344# 0.01fF
C58855 POR2X1_57/A PAND2X1_211/A 0.03fF
C58856 POR2X1_65/A PAND2X1_724/O 0.01fF
C58857 POR2X1_121/B POR2X1_101/Y 0.05fF
C58858 POR2X1_38/B POR2X1_226/Y 0.02fF
C58859 POR2X1_356/A PAND2X1_524/a_56_28# 0.00fF
C58860 POR2X1_564/Y POR2X1_366/Y 0.07fF
C58861 POR2X1_287/B POR2X1_68/B 0.19fF
C58862 POR2X1_83/B PAND2X1_196/O 0.01fF
C58863 POR2X1_416/B PAND2X1_464/B 0.07fF
C58864 PAND2X1_6/Y PAND2X1_627/O 0.03fF
C58865 POR2X1_68/A POR2X1_471/O 0.02fF
C58866 POR2X1_596/A PAND2X1_597/O 0.02fF
C58867 POR2X1_278/Y PAND2X1_798/B 0.07fF
C58868 POR2X1_130/A POR2X1_712/Y 0.07fF
C58869 POR2X1_814/B PAND2X1_757/CTRL 0.01fF
C58870 PAND2X1_65/B POR2X1_341/Y 0.01fF
C58871 PAND2X1_129/CTRL POR2X1_68/B 0.01fF
C58872 POR2X1_857/B POR2X1_294/B 0.05fF
C58873 POR2X1_513/Y VDD 0.41fF
C58874 POR2X1_814/A POR2X1_768/A 0.03fF
C58875 POR2X1_158/O POR2X1_257/A 0.01fF
C58876 PAND2X1_85/Y POR2X1_532/A 0.00fF
C58877 PAND2X1_633/O POR2X1_278/A 0.00fF
C58878 POR2X1_52/A POR2X1_617/a_56_344# 0.00fF
C58879 POR2X1_734/B PAND2X1_48/A 0.01fF
C58880 POR2X1_60/A PAND2X1_301/CTRL2 0.00fF
C58881 POR2X1_546/A POR2X1_844/B 0.28fF
C58882 PAND2X1_324/O VDD 0.00fF
C58883 POR2X1_761/Y PAND2X1_687/Y 0.06fF
C58884 POR2X1_219/B VDD 0.54fF
C58885 POR2X1_614/A POR2X1_786/a_16_28# 0.09fF
C58886 POR2X1_60/O POR2X1_497/Y 0.01fF
C58887 POR2X1_46/Y PAND2X1_546/CTRL2 0.01fF
C58888 POR2X1_66/A PAND2X1_18/B 0.01fF
C58889 POR2X1_811/CTRL POR2X1_294/A 0.08fF
C58890 POR2X1_270/Y POR2X1_370/a_76_344# 0.00fF
C58891 POR2X1_230/O PAND2X1_338/B 0.01fF
C58892 PAND2X1_684/a_16_344# POR2X1_296/B 0.05fF
C58893 POR2X1_334/B PAND2X1_55/Y 0.26fF
C58894 POR2X1_68/A POR2X1_555/a_16_28# 0.02fF
C58895 POR2X1_68/B PAND2X1_8/Y 1.75fF
C58896 POR2X1_480/A POR2X1_478/B 0.07fF
C58897 POR2X1_567/B POR2X1_188/Y 0.05fF
C58898 PAND2X1_643/Y PAND2X1_719/O 0.07fF
C58899 POR2X1_140/B POR2X1_193/A 0.03fF
C58900 PAND2X1_483/O POR2X1_482/Y 0.01fF
C58901 POR2X1_220/Y POR2X1_556/Y 0.09fF
C58902 POR2X1_550/A POR2X1_5/Y 0.02fF
C58903 POR2X1_205/A VDD 0.00fF
C58904 POR2X1_280/a_16_28# POR2X1_236/Y 0.04fF
C58905 PAND2X1_96/B POR2X1_190/Y 0.15fF
C58906 POR2X1_41/B POR2X1_111/CTRL2 0.03fF
C58907 PAND2X1_90/A POR2X1_559/Y 0.01fF
C58908 POR2X1_236/Y PAND2X1_656/A 0.07fF
C58909 PAND2X1_48/B PAND2X1_146/a_56_28# 0.00fF
C58910 POR2X1_37/Y PAND2X1_500/CTRL2 0.03fF
C58911 POR2X1_614/A POR2X1_565/B -0.02fF
C58912 POR2X1_660/Y POR2X1_512/CTRL2 0.01fF
C58913 POR2X1_20/CTRL2 POR2X1_68/B 0.01fF
C58914 POR2X1_215/a_76_344# PAND2X1_88/Y 0.00fF
C58915 POR2X1_57/A POR2X1_96/A 0.30fF
C58916 PAND2X1_90/Y POR2X1_741/m4_208_n4# 0.05fF
C58917 POR2X1_859/A POR2X1_750/O 0.10fF
C58918 POR2X1_78/A POR2X1_620/B 0.03fF
C58919 PAND2X1_651/Y PAND2X1_242/CTRL2 0.00fF
C58920 PAND2X1_682/CTRL POR2X1_68/A 0.00fF
C58921 VDD POR2X1_366/A 0.40fF
C58922 PAND2X1_20/A PAND2X1_527/CTRL 0.02fF
C58923 POR2X1_565/B POR2X1_38/B 0.15fF
C58924 PAND2X1_117/a_16_344# PAND2X1_32/B 0.02fF
C58925 POR2X1_853/A POR2X1_364/A 0.03fF
C58926 POR2X1_43/B POR2X1_56/Y 0.06fF
C58927 POR2X1_236/Y PAND2X1_124/CTRL2 0.10fF
C58928 POR2X1_556/A PAND2X1_135/O 0.08fF
C58929 POR2X1_13/A PAND2X1_175/B 0.03fF
C58930 POR2X1_730/Y PAND2X1_90/Y 0.12fF
C58931 POR2X1_519/Y PAND2X1_642/B 0.00fF
C58932 POR2X1_567/A POR2X1_590/A 0.09fF
C58933 PAND2X1_373/CTRL VDD -0.00fF
C58934 PAND2X1_217/B POR2X1_129/Y 0.05fF
C58935 POR2X1_492/O POR2X1_394/A 0.05fF
C58936 POR2X1_256/O POR2X1_7/A 0.01fF
C58937 POR2X1_416/Y PAND2X1_642/B 0.01fF
C58938 PAND2X1_353/O VDD 0.00fF
C58939 PAND2X1_794/B PAND2X1_365/B 0.00fF
C58940 POR2X1_7/A PAND2X1_515/CTRL 0.00fF
C58941 POR2X1_697/Y POR2X1_511/CTRL2 0.01fF
C58942 POR2X1_96/A POR2X1_229/Y 0.64fF
C58943 POR2X1_186/Y POR2X1_186/B 0.36fF
C58944 POR2X1_219/B POR2X1_741/Y 0.10fF
C58945 POR2X1_198/B PAND2X1_88/Y 0.00fF
C58946 POR2X1_465/A POR2X1_569/A 0.05fF
C58947 PAND2X1_678/CTRL2 PAND2X1_860/A 0.01fF
C58948 POR2X1_809/A POR2X1_864/a_76_344# 0.00fF
C58949 POR2X1_174/CTRL2 VDD 0.00fF
C58950 POR2X1_614/A POR2X1_407/A 2.50fF
C58951 PAND2X1_844/Y PAND2X1_338/B 0.00fF
C58952 POR2X1_78/A POR2X1_374/CTRL 0.01fF
C58953 PAND2X1_794/B POR2X1_759/A 0.02fF
C58954 PAND2X1_95/B INPUT_6 0.04fF
C58955 PAND2X1_6/A POR2X1_90/Y 0.07fF
C58956 VDD PAND2X1_124/O 0.00fF
C58957 PAND2X1_244/B POR2X1_230/Y 0.06fF
C58958 PAND2X1_467/Y PAND2X1_707/O 0.02fF
C58959 PAND2X1_6/Y POR2X1_196/Y 0.02fF
C58960 POR2X1_578/Y POR2X1_577/m4_208_n4# 0.12fF
C58961 PAND2X1_743/CTRL2 PAND2X1_32/B 0.03fF
C58962 POR2X1_68/A POR2X1_596/A 0.03fF
C58963 POR2X1_513/Y PAND2X1_32/B 0.03fF
C58964 PAND2X1_659/Y PAND2X1_217/B 0.05fF
C58965 POR2X1_36/B POR2X1_581/CTRL2 0.01fF
C58966 PAND2X1_824/B POR2X1_207/CTRL 0.06fF
C58967 PAND2X1_691/Y POR2X1_829/A 0.05fF
C58968 POR2X1_330/Y POR2X1_330/CTRL2 0.05fF
C58969 PAND2X1_96/B POR2X1_702/A 0.07fF
C58970 POR2X1_66/B PAND2X1_665/CTRL 0.12fF
C58971 POR2X1_539/A POR2X1_662/Y 0.20fF
C58972 POR2X1_590/A POR2X1_532/a_76_344# 0.03fF
C58973 PAND2X1_94/A PAND2X1_92/a_16_344# 0.01fF
C58974 POR2X1_324/O VDD 0.00fF
C58975 PAND2X1_620/O POR2X1_13/A 0.02fF
C58976 POR2X1_13/A PAND2X1_777/CTRL 0.01fF
C58977 POR2X1_129/Y VDD 0.90fF
C58978 POR2X1_7/A PAND2X1_506/a_16_344# 0.02fF
C58979 PAND2X1_579/A POR2X1_46/Y 0.16fF
C58980 POR2X1_687/A POR2X1_730/CTRL2 0.01fF
C58981 PAND2X1_48/B PAND2X1_94/A 2.96fF
C58982 INPUT_1 PAND2X1_243/B 0.03fF
C58983 POR2X1_500/Y POR2X1_573/A 0.02fF
C58984 PAND2X1_41/B PAND2X1_41/Y 0.04fF
C58985 POR2X1_272/Y POR2X1_75/Y 0.04fF
C58986 POR2X1_112/Y POR2X1_318/A 0.07fF
C58987 PAND2X1_605/O POR2X1_7/B 0.01fF
C58988 PAND2X1_723/CTRL2 POR2X1_7/A 0.01fF
C58989 POR2X1_760/A POR2X1_329/A 2.80fF
C58990 PAND2X1_552/B PAND2X1_569/Y 2.73fF
C58991 PAND2X1_551/Y POR2X1_765/Y 0.02fF
C58992 PAND2X1_397/O POR2X1_35/Y 0.02fF
C58993 PAND2X1_65/Y POR2X1_4/Y 0.01fF
C58994 POR2X1_403/Y POR2X1_294/A 0.01fF
C58995 PAND2X1_81/O PAND2X1_60/B 0.02fF
C58996 PAND2X1_777/CTRL2 POR2X1_293/Y 0.01fF
C58997 PAND2X1_357/Y POR2X1_103/Y 0.05fF
C58998 POR2X1_164/Y POR2X1_238/Y 0.52fF
C58999 POR2X1_292/O POR2X1_411/B 0.02fF
C59000 POR2X1_41/B POR2X1_394/A 0.41fF
C59001 POR2X1_786/Y POR2X1_222/A 0.01fF
C59002 POR2X1_339/O POR2X1_785/A 0.02fF
C59003 POR2X1_327/Y POR2X1_115/O 0.01fF
C59004 POR2X1_762/CTRL2 INPUT_4 0.01fF
C59005 PAND2X1_476/A POR2X1_5/Y 0.02fF
C59006 POR2X1_614/A PAND2X1_315/CTRL 0.01fF
C59007 POR2X1_366/A PAND2X1_32/B 0.03fF
C59008 PAND2X1_702/CTRL POR2X1_7/A 0.00fF
C59009 POR2X1_730/Y POR2X1_732/CTRL2 0.01fF
C59010 POR2X1_78/B POR2X1_188/Y 0.03fF
C59011 PAND2X1_54/CTRL POR2X1_4/Y 0.07fF
C59012 PAND2X1_659/Y VDD 0.60fF
C59013 PAND2X1_243/B POR2X1_153/Y 0.07fF
C59014 PAND2X1_553/B PAND2X1_853/B 0.07fF
C59015 PAND2X1_858/O POR2X1_13/A 0.01fF
C59016 PAND2X1_631/A POR2X1_236/Y 0.03fF
C59017 PAND2X1_90/Y POR2X1_542/CTRL 0.15fF
C59018 POR2X1_502/A POR2X1_294/A 0.15fF
C59019 POR2X1_448/Y POR2X1_532/O 0.01fF
C59020 PAND2X1_644/CTRL POR2X1_597/Y 0.00fF
C59021 POR2X1_57/A POR2X1_7/A 0.00fF
C59022 POR2X1_783/A POR2X1_294/A 0.02fF
C59023 POR2X1_68/A POR2X1_782/CTRL2 0.03fF
C59024 PAND2X1_474/Y PAND2X1_500/CTRL 0.00fF
C59025 PAND2X1_774/O PAND2X1_568/B 0.02fF
C59026 PAND2X1_519/O POR2X1_260/A 0.04fF
C59027 POR2X1_540/A POR2X1_181/B 0.37fF
C59028 PAND2X1_455/CTRL POR2X1_77/Y 0.01fF
C59029 POR2X1_149/Y POR2X1_209/O 0.00fF
C59030 POR2X1_566/A POR2X1_566/a_16_28# 0.03fF
C59031 PAND2X1_143/O PAND2X1_8/Y 0.17fF
C59032 POR2X1_96/Y VDD 0.25fF
C59033 POR2X1_57/A PAND2X1_130/O 0.08fF
C59034 POR2X1_375/O PAND2X1_32/B 0.18fF
C59035 PAND2X1_687/B VDD 0.16fF
C59036 POR2X1_79/A POR2X1_767/a_16_28# 0.03fF
C59037 INPUT_0 PAND2X1_729/O 0.01fF
C59038 POR2X1_68/A POR2X1_449/A 0.07fF
C59039 PAND2X1_691/Y POR2X1_761/Y 0.03fF
C59040 POR2X1_697/Y PAND2X1_708/O 0.00fF
C59041 PAND2X1_555/A PAND2X1_345/Y 0.09fF
C59042 INPUT_0 POR2X1_371/m4_208_n4# 0.08fF
C59043 POR2X1_835/B POR2X1_776/A 0.01fF
C59044 PAND2X1_427/a_56_28# PAND2X1_72/A 0.00fF
C59045 PAND2X1_140/A POR2X1_103/Y 0.00fF
C59046 PAND2X1_837/a_16_344# POR2X1_826/Y 0.04fF
C59047 PAND2X1_501/a_76_28# POR2X1_72/B 0.01fF
C59048 PAND2X1_28/CTRL2 PAND2X1_63/B 0.01fF
C59049 POR2X1_216/O POR2X1_276/Y 0.01fF
C59050 PAND2X1_698/a_16_344# POR2X1_532/A 0.02fF
C59051 POR2X1_130/A POR2X1_561/B 0.04fF
C59052 POR2X1_294/B POR2X1_788/CTRL2 0.05fF
C59053 POR2X1_383/A POR2X1_101/Y 0.40fF
C59054 POR2X1_62/Y POR2X1_620/CTRL 0.01fF
C59055 PAND2X1_482/O POR2X1_786/Y 0.31fF
C59056 PAND2X1_122/a_16_344# POR2X1_121/Y 0.02fF
C59057 PAND2X1_856/B PAND2X1_854/A 0.01fF
C59058 PAND2X1_274/CTRL POR2X1_39/B 0.01fF
C59059 PAND2X1_849/B PAND2X1_63/B 0.12fF
C59060 POR2X1_508/A D_GATE_741 0.03fF
C59061 POR2X1_351/Y POR2X1_502/Y 0.03fF
C59062 VDD PAND2X1_333/Y 0.13fF
C59063 POR2X1_111/Y POR2X1_7/A 0.02fF
C59064 PAND2X1_6/Y POR2X1_447/B 0.03fF
C59065 PAND2X1_655/Y POR2X1_690/O 0.01fF
C59066 PAND2X1_6/Y POR2X1_552/a_16_28# 0.03fF
C59067 POR2X1_326/A POR2X1_209/A 0.03fF
C59068 POR2X1_86/Y POR2X1_88/Y 0.01fF
C59069 POR2X1_52/A POR2X1_305/CTRL 0.01fF
C59070 POR2X1_272/Y PAND2X1_332/Y 0.40fF
C59071 POR2X1_732/B PAND2X1_179/O 0.07fF
C59072 POR2X1_119/Y POR2X1_90/Y 0.07fF
C59073 INPUT_1 POR2X1_376/CTRL2 0.00fF
C59074 POR2X1_675/Y POR2X1_737/O 0.01fF
C59075 PAND2X1_857/A POR2X1_153/Y 0.07fF
C59076 POR2X1_191/B POR2X1_319/Y 0.03fF
C59077 POR2X1_681/CTRL2 POR2X1_32/A 0.01fF
C59078 POR2X1_52/A PAND2X1_440/O 0.01fF
C59079 POR2X1_385/Y PAND2X1_389/a_76_28# 0.05fF
C59080 POR2X1_110/a_76_344# POR2X1_73/Y 0.00fF
C59081 INPUT_1 POR2X1_260/A 0.06fF
C59082 POR2X1_305/O POR2X1_55/Y 0.01fF
C59083 POR2X1_525/Y POR2X1_416/B 0.05fF
C59084 D_GATE_741 POR2X1_568/B 0.02fF
C59085 POR2X1_863/A POR2X1_552/Y 0.01fF
C59086 POR2X1_517/CTRL2 POR2X1_73/Y 0.03fF
C59087 POR2X1_510/Y POR2X1_553/a_16_28# 0.03fF
C59088 POR2X1_719/O POR2X1_294/A 0.01fF
C59089 PAND2X1_631/A PAND2X1_344/CTRL 0.06fF
C59090 POR2X1_523/Y POR2X1_39/B 0.03fF
C59091 PAND2X1_640/B POR2X1_411/B 0.03fF
C59092 PAND2X1_403/B POR2X1_399/Y 0.04fF
C59093 PAND2X1_96/B PAND2X1_759/O 0.02fF
C59094 POR2X1_390/B POR2X1_327/Y 0.03fF
C59095 POR2X1_782/O POR2X1_260/A 0.01fF
C59096 POR2X1_101/Y PAND2X1_71/Y 0.05fF
C59097 POR2X1_257/A POR2X1_23/Y 0.52fF
C59098 POR2X1_14/CTRL INPUT_3 0.01fF
C59099 POR2X1_507/O POR2X1_507/B 0.04fF
C59100 POR2X1_394/A PAND2X1_308/Y 0.03fF
C59101 POR2X1_150/Y POR2X1_32/A 0.31fF
C59102 PAND2X1_341/A POR2X1_39/B 0.01fF
C59103 POR2X1_666/CTRL POR2X1_411/B 0.01fF
C59104 POR2X1_760/A PAND2X1_361/O 0.06fF
C59105 POR2X1_54/Y PAND2X1_68/CTRL 0.02fF
C59106 POR2X1_137/B POR2X1_78/A 0.07fF
C59107 POR2X1_48/A POR2X1_815/A 0.01fF
C59108 PAND2X1_50/CTRL D_INPUT_7 0.01fF
C59109 POR2X1_93/A POR2X1_39/B 3.52fF
C59110 POR2X1_39/B POR2X1_91/Y 0.06fF
C59111 POR2X1_119/Y PAND2X1_123/a_76_28# 0.03fF
C59112 POR2X1_537/Y POR2X1_733/Y 0.08fF
C59113 PAND2X1_74/CTRL2 POR2X1_341/A 0.06fF
C59114 POR2X1_411/B POR2X1_272/CTRL2 0.02fF
C59115 POR2X1_14/Y PAND2X1_407/CTRL 0.01fF
C59116 POR2X1_284/a_16_28# POR2X1_325/A 0.01fF
C59117 POR2X1_416/B PAND2X1_551/O 0.04fF
C59118 POR2X1_416/B POR2X1_283/A 18.85fF
C59119 PAND2X1_631/A POR2X1_271/A 0.07fF
C59120 D_INPUT_0 POR2X1_218/Y 0.07fF
C59121 PAND2X1_637/O POR2X1_586/Y 0.00fF
C59122 POR2X1_97/A POR2X1_66/A 0.03fF
C59123 PAND2X1_93/B POR2X1_78/A 0.06fF
C59124 PAND2X1_452/A POR2X1_416/B 0.04fF
C59125 POR2X1_257/A POR2X1_312/Y 0.03fF
C59126 POR2X1_49/Y PAND2X1_796/B 0.01fF
C59127 PAND2X1_239/O POR2X1_590/A 0.02fF
C59128 POR2X1_703/Y POR2X1_169/A 0.01fF
C59129 POR2X1_333/A POR2X1_212/a_16_28# 0.04fF
C59130 POR2X1_257/A POR2X1_764/Y 0.03fF
C59131 POR2X1_49/Y PAND2X1_454/B 0.00fF
C59132 POR2X1_110/Y POR2X1_119/Y 0.10fF
C59133 POR2X1_855/B PAND2X1_72/A 0.03fF
C59134 PAND2X1_221/Y PAND2X1_365/B 0.04fF
C59135 POR2X1_815/O INPUT_0 0.24fF
C59136 PAND2X1_57/B PAND2X1_45/CTRL 0.01fF
C59137 POR2X1_169/B POR2X1_192/B 0.18fF
C59138 POR2X1_180/A POR2X1_181/Y 0.42fF
C59139 POR2X1_399/O POR2X1_20/B 0.02fF
C59140 POR2X1_352/CTRL PAND2X1_52/B 0.03fF
C59141 PAND2X1_623/O POR2X1_669/B 0.18fF
C59142 POR2X1_846/A POR2X1_793/A 0.03fF
C59143 POR2X1_814/A POR2X1_575/B 0.19fF
C59144 POR2X1_438/Y POR2X1_40/Y 0.03fF
C59145 POR2X1_383/A POR2X1_579/O 0.01fF
C59146 POR2X1_352/CTRL POR2X1_212/B 0.01fF
C59147 POR2X1_260/B POR2X1_752/Y 0.02fF
C59148 PAND2X1_48/B POR2X1_462/CTRL2 0.01fF
C59149 POR2X1_394/A POR2X1_77/Y 0.35fF
C59150 POR2X1_812/A POR2X1_801/B 0.05fF
C59151 POR2X1_593/a_16_28# POR2X1_592/Y 0.05fF
C59152 POR2X1_287/B POR2X1_458/CTRL2 0.01fF
C59153 POR2X1_856/B POR2X1_436/O 0.06fF
C59154 PAND2X1_443/O PAND2X1_803/A 0.00fF
C59155 POR2X1_49/Y POR2X1_23/Y 3.25fF
C59156 POR2X1_56/a_16_28# POR2X1_669/B 0.03fF
C59157 POR2X1_130/A PAND2X1_39/B 0.19fF
C59158 POR2X1_734/B POR2X1_288/A 0.02fF
C59159 POR2X1_812/CTRL2 POR2X1_452/Y 0.01fF
C59160 POR2X1_137/B PAND2X1_132/CTRL 0.01fF
C59161 PAND2X1_841/CTRL2 POR2X1_271/B 0.01fF
C59162 POR2X1_43/B PAND2X1_97/Y 0.03fF
C59163 POR2X1_634/A POR2X1_805/Y 0.05fF
C59164 POR2X1_590/A POR2X1_643/A 0.12fF
C59165 POR2X1_411/B POR2X1_7/B 0.10fF
C59166 POR2X1_45/CTRL2 POR2X1_23/Y 0.03fF
C59167 POR2X1_39/B POR2X1_397/O 0.18fF
C59168 POR2X1_83/B PAND2X1_249/CTRL 0.01fF
C59169 PAND2X1_282/O PAND2X1_41/B 0.04fF
C59170 PAND2X1_231/a_16_344# POR2X1_263/Y 0.00fF
C59171 POR2X1_833/CTRL2 POR2X1_541/B 0.05fF
C59172 POR2X1_465/B POR2X1_341/A 0.03fF
C59173 POR2X1_679/A PAND2X1_804/B 0.01fF
C59174 PAND2X1_20/A POR2X1_634/A 0.05fF
C59175 POR2X1_274/a_16_28# POR2X1_330/Y 0.01fF
C59176 POR2X1_189/Y POR2X1_150/Y 0.06fF
C59177 POR2X1_748/A POR2X1_102/Y 0.01fF
C59178 PAND2X1_476/CTRL POR2X1_102/Y 0.00fF
C59179 POR2X1_597/Y POR2X1_761/CTRL 0.01fF
C59180 PAND2X1_94/A PAND2X1_233/CTRL2 0.02fF
C59181 POR2X1_603/Y POR2X1_40/Y 0.03fF
C59182 POR2X1_329/A POR2X1_38/Y 0.10fF
C59183 POR2X1_96/A POR2X1_271/CTRL2 0.03fF
C59184 PAND2X1_128/O POR2X1_411/B 0.01fF
C59185 POR2X1_376/B PAND2X1_796/CTRL 0.00fF
C59186 POR2X1_150/Y POR2X1_184/Y 0.03fF
C59187 POR2X1_20/B POR2X1_619/O 0.01fF
C59188 PAND2X1_20/A POR2X1_489/CTRL2 0.02fF
C59189 POR2X1_801/CTRL POR2X1_121/B 0.04fF
C59190 POR2X1_296/CTRL2 PAND2X1_69/A 0.03fF
C59191 POR2X1_60/A PAND2X1_140/CTRL 0.00fF
C59192 POR2X1_807/A POR2X1_590/A 0.09fF
C59193 POR2X1_48/A POR2X1_481/CTRL2 0.01fF
C59194 PAND2X1_407/CTRL POR2X1_55/Y 0.01fF
C59195 POR2X1_447/B PAND2X1_52/B 0.12fF
C59196 POR2X1_193/Y POR2X1_555/B 0.03fF
C59197 POR2X1_338/CTRL2 POR2X1_814/A 0.06fF
C59198 PAND2X1_58/A POR2X1_585/CTRL 0.27fF
C59199 POR2X1_37/Y VDD 5.10fF
C59200 POR2X1_57/A POR2X1_760/A 0.07fF
C59201 PAND2X1_410/O POR2X1_290/Y 0.37fF
C59202 POR2X1_817/CTRL POR2X1_817/A 0.01fF
C59203 PAND2X1_23/Y POR2X1_446/B 0.03fF
C59204 PAND2X1_73/Y POR2X1_573/O 0.02fF
C59205 PAND2X1_463/CTRL POR2X1_94/A 0.01fF
C59206 POR2X1_196/a_56_344# PAND2X1_48/Y 0.00fF
C59207 PAND2X1_35/A POR2X1_42/Y 0.03fF
C59208 PAND2X1_75/O PAND2X1_60/B 0.17fF
C59209 POR2X1_83/B PAND2X1_803/A 0.08fF
C59210 POR2X1_814/B POR2X1_634/A 0.05fF
C59211 PAND2X1_99/B PAND2X1_99/CTRL 0.01fF
C59212 PAND2X1_58/A POR2X1_830/A 0.12fF
C59213 POR2X1_13/A POR2X1_409/B 0.03fF
C59214 POR2X1_32/A POR2X1_701/Y 0.01fF
C59215 POR2X1_188/A POR2X1_389/Y 0.03fF
C59216 PAND2X1_612/B PAND2X1_283/CTRL2 0.00fF
C59217 POR2X1_52/A PAND2X1_640/B 0.03fF
C59218 POR2X1_777/B PAND2X1_41/B 0.03fF
C59219 POR2X1_20/B POR2X1_68/B 0.03fF
C59220 POR2X1_231/CTRL2 POR2X1_66/A 0.01fF
C59221 PAND2X1_492/O POR2X1_78/A 0.04fF
C59222 D_INPUT_0 POR2X1_46/Y 2.91fF
C59223 POR2X1_836/CTRL2 POR2X1_578/Y 0.03fF
C59224 PAND2X1_695/CTRL POR2X1_634/A 0.13fF
C59225 POR2X1_567/B POR2X1_466/CTRL 0.00fF
C59226 POR2X1_194/A PAND2X1_41/B 0.19fF
C59227 POR2X1_582/CTRL2 POR2X1_257/A 0.03fF
C59228 POR2X1_130/A POR2X1_805/Y 0.02fF
C59229 POR2X1_92/CTRL2 INPUT_3 0.11fF
C59230 POR2X1_210/CTRL POR2X1_220/Y 0.00fF
C59231 POR2X1_865/B POR2X1_475/CTRL 0.08fF
C59232 POR2X1_65/A POR2X1_503/A 0.04fF
C59233 POR2X1_638/O POR2X1_66/A 0.01fF
C59234 POR2X1_722/B POR2X1_66/A 0.02fF
C59235 POR2X1_323/CTRL2 POR2X1_65/A 0.03fF
C59236 POR2X1_813/O POR2X1_38/Y 0.03fF
C59237 POR2X1_296/B POR2X1_722/Y 0.01fF
C59238 POR2X1_41/B POR2X1_669/B 0.28fF
C59239 PAND2X1_9/Y POR2X1_205/A 0.03fF
C59240 PAND2X1_20/A POR2X1_130/A 0.29fF
C59241 PAND2X1_39/B POR2X1_573/A 0.03fF
C59242 POR2X1_366/Y POR2X1_66/A 0.07fF
C59243 POR2X1_83/B PAND2X1_673/Y 4.91fF
C59244 POR2X1_66/A POR2X1_294/B 2.27fF
C59245 PAND2X1_48/B POR2X1_477/Y 0.07fF
C59246 POR2X1_76/A POR2X1_804/A 2.14fF
C59247 PAND2X1_778/Y PAND2X1_796/B 0.10fF
C59248 POR2X1_32/A PAND2X1_364/B 0.07fF
C59249 POR2X1_266/CTRL PAND2X1_69/A 0.01fF
C59250 PAND2X1_65/B PAND2X1_41/B 1.78fF
C59251 POR2X1_429/CTRL VDD 0.00fF
C59252 POR2X1_805/a_16_28# POR2X1_805/A 0.00fF
C59253 POR2X1_566/A PAND2X1_20/A 0.05fF
C59254 POR2X1_654/B POR2X1_476/Y 0.03fF
C59255 POR2X1_490/CTRL POR2X1_7/A 0.01fF
C59256 POR2X1_640/CTRL INPUT_0 0.01fF
C59257 PAND2X1_73/O PAND2X1_8/Y 0.07fF
C59258 POR2X1_523/Y POR2X1_48/A 0.00fF
C59259 POR2X1_485/Y PAND2X1_550/B 0.04fF
C59260 PAND2X1_246/m4_208_n4# POR2X1_101/Y 0.05fF
C59261 POR2X1_590/A POR2X1_546/B 0.01fF
C59262 POR2X1_565/B POR2X1_590/A 0.02fF
C59263 POR2X1_502/A POR2X1_638/A 0.01fF
C59264 POR2X1_102/Y PAND2X1_598/a_76_28# 0.02fF
C59265 POR2X1_329/A POR2X1_153/Y 0.10fF
C59266 POR2X1_68/A D_INPUT_0 0.11fF
C59267 PAND2X1_453/CTRL2 POR2X1_14/Y 0.00fF
C59268 POR2X1_378/Y PAND2X1_459/CTRL2 0.01fF
C59269 POR2X1_244/O POR2X1_243/Y 0.05fF
C59270 PAND2X1_205/A POR2X1_498/A 0.02fF
C59271 POR2X1_13/A PAND2X1_244/a_56_28# 0.00fF
C59272 PAND2X1_48/B PAND2X1_11/Y 0.00fF
C59273 PAND2X1_248/CTRL POR2X1_532/A 0.01fF
C59274 POR2X1_509/B VDD 0.11fF
C59275 POR2X1_482/Y POR2X1_252/CTRL2 0.01fF
C59276 POR2X1_744/Y POR2X1_158/B 0.39fF
C59277 POR2X1_43/B POR2X1_754/Y 0.12fF
C59278 POR2X1_330/Y PAND2X1_516/O 0.04fF
C59279 PAND2X1_862/B POR2X1_72/B 0.03fF
C59280 PAND2X1_23/Y POR2X1_121/B 0.06fF
C59281 POR2X1_186/Y PAND2X1_321/a_76_28# 0.02fF
C59282 POR2X1_297/A PAND2X1_768/Y 0.02fF
C59283 PAND2X1_859/A POR2X1_224/O 0.01fF
C59284 POR2X1_181/m4_208_n4# POR2X1_181/A 0.01fF
C59285 POR2X1_432/O PAND2X1_658/B 0.01fF
C59286 POR2X1_416/B POR2X1_32/CTRL 0.01fF
C59287 POR2X1_647/CTRL2 PAND2X1_60/B 0.10fF
C59288 POR2X1_814/B POR2X1_130/A 0.38fF
C59289 PAND2X1_96/B POR2X1_499/O 0.16fF
C59290 PAND2X1_661/B POR2X1_409/B 0.96fF
C59291 POR2X1_859/A POR2X1_720/A 0.03fF
C59292 PAND2X1_139/O PAND2X1_137/Y 0.00fF
C59293 POR2X1_407/A POR2X1_590/A 0.13fF
C59294 POR2X1_566/A POR2X1_814/B 0.10fF
C59295 POR2X1_48/A POR2X1_93/A 0.08fF
C59296 POR2X1_29/A POR2X1_409/CTRL2 0.01fF
C59297 PAND2X1_725/Y POR2X1_763/Y 0.02fF
C59298 POR2X1_734/A POR2X1_784/A 0.07fF
C59299 POR2X1_2/CTRL VDD -0.00fF
C59300 POR2X1_48/A POR2X1_91/Y 0.03fF
C59301 POR2X1_54/Y PAND2X1_819/O 0.07fF
C59302 POR2X1_528/O POR2X1_14/Y 0.17fF
C59303 POR2X1_66/CTRL2 PAND2X1_58/A 0.01fF
C59304 PAND2X1_787/CTRL2 POR2X1_7/B 0.00fF
C59305 PAND2X1_47/B PAND2X1_587/CTRL 0.01fF
C59306 POR2X1_330/Y PAND2X1_369/a_16_344# 0.06fF
C59307 POR2X1_54/Y POR2X1_773/B 0.12fF
C59308 POR2X1_681/a_16_28# POR2X1_153/Y 0.07fF
C59309 POR2X1_528/O PAND2X1_453/A 0.01fF
C59310 POR2X1_379/O POR2X1_260/B 0.01fF
C59311 POR2X1_83/B PAND2X1_365/B 0.01fF
C59312 POR2X1_141/Y POR2X1_276/O 0.18fF
C59313 POR2X1_356/A POR2X1_439/Y 0.05fF
C59314 POR2X1_33/CTRL POR2X1_68/B 0.01fF
C59315 POR2X1_406/Y VDD 0.16fF
C59316 POR2X1_231/A POR2X1_231/B 0.02fF
C59317 PAND2X1_20/A POR2X1_844/B 0.04fF
C59318 PAND2X1_454/a_16_344# POR2X1_72/B 0.02fF
C59319 POR2X1_66/A PAND2X1_111/B 0.00fF
C59320 PAND2X1_55/Y POR2X1_593/B 0.01fF
C59321 PAND2X1_797/O PAND2X1_782/Y -0.00fF
C59322 POR2X1_93/A POR2X1_225/CTRL2 0.03fF
C59323 POR2X1_218/Y POR2X1_361/O 0.02fF
C59324 POR2X1_13/A POR2X1_272/Y 0.07fF
C59325 POR2X1_376/B POR2X1_7/B 2.15fF
C59326 PAND2X1_859/B PAND2X1_61/Y 0.06fF
C59327 PAND2X1_471/B POR2X1_236/Y 0.20fF
C59328 POR2X1_776/A POR2X1_566/CTRL2 0.01fF
C59329 POR2X1_835/B POR2X1_191/Y 0.05fF
C59330 PAND2X1_414/O POR2X1_4/Y 0.06fF
C59331 POR2X1_468/a_16_28# PAND2X1_41/B 0.01fF
C59332 POR2X1_96/A PAND2X1_84/Y 0.02fF
C59333 POR2X1_730/B POR2X1_330/Y 0.03fF
C59334 PAND2X1_741/B PAND2X1_364/B 0.07fF
C59335 POR2X1_48/A POR2X1_416/O 0.01fF
C59336 POR2X1_596/A PAND2X1_58/A 0.03fF
C59337 POR2X1_60/A PAND2X1_509/CTRL 0.04fF
C59338 PAND2X1_129/CTRL PAND2X1_90/A 0.01fF
C59339 PAND2X1_6/Y POR2X1_141/Y 0.03fF
C59340 POR2X1_78/A PAND2X1_173/CTRL 0.01fF
C59341 PAND2X1_771/Y PAND2X1_552/O 0.34fF
C59342 POR2X1_57/A POR2X1_311/Y 0.03fF
C59343 POR2X1_813/Y POR2X1_37/Y 0.02fF
C59344 POR2X1_136/O POR2X1_40/Y 0.04fF
C59345 PAND2X1_6/Y PAND2X1_423/CTRL2 0.00fF
C59346 POR2X1_814/B POR2X1_204/CTRL 0.00fF
C59347 PAND2X1_738/Y PAND2X1_182/A 0.03fF
C59348 PAND2X1_655/Y INPUT_0 0.03fF
C59349 POR2X1_130/A POR2X1_513/B 0.04fF
C59350 POR2X1_13/A PAND2X1_351/Y 0.01fF
C59351 POR2X1_293/Y VDD 2.41fF
C59352 POR2X1_566/A PAND2X1_176/CTRL2 0.01fF
C59353 POR2X1_842/CTRL POR2X1_675/Y 0.01fF
C59354 PAND2X1_60/CTRL2 PAND2X1_58/A 0.01fF
C59355 PAND2X1_115/a_56_28# PAND2X1_787/Y 0.00fF
C59356 PAND2X1_555/A VDD 0.11fF
C59357 PAND2X1_48/B POR2X1_215/CTRL2 0.01fF
C59358 PAND2X1_90/A PAND2X1_8/Y 1.91fF
C59359 POR2X1_66/B POR2X1_318/A 0.06fF
C59360 POR2X1_655/A POR2X1_774/A 0.03fF
C59361 POR2X1_416/B POR2X1_399/Y 0.01fF
C59362 POR2X1_865/m4_208_n4# PAND2X1_48/A 0.09fF
C59363 POR2X1_832/B VDD 0.29fF
C59364 POR2X1_68/A PAND2X1_90/Y 0.16fF
C59365 POR2X1_12/A POR2X1_762/O 0.01fF
C59366 PAND2X1_450/a_16_344# POR2X1_427/Y 0.02fF
C59367 PAND2X1_81/B POR2X1_786/CTRL 0.04fF
C59368 PAND2X1_62/O PAND2X1_6/A 0.09fF
C59369 POR2X1_72/O PAND2X1_651/Y 0.02fF
C59370 POR2X1_812/B POR2X1_750/B 0.01fF
C59371 PAND2X1_849/B POR2X1_32/A 0.02fF
C59372 POR2X1_96/Y PAND2X1_9/Y 0.03fF
C59373 POR2X1_66/B POR2X1_713/B 0.05fF
C59374 PAND2X1_659/O PAND2X1_575/A 0.02fF
C59375 PAND2X1_96/B POR2X1_653/B 0.13fF
C59376 PAND2X1_96/B PAND2X1_323/m4_208_n4# 0.07fF
C59377 POR2X1_52/A POR2X1_7/B 6.69fF
C59378 PAND2X1_675/A PAND2X1_740/Y 1.15fF
C59379 POR2X1_461/B POR2X1_793/A 0.02fF
C59380 PAND2X1_197/CTRL2 PAND2X1_364/B 0.03fF
C59381 POR2X1_463/O PAND2X1_52/B 0.02fF
C59382 POR2X1_186/Y POR2X1_736/O 0.01fF
C59383 POR2X1_403/B POR2X1_35/Y 0.03fF
C59384 PAND2X1_73/Y POR2X1_456/B 0.00fF
C59385 PAND2X1_96/B POR2X1_640/A 0.00fF
C59386 POR2X1_502/A PAND2X1_95/a_16_344# 0.01fF
C59387 POR2X1_188/A POR2X1_713/B 0.05fF
C59388 PAND2X1_817/CTRL2 POR2X1_750/Y 0.04fF
C59389 POR2X1_537/CTRL POR2X1_590/A 0.01fF
C59390 POR2X1_655/Y POR2X1_725/Y 0.12fF
C59391 POR2X1_78/B POR2X1_243/CTRL2 0.03fF
C59392 PAND2X1_6/A INPUT_0 0.46fF
C59393 POR2X1_669/B PAND2X1_308/Y 0.03fF
C59394 POR2X1_57/A POR2X1_485/CTRL2 0.01fF
C59395 POR2X1_83/Y PAND2X1_404/Y 0.02fF
C59396 PAND2X1_417/O POR2X1_736/A 0.12fF
C59397 POR2X1_697/Y POR2X1_531/O 0.01fF
C59398 POR2X1_296/B POR2X1_244/Y 0.06fF
C59399 POR2X1_558/B PAND2X1_48/A 0.07fF
C59400 PAND2X1_65/B POR2X1_686/O 0.01fF
C59401 POR2X1_66/B POR2X1_61/CTRL 0.01fF
C59402 POR2X1_480/A POR2X1_209/A 0.07fF
C59403 PAND2X1_55/O PAND2X1_60/B 0.03fF
C59404 PAND2X1_467/Y POR2X1_40/Y 0.03fF
C59405 POR2X1_277/a_16_28# POR2X1_46/Y 0.02fF
C59406 POR2X1_325/A POR2X1_573/A 0.03fF
C59407 POR2X1_805/B PAND2X1_60/B 0.04fF
C59408 PAND2X1_6/Y POR2X1_220/Y 0.13fF
C59409 PAND2X1_631/CTRL POR2X1_625/Y 0.03fF
C59410 POR2X1_305/a_16_28# POR2X1_305/Y 0.03fF
C59411 POR2X1_671/O POR2X1_38/B 0.02fF
C59412 PAND2X1_65/B PAND2X1_518/a_76_28# 0.02fF
C59413 POR2X1_353/Y POR2X1_319/Y 0.03fF
C59414 POR2X1_71/Y POR2X1_43/B 0.04fF
C59415 PAND2X1_65/B POR2X1_228/Y 0.03fF
C59416 PAND2X1_192/Y POR2X1_283/A 0.03fF
C59417 POR2X1_234/Y POR2X1_232/Y 0.03fF
C59418 POR2X1_222/Y POR2X1_294/B 0.06fF
C59419 PAND2X1_739/B PAND2X1_739/O 0.02fF
C59420 POR2X1_57/A PAND2X1_719/CTRL 0.01fF
C59421 POR2X1_296/B PAND2X1_527/CTRL2 0.00fF
C59422 POR2X1_860/A POR2X1_218/O 0.01fF
C59423 PAND2X1_56/Y PAND2X1_23/Y 0.15fF
C59424 POR2X1_119/Y POR2X1_265/a_16_28# 0.08fF
C59425 PAND2X1_35/Y POR2X1_229/O 0.01fF
C59426 POR2X1_52/A PAND2X1_477/B 0.03fF
C59427 PAND2X1_6/Y POR2X1_404/Y 0.03fF
C59428 POR2X1_807/A POR2X1_590/a_56_344# 0.00fF
C59429 PAND2X1_651/Y PAND2X1_364/B 0.10fF
C59430 POR2X1_43/B POR2X1_42/Y 1.14fF
C59431 POR2X1_567/A POR2X1_66/A 0.24fF
C59432 POR2X1_192/Y POR2X1_190/O 0.04fF
C59433 POR2X1_78/B POR2X1_510/Y 0.08fF
C59434 POR2X1_38/B POR2X1_817/A 0.09fF
C59435 POR2X1_66/B POR2X1_574/Y 0.03fF
C59436 POR2X1_84/a_16_28# POR2X1_294/B 0.02fF
C59437 PAND2X1_535/O POR2X1_236/Y 0.04fF
C59438 POR2X1_111/CTRL POR2X1_46/Y 0.25fF
C59439 POR2X1_809/A POR2X1_121/B 0.04fF
C59440 POR2X1_408/Y VDD 7.15fF
C59441 PAND2X1_484/a_56_28# PAND2X1_73/Y 0.00fF
C59442 POR2X1_389/A POR2X1_502/A 0.03fF
C59443 POR2X1_180/B PAND2X1_90/Y 0.03fF
C59444 POR2X1_802/CTRL2 POR2X1_435/Y 0.03fF
C59445 POR2X1_72/B PAND2X1_704/CTRL 0.06fF
C59446 POR2X1_569/a_16_28# POR2X1_569/A -0.00fF
C59447 POR2X1_32/A POR2X1_150/O 0.01fF
C59448 PAND2X1_6/Y PAND2X1_273/CTRL 0.07fF
C59449 POR2X1_437/Y PAND2X1_798/B 0.04fF
C59450 POR2X1_573/CTRL2 POR2X1_456/B 0.01fF
C59451 POR2X1_43/B POR2X1_309/Y 0.05fF
C59452 PAND2X1_65/B POR2X1_502/CTRL 0.01fF
C59453 PAND2X1_95/B POR2X1_638/Y 0.28fF
C59454 POR2X1_859/A POR2X1_713/B 0.07fF
C59455 PAND2X1_845/a_16_344# POR2X1_55/Y 0.04fF
C59456 PAND2X1_119/O POR2X1_294/B 0.03fF
C59457 PAND2X1_633/CTRL2 POR2X1_153/Y 0.05fF
C59458 POR2X1_708/m4_208_n4# PAND2X1_743/m4_208_n4# 0.05fF
C59459 PAND2X1_807/a_16_344# POR2X1_7/B 0.02fF
C59460 PAND2X1_614/O POR2X1_129/Y 0.02fF
C59461 POR2X1_38/B POR2X1_42/Y 0.12fF
C59462 POR2X1_532/A POR2X1_294/B 4.80fF
C59463 PAND2X1_341/A PAND2X1_197/Y 0.01fF
C59464 PAND2X1_48/B POR2X1_98/B 0.00fF
C59465 PAND2X1_726/B POR2X1_763/CTRL 0.04fF
C59466 POR2X1_569/a_16_28# POR2X1_570/Y 0.07fF
C59467 POR2X1_192/Y POR2X1_569/A 0.12fF
C59468 PAND2X1_347/Y PAND2X1_343/CTRL2 0.01fF
C59469 INPUT_0 POR2X1_385/CTRL 0.01fF
C59470 POR2X1_264/Y POR2X1_68/B 0.03fF
C59471 POR2X1_96/B POR2X1_96/A 0.00fF
C59472 POR2X1_83/CTRL2 PAND2X1_734/B 0.01fF
C59473 PAND2X1_453/a_16_344# PAND2X1_241/Y 0.03fF
C59474 POR2X1_83/B PAND2X1_352/O 0.06fF
C59475 POR2X1_237/Y POR2X1_90/Y 0.02fF
C59476 PAND2X1_569/CTRL VDD 0.00fF
C59477 POR2X1_72/B PAND2X1_716/B 0.03fF
C59478 PAND2X1_530/a_76_28# PAND2X1_32/B 0.01fF
C59479 PAND2X1_686/CTRL2 POR2X1_13/A 0.00fF
C59480 PAND2X1_216/a_56_28# PAND2X1_656/A 0.00fF
C59481 PAND2X1_651/Y POR2X1_229/O 0.04fF
C59482 POR2X1_192/Y POR2X1_570/Y 0.10fF
C59483 POR2X1_356/A POR2X1_568/Y 0.10fF
C59484 PAND2X1_849/B PAND2X1_35/Y 0.03fF
C59485 PAND2X1_23/Y POR2X1_383/A 0.22fF
C59486 POR2X1_700/Y PAND2X1_711/A 0.90fF
C59487 POR2X1_68/A POR2X1_348/CTRL2 0.32fF
C59488 POR2X1_43/B PAND2X1_99/Y 0.02fF
C59489 PAND2X1_7/O POR2X1_510/Y 0.05fF
C59490 POR2X1_697/Y POR2X1_527/Y 0.31fF
C59491 POR2X1_703/A PAND2X1_176/CTRL 0.01fF
C59492 POR2X1_669/B POR2X1_77/Y 0.27fF
C59493 POR2X1_590/Y POR2X1_722/Y 0.09fF
C59494 POR2X1_199/CTRL PAND2X1_824/B 0.07fF
C59495 POR2X1_121/B POR2X1_711/Y 0.07fF
C59496 POR2X1_57/A POR2X1_38/Y 0.07fF
C59497 POR2X1_51/CTRL INPUT_7 0.01fF
C59498 PAND2X1_474/Y POR2X1_150/CTRL 0.00fF
C59499 POR2X1_416/B POR2X1_14/Y 0.83fF
C59500 POR2X1_390/B POR2X1_335/A 0.00fF
C59501 POR2X1_532/A PAND2X1_111/B 0.03fF
C59502 POR2X1_222/A POR2X1_556/Y 0.04fF
C59503 PAND2X1_533/O POR2X1_802/B 0.05fF
C59504 POR2X1_416/B PAND2X1_453/A 0.03fF
C59505 POR2X1_366/CTRL PAND2X1_6/Y 0.06fF
C59506 PAND2X1_319/B PAND2X1_388/Y 0.07fF
C59507 POR2X1_16/A PAND2X1_798/B 2.22fF
C59508 PAND2X1_115/O PAND2X1_348/A 0.04fF
C59509 POR2X1_776/B POR2X1_566/CTRL 0.01fF
C59510 POR2X1_123/A PAND2X1_518/O 0.03fF
C59511 PAND2X1_608/CTRL2 POR2X1_411/B 0.01fF
C59512 POR2X1_346/B POR2X1_61/B 0.00fF
C59513 POR2X1_38/Y POR2X1_229/Y 0.08fF
C59514 POR2X1_96/A PAND2X1_507/a_76_28# 0.04fF
C59515 POR2X1_119/Y INPUT_0 0.10fF
C59516 POR2X1_464/Y POR2X1_543/a_16_28# 0.07fF
C59517 POR2X1_7/B POR2X1_376/m4_208_n4# 0.09fF
C59518 POR2X1_51/A POR2X1_328/CTRL 0.01fF
C59519 POR2X1_110/Y POR2X1_693/CTRL2 0.02fF
C59520 POR2X1_557/A PAND2X1_6/Y 0.01fF
C59521 POR2X1_411/B PAND2X1_206/B 0.07fF
C59522 POR2X1_96/A PAND2X1_858/a_16_344# 0.01fF
C59523 POR2X1_65/A PAND2X1_169/O 0.01fF
C59524 POR2X1_478/B POR2X1_319/Y 0.06fF
C59525 POR2X1_510/B PAND2X1_824/CTRL 0.00fF
C59526 POR2X1_366/a_16_28# POR2X1_68/A 0.06fF
C59527 PAND2X1_90/Y POR2X1_169/A 0.15fF
C59528 PAND2X1_284/O POR2X1_394/A 0.02fF
C59529 POR2X1_220/A POR2X1_568/Y 0.05fF
C59530 POR2X1_409/Y POR2X1_409/O 0.01fF
C59531 VDD POR2X1_330/O 0.00fF
C59532 POR2X1_369/O POR2X1_43/B -0.01fF
C59533 POR2X1_41/B PAND2X1_353/Y 0.01fF
C59534 POR2X1_790/A POR2X1_720/CTRL2 0.06fF
C59535 POR2X1_41/B POR2X1_41/Y 0.01fF
C59536 POR2X1_637/B PAND2X1_56/A 0.01fF
C59537 POR2X1_556/A POR2X1_658/O 0.02fF
C59538 POR2X1_57/A INPUT_1 0.03fF
C59539 PAND2X1_292/O PAND2X1_41/B 0.01fF
C59540 PAND2X1_96/B POR2X1_449/A 0.03fF
C59541 POR2X1_75/O POR2X1_271/A 0.08fF
C59542 PAND2X1_187/O POR2X1_568/Y 0.04fF
C59543 POR2X1_85/Y POR2X1_230/O 0.00fF
C59544 POR2X1_528/Y POR2X1_527/Y 0.01fF
C59545 POR2X1_383/A POR2X1_520/A 0.15fF
C59546 POR2X1_439/Y PAND2X1_72/A 0.03fF
C59547 POR2X1_158/Y PAND2X1_712/CTRL 0.00fF
C59548 POR2X1_416/B POR2X1_48/O 0.04fF
C59549 POR2X1_532/A PAND2X1_533/O 0.02fF
C59550 POR2X1_150/Y PAND2X1_211/CTRL 0.10fF
C59551 POR2X1_326/CTRL2 POR2X1_854/B 0.00fF
C59552 POR2X1_416/B POR2X1_488/a_16_28# 0.01fF
C59553 POR2X1_505/CTRL POR2X1_245/Y 0.03fF
C59554 POR2X1_57/A POR2X1_153/Y 0.07fF
C59555 POR2X1_220/Y POR2X1_632/Y 25.08fF
C59556 POR2X1_119/Y POR2X1_234/CTRL2 0.01fF
C59557 POR2X1_62/Y PAND2X1_69/A 0.10fF
C59558 POR2X1_294/B POR2X1_510/CTRL2 0.01fF
C59559 POR2X1_728/CTRL2 PAND2X1_52/B 0.13fF
C59560 POR2X1_62/Y PAND2X1_341/A 0.07fF
C59561 POR2X1_88/CTRL POR2X1_88/A 0.01fF
C59562 POR2X1_766/Y POR2X1_73/Y 0.01fF
C59563 PAND2X1_691/Y POR2X1_16/A 0.03fF
C59564 POR2X1_571/CTRL2 POR2X1_569/A 0.02fF
C59565 POR2X1_416/B PAND2X1_472/B 0.10fF
C59566 POR2X1_49/O POR2X1_236/Y 0.29fF
C59567 POR2X1_443/A POR2X1_443/a_16_28# 0.11fF
C59568 POR2X1_229/Y POR2X1_153/Y 0.26fF
C59569 POR2X1_760/A POR2X1_674/a_56_344# 0.00fF
C59570 POR2X1_62/Y POR2X1_91/Y 0.07fF
C59571 POR2X1_41/B PAND2X1_327/O 0.00fF
C59572 POR2X1_192/Y PAND2X1_72/A 0.14fF
C59573 POR2X1_220/Y PAND2X1_52/B 0.01fF
C59574 POR2X1_748/A POR2X1_9/Y 0.07fF
C59575 POR2X1_43/B PAND2X1_860/a_56_28# 0.00fF
C59576 POR2X1_848/A POR2X1_20/B 0.07fF
C59577 PAND2X1_224/m4_208_n4# POR2X1_590/A 0.07fF
C59578 POR2X1_567/A POR2X1_532/A 0.28fF
C59579 PAND2X1_174/CTRL POR2X1_77/Y 0.02fF
C59580 PAND2X1_209/A PAND2X1_797/Y 0.03fF
C59581 POR2X1_416/B POR2X1_55/Y 2.43fF
C59582 PAND2X1_837/CTRL2 POR2X1_39/B 0.00fF
C59583 POR2X1_865/a_16_28# POR2X1_862/Y 0.03fF
C59584 PAND2X1_850/Y PAND2X1_858/Y 0.01fF
C59585 POR2X1_140/B POR2X1_554/a_16_28# 0.04fF
C59586 POR2X1_496/a_56_344# POR2X1_260/B 0.00fF
C59587 PAND2X1_56/Y POR2X1_711/Y 0.09fF
C59588 POR2X1_738/A POR2X1_726/CTRL2 0.00fF
C59589 PAND2X1_242/Y VDD 2.55fF
C59590 POR2X1_27/CTRL POR2X1_27/Y 0.00fF
C59591 PAND2X1_9/Y POR2X1_37/Y 0.03fF
C59592 POR2X1_228/CTRL2 POR2X1_260/A 0.03fF
C59593 POR2X1_459/Y PAND2X1_58/A 0.01fF
C59594 POR2X1_158/Y POR2X1_426/O 0.00fF
C59595 POR2X1_276/Y POR2X1_294/A 0.03fF
C59596 POR2X1_362/A PAND2X1_48/A 0.04fF
C59597 PAND2X1_139/CTRL PAND2X1_349/A 0.01fF
C59598 PAND2X1_853/B POR2X1_7/a_16_28# 0.00fF
C59599 PAND2X1_26/A PAND2X1_59/B 0.19fF
C59600 POR2X1_16/A POR2X1_599/a_76_344# -0.01fF
C59601 POR2X1_475/a_16_28# POR2X1_734/B 0.06fF
C59602 POR2X1_814/A PAND2X1_41/B 0.13fF
C59603 POR2X1_737/A POR2X1_675/Y 2.21fF
C59604 POR2X1_502/Y POR2X1_502/O 0.00fF
C59605 POR2X1_768/CTRL2 POR2X1_294/A 0.01fF
C59606 PAND2X1_674/a_16_344# PAND2X1_72/A 0.02fF
C59607 POR2X1_38/Y PAND2X1_339/CTRL 0.07fF
C59608 PAND2X1_623/Y POR2X1_90/O 0.01fF
C59609 PAND2X1_93/B POR2X1_84/A 0.03fF
C59610 POR2X1_791/B PAND2X1_56/A 0.35fF
C59611 PAND2X1_601/O D_INPUT_0 0.04fF
C59612 POR2X1_67/Y POR2X1_849/O 0.01fF
C59613 PAND2X1_338/B POR2X1_39/B 0.00fF
C59614 PAND2X1_29/a_16_344# PAND2X1_52/B 0.03fF
C59615 POR2X1_376/B PAND2X1_206/B 0.09fF
C59616 PAND2X1_224/O VDD 0.00fF
C59617 POR2X1_129/Y PAND2X1_851/CTRL2 0.01fF
C59618 PAND2X1_23/Y POR2X1_354/O 0.11fF
C59619 D_INPUT_5 PAND2X1_11/Y 0.22fF
C59620 PAND2X1_834/O PAND2X1_349/A 0.02fF
C59621 POR2X1_542/B POR2X1_717/B 0.01fF
C59622 PAND2X1_609/O POR2X1_608/Y 0.00fF
C59623 PAND2X1_217/B POR2X1_275/A 0.03fF
C59624 POR2X1_383/A POR2X1_711/Y 0.17fF
C59625 POR2X1_817/CTRL2 POR2X1_32/A 0.02fF
C59626 PAND2X1_732/A PAND2X1_326/B 0.12fF
C59627 D_INPUT_7 INPUT_5 1.59fF
C59628 POR2X1_54/Y PAND2X1_817/a_16_344# 0.06fF
C59629 POR2X1_113/CTRL2 POR2X1_768/A 0.03fF
C59630 POR2X1_776/A POR2X1_186/Y 0.03fF
C59631 PAND2X1_220/Y POR2X1_411/B 0.03fF
C59632 POR2X1_97/A POR2X1_220/B 0.03fF
C59633 POR2X1_362/Y PAND2X1_93/B 0.03fF
C59634 POR2X1_721/O POR2X1_383/Y 0.00fF
C59635 PAND2X1_253/a_16_344# POR2X1_78/A 0.02fF
C59636 PAND2X1_789/CTRL2 POR2X1_39/B 0.00fF
C59637 POR2X1_409/B POR2X1_29/A 0.80fF
C59638 POR2X1_399/CTRL2 POR2X1_411/B 0.01fF
C59639 POR2X1_281/O POR2X1_416/B 0.01fF
C59640 POR2X1_260/B POR2X1_605/a_16_28# 0.02fF
C59641 PAND2X1_60/B PAND2X1_135/O 0.03fF
C59642 POR2X1_105/Y PAND2X1_39/B 0.25fF
C59643 POR2X1_847/B POR2X1_415/A 0.02fF
C59644 POR2X1_412/O VDD 0.00fF
C59645 PAND2X1_759/CTRL PAND2X1_48/A 0.13fF
C59646 POR2X1_490/Y POR2X1_72/B 0.03fF
C59647 PAND2X1_58/A D_INPUT_0 3.16fF
C59648 POR2X1_609/Y PAND2X1_404/CTRL 0.00fF
C59649 PAND2X1_644/Y POR2X1_40/Y 0.01fF
C59650 D_INPUT_5 POR2X1_25/CTRL 0.03fF
C59651 POR2X1_41/B POR2X1_603/CTRL2 0.02fF
C59652 PAND2X1_798/Y PAND2X1_366/a_16_344# 0.03fF
C59653 PAND2X1_487/O POR2X1_287/B 0.02fF
C59654 POR2X1_78/A POR2X1_285/Y 0.03fF
C59655 PAND2X1_65/B POR2X1_454/A 0.03fF
C59656 POR2X1_366/Y PAND2X1_417/CTRL2 0.04fF
C59657 PAND2X1_224/O PAND2X1_32/B 0.03fF
C59658 PAND2X1_577/B VDD 0.05fF
C59659 POR2X1_864/A POR2X1_828/CTRL2 0.00fF
C59660 POR2X1_856/B POR2X1_186/Y 0.10fF
C59661 POR2X1_76/B POR2X1_569/A 0.06fF
C59662 POR2X1_150/Y PAND2X1_335/CTRL 0.14fF
C59663 PAND2X1_20/A POR2X1_241/B 0.06fF
C59664 PAND2X1_449/Y POR2X1_329/A 0.00fF
C59665 POR2X1_23/Y POR2X1_278/CTRL 0.01fF
C59666 POR2X1_814/B POR2X1_805/a_16_28# 0.03fF
C59667 PAND2X1_93/B PAND2X1_65/Y 0.12fF
C59668 PAND2X1_402/O D_INPUT_0 0.05fF
C59669 PAND2X1_48/B POR2X1_705/B 0.03fF
C59670 PAND2X1_65/B POR2X1_644/a_16_28# 0.01fF
C59671 PAND2X1_613/CTRL PAND2X1_8/Y 0.05fF
C59672 POR2X1_260/B PAND2X1_380/O 0.02fF
C59673 POR2X1_445/a_56_344# POR2X1_341/A 0.01fF
C59674 PAND2X1_20/A POR2X1_719/A 0.00fF
C59675 PAND2X1_9/Y POR2X1_293/Y 0.03fF
C59676 POR2X1_416/B PAND2X1_199/B 0.05fF
C59677 PAND2X1_331/O POR2X1_330/Y 0.01fF
C59678 POR2X1_666/a_16_28# PAND2X1_718/Y 0.03fF
C59679 PAND2X1_839/CTRL2 POR2X1_411/B 0.01fF
C59680 POR2X1_241/B POR2X1_254/CTRL 0.01fF
C59681 PAND2X1_8/CTRL2 INPUT_3 0.02fF
C59682 POR2X1_445/A POR2X1_445/CTRL 0.01fF
C59683 POR2X1_157/CTRL POR2X1_257/A 0.01fF
C59684 PAND2X1_216/B PAND2X1_860/A 0.03fF
C59685 POR2X1_427/Y POR2X1_32/A 0.03fF
C59686 POR2X1_760/A POR2X1_594/A 0.02fF
C59687 POR2X1_430/a_16_28# POR2X1_430/A 0.05fF
C59688 PAND2X1_94/A PAND2X1_54/a_76_28# 0.02fF
C59689 POR2X1_819/a_16_28# POR2X1_94/A 0.00fF
C59690 PAND2X1_217/B POR2X1_60/A 0.05fF
C59691 POR2X1_567/A POR2X1_567/a_16_28# 0.03fF
C59692 PAND2X1_656/B VDD 0.04fF
C59693 POR2X1_730/Y POR2X1_440/CTRL2 0.01fF
C59694 POR2X1_566/A PAND2X1_258/CTRL2 0.14fF
C59695 PAND2X1_23/Y PAND2X1_67/CTRL2 0.01fF
C59696 PAND2X1_459/CTRL2 POR2X1_750/B 0.01fF
C59697 POR2X1_814/A POR2X1_228/Y 2.30fF
C59698 POR2X1_29/CTRL2 POR2X1_29/A 0.01fF
C59699 D_INPUT_0 PAND2X1_206/O 0.03fF
C59700 POR2X1_490/Y PAND2X1_216/CTRL 0.01fF
C59701 POR2X1_257/A POR2X1_238/Y 0.03fF
C59702 POR2X1_257/A PAND2X1_658/B 0.01fF
C59703 PAND2X1_211/CTRL2 PAND2X1_357/Y 0.01fF
C59704 D_INPUT_0 POR2X1_435/Y 0.03fF
C59705 POR2X1_818/Y POR2X1_415/a_16_28# 0.02fF
C59706 POR2X1_42/O POR2X1_20/B 0.02fF
C59707 PAND2X1_58/A PAND2X1_90/Y 0.10fF
C59708 PAND2X1_286/O POR2X1_283/Y 0.01fF
C59709 PAND2X1_405/O PAND2X1_737/B 0.02fF
C59710 PAND2X1_93/B POR2X1_661/B 0.03fF
C59711 PAND2X1_661/Y POR2X1_681/CTRL 0.03fF
C59712 PAND2X1_205/Y POR2X1_72/B 0.03fF
C59713 POR2X1_83/B POR2X1_250/CTRL2 0.01fF
C59714 POR2X1_466/A POR2X1_724/a_16_28# 0.08fF
C59715 PAND2X1_803/A PAND2X1_444/Y 0.02fF
C59716 POR2X1_614/A POR2X1_676/CTRL 0.01fF
C59717 PAND2X1_139/a_56_28# POR2X1_40/Y 0.00fF
C59718 POR2X1_852/B PAND2X1_41/B 0.07fF
C59719 PAND2X1_340/B PAND2X1_6/A 0.03fF
C59720 PAND2X1_212/CTRL2 PAND2X1_357/Y 0.01fF
C59721 PAND2X1_691/Y PAND2X1_644/O 0.01fF
C59722 PAND2X1_73/Y PAND2X1_57/B 0.17fF
C59723 POR2X1_66/A POR2X1_546/B 0.03fF
C59724 POR2X1_473/CTRL PAND2X1_32/B 0.05fF
C59725 POR2X1_60/A VDD 5.96fF
C59726 POR2X1_60/A PAND2X1_788/CTRL 0.09fF
C59727 POR2X1_824/Y POR2X1_411/B 0.03fF
C59728 PAND2X1_678/CTRL PAND2X1_175/B 0.01fF
C59729 PAND2X1_276/CTRL PAND2X1_390/Y 0.01fF
C59730 POR2X1_296/B POR2X1_723/a_16_28# 0.09fF
C59731 POR2X1_645/CTRL POR2X1_330/Y 0.15fF
C59732 PAND2X1_92/m4_208_n4# POR2X1_66/A 0.06fF
C59733 PAND2X1_540/O POR2X1_106/Y 0.02fF
C59734 POR2X1_624/Y POR2X1_68/B 0.03fF
C59735 POR2X1_634/A VDD 4.37fF
C59736 POR2X1_814/B POR2X1_105/Y 0.04fF
C59737 POR2X1_66/B PAND2X1_131/O 0.03fF
C59738 PAND2X1_6/Y POR2X1_841/B 0.12fF
C59739 POR2X1_591/A VDD 0.09fF
C59740 PAND2X1_9/Y POR2X1_408/Y 0.03fF
C59741 POR2X1_260/B POR2X1_702/A 0.04fF
C59742 PAND2X1_95/B PAND2X1_64/a_76_28# 0.05fF
C59743 POR2X1_76/A PAND2X1_311/O 0.08fF
C59744 PAND2X1_859/A POR2X1_236/Y 0.05fF
C59745 PAND2X1_783/Y PAND2X1_803/A 0.17fF
C59746 PAND2X1_556/B POR2X1_40/Y 0.02fF
C59747 PAND2X1_211/A POR2X1_236/Y 0.02fF
C59748 POR2X1_467/Y POR2X1_220/Y 0.02fF
C59749 POR2X1_65/A POR2X1_122/Y 0.03fF
C59750 POR2X1_822/a_16_28# POR2X1_40/Y 0.03fF
C59751 POR2X1_186/Y POR2X1_776/a_16_28# 0.02fF
C59752 POR2X1_208/A PAND2X1_39/B 0.03fF
C59753 POR2X1_623/B POR2X1_55/Y 0.00fF
C59754 POR2X1_407/A POR2X1_66/A 0.03fF
C59755 POR2X1_102/Y PAND2X1_215/B 0.00fF
C59756 POR2X1_287/CTRL POR2X1_733/A 0.13fF
C59757 PAND2X1_790/CTRL2 POR2X1_7/A 0.08fF
C59758 PAND2X1_73/Y POR2X1_285/A 0.07fF
C59759 PAND2X1_653/Y POR2X1_23/Y 0.03fF
C59760 POR2X1_116/A POR2X1_276/Y 0.05fF
C59761 POR2X1_269/O POR2X1_741/Y 0.01fF
C59762 POR2X1_383/A PAND2X1_271/CTRL2 0.03fF
C59763 POR2X1_477/A POR2X1_174/A 0.00fF
C59764 POR2X1_404/a_16_28# POR2X1_403/Y 0.11fF
C59765 PAND2X1_48/B POR2X1_489/B 0.01fF
C59766 POR2X1_121/B POR2X1_733/A 0.05fF
C59767 PAND2X1_792/CTRL2 POR2X1_759/Y 0.00fF
C59768 PAND2X1_859/CTRL VDD -0.00fF
C59769 POR2X1_462/O POR2X1_559/A 0.18fF
C59770 POR2X1_41/B PAND2X1_35/B 0.00fF
C59771 PAND2X1_230/O POR2X1_785/A 0.15fF
C59772 POR2X1_556/A POR2X1_260/A 1.61fF
C59773 PAND2X1_208/O PAND2X1_198/Y 0.02fF
C59774 PAND2X1_456/O POR2X1_516/B 0.00fF
C59775 PAND2X1_6/Y PAND2X1_603/O 0.06fF
C59776 POR2X1_121/O POR2X1_260/B 0.02fF
C59777 POR2X1_52/A POR2X1_750/B 0.05fF
C59778 PAND2X1_96/B D_INPUT_0 0.03fF
C59779 POR2X1_48/A POR2X1_425/Y 0.00fF
C59780 PAND2X1_94/A POR2X1_628/Y 0.00fF
C59781 PAND2X1_3/A D_INPUT_6 0.04fF
C59782 PAND2X1_733/CTRL POR2X1_7/B 0.01fF
C59783 POR2X1_274/CTRL POR2X1_573/A 0.01fF
C59784 POR2X1_496/O POR2X1_789/B 0.09fF
C59785 POR2X1_435/Y PAND2X1_90/Y 0.10fF
C59786 POR2X1_102/Y PAND2X1_6/A 0.07fF
C59787 PAND2X1_73/Y POR2X1_828/A 0.39fF
C59788 POR2X1_860/O PAND2X1_39/B 0.01fF
C59789 PAND2X1_204/CTRL PAND2X1_735/Y 0.04fF
C59790 POR2X1_821/CTRL POR2X1_236/Y 0.05fF
C59791 POR2X1_514/O PAND2X1_20/A 0.01fF
C59792 POR2X1_667/A POR2X1_518/Y 0.01fF
C59793 POR2X1_296/B POR2X1_501/B 0.09fF
C59794 PAND2X1_6/Y PAND2X1_626/CTRL 0.01fF
C59795 POR2X1_614/A POR2X1_806/CTRL 0.00fF
C59796 POR2X1_651/Y POR2X1_725/CTRL 0.02fF
C59797 POR2X1_20/B PAND2X1_853/B 0.09fF
C59798 POR2X1_130/A VDD 6.38fF
C59799 POR2X1_599/A POR2X1_40/Y 0.05fF
C59800 POR2X1_642/O POR2X1_734/A 0.03fF
C59801 POR2X1_76/B PAND2X1_72/A 0.03fF
C59802 POR2X1_96/A POR2X1_236/Y 0.44fF
C59803 POR2X1_54/Y POR2X1_753/CTRL 0.02fF
C59804 POR2X1_272/a_16_28# POR2X1_42/Y 0.03fF
C59805 POR2X1_630/a_16_28# POR2X1_510/Y 0.01fF
C59806 POR2X1_41/B PAND2X1_499/Y 0.04fF
C59807 POR2X1_688/a_56_344# POR2X1_294/A 0.00fF
C59808 POR2X1_49/Y POR2X1_238/Y 0.07fF
C59809 POR2X1_566/A VDD 5.97fF
C59810 POR2X1_814/A PAND2X1_122/O 0.05fF
C59811 PAND2X1_241/Y POR2X1_669/B 0.03fF
C59812 PAND2X1_821/O PAND2X1_41/B 0.08fF
C59813 POR2X1_628/Y PAND2X1_507/O 0.00fF
C59814 PAND2X1_453/CTRL2 POR2X1_511/Y 0.03fF
C59815 POR2X1_634/A PAND2X1_32/B 0.02fF
C59816 POR2X1_114/B POR2X1_405/O 0.01fF
C59817 POR2X1_661/a_16_28# POR2X1_661/B 0.03fF
C59818 POR2X1_244/B POR2X1_192/Y 0.05fF
C59819 PAND2X1_231/a_76_28# POR2X1_293/Y 0.02fF
C59820 PAND2X1_401/CTRL2 POR2X1_5/Y 0.00fF
C59821 POR2X1_448/CTRL2 PAND2X1_60/B 0.00fF
C59822 POR2X1_66/B POR2X1_194/CTRL 0.00fF
C59823 PAND2X1_651/Y PAND2X1_465/O 0.00fF
C59824 POR2X1_647/B POR2X1_774/A 0.03fF
C59825 POR2X1_278/Y POR2X1_79/Y 0.12fF
C59826 POR2X1_720/B POR2X1_720/A 0.00fF
C59827 POR2X1_271/CTRL2 POR2X1_153/Y 0.00fF
C59828 POR2X1_13/A PAND2X1_768/O 0.15fF
C59829 POR2X1_634/A POR2X1_711/O 0.08fF
C59830 POR2X1_707/A POR2X1_407/Y 0.01fF
C59831 PAND2X1_735/Y POR2X1_46/Y 0.10fF
C59832 POR2X1_333/A POR2X1_478/B 0.19fF
C59833 POR2X1_325/CTRL POR2X1_78/A 0.01fF
C59834 PAND2X1_717/A POR2X1_39/B 0.03fF
C59835 PAND2X1_809/A VDD 0.08fF
C59836 PAND2X1_697/CTRL2 PAND2X1_65/B 0.01fF
C59837 POR2X1_388/CTRL POR2X1_814/B 0.01fF
C59838 POR2X1_379/CTRL2 PAND2X1_20/A 0.00fF
C59839 POR2X1_634/A PAND2X1_764/CTRL2 0.06fF
C59840 POR2X1_114/O POR2X1_475/A 0.01fF
C59841 POR2X1_210/Y POR2X1_750/B 0.06fF
C59842 POR2X1_48/A PAND2X1_341/Y 0.03fF
C59843 PAND2X1_568/a_16_344# POR2X1_7/B 0.02fF
C59844 PAND2X1_738/Y POR2X1_55/Y 0.05fF
C59845 PAND2X1_207/CTRL PAND2X1_123/Y 0.01fF
C59846 POR2X1_51/A POR2X1_408/O 0.01fF
C59847 POR2X1_567/B POR2X1_317/B 0.05fF
C59848 POR2X1_154/CTRL POR2X1_803/A 0.01fF
C59849 POR2X1_332/B PAND2X1_111/CTRL2 0.01fF
C59850 POR2X1_616/O POR2X1_129/Y 0.01fF
C59851 POR2X1_201/CTRL2 POR2X1_201/Y 0.02fF
C59852 POR2X1_46/Y PAND2X1_493/Y 0.05fF
C59853 POR2X1_579/Y POR2X1_776/B 0.03fF
C59854 POR2X1_641/m4_208_n4# PAND2X1_60/B 0.09fF
C59855 POR2X1_624/Y PAND2X1_143/O 0.01fF
C59856 VDD PAND2X1_111/O 0.00fF
C59857 POR2X1_78/B POR2X1_712/A 0.03fF
C59858 PAND2X1_218/a_76_28# PAND2X1_741/B 0.02fF
C59859 POR2X1_83/B PAND2X1_593/Y 0.12fF
C59860 POR2X1_493/O PAND2X1_41/B 0.07fF
C59861 PAND2X1_96/B PAND2X1_90/Y 0.21fF
C59862 POR2X1_566/A POR2X1_741/Y 0.04fF
C59863 POR2X1_614/A POR2X1_549/a_16_28# 0.08fF
C59864 PAND2X1_844/O D_INPUT_0 0.18fF
C59865 PAND2X1_842/CTRL PAND2X1_389/Y 0.01fF
C59866 POR2X1_131/CTRL PAND2X1_140/Y 0.01fF
C59867 PAND2X1_90/Y POR2X1_736/CTRL2 0.16fF
C59868 POR2X1_786/A POR2X1_294/B 0.05fF
C59869 VDD POR2X1_844/B 0.04fF
C59870 PAND2X1_857/A POR2X1_72/B 0.03fF
C59871 POR2X1_311/a_16_28# POR2X1_102/Y 0.12fF
C59872 POR2X1_448/A POR2X1_788/B 0.01fF
C59873 PAND2X1_793/Y POR2X1_45/Y 0.03fF
C59874 POR2X1_78/A PAND2X1_528/a_76_28# 0.02fF
C59875 PAND2X1_819/CTRL2 POR2X1_750/B 0.03fF
C59876 POR2X1_272/a_76_344# PAND2X1_349/A 0.00fF
C59877 POR2X1_496/Y PAND2X1_748/m4_208_n4# 0.15fF
C59878 POR2X1_368/Y POR2X1_13/A 0.01fF
C59879 POR2X1_68/A PAND2X1_524/O 0.04fF
C59880 POR2X1_72/B PAND2X1_374/O 0.03fF
C59881 POR2X1_130/A PAND2X1_32/B 0.28fF
C59882 POR2X1_38/Y PAND2X1_84/Y 0.03fF
C59883 PAND2X1_90/A POR2X1_264/Y 0.03fF
C59884 POR2X1_807/a_56_344# PAND2X1_48/A 0.00fF
C59885 POR2X1_166/CTRL2 PAND2X1_738/Y 0.06fF
C59886 POR2X1_16/A PAND2X1_195/O 0.11fF
C59887 PAND2X1_540/O PAND2X1_114/B 0.16fF
C59888 VDD POR2X1_573/A 0.58fF
C59889 POR2X1_303/a_76_344# POR2X1_274/A 0.01fF
C59890 POR2X1_516/B POR2X1_73/Y 0.03fF
C59891 POR2X1_186/Y POR2X1_151/CTRL2 0.04fF
C59892 POR2X1_566/A PAND2X1_32/B 0.05fF
C59893 PAND2X1_232/CTRL2 PAND2X1_41/B 0.01fF
C59894 PAND2X1_56/Y POR2X1_733/A 0.10fF
C59895 PAND2X1_803/CTRL POR2X1_60/A 0.11fF
C59896 POR2X1_72/B POR2X1_260/A 0.03fF
C59897 POR2X1_494/Y POR2X1_56/Y 0.03fF
C59898 POR2X1_683/Y POR2X1_42/Y 0.12fF
C59899 POR2X1_7/A POR2X1_236/Y 0.12fF
C59900 POR2X1_332/Y POR2X1_241/B 0.02fF
C59901 PAND2X1_230/O POR2X1_186/B 0.01fF
C59902 POR2X1_327/Y POR2X1_806/O 0.02fF
C59903 PAND2X1_718/Y POR2X1_394/A 0.00fF
C59904 PAND2X1_350/CTRL INPUT_0 0.05fF
C59905 PAND2X1_254/O POR2X1_253/Y 0.53fF
C59906 PAND2X1_20/A PAND2X1_586/O 0.00fF
C59907 POR2X1_532/A PAND2X1_386/Y 0.03fF
C59908 POR2X1_135/O D_INPUT_0 0.02fF
C59909 PAND2X1_852/B POR2X1_293/Y 0.01fF
C59910 POR2X1_515/O POR2X1_276/A 0.09fF
C59911 PAND2X1_494/O POR2X1_264/Y 0.04fF
C59912 PAND2X1_496/O D_INPUT_1 0.05fF
C59913 POR2X1_566/A POR2X1_336/a_16_28# 0.02fF
C59914 POR2X1_774/O VDD 0.00fF
C59915 POR2X1_68/A D_GATE_222 0.03fF
C59916 PAND2X1_55/Y POR2X1_702/A 0.03fF
C59917 POR2X1_101/a_16_28# POR2X1_814/B 0.03fF
C59918 PAND2X1_318/CTRL2 PAND2X1_787/A 0.03fF
C59919 PAND2X1_358/A POR2X1_40/Y 0.03fF
C59920 PAND2X1_521/m4_208_n4# INPUT_0 0.06fF
C59921 POR2X1_414/CTRL POR2X1_4/Y 0.01fF
C59922 PAND2X1_523/O PAND2X1_844/B 0.03fF
C59923 POR2X1_40/Y POR2X1_599/O 0.02fF
C59924 POR2X1_193/O POR2X1_631/B 0.03fF
C59925 PAND2X1_6/Y POR2X1_114/B 0.03fF
C59926 POR2X1_16/A POR2X1_666/A 0.03fF
C59927 POR2X1_52/A POR2X1_824/Y 0.01fF
C59928 POR2X1_119/Y POR2X1_102/Y 3.02fF
C59929 POR2X1_16/A POR2X1_177/Y 0.00fF
C59930 POR2X1_54/Y POR2X1_8/CTRL2 0.01fF
C59931 INPUT_0 POR2X1_520/A 0.05fF
C59932 POR2X1_61/A PAND2X1_58/A 0.02fF
C59933 POR2X1_501/O POR2X1_501/B 0.02fF
C59934 POR2X1_501/CTRL2 POR2X1_573/A 0.01fF
C59935 POR2X1_593/O POR2X1_593/B 0.00fF
C59936 POR2X1_272/Y PAND2X1_301/CTRL2 0.01fF
C59937 POR2X1_744/CTRL VDD 0.00fF
C59938 POR2X1_456/B POR2X1_552/Y 0.01fF
C59939 PAND2X1_684/O PAND2X1_90/Y 0.18fF
C59940 POR2X1_582/m4_208_n4# INPUT_4 0.09fF
C59941 PAND2X1_664/CTRL2 PAND2X1_645/B 0.05fF
C59942 PAND2X1_111/O PAND2X1_32/B 0.04fF
C59943 PAND2X1_445/a_16_344# POR2X1_90/Y 0.01fF
C59944 POR2X1_741/Y POR2X1_573/A 0.03fF
C59945 POR2X1_596/CTRL VDD 0.00fF
C59946 POR2X1_800/A POR2X1_783/Y 0.00fF
C59947 POR2X1_149/B POR2X1_788/B 0.09fF
C59948 POR2X1_140/B POR2X1_532/A 0.00fF
C59949 POR2X1_121/O PAND2X1_55/Y 0.02fF
C59950 POR2X1_136/Y POR2X1_55/Y 0.34fF
C59951 POR2X1_844/B PAND2X1_32/B 0.03fF
C59952 POR2X1_65/A PAND2X1_508/Y 0.03fF
C59953 POR2X1_154/a_76_344# POR2X1_855/B 0.00fF
C59954 POR2X1_804/A PAND2X1_69/A 0.05fF
C59955 POR2X1_407/A POR2X1_532/A 0.03fF
C59956 POR2X1_566/A PAND2X1_253/O 0.24fF
C59957 POR2X1_413/A PAND2X1_647/O 0.02fF
C59958 PAND2X1_865/Y PAND2X1_575/B 0.00fF
C59959 PAND2X1_499/Y PAND2X1_861/a_76_28# 0.03fF
C59960 POR2X1_257/Y POR2X1_258/Y 0.18fF
C59961 PAND2X1_69/O PAND2X1_69/A -0.00fF
C59962 PAND2X1_6/Y PAND2X1_424/CTRL 0.01fF
C59963 POR2X1_383/A POR2X1_733/A 0.10fF
C59964 POR2X1_853/A POR2X1_578/a_16_28# 0.03fF
C59965 POR2X1_334/B POR2X1_383/A 0.05fF
C59966 PAND2X1_299/CTRL POR2X1_188/Y 0.01fF
C59967 POR2X1_327/Y POR2X1_78/B 0.07fF
C59968 PAND2X1_546/O POR2X1_526/Y -0.00fF
C59969 POR2X1_344/Y VDD 0.10fF
C59970 PAND2X1_94/A POR2X1_247/O 0.01fF
C59971 POR2X1_573/A PAND2X1_32/B 0.03fF
C59972 POR2X1_740/Y POR2X1_738/A 0.02fF
C59973 POR2X1_16/A POR2X1_669/O 0.01fF
C59974 POR2X1_857/B PAND2X1_503/O 0.02fF
C59975 PAND2X1_691/Y POR2X1_761/O 0.01fF
C59976 PAND2X1_675/O PAND2X1_557/A 0.08fF
C59977 POR2X1_529/Y POR2X1_816/A 0.02fF
C59978 PAND2X1_6/Y POR2X1_222/A 0.02fF
C59979 POR2X1_283/A POR2X1_248/CTRL2 0.01fF
C59980 POR2X1_406/a_16_28# PAND2X1_737/B 0.01fF
C59981 POR2X1_113/Y PAND2X1_153/CTRL 0.01fF
C59982 POR2X1_16/A PAND2X1_552/B 0.03fF
C59983 PAND2X1_140/A PAND2X1_113/CTRL2 0.01fF
C59984 POR2X1_539/O POR2X1_741/Y 0.00fF
C59985 POR2X1_220/B POR2X1_161/a_76_344# 0.01fF
C59986 POR2X1_39/Y POR2X1_42/Y 0.02fF
C59987 POR2X1_255/CTRL PAND2X1_840/Y 0.06fF
C59988 POR2X1_709/CTRL PAND2X1_69/A 0.01fF
C59989 POR2X1_130/A POR2X1_557/CTRL 0.01fF
C59990 PAND2X1_814/O POR2X1_283/A -0.00fF
C59991 POR2X1_278/Y PAND2X1_730/A 0.03fF
C59992 POR2X1_132/CTRL2 POR2X1_7/B 0.03fF
C59993 POR2X1_754/Y POR2X1_90/CTRL -0.02fF
C59994 POR2X1_416/B PAND2X1_733/CTRL2 0.05fF
C59995 VDD PAND2X1_167/CTRL 0.00fF
C59996 PAND2X1_804/CTRL PAND2X1_860/A 0.01fF
C59997 POR2X1_825/Y D_INPUT_0 0.03fF
C59998 POR2X1_673/Y POR2X1_844/B 0.03fF
C59999 PAND2X1_6/Y PAND2X1_300/a_76_28# 0.03fF
C60000 INPUT_1 POR2X1_409/CTRL 0.01fF
C60001 POR2X1_61/B POR2X1_507/A 0.03fF
C60002 PAND2X1_639/Y POR2X1_13/A 0.13fF
C60003 POR2X1_7/B PAND2X1_716/B 0.03fF
C60004 PAND2X1_414/O INPUT_3 0.03fF
C60005 PAND2X1_562/O POR2X1_394/A 0.02fF
C60006 PAND2X1_41/B POR2X1_180/Y 0.01fF
C60007 POR2X1_334/B PAND2X1_71/Y 0.03fF
C60008 POR2X1_579/Y POR2X1_192/B 0.14fF
C60009 POR2X1_711/a_16_28# POR2X1_710/Y 0.05fF
C60010 PAND2X1_21/CTRL D_INPUT_4 0.00fF
C60011 POR2X1_572/B PAND2X1_48/A 0.06fF
C60012 POR2X1_509/A POR2X1_227/O 0.01fF
C60013 POR2X1_141/CTRL POR2X1_343/Y -0.00fF
C60014 POR2X1_258/Y PAND2X1_854/A 0.02fF
C60015 PAND2X1_390/Y PAND2X1_332/Y 0.03fF
C60016 POR2X1_814/A POR2X1_454/A 0.07fF
C60017 POR2X1_71/Y PAND2X1_865/Y 0.00fF
C60018 PAND2X1_6/Y PAND2X1_482/O 0.08fF
C60019 POR2X1_346/CTRL POR2X1_507/A 0.04fF
C60020 POR2X1_62/Y PAND2X1_341/a_56_28# 0.00fF
C60021 POR2X1_264/Y POR2X1_572/Y 0.01fF
C60022 POR2X1_447/B PAND2X1_625/CTRL2 0.04fF
C60023 POR2X1_545/A POR2X1_192/B 0.12fF
C60024 PAND2X1_865/Y POR2X1_42/Y 0.07fF
C60025 POR2X1_702/O POR2X1_260/A 0.02fF
C60026 POR2X1_614/A PAND2X1_48/A 0.03fF
C60027 PAND2X1_771/B PAND2X1_769/Y 0.02fF
C60028 POR2X1_10/CTRL2 PAND2X1_63/B 0.01fF
C60029 POR2X1_48/A PAND2X1_717/A 0.03fF
C60030 POR2X1_96/B INPUT_1 0.06fF
C60031 POR2X1_41/B POR2X1_39/B 21.97fF
C60032 POR2X1_119/Y POR2X1_531/Y 0.10fF
C60033 POR2X1_317/Y POR2X1_192/B 0.03fF
C60034 POR2X1_108/Y PAND2X1_114/O -0.00fF
C60035 POR2X1_804/A POR2X1_512/CTRL 0.00fF
C60036 PAND2X1_139/CTRL POR2X1_184/Y 0.00fF
C60037 POR2X1_265/Y POR2X1_73/Y 0.03fF
C60038 POR2X1_560/CTRL POR2X1_844/B 0.01fF
C60039 PAND2X1_440/CTRL PAND2X1_793/Y 0.01fF
C60040 POR2X1_730/Y POR2X1_727/a_16_28# 0.02fF
C60041 POR2X1_290/O POR2X1_234/A 0.01fF
C60042 PAND2X1_352/O PAND2X1_357/Y 0.02fF
C60043 POR2X1_271/A POR2X1_7/A 3.11fF
C60044 POR2X1_394/A PAND2X1_349/A 0.05fF
C60045 POR2X1_334/Y POR2X1_510/Y 0.07fF
C60046 POR2X1_394/A PAND2X1_63/B 0.05fF
C60047 POR2X1_703/A POR2X1_543/CTRL 0.03fF
C60048 POR2X1_416/B POR2X1_628/CTRL2 0.01fF
C60049 POR2X1_96/B POR2X1_153/Y 0.05fF
C60050 POR2X1_72/CTRL2 POR2X1_816/A 0.03fF
C60051 POR2X1_62/Y PAND2X1_338/B 0.03fF
C60052 POR2X1_740/Y POR2X1_731/Y 0.00fF
C60053 PAND2X1_501/O POR2X1_494/Y 0.00fF
C60054 POR2X1_446/B POR2X1_222/CTRL2 0.01fF
C60055 PAND2X1_98/O POR2X1_93/Y 0.08fF
C60056 POR2X1_23/Y POR2X1_20/B 0.29fF
C60057 POR2X1_172/Y POR2X1_171/Y 0.00fF
C60058 POR2X1_628/a_76_344# POR2X1_39/B 0.00fF
C60059 PAND2X1_787/Y POR2X1_173/Y 0.23fF
C60060 POR2X1_303/CTRL POR2X1_228/Y 0.01fF
C60061 PAND2X1_6/Y POR2X1_513/A 0.03fF
C60062 POR2X1_43/B PAND2X1_840/Y 0.20fF
C60063 POR2X1_145/a_16_28# POR2X1_77/Y 0.02fF
C60064 PAND2X1_82/a_16_344# POR2X1_84/A 0.02fF
C60065 POR2X1_186/CTRL POR2X1_186/B 0.00fF
C60066 POR2X1_68/B PAND2X1_517/a_56_28# 0.00fF
C60067 POR2X1_260/B PAND2X1_609/O 0.01fF
C60068 POR2X1_341/Y POR2X1_568/B 0.03fF
C60069 POR2X1_329/A POR2X1_72/B 0.13fF
C60070 POR2X1_452/Y POR2X1_809/a_16_28# 0.03fF
C60071 POR2X1_130/a_76_344# POR2X1_244/Y 0.01fF
C60072 PAND2X1_59/CTRL D_INPUT_4 0.01fF
C60073 POR2X1_184/CTRL POR2X1_91/Y 0.09fF
C60074 PAND2X1_619/CTRL2 POR2X1_29/A 0.03fF
C60075 POR2X1_83/B PAND2X1_201/O 0.04fF
C60076 POR2X1_532/CTRL PAND2X1_60/B 0.00fF
C60077 POR2X1_114/B PAND2X1_52/B 0.06fF
C60078 POR2X1_652/CTRL2 PAND2X1_72/A 0.01fF
C60079 POR2X1_416/B PAND2X1_324/O 0.05fF
C60080 POR2X1_451/A INPUT_4 0.25fF
C60081 POR2X1_99/B POR2X1_259/O 0.00fF
C60082 POR2X1_62/Y PAND2X1_341/Y 0.01fF
C60083 POR2X1_440/Y POR2X1_726/a_16_28# 0.08fF
C60084 POR2X1_866/A POR2X1_807/CTRL 0.07fF
C60085 POR2X1_326/A POR2X1_186/B 0.15fF
C60086 POR2X1_60/A PAND2X1_9/Y 0.03fF
C60087 D_INPUT_7 PAND2X1_587/Y 0.04fF
C60088 POR2X1_441/Y POR2X1_40/Y 4.35fF
C60089 POR2X1_222/A POR2X1_632/Y 0.03fF
C60090 POR2X1_327/Y POR2X1_294/A 0.03fF
C60091 PAND2X1_43/CTRL2 POR2X1_330/Y 0.03fF
C60092 POR2X1_326/A POR2X1_802/A 0.03fF
C60093 POR2X1_99/CTRL2 PAND2X1_65/Y 0.01fF
C60094 POR2X1_73/Y POR2X1_167/Y 0.01fF
C60095 POR2X1_633/a_16_28# POR2X1_734/A 0.06fF
C60096 POR2X1_20/B POR2X1_312/Y 0.04fF
C60097 POR2X1_800/O POR2X1_452/Y 0.01fF
C60098 POR2X1_383/A POR2X1_343/a_16_28# 0.01fF
C60099 POR2X1_41/B POR2X1_827/O 0.01fF
C60100 POR2X1_577/O POR2X1_568/A 0.10fF
C60101 PAND2X1_72/A POR2X1_704/CTRL2 0.00fF
C60102 POR2X1_612/Y POR2X1_413/CTRL 0.08fF
C60103 INPUT_3 POR2X1_293/CTRL 0.00fF
C60104 POR2X1_270/Y POR2X1_269/A 0.01fF
C60105 POR2X1_291/O POR2X1_39/B 0.18fF
C60106 POR2X1_466/A POR2X1_436/B 0.63fF
C60107 POR2X1_864/A POR2X1_855/A 0.44fF
C60108 PAND2X1_58/A PAND2X1_591/CTRL2 0.01fF
C60109 POR2X1_48/A POR2X1_484/m4_208_n4# 0.08fF
C60110 PAND2X1_60/B POR2X1_343/B 0.07fF
C60111 POR2X1_360/A POR2X1_814/A 0.02fF
C60112 POR2X1_661/A POR2X1_513/Y 0.02fF
C60113 PAND2X1_810/B VDD 0.20fF
C60114 POR2X1_119/Y POR2X1_74/Y 0.03fF
C60115 POR2X1_9/Y PAND2X1_6/A 0.61fF
C60116 PAND2X1_628/CTRL2 POR2X1_532/A 0.01fF
C60117 POR2X1_455/O POR2X1_341/A 0.05fF
C60118 POR2X1_37/CTRL2 D_INPUT_0 0.00fF
C60119 PAND2X1_466/B POR2X1_236/Y 0.03fF
C60120 POR2X1_66/B PAND2X1_3/A 0.01fF
C60121 PAND2X1_47/B PAND2X1_25/CTRL 0.13fF
C60122 POR2X1_78/B POR2X1_240/CTRL2 0.04fF
C60123 PAND2X1_120/CTRL POR2X1_77/Y 0.01fF
C60124 POR2X1_666/a_16_28# POR2X1_32/A 0.00fF
C60125 POR2X1_416/B POR2X1_129/Y 0.02fF
C60126 POR2X1_814/B POR2X1_240/a_16_28# 0.04fF
C60127 POR2X1_254/Y POR2X1_341/A 2.22fF
C60128 POR2X1_640/A POR2X1_260/B -0.00fF
C60129 POR2X1_81/O PAND2X1_573/B 0.01fF
C60130 PAND2X1_841/B POR2X1_271/B 0.49fF
C60131 POR2X1_482/Y POR2X1_669/B 0.05fF
C60132 PAND2X1_48/B PAND2X1_417/a_16_344# 0.02fF
C60133 POR2X1_655/Y POR2X1_296/B 0.01fF
C60134 PAND2X1_699/O POR2X1_43/B 0.01fF
C60135 POR2X1_698/Y POR2X1_158/B 0.03fF
C60136 PAND2X1_659/Y POR2X1_416/B 0.18fF
C60137 POR2X1_96/A POR2X1_679/Y 0.01fF
C60138 POR2X1_855/O POR2X1_855/A 0.01fF
C60139 POR2X1_319/A POR2X1_192/Y 0.05fF
C60140 POR2X1_536/m4_208_n4# POR2X1_250/A 0.12fF
C60141 PAND2X1_853/B POR2X1_589/Y 0.05fF
C60142 POR2X1_660/Y POR2X1_807/A 0.02fF
C60143 POR2X1_341/A POR2X1_575/B 0.03fF
C60144 POR2X1_168/A POR2X1_191/Y 0.05fF
C60145 POR2X1_69/m4_208_n4# PAND2X1_58/A 0.15fF
C60146 POR2X1_56/a_76_344# POR2X1_423/Y 0.01fF
C60147 PAND2X1_39/B POR2X1_198/B 0.03fF
C60148 PAND2X1_90/A POR2X1_624/Y 0.13fF
C60149 PAND2X1_9/Y POR2X1_204/CTRL 0.05fF
C60150 PAND2X1_246/CTRL2 POR2X1_205/A -0.02fF
C60151 PAND2X1_810/A PAND2X1_866/A 0.01fF
C60152 POR2X1_608/Y PAND2X1_90/Y 0.05fF
C60153 PAND2X1_666/CTRL POR2X1_130/A 0.03fF
C60154 PAND2X1_224/a_16_344# POR2X1_566/B 0.04fF
C60155 PAND2X1_75/O POR2X1_318/A 0.03fF
C60156 POR2X1_66/B POR2X1_654/B 0.03fF
C60157 PAND2X1_836/O POR2X1_20/B 0.04fF
C60158 POR2X1_60/A POR2X1_609/a_16_28# 0.02fF
C60159 POR2X1_278/Y POR2X1_263/Y 0.05fF
C60160 PAND2X1_236/O POR2X1_29/A -0.00fF
C60161 POR2X1_846/a_56_344# POR2X1_129/Y 0.00fF
C60162 POR2X1_68/A POR2X1_54/Y 0.76fF
C60163 POR2X1_41/B POR2X1_48/A 0.54fF
C60164 POR2X1_96/A POR2X1_626/CTRL 0.01fF
C60165 POR2X1_206/A POR2X1_296/B 0.07fF
C60166 POR2X1_188/A POR2X1_654/B 0.03fF
C60167 POR2X1_77/Y POR2X1_39/B 0.24fF
C60168 POR2X1_232/CTRL2 POR2X1_37/Y 0.03fF
C60169 POR2X1_241/B VDD 0.84fF
C60170 POR2X1_632/CTRL POR2X1_222/Y 0.00fF
C60171 POR2X1_68/A POR2X1_202/A 0.00fF
C60172 POR2X1_658/O PAND2X1_60/B 0.09fF
C60173 POR2X1_41/B POR2X1_225/CTRL2 0.03fF
C60174 POR2X1_130/A POR2X1_267/A 0.37fF
C60175 POR2X1_514/Y PAND2X1_93/B 0.06fF
C60176 PAND2X1_556/O VDD 0.00fF
C60177 PAND2X1_853/CTRL2 POR2X1_23/Y 0.01fF
C60178 POR2X1_719/A VDD 0.00fF
C60179 PAND2X1_644/Y POR2X1_759/m4_208_n4# 0.08fF
C60180 POR2X1_174/A POR2X1_190/Y 0.07fF
C60181 POR2X1_261/O PAND2X1_569/Y 0.02fF
C60182 POR2X1_471/A POR2X1_724/A 0.03fF
C60183 PAND2X1_654/O POR2X1_409/B 0.02fF
C60184 PAND2X1_6/Y POR2X1_629/CTRL 0.01fF
C60185 PAND2X1_118/CTRL2 POR2X1_66/A 0.03fF
C60186 PAND2X1_476/CTRL2 PAND2X1_473/Y 0.03fF
C60187 POR2X1_590/A POR2X1_776/B 0.03fF
C60188 PAND2X1_443/O POR2X1_90/Y 0.15fF
C60189 POR2X1_499/A POR2X1_569/A 0.03fF
C60190 POR2X1_297/CTRL2 PAND2X1_347/Y 0.01fF
C60191 POR2X1_750/A VDD 0.39fF
C60192 PAND2X1_333/CTRL2 POR2X1_5/Y 0.03fF
C60193 POR2X1_43/B PAND2X1_61/CTRL2 0.03fF
C60194 POR2X1_334/B PAND2X1_15/CTRL2 0.10fF
C60195 POR2X1_119/Y POR2X1_677/Y 0.03fF
C60196 POR2X1_407/A POR2X1_858/CTRL2 0.01fF
C60197 PAND2X1_478/Y POR2X1_236/Y 0.01fF
C60198 POR2X1_257/A POR2X1_387/Y 0.07fF
C60199 POR2X1_257/A POR2X1_695/CTRL 0.01fF
C60200 PAND2X1_56/CTRL2 POR2X1_330/Y 0.30fF
C60201 POR2X1_83/B PAND2X1_364/CTRL 0.01fF
C60202 POR2X1_322/CTRL2 POR2X1_83/B 0.03fF
C60203 POR2X1_306/Y VDD 0.21fF
C60204 POR2X1_389/A PAND2X1_609/CTRL2 0.01fF
C60205 PAND2X1_20/A POR2X1_465/B 0.03fF
C60206 POR2X1_632/CTRL POR2X1_532/A 0.01fF
C60207 PAND2X1_777/m4_208_n4# POR2X1_55/Y 0.12fF
C60208 POR2X1_596/A POR2X1_260/B 4.39fF
C60209 POR2X1_814/A POR2X1_579/B 0.16fF
C60210 PAND2X1_116/CTRL2 VDD 0.00fF
C60211 POR2X1_68/A POR2X1_346/A 0.00fF
C60212 POR2X1_13/A POR2X1_272/O 0.02fF
C60213 POR2X1_185/CTRL2 PAND2X1_73/Y 0.05fF
C60214 POR2X1_60/A PAND2X1_714/O 0.01fF
C60215 POR2X1_666/Y PAND2X1_719/O 0.08fF
C60216 PAND2X1_42/O POR2X1_547/B 0.00fF
C60217 POR2X1_303/a_16_28# POR2X1_325/A 0.03fF
C60218 POR2X1_13/A PAND2X1_390/Y 0.07fF
C60219 POR2X1_48/A POR2X1_256/Y 0.01fF
C60220 PAND2X1_473/B PAND2X1_736/CTRL 0.00fF
C60221 POR2X1_821/a_56_344# POR2X1_72/B 0.01fF
C60222 GATE_479 VDD 0.36fF
C60223 POR2X1_774/Y VDD 0.44fF
C60224 PAND2X1_403/B POR2X1_293/Y 0.17fF
C60225 POR2X1_590/A POR2X1_565/CTRL 0.01fF
C60226 POR2X1_105/Y VDD 0.21fF
C60227 POR2X1_102/Y PAND2X1_219/O 0.02fF
C60228 POR2X1_242/CTRL POR2X1_578/Y 0.00fF
C60229 POR2X1_502/A PAND2X1_278/O 0.01fF
C60230 POR2X1_728/a_16_28# POR2X1_330/Y 0.04fF
C60231 POR2X1_405/O POR2X1_405/Y 0.00fF
C60232 PAND2X1_40/CTRL2 PAND2X1_11/Y 0.01fF
C60233 POR2X1_569/CTRL POR2X1_355/B 0.03fF
C60234 POR2X1_413/A POR2X1_607/CTRL 0.01fF
C60235 POR2X1_65/A PAND2X1_564/a_16_344# 0.02fF
C60236 POR2X1_83/A POR2X1_83/B 0.89fF
C60237 PAND2X1_422/a_16_344# POR2X1_260/B 0.01fF
C60238 POR2X1_853/O PAND2X1_41/B 0.01fF
C60239 POR2X1_76/A POR2X1_569/A 0.09fF
C60240 POR2X1_511/Y PAND2X1_512/Y 0.01fF
C60241 PAND2X1_738/Y PAND2X1_180/CTRL 0.14fF
C60242 PAND2X1_671/CTRL POR2X1_54/Y 0.01fF
C60243 PAND2X1_859/a_56_28# INPUT_0 0.00fF
C60244 POR2X1_305/Y POR2X1_14/Y 0.00fF
C60245 POR2X1_237/Y POR2X1_102/Y 1.18fF
C60246 POR2X1_99/B POR2X1_814/A 0.03fF
C60247 POR2X1_855/B POR2X1_796/Y 0.01fF
C60248 POR2X1_327/Y POR2X1_116/A 0.08fF
C60249 POR2X1_267/A POR2X1_844/B 0.03fF
C60250 PAND2X1_245/CTRL2 POR2X1_68/B 0.00fF
C60251 POR2X1_355/a_16_28# POR2X1_192/Y 0.05fF
C60252 POR2X1_241/B PAND2X1_32/B 0.06fF
C60253 POR2X1_114/a_16_28# POR2X1_590/A 0.03fF
C60254 PAND2X1_23/Y PAND2X1_23/O 0.00fF
C60255 POR2X1_449/m4_208_n4# PAND2X1_90/Y 0.03fF
C60256 PAND2X1_824/O POR2X1_856/B 0.06fF
C60257 POR2X1_83/B POR2X1_90/Y 0.17fF
C60258 POR2X1_5/Y POR2X1_395/CTRL 0.01fF
C60259 POR2X1_708/B PAND2X1_90/Y 0.05fF
C60260 POR2X1_810/CTRL POR2X1_750/B 0.01fF
C60261 POR2X1_254/Y PAND2X1_48/CTRL 0.04fF
C60262 PAND2X1_438/CTRL2 VDD 0.00fF
C60263 PAND2X1_3/a_76_28# D_INPUT_5 0.01fF
C60264 POR2X1_843/CTRL2 PAND2X1_60/B 0.00fF
C60265 PAND2X1_616/O PAND2X1_6/A 0.02fF
C60266 PAND2X1_853/O POR2X1_40/Y 0.01fF
C60267 POR2X1_185/O POR2X1_188/A 0.00fF
C60268 PAND2X1_6/Y POR2X1_783/O 0.17fF
C60269 PAND2X1_56/Y POR2X1_593/B 0.01fF
C60270 POR2X1_164/CTRL POR2X1_40/Y 0.01fF
C60271 POR2X1_79/Y PAND2X1_730/B 0.00fF
C60272 PAND2X1_771/Y PAND2X1_578/O 0.02fF
C60273 POR2X1_304/CTRL POR2X1_329/A 0.03fF
C60274 PAND2X1_118/O PAND2X1_41/B 0.22fF
C60275 PAND2X1_55/Y POR2X1_830/A 0.03fF
C60276 POR2X1_67/A PAND2X1_154/CTRL2 0.13fF
C60277 POR2X1_49/Y POR2X1_90/a_16_28# 0.07fF
C60278 PAND2X1_658/CTRL POR2X1_816/A 0.01fF
C60279 PAND2X1_96/B POR2X1_634/CTRL 0.01fF
C60280 POR2X1_97/A POR2X1_854/B 0.05fF
C60281 PAND2X1_94/A POR2X1_558/B 0.35fF
C60282 PAND2X1_140/A PAND2X1_577/Y 0.10fF
C60283 POR2X1_120/CTRL2 POR2X1_294/B 0.03fF
C60284 POR2X1_639/Y POR2X1_634/A 0.07fF
C60285 POR2X1_748/A POR2X1_748/CTRL 0.01fF
C60286 POR2X1_504/Y POR2X1_628/a_16_28# 0.02fF
C60287 PAND2X1_632/B POR2X1_482/CTRL2 0.01fF
C60288 PAND2X1_651/Y PAND2X1_455/CTRL 0.02fF
C60289 POR2X1_734/A POR2X1_705/CTRL2 0.13fF
C60290 POR2X1_96/A POR2X1_230/Y 0.05fF
C60291 POR2X1_775/A PAND2X1_65/B 0.03fF
C60292 POR2X1_669/B PAND2X1_63/B 0.03fF
C60293 POR2X1_30/CTRL INPUT_7 0.01fF
C60294 POR2X1_83/CTRL D_INPUT_0 0.03fF
C60295 PAND2X1_669/CTRL POR2X1_750/Y 0.25fF
C60296 POR2X1_60/A PAND2X1_370/m4_208_n4# 0.05fF
C60297 POR2X1_599/A POR2X1_5/Y 0.05fF
C60298 POR2X1_741/Y POR2X1_733/O 0.00fF
C60299 POR2X1_786/A POR2X1_786/a_16_28# 0.03fF
C60300 POR2X1_277/CTRL2 POR2X1_46/Y 0.01fF
C60301 POR2X1_89/O POR2X1_394/A 0.04fF
C60302 POR2X1_83/B PAND2X1_154/CTRL 0.01fF
C60303 PAND2X1_97/CTRL POR2X1_394/A 0.08fF
C60304 POR2X1_278/Y PAND2X1_215/B 0.05fF
C60305 POR2X1_614/A POR2X1_193/Y 0.03fF
C60306 POR2X1_57/A POR2X1_72/B 0.27fF
C60307 POR2X1_537/Y POR2X1_841/a_16_28# 0.02fF
C60308 PAND2X1_638/B POR2X1_588/Y 0.07fF
C60309 PAND2X1_585/O PAND2X1_60/B 0.01fF
C60310 POR2X1_334/B INPUT_0 0.10fF
C60311 POR2X1_774/Y PAND2X1_32/B 0.03fF
C60312 PAND2X1_834/a_16_344# PAND2X1_658/B 0.02fF
C60313 PAND2X1_575/A INPUT_0 0.03fF
C60314 PAND2X1_417/CTRL POR2X1_169/A 0.00fF
C60315 POR2X1_865/B PAND2X1_41/B 0.03fF
C60316 POR2X1_65/A PAND2X1_640/a_16_344# 0.02fF
C60317 PAND2X1_41/B PAND2X1_88/Y 0.01fF
C60318 POR2X1_232/CTRL2 POR2X1_293/Y 0.01fF
C60319 GATE_479 POR2X1_694/a_16_28# 0.02fF
C60320 POR2X1_10/CTRL2 POR2X1_32/A 0.01fF
C60321 POR2X1_860/CTRL POR2X1_296/B 0.09fF
C60322 POR2X1_43/Y POR2X1_827/CTRL 0.00fF
C60323 POR2X1_502/A POR2X1_740/Y 0.03fF
C60324 POR2X1_497/Y POR2X1_56/Y 0.03fF
C60325 POR2X1_483/A POR2X1_786/Y 0.04fF
C60326 POR2X1_493/A POR2X1_557/B 0.03fF
C60327 INPUT_1 POR2X1_296/B 0.05fF
C60328 POR2X1_52/A PAND2X1_776/CTRL 0.01fF
C60329 PAND2X1_253/O POR2X1_241/B 0.03fF
C60330 POR2X1_78/A POR2X1_773/B 0.12fF
C60331 PAND2X1_57/B POR2X1_715/a_16_28# 0.03fF
C60332 POR2X1_71/Y POR2X1_494/Y 0.03fF
C60333 POR2X1_97/O POR2X1_78/A 0.01fF
C60334 PAND2X1_651/Y PAND2X1_84/CTRL 0.01fF
C60335 POR2X1_514/O VDD 0.00fF
C60336 POR2X1_505/O POR2X1_669/B 0.03fF
C60337 POR2X1_634/A POR2X1_769/Y 0.02fF
C60338 POR2X1_267/CTRL POR2X1_260/A 0.00fF
C60339 PAND2X1_217/B PAND2X1_175/B 0.05fF
C60340 POR2X1_334/B POR2X1_137/CTRL2 0.13fF
C60341 POR2X1_833/A PAND2X1_73/Y 0.07fF
C60342 PAND2X1_490/a_16_344# PAND2X1_85/Y 0.04fF
C60343 PAND2X1_57/B POR2X1_35/Y 0.03fF
C60344 PAND2X1_661/Y POR2X1_39/CTRL2 0.01fF
C60345 PAND2X1_286/O PAND2X1_568/B 0.05fF
C60346 PAND2X1_183/O POR2X1_732/B 0.02fF
C60347 PAND2X1_58/A POR2X1_592/A 0.01fF
C60348 POR2X1_83/B PAND2X1_732/A 0.03fF
C60349 POR2X1_283/A POR2X1_503/A 0.04fF
C60350 PAND2X1_435/O POR2X1_433/Y 0.01fF
C60351 POR2X1_673/CTRL2 POR2X1_260/A 0.03fF
C60352 POR2X1_579/Y PAND2X1_111/CTRL2 0.00fF
C60353 POR2X1_38/Y POR2X1_236/Y 0.12fF
C60354 PAND2X1_418/CTRL PAND2X1_52/B 0.01fF
C60355 PAND2X1_468/O PAND2X1_798/B 0.03fF
C60356 PAND2X1_76/Y POR2X1_91/Y 0.17fF
C60357 POR2X1_32/A POR2X1_394/A 5.01fF
C60358 POR2X1_65/A PAND2X1_551/O 0.01fF
C60359 POR2X1_29/A POR2X1_720/CTRL2 0.03fF
C60360 POR2X1_57/A PAND2X1_756/O 0.01fF
C60361 POR2X1_65/A POR2X1_283/A 0.07fF
C60362 POR2X1_52/A POR2X1_823/CTRL 0.01fF
C60363 POR2X1_57/A PAND2X1_520/CTRL2 0.02fF
C60364 PAND2X1_228/O PAND2X1_197/Y 0.00fF
C60365 PAND2X1_716/O PAND2X1_364/B 0.06fF
C60366 POR2X1_144/O POR2X1_669/B 0.03fF
C60367 POR2X1_786/O PAND2X1_60/B 0.03fF
C60368 POR2X1_515/O PAND2X1_60/B 0.01fF
C60369 POR2X1_305/Y POR2X1_55/Y 0.67fF
C60370 POR2X1_719/CTRL VDD 0.00fF
C60371 POR2X1_750/B PAND2X1_1/a_76_28# 0.01fF
C60372 VDD POR2X1_142/Y 0.32fF
C60373 POR2X1_499/A PAND2X1_72/A 0.03fF
C60374 PAND2X1_241/CTRL2 POR2X1_90/Y 0.01fF
C60375 POR2X1_335/B PAND2X1_57/B 0.03fF
C60376 POR2X1_549/a_76_344# POR2X1_383/A 0.01fF
C60377 POR2X1_590/A PAND2X1_48/A 0.16fF
C60378 POR2X1_52/A PAND2X1_814/CTRL 0.01fF
C60379 POR2X1_853/A POR2X1_170/CTRL 0.01fF
C60380 POR2X1_475/A POR2X1_276/Y 0.01fF
C60381 POR2X1_807/A POR2X1_308/B 0.02fF
C60382 POR2X1_208/A VDD 0.00fF
C60383 PAND2X1_175/B VDD 0.08fF
C60384 POR2X1_590/A POR2X1_192/B 0.16fF
C60385 POR2X1_57/A POR2X1_399/m4_208_n4# 0.07fF
C60386 PAND2X1_6/Y POR2X1_732/B 0.03fF
C60387 POR2X1_417/Y POR2X1_394/A 0.03fF
C60388 POR2X1_614/A PAND2X1_111/CTRL2 0.03fF
C60389 POR2X1_356/A POR2X1_540/A 0.05fF
C60390 POR2X1_684/Y POR2X1_669/B 0.02fF
C60391 PAND2X1_787/A POR2X1_46/Y 0.10fF
C60392 POR2X1_49/Y POR2X1_419/a_16_28# 0.06fF
C60393 POR2X1_700/O PAND2X1_711/A 0.01fF
C60394 POR2X1_68/A PAND2X1_29/CTRL 0.01fF
C60395 POR2X1_110/Y POR2X1_83/B 0.11fF
C60396 POR2X1_52/A POR2X1_92/O 0.01fF
C60397 POR2X1_343/Y PAND2X1_251/CTRL2 0.01fF
C60398 PAND2X1_137/a_56_28# POR2X1_132/Y 0.00fF
C60399 POR2X1_840/a_16_28# POR2X1_307/Y 0.03fF
C60400 POR2X1_57/A POR2X1_323/Y 0.01fF
C60401 POR2X1_5/Y POR2X1_6/CTRL 0.01fF
C60402 PAND2X1_553/B POR2X1_387/Y 0.10fF
C60403 PAND2X1_20/A POR2X1_557/O 0.01fF
C60404 INPUT_1 POR2X1_236/Y 0.12fF
C60405 PAND2X1_118/CTRL2 POR2X1_532/A 0.01fF
C60406 POR2X1_163/CTRL POR2X1_394/A 0.01fF
C60407 INPUT_1 PAND2X1_721/m4_208_n4# 0.15fF
C60408 PAND2X1_57/B PAND2X1_765/O 0.17fF
C60409 PAND2X1_96/B D_GATE_222 1.23fF
C60410 INPUT_1 POR2X1_547/B 0.03fF
C60411 POR2X1_296/B PAND2X1_136/CTRL 0.01fF
C60412 PAND2X1_20/A POR2X1_560/O 0.01fF
C60413 POR2X1_45/Y PAND2X1_702/O 0.02fF
C60414 INPUT_2 PAND2X1_6/A 5.96fF
C60415 POR2X1_514/O PAND2X1_32/B 0.01fF
C60416 POR2X1_48/A POR2X1_77/Y 0.11fF
C60417 PAND2X1_57/B PAND2X1_368/O 0.01fF
C60418 PAND2X1_865/Y PAND2X1_78/CTRL 0.01fF
C60419 POR2X1_57/A PAND2X1_547/CTRL2 0.01fF
C60420 POR2X1_16/A POR2X1_79/A 0.01fF
C60421 PAND2X1_388/Y PAND2X1_552/B 0.01fF
C60422 POR2X1_590/A PAND2X1_102/CTRL2 0.00fF
C60423 POR2X1_416/B POR2X1_37/Y 0.56fF
C60424 POR2X1_138/a_16_28# POR2X1_318/A 0.07fF
C60425 POR2X1_366/Y POR2X1_854/B 0.10fF
C60426 POR2X1_236/Y POR2X1_153/Y 0.12fF
C60427 D_GATE_366 POR2X1_319/Y 0.12fF
C60428 POR2X1_79/CTRL2 PAND2X1_798/B 0.01fF
C60429 POR2X1_750/B POR2X1_540/Y 0.03fF
C60430 POR2X1_383/A PAND2X1_530/CTRL 0.00fF
C60431 POR2X1_16/A PAND2X1_468/CTRL2 0.07fF
C60432 POR2X1_572/O POR2X1_260/A 0.01fF
C60433 POR2X1_16/A POR2X1_79/Y 0.03fF
C60434 POR2X1_384/A POR2X1_236/Y 0.03fF
C60435 PAND2X1_69/A PAND2X1_311/O 0.06fF
C60436 PAND2X1_57/B PAND2X1_701/CTRL 0.02fF
C60437 POR2X1_57/A PAND2X1_835/Y 0.00fF
C60438 PAND2X1_76/Y POR2X1_109/Y 0.00fF
C60439 PAND2X1_41/B PAND2X1_165/a_16_344# 0.02fF
C60440 POR2X1_130/A POR2X1_558/Y 0.04fF
C60441 POR2X1_7/B POR2X1_260/A 0.04fF
C60442 VDD PAND2X1_156/B 0.07fF
C60443 POR2X1_596/A POR2X1_407/Y 0.03fF
C60444 POR2X1_3/A PAND2X1_711/A 0.03fF
C60445 POR2X1_283/A PAND2X1_190/Y 0.05fF
C60446 POR2X1_68/B PAND2X1_79/Y 0.03fF
C60447 PAND2X1_661/Y POR2X1_43/B 0.03fF
C60448 POR2X1_480/A POR2X1_802/A 0.02fF
C60449 POR2X1_209/A POR2X1_788/B 0.04fF
C60450 POR2X1_346/B POR2X1_785/A 0.03fF
C60451 PAND2X1_84/Y POR2X1_150/CTRL2 0.04fF
C60452 POR2X1_719/CTRL PAND2X1_32/B 0.03fF
C60453 POR2X1_213/O POR2X1_568/Y 0.04fF
C60454 PAND2X1_35/Y POR2X1_394/A 0.03fF
C60455 PAND2X1_63/Y PAND2X1_60/B 0.14fF
C60456 POR2X1_651/Y POR2X1_655/A 0.03fF
C60457 PAND2X1_23/Y POR2X1_332/CTRL2 0.01fF
C60458 POR2X1_773/A VDD 0.04fF
C60459 POR2X1_502/A POR2X1_774/A 0.07fF
C60460 PAND2X1_194/O POR2X1_73/Y 0.05fF
C60461 POR2X1_124/CTRL2 POR2X1_78/A 0.01fF
C60462 POR2X1_190/Y PAND2X1_189/O 0.17fF
C60463 POR2X1_38/B PAND2X1_670/O 0.04fF
C60464 PAND2X1_343/O POR2X1_42/Y 0.03fF
C60465 PAND2X1_585/CTRL PAND2X1_56/A 0.01fF
C60466 POR2X1_218/A POR2X1_276/Y 0.07fF
C60467 POR2X1_447/O POR2X1_510/Y 0.01fF
C60468 PAND2X1_495/O PAND2X1_60/B 0.01fF
C60469 POR2X1_553/Y POR2X1_186/B 0.01fF
C60470 PAND2X1_778/Y POR2X1_387/Y 0.06fF
C60471 PAND2X1_41/B POR2X1_568/B 0.04fF
C60472 PAND2X1_580/B POR2X1_767/O 0.00fF
C60473 POR2X1_664/CTRL2 POR2X1_712/Y 0.03fF
C60474 PAND2X1_460/O POR2X1_380/Y -0.00fF
C60475 PAND2X1_341/B PAND2X1_206/a_16_344# 0.01fF
C60476 PAND2X1_115/B PAND2X1_853/B 2.31fF
C60477 PAND2X1_47/B PAND2X1_72/A 0.08fF
C60478 PAND2X1_555/Y PAND2X1_854/A 1.08fF
C60479 POR2X1_789/A POR2X1_789/B 0.15fF
C60480 PAND2X1_90/A POR2X1_186/B 0.07fF
C60481 POR2X1_278/Y POR2X1_119/Y 0.10fF
C60482 PAND2X1_674/CTRL2 POR2X1_186/B 0.01fF
C60483 POR2X1_347/A POR2X1_68/A 0.01fF
C60484 POR2X1_327/Y POR2X1_861/CTRL2 0.01fF
C60485 PAND2X1_470/O PAND2X1_467/Y 0.01fF
C60486 PAND2X1_726/B PAND2X1_546/O 0.06fF
C60487 PAND2X1_631/A POR2X1_516/B 0.01fF
C60488 PAND2X1_458/m4_208_n4# PAND2X1_785/m4_208_n4# 0.05fF
C60489 POR2X1_783/O PAND2X1_52/B 0.01fF
C60490 POR2X1_717/O POR2X1_101/Y 0.07fF
C60491 POR2X1_315/Y POR2X1_91/Y 0.06fF
C60492 PAND2X1_127/CTRL2 POR2X1_532/A 0.01fF
C60493 POR2X1_184/Y POR2X1_394/A 0.05fF
C60494 POR2X1_569/CTRL2 PAND2X1_52/B 0.04fF
C60495 PAND2X1_513/O POR2X1_77/Y 0.09fF
C60496 POR2X1_462/B POR2X1_753/CTRL 0.03fF
C60497 PAND2X1_701/CTRL2 PAND2X1_69/A 0.00fF
C60498 POR2X1_62/Y PAND2X1_228/O 0.02fF
C60499 POR2X1_713/A POR2X1_711/Y 0.02fF
C60500 POR2X1_100/O PAND2X1_86/Y 0.04fF
C60501 PAND2X1_651/Y POR2X1_394/A 0.10fF
C60502 POR2X1_523/Y POR2X1_523/B 0.04fF
C60503 POR2X1_163/O POR2X1_158/Y 0.00fF
C60504 POR2X1_740/Y POR2X1_188/Y 0.03fF
C60505 PAND2X1_60/B POR2X1_260/A 3.12fF
C60506 POR2X1_554/B POR2X1_446/B 0.02fF
C60507 PAND2X1_661/O POR2X1_761/A 0.02fF
C60508 POR2X1_737/A POR2X1_513/Y 0.03fF
C60509 POR2X1_257/A POR2X1_431/Y 0.04fF
C60510 POR2X1_326/A POR2X1_542/B -0.00fF
C60511 POR2X1_78/B POR2X1_147/CTRL 0.03fF
C60512 POR2X1_773/A PAND2X1_32/B 0.03fF
C60513 POR2X1_68/A POR2X1_4/Y 0.07fF
C60514 PAND2X1_652/O POR2X1_594/Y 0.00fF
C60515 POR2X1_376/A POR2X1_376/a_16_28# 0.05fF
C60516 PAND2X1_30/CTRL2 POR2X1_750/B 0.01fF
C60517 PAND2X1_48/B POR2X1_486/B 0.31fF
C60518 PAND2X1_172/m4_208_n4# POR2X1_854/B 0.04fF
C60519 POR2X1_309/Y PAND2X1_352/Y 0.05fF
C60520 POR2X1_391/Y PAND2X1_134/CTRL 0.03fF
C60521 POR2X1_119/Y INPUT_2 0.01fF
C60522 POR2X1_136/Y POR2X1_129/Y 0.03fF
C60523 PAND2X1_607/O PAND2X1_58/A 0.02fF
C60524 POR2X1_850/CTRL2 POR2X1_737/A 0.01fF
C60525 PAND2X1_90/O POR2X1_38/B 0.21fF
C60526 POR2X1_394/A POR2X1_503/Y 0.05fF
C60527 POR2X1_302/Y POR2X1_717/B 0.02fF
C60528 POR2X1_361/CTRL2 POR2X1_294/A 0.00fF
C60529 POR2X1_361/CTRL PAND2X1_48/A 0.01fF
C60530 POR2X1_101/CTRL POR2X1_334/Y 0.01fF
C60531 POR2X1_416/B POR2X1_293/Y 0.27fF
C60532 POR2X1_54/Y POR2X1_126/CTRL 0.01fF
C60533 POR2X1_278/Y PAND2X1_349/CTRL2 0.00fF
C60534 POR2X1_405/Y PAND2X1_52/B 0.03fF
C60535 POR2X1_537/a_16_28# POR2X1_537/A 0.09fF
C60536 PAND2X1_20/A PAND2X1_85/CTRL 0.00fF
C60537 POR2X1_566/A POR2X1_568/A 0.07fF
C60538 POR2X1_784/A PAND2X1_52/B 0.03fF
C60539 PAND2X1_809/B PAND2X1_794/B 0.03fF
C60540 POR2X1_189/CTRL2 POR2X1_816/A 0.01fF
C60541 POR2X1_616/Y PAND2X1_154/CTRL2 0.01fF
C60542 POR2X1_129/CTRL2 POR2X1_411/B 0.01fF
C60543 PAND2X1_350/O POR2X1_4/Y 0.02fF
C60544 POR2X1_62/Y PAND2X1_100/CTRL2 0.01fF
C60545 PAND2X1_39/B POR2X1_807/CTRL2 0.00fF
C60546 PAND2X1_604/O PAND2X1_72/A 0.05fF
C60547 POR2X1_557/B POR2X1_768/CTRL2 0.00fF
C60548 POR2X1_567/A POR2X1_854/B 0.00fF
C60549 POR2X1_234/A POR2X1_233/O 0.00fF
C60550 POR2X1_77/Y PAND2X1_359/O 0.05fF
C60551 POR2X1_271/A POR2X1_153/Y 0.03fF
C60552 POR2X1_36/O POR2X1_39/B 0.20fF
C60553 POR2X1_7/CTRL POR2X1_7/Y 0.01fF
C60554 POR2X1_814/B PAND2X1_85/CTRL 0.00fF
C60555 POR2X1_461/Y POR2X1_590/A 0.05fF
C60556 POR2X1_271/B POR2X1_516/Y 0.03fF
C60557 PAND2X1_220/Y POR2X1_250/Y 0.63fF
C60558 POR2X1_862/A POR2X1_286/CTRL 0.00fF
C60559 PAND2X1_23/Y POR2X1_863/A 0.03fF
C60560 PAND2X1_48/B POR2X1_76/B 0.03fF
C60561 POR2X1_78/A POR2X1_471/A 0.17fF
C60562 POR2X1_191/Y POR2X1_545/O 0.05fF
C60563 POR2X1_260/B D_INPUT_0 0.13fF
C60564 PAND2X1_407/O POR2X1_29/A 0.02fF
C60565 POR2X1_850/B PAND2X1_39/B 0.04fF
C60566 POR2X1_54/Y PAND2X1_58/A 1.03fF
C60567 POR2X1_119/Y POR2X1_122/CTRL2 0.01fF
C60568 POR2X1_66/B PAND2X1_416/CTRL2 0.01fF
C60569 POR2X1_540/A PAND2X1_72/A 4.84fF
C60570 POR2X1_411/B POR2X1_40/Y 9.33fF
C60571 PAND2X1_827/O POR2X1_294/Y 0.00fF
C60572 PAND2X1_678/O POR2X1_72/B 0.16fF
C60573 POR2X1_416/B POR2X1_408/Y 0.04fF
C60574 POR2X1_122/O PAND2X1_659/Y 0.11fF
C60575 PAND2X1_58/A POR2X1_202/A 0.10fF
C60576 PAND2X1_11/CTRL INPUT_5 0.01fF
C60577 POR2X1_65/A PAND2X1_449/a_76_28# 0.01fF
C60578 POR2X1_848/A POR2X1_753/Y 0.09fF
C60579 POR2X1_796/A POR2X1_711/Y 0.07fF
C60580 POR2X1_479/B POR2X1_66/A 0.02fF
C60581 PAND2X1_237/CTRL2 POR2X1_241/B 0.01fF
C60582 POR2X1_66/A PAND2X1_595/O 0.01fF
C60583 PAND2X1_67/CTRL POR2X1_330/Y 0.03fF
C60584 PAND2X1_173/a_16_344# PAND2X1_72/A 0.02fF
C60585 POR2X1_165/Y PAND2X1_326/B 0.12fF
C60586 PAND2X1_650/A POR2X1_77/Y 0.01fF
C60587 POR2X1_274/CTRL2 POR2X1_296/B 0.03fF
C60588 PAND2X1_65/B POR2X1_541/B 0.00fF
C60589 POR2X1_445/A POR2X1_750/B 0.10fF
C60590 POR2X1_456/B POR2X1_736/A 0.03fF
C60591 POR2X1_357/a_16_28# POR2X1_357/B -0.00fF
C60592 POR2X1_329/A POR2X1_7/B 0.17fF
C60593 PAND2X1_93/B POR2X1_201/CTRL2 0.00fF
C60594 PAND2X1_48/B POR2X1_486/CTRL2 0.03fF
C60595 POR2X1_87/CTRL2 POR2X1_260/A 0.03fF
C60596 POR2X1_210/A POR2X1_330/O 0.01fF
C60597 POR2X1_150/Y POR2X1_481/A 0.03fF
C60598 POR2X1_259/A POR2X1_454/A 0.24fF
C60599 POR2X1_669/B POR2X1_32/A 4.05fF
C60600 PAND2X1_666/O PAND2X1_20/A 0.23fF
C60601 POR2X1_191/a_16_28# POR2X1_191/B 0.03fF
C60602 POR2X1_68/A POR2X1_458/Y 0.10fF
C60603 POR2X1_346/A PAND2X1_58/A 0.00fF
C60604 POR2X1_614/Y POR2X1_590/A 0.02fF
C60605 POR2X1_537/Y POR2X1_840/Y 0.00fF
C60606 POR2X1_102/Y POR2X1_268/O 0.02fF
C60607 POR2X1_859/O PAND2X1_57/B 0.02fF
C60608 POR2X1_691/O POR2X1_814/A 0.02fF
C60609 PAND2X1_217/O INPUT_0 0.02fF
C60610 PAND2X1_633/CTRL2 PAND2X1_640/B 0.03fF
C60611 POR2X1_329/a_16_28# POR2X1_760/A 0.03fF
C60612 POR2X1_260/B PAND2X1_90/Y 0.42fF
C60613 PAND2X1_52/O POR2X1_35/Y 0.02fF
C60614 POR2X1_692/CTRL2 POR2X1_692/Y 0.01fF
C60615 POR2X1_62/Y POR2X1_77/Y 0.03fF
C60616 POR2X1_290/Y POR2X1_20/B 0.14fF
C60617 PAND2X1_477/B POR2X1_329/A 0.02fF
C60618 POR2X1_188/A PAND2X1_282/O 0.02fF
C60619 POR2X1_13/A POR2X1_604/a_56_344# 0.00fF
C60620 POR2X1_102/Y POR2X1_251/CTRL2 0.01fF
C60621 PAND2X1_10/CTRL PAND2X1_41/B 0.03fF
C60622 POR2X1_48/A PAND2X1_712/CTRL2 0.01fF
C60623 PAND2X1_56/Y POR2X1_554/B 0.03fF
C60624 POR2X1_189/Y POR2X1_679/O 0.01fF
C60625 PAND2X1_390/Y POR2X1_29/A 0.85fF
C60626 PAND2X1_231/CTRL POR2X1_32/A 0.01fF
C60627 POR2X1_163/A POR2X1_257/A 0.01fF
C60628 PAND2X1_472/A PAND2X1_608/m4_208_n4# 0.08fF
C60629 POR2X1_288/A POR2X1_590/A 0.03fF
C60630 POR2X1_846/O POR2X1_260/A 0.09fF
C60631 POR2X1_20/B POR2X1_238/Y 0.03fF
C60632 PAND2X1_124/Y INPUT_0 0.01fF
C60633 POR2X1_23/Y PAND2X1_735/CTRL 0.01fF
C60634 POR2X1_20/B PAND2X1_658/B 0.05fF
C60635 PAND2X1_58/A PAND2X1_23/CTRL 0.01fF
C60636 POR2X1_13/A POR2X1_265/O 0.02fF
C60637 POR2X1_23/Y PAND2X1_579/B 0.23fF
C60638 PAND2X1_485/CTRL2 POR2X1_546/A 0.10fF
C60639 POR2X1_832/Y POR2X1_722/Y 0.01fF
C60640 POR2X1_590/A POR2X1_193/Y 0.03fF
C60641 POR2X1_230/O POR2X1_32/A 0.00fF
C60642 PAND2X1_848/B POR2X1_411/B 0.03fF
C60643 POR2X1_257/A PAND2X1_162/CTRL2 0.00fF
C60644 POR2X1_12/A POR2X1_700/CTRL 0.08fF
C60645 POR2X1_66/B POR2X1_777/B 0.03fF
C60646 POR2X1_409/B VDD 0.03fF
C60647 PAND2X1_793/Y PAND2X1_287/Y 3.06fF
C60648 POR2X1_454/A POR2X1_231/B 0.03fF
C60649 POR2X1_65/A POR2X1_14/Y 0.08fF
C60650 POR2X1_814/A POR2X1_162/Y 0.08fF
C60651 POR2X1_49/Y PAND2X1_476/CTRL2 0.00fF
C60652 POR2X1_567/B PAND2X1_524/CTRL2 0.49fF
C60653 POR2X1_66/A POR2X1_194/B 0.01fF
C60654 PAND2X1_20/A POR2X1_231/A 0.01fF
C60655 POR2X1_105/CTRL POR2X1_814/B 0.01fF
C60656 POR2X1_66/B POR2X1_194/A 0.23fF
C60657 PAND2X1_267/CTRL PAND2X1_215/B 0.03fF
C60658 POR2X1_779/A PAND2X1_39/B 0.03fF
C60659 PAND2X1_9/Y POR2X1_409/CTRL2 0.01fF
C60660 PAND2X1_65/B POR2X1_390/O 0.04fF
C60661 POR2X1_862/A POR2X1_294/B 0.03fF
C60662 POR2X1_188/A POR2X1_777/B 0.05fF
C60663 PAND2X1_23/Y POR2X1_274/A 0.08fF
C60664 PAND2X1_437/CTRL2 POR2X1_186/B 0.01fF
C60665 PAND2X1_217/B PAND2X1_659/A 0.01fF
C60666 POR2X1_389/O POR2X1_260/B 0.02fF
C60667 POR2X1_23/Y POR2X1_763/Y 0.14fF
C60668 POR2X1_66/B PAND2X1_65/B 0.16fF
C60669 PAND2X1_114/Y POR2X1_48/A 0.01fF
C60670 POR2X1_188/A POR2X1_660/A 0.03fF
C60671 POR2X1_466/A PAND2X1_183/O 0.15fF
C60672 POR2X1_376/B POR2X1_40/Y 2.94fF
C60673 POR2X1_45/Y PAND2X1_267/Y 0.03fF
C60674 POR2X1_590/A POR2X1_723/a_56_344# 0.00fF
C60675 PAND2X1_808/Y PAND2X1_773/Y 1.27fF
C60676 POR2X1_96/A PAND2X1_223/B 0.03fF
C60677 POR2X1_83/B INPUT_0 5.18fF
C60678 POR2X1_669/B PAND2X1_35/Y 0.03fF
C60679 POR2X1_383/A POR2X1_554/B 0.01fF
C60680 POR2X1_20/B POR2X1_299/a_76_344# 0.01fF
C60681 POR2X1_54/Y PAND2X1_96/B 0.03fF
C60682 PAND2X1_209/A PAND2X1_213/CTRL 0.01fF
C60683 PAND2X1_809/a_76_28# PAND2X1_539/Y 0.05fF
C60684 POR2X1_486/O POR2X1_260/A 0.01fF
C60685 POR2X1_188/A PAND2X1_65/B 0.03fF
C60686 POR2X1_16/A POR2X1_600/CTRL 0.01fF
C60687 PAND2X1_658/A POR2X1_23/Y 0.03fF
C60688 PAND2X1_655/O PAND2X1_655/B 0.07fF
C60689 POR2X1_814/A POR2X1_734/O 0.01fF
C60690 PAND2X1_55/Y D_INPUT_0 1.63fF
C60691 PAND2X1_786/O PAND2X1_84/Y 0.02fF
C60692 POR2X1_24/Y POR2X1_38/Y 0.03fF
C60693 PAND2X1_40/CTRL PAND2X1_59/B 0.01fF
C60694 POR2X1_44/O INPUT_7 0.16fF
C60695 POR2X1_49/Y PAND2X1_596/CTRL 0.01fF
C60696 POR2X1_646/CTRL POR2X1_121/B 0.20fF
C60697 POR2X1_568/A POR2X1_568/CTRL2 0.01fF
C60698 PAND2X1_826/a_16_344# PAND2X1_96/B 0.02fF
C60699 PAND2X1_96/B POR2X1_202/A 0.00fF
C60700 POR2X1_643/O POR2X1_294/A 0.50fF
C60701 POR2X1_341/A POR2X1_228/Y 0.10fF
C60702 PAND2X1_217/B POR2X1_272/Y 0.09fF
C60703 PAND2X1_84/Y POR2X1_72/B 0.02fF
C60704 PAND2X1_90/A PAND2X1_245/CTRL2 0.03fF
C60705 PAND2X1_391/O POR2X1_42/Y 0.09fF
C60706 POR2X1_865/CTRL POR2X1_260/B 0.00fF
C60707 PAND2X1_73/Y POR2X1_294/B 0.37fF
C60708 POR2X1_674/Y PAND2X1_592/Y 0.03fF
C60709 PAND2X1_791/O POR2X1_755/Y 0.01fF
C60710 POR2X1_454/A PAND2X1_88/Y 0.02fF
C60711 POR2X1_376/B PAND2X1_185/a_76_28# 0.03fF
C60712 POR2X1_607/A POR2X1_411/O 0.00fF
C60713 PAND2X1_247/a_56_28# POR2X1_7/A 0.00fF
C60714 POR2X1_509/A POR2X1_97/A 0.01fF
C60715 POR2X1_821/Y PAND2X1_852/A 0.03fF
C60716 POR2X1_499/CTRL POR2X1_576/Y 0.02fF
C60717 POR2X1_52/A PAND2X1_512/CTRL2 0.03fF
C60718 PAND2X1_863/B POR2X1_595/a_16_28# 0.02fF
C60719 POR2X1_814/B PAND2X1_236/O 0.06fF
C60720 POR2X1_63/CTRL POR2X1_669/B 0.01fF
C60721 PAND2X1_6/Y POR2X1_466/A 1.91fF
C60722 POR2X1_23/Y POR2X1_73/Y 1.11fF
C60723 POR2X1_72/B POR2X1_531/CTRL2 0.01fF
C60724 POR2X1_422/CTRL POR2X1_93/A 0.00fF
C60725 PAND2X1_39/B POR2X1_598/CTRL2 0.02fF
C60726 D_INPUT_3 POR2X1_612/B 0.01fF
C60727 PAND2X1_216/B POR2X1_150/Y 0.06fF
C60728 POR2X1_863/A POR2X1_711/Y 0.07fF
C60729 POR2X1_218/Y D_INPUT_1 0.07fF
C60730 POR2X1_52/A POR2X1_40/Y 1.98fF
C60731 POR2X1_41/B PAND2X1_842/CTRL2 0.03fF
C60732 POR2X1_57/A PAND2X1_640/B 0.03fF
C60733 POR2X1_270/CTRL2 POR2X1_66/A 0.09fF
C60734 POR2X1_264/CTRL POR2X1_294/B 0.05fF
C60735 POR2X1_264/Y POR2X1_264/CTRL2 0.01fF
C60736 PAND2X1_554/a_56_28# POR2X1_7/B 0.00fF
C60737 D_INPUT_0 POR2X1_407/Y 0.03fF
C60738 POR2X1_760/A POR2X1_594/CTRL2 0.03fF
C60739 PAND2X1_89/CTRL2 POR2X1_61/Y 0.03fF
C60740 PAND2X1_651/Y POR2X1_669/B 0.03fF
C60741 POR2X1_346/A PAND2X1_96/B 0.00fF
C60742 POR2X1_558/a_16_28# POR2X1_590/A 0.01fF
C60743 POR2X1_278/Y PAND2X1_204/CTRL2 0.05fF
C60744 POR2X1_709/A PAND2X1_748/O 0.11fF
C60745 POR2X1_102/Y PAND2X1_794/B 0.03fF
C60746 POR2X1_60/A POR2X1_289/CTRL 0.01fF
C60747 PAND2X1_65/B POR2X1_859/A 0.07fF
C60748 D_INPUT_0 POR2X1_783/Y 0.00fF
C60749 POR2X1_272/Y VDD 0.14fF
C60750 POR2X1_40/Y POR2X1_152/A 0.03fF
C60751 POR2X1_567/B POR2X1_714/O 0.02fF
C60752 POR2X1_218/Y POR2X1_724/A 0.08fF
C60753 PAND2X1_47/CTRL2 PAND2X1_11/Y 0.04fF
C60754 POR2X1_763/Y POR2X1_764/Y 0.03fF
C60755 POR2X1_625/Y POR2X1_5/Y 0.03fF
C60756 PAND2X1_738/Y PAND2X1_544/CTRL 0.32fF
C60757 POR2X1_811/A POR2X1_783/Y 0.00fF
C60758 INPUT_1 POR2X1_24/Y 0.04fF
C60759 PAND2X1_408/Y PAND2X1_11/Y 0.12fF
C60760 POR2X1_43/B PAND2X1_639/CTRL2 0.03fF
C60761 POR2X1_781/O VDD 0.00fF
C60762 PAND2X1_620/Y POR2X1_55/Y 0.03fF
C60763 POR2X1_102/Y PAND2X1_723/O 0.02fF
C60764 POR2X1_66/A POR2X1_537/B 0.01fF
C60765 POR2X1_57/A POR2X1_666/CTRL 0.01fF
C60766 POR2X1_69/A PAND2X1_6/A 0.02fF
C60767 POR2X1_646/O PAND2X1_90/Y 0.02fF
C60768 POR2X1_65/A POR2X1_55/Y 0.14fF
C60769 POR2X1_135/Y POR2X1_46/Y 1.08fF
C60770 PAND2X1_280/a_16_344# PAND2X1_90/Y 0.07fF
C60771 PAND2X1_11/Y PAND2X1_26/CTRL 0.03fF
C60772 PAND2X1_65/B POR2X1_828/CTRL 0.01fF
C60773 D_GATE_222 POR2X1_355/A 0.02fF
C60774 POR2X1_23/Y PAND2X1_244/B 0.04fF
C60775 PAND2X1_795/B INPUT_0 0.03fF
C60776 POR2X1_814/B PAND2X1_385/O 0.01fF
C60777 PAND2X1_74/CTRL2 PAND2X1_32/B 0.01fF
C60778 PAND2X1_48/Y PAND2X1_23/Y 0.02fF
C60779 PAND2X1_845/a_16_344# POR2X1_60/A 0.00fF
C60780 POR2X1_399/CTRL POR2X1_293/Y 0.01fF
C60781 VDD PAND2X1_351/Y 0.11fF
C60782 PAND2X1_444/Y POR2X1_90/Y 0.03fF
C60783 PAND2X1_340/O POR2X1_42/Y 0.02fF
C60784 POR2X1_71/Y POR2X1_497/Y 0.16fF
C60785 D_INPUT_2 POR2X1_611/O 0.01fF
C60786 PAND2X1_73/Y PAND2X1_111/B 0.15fF
C60787 INPUT_7 POR2X1_587/CTRL 0.01fF
C60788 POR2X1_423/Y POR2X1_56/Y 0.14fF
C60789 PAND2X1_55/Y PAND2X1_90/Y 0.17fF
C60790 POR2X1_302/B POR2X1_513/Y 0.03fF
C60791 POR2X1_416/B PAND2X1_405/CTRL 0.01fF
C60792 POR2X1_590/A PAND2X1_670/O 0.00fF
C60793 PAND2X1_423/m4_208_n4# PAND2X1_56/m4_208_n4# 0.13fF
C60794 PAND2X1_423/a_56_28# PAND2X1_55/Y 0.00fF
C60795 POR2X1_465/B VDD 0.00fF
C60796 POR2X1_68/A PAND2X1_52/Y 0.01fF
C60797 D_INPUT_0 PAND2X1_28/O 0.03fF
C60798 POR2X1_848/A POR2X1_754/O 0.02fF
C60799 PAND2X1_512/Y POR2X1_293/Y 0.07fF
C60800 POR2X1_72/B POR2X1_594/A 0.01fF
C60801 POR2X1_121/O POR2X1_121/B 0.02fF
C60802 POR2X1_266/A POR2X1_624/Y 0.03fF
C60803 POR2X1_707/B INPUT_6 0.01fF
C60804 PAND2X1_848/B POR2X1_376/B 0.02fF
C60805 POR2X1_496/Y PAND2X1_748/CTRL2 0.11fF
C60806 PAND2X1_41/B PAND2X1_767/O 0.01fF
C60807 POR2X1_16/A POR2X1_263/Y 0.03fF
C60808 PAND2X1_308/B POR2X1_56/B 0.07fF
C60809 POR2X1_490/Y PAND2X1_560/B 0.03fF
C60810 PAND2X1_460/CTRL POR2X1_94/A 0.01fF
C60811 POR2X1_198/B VDD 0.16fF
C60812 POR2X1_651/CTRL PAND2X1_386/Y 0.01fF
C60813 POR2X1_25/Y D_INPUT_5 0.03fF
C60814 POR2X1_539/CTRL2 POR2X1_590/A 0.03fF
C60815 PAND2X1_480/B PAND2X1_303/CTRL 0.30fF
C60816 POR2X1_764/Y POR2X1_73/Y 0.01fF
C60817 PAND2X1_42/CTRL POR2X1_38/B 0.05fF
C60818 POR2X1_844/O POR2X1_94/A 0.02fF
C60819 POR2X1_65/A POR2X1_166/CTRL2 0.03fF
C60820 PAND2X1_783/Y POR2X1_90/Y 0.03fF
C60821 VDD POR2X1_501/CTRL 0.00fF
C60822 PAND2X1_425/CTRL INPUT_6 0.01fF
C60823 POR2X1_41/B POR2X1_597/A 0.08fF
C60824 PAND2X1_526/O PAND2X1_32/B 0.15fF
C60825 POR2X1_687/Y POR2X1_800/O 0.00fF
C60826 POR2X1_680/Y POR2X1_79/Y 0.04fF
C60827 POR2X1_323/CTRL POR2X1_73/Y 0.01fF
C60828 POR2X1_686/A POR2X1_596/A 0.02fF
C60829 POR2X1_78/A POR2X1_116/Y 0.05fF
C60830 PAND2X1_449/Y POR2X1_236/Y 0.01fF
C60831 D_GATE_741 VDD -0.00fF
C60832 PAND2X1_20/A PAND2X1_297/CTRL2 0.00fF
C60833 POR2X1_708/CTRL2 POR2X1_407/A 0.00fF
C60834 POR2X1_748/A POR2X1_245/a_76_344# 0.00fF
C60835 POR2X1_49/Y D_INPUT_3 0.05fF
C60836 PAND2X1_65/B POR2X1_705/a_56_344# 0.00fF
C60837 POR2X1_346/B PAND2X1_39/CTRL 0.00fF
C60838 PAND2X1_810/A GATE_811 0.12fF
C60839 POR2X1_311/Y PAND2X1_336/CTRL2 0.01fF
C60840 POR2X1_41/B POR2X1_48/Y 1.68fF
C60841 POR2X1_730/Y POR2X1_78/A 0.03fF
C60842 POR2X1_437/CTRL POR2X1_385/Y 0.13fF
C60843 POR2X1_407/Y PAND2X1_90/Y 0.04fF
C60844 POR2X1_126/CTRL POR2X1_4/Y 0.01fF
C60845 POR2X1_855/B POR2X1_330/Y 0.05fF
C60846 POR2X1_614/A POR2X1_284/B 0.03fF
C60847 PAND2X1_20/A POR2X1_664/CTRL2 0.00fF
C60848 PAND2X1_65/B PAND2X1_59/O 0.03fF
C60849 POR2X1_128/O POR2X1_222/Y 0.05fF
C60850 PAND2X1_58/A PAND2X1_748/O 0.32fF
C60851 POR2X1_326/A POR2X1_856/B 0.03fF
C60852 PAND2X1_839/CTRL POR2X1_293/Y 0.01fF
C60853 POR2X1_41/B PAND2X1_652/A 7.24fF
C60854 POR2X1_685/A POR2X1_750/B 1.92fF
C60855 POR2X1_93/O VDD 0.00fF
C60856 PAND2X1_498/O POR2X1_733/A 0.04fF
C60857 POR2X1_718/A PAND2X1_60/B 0.06fF
C60858 POR2X1_101/CTRL2 POR2X1_814/B 0.01fF
C60859 PAND2X1_562/B PAND2X1_348/Y 0.01fF
C60860 POR2X1_502/A POR2X1_459/B 0.01fF
C60861 PAND2X1_88/CTRL2 POR2X1_260/A 0.03fF
C60862 PAND2X1_441/a_76_28# PAND2X1_52/B 0.02fF
C60863 POR2X1_591/Y POR2X1_236/Y 0.07fF
C60864 POR2X1_347/A PAND2X1_58/A 0.01fF
C60865 VDD POR2X1_685/B 0.00fF
C60866 POR2X1_66/A PAND2X1_48/A 0.51fF
C60867 POR2X1_22/A POR2X1_22/a_76_344# 0.00fF
C60868 POR2X1_294/B PAND2X1_144/CTRL 0.03fF
C60869 POR2X1_779/A POR2X1_513/B 0.01fF
C60870 POR2X1_46/Y POR2X1_816/A 0.03fF
C60871 POR2X1_311/Y PAND2X1_182/B 0.05fF
C60872 POR2X1_502/A POR2X1_638/Y 0.03fF
C60873 POR2X1_34/B POR2X1_294/A 0.01fF
C60874 POR2X1_844/CTRL2 POR2X1_546/A 0.01fF
C60875 PAND2X1_696/CTRL PAND2X1_93/B 0.03fF
C60876 POR2X1_686/B POR2X1_686/O 0.01fF
C60877 PAND2X1_38/CTRL POR2X1_68/B 0.02fF
C60878 POR2X1_582/CTRL2 INPUT_4 0.10fF
C60879 POR2X1_750/B POR2X1_260/A 0.14fF
C60880 PAND2X1_793/Y PAND2X1_575/CTRL2 0.01fF
C60881 PAND2X1_499/Y PAND2X1_349/A 0.03fF
C60882 POR2X1_230/Y POR2X1_38/Y 0.05fF
C60883 POR2X1_356/A PAND2X1_69/A 0.05fF
C60884 PAND2X1_209/A PAND2X1_213/B 0.57fF
C60885 POR2X1_465/B PAND2X1_32/B 0.37fF
C60886 POR2X1_68/A D_GATE_662 0.07fF
C60887 POR2X1_740/Y POR2X1_731/CTRL2 0.00fF
C60888 PAND2X1_689/CTRL2 POR2X1_691/A 0.01fF
C60889 PAND2X1_90/A PAND2X1_110/m4_208_n4# 0.07fF
C60890 POR2X1_505/Y PAND2X1_507/CTRL 0.00fF
C60891 PAND2X1_6/Y POR2X1_691/CTRL2 0.00fF
C60892 POR2X1_101/Y POR2X1_573/O 0.02fF
C60893 POR2X1_8/Y PAND2X1_859/A 0.03fF
C60894 POR2X1_294/B POR2X1_631/B 10.58fF
C60895 POR2X1_52/Y PAND2X1_197/Y 0.03fF
C60896 POR2X1_367/O POR2X1_568/Y 0.04fF
C60897 POR2X1_57/A PAND2X1_830/Y 1.40fF
C60898 POR2X1_754/A POR2X1_93/A 0.03fF
C60899 POR2X1_532/A POR2X1_776/B 0.03fF
C60900 D_INPUT_6 INPUT_5 0.07fF
C60901 PAND2X1_90/O POR2X1_590/A 0.04fF
C60902 POR2X1_858/B POR2X1_850/A 0.01fF
C60903 POR2X1_41/B POR2X1_152/Y 0.04fF
C60904 POR2X1_360/A PAND2X1_88/Y 2.23fF
C60905 PAND2X1_290/O POR2X1_84/A 0.02fF
C60906 POR2X1_94/A POR2X1_394/A 0.07fF
C60907 POR2X1_57/A POR2X1_7/B 0.13fF
C60908 POR2X1_125/Y POR2X1_127/Y 0.18fF
C60909 POR2X1_13/A PAND2X1_348/Y 0.57fF
C60910 POR2X1_567/A PAND2X1_73/Y 0.05fF
C60911 POR2X1_234/A POR2X1_411/A 0.01fF
C60912 POR2X1_88/Y POR2X1_7/A 0.04fF
C60913 POR2X1_558/CTRL PAND2X1_32/B 0.01fF
C60914 POR2X1_738/Y POR2X1_319/Y 0.01fF
C60915 PAND2X1_90/A PAND2X1_79/Y 0.03fF
C60916 POR2X1_102/a_16_28# POR2X1_48/A 0.01fF
C60917 PAND2X1_20/A PAND2X1_692/O 0.04fF
C60918 PAND2X1_6/Y POR2X1_149/B 0.03fF
C60919 POR2X1_575/B POR2X1_500/Y 0.12fF
C60920 PAND2X1_649/A POR2X1_32/A 0.00fF
C60921 PAND2X1_73/Y PAND2X1_323/O 0.04fF
C60922 POR2X1_501/CTRL PAND2X1_32/B 0.03fF
C60923 POR2X1_327/Y PAND2X1_299/CTRL 0.01fF
C60924 PAND2X1_56/Y POR2X1_702/A 0.04fF
C60925 PAND2X1_682/O POR2X1_614/A 0.15fF
C60926 POR2X1_502/A POR2X1_169/Y 0.00fF
C60927 POR2X1_247/a_16_28# POR2X1_532/A 0.02fF
C60928 POR2X1_806/a_16_28# POR2X1_737/A 0.02fF
C60929 POR2X1_68/A D_INPUT_1 0.13fF
C60930 PAND2X1_58/A POR2X1_4/Y 0.07fF
C60931 POR2X1_823/Y POR2X1_293/Y 0.00fF
C60932 INPUT_6 POR2X1_408/O 0.00fF
C60933 PAND2X1_551/Y POR2X1_73/Y 0.03fF
C60934 PAND2X1_148/Y PAND2X1_209/A 0.01fF
C60935 PAND2X1_48/B POR2X1_215/Y 0.04fF
C60936 PAND2X1_594/CTRL2 POR2X1_711/Y 0.03fF
C60937 POR2X1_407/CTRL POR2X1_513/B 0.23fF
C60938 PAND2X1_6/Y POR2X1_644/A 0.03fF
C60939 POR2X1_740/Y POR2X1_510/Y 0.02fF
C60940 POR2X1_38/B POR2X1_380/O 0.01fF
C60941 POR2X1_260/B POR2X1_715/O 0.01fF
C60942 POR2X1_417/Y PAND2X1_353/Y 0.03fF
C60943 POR2X1_463/Y PAND2X1_57/B 5.87fF
C60944 PAND2X1_491/O PAND2X1_32/B 0.06fF
C60945 PAND2X1_632/B POR2X1_252/O 0.02fF
C60946 POR2X1_49/Y POR2X1_83/Y 0.02fF
C60947 PAND2X1_32/B POR2X1_685/B 0.01fF
C60948 POR2X1_99/B POR2X1_259/A 0.00fF
C60949 POR2X1_383/A POR2X1_205/CTRL 0.06fF
C60950 POR2X1_268/a_16_28# POR2X1_39/B 0.01fF
C60951 PAND2X1_57/B POR2X1_756/Y 0.01fF
C60952 POR2X1_94/a_16_28# POR2X1_38/Y 0.02fF
C60953 PAND2X1_865/Y PAND2X1_579/CTRL2 0.00fF
C60954 PAND2X1_363/O POR2X1_42/Y 0.05fF
C60955 POR2X1_370/a_16_28# POR2X1_543/A 0.05fF
C60956 PAND2X1_703/CTRL2 POR2X1_236/Y 0.01fF
C60957 POR2X1_840/B POR2X1_573/A 0.03fF
C60958 POR2X1_544/A POR2X1_544/B 0.01fF
C60959 PAND2X1_216/B PAND2X1_364/B 0.01fF
C60960 POR2X1_860/CTRL2 POR2X1_572/B 0.01fF
C60961 POR2X1_16/A PAND2X1_215/B 0.10fF
C60962 POR2X1_158/Y POR2X1_163/Y 0.04fF
C60963 POR2X1_51/A POR2X1_394/A 0.03fF
C60964 PAND2X1_709/a_16_344# POR2X1_158/B 0.00fF
C60965 PAND2X1_373/a_16_344# POR2X1_732/B 0.09fF
C60966 POR2X1_111/Y POR2X1_7/B 0.02fF
C60967 POR2X1_38/Y POR2X1_619/Y 0.44fF
C60968 POR2X1_356/A PAND2X1_824/B 1.68fF
C60969 PAND2X1_140/A POR2X1_90/Y 0.03fF
C60970 POR2X1_334/B PAND2X1_184/CTRL2 0.31fF
C60971 POR2X1_482/Y POR2X1_39/B 0.02fF
C60972 PAND2X1_308/O POR2X1_56/B 0.06fF
C60973 POR2X1_199/a_16_28# POR2X1_260/A 0.01fF
C60974 POR2X1_416/B POR2X1_60/A 2.84fF
C60975 POR2X1_327/Y POR2X1_327/CTRL 0.01fF
C60976 POR2X1_383/A POR2X1_702/A 2.23fF
C60977 PAND2X1_94/A POR2X1_43/B 0.03fF
C60978 POR2X1_528/Y POR2X1_90/Y 0.22fF
C60979 POR2X1_98/A PAND2X1_39/B 0.03fF
C60980 PAND2X1_319/B PAND2X1_803/Y 0.02fF
C60981 POR2X1_846/A POR2X1_496/O 0.18fF
C60982 POR2X1_785/A POR2X1_507/A 0.07fF
C60983 POR2X1_309/Y POR2X1_310/Y 0.01fF
C60984 POR2X1_550/CTRL POR2X1_550/Y 0.01fF
C60985 PAND2X1_382/a_16_344# PAND2X1_69/A 0.02fF
C60986 PAND2X1_846/CTRL POR2X1_750/A 0.06fF
C60987 PAND2X1_90/Y POR2X1_741/O 0.02fF
C60988 POR2X1_315/Y POR2X1_299/CTRL 0.01fF
C60989 POR2X1_614/A PAND2X1_94/A 0.07fF
C60990 POR2X1_16/A PAND2X1_6/A 0.10fF
C60991 POR2X1_122/O POR2X1_293/Y 0.16fF
C60992 POR2X1_717/m4_208_n4# POR2X1_114/m4_208_n4# 0.13fF
C60993 POR2X1_241/B POR2X1_568/A 0.03fF
C60994 PAND2X1_751/CTRL POR2X1_294/A 0.01fF
C60995 POR2X1_96/A POR2X1_385/Y 0.05fF
C60996 POR2X1_542/B POR2X1_787/CTRL 0.01fF
C60997 PAND2X1_108/CTRL POR2X1_862/B 0.00fF
C60998 POR2X1_110/CTRL POR2X1_372/Y 0.06fF
C60999 PAND2X1_20/A POR2X1_768/A 0.00fF
C61000 POR2X1_717/CTRL2 POR2X1_390/B 0.00fF
C61001 POR2X1_276/A POR2X1_140/a_16_28# 0.07fF
C61002 PAND2X1_476/A POR2X1_13/A 0.02fF
C61003 PAND2X1_94/A POR2X1_38/B 0.10fF
C61004 INPUT_3 PAND2X1_87/a_76_28# 0.05fF
C61005 PAND2X1_504/O POR2X1_507/A 0.05fF
C61006 POR2X1_725/Y PAND2X1_60/B 0.26fF
C61007 POR2X1_234/A POR2X1_32/A 0.12fF
C61008 POR2X1_845/CTRL POR2X1_7/A 0.01fF
C61009 POR2X1_617/Y POR2X1_617/O 0.01fF
C61010 POR2X1_680/Y PAND2X1_730/A 0.07fF
C61011 PAND2X1_333/O POR2X1_77/Y 0.06fF
C61012 POR2X1_327/Y POR2X1_218/A 0.57fF
C61013 POR2X1_866/A POR2X1_655/a_16_28# 0.03fF
C61014 POR2X1_750/B PAND2X1_681/O 0.02fF
C61015 PAND2X1_569/B PAND2X1_168/CTRL 0.01fF
C61016 POR2X1_3/B POR2X1_587/Y 0.03fF
C61017 POR2X1_686/CTRL2 POR2X1_260/A 0.01fF
C61018 POR2X1_347/A PAND2X1_96/B 0.01fF
C61019 PAND2X1_360/Y PAND2X1_357/Y 0.03fF
C61020 POR2X1_119/Y PAND2X1_462/B 0.01fF
C61021 POR2X1_627/a_16_28# POR2X1_39/B 0.03fF
C61022 POR2X1_119/Y PAND2X1_478/CTRL2 0.00fF
C61023 POR2X1_294/Y POR2X1_837/A 0.03fF
C61024 POR2X1_711/B POR2X1_805/A 0.03fF
C61025 PAND2X1_632/B POR2X1_245/Y 0.03fF
C61026 INPUT_0 PAND2X1_841/Y 0.02fF
C61027 POR2X1_361/a_16_28# POR2X1_276/Y 0.02fF
C61028 PAND2X1_717/A PAND2X1_205/A 0.03fF
C61029 POR2X1_62/Y POR2X1_52/Y 0.01fF
C61030 POR2X1_130/A PAND2X1_56/A 0.19fF
C61031 POR2X1_68/B PAND2X1_527/CTRL2 0.00fF
C61032 POR2X1_8/Y POR2X1_7/A 0.62fF
C61033 POR2X1_322/Y POR2X1_165/Y 0.02fF
C61034 POR2X1_614/A PAND2X1_680/CTRL2 0.00fF
C61035 POR2X1_725/Y POR2X1_353/A 0.17fF
C61036 PAND2X1_659/Y PAND2X1_473/CTRL2 0.11fF
C61037 POR2X1_101/Y POR2X1_456/B 0.05fF
C61038 POR2X1_16/A POR2X1_280/Y 0.13fF
C61039 POR2X1_532/A PAND2X1_48/A 0.10fF
C61040 PAND2X1_20/A POR2X1_98/A 0.02fF
C61041 POR2X1_532/A POR2X1_192/B 0.05fF
C61042 PAND2X1_35/Y PAND2X1_327/O 0.02fF
C61043 POR2X1_458/Y PAND2X1_58/A 0.26fF
C61044 POR2X1_313/Y PAND2X1_317/CTRL2 0.01fF
C61045 PAND2X1_771/O PAND2X1_771/Y 0.02fF
C61046 PAND2X1_809/A POR2X1_416/B 0.12fF
C61047 POR2X1_263/CTRL2 POR2X1_37/Y 0.01fF
C61048 POR2X1_283/A PAND2X1_508/Y 0.03fF
C61049 POR2X1_566/B POR2X1_580/m4_208_n4# 0.08fF
C61050 POR2X1_760/A PAND2X1_223/B 0.03fF
C61051 POR2X1_540/Y POR2X1_318/A 0.02fF
C61052 PAND2X1_651/O POR2X1_260/A 0.08fF
C61053 PAND2X1_155/O POR2X1_153/Y 0.00fF
C61054 PAND2X1_358/A PAND2X1_100/CTRL 0.04fF
C61055 POR2X1_463/Y PAND2X1_701/O 0.07fF
C61056 POR2X1_703/Y POR2X1_704/Y 0.03fF
C61057 POR2X1_66/B POR2X1_814/A 0.14fF
C61058 POR2X1_66/B PAND2X1_75/CTRL 0.01fF
C61059 POR2X1_537/Y POR2X1_537/A 0.01fF
C61060 POR2X1_539/A POR2X1_537/Y 0.05fF
C61061 POR2X1_461/Y POR2X1_66/A 0.51fF
C61062 PAND2X1_474/O POR2X1_37/Y 0.03fF
C61063 POR2X1_691/CTRL2 PAND2X1_52/B 0.03fF
C61064 PAND2X1_9/Y POR2X1_409/B 0.01fF
C61065 D_INPUT_1 PAND2X1_529/CTRL 0.01fF
C61066 POR2X1_441/O POR2X1_40/Y 0.01fF
C61067 POR2X1_188/A POR2X1_814/A 0.05fF
C61068 PAND2X1_838/B POR2X1_37/Y 0.11fF
C61069 POR2X1_813/CTRL2 POR2X1_669/B 0.01fF
C61070 POR2X1_556/A POR2X1_296/B 0.08fF
C61071 POR2X1_343/Y POR2X1_786/Y 0.10fF
C61072 POR2X1_333/O POR2X1_192/B 0.07fF
C61073 POR2X1_333/CTRL POR2X1_191/Y 0.11fF
C61074 POR2X1_317/a_16_28# PAND2X1_52/B 0.01fF
C61075 POR2X1_130/A POR2X1_661/A 0.10fF
C61076 PAND2X1_348/A PAND2X1_853/B 0.07fF
C61077 PAND2X1_126/a_76_28# POR2X1_62/Y 0.01fF
C61078 PAND2X1_23/Y PAND2X1_96/O 0.00fF
C61079 POR2X1_66/B POR2X1_846/Y 0.03fF
C61080 POR2X1_8/Y POR2X1_384/Y 0.01fF
C61081 POR2X1_593/O POR2X1_449/A 0.01fF
C61082 POR2X1_38/Y PAND2X1_379/m4_208_n4# 0.12fF
C61083 POR2X1_559/Y PAND2X1_52/B 0.01fF
C61084 POR2X1_78/B PAND2X1_607/CTRL2 0.03fF
C61085 POR2X1_383/A PAND2X1_759/O 0.02fF
C61086 PAND2X1_123/a_76_28# POR2X1_117/Y 0.01fF
C61087 POR2X1_119/Y POR2X1_16/A 0.37fF
C61088 PAND2X1_323/CTRL2 POR2X1_456/B 0.01fF
C61089 POR2X1_458/Y POR2X1_457/B 0.04fF
C61090 POR2X1_820/Y POR2X1_9/Y 0.11fF
C61091 PAND2X1_535/CTRL2 POR2X1_533/Y 0.00fF
C61092 PAND2X1_438/CTRL POR2X1_192/Y 0.15fF
C61093 POR2X1_649/CTRL PAND2X1_52/B 0.01fF
C61094 PAND2X1_33/CTRL2 POR2X1_94/A 0.01fF
C61095 PAND2X1_69/A PAND2X1_72/A 0.13fF
C61096 POR2X1_644/A PAND2X1_52/B 0.03fF
C61097 PAND2X1_349/A POR2X1_39/B 0.10fF
C61098 POR2X1_298/CTRL2 POR2X1_32/A 0.01fF
C61099 PAND2X1_63/B POR2X1_39/B 0.05fF
C61100 PAND2X1_93/B POR2X1_218/Y 0.07fF
C61101 POR2X1_112/Y PAND2X1_135/CTRL2 0.00fF
C61102 POR2X1_4/O POR2X1_4/Y 0.01fF
C61103 PAND2X1_85/CTRL VDD -0.00fF
C61104 POR2X1_83/B PAND2X1_340/B 0.01fF
C61105 POR2X1_16/A POR2X1_85/CTRL 0.11fF
C61106 PAND2X1_61/Y POR2X1_262/Y 0.03fF
C61107 PAND2X1_207/O POR2X1_32/A 0.04fF
C61108 POR2X1_502/A POR2X1_463/O 0.01fF
C61109 PAND2X1_600/CTRL2 PAND2X1_20/A 0.00fF
C61110 POR2X1_102/Y PAND2X1_124/Y 0.06fF
C61111 POR2X1_624/B PAND2X1_8/Y 0.21fF
C61112 POR2X1_634/CTRL POR2X1_260/B 0.01fF
C61113 POR2X1_257/A PAND2X1_541/O 0.03fF
C61114 POR2X1_634/A POR2X1_610/O 0.00fF
C61115 POR2X1_866/A POR2X1_866/O 0.10fF
C61116 POR2X1_411/B POR2X1_5/Y 0.16fF
C61117 POR2X1_417/Y POR2X1_298/CTRL2 0.01fF
C61118 POR2X1_862/A POR2X1_643/A 0.02fF
C61119 POR2X1_558/B POR2X1_474/CTRL2 0.02fF
C61120 POR2X1_78/B PAND2X1_418/m4_208_n4# 0.06fF
C61121 POR2X1_29/CTRL2 PAND2X1_9/Y 0.01fF
C61122 POR2X1_78/A POR2X1_218/Y 0.01fF
C61123 POR2X1_846/Y POR2X1_859/A 0.07fF
C61124 POR2X1_852/CTRL2 POR2X1_776/A 0.03fF
C61125 PAND2X1_580/a_76_28# PAND2X1_580/B 0.04fF
C61126 POR2X1_48/A POR2X1_482/Y 1.80fF
C61127 POR2X1_78/B POR2X1_663/B 0.04fF
C61128 POR2X1_96/A POR2X1_679/CTRL 0.01fF
C61129 PAND2X1_639/a_76_28# POR2X1_408/Y 0.05fF
C61130 POR2X1_475/CTRL VDD 0.00fF
C61131 POR2X1_62/Y PAND2X1_358/CTRL2 0.01fF
C61132 PAND2X1_318/a_16_344# PAND2X1_464/B 0.02fF
C61133 POR2X1_848/A POR2X1_615/CTRL -0.01fF
C61134 POR2X1_311/Y PAND2X1_223/B 0.01fF
C61135 PAND2X1_669/CTRL2 POR2X1_750/B 0.01fF
C61136 POR2X1_864/O POR2X1_801/B 0.01fF
C61137 PAND2X1_115/CTRL2 POR2X1_150/Y 0.03fF
C61138 POR2X1_805/CTRL2 PAND2X1_90/Y 0.12fF
C61139 PAND2X1_285/O PAND2X1_805/A 0.02fF
C61140 POR2X1_679/A VDD 0.04fF
C61141 POR2X1_83/B POR2X1_102/Y 0.16fF
C61142 POR2X1_62/Y PAND2X1_529/O 0.03fF
C61143 POR2X1_69/O POR2X1_29/A 0.01fF
C61144 POR2X1_456/B POR2X1_579/O 0.01fF
C61145 PAND2X1_48/B POR2X1_499/A 0.09fF
C61146 PAND2X1_73/Y POR2X1_643/A 0.30fF
C61147 POR2X1_115/CTRL2 POR2X1_76/A 0.01fF
C61148 POR2X1_77/CTRL2 POR2X1_13/A 0.01fF
C61149 PAND2X1_240/O D_INPUT_0 0.05fF
C61150 PAND2X1_474/O POR2X1_293/Y 0.03fF
C61151 POR2X1_669/B POR2X1_94/A 0.05fF
C61152 POR2X1_48/A POR2X1_106/Y 0.01fF
C61153 POR2X1_669/B PAND2X1_731/B 0.02fF
C61154 POR2X1_4/Y POR2X1_342/B 0.01fF
C61155 POR2X1_150/Y PAND2X1_717/CTRL 0.01fF
C61156 POR2X1_202/O POR2X1_296/B 0.31fF
C61157 POR2X1_49/CTRL2 POR2X1_14/Y 0.03fF
C61158 POR2X1_504/Y POR2X1_496/Y 0.02fF
C61159 POR2X1_496/Y PAND2X1_513/CTRL2 0.00fF
C61160 POR2X1_29/A PAND2X1_41/B 0.06fF
C61161 PAND2X1_436/A POR2X1_83/B 0.08fF
C61162 POR2X1_13/A PAND2X1_436/CTRL 0.01fF
C61163 PAND2X1_318/a_56_28# POR2X1_20/B 0.00fF
C61164 POR2X1_856/B POR2X1_480/A 0.10fF
C61165 POR2X1_23/Y PAND2X1_804/A 0.01fF
C61166 PAND2X1_237/CTRL VDD -0.00fF
C61167 POR2X1_665/CTRL2 PAND2X1_645/B 0.05fF
C61168 PAND2X1_137/a_76_28# POR2X1_20/B 0.01fF
C61169 POR2X1_273/Y POR2X1_275/A 0.03fF
C61170 POR2X1_18/a_56_344# D_INPUT_6 0.00fF
C61171 PAND2X1_711/B POR2X1_763/A 0.06fF
C61172 PAND2X1_39/B POR2X1_575/B 0.04fF
C61173 POR2X1_376/B PAND2X1_68/a_76_28# 0.02fF
C61174 POR2X1_848/CTRL POR2X1_713/B 0.30fF
C61175 POR2X1_688/CTRL PAND2X1_32/B 0.01fF
C61176 POR2X1_650/a_16_28# POR2X1_640/Y -0.00fF
C61177 POR2X1_515/a_76_344# PAND2X1_93/B 0.01fF
C61178 D_INPUT_2 POR2X1_612/O 0.02fF
C61179 D_GATE_865 POR2X1_801/B 0.03fF
C61180 POR2X1_23/Y PAND2X1_785/Y 0.03fF
C61181 POR2X1_814/B POR2X1_267/O 0.04fF
C61182 POR2X1_270/Y PAND2X1_57/B 0.06fF
C61183 PAND2X1_277/CTRL POR2X1_546/A 0.02fF
C61184 PAND2X1_48/B POR2X1_76/A 6.39fF
C61185 PAND2X1_16/CTRL2 POR2X1_630/A 0.01fF
C61186 PAND2X1_90/Y POR2X1_174/A 0.03fF
C61187 POR2X1_804/O POR2X1_435/Y 0.05fF
C61188 POR2X1_66/B POR2X1_852/B 0.07fF
C61189 PAND2X1_673/CTRL2 POR2X1_14/Y 0.03fF
C61190 POR2X1_43/CTRL2 POR2X1_39/B 0.00fF
C61191 PAND2X1_816/CTRL2 POR2X1_862/A 0.02fF
C61192 POR2X1_814/B POR2X1_673/CTRL 0.00fF
C61193 POR2X1_411/B PAND2X1_570/a_56_28# 0.00fF
C61194 POR2X1_411/B POR2X1_310/O 0.02fF
C61195 POR2X1_114/B POR2X1_647/B 0.03fF
C61196 POR2X1_821/CTRL2 POR2X1_669/B 0.01fF
C61197 POR2X1_315/Y PAND2X1_717/A 0.07fF
C61198 POR2X1_49/Y POR2X1_60/Y 0.02fF
C61199 PAND2X1_464/B POR2X1_283/A 0.03fF
C61200 PAND2X1_750/a_16_344# POR2X1_816/A 0.01fF
C61201 PAND2X1_55/Y PAND2X1_591/CTRL2 0.03fF
C61202 POR2X1_596/A POR2X1_678/CTRL 0.01fF
C61203 POR2X1_102/Y PAND2X1_140/Y 0.01fF
C61204 POR2X1_658/O POR2X1_318/A 0.03fF
C61205 POR2X1_461/Y POR2X1_532/A 0.10fF
C61206 PAND2X1_849/CTRL2 PAND2X1_61/Y 0.01fF
C61207 POR2X1_467/Y POR2X1_448/A 0.01fF
C61208 POR2X1_260/B D_GATE_222 0.65fF
C61209 POR2X1_835/B POR2X1_566/B 0.05fF
C61210 POR2X1_850/B VDD 0.00fF
C61211 POR2X1_105/CTRL VDD 0.00fF
C61212 POR2X1_441/Y PAND2X1_551/CTRL 0.03fF
C61213 POR2X1_126/CTRL D_INPUT_1 0.01fF
C61214 POR2X1_102/Y PAND2X1_795/B 0.02fF
C61215 POR2X1_20/B POR2X1_387/Y 0.19fF
C61216 POR2X1_647/B POR2X1_649/B 0.15fF
C61217 POR2X1_76/CTRL2 POR2X1_573/A 0.01fF
C61218 POR2X1_260/B POR2X1_140/A 0.01fF
C61219 POR2X1_60/A PAND2X1_738/Y 0.05fF
C61220 POR2X1_174/B POR2X1_355/B 0.07fF
C61221 PAND2X1_41/B POR2X1_213/B 0.00fF
C61222 POR2X1_68/A PAND2X1_93/B 0.18fF
C61223 PAND2X1_203/O POR2X1_91/Y 0.07fF
C61224 PAND2X1_630/CTRL POR2X1_48/A 0.00fF
C61225 PAND2X1_58/A POR2X1_459/O 0.16fF
C61226 PAND2X1_95/O POR2X1_66/A 0.01fF
C61227 POR2X1_72/B POR2X1_236/Y 1.55fF
C61228 PAND2X1_104/CTRL INPUT_0 0.01fF
C61229 PAND2X1_465/CTRL VDD -0.00fF
C61230 PAND2X1_651/Y PAND2X1_436/O 0.45fF
C61231 POR2X1_686/A PAND2X1_90/Y 0.03fF
C61232 PAND2X1_607/CTRL2 POR2X1_294/A 0.09fF
C61233 PAND2X1_241/CTRL2 POR2X1_102/Y 0.01fF
C61234 POR2X1_14/Y POR2X1_395/CTRL2 0.01fF
C61235 POR2X1_376/B POR2X1_5/Y 8.25fF
C61236 POR2X1_65/A POR2X1_511/Y 0.03fF
C61237 POR2X1_445/A POR2X1_318/A 0.29fF
C61238 POR2X1_20/B PAND2X1_121/O 0.04fF
C61239 PAND2X1_795/O INPUT_0 0.05fF
C61240 PAND2X1_90/A PAND2X1_77/CTRL 0.01fF
C61241 POR2X1_416/Y POR2X1_609/Y 0.03fF
C61242 POR2X1_645/CTRL2 PAND2X1_90/Y 0.06fF
C61243 POR2X1_66/B INPUT_5 0.05fF
C61244 POR2X1_175/A POR2X1_192/Y 0.03fF
C61245 POR2X1_629/A POR2X1_629/B 0.00fF
C61246 POR2X1_302/a_16_28# POR2X1_302/B 0.02fF
C61247 POR2X1_42/CTRL2 POR2X1_37/Y 0.01fF
C61248 PAND2X1_59/B POR2X1_407/Y 0.02fF
C61249 POR2X1_178/Y POR2X1_411/B 0.02fF
C61250 POR2X1_333/A POR2X1_785/A 0.05fF
C61251 PAND2X1_159/CTRL POR2X1_55/Y 0.01fF
C61252 POR2X1_257/A PAND2X1_112/CTRL 0.07fF
C61253 POR2X1_614/A POR2X1_801/B 0.08fF
C61254 POR2X1_212/A POR2X1_568/Y 0.05fF
C61255 POR2X1_68/A POR2X1_78/A 0.40fF
C61256 POR2X1_407/A PAND2X1_73/Y 0.04fF
C61257 POR2X1_850/B POR2X1_741/Y 0.03fF
C61258 POR2X1_49/CTRL2 POR2X1_55/Y 0.00fF
C61259 POR2X1_472/O POR2X1_862/A 0.06fF
C61260 PAND2X1_520/CTRL2 POR2X1_236/Y 0.01fF
C61261 POR2X1_192/Y POR2X1_776/O 0.01fF
C61262 PAND2X1_736/A PAND2X1_557/A 0.11fF
C61263 POR2X1_96/A POR2X1_230/CTRL 0.01fF
C61264 PAND2X1_9/CTRL PAND2X1_6/A 0.01fF
C61265 INPUT_3 POR2X1_376/O 0.04fF
C61266 PAND2X1_20/A POR2X1_574/O 0.01fF
C61267 PAND2X1_845/CTRL POR2X1_83/B 0.01fF
C61268 POR2X1_94/CTRL2 POR2X1_94/A 0.03fF
C61269 POR2X1_23/Y PAND2X1_656/A 0.06fF
C61270 PAND2X1_831/Y POR2X1_271/a_16_28# 0.03fF
C61271 POR2X1_201/CTRL POR2X1_35/Y 0.01fF
C61272 POR2X1_423/Y POR2X1_42/Y 0.15fF
C61273 POR2X1_149/B POR2X1_467/Y 0.03fF
C61274 POR2X1_41/B PAND2X1_76/Y 0.07fF
C61275 POR2X1_462/B PAND2X1_58/A 0.24fF
C61276 PAND2X1_51/CTRL POR2X1_635/A 0.01fF
C61277 POR2X1_400/A POR2X1_214/CTRL2 0.00fF
C61278 POR2X1_590/A POR2X1_447/CTRL 0.01fF
C61279 POR2X1_436/a_16_28# POR2X1_802/B 0.03fF
C61280 PAND2X1_58/A D_INPUT_1 1.03fF
C61281 POR2X1_480/A POR2X1_722/Y 0.03fF
C61282 POR2X1_760/A POR2X1_385/Y 0.03fF
C61283 POR2X1_48/A PAND2X1_349/A 0.00fF
C61284 POR2X1_52/A POR2X1_5/Y 2.11fF
C61285 POR2X1_48/A PAND2X1_63/B 0.03fF
C61286 POR2X1_446/B POR2X1_703/Y 1.23fF
C61287 POR2X1_61/Y POR2X1_294/B 0.07fF
C61288 POR2X1_130/CTRL2 POR2X1_260/B 0.01fF
C61289 POR2X1_383/A PAND2X1_237/a_76_28# 0.02fF
C61290 POR2X1_73/CTRL2 D_INPUT_0 0.01fF
C61291 POR2X1_596/A POR2X1_121/B 0.03fF
C61292 POR2X1_124/m4_208_n4# PAND2X1_41/B 0.09fF
C61293 POR2X1_52/A PAND2X1_209/CTRL2 0.03fF
C61294 POR2X1_852/O POR2X1_776/B 0.11fF
C61295 POR2X1_341/A POR2X1_579/B 0.02fF
C61296 PAND2X1_64/CTRL2 POR2X1_260/A 0.01fF
C61297 POR2X1_483/A POR2X1_795/CTRL2 0.04fF
C61298 PAND2X1_20/A POR2X1_844/CTRL2 0.01fF
C61299 PAND2X1_862/B PAND2X1_659/B 0.00fF
C61300 POR2X1_48/A PAND2X1_114/B 1.39fF
C61301 POR2X1_590/A POR2X1_307/A 0.03fF
C61302 PAND2X1_20/A POR2X1_341/Y 0.06fF
C61303 PAND2X1_6/Y POR2X1_244/O 0.08fF
C61304 PAND2X1_275/O POR2X1_274/Y 0.03fF
C61305 POR2X1_355/B POR2X1_544/A 0.01fF
C61306 PAND2X1_573/O PAND2X1_735/Y 0.05fF
C61307 POR2X1_440/Y POR2X1_477/Y 0.03fF
C61308 PAND2X1_621/Y VDD 0.17fF
C61309 POR2X1_653/CTRL POR2X1_661/B 0.01fF
C61310 POR2X1_51/A POR2X1_22/CTRL 0.01fF
C61311 POR2X1_751/A POR2X1_283/A 0.01fF
C61312 POR2X1_502/A POR2X1_220/Y 0.03fF
C61313 PAND2X1_56/Y POR2X1_830/A 0.05fF
C61314 POR2X1_774/Y PAND2X1_583/CTRL2 0.01fF
C61315 PAND2X1_864/B VDD 0.22fF
C61316 POR2X1_639/Y POR2X1_639/CTRL 0.00fF
C61317 POR2X1_276/A POR2X1_296/B 0.01fF
C61318 POR2X1_811/B PAND2X1_60/B 0.03fF
C61319 POR2X1_341/A POR2X1_571/Y 0.03fF
C61320 POR2X1_338/CTRL2 PAND2X1_20/A 0.00fF
C61321 POR2X1_41/B PAND2X1_863/B 0.03fF
C61322 PAND2X1_76/O POR2X1_91/Y 0.01fF
C61323 POR2X1_505/O POR2X1_48/A 0.01fF
C61324 PAND2X1_94/A POR2X1_55/CTRL2 0.00fF
C61325 PAND2X1_385/O VDD 0.00fF
C61326 PAND2X1_216/CTRL2 PAND2X1_364/B 0.03fF
C61327 POR2X1_43/B POR2X1_421/CTRL 0.01fF
C61328 POR2X1_231/A PAND2X1_32/B 0.01fF
C61329 POR2X1_502/A PAND2X1_322/a_76_28# 0.07fF
C61330 PAND2X1_96/B PAND2X1_52/Y 0.03fF
C61331 POR2X1_180/B POR2X1_78/A 0.03fF
C61332 PAND2X1_90/A PAND2X1_38/CTRL 0.01fF
C61333 POR2X1_459/CTRL2 POR2X1_459/A 0.00fF
C61334 POR2X1_362/B POR2X1_513/Y 0.03fF
C61335 PAND2X1_94/A POR2X1_590/A 0.49fF
C61336 PAND2X1_6/Y POR2X1_483/A 0.03fF
C61337 PAND2X1_554/O PAND2X1_348/Y 0.10fF
C61338 PAND2X1_76/Y POR2X1_256/Y 0.00fF
C61339 POR2X1_631/m4_208_n4# POR2X1_219/m4_208_n4# 0.13fF
C61340 POR2X1_262/CTRL PAND2X1_215/B 0.01fF
C61341 POR2X1_32/A PAND2X1_514/O 0.01fF
C61342 PAND2X1_823/CTRL2 POR2X1_836/A 0.01fF
C61343 POR2X1_57/A PAND2X1_220/Y 0.06fF
C61344 POR2X1_305/a_16_28# POR2X1_55/Y 0.02fF
C61345 POR2X1_779/A VDD -0.00fF
C61346 POR2X1_817/a_16_28# POR2X1_394/A 0.04fF
C61347 POR2X1_193/Y POR2X1_532/A 0.03fF
C61348 POR2X1_113/Y POR2X1_389/Y 0.09fF
C61349 POR2X1_368/Y VDD 0.15fF
C61350 PAND2X1_387/CTRL2 PAND2X1_60/B 0.01fF
C61351 PAND2X1_6/Y PAND2X1_8/Y 0.03fF
C61352 POR2X1_474/CTRL2 POR2X1_362/A 0.03fF
C61353 POR2X1_474/CTRL POR2X1_276/Y 0.01fF
C61354 POR2X1_278/Y PAND2X1_794/B 0.03fF
C61355 POR2X1_594/Y PAND2X1_592/Y 0.01fF
C61356 POR2X1_66/B PAND2X1_232/CTRL2 0.01fF
C61357 POR2X1_567/B POR2X1_564/CTRL2 0.03fF
C61358 POR2X1_750/B POR2X1_725/Y 0.07fF
C61359 POR2X1_57/A POR2X1_399/CTRL2 0.09fF
C61360 POR2X1_16/A POR2X1_279/a_16_28# 0.03fF
C61361 POR2X1_850/CTRL2 POR2X1_362/B 0.00fF
C61362 PAND2X1_52/a_16_344# PAND2X1_72/A 0.01fF
C61363 PAND2X1_473/O PAND2X1_741/B 0.01fF
C61364 POR2X1_366/Y POR2X1_317/CTRL 0.08fF
C61365 PAND2X1_218/O PAND2X1_364/B 0.04fF
C61366 PAND2X1_41/B PAND2X1_670/a_56_28# 0.00fF
C61367 PAND2X1_480/B POR2X1_310/CTRL -0.01fF
C61368 POR2X1_294/B POR2X1_193/CTRL 0.03fF
C61369 POR2X1_775/A POR2X1_231/B 0.50fF
C61370 POR2X1_243/O INPUT_0 0.18fF
C61371 POR2X1_43/B PAND2X1_351/O 0.08fF
C61372 POR2X1_294/Y POR2X1_294/A 0.00fF
C61373 POR2X1_832/A PAND2X1_65/B 0.07fF
C61374 POR2X1_43/B POR2X1_275/O 0.15fF
C61375 POR2X1_165/Y POR2X1_83/B 0.04fF
C61376 POR2X1_115/O POR2X1_804/A 0.02fF
C61377 POR2X1_388/O POR2X1_220/Y 0.05fF
C61378 POR2X1_305/Y POR2X1_293/Y 0.01fF
C61379 POR2X1_52/A POR2X1_526/CTRL2 0.03fF
C61380 PAND2X1_652/A PAND2X1_742/B 0.05fF
C61381 POR2X1_220/B POR2X1_192/B 0.05fF
C61382 POR2X1_290/Y PAND2X1_334/a_76_28# 0.01fF
C61383 PAND2X1_631/A POR2X1_23/Y 0.27fF
C61384 PAND2X1_821/CTRL2 POR2X1_510/A 0.00fF
C61385 POR2X1_38/Y POR2X1_88/Y 0.08fF
C61386 POR2X1_35/Y POR2X1_294/B 0.03fF
C61387 PAND2X1_451/O POR2X1_430/Y 0.00fF
C61388 POR2X1_517/Y PAND2X1_642/B 0.02fF
C61389 PAND2X1_658/A PAND2X1_658/B 0.18fF
C61390 POR2X1_239/CTRL POR2X1_7/B 0.01fF
C61391 POR2X1_858/B POR2X1_660/A 0.03fF
C61392 POR2X1_389/Y POR2X1_260/A 0.02fF
C61393 PAND2X1_23/Y POR2X1_249/CTRL 0.01fF
C61394 POR2X1_397/Y PAND2X1_720/CTRL 0.00fF
C61395 POR2X1_141/O POR2X1_141/A 0.02fF
C61396 POR2X1_290/Y POR2X1_73/Y 0.07fF
C61397 POR2X1_537/a_56_344# POR2X1_188/A 0.00fF
C61398 POR2X1_313/Y PAND2X1_714/A 0.03fF
C61399 PAND2X1_41/B POR2X1_520/B 0.01fF
C61400 PAND2X1_784/CTRL2 PAND2X1_778/Y 0.01fF
C61401 POR2X1_468/CTRL POR2X1_478/B 0.00fF
C61402 POR2X1_16/A PAND2X1_204/CTRL2 0.20fF
C61403 POR2X1_186/Y PAND2X1_746/CTRL2 0.37fF
C61404 PAND2X1_383/a_76_28# POR2X1_236/Y 0.02fF
C61405 POR2X1_16/A POR2X1_238/CTRL 0.01fF
C61406 POR2X1_43/B POR2X1_584/O 0.08fF
C61407 PAND2X1_48/B POR2X1_540/A 0.03fF
C61408 PAND2X1_476/A POR2X1_29/A 0.02fF
C61409 PAND2X1_650/O POR2X1_46/Y 0.02fF
C61410 POR2X1_347/CTRL2 POR2X1_296/B 0.00fF
C61411 POR2X1_136/a_16_28# POR2X1_42/Y 0.01fF
C61412 VDD POR2X1_317/A 0.00fF
C61413 POR2X1_57/A PAND2X1_839/CTRL2 0.02fF
C61414 POR2X1_853/A POR2X1_570/B 0.03fF
C61415 POR2X1_853/CTRL2 POR2X1_854/B 0.16fF
C61416 POR2X1_853/A POR2X1_211/a_16_28# 0.12fF
C61417 POR2X1_130/A POR2X1_561/CTRL2 0.01fF
C61418 POR2X1_301/O PAND2X1_6/Y 0.02fF
C61419 PAND2X1_620/Y POR2X1_129/Y 0.03fF
C61420 POR2X1_3/A PAND2X1_709/CTRL 0.01fF
C61421 PAND2X1_658/B POR2X1_73/Y 0.05fF
C61422 POR2X1_469/O POR2X1_478/B 0.01fF
C61423 POR2X1_481/A PAND2X1_336/CTRL 0.01fF
C61424 PAND2X1_90/Y POR2X1_704/Y 0.01fF
C61425 PAND2X1_858/CTRL PAND2X1_390/Y 0.01fF
C61426 POR2X1_779/A PAND2X1_32/B 0.03fF
C61427 PAND2X1_57/B POR2X1_101/Y 0.03fF
C61428 PAND2X1_824/B POR2X1_632/A 0.04fF
C61429 PAND2X1_651/Y POR2X1_521/O 0.02fF
C61430 POR2X1_41/B POR2X1_315/Y 0.07fF
C61431 PAND2X1_126/CTRL2 PAND2X1_90/A 0.01fF
C61432 POR2X1_327/Y POR2X1_449/Y 0.30fF
C61433 POR2X1_339/CTRL VDD -0.00fF
C61434 POR2X1_500/A POR2X1_571/Y 0.00fF
C61435 POR2X1_96/B POR2X1_7/B 1.13fF
C61436 POR2X1_668/Y POR2X1_750/Y 0.13fF
C61437 PAND2X1_794/B POR2X1_761/Y 0.03fF
C61438 POR2X1_3/A POR2X1_22/A 0.03fF
C61439 POR2X1_725/Y POR2X1_777/CTRL2 0.05fF
C61440 PAND2X1_318/CTRL POR2X1_315/Y 0.02fF
C61441 INPUT_1 POR2X1_88/Y 0.03fF
C61442 POR2X1_663/O POR2X1_544/B 0.01fF
C61443 PAND2X1_319/B POR2X1_309/Y 0.07fF
C61444 POR2X1_218/A POR2X1_361/CTRL2 0.00fF
C61445 PAND2X1_96/B D_INPUT_1 0.03fF
C61446 POR2X1_78/A POR2X1_169/A 0.03fF
C61447 POR2X1_32/A POR2X1_39/B 0.96fF
C61448 PAND2X1_644/Y POR2X1_759/CTRL2 0.00fF
C61449 POR2X1_49/Y POR2X1_144/a_16_28# 0.03fF
C61450 PAND2X1_844/B POR2X1_521/O 0.01fF
C61451 POR2X1_515/O POR2X1_574/Y 0.01fF
C61452 D_INPUT_3 PAND2X1_341/a_76_28# 0.03fF
C61453 POR2X1_383/A PAND2X1_519/CTRL2 0.01fF
C61454 POR2X1_68/A PAND2X1_306/O 0.01fF
C61455 POR2X1_65/A PAND2X1_659/Y 0.03fF
C61456 POR2X1_243/Y POR2X1_244/Y 0.01fF
C61457 PAND2X1_20/A POR2X1_554/a_56_344# 0.00fF
C61458 POR2X1_68/B POR2X1_501/B 0.15fF
C61459 PAND2X1_153/O PAND2X1_32/B 0.07fF
C61460 PAND2X1_169/Y PAND2X1_326/B 0.01fF
C61461 POR2X1_428/Y POR2X1_698/Y 0.00fF
C61462 PAND2X1_96/B POR2X1_724/A 0.10fF
C61463 POR2X1_675/A POR2X1_188/Y 0.00fF
C61464 PAND2X1_63/Y POR2X1_318/A 0.10fF
C61465 POR2X1_38/B POR2X1_382/Y 0.02fF
C61466 POR2X1_219/a_76_344# PAND2X1_88/Y 0.00fF
C61467 PAND2X1_631/A PAND2X1_513/CTRL 0.01fF
C61468 PAND2X1_6/A PAND2X1_549/B 0.07fF
C61469 PAND2X1_244/B PAND2X1_658/B 0.07fF
C61470 POR2X1_65/A POR2X1_96/Y 0.03fF
C61471 POR2X1_498/O POR2X1_394/A 0.02fF
C61472 POR2X1_315/a_16_28# POR2X1_91/Y 0.02fF
C61473 PAND2X1_23/Y POR2X1_456/B 0.06fF
C61474 POR2X1_833/CTRL2 POR2X1_260/A 0.01fF
C61475 POR2X1_245/Y POR2X1_90/Y 0.43fF
C61476 VDD POR2X1_113/B 0.45fF
C61477 POR2X1_417/Y POR2X1_39/B 0.03fF
C61478 POR2X1_57/A POR2X1_824/Y 0.03fF
C61479 POR2X1_416/B PAND2X1_556/O 0.02fF
C61480 POR2X1_709/B POR2X1_502/A 0.08fF
C61481 PAND2X1_800/a_56_28# POR2X1_96/A 0.00fF
C61482 PAND2X1_213/Y POR2X1_142/Y 0.03fF
C61483 POR2X1_135/Y POR2X1_135/O 0.01fF
C61484 POR2X1_68/A PAND2X1_6/CTRL 0.00fF
C61485 POR2X1_23/Y PAND2X1_193/Y 0.02fF
C61486 POR2X1_96/A POR2X1_265/Y 0.41fF
C61487 PAND2X1_639/Y VDD 0.10fF
C61488 POR2X1_743/Y POR2X1_153/Y 0.04fF
C61489 POR2X1_192/Y POR2X1_337/Y 0.10fF
C61490 POR2X1_390/B POR2X1_804/A 0.05fF
C61491 PAND2X1_653/Y POR2X1_7/CTRL 0.03fF
C61492 PAND2X1_90/A PAND2X1_527/CTRL2 0.07fF
C61493 POR2X1_327/Y POR2X1_740/Y 0.10fF
C61494 POR2X1_579/Y PAND2X1_171/CTRL 0.01fF
C61495 POR2X1_554/Y POR2X1_735/CTRL 0.01fF
C61496 POR2X1_7/B PAND2X1_507/a_76_28# 0.02fF
C61497 POR2X1_567/B PAND2X1_437/CTRL 0.01fF
C61498 POR2X1_687/A POR2X1_685/B 0.02fF
C61499 POR2X1_220/Y POR2X1_188/Y 0.03fF
C61500 POR2X1_760/Y VDD 0.05fF
C61501 PAND2X1_508/Y POR2X1_55/Y 0.02fF
C61502 POR2X1_43/Y PAND2X1_195/CTRL2 0.01fF
C61503 POR2X1_265/Y POR2X1_406/CTRL 0.01fF
C61504 POR2X1_545/A POR2X1_545/a_16_28# 0.03fF
C61505 POR2X1_257/A POR2X1_431/CTRL 0.01fF
C61506 POR2X1_25/Y POR2X1_47/CTRL2 0.01fF
C61507 POR2X1_43/B PAND2X1_200/B 0.02fF
C61508 POR2X1_772/O PAND2X1_32/B 0.01fF
C61509 PAND2X1_298/O PAND2X1_32/B 0.03fF
C61510 POR2X1_416/B POR2X1_255/a_16_28# 0.02fF
C61511 POR2X1_358/O POR2X1_192/B 0.07fF
C61512 POR2X1_358/CTRL2 POR2X1_191/Y 0.13fF
C61513 PAND2X1_349/A PAND2X1_840/O 0.02fF
C61514 POR2X1_183/Y PAND2X1_853/B 0.03fF
C61515 POR2X1_567/A POR2X1_652/Y 0.19fF
C61516 POR2X1_49/Y PAND2X1_351/A 0.01fF
C61517 PAND2X1_76/Y POR2X1_77/Y 0.12fF
C61518 POR2X1_786/Y POR2X1_186/B 0.18fF
C61519 POR2X1_8/Y POR2X1_38/Y 0.08fF
C61520 POR2X1_712/A POR2X1_774/A 0.03fF
C61521 PAND2X1_476/A POR2X1_406/O 0.00fF
C61522 POR2X1_467/CTRL POR2X1_210/A 0.01fF
C61523 POR2X1_502/A PAND2X1_109/CTRL2 0.10fF
C61524 POR2X1_416/B POR2X1_485/O 0.06fF
C61525 POR2X1_25/Y POR2X1_22/A 0.03fF
C61526 POR2X1_318/A POR2X1_260/A 0.07fF
C61527 POR2X1_297/A POR2X1_77/Y 0.01fF
C61528 POR2X1_287/B PAND2X1_52/B 0.03fF
C61529 POR2X1_16/A PAND2X1_350/CTRL 0.00fF
C61530 PAND2X1_844/Y PAND2X1_338/O 0.02fF
C61531 PAND2X1_530/O POR2X1_4/Y 0.06fF
C61532 PAND2X1_715/B POR2X1_387/Y 0.05fF
C61533 POR2X1_713/B POR2X1_260/A 0.01fF
C61534 PAND2X1_94/Y POR2X1_296/B 0.02fF
C61535 PAND2X1_612/B PAND2X1_612/O 0.01fF
C61536 POR2X1_567/A POR2X1_231/a_16_28# 0.05fF
C61537 POR2X1_57/A PAND2X1_560/B 0.03fF
C61538 POR2X1_76/B POR2X1_330/Y 0.03fF
C61539 POR2X1_569/A POR2X1_576/CTRL 0.02fF
C61540 POR2X1_83/B POR2X1_677/Y 0.04fF
C61541 PAND2X1_35/Y POR2X1_39/B 0.05fF
C61542 PAND2X1_503/O POR2X1_854/B 0.06fF
C61543 POR2X1_567/A POR2X1_35/Y 0.05fF
C61544 PAND2X1_793/Y POR2X1_184/a_16_28# 0.02fF
C61545 POR2X1_765/Y PAND2X1_569/O 0.01fF
C61546 POR2X1_113/B PAND2X1_32/B 0.03fF
C61547 POR2X1_537/Y PAND2X1_69/A 0.03fF
C61548 PAND2X1_657/B POR2X1_73/Y 0.03fF
C61549 POR2X1_83/B POR2X1_9/Y 1.02fF
C61550 POR2X1_209/a_56_344# POR2X1_209/A 0.00fF
C61551 POR2X1_527/a_56_344# PAND2X1_550/B 0.00fF
C61552 PAND2X1_8/Y PAND2X1_52/B 0.19fF
C61553 POR2X1_648/Y POR2X1_807/a_76_344# 0.01fF
C61554 POR2X1_62/Y POR2X1_15/CTRL 0.01fF
C61555 POR2X1_13/A POR2X1_80/CTRL 0.01fF
C61556 PAND2X1_641/Y POR2X1_83/CTRL2 0.04fF
C61557 POR2X1_315/Y PAND2X1_308/Y 0.11fF
C61558 POR2X1_48/A POR2X1_411/A 0.03fF
C61559 POR2X1_510/a_16_28# PAND2X1_72/A 0.00fF
C61560 POR2X1_529/CTRL POR2X1_39/B 0.15fF
C61561 VDD POR2X1_768/A 0.04fF
C61562 POR2X1_327/Y POR2X1_361/a_16_28# 0.02fF
C61563 PAND2X1_639/Y POR2X1_584/a_76_344# 0.00fF
C61564 POR2X1_566/B POR2X1_566/CTRL2 0.01fF
C61565 POR2X1_775/A POR2X1_568/B 0.03fF
C61566 POR2X1_36/B POR2X1_328/CTRL 0.13fF
C61567 POR2X1_8/Y INPUT_1 1.30fF
C61568 POR2X1_83/B POR2X1_827/a_16_28# 0.01fF
C61569 PAND2X1_96/B PAND2X1_134/O 0.03fF
C61570 PAND2X1_798/Y PAND2X1_365/B 0.03fF
C61571 POR2X1_54/Y POR2X1_260/B 0.06fF
C61572 POR2X1_184/Y POR2X1_39/B 0.05fF
C61573 POR2X1_62/Y PAND2X1_63/B 0.10fF
C61574 POR2X1_265/Y POR2X1_7/A 0.12fF
C61575 POR2X1_840/O POR2X1_840/Y 0.00fF
C61576 POR2X1_447/B POR2X1_510/Y 0.00fF
C61577 POR2X1_540/A POR2X1_181/CTRL 0.01fF
C61578 POR2X1_380/Y POR2X1_4/Y 0.03fF
C61579 POR2X1_774/B POR2X1_774/A 0.00fF
C61580 PAND2X1_165/CTRL POR2X1_854/B 0.32fF
C61581 PAND2X1_271/CTRL PAND2X1_93/B 0.01fF
C61582 POR2X1_119/Y PAND2X1_549/B 0.07fF
C61583 PAND2X1_651/Y POR2X1_39/B 1.70fF
C61584 POR2X1_299/a_16_28# PAND2X1_776/Y 0.03fF
C61585 POR2X1_842/O PAND2X1_39/B 0.01fF
C61586 PAND2X1_566/Y POR2X1_77/Y 0.16fF
C61587 POR2X1_8/Y POR2X1_384/A 0.01fF
C61588 PAND2X1_723/A POR2X1_7/Y 0.00fF
C61589 PAND2X1_717/A PAND2X1_558/Y 0.00fF
C61590 POR2X1_309/O POR2X1_150/Y 0.13fF
C61591 POR2X1_188/Y POR2X1_737/CTRL2 0.01fF
C61592 PAND2X1_601/O PAND2X1_93/B 0.02fF
C61593 POR2X1_502/A POR2X1_651/Y 0.03fF
C61594 PAND2X1_407/CTRL POR2X1_409/B 0.01fF
C61595 PAND2X1_446/Y POR2X1_669/B 0.07fF
C61596 POR2X1_278/Y PAND2X1_221/Y 0.07fF
C61597 POR2X1_446/B D_INPUT_0 0.12fF
C61598 PAND2X1_72/A POR2X1_723/B 0.03fF
C61599 POR2X1_316/O POR2X1_129/Y 0.01fF
C61600 D_GATE_741 POR2X1_568/A 0.02fF
C61601 POR2X1_9/Y POR2X1_415/CTRL2 0.05fF
C61602 POR2X1_387/Y POR2X1_372/CTRL2 0.04fF
C61603 PAND2X1_593/Y PAND2X1_643/A 0.01fF
C61604 POR2X1_477/A POR2X1_863/A 0.03fF
C61605 POR2X1_376/B POR2X1_27/O 0.04fF
C61606 POR2X1_165/a_16_28# PAND2X1_326/B 0.02fF
C61607 POR2X1_568/B POR2X1_162/Y 0.05fF
C61608 POR2X1_98/A VDD 0.28fF
C61609 PAND2X1_469/CTRL2 POR2X1_32/A 0.03fF
C61610 POR2X1_257/A POR2X1_279/a_56_344# 0.00fF
C61611 INPUT_3 PAND2X1_58/A 0.08fF
C61612 POR2X1_644/B POR2X1_260/B 0.01fF
C61613 POR2X1_96/A PAND2X1_630/B 0.17fF
C61614 POR2X1_711/Y POR2X1_513/CTRL 0.02fF
C61615 POR2X1_612/Y POR2X1_37/Y 0.03fF
C61616 POR2X1_474/a_16_28# POR2X1_556/A 0.02fF
C61617 POR2X1_416/B POR2X1_142/Y 0.00fF
C61618 POR2X1_768/A PAND2X1_32/B 0.01fF
C61619 PAND2X1_467/Y PAND2X1_452/B 0.01fF
C61620 POR2X1_16/A PAND2X1_326/B 0.00fF
C61621 PAND2X1_65/B PAND2X1_256/O 0.17fF
C61622 POR2X1_161/CTRL2 POR2X1_162/Y 0.01fF
C61623 PAND2X1_480/B PAND2X1_717/A 0.07fF
C61624 POR2X1_48/A POR2X1_32/A 3.65fF
C61625 PAND2X1_47/B PAND2X1_31/CTRL 0.00fF
C61626 POR2X1_333/A PAND2X1_91/a_16_344# 0.04fF
C61627 PAND2X1_39/B PAND2X1_41/B 0.15fF
C61628 PAND2X1_850/Y PAND2X1_853/B 0.46fF
C61629 PAND2X1_510/B POR2X1_80/CTRL 0.01fF
C61630 PAND2X1_93/B PAND2X1_58/A 0.03fF
C61631 PAND2X1_472/CTRL2 POR2X1_77/Y 0.00fF
C61632 POR2X1_490/Y POR2X1_40/Y 0.10fF
C61633 POR2X1_43/B POR2X1_846/A 0.03fF
C61634 D_INPUT_0 POR2X1_121/B 0.06fF
C61635 PAND2X1_384/O POR2X1_383/Y 0.00fF
C61636 POR2X1_846/A POR2X1_789/A 0.12fF
C61637 POR2X1_48/A POR2X1_419/Y 0.06fF
C61638 POR2X1_446/B PAND2X1_90/Y 0.00fF
C61639 POR2X1_483/O POR2X1_556/A 0.01fF
C61640 PAND2X1_435/O POR2X1_411/B 0.02fF
C61641 PAND2X1_698/a_76_28# PAND2X1_52/B 0.01fF
C61642 POR2X1_804/a_56_344# POR2X1_330/Y 0.03fF
C61643 POR2X1_66/B POR2X1_496/Y 0.07fF
C61644 POR2X1_78/A PAND2X1_58/A 0.18fF
C61645 POR2X1_416/B PAND2X1_156/B 0.01fF
C61646 PAND2X1_417/CTRL PAND2X1_55/Y 0.03fF
C61647 POR2X1_257/A PAND2X1_151/O 0.07fF
C61648 PAND2X1_6/Y POR2X1_630/B 0.72fF
C61649 POR2X1_830/Y POR2X1_850/B 0.04fF
C61650 POR2X1_389/A PAND2X1_607/CTRL2 0.10fF
C61651 POR2X1_49/Y PAND2X1_443/m4_208_n4# 0.15fF
C61652 POR2X1_866/A POR2X1_480/A 0.10fF
C61653 POR2X1_400/O POR2X1_400/B 0.00fF
C61654 POR2X1_66/A PAND2X1_16/O 0.02fF
C61655 POR2X1_499/A POR2X1_717/Y 0.03fF
C61656 POR2X1_66/B PAND2X1_39/O 0.01fF
C61657 PAND2X1_865/CTRL PAND2X1_860/A 0.01fF
C61658 POR2X1_65/A POR2X1_37/Y 0.07fF
C61659 PAND2X1_859/a_76_28# POR2X1_93/Y 0.01fF
C61660 POR2X1_816/Y INPUT_0 0.02fF
C61661 POR2X1_708/a_76_344# PAND2X1_39/B 0.01fF
C61662 PAND2X1_414/a_16_344# PAND2X1_6/A 0.01fF
C61663 PAND2X1_630/B POR2X1_7/A 0.04fF
C61664 POR2X1_614/A PAND2X1_426/O 0.17fF
C61665 POR2X1_287/A POR2X1_249/CTRL2 0.01fF
C61666 PAND2X1_319/O POR2X1_48/A 0.04fF
C61667 PAND2X1_657/CTRL PAND2X1_217/B 0.01fF
C61668 POR2X1_566/A POR2X1_447/A 0.05fF
C61669 POR2X1_647/B POR2X1_784/A 0.03fF
C61670 PAND2X1_640/B POR2X1_236/Y 0.03fF
C61671 POR2X1_39/O POR2X1_669/B 0.01fF
C61672 PAND2X1_831/CTRL POR2X1_102/Y 0.00fF
C61673 POR2X1_49/Y PAND2X1_443/Y 0.00fF
C61674 D_INPUT_2 POR2X1_411/B 0.03fF
C61675 POR2X1_102/Y PAND2X1_795/O 0.03fF
C61676 POR2X1_830/a_16_28# PAND2X1_58/A 0.03fF
C61677 POR2X1_159/a_16_28# POR2X1_32/A 0.03fF
C61678 POR2X1_294/CTRL2 POR2X1_294/B 0.00fF
C61679 PAND2X1_629/a_16_344# POR2X1_496/Y 0.00fF
C61680 POR2X1_805/Y PAND2X1_41/B 1.73fF
C61681 PAND2X1_93/B POR2X1_435/Y 0.07fF
C61682 POR2X1_678/A POR2X1_330/Y 0.28fF
C61683 POR2X1_54/Y PAND2X1_55/Y 0.08fF
C61684 POR2X1_495/Y POR2X1_257/A 0.12fF
C61685 PAND2X1_20/A PAND2X1_41/B 0.16fF
C61686 POR2X1_460/Y PAND2X1_752/Y 0.02fF
C61687 POR2X1_775/A POR2X1_341/A 0.02fF
C61688 PAND2X1_404/Y PAND2X1_364/B 0.07fF
C61689 POR2X1_32/A PAND2X1_199/A 0.03fF
C61690 PAND2X1_71/a_56_28# PAND2X1_39/B 0.00fF
C61691 POR2X1_96/A PAND2X1_776/Y 0.29fF
C61692 POR2X1_814/A POR2X1_780/B 0.05fF
C61693 POR2X1_774/Y POR2X1_866/CTRL2 0.01fF
C61694 POR2X1_254/A POR2X1_254/O 0.01fF
C61695 PAND2X1_55/Y POR2X1_202/A 0.11fF
C61696 POR2X1_121/B PAND2X1_90/Y 0.10fF
C61697 PAND2X1_621/Y POR2X1_818/Y 0.01fF
C61698 PAND2X1_217/B POR2X1_272/O 0.03fF
C61699 POR2X1_137/B PAND2X1_96/B 0.08fF
C61700 PAND2X1_217/B PAND2X1_390/Y 0.05fF
C61701 POR2X1_23/Y PAND2X1_775/CTRL 0.10fF
C61702 POR2X1_254/O POR2X1_750/B 0.02fF
C61703 POR2X1_730/B POR2X1_452/Y 0.76fF
C61704 PAND2X1_205/Y POR2X1_40/Y 0.05fF
C61705 POR2X1_492/O PAND2X1_558/Y 0.17fF
C61706 POR2X1_800/A POR2X1_808/O 0.00fF
C61707 POR2X1_341/A POR2X1_112/Y 0.11fF
C61708 POR2X1_634/O POR2X1_640/A 0.01fF
C61709 PAND2X1_23/Y PAND2X1_94/CTRL2 0.00fF
C61710 POR2X1_416/Y PAND2X1_606/CTRL 0.01fF
C61711 D_INPUT_0 PAND2X1_351/CTRL 0.11fF
C61712 PAND2X1_392/B PAND2X1_390/Y 0.07fF
C61713 POR2X1_402/A POR2X1_202/A 0.12fF
C61714 D_INPUT_3 POR2X1_20/B 0.03fF
C61715 POR2X1_78/A POR2X1_435/Y 0.07fF
C61716 POR2X1_814/B PAND2X1_41/B 0.72fF
C61717 POR2X1_188/A POR2X1_285/CTRL2 0.01fF
C61718 POR2X1_453/a_16_28# POR2X1_449/Y 0.04fF
C61719 PAND2X1_254/Y POR2X1_496/Y 0.03fF
C61720 POR2X1_96/A POR2X1_283/a_16_28# 0.02fF
C61721 PAND2X1_20/A POR2X1_402/B 0.01fF
C61722 PAND2X1_787/A PAND2X1_211/CTRL2 0.00fF
C61723 POR2X1_13/A POR2X1_603/Y 0.01fF
C61724 POR2X1_814/B POR2X1_461/a_56_344# 0.00fF
C61725 POR2X1_673/CTRL VDD 0.00fF
C61726 PAND2X1_272/O POR2X1_193/A 0.02fF
C61727 PAND2X1_676/O POR2X1_257/A 0.02fF
C61728 PAND2X1_659/CTRL2 POR2X1_72/B 0.03fF
C61729 POR2X1_272/CTRL POR2X1_272/Y 0.06fF
C61730 POR2X1_692/a_16_28# POR2X1_763/Y 0.04fF
C61731 PAND2X1_695/CTRL PAND2X1_41/B 0.01fF
C61732 POR2X1_686/O PAND2X1_39/B 0.07fF
C61733 POR2X1_346/A PAND2X1_55/Y 0.05fF
C61734 POR2X1_609/CTRL2 POR2X1_609/A 0.01fF
C61735 POR2X1_48/A POR2X1_184/Y 0.03fF
C61736 POR2X1_617/Y POR2X1_9/Y 0.03fF
C61737 POR2X1_669/B POR2X1_252/a_16_28# 0.11fF
C61738 POR2X1_222/CTRL POR2X1_724/A 0.02fF
C61739 PAND2X1_390/Y VDD 0.99fF
C61740 POR2X1_457/CTRL POR2X1_220/Y 0.02fF
C61741 PAND2X1_600/CTRL2 PAND2X1_32/B 0.03fF
C61742 PAND2X1_48/B POR2X1_247/Y 0.01fF
C61743 POR2X1_625/CTRL POR2X1_5/Y 0.01fF
C61744 PAND2X1_675/A PAND2X1_352/A 0.10fF
C61745 POR2X1_661/Y PAND2X1_55/Y 0.00fF
C61746 POR2X1_423/Y PAND2X1_139/Y 0.00fF
C61747 POR2X1_434/O POR2X1_209/A 0.01fF
C61748 PAND2X1_651/Y POR2X1_48/A 1.60fF
C61749 PAND2X1_118/CTRL2 PAND2X1_73/Y 0.09fF
C61750 PAND2X1_93/B PAND2X1_96/B 0.06fF
C61751 POR2X1_445/A POR2X1_540/a_16_28# -0.00fF
C61752 POR2X1_857/O POR2X1_785/A 0.16fF
C61753 PAND2X1_68/O PAND2X1_6/A 0.08fF
C61754 PAND2X1_260/O POR2X1_13/A -0.00fF
C61755 POR2X1_411/B PAND2X1_346/Y 0.03fF
C61756 POR2X1_389/O POR2X1_121/B 0.01fF
C61757 POR2X1_23/Y PAND2X1_243/O 0.02fF
C61758 POR2X1_52/A POR2X1_491/CTRL 0.01fF
C61759 POR2X1_72/a_16_28# PAND2X1_499/Y 0.13fF
C61760 POR2X1_750/B PAND2X1_176/CTRL 0.01fF
C61761 POR2X1_644/B POR2X1_407/Y 0.03fF
C61762 PAND2X1_57/B PAND2X1_597/CTRL 0.01fF
C61763 POR2X1_801/B PAND2X1_583/O 0.01fF
C61764 POR2X1_362/Y POR2X1_68/A 0.36fF
C61765 POR2X1_96/A PAND2X1_192/CTRL 0.01fF
C61766 PAND2X1_564/B PAND2X1_551/Y 0.00fF
C61767 PAND2X1_862/B POR2X1_5/Y 0.23fF
C61768 PAND2X1_620/Y POR2X1_293/Y 0.07fF
C61769 POR2X1_677/Y PAND2X1_841/Y 0.02fF
C61770 PAND2X1_798/B PAND2X1_575/B 0.89fF
C61771 INPUT_0 POR2X1_372/O 0.04fF
C61772 POR2X1_794/CTRL VDD 0.00fF
C61773 PAND2X1_23/CTRL PAND2X1_55/Y 0.01fF
C61774 POR2X1_66/A POR2X1_307/A 0.07fF
C61775 POR2X1_65/A POR2X1_293/Y 0.11fF
C61776 PAND2X1_96/B POR2X1_78/A 0.19fF
C61777 POR2X1_66/B POR2X1_790/A 0.03fF
C61778 POR2X1_263/Y POR2X1_235/CTRL2 0.01fF
C61779 POR2X1_865/O POR2X1_590/A 0.02fF
C61780 PAND2X1_658/A PAND2X1_185/CTRL 0.01fF
C61781 POR2X1_254/Y VDD 1.24fF
C61782 POR2X1_121/B PAND2X1_583/a_16_344# 0.04fF
C61783 POR2X1_41/B PAND2X1_596/O 0.15fF
C61784 POR2X1_411/B PAND2X1_502/O 0.02fF
C61785 POR2X1_467/Y POR2X1_535/a_16_28# 0.02fF
C61786 POR2X1_98/B POR2X1_590/A 0.02fF
C61787 PAND2X1_7/CTRL PAND2X1_52/Y 0.01fF
C61788 POR2X1_383/A D_INPUT_0 0.17fF
C61789 PAND2X1_659/O PAND2X1_735/Y 0.07fF
C61790 POR2X1_78/A POR2X1_216/CTRL2 0.01fF
C61791 PAND2X1_50/O INPUT_5 0.01fF
C61792 POR2X1_278/Y PAND2X1_795/B 0.07fF
C61793 POR2X1_7/B POR2X1_236/Y 0.17fF
C61794 PAND2X1_621/CTRL POR2X1_818/Y 0.01fF
C61795 POR2X1_498/CTRL2 PAND2X1_735/Y 0.03fF
C61796 POR2X1_840/B POR2X1_287/a_16_28# 0.05fF
C61797 POR2X1_346/B POR2X1_195/A 0.02fF
C61798 POR2X1_296/B PAND2X1_60/B 1.21fF
C61799 PAND2X1_651/Y PAND2X1_512/O 0.00fF
C61800 POR2X1_814/B PAND2X1_411/CTRL 0.01fF
C61801 POR2X1_558/A POR2X1_78/A 0.03fF
C61802 PAND2X1_416/m4_208_n4# POR2X1_260/A 0.15fF
C61803 POR2X1_844/m4_208_n4# POR2X1_590/A 0.15fF
C61804 POR2X1_614/A PAND2X1_279/a_76_28# 0.02fF
C61805 POR2X1_66/B PAND2X1_88/Y 0.04fF
C61806 POR2X1_631/a_16_28# POR2X1_631/B 0.01fF
C61807 POR2X1_829/O POR2X1_761/Y 0.01fF
C61808 POR2X1_41/B PAND2X1_480/B 0.10fF
C61809 POR2X1_467/Y POR2X1_209/A 0.03fF
C61810 PAND2X1_94/A POR2X1_66/A 0.15fF
C61811 PAND2X1_58/A PAND2X1_306/O 0.05fF
C61812 POR2X1_83/Y POR2X1_20/B 2.05fF
C61813 POR2X1_630/B POR2X1_632/Y 0.09fF
C61814 PAND2X1_687/Y POR2X1_42/Y 0.03fF
C61815 PAND2X1_23/Y PAND2X1_131/CTRL2 0.01fF
C61816 PAND2X1_137/Y POR2X1_96/A 0.12fF
C61817 PAND2X1_20/A POR2X1_228/Y 0.03fF
C61818 PAND2X1_140/A POR2X1_102/Y 0.12fF
C61819 PAND2X1_226/O POR2X1_241/Y 0.01fF
C61820 D_GATE_222 PAND2X1_164/CTRL2 0.03fF
C61821 PAND2X1_185/CTRL POR2X1_73/Y 0.01fF
C61822 POR2X1_575/B VDD 0.47fF
C61823 POR2X1_302/CTRL2 POR2X1_114/B 0.01fF
C61824 POR2X1_41/B POR2X1_754/A 0.02fF
C61825 POR2X1_325/A POR2X1_130/Y 0.03fF
C61826 POR2X1_528/Y POR2X1_102/Y 0.03fF
C61827 PAND2X1_857/B POR2X1_83/B 0.04fF
C61828 POR2X1_549/CTRL2 POR2X1_68/B 0.01fF
C61829 PAND2X1_778/a_76_28# POR2X1_55/Y 0.01fF
C61830 PAND2X1_652/A PAND2X1_580/B 0.00fF
C61831 POR2X1_65/A PAND2X1_553/CTRL 0.00fF
C61832 PAND2X1_23/Y PAND2X1_57/B 12.35fF
C61833 PAND2X1_42/O POR2X1_68/B 0.02fF
C61834 PAND2X1_434/O POR2X1_129/Y 0.02fF
C61835 PAND2X1_48/B POR2X1_663/m4_208_n4# 0.09fF
C61836 POR2X1_254/CTRL POR2X1_228/Y 0.01fF
C61837 PAND2X1_182/A POR2X1_55/Y 0.00fF
C61838 POR2X1_614/A POR2X1_549/B 0.02fF
C61839 POR2X1_174/B POR2X1_174/CTRL2 0.03fF
C61840 POR2X1_254/Y POR2X1_741/Y 0.07fF
C61841 PAND2X1_96/B POR2X1_573/CTRL 0.01fF
C61842 POR2X1_217/a_16_28# POR2X1_572/B 0.03fF
C61843 POR2X1_417/CTRL POR2X1_5/Y 0.01fF
C61844 PAND2X1_654/A POR2X1_409/B 0.06fF
C61845 POR2X1_574/O VDD -0.00fF
C61846 POR2X1_141/Y POR2X1_510/Y 0.14fF
C61847 POR2X1_113/O POR2X1_640/Y 0.02fF
C61848 POR2X1_230/CTRL POR2X1_38/Y 0.04fF
C61849 POR2X1_350/Y VDD 0.10fF
C61850 PAND2X1_48/B PAND2X1_371/CTRL 0.00fF
C61851 GATE_741 PAND2X1_794/B 0.03fF
C61852 PAND2X1_857/A POR2X1_40/Y 1.51fF
C61853 POR2X1_159/a_56_344# POR2X1_408/Y 0.03fF
C61854 POR2X1_491/Y POR2X1_411/B 0.01fF
C61855 POR2X1_742/a_16_28# POR2X1_741/Y 0.11fF
C61856 PAND2X1_254/Y PAND2X1_514/Y 0.00fF
C61857 PAND2X1_349/A PAND2X1_349/B 0.07fF
C61858 POR2X1_593/B POR2X1_592/CTRL 0.01fF
C61859 POR2X1_343/Y PAND2X1_256/a_16_344# 0.02fF
C61860 POR2X1_813/CTRL2 POR2X1_39/B 0.24fF
C61861 POR2X1_38/B POR2X1_549/B 0.03fF
C61862 POR2X1_502/A POR2X1_114/B 0.15fF
C61863 POR2X1_814/B POR2X1_228/Y 2.22fF
C61864 POR2X1_859/A POR2X1_790/A 0.09fF
C61865 POR2X1_850/CTRL POR2X1_850/A 0.01fF
C61866 PAND2X1_434/CTRL2 POR2X1_72/B 0.01fF
C61867 PAND2X1_58/O PAND2X1_69/A 0.05fF
C61868 POR2X1_795/O POR2X1_294/B 0.01fF
C61869 PAND2X1_374/O POR2X1_40/Y 0.04fF
C61870 POR2X1_356/A POR2X1_853/A 0.05fF
C61871 PAND2X1_684/O POR2X1_78/A 0.01fF
C61872 POR2X1_841/B POR2X1_188/Y 0.03fF
C61873 PAND2X1_391/m4_208_n4# POR2X1_384/m4_208_n4# 0.04fF
C61874 PAND2X1_391/CTRL POR2X1_384/Y 0.00fF
C61875 POR2X1_590/A POR2X1_733/Y 0.01fF
C61876 POR2X1_389/Y POR2X1_725/Y 0.02fF
C61877 POR2X1_62/Y PAND2X1_10/CTRL2 0.00fF
C61878 PAND2X1_340/CTRL2 POR2X1_7/A 0.01fF
C61879 POR2X1_550/A PAND2X1_525/CTRL 0.01fF
C61880 POR2X1_71/Y PAND2X1_798/B 0.00fF
C61881 POR2X1_66/B PAND2X1_376/O 0.01fF
C61882 POR2X1_802/a_76_344# POR2X1_750/B 0.01fF
C61883 POR2X1_49/Y PAND2X1_723/A 0.07fF
C61884 POR2X1_844/CTRL2 VDD 0.00fF
C61885 POR2X1_254/Y PAND2X1_32/B 0.29fF
C61886 POR2X1_341/Y VDD -0.00fF
C61887 PAND2X1_672/O D_INPUT_0 0.06fF
C61888 POR2X1_575/B POR2X1_501/CTRL2 0.10fF
C61889 POR2X1_141/Y POR2X1_276/Y 0.01fF
C61890 PAND2X1_643/CTRL2 POR2X1_13/Y 0.01fF
C61891 PAND2X1_94/A PAND2X1_88/a_16_344# 0.02fF
C61892 POR2X1_397/Y PAND2X1_338/B 0.02fF
C61893 POR2X1_717/m4_208_n4# POR2X1_475/A 0.15fF
C61894 PAND2X1_836/CTRL2 POR2X1_293/Y 0.00fF
C61895 PAND2X1_798/B POR2X1_42/Y 0.07fF
C61896 POR2X1_335/A POR2X1_740/Y 0.21fF
C61897 POR2X1_325/A POR2X1_228/Y 0.03fF
C61898 POR2X1_383/A PAND2X1_90/Y 0.92fF
C61899 PAND2X1_283/O POR2X1_294/B 0.02fF
C61900 POR2X1_62/Y POR2X1_32/A 0.12fF
C61901 PAND2X1_453/O PAND2X1_449/Y 0.00fF
C61902 POR2X1_547/B PAND2X1_60/B 0.03fF
C61903 POR2X1_35/B POR2X1_260/A 0.00fF
C61904 PAND2X1_55/Y PAND2X1_29/CTRL 0.00fF
C61905 PAND2X1_149/a_76_28# PAND2X1_148/Y 0.01fF
C61906 POR2X1_697/Y POR2X1_531/Y 0.01fF
C61907 POR2X1_43/B POR2X1_45/Y 0.03fF
C61908 PAND2X1_48/B POR2X1_219/CTRL2 0.01fF
C61909 PAND2X1_6/Y PAND2X1_599/CTRL 0.01fF
C61910 POR2X1_556/A POR2X1_717/B 0.03fF
C61911 PAND2X1_808/Y PAND2X1_357/Y 0.03fF
C61912 POR2X1_488/a_16_28# POR2X1_283/A 0.07fF
C61913 PAND2X1_793/Y POR2X1_93/A 0.03fF
C61914 PAND2X1_429/Y INPUT_6 0.00fF
C61915 POR2X1_785/A POR2X1_556/Y 0.03fF
C61916 POR2X1_741/Y POR2X1_574/O 0.10fF
C61917 PAND2X1_48/B PAND2X1_69/A 5.53fF
C61918 POR2X1_437/CTRL2 PAND2X1_580/B 0.00fF
C61919 PAND2X1_284/O PAND2X1_566/Y 0.00fF
C61920 PAND2X1_793/Y POR2X1_91/Y 0.03fF
C61921 POR2X1_437/Y PAND2X1_794/B 0.01fF
C61922 POR2X1_575/B PAND2X1_32/B 0.07fF
C61923 PAND2X1_472/A PAND2X1_401/O 0.05fF
C61924 POR2X1_220/Y POR2X1_510/Y 0.03fF
C61925 PAND2X1_625/CTRL PAND2X1_69/A 0.01fF
C61926 PAND2X1_211/A PAND2X1_853/B 0.01fF
C61927 POR2X1_111/Y PAND2X1_332/O 0.07fF
C61928 POR2X1_631/A POR2X1_294/B 0.10fF
C61929 POR2X1_278/Y POR2X1_187/CTRL 0.08fF
C61930 POR2X1_48/A POR2X1_524/a_16_28# 0.01fF
C61931 PAND2X1_115/B POR2X1_387/Y 0.29fF
C61932 PAND2X1_94/A PAND2X1_293/O 0.03fF
C61933 PAND2X1_804/B PAND2X1_175/CTRL2 0.01fF
C61934 POR2X1_776/B POR2X1_854/B 1.47fF
C61935 POR2X1_139/Y POR2X1_383/A 0.01fF
C61936 PAND2X1_106/CTRL PAND2X1_48/B 0.01fF
C61937 POR2X1_335/a_16_28# POR2X1_337/A 0.07fF
C61938 PAND2X1_458/O PAND2X1_464/B 0.00fF
C61939 POR2X1_707/CTRL PAND2X1_57/B 0.01fF
C61940 POR2X1_764/CTRL VDD 0.00fF
C61941 POR2X1_416/B POR2X1_409/B 0.14fF
C61942 POR2X1_283/A POR2X1_55/Y 0.17fF
C61943 PAND2X1_252/O POR2X1_556/Y 0.17fF
C61944 VDD POR2X1_731/A 0.00fF
C61945 PAND2X1_79/Y POR2X1_786/Y 0.17fF
C61946 POR2X1_574/CTRL2 POR2X1_574/A 0.01fF
C61947 POR2X1_533/A POR2X1_533/a_16_28# 0.12fF
C61948 POR2X1_528/CTRL2 POR2X1_528/Y 0.01fF
C61949 POR2X1_257/A PAND2X1_860/A 0.03fF
C61950 POR2X1_404/Y POR2X1_276/Y 0.12fF
C61951 POR2X1_324/A POR2X1_324/Y 0.01fF
C61952 PAND2X1_480/B PAND2X1_308/Y 0.05fF
C61953 POR2X1_511/Y PAND2X1_508/Y 0.03fF
C61954 POR2X1_853/A POR2X1_569/A 0.08fF
C61955 POR2X1_5/Y PAND2X1_716/B 0.03fF
C61956 POR2X1_532/A POR2X1_140/CTRL2 0.01fF
C61957 POR2X1_314/CTRL POR2X1_16/A 0.01fF
C61958 POR2X1_23/Y POR2X1_49/O 0.01fF
C61959 POR2X1_57/A PAND2X1_724/CTRL 0.01fF
C61960 PAND2X1_691/Y POR2X1_42/Y 0.06fF
C61961 PAND2X1_356/a_16_344# POR2X1_42/Y 0.02fF
C61962 PAND2X1_575/B POR2X1_184/O 0.01fF
C61963 POR2X1_261/A PAND2X1_345/Y 0.03fF
C61964 POR2X1_800/A POR2X1_796/A -0.00fF
C61965 D_INPUT_1 POR2X1_380/Y 0.03fF
C61966 POR2X1_355/B POR2X1_544/B 0.03fF
C61967 INPUT_1 POR2X1_618/a_56_344# 0.00fF
C61968 POR2X1_192/Y POR2X1_566/CTRL 0.13fF
C61969 POR2X1_96/A PAND2X1_853/B 0.03fF
C61970 PAND2X1_763/O PAND2X1_48/A 0.09fF
C61971 POR2X1_387/Y POR2X1_73/Y 0.07fF
C61972 POR2X1_614/A POR2X1_855/B 0.03fF
C61973 POR2X1_853/A POR2X1_570/Y 0.48fF
C61974 POR2X1_711/B VDD 0.06fF
C61975 PAND2X1_48/B PAND2X1_824/B 0.02fF
C61976 POR2X1_347/A PAND2X1_55/Y 1.87fF
C61977 POR2X1_60/A POR2X1_80/CTRL2 0.03fF
C61978 PAND2X1_6/Y POR2X1_259/CTRL 0.01fF
C61979 POR2X1_383/A POR2X1_865/CTRL 0.01fF
C61980 POR2X1_41/B POR2X1_373/Y 0.04fF
C61981 PAND2X1_546/Y PAND2X1_726/B 0.02fF
C61982 POR2X1_94/A POR2X1_39/B 0.07fF
C61983 PAND2X1_367/CTRL2 VDD 0.00fF
C61984 POR2X1_802/CTRL POR2X1_532/A 0.01fF
C61985 PAND2X1_731/B POR2X1_39/B 0.12fF
C61986 PAND2X1_691/Y PAND2X1_664/O 0.01fF
C61987 POR2X1_313/Y PAND2X1_675/A 0.01fF
C61988 PAND2X1_206/A POR2X1_9/Y 0.01fF
C61989 POR2X1_52/A PAND2X1_123/Y 0.03fF
C61990 POR2X1_509/A PAND2X1_503/O 0.00fF
C61991 PAND2X1_295/CTRL POR2X1_837/B 0.00fF
C61992 POR2X1_316/O POR2X1_293/Y 0.02fF
C61993 POR2X1_52/A PAND2X1_502/O 0.04fF
C61994 POR2X1_16/A PAND2X1_794/B 0.00fF
C61995 PAND2X1_23/Y PAND2X1_701/O 0.00fF
C61996 POR2X1_537/Y POR2X1_121/Y 0.23fF
C61997 POR2X1_24/O POR2X1_77/Y 0.02fF
C61998 POR2X1_62/Y PAND2X1_197/CTRL2 0.01fF
C61999 POR2X1_347/A POR2X1_402/A 0.04fF
C62000 POR2X1_180/B POR2X1_540/CTRL 0.00fF
C62001 POR2X1_130/A PAND2X1_304/CTRL2 0.01fF
C62002 PAND2X1_23/Y POR2X1_227/O 0.08fF
C62003 POR2X1_16/A PAND2X1_723/O 0.01fF
C62004 PAND2X1_386/a_56_28# D_INPUT_4 0.00fF
C62005 POR2X1_57/A POR2X1_527/CTRL2 0.01fF
C62006 POR2X1_383/A POR2X1_361/O 0.01fF
C62007 PAND2X1_119/O PAND2X1_94/A 0.00fF
C62008 POR2X1_730/Y POR2X1_156/B 0.03fF
C62009 POR2X1_390/B PAND2X1_311/O 0.00fF
C62010 PAND2X1_787/O POR2X1_77/Y 0.03fF
C62011 PAND2X1_94/A POR2X1_532/A 0.13fF
C62012 POR2X1_137/Y POR2X1_101/Y 0.05fF
C62013 POR2X1_502/A PAND2X1_665/CTRL2 0.01fF
C62014 POR2X1_447/B POR2X1_578/Y 0.03fF
C62015 INPUT_1 POR2X1_68/B 0.17fF
C62016 POR2X1_590/A POR2X1_303/B 0.01fF
C62017 PAND2X1_801/CTRL2 PAND2X1_863/B 0.01fF
C62018 POR2X1_545/A POR2X1_564/B 0.17fF
C62019 PAND2X1_661/Y PAND2X1_194/a_16_344# 0.02fF
C62020 POR2X1_814/A POR2X1_647/CTRL2 0.04fF
C62021 PAND2X1_530/O POR2X1_620/B 0.02fF
C62022 POR2X1_821/CTRL2 POR2X1_39/B 0.00fF
C62023 PAND2X1_55/Y POR2X1_4/Y 0.03fF
C62024 POR2X1_828/Y PAND2X1_72/A 0.03fF
C62025 POR2X1_189/CTRL PAND2X1_480/B 0.29fF
C62026 POR2X1_394/A PAND2X1_645/B 0.07fF
C62027 POR2X1_145/CTRL PAND2X1_797/Y 0.01fF
C62028 POR2X1_845/CTRL2 POR2X1_673/Y 0.03fF
C62029 PAND2X1_632/A PAND2X1_508/CTRL2 0.01fF
C62030 POR2X1_541/B POR2X1_341/A 0.08fF
C62031 POR2X1_809/A POR2X1_828/A 0.03fF
C62032 POR2X1_51/A POR2X1_39/B 0.05fF
C62033 POR2X1_566/B POR2X1_192/CTRL2 0.02fF
C62034 POR2X1_778/B PAND2X1_48/A 0.08fF
C62035 POR2X1_62/Y PAND2X1_651/Y 0.03fF
C62036 PAND2X1_629/a_76_28# POR2X1_626/Y 0.02fF
C62037 POR2X1_410/CTRL2 PAND2X1_52/B 0.01fF
C62038 POR2X1_52/A POR2X1_491/Y 0.54fF
C62039 POR2X1_114/B POR2X1_188/Y 1.75fF
C62040 POR2X1_366/CTRL POR2X1_276/Y 0.04fF
C62041 PAND2X1_308/Y PAND2X1_303/B 0.01fF
C62042 PAND2X1_631/A PAND2X1_658/B 0.16fF
C62043 POR2X1_257/A POR2X1_253/CTRL2 0.01fF
C62044 PAND2X1_57/B POR2X1_711/Y 0.07fF
C62045 POR2X1_68/B POR2X1_768/Y 0.01fF
C62046 PAND2X1_480/B POR2X1_77/Y 0.05fF
C62047 POR2X1_554/B POR2X1_274/A 0.03fF
C62048 PAND2X1_326/B PAND2X1_324/Y 0.17fF
C62049 POR2X1_773/B POR2X1_116/Y 0.27fF
C62050 POR2X1_462/CTRL2 POR2X1_66/A 0.01fF
C62051 POR2X1_304/CTRL2 POR2X1_43/B 0.03fF
C62052 POR2X1_814/A POR2X1_210/CTRL2 0.02fF
C62053 PAND2X1_9/Y PAND2X1_407/O 0.02fF
C62054 POR2X1_62/Y PAND2X1_844/B 0.10fF
C62055 POR2X1_65/A PAND2X1_242/Y 0.03fF
C62056 POR2X1_571/Y POR2X1_500/Y 0.01fF
C62057 POR2X1_265/Y POR2X1_38/Y 0.02fF
C62058 POR2X1_317/O POR2X1_169/A 0.00fF
C62059 POR2X1_833/A POR2X1_101/Y 0.10fF
C62060 POR2X1_7/A PAND2X1_853/B 0.05fF
C62061 PAND2X1_65/B POR2X1_535/CTRL 0.01fF
C62062 PAND2X1_831/CTRL POR2X1_677/Y 0.00fF
C62063 POR2X1_332/Y POR2X1_228/Y 0.34fF
C62064 POR2X1_591/Y POR2X1_385/Y 0.12fF
C62065 POR2X1_76/Y POR2X1_715/CTRL 0.01fF
C62066 POR2X1_366/Y POR2X1_736/A 0.10fF
C62067 PAND2X1_634/CTRL2 POR2X1_37/Y 0.03fF
C62068 POR2X1_614/A PAND2X1_143/a_76_28# 0.01fF
C62069 PAND2X1_426/CTRL2 POR2X1_121/B 0.01fF
C62070 PAND2X1_469/B POR2X1_589/a_56_344# 0.00fF
C62071 POR2X1_57/A PAND2X1_352/B 0.04fF
C62072 PAND2X1_737/B POR2X1_394/A 0.03fF
C62073 POR2X1_673/Y POR2X1_546/a_76_344# 0.01fF
C62074 POR2X1_249/Y POR2X1_774/A 0.03fF
C62075 POR2X1_59/CTRL POR2X1_394/A 0.01fF
C62076 POR2X1_191/Y POR2X1_319/Y 0.03fF
C62077 PAND2X1_216/B POR2X1_394/A 0.03fF
C62078 PAND2X1_599/CTRL PAND2X1_52/B 0.01fF
C62079 PAND2X1_63/O PAND2X1_9/Y 0.17fF
C62080 PAND2X1_222/A PAND2X1_267/Y 0.01fF
C62081 PAND2X1_508/Y PAND2X1_861/CTRL 0.00fF
C62082 POR2X1_188/a_16_28# POR2X1_737/A 0.01fF
C62083 POR2X1_705/B POR2X1_590/A 0.01fF
C62084 POR2X1_329/A POR2X1_40/Y 0.10fF
C62085 POR2X1_264/Y PAND2X1_52/B 0.03fF
C62086 PAND2X1_109/O PAND2X1_32/B 0.01fF
C62087 PAND2X1_6/Y POR2X1_343/Y 0.03fF
C62088 PAND2X1_308/Y PAND2X1_727/a_76_28# 0.01fF
C62089 POR2X1_817/O PAND2X1_340/B 0.01fF
C62090 POR2X1_853/A PAND2X1_72/A 0.03fF
C62091 PAND2X1_221/Y PAND2X1_730/B 0.00fF
C62092 PAND2X1_289/O POR2X1_220/B 0.01fF
C62093 PAND2X1_221/Y GATE_741 0.03fF
C62094 POR2X1_510/Y POR2X1_554/CTRL 0.01fF
C62095 POR2X1_182/CTRL POR2X1_854/B 0.33fF
C62096 POR2X1_23/Y POR2X1_437/CTRL 0.01fF
C62097 POR2X1_772/CTRL POR2X1_113/B 0.01fF
C62098 POR2X1_51/CTRL POR2X1_51/B 0.01fF
C62099 PAND2X1_535/Y POR2X1_533/Y 0.06fF
C62100 PAND2X1_56/Y POR2X1_715/O 0.03fF
C62101 POR2X1_66/B POR2X1_658/CTRL2 0.01fF
C62102 POR2X1_21/O D_INPUT_4 0.00fF
C62103 POR2X1_434/CTRL2 POR2X1_434/A 0.01fF
C62104 POR2X1_93/m4_208_n4# POR2X1_39/B 0.05fF
C62105 PAND2X1_508/Y POR2X1_129/Y 0.03fF
C62106 D_INPUT_7 VDD 0.64fF
C62107 POR2X1_90/Y PAND2X1_326/a_16_344# 0.02fF
C62108 POR2X1_343/Y POR2X1_575/CTRL2 0.13fF
C62109 POR2X1_648/Y PAND2X1_90/Y 0.09fF
C62110 POR2X1_464/a_16_28# POR2X1_458/Y -0.00fF
C62111 POR2X1_66/B POR2X1_341/A 0.07fF
C62112 PAND2X1_206/B POR2X1_236/Y 0.10fF
C62113 POR2X1_60/Y POR2X1_20/B 2.13fF
C62114 POR2X1_411/B PAND2X1_354/A 0.03fF
C62115 PAND2X1_41/CTRL POR2X1_330/Y 0.09fF
C62116 PAND2X1_202/CTRL2 POR2X1_69/Y 0.03fF
C62117 POR2X1_585/Y POR2X1_260/B 0.02fF
C62118 PAND2X1_737/B PAND2X1_198/CTRL2 0.01fF
C62119 PAND2X1_659/B POR2X1_329/A 0.03fF
C62120 POR2X1_20/B PAND2X1_541/O 0.04fF
C62121 PAND2X1_264/CTRL2 POR2X1_77/Y 0.01fF
C62122 PAND2X1_628/CTRL2 POR2X1_35/Y 0.01fF
C62123 PAND2X1_20/A POR2X1_454/A 0.12fF
C62124 POR2X1_168/A POR2X1_566/B 0.05fF
C62125 POR2X1_150/Y PAND2X1_736/O 0.02fF
C62126 POR2X1_458/Y PAND2X1_369/O 0.06fF
C62127 POR2X1_76/A POR2X1_330/Y 0.05fF
C62128 PAND2X1_837/O POR2X1_13/A 0.01fF
C62129 PAND2X1_11/Y POR2X1_66/A 0.41fF
C62130 POR2X1_83/B PAND2X1_392/CTRL 0.00fF
C62131 PAND2X1_266/CTRL PAND2X1_215/B 0.01fF
C62132 POR2X1_811/a_16_28# PAND2X1_73/Y 0.02fF
C62133 POR2X1_260/B PAND2X1_13/CTRL2 0.00fF
C62134 POR2X1_604/CTRL POR2X1_236/Y 0.03fF
C62135 POR2X1_99/A PAND2X1_93/B 0.62fF
C62136 POR2X1_78/A POR2X1_608/Y 0.00fF
C62137 POR2X1_834/Y PAND2X1_72/A 0.03fF
C62138 POR2X1_632/CTRL POR2X1_61/Y 0.03fF
C62139 POR2X1_48/A POR2X1_94/A 0.00fF
C62140 POR2X1_48/A PAND2X1_731/B 0.04fF
C62141 D_INPUT_7 PAND2X1_32/B 0.01fF
C62142 PAND2X1_55/Y PAND2X1_45/O 0.03fF
C62143 POR2X1_474/CTRL2 POR2X1_590/A 0.00fF
C62144 POR2X1_373/Y POR2X1_77/Y 0.54fF
C62145 PAND2X1_56/Y POR2X1_260/O 0.02fF
C62146 POR2X1_38/CTRL POR2X1_5/Y 0.00fF
C62147 POR2X1_23/Y PAND2X1_579/O 0.01fF
C62148 POR2X1_68/A PAND2X1_52/CTRL 0.01fF
C62149 POR2X1_490/Y POR2X1_5/Y 0.02fF
C62150 POR2X1_846/A POR2X1_789/CTRL 0.01fF
C62151 PAND2X1_673/a_16_344# POR2X1_672/Y 0.01fF
C62152 POR2X1_302/Y POR2X1_831/a_16_28# 0.02fF
C62153 PAND2X1_458/CTRL2 POR2X1_387/Y 0.06fF
C62154 POR2X1_96/A PAND2X1_796/B 0.03fF
C62155 POR2X1_609/Y PAND2X1_240/CTRL 0.00fF
C62156 POR2X1_607/A POR2X1_102/Y 0.01fF
C62157 POR2X1_416/B PAND2X1_703/O 0.01fF
C62158 PAND2X1_475/CTRL POR2X1_102/Y 0.01fF
C62159 PAND2X1_578/Y VDD 0.17fF
C62160 POR2X1_20/B POR2X1_628/CTRL 0.01fF
C62161 POR2X1_96/A PAND2X1_454/B 0.01fF
C62162 POR2X1_14/Y PAND2X1_453/A 2.69fF
C62163 POR2X1_750/B POR2X1_296/B 0.07fF
C62164 POR2X1_360/A PAND2X1_39/B 0.75fF
C62165 POR2X1_411/B PAND2X1_724/B 0.01fF
C62166 POR2X1_638/Y PAND2X1_53/CTRL 0.04fF
C62167 POR2X1_83/B PAND2X1_169/Y 0.03fF
C62168 POR2X1_567/A POR2X1_736/A 0.07fF
C62169 POR2X1_814/A POR2X1_210/Y 0.03fF
C62170 PAND2X1_657/O POR2X1_72/B 0.20fF
C62171 PAND2X1_458/O POR2X1_283/A 0.01fF
C62172 POR2X1_843/O POR2X1_343/A 0.01fF
C62173 POR2X1_843/CTRL POR2X1_287/B 0.01fF
C62174 PAND2X1_62/O D_INPUT_0 0.04fF
C62175 POR2X1_24/Y POR2X1_7/B 0.05fF
C62176 POR2X1_260/B POR2X1_459/O 0.01fF
C62177 POR2X1_48/A POR2X1_256/CTRL2 0.01fF
C62178 PAND2X1_23/Y POR2X1_294/O 0.01fF
C62179 POR2X1_41/B POR2X1_692/CTRL2 0.01fF
C62180 PAND2X1_65/B POR2X1_448/CTRL2 0.01fF
C62181 POR2X1_841/B POR2X1_284/CTRL2 0.01fF
C62182 PAND2X1_557/A POR2X1_331/Y 0.03fF
C62183 POR2X1_569/a_76_344# POR2X1_174/A 0.01fF
C62184 POR2X1_51/A POR2X1_48/A 0.03fF
C62185 POR2X1_96/A POR2X1_23/Y 0.22fF
C62186 POR2X1_65/A POR2X1_60/A 0.24fF
C62187 D_INPUT_0 INPUT_0 0.17fF
C62188 POR2X1_251/A PAND2X1_540/CTRL 0.01fF
C62189 PAND2X1_438/O POR2X1_456/B 0.04fF
C62190 POR2X1_708/B PAND2X1_93/B 0.02fF
C62191 POR2X1_200/O PAND2X1_41/B 0.01fF
C62192 PAND2X1_550/O POR2X1_32/A 0.01fF
C62193 POR2X1_341/A PAND2X1_316/a_16_344# 0.05fF
C62194 POR2X1_383/A POR2X1_260/O 0.10fF
C62195 POR2X1_97/CTRL2 POR2X1_814/A 0.03fF
C62196 POR2X1_65/A POR2X1_591/A 0.00fF
C62197 POR2X1_833/A PAND2X1_255/CTRL 0.06fF
C62198 PAND2X1_580/CTRL2 PAND2X1_578/Y 0.01fF
C62199 PAND2X1_10/a_16_344# PAND2X1_8/Y 0.06fF
C62200 PAND2X1_679/CTRL2 POR2X1_750/B 0.01fF
C62201 PAND2X1_6/Y POR2X1_624/Y 0.23fF
C62202 PAND2X1_719/Y POR2X1_666/A 0.09fF
C62203 PAND2X1_235/O PAND2X1_85/Y 0.03fF
C62204 POR2X1_66/B PAND2X1_815/O 0.06fF
C62205 PAND2X1_435/Y INPUT_0 0.05fF
C62206 POR2X1_41/B POR2X1_484/O 0.02fF
C62207 POR2X1_366/Y POR2X1_270/Y 0.95fF
C62208 POR2X1_23/Y PAND2X1_445/CTRL2 0.30fF
C62209 POR2X1_83/B PAND2X1_730/B 0.03fF
C62210 POR2X1_632/CTRL POR2X1_35/Y 0.01fF
C62211 POR2X1_750/B PAND2X1_526/a_16_344# 0.01fF
C62212 D_INPUT_5 PAND2X1_69/A 0.03fF
C62213 PAND2X1_404/A PAND2X1_404/O 0.02fF
C62214 POR2X1_647/B POR2X1_649/CTRL 0.01fF
C62215 PAND2X1_30/O PAND2X1_3/B 0.04fF
C62216 PAND2X1_771/Y PAND2X1_552/B 0.05fF
C62217 POR2X1_139/a_16_28# POR2X1_624/Y 0.03fF
C62218 POR2X1_324/B PAND2X1_320/CTRL 0.01fF
C62219 PAND2X1_77/a_76_28# PAND2X1_8/Y 0.01fF
C62220 POR2X1_260/B POR2X1_816/A 0.03fF
C62221 POR2X1_842/O POR2X1_741/Y 0.02fF
C62222 POR2X1_697/O POR2X1_72/B 0.01fF
C62223 POR2X1_462/B POR2X1_260/B 0.03fF
C62224 PAND2X1_733/CTRL PAND2X1_723/Y 0.02fF
C62225 PAND2X1_860/A PAND2X1_865/A 0.01fF
C62226 POR2X1_311/Y PAND2X1_137/Y 0.03fF
C62227 INPUT_3 POR2X1_380/Y -0.02fF
C62228 PAND2X1_471/a_16_344# POR2X1_83/B 0.02fF
C62229 POR2X1_260/B D_INPUT_1 0.06fF
C62230 POR2X1_343/Y PAND2X1_52/B 0.00fF
C62231 PAND2X1_472/B POR2X1_14/Y 0.49fF
C62232 POR2X1_791/Y POR2X1_637/B 0.01fF
C62233 POR2X1_796/Y PAND2X1_69/A 0.03fF
C62234 POR2X1_96/A PAND2X1_221/O 0.04fF
C62235 POR2X1_360/A PAND2X1_20/A 0.12fF
C62236 POR2X1_48/Y POR2X1_32/A 0.01fF
C62237 PAND2X1_71/a_16_344# POR2X1_296/B 0.01fF
C62238 POR2X1_68/CTRL2 POR2X1_402/A 0.01fF
C62239 POR2X1_814/A PAND2X1_310/CTRL 0.09fF
C62240 POR2X1_52/A POR2X1_421/Y 0.12fF
C62241 PAND2X1_319/B PAND2X1_212/CTRL 0.03fF
C62242 PAND2X1_56/Y POR2X1_842/a_16_28# 0.06fF
C62243 PAND2X1_41/B VDD 3.30fF
C62244 POR2X1_783/A POR2X1_783/O 0.03fF
C62245 POR2X1_447/a_16_28# POR2X1_447/A 0.00fF
C62246 POR2X1_260/B POR2X1_724/A 0.03fF
C62247 PAND2X1_652/A POR2X1_32/A 0.12fF
C62248 PAND2X1_6/Y PAND2X1_689/CTRL2 0.00fF
C62249 POR2X1_448/O POR2X1_294/B 0.03fF
C62250 POR2X1_14/Y POR2X1_55/Y 3.30fF
C62251 PAND2X1_137/Y PAND2X1_140/CTRL2 0.03fF
C62252 PAND2X1_220/CTRL POR2X1_83/B 0.01fF
C62253 POR2X1_503/CTRL POR2X1_411/B 0.10fF
C62254 PAND2X1_220/A PAND2X1_566/Y 0.02fF
C62255 POR2X1_760/A PAND2X1_853/B 0.07fF
C62256 PAND2X1_362/A PAND2X1_354/CTRL2 0.01fF
C62257 POR2X1_856/B POR2X1_788/B 0.02fF
C62258 POR2X1_48/A PAND2X1_113/O 0.08fF
C62259 POR2X1_781/A VDD -0.00fF
C62260 POR2X1_404/CTRL2 POR2X1_404/Y 0.01fF
C62261 POR2X1_356/A POR2X1_439/O 0.03fF
C62262 PAND2X1_90/Y INPUT_0 0.08fF
C62263 POR2X1_43/B POR2X1_420/Y 0.03fF
C62264 POR2X1_98/B POR2X1_66/A 0.01fF
C62265 PAND2X1_798/B PAND2X1_78/CTRL 0.01fF
C62266 POR2X1_60/A PAND2X1_190/Y 0.12fF
C62267 POR2X1_661/O POR2X1_722/Y 0.00fF
C62268 PAND2X1_20/A POR2X1_713/O 0.01fF
C62269 POR2X1_119/Y PAND2X1_266/CTRL 0.13fF
C62270 POR2X1_360/A POR2X1_814/B 0.39fF
C62271 POR2X1_261/A VDD 0.00fF
C62272 D_INPUT_0 POR2X1_780/A 0.48fF
C62273 PAND2X1_180/CTRL PAND2X1_182/A 0.00fF
C62274 POR2X1_630/A D_GATE_222 0.03fF
C62275 PAND2X1_660/CTRL2 POR2X1_413/A 0.01fF
C62276 POR2X1_660/CTRL POR2X1_840/B 0.14fF
C62277 POR2X1_68/A POR2X1_244/CTRL2 0.10fF
C62278 POR2X1_346/B PAND2X1_60/O 0.00fF
C62279 POR2X1_23/Y POR2X1_7/A 1.61fF
C62280 POR2X1_448/Y POR2X1_802/B 0.07fF
C62281 POR2X1_669/B PAND2X1_645/B 0.03fF
C62282 POR2X1_825/a_16_28# POR2X1_42/Y 0.03fF
C62283 POR2X1_402/B VDD 0.15fF
C62284 PAND2X1_204/O POR2X1_79/Y 0.02fF
C62285 POR2X1_805/Y POR2X1_758/CTRL2 0.01fF
C62286 POR2X1_66/B POR2X1_460/a_76_344# 0.01fF
C62287 PAND2X1_248/CTRL POR2X1_101/Y 0.03fF
C62288 PAND2X1_23/Y POR2X1_343/A 0.06fF
C62289 PAND2X1_90/A PAND2X1_42/O 0.05fF
C62290 POR2X1_814/B POR2X1_756/O 0.04fF
C62291 POR2X1_702/B POR2X1_205/Y 0.06fF
C62292 POR2X1_41/B PAND2X1_473/B 0.08fF
C62293 PAND2X1_96/B POR2X1_285/Y 0.03fF
C62294 PAND2X1_230/CTRL PAND2X1_32/B 0.01fF
C62295 POR2X1_806/O POR2X1_804/A 0.17fF
C62296 PAND2X1_243/B POR2X1_5/Y 0.02fF
C62297 PAND2X1_474/a_16_344# POR2X1_153/Y 0.02fF
C62298 POR2X1_16/A PAND2X1_443/O 0.04fF
C62299 POR2X1_702/B PAND2X1_55/Y 0.01fF
C62300 PAND2X1_41/B POR2X1_741/Y 0.05fF
C62301 POR2X1_866/CTRL PAND2X1_32/B 0.01fF
C62302 POR2X1_333/A POR2X1_577/CTRL 0.01fF
C62303 POR2X1_66/B PAND2X1_767/O 0.04fF
C62304 POR2X1_122/Y POR2X1_293/Y 0.01fF
C62305 POR2X1_41/CTRL PAND2X1_852/A 0.01fF
C62306 PAND2X1_39/B POR2X1_579/B 0.12fF
C62307 PAND2X1_48/B POR2X1_778/CTRL2 0.02fF
C62308 PAND2X1_284/a_56_28# POR2X1_279/Y 0.00fF
C62309 POR2X1_16/A PAND2X1_124/Y 0.09fF
C62310 PAND2X1_576/O POR2X1_599/A 0.02fF
C62311 PAND2X1_653/Y PAND2X1_557/A 0.01fF
C62312 POR2X1_114/B POR2X1_862/B 0.05fF
C62313 POR2X1_113/Y POR2X1_390/CTRL2 0.05fF
C62314 POR2X1_257/A PAND2X1_156/A 0.12fF
C62315 PAND2X1_592/Y VDD 0.50fF
C62316 PAND2X1_412/O POR2X1_391/Y 0.02fF
C62317 PAND2X1_702/CTRL POR2X1_40/Y 0.00fF
C62318 POR2X1_27/Y POR2X1_38/Y 1.01fF
C62319 PAND2X1_421/a_56_28# PAND2X1_90/Y 0.00fF
C62320 PAND2X1_41/B PAND2X1_32/B 0.82fF
C62321 PAND2X1_455/Y PAND2X1_465/B 0.14fF
C62322 POR2X1_57/A POR2X1_40/Y 65.54fF
C62323 PAND2X1_635/CTRL INPUT_7 0.00fF
C62324 POR2X1_192/Y POR2X1_579/Y 0.03fF
C62325 POR2X1_135/CTRL2 POR2X1_257/A 0.01fF
C62326 PAND2X1_63/Y PAND2X1_262/O 0.00fF
C62327 POR2X1_40/O POR2X1_32/A 0.01fF
C62328 PAND2X1_433/a_76_28# PAND2X1_65/B 0.02fF
C62329 POR2X1_52/A INPUT_5 0.16fF
C62330 POR2X1_273/Y POR2X1_272/Y 0.28fF
C62331 POR2X1_130/Y VDD 0.26fF
C62332 PAND2X1_41/B POR2X1_711/O 0.01fF
C62333 PAND2X1_48/B POR2X1_121/Y 0.00fF
C62334 PAND2X1_57/B POR2X1_733/A 0.15fF
C62335 POR2X1_119/Y PAND2X1_203/a_76_28# 0.03fF
C62336 POR2X1_56/B POR2X1_372/Y 0.10fF
C62337 POR2X1_334/B PAND2X1_57/B 0.05fF
C62338 PAND2X1_411/m4_208_n4# PAND2X1_90/Y 0.06fF
C62339 POR2X1_502/A POR2X1_732/B 0.03fF
C62340 POR2X1_448/Y POR2X1_532/A 0.03fF
C62341 POR2X1_220/Y POR2X1_803/A 0.03fF
C62342 PAND2X1_69/A PAND2X1_396/m4_208_n4# 0.15fF
C62343 POR2X1_791/B POR2X1_637/B 0.03fF
C62344 POR2X1_113/Y POR2X1_654/B 0.01fF
C62345 POR2X1_186/Y PAND2X1_60/B 0.07fF
C62346 POR2X1_13/A POR2X1_599/A 0.02fF
C62347 POR2X1_192/Y POR2X1_545/A 0.58fF
C62348 POR2X1_390/CTRL2 POR2X1_260/A 0.00fF
C62349 POR2X1_65/A PAND2X1_113/a_76_28# 0.01fF
C62350 POR2X1_16/A POR2X1_83/B 1.55fF
C62351 PAND2X1_72/CTRL VDD 0.00fF
C62352 POR2X1_278/Y PAND2X1_357/Y 0.03fF
C62353 POR2X1_10/a_16_28# POR2X1_669/B 0.02fF
C62354 POR2X1_37/Y PAND2X1_508/Y 0.03fF
C62355 PAND2X1_824/B POR2X1_632/B 0.04fF
C62356 POR2X1_526/Y POR2X1_692/Y 0.07fF
C62357 POR2X1_614/A POR2X1_192/Y 0.02fF
C62358 POR2X1_113/CTRL PAND2X1_65/B 0.01fF
C62359 POR2X1_763/Y PAND2X1_726/O 0.09fF
C62360 PAND2X1_691/Y POR2X1_829/a_76_344# 0.01fF
C62361 POR2X1_866/A POR2X1_691/A 0.05fF
C62362 PAND2X1_592/Y PAND2X1_850/CTRL 0.01fF
C62363 POR2X1_210/a_16_28# POR2X1_210/B 0.07fF
C62364 POR2X1_124/B PAND2X1_57/B 0.00fF
C62365 PAND2X1_635/CTRL INPUT_4 0.01fF
C62366 PAND2X1_202/O D_INPUT_1 0.14fF
C62367 VDD PAND2X1_314/CTRL 0.00fF
C62368 POR2X1_532/A POR2X1_215/CTRL2 0.01fF
C62369 PAND2X1_94/A PAND2X1_23/CTRL2 0.01fF
C62370 POR2X1_728/B PAND2X1_69/A 0.01fF
C62371 INPUT_1 PAND2X1_73/O 0.04fF
C62372 POR2X1_824/Y POR2X1_236/Y 0.01fF
C62373 PAND2X1_76/Y PAND2X1_349/A 0.03fF
C62374 POR2X1_624/Y POR2X1_632/Y 0.00fF
C62375 VDD POR2X1_714/CTRL 0.00fF
C62376 PAND2X1_620/a_76_28# POR2X1_422/Y 0.02fF
C62377 POR2X1_664/Y POR2X1_712/Y 0.03fF
C62378 PAND2X1_48/B POR2X1_723/B 0.03fF
C62379 PAND2X1_785/CTRL2 POR2X1_7/B 0.00fF
C62380 PAND2X1_824/B POR2X1_631/O 0.06fF
C62381 PAND2X1_474/A POR2X1_171/O 0.16fF
C62382 POR2X1_283/A POR2X1_511/Y 0.03fF
C62383 POR2X1_502/A POR2X1_578/CTRL2 0.01fF
C62384 PAND2X1_6/Y POR2X1_785/A 0.18fF
C62385 PAND2X1_73/Y PAND2X1_48/A 0.32fF
C62386 POR2X1_52/A PAND2X1_186/CTRL2 0.00fF
C62387 POR2X1_65/A POR2X1_744/CTRL 0.01fF
C62388 VDD POR2X1_228/Y 3.49fF
C62389 POR2X1_20/B PAND2X1_351/A 0.01fF
C62390 PAND2X1_839/B VDD 0.04fF
C62391 VDD PAND2X1_348/Y 0.96fF
C62392 D_GATE_222 POR2X1_795/B 0.07fF
C62393 POR2X1_532/A POR2X1_794/a_16_28# 0.02fF
C62394 POR2X1_186/Y POR2X1_353/A 0.71fF
C62395 POR2X1_197/Y POR2X1_243/Y 0.04fF
C62396 PAND2X1_808/Y PAND2X1_773/CTRL2 0.01fF
C62397 POR2X1_32/A PAND2X1_506/Y 0.05fF
C62398 POR2X1_550/A VDD 0.25fF
C62399 PAND2X1_55/Y D_INPUT_1 0.09fF
C62400 POR2X1_49/Y PAND2X1_844/CTRL2 0.00fF
C62401 PAND2X1_785/Y POR2X1_387/Y 0.03fF
C62402 PAND2X1_754/m4_208_n4# PAND2X1_69/A 0.15fF
C62403 POR2X1_787/CTRL2 POR2X1_325/A 0.01fF
C62404 POR2X1_326/A POR2X1_436/CTRL2 0.00fF
C62405 POR2X1_327/Y POR2X1_141/Y 0.00fF
C62406 PAND2X1_562/O PAND2X1_566/Y 0.14fF
C62407 POR2X1_720/B POR2X1_790/A 0.44fF
C62408 POR2X1_624/Y PAND2X1_52/B 0.05fF
C62409 PAND2X1_20/A POR2X1_571/Y 0.04fF
C62410 POR2X1_83/B PAND2X1_336/Y 0.90fF
C62411 POR2X1_502/A PAND2X1_306/a_76_28# 0.02fF
C62412 PAND2X1_215/CTRL POR2X1_7/Y 0.01fF
C62413 POR2X1_370/Y PAND2X1_368/CTRL 0.01fF
C62414 POR2X1_447/B POR2X1_629/B 0.06fF
C62415 POR2X1_334/Y PAND2X1_7/Y 0.03fF
C62416 POR2X1_66/B POR2X1_735/O 0.03fF
C62417 PAND2X1_55/Y POR2X1_724/A 0.07fF
C62418 POR2X1_244/B POR2X1_259/CTRL2 0.01fF
C62419 POR2X1_765/CTRL POR2X1_73/Y 0.08fF
C62420 PAND2X1_661/B POR2X1_599/A 0.04fF
C62421 PAND2X1_852/CTRL POR2X1_821/Y 0.00fF
C62422 POR2X1_675/CTRL2 POR2X1_188/Y 0.01fF
C62423 POR2X1_346/B POR2X1_206/A 0.02fF
C62424 POR2X1_99/B PAND2X1_20/A 0.01fF
C62425 PAND2X1_63/Y PAND2X1_316/CTRL 0.04fF
C62426 POR2X1_38/B POR2X1_382/O 0.01fF
C62427 PAND2X1_317/Y POR2X1_258/a_16_28# 0.03fF
C62428 PAND2X1_390/Y PAND2X1_851/CTRL2 0.01fF
C62429 POR2X1_156/B POR2X1_68/A 0.14fF
C62430 POR2X1_49/Y PAND2X1_156/A 0.10fF
C62431 POR2X1_62/Y POR2X1_94/A 0.07fF
C62432 POR2X1_810/CTRL2 POR2X1_809/Y 0.01fF
C62433 PAND2X1_550/B PAND2X1_549/a_16_344# 0.01fF
C62434 PAND2X1_56/Y POR2X1_702/CTRL2 0.13fF
C62435 PAND2X1_566/Y PAND2X1_347/O 0.19fF
C62436 POR2X1_416/B POR2X1_626/CTRL2 0.01fF
C62437 D_INPUT_0 POR2X1_522/CTRL2 0.06fF
C62438 POR2X1_72/B POR2X1_385/Y 0.37fF
C62439 POR2X1_356/A PAND2X1_315/O 0.06fF
C62440 PAND2X1_385/a_16_344# PAND2X1_60/B 0.02fF
C62441 PAND2X1_215/B PAND2X1_717/Y 0.07fF
C62442 POR2X1_38/B PAND2X1_29/O 0.06fF
C62443 PAND2X1_793/Y PAND2X1_574/O 0.02fF
C62444 PAND2X1_553/B PAND2X1_114/CTRL2 0.05fF
C62445 POR2X1_322/CTRL2 PAND2X1_569/B 0.01fF
C62446 POR2X1_741/Y POR2X1_228/Y 0.03fF
C62447 POR2X1_578/Y POR2X1_577/Y 0.00fF
C62448 POR2X1_7/B PAND2X1_336/CTRL2 0.00fF
C62449 POR2X1_121/A PAND2X1_60/B 0.01fF
C62450 PAND2X1_403/O POR2X1_20/B 0.16fF
C62451 PAND2X1_118/CTRL2 POR2X1_123/A 0.01fF
C62452 POR2X1_81/A PAND2X1_244/O 0.12fF
C62453 POR2X1_300/O PAND2X1_349/A 0.01fF
C62454 POR2X1_503/CTRL POR2X1_52/A 0.01fF
C62455 POR2X1_7/B PAND2X1_155/O 0.01fF
C62456 PAND2X1_284/CTRL POR2X1_258/Y 0.01fF
C62457 POR2X1_101/Y POR2X1_294/B 0.03fF
C62458 PAND2X1_81/O POR2X1_84/Y 0.03fF
C62459 POR2X1_166/CTRL POR2X1_73/Y 0.01fF
C62460 POR2X1_383/A D_GATE_222 0.07fF
C62461 PAND2X1_689/CTRL2 PAND2X1_52/B 0.02fF
C62462 POR2X1_41/CTRL2 POR2X1_42/Y 0.01fF
C62463 POR2X1_634/A D_INPUT_4 0.05fF
C62464 PAND2X1_365/B PAND2X1_854/A 0.02fF
C62465 POR2X1_297/Y PAND2X1_359/Y 0.04fF
C62466 PAND2X1_90/A INPUT_1 0.22fF
C62467 POR2X1_327/Y POR2X1_220/Y 0.10fF
C62468 POR2X1_477/A POR2X1_456/B 0.03fF
C62469 PAND2X1_65/B POR2X1_540/Y 0.02fF
C62470 POR2X1_228/Y PAND2X1_32/B 0.02fF
C62471 POR2X1_13/A POR2X1_599/O 0.17fF
C62472 POR2X1_55/Y PAND2X1_508/O 0.05fF
C62473 PAND2X1_182/B POR2X1_7/B 0.03fF
C62474 PAND2X1_383/a_16_344# POR2X1_90/Y 0.02fF
C62475 POR2X1_355/B POR2X1_209/O 0.01fF
C62476 POR2X1_100/a_56_344# PAND2X1_88/Y 0.00fF
C62477 POR2X1_364/A POR2X1_169/Y 0.10fF
C62478 PAND2X1_805/A PAND2X1_367/a_16_344# 0.02fF
C62479 POR2X1_706/B PAND2X1_692/m4_208_n4# 0.03fF
C62480 POR2X1_564/Y POR2X1_564/B 0.07fF
C62481 POR2X1_417/CTRL2 POR2X1_283/A 0.03fF
C62482 POR2X1_38/Y PAND2X1_194/O 0.01fF
C62483 PAND2X1_83/O PAND2X1_82/Y 0.03fF
C62484 POR2X1_731/O POR2X1_854/B 0.01fF
C62485 POR2X1_327/Y POR2X1_404/Y 0.03fF
C62486 POR2X1_203/CTRL PAND2X1_111/B 0.01fF
C62487 POR2X1_795/CTRL2 POR2X1_186/B 0.01fF
C62488 POR2X1_318/A POR2X1_140/a_16_28# 0.07fF
C62489 POR2X1_41/B POR2X1_131/A 0.01fF
C62490 POR2X1_3/B INPUT_5 0.00fF
C62491 POR2X1_541/O POR2X1_366/A 0.01fF
C62492 PAND2X1_684/CTRL2 POR2X1_149/B 0.01fF
C62493 PAND2X1_422/CTRL2 PAND2X1_60/B 0.00fF
C62494 PAND2X1_569/B POR2X1_90/Y 0.08fF
C62495 PAND2X1_476/A VDD 0.89fF
C62496 POR2X1_9/Y PAND2X1_66/CTRL2 0.03fF
C62497 PAND2X1_508/Y POR2X1_293/Y 0.03fF
C62498 POR2X1_349/O PAND2X1_57/B 0.01fF
C62499 PAND2X1_224/CTRL2 POR2X1_191/Y 0.22fF
C62500 PAND2X1_141/a_76_28# POR2X1_39/B 0.02fF
C62501 INPUT_0 PAND2X1_643/A 0.04fF
C62502 POR2X1_596/A POR2X1_796/A 0.03fF
C62503 POR2X1_705/CTRL POR2X1_260/A 0.01fF
C62504 INPUT_1 POR2X1_248/CTRL 0.01fF
C62505 POR2X1_553/A POR2X1_573/A 0.00fF
C62506 PAND2X1_840/B POR2X1_153/Y 0.04fF
C62507 PAND2X1_481/O D_GATE_741 0.07fF
C62508 POR2X1_300/CTRL POR2X1_300/Y 0.01fF
C62509 VDD PAND2X1_122/O 0.00fF
C62510 POR2X1_222/A POR2X1_510/Y 0.03fF
C62511 POR2X1_532/A PAND2X1_133/O 0.02fF
C62512 POR2X1_345/O PAND2X1_6/Y 0.17fF
C62513 POR2X1_135/CTRL2 PAND2X1_553/B 0.01fF
C62514 POR2X1_722/B POR2X1_722/O 0.01fF
C62515 PAND2X1_584/CTRL PAND2X1_52/B 0.01fF
C62516 PAND2X1_23/Y PAND2X1_18/B 0.03fF
C62517 POR2X1_260/m4_208_n4# PAND2X1_45/m4_208_n4# 0.13fF
C62518 POR2X1_786/Y POR2X1_244/Y 0.07fF
C62519 POR2X1_350/B POR2X1_351/O 0.05fF
C62520 POR2X1_52/A POR2X1_824/O 0.02fF
C62521 VDD POR2X1_769/B 0.09fF
C62522 PAND2X1_833/CTRL POR2X1_39/B 0.01fF
C62523 PAND2X1_510/O POR2X1_73/Y 0.17fF
C62524 POR2X1_294/B POR2X1_722/O 0.01fF
C62525 PAND2X1_218/A PAND2X1_853/B 0.05fF
C62526 POR2X1_566/A PAND2X1_179/CTRL 0.03fF
C62527 POR2X1_101/Y PAND2X1_111/B 0.05fF
C62528 PAND2X1_72/Y POR2X1_203/Y 0.04fF
C62529 POR2X1_554/B POR2X1_276/B 0.03fF
C62530 PAND2X1_6/Y POR2X1_186/B 0.10fF
C62531 POR2X1_248/CTRL POR2X1_153/Y 0.28fF
C62532 POR2X1_513/B PAND2X1_304/CTRL 0.00fF
C62533 POR2X1_777/B POR2X1_343/B 0.05fF
C62534 PAND2X1_357/Y PAND2X1_357/O 0.03fF
C62535 PAND2X1_865/O PAND2X1_175/B 0.01fF
C62536 POR2X1_732/B POR2X1_188/Y 0.05fF
C62537 POR2X1_378/A PAND2X1_94/A 0.01fF
C62538 PAND2X1_661/B POR2X1_599/O 0.01fF
C62539 PAND2X1_437/a_16_344# POR2X1_174/A 0.03fF
C62540 POR2X1_38/Y PAND2X1_853/B 0.03fF
C62541 POR2X1_550/A POR2X1_673/Y 0.07fF
C62542 POR2X1_7/B POR2X1_767/Y 0.09fF
C62543 PAND2X1_678/a_16_344# POR2X1_257/A 0.02fF
C62544 PAND2X1_865/Y POR2X1_45/Y 0.03fF
C62545 PAND2X1_348/A POR2X1_387/Y 0.10fF
C62546 POR2X1_383/A POR2X1_561/a_16_28# 0.01fF
C62547 PAND2X1_90/CTRL D_INPUT_1 0.04fF
C62548 PAND2X1_470/CTRL2 POR2X1_119/Y 0.00fF
C62549 POR2X1_3/A POR2X1_762/CTRL 0.01fF
C62550 PAND2X1_778/Y PAND2X1_156/A 0.05fF
C62551 PAND2X1_651/Y PAND2X1_506/Y 0.02fF
C62552 POR2X1_760/A POR2X1_23/Y 0.01fF
C62553 POR2X1_775/O POR2X1_191/Y -0.01fF
C62554 PAND2X1_607/CTRL POR2X1_606/Y 0.01fF
C62555 PAND2X1_732/A PAND2X1_569/B 0.07fF
C62556 POR2X1_137/B POR2X1_260/B 0.46fF
C62557 POR2X1_83/Y POR2X1_73/Y 0.02fF
C62558 POR2X1_283/A POR2X1_129/Y 0.09fF
C62559 POR2X1_461/Y POR2X1_862/A 0.01fF
C62560 PAND2X1_373/CTRL POR2X1_544/B 0.01fF
C62561 POR2X1_576/O POR2X1_260/A 0.01fF
C62562 POR2X1_673/Y POR2X1_721/CTRL 0.02fF
C62563 POR2X1_499/A POR2X1_558/B 1.88fF
C62564 INPUT_3 POR2X1_260/B 0.06fF
C62565 POR2X1_244/Y POR2X1_575/m4_208_n4# 0.09fF
C62566 POR2X1_705/B POR2X1_66/A 0.03fF
C62567 POR2X1_245/a_16_28# PAND2X1_156/A 0.02fF
C62568 POR2X1_318/m4_208_n4# POR2X1_454/m4_208_n4# 0.13fF
C62569 PAND2X1_27/CTRL POR2X1_294/A 0.01fF
C62570 POR2X1_446/B POR2X1_446/O 0.04fF
C62571 POR2X1_785/A PAND2X1_52/B 0.03fF
C62572 PAND2X1_816/O PAND2X1_52/B 0.02fF
C62573 POR2X1_635/B VDD 0.21fF
C62574 POR2X1_48/A PAND2X1_415/CTRL 0.01fF
C62575 PAND2X1_448/a_16_344# POR2X1_20/B 0.01fF
C62576 POR2X1_485/m4_208_n4# POR2X1_236/Y 0.07fF
C62577 POR2X1_416/B PAND2X1_547/CTRL 0.02fF
C62578 POR2X1_368/Y POR2X1_416/B 0.00fF
C62579 POR2X1_154/m4_208_n4# PAND2X1_72/A 0.15fF
C62580 POR2X1_648/O D_INPUT_0 0.08fF
C62581 PAND2X1_73/Y POR2X1_461/Y 0.03fF
C62582 POR2X1_452/Y POR2X1_801/B 0.02fF
C62583 PAND2X1_93/B POR2X1_260/B 0.11fF
C62584 POR2X1_514/Y POR2X1_138/A 0.01fF
C62585 POR2X1_276/Y POR2X1_362/O 0.01fF
C62586 POR2X1_172/Y POR2X1_39/B 0.04fF
C62587 POR2X1_54/Y POR2X1_55/O 0.01fF
C62588 POR2X1_99/A POR2X1_99/CTRL2 0.01fF
C62589 POR2X1_329/A POR2X1_5/Y 0.08fF
C62590 POR2X1_350/Y POR2X1_568/A 0.01fF
C62591 POR2X1_411/B PAND2X1_733/A 0.00fF
C62592 POR2X1_65/A POR2X1_329/Y 0.05fF
C62593 POR2X1_490/CTRL POR2X1_40/Y 0.01fF
C62594 POR2X1_313/CTRL POR2X1_167/Y 0.01fF
C62595 POR2X1_250/Y PAND2X1_347/Y 0.11fF
C62596 POR2X1_661/A PAND2X1_385/O 0.07fF
C62597 POR2X1_477/CTRL POR2X1_186/Y 0.14fF
C62598 POR2X1_493/CTRL2 PAND2X1_72/A 0.00fF
C62599 POR2X1_864/A POR2X1_774/Y 0.04fF
C62600 POR2X1_78/A POR2X1_260/B 2.51fF
C62601 POR2X1_477/Y POR2X1_220/B 0.01fF
C62602 PAND2X1_9/Y PAND2X1_41/B 0.03fF
C62603 POR2X1_856/B POR2X1_436/B 1.26fF
C62604 PAND2X1_717/A PAND2X1_151/a_16_344# 0.02fF
C62605 PAND2X1_60/B POR2X1_717/B 0.03fF
C62606 POR2X1_472/B POR2X1_734/A -0.01fF
C62607 POR2X1_485/Y POR2X1_692/Y 0.10fF
C62608 PAND2X1_497/O POR2X1_267/A 0.05fF
C62609 POR2X1_416/B PAND2X1_155/CTRL 0.01fF
C62610 PAND2X1_793/Y PAND2X1_717/A 0.03fF
C62611 POR2X1_394/A PAND2X1_379/O 0.09fF
C62612 POR2X1_635/B PAND2X1_32/B 0.01fF
C62613 POR2X1_842/CTRL POR2X1_850/B 0.01fF
C62614 PAND2X1_72/A PAND2X1_315/O 0.04fF
C62615 POR2X1_263/CTRL VDD 0.00fF
C62616 POR2X1_49/Y PAND2X1_443/CTRL 0.00fF
C62617 POR2X1_83/B PAND2X1_214/O 0.04fF
C62618 PAND2X1_246/a_76_28# INPUT_0 0.02fF
C62619 POR2X1_62/Y POR2X1_150/a_16_28# 0.10fF
C62620 POR2X1_102/Y D_INPUT_0 0.18fF
C62621 POR2X1_816/O INPUT_0 -0.00fF
C62622 PAND2X1_694/CTRL2 PAND2X1_425/Y 0.03fF
C62623 POR2X1_657/Y VDD 0.22fF
C62624 POR2X1_390/B PAND2X1_72/A 0.03fF
C62625 POR2X1_632/Y POR2X1_186/B 0.03fF
C62626 PAND2X1_464/B POR2X1_293/Y 0.02fF
C62627 POR2X1_648/O PAND2X1_90/Y 0.09fF
C62628 PAND2X1_652/CTRL POR2X1_385/Y 0.00fF
C62629 POR2X1_445/A PAND2X1_65/B 0.03fF
C62630 PAND2X1_414/CTRL POR2X1_42/Y 0.26fF
C62631 POR2X1_20/B PAND2X1_151/O 0.15fF
C62632 PAND2X1_213/Y PAND2X1_147/O 0.02fF
C62633 POR2X1_110/Y POR2X1_316/Y 0.03fF
C62634 POR2X1_634/a_56_344# POR2X1_66/A 0.00fF
C62635 POR2X1_814/A POR2X1_790/B 0.06fF
C62636 POR2X1_411/B PAND2X1_804/B 0.03fF
C62637 POR2X1_241/O POR2X1_241/B 0.01fF
C62638 PAND2X1_226/O POR2X1_227/A 0.00fF
C62639 PAND2X1_493/a_76_28# POR2X1_491/Y 0.05fF
C62640 POR2X1_78/B POR2X1_602/O 0.35fF
C62641 POR2X1_846/Y POR2X1_790/B 0.00fF
C62642 POR2X1_454/A VDD 0.48fF
C62643 PAND2X1_436/A PAND2X1_435/Y 0.07fF
C62644 PAND2X1_46/O POR2X1_296/B 0.00fF
C62645 PAND2X1_736/A POR2X1_150/Y 0.27fF
C62646 POR2X1_850/A POR2X1_656/CTRL2 0.08fF
C62647 POR2X1_728/a_16_28# POR2X1_452/Y 0.03fF
C62648 PAND2X1_207/CTRL VDD 0.00fF
C62649 POR2X1_9/Y POR2X1_245/Y 0.04fF
C62650 POR2X1_863/A POR2X1_703/Y 0.03fF
C62651 PAND2X1_48/B PAND2X1_268/CTRL2 0.01fF
C62652 PAND2X1_807/B PAND2X1_354/A 0.03fF
C62653 POR2X1_427/a_16_28# POR2X1_72/B 0.02fF
C62654 POR2X1_652/A PAND2X1_72/A 0.10fF
C62655 POR2X1_664/O POR2X1_651/Y 0.01fF
C62656 PAND2X1_865/Y PAND2X1_440/CTRL 0.01fF
C62657 POR2X1_376/B POR2X1_496/Y 0.10fF
C62658 POR2X1_518/CTRL POR2X1_77/Y 0.01fF
C62659 POR2X1_439/Y POR2X1_590/A 0.03fF
C62660 POR2X1_864/CTRL2 POR2X1_750/B 0.01fF
C62661 POR2X1_267/A PAND2X1_41/B 0.07fF
C62662 PAND2X1_638/B POR2X1_585/CTRL 0.01fF
C62663 POR2X1_586/Y POR2X1_585/O 0.02fF
C62664 POR2X1_48/A PAND2X1_818/CTRL 0.01fF
C62665 PAND2X1_76/Y POR2X1_32/A 0.03fF
C62666 POR2X1_376/Y POR2X1_29/A 0.17fF
C62667 POR2X1_63/Y POR2X1_43/B 0.05fF
C62668 POR2X1_760/Y POR2X1_416/B 0.01fF
C62669 PAND2X1_392/a_16_344# POR2X1_236/Y 0.01fF
C62670 POR2X1_689/CTRL POR2X1_32/A 0.01fF
C62671 POR2X1_116/A POR2X1_804/A 0.03fF
C62672 POR2X1_260/B PAND2X1_132/CTRL 0.01fF
C62673 POR2X1_692/CTRL POR2X1_46/Y 0.01fF
C62674 POR2X1_254/A POR2X1_186/Y 0.05fF
C62675 PAND2X1_400/O VDD 0.00fF
C62676 POR2X1_68/A POR2X1_471/A 0.03fF
C62677 PAND2X1_256/CTRL POR2X1_205/A 0.06fF
C62678 PAND2X1_242/Y PAND2X1_508/Y 0.05fF
C62679 POR2X1_705/B POR2X1_532/A 0.05fF
C62680 POR2X1_502/A POR2X1_466/A 0.03fF
C62681 POR2X1_540/Y PAND2X1_178/CTRL2 0.01fF
C62682 POR2X1_186/Y POR2X1_750/B 0.03fF
C62683 POR2X1_556/A POR2X1_68/B 0.03fF
C62684 PAND2X1_48/B PAND2X1_248/O 0.02fF
C62685 POR2X1_14/Y POR2X1_511/Y 0.03fF
C62686 PAND2X1_93/B POR2X1_205/Y 0.09fF
C62687 POR2X1_614/A POR2X1_841/a_16_28# 0.03fF
C62688 PAND2X1_93/B PAND2X1_55/Y 0.19fF
C62689 PAND2X1_276/CTRL POR2X1_271/Y 0.02fF
C62690 PAND2X1_675/a_16_344# POR2X1_416/B 0.02fF
C62691 POR2X1_66/A PAND2X1_385/CTRL2 0.01fF
C62692 POR2X1_859/A POR2X1_29/A 0.03fF
C62693 POR2X1_825/Y POR2X1_397/CTRL2 0.00fF
C62694 PAND2X1_766/CTRL2 PAND2X1_90/Y 0.04fF
C62695 POR2X1_417/Y PAND2X1_76/Y 0.02fF
C62696 POR2X1_192/Y POR2X1_590/A 0.09fF
C62697 POR2X1_99/A PAND2X1_65/Y 0.03fF
C62698 PAND2X1_863/B POR2X1_32/A 0.01fF
C62699 POR2X1_484/CTRL POR2X1_763/Y 0.08fF
C62700 POR2X1_347/B POR2X1_296/B 0.09fF
C62701 POR2X1_348/A POR2X1_244/a_16_28# 0.05fF
C62702 POR2X1_341/A POR2X1_541/a_56_344# 0.01fF
C62703 PAND2X1_48/B PAND2X1_282/CTRL2 0.09fF
C62704 POR2X1_65/A GATE_479 0.03fF
C62705 POR2X1_52/A POR2X1_496/Y 0.07fF
C62706 POR2X1_43/m4_208_n4# POR2X1_77/Y 0.07fF
C62707 PAND2X1_93/B POR2X1_788/Y 0.01fF
C62708 POR2X1_93/A POR2X1_628/Y 0.03fF
C62709 POR2X1_854/CTRL2 POR2X1_776/A 0.01fF
C62710 POR2X1_294/Y POR2X1_740/Y 0.05fF
C62711 POR2X1_295/CTRL POR2X1_481/A 0.01fF
C62712 POR2X1_634/CTRL INPUT_0 0.01fF
C62713 POR2X1_78/A POR2X1_646/O 0.01fF
C62714 POR2X1_454/A PAND2X1_32/B 0.03fF
C62715 PAND2X1_259/O POR2X1_258/Y 0.02fF
C62716 PAND2X1_205/Y PAND2X1_723/Y 0.00fF
C62717 POR2X1_105/Y POR2X1_362/B 0.10fF
C62718 POR2X1_65/A POR2X1_485/O 0.01fF
C62719 POR2X1_180/Y POR2X1_181/Y 0.02fF
C62720 POR2X1_300/O POR2X1_32/A 0.01fF
C62721 POR2X1_78/A PAND2X1_55/Y 0.18fF
C62722 POR2X1_490/Y PAND2X1_572/CTRL2 0.03fF
C62723 POR2X1_499/A POR2X1_362/A 0.19fF
C62724 PAND2X1_23/Y POR2X1_838/B 0.01fF
C62725 POR2X1_224/m4_208_n4# PAND2X1_502/m4_208_n4# 0.13fF
C62726 POR2X1_40/Y POR2X1_531/CTRL2 0.01fF
C62727 PAND2X1_20/A POR2X1_664/Y 0.02fF
C62728 D_GATE_662 POR2X1_174/A 0.07fF
C62729 INPUT_3 PAND2X1_28/O 0.07fF
C62730 POR2X1_846/Y POR2X1_754/a_76_344# 0.00fF
C62731 PAND2X1_57/B POR2X1_593/B 0.04fF
C62732 POR2X1_180/B POR2X1_471/A 0.03fF
C62733 POR2X1_23/Y POR2X1_38/Y 11.74fF
C62734 POR2X1_657/O POR2X1_741/Y 0.01fF
C62735 POR2X1_346/B PAND2X1_43/O 0.00fF
C62736 POR2X1_445/a_76_344# POR2X1_750/B 0.03fF
C62737 POR2X1_775/A PAND2X1_20/A 0.03fF
C62738 PAND2X1_416/CTRL2 POR2X1_260/A 0.01fF
C62739 POR2X1_353/Y POR2X1_502/A 0.03fF
C62740 POR2X1_748/A POR2X1_42/Y 0.05fF
C62741 POR2X1_800/A POR2X1_783/CTRL2 0.00fF
C62742 POR2X1_49/Y POR2X1_58/Y 0.82fF
C62743 POR2X1_862/B POR2X1_784/A 0.02fF
C62744 POR2X1_223/a_16_28# POR2X1_186/Y 0.03fF
C62745 POR2X1_814/A POR2X1_540/Y 0.05fF
C62746 POR2X1_197/CTRL VDD 0.00fF
C62747 PAND2X1_612/B POR2X1_249/Y 0.45fF
C62748 POR2X1_614/A POR2X1_788/A 0.19fF
C62749 POR2X1_81/Y PAND2X1_500/a_76_28# 0.03fF
C62750 PAND2X1_116/CTRL PAND2X1_553/B 0.03fF
C62751 POR2X1_16/A PAND2X1_206/A 0.75fF
C62752 POR2X1_814/A POR2X1_383/a_16_28# 0.02fF
C62753 POR2X1_66/A PAND2X1_393/CTRL 0.00fF
C62754 INPUT_2 POR2X1_104/CTRL 0.01fF
C62755 POR2X1_569/a_16_28# POR2X1_564/Y -0.00fF
C62756 PAND2X1_622/a_16_344# PAND2X1_621/Y 0.04fF
C62757 PAND2X1_20/A POR2X1_112/Y 0.03fF
C62758 POR2X1_188/A POR2X1_805/A 0.03fF
C62759 POR2X1_417/Y PAND2X1_566/Y 0.07fF
C62760 PAND2X1_798/B PAND2X1_579/CTRL2 0.01fF
C62761 PAND2X1_796/B POR2X1_153/Y 0.05fF
C62762 POR2X1_614/A POR2X1_678/A 0.01fF
C62763 POR2X1_37/Y POR2X1_283/A 0.06fF
C62764 PAND2X1_454/O POR2X1_376/B 0.05fF
C62765 PAND2X1_735/Y INPUT_0 0.07fF
C62766 POR2X1_235/Y POR2X1_263/Y 0.01fF
C62767 PAND2X1_479/B VDD 0.11fF
C62768 PAND2X1_454/B POR2X1_153/Y 0.03fF
C62769 POR2X1_296/B POR2X1_318/A 0.08fF
C62770 PAND2X1_807/B PAND2X1_807/O 0.00fF
C62771 PAND2X1_784/A POR2X1_90/Y 0.03fF
C62772 PAND2X1_190/Y PAND2X1_140/O 0.11fF
C62773 POR2X1_751/A POR2X1_408/Y 0.02fF
C62774 POR2X1_859/A POR2X1_546/A 0.05fF
C62775 POR2X1_29/Y POR2X1_159/O 0.09fF
C62776 PAND2X1_643/CTRL POR2X1_595/Y 0.01fF
C62777 POR2X1_360/A VDD 0.34fF
C62778 PAND2X1_225/CTRL POR2X1_38/B -0.03fF
C62779 D_INPUT_0 POR2X1_796/A 0.06fF
C62780 PAND2X1_69/A POR2X1_330/Y 0.08fF
C62781 POR2X1_511/Y POR2X1_55/Y 0.03fF
C62782 POR2X1_348/m4_208_n4# PAND2X1_93/B 0.12fF
C62783 POR2X1_239/CTRL POR2X1_40/Y 0.04fF
C62784 POR2X1_564/Y POR2X1_192/Y 0.03fF
C62785 POR2X1_40/Y POR2X1_594/A 0.02fF
C62786 POR2X1_811/A POR2X1_796/A 0.03fF
C62787 INPUT_1 POR2X1_23/Y 0.12fF
C62788 POR2X1_83/B PAND2X1_388/Y 0.03fF
C62789 POR2X1_334/B PAND2X1_85/Y 0.83fF
C62790 PAND2X1_6/A POR2X1_226/Y 0.03fF
C62791 PAND2X1_404/Y POR2X1_394/A 0.07fF
C62792 PAND2X1_659/B PAND2X1_659/a_76_28# 0.01fF
C62793 POR2X1_37/Y PAND2X1_100/O 0.04fF
C62794 POR2X1_315/Y POR2X1_32/A 0.07fF
C62795 POR2X1_83/B POR2X1_245/a_76_344# 0.02fF
C62796 POR2X1_780/CTRL POR2X1_532/A 0.01fF
C62797 POR2X1_780/CTRL2 POR2X1_780/A 0.01fF
C62798 PAND2X1_76/Y POR2X1_184/Y 0.03fF
C62799 POR2X1_860/A D_INPUT_1 0.03fF
C62800 POR2X1_41/B PAND2X1_793/Y 0.03fF
C62801 POR2X1_83/B PAND2X1_720/CTRL2 -0.00fF
C62802 PAND2X1_859/B INPUT_0 0.21fF
C62803 POR2X1_83/B PAND2X1_549/B 0.03fF
C62804 INPUT_0 PAND2X1_493/Y 0.04fF
C62805 PAND2X1_478/O POR2X1_236/Y 0.01fF
C62806 D_INPUT_5 PAND2X1_3/B 0.05fF
C62807 PAND2X1_218/CTRL2 INPUT_0 0.01fF
C62808 POR2X1_197/O POR2X1_740/Y 0.02fF
C62809 PAND2X1_476/A PAND2X1_9/Y 0.02fF
C62810 POR2X1_639/Y PAND2X1_41/B 0.03fF
C62811 POR2X1_327/Y POR2X1_841/B 0.03fF
C62812 POR2X1_23/Y POR2X1_153/Y 0.32fF
C62813 POR2X1_823/CTRL POR2X1_236/Y 0.01fF
C62814 PAND2X1_645/O PAND2X1_602/Y 0.07fF
C62815 POR2X1_631/A POR2X1_631/a_16_28# 0.01fF
C62816 D_INPUT_0 PAND2X1_514/a_56_28# 0.00fF
C62817 PAND2X1_422/CTRL2 POR2X1_750/B 0.01fF
C62818 POR2X1_453/a_76_344# PAND2X1_60/B 0.01fF
C62819 PAND2X1_63/Y PAND2X1_65/B 0.42fF
C62820 POR2X1_335/a_76_344# POR2X1_740/Y 0.02fF
C62821 POR2X1_65/A PAND2X1_509/O 0.01fF
C62822 POR2X1_113/Y POR2X1_777/B 0.10fF
C62823 POR2X1_79/Y POR2X1_42/Y 0.03fF
C62824 PAND2X1_95/B INPUT_4 0.01fF
C62825 POR2X1_539/A POR2X1_457/O 0.01fF
C62826 PAND2X1_357/Y PAND2X1_730/B 0.03fF
C62827 POR2X1_628/CTRL2 POR2X1_55/Y 0.01fF
C62828 POR2X1_496/Y PAND2X1_508/a_16_344# 0.06fF
C62829 PAND2X1_71/O POR2X1_579/Y 0.00fF
C62830 POR2X1_96/A POR2X1_238/Y 0.03fF
C62831 GATE_741 PAND2X1_357/Y 0.01fF
C62832 PAND2X1_31/O PAND2X1_18/B 0.01fF
C62833 POR2X1_83/B POR2X1_428/O 0.18fF
C62834 POR2X1_96/B POR2X1_40/Y 0.03fF
C62835 POR2X1_483/A POR2X1_203/Y 0.02fF
C62836 POR2X1_7/B POR2X1_743/Y 0.01fF
C62837 POR2X1_65/A POR2X1_142/Y 0.03fF
C62838 POR2X1_57/A POR2X1_5/Y 0.01fF
C62839 PAND2X1_342/a_76_28# POR2X1_5/Y 0.00fF
C62840 PAND2X1_694/CTRL2 POR2X1_614/A 0.00fF
C62841 PAND2X1_236/CTRL2 POR2X1_68/B 0.10fF
C62842 POR2X1_315/Y POR2X1_417/Y 0.18fF
C62843 POR2X1_666/CTRL2 POR2X1_394/A 0.10fF
C62844 POR2X1_257/A POR2X1_524/O 0.18fF
C62845 POR2X1_814/A POR2X1_343/B 0.03fF
C62846 POR2X1_38/Y PAND2X1_558/O 0.03fF
C62847 POR2X1_471/A POR2X1_181/O 0.01fF
C62848 PAND2X1_472/O POR2X1_83/B 0.01fF
C62849 POR2X1_547/a_56_344# POR2X1_502/A 0.00fF
C62850 PAND2X1_308/CTRL2 POR2X1_14/Y 0.00fF
C62851 POR2X1_366/Y PAND2X1_23/Y 0.01fF
C62852 PAND2X1_23/Y POR2X1_294/B 3.05fF
C62853 PAND2X1_69/A POR2X1_585/m4_208_n4# 0.08fF
C62854 POR2X1_471/A POR2X1_169/A 0.03fF
C62855 POR2X1_60/Y PAND2X1_244/B 0.03fF
C62856 PAND2X1_652/Y PAND2X1_652/A -0.02fF
C62857 POR2X1_296/B POR2X1_574/Y 0.03fF
C62858 POR2X1_113/Y PAND2X1_65/B 1.56fF
C62859 PAND2X1_308/CTRL2 PAND2X1_453/A 0.01fF
C62860 POR2X1_35/Y POR2X1_776/B 9.85fF
C62861 POR2X1_539/A POR2X1_543/A 0.03fF
C62862 POR2X1_333/Y POR2X1_78/A 0.00fF
C62863 POR2X1_16/A PAND2X1_444/Y 0.00fF
C62864 PAND2X1_65/B PAND2X1_534/CTRL 0.01fF
C62865 POR2X1_72/B POR2X1_172/O 0.07fF
C62866 POR2X1_57/A PAND2X1_549/CTRL2 0.01fF
C62867 D_INPUT_0 POR2X1_5/O 0.18fF
C62868 POR2X1_274/Y POR2X1_569/A 0.08fF
C62869 PAND2X1_159/m4_208_n4# PAND2X1_460/m4_208_n4# 0.13fF
C62870 POR2X1_806/a_16_28# POR2X1_675/Y 0.04fF
C62871 POR2X1_706/A POR2X1_383/A 0.01fF
C62872 PAND2X1_388/Y PAND2X1_140/Y 0.03fF
C62873 POR2X1_466/A POR2X1_188/Y 0.05fF
C62874 PAND2X1_715/CTRL2 POR2X1_387/Y 0.06fF
C62875 POR2X1_777/B POR2X1_260/A 0.06fF
C62876 POR2X1_614/A PAND2X1_71/O 0.03fF
C62877 POR2X1_717/Y POR2X1_723/B 0.21fF
C62878 PAND2X1_793/Y PAND2X1_548/O 0.02fF
C62879 PAND2X1_194/CTRL VDD -0.00fF
C62880 PAND2X1_41/B POR2X1_352/O 0.02fF
C62881 POR2X1_444/A POR2X1_551/A 0.15fF
C62882 PAND2X1_824/B POR2X1_330/Y 0.07fF
C62883 POR2X1_107/O POR2X1_107/Y 0.00fF
C62884 PAND2X1_90/Y POR2X1_796/A 0.07fF
C62885 POR2X1_300/O POR2X1_184/Y 0.00fF
C62886 PAND2X1_803/Y PAND2X1_543/a_76_28# 0.03fF
C62887 PAND2X1_716/O PAND2X1_197/Y 0.00fF
C62888 POR2X1_60/A PAND2X1_337/a_16_344# 0.06fF
C62889 POR2X1_483/CTRL2 POR2X1_228/Y 0.08fF
C62890 POR2X1_60/A PAND2X1_508/Y 0.06fF
C62891 POR2X1_411/B PAND2X1_332/Y 0.03fF
C62892 POR2X1_850/B POR2X1_737/A 0.01fF
C62893 VDD POR2X1_727/CTRL 0.00fF
C62894 PAND2X1_620/O PAND2X1_620/Y 0.01fF
C62895 POR2X1_283/A PAND2X1_715/O 0.05fF
C62896 POR2X1_185/a_56_344# POR2X1_805/A 0.00fF
C62897 PAND2X1_65/B POR2X1_260/A 4.71fF
C62898 POR2X1_372/Y POR2X1_91/Y 0.03fF
C62899 PAND2X1_839/O PAND2X1_852/B 0.00fF
C62900 POR2X1_814/a_16_28# POR2X1_814/A 0.04fF
C62901 POR2X1_440/O POR2X1_440/B 0.01fF
C62902 PAND2X1_480/B PAND2X1_349/A 0.05fF
C62903 PAND2X1_6/A POR2X1_56/Y 0.02fF
C62904 POR2X1_360/A PAND2X1_82/O 0.02fF
C62905 PAND2X1_726/B POR2X1_692/Y 0.01fF
C62906 PAND2X1_17/CTRL INPUT_6 0.01fF
C62907 POR2X1_291/Y POR2X1_42/Y 0.01fF
C62908 POR2X1_111/Y POR2X1_5/Y 0.01fF
C62909 POR2X1_102/Y PAND2X1_643/A 0.32fF
C62910 POR2X1_66/B PAND2X1_281/a_16_344# 0.02fF
C62911 PAND2X1_260/O PAND2X1_345/Y 0.04fF
C62912 POR2X1_176/Y VDD 0.23fF
C62913 POR2X1_804/B POR2X1_804/A 0.36fF
C62914 POR2X1_96/A PAND2X1_356/O 0.01fF
C62915 POR2X1_383/A PAND2X1_322/O 0.04fF
C62916 POR2X1_96/Y POR2X1_14/Y 0.03fF
C62917 POR2X1_334/B POR2X1_137/Y 0.09fF
C62918 POR2X1_265/Y POR2X1_72/B 2.00fF
C62919 POR2X1_330/Y POR2X1_512/CTRL 0.43fF
C62920 POR2X1_549/CTRL2 POR2X1_266/A 0.01fF
C62921 PAND2X1_63/Y PAND2X1_81/CTRL 0.02fF
C62922 POR2X1_283/A POR2X1_293/Y 0.17fF
C62923 POR2X1_306/O POR2X1_43/B 0.01fF
C62924 POR2X1_566/A PAND2X1_313/CTRL2 0.13fF
C62925 PAND2X1_411/O POR2X1_410/Y -0.00fF
C62926 PAND2X1_860/A POR2X1_20/B 0.02fF
C62927 PAND2X1_450/CTRL POR2X1_425/Y 0.01fF
C62928 POR2X1_85/a_16_28# POR2X1_37/Y 0.00fF
C62929 POR2X1_276/CTRL POR2X1_366/A 0.01fF
C62930 POR2X1_327/Y POR2X1_217/CTRL2 0.01fF
C62931 POR2X1_71/Y PAND2X1_574/CTRL2 0.01fF
C62932 POR2X1_78/CTRL2 PAND2X1_79/Y 0.00fF
C62933 POR2X1_786/Y PAND2X1_150/CTRL2 0.01fF
C62934 POR2X1_486/B POR2X1_590/A 0.01fF
C62935 POR2X1_346/a_16_28# PAND2X1_55/Y 0.02fF
C62936 POR2X1_206/A POR2X1_507/A 0.01fF
C62937 POR2X1_41/B PAND2X1_374/a_16_344# 0.01fF
C62938 PAND2X1_866/O VDD 0.00fF
C62939 POR2X1_860/A POR2X1_362/CTRL2 0.02fF
C62940 POR2X1_345/CTRL POR2X1_244/B 0.01fF
C62941 POR2X1_333/A POR2X1_738/a_16_28# 0.07fF
C62942 POR2X1_619/A POR2X1_816/A 0.03fF
C62943 POR2X1_267/Y POR2X1_318/A 0.03fF
C62944 PAND2X1_319/B PAND2X1_182/CTRL 0.06fF
C62945 PAND2X1_658/B POR2X1_7/A 0.10fF
C62946 POR2X1_519/CTRL POR2X1_42/Y 0.01fF
C62947 POR2X1_315/Y PAND2X1_302/CTRL 0.01fF
C62948 POR2X1_183/Y POR2X1_387/Y 0.03fF
C62949 PAND2X1_264/CTRL POR2X1_42/Y 0.00fF
C62950 POR2X1_68/B PAND2X1_153/CTRL 0.09fF
C62951 POR2X1_669/B POR2X1_747/CTRL 0.01fF
C62952 PAND2X1_69/A POR2X1_148/A 0.19fF
C62953 POR2X1_124/B POR2X1_137/Y 0.00fF
C62954 POR2X1_579/B VDD 0.00fF
C62955 PAND2X1_148/CTRL2 PAND2X1_209/A 0.01fF
C62956 PAND2X1_148/O PAND2X1_148/Y 0.01fF
C62957 POR2X1_8/Y POR2X1_7/B 0.06fF
C62958 POR2X1_741/Y POR2X1_787/CTRL2 0.09fF
C62959 PAND2X1_72/a_76_28# POR2X1_532/A 0.01fF
C62960 PAND2X1_80/O PAND2X1_71/Y 0.02fF
C62961 PAND2X1_738/Y PAND2X1_343/m4_208_n4# 0.04fF
C62962 POR2X1_57/A POR2X1_165/CTRL 0.01fF
C62963 POR2X1_545/A POR2X1_551/CTRL 0.01fF
C62964 POR2X1_327/Y PAND2X1_421/CTRL2 0.00fF
C62965 POR2X1_407/A POR2X1_101/Y 0.03fF
C62966 VDD POR2X1_571/Y 0.34fF
C62967 PAND2X1_737/O PAND2X1_733/Y 0.00fF
C62968 POR2X1_8/Y POR2X1_143/a_16_28# 0.02fF
C62969 PAND2X1_658/A PAND2X1_861/O 0.01fF
C62970 PAND2X1_493/a_16_344# PAND2X1_480/B 0.01fF
C62971 POR2X1_730/Y POR2X1_68/A 0.03fF
C62972 POR2X1_364/A POR2X1_577/Y 0.01fF
C62973 PAND2X1_241/Y POR2X1_239/Y 0.01fF
C62974 POR2X1_99/B VDD 0.05fF
C62975 PAND2X1_671/O PAND2X1_6/A 0.02fF
C62976 POR2X1_16/A PAND2X1_357/Y 0.07fF
C62977 POR2X1_562/CTRL2 POR2X1_186/B 0.02fF
C62978 POR2X1_55/Y POR2X1_129/Y 0.05fF
C62979 POR2X1_289/CTRL2 POR2X1_394/A 0.03fF
C62980 POR2X1_738/A POR2X1_209/A 0.00fF
C62981 PAND2X1_790/Y PAND2X1_156/A 0.18fF
C62982 POR2X1_456/B POR2X1_702/A 0.03fF
C62983 POR2X1_579/B POR2X1_501/CTRL2 0.00fF
C62984 POR2X1_814/A POR2X1_220/CTRL2 0.02fF
C62985 POR2X1_108/O POR2X1_108/Y 0.01fF
C62986 POR2X1_809/A POR2X1_294/B 0.03fF
C62987 POR2X1_343/A POR2X1_343/a_16_28# 0.05fF
C62988 POR2X1_287/B POR2X1_343/a_76_344# 0.00fF
C62989 PAND2X1_364/B POR2X1_7/Y 0.01fF
C62990 POR2X1_271/Y PAND2X1_332/Y 0.03fF
C62991 POR2X1_283/A POR2X1_408/Y 0.02fF
C62992 POR2X1_137/Y POR2X1_218/O 0.00fF
C62993 POR2X1_68/B POR2X1_772/CTRL2 0.09fF
C62994 POR2X1_327/Y POR2X1_114/B 0.07fF
C62995 POR2X1_96/Y PAND2X1_472/B 0.02fF
C62996 PAND2X1_281/a_76_28# POR2X1_121/Y 0.01fF
C62997 POR2X1_677/Y D_INPUT_0 0.03fF
C62998 POR2X1_775/A POR2X1_332/Y 0.34fF
C62999 PAND2X1_473/O PAND2X1_216/B 0.16fF
C63000 PAND2X1_730/A POR2X1_42/Y 1.26fF
C63001 POR2X1_316/Y INPUT_0 0.14fF
C63002 PAND2X1_76/Y PAND2X1_858/B 0.01fF
C63003 POR2X1_394/A PAND2X1_565/A 0.05fF
C63004 POR2X1_837/B PAND2X1_419/O 0.01fF
C63005 PAND2X1_641/a_16_344# POR2X1_38/Y 0.02fF
C63006 POR2X1_172/Y POR2X1_530/O 0.02fF
C63007 POR2X1_72/B POR2X1_167/Y 0.03fF
C63008 POR2X1_96/A POR2X1_184/CTRL2 0.04fF
C63009 POR2X1_66/O PAND2X1_39/B 0.02fF
C63010 POR2X1_548/B PAND2X1_143/O 0.01fF
C63011 POR2X1_9/Y D_INPUT_0 0.58fF
C63012 POR2X1_481/A POR2X1_39/B 0.01fF
C63013 PAND2X1_23/Y POR2X1_567/A 0.14fF
C63014 POR2X1_333/CTRL POR2X1_566/B 0.16fF
C63015 POR2X1_712/O POR2X1_260/A 0.01fF
C63016 PAND2X1_41/B POR2X1_568/A 19.36fF
C63017 POR2X1_653/O POR2X1_711/Y 0.03fF
C63018 POR2X1_96/Y POR2X1_55/Y 0.08fF
C63019 PAND2X1_140/A POR2X1_16/A 0.03fF
C63020 POR2X1_579/B PAND2X1_32/B 0.02fF
C63021 PAND2X1_435/Y POR2X1_677/Y 0.06fF
C63022 POR2X1_257/A POR2X1_150/Y 0.07fF
C63023 POR2X1_99/B POR2X1_741/Y 0.03fF
C63024 POR2X1_541/B PAND2X1_39/B 0.09fF
C63025 PAND2X1_48/B PAND2X1_696/O 0.01fF
C63026 POR2X1_57/A PAND2X1_779/CTRL2 0.01fF
C63027 POR2X1_781/A POR2X1_568/A 0.03fF
C63028 PAND2X1_69/A POR2X1_703/O 0.01fF
C63029 PAND2X1_610/CTRL D_INPUT_2 0.02fF
C63030 POR2X1_249/Y POR2X1_773/CTRL 0.01fF
C63031 D_INPUT_3 POR2X1_4/a_16_28# 0.01fF
C63032 POR2X1_356/A PAND2X1_167/a_76_28# 0.10fF
C63033 POR2X1_365/Y POR2X1_169/A 0.01fF
C63034 POR2X1_571/Y PAND2X1_32/B 0.01fF
C63035 PAND2X1_69/A POR2X1_337/Y 0.12fF
C63036 PAND2X1_793/Y POR2X1_77/Y 0.08fF
C63037 POR2X1_259/O POR2X1_260/A 0.01fF
C63038 POR2X1_493/B POR2X1_773/B 0.04fF
C63039 PAND2X1_321/a_76_28# PAND2X1_52/B 0.02fF
C63040 PAND2X1_194/a_76_28# POR2X1_39/Y 0.07fF
C63041 PAND2X1_856/B PAND2X1_856/CTRL2 0.00fF
C63042 POR2X1_34/m4_208_n4# PAND2X1_32/m4_208_n4# 0.05fF
C63043 POR2X1_863/A PAND2X1_90/Y 0.06fF
C63044 POR2X1_416/B POR2X1_232/CTRL 0.01fF
C63045 PAND2X1_48/B POR2X1_342/Y 0.01fF
C63046 POR2X1_294/B POR2X1_711/Y 0.03fF
C63047 PAND2X1_691/Y PAND2X1_686/a_16_344# 0.01fF
C63048 PAND2X1_633/Y POR2X1_153/Y -0.01fF
C63049 POR2X1_847/CTRL POR2X1_67/A 0.15fF
C63050 PAND2X1_193/Y PAND2X1_596/CTRL 0.01fF
C63051 POR2X1_52/A PAND2X1_332/Y 0.03fF
C63052 POR2X1_20/B POR2X1_268/CTRL2 0.03fF
C63053 POR2X1_83/Y PAND2X1_656/A 0.02fF
C63054 POR2X1_639/Y POR2X1_769/B 0.00fF
C63055 PAND2X1_742/B POR2X1_331/CTRL 0.01fF
C63056 POR2X1_68/A POR2X1_555/O 0.01fF
C63057 PAND2X1_680/O POR2X1_162/Y 0.02fF
C63058 POR2X1_383/A POR2X1_4/Y 0.09fF
C63059 PAND2X1_659/Y POR2X1_7/CTRL2 0.10fF
C63060 POR2X1_86/a_16_28# POR2X1_73/Y 0.02fF
C63061 POR2X1_210/Y POR2X1_568/B 0.05fF
C63062 POR2X1_9/Y PAND2X1_90/Y 0.03fF
C63063 PAND2X1_118/CTRL PAND2X1_72/A 0.01fF
C63064 PAND2X1_317/O POR2X1_314/Y -0.00fF
C63065 POR2X1_294/Y PAND2X1_67/O 0.00fF
C63066 POR2X1_439/Y POR2X1_440/B 0.03fF
C63067 PAND2X1_169/O POR2X1_142/Y 0.02fF
C63068 POR2X1_736/A POR2X1_736/CTRL 0.04fF
C63069 POR2X1_67/Y POR2X1_668/CTRL 0.00fF
C63070 POR2X1_827/CTRL2 VDD 0.00fF
C63071 POR2X1_168/a_76_344# POR2X1_566/B 0.03fF
C63072 POR2X1_760/A POR2X1_250/A 2.30fF
C63073 PAND2X1_79/Y POR2X1_500/CTRL 0.00fF
C63074 POR2X1_411/B POR2X1_226/a_16_28# 0.04fF
C63075 POR2X1_441/Y PAND2X1_545/a_16_344# 0.02fF
C63076 PAND2X1_659/Y PAND2X1_557/CTRL2 0.12fF
C63077 POR2X1_329/A PAND2X1_723/Y 0.03fF
C63078 POR2X1_610/CTRL2 POR2X1_590/A 0.03fF
C63079 POR2X1_394/A POR2X1_701/O 0.01fF
C63080 PAND2X1_73/CTRL PAND2X1_9/Y 0.01fF
C63081 PAND2X1_404/Y POR2X1_669/B 0.02fF
C63082 POR2X1_846/Y POR2X1_615/a_56_344# 0.00fF
C63083 POR2X1_66/B PAND2X1_39/B 2.39fF
C63084 POR2X1_61/a_16_28# POR2X1_61/A 0.03fF
C63085 POR2X1_301/A POR2X1_590/A 0.02fF
C63086 PAND2X1_466/A PAND2X1_803/A 0.00fF
C63087 PAND2X1_261/O POR2X1_814/A 0.13fF
C63088 POR2X1_150/Y PAND2X1_558/CTRL2 0.01fF
C63089 POR2X1_440/B POR2X1_192/Y 0.28fF
C63090 POR2X1_260/B POR2X1_285/Y 0.01fF
C63091 POR2X1_23/Y PAND2X1_794/CTRL2 0.03fF
C63092 POR2X1_188/A PAND2X1_39/B 0.03fF
C63093 POR2X1_99/B POR2X1_228/CTRL 0.00fF
C63094 PAND2X1_206/B POR2X1_88/Y 0.00fF
C63095 POR2X1_48/A POR2X1_819/CTRL2 0.03fF
C63096 POR2X1_411/B PAND2X1_562/B 0.15fF
C63097 POR2X1_294/CTRL POR2X1_355/A 0.01fF
C63098 PAND2X1_86/O POR2X1_243/Y 0.06fF
C63099 POR2X1_399/Y POR2X1_293/Y 0.01fF
C63100 POR2X1_782/B POR2X1_568/B 0.02fF
C63101 POR2X1_681/Y PAND2X1_733/A 0.03fF
C63102 POR2X1_479/B POR2X1_479/CTRL 0.01fF
C63103 PAND2X1_212/B PAND2X1_352/A 0.34fF
C63104 POR2X1_56/CTRL2 POR2X1_496/Y 0.06fF
C63105 PAND2X1_244/B PAND2X1_351/A 0.03fF
C63106 PAND2X1_56/Y POR2X1_458/Y 0.10fF
C63107 POR2X1_96/A PAND2X1_447/CTRL 0.01fF
C63108 POR2X1_14/Y PAND2X1_448/CTRL 0.01fF
C63109 POR2X1_554/B PAND2X1_57/B 0.08fF
C63110 POR2X1_14/Y POR2X1_37/Y 0.08fF
C63111 POR2X1_23/Y PAND2X1_214/A 0.12fF
C63112 POR2X1_411/B PAND2X1_715/CTRL 0.01fF
C63113 PAND2X1_448/O POR2X1_421/Y 0.02fF
C63114 POR2X1_82/O PAND2X1_9/Y 0.01fF
C63115 PAND2X1_477/CTRL2 PAND2X1_803/A 0.00fF
C63116 PAND2X1_58/A PAND2X1_37/CTRL 0.00fF
C63117 POR2X1_650/A POR2X1_473/a_16_28# 0.02fF
C63118 PAND2X1_242/Y POR2X1_283/A 0.05fF
C63119 POR2X1_13/A POR2X1_411/B 0.10fF
C63120 POR2X1_174/B POR2X1_241/B 0.16fF
C63121 POR2X1_294/Y POR2X1_202/CTRL 0.01fF
C63122 POR2X1_54/Y INPUT_0 0.12fF
C63123 POR2X1_150/Y PAND2X1_553/B 0.07fF
C63124 PAND2X1_58/A PAND2X1_752/a_16_344# 0.03fF
C63125 POR2X1_65/Y POR2X1_88/Y 0.29fF
C63126 PAND2X1_138/O POR2X1_39/B 0.01fF
C63127 POR2X1_89/a_76_344# POR2X1_376/B 0.04fF
C63128 POR2X1_600/Y VDD 0.00fF
C63129 POR2X1_748/A POR2X1_67/A 0.07fF
C63130 PAND2X1_56/Y PAND2X1_45/O 0.03fF
C63131 POR2X1_66/B POR2X1_805/Y 0.01fF
C63132 POR2X1_360/A PAND2X1_9/Y 0.15fF
C63133 POR2X1_65/A POR2X1_409/B 0.03fF
C63134 PAND2X1_90/A POR2X1_556/A 0.03fF
C63135 POR2X1_450/Y VDD 0.10fF
C63136 POR2X1_463/CTRL POR2X1_532/A 0.03fF
C63137 POR2X1_499/A POR2X1_572/B 0.03fF
C63138 PAND2X1_558/Y POR2X1_32/A 0.01fF
C63139 POR2X1_289/Y VDD 0.01fF
C63140 POR2X1_66/B PAND2X1_20/A 1.83fF
C63141 POR2X1_450/A POR2X1_121/B 0.04fF
C63142 PAND2X1_65/B PAND2X1_65/O 0.16fF
C63143 POR2X1_503/a_16_28# POR2X1_503/A 0.07fF
C63144 POR2X1_35/B POR2X1_296/B 0.03fF
C63145 PAND2X1_798/O PAND2X1_354/A 0.01fF
C63146 POR2X1_567/A POR2X1_711/Y 0.07fF
C63147 PAND2X1_594/CTRL2 PAND2X1_90/Y 0.14fF
C63148 PAND2X1_39/B POR2X1_828/CTRL 0.06fF
C63149 POR2X1_102/Y POR2X1_609/O 0.01fF
C63150 PAND2X1_73/Y PAND2X1_42/CTRL 0.03fF
C63151 POR2X1_438/Y VDD 0.17fF
C63152 POR2X1_32/O INPUT_3 0.04fF
C63153 PAND2X1_603/CTRL2 PAND2X1_90/Y 0.02fF
C63154 POR2X1_188/A PAND2X1_20/A 0.03fF
C63155 POR2X1_366/Y PAND2X1_271/CTRL2 0.01fF
C63156 POR2X1_686/A POR2X1_78/A 0.01fF
C63157 POR2X1_78/A POR2X1_860/A 1.79fF
C63158 POR2X1_383/A POR2X1_458/Y 0.03fF
C63159 POR2X1_66/B POR2X1_254/CTRL 0.11fF
C63160 POR2X1_41/B POR2X1_827/Y 0.00fF
C63161 POR2X1_753/Y POR2X1_625/O 0.01fF
C63162 POR2X1_168/O POR2X1_168/A 0.01fF
C63163 POR2X1_333/A POR2X1_324/A 0.03fF
C63164 PAND2X1_601/CTRL POR2X1_294/B 0.01fF
C63165 POR2X1_102/Y PAND2X1_805/A 11.57fF
C63166 POR2X1_32/A PAND2X1_596/O 0.01fF
C63167 POR2X1_552/A PAND2X1_72/A 0.01fF
C63168 POR2X1_492/a_16_28# POR2X1_60/A 0.01fF
C63169 INPUT_3 POR2X1_380/CTRL 0.07fF
C63170 POR2X1_109/O POR2X1_7/B 0.17fF
C63171 PAND2X1_47/O PAND2X1_32/B 0.02fF
C63172 POR2X1_278/Y D_INPUT_0 0.17fF
C63173 POR2X1_66/B POR2X1_814/B 0.82fF
C63174 POR2X1_685/A POR2X1_814/A 0.01fF
C63175 POR2X1_52/A PAND2X1_97/O 0.01fF
C63176 POR2X1_115/CTRL POR2X1_218/Y 0.01fF
C63177 POR2X1_10/O POR2X1_9/Y 0.13fF
C63178 POR2X1_796/Y PAND2X1_599/CTRL2 0.01fF
C63179 PAND2X1_643/Y POR2X1_411/B 0.03fF
C63180 PAND2X1_472/B POR2X1_37/Y 0.07fF
C63181 POR2X1_84/A PAND2X1_55/Y 0.03fF
C63182 POR2X1_52/A PAND2X1_448/CTRL2 0.01fF
C63183 POR2X1_20/Y POR2X1_24/Y 0.01fF
C63184 POR2X1_188/A POR2X1_814/B 0.06fF
C63185 PAND2X1_480/B POR2X1_32/A 0.11fF
C63186 PAND2X1_255/CTRL2 POR2X1_186/B 0.01fF
C63187 POR2X1_335/m4_208_n4# POR2X1_66/A 0.09fF
C63188 POR2X1_603/Y VDD 0.09fF
C63189 PAND2X1_413/a_16_344# PAND2X1_57/B 0.01fF
C63190 POR2X1_568/B POR2X1_181/Y 0.03fF
C63191 POR2X1_374/a_16_28# POR2X1_325/B 0.02fF
C63192 PAND2X1_573/CTRL2 PAND2X1_573/B 0.01fF
C63193 POR2X1_66/B POR2X1_325/A 0.03fF
C63194 POR2X1_814/A POR2X1_260/A 2.30fF
C63195 INPUT_3 POR2X1_619/A 0.22fF
C63196 POR2X1_188/A POR2X1_733/CTRL 0.01fF
C63197 POR2X1_37/Y POR2X1_55/Y 0.17fF
C63198 POR2X1_262/Y PAND2X1_560/a_16_344# 0.01fF
C63199 POR2X1_102/Y PAND2X1_735/Y 0.07fF
C63200 POR2X1_221/CTRL POR2X1_186/Y 0.01fF
C63201 POR2X1_855/Y PAND2X1_73/Y 1.32fF
C63202 POR2X1_416/B POR2X1_158/Y 0.01fF
C63203 POR2X1_40/Y POR2X1_236/Y 0.22fF
C63204 PAND2X1_20/A POR2X1_859/A 0.01fF
C63205 POR2X1_418/Y POR2X1_418/O 0.02fF
C63206 POR2X1_130/A POR2X1_288/a_16_28# 0.05fF
C63207 POR2X1_360/A PAND2X1_15/O 0.08fF
C63208 POR2X1_14/Y PAND2X1_377/a_16_344# 0.05fF
C63209 POR2X1_193/Y POR2X1_61/Y 0.07fF
C63210 POR2X1_41/B POR2X1_516/Y 0.07fF
C63211 POR2X1_43/B POR2X1_420/CTRL 0.01fF
C63212 POR2X1_460/A PAND2X1_26/A 0.25fF
C63213 PAND2X1_93/CTRL POR2X1_66/A 0.01fF
C63214 POR2X1_683/a_16_28# POR2X1_669/B 0.02fF
C63215 POR2X1_446/B POR2X1_724/A 0.07fF
C63216 PAND2X1_294/CTRL2 POR2X1_387/Y 0.06fF
C63217 POR2X1_596/A POR2X1_644/CTRL2 0.01fF
C63218 PAND2X1_275/CTRL2 POR2X1_296/B 0.02fF
C63219 POR2X1_718/O PAND2X1_65/B 0.07fF
C63220 POR2X1_13/A POR2X1_271/Y 0.03fF
C63221 D_INPUT_0 PAND2X1_744/CTRL 0.09fF
C63222 POR2X1_846/Y POR2X1_260/A 0.03fF
C63223 POR2X1_814/A POR2X1_363/A 0.04fF
C63224 PAND2X1_57/CTRL PAND2X1_41/B 0.01fF
C63225 POR2X1_707/A PAND2X1_57/B 0.01fF
C63226 PAND2X1_44/O PAND2X1_587/Y 0.00fF
C63227 POR2X1_417/Y PAND2X1_480/B 0.03fF
C63228 POR2X1_68/A POR2X1_218/Y 0.10fF
C63229 PAND2X1_6/Y POR2X1_856/B 0.05fF
C63230 POR2X1_556/A POR2X1_787/CTRL 0.01fF
C63231 POR2X1_14/Y POR2X1_293/Y 0.11fF
C63232 POR2X1_855/B POR2X1_452/Y 0.02fF
C63233 PAND2X1_863/B PAND2X1_249/O 0.02fF
C63234 POR2X1_102/Y PAND2X1_493/Y 0.10fF
C63235 POR2X1_683/CTRL2 POR2X1_72/B 0.03fF
C63236 POR2X1_41/B PAND2X1_361/a_16_344# 0.02fF
C63237 PAND2X1_55/Y POR2X1_285/Y 0.03fF
C63238 POR2X1_754/Y PAND2X1_6/A 0.07fF
C63239 PAND2X1_854/O POR2X1_102/Y 0.05fF
C63240 PAND2X1_846/m4_208_n4# POR2X1_750/A 0.09fF
C63241 POR2X1_720/B POR2X1_29/A 0.03fF
C63242 PAND2X1_462/B POR2X1_607/A 0.07fF
C63243 POR2X1_102/Y PAND2X1_174/O 0.02fF
C63244 POR2X1_23/Y POR2X1_591/Y 0.05fF
C63245 INPUT_2 D_INPUT_0 0.02fF
C63246 POR2X1_48/A PAND2X1_645/B 0.00fF
C63247 PAND2X1_84/Y POR2X1_5/Y 0.01fF
C63248 POR2X1_855/B POR2X1_808/CTRL2 0.01fF
C63249 PAND2X1_630/a_16_344# POR2X1_496/Y 0.03fF
C63250 POR2X1_355/B POR2X1_509/B 0.14fF
C63251 POR2X1_407/A POR2X1_843/O 0.01fF
C63252 POR2X1_567/B POR2X1_190/O 0.34fF
C63253 POR2X1_632/a_76_344# PAND2X1_88/Y 0.00fF
C63254 PAND2X1_80/a_76_28# PAND2X1_41/B 0.01fF
C63255 POR2X1_708/CTRL PAND2X1_90/Y 0.05fF
C63256 POR2X1_254/Y PAND2X1_13/a_16_344# 0.01fF
C63257 PAND2X1_108/a_76_28# POR2X1_862/B 0.07fF
C63258 PAND2X1_340/a_16_344# INPUT_0 0.04fF
C63259 POR2X1_502/A POR2X1_287/B 0.21fF
C63260 POR2X1_48/A INPUT_6 0.02fF
C63261 POR2X1_49/Y PAND2X1_364/B 0.07fF
C63262 PAND2X1_844/CTRL2 POR2X1_20/B 0.01fF
C63263 POR2X1_13/A POR2X1_376/B 0.11fF
C63264 PAND2X1_473/B PAND2X1_580/B 0.03fF
C63265 POR2X1_631/a_56_344# POR2X1_294/B 0.00fF
C63266 POR2X1_716/O POR2X1_303/B 0.01fF
C63267 POR2X1_13/A PAND2X1_596/CTRL2 0.00fF
C63268 PAND2X1_73/Y POR2X1_576/Y 0.00fF
C63269 PAND2X1_129/CTRL POR2X1_502/A 0.47fF
C63270 POR2X1_51/a_16_28# POR2X1_51/A 0.07fF
C63271 POR2X1_834/Y PAND2X1_601/CTRL2 0.15fF
C63272 PAND2X1_12/CTRL2 POR2X1_260/A 0.02fF
C63273 POR2X1_638/A POR2X1_638/B 0.00fF
C63274 INPUT_0 POR2X1_572/CTRL2 0.04fF
C63275 PAND2X1_531/O PAND2X1_32/B 0.08fF
C63276 PAND2X1_94/A POR2X1_862/A 0.68fF
C63277 PAND2X1_404/A POR2X1_233/CTRL2 0.00fF
C63278 PAND2X1_13/CTRL2 POR2X1_795/B 0.01fF
C63279 POR2X1_567/B POR2X1_569/A 0.10fF
C63280 PAND2X1_274/a_16_344# POR2X1_272/Y 0.01fF
C63281 PAND2X1_478/Y POR2X1_238/Y 0.03fF
C63282 PAND2X1_479/A PAND2X1_579/B 0.02fF
C63283 POR2X1_20/B PAND2X1_156/A 2.49fF
C63284 POR2X1_651/O PAND2X1_90/Y 0.01fF
C63285 POR2X1_502/A PAND2X1_8/Y 0.01fF
C63286 PAND2X1_483/CTRL2 POR2X1_23/Y 0.02fF
C63287 PAND2X1_105/CTRL2 PAND2X1_562/B 0.03fF
C63288 POR2X1_245/Y PAND2X1_777/O -0.00fF
C63289 POR2X1_280/Y PAND2X1_771/Y 0.08fF
C63290 PAND2X1_288/A PAND2X1_366/Y 0.54fF
C63291 POR2X1_13/A PAND2X1_735/a_16_344# 0.02fF
C63292 POR2X1_356/A POR2X1_78/B 0.10fF
C63293 POR2X1_52/A PAND2X1_474/Y 0.03fF
C63294 PAND2X1_583/CTRL POR2X1_750/B 0.01fF
C63295 POR2X1_614/A POR2X1_264/a_56_344# 0.00fF
C63296 POR2X1_516/O POR2X1_423/Y 0.01fF
C63297 POR2X1_113/Y POR2X1_650/O 0.18fF
C63298 PAND2X1_553/A PAND2X1_553/B 0.09fF
C63299 POR2X1_673/Y POR2X1_623/CTRL2 0.04fF
C63300 PAND2X1_137/Y PAND2X1_768/CTRL 0.01fF
C63301 POR2X1_57/A POR2X1_825/CTRL2 0.03fF
C63302 POR2X1_567/B POR2X1_570/Y 0.59fF
C63303 POR2X1_502/A POR2X1_170/B 0.03fF
C63304 POR2X1_193/Y POR2X1_35/Y 0.03fF
C63305 POR2X1_499/O POR2X1_456/B 0.01fF
C63306 PAND2X1_735/O POR2X1_293/Y 0.03fF
C63307 PAND2X1_216/B POR2X1_48/A 0.01fF
C63308 POR2X1_664/Y VDD 0.14fF
C63309 POR2X1_52/A POR2X1_13/A 3.47fF
C63310 POR2X1_14/Y POR2X1_408/Y 0.05fF
C63311 PAND2X1_824/B POR2X1_630/CTRL 0.07fF
C63312 PAND2X1_151/CTRL2 POR2X1_55/Y 0.03fF
C63313 POR2X1_404/B POR2X1_404/Y 0.01fF
C63314 POR2X1_471/CTRL2 POR2X1_732/B 0.08fF
C63315 PAND2X1_635/CTRL POR2X1_763/A 0.09fF
C63316 POR2X1_96/A PAND2X1_191/CTRL 0.01fF
C63317 POR2X1_41/B POR2X1_821/a_16_28# 0.09fF
C63318 D_INPUT_5 PAND2X1_2/O 0.01fF
C63319 PAND2X1_275/CTRL VDD -0.00fF
C63320 POR2X1_65/A POR2X1_93/O 0.21fF
C63321 PAND2X1_714/A POR2X1_90/Y 0.07fF
C63322 PAND2X1_261/O POR2X1_260/Y 0.03fF
C63323 POR2X1_124/B POR2X1_650/A 0.01fF
C63324 POR2X1_13/Y INPUT_0 0.03fF
C63325 POR2X1_573/CTRL2 POR2X1_576/Y 0.01fF
C63326 POR2X1_60/A POR2X1_283/A 0.10fF
C63327 PAND2X1_679/O PAND2X1_69/A 0.02fF
C63328 POR2X1_515/CTRL2 PAND2X1_6/Y 0.17fF
C63329 PAND2X1_317/Y POR2X1_13/A 0.13fF
C63330 POR2X1_52/A PAND2X1_214/B 0.25fF
C63331 POR2X1_775/A VDD 0.01fF
C63332 PAND2X1_94/A PAND2X1_73/Y 1.01fF
C63333 PAND2X1_48/B POR2X1_115/O 0.09fF
C63334 POR2X1_392/B PAND2X1_153/O 0.08fF
C63335 POR2X1_49/Y PAND2X1_560/CTRL 0.01fF
C63336 POR2X1_566/A POR2X1_563/Y 0.03fF
C63337 POR2X1_186/Y POR2X1_318/A 0.19fF
C63338 POR2X1_536/CTRL POR2X1_102/Y 0.01fF
C63339 POR2X1_121/B PAND2X1_300/O 0.01fF
C63340 POR2X1_433/Y VDD 0.30fF
C63341 POR2X1_463/Y POR2X1_792/O 0.02fF
C63342 POR2X1_192/Y POR2X1_222/Y 0.03fF
C63343 POR2X1_220/Y POR2X1_221/Y -0.00fF
C63344 PAND2X1_264/O POR2X1_83/B 0.09fF
C63345 POR2X1_199/CTRL POR2X1_740/Y 0.00fF
C63346 POR2X1_199/CTRL2 POR2X1_741/Y 0.04fF
C63347 PAND2X1_824/CTRL PAND2X1_41/B 0.00fF
C63348 POR2X1_62/Y POR2X1_614/O 0.06fF
C63349 PAND2X1_836/CTRL VDD 0.00fF
C63350 POR2X1_55/Y POR2X1_293/Y 5.33fF
C63351 POR2X1_515/a_76_344# POR2X1_68/A 0.03fF
C63352 PAND2X1_480/B POR2X1_184/Y 0.05fF
C63353 POR2X1_136/O VDD 0.00fF
C63354 POR2X1_548/B PAND2X1_90/A 0.06fF
C63355 POR2X1_302/a_76_344# PAND2X1_6/Y 0.01fF
C63356 POR2X1_102/Y POR2X1_172/a_16_28# 0.03fF
C63357 POR2X1_48/A POR2X1_749/m4_208_n4# 0.09fF
C63358 PAND2X1_140/A POR2X1_127/Y 0.04fF
C63359 PAND2X1_23/Y PAND2X1_816/CTRL2 0.13fF
C63360 POR2X1_718/CTRL POR2X1_832/A 0.01fF
C63361 POR2X1_809/A POR2X1_809/a_16_28# 0.05fF
C63362 VDD POR2X1_112/Y 0.40fF
C63363 POR2X1_502/A POR2X1_705/CTRL2 0.01fF
C63364 POR2X1_57/A PAND2X1_723/Y 0.03fF
C63365 POR2X1_401/CTRL POR2X1_68/B 0.01fF
C63366 POR2X1_167/CTRL2 PAND2X1_714/A 0.02fF
C63367 PAND2X1_6/A POR2X1_817/A 0.03fF
C63368 POR2X1_334/B POR2X1_294/B 0.14fF
C63369 PAND2X1_6/Y POR2X1_722/Y 0.03fF
C63370 PAND2X1_252/m4_208_n4# POR2X1_254/m4_208_n4# 0.05fF
C63371 PAND2X1_859/CTRL POR2X1_283/A 0.00fF
C63372 PAND2X1_58/A POR2X1_753/CTRL 0.18fF
C63373 POR2X1_471/CTRL POR2X1_540/A 0.00fF
C63374 POR2X1_57/A PAND2X1_347/Y 2.39fF
C63375 POR2X1_56/B POR2X1_43/B 0.14fF
C63376 POR2X1_25/a_56_344# D_INPUT_6 0.00fF
C63377 POR2X1_702/B POR2X1_383/A 0.03fF
C63378 POR2X1_355/B POR2X1_508/a_16_28# 0.00fF
C63379 POR2X1_660/A POR2X1_725/Y 0.06fF
C63380 PAND2X1_865/Y PAND2X1_287/Y 0.46fF
C63381 PAND2X1_57/B POR2X1_702/A 0.03fF
C63382 PAND2X1_209/A PAND2X1_209/a_76_28# 0.05fF
C63383 PAND2X1_783/Y PAND2X1_549/B 0.18fF
C63384 D_INPUT_6 VDD 0.66fF
C63385 POR2X1_51/B POR2X1_44/O 0.03fF
C63386 PAND2X1_488/CTRL2 POR2X1_260/A 0.01fF
C63387 INPUT_1 POR2X1_49/CTRL 0.01fF
C63388 POR2X1_196/O POR2X1_334/Y 0.06fF
C63389 PAND2X1_23/Y PAND2X1_504/CTRL 0.01fF
C63390 POR2X1_49/Y PAND2X1_849/B 0.00fF
C63391 POR2X1_256/a_76_344# POR2X1_255/Y 0.02fF
C63392 POR2X1_447/B POR2X1_294/Y 0.02fF
C63393 POR2X1_192/Y POR2X1_532/A 0.05fF
C63394 PAND2X1_23/Y POR2X1_140/B 0.03fF
C63395 POR2X1_376/B PAND2X1_510/B 0.03fF
C63396 PAND2X1_293/CTRL2 PAND2X1_60/B 0.01fF
C63397 PAND2X1_23/Y POR2X1_407/A 0.07fF
C63398 PAND2X1_661/Y POR2X1_666/A 0.04fF
C63399 PAND2X1_6/A POR2X1_42/Y 0.29fF
C63400 POR2X1_861/A POR2X1_218/Y 0.04fF
C63401 POR2X1_52/A PAND2X1_661/B 0.03fF
C63402 POR2X1_307/B POR2X1_590/O 0.03fF
C63403 POR2X1_852/B POR2X1_260/A 0.07fF
C63404 PAND2X1_281/CTRL POR2X1_285/Y 0.00fF
C63405 VDD POR2X1_162/Y -0.00fF
C63406 POR2X1_124/B POR2X1_294/B 0.02fF
C63407 POR2X1_68/B POR2X1_7/B 0.31fF
C63408 POR2X1_776/A PAND2X1_52/B 0.09fF
C63409 PAND2X1_217/CTRL2 PAND2X1_364/B 0.03fF
C63410 POR2X1_78/B POR2X1_569/A 0.17fF
C63411 POR2X1_316/Y PAND2X1_436/a_56_28# 0.00fF
C63412 PAND2X1_41/B POR2X1_444/Y 0.25fF
C63413 POR2X1_578/Y POR2X1_578/CTRL2 0.00fF
C63414 POR2X1_123/B POR2X1_123/CTRL2 0.03fF
C63415 POR2X1_790/B POR2X1_790/A 0.12fF
C63416 POR2X1_192/Y POR2X1_714/a_56_344# 0.00fF
C63417 POR2X1_590/A POR2X1_362/CTRL 0.01fF
C63418 POR2X1_96/A POR2X1_387/Y 0.14fF
C63419 POR2X1_120/a_16_28# PAND2X1_60/B 0.03fF
C63420 POR2X1_72/B PAND2X1_853/B 0.03fF
C63421 POR2X1_267/A POR2X1_571/Y 0.03fF
C63422 POR2X1_614/A D_GATE_811 0.01fF
C63423 POR2X1_23/CTRL2 POR2X1_4/Y 0.10fF
C63424 PAND2X1_631/A POR2X1_56/CTRL 0.01fF
C63425 PAND2X1_170/O PAND2X1_169/Y 0.15fF
C63426 PAND2X1_6/Y PAND2X1_7/a_16_344# 0.03fF
C63427 POR2X1_596/A PAND2X1_604/CTRL 0.01fF
C63428 POR2X1_800/A POR2X1_828/A 0.03fF
C63429 POR2X1_827/Y POR2X1_77/Y 0.03fF
C63430 POR2X1_788/A POR2X1_788/CTRL2 0.01fF
C63431 POR2X1_640/a_76_344# POR2X1_559/A 0.10fF
C63432 POR2X1_741/Y POR2X1_112/Y 0.03fF
C63433 PAND2X1_741/B POR2X1_7/O 0.13fF
C63434 PAND2X1_467/Y VDD 0.31fF
C63435 POR2X1_775/A PAND2X1_32/B 0.87fF
C63436 POR2X1_840/B POR2X1_130/Y 0.10fF
C63437 POR2X1_401/A PAND2X1_69/A 0.01fF
C63438 PAND2X1_844/O PAND2X1_61/Y 0.02fF
C63439 POR2X1_94/A POR2X1_523/B 0.02fF
C63440 POR2X1_791/O POR2X1_791/A 0.01fF
C63441 INPUT_1 POR2X1_372/A 0.00fF
C63442 POR2X1_334/CTRL2 INPUT_0 0.03fF
C63443 PAND2X1_408/CTRL PAND2X1_408/Y 0.00fF
C63444 POR2X1_119/Y PAND2X1_575/B 0.05fF
C63445 POR2X1_78/B PAND2X1_232/a_56_28# 0.00fF
C63446 POR2X1_840/Y POR2X1_590/A 0.03fF
C63447 PAND2X1_86/Y VDD 0.14fF
C63448 POR2X1_297/O PAND2X1_359/Y 0.01fF
C63449 POR2X1_96/A POR2X1_134/O 0.01fF
C63450 POR2X1_616/Y POR2X1_748/A 0.03fF
C63451 PAND2X1_65/B POR2X1_559/A 4.21fF
C63452 PAND2X1_56/Y POR2X1_724/A 0.10fF
C63453 POR2X1_90/Y POR2X1_816/A 0.12fF
C63454 POR2X1_52/CTRL2 POR2X1_102/Y 0.01fF
C63455 POR2X1_408/Y POR2X1_55/Y 0.15fF
C63456 PAND2X1_835/a_76_28# PAND2X1_852/B 0.02fF
C63457 PAND2X1_649/A POR2X1_394/Y 0.01fF
C63458 POR2X1_334/B PAND2X1_111/B 0.03fF
C63459 POR2X1_730/Y POR2X1_435/Y 0.07fF
C63460 PAND2X1_812/CTRL2 PAND2X1_811/Y 0.00fF
C63461 PAND2X1_441/CTRL POR2X1_854/B 0.32fF
C63462 POR2X1_52/A PAND2X1_510/B 0.02fF
C63463 POR2X1_187/O POR2X1_79/Y 0.01fF
C63464 POR2X1_325/CTRL PAND2X1_55/Y 0.08fF
C63465 POR2X1_41/B PAND2X1_114/CTRL 0.02fF
C63466 PAND2X1_276/O POR2X1_129/Y 0.02fF
C63467 POR2X1_112/Y PAND2X1_32/B 0.03fF
C63468 POR2X1_465/B POR2X1_553/A 0.09fF
C63469 POR2X1_614/A POR2X1_540/A 0.03fF
C63470 POR2X1_697/Y PAND2X1_549/B 0.01fF
C63471 POR2X1_372/A POR2X1_153/Y 0.05fF
C63472 POR2X1_306/CTRL2 POR2X1_90/Y 0.01fF
C63473 POR2X1_588/Y POR2X1_42/Y 0.07fF
C63474 POR2X1_644/A POR2X1_796/m4_208_n4# 0.07fF
C63475 POR2X1_567/B PAND2X1_72/A 0.38fF
C63476 POR2X1_133/CTRL2 POR2X1_384/A 0.01fF
C63477 PAND2X1_388/Y PAND2X1_357/Y 0.03fF
C63478 PAND2X1_824/B POR2X1_214/CTRL 0.07fF
C63479 POR2X1_419/CTRL2 POR2X1_42/Y 0.02fF
C63480 INPUT_5 POR2X1_260/A 0.18fF
C63481 D_INPUT_6 PAND2X1_32/B 0.71fF
C63482 POR2X1_51/B POR2X1_587/CTRL 0.01fF
C63483 POR2X1_390/B PAND2X1_48/B 0.03fF
C63484 POR2X1_287/B POR2X1_188/Y 0.07fF
C63485 POR2X1_466/Y POR2X1_568/B 0.03fF
C63486 POR2X1_96/A POR2X1_419/a_16_28# 0.02fF
C63487 PAND2X1_384/CTRL2 POR2X1_546/A 0.12fF
C63488 VDD POR2X1_339/Y -0.00fF
C63489 POR2X1_8/Y POR2X1_618/CTRL 0.01fF
C63490 POR2X1_703/A PAND2X1_178/CTRL 0.00fF
C63491 PAND2X1_404/Y POR2X1_234/A 0.47fF
C63492 PAND2X1_72/O PAND2X1_60/B 0.01fF
C63493 PAND2X1_63/Y POR2X1_493/O 0.04fF
C63494 POR2X1_316/Y PAND2X1_436/A 0.11fF
C63495 POR2X1_844/a_16_28# D_INPUT_1 0.02fF
C63496 PAND2X1_737/B PAND2X1_197/Y 0.00fF
C63497 PAND2X1_291/CTRL2 PAND2X1_88/Y 0.01fF
C63498 POR2X1_513/Y POR2X1_366/A 0.03fF
C63499 POR2X1_67/Y POR2X1_816/CTRL2 0.03fF
C63500 POR2X1_614/A POR2X1_539/A 0.03fF
C63501 POR2X1_327/Y POR2X1_405/Y 0.01fF
C63502 POR2X1_13/A POR2X1_3/B 0.01fF
C63503 POR2X1_383/A D_INPUT_1 0.10fF
C63504 POR2X1_68/B PAND2X1_60/B 0.11fF
C63505 PAND2X1_816/a_16_344# POR2X1_260/A 0.02fF
C63506 PAND2X1_854/A POR2X1_90/Y 0.01fF
C63507 POR2X1_538/A PAND2X1_69/A 0.02fF
C63508 POR2X1_114/B POR2X1_249/Y 0.03fF
C63509 PAND2X1_344/O POR2X1_91/Y 0.07fF
C63510 D_GATE_222 POR2X1_332/CTRL2 0.01fF
C63511 PAND2X1_109/CTRL PAND2X1_41/B 0.00fF
C63512 POR2X1_583/Y POR2X1_42/Y -0.02fF
C63513 POR2X1_567/B POR2X1_535/O 0.00fF
C63514 POR2X1_722/A PAND2X1_48/B 0.32fF
C63515 PAND2X1_71/CTRL PAND2X1_71/Y 0.01fF
C63516 POR2X1_377/a_16_28# PAND2X1_94/A 0.01fF
C63517 POR2X1_21/a_16_28# POR2X1_460/A 0.03fF
C63518 POR2X1_260/Y POR2X1_363/A 0.03fF
C63519 POR2X1_334/A POR2X1_198/B 0.01fF
C63520 INPUT_0 POR2X1_4/Y 0.14fF
C63521 POR2X1_407/Y PAND2X1_765/a_16_344# 0.00fF
C63522 POR2X1_532/A POR2X1_568/Y 0.05fF
C63523 PAND2X1_467/Y POR2X1_694/a_16_28# 0.01fF
C63524 PAND2X1_41/B PAND2X1_56/A 0.03fF
C63525 PAND2X1_6/Y POR2X1_799/a_16_28# 0.00fF
C63526 PAND2X1_658/B POR2X1_153/Y 0.10fF
C63527 POR2X1_610/Y POR2X1_814/A 0.19fF
C63528 POR2X1_7/A POR2X1_387/Y 1.45fF
C63529 PAND2X1_633/CTRL POR2X1_77/Y 0.01fF
C63530 PAND2X1_496/CTRL PAND2X1_48/A 0.00fF
C63531 POR2X1_648/A POR2X1_648/a_16_28# 0.03fF
C63532 POR2X1_87/CTRL PAND2X1_41/B 0.01fF
C63533 POR2X1_807/A POR2X1_711/Y 0.02fF
C63534 POR2X1_68/B POR2X1_773/O 0.16fF
C63535 POR2X1_730/Y PAND2X1_96/B 10.08fF
C63536 PAND2X1_6/Y POR2X1_244/Y 0.06fF
C63537 POR2X1_78/B PAND2X1_290/CTRL 0.00fF
C63538 POR2X1_216/CTRL POR2X1_101/Y 0.03fF
C63539 POR2X1_71/Y POR2X1_119/Y 0.14fF
C63540 POR2X1_32/A POR2X1_386/Y 0.36fF
C63541 PAND2X1_61/Y PAND2X1_339/a_76_28# 0.02fF
C63542 PAND2X1_569/O POR2X1_73/Y 0.01fF
C63543 POR2X1_516/A POR2X1_283/A 0.03fF
C63544 PAND2X1_514/Y PAND2X1_716/B 0.05fF
C63545 POR2X1_41/B PAND2X1_797/Y 0.07fF
C63546 POR2X1_119/Y POR2X1_42/Y 0.05fF
C63547 POR2X1_809/A POR2X1_407/A 0.03fF
C63548 PAND2X1_283/CTRL POR2X1_294/A 0.00fF
C63549 POR2X1_7/B PAND2X1_539/a_16_344# 0.02fF
C63550 POR2X1_68/B POR2X1_571/O 0.01fF
C63551 POR2X1_493/O POR2X1_260/A 0.01fF
C63552 POR2X1_461/Y POR2X1_859/O 0.01fF
C63553 POR2X1_85/Y PAND2X1_206/CTRL2 0.01fF
C63554 PAND2X1_469/B POR2X1_183/a_56_344# 0.00fF
C63555 POR2X1_188/O POR2X1_456/B 0.17fF
C63556 POR2X1_244/Y POR2X1_575/CTRL2 0.10fF
C63557 D_INPUT_1 PAND2X1_71/Y 0.03fF
C63558 POR2X1_862/a_76_344# POR2X1_480/A 0.03fF
C63559 PAND2X1_359/Y PAND2X1_359/O 0.01fF
C63560 POR2X1_709/CTRL2 INPUT_1 0.01fF
C63561 POR2X1_618/a_16_28# POR2X1_4/Y 0.02fF
C63562 POR2X1_411/B PAND2X1_562/Y 0.72fF
C63563 POR2X1_814/A PAND2X1_65/O 0.02fF
C63564 PAND2X1_672/O D_INPUT_1 0.01fF
C63565 POR2X1_69/Y POR2X1_66/A 0.05fF
C63566 PAND2X1_294/CTRL POR2X1_411/B 0.01fF
C63567 PAND2X1_593/Y PAND2X1_537/CTRL2 0.01fF
C63568 POR2X1_252/Y PAND2X1_6/A 0.03fF
C63569 PAND2X1_211/O POR2X1_411/B 0.01fF
C63570 POR2X1_78/B PAND2X1_72/A 0.16fF
C63571 PAND2X1_69/A POR2X1_342/O 0.02fF
C63572 POR2X1_192/Y POR2X1_567/a_16_28# 0.02fF
C63573 PAND2X1_847/O POR2X1_820/Y 0.03fF
C63574 PAND2X1_232/CTRL2 POR2X1_260/A 0.03fF
C63575 POR2X1_257/A PAND2X1_213/CTRL2 0.00fF
C63576 POR2X1_416/B POR2X1_425/O 0.18fF
C63577 PAND2X1_613/CTRL2 PAND2X1_9/Y 0.01fF
C63578 POR2X1_523/Y POR2X1_560/a_16_28# -0.00fF
C63579 PAND2X1_193/Y PAND2X1_733/O 0.05fF
C63580 POR2X1_383/A POR2X1_734/m4_208_n4# 0.12fF
C63581 POR2X1_846/a_16_28# POR2X1_750/B 0.03fF
C63582 PAND2X1_134/CTRL2 PAND2X1_32/B 0.00fF
C63583 POR2X1_326/A PAND2X1_60/B 0.03fF
C63584 POR2X1_745/Y POR2X1_746/CTRL2 0.00fF
C63585 POR2X1_154/CTRL PAND2X1_72/A 0.11fF
C63586 POR2X1_669/B POR2X1_67/Y 0.05fF
C63587 PAND2X1_38/CTRL PAND2X1_52/B 0.01fF
C63588 POR2X1_52/A POR2X1_387/O 0.02fF
C63589 PAND2X1_96/B PAND2X1_323/CTRL 0.00fF
C63590 PAND2X1_508/Y PAND2X1_175/B 0.03fF
C63591 PAND2X1_865/Y PAND2X1_575/CTRL2 0.00fF
C63592 POR2X1_165/Y PAND2X1_569/B 0.05fF
C63593 POR2X1_566/A PAND2X1_292/a_16_344# 0.04fF
C63594 POR2X1_456/B POR2X1_703/Y 0.01fF
C63595 POR2X1_209/A POR2X1_726/a_56_344# 0.00fF
C63596 POR2X1_1/CTRL PAND2X1_18/B 0.06fF
C63597 POR2X1_164/Y POR2X1_394/A 0.03fF
C63598 PAND2X1_349/A POR2X1_131/A 0.00fF
C63599 PAND2X1_171/CTRL POR2X1_854/B 0.30fF
C63600 POR2X1_186/CTRL POR2X1_353/A 0.01fF
C63601 POR2X1_218/a_16_28# POR2X1_216/Y -0.00fF
C63602 POR2X1_623/CTRL2 PAND2X1_9/Y 0.01fF
C63603 POR2X1_383/A POR2X1_620/B 0.03fF
C63604 POR2X1_326/A POR2X1_737/CTRL 0.14fF
C63605 POR2X1_569/A POR2X1_294/A 0.07fF
C63606 POR2X1_407/A POR2X1_711/Y 0.07fF
C63607 PAND2X1_439/CTRL POR2X1_72/B 0.01fF
C63608 PAND2X1_404/CTRL POR2X1_411/A 0.01fF
C63609 PAND2X1_93/B POR2X1_446/B 0.03fF
C63610 POR2X1_486/B POR2X1_532/A 0.10fF
C63611 POR2X1_499/A POR2X1_590/A 7.73fF
C63612 POR2X1_411/B PAND2X1_722/O 0.02fF
C63613 POR2X1_814/A POR2X1_489/CTRL 0.01fF
C63614 POR2X1_411/B POR2X1_29/A 0.06fF
C63615 POR2X1_326/A POR2X1_353/A 0.03fF
C63616 POR2X1_270/Y POR2X1_222/O 0.01fF
C63617 PAND2X1_631/O POR2X1_416/B 0.02fF
C63618 POR2X1_407/A POR2X1_728/A 0.00fF
C63619 POR2X1_669/B POR2X1_604/CTRL2 0.01fF
C63620 POR2X1_122/CTRL POR2X1_394/A 0.03fF
C63621 POR2X1_565/O PAND2X1_52/B 0.05fF
C63622 POR2X1_87/CTRL2 POR2X1_68/B 0.05fF
C63623 POR2X1_462/O POR2X1_734/A 0.03fF
C63624 PAND2X1_242/Y POR2X1_55/Y 0.03fF
C63625 PAND2X1_641/Y PAND2X1_341/B 0.01fF
C63626 POR2X1_863/A D_GATE_222 0.02fF
C63627 POR2X1_88/CTRL POR2X1_669/B 0.02fF
C63628 POR2X1_180/B POR2X1_181/O 0.00fF
C63629 POR2X1_13/A PAND2X1_458/a_16_344# 0.01fF
C63630 POR2X1_78/A POR2X1_446/B 0.03fF
C63631 POR2X1_76/A POR2X1_590/A 0.19fF
C63632 PAND2X1_48/B PAND2X1_628/CTRL 0.01fF
C63633 PAND2X1_630/B POR2X1_7/B 0.03fF
C63634 POR2X1_180/B POR2X1_169/A 0.00fF
C63635 PAND2X1_58/A PAND2X1_24/a_16_344# 0.02fF
C63636 PAND2X1_658/A PAND2X1_860/A 0.44fF
C63637 PAND2X1_139/O POR2X1_150/Y 0.01fF
C63638 POR2X1_75/Y PAND2X1_716/B 0.56fF
C63639 PAND2X1_458/O POR2X1_293/Y 0.12fF
C63640 POR2X1_411/B POR2X1_820/A 0.07fF
C63641 POR2X1_9/Y POR2X1_617/CTRL 0.04fF
C63642 POR2X1_416/B PAND2X1_181/CTRL 0.12fF
C63643 POR2X1_865/B POR2X1_343/B 0.03fF
C63644 POR2X1_750/Y POR2X1_39/B 0.03fF
C63645 POR2X1_505/a_16_28# PAND2X1_631/A 0.03fF
C63646 PAND2X1_796/B POR2X1_72/B 0.01fF
C63647 POR2X1_629/CTRL POR2X1_629/B 0.01fF
C63648 PAND2X1_109/a_76_28# POR2X1_854/B 0.03fF
C63649 PAND2X1_643/A PAND2X1_538/CTRL 0.01fF
C63650 POR2X1_814/a_56_344# POR2X1_790/B 0.00fF
C63651 PAND2X1_454/B POR2X1_72/B 0.01fF
C63652 PAND2X1_93/B POR2X1_121/B 0.10fF
C63653 POR2X1_612/A POR2X1_293/Y 0.01fF
C63654 PAND2X1_651/Y POR2X1_386/Y 0.03fF
C63655 POR2X1_54/Y PAND2X1_23/O 0.05fF
C63656 POR2X1_329/A INPUT_5 0.00fF
C63657 POR2X1_257/A POR2X1_427/Y 0.03fF
C63658 POR2X1_76/B POR2X1_532/A 0.03fF
C63659 PAND2X1_624/O POR2X1_20/B 0.05fF
C63660 POR2X1_479/B POR2X1_288/O 0.01fF
C63661 PAND2X1_223/B POR2X1_283/O 0.00fF
C63662 PAND2X1_860/A POR2X1_73/Y 0.43fF
C63663 PAND2X1_717/A POR2X1_372/Y 0.00fF
C63664 PAND2X1_72/A POR2X1_141/A 0.01fF
C63665 POR2X1_788/A POR2X1_66/A 0.04fF
C63666 POR2X1_846/Y POR2X1_790/CTRL2 0.01fF
C63667 POR2X1_541/B VDD 0.14fF
C63668 PAND2X1_798/Y PAND2X1_354/Y 1.68fF
C63669 POR2X1_856/B POR2X1_467/Y 0.03fF
C63670 POR2X1_610/O PAND2X1_41/B 0.01fF
C63671 POR2X1_597/Y INPUT_0 0.00fF
C63672 POR2X1_23/Y POR2X1_72/B 0.23fF
C63673 POR2X1_811/A POR2X1_783/CTRL2 0.00fF
C63674 POR2X1_69/A D_INPUT_0 0.01fF
C63675 POR2X1_49/CTRL2 POR2X1_409/B 0.03fF
C63676 PAND2X1_340/B PAND2X1_340/a_16_344# 0.01fF
C63677 POR2X1_241/Y POR2X1_776/A 0.07fF
C63678 POR2X1_78/A POR2X1_121/B 0.03fF
C63679 POR2X1_837/B PAND2X1_505/CTRL2 0.02fF
C63680 POR2X1_67/Y POR2X1_619/a_56_344# 0.00fF
C63681 POR2X1_266/a_16_28# PAND2X1_41/B 0.01fF
C63682 POR2X1_478/O POR2X1_480/A 0.04fF
C63683 PAND2X1_142/CTRL2 PAND2X1_72/A 0.01fF
C63684 PAND2X1_404/Y PAND2X1_499/Y 0.41fF
C63685 PAND2X1_23/Y POR2X1_287/A 0.23fF
C63686 POR2X1_354/O POR2X1_356/B 0.01fF
C63687 POR2X1_848/Y VDD 0.09fF
C63688 POR2X1_49/Y POR2X1_626/O 0.09fF
C63689 POR2X1_60/A POR2X1_14/Y 0.08fF
C63690 POR2X1_24/CTRL2 POR2X1_29/A 0.01fF
C63691 POR2X1_291/CTRL2 POR2X1_825/Y 0.00fF
C63692 POR2X1_456/O POR2X1_66/A 0.01fF
C63693 POR2X1_625/CTRL2 POR2X1_37/Y 0.00fF
C63694 POR2X1_60/A PAND2X1_453/A 0.05fF
C63695 PAND2X1_73/Y PAND2X1_278/CTRL 0.00fF
C63696 POR2X1_32/A PAND2X1_733/a_16_344# 0.02fF
C63697 PAND2X1_603/m4_208_n4# POR2X1_750/B 0.08fF
C63698 PAND2X1_436/a_76_28# PAND2X1_499/Y 0.01fF
C63699 PAND2X1_644/Y VDD 0.15fF
C63700 POR2X1_548/O POR2X1_66/A 0.05fF
C63701 POR2X1_37/Y POR2X1_511/Y 0.00fF
C63702 POR2X1_294/A PAND2X1_72/A 0.06fF
C63703 PAND2X1_262/O POR2X1_296/B 0.01fF
C63704 PAND2X1_622/O POR2X1_669/B 0.04fF
C63705 POR2X1_119/Y PAND2X1_339/m4_208_n4# 0.04fF
C63706 POR2X1_376/B POR2X1_29/A 0.14fF
C63707 PAND2X1_716/B PAND2X1_332/Y 22.29fF
C63708 PAND2X1_797/Y POR2X1_77/Y 0.03fF
C63709 POR2X1_866/O POR2X1_750/B 0.01fF
C63710 POR2X1_191/Y PAND2X1_52/B 0.05fF
C63711 POR2X1_20/B POR2X1_396/O 0.01fF
C63712 POR2X1_41/B PAND2X1_267/Y 2.36fF
C63713 POR2X1_567/B POR2X1_244/B 0.05fF
C63714 POR2X1_296/B POR2X1_5/Y 0.16fF
C63715 POR2X1_498/O PAND2X1_205/A 0.00fF
C63716 POR2X1_672/A POR2X1_672/a_16_28# 0.10fF
C63717 POR2X1_32/A PAND2X1_473/B 0.03fF
C63718 PAND2X1_626/a_76_28# POR2X1_750/B 0.04fF
C63719 PAND2X1_208/CTRL POR2X1_40/Y 0.01fF
C63720 PAND2X1_571/A POR2X1_46/Y 0.03fF
C63721 POR2X1_856/B POR2X1_570/O 0.55fF
C63722 POR2X1_814/A POR2X1_725/Y 0.10fF
C63723 POR2X1_330/CTRL PAND2X1_52/B 0.01fF
C63724 PAND2X1_776/Y POR2X1_7/B 0.00fF
C63725 PAND2X1_268/m4_208_n4# POR2X1_193/A 0.09fF
C63726 PAND2X1_464/B PAND2X1_785/a_76_28# 0.02fF
C63727 POR2X1_192/Y POR2X1_220/B 0.07fF
C63728 PAND2X1_65/B POR2X1_811/B 0.03fF
C63729 POR2X1_294/Y POR2X1_220/Y 0.00fF
C63730 PAND2X1_48/B POR2X1_632/O 0.01fF
C63731 POR2X1_850/B POR2X1_362/B 0.33fF
C63732 PAND2X1_215/CTRL2 PAND2X1_723/Y 0.00fF
C63733 PAND2X1_619/a_16_344# PAND2X1_69/A 0.02fF
C63734 POR2X1_48/O POR2X1_60/A 0.01fF
C63735 PAND2X1_23/Y PAND2X1_827/CTRL 0.01fF
C63736 POR2X1_41/B POR2X1_674/a_16_28# 0.02fF
C63737 PAND2X1_659/O POR2X1_498/Y 0.03fF
C63738 POR2X1_675/a_16_28# POR2X1_675/A 0.10fF
C63739 POR2X1_43/B PAND2X1_477/CTRL 0.01fF
C63740 PAND2X1_6/Y PAND2X1_27/O 0.03fF
C63741 POR2X1_83/B PAND2X1_435/CTRL2 0.03fF
C63742 POR2X1_186/Y POR2X1_798/O 0.11fF
C63743 POR2X1_855/CTRL2 POR2X1_803/A 0.01fF
C63744 POR2X1_428/Y POR2X1_90/Y 0.00fF
C63745 PAND2X1_57/B PAND2X1_591/m4_208_n4# 0.07fF
C63746 PAND2X1_56/Y PAND2X1_93/B 0.05fF
C63747 PAND2X1_462/B D_INPUT_0 0.08fF
C63748 POR2X1_43/B POR2X1_118/Y 0.03fF
C63749 POR2X1_88/A POR2X1_7/A 0.02fF
C63750 PAND2X1_65/B POR2X1_254/O 0.18fF
C63751 POR2X1_66/B VDD 2.06fF
C63752 POR2X1_52/A POR2X1_29/A 0.03fF
C63753 PAND2X1_6/Y POR2X1_866/A 0.05fF
C63754 POR2X1_72/B PAND2X1_558/O 0.07fF
C63755 POR2X1_60/A PAND2X1_598/CTRL 0.01fF
C63756 PAND2X1_863/O PAND2X1_805/A 0.02fF
C63757 PAND2X1_784/CTRL POR2X1_32/A 0.01fF
C63758 PAND2X1_61/O POR2X1_55/Y 0.27fF
C63759 POR2X1_864/A POR2X1_598/CTRL2 0.00fF
C63760 POR2X1_49/Y POR2X1_58/O 0.18fF
C63761 POR2X1_610/CTRL2 POR2X1_532/A 0.07fF
C63762 POR2X1_41/B PAND2X1_215/O 0.06fF
C63763 POR2X1_814/A POR2X1_559/A 0.14fF
C63764 POR2X1_188/A VDD 1.08fF
C63765 PAND2X1_287/O PAND2X1_577/Y 0.02fF
C63766 PAND2X1_39/B POR2X1_780/B 0.59fF
C63767 POR2X1_16/A PAND2X1_201/CTRL 0.00fF
C63768 POR2X1_71/Y POR2X1_497/CTRL 0.07fF
C63769 POR2X1_863/O PAND2X1_73/Y 0.01fF
C63770 POR2X1_76/m4_208_n4# POR2X1_724/A 0.01fF
C63771 PAND2X1_333/CTRL2 VDD 0.00fF
C63772 POR2X1_62/m4_208_n4# PAND2X1_28/m4_208_n4# 0.05fF
C63773 PAND2X1_82/Y PAND2X1_39/B 0.04fF
C63774 POR2X1_5/Y POR2X1_236/Y 0.17fF
C63775 POR2X1_611/O VDD 0.00fF
C63776 POR2X1_97/A POR2X1_562/B 0.02fF
C63777 POR2X1_60/A POR2X1_55/Y 4.19fF
C63778 PAND2X1_480/B PAND2X1_579/CTRL 0.28fF
C63779 POR2X1_407/A POR2X1_656/O 0.02fF
C63780 POR2X1_344/O POR2X1_344/A 0.01fF
C63781 PAND2X1_20/A POR2X1_231/a_56_344# 0.00fF
C63782 POR2X1_13/Y POR2X1_102/Y 0.02fF
C63783 POR2X1_155/a_16_28# POR2X1_467/Y 0.03fF
C63784 POR2X1_78/A POR2X1_795/B 0.10fF
C63785 PAND2X1_56/Y POR2X1_78/A 0.03fF
C63786 POR2X1_5/Y POR2X1_547/B 0.00fF
C63787 PAND2X1_473/B PAND2X1_741/B 2.46fF
C63788 POR2X1_376/Y VDD 0.17fF
C63789 PAND2X1_49/O POR2X1_29/A 0.01fF
C63790 POR2X1_174/B D_GATE_741 0.02fF
C63791 POR2X1_857/a_16_28# POR2X1_579/Y 0.01fF
C63792 POR2X1_316/Y POR2X1_677/Y 0.03fF
C63793 PAND2X1_693/O PAND2X1_20/A 0.07fF
C63794 POR2X1_614/A POR2X1_450/O 0.01fF
C63795 POR2X1_43/B PAND2X1_573/B 0.03fF
C63796 POR2X1_692/O POR2X1_526/Y 0.01fF
C63797 PAND2X1_577/Y PAND2X1_578/A 0.13fF
C63798 POR2X1_422/CTRL2 POR2X1_7/A 0.09fF
C63799 POR2X1_315/Y PAND2X1_444/CTRL2 0.05fF
C63800 PAND2X1_550/CTRL VDD 0.00fF
C63801 PAND2X1_599/CTRL2 POR2X1_330/Y 0.31fF
C63802 POR2X1_68/A PAND2X1_58/A 0.77fF
C63803 PAND2X1_816/a_56_28# POR2X1_634/A 0.00fF
C63804 POR2X1_387/CTRL POR2X1_386/Y 0.00fF
C63805 POR2X1_830/CTRL POR2X1_741/Y 0.00fF
C63806 PAND2X1_57/B POR2X1_830/A 0.01fF
C63807 POR2X1_66/B POR2X1_741/Y 0.08fF
C63808 POR2X1_49/Y PAND2X1_523/O 0.17fF
C63809 PAND2X1_741/O PAND2X1_473/B 0.05fF
C63810 POR2X1_525/CTRL2 POR2X1_763/Y 0.05fF
C63811 POR2X1_525/O POR2X1_46/Y 0.01fF
C63812 PAND2X1_36/CTRL D_INPUT_6 0.01fF
C63813 POR2X1_502/A POR2X1_663/CTRL 0.01fF
C63814 POR2X1_673/A INPUT_0 0.00fF
C63815 POR2X1_383/A PAND2X1_93/B 2.20fF
C63816 PAND2X1_470/CTRL2 POR2X1_83/B 0.00fF
C63817 POR2X1_315/a_16_28# POR2X1_32/A 0.01fF
C63818 POR2X1_525/Y GATE_479 0.03fF
C63819 PAND2X1_556/B VDD 0.71fF
C63820 POR2X1_78/B POR2X1_244/B 0.05fF
C63821 PAND2X1_192/Y PAND2X1_592/Y 0.01fF
C63822 PAND2X1_287/Y PAND2X1_578/O 0.15fF
C63823 POR2X1_66/B POR2X1_389/a_16_28# 0.02fF
C63824 POR2X1_465/B POR2X1_563/CTRL2 0.00fF
C63825 PAND2X1_787/Y PAND2X1_592/a_16_344# 0.06fF
C63826 POR2X1_590/A POR2X1_206/CTRL 0.01fF
C63827 POR2X1_188/A POR2X1_741/Y 0.02fF
C63828 POR2X1_81/Y POR2X1_5/Y 0.00fF
C63829 PAND2X1_65/B PAND2X1_176/CTRL 0.01fF
C63830 POR2X1_221/a_16_28# POR2X1_220/Y 0.00fF
C63831 POR2X1_45/Y POR2X1_423/Y 0.00fF
C63832 PAND2X1_593/a_16_344# INPUT_0 0.01fF
C63833 POR2X1_859/A VDD 0.87fF
C63834 PAND2X1_65/B POR2X1_783/B 0.01fF
C63835 POR2X1_260/B POR2X1_773/B 0.02fF
C63836 PAND2X1_433/CTRL POR2X1_807/A 0.01fF
C63837 POR2X1_807/A POR2X1_733/A 0.03fF
C63838 POR2X1_460/A PAND2X1_58/A 0.02fF
C63839 PAND2X1_13/CTRL POR2X1_222/Y 0.00fF
C63840 POR2X1_108/CTRL POR2X1_102/Y 0.01fF
C63841 POR2X1_511/Y POR2X1_293/Y 0.07fF
C63842 PAND2X1_267/Y POR2X1_385/a_56_344# 0.00fF
C63843 POR2X1_615/CTRL2 PAND2X1_6/A 0.03fF
C63844 POR2X1_66/B PAND2X1_32/B 8.84fF
C63845 PAND2X1_653/CTRL2 POR2X1_329/A 0.00fF
C63846 POR2X1_114/CTRL POR2X1_777/B 0.26fF
C63847 POR2X1_278/Y PAND2X1_735/Y 2.13fF
C63848 PAND2X1_88/CTRL2 POR2X1_68/B 0.03fF
C63849 PAND2X1_254/Y VDD 0.01fF
C63850 PAND2X1_793/Y PAND2X1_580/B 3.77fF
C63851 POR2X1_43/B PAND2X1_849/CTRL 0.01fF
C63852 PAND2X1_63/Y POR2X1_641/a_76_344# 0.03fF
C63853 POR2X1_16/A PAND2X1_590/CTRL 0.01fF
C63854 POR2X1_220/B POR2X1_568/Y 0.64fF
C63855 POR2X1_48/A PAND2X1_348/O 0.01fF
C63856 PAND2X1_382/O PAND2X1_381/Y 0.15fF
C63857 POR2X1_355/B POR2X1_566/A 0.07fF
C63858 INPUT_2 POR2X1_609/O 0.01fF
C63859 POR2X1_555/A D_GATE_741 0.02fF
C63860 PAND2X1_6/Y POR2X1_457/a_16_28# 0.03fF
C63861 POR2X1_805/B POR2X1_805/A 0.13fF
C63862 POR2X1_65/A PAND2X1_547/CTRL 0.01fF
C63863 POR2X1_188/A PAND2X1_32/B 0.03fF
C63864 POR2X1_189/Y PAND2X1_473/B 0.03fF
C63865 PAND2X1_341/B POR2X1_63/Y 0.75fF
C63866 POR2X1_590/A POR2X1_537/A 0.06fF
C63867 POR2X1_539/A POR2X1_590/A 0.00fF
C63868 POR2X1_383/A POR2X1_78/A 0.31fF
C63869 POR2X1_68/B POR2X1_750/B 0.07fF
C63870 POR2X1_488/Y VDD 0.03fF
C63871 PAND2X1_830/Y PAND2X1_137/Y 0.19fF
C63872 POR2X1_649/B POR2X1_476/O 0.02fF
C63873 POR2X1_16/A D_INPUT_0 0.06fF
C63874 POR2X1_259/CTRL2 POR2X1_555/B 0.01fF
C63875 POR2X1_220/Y POR2X1_554/Y 0.03fF
C63876 POR2X1_57/A PAND2X1_354/A 0.01fF
C63877 PAND2X1_771/Y PAND2X1_569/a_16_344# 0.07fF
C63878 POR2X1_41/B POR2X1_372/Y 0.19fF
C63879 PAND2X1_41/B PAND2X1_177/O 0.15fF
C63880 POR2X1_55/Y PAND2X1_515/CTRL2 0.00fF
C63881 POR2X1_419/Y POR2X1_239/Y 0.00fF
C63882 PAND2X1_763/O PAND2X1_762/Y -0.00fF
C63883 PAND2X1_20/A PAND2X1_82/Y 0.06fF
C63884 POR2X1_599/A VDD 1.95fF
C63885 POR2X1_496/Y POR2X1_260/A 0.09fF
C63886 POR2X1_378/Y PAND2X1_90/A 0.03fF
C63887 PAND2X1_140/CTRL2 POR2X1_387/Y 0.13fF
C63888 D_INPUT_3 PAND2X1_859/A 0.03fF
C63889 PAND2X1_592/O POR2X1_42/Y 0.03fF
C63890 D_GATE_366 POR2X1_502/A 0.00fF
C63891 POR2X1_344/CTRL2 POR2X1_383/A 0.06fF
C63892 POR2X1_502/A POR2X1_264/Y 0.05fF
C63893 POR2X1_603/O POR2X1_761/A 0.03fF
C63894 PAND2X1_7/O POR2X1_244/B 0.02fF
C63895 POR2X1_723/CTRL2 POR2X1_723/B 0.01fF
C63896 POR2X1_357/CTRL2 POR2X1_220/B 0.01fF
C63897 POR2X1_538/CTRL POR2X1_566/A 0.01fF
C63898 POR2X1_186/Y POR2X1_540/a_16_28# 0.03fF
C63899 PAND2X1_90/A POR2X1_7/B 0.03fF
C63900 POR2X1_750/B POR2X1_750/a_16_28# 0.07fF
C63901 POR2X1_596/A POR2X1_448/B 0.03fF
C63902 POR2X1_68/A POR2X1_435/Y 0.07fF
C63903 PAND2X1_340/B POR2X1_4/Y 0.03fF
C63904 POR2X1_208/A POR2X1_201/a_16_28# 0.03fF
C63905 POR2X1_37/Y POR2X1_129/Y 5.42fF
C63906 POR2X1_210/Y POR2X1_213/B 0.05fF
C63907 POR2X1_356/A POR2X1_340/O 0.11fF
C63908 PAND2X1_6/Y POR2X1_302/Y 0.02fF
C63909 INPUT_0 POR2X1_816/A 0.22fF
C63910 PAND2X1_309/CTRL2 POR2X1_68/A 0.01fF
C63911 POR2X1_52/A PAND2X1_506/O 0.01fF
C63912 POR2X1_462/B INPUT_0 0.03fF
C63913 POR2X1_842/O POR2X1_737/A 0.01fF
C63914 POR2X1_304/CTRL PAND2X1_454/B 0.01fF
C63915 D_INPUT_1 INPUT_0 0.63fF
C63916 PAND2X1_496/O PAND2X1_55/Y -0.00fF
C63917 PAND2X1_116/CTRL2 POR2X1_283/A 0.11fF
C63918 POR2X1_84/Y POR2X1_786/O 0.02fF
C63919 PAND2X1_161/Y VDD 0.18fF
C63920 PAND2X1_388/O POR2X1_236/Y 0.02fF
C63921 PAND2X1_56/CTRL POR2X1_804/A 0.30fF
C63922 POR2X1_294/B POR2X1_565/CTRL2 0.00fF
C63923 PAND2X1_3/O POR2X1_750/B 0.02fF
C63924 POR2X1_76/Y POR2X1_804/A 0.11fF
C63925 POR2X1_130/A POR2X1_791/B 0.04fF
C63926 POR2X1_859/A PAND2X1_32/B 0.03fF
C63927 POR2X1_72/B POR2X1_530/CTRL 0.04fF
C63928 PAND2X1_93/B POR2X1_788/CTRL 0.01fF
C63929 PAND2X1_8/Y PAND2X1_670/CTRL2 0.05fF
C63930 POR2X1_13/A POR2X1_417/CTRL 0.01fF
C63931 POR2X1_480/A PAND2X1_60/B 0.10fF
C63932 PAND2X1_334/CTRL POR2X1_42/Y 0.01fF
C63933 PAND2X1_91/CTRL2 POR2X1_169/A 0.03fF
C63934 PAND2X1_774/CTRL VDD 0.00fF
C63935 PAND2X1_140/A POR2X1_107/O 0.01fF
C63936 POR2X1_840/Y POR2X1_851/A 0.03fF
C63937 POR2X1_596/A PAND2X1_57/B 0.10fF
C63938 POR2X1_49/Y PAND2X1_155/a_16_344# 0.02fF
C63939 POR2X1_116/A PAND2X1_72/A 0.03fF
C63940 POR2X1_259/A POR2X1_260/A 0.01fF
C63941 POR2X1_288/O PAND2X1_48/A 0.06fF
C63942 POR2X1_407/A POR2X1_733/A 3.79fF
C63943 POR2X1_40/Y POR2X1_171/a_16_28# 0.03fF
C63944 PAND2X1_320/CTRL POR2X1_568/Y 0.01fF
C63945 POR2X1_63/Y PAND2X1_327/a_16_344# 0.03fF
C63946 POR2X1_97/A POR2X1_357/B 0.04fF
C63947 POR2X1_417/CTRL2 POR2X1_293/Y 0.01fF
C63948 PAND2X1_549/B POR2X1_372/O 0.01fF
C63949 POR2X1_96/Y POR2X1_37/Y 0.11fF
C63950 POR2X1_243/Y PAND2X1_60/B 0.07fF
C63951 PAND2X1_404/Y POR2X1_39/B 0.02fF
C63952 POR2X1_416/B POR2X1_77/CTRL2 0.21fF
C63953 PAND2X1_182/B POR2X1_40/Y 0.01fF
C63954 PAND2X1_710/CTRL POR2X1_701/Y 0.00fF
C63955 POR2X1_96/A D_INPUT_3 0.01fF
C63956 POR2X1_202/O POR2X1_507/A 0.03fF
C63957 POR2X1_41/B POR2X1_526/Y 0.05fF
C63958 POR2X1_804/A POR2X1_740/Y 0.10fF
C63959 POR2X1_562/a_76_344# POR2X1_562/B 0.00fF
C63960 POR2X1_730/B POR2X1_730/O 0.01fF
C63961 POR2X1_68/A POR2X1_782/A 0.00fF
C63962 POR2X1_60/A PAND2X1_199/B 0.02fF
C63963 PAND2X1_90/Y POR2X1_456/B 1.43fF
C63964 POR2X1_831/O POR2X1_717/B 0.01fF
C63965 POR2X1_52/A POR2X1_583/O 0.01fF
C63966 PAND2X1_175/CTRL2 VDD 0.00fF
C63967 PAND2X1_738/Y PAND2X1_181/CTRL 0.28fF
C63968 POR2X1_84/CTRL POR2X1_532/A 0.01fF
C63969 POR2X1_373/Y PAND2X1_731/B 0.02fF
C63970 PAND2X1_442/m4_208_n4# POR2X1_568/Y 0.06fF
C63971 POR2X1_78/A POR2X1_788/CTRL 0.09fF
C63972 POR2X1_57/A PAND2X1_724/B 0.05fF
C63973 PAND2X1_675/A POR2X1_90/Y 0.01fF
C63974 POR2X1_832/A POR2X1_513/B 0.03fF
C63975 POR2X1_496/Y PAND2X1_508/B 0.04fF
C63976 PAND2X1_862/B PAND2X1_510/B 1.67fF
C63977 POR2X1_547/B POR2X1_6/CTRL2 0.01fF
C63978 POR2X1_740/Y PAND2X1_306/CTRL2 0.00fF
C63979 POR2X1_789/A PAND2X1_69/A 0.03fF
C63980 PAND2X1_48/B POR2X1_359/Y 0.01fF
C63981 POR2X1_43/B PAND2X1_341/A 0.10fF
C63982 POR2X1_68/A PAND2X1_96/B 3.67fF
C63983 PAND2X1_90/A PAND2X1_60/B 0.03fF
C63984 PAND2X1_674/CTRL2 PAND2X1_60/B 0.00fF
C63985 POR2X1_271/A POR2X1_5/Y 0.02fF
C63986 POR2X1_41/B POR2X1_83/CTRL2 0.00fF
C63987 POR2X1_614/A PAND2X1_69/A 32.67fF
C63988 PAND2X1_440/O POR2X1_23/Y 0.01fF
C63989 PAND2X1_442/a_16_344# POR2X1_444/Y 0.01fF
C63990 POR2X1_866/A PAND2X1_52/B 0.05fF
C63991 PAND2X1_744/O POR2X1_532/A 0.01fF
C63992 PAND2X1_587/Y POR2X1_260/A 0.03fF
C63993 POR2X1_89/a_16_28# PAND2X1_333/Y 0.03fF
C63994 POR2X1_394/A PAND2X1_713/B 0.00fF
C63995 POR2X1_208/A POR2X1_208/a_16_28# 0.02fF
C63996 POR2X1_43/B POR2X1_91/Y 0.59fF
C63997 PAND2X1_56/Y PAND2X1_306/O 0.01fF
C63998 PAND2X1_428/m4_208_n4# PAND2X1_48/A 0.04fF
C63999 POR2X1_30/O POR2X1_3/A 0.02fF
C64000 INPUT_6 PAND2X1_587/CTRL 0.01fF
C64001 POR2X1_249/Y POR2X1_784/A 0.03fF
C64002 POR2X1_516/A POR2X1_55/Y 0.01fF
C64003 POR2X1_38/B PAND2X1_69/A 0.39fF
C64004 INPUT_1 POR2X1_669/CTRL2 0.12fF
C64005 PAND2X1_108/CTRL POR2X1_646/Y 0.01fF
C64006 PAND2X1_696/a_16_344# POR2X1_811/B 0.02fF
C64007 POR2X1_37/Y PAND2X1_333/Y 0.04fF
C64008 POR2X1_309/O POR2X1_39/B 0.01fF
C64009 POR2X1_416/B POR2X1_420/a_16_28# 0.03fF
C64010 PAND2X1_473/Y POR2X1_394/A 0.03fF
C64011 POR2X1_207/A POR2X1_195/O 0.01fF
C64012 PAND2X1_63/Y POR2X1_84/Y 0.08fF
C64013 POR2X1_822/Y POR2X1_821/Y 0.02fF
C64014 PAND2X1_55/Y POR2X1_576/CTRL2 0.04fF
C64015 POR2X1_863/A POR2X1_446/O 0.02fF
C64016 PAND2X1_847/CTRL2 POR2X1_32/A 0.04fF
C64017 PAND2X1_438/CTRL2 POR2X1_544/B 0.02fF
C64018 PAND2X1_6/Y POR2X1_774/CTRL2 0.00fF
C64019 POR2X1_281/O PAND2X1_809/A 0.01fF
C64020 POR2X1_390/B POR2X1_717/Y 0.00fF
C64021 PAND2X1_651/Y POR2X1_239/Y 0.20fF
C64022 PAND2X1_785/CTRL POR2X1_91/Y 0.11fF
C64023 POR2X1_93/A POR2X1_38/B 1.14fF
C64024 POR2X1_78/B POR2X1_537/Y 0.03fF
C64025 POR2X1_65/A POR2X1_760/Y 0.01fF
C64026 PAND2X1_474/Y PAND2X1_716/B 0.03fF
C64027 POR2X1_865/B POR2X1_113/Y 0.19fF
C64028 POR2X1_54/Y POR2X1_9/Y 0.40fF
C64029 POR2X1_674/Y POR2X1_331/CTRL2 0.01fF
C64030 POR2X1_538/a_16_28# POR2X1_538/A 0.03fF
C64031 POR2X1_7/B PAND2X1_853/B 0.16fF
C64032 POR2X1_538/O POR2X1_703/A 0.03fF
C64033 PAND2X1_216/B PAND2X1_652/A 0.03fF
C64034 POR2X1_383/A POR2X1_784/CTRL 0.00fF
C64035 POR2X1_532/A POR2X1_215/Y 0.01fF
C64036 POR2X1_356/A POR2X1_334/Y 0.10fF
C64037 POR2X1_129/Y POR2X1_293/Y 0.09fF
C64038 POR2X1_13/A PAND2X1_716/B 26.21fF
C64039 POR2X1_145/O POR2X1_394/A 0.01fF
C64040 PAND2X1_6/Y POR2X1_703/A 0.02fF
C64041 PAND2X1_358/A PAND2X1_101/CTRL2 0.05fF
C64042 PAND2X1_553/B POR2X1_183/CTRL2 0.03fF
C64043 PAND2X1_730/B PAND2X1_643/A 0.08fF
C64044 POR2X1_790/A POR2X1_260/A 0.03fF
C64045 POR2X1_180/B PAND2X1_96/B 0.03fF
C64046 D_INPUT_3 POR2X1_7/A 0.03fF
C64047 POR2X1_828/A POR2X1_598/O 0.01fF
C64048 PAND2X1_297/O PAND2X1_69/A 0.01fF
C64049 PAND2X1_724/CTRL2 PAND2X1_714/Y 0.01fF
C64050 POR2X1_187/Y POR2X1_96/A 0.07fF
C64051 POR2X1_38/Y PAND2X1_121/O 0.01fF
C64052 POR2X1_638/A PAND2X1_72/A 0.01fF
C64053 POR2X1_83/Y POR2X1_96/A 0.02fF
C64054 POR2X1_317/a_16_28# POR2X1_317/B -0.00fF
C64055 PAND2X1_403/CTRL2 POR2X1_37/Y 0.08fF
C64056 PAND2X1_835/O POR2X1_394/A 0.05fF
C64057 POR2X1_242/O PAND2X1_52/B 0.01fF
C64058 VDD POR2X1_199/B 0.10fF
C64059 POR2X1_687/Y POR2X1_855/B 0.00fF
C64060 POR2X1_12/A POR2X1_18/CTRL2 0.01fF
C64061 D_INPUT_5 POR2X1_18/CTRL 0.02fF
C64062 PAND2X1_659/Y POR2X1_293/Y 0.03fF
C64063 PAND2X1_23/Y POR2X1_507/B 0.01fF
C64064 POR2X1_48/A PAND2X1_635/Y 0.35fF
C64065 POR2X1_327/Y POR2X1_149/B 0.03fF
C64066 PAND2X1_675/A PAND2X1_360/Y 0.03fF
C64067 PAND2X1_48/B POR2X1_359/CTRL 0.01fF
C64068 PAND2X1_23/Y POR2X1_359/CTRL2 0.01fF
C64069 POR2X1_135/O POR2X1_46/Y 0.25fF
C64070 POR2X1_491/Y PAND2X1_84/Y 0.05fF
C64071 POR2X1_596/A POR2X1_771/A 0.03fF
C64072 POR2X1_865/B POR2X1_260/A 0.03fF
C64073 PAND2X1_88/Y POR2X1_260/A 0.07fF
C64074 PAND2X1_723/A PAND2X1_656/A 1.57fF
C64075 POR2X1_578/a_16_28# POR2X1_577/Y 0.04fF
C64076 POR2X1_150/Y POR2X1_20/B 0.00fF
C64077 PAND2X1_824/B POR2X1_38/B 0.01fF
C64078 POR2X1_184/Y POR2X1_131/A 0.02fF
C64079 POR2X1_346/B PAND2X1_60/B 0.03fF
C64080 PAND2X1_48/B POR2X1_552/A 0.01fF
C64081 INPUT_1 POR2X1_387/Y 0.16fF
C64082 PAND2X1_93/B PAND2X1_86/CTRL2 0.01fF
C64083 PAND2X1_732/A PAND2X1_731/A 0.09fF
C64084 POR2X1_203/Y POR2X1_186/B 0.02fF
C64085 PAND2X1_93/B POR2X1_648/Y 0.07fF
C64086 PAND2X1_864/a_16_344# PAND2X1_568/B 0.01fF
C64087 POR2X1_92/O POR2X1_8/Y 0.16fF
C64088 PAND2X1_310/O POR2X1_501/B 0.02fF
C64089 POR2X1_616/Y PAND2X1_6/A 0.03fF
C64090 PAND2X1_63/B POR2X1_376/CTRL 0.01fF
C64091 PAND2X1_73/Y POR2X1_846/A 0.03fF
C64092 POR2X1_614/A POR2X1_512/CTRL 0.00fF
C64093 POR2X1_119/Y PAND2X1_642/B 0.12fF
C64094 PAND2X1_658/A PAND2X1_860/CTRL2 0.01fF
C64095 PAND2X1_785/CTRL POR2X1_109/Y 0.01fF
C64096 PAND2X1_860/A PAND2X1_360/a_16_344# 0.01fF
C64097 POR2X1_387/Y POR2X1_153/Y 0.10fF
C64098 POR2X1_451/A POR2X1_750/B 3.07fF
C64099 POR2X1_727/O POR2X1_353/A 0.16fF
C64100 POR2X1_375/CTRL POR2X1_260/A 0.03fF
C64101 PAND2X1_26/O PAND2X1_18/B 0.02fF
C64102 POR2X1_71/Y PAND2X1_501/CTRL 0.09fF
C64103 POR2X1_188/a_16_28# POR2X1_675/Y 0.02fF
C64104 POR2X1_408/Y POR2X1_129/Y 0.03fF
C64105 PAND2X1_79/Y PAND2X1_527/O 0.01fF
C64106 PAND2X1_290/O PAND2X1_55/Y 0.01fF
C64107 PAND2X1_659/Y PAND2X1_676/CTRL2 0.00fF
C64108 POR2X1_394/A POR2X1_765/Y 0.03fF
C64109 POR2X1_203/CTRL PAND2X1_48/A 0.02fF
C64110 POR2X1_372/Y POR2X1_77/Y 0.50fF
C64111 POR2X1_445/A POR2X1_341/A 0.02fF
C64112 POR2X1_518/O POR2X1_518/Y 0.00fF
C64113 PAND2X1_48/B POR2X1_342/A 0.04fF
C64114 POR2X1_38/Y PAND2X1_737/CTRL2 0.00fF
C64115 PAND2X1_39/B POR2X1_647/CTRL2 0.01fF
C64116 POR2X1_78/A POR2X1_648/Y 0.03fF
C64117 POR2X1_692/O POR2X1_485/Y 0.18fF
C64118 POR2X1_725/Y POR2X1_151/Y 0.02fF
C64119 POR2X1_73/Y PAND2X1_860/CTRL2 0.00fF
C64120 POR2X1_439/Y PAND2X1_437/O 0.01fF
C64121 POR2X1_96/A POR2X1_759/O 0.01fF
C64122 PAND2X1_338/B PAND2X1_338/CTRL2 0.07fF
C64123 POR2X1_123/CTRL2 PAND2X1_72/A 0.02fF
C64124 POR2X1_74/CTRL POR2X1_271/A 0.04fF
C64125 PAND2X1_501/O PAND2X1_575/A 0.02fF
C64126 POR2X1_334/Y POR2X1_97/CTRL 0.08fF
C64127 POR2X1_519/Y POR2X1_77/Y 0.03fF
C64128 PAND2X1_860/A PAND2X1_804/A 0.00fF
C64129 POR2X1_44/a_56_344# PAND2X1_635/Y 0.00fF
C64130 POR2X1_83/Y POR2X1_7/A 0.02fF
C64131 POR2X1_101/Y PAND2X1_48/A 0.22fF
C64132 POR2X1_23/Y PAND2X1_407/CTRL2 0.03fF
C64133 POR2X1_383/CTRL2 POR2X1_520/A 0.01fF
C64134 PAND2X1_565/A POR2X1_39/B 0.01fF
C64135 PAND2X1_96/B POR2X1_169/A 0.03fF
C64136 PAND2X1_41/CTRL POR2X1_66/A 0.01fF
C64137 PAND2X1_73/Y POR2X1_705/B 0.03fF
C64138 POR2X1_340/O PAND2X1_72/A 0.02fF
C64139 POR2X1_84/A POR2X1_240/O 0.01fF
C64140 PAND2X1_483/CTRL PAND2X1_508/Y 0.00fF
C64141 POR2X1_861/CTRL2 PAND2X1_72/A 0.01fF
C64142 POR2X1_253/Y POR2X1_77/Y 0.05fF
C64143 PAND2X1_462/O PAND2X1_472/A 0.02fF
C64144 POR2X1_119/Y PAND2X1_550/B 0.03fF
C64145 PAND2X1_860/A PAND2X1_785/Y 0.03fF
C64146 PAND2X1_372/m4_208_n4# POR2X1_717/B 0.01fF
C64147 POR2X1_319/A POR2X1_567/B 0.05fF
C64148 POR2X1_73/Y PAND2X1_339/O 0.07fF
C64149 POR2X1_775/A POR2X1_568/A 0.05fF
C64150 POR2X1_76/A POR2X1_66/A 0.03fF
C64151 PAND2X1_437/O POR2X1_192/Y 0.17fF
C64152 POR2X1_36/B POR2X1_39/B 0.29fF
C64153 PAND2X1_206/B PAND2X1_340/CTRL2 0.00fF
C64154 POR2X1_491/CTRL2 POR2X1_150/Y 0.01fF
C64155 PAND2X1_773/Y PAND2X1_771/Y 0.23fF
C64156 PAND2X1_63/B PAND2X1_529/CTRL2 0.01fF
C64157 POR2X1_137/B POR2X1_634/O 0.14fF
C64158 PAND2X1_809/B PAND2X1_854/A 0.02fF
C64159 PAND2X1_403/CTRL2 POR2X1_293/Y 0.00fF
C64160 POR2X1_610/m4_208_n4# POR2X1_862/A 0.01fF
C64161 POR2X1_709/A PAND2X1_58/A 0.05fF
C64162 PAND2X1_60/B POR2X1_716/CTRL 0.00fF
C64163 POR2X1_265/Y PAND2X1_560/B 0.03fF
C64164 POR2X1_71/a_56_344# POR2X1_62/Y 0.00fF
C64165 POR2X1_394/A POR2X1_7/Y 0.03fF
C64166 POR2X1_428/Y POR2X1_430/Y 0.01fF
C64167 POR2X1_271/B POR2X1_423/Y 0.00fF
C64168 POR2X1_378/CTRL2 PAND2X1_9/Y 0.01fF
C64169 POR2X1_359/O POR2X1_363/A 0.25fF
C64170 POR2X1_825/Y PAND2X1_334/O 0.00fF
C64171 POR2X1_389/A PAND2X1_72/A 0.12fF
C64172 POR2X1_632/B POR2X1_632/O 0.02fF
C64173 POR2X1_774/CTRL2 PAND2X1_52/B 0.03fF
C64174 POR2X1_849/A D_INPUT_0 0.03fF
C64175 PAND2X1_617/O VDD 0.00fF
C64176 PAND2X1_23/Y POR2X1_837/B 0.13fF
C64177 POR2X1_568/B POR2X1_260/A 0.05fF
C64178 PAND2X1_761/O POR2X1_750/B 0.02fF
C64179 POR2X1_101/Y POR2X1_514/m4_208_n4# 0.03fF
C64180 PAND2X1_806/CTRL PAND2X1_362/A 0.01fF
C64181 PAND2X1_3/A PAND2X1_36/O 0.02fF
C64182 POR2X1_416/B PAND2X1_514/CTRL 0.01fF
C64183 PAND2X1_492/CTRL2 POR2X1_556/A 0.01fF
C64184 POR2X1_477/CTRL POR2X1_480/A 0.08fF
C64185 POR2X1_568/A POR2X1_162/Y 0.03fF
C64186 POR2X1_376/Y PAND2X1_9/Y 0.02fF
C64187 POR2X1_814/A POR2X1_783/B 0.22fF
C64188 POR2X1_48/A POR2X1_394/Y 0.20fF
C64189 POR2X1_66/B POR2X1_818/Y 0.56fF
C64190 POR2X1_567/B POR2X1_439/CTRL2 0.18fF
C64191 POR2X1_441/Y VDD 0.56fF
C64192 PAND2X1_9/CTRL D_INPUT_0 0.05fF
C64193 POR2X1_137/B INPUT_0 0.10fF
C64194 POR2X1_450/CTRL2 POR2X1_121/B 0.05fF
C64195 POR2X1_848/A POR2X1_750/B 0.07fF
C64196 POR2X1_24/Y POR2X1_5/Y 0.04fF
C64197 PAND2X1_817/CTRL2 PAND2X1_381/Y 0.00fF
C64198 POR2X1_41/B POR2X1_485/Y 0.03fF
C64199 INPUT_3 INPUT_0 0.10fF
C64200 POR2X1_126/m4_208_n4# POR2X1_94/A 0.12fF
C64201 POR2X1_456/B POR2X1_715/O 0.09fF
C64202 PAND2X1_818/O POR2X1_411/B 0.07fF
C64203 PAND2X1_437/CTRL2 PAND2X1_60/B 0.00fF
C64204 PAND2X1_416/CTRL VDD -0.00fF
C64205 POR2X1_41/B PAND2X1_838/CTRL 0.01fF
C64206 POR2X1_83/B PAND2X1_721/B 0.01fF
C64207 POR2X1_661/A PAND2X1_305/CTRL 0.03fF
C64208 PAND2X1_601/m4_208_n4# POR2X1_718/A 0.01fF
C64209 POR2X1_96/A PAND2X1_203/CTRL 0.04fF
C64210 PAND2X1_7/m4_208_n4# PAND2X1_257/m4_208_n4# 0.13fF
C64211 POR2X1_102/Y PAND2X1_219/A 0.09fF
C64212 POR2X1_78/B POR2X1_319/A 0.12fF
C64213 POR2X1_830/CTRL POR2X1_830/Y 0.01fF
C64214 POR2X1_502/A POR2X1_624/Y 1.54fF
C64215 PAND2X1_860/A PAND2X1_861/CTRL2 0.01fF
C64216 POR2X1_448/a_16_28# POR2X1_296/B 0.11fF
C64217 POR2X1_334/Y PAND2X1_72/A 0.12fF
C64218 POR2X1_66/B POR2X1_267/A 1.57fF
C64219 PAND2X1_73/Y POR2X1_780/CTRL 0.01fF
C64220 POR2X1_322/O POR2X1_441/Y 0.07fF
C64221 POR2X1_654/CTRL2 POR2X1_121/B 0.02fF
C64222 POR2X1_777/B POR2X1_296/B 0.10fF
C64223 PAND2X1_699/O PAND2X1_6/A 0.03fF
C64224 PAND2X1_796/B POR2X1_7/B 0.02fF
C64225 POR2X1_14/Y POR2X1_750/A 0.05fF
C64226 POR2X1_288/A POR2X1_288/O 0.00fF
C64227 POR2X1_188/A POR2X1_830/Y 0.01fF
C64228 POR2X1_93/Y INPUT_0 0.21fF
C64229 POR2X1_490/Y POR2X1_13/A 0.02fF
C64230 PAND2X1_93/B INPUT_0 0.04fF
C64231 POR2X1_306/Y POR2X1_14/Y 0.05fF
C64232 PAND2X1_219/B POR2X1_32/A 0.01fF
C64233 POR2X1_60/A PAND2X1_541/CTRL 0.01fF
C64234 POR2X1_306/Y PAND2X1_453/A 0.06fF
C64235 PAND2X1_466/A POR2X1_90/Y 0.02fF
C64236 PAND2X1_474/A PAND2X1_573/B 0.09fF
C64237 PAND2X1_304/CTRL PAND2X1_56/A 0.01fF
C64238 POR2X1_859/A POR2X1_818/Y 0.11fF
C64239 PAND2X1_65/B POR2X1_296/B 0.13fF
C64240 PAND2X1_201/CTRL2 PAND2X1_341/A 0.01fF
C64241 PAND2X1_242/Y POR2X1_129/Y 0.03fF
C64242 POR2X1_556/A POR2X1_786/Y 0.05fF
C64243 POR2X1_630/B POR2X1_510/Y 0.02fF
C64244 POR2X1_805/Y POR2X1_805/B 0.11fF
C64245 POR2X1_158/CTRL POR2X1_416/B 0.01fF
C64246 POR2X1_669/B PAND2X1_713/B 0.04fF
C64247 PAND2X1_20/A POR2X1_849/CTRL 0.01fF
C64248 POR2X1_68/A POR2X1_676/CTRL2 0.08fF
C64249 POR2X1_263/Y PAND2X1_734/B 0.00fF
C64250 PAND2X1_57/B D_INPUT_0 0.03fF
C64251 PAND2X1_234/O POR2X1_260/A 0.05fF
C64252 POR2X1_23/Y POR2X1_7/B 0.20fF
C64253 PAND2X1_852/A POR2X1_42/Y 0.99fF
C64254 PAND2X1_97/a_16_344# POR2X1_293/Y 0.01fF
C64255 PAND2X1_63/Y POR2X1_341/A 1.42fF
C64256 POR2X1_490/O POR2X1_73/Y 0.01fF
C64257 POR2X1_60/A POR2X1_511/Y 0.13fF
C64258 POR2X1_682/Y POR2X1_32/A 0.01fF
C64259 POR2X1_66/B POR2X1_472/Y 0.37fF
C64260 PAND2X1_48/B POR2X1_567/B 0.05fF
C64261 POR2X1_78/A INPUT_0 0.13fF
C64262 PAND2X1_73/Y POR2X1_465/A 0.01fF
C64263 PAND2X1_862/B POR2X1_29/A 0.00fF
C64264 POR2X1_37/Y POR2X1_293/Y 0.29fF
C64265 INPUT_2 POR2X1_54/Y 0.13fF
C64266 PAND2X1_657/O PAND2X1_659/B 0.00fF
C64267 POR2X1_198/O PAND2X1_93/B 0.19fF
C64268 PAND2X1_793/Y POR2X1_32/A 0.03fF
C64269 PAND2X1_58/A POR2X1_435/Y 0.07fF
C64270 POR2X1_114/B POR2X1_458/CTRL 0.12fF
C64271 POR2X1_355/B POR2X1_241/B 0.03fF
C64272 PAND2X1_794/a_76_28# PAND2X1_473/B 0.02fF
C64273 POR2X1_697/O POR2X1_40/Y 0.02fF
C64274 POR2X1_480/A POR2X1_750/B 0.07fF
C64275 PAND2X1_841/B POR2X1_32/A 0.03fF
C64276 PAND2X1_309/CTRL2 PAND2X1_58/A 0.01fF
C64277 POR2X1_814/B POR2X1_805/B 0.05fF
C64278 POR2X1_145/Y POR2X1_257/A 0.03fF
C64279 PAND2X1_267/Y POR2X1_52/Y 0.02fF
C64280 POR2X1_72/B POR2X1_372/A 0.01fF
C64281 POR2X1_674/a_16_28# PAND2X1_742/B 0.02fF
C64282 INPUT_1 POR2X1_624/B 0.22fF
C64283 POR2X1_76/A POR2X1_532/A 0.00fF
C64284 PAND2X1_23/Y POR2X1_792/O 0.06fF
C64285 POR2X1_448/B PAND2X1_90/Y 0.03fF
C64286 POR2X1_88/Y POR2X1_40/Y 0.03fF
C64287 POR2X1_78/B PAND2X1_597/CTRL2 0.02fF
C64288 POR2X1_66/B POR2X1_445/O 0.01fF
C64289 PAND2X1_223/CTRL VDD 0.00fF
C64290 POR2X1_458/CTRL POR2X1_458/B 0.04fF
C64291 POR2X1_482/O PAND2X1_6/A 0.05fF
C64292 POR2X1_236/O POR2X1_5/Y 0.02fF
C64293 PAND2X1_58/A PAND2X1_377/Y 0.01fF
C64294 PAND2X1_849/B POR2X1_20/B 0.05fF
C64295 POR2X1_115/O POR2X1_330/Y 0.07fF
C64296 POR2X1_196/O POR2X1_740/Y 0.04fF
C64297 PAND2X1_412/CTRL POR2X1_546/A 0.03fF
C64298 PAND2X1_833/O POR2X1_376/B 0.08fF
C64299 POR2X1_9/Y POR2X1_4/Y 0.03fF
C64300 PAND2X1_685/a_16_344# POR2X1_32/A 0.02fF
C64301 PAND2X1_192/Y PAND2X1_739/O 0.03fF
C64302 POR2X1_348/A POR2X1_244/B 0.10fF
C64303 POR2X1_61/Y POR2X1_215/CTRL2 0.03fF
C64304 POR2X1_220/Y PAND2X1_7/Y 0.01fF
C64305 POR2X1_811/A POR2X1_828/A 0.03fF
C64306 POR2X1_523/Y POR2X1_590/A 0.03fF
C64307 PAND2X1_805/A GATE_741 0.03fF
C64308 PAND2X1_812/a_76_28# PAND2X1_811/A 0.04fF
C64309 POR2X1_96/A PAND2X1_541/O 0.04fF
C64310 PAND2X1_213/Y POR2X1_438/Y 0.15fF
C64311 POR2X1_66/A POR2X1_540/A 0.03fF
C64312 PAND2X1_137/Y PAND2X1_220/Y 0.03fF
C64313 PAND2X1_65/CTRL POR2X1_205/A 0.06fF
C64314 D_INPUT_5 PAND2X1_1/a_16_344# 0.01fF
C64315 PAND2X1_818/O POR2X1_376/B 0.03fF
C64316 POR2X1_60/O D_INPUT_0 0.06fF
C64317 POR2X1_341/A POR2X1_260/A 0.07fF
C64318 PAND2X1_575/A PAND2X1_575/B 0.17fF
C64319 PAND2X1_540/O PAND2X1_553/B 0.11fF
C64320 POR2X1_312/Y POR2X1_7/B 0.00fF
C64321 POR2X1_740/Y POR2X1_794/B 0.03fF
C64322 POR2X1_40/Y POR2X1_743/Y 0.01fF
C64323 PAND2X1_50/O VDD 0.00fF
C64324 PAND2X1_387/O PAND2X1_386/Y 0.01fF
C64325 PAND2X1_57/B PAND2X1_90/Y 0.17fF
C64326 POR2X1_590/A PAND2X1_69/A 2.76fF
C64327 POR2X1_275/A POR2X1_129/Y 0.60fF
C64328 POR2X1_102/Y POR2X1_816/A 0.03fF
C64329 POR2X1_763/CTRL2 POR2X1_46/Y 0.01fF
C64330 PAND2X1_208/CTRL2 POR2X1_599/A 0.32fF
C64331 POR2X1_102/Y D_INPUT_1 0.01fF
C64332 POR2X1_257/A POR2X1_764/O 0.09fF
C64333 POR2X1_483/A POR2X1_483/a_56_344# 0.00fF
C64334 PAND2X1_116/O PAND2X1_115/Y 0.00fF
C64335 POR2X1_186/Y PAND2X1_145/CTRL 0.01fF
C64336 POR2X1_72/B PAND2X1_658/B 0.08fF
C64337 POR2X1_37/Y POR2X1_408/Y 0.01fF
C64338 POR2X1_306/CTRL2 POR2X1_102/Y 0.01fF
C64339 PAND2X1_96/B PAND2X1_58/A 2.71fF
C64340 PAND2X1_20/A POR2X1_139/a_76_344# 0.00fF
C64341 POR2X1_110/Y PAND2X1_466/A 0.00fF
C64342 POR2X1_257/A POR2X1_394/A 0.34fF
C64343 POR2X1_730/Y POR2X1_260/B 0.03fF
C64344 POR2X1_243/A PAND2X1_88/Y 0.12fF
C64345 POR2X1_625/Y VDD 0.24fF
C64346 POR2X1_832/B PAND2X1_589/CTRL2 0.01fF
C64347 POR2X1_539/A POR2X1_66/A 0.01fF
C64348 INPUT_1 POR2X1_422/CTRL2 0.01fF
C64349 POR2X1_463/Y POR2X1_805/CTRL 0.00fF
C64350 PAND2X1_425/Y PAND2X1_3/B 0.05fF
C64351 POR2X1_411/B PAND2X1_345/Y 0.02fF
C64352 PAND2X1_805/a_16_344# PAND2X1_793/Y 0.01fF
C64353 PAND2X1_661/CTRL2 POR2X1_13/A 0.00fF
C64354 PAND2X1_633/Y PAND2X1_640/B -0.01fF
C64355 POR2X1_43/B POR2X1_278/CTRL2 0.17fF
C64356 POR2X1_192/Y POR2X1_223/CTRL 0.01fF
C64357 POR2X1_221/CTRL2 POR2X1_221/Y 0.03fF
C64358 POR2X1_290/CTRL2 PAND2X1_642/B 0.01fF
C64359 POR2X1_273/CTRL POR2X1_153/Y 0.01fF
C64360 POR2X1_288/m4_208_n4# PAND2X1_32/B 0.08fF
C64361 POR2X1_657/CTRL POR2X1_228/Y 0.03fF
C64362 PAND2X1_287/CTRL2 VDD 0.00fF
C64363 POR2X1_300/CTRL2 POR2X1_272/Y 0.01fF
C64364 PAND2X1_803/Y POR2X1_83/B 0.04fF
C64365 PAND2X1_63/Y POR2X1_500/A 0.05fF
C64366 PAND2X1_216/B PAND2X1_205/A 0.03fF
C64367 PAND2X1_48/B PAND2X1_48/CTRL2 0.04fF
C64368 POR2X1_503/a_16_28# POR2X1_283/A 0.07fF
C64369 POR2X1_78/B PAND2X1_48/B 0.35fF
C64370 POR2X1_614/A PAND2X1_262/CTRL 0.06fF
C64371 POR2X1_178/CTRL PAND2X1_562/B 0.06fF
C64372 PAND2X1_715/O POR2X1_293/Y 0.03fF
C64373 POR2X1_809/A POR2X1_676/CTRL 0.01fF
C64374 POR2X1_67/Y POR2X1_39/B 0.06fF
C64375 POR2X1_444/O POR2X1_191/Y 0.01fF
C64376 POR2X1_654/a_16_28# POR2X1_651/Y 0.03fF
C64377 PAND2X1_567/CTRL VDD -0.00fF
C64378 PAND2X1_624/a_16_344# PAND2X1_623/Y 0.01fF
C64379 POR2X1_692/O PAND2X1_726/B 0.03fF
C64380 PAND2X1_46/O POR2X1_68/B 0.17fF
C64381 POR2X1_57/A PAND2X1_733/A -0.00fF
C64382 POR2X1_102/Y PAND2X1_854/A 0.07fF
C64383 POR2X1_13/A PAND2X1_243/B 0.03fF
C64384 POR2X1_362/Y POR2X1_383/A 0.52fF
C64385 POR2X1_516/Y PAND2X1_349/A 0.03fF
C64386 POR2X1_383/A POR2X1_285/Y 0.03fF
C64387 POR2X1_68/B POR2X1_389/Y 0.03fF
C64388 POR2X1_83/B POR2X1_235/Y 0.00fF
C64389 POR2X1_481/a_16_28# POR2X1_7/B 0.03fF
C64390 PAND2X1_653/O POR2X1_760/A 0.01fF
C64391 POR2X1_502/A POR2X1_785/A 0.03fF
C64392 PAND2X1_695/a_76_28# PAND2X1_23/Y 0.02fF
C64393 POR2X1_46/Y POR2X1_531/O 0.05fF
C64394 POR2X1_244/B POR2X1_340/O 0.01fF
C64395 POR2X1_672/O POR2X1_5/Y 0.01fF
C64396 PAND2X1_217/B PAND2X1_572/O 0.09fF
C64397 POR2X1_652/CTRL POR2X1_480/A 0.04fF
C64398 POR2X1_62/Y PAND2X1_404/Y 0.03fF
C64399 POR2X1_847/A POR2X1_283/A 0.07fF
C64400 POR2X1_13/A PAND2X1_639/B 0.03fF
C64401 PAND2X1_360/O PAND2X1_843/Y 0.02fF
C64402 POR2X1_97/CTRL2 PAND2X1_20/A 0.00fF
C64403 POR2X1_646/CTRL POR2X1_294/B 0.00fF
C64404 POR2X1_215/CTRL2 POR2X1_35/Y 0.01fF
C64405 POR2X1_720/B VDD 0.14fF
C64406 PAND2X1_226/O POR2X1_578/Y 0.03fF
C64407 PAND2X1_362/B PAND2X1_357/Y 0.03fF
C64408 POR2X1_426/Y POR2X1_427/Y 0.00fF
C64409 POR2X1_597/Y POR2X1_761/A 0.33fF
C64410 POR2X1_519/O POR2X1_667/A 0.07fF
C64411 PAND2X1_23/Y POR2X1_776/B 0.03fF
C64412 POR2X1_49/Y PAND2X1_469/Y 0.02fF
C64413 POR2X1_402/CTRL2 PAND2X1_60/B 0.01fF
C64414 POR2X1_445/A POR2X1_703/m4_208_n4# 0.03fF
C64415 PAND2X1_269/CTRL2 POR2X1_55/Y 0.00fF
C64416 POR2X1_777/O POR2X1_784/A 0.11fF
C64417 POR2X1_465/B POR2X1_563/Y 0.10fF
C64418 PAND2X1_90/Y POR2X1_540/O 0.01fF
C64419 POR2X1_71/Y PAND2X1_575/A 0.03fF
C64420 PAND2X1_824/B POR2X1_590/A 0.05fF
C64421 POR2X1_265/Y PAND2X1_267/a_16_344# 0.02fF
C64422 POR2X1_193/A POR2X1_556/O 0.04fF
C64423 POR2X1_346/B PAND2X1_626/O 0.00fF
C64424 PAND2X1_81/O VDD 0.00fF
C64425 PAND2X1_541/O POR2X1_7/A 0.01fF
C64426 POR2X1_78/A POR2X1_502/a_76_344# 0.01fF
C64427 PAND2X1_525/CTRL POR2X1_550/Y 0.01fF
C64428 POR2X1_193/A POR2X1_795/a_16_28# 0.03fF
C64429 PAND2X1_793/Y POR2X1_184/Y 0.03fF
C64430 PAND2X1_424/O POR2X1_480/A 0.06fF
C64431 POR2X1_614/A POR2X1_812/CTRL 0.01fF
C64432 POR2X1_333/a_16_28# POR2X1_333/A 0.03fF
C64433 POR2X1_390/B POR2X1_330/Y 0.05fF
C64434 POR2X1_41/B POR2X1_152/O 0.03fF
C64435 POR2X1_288/A POR2X1_101/Y 0.05fF
C64436 PAND2X1_96/B POR2X1_435/Y 0.15fF
C64437 POR2X1_383/A PAND2X1_65/Y 0.03fF
C64438 PAND2X1_492/a_16_344# POR2X1_532/A 0.06fF
C64439 POR2X1_245/CTRL VDD 0.00fF
C64440 D_INPUT_0 POR2X1_512/CTRL2 0.03fF
C64441 PAND2X1_84/O POR2X1_91/Y 0.15fF
C64442 PAND2X1_651/Y PAND2X1_793/Y 0.05fF
C64443 POR2X1_812/B VDD 0.10fF
C64444 POR2X1_346/B POR2X1_750/B 0.05fF
C64445 POR2X1_52/A POR2X1_239/CTRL2 0.03fF
C64446 PAND2X1_803/Y PAND2X1_140/Y 0.01fF
C64447 INPUT_1 POR2X1_24/CTRL 0.01fF
C64448 PAND2X1_241/O POR2X1_237/Y 0.02fF
C64449 POR2X1_142/O POR2X1_394/A 0.06fF
C64450 POR2X1_60/A POR2X1_129/Y 0.10fF
C64451 PAND2X1_794/B POR2X1_42/Y 0.03fF
C64452 POR2X1_345/CTRL POR2X1_330/Y 0.03fF
C64453 POR2X1_347/B POR2X1_68/B 0.19fF
C64454 POR2X1_8/Y POR2X1_40/Y 0.43fF
C64455 POR2X1_45/Y PAND2X1_798/B 0.03fF
C64456 POR2X1_57/A PAND2X1_804/B 0.07fF
C64457 POR2X1_409/CTRL2 POR2X1_55/Y 0.00fF
C64458 POR2X1_38/Y PAND2X1_598/a_16_344# 0.01fF
C64459 POR2X1_599/A PAND2X1_717/O 0.02fF
C64460 POR2X1_832/A VDD 0.16fF
C64461 POR2X1_106/Y PAND2X1_114/CTRL 0.01fF
C64462 PAND2X1_90/Y POR2X1_707/Y 0.02fF
C64463 POR2X1_780/B VDD 0.43fF
C64464 POR2X1_614/A POR2X1_556/O 0.01fF
C64465 POR2X1_294/B POR2X1_702/A 0.04fF
C64466 POR2X1_863/A POR2X1_453/Y 0.01fF
C64467 POR2X1_751/CTRL POR2X1_7/B 0.01fF
C64468 GATE_811 VDD 0.00fF
C64469 POR2X1_613/Y POR2X1_32/A 0.02fF
C64470 POR2X1_96/Y PAND2X1_61/O 0.01fF
C64471 PAND2X1_243/B PAND2X1_243/a_16_344# 0.02fF
C64472 PAND2X1_82/Y VDD 0.07fF
C64473 PAND2X1_486/O POR2X1_526/Y 0.05fF
C64474 POR2X1_49/Y POR2X1_394/A 0.28fF
C64475 POR2X1_316/O PAND2X1_390/Y 0.01fF
C64476 POR2X1_812/A POR2X1_294/A 0.03fF
C64477 PAND2X1_857/A POR2X1_13/A 0.12fF
C64478 PAND2X1_651/Y PAND2X1_197/m4_208_n4# 0.06fF
C64479 POR2X1_192/Y POR2X1_854/B 0.12fF
C64480 PAND2X1_659/Y POR2X1_60/A 0.06fF
C64481 POR2X1_55/Y PAND2X1_509/O 0.29fF
C64482 PAND2X1_672/CTRL2 POR2X1_35/B 0.01fF
C64483 PAND2X1_212/B PAND2X1_352/O 0.02fF
C64484 PAND2X1_209/A PAND2X1_162/O 0.03fF
C64485 INPUT_0 PAND2X1_537/CTRL2 0.01fF
C64486 POR2X1_840/Y POR2X1_660/Y 0.01fF
C64487 POR2X1_394/A PAND2X1_558/CTRL2 0.11fF
C64488 POR2X1_858/B VDD 0.05fF
C64489 PAND2X1_65/B POR2X1_590/Y 0.03fF
C64490 POR2X1_693/CTRL2 PAND2X1_550/B 0.01fF
C64491 POR2X1_408/Y POR2X1_293/Y 0.10fF
C64492 POR2X1_316/a_16_28# PAND2X1_436/A 0.04fF
C64493 POR2X1_55/Y POR2X1_142/Y 0.03fF
C64494 POR2X1_72/B PAND2X1_657/B 0.00fF
C64495 POR2X1_22/A POR2X1_36/O 0.04fF
C64496 POR2X1_222/A POR2X1_554/Y 0.09fF
C64497 POR2X1_96/Y POR2X1_60/A 0.03fF
C64498 PAND2X1_48/CTRL POR2X1_260/A 0.01fF
C64499 POR2X1_840/CTRL2 POR2X1_513/Y 0.04fF
C64500 POR2X1_686/B POR2X1_260/A 0.66fF
C64501 POR2X1_12/O POR2X1_3/B 0.19fF
C64502 PAND2X1_96/O POR2X1_202/A 0.06fF
C64503 POR2X1_16/A PAND2X1_735/Y 0.10fF
C64504 POR2X1_336/CTRL2 PAND2X1_69/A 0.01fF
C64505 POR2X1_42/Y PAND2X1_842/Y 0.04fF
C64506 POR2X1_124/B POR2X1_123/Y 0.00fF
C64507 PAND2X1_808/a_16_344# PAND2X1_803/Y 0.02fF
C64508 D_GATE_222 PAND2X1_173/O 0.03fF
C64509 PAND2X1_6/Y POR2X1_140/O 0.01fF
C64510 POR2X1_43/B PAND2X1_338/B 0.07fF
C64511 PAND2X1_808/Y PAND2X1_854/A 0.02fF
C64512 PAND2X1_524/O POR2X1_456/B 0.09fF
C64513 POR2X1_257/Y PAND2X1_569/Y 0.03fF
C64514 POR2X1_646/a_16_28# POR2X1_646/A 0.03fF
C64515 POR2X1_41/B PAND2X1_726/B 0.02fF
C64516 POR2X1_236/Y PAND2X1_123/Y 0.18fF
C64517 PAND2X1_716/a_76_28# POR2X1_73/Y 0.01fF
C64518 PAND2X1_96/B POR2X1_736/CTRL2 0.01fF
C64519 PAND2X1_90/Y PAND2X1_384/a_76_28# 0.01fF
C64520 PAND2X1_6/Y POR2X1_197/Y 1.04fF
C64521 PAND2X1_411/O POR2X1_713/B 0.32fF
C64522 GATE_662 PAND2X1_660/B 0.05fF
C64523 PAND2X1_823/O POR2X1_857/B 0.05fF
C64524 POR2X1_297/A PAND2X1_359/Y 0.01fF
C64525 PAND2X1_61/Y PAND2X1_338/CTRL 0.01fF
C64526 PAND2X1_111/O POR2X1_366/A 0.06fF
C64527 POR2X1_303/O POR2X1_814/B 0.01fF
C64528 POR2X1_256/Y PAND2X1_344/O 0.00fF
C64529 POR2X1_786/Y POR2X1_702/O 0.26fF
C64530 PAND2X1_111/B POR2X1_702/A 0.04fF
C64531 D_INPUT_3 PAND2X1_509/CTRL2 0.04fF
C64532 PAND2X1_410/O POR2X1_234/A 0.02fF
C64533 INPUT_1 PAND2X1_341/CTRL 0.00fF
C64534 POR2X1_730/Y PAND2X1_55/Y 0.00fF
C64535 POR2X1_502/A POR2X1_186/B 0.03fF
C64536 PAND2X1_6/Y POR2X1_802/O 0.01fF
C64537 D_INPUT_3 POR2X1_38/Y 0.10fF
C64538 POR2X1_502/m4_208_n4# POR2X1_854/B 0.06fF
C64539 PAND2X1_56/Y PAND2X1_368/a_16_344# 0.04fF
C64540 PAND2X1_553/B POR2X1_394/A 0.03fF
C64541 POR2X1_93/O POR2X1_283/A 0.01fF
C64542 POR2X1_49/Y PAND2X1_198/CTRL2 0.03fF
C64543 POR2X1_356/A POR2X1_724/B 0.33fF
C64544 PAND2X1_777/CTRL POR2X1_55/Y 0.09fF
C64545 PAND2X1_94/A PAND2X1_283/O 0.22fF
C64546 PAND2X1_714/B VDD 0.23fF
C64547 POR2X1_417/O POR2X1_7/A 0.05fF
C64548 PAND2X1_824/B POR2X1_214/B 0.06fF
C64549 POR2X1_343/Y PAND2X1_74/O 0.24fF
C64550 POR2X1_60/A PAND2X1_333/Y 0.98fF
C64551 POR2X1_862/CTRL2 POR2X1_389/Y 0.03fF
C64552 POR2X1_366/A POR2X1_573/A 0.03fF
C64553 PAND2X1_242/Y POR2X1_37/Y 0.05fF
C64554 POR2X1_394/A PAND2X1_188/O 0.15fF
C64555 POR2X1_46/Y PAND2X1_325/O 0.02fF
C64556 PAND2X1_6/Y INPUT_1 0.03fF
C64557 POR2X1_93/A POR2X1_384/O 0.01fF
C64558 POR2X1_416/B PAND2X1_260/O 0.00fF
C64559 POR2X1_328/CTRL INPUT_4 0.01fF
C64560 POR2X1_328/CTRL2 INPUT_5 0.00fF
C64561 PAND2X1_150/a_76_28# PAND2X1_63/B 0.01fF
C64562 PAND2X1_118/O POR2X1_559/A 0.18fF
C64563 POR2X1_504/Y POR2X1_416/B 2.25fF
C64564 PAND2X1_23/Y PAND2X1_48/A 0.07fF
C64565 PAND2X1_48/B POR2X1_294/A 0.13fF
C64566 PAND2X1_495/CTRL POR2X1_260/A 0.01fF
C64567 POR2X1_416/B PAND2X1_740/CTRL 0.10fF
C64568 PAND2X1_850/Y PAND2X1_592/CTRL2 0.01fF
C64569 PAND2X1_649/A POR2X1_393/a_16_28# 0.02fF
C64570 POR2X1_278/Y POR2X1_680/CTRL 0.06fF
C64571 PAND2X1_631/A PAND2X1_515/O 0.10fF
C64572 PAND2X1_23/Y POR2X1_192/B 0.09fF
C64573 POR2X1_549/CTRL2 PAND2X1_52/B 0.31fF
C64574 POR2X1_327/Y POR2X1_276/a_16_28# 0.02fF
C64575 PAND2X1_630/O PAND2X1_156/A 0.05fF
C64576 PAND2X1_798/Y GATE_741 0.03fF
C64577 POR2X1_568/Y POR2X1_854/B 0.03fF
C64578 D_INPUT_3 INPUT_1 0.26fF
C64579 PAND2X1_625/CTRL POR2X1_294/A 0.01fF
C64580 PAND2X1_843/m4_208_n4# POR2X1_416/B 0.12fF
C64581 PAND2X1_658/A POR2X1_171/Y 0.02fF
C64582 POR2X1_83/A POR2X1_397/CTRL2 0.01fF
C64583 POR2X1_726/Y POR2X1_738/A 0.01fF
C64584 POR2X1_265/Y PAND2X1_734/CTRL2 0.01fF
C64585 POR2X1_622/CTRL2 POR2X1_29/A 0.03fF
C64586 POR2X1_763/Y POR2X1_524/O 0.00fF
C64587 POR2X1_353/A POR2X1_319/Y 0.03fF
C64588 POR2X1_344/Y POR2X1_205/A 0.02fF
C64589 POR2X1_48/A POR2X1_67/Y 0.03fF
C64590 POR2X1_507/A PAND2X1_60/B 0.07fF
C64591 D_INPUT_3 POR2X1_153/Y 0.03fF
C64592 D_INPUT_3 POR2X1_384/A 0.00fF
C64593 POR2X1_540/A POR2X1_552/CTRL 0.02fF
C64594 POR2X1_778/O POR2X1_717/B 0.01fF
C64595 PAND2X1_531/CTRL PAND2X1_111/B 0.02fF
C64596 PAND2X1_824/B PAND2X1_824/a_16_344# 0.01fF
C64597 POR2X1_613/Y PAND2X1_651/Y 0.00fF
C64598 PAND2X1_94/A POR2X1_463/Y 0.07fF
C64599 PAND2X1_787/A PAND2X1_357/O 0.02fF
C64600 INPUT_2 POR2X1_4/Y 0.04fF
C64601 POR2X1_814/A POR2X1_296/B 0.09fF
C64602 PAND2X1_323/O POR2X1_702/A 0.00fF
C64603 POR2X1_210/A POR2X1_162/Y 0.01fF
C64604 POR2X1_246/CTRL2 POR2X1_39/B 0.03fF
C64605 POR2X1_83/Y POR2X1_38/Y 0.02fF
C64606 PAND2X1_109/CTRL POR2X1_775/A 0.01fF
C64607 POR2X1_316/Y PAND2X1_457/CTRL2 0.01fF
C64608 POR2X1_841/O POR2X1_841/B 0.07fF
C64609 POR2X1_327/CTRL PAND2X1_72/A 0.01fF
C64610 POR2X1_455/A POR2X1_632/Y 0.03fF
C64611 POR2X1_132/a_56_344# PAND2X1_140/A 0.00fF
C64612 PAND2X1_440/CTRL PAND2X1_798/B 0.03fF
C64613 PAND2X1_865/Y POR2X1_91/Y 0.03fF
C64614 POR2X1_20/B POR2X1_626/O 0.01fF
C64615 POR2X1_86/Y PAND2X1_101/O 0.03fF
C64616 POR2X1_55/a_76_344# POR2X1_624/B 0.03fF
C64617 POR2X1_799/O POR2X1_652/A 0.00fF
C64618 POR2X1_447/A POR2X1_454/A 0.03fF
C64619 PAND2X1_661/Y POR2X1_119/Y 0.05fF
C64620 POR2X1_866/A POR2X1_655/A 0.06fF
C64621 POR2X1_707/CTRL PAND2X1_48/A 0.01fF
C64622 PAND2X1_789/O POR2X1_751/Y 0.00fF
C64623 POR2X1_416/B POR2X1_136/O 0.01fF
C64624 POR2X1_390/B POR2X1_337/Y 0.00fF
C64625 PAND2X1_301/O POR2X1_75/Y 0.02fF
C64626 PAND2X1_301/CTRL2 PAND2X1_716/B 0.01fF
C64627 POR2X1_23/Y POR2X1_265/CTRL2 0.01fF
C64628 POR2X1_218/A PAND2X1_72/A 0.01fF
C64629 POR2X1_57/A POR2X1_43/O 0.01fF
C64630 POR2X1_750/CTRL POR2X1_39/B 0.03fF
C64631 PAND2X1_242/Y POR2X1_293/Y 0.07fF
C64632 POR2X1_257/A POR2X1_669/B 0.38fF
C64633 PAND2X1_737/B PAND2X1_737/CTRL 0.02fF
C64634 POR2X1_435/CTRL PAND2X1_72/A 0.01fF
C64635 POR2X1_611/a_16_28# POR2X1_293/Y 0.03fF
C64636 POR2X1_228/Y POR2X1_716/CTRL2 0.01fF
C64637 PAND2X1_663/a_56_28# PAND2X1_659/Y 0.00fF
C64638 D_GATE_662 POR2X1_863/A 0.07fF
C64639 PAND2X1_605/m4_208_n4# POR2X1_604/m4_208_n4# 0.05fF
C64640 POR2X1_820/O POR2X1_411/B 0.02fF
C64641 POR2X1_537/B POR2X1_711/Y 0.03fF
C64642 POR2X1_11/CTRL2 INPUT_7 0.03fF
C64643 PAND2X1_474/Y POR2X1_329/A 0.03fF
C64644 PAND2X1_439/CTRL2 PAND2X1_738/Y 0.14fF
C64645 PAND2X1_221/Y POR2X1_42/Y 0.03fF
C64646 PAND2X1_217/B POR2X1_411/B 0.12fF
C64647 POR2X1_188/Y POR2X1_186/B 0.03fF
C64648 POR2X1_666/Y POR2X1_411/B 0.04fF
C64649 PAND2X1_856/O PAND2X1_854/Y 0.02fF
C64650 POR2X1_54/Y POR2X1_69/A 0.06fF
C64651 PAND2X1_798/Y PAND2X1_356/a_56_28# 0.00fF
C64652 POR2X1_514/a_16_28# POR2X1_138/A 0.09fF
C64653 POR2X1_106/CTRL2 POR2X1_48/A 0.01fF
C64654 POR2X1_67/a_16_28# POR2X1_67/A 0.02fF
C64655 POR2X1_777/B POR2X1_475/O 0.04fF
C64656 POR2X1_371/a_16_28# POR2X1_153/Y 0.08fF
C64657 POR2X1_13/A POR2X1_329/A 0.07fF
C64658 POR2X1_567/A POR2X1_566/O 0.03fF
C64659 PAND2X1_68/O D_INPUT_0 0.08fF
C64660 POR2X1_411/B PAND2X1_392/B 0.03fF
C64661 PAND2X1_467/Y POR2X1_416/B 0.03fF
C64662 POR2X1_16/A PAND2X1_440/CTRL2 0.02fF
C64663 PAND2X1_631/A PAND2X1_156/A 0.03fF
C64664 POR2X1_343/Y POR2X1_276/Y 0.05fF
C64665 POR2X1_685/A PAND2X1_681/CTRL 0.00fF
C64666 POR2X1_144/O PAND2X1_797/Y 0.01fF
C64667 PAND2X1_849/B POR2X1_86/Y 0.00fF
C64668 POR2X1_89/a_16_28# POR2X1_60/A 0.01fF
C64669 POR2X1_14/Y POR2X1_409/B 0.03fF
C64670 POR2X1_150/Y PAND2X1_579/B 0.03fF
C64671 POR2X1_60/A POR2X1_37/Y 0.18fF
C64672 POR2X1_257/A PAND2X1_210/CTRL 0.01fF
C64673 POR2X1_11/CTRL2 INPUT_4 0.02fF
C64674 POR2X1_9/Y POR2X1_816/A 0.10fF
C64675 POR2X1_411/B VDD 2.53fF
C64676 POR2X1_91/O POR2X1_91/Y 0.02fF
C64677 INPUT_1 PAND2X1_52/B 0.08fF
C64678 PAND2X1_827/CTRL2 POR2X1_355/A 0.01fF
C64679 POR2X1_590/A POR2X1_720/O 0.01fF
C64680 PAND2X1_434/O PAND2X1_390/Y 0.02fF
C64681 POR2X1_32/A POR2X1_516/Y 0.06fF
C64682 PAND2X1_58/A POR2X1_608/Y 0.01fF
C64683 POR2X1_567/A POR2X1_741/CTRL 0.01fF
C64684 POR2X1_585/Y PAND2X1_638/B 0.01fF
C64685 PAND2X1_678/O PAND2X1_804/B 0.02fF
C64686 POR2X1_260/B PAND2X1_597/O 0.02fF
C64687 POR2X1_43/B PAND2X1_717/A 0.06fF
C64688 PAND2X1_777/O PAND2X1_784/A 0.02fF
C64689 POR2X1_142/O POR2X1_669/B 0.03fF
C64690 POR2X1_78/B PAND2X1_601/CTRL2 0.02fF
C64691 PAND2X1_75/O POR2X1_741/Y 0.08fF
C64692 PAND2X1_486/O POR2X1_485/Y 0.00fF
C64693 POR2X1_506/B POR2X1_590/A 0.06fF
C64694 PAND2X1_301/O PAND2X1_332/Y 0.03fF
C64695 POR2X1_23/Y PAND2X1_220/Y 0.05fF
C64696 PAND2X1_420/O POR2X1_590/A 0.17fF
C64697 POR2X1_597/Y POR2X1_829/A 0.03fF
C64698 PAND2X1_48/A POR2X1_711/Y 0.07fF
C64699 POR2X1_150/Y PAND2X1_592/m4_208_n4# 0.08fF
C64700 PAND2X1_586/CTRL2 PAND2X1_72/A 0.01fF
C64701 POR2X1_347/A PAND2X1_96/O 0.02fF
C64702 PAND2X1_622/O POR2X1_48/A 0.01fF
C64703 PAND2X1_48/B POR2X1_116/A 0.03fF
C64704 PAND2X1_65/B PAND2X1_237/O 0.15fF
C64705 PAND2X1_859/CTRL POR2X1_37/Y 0.04fF
C64706 POR2X1_603/a_16_28# POR2X1_597/A 0.04fF
C64707 POR2X1_368/Y PAND2X1_464/B 0.02fF
C64708 POR2X1_347/B POR2X1_68/Y 0.08fF
C64709 POR2X1_557/B PAND2X1_72/A 0.07fF
C64710 PAND2X1_420/CTRL2 POR2X1_630/A 0.02fF
C64711 POR2X1_49/Y POR2X1_669/B 1.73fF
C64712 POR2X1_554/B POR2X1_140/B 0.00fF
C64713 PAND2X1_23/Y POR2X1_461/Y 0.05fF
C64714 PAND2X1_633/CTRL POR2X1_32/A 0.01fF
C64715 POR2X1_852/B POR2X1_296/B 0.09fF
C64716 POR2X1_84/A INPUT_0 0.03fF
C64717 POR2X1_41/B PAND2X1_35/A 0.00fF
C64718 PAND2X1_294/O POR2X1_293/Y 0.00fF
C64719 PAND2X1_443/Y PAND2X1_211/A 0.72fF
C64720 POR2X1_312/CTRL POR2X1_20/B 0.01fF
C64721 POR2X1_660/O POR2X1_660/A 0.14fF
C64722 PAND2X1_738/Y POR2X1_438/Y 0.10fF
C64723 POR2X1_726/a_16_28# POR2X1_711/Y 0.07fF
C64724 POR2X1_428/Y POR2X1_700/CTRL 0.01fF
C64725 PAND2X1_57/B PAND2X1_59/B 0.18fF
C64726 PAND2X1_807/B PAND2X1_363/Y 0.02fF
C64727 PAND2X1_52/B PAND2X1_680/CTRL 0.04fF
C64728 PAND2X1_217/B POR2X1_271/Y 0.05fF
C64729 PAND2X1_200/a_16_344# POR2X1_72/B 0.05fF
C64730 POR2X1_568/B POR2X1_568/CTRL 0.05fF
C64731 D_GATE_811 POR2X1_452/Y 0.07fF
C64732 PAND2X1_221/O PAND2X1_220/Y 0.09fF
C64733 PAND2X1_221/CTRL PAND2X1_192/Y 0.01fF
C64734 POR2X1_801/A POR2X1_121/B 0.15fF
C64735 POR2X1_514/Y POR2X1_446/B 0.04fF
C64736 PAND2X1_609/O POR2X1_294/B 0.01fF
C64737 PAND2X1_838/CTRL2 POR2X1_73/Y 0.03fF
C64738 POR2X1_840/B POR2X1_541/B 0.04fF
C64739 PAND2X1_81/O PAND2X1_9/Y 0.15fF
C64740 POR2X1_487/O PAND2X1_738/Y 0.02fF
C64741 PAND2X1_65/B POR2X1_633/A 0.02fF
C64742 PAND2X1_640/B POR2X1_290/Y 0.08fF
C64743 POR2X1_820/O POR2X1_376/B 0.07fF
C64744 PAND2X1_277/a_76_28# PAND2X1_57/B 0.05fF
C64745 POR2X1_864/A POR2X1_686/O 0.00fF
C64746 POR2X1_689/A PAND2X1_590/O 0.02fF
C64747 POR2X1_706/a_16_28# POR2X1_706/A 0.03fF
C64748 POR2X1_498/Y INPUT_0 0.15fF
C64749 POR2X1_423/O INPUT_0 0.02fF
C64750 PAND2X1_73/Y POR2X1_192/Y 0.03fF
C64751 POR2X1_760/A POR2X1_385/CTRL2 0.00fF
C64752 POR2X1_809/B POR2X1_121/B 0.03fF
C64753 POR2X1_68/A POR2X1_260/B 0.10fF
C64754 POR2X1_13/O POR2X1_102/Y 0.05fF
C64755 POR2X1_406/Y POR2X1_60/A 0.68fF
C64756 POR2X1_42/a_16_28# INPUT_3 0.13fF
C64757 POR2X1_278/Y POR2X1_487/m4_208_n4# 0.07fF
C64758 POR2X1_590/A POR2X1_121/Y 0.01fF
C64759 POR2X1_409/B POR2X1_55/Y 1.47fF
C64760 POR2X1_642/CTRL POR2X1_66/A 0.01fF
C64761 PAND2X1_65/B POR2X1_186/Y 0.06fF
C64762 POR2X1_41/B PAND2X1_804/a_76_28# 0.01fF
C64763 PAND2X1_221/CTRL PAND2X1_738/Y 0.31fF
C64764 POR2X1_362/B PAND2X1_41/B 0.07fF
C64765 PAND2X1_448/m4_208_n4# POR2X1_421/m4_208_n4# 0.05fF
C64766 POR2X1_343/O POR2X1_343/B 0.02fF
C64767 POR2X1_702/B PAND2X1_48/Y 1.39fF
C64768 POR2X1_3/A POR2X1_582/Y 0.00fF
C64769 PAND2X1_795/B PAND2X1_575/B 0.03fF
C64770 POR2X1_480/A POR2X1_389/Y 4.34fF
C64771 PAND2X1_814/a_76_28# INPUT_3 0.05fF
C64772 POR2X1_673/O PAND2X1_8/Y 0.03fF
C64773 POR2X1_78/A PAND2X1_322/a_16_344# 0.00fF
C64774 PAND2X1_668/O POR2X1_83/B 0.17fF
C64775 POR2X1_459/CTRL2 POR2X1_750/B 0.01fF
C64776 POR2X1_523/Y POR2X1_66/A 0.03fF
C64777 POR2X1_856/B POR2X1_340/a_16_28# 0.09fF
C64778 PAND2X1_58/A POR2X1_791/CTRL2 0.00fF
C64779 PAND2X1_139/B POR2X1_423/Y 0.01fF
C64780 POR2X1_460/A POR2X1_260/B 0.00fF
C64781 POR2X1_96/A PAND2X1_557/A 0.07fF
C64782 PAND2X1_787/CTRL2 VDD 0.00fF
C64783 POR2X1_411/Y POR2X1_102/Y 0.01fF
C64784 POR2X1_175/A POR2X1_175/a_16_28# 0.01fF
C64785 POR2X1_60/A POR2X1_293/Y 0.28fF
C64786 POR2X1_226/CTRL2 POR2X1_42/Y 0.03fF
C64787 PAND2X1_573/B POR2X1_494/Y 0.02fF
C64788 POR2X1_836/A POR2X1_579/Y 0.01fF
C64789 PAND2X1_84/CTRL2 POR2X1_5/Y 0.00fF
C64790 PAND2X1_699/a_76_28# POR2X1_260/A 0.02fF
C64791 POR2X1_653/O POR2X1_653/B 0.01fF
C64792 PAND2X1_159/O POR2X1_7/B 0.03fF
C64793 POR2X1_83/B POR2X1_42/Y 0.22fF
C64794 PAND2X1_217/B PAND2X1_598/O 0.04fF
C64795 POR2X1_417/Y PAND2X1_515/a_16_344# 0.02fF
C64796 PAND2X1_614/O POR2X1_625/Y 0.07fF
C64797 POR2X1_66/A PAND2X1_69/A 1.64fF
C64798 POR2X1_23/Y PAND2X1_575/CTRL 0.01fF
C64799 POR2X1_376/B VDD 4.37fF
C64800 POR2X1_805/B VDD 0.02fF
C64801 POR2X1_590/A POR2X1_723/B 0.07fF
C64802 PAND2X1_675/A POR2X1_102/Y 0.03fF
C64803 POR2X1_52/A PAND2X1_217/B 0.05fF
C64804 POR2X1_76/CTRL POR2X1_553/A 0.02fF
C64805 POR2X1_493/CTRL POR2X1_493/A 0.01fF
C64806 POR2X1_493/CTRL2 POR2X1_558/B 0.00fF
C64807 PAND2X1_793/Y PAND2X1_579/CTRL 0.01fF
C64808 PAND2X1_96/B PAND2X1_595/CTRL 0.01fF
C64809 PAND2X1_859/O POR2X1_13/A 0.05fF
C64810 PAND2X1_467/Y PAND2X1_452/CTRL2 0.01fF
C64811 PAND2X1_469/B POR2X1_102/Y 0.03fF
C64812 POR2X1_430/A VDD 0.00fF
C64813 POR2X1_17/CTRL INPUT_5 0.01fF
C64814 POR2X1_516/Y POR2X1_184/Y 0.03fF
C64815 POR2X1_174/B POR2X1_350/Y 0.01fF
C64816 POR2X1_88/Y POR2X1_5/Y 0.03fF
C64817 POR2X1_83/B POR2X1_309/Y 0.03fF
C64818 PAND2X1_689/O PAND2X1_32/B 0.05fF
C64819 POR2X1_49/Y PAND2X1_844/Y 0.01fF
C64820 PAND2X1_90/A PAND2X1_46/O 0.01fF
C64821 POR2X1_798/O POR2X1_468/B 0.04fF
C64822 PAND2X1_54/CTRL INPUT_0 0.01fF
C64823 PAND2X1_65/B POR2X1_483/O 0.17fF
C64824 POR2X1_7/B POR2X1_250/A 0.03fF
C64825 PAND2X1_78/CTRL PAND2X1_794/B 0.01fF
C64826 PAND2X1_803/A POR2X1_46/Y 0.03fF
C64827 PAND2X1_16/CTRL2 POR2X1_294/B 0.01fF
C64828 PAND2X1_341/B POR2X1_65/CTRL2 0.01fF
C64829 POR2X1_383/A POR2X1_647/a_76_344# 0.01fF
C64830 POR2X1_41/B PAND2X1_499/O 0.08fF
C64831 POR2X1_366/CTRL2 PAND2X1_93/B 0.01fF
C64832 POR2X1_57/A POR2X1_279/CTRL2 0.02fF
C64833 POR2X1_752/Y POR2X1_42/Y 0.07fF
C64834 POR2X1_196/O POR2X1_196/Y 0.01fF
C64835 PAND2X1_242/a_76_28# POR2X1_60/A 0.02fF
C64836 PAND2X1_25/CTRL INPUT_6 0.01fF
C64837 POR2X1_247/Y POR2X1_532/A 0.01fF
C64838 PAND2X1_37/O POR2X1_38/B 0.05fF
C64839 POR2X1_862/B PAND2X1_536/CTRL2 0.00fF
C64840 PAND2X1_93/B POR2X1_796/A 0.07fF
C64841 POR2X1_23/Y PAND2X1_713/A 0.04fF
C64842 PAND2X1_225/CTRL2 D_INPUT_1 0.00fF
C64843 POR2X1_685/A POR2X1_678/Y 0.00fF
C64844 D_INPUT_7 D_INPUT_4 0.12fF
C64845 POR2X1_232/O POR2X1_5/Y 0.09fF
C64846 D_INPUT_0 POR2X1_575/O 0.01fF
C64847 POR2X1_690/a_16_28# INPUT_0 0.00fF
C64848 POR2X1_662/O POR2X1_353/A 0.01fF
C64849 POR2X1_856/B POR2X1_738/A 0.03fF
C64850 POR2X1_260/B POR2X1_391/B 0.04fF
C64851 PAND2X1_425/Y PAND2X1_2/O 0.05fF
C64852 POR2X1_322/O POR2X1_376/B 0.18fF
C64853 POR2X1_29/CTRL2 POR2X1_55/Y 0.00fF
C64854 POR2X1_66/B POR2X1_840/B 0.05fF
C64855 POR2X1_227/A POR2X1_191/Y 0.05fF
C64856 POR2X1_814/B POR2X1_790/B 0.04fF
C64857 POR2X1_390/B POR2X1_558/B 0.00fF
C64858 POR2X1_52/A VDD 4.53fF
C64859 POR2X1_141/Y POR2X1_804/A 0.03fF
C64860 PAND2X1_724/B POR2X1_236/Y 0.03fF
C64861 POR2X1_678/Y POR2X1_260/A 0.03fF
C64862 POR2X1_502/A POR2X1_853/CTRL 0.15fF
C64863 POR2X1_188/A POR2X1_840/B 0.05fF
C64864 POR2X1_669/B PAND2X1_720/O 0.10fF
C64865 PAND2X1_269/a_16_344# POR2X1_39/B 0.02fF
C64866 POR2X1_634/A PAND2X1_757/CTRL 0.13fF
C64867 PAND2X1_478/B POR2X1_91/Y 0.03fF
C64868 POR2X1_669/B PAND2X1_559/CTRL 0.01fF
C64869 PAND2X1_317/Y VDD 0.05fF
C64870 POR2X1_35/B POR2X1_68/B 0.24fF
C64871 POR2X1_152/A VDD 0.27fF
C64872 POR2X1_13/Y PAND2X1_730/B 0.06fF
C64873 POR2X1_78/A POR2X1_796/A 0.03fF
C64874 POR2X1_750/B POR2X1_194/a_76_344# 0.04fF
C64875 PAND2X1_41/B POR2X1_194/O 0.01fF
C64876 POR2X1_38/Y PAND2X1_733/O 0.16fF
C64877 POR2X1_62/Y POR2X1_88/CTRL 0.01fF
C64878 POR2X1_23/Y PAND2X1_560/B 0.03fF
C64879 POR2X1_251/A POR2X1_387/Y 0.25fF
C64880 PAND2X1_824/B POR2X1_66/A 2.63fF
C64881 POR2X1_316/Y PAND2X1_464/CTRL2 0.01fF
C64882 PAND2X1_42/CTRL2 PAND2X1_111/B 0.01fF
C64883 POR2X1_407/Y PAND2X1_597/O 0.02fF
C64884 PAND2X1_768/Y PAND2X1_359/a_16_344# 0.03fF
C64885 POR2X1_72/B POR2X1_387/Y 0.08fF
C64886 POR2X1_408/CTRL INPUT_5 0.01fF
C64887 POR2X1_29/A POR2X1_260/A 0.10fF
C64888 POR2X1_57/A PAND2X1_562/B 0.07fF
C64889 POR2X1_730/Y POR2X1_174/A 0.02fF
C64890 PAND2X1_856/B POR2X1_102/Y 0.03fF
C64891 PAND2X1_855/CTRL POR2X1_236/Y 0.02fF
C64892 POR2X1_502/A POR2X1_459/A 0.04fF
C64893 PAND2X1_550/Y POR2X1_40/Y 0.02fF
C64894 POR2X1_96/a_16_28# POR2X1_37/Y 0.05fF
C64895 POR2X1_356/A POR2X1_740/Y 0.05fF
C64896 POR2X1_355/B D_GATE_741 0.02fF
C64897 PAND2X1_181/O POR2X1_40/Y 0.17fF
C64898 PAND2X1_48/B PAND2X1_280/a_56_28# 0.00fF
C64899 PAND2X1_445/Y POR2X1_237/Y 0.01fF
C64900 PAND2X1_7/Y POR2X1_222/A 0.06fF
C64901 POR2X1_850/B POR2X1_675/Y 1.24fF
C64902 POR2X1_41/B POR2X1_43/B 0.63fF
C64903 PAND2X1_429/m4_208_n4# POR2X1_260/A 0.01fF
C64904 POR2X1_278/Y POR2X1_816/A 0.07fF
C64905 POR2X1_826/Y POR2X1_39/B 0.00fF
C64906 POR2X1_237/a_76_344# POR2X1_90/Y -0.00fF
C64907 POR2X1_333/A POR2X1_353/A 0.05fF
C64908 POR2X1_32/A PAND2X1_708/CTRL 0.01fF
C64909 POR2X1_210/Y VDD 0.23fF
C64910 POR2X1_409/B PAND2X1_199/B 0.01fF
C64911 PAND2X1_492/CTRL2 PAND2X1_60/B 0.01fF
C64912 POR2X1_410/Y POR2X1_410/O 0.00fF
C64913 POR2X1_364/A POR2X1_170/B 0.03fF
C64914 PAND2X1_543/CTRL POR2X1_142/Y 0.00fF
C64915 POR2X1_845/CTRL POR2X1_5/Y 0.04fF
C64916 POR2X1_502/A POR2X1_542/B 1.84fF
C64917 POR2X1_128/CTRL PAND2X1_96/B 0.01fF
C64918 POR2X1_773/O POR2X1_734/A 0.03fF
C64919 POR2X1_52/A POR2X1_93/CTRL 0.01fF
C64920 POR2X1_860/A POR2X1_116/Y 0.12fF
C64921 POR2X1_68/A PAND2X1_55/Y 0.28fF
C64922 POR2X1_43/B PAND2X1_228/O 0.20fF
C64923 PAND2X1_216/B PAND2X1_558/Y 0.09fF
C64924 POR2X1_66/B PAND2X1_748/a_76_28# 0.01fF
C64925 PAND2X1_808/Y PAND2X1_675/A 0.05fF
C64926 POR2X1_57/A POR2X1_13/A 0.26fF
C64927 PAND2X1_254/O PAND2X1_6/A -0.01fF
C64928 POR2X1_287/B POR2X1_249/Y 0.02fF
C64929 INPUT_4 POR2X1_3/O 0.05fF
C64930 POR2X1_730/Y POR2X1_686/A 0.01fF
C64931 POR2X1_73/Y PAND2X1_364/B 0.07fF
C64932 PAND2X1_661/Y PAND2X1_688/CTRL 0.09fF
C64933 POR2X1_856/B PAND2X1_167/O 0.02fF
C64934 VDD POR2X1_550/Y 0.00fF
C64935 POR2X1_407/A POR2X1_800/A 0.03fF
C64936 PAND2X1_803/A PAND2X1_727/CTRL2 0.00fF
C64937 POR2X1_93/O POR2X1_55/Y 0.02fF
C64938 POR2X1_853/A POR2X1_614/A 0.03fF
C64939 POR2X1_301/O POR2X1_335/A 0.01fF
C64940 PAND2X1_428/CTRL2 PAND2X1_48/A 0.17fF
C64941 POR2X1_60/Y POR2X1_153/Y 0.05fF
C64942 PAND2X1_477/B POR2X1_238/Y 0.02fF
C64943 POR2X1_70/m4_208_n4# POR2X1_90/Y 0.15fF
C64944 PAND2X1_857/A POR2X1_821/O 0.02fF
C64945 POR2X1_68/A POR2X1_402/A 0.07fF
C64946 INPUT_1 POR2X1_625/O 0.01fF
C64947 POR2X1_278/Y PAND2X1_854/A 0.02fF
C64948 POR2X1_222/Y PAND2X1_69/A 0.03fF
C64949 POR2X1_679/B VDD 0.10fF
C64950 POR2X1_596/A POR2X1_294/B 0.03fF
C64951 POR2X1_396/Y POR2X1_669/O 0.02fF
C64952 PAND2X1_63/Y POR2X1_204/CTRL2 0.01fF
C64953 POR2X1_503/CTRL POR2X1_236/Y 0.15fF
C64954 POR2X1_8/Y POR2X1_5/Y 0.10fF
C64955 POR2X1_494/Y POR2X1_91/Y 0.03fF
C64956 PAND2X1_229/CTRL POR2X1_186/B 0.01fF
C64957 POR2X1_389/A PAND2X1_48/B 0.01fF
C64958 PAND2X1_6/Y POR2X1_796/O 0.18fF
C64959 PAND2X1_390/Y PAND2X1_508/Y 0.03fF
C64960 POR2X1_122/a_56_344# POR2X1_40/Y 0.01fF
C64961 POR2X1_390/B POR2X1_723/CTRL2 0.00fF
C64962 PAND2X1_20/A POR2X1_540/Y 0.05fF
C64963 PAND2X1_90/A POR2X1_318/A 0.07fF
C64964 POR2X1_76/Y POR2X1_569/A 0.02fF
C64965 POR2X1_391/a_16_28# POR2X1_546/A 0.07fF
C64966 POR2X1_96/A PAND2X1_723/A 0.06fF
C64967 POR2X1_265/Y POR2X1_40/Y 0.04fF
C64968 POR2X1_777/Y POR2X1_784/A 0.01fF
C64969 PAND2X1_96/B PAND2X1_767/CTRL2 0.01fF
C64970 PAND2X1_144/CTRL2 PAND2X1_60/B 0.00fF
C64971 POR2X1_147/A POR2X1_532/A 0.02fF
C64972 POR2X1_122/A POR2X1_394/A 0.02fF
C64973 POR2X1_141/CTRL POR2X1_574/Y 0.01fF
C64974 POR2X1_785/A POR2X1_510/Y 0.10fF
C64975 POR2X1_523/Y POR2X1_532/A 0.03fF
C64976 POR2X1_65/A PAND2X1_800/a_16_344# 0.02fF
C64977 PAND2X1_392/O POR2X1_39/B 0.04fF
C64978 POR2X1_299/CTRL2 POR2X1_90/Y 0.01fF
C64979 POR2X1_326/A POR2X1_798/O 0.18fF
C64980 POR2X1_96/CTRL2 PAND2X1_472/B 0.03fF
C64981 POR2X1_502/A PAND2X1_376/CTRL 0.01fF
C64982 INPUT_2 D_INPUT_1 2.21fF
C64983 POR2X1_546/A POR2X1_260/A 0.06fF
C64984 POR2X1_865/B POR2X1_114/CTRL 0.00fF
C64985 POR2X1_489/O POR2X1_294/A 0.05fF
C64986 POR2X1_782/B VDD 0.13fF
C64987 POR2X1_532/A POR2X1_219/CTRL2 0.01fF
C64988 POR2X1_25/CTRL2 PAND2X1_18/B 0.03fF
C64989 PAND2X1_63/Y POR2X1_500/Y 0.21fF
C64990 POR2X1_260/B POR2X1_138/A 0.03fF
C64991 POR2X1_13/A PAND2X1_301/O 0.04fF
C64992 POR2X1_356/A PAND2X1_824/a_76_28# 0.02fF
C64993 PAND2X1_803/Y PAND2X1_357/Y 0.02fF
C64994 POR2X1_464/O POR2X1_186/B 0.01fF
C64995 POR2X1_740/Y POR2X1_569/A 0.10fF
C64996 POR2X1_532/A PAND2X1_69/A 0.21fF
C64997 PAND2X1_557/CTRL VDD 0.00fF
C64998 POR2X1_514/Y POR2X1_383/A 0.03fF
C64999 POR2X1_174/B PAND2X1_109/O 0.13fF
C65000 PAND2X1_632/a_76_28# INPUT_0 0.04fF
C65001 POR2X1_180/B PAND2X1_55/Y 0.00fF
C65002 POR2X1_81/a_16_28# POR2X1_81/A 0.03fF
C65003 POR2X1_326/O POR2X1_468/B 0.02fF
C65004 PAND2X1_341/Y PAND2X1_350/A 0.00fF
C65005 POR2X1_564/B POR2X1_552/Y 0.00fF
C65006 POR2X1_57/A PAND2X1_643/Y 0.03fF
C65007 POR2X1_814/B POR2X1_540/Y 0.05fF
C65008 POR2X1_786/Y PAND2X1_60/B 0.12fF
C65009 POR2X1_751/a_56_344# POR2X1_816/A 0.00fF
C65010 PAND2X1_486/O PAND2X1_726/B 0.10fF
C65011 POR2X1_567/A POR2X1_653/B 0.03fF
C65012 POR2X1_452/A POR2X1_452/a_16_28# 0.11fF
C65013 POR2X1_637/CTRL PAND2X1_72/A 0.01fF
C65014 POR2X1_65/A PAND2X1_476/A 0.03fF
C65015 PAND2X1_483/CTRL POR2X1_55/Y 0.01fF
C65016 POR2X1_3/B VDD 0.48fF
C65017 PAND2X1_569/B PAND2X1_324/Y 0.01fF
C65018 POR2X1_136/O POR2X1_136/Y 0.04fF
C65019 POR2X1_750/B PAND2X1_179/O 0.04fF
C65020 PAND2X1_213/Y PAND2X1_161/Y 0.06fF
C65021 POR2X1_368/Y POR2X1_283/A 0.02fF
C65022 INPUT_3 POR2X1_9/Y 0.26fF
C65023 PAND2X1_60/B POR2X1_788/B 1.74fF
C65024 POR2X1_29/Y PAND2X1_63/B 0.03fF
C65025 POR2X1_824/O POR2X1_236/Y 0.01fF
C65026 POR2X1_366/Y POR2X1_703/Y 0.02fF
C65027 POR2X1_567/A POR2X1_542/m4_208_n4# 0.03fF
C65028 PAND2X1_348/Y PAND2X1_359/B 0.14fF
C65029 POR2X1_183/Y PAND2X1_114/CTRL2 0.00fF
C65030 PAND2X1_838/B POR2X1_827/CTRL2 0.01fF
C65031 POR2X1_66/B PAND2X1_56/A 0.03fF
C65032 PAND2X1_863/B POR2X1_595/CTRL2 0.01fF
C65033 POR2X1_204/CTRL2 POR2X1_260/A 0.01fF
C65034 PAND2X1_94/A PAND2X1_6/A 4.15fF
C65035 POR2X1_761/Y PAND2X1_854/A 0.02fF
C65036 POR2X1_137/Y POR2X1_361/O 0.01fF
C65037 POR2X1_101/Y POR2X1_576/Y 0.05fF
C65038 PAND2X1_41/B D_INPUT_4 0.12fF
C65039 POR2X1_778/B PAND2X1_103/CTRL 0.00fF
C65040 POR2X1_712/Y POR2X1_260/A 0.01fF
C65041 PAND2X1_824/B POR2X1_222/Y 0.07fF
C65042 PAND2X1_48/B POR2X1_334/Y 0.07fF
C65043 POR2X1_322/Y PAND2X1_168/O 0.00fF
C65044 PAND2X1_801/CTRL POR2X1_236/Y 0.02fF
C65045 POR2X1_40/Y PAND2X1_327/CTRL 0.01fF
C65046 POR2X1_502/A POR2X1_383/O 0.04fF
C65047 POR2X1_43/B PAND2X1_308/Y 1.38fF
C65048 POR2X1_322/CTRL POR2X1_373/Y 0.01fF
C65049 D_GATE_222 POR2X1_259/B 0.06fF
C65050 POR2X1_327/Y POR2X1_264/Y 0.00fF
C65051 PAND2X1_317/Y PAND2X1_703/CTRL 0.08fF
C65052 POR2X1_78/A POR2X1_863/A 0.06fF
C65053 PAND2X1_686/CTRL POR2X1_73/Y 0.00fF
C65054 PAND2X1_73/Y POR2X1_76/B 0.01fF
C65055 POR2X1_567/B PAND2X1_438/CTRL 0.13fF
C65056 PAND2X1_432/O PAND2X1_72/A 0.03fF
C65057 PAND2X1_714/O PAND2X1_714/B 0.00fF
C65058 POR2X1_500/Y POR2X1_260/A 0.03fF
C65059 POR2X1_334/B PAND2X1_48/A 0.05fF
C65060 PAND2X1_150/CTRL POR2X1_260/A 0.01fF
C65061 POR2X1_553/A POR2X1_228/Y 0.03fF
C65062 POR2X1_777/B POR2X1_717/B 0.48fF
C65063 POR2X1_40/Y POR2X1_167/Y 0.53fF
C65064 POR2X1_416/B POR2X1_376/Y 0.23fF
C65065 PAND2X1_723/A POR2X1_7/A 0.15fF
C65066 PAND2X1_6/Y POR2X1_228/CTRL2 0.00fF
C65067 POR2X1_60/A PAND2X1_242/Y 0.05fF
C65068 POR2X1_168/A PAND2X1_65/B 0.01fF
C65069 POR2X1_406/Y PAND2X1_339/CTRL2 0.03fF
C65070 PAND2X1_175/B PAND2X1_861/CTRL 0.01fF
C65071 POR2X1_110/Y POR2X1_693/Y 0.03fF
C65072 POR2X1_411/B PAND2X1_9/Y 0.03fF
C65073 POR2X1_655/CTRL POR2X1_646/Y 0.00fF
C65074 POR2X1_390/B POR2X1_538/A 0.44fF
C65075 POR2X1_551/CTRL POR2X1_854/B 0.15fF
C65076 POR2X1_725/Y POR2X1_151/CTRL 0.03fF
C65077 PAND2X1_704/CTRL2 POR2X1_142/Y 0.10fF
C65078 POR2X1_814/B POR2X1_343/B 0.01fF
C65079 POR2X1_383/A POR2X1_773/B 0.03fF
C65080 POR2X1_673/Y POR2X1_550/Y 0.03fF
C65081 POR2X1_219/B PAND2X1_394/CTRL2 0.09fF
C65082 POR2X1_416/B PAND2X1_556/B 0.00fF
C65083 POR2X1_119/Y PAND2X1_716/CTRL 0.12fF
C65084 POR2X1_509/CTRL VDD 0.00fF
C65085 PAND2X1_358/a_16_344# PAND2X1_351/Y 0.02fF
C65086 POR2X1_66/B POR2X1_661/A 0.10fF
C65087 PAND2X1_23/Y POR2X1_343/CTRL2 0.03fF
C65088 PAND2X1_683/CTRL2 POR2X1_596/A 0.01fF
C65089 VDD POR2X1_181/Y 0.00fF
C65090 PAND2X1_55/Y POR2X1_169/A 2.23fF
C65091 POR2X1_510/Y POR2X1_186/B 0.06fF
C65092 PAND2X1_84/Y PAND2X1_332/Y 0.03fF
C65093 POR2X1_346/B POR2X1_61/CTRL 0.00fF
C65094 POR2X1_416/B PAND2X1_254/Y 0.05fF
C65095 PAND2X1_341/B PAND2X1_341/A 0.12fF
C65096 POR2X1_471/A POR2X1_446/B 0.03fF
C65097 POR2X1_16/A PAND2X1_317/CTRL2 0.03fF
C65098 POR2X1_76/Y PAND2X1_72/A 0.02fF
C65099 VDD PAND2X1_135/O 0.00fF
C65100 POR2X1_661/CTRL POR2X1_661/A 0.06fF
C65101 PAND2X1_490/a_56_28# POR2X1_4/Y 0.00fF
C65102 POR2X1_709/A POR2X1_260/B 1.05fF
C65103 POR2X1_110/O POR2X1_387/Y 0.05fF
C65104 POR2X1_736/O POR2X1_188/Y 0.02fF
C65105 POR2X1_329/A PAND2X1_361/CTRL 0.01fF
C65106 VDD POR2X1_535/CTRL 0.00fF
C65107 POR2X1_614/A POR2X1_383/Y 0.03fF
C65108 POR2X1_647/B POR2X1_866/A 0.01fF
C65109 POR2X1_832/CTRL2 POR2X1_661/A 0.05fF
C65110 POR2X1_43/B POR2X1_77/Y 0.13fF
C65111 PAND2X1_217/O PAND2X1_576/B 0.05fF
C65112 POR2X1_312/O POR2X1_77/Y 0.01fF
C65113 POR2X1_416/B POR2X1_599/A 0.10fF
C65114 POR2X1_624/Y POR2X1_499/CTRL2 0.01fF
C65115 PAND2X1_93/B POR2X1_243/B 0.02fF
C65116 PAND2X1_563/A POR2X1_394/A 0.05fF
C65117 POR2X1_740/Y PAND2X1_72/A 0.08fF
C65118 PAND2X1_466/A POR2X1_102/Y 0.02fF
C65119 POR2X1_447/B PAND2X1_823/CTRL2 -0.00fF
C65120 PAND2X1_94/CTRL2 POR2X1_202/A 0.02fF
C65121 PAND2X1_551/A PAND2X1_326/O 0.02fF
C65122 POR2X1_814/A POR2X1_186/Y 0.07fF
C65123 PAND2X1_641/CTRL2 PAND2X1_341/B 0.00fF
C65124 POR2X1_274/A PAND2X1_93/B 0.03fF
C65125 POR2X1_760/A PAND2X1_557/A 0.06fF
C65126 POR2X1_96/A PAND2X1_860/A 0.03fF
C65127 PAND2X1_785/CTRL POR2X1_77/Y 0.01fF
C65128 POR2X1_262/Y POR2X1_102/Y 0.03fF
C65129 POR2X1_796/O PAND2X1_52/B 0.01fF
C65130 POR2X1_38/B POR2X1_77/Y 0.03fF
C65131 PAND2X1_212/CTRL2 PAND2X1_352/A 0.01fF
C65132 PAND2X1_124/Y PAND2X1_576/B 0.08fF
C65133 POR2X1_16/A POR2X1_4/Y 0.03fF
C65134 PAND2X1_641/O PAND2X1_476/A 0.00fF
C65135 PAND2X1_858/O POR2X1_129/Y 0.02fF
C65136 PAND2X1_459/CTRL2 PAND2X1_9/Y 0.03fF
C65137 PAND2X1_351/m4_208_n4# POR2X1_153/Y 0.04fF
C65138 POR2X1_864/A POR2X1_783/a_16_28# 0.02fF
C65139 PAND2X1_675/a_16_344# POR2X1_283/A 0.01fF
C65140 POR2X1_41/O POR2X1_41/Y 0.01fF
C65141 PAND2X1_294/O POR2X1_60/A 0.20fF
C65142 POR2X1_24/CTRL2 PAND2X1_9/Y 0.01fF
C65143 PAND2X1_20/A POR2X1_445/A 7.21fF
C65144 PAND2X1_217/B PAND2X1_203/CTRL2 0.01fF
C65145 PAND2X1_488/O POR2X1_556/A 0.04fF
C65146 POR2X1_634/A PAND2X1_59/a_56_28# 0.00fF
C65147 INPUT_6 PAND2X1_72/A 0.03fF
C65148 D_INPUT_5 POR2X1_638/A 0.00fF
C65149 PAND2X1_93/B POR2X1_269/A 0.01fF
C65150 PAND2X1_472/A POR2X1_825/Y 0.03fF
C65151 POR2X1_818/CTRL POR2X1_734/A 0.14fF
C65152 POR2X1_741/CTRL2 POR2X1_186/B 0.01fF
C65153 POR2X1_260/B PAND2X1_58/A 0.14fF
C65154 POR2X1_411/B POR2X1_609/a_16_28# 0.02fF
C65155 PAND2X1_93/B POR2X1_602/A 0.01fF
C65156 POR2X1_20/B POR2X1_432/Y 0.01fF
C65157 POR2X1_77/CTRL POR2X1_40/Y 0.03fF
C65158 POR2X1_66/B POR2X1_610/O 0.16fF
C65159 PAND2X1_282/CTRL2 POR2X1_590/A 0.01fF
C65160 POR2X1_78/B POR2X1_318/O 0.03fF
C65161 POR2X1_863/A PAND2X1_173/CTRL 0.05fF
C65162 POR2X1_150/Y PAND2X1_804/A 0.01fF
C65163 PAND2X1_603/CTRL2 POR2X1_78/A 0.03fF
C65164 POR2X1_422/CTRL2 POR2X1_72/B 0.03fF
C65165 POR2X1_445/A POR2X1_814/B 3.01fF
C65166 POR2X1_594/Y POR2X1_329/A 0.00fF
C65167 PAND2X1_245/CTRL POR2X1_296/B 0.00fF
C65168 POR2X1_859/a_56_344# INPUT_0 0.03fF
C65169 PAND2X1_61/O POR2X1_60/A 0.06fF
C65170 PAND2X1_98/O INPUT_0 0.09fF
C65171 POR2X1_83/B POR2X1_67/A 0.12fF
C65172 POR2X1_175/A POR2X1_567/B 0.05fF
C65173 POR2X1_327/Y POR2X1_343/Y 0.05fF
C65174 POR2X1_477/B POR2X1_477/Y 0.00fF
C65175 POR2X1_283/A POR2X1_310/CTRL2 0.05fF
C65176 PAND2X1_746/CTRL2 PAND2X1_52/B 0.04fF
C65177 POR2X1_153/Y PAND2X1_351/A 0.05fF
C65178 POR2X1_591/A PAND2X1_722/a_16_344# 0.03fF
C65179 POR2X1_411/B PAND2X1_216/O 0.03fF
C65180 POR2X1_669/B PAND2X1_706/CTRL 0.08fF
C65181 POR2X1_54/Y PAND2X1_57/B 0.03fF
C65182 PAND2X1_267/Y PAND2X1_741/B 0.03fF
C65183 POR2X1_23/a_16_28# POR2X1_14/Y 0.03fF
C65184 POR2X1_860/A POR2X1_218/Y 0.02fF
C65185 POR2X1_116/A POR2X1_717/Y 0.01fF
C65186 POR2X1_23/Y PAND2X1_332/O 0.01fF
C65187 POR2X1_51/A D_INPUT_5 0.00fF
C65188 POR2X1_774/A PAND2X1_72/A 0.03fF
C65189 POR2X1_416/Y POR2X1_411/A 0.09fF
C65190 POR2X1_43/B PAND2X1_449/O 0.04fF
C65191 POR2X1_83/B PAND2X1_215/a_76_28# 0.02fF
C65192 POR2X1_311/Y PAND2X1_557/A 0.03fF
C65193 POR2X1_807/A POR2X1_807/a_76_344# 0.01fF
C65194 POR2X1_48/A PAND2X1_713/B 0.33fF
C65195 PAND2X1_838/O POR2X1_42/Y 0.02fF
C65196 PAND2X1_57/B POR2X1_202/A 0.08fF
C65197 POR2X1_682/O POR2X1_32/A 0.02fF
C65198 POR2X1_517/O POR2X1_669/B 0.16fF
C65199 POR2X1_174/B PAND2X1_41/B 0.07fF
C65200 POR2X1_333/A POR2X1_750/B 0.16fF
C65201 PAND2X1_73/Y POR2X1_456/O 0.02fF
C65202 POR2X1_97/A PAND2X1_90/Y 4.80fF
C65203 POR2X1_76/A PAND2X1_131/a_76_28# 0.02fF
C65204 POR2X1_54/Y POR2X1_642/CTRL2 0.03fF
C65205 POR2X1_707/B PAND2X1_428/O 0.03fF
C65206 POR2X1_484/CTRL2 VDD 0.00fF
C65207 PAND2X1_6/Y POR2X1_556/A 0.06fF
C65208 POR2X1_499/A POR2X1_778/B 0.03fF
C65209 POR2X1_496/Y POR2X1_236/Y 0.07fF
C65210 PAND2X1_790/O POR2X1_42/Y 0.15fF
C65211 POR2X1_65/A POR2X1_295/CTRL2 0.03fF
C65212 POR2X1_502/A POR2X1_856/B 0.03fF
C65213 POR2X1_66/B POR2X1_461/O 0.15fF
C65214 POR2X1_127/O VDD 0.00fF
C65215 PAND2X1_793/Y PAND2X1_489/O 0.03fF
C65216 POR2X1_620/A PAND2X1_8/Y 0.04fF
C65217 POR2X1_814/B PAND2X1_585/O 0.04fF
C65218 POR2X1_644/B PAND2X1_57/B 0.01fF
C65219 POR2X1_78/B POR2X1_555/B 0.05fF
C65220 POR2X1_451/O POR2X1_750/B 0.01fF
C65221 POR2X1_14/Y POR2X1_236/CTRL 0.01fF
C65222 POR2X1_413/A PAND2X1_646/CTRL 0.01fF
C65223 POR2X1_83/B PAND2X1_733/Y 0.01fF
C65224 POR2X1_66/A POR2X1_121/Y 0.03fF
C65225 PAND2X1_852/B POR2X1_411/B 0.01fF
C65226 POR2X1_355/CTRL2 POR2X1_355/A 0.01fF
C65227 PAND2X1_117/CTRL POR2X1_558/B 0.00fF
C65228 PAND2X1_117/O POR2X1_493/A 0.02fF
C65229 INPUT_2 INPUT_3 0.29fF
C65230 PAND2X1_169/Y PAND2X1_714/A 0.19fF
C65231 POR2X1_602/B POR2X1_718/A 0.03fF
C65232 POR2X1_852/B POR2X1_186/Y 0.07fF
C65233 POR2X1_729/a_16_28# POR2X1_452/Y 0.02fF
C65234 PAND2X1_213/Y POR2X1_441/Y 0.03fF
C65235 PAND2X1_807/B VDD 0.30fF
C65236 POR2X1_515/O PAND2X1_20/A 0.01fF
C65237 PAND2X1_239/a_16_344# POR2X1_578/Y 0.01fF
C65238 POR2X1_661/Y PAND2X1_57/B 0.14fF
C65239 POR2X1_626/CTRL2 POR2X1_55/Y 0.01fF
C65240 POR2X1_760/A PAND2X1_723/A 0.07fF
C65241 POR2X1_466/Y VDD 0.10fF
C65242 POR2X1_555/A PAND2X1_41/B 0.03fF
C65243 D_INPUT_0 POR2X1_294/B 0.96fF
C65244 POR2X1_808/B POR2X1_800/A 0.07fF
C65245 PAND2X1_733/A POR2X1_236/Y 0.07fF
C65246 POR2X1_83/B PAND2X1_198/Y 0.00fF
C65247 PAND2X1_48/CTRL2 POR2X1_330/Y 0.02fF
C65248 POR2X1_148/O PAND2X1_69/A 0.01fF
C65249 POR2X1_78/B POR2X1_330/Y 0.13fF
C65250 POR2X1_457/O POR2X1_370/Y 0.16fF
C65251 POR2X1_118/CTRL2 POR2X1_118/Y 0.01fF
C65252 PAND2X1_660/O PAND2X1_660/B 0.02fF
C65253 POR2X1_814/B PAND2X1_395/a_16_344# 0.02fF
C65254 POR2X1_47/CTRL2 POR2X1_32/A 0.02fF
C65255 POR2X1_590/A POR2X1_208/O 0.16fF
C65256 POR2X1_841/B POR2X1_804/A 3.35fF
C65257 INPUT_1 POR2X1_623/Y 0.04fF
C65258 PAND2X1_96/B POR2X1_260/B 0.73fF
C65259 POR2X1_820/B POR2X1_820/A 0.59fF
C65260 POR2X1_458/O PAND2X1_69/A 0.25fF
C65261 PAND2X1_580/a_16_344# PAND2X1_771/Y 0.07fF
C65262 POR2X1_857/B POR2X1_836/A 0.03fF
C65263 PAND2X1_206/A PAND2X1_99/Y 0.00fF
C65264 PAND2X1_241/O POR2X1_83/B 0.00fF
C65265 POR2X1_683/CTRL2 POR2X1_40/Y 0.01fF
C65266 POR2X1_143/CTRL POR2X1_40/Y 0.01fF
C65267 PAND2X1_392/CTRL POR2X1_816/A 0.01fF
C65268 POR2X1_370/Y POR2X1_543/A 0.01fF
C65269 PAND2X1_58/A PAND2X1_369/O 0.03fF
C65270 POR2X1_544/A PAND2X1_41/B 0.01fF
C65271 PAND2X1_862/B PAND2X1_217/B 0.03fF
C65272 PAND2X1_137/Y POR2X1_40/Y 0.05fF
C65273 POR2X1_22/A POR2X1_32/A 0.14fF
C65274 PAND2X1_58/A PAND2X1_55/Y 1.14fF
C65275 PAND2X1_7/O POR2X1_555/B 0.04fF
C65276 PAND2X1_650/A POR2X1_826/Y 0.01fF
C65277 POR2X1_602/CTRL PAND2X1_60/B 0.01fF
C65278 POR2X1_788/A PAND2X1_144/CTRL 0.01fF
C65279 POR2X1_63/CTRL2 POR2X1_83/B 0.00fF
C65280 POR2X1_625/CTRL VDD 0.00fF
C65281 POR2X1_417/Y POR2X1_372/Y 0.20fF
C65282 POR2X1_558/A POR2X1_260/B 0.01fF
C65283 PAND2X1_543/CTRL2 POR2X1_236/Y 0.01fF
C65284 POR2X1_220/B PAND2X1_69/A 0.03fF
C65285 PAND2X1_425/Y PAND2X1_157/CTRL2 0.01fF
C65286 PAND2X1_808/Y PAND2X1_772/O 0.02fF
C65287 PAND2X1_73/Y PAND2X1_744/O 0.02fF
C65288 POR2X1_68/A POR2X1_174/A 0.03fF
C65289 POR2X1_828/Y PAND2X1_760/CTRL 0.01fF
C65290 POR2X1_590/A POR2X1_391/Y 0.03fF
C65291 POR2X1_300/a_56_344# POR2X1_102/Y 0.00fF
C65292 POR2X1_487/Y POR2X1_488/Y 0.02fF
C65293 POR2X1_150/Y PAND2X1_348/A 0.07fF
C65294 PAND2X1_58/A POR2X1_788/Y 0.01fF
C65295 POR2X1_814/B POR2X1_114/Y 0.13fF
C65296 POR2X1_56/B POR2X1_423/Y 0.10fF
C65297 POR2X1_29/Y POR2X1_32/A 0.04fF
C65298 PAND2X1_667/CTRL2 POR2X1_546/A 0.01fF
C65299 POR2X1_660/Y PAND2X1_69/A 0.03fF
C65300 PAND2X1_94/A PAND2X1_24/O 0.17fF
C65301 PAND2X1_309/CTRL POR2X1_543/A 0.01fF
C65302 POR2X1_344/A PAND2X1_65/B 0.54fF
C65303 PAND2X1_58/A POR2X1_402/A 0.64fF
C65304 PAND2X1_39/B POR2X1_260/A 0.20fF
C65305 PAND2X1_474/Y PAND2X1_84/Y 0.03fF
C65306 POR2X1_504/O POR2X1_20/B 0.01fF
C65307 PAND2X1_128/CTRL2 POR2X1_127/Y 0.01fF
C65308 POR2X1_83/B PAND2X1_642/B 0.02fF
C65309 POR2X1_20/B POR2X1_394/A 0.25fF
C65310 PAND2X1_223/O POR2X1_7/B 0.04fF
C65311 POR2X1_657/CTRL POR2X1_112/Y 0.01fF
C65312 PAND2X1_140/A PAND2X1_771/Y 0.17fF
C65313 PAND2X1_140/Y PAND2X1_139/Y 0.01fF
C65314 POR2X1_57/A PAND2X1_722/O 0.01fF
C65315 PAND2X1_558/Y PAND2X1_717/CTRL 0.00fF
C65316 PAND2X1_865/Y PAND2X1_717/A 0.03fF
C65317 POR2X1_509/m4_208_n4# PAND2X1_41/B 0.07fF
C65318 POR2X1_383/A POR2X1_286/CTRL2 0.01fF
C65319 POR2X1_674/Y POR2X1_594/A 0.02fF
C65320 POR2X1_48/A POR2X1_765/Y 0.03fF
C65321 POR2X1_83/B PAND2X1_243/CTRL2 0.03fF
C65322 POR2X1_68/B POR2X1_390/CTRL2 0.01fF
C65323 POR2X1_49/Y PAND2X1_466/O 0.17fF
C65324 PAND2X1_63/Y PAND2X1_20/A 0.06fF
C65325 POR2X1_278/Y PAND2X1_740/Y -0.01fF
C65326 POR2X1_32/A POR2X1_526/Y 0.01fF
C65327 PAND2X1_48/B POR2X1_475/A 0.07fF
C65328 POR2X1_493/B POR2X1_260/B 0.01fF
C65329 PAND2X1_695/CTRL2 PAND2X1_48/B 0.03fF
C65330 POR2X1_763/A PAND2X1_709/CTRL2 -0.01fF
C65331 PAND2X1_862/B VDD 0.53fF
C65332 PAND2X1_129/CTRL2 POR2X1_814/A 0.01fF
C65333 POR2X1_366/Y PAND2X1_90/Y 0.07fF
C65334 PAND2X1_687/CTRL POR2X1_597/Y 0.03fF
C65335 PAND2X1_90/Y POR2X1_294/B 0.46fF
C65336 POR2X1_327/Y POR2X1_624/Y 0.00fF
C65337 PAND2X1_495/O PAND2X1_20/A 0.02fF
C65338 POR2X1_662/Y POR2X1_741/a_16_28# 0.01fF
C65339 POR2X1_686/A POR2X1_68/A 0.00fF
C65340 PAND2X1_668/CTRL PAND2X1_673/Y 0.01fF
C65341 PAND2X1_684/O POR2X1_260/B 0.03fF
C65342 PAND2X1_3/O PAND2X1_3/A 0.08fF
C65343 POR2X1_315/CTRL2 PAND2X1_803/A 0.00fF
C65344 POR2X1_49/Y POR2X1_521/O 0.18fF
C65345 POR2X1_502/A POR2X1_722/Y 0.04fF
C65346 POR2X1_319/A POR2X1_724/B 0.12fF
C65347 PAND2X1_44/O PAND2X1_32/B 0.03fF
C65348 PAND2X1_345/CTRL2 PAND2X1_555/A 0.01fF
C65349 POR2X1_83/B PAND2X1_168/O 0.01fF
C65350 POR2X1_347/A PAND2X1_94/CTRL2 0.04fF
C65351 PAND2X1_116/CTRL POR2X1_183/Y 0.00fF
C65352 PAND2X1_57/B PAND2X1_322/O 0.00fF
C65353 POR2X1_590/A PAND2X1_528/CTRL2 0.05fF
C65354 PAND2X1_119/CTRL POR2X1_654/B 0.01fF
C65355 POR2X1_750/B POR2X1_788/B 0.03fF
C65356 PAND2X1_23/Y POR2X1_284/B 0.02fF
C65357 POR2X1_689/A INPUT_0 0.03fF
C65358 PAND2X1_48/B POR2X1_349/Y 0.04fF
C65359 PAND2X1_412/CTRL PAND2X1_32/B 0.01fF
C65360 PAND2X1_731/O PAND2X1_738/B 0.03fF
C65361 POR2X1_102/Y PAND2X1_572/m4_208_n4# 0.12fF
C65362 PAND2X1_496/O INPUT_0 0.09fF
C65363 POR2X1_640/Y POR2X1_532/A 0.05fF
C65364 PAND2X1_63/Y POR2X1_814/B 0.03fF
C65365 POR2X1_65/CTRL POR2X1_39/B 0.13fF
C65366 POR2X1_654/B POR2X1_68/B 0.02fF
C65367 POR2X1_309/a_16_28# POR2X1_283/A 0.03fF
C65368 PAND2X1_521/O POR2X1_750/A 0.03fF
C65369 POR2X1_351/Y PAND2X1_65/B 0.02fF
C65370 POR2X1_244/B POR2X1_740/Y 0.05fF
C65371 POR2X1_83/B PAND2X1_550/B 0.06fF
C65372 PAND2X1_341/a_16_344# INPUT_0 0.03fF
C65373 POR2X1_790/B VDD 0.15fF
C65374 POR2X1_516/A POR2X1_60/A 0.00fF
C65375 POR2X1_734/A PAND2X1_518/a_56_28# 0.00fF
C65376 POR2X1_49/Y PAND2X1_814/a_16_344# 0.02fF
C65377 PAND2X1_94/A POR2X1_35/a_16_28# 0.03fF
C65378 PAND2X1_58/A PAND2X1_28/O 0.05fF
C65379 PAND2X1_495/O POR2X1_814/B 0.01fF
C65380 POR2X1_356/A PAND2X1_524/a_76_28# 0.04fF
C65381 POR2X1_278/Y PAND2X1_675/A 0.07fF
C65382 POR2X1_174/B POR2X1_502/CTRL 0.02fF
C65383 POR2X1_298/Y PAND2X1_308/Y 0.00fF
C65384 POR2X1_435/Y POR2X1_788/Y 0.09fF
C65385 POR2X1_68/B POR2X1_5/Y 0.03fF
C65386 POR2X1_578/Y POR2X1_785/A 0.03fF
C65387 PAND2X1_580/O PAND2X1_580/B 0.00fF
C65388 POR2X1_625/a_16_28# POR2X1_90/Y 0.05fF
C65389 POR2X1_788/O PAND2X1_60/B 0.17fF
C65390 PAND2X1_59/B PAND2X1_18/B 0.81fF
C65391 PAND2X1_639/O POR2X1_408/Y 0.19fF
C65392 POR2X1_192/Y POR2X1_35/Y 0.05fF
C65393 POR2X1_814/A POR2X1_717/B 0.07fF
C65394 POR2X1_327/Y PAND2X1_431/a_76_28# 0.05fF
C65395 POR2X1_113/Y POR2X1_814/B 0.07fF
C65396 PAND2X1_743/CTRL VDD 0.00fF
C65397 POR2X1_556/A POR2X1_632/Y 0.03fF
C65398 PAND2X1_94/A PAND2X1_235/O 0.18fF
C65399 POR2X1_502/A POR2X1_565/O 0.02fF
C65400 PAND2X1_20/A POR2X1_260/A 17.01fF
C65401 PAND2X1_115/a_16_344# PAND2X1_115/B 0.02fF
C65402 POR2X1_52/A PAND2X1_717/O 0.15fF
C65403 POR2X1_60/A PAND2X1_301/CTRL 0.01fF
C65404 POR2X1_46/Y PAND2X1_546/CTRL 0.01fF
C65405 POR2X1_416/B POR2X1_441/Y 0.03fF
C65406 POR2X1_567/B POR2X1_337/Y 0.10fF
C65407 POR2X1_811/O POR2X1_294/A 0.05fF
C65408 POR2X1_270/Y POR2X1_370/a_16_28# 0.00fF
C65409 PAND2X1_700/O POR2X1_532/A 0.06fF
C65410 PAND2X1_864/O PAND2X1_810/A 0.02fF
C65411 POR2X1_497/Y POR2X1_91/Y 0.07fF
C65412 POR2X1_627/CTRL2 POR2X1_7/A 0.03fF
C65413 POR2X1_131/Y PAND2X1_140/CTRL2 0.01fF
C65414 POR2X1_257/A POR2X1_39/B 0.79fF
C65415 POR2X1_856/B POR2X1_188/Y 0.03fF
C65416 PAND2X1_96/B PAND2X1_516/CTRL 0.01fF
C65417 POR2X1_134/Y PAND2X1_137/Y 0.01fF
C65418 PAND2X1_651/Y POR2X1_372/Y 0.10fF
C65419 POR2X1_13/A POR2X1_9/CTRL2 0.01fF
C65420 POR2X1_65/A POR2X1_527/CTRL 0.01fF
C65421 PAND2X1_357/Y POR2X1_42/Y 0.03fF
C65422 POR2X1_66/B PAND2X1_481/O 0.10fF
C65423 PAND2X1_755/CTRL2 PAND2X1_60/B 0.01fF
C65424 POR2X1_376/B PAND2X1_155/CTRL2 0.00fF
C65425 POR2X1_786/A PAND2X1_69/A 0.16fF
C65426 POR2X1_327/O PAND2X1_63/Y 0.16fF
C65427 PAND2X1_48/B PAND2X1_146/a_76_28# 0.01fF
C65428 POR2X1_37/Y PAND2X1_500/CTRL 0.03fF
C65429 POR2X1_660/Y POR2X1_512/CTRL 0.01fF
C65430 POR2X1_96/Y POR2X1_409/B 0.07fF
C65431 POR2X1_20/CTRL POR2X1_68/B 0.00fF
C65432 POR2X1_814/B POR2X1_260/A 20.29fF
C65433 POR2X1_529/Y INPUT_0 0.07fF
C65434 POR2X1_16/A PAND2X1_714/A 0.04fF
C65435 POR2X1_5/Y POR2X1_172/O 0.34fF
C65436 PAND2X1_682/CTRL POR2X1_407/A -0.02fF
C65437 GATE_741 PAND2X1_854/A 0.02fF
C65438 POR2X1_40/Y PAND2X1_853/B 0.09fF
C65439 POR2X1_124/a_76_344# PAND2X1_96/B 0.01fF
C65440 PAND2X1_64/CTRL D_INPUT_4 0.01fF
C65441 PAND2X1_852/CTRL2 POR2X1_73/Y 0.03fF
C65442 PAND2X1_96/B PAND2X1_55/Y 0.30fF
C65443 PAND2X1_357/Y POR2X1_309/Y 0.03fF
C65444 POR2X1_616/Y POR2X1_83/B 0.35fF
C65445 POR2X1_236/Y PAND2X1_124/CTRL 0.04fF
C65446 POR2X1_16/A PAND2X1_645/CTRL2 0.01fF
C65447 POR2X1_43/B POR2X1_52/Y 0.14fF
C65448 PAND2X1_659/Y PAND2X1_473/m4_208_n4# 0.22fF
C65449 PAND2X1_484/CTRL PAND2X1_41/B 0.00fF
C65450 POR2X1_516/O PAND2X1_6/A 0.04fF
C65451 POR2X1_65/A PAND2X1_120/CTRL2 0.03fF
C65452 POR2X1_677/CTRL2 POR2X1_129/Y 0.01fF
C65453 POR2X1_49/Y POR2X1_177/CTRL 0.01fF
C65454 POR2X1_712/Y POR2X1_713/Y 0.03fF
C65455 POR2X1_7/B POR2X1_387/Y 0.09fF
C65456 POR2X1_114/B POR2X1_804/A 0.03fF
C65457 PAND2X1_216/B PAND2X1_473/B 0.41fF
C65458 POR2X1_7/A PAND2X1_515/O 0.08fF
C65459 POR2X1_186/Y POR2X1_151/Y 0.18fF
C65460 PAND2X1_798/B PAND2X1_575/CTRL2 0.01fF
C65461 PAND2X1_639/Y POR2X1_14/Y 0.02fF
C65462 POR2X1_325/A POR2X1_260/A 0.03fF
C65463 POR2X1_814/B POR2X1_363/A 0.01fF
C65464 PAND2X1_364/B PAND2X1_656/A 0.02fF
C65465 POR2X1_493/CTRL2 POR2X1_572/B 0.02fF
C65466 POR2X1_330/Y POR2X1_294/A 0.03fF
C65467 POR2X1_188/A POR2X1_737/A 0.02fF
C65468 PAND2X1_344/CTRL PAND2X1_514/Y 0.01fF
C65469 PAND2X1_175/B POR2X1_293/Y 0.03fF
C65470 POR2X1_773/B INPUT_0 0.12fF
C65471 POR2X1_83/CTRL2 PAND2X1_35/Y 0.01fF
C65472 POR2X1_861/a_76_344# POR2X1_501/B 0.00fF
C65473 PAND2X1_90/Y PAND2X1_533/O 0.29fF
C65474 POR2X1_334/CTRL2 PAND2X1_57/B 0.04fF
C65475 PAND2X1_96/B POR2X1_402/A 0.00fF
C65476 POR2X1_78/A PAND2X1_134/a_16_344# 0.01fF
C65477 PAND2X1_480/CTRL POR2X1_236/Y 0.01fF
C65478 POR2X1_164/O PAND2X1_565/A 0.00fF
C65479 PAND2X1_217/B PAND2X1_716/B 0.03fF
C65480 POR2X1_593/B PAND2X1_48/A 0.05fF
C65481 PAND2X1_308/CTRL VDD 0.00fF
C65482 PAND2X1_743/CTRL PAND2X1_32/B 0.03fF
C65483 POR2X1_407/A POR2X1_596/A 0.07fF
C65484 POR2X1_174/A POR2X1_169/A 0.03fF
C65485 POR2X1_3/A POR2X1_581/O 0.03fF
C65486 POR2X1_36/B POR2X1_581/CTRL 0.01fF
C65487 PAND2X1_651/Y POR2X1_239/O 0.00fF
C65488 POR2X1_528/Y POR2X1_42/Y 0.10fF
C65489 PAND2X1_824/B POR2X1_207/O 0.06fF
C65490 POR2X1_276/A POR2X1_276/O 0.02fF
C65491 PAND2X1_101/a_16_344# PAND2X1_99/Y 0.01fF
C65492 POR2X1_760/A PAND2X1_405/O 0.01fF
C65493 POR2X1_347/A PAND2X1_57/B 0.07fF
C65494 PAND2X1_94/A PAND2X1_92/a_56_28# 0.00fF
C65495 VDD POR2X1_673/B 0.01fF
C65496 POR2X1_414/Y POR2X1_4/Y 0.01fF
C65497 POR2X1_265/Y POR2X1_5/Y 0.79fF
C65498 POR2X1_861/A POR2X1_860/A 0.06fF
C65499 POR2X1_369/a_16_28# POR2X1_236/Y 0.02fF
C65500 PAND2X1_797/Y PAND2X1_731/B 0.03fF
C65501 POR2X1_327/O POR2X1_260/A 0.01fF
C65502 PAND2X1_23/Y PAND2X1_94/A 0.23fF
C65503 D_INPUT_4 GND 0.41fF
C65504 PAND2X1_2/m4_208_n4# GND 0.00fF
C65505 POR2X1_673/B GND 0.21fF
C65506 PAND2X1_54/m4_208_n4# GND -0.00fF
C65507 PAND2X1_670/CTRL GND 0.02fF
C65508 POR2X1_685/B GND 0.16fF
C65509 PAND2X1_32/B GND 2.06fF
C65510 PAND2X1_681/m4_208_n4# GND 0.00fF
C65511 PAND2X1_692/m4_208_n4# GND -0.00fF
C65512 POR2X1_91/Y GND 1.00fF
C65513 POR2X1_80/CTRL GND 0.02fF
C65514 POR2X1_210/B GND 0.21fF
C65515 POR2X1_156/Y GND 0.18fF
C65516 POR2X1_260/A GND 1.66fF
C65517 PAND2X1_158/m4_208_n4# GND 0.00fF
C65518 PAND2X1_149/A GND 0.46fF
C65519 POR2X1_142/Y GND 0.26fF
C65520 PAND2X1_147/m4_208_n4# GND 0.00fF
C65521 POR2X1_166/Y GND 0.17fF
C65522 POR2X1_167/Y GND 0.03fF
C65523 PAND2X1_169/CTRL GND 0.02fF
C65524 PAND2X1_114/m4_208_n4# GND -0.00fF
C65525 POR2X1_128/B GND 0.23fF
C65526 PAND2X1_125/m4_208_n4# GND 0.00fF
C65527 POR2X1_138/A GND 0.38fF
C65528 POR2X1_514/m4_208_n4# GND -0.00fF
C65529 POR2X1_113/B GND 0.14fF
C65530 PAND2X1_103/m4_208_n4# GND 0.00fF
C65531 POR2X1_162/Y GND -0.26fF
C65532 POR2X1_161/Y GND -0.15fF
C65533 POR2X1_162/m4_208_n4# GND 0.00fF
C65534 POR2X1_173/Y GND 0.17fF
C65535 POR2X1_173/CTRL GND 0.02fF
C65536 POR2X1_199/B GND 0.08fF
C65537 PAND2X1_41/Y GND 0.13fF
C65538 POR2X1_195/m4_208_n4# GND 0.00fF
C65539 POR2X1_151/Y GND 0.18fF
C65540 POR2X1_186/B GND 0.81fF
C65541 POR2X1_141/A GND 0.29fF
C65542 PAND2X1_858/Y GND -0.10fF
C65543 PAND2X1_862/m4_208_n4# GND -0.00fF
C65544 PAND2X1_858/B GND 0.20fF
C65545 PAND2X1_840/Y GND 0.35fF
C65546 PAND2X1_841/Y GND 0.12fF
C65547 PAND2X1_851/m4_208_n4# GND 0.00fF
C65548 PAND2X1_840/m4_208_n4# GND 0.00fF
C65549 PAND2X1_332/Y GND 0.19fF
C65550 PAND2X1_339/m4_208_n4# GND -0.00fF
C65551 POR2X1_314/Y GND 0.16fF
C65552 POR2X1_308/B GND 0.29fF
C65553 POR2X1_386/Y GND -0.00fF
C65554 POR2X1_387/m4_208_n4# GND 0.00fF
C65555 POR2X1_356/B GND 0.24fF
C65556 POR2X1_854/B GND 2.39fF
C65557 POR2X1_319/Y GND -1.17fF
C65558 POR2X1_354/m4_208_n4# GND 0.00fF
C65559 POR2X1_356/Y GND 0.34fF
C65560 POR2X1_365/CTRL2 GND 0.02fF
C65561 POR2X1_321/Y GND 0.20fF
C65562 POR2X1_320/m4_208_n4# GND -0.01fF
C65563 POR2X1_343/B GND 0.09fF
C65564 POR2X1_343/m4_208_n4# GND 0.00fF
C65565 POR2X1_332/m4_208_n4# GND 0.00fF
C65566 POR2X1_310/Y GND 0.33fF
C65567 POR2X1_310/CTRL GND 0.02fF
C65568 PAND2X1_510/B GND -0.74fF
C65569 POR2X1_503/Y GND 0.23fF
C65570 PAND2X1_509/m4_208_n4# GND -0.00fF
C65571 POR2X1_576/Y GND 0.14fF
C65572 POR2X1_579/m4_208_n4# GND 0.00fF
C65573 POR2X1_579/CTRL GND 0.02fF
C65574 POR2X1_568/m4_208_n4# GND 0.00fF
C65575 POR2X1_561/B GND 0.19fF
C65576 POR2X1_558/m4_208_n4# GND -0.01fF
C65577 POR2X1_550/B GND 0.33fF
C65578 POR2X1_513/m4_208_n4# GND 0.00fF
C65579 POR2X1_535/A GND 0.13fF
C65580 POR2X1_788/B GND 0.35fF
C65581 POR2X1_535/m4_208_n4# GND 0.00fF
C65582 POR2X1_731/Y GND 0.14fF
C65583 POR2X1_749/Y GND 0.26fF
C65584 POR2X1_749/m4_208_n4# GND 0.00fF
C65585 POR2X1_731/A GND 0.17fF
C65586 POR2X1_444/Y GND 0.50fF
C65587 POR2X1_353/A GND -1.08fF
C65588 POR2X1_727/CTRL GND 0.01fF
C65589 POR2X1_713/B GND 0.58fF
C65590 POR2X1_705/m4_208_n4# GND 0.00fF
C65591 POR2X1_723/B GND 0.29fF
C65592 POR2X1_303/B GND 0.34fF
C65593 POR2X1_301/m4_208_n4# GND -0.01fF
C65594 POR2X1_689/Y GND 0.20fF
C65595 POR2X1_728/A GND 0.43fF
C65596 PAND2X1_680/m4_208_n4# GND 0.00fF
C65597 POR2X1_90/m4_208_n4# GND 0.00fF
C65598 POR2X1_90/CTRL GND 0.02fF
C65599 PAND2X1_3/B GND -1.03fF
C65600 PAND2X1_18/B GND 0.40fF
C65601 PAND2X1_157/m4_208_n4# GND 0.00fF
C65602 POR2X1_148/A GND 0.21fF
C65603 POR2X1_181/A GND 0.22fF
C65604 PAND2X1_123/Y GND 0.20fF
C65605 PAND2X1_124/m4_208_n4# GND -0.00fF
C65606 PAND2X1_114/B GND 0.08fF
C65607 POR2X1_103/Y GND 0.22fF
C65608 POR2X1_107/Y GND -0.18fF
C65609 POR2X1_702/A GND 0.60fF
C65610 PAND2X1_135/m4_208_n4# GND 0.00fF
C65611 POR2X1_183/m4_208_n4# GND -0.01fF
C65612 POR2X1_200/A GND 0.16fF
C65613 POR2X1_194/m4_208_n4# GND -0.00fF
C65614 POR2X1_194/O GND 0.01fF
C65615 POR2X1_161/m4_208_n4# GND 0.00fF
C65616 POR2X1_150/O GND 0.02fF
C65617 PAND2X1_865/A GND 0.13fF
C65618 PAND2X1_842/Y GND 0.20fF
C65619 PAND2X1_843/Y GND -0.10fF
C65620 PAND2X1_850/CTRL GND 0.02fF
C65621 PAND2X1_359/B GND 0.14fF
C65622 PAND2X1_349/O GND 0.02fF
C65623 PAND2X1_351/A GND 0.26fF
C65624 PAND2X1_333/Y GND 0.19fF
C65625 PAND2X1_305/m4_208_n4# GND -0.00fF
C65626 POR2X1_318/A GND 0.72fF
C65627 PAND2X1_327/CTRL2 GND 0.02fF
C65628 POR2X1_397/m4_208_n4# GND 0.00fF
C65629 POR2X1_397/CTRL2 GND 0.02fF
C65630 POR2X1_22/m4_208_n4# GND -0.01fF
C65631 POR2X1_386/m4_208_n4# GND 0.00fF
C65632 POR2X1_365/A GND 0.19fF
C65633 POR2X1_357/Y GND 0.23fF
C65634 POR2X1_364/CTRL2 GND 0.02fF
C65635 POR2X1_320/Y GND 0.19fF
C65636 POR2X1_39/B GND 1.78fF
C65637 POR2X1_353/m4_208_n4# GND 0.00fF
C65638 POR2X1_594/A GND 0.60fF
C65639 POR2X1_331/m4_208_n4# GND 0.00fF
C65640 POR2X1_342/A GND 0.13fF
C65641 POR2X1_342/B GND 0.26fF
C65642 POR2X1_342/m4_208_n4# GND 0.00fF
C65643 PAND2X1_506/Y GND 0.29fF
C65644 PAND2X1_508/m4_208_n4# GND 0.00fF
C65645 POR2X1_520/A GND 0.29fF
C65646 PAND2X1_492/m4_208_n4# GND -0.01fF
C65647 POR2X1_589/Y GND 0.19fF
C65648 POR2X1_589/m4_208_n4# GND 0.00fF
C65649 POR2X1_551/A GND 0.18fF
C65650 POR2X1_545/m4_208_n4# GND 0.00fF
C65651 POR2X1_577/Y GND -0.16fF
C65652 POR2X1_568/Y GND 2.31fF
C65653 POR2X1_578/m4_208_n4# GND 0.00fF
C65654 POR2X1_631/B GND 0.46fF
C65655 POR2X1_556/m4_208_n4# GND 0.00fF
C65656 POR2X1_568/A GND 0.45fF
C65657 POR2X1_567/m4_208_n4# GND -0.01fF
C65658 POR2X1_513/A GND 0.30fF
C65659 POR2X1_512/m4_208_n4# GND 0.00fF
C65660 POR2X1_512/CTRL GND 0.01fF
C65661 POR2X1_523/B GND 0.28fF
C65662 POR2X1_523/O GND 0.02fF
C65663 POR2X1_534/Y GND 0.14fF
C65664 POR2X1_829/m4_208_n4# GND -0.01fF
C65665 POR2X1_573/A GND 0.48fF
C65666 POR2X1_500/Y GND 0.12fF
C65667 POR2X1_501/B GND 0.19fF
C65668 POR2X1_501/m4_208_n4# GND 0.00fF
C65669 POR2X1_741/A GND 0.11fF
C65670 POR2X1_733/Y GND 0.04fF
C65671 POR2X1_737/m4_208_n4# GND 0.00fF
C65672 POR2X1_748/Y GND 0.18fF
C65673 POR2X1_748/m4_208_n4# GND 0.00fF
C65674 POR2X1_759/Y GND 0.27fF
C65675 POR2X1_711/Y GND -4.38fF
C65676 POR2X1_726/CTRL GND 0.01fF
C65677 POR2X1_317/B GND 0.30fF
C65678 POR2X1_704/m4_208_n4# GND 0.00fF
C65679 POR2X1_724/A GND 0.31fF
C65680 POR2X1_112/Y GND 0.56fF
C65681 POR2X1_691/A GND -0.10fF
C65682 POR2X1_188/Y GND 0.24fF
C65683 PAND2X1_189/m4_208_n4# GND 0.00fF
C65684 POR2X1_158/B GND 0.32fF
C65685 PAND2X1_178/m4_208_n4# GND 0.00fF
C65686 POR2X1_117/Y GND 0.20fF
C65687 POR2X1_117/m4_208_n4# GND -0.01fF
C65688 POR2X1_148/B GND 0.20fF
C65689 PAND2X1_146/m4_208_n4# GND -0.01fF
C65690 POR2X1_768/A GND 0.56fF
C65691 PAND2X1_107/m4_208_n4# GND -0.01fF
C65692 POR2X1_109/Y GND 0.43fF
C65693 PAND2X1_112/m4_208_n4# GND 0.00fF
C65694 PAND2X1_656/A GND 0.50fF
C65695 PAND2X1_99/Y GND 0.17fF
C65696 POR2X1_212/B GND 0.31fF
C65697 POR2X1_181/Y GND 0.03fF
C65698 POR2X1_180/Y GND 0.13fF
C65699 POR2X1_182/CTRL GND 0.02fF
C65700 POR2X1_171/Y GND 0.54fF
C65701 POR2X1_193/O GND 0.02fF
C65702 POR2X1_162/B GND 0.32fF
C65703 POR2X1_356/m4_208_n4# GND -0.01fF
C65704 PAND2X1_861/B GND 0.20fF
C65705 PAND2X1_860/CTRL GND 0.02fF
C65706 PAND2X1_345/Y GND 0.15fF
C65707 PAND2X1_348/Y GND 0.45fF
C65708 PAND2X1_359/O GND 0.02fF
C65709 PAND2X1_324/Y GND 0.16fF
C65710 PAND2X1_326/CTRL GND 0.02fF
C65711 PAND2X1_56/A GND 0.20fF
C65712 PAND2X1_304/CTRL GND 0.02fF
C65713 PAND2X1_352/B GND 0.18fF
C65714 PAND2X1_336/Y GND 0.07fF
C65715 POR2X1_396/m4_208_n4# GND 0.00fF
C65716 POR2X1_396/CTRL GND 0.02fF
C65717 POR2X1_717/B GND 0.46fF
C65718 POR2X1_325/B GND 0.35fF
C65719 POR2X1_374/CTRL2 GND 0.01fF
C65720 POR2X1_385/m4_208_n4# GND -0.01fF
C65721 POR2X1_366/A GND -0.55fF
C65722 POR2X1_359/Y GND -0.22fF
C65723 POR2X1_205/m4_208_n4# GND -0.01fF
C65724 PAND2X1_72/A GND 1.16fF
C65725 PAND2X1_52/B GND -20.32fF
C65726 POR2X1_330/m4_208_n4# GND 0.00fF
C65727 POR2X1_357/B GND 0.21fF
C65728 POR2X1_337/Y GND -1.52fF
C65729 POR2X1_352/m4_208_n4# GND 0.00fF
C65730 POR2X1_228/Y GND 0.83fF
C65731 PAND2X1_508/B GND 0.19fF
C65732 PAND2X1_518/m4_208_n4# GND 0.00fF
C65733 PAND2X1_518/CTRL GND 0.01fF
C65734 POR2X1_587/Y GND 0.15fF
C65735 POR2X1_588/m4_208_n4# GND 0.00fF
C65736 POR2X1_761/A GND 0.35fF
C65737 POR2X1_570/Y GND -0.31fF
C65738 POR2X1_569/Y GND -0.01fF
C65739 POR2X1_562/B GND 0.32fF
C65740 POR2X1_555/CTRL GND 0.02fF
C65741 POR2X1_568/B GND 1.26fF
C65742 POR2X1_566/m4_208_n4# GND 0.00fF
C65743 POR2X1_544/m4_208_n4# GND -0.01fF
C65744 POR2X1_522/CTRL GND 0.02fF
C65745 POR2X1_533/Y GND 0.25fF
C65746 POR2X1_533/O GND 0.02fF
C65747 POR2X1_511/O GND 0.02fF
C65748 POR2X1_844/B GND 0.35fF
C65749 POR2X1_7/Y GND 0.34fF
C65750 POR2X1_758/Y GND 0.19fF
C65751 POR2X1_758/O GND 0.02fF
C65752 POR2X1_747/Y GND 0.33fF
C65753 POR2X1_747/m4_208_n4# GND 0.00fF
C65754 POR2X1_769/B GND 0.02fF
C65755 POR2X1_741/B GND 0.18fF
C65756 POR2X1_675/Y GND 0.48fF
C65757 POR2X1_741/m4_208_n4# GND -0.01fF
C65758 POR2X1_713/Y GND 0.09fF
C65759 POR2X1_712/Y GND 0.06fF
C65760 POR2X1_725/m4_208_n4# GND 0.00fF
C65761 POR2X1_169/A GND 0.38fF
C65762 POR2X1_703/m4_208_n4# GND -0.00fF
C65763 POR2X1_724/B GND 0.19fF
C65764 POR2X1_704/Y GND 0.17fF
C65765 POR2X1_703/Y GND 0.20fF
C65766 POR2X1_714/m4_208_n4# GND 0.00fF
C65767 PAND2X1_207/A GND 0.24fF
C65768 PAND2X1_199/m4_208_n4# GND 0.00fF
C65769 PAND2X1_156/B GND 0.20fF
C65770 POR2X1_153/Y GND 2.30fF
C65771 POR2X1_180/A GND 0.33fF
C65772 POR2X1_498/A GND -0.22fF
C65773 POR2X1_816/A GND 0.28fF
C65774 PAND2X1_133/CTRL2 GND 0.02fF
C65775 PAND2X1_60/B GND 1.65fF
C65776 PAND2X1_144/m4_208_n4# GND -0.01fF
C65777 POR2X1_121/Y GND 0.21fF
C65778 PAND2X1_122/m4_208_n4# GND 0.00fF
C65779 PAND2X1_122/CTRL2 GND 0.02fF
C65780 PAND2X1_101/B GND 0.16fF
C65781 PAND2X1_100/m4_208_n4# GND 0.00fF
C65782 PAND2X1_111/m4_208_n4# GND 0.00fF
C65783 POR2X1_181/m4_208_n4# GND -0.00fF
C65784 POR2X1_191/Y GND 0.79fF
C65785 POR2X1_192/B GND 1.26fF
C65786 POR2X1_580/m4_208_n4# GND -0.01fF
C65787 POR2X1_566/B GND 1.64fF
C65788 POR2X1_169/Y GND 0.14fF
C65789 POR2X1_170/m4_208_n4# GND -0.01fF
C65790 PAND2X1_346/Y GND 0.16fF
C65791 PAND2X1_369/m4_208_n4# GND 0.00fF
C65792 PAND2X1_369/CTRL2 GND 0.02fF
C65793 PAND2X1_364/B GND 0.36fF
C65794 PAND2X1_351/Y GND 0.17fF
C65795 PAND2X1_326/B GND 0.33fF
C65796 PAND2X1_565/m4_208_n4# GND -0.01fF
C65797 POR2X1_317/A GND 0.18fF
C65798 PAND2X1_303/O GND 0.02fF
C65799 POR2X1_77/Y GND 1.52fF
C65800 POR2X1_384/Y GND 0.29fF
C65801 POR2X1_384/m4_208_n4# GND 0.00fF
C65802 POR2X1_395/Y GND -0.11fF
C65803 POR2X1_395/m4_208_n4# GND 0.00fF
C65804 POR2X1_362/m4_208_n4# GND 0.00fF
C65805 POR2X1_339/Y GND 0.25fF
C65806 POR2X1_351/m4_208_n4# GND -0.01fF
C65807 POR2X1_350/B GND 0.22fF
C65808 PAND2X1_88/Y GND -1.29fF
C65809 POR2X1_340/m4_208_n4# GND 0.00fF
C65810 POR2X1_620/B GND 0.15fF
C65811 POR2X1_239/Y GND 0.29fF
C65812 PAND2X1_506/m4_208_n4# GND 0.00fF
C65813 PAND2X1_506/O GND 0.02fF
C65814 PAND2X1_517/m4_208_n4# GND 0.00fF
C65815 POR2X1_294/A GND 1.53fF
C65816 PAND2X1_48/A GND 0.96fF
C65817 POR2X1_598/m4_208_n4# GND -0.01fF
C65818 POR2X1_554/O GND 0.02fF
C65819 POR2X1_572/Y GND 0.19fF
C65820 POR2X1_571/Y GND 0.09fF
C65821 POR2X1_569/A GND 0.73fF
C65822 POR2X1_550/Y GND 0.13fF
C65823 POR2X1_565/m4_208_n4# GND 0.00fF
C65824 POR2X1_532/Y GND 0.22fF
C65825 POR2X1_532/m4_208_n4# GND 0.00fF
C65826 POR2X1_552/A GND -0.35fF
C65827 POR2X1_521/Y GND 0.18fF
C65828 PAND2X1_52/m4_208_n4# GND -0.01fF
C65829 POR2X1_4/Y GND 1.00fF
C65830 POR2X1_6/m4_208_n4# GND 0.00fF
C65831 PAND2X1_711/A GND -0.08fF
C65832 PAND2X1_709/CTRL GND 0.02fF
C65833 POR2X1_783/B GND 0.26fF
C65834 POR2X1_513/B GND 0.86fF
C65835 POR2X1_779/CTRL GND 0.02fF
C65836 POR2X1_746/Y GND 0.21fF
C65837 POR2X1_746/m4_208_n4# GND 0.00fF
C65838 POR2X1_768/m4_208_n4# GND 0.00fF
C65839 POR2X1_757/Y GND 0.20fF
C65840 POR2X1_755/m4_208_n4# GND -0.01fF
C65841 POR2X1_713/m4_208_n4# GND 0.00fF
C65842 POR2X1_732/B GND 0.50fF
C65843 POR2X1_724/m4_208_n4# GND 0.00fF
C65844 POR2X1_736/A GND 1.07fF
C65845 POR2X1_632/Y GND 0.45fF
C65846 POR2X1_735/m4_208_n4# GND 0.00fF
C65847 POR2X1_715/A GND 0.35fF
C65848 POR2X1_702/m4_208_n4# GND 0.00fF
C65849 POR2X1_57/Y GND 0.16fF
C65850 PAND2X1_197/Y GND 0.27fF
C65851 PAND2X1_198/CTRL2 GND 0.02fF
C65852 POR2X1_191/B GND 0.12fF
C65853 PAND2X1_176/m4_208_n4# GND 0.00fF
C65854 PAND2X1_176/CTRL2 GND 0.02fF
C65855 PAND2X1_165/m4_208_n4# GND 0.00fF
C65856 PAND2X1_156/A GND 0.48fF
C65857 PAND2X1_154/CTRL GND 0.02fF
C65858 PAND2X1_8/Y GND 0.64fF
C65859 PAND2X1_143/CTRL2 GND 0.02fF
C65860 PAND2X1_121/m4_208_n4# GND 0.00fF
C65861 PAND2X1_111/B GND 0.03fF
C65862 PAND2X1_110/m4_208_n4# GND 0.00fF
C65863 PAND2X1_110/CTRL2 GND 0.02fF
C65864 POR2X1_190/Y GND 0.25fF
C65865 POR2X1_191/m4_208_n4# GND -0.01fF
C65866 POR2X1_180/CTRL GND 0.02fF
C65867 PAND2X1_379/m4_208_n4# GND 0.00fF
C65868 PAND2X1_352/Y GND -0.43fF
C65869 PAND2X1_353/Y GND 0.20fF
C65870 PAND2X1_357/CTRL GND 0.02fF
C65871 PAND2X1_368/m4_208_n4# GND 0.00fF
C65872 PAND2X1_337/A GND -0.27fF
C65873 POR2X1_309/Y GND 0.33fF
C65874 PAND2X1_335/O GND 0.02fF
C65875 POR2X1_295/Y GND 0.83fF
C65876 POR2X1_481/m4_208_n4# GND -0.01fF
C65877 PAND2X1_313/m4_208_n4# GND 0.00fF
C65878 PAND2X1_303/B GND 0.20fF
C65879 PAND2X1_302/CTRL2 GND 0.02fF
C65880 POR2X1_372/Y GND 0.67fF
C65881 POR2X1_372/m4_208_n4# GND -0.00fF
C65882 POR2X1_383/Y GND 0.30fF
C65883 POR2X1_383/m4_208_n4# GND -0.01fF
C65884 POR2X1_394/CTRL GND 0.02fF
C65885 POR2X1_362/A GND 0.33fF
C65886 POR2X1_276/Y GND 0.54fF
C65887 POR2X1_361/m4_208_n4# GND 0.00fF
C65888 POR2X1_361/CTRL GND 0.01fF
C65889 POR2X1_341/Y GND -0.17fF
C65890 POR2X1_502/m4_208_n4# GND -0.01fF
C65891 PAND2X1_565/A GND 0.38fF
C65892 POR2X1_531/Y GND 0.20fF
C65893 PAND2X1_549/CTRL GND 0.02fF
C65894 PAND2X1_539/B GND 0.20fF
C65895 PAND2X1_802/m4_208_n4# GND -0.01fF
C65896 POR2X1_507/A GND 0.84fF
C65897 PAND2X1_505/m4_208_n4# GND 0.00fF
C65898 PAND2X1_505/CTRL2 GND 0.02fF
C65899 POR2X1_513/Y GND 0.20fF
C65900 POR2X1_515/Y GND 0.17fF
C65901 POR2X1_547/B GND 0.46fF
C65902 PAND2X1_527/m4_208_n4# GND 0.00fF
C65903 POR2X1_597/CTRL GND 0.02fF
C65904 POR2X1_586/m4_208_n4# GND -0.00fF
C65905 POR2X1_552/Y GND 0.13fF
C65906 POR2X1_564/CTRL GND 0.02fF
C65907 POR2X1_579/B GND 0.29fF
C65908 POR2X1_574/Y GND 0.33fF
C65909 POR2X1_575/m4_208_n4# GND 0.00fF
C65910 POR2X1_73/Y GND 1.85fF
C65911 POR2X1_531/CTRL GND 0.02fF
C65912 POR2X1_542/m4_208_n4# GND 0.00fF
C65913 POR2X1_540/Y GND -3.37fF
C65914 POR2X1_553/m4_208_n4# GND 0.00fF
C65915 POR2X1_559/A GND 0.69fF
C65916 POR2X1_520/B GND 0.29fF
C65917 POR2X1_520/m4_208_n4# GND 0.00fF
C65918 POR2X1_520/CTRL GND 0.01fF
C65919 POR2X1_5/m4_208_n4# GND 0.00fF
C65920 POR2X1_665/Y GND 0.07fF
C65921 PAND2X1_719/m4_208_n4# GND 0.00fF
C65922 PAND2X1_712/B GND 0.30fF
C65923 PAND2X1_708/CTRL GND 0.02fF
C65924 POR2X1_789/B GND 0.15fF
C65925 POR2X1_789/m4_208_n4# GND 0.00fF
C65926 POR2X1_784/A GND 0.30fF
C65927 POR2X1_778/m4_208_n4# GND 0.00fF
C65928 POR2X1_778/CTRL2 GND 0.02fF
C65929 POR2X1_767/Y GND 0.23fF
C65930 POR2X1_767/m4_208_n4# GND 0.00fF
C65931 POR2X1_737/A GND 0.31fF
C65932 POR2X1_734/m4_208_n4# GND 0.00fF
C65933 POR2X1_707/Y GND 0.21fF
C65934 POR2X1_745/Y GND 0.24fF
C65935 POR2X1_733/A GND 0.67fF
C65936 POR2X1_717/Y GND 0.18fF
C65937 POR2X1_723/m4_208_n4# GND -0.01fF
C65938 POR2X1_701/Y GND 0.15fF
C65939 POR2X1_236/Y GND 2.58fF
C65940 POR2X1_701/m4_208_n4# GND -0.00fF
C65941 POR2X1_701/CTRL GND 0.02fF
C65942 PAND2X1_853/B GND -1.58fF
C65943 POR2X1_52/Y GND 0.24fF
C65944 POR2X1_56/Y GND 0.36fF
C65945 POR2X1_776/B GND 0.60fF
C65946 PAND2X1_164/m4_208_n4# GND 0.00fF
C65947 POR2X1_830/A GND 0.60fF
C65948 PAND2X1_142/O GND 0.02fF
C65949 PAND2X1_153/CTRL GND 0.02fF
C65950 POR2X1_140/A GND 0.16fF
C65951 POR2X1_130/Y GND 0.12fF
C65952 POR2X1_666/A GND 0.42fF
C65953 PAND2X1_120/m4_208_n4# GND 0.00fF
C65954 POR2X1_456/B GND 0.55fF
C65955 POR2X1_190/m4_208_n4# GND 0.00fF
C65956 POR2X1_387/Y GND 0.62fF
C65957 PAND2X1_389/m4_208_n4# GND 0.00fF
C65958 POR2X1_459/A GND 0.26fF
C65959 POR2X1_42/Y GND -19.68fF
C65960 PAND2X1_377/Y GND 0.16fF
C65961 PAND2X1_378/m4_208_n4# GND 0.00fF
C65962 GATE_366 GND 0.17fF
C65963 PAND2X1_366/Y GND 0.14fF
C65964 PAND2X1_365/A GND 0.20fF
C65965 PAND2X1_354/Y GND 0.25fF
C65966 PAND2X1_356/O GND 0.02fF
C65967 PAND2X1_338/B GND -0.45fF
C65968 POR2X1_291/Y GND 0.08fF
C65969 PAND2X1_334/m4_208_n4# GND 0.00fF
C65970 PAND2X1_555/A GND 0.28fF
C65971 PAND2X1_345/m4_208_n4# GND 0.00fF
C65972 POR2X1_325/A GND 0.35fF
C65973 PAND2X1_323/m4_208_n4# GND 0.00fF
C65974 PAND2X1_323/O GND 0.01fF
C65975 PAND2X1_716/B GND 0.36fF
C65976 POR2X1_75/Y GND 0.34fF
C65977 POR2X1_300/Y GND -0.20fF
C65978 PAND2X1_301/CTRL2 GND 0.02fF
C65979 POR2X1_703/A GND 0.85fF
C65980 POR2X1_382/Y GND 0.43fF
C65981 POR2X1_382/CTRL GND 0.02fF
C65982 POR2X1_372/A GND 0.28fF
C65983 POR2X1_5/Y GND 1.65fF
C65984 POR2X1_371/m4_208_n4# GND 0.00fF
C65985 POR2X1_363/A GND 0.08fF
C65986 POR2X1_244/Y GND -1.03fF
C65987 POR2X1_360/CTRL2 GND 0.02fF
C65988 PAND2X1_560/B GND 0.53fF
C65989 PAND2X1_559/m4_208_n4# GND 0.00fF
C65990 PAND2X1_549/B GND 0.35fF
C65991 POR2X1_530/Y GND 0.21fF
C65992 PAND2X1_548/m4_208_n4# GND 0.00fF
C65993 PAND2X1_514/Y GND 0.08fF
C65994 PAND2X1_515/m4_208_n4# GND 0.00fF
C65995 POR2X1_546/A GND 0.44fF
C65996 PAND2X1_643/A GND 0.41fF
C65997 POR2X1_385/Y GND 0.54fF
C65998 PAND2X1_537/CTRL GND 0.02fF
C65999 PAND2X1_504/CTRL GND 0.02fF
C66000 POR2X1_293/Y GND -12.05fF
C66001 POR2X1_585/m4_208_n4# GND 0.00fF
C66002 POR2X1_574/A GND 0.04fF
C66003 POR2X1_510/Y GND 0.67fF
C66004 POR2X1_574/m4_208_n4# GND 0.00fF
C66005 POR2X1_554/Y GND 0.21fF
C66006 POR2X1_553/Y GND 0.07fF
C66007 POR2X1_563/m4_208_n4# GND 0.00fF
C66008 POR2X1_542/Y GND 0.17fF
C66009 POR2X1_552/m4_208_n4# GND 0.00fF
C66010 POR2X1_530/m4_208_n4# GND 0.00fF
C66011 POR2X1_553/A GND -0.29fF
C66012 POR2X1_274/B GND 0.46fF
C66013 POR2X1_541/m4_208_n4# GND 0.00fF
C66014 POR2X1_4/m4_208_n4# GND 0.00fF
C66015 POR2X1_4/CTRL GND 0.02fF
C66016 POR2X1_591/Y GND 0.49fF
C66017 PAND2X1_645/B GND 0.26fF
C66018 PAND2X1_730/B GND 0.39fF
C66019 PAND2X1_687/Y GND 0.41fF
C66020 PAND2X1_729/m4_208_n4# GND -0.00fF
C66021 POR2X1_802/A GND 0.46fF
C66022 POR2X1_652/A GND 0.50fF
C66023 POR2X1_593/m4_208_n4# GND -0.01fF
C66024 POR2X1_307/A GND -0.23fF
C66025 POR2X1_777/m4_208_n4# GND 0.00fF
C66026 POR2X1_788/CTRL2 GND 0.02fF
C66027 POR2X1_766/Y GND 0.13fF
C66028 POR2X1_766/m4_208_n4# GND 0.00fF
C66029 POR2X1_755/Y GND 0.14fF
C66030 POR2X1_665/A GND -0.05fF
C66031 POR2X1_722/Y GND 0.36fF
C66032 POR2X1_744/O GND 0.02fF
C66033 POR2X1_710/Y GND 0.16fF
C66034 POR2X1_711/m4_208_n4# GND 0.00fF
C66035 POR2X1_700/Y GND -0.13fF
C66036 POR2X1_90/Y GND 1.01fF
C66037 POR2X1_700/m4_208_n4# GND 0.00fF
C66038 PAND2X1_199/B GND 0.30fF
C66039 PAND2X1_196/CTRL2 GND 0.02fF
C66040 PAND2X1_175/B GND 0.32fF
C66041 POR2X1_172/Y GND 0.15fF
C66042 PAND2X1_185/CTRL GND 0.02fF
C66043 POR2X1_210/A GND 0.16fF
C66044 POR2X1_209/A GND 0.48fF
C66045 PAND2X1_139/Y GND 0.20fF
C66046 PAND2X1_140/Y GND 0.12fF
C66047 POR2X1_131/A GND 0.25fF
C66048 POR2X1_129/Y GND 0.67fF
C66049 POR2X1_398/Y GND -0.02fF
C66050 PAND2X1_399/CTRL2 GND 0.02fF
C66051 POR2X1_176/Y GND 0.35fF
C66052 PAND2X1_439/m4_208_n4# GND -0.01fF
C66053 PAND2X1_376/m4_208_n4# GND -0.00fF
C66054 PAND2X1_363/Y GND 0.45fF
C66055 PAND2X1_348/A GND -3.05fF
C66056 PAND2X1_322/CTRL2 GND 0.01fF
C66057 PAND2X1_333/O GND 0.02fF
C66058 PAND2X1_356/B GND 0.14fF
C66059 POR2X1_331/Y GND 0.14fF
C66060 PAND2X1_355/O GND 0.02fF
C66061 PAND2X1_300/m4_208_n4# GND 0.00fF
C66062 PAND2X1_311/m4_208_n4# GND 0.00fF
C66063 PAND2X1_311/CTRL2 GND 0.02fF
C66064 POR2X1_391/Y GND 0.40fF
C66065 POR2X1_392/CTRL GND 0.02fF
C66066 POR2X1_817/A GND 0.09fF
C66067 POR2X1_381/CTRL GND 0.02fF
C66068 POR2X1_543/A GND -0.32fF
C66069 POR2X1_370/m4_208_n4# GND 0.00fF
C66070 PAND2X1_770/m4_208_n4# GND -0.01fF
C66071 PAND2X1_550/B GND 0.29fF
C66072 POR2X1_527/Y GND -0.07fF
C66073 PAND2X1_493/Y GND 0.27fF
C66074 POR2X1_494/Y GND 0.31fF
C66075 POR2X1_537/A GND 0.21fF
C66076 PAND2X1_536/m4_208_n4# GND 0.00fF
C66077 POR2X1_546/B GND 0.17fF
C66078 POR2X1_546/m4_208_n4# GND -0.01fF
C66079 POR2X1_502/Y GND 0.29fF
C66080 POR2X1_584/Y GND 0.00fF
C66081 POR2X1_7/A GND -7.67fF
C66082 POR2X1_575/B GND 0.20fF
C66083 POR2X1_404/Y GND 0.39fF
C66084 POR2X1_573/m4_208_n4# GND 0.00fF
C66085 POR2X1_595/Y GND 0.34fF
C66086 POR2X1_250/A GND 0.55fF
C66087 POR2X1_564/B GND 0.16fF
C66088 POR2X1_544/Y GND 0.13fF
C66089 POR2X1_551/CTRL GND 0.02fF
C66090 POR2X1_181/B GND 0.19fF
C66091 POR2X1_540/m4_208_n4# GND 0.00fF
C66092 POR2X1_570/B GND 0.21fF
C66093 POR2X1_556/Y GND -0.09fF
C66094 POR2X1_562/m4_208_n4# GND 0.00fF
C66095 PAND2X1_739/CTRL GND 0.02fF
C66096 PAND2X1_713/B GND 0.31fF
C66097 POR2X1_692/Y GND 0.20fF
C66098 PAND2X1_706/m4_208_n4# GND 0.00fF
C66099 PAND2X1_730/A GND 0.49fF
C66100 PAND2X1_728/O GND 0.02fF
C66101 PAND2X1_717/CTRL2 GND 0.02fF
C66102 POR2X1_802/B GND 0.52fF
C66103 POR2X1_468/B GND -0.04fF
C66104 POR2X1_798/m4_208_n4# GND 0.00fF
C66105 POR2X1_794/B GND 0.47fF
C66106 POR2X1_787/m4_208_n4# GND 0.00fF
C66107 POR2X1_765/Y GND 0.26fF
C66108 POR2X1_765/m4_208_n4# GND -0.01fF
C66109 POR2X1_785/A GND 0.32fF
C66110 POR2X1_776/CTRL GND 0.02fF
C66111 POR2X1_754/m4_208_n4# GND 0.00fF
C66112 POR2X1_738/A GND 0.23fF
C66113 POR2X1_725/Y GND -3.84fF
C66114 POR2X1_732/m4_208_n4# GND 0.00fF
C66115 POR2X1_743/Y GND 0.23fF
C66116 POR2X1_7/B GND 1.07fF
C66117 POR2X1_734/A GND -7.09fF
C66118 POR2X1_720/Y GND 0.13fF
C66119 POR2X1_721/m4_208_n4# GND 0.00fF
C66120 POR2X1_710/B GND 0.16fF
C66121 POR2X1_213/B GND 0.17fF
C66122 POR2X1_209/m4_208_n4# GND 0.00fF
C66123 PAND2X1_199/A GND 0.08fF
C66124 PAND2X1_195/CTRL GND 0.02fF
C66125 PAND2X1_71/Y GND -0.04fF
C66126 PAND2X1_184/m4_208_n4# GND 0.00fF
C66127 POR2X1_175/B GND 0.14fF
C66128 PAND2X1_173/m4_208_n4# GND 0.00fF
C66129 PAND2X1_161/Y GND -0.20fF
C66130 PAND2X1_162/m4_208_n4# GND 0.00fF
C66131 POR2X1_152/A GND -0.23fF
C66132 POR2X1_55/Y GND 2.20fF
C66133 PAND2X1_151/m4_208_n4# GND 0.00fF
C66134 PAND2X1_140/m4_208_n4# GND 0.00fF
C66135 PAND2X1_398/m4_208_n4# GND 0.00fF
C66136 PAND2X1_386/Y GND -0.04fF
C66137 PAND2X1_387/m4_208_n4# GND 0.00fF
C66138 POR2X1_375/Y GND -0.15fF
C66139 PAND2X1_367/A GND 0.20fF
C66140 PAND2X1_349/B GND 0.19fF
C66141 PAND2X1_343/m4_208_n4# GND 0.00fF
C66142 PAND2X1_854/A GND 0.71fF
C66143 POR2X1_294/B GND 2.32fF
C66144 PAND2X1_321/m4_208_n4# GND 0.00fF
C66145 PAND2X1_310/CTRL GND 0.02fF
C66146 POR2X1_391/B GND 0.21fF
C66147 POR2X1_391/CTRL GND 0.02fF
C66148 POR2X1_380/Y GND -0.23fF
C66149 POR2X1_380/A GND 0.13fF
C66150 POR2X1_380/m4_208_n4# GND 0.00fF
C66151 PAND2X1_578/A GND 0.18fF
C66152 PAND2X1_566/Y GND 1.02fF
C66153 PAND2X1_347/m4_208_n4# GND -0.01fF
C66154 PAND2X1_580/B GND 0.45fF
C66155 PAND2X1_579/m4_208_n4# GND 0.00fF
C66156 PAND2X1_561/A GND 0.23fF
C66157 PAND2X1_473/m4_208_n4# GND -0.01fF
C66158 PAND2X1_855/m4_208_n4# GND -0.01fF
C66159 POR2X1_526/Y GND 0.23fF
C66160 PAND2X1_546/m4_208_n4# GND 0.00fF
C66161 POR2X1_545/A GND 0.29fF
C66162 PAND2X1_524/m4_208_n4# GND 0.00fF
C66163 POR2X1_516/B GND 0.16fF
C66164 PAND2X1_512/Y GND 0.28fF
C66165 POR2X1_503/A GND 0.21fF
C66166 PAND2X1_502/O GND 0.02fF
C66167 POR2X1_583/Y GND 0.03fF
C66168 POR2X1_583/m4_208_n4# GND 0.00fF
C66169 POR2X1_267/Y GND -0.20fF
C66170 POR2X1_572/CTRL GND 0.02fF
C66171 POR2X1_558/Y GND 0.25fF
C66172 POR2X1_550/m4_208_n4# GND 0.00fF
C66173 INPUT_5 GND 0.44fF
C66174 INPUT_4 GND 0.62fF
C66175 POR2X1_2/m4_208_n4# GND 0.00fF
C66176 POR2X1_750/A GND 0.30fF
C66177 PAND2X1_749/m4_208_n4# GND 0.00fF
C66178 PAND2X1_749/CTRL2 GND 0.02fF
C66179 PAND2X1_713/A GND 0.16fF
C66180 PAND2X1_705/m4_208_n4# GND 0.00fF
C66181 PAND2X1_738/CTRL GND 0.02fF
C66182 PAND2X1_731/B GND -0.84fF
C66183 PAND2X1_444/Y GND 0.42fF
C66184 PAND2X1_727/CTRL2 GND 0.02fF
C66185 PAND2X1_723/A GND 0.68fF
C66186 POR2X1_803/A GND 0.28fF
C66187 POR2X1_149/Y GND -0.24fF
C66188 POR2X1_797/O GND 0.02fF
C66189 POR2X1_764/Y GND 0.20fF
C66190 POR2X1_40/Y GND 1.68fF
C66191 POR2X1_785/B GND 0.26fF
C66192 POR2X1_785/m4_208_n4# GND -0.01fF
C66193 POR2X1_786/m4_208_n4# GND 0.00fF
C66194 POR2X1_752/Y GND -0.69fF
C66195 POR2X1_726/Y GND 0.13fF
C66196 POR2X1_731/CTRL GND 0.01fF
C66197 D_GATE_741 GND 0.43fF
C66198 POR2X1_741/Y GND 1.71fF
C66199 POR2X1_740/Y GND 2.36fF
C66200 POR2X1_742/m4_208_n4# GND 0.00fF
C66201 POR2X1_720/A GND 0.16fF
C66202 POR2X1_720/m4_208_n4# GND 0.00fF
C66203 POR2X1_222/A GND 0.46fF
C66204 POR2X1_215/Y GND 0.14fF
C66205 POR2X1_219/O GND 0.02fF
C66206 POR2X1_35/Y GND 0.35fF
C66207 PAND2X1_200/B GND 0.30fF
C66208 POR2X1_16/Y GND 0.16fF
C66209 POR2X1_39/Y GND 0.22fF
C66210 PAND2X1_194/m4_208_n4# GND -0.00fF
C66211 POR2X1_540/A GND -0.78fF
C66212 PAND2X1_161/m4_208_n4# GND 0.00fF
C66213 POR2X1_174/A GND 0.51fF
C66214 PAND2X1_63/B GND 0.39fF
C66215 PAND2X1_150/m4_208_n4# GND 0.00fF
C66216 POR2X1_398/m4_208_n4# GND -0.01fF
C66217 POR2X1_376/A GND 0.10fF
C66218 PAND2X1_386/m4_208_n4# GND 0.00fF
C66219 POR2X1_355/A GND -0.26fF
C66220 POR2X1_330/Y GND 2.49fF
C66221 PAND2X1_331/m4_208_n4# GND 0.00fF
C66222 PAND2X1_303/Y GND 0.19fF
C66223 PAND2X1_308/Y GND 0.29fF
C66224 PAND2X1_353/CTRL GND 0.02fF
C66225 PAND2X1_349/A GND 0.34fF
C66226 POR2X1_248/Y GND 0.16fF
C66227 PAND2X1_342/CTRL GND 0.02fF
C66228 PAND2X1_365/B GND 0.22fF
C66229 PAND2X1_357/Y GND 0.53fF
C66230 PAND2X1_364/m4_208_n4# GND 0.00fF
C66231 PAND2X1_320/m4_208_n4# GND 0.00fF
C66232 POR2X1_392/B GND 0.51fF
C66233 POR2X1_389/Y GND 0.35fF
C66234 POR2X1_390/m4_208_n4# GND -0.00fF
C66235 POR2X1_390/O GND 0.02fF
C66236 PAND2X1_589/m4_208_n4# GND 0.00fF
C66237 PAND2X1_562/B GND 0.62fF
C66238 PAND2X1_577/Y GND 0.39fF
C66239 PAND2X1_287/m4_208_n4# GND -0.01fF
C66240 PAND2X1_568/B GND 0.45fF
C66241 POR2X1_524/Y GND 0.31fF
C66242 POR2X1_296/B GND 1.94fF
C66243 PAND2X1_534/m4_208_n4# GND 0.00fF
C66244 PAND2X1_844/B GND 0.42fF
C66245 POR2X1_522/Y GND -0.19fF
C66246 PAND2X1_523/CTRL GND 0.02fF
C66247 INPUT_0 GND 2.78fF
C66248 PAND2X1_512/m4_208_n4# GND 0.00fF
C66249 PAND2X1_573/B GND -0.51fF
C66250 POR2X1_498/Y GND 0.17fF
C66251 POR2X1_592/Y GND 0.09fF
C66252 POR2X1_559/Y GND 0.23fF
C66253 POR2X1_523/Y GND 0.31fF
C66254 POR2X1_561/Y GND -0.20fF
C66255 POR2X1_560/Y GND 0.13fF
C66256 POR2X1_571/m4_208_n4# GND 0.00fF
C66257 POR2X1_3/B GND 0.46fF
C66258 POR2X1_792/B GND 0.21fF
C66259 PAND2X1_731/A GND 0.24fF
C66260 POR2X1_152/Y GND 0.30fF
C66261 PAND2X1_724/B GND 0.33fF
C66262 PAND2X1_115/B GND 0.23fF
C66263 PAND2X1_715/m4_208_n4# GND 0.00fF
C66264 PAND2X1_741/B GND 0.41fF
C66265 PAND2X1_733/Y GND -0.24fF
C66266 PAND2X1_737/CTRL2 GND 0.02fF
C66267 PAND2X1_714/B GND -0.16fF
C66268 POR2X1_774/m4_208_n4# GND 0.00fF
C66269 POR2X1_774/CTRL GND 0.02fF
C66270 POR2X1_783/Y GND 0.13fF
C66271 POR2X1_795/B GND 0.45fF
C66272 POR2X1_729/Y GND 0.19fF
C66273 POR2X1_730/m4_208_n4# GND 0.00fF
C66274 POR2X1_763/Y GND 1.20fF
C66275 POR2X1_46/Y GND 1.74fF
C66276 POR2X1_216/Y GND 0.13fF
C66277 POR2X1_218/m4_208_n4# GND 0.00fF
C66278 POR2X1_218/CTRL GND 0.01fF
C66279 POR2X1_229/Y GND -0.18fF
C66280 POR2X1_229/m4_208_n4# GND -0.01fF
C66281 POR2X1_214/B GND 0.22fF
C66282 POR2X1_207/O GND 0.02fF
C66283 PAND2X1_182/O GND 0.02fF
C66284 PAND2X1_193/CTRL2 GND 0.02fF
C66285 PAND2X1_162/A GND 0.32fF
C66286 POR2X1_394/A GND 3.17fF
C66287 PAND2X1_160/m4_208_n4# GND 0.00fF
C66288 PAND2X1_160/CTRL GND 0.02fF
C66289 PAND2X1_396/m4_208_n4# GND 0.00fF
C66290 POR2X1_373/Y GND 0.28fF
C66291 PAND2X1_374/CTRL GND 0.02fF
C66292 POR2X1_537/B GND 0.36fF
C66293 PAND2X1_352/O GND 0.02fF
C66294 PAND2X1_359/Y GND -0.32fF
C66295 PAND2X1_360/Y GND 0.10fF
C66296 PAND2X1_363/O GND 0.02fF
C66297 PAND2X1_341/m4_208_n4# GND 0.00fF
C66298 POR2X1_331/A GND -0.26fF
C66299 PAND2X1_330/m4_208_n4# GND 0.00fF
C66300 POR2X1_644/A GND 0.25fF
C66301 PAND2X1_69/A GND 1.65fF
C66302 POR2X1_828/A GND 0.53fF
C66303 PAND2X1_587/Y GND 0.13fF
C66304 PAND2X1_588/m4_208_n4# GND 0.00fF
C66305 PAND2X1_211/A GND 0.49fF
C66306 PAND2X1_566/O GND 0.02fF
C66307 PAND2X1_569/Y GND 0.18fF
C66308 PAND2X1_551/A GND 0.24fF
C66309 PAND2X1_544/CTRL2 GND 0.02fF
C66310 PAND2X1_555/m4_208_n4# GND 0.00fF
C66311 PAND2X1_501/B GND 0.25fF
C66312 POR2X1_497/Y GND -1.13fF
C66313 PAND2X1_499/Y GND -3.31fF
C66314 POR2X1_523/A GND 0.16fF
C66315 PAND2X1_522/O GND 0.02fF
C66316 POR2X1_592/A GND 0.13fF
C66317 POR2X1_582/A GND 0.14fF
C66318 D_INPUT_6 GND 0.16fF
C66319 POR2X1_581/m4_208_n4# GND 0.00fF
C66320 POR2X1_581/CTRL GND 0.01fF
C66321 POR2X1_563/Y GND 0.13fF
C66322 POR2X1_570/m4_208_n4# GND 0.00fF
C66323 POR2X1_759/A GND 0.19fF
C66324 PAND2X1_758/m4_208_n4# GND 0.00fF
C66325 POR2X1_782/B GND 0.16fF
C66326 PAND2X1_747/CTRL GND 0.02fF
C66327 PAND2X1_735/Y GND 0.64fF
C66328 PAND2X1_714/A GND 0.19fF
C66329 POR2X1_312/Y GND 0.32fF
C66330 PAND2X1_317/m4_208_n4# GND -0.01fF
C66331 POR2X1_774/A GND 0.29fF
C66332 POR2X1_773/m4_208_n4# GND 0.00fF
C66333 POR2X1_796/A GND 0.28fF
C66334 POR2X1_777/Y GND -0.27fF
C66335 POR2X1_784/m4_208_n4# GND 0.00fF
C66336 POR2X1_804/A GND 1.75fF
C66337 POR2X1_786/Y GND -2.78fF
C66338 POR2X1_795/m4_208_n4# GND 0.00fF
C66339 POR2X1_738/Y GND 0.13fF
C66340 POR2X1_740/m4_208_n4# GND 0.00fF
C66341 POR2X1_763/A GND 0.62fF
C66342 POR2X1_751/Y GND 0.27fF
C66343 POR2X1_239/m4_208_n4# GND 0.00fF
C66344 POR2X1_218/A GND 0.46fF
C66345 POR2X1_572/B GND 0.24fF
C66346 PAND2X1_52/Y GND 0.29fF
C66347 PAND2X1_7/Y GND -0.22fF
C66348 POR2X1_228/m4_208_n4# GND 0.00fF
C66349 POR2X1_215/A GND 0.27fF
C66350 POR2X1_201/Y GND 0.21fF
C66351 POR2X1_408/Y GND -16.98fF
C66352 POR2X1_409/CTRL GND 0.02fF
C66353 PAND2X1_191/Y GND -0.28fF
C66354 PAND2X1_192/CTRL GND 0.02fF
C66355 PAND2X1_168/Y GND 0.21fF
C66356 PAND2X1_169/Y GND -0.45fF
C66357 PAND2X1_170/CTRL GND 0.02fF
C66358 PAND2X1_182/B GND -0.21fF
C66359 POR2X1_401/B GND 0.35fF
C66360 PAND2X1_395/m4_208_n4# GND 0.00fF
C66361 PAND2X1_395/CTRL2 GND 0.02fF
C66362 POR2X1_391/A GND 0.27fF
C66363 POR2X1_544/B GND 0.41fF
C66364 PAND2X1_366/A GND 0.19fF
C66365 PAND2X1_806/m4_208_n4# GND -0.01fF
C66366 PAND2X1_339/Y GND 0.09fF
C66367 PAND2X1_350/A GND 0.21fF
C66368 POR2X1_88/Y GND 0.16fF
C66369 PAND2X1_587/m4_208_n4# GND 0.00fF
C66370 POR2X1_599/A GND -5.98fF
C66371 PAND2X1_598/CTRL GND 0.02fF
C66372 PAND2X1_579/B GND 0.33fF
C66373 PAND2X1_571/Y GND 0.13fF
C66374 POR2X1_533/A GND 0.32fF
C66375 PAND2X1_791/m4_208_n4# GND -0.01fF
C66376 PAND2X1_569/B GND 1.44fF
C66377 PAND2X1_550/Y GND 0.14fF
C66378 PAND2X1_552/B GND 0.23fF
C66379 PAND2X1_563/B GND 0.20fF
C66380 POR2X1_106/Y GND 0.50fF
C66381 PAND2X1_657/B GND 0.32fF
C66382 PAND2X1_508/Y GND 0.58fF
C66383 PAND2X1_510/CTRL GND 0.02fF
C66384 PAND2X1_521/m4_208_n4# GND 0.00fF
C66385 POR2X1_591/O GND 0.02fF
C66386 D_GATE_579 GND 0.26fF
C66387 POR2X1_579/Y GND 0.09fF
C66388 POR2X1_578/Y GND 0.55fF
C66389 POR2X1_511/Y GND 0.20fF
C66390 PAND2X1_779/m4_208_n4# GND 0.00fF
C66391 POR2X1_756/Y GND 0.16fF
C66392 PAND2X1_757/CTRL GND 0.02fF
C66393 PAND2X1_768/CTRL GND 0.02fF
C66394 POR2X1_781/A GND 0.22fF
C66395 PAND2X1_746/CTRL GND 0.02fF
C66396 PAND2X1_732/A GND -0.07fF
C66397 PAND2X1_714/Y GND -0.51fF
C66398 PAND2X1_724/CTRL GND 0.02fF
C66399 PAND2X1_658/B GND 0.33fF
C66400 PAND2X1_735/O GND 0.02fF
C66401 PAND2X1_725/B GND 0.24fF
C66402 PAND2X1_713/m4_208_n4# GND 0.00fF
C66403 PAND2X1_715/B GND 0.30fF
C66404 PAND2X1_702/O GND 0.02fF
C66405 POR2X1_804/B GND 0.21fF
C66406 POR2X1_788/Y GND 0.32fF
C66407 POR2X1_783/m4_208_n4# GND -0.00fF
C66408 POR2X1_773/A GND 0.33fF
C66409 POR2X1_768/Y GND 0.14fF
C66410 POR2X1_557/B GND 0.33fF
C66411 POR2X1_772/m4_208_n4# GND 0.00fF
C66412 POR2X1_750/Y GND -2.06fF
C66413 POR2X1_750/m4_208_n4# GND -0.00fF
C66414 POR2X1_761/Y GND 0.28fF
C66415 POR2X1_761/m4_208_n4# GND 0.00fF
C66416 POR2X1_249/Y GND 0.35fF
C66417 POR2X1_249/m4_208_n4# GND 0.00fF
C66418 POR2X1_238/Y GND -0.65fF
C66419 POR2X1_238/CTRL GND 0.02fF
C66420 POR2X1_509/B GND 0.34fF
C66421 POR2X1_227/m4_208_n4# GND -0.01fF
C66422 POR2X1_116/Y GND -0.27fF
C66423 POR2X1_101/Y GND 1.19fF
C66424 POR2X1_216/m4_208_n4# GND 0.00fF
C66425 POR2X1_216/CTRL GND 0.01fF
C66426 POR2X1_203/Y GND 0.21fF
C66427 POR2X1_419/Y GND 0.26fF
C66428 POR2X1_419/O GND 0.02fF
C66429 POR2X1_408/m4_208_n4# GND -0.00fF
C66430 PAND2X1_190/Y GND 0.36fF
C66431 PAND2X1_182/A GND 0.02fF
C66432 PAND2X1_180/m4_208_n4# GND 0.00fF
C66433 PAND2X1_394/m4_208_n4# GND 0.00fF
C66434 POR2X1_384/A GND 0.50fF
C66435 PAND2X1_383/m4_208_n4# GND 0.00fF
C66436 POR2X1_458/B GND 0.21fF
C66437 D_INPUT_1 GND 1.39fF
C66438 POR2X1_778/B GND 0.25fF
C66439 PAND2X1_372/m4_208_n4# GND -0.00fF
C66440 PAND2X1_362/B GND 0.27fF
C66441 PAND2X1_473/B GND -1.04fF
C66442 PAND2X1_358/A GND 0.59fF
C66443 PAND2X1_341/Y GND -0.22fF
C66444 PAND2X1_350/m4_208_n4# GND 0.00fF
C66445 POR2X1_596/Y GND 0.16fF
C66446 PAND2X1_597/O GND 0.02fF
C66447 POR2X1_637/A GND 0.16fF
C66448 PAND2X1_586/m4_208_n4# GND 0.00fF
C66449 PAND2X1_579/A GND 0.16fF
C66450 PAND2X1_575/m4_208_n4# GND 0.00fF
C66451 PAND2X1_569/A GND 0.19fF
C66452 PAND2X1_551/Y GND 0.26fF
C66453 PAND2X1_564/O GND 0.02fF
C66454 PAND2X1_552/A GND 0.20fF
C66455 PAND2X1_563/A GND 0.27fF
C66456 PAND2X1_642/B GND 0.36fF
C66457 POR2X1_518/Y GND 0.19fF
C66458 POR2X1_519/Y GND 0.14fF
C66459 POR2X1_549/B GND 0.25fF
C66460 POR2X1_590/Y GND 0.29fF
C66461 POR2X1_590/CTRL GND 0.02fF
C66462 PAND2X1_778/m4_208_n4# GND 0.00fF
C66463 PAND2X1_778/O GND 0.02fF
C66464 PAND2X1_793/A GND -0.13fF
C66465 PAND2X1_793/m4_208_n4# GND -0.01fF
C66466 POR2X1_773/B GND -4.10fF
C66467 PAND2X1_491/m4_208_n4# GND -0.01fF
C66468 POR2X1_757/A GND 0.16fF
C66469 PAND2X1_756/CTRL GND 0.02fF
C66470 POR2X1_781/B GND 0.17fF
C66471 PAND2X1_41/B GND 1.65fF
C66472 POR2X1_750/B GND 3.45fF
C66473 PAND2X1_737/B GND 0.26fF
C66474 PAND2X1_734/m4_208_n4# GND 0.00fF
C66475 PAND2X1_725/A GND 0.30fF
C66476 PAND2X1_707/Y GND 0.19fF
C66477 PAND2X1_712/m4_208_n4# GND 0.00fF
C66478 PAND2X1_712/CTRL GND 0.02fF
C66479 POR2X1_710/A GND -0.25fF
C66480 PAND2X1_701/m4_208_n4# GND 0.00fF
C66481 PAND2X1_717/Y GND 0.35fF
C66482 PAND2X1_216/m4_208_n4# GND -0.01fF
C66483 POR2X1_805/A GND 0.41fF
C66484 POR2X1_789/Y GND -0.10fF
C66485 POR2X1_793/m4_208_n4# GND 0.00fF
C66486 POR2X1_797/A GND 0.10fF
C66487 POR2X1_782/O GND 0.02fF
C66488 POR2X1_774/B GND -0.21fF
C66489 POR2X1_769/Y GND -0.01fF
C66490 POR2X1_771/m4_208_n4# GND -0.01fF
C66491 POR2X1_226/Y GND 0.35fF
C66492 POR2X1_226/CTRL GND 0.02fF
C66493 POR2X1_555/B GND 0.29fF
C66494 POR2X1_259/B GND -0.29fF
C66495 PAND2X1_89/m4_208_n4# GND -0.01fF
C66496 POR2X1_205/A GND 0.22fF
C66497 POR2X1_84/Y GND 0.30fF
C66498 PAND2X1_79/Y GND 0.33fF
C66499 POR2X1_205/Y GND 0.18fF
C66500 POR2X1_215/CTRL GND 0.02fF
C66501 POR2X1_418/CTRL2 GND 0.02fF
C66502 POR2X1_430/A GND 0.16fF
C66503 INPUT_7 GND 0.28fF
C66504 POR2X1_407/m4_208_n4# GND 0.00fF
C66505 POR2X1_183/Y GND -0.77fF
C66506 POR2X1_184/Y GND -1.77fF
C66507 PAND2X1_19/m4_208_n4# GND 0.00fF
C66508 POR2X1_400/B GND 0.16fF
C66509 PAND2X1_393/m4_208_n4# GND 0.00fF
C66510 POR2X1_68/B GND 1.17fF
C66511 PAND2X1_371/m4_208_n4# GND 0.00fF
C66512 PAND2X1_371/CTRL GND 0.02fF
C66513 PAND2X1_347/Y GND 0.20fF
C66514 PAND2X1_360/m4_208_n4# GND 0.00fF
C66515 POR2X1_29/A GND -2.62fF
C66516 PAND2X1_381/Y GND 0.22fF
C66517 PAND2X1_382/CTRL GND 0.02fF
C66518 POR2X1_597/A GND 0.31fF
C66519 PAND2X1_596/m4_208_n4# GND 0.00fF
C66520 POR2X1_637/B GND 0.32fF
C66521 PAND2X1_585/m4_208_n4# GND 0.00fF
C66522 PAND2X1_564/B GND 0.08fF
C66523 PAND2X1_570/B GND 0.21fF
C66524 PAND2X1_562/m4_208_n4# GND -0.01fF
C66525 PAND2X1_553/B GND 0.48fF
C66526 PAND2X1_344/m4_208_n4# GND -0.01fF
C66527 PAND2X1_575/B GND 0.30fF
C66528 POR2X1_516/Y GND 0.38fF
C66529 PAND2X1_574/CTRL GND 0.02fF
C66530 POR2X1_548/A GND -0.18fF
C66531 POR2X1_548/m4_208_n4# GND -0.01fF
C66532 PAND2X1_794/B GND 0.30fF
C66533 POR2X1_770/A GND -0.15fF
C66534 PAND2X1_90/Y GND 1.57fF
C66535 PAND2X1_766/m4_208_n4# GND 0.00fF
C66536 PAND2X1_784/A GND 0.22fF
C66537 PAND2X1_777/m4_208_n4# GND 0.00fF
C66538 PAND2X1_802/B GND 0.14fF
C66539 PAND2X1_539/Y GND 0.26fF
C66540 PAND2X1_593/Y GND 0.15fF
C66541 POR2X1_780/A GND 0.24fF
C66542 POR2X1_532/A GND -16.53fF
C66543 POR2X1_664/Y GND 0.32fF
C66544 PAND2X1_723/Y GND 0.18fF
C66545 PAND2X1_733/CTRL2 GND 0.02fF
C66546 PAND2X1_733/A GND -0.51fF
C66547 PAND2X1_718/Y GND 0.16fF
C66548 PAND2X1_719/Y GND 0.20fF
C66549 PAND2X1_722/m4_208_n4# GND 0.00fF
C66550 PAND2X1_726/B GND 0.61fF
C66551 PAND2X1_700/CTRL GND 0.02fF
C66552 POR2X1_805/B GND 0.27fF
C66553 POR2X1_791/Y GND 0.21fF
C66554 POR2X1_792/CTRL GND 0.02fF
C66555 POR2X1_771/A GND -0.06fF
C66556 POR2X1_770/m4_208_n4# GND 0.00fF
C66557 POR2X1_782/A GND -0.23fF
C66558 POR2X1_269/Y GND -0.05fF
C66559 POR2X1_258/Y GND 0.24fF
C66560 POR2X1_258/O GND 0.02fF
C66561 POR2X1_247/CTRL GND 0.02fF
C66562 POR2X1_225/m4_208_n4# GND 0.00fF
C66563 PAND2X1_72/Y GND 0.08fF
C66564 POR2X1_203/m4_208_n4# GND 0.00fF
C66565 POR2X1_219/B GND 0.25fF
C66566 POR2X1_208/Y GND 0.38fF
C66567 POR2X1_544/A GND 0.36fF
C66568 POR2X1_32/A GND 1.90fF
C66569 POR2X1_428/m4_208_n4# GND -0.01fF
C66570 POR2X1_283/A GND 1.59fF
C66571 POR2X1_417/m4_208_n4# GND 0.00fF
C66572 POR2X1_406/A GND 0.16fF
C66573 POR2X1_406/CTRL2 GND 0.02fF
C66574 POR2X1_609/A GND 0.21fF
C66575 PAND2X1_29/m4_208_n4# GND 0.00fF
C66576 PAND2X1_29/CTRL2 GND 0.02fF
C66577 PAND2X1_18/O GND 0.02fF
C66578 PAND2X1_474/A GND 0.28fF
C66579 PAND2X1_390/Y GND 0.18fF
C66580 PAND2X1_370/m4_208_n4# GND 0.00fF
C66581 POR2X1_636/A GND 0.16fF
C66582 POR2X1_643/A GND -0.11fF
C66583 PAND2X1_595/m4_208_n4# GND -0.00fF
C66584 PAND2X1_545/Y GND 0.14fF
C66585 PAND2X1_555/Y GND 0.26fF
C66586 PAND2X1_575/A GND 0.48fF
C66587 POR2X1_72/m4_208_n4# GND -0.01fF
C66588 PAND2X1_553/A GND 0.18fF
C66589 PAND2X1_540/CTRL GND 0.02fF
C66590 PAND2X1_556/B GND 0.29fF
C66591 PAND2X1_787/O GND 0.02fF
C66592 PAND2X1_354/A GND 0.17fF
C66593 PAND2X1_798/m4_208_n4# GND 0.00fF
C66594 POR2X1_770/B GND 0.20fF
C66595 PAND2X1_765/m4_208_n4# GND 0.00fF
C66596 POR2X1_780/B GND 0.04fF
C66597 PAND2X1_743/CTRL2 GND 0.02fF
C66598 POR2X1_790/A GND 0.29fF
C66599 PAND2X1_734/B GND 0.24fF
C66600 PAND2X1_673/Y GND 0.79fF
C66601 PAND2X1_738/B GND 0.22fF
C66602 PAND2X1_725/Y GND -0.69fF
C66603 PAND2X1_711/B GND -0.13fF
C66604 PAND2X1_710/CTRL GND 0.02fF
C66605 POR2X1_791/A GND 0.15fF
C66606 POR2X1_791/B GND 0.10fF
C66607 POR2X1_791/CTRL GND 0.02fF
C66608 POR2X1_783/A GND -0.29fF
C66609 PAND2X1_213/A GND -0.01fF
C66610 PAND2X1_209/m4_208_n4# GND 0.00fF
C66611 POR2X1_279/Y GND 0.16fF
C66612 POR2X1_279/CTRL2 GND 0.02fF
C66613 POR2X1_246/Y GND 0.14fF
C66614 POR2X1_245/Y GND 0.68fF
C66615 POR2X1_246/m4_208_n4# GND 0.00fF
C66616 POR2X1_257/Y GND 0.17fF
C66617 POR2X1_257/m4_208_n4# GND 0.00fF
C66618 POR2X1_268/Y GND 0.13fF
C66619 POR2X1_220/A GND 0.33fF
C66620 POR2X1_210/Y GND 0.21fF
C66621 POR2X1_213/O GND 0.02fF
C66622 POR2X1_224/Y GND 0.16fF
C66623 POR2X1_224/m4_208_n4# GND 0.00fF
C66624 POR2X1_206/A GND 0.11fF
C66625 POR2X1_202/m4_208_n4# GND 0.00fF
C66626 POR2X1_832/B GND 0.43fF
C66627 POR2X1_427/Y GND 0.28fF
C66628 POR2X1_72/B GND -7.12fF
C66629 POR2X1_438/Y GND 0.22fF
C66630 POR2X1_438/CTRL GND 0.02fF
C66631 POR2X1_405/Y GND 0.22fF
C66632 POR2X1_405/m4_208_n4# GND -0.00fF
C66633 POR2X1_416/m4_208_n4# GND 0.00fF
C66634 POR2X1_619/Y GND 0.02fF
C66635 POR2X1_608/O GND 0.02fF
C66636 POR2X1_194/A GND 0.23fF
C66637 PAND2X1_39/m4_208_n4# GND 0.00fF
C66638 PAND2X1_39/O GND 0.01fF
C66639 PAND2X1_28/CTRL2 GND 0.02fF
C66640 INPUT_6 GND 0.51fF
C66641 PAND2X1_17/m4_208_n4# GND 0.00fF
C66642 PAND2X1_17/CTRL GND 0.01fF
C66643 POR2X1_460/B GND 0.13fF
C66644 PAND2X1_392/B GND 0.19fF
C66645 POR2X1_653/B GND -0.05fF
C66646 POR2X1_186/Y GND 1.31fF
C66647 POR2X1_636/B GND 0.32fF
C66648 PAND2X1_583/m4_208_n4# GND 0.00fF
C66649 PAND2X1_546/Y GND 0.21fF
C66650 PAND2X1_550/m4_208_n4# GND 0.00fF
C66651 PAND2X1_558/Y GND 0.25fF
C66652 PAND2X1_576/B GND 0.30fF
C66653 PAND2X1_124/Y GND 0.36fF
C66654 PAND2X1_267/Y GND -0.45fF
C66655 PAND2X1_782/Y GND -0.01fF
C66656 PAND2X1_797/m4_208_n4# GND 0.00fF
C66657 PAND2X1_785/A GND 0.21fF
C66658 PAND2X1_795/B GND 0.21fF
C66659 PAND2X1_84/Y GND 0.31fF
C66660 PAND2X1_786/m4_208_n4# GND 0.00fF
C66661 POR2X1_769/A GND 0.12fF
C66662 PAND2X1_752/Y GND 0.25fF
C66663 PAND2X1_753/m4_208_n4# GND -0.00fF
C66664 GATE_741 GND 0.19fF
C66665 PAND2X1_740/Y GND 0.57fF
C66666 PAND2X1_675/m4_208_n4# GND -0.01fF
C66667 PAND2X1_721/B GND 0.29fF
C66668 POR2X1_667/Y GND 0.19fF
C66669 PAND2X1_720/m4_208_n4# GND 0.00fF
C66670 PAND2X1_720/CTRL2 GND 0.02fF
C66671 PAND2X1_738/A GND 0.20fF
C66672 PAND2X1_731/O GND 0.02fF
C66673 POR2X1_793/A GND 0.28fF
C66674 POR2X1_790/B GND 0.08fF
C66675 PAND2X1_222/B GND 0.31fF
C66676 PAND2X1_219/m4_208_n4# GND 0.00fF
C66677 PAND2X1_214/B GND 0.21fF
C66678 PAND2X1_35/Y GND 0.60fF
C66679 PAND2X1_198/Y GND 0.19fF
C66680 PAND2X1_208/CTRL2 GND 0.02fF
C66681 POR2X1_289/Y GND 0.26fF
C66682 POR2X1_289/CTRL GND 0.02fF
C66683 POR2X1_278/O GND 0.02fF
C66684 POR2X1_37/Y GND 1.07fF
C66685 POR2X1_245/m4_208_n4# GND 0.00fF
C66686 POR2X1_256/Y GND 0.19fF
C66687 POR2X1_255/Y GND 0.48fF
C66688 PAND2X1_6/A GND 1.09fF
C66689 POR2X1_256/m4_208_n4# GND 0.00fF
C66690 POR2X1_267/CTRL GND 0.02fF
C66691 POR2X1_220/B GND 0.36fF
C66692 POR2X1_234/m4_208_n4# GND 0.00fF
C66693 D_GATE_222 GND 0.61fF
C66694 POR2X1_222/Y GND -1.48fF
C66695 POR2X1_221/Y GND 0.12fF
C66696 POR2X1_223/m4_208_n4# GND 0.00fF
C66697 POR2X1_223/CTRL GND 0.02fF
C66698 PAND2X1_65/Y GND 0.28fF
C66699 POR2X1_61/Y GND 0.32fF
C66700 POR2X1_459/B GND 0.13fF
C66701 POR2X1_459/O GND 0.02fF
C66702 POR2X1_448/A GND 0.08fF
C66703 POR2X1_448/B GND 0.12fF
C66704 POR2X1_448/CTRL GND 0.02fF
C66705 POR2X1_437/CTRL2 GND 0.02fF
C66706 POR2X1_426/Y GND 0.17fF
C66707 POR2X1_425/Y GND 0.36fF
C66708 POR2X1_426/m4_208_n4# GND 0.00fF
C66709 POR2X1_415/Y GND 0.20fF
C66710 POR2X1_415/m4_208_n4# GND 0.00fF
C66711 POR2X1_403/Y GND 0.20fF
C66712 POR2X1_404/CTRL2 GND 0.02fF
C66713 POR2X1_630/A GND 0.42fF
C66714 POR2X1_629/B GND 0.12fF
C66715 POR2X1_619/A GND 0.31fF
C66716 POR2X1_38/B GND 0.69fF
C66717 POR2X1_618/m4_208_n4# GND 0.00fF
C66718 POR2X1_607/Y GND 0.16fF
C66719 POR2X1_607/m4_208_n4# GND 0.00fF
C66720 PAND2X1_49/m4_208_n4# GND -0.01fF
C66721 PAND2X1_49/CTRL GND 0.02fF
C66722 POR2X1_194/B GND 0.22fF
C66723 PAND2X1_16/m4_208_n4# GND 0.00fF
C66724 PAND2X1_16/O GND 0.01fF
C66725 PAND2X1_388/Y GND 0.06fF
C66726 PAND2X1_389/Y GND 0.08fF
C66727 PAND2X1_390/m4_208_n4# GND 0.00fF
C66728 PAND2X1_592/Y GND 0.19fF
C66729 PAND2X1_593/O GND 0.02fF
C66730 PAND2X1_581/Y GND 0.16fF
C66731 PAND2X1_582/m4_208_n4# GND 0.00fF
C66732 PAND2X1_561/Y GND 0.20fF
C66733 PAND2X1_571/A GND 0.38fF
C66734 PAND2X1_803/A GND -0.47fF
C66735 PAND2X1_783/Y GND 0.15fF
C66736 PAND2X1_776/Y GND 0.24fF
C66737 PAND2X1_785/CTRL2 GND 0.02fF
C66738 PAND2X1_762/Y GND 0.08fF
C66739 PAND2X1_763/m4_208_n4# GND 0.00fF
C66740 PAND2X1_771/Y GND 1.01fF
C66741 PAND2X1_773/Y GND 0.28fF
C66742 PAND2X1_580/m4_208_n4# GND -0.01fF
C66743 PAND2X1_739/B GND -0.04fF
C66744 PAND2X1_730/CTRL GND 0.02fF
C66745 PAND2X1_742/B GND -0.40fF
C66746 PAND2X1_736/Y GND 0.17fF
C66747 POR2X1_231/B GND 0.29fF
C66748 PAND2X1_214/A GND 0.19fF
C66749 PAND2X1_200/Y GND 0.16fF
C66750 PAND2X1_222/A GND 0.53fF
C66751 POR2X1_7/m4_208_n4# GND -0.01fF
C66752 POR2X1_362/B GND -0.93fF
C66753 POR2X1_286/Y GND 0.01fF
C66754 POR2X1_288/m4_208_n4# GND -0.00fF
C66755 POR2X1_299/Y GND -0.07fF
C66756 POR2X1_299/O GND 0.02fF
C66757 POR2X1_255/m4_208_n4# GND 0.00fF
C66758 POR2X1_267/A GND 0.30fF
C66759 POR2X1_266/m4_208_n4# GND 0.00fF
C66760 POR2X1_278/A GND 0.17fF
C66761 POR2X1_277/m4_208_n4# GND 0.00fF
C66762 POR2X1_243/Y GND -1.70fF
C66763 POR2X1_244/m4_208_n4# GND 0.00fF
C66764 POR2X1_218/Y GND 0.17fF
C66765 POR2X1_222/m4_208_n4# GND 0.00fF
C66766 POR2X1_212/A GND 0.39fF
C66767 POR2X1_211/m4_208_n4# GND 0.00fF
C66768 POR2X1_233/m4_208_n4# GND 0.00fF
C66769 POR2X1_207/A GND 0.28fF
C66770 POR2X1_193/Y GND 0.30fF
C66771 POR2X1_200/m4_208_n4# GND 0.00fF
C66772 POR2X1_478/B GND 0.39fF
C66773 POR2X1_468/Y GND 0.14fF
C66774 POR2X1_469/O GND 0.02fF
C66775 POR2X1_435/Y GND 0.56fF
C66776 POR2X1_458/m4_208_n4# GND -0.00fF
C66777 POR2X1_458/CTRL2 GND 0.02fF
C66778 POR2X1_454/A GND 0.36fF
C66779 POR2X1_447/A GND -0.14fF
C66780 POR2X1_447/CTRL GND 0.02fF
C66781 POR2X1_425/m4_208_n4# GND 0.00fF
C66782 POR2X1_403/B GND -0.53fF
C66783 POR2X1_403/m4_208_n4# GND -0.00fF
C66784 POR2X1_414/Y GND 0.35fF
C66785 POR2X1_414/m4_208_n4# GND 0.00fF
C66786 POR2X1_628/Y GND 0.35fF
C66787 POR2X1_93/A GND 0.71fF
C66788 POR2X1_628/m4_208_n4# GND 0.00fF
C66789 POR2X1_635/Y GND 0.12fF
C66790 POR2X1_639/m4_208_n4# GND 0.00fF
C66791 POR2X1_606/Y GND 0.19fF
C66792 POR2X1_121/B GND 1.46fF
C66793 POR2X1_590/A GND 1.33fF
C66794 POR2X1_606/m4_208_n4# GND 0.00fF
C66795 POR2X1_38/Y GND -7.07fF
C66796 POR2X1_617/CTRL2 GND 0.02fF
C66797 PAND2X1_37/m4_208_n4# GND 0.00fF
C66798 PAND2X1_59/CTRL GND 0.02fF
C66799 PAND2X1_48/m4_208_n4# GND 0.00fF
C66800 PAND2X1_15/m4_208_n4# GND 0.00fF
C66801 POR2X1_66/A GND -0.54fF
C66802 PAND2X1_26/CTRL GND 0.02fF
C66803 POR2X1_809/m4_208_n4# GND 0.00fF
C66804 PAND2X1_581/m4_208_n4# GND 0.00fF
C66805 PAND2X1_577/B GND 0.20fF
C66806 PAND2X1_562/Y GND 0.27fF
C66807 PAND2X1_592/m4_208_n4# GND 0.00fF
C66808 PAND2X1_796/B GND 0.39fF
C66809 PAND2X1_778/Y GND 0.12fF
C66810 PAND2X1_784/m4_208_n4# GND 0.00fF
C66811 PAND2X1_804/B GND 0.50fF
C66812 PAND2X1_785/Y GND 0.34fF
C66813 PAND2X1_795/O GND 0.02fF
C66814 PAND2X1_11/Y GND -1.31fF
C66815 PAND2X1_762/m4_208_n4# GND 0.00fF
C66816 PAND2X1_773/O GND 0.02fF
C66817 POR2X1_789/A GND 0.21fF
C66818 PAND2X1_738/Y GND -12.84fF
C66819 PAND2X1_739/Y GND 0.07fF
C66820 PAND2X1_740/m4_208_n4# GND 0.00fF
C66821 POR2X1_506/B GND 0.46fF
C66822 PAND2X1_239/m4_208_n4# GND 0.00fF
C66823 PAND2X1_218/B GND 0.19fF
C66824 PAND2X1_341/A GND 0.37fF
C66825 PAND2X1_228/m4_208_n4# GND 0.00fF
C66826 PAND2X1_215/B GND 0.64fF
C66827 PAND2X1_206/CTRL GND 0.02fF
C66828 POR2X1_288/A GND 0.32fF
C66829 POR2X1_298/Y GND 0.14fF
C66830 POR2X1_298/CTRL2 GND 0.02fF
C66831 POR2X1_276/B GND 0.25fF
C66832 POR2X1_366/m4_208_n4# GND -0.01fF
C66833 POR2X1_483/B GND 0.19fF
C66834 POR2X1_254/CTRL2 GND 0.02fF
C66835 POR2X1_667/A GND 0.69fF
C66836 POR2X1_265/CTRL2 GND 0.02fF
C66837 POR2X1_243/B GND 0.17fF
C66838 POR2X1_243/m4_208_n4# GND 0.00fF
C66839 POR2X1_232/Y GND 0.08fF
C66840 POR2X1_232/m4_208_n4# GND 0.00fF
C66841 POR2X1_232/CTRL GND 0.02fF
C66842 POR2X1_220/Y GND -2.51fF
C66843 POR2X1_192/Y GND -19.08fF
C66844 POR2X1_294/m4_208_n4# GND -0.01fF
C66845 POR2X1_210/m4_208_n4# GND 0.00fF
C66846 POR2X1_407/Y GND 0.30fF
C66847 PAND2X1_408/Y GND 0.15fF
C66848 POR2X1_480/A GND -6.18fF
C66849 POR2X1_476/Y GND 0.18fF
C66850 POR2X1_479/m4_208_n4# GND 0.00fF
C66851 POR2X1_468/O GND 0.02fF
C66852 POR2X1_370/Y GND 0.31fF
C66853 POR2X1_457/B GND 0.17fF
C66854 POR2X1_457/m4_208_n4# GND 0.00fF
C66855 POR2X1_457/CTRL2 GND 0.02fF
C66856 POR2X1_454/B GND 0.18fF
C66857 POR2X1_446/CTRL GND 0.02fF
C66858 POR2X1_435/B GND 0.13fF
C66859 POR2X1_722/m4_208_n4# GND -0.01fF
C66860 POR2X1_424/m4_208_n4# GND -0.00fF
C66861 POR2X1_404/B GND -0.41fF
C66862 POR2X1_402/B GND 0.13fF
C66863 POR2X1_402/m4_208_n4# GND 0.00fF
C66864 POR2X1_413/m4_208_n4# GND 0.00fF
C66865 POR2X1_655/A GND 0.26fF
C66866 POR2X1_643/Y GND 0.29fF
C66867 POR2X1_649/m4_208_n4# GND 0.00fF
C66868 POR2X1_638/B GND 0.15fF
C66869 POR2X1_638/m4_208_n4# GND 0.00fF
C66870 POR2X1_627/Y GND 0.13fF
C66871 POR2X1_718/A GND 0.76fF
C66872 POR2X1_605/CTRL GND 0.02fF
C66873 POR2X1_616/CTRL GND 0.02fF
C66874 POR2X1_202/A GND -2.62fF
C66875 POR2X1_68/Y GND 0.13fF
C66876 PAND2X1_69/m4_208_n4# GND 0.00fF
C66877 PAND2X1_69/CTRL2 GND 0.02fF
C66878 POR2X1_61/B GND 0.08fF
C66879 PAND2X1_58/m4_208_n4# GND 0.00fF
C66880 PAND2X1_36/m4_208_n4# GND -0.00fF
C66881 PAND2X1_59/B GND 0.19fF
C66882 PAND2X1_25/m4_208_n4# GND 0.00fF
C66883 POR2X1_820/A GND -0.06fF
C66884 POR2X1_94/A GND 1.03fF
C66885 POR2X1_819/m4_208_n4# GND 0.00fF
C66886 POR2X1_811/A GND 0.59fF
C66887 POR2X1_593/B GND 0.30fF
C66888 PAND2X1_591/m4_208_n4# GND 0.00fF
C66889 GATE_579 GND 0.17fF
C66890 PAND2X1_578/Y GND 0.00fF
C66891 PAND2X1_804/A GND 0.23fF
C66892 PAND2X1_787/Y GND 1.17fF
C66893 PAND2X1_794/CTRL GND 0.02fF
C66894 POR2X1_801/B GND 0.31fF
C66895 D_INPUT_0 GND 1.92fF
C66896 PAND2X1_779/Y GND 0.17fF
C66897 PAND2X1_783/m4_208_n4# GND 0.00fF
C66898 PAND2X1_773/B GND 0.20fF
C66899 PAND2X1_768/Y GND 0.17fF
C66900 PAND2X1_772/O GND 0.02fF
C66901 POR2X1_751/A GND 0.14fF
C66902 POR2X1_776/A GND 0.52fF
C66903 POR2X1_241/m4_208_n4# GND -0.01fF
C66904 PAND2X1_249/CTRL2 GND 0.02fF
C66905 PAND2X1_205/m4_208_n4# GND 0.00fF
C66906 PAND2X1_340/B GND -0.48fF
C66907 POR2X1_503/m4_208_n4# GND -0.01fF
C66908 PAND2X1_218/A GND 0.20fF
C66909 POR2X1_297/Y GND 0.28fF
C66910 POR2X1_297/m4_208_n4# GND 0.00fF
C66911 POR2X1_285/Y GND -0.21fF
C66912 POR2X1_286/m4_208_n4# GND 0.00fF
C66913 POR2X1_56/m4_208_n4# GND -0.01fF
C66914 POR2X1_275/Y GND 0.17fF
C66915 POR2X1_275/A GND 0.14fF
C66916 POR2X1_264/O GND 0.02fF
C66917 POR2X1_220/m4_208_n4# GND 0.00fF
C66918 POR2X1_341/A GND -4.32fF
C66919 POR2X1_244/B GND 0.49fF
C66920 POR2X1_241/Y GND 0.33fF
C66921 POR2X1_242/m4_208_n4# GND 0.00fF
C66922 PAND2X1_419/m4_208_n4# GND 0.00fF
C66923 PAND2X1_419/CTRL GND 0.02fF
C66924 PAND2X1_26/A GND -0.21fF
C66925 POR2X1_489/A GND 0.13fF
C66926 POR2X1_489/m4_208_n4# GND -0.01fF
C66927 POR2X1_477/Y GND 0.13fF
C66928 POR2X1_478/m4_208_n4# GND 0.00fF
C66929 POR2X1_452/Y GND -0.46fF
C66930 POR2X1_467/m4_208_n4# GND 0.00fF
C66931 POR2X1_455/A GND -0.36fF
C66932 POR2X1_445/m4_208_n4# GND 0.00fF
C66933 POR2X1_445/CTRL GND 0.02fF
C66934 POR2X1_465/A GND 0.17fF
C66935 POR2X1_456/m4_208_n4# GND 0.00fF
C66936 POR2X1_456/CTRL GND 0.02fF
C66937 POR2X1_423/Y GND 0.73fF
C66938 POR2X1_423/m4_208_n4# GND -0.00fF
C66939 POR2X1_436/B GND 0.29fF
C66940 POR2X1_434/A GND 0.19fF
C66941 POR2X1_434/CTRL GND 0.02fF
C66942 POR2X1_412/m4_208_n4# GND 0.00fF
C66943 POR2X1_412/CTRL2 GND 0.02fF
C66944 POR2X1_402/A GND 0.42fF
C66945 POR2X1_401/A GND 0.16fF
C66946 POR2X1_401/m4_208_n4# GND 0.00fF
C66947 POR2X1_638/A GND 0.20fF
C66948 POR2X1_637/m4_208_n4# GND 0.00fF
C66949 POR2X1_644/Y GND 0.22fF
C66950 POR2X1_648/CTRL GND 0.02fF
C66951 POR2X1_663/B GND 0.28fF
C66952 POR2X1_657/Y GND -0.20fF
C66953 POR2X1_615/Y GND 0.17fF
C66954 POR2X1_754/A GND 0.27fF
C66955 POR2X1_615/m4_208_n4# GND 0.00fF
C66956 POR2X1_615/CTRL GND 0.02fF
C66957 POR2X1_626/Y GND 0.06fF
C66958 POR2X1_626/m4_208_n4# GND 0.00fF
C66959 POR2X1_604/CTRL2 GND 0.02fF
C66960 POR2X1_78/Y GND -0.61fF
C66961 PAND2X1_79/CTRL GND 0.02fF
C66962 POR2X1_198/B GND 0.23fF
C66963 PAND2X1_57/m4_208_n4# GND 0.00fF
C66964 PAND2X1_46/m4_208_n4# GND 0.00fF
C66965 POR2X1_69/A GND -0.47fF
C66966 PAND2X1_68/m4_208_n4# GND 0.00fF
C66967 POR2X1_33/A GND 0.31fF
C66968 PAND2X1_24/m4_208_n4# GND 0.00fF
C66969 POR2X1_193/A GND -0.77fF
C66970 POR2X1_829/Y GND 0.10fF
C66971 POR2X1_811/B GND 0.43fF
C66972 POR2X1_805/Y GND 0.14fF
C66973 POR2X1_807/m4_208_n4# GND -0.00fF
C66974 POR2X1_818/Y GND -0.45fF
C66975 POR2X1_818/m4_208_n4# GND 0.00fF
C66976 POR2X1_591/A GND 0.11fF
C66977 PAND2X1_790/Y GND 0.16fF
C66978 PAND2X1_781/Y GND 0.15fF
C66979 PAND2X1_769/Y GND 0.18fF
C66980 POR2X1_800/A GND 0.32fF
C66981 PAND2X1_760/CTRL GND 0.02fF
C66982 POR2X1_247/Y GND 0.18fF
C66983 PAND2X1_248/CTRL GND 0.02fF
C66984 PAND2X1_259/m4_208_n4# GND 0.00fF
C66985 POR2X1_227/A GND 0.27fF
C66986 PAND2X1_226/m4_208_n4# GND 0.00fF
C66987 PAND2X1_205/B GND 0.22fF
C66988 POR2X1_79/Y GND 0.31fF
C66989 POR2X1_679/m4_208_n4# GND -0.01fF
C66990 PAND2X1_219/B GND 0.21fF
C66991 PAND2X1_205/Y GND 0.52fF
C66992 POR2X1_241/B GND 0.33fF
C66993 POR2X1_296/m4_208_n4# GND 0.00fF
C66994 POR2X1_285/A GND 0.08fF
C66995 POR2X1_274/Y GND 0.20fF
C66996 POR2X1_274/m4_208_n4# GND -0.00fF
C66997 POR2X1_274/O GND 0.01fF
C66998 POR2X1_63/m4_208_n4# GND -0.01fF
C66999 POR2X1_252/m4_208_n4# GND 0.00fF
C67000 POR2X1_252/CTRL2 GND 0.02fF
C67001 POR2X1_230/Y GND 0.16fF
C67002 PAND2X1_429/m4_208_n4# GND -0.00fF
C67003 POR2X1_409/B GND 0.50fF
C67004 PAND2X1_407/m4_208_n4# GND 0.00fF
C67005 POR2X1_446/A GND -0.00fF
C67006 POR2X1_488/Y GND 0.27fF
C67007 POR2X1_488/O GND 0.02fF
C67008 POR2X1_500/A GND 0.30fF
C67009 POR2X1_499/m4_208_n4# GND -0.00fF
C67010 POR2X1_477/m4_208_n4# GND 0.00fF
C67011 POR2X1_453/Y GND 0.13fF
C67012 POR2X1_466/CTRL GND 0.02fF
C67013 POR2X1_465/B GND 0.22fF
C67014 POR2X1_76/Y GND 0.27fF
C67015 POR2X1_455/m4_208_n4# GND 0.00fF
C67016 POR2X1_433/m4_208_n4# GND 0.00fF
C67017 POR2X1_422/Y GND 0.31fF
C67018 POR2X1_422/m4_208_n4# GND 0.00fF
C67019 POR2X1_422/O GND 0.02fF
C67020 POR2X1_444/B GND 0.21fF
C67021 POR2X1_444/m4_208_n4# GND 0.00fF
C67022 POR2X1_411/A GND 0.32fF
C67023 POR2X1_411/m4_208_n4# GND 0.00fF
C67024 POR2X1_403/A GND 0.00fF
C67025 POR2X1_400/A GND 0.32fF
C67026 POR2X1_400/m4_208_n4# GND 0.00fF
C67027 POR2X1_646/Y GND 0.15fF
C67028 POR2X1_647/m4_208_n4# GND 0.00fF
C67029 POR2X1_659/A GND 0.20fF
C67030 POR2X1_624/Y GND 0.43fF
C67031 POR2X1_658/m4_208_n4# GND 0.00fF
C67032 POR2X1_669/Y GND 0.20fF
C67033 POR2X1_669/m4_208_n4# GND 0.00fF
C67034 POR2X1_625/Y GND 0.19fF
C67035 POR2X1_625/m4_208_n4# GND -0.01fF
C67036 POR2X1_639/A GND 0.19fF
C67037 POR2X1_614/Y GND 0.31fF
C67038 POR2X1_614/m4_208_n4# GND 0.00fF
C67039 POR2X1_603/CTRL GND 0.02fF
C67040 POR2X1_79/A GND 0.18fF
C67041 PAND2X1_78/m4_208_n4# GND 0.00fF
C67042 POR2X1_202/B GND 0.19fF
C67043 PAND2X1_67/m4_208_n4# GND 0.00fF
C67044 PAND2X1_45/O GND 0.02fF
C67045 PAND2X1_55/Y GND 1.57fF
C67046 PAND2X1_56/m4_208_n4# GND 0.00fF
C67047 PAND2X1_23/m4_208_n4# GND 0.00fF
C67048 PAND2X1_35/B GND 0.19fF
C67049 POR2X1_27/Y GND 0.19fF
C67050 PAND2X1_3/A GND 0.29fF
C67051 POR2X1_808/m4_208_n4# GND -0.01fF
C67052 POR2X1_852/A GND 0.13fF
C67053 POR2X1_836/Y GND 0.20fF
C67054 POR2X1_835/Y GND 0.08fF
C67055 POR2X1_836/m4_208_n4# GND -0.00fF
C67056 POR2X1_839/CTRL GND 0.02fF
C67057 POR2X1_807/A GND 0.47fF
C67058 POR2X1_806/m4_208_n4# GND 0.00fF
C67059 PAND2X1_805/A GND 0.28fF
C67060 PAND2X1_792/m4_208_n4# GND 0.00fF
C67061 PAND2X1_781/m4_208_n4# GND 0.00fF
C67062 PAND2X1_771/B GND 0.18fF
C67063 POR2X1_259/A GND 0.21fF
C67064 PAND2X1_258/O GND 0.02fF
C67065 POR2X1_248/A GND 0.19fF
C67066 POR2X1_271/B GND 0.25fF
C67067 PAND2X1_236/m4_208_n4# GND 0.00fF
C67068 PAND2X1_225/m4_208_n4# GND 0.00fF
C67069 PAND2X1_219/A GND -0.45fF
C67070 PAND2X1_214/CTRL2 GND 0.02fF
C67071 PAND2X1_205/A GND 0.55fF
C67072 POR2X1_287/A GND 0.34fF
C67073 POR2X1_284/m4_208_n4# GND 0.00fF
C67074 POR2X1_284/CTRL GND 0.01fF
C67075 POR2X1_481/A GND 0.33fF
C67076 POR2X1_273/m4_208_n4# GND 0.00fF
C67077 POR2X1_262/m4_208_n4# GND 0.00fF
C67078 POR2X1_251/m4_208_n4# GND 0.00fF
C67079 POR2X1_243/A GND -0.06fF
C67080 POR2X1_240/m4_208_n4# GND 0.00fF
C67081 PAND2X1_428/m4_208_n4# GND 0.00fF
C67082 PAND2X1_406/m4_208_n4# GND 0.00fF
C67083 POR2X1_446/B GND 0.26fF
C67084 POR2X1_472/Y GND -0.17fF
C67085 POR2X1_476/m4_208_n4# GND 0.00fF
C67086 POR2X1_487/Y GND 0.15fF
C67087 POR2X1_487/m4_208_n4# GND 0.00fF
C67088 POR2X1_466/A GND -8.92fF
C67089 POR2X1_454/O GND 0.02fF
C67090 POR2X1_471/A GND 0.63fF
C67091 POR2X1_329/A GND 0.86fF
C67092 POR2X1_421/CTRL2 GND 0.02fF
C67093 POR2X1_432/Y GND 0.17fF
C67094 POR2X1_444/A GND 0.48fF
C67095 POR2X1_443/O GND 0.02fF
C67096 POR2X1_608/Y GND 0.10fF
C67097 PAND2X1_609/m4_208_n4# GND 0.00fF
C67098 POR2X1_679/Y GND 0.17fF
C67099 POR2X1_679/A GND 0.26fF
C67100 POR2X1_646/A GND -0.19fF
C67101 POR2X1_646/B GND 0.03fF
C67102 POR2X1_646/m4_208_n4# GND 0.00fF
C67103 POR2X1_668/Y GND 0.20fF
C67104 POR2X1_668/m4_208_n4# GND 0.00fF
C67105 POR2X1_141/Y GND 0.08fF
C67106 POR2X1_613/m4_208_n4# GND 0.00fF
C67107 POR2X1_613/CTRL GND 0.02fF
C67108 POR2X1_635/A GND 0.14fF
C67109 POR2X1_635/m4_208_n4# GND 0.00fF
C67110 POR2X1_623/Y GND 0.20fF
C67111 POR2X1_87/Y GND 0.12fF
C67112 PAND2X1_88/m4_208_n4# GND 0.00fF
C67113 POR2X1_788/A GND 0.28fF
C67114 POR2X1_602/A GND 0.13fF
C67115 POR2X1_602/m4_208_n4# GND 0.00fF
C67116 POR2X1_20/A GND 0.19fF
C67117 POR2X1_19/m4_208_n4# GND 0.00fF
C67118 PAND2X1_97/Y GND 0.02fF
C67119 PAND2X1_55/m4_208_n4# GND 0.00fF
C67120 PAND2X1_77/CTRL GND 0.02fF
C67121 POR2X1_67/A GND -1.34fF
C67122 PAND2X1_66/CTRL GND 0.02fF
C67123 PAND2X1_35/A GND 0.42fF
C67124 POR2X1_24/Y GND 0.24fF
C67125 PAND2X1_33/CTRL GND 0.02fF
C67126 PAND2X1_11/m4_208_n4# GND 0.00fF
C67127 PAND2X1_57/B GND 1.58fF
C67128 PAND2X1_44/m4_208_n4# GND 0.00fF
C67129 PAND2X1_58/A GND 1.64fF
C67130 POR2X1_859/A GND 0.32fF
C67131 POR2X1_852/B GND 0.33fF
C67132 POR2X1_837/Y GND 0.16fF
C67133 POR2X1_838/m4_208_n4# GND 0.00fF
C67134 POR2X1_805/CTRL GND 0.02fF
C67135 POR2X1_816/Y GND -0.40fF
C67136 POR2X1_816/m4_208_n4# GND 0.00fF
C67137 POR2X1_827/m4_208_n4# GND 0.00fF
C67138 PAND2X1_792/B GND 0.15fF
C67139 PAND2X1_783/B GND 0.23fF
C67140 POR2X1_744/Y GND 0.14fF
C67141 PAND2X1_257/m4_208_n4# GND 0.00fF
C67142 POR2X1_284/B GND 0.30fF
C67143 POR2X1_269/A GND 0.27fF
C67144 POR2X1_227/B GND 0.17fF
C67145 PAND2X1_224/m4_208_n4# GND 0.00fF
C67146 PAND2X1_85/Y GND -0.73fF
C67147 PAND2X1_213/m4_208_n4# GND 0.00fF
C67148 PAND2X1_9/Y GND 0.37fF
C67149 PAND2X1_206/B GND 1.11fF
C67150 POR2X1_67/Y GND 0.12fF
C67151 POR2X1_69/Y GND 0.09fF
C67152 POR2X1_272/Y GND -0.72fF
C67153 POR2X1_272/O GND 0.02fF
C67154 POR2X1_283/Y GND 0.30fF
C67155 POR2X1_283/m4_208_n4# GND 0.00fF
C67156 POR2X1_261/Y GND 0.21fF
C67157 POR2X1_411/B GND 2.19fF
C67158 POR2X1_261/m4_208_n4# GND 0.00fF
C67159 POR2X1_250/Y GND 0.59fF
C67160 POR2X1_250/CTRL GND 0.02fF
C67161 POR2X1_424/Y GND 0.15fF
C67162 PAND2X1_438/m4_208_n4# GND 0.00fF
C67163 PAND2X1_416/m4_208_n4# GND 0.00fF
C67164 PAND2X1_405/CTRL2 GND 0.02fF
C67165 POR2X1_479/B GND 0.26fF
C67166 POR2X1_734/B GND 0.32fF
C67167 POR2X1_475/m4_208_n4# GND 0.00fF
C67168 POR2X1_556/A GND -2.29fF
C67169 POR2X1_705/B GND 0.28fF
C67170 POR2X1_486/CTRL2 GND 0.02fF
C67171 POR2X1_458/Y GND 0.27fF
C67172 POR2X1_457/Y GND 0.13fF
C67173 POR2X1_464/m4_208_n4# GND 0.00fF
C67174 POR2X1_449/Y GND -0.14fF
C67175 POR2X1_448/Y GND -0.13fF
C67176 POR2X1_453/O GND 0.02fF
C67177 POR2X1_420/Y GND 0.13fF
C67178 POR2X1_102/Y GND 1.88fF
C67179 POR2X1_420/m4_208_n4# GND 0.00fF
C67180 POR2X1_431/Y GND 0.19fF
C67181 POR2X1_431/CTRL GND 0.02fF
C67182 PAND2X1_618/Y GND 0.08fF
C67183 PAND2X1_608/m4_208_n4# GND 0.00fF
C67184 POR2X1_689/CTRL GND 0.02fF
C67185 POR2X1_660/A GND 0.35fF
C67186 POR2X1_647/Y GND 0.16fF
C67187 POR2X1_656/m4_208_n4# GND 0.00fF
C67188 POR2X1_678/Y GND 0.28fF
C67189 POR2X1_260/B GND 1.45fF
C67190 POR2X1_678/CTRL2 GND 0.02fF
C67191 POR2X1_667/m4_208_n4# GND 0.00fF
C67192 POR2X1_667/CTRL2 GND 0.02fF
C67193 POR2X1_648/A GND 0.13fF
C67194 POR2X1_645/O GND 0.02fF
C67195 POR2X1_640/A GND 0.03fF
C67196 POR2X1_623/B GND 0.24fF
C67197 POR2X1_623/CTRL2 GND 0.02fF
C67198 POR2X1_612/Y GND 0.71fF
C67199 POR2X1_612/B GND 0.20fF
C67200 POR2X1_612/m4_208_n4# GND 0.00fF
C67201 POR2X1_20/B GND 1.54fF
C67202 POR2X1_18/m4_208_n4# GND 0.00fF
C67203 POR2X1_601/m4_208_n4# GND 0.00fF
C67204 PAND2X1_99/B GND 0.20fF
C67205 POR2X1_93/Y GND 0.24fF
C67206 POR2X1_88/A GND 0.14fF
C67207 PAND2X1_87/CTRL GND 0.02fF
C67208 PAND2X1_54/CTRL GND 0.02fF
C67209 PAND2X1_76/Y GND -1.42fF
C67210 PAND2X1_76/CTRL2 GND 0.02fF
C67211 PAND2X1_65/O GND 0.02fF
C67212 POR2X1_195/A GND 0.20fF
C67213 PAND2X1_43/m4_208_n4# GND 0.00fF
C67214 PAND2X1_43/CTRL2 GND 0.02fF
C67215 PAND2X1_32/CTRL2 GND 0.02fF
C67216 POR2X1_862/A GND -1.64fF
C67217 POR2X1_848/Y GND 0.12fF
C67218 POR2X1_859/m4_208_n4# GND 0.00fF
C67219 POR2X1_859/O GND 0.02fF
C67220 POR2X1_846/Y GND 0.17fF
C67221 POR2X1_848/m4_208_n4# GND 0.00fF
C67222 POR2X1_848/O GND 0.02fF
C67223 POR2X1_837/A GND 0.30fF
C67224 POR2X1_837/B GND 0.12fF
C67225 POR2X1_837/m4_208_n4# GND 0.00fF
C67226 POR2X1_808/A GND 0.48fF
C67227 POR2X1_815/Y GND 0.17fF
C67228 POR2X1_815/A GND 0.15fF
C67229 POR2X1_753/Y GND 0.29fF
C67230 POR2X1_754/Y GND 0.14fF
C67231 PAND2X1_289/m4_208_n4# GND 0.00fF
C67232 POR2X1_9/Y GND 1.27fF
C67233 POR2X1_240/A GND 0.19fF
C67234 PAND2X1_234/m4_208_n4# GND 0.00fF
C67235 GATE_222 GND 0.09fF
C67236 PAND2X1_221/Y GND 0.55fF
C67237 PAND2X1_365/m4_208_n4# GND -0.01fF
C67238 POR2X1_777/B GND 1.54fF
C67239 PAND2X1_245/m4_208_n4# GND 0.00fF
C67240 PAND2X1_220/A GND 0.14fF
C67241 PAND2X1_352/A GND 0.19fF
C67242 PAND2X1_212/m4_208_n4# GND 0.00fF
C67243 PAND2X1_206/A GND 0.54fF
C67244 POR2X1_65/m4_208_n4# GND -0.00fF
C67245 PAND2X1_201/CTRL GND 0.02fF
C67246 POR2X1_282/Y GND 0.06fF
C67247 POR2X1_282/m4_208_n4# GND 0.00fF
C67248 POR2X1_293/m4_208_n4# GND 0.00fF
C67249 POR2X1_271/Y GND 0.36fF
C67250 POR2X1_271/O GND 0.02fF
C67251 POR2X1_260/m4_208_n4# GND 0.00fF
C67252 POR2X1_376/Y GND 0.14fF
C67253 PAND2X1_459/CTRL GND 0.02fF
C67254 PAND2X1_453/A GND 0.44fF
C67255 POR2X1_421/Y GND 0.16fF
C67256 PAND2X1_448/CTRL2 GND 0.02fF
C67257 POR2X1_416/A GND 0.19fF
C67258 PAND2X1_415/m4_208_n4# GND 0.00fF
C67259 PAND2X1_415/CTRL2 GND 0.02fF
C67260 PAND2X1_425/Y GND -0.44fF
C67261 PAND2X1_426/m4_208_n4# GND 0.00fF
C67262 POR2X1_440/B GND 0.08fF
C67263 PAND2X1_403/Y GND 0.11fF
C67264 PAND2X1_404/m4_208_n4# GND -0.01fF
C67265 POR2X1_496/Y GND -5.54fF
C67266 POR2X1_460/Y GND 0.00fF
C67267 POR2X1_459/Y GND 0.17fF
C67268 POR2X1_475/A GND 0.20fF
C67269 POR2X1_860/A GND 0.07fF
C67270 POR2X1_474/m4_208_n4# GND 0.00fF
C67271 POR2X1_430/Y GND 0.16fF
C67272 POR2X1_669/B GND 3.36fF
C67273 POR2X1_450/Y GND 0.14fF
C67274 POR2X1_441/Y GND -0.45fF
C67275 POR2X1_441/m4_208_n4# GND 0.00fF
C67276 PAND2X1_607/O GND 0.02fF
C67277 PAND2X1_630/B GND 0.20fF
C67278 POR2X1_748/A GND 0.54fF
C67279 POR2X1_14/Y GND 0.80fF
C67280 POR2X1_699/O GND 0.02fF
C67281 POR2X1_688/Y GND 0.26fF
C67282 PAND2X1_39/B GND 1.46fF
C67283 POR2X1_688/m4_208_n4# GND 0.00fF
C67284 POR2X1_648/Y GND 0.28fF
C67285 POR2X1_655/m4_208_n4# GND 0.00fF
C67286 POR2X1_677/Y GND 0.38fF
C67287 POR2X1_677/CTRL GND 0.02fF
C67288 POR2X1_666/Y GND -0.13fF
C67289 POR2X1_644/B GND 0.13fF
C67290 POR2X1_644/CTRL GND 0.02fF
C67291 POR2X1_624/B GND 0.21fF
C67292 POR2X1_622/B GND -0.15fF
C67293 POR2X1_622/CTRL2 GND 0.02fF
C67294 POR2X1_39/m4_208_n4# GND 0.00fF
C67295 POR2X1_28/m4_208_n4# GND 0.00fF
C67296 POR2X1_28/CTRL GND 0.02fF
C67297 POR2X1_600/Y GND 0.33fF
C67298 POR2X1_612/A GND 0.39fF
C67299 POR2X1_611/m4_208_n4# GND 0.00fF
C67300 PAND2X1_97/m4_208_n4# GND -0.01fF
C67301 PAND2X1_86/CTRL GND 0.02fF
C67302 D_INPUT_7 GND -1.40fF
C67303 POR2X1_17/m4_208_n4# GND 0.00fF
C67304 POR2X1_17/CTRL GND 0.01fF
C67305 POR2X1_76/A GND 0.52fF
C67306 PAND2X1_75/O GND 0.02fF
C67307 PAND2X1_19/Y GND 0.01fF
C67308 PAND2X1_20/m4_208_n4# GND 0.00fF
C67309 PAND2X1_53/m4_208_n4# GND 0.00fF
C67310 PAND2X1_42/m4_208_n4# GND -0.00fF
C67311 PAND2X1_42/O GND 0.01fF
C67312 POR2X1_862/B GND 0.32fF
C67313 POR2X1_858/m4_208_n4# GND 0.00fF
C67314 POR2X1_848/A GND 0.21fF
C67315 POR2X1_847/m4_208_n4# GND -0.00fF
C67316 POR2X1_847/CTRL GND 0.02fF
C67317 POR2X1_814/Y GND 0.13fF
C67318 POR2X1_814/A GND 3.18fF
C67319 POR2X1_825/Y GND 0.39fF
C67320 POR2X1_825/m4_208_n4# GND 0.00fF
C67321 POR2X1_836/A GND 0.03fF
C67322 POR2X1_836/B GND 0.14fF
C67323 POR2X1_836/CTRL GND 0.02fF
C67324 POR2X1_808/B GND 0.13fF
C67325 POR2X1_796/Y GND 0.09fF
C67326 PAND2X1_299/m4_208_n4# GND 0.00fF
C67327 POR2X1_633/A GND -0.30fF
C67328 PAND2X1_277/m4_208_n4# GND 0.00fF
C67329 PAND2X1_287/Y GND 0.30fF
C67330 PAND2X1_267/B GND 0.21fF
C67331 POR2X1_262/Y GND 0.41fF
C67332 PAND2X1_716/m4_208_n4# GND -0.01fF
C67333 PAND2X1_860/A GND -0.86fF
C67334 PAND2X1_242/Y GND 1.04fF
C67335 PAND2X1_223/B GND 0.30fF
C67336 PAND2X1_799/m4_208_n4# GND -0.01fF
C67337 POR2X1_541/B GND 0.46fF
C67338 PAND2X1_255/m4_208_n4# GND 0.00fF
C67339 PAND2X1_193/Y GND -0.38fF
C67340 PAND2X1_200/m4_208_n4# GND 0.00fF
C67341 PAND2X1_212/B GND 0.34fF
C67342 PAND2X1_211/m4_208_n4# GND 0.00fF
C67343 POR2X1_292/Y GND 0.16fF
C67344 POR2X1_150/Y GND 0.81fF
C67345 POR2X1_295/m4_208_n4# GND -0.01fF
C67346 POR2X1_281/Y GND 0.19fF
C67347 POR2X1_281/CTRL GND 0.02fF
C67348 PAND2X1_469/O GND 0.02fF
C67349 PAND2X1_454/B GND 0.30fF
C67350 PAND2X1_447/m4_208_n4# GND 0.00fF
C67351 PAND2X1_464/B GND 0.19fF
C67352 PAND2X1_717/A GND 0.34fF
C67353 PAND2X1_458/CTRL2 GND 0.02fF
C67354 PAND2X1_425/m4_208_n4# GND 0.00fF
C67355 PAND2X1_425/CTRL GND 0.01fF
C67356 PAND2X1_435/Y GND -0.17fF
C67357 PAND2X1_436/m4_208_n4# GND 0.00fF
C67358 POR2X1_415/A GND -1.52fF
C67359 INPUT_3 GND -12.76fF
C67360 PAND2X1_414/m4_208_n4# GND 0.00fF
C67361 POR2X1_399/Y GND 0.17fF
C67362 PAND2X1_403/m4_208_n4# GND 0.00fF
C67363 POR2X1_484/m4_208_n4# GND 0.00fF
C67364 POR2X1_476/A GND 0.29fF
C67365 POR2X1_472/B GND 0.27fF
C67366 POR2X1_461/Y GND 0.18fF
C67367 POR2X1_462/m4_208_n4# GND 0.00fF
C67368 POR2X1_440/CTRL GND 0.01fF
C67369 POR2X1_452/A GND 0.16fF
C67370 POR2X1_451/A GND 0.21fF
C67371 POR2X1_635/B GND 0.32fF
C67372 POR2X1_451/m4_208_n4# GND 0.00fF
C67373 PAND2X1_635/Y GND 0.19fF
C67374 PAND2X1_639/O GND 0.02fF
C67375 POR2X1_607/A GND 0.50fF
C67376 PAND2X1_606/m4_208_n4# GND -0.00fF
C67377 PAND2X1_606/CTRL2 GND 0.02fF
C67378 POR2X1_621/A GND 0.39fF
C67379 POR2X1_630/B GND 0.28fF
C67380 PAND2X1_628/m4_208_n4# GND 0.00fF
C67381 POR2X1_698/Y GND -0.20fF
C67382 POR2X1_698/m4_208_n4# GND -0.00fF
C67383 POR2X1_698/CTRL GND 0.02fF
C67384 POR2X1_687/m4_208_n4# GND 0.00fF
C67385 POR2X1_676/m4_208_n4# GND 0.00fF
C67386 POR2X1_676/O GND 0.02fF
C67387 POR2X1_665/CTRL GND 0.02fF
C67388 POR2X1_643/m4_208_n4# GND 0.00fF
C67389 POR2X1_661/A GND 0.49fF
C67390 POR2X1_651/Y GND 0.29fF
C67391 POR2X1_654/m4_208_n4# GND 0.00fF
C67392 POR2X1_632/CTRL GND 0.02fF
C67393 POR2X1_622/A GND 0.17fF
C67394 POR2X1_621/CTRL2 GND 0.02fF
C67395 POR2X1_98/A GND -0.46fF
C67396 PAND2X1_94/Y GND -0.23fF
C67397 POR2X1_610/m4_208_n4# GND 0.00fF
C67398 POR2X1_610/O GND 0.02fF
C67399 POR2X1_49/CTRL GND 0.02fF
C67400 POR2X1_38/CTRL GND 0.02fF
C67401 PAND2X1_85/m4_208_n4# GND 0.00fF
C67402 POR2X1_16/m4_208_n4# GND -0.01fF
C67403 POR2X1_76/B GND -0.36fF
C67404 PAND2X1_41/m4_208_n4# GND 0.00fF
C67405 PAND2X1_30/m4_208_n4# GND 0.00fF
C67406 PAND2X1_810/B GND 0.28fF
C67407 POR2X1_846/A GND 0.13fF
C67408 POR2X1_846/m4_208_n4# GND 0.00fF
C67409 POR2X1_863/A GND 0.63fF
C67410 POR2X1_857/m4_208_n4# GND 0.00fF
C67411 POR2X1_263/Y GND -0.54fF
C67412 POR2X1_813/CTRL GND 0.02fF
C67413 POR2X1_835/A GND 0.18fF
C67414 POR2X1_835/B GND 0.12fF
C67415 POR2X1_234/A GND 0.26fF
C67416 POR2X1_824/m4_208_n4# GND 0.00fF
C67417 POR2X1_809/A GND 0.51fF
C67418 POR2X1_802/m4_208_n4# GND 0.00fF
C67419 POR2X1_302/B GND 0.24fF
C67420 PAND2X1_284/Y GND 0.20fF
C67421 PAND2X1_276/m4_208_n4# GND 0.00fF
C67422 POR2X1_267/B GND 0.33fF
C67423 PAND2X1_265/m4_208_n4# GND 0.00fF
C67424 POR2X1_240/B GND 0.35fF
C67425 PAND2X1_232/m4_208_n4# GND 0.00fF
C67426 PAND2X1_244/B GND 0.28fF
C67427 POR2X1_235/Y GND 0.17fF
C67428 POR2X1_230/m4_208_n4# GND -0.01fF
C67429 POR2X1_253/Y GND -0.53fF
C67430 PAND2X1_254/m4_208_n4# GND 0.00fF
C67431 PAND2X1_213/B GND 0.21fF
C67432 PAND2X1_210/m4_208_n4# GND 0.00fF
C67433 PAND2X1_192/Y GND -0.16fF
C67434 PAND2X1_220/Y GND 0.54fF
C67435 PAND2X1_221/m4_208_n4# GND 0.00fF
C67436 POR2X1_291/m4_208_n4# GND 0.00fF
C67437 POR2X1_280/Y GND 0.33fF
C67438 PAND2X1_787/A GND 0.44fF
C67439 PAND2X1_457/O GND 0.02fF
C67440 PAND2X1_469/B GND 0.45fF
C67441 PAND2X1_798/B GND -2.85fF
C67442 PAND2X1_652/A GND 0.74fF
C67443 PAND2X1_468/CTRL GND 0.02fF
C67444 PAND2X1_480/B GND 2.33fF
C67445 POR2X1_417/Y GND 0.43fF
C67446 POR2X1_418/Y GND 0.09fF
C67447 PAND2X1_446/CTRL2 GND 0.02fF
C67448 POR2X1_449/A GND -0.14fF
C67449 POR2X1_592/m4_208_n4# GND -0.01fF
C67450 POR2X1_433/Y GND 0.15fF
C67451 PAND2X1_404/A GND 0.42fF
C67452 POR2X1_397/Y GND 0.25fF
C67453 PAND2X1_402/m4_208_n4# GND 0.00fF
C67454 POR2X1_461/A GND 0.19fF
C67455 POR2X1_634/A GND 0.99fF
C67456 PAND2X1_413/m4_208_n4# GND 0.00fF
C67457 PAND2X1_413/O GND 0.02fF
C67458 POR2X1_463/Y GND 0.27fF
C67459 POR2X1_472/m4_208_n4# GND 0.00fF
C67460 POR2X1_494/CTRL GND 0.02fF
C67461 POR2X1_483/m4_208_n4# GND 0.00fF
C67462 POR2X1_461/B GND 0.20fF
C67463 POR2X1_450/A GND -0.23fF
C67464 POR2X1_450/B GND -0.52fF
C67465 PAND2X1_655/B GND -0.13fF
C67466 PAND2X1_643/Y GND 0.18fF
C67467 PAND2X1_649/CTRL GND 0.02fF
C67468 POR2X1_629/A GND 0.16fF
C67469 PAND2X1_627/m4_208_n4# GND 0.00fF
C67470 POR2X1_621/B GND 0.21fF
C67471 POR2X1_603/Y GND 0.33fF
C67472 POR2X1_604/Y GND 0.69fF
C67473 PAND2X1_605/CTRL2 GND 0.02fF
C67474 PAND2X1_651/A GND 0.09fF
C67475 POR2X1_588/Y GND 0.03fF
C67476 PAND2X1_638/m4_208_n4# GND 0.00fF
C67477 POR2X1_697/Y GND 0.35fF
C67478 POR2X1_675/A GND 0.15fF
C67479 POR2X1_439/Y GND 0.44fF
C67480 POR2X1_675/CTRL2 GND 0.01fF
C67481 POR2X1_78/A GND 1.21fF
C67482 PAND2X1_73/Y GND -10.52fF
C67483 POR2X1_664/O GND 0.02fF
C67484 POR2X1_687/A GND 0.37fF
C67485 POR2X1_686/m4_208_n4# GND -0.00fF
C67486 POR2X1_649/B GND 0.20fF
C67487 POR2X1_462/B GND 0.09fF
C67488 POR2X1_642/m4_208_n4# GND 0.00fF
C67489 POR2X1_661/B GND 0.18fF
C67490 POR2X1_652/Y GND 0.22fF
C67491 POR2X1_632/A GND 0.21fF
C67492 POR2X1_631/m4_208_n4# GND 0.00fF
C67493 POR2X1_60/A GND 2.23fF
C67494 POR2X1_59/m4_208_n4# GND 0.00fF
C67495 POR2X1_623/A GND 0.22fF
C67496 POR2X1_48/Y GND 0.18fF
C67497 POR2X1_48/CTRL2 GND 0.02fF
C67498 POR2X1_37/m4_208_n4# GND 0.00fF
C67499 POR2X1_83/B GND -3.81fF
C67500 POR2X1_26/m4_208_n4# GND 0.00fF
C67501 POR2X1_15/m4_208_n4# GND 0.00fF
C67502 PAND2X1_96/B GND 1.23fF
C67503 PAND2X1_95/O GND 0.02fF
C67504 POR2X1_81/Y GND 0.00fF
C67505 PAND2X1_84/m4_208_n4# GND -0.01fF
C67506 PAND2X1_73/m4_208_n4# GND 0.00fF
C67507 PAND2X1_47/B GND -0.28fF
C67508 PAND2X1_51/m4_208_n4# GND 0.00fF
C67509 PAND2X1_62/m4_208_n4# GND 0.00fF
C67510 PAND2X1_62/CTRL GND 0.02fF
C67511 POR2X1_108/Y GND 0.03fF
C67512 POR2X1_108/O GND 0.02fF
C67513 POR2X1_236/m4_208_n4# GND -0.01fF
C67514 PAND2X1_820/B GND 0.07fF
C67515 PAND2X1_803/Y GND -1.38fF
C67516 PAND2X1_808/CTRL2 GND 0.02fF
C67517 POR2X1_863/B GND 0.06fF
C67518 POR2X1_855/Y GND -0.19fF
C67519 POR2X1_856/m4_208_n4# GND 0.00fF
C67520 POR2X1_678/A GND 0.22fF
C67521 POR2X1_834/m4_208_n4# GND -0.00fF
C67522 POR2X1_849/A GND 0.38fF
C67523 POR2X1_673/Y GND 0.61fF
C67524 POR2X1_845/m4_208_n4# GND -0.00fF
C67525 POR2X1_845/CTRL GND 0.02fF
C67526 POR2X1_823/CTRL2 GND 0.02fF
C67527 D_GATE_811 GND 0.09fF
C67528 POR2X1_812/m4_208_n4# GND 0.00fF
C67529 POR2X1_809/B GND 0.12fF
C67530 POR2X1_801/m4_208_n4# GND 0.00fF
C67531 POR2X1_296/Y GND 0.12fF
C67532 PAND2X1_297/m4_208_n4# GND 0.00fF
C67533 PAND2X1_297/CTRL2 GND 0.02fF
C67534 POR2X1_276/A GND 0.11fF
C67535 PAND2X1_288/A GND 0.23fF
C67536 PAND2X1_264/m4_208_n4# GND 0.00fF
C67537 PAND2X1_241/Y GND 0.22fF
C67538 PAND2X1_231/O GND 0.02fF
C67539 POR2X1_254/A GND 0.27fF
C67540 PAND2X1_253/m4_208_n4# GND 0.00fF
C67541 PAND2X1_213/Y GND 0.34fF
C67542 PAND2X1_220/m4_208_n4# GND 0.00fF
C67543 POR2X1_290/Y GND -1.84fF
C67544 POR2X1_163/Y GND 0.35fF
C67545 PAND2X1_467/m4_208_n4# GND 0.00fF
C67546 PAND2X1_469/Y GND 0.19fF
C67547 PAND2X1_465/B GND -0.32fF
C67548 PAND2X1_254/Y GND 0.37fF
C67549 PAND2X1_557/A GND 0.63fF
C67550 PAND2X1_489/m4_208_n4# GND 0.00fF
C67551 PAND2X1_445/m4_208_n4# GND 0.00fF
C67552 PAND2X1_423/O GND 0.02fF
C67553 PAND2X1_436/A GND -0.60fF
C67554 PAND2X1_434/CTRL GND 0.02fF
C67555 PAND2X1_402/B GND -0.21fF
C67556 POR2X1_396/Y GND 0.15fF
C67557 PAND2X1_401/m4_208_n4# GND 0.00fF
C67558 PAND2X1_412/O GND 0.02fF
C67559 POR2X1_482/Y GND 0.22fF
C67560 POR2X1_482/m4_208_n4# GND 0.00fF
C67561 POR2X1_482/CTRL GND 0.02fF
C67562 POR2X1_558/B GND 0.33fF
C67563 POR2X1_493/A GND -0.11fF
C67564 POR2X1_493/m4_208_n4# GND 0.00fF
C67565 POR2X1_493/CTRL GND 0.01fF
C67566 POR2X1_460/A GND -0.55fF
C67567 POR2X1_477/A GND 0.35fF
C67568 POR2X1_464/Y GND 0.20fF
C67569 PAND2X1_644/Y GND 0.51fF
C67570 PAND2X1_645/Y GND 0.21fF
C67571 PAND2X1_648/m4_208_n4# GND 0.00fF
C67572 PAND2X1_203/m4_208_n4# GND -0.01fF
C67573 PAND2X1_626/m4_208_n4# GND 0.00fF
C67574 PAND2X1_626/O GND 0.01fF
C67575 PAND2X1_638/B GND 0.23fF
C67576 POR2X1_585/Y GND 0.16fF
C67577 POR2X1_586/Y GND 0.12fF
C67578 PAND2X1_637/m4_208_n4# GND 0.00fF
C67579 POR2X1_605/A GND 0.24fF
C67580 PAND2X1_604/m4_208_n4# GND 0.00fF
C67581 POR2X1_687/B GND 0.13fF
C67582 POR2X1_685/m4_208_n4# GND 0.00fF
C67583 POR2X1_696/Y GND 0.18fF
C67584 POR2X1_376/B GND 1.20fF
C67585 POR2X1_696/CTRL GND 0.02fF
C67586 POR2X1_674/Y GND -0.37fF
C67587 POR2X1_674/CTRL GND 0.02fF
C67588 POR2X1_440/Y GND -0.44fF
C67589 D_GATE_662 GND 0.11fF
C67590 POR2X1_662/Y GND -0.54fF
C67591 POR2X1_650/A GND 0.33fF
C67592 POR2X1_641/m4_208_n4# GND 0.00fF
C67593 POR2X1_632/B GND 0.04fF
C67594 POR2X1_630/CTRL GND 0.02fF
C67595 POR2X1_36/m4_208_n4# GND -0.00fF
C67596 POR2X1_47/m4_208_n4# GND 0.00fF
C67597 POR2X1_58/Y GND 0.04fF
C67598 POR2X1_58/CTRL GND 0.02fF
C67599 POR2X1_69/m4_208_n4# GND 0.00fF
C67600 POR2X1_84/A GND 0.34fF
C67601 PAND2X1_82/Y GND 0.29fF
C67602 PAND2X1_83/CTRL2 GND 0.02fF
C67603 POR2X1_14/m4_208_n4# GND -0.00fF
C67604 PAND2X1_72/m4_208_n4# GND 0.00fF
C67605 PAND2X1_50/m4_208_n4# GND 0.00fF
C67606 PAND2X1_61/Y GND 0.63fF
C67607 POR2X1_60/Y GND -0.33fF
C67608 POR2X1_118/Y GND 0.24fF
C67609 POR2X1_118/m4_208_n4# GND 0.00fF
C67610 POR2X1_107/CTRL GND 0.02fF
C67611 POR2X1_855/A GND 0.25fF
C67612 PAND2X1_65/B GND 1.46fF
C67613 POR2X1_828/Y GND 0.20fF
C67614 PAND2X1_829/O GND 0.02fF
C67615 PAND2X1_811/A GND 0.25fF
C67616 PAND2X1_805/Y GND 0.18fF
C67617 PAND2X1_818/CTRL GND 0.02fF
C67618 D_GATE_865 GND -0.18fF
C67619 POR2X1_866/m4_208_n4# GND 0.00fF
C67620 POR2X1_855/m4_208_n4# GND 0.00fF
C67621 POR2X1_849/B GND 0.13fF
C67622 POR2X1_844/CTRL GND 0.02fF
C67623 POR2X1_840/B GND 0.47fF
C67624 POR2X1_833/m4_208_n4# GND 0.00fF
C67625 POR2X1_822/O GND 0.02fF
C67626 POR2X1_801/A GND 0.18fF
C67627 POR2X1_800/m4_208_n4# GND 0.00fF
C67628 POR2X1_812/A GND 0.34fF
C67629 POR2X1_811/m4_208_n4# GND 0.00fF
C67630 POR2X1_273/Y GND 0.26fF
C67631 PAND2X1_274/m4_208_n4# GND 0.00fF
C67632 POR2X1_297/A GND 0.16fF
C67633 PAND2X1_296/m4_208_n4# GND 0.00fF
C67634 PAND2X1_286/B GND 0.30fF
C67635 PAND2X1_567/m4_208_n4# GND -0.01fF
C67636 PAND2X1_252/CTRL2 GND 0.02fF
C67637 POR2X1_237/Y GND 0.30fF
C67638 PAND2X1_241/m4_208_n4# GND 0.00fF
C67639 PAND2X1_263/m4_208_n4# GND -0.00fF
C67640 POR2X1_231/A GND 0.16fF
C67641 PAND2X1_478/B GND 0.34fF
C67642 PAND2X1_477/CTRL GND 0.02fF
C67643 PAND2X1_470/A GND 0.18fF
C67644 PAND2X1_466/CTRL2 GND 0.02fF
C67645 PAND2X1_488/CTRL2 GND 0.02fF
C67646 POR2X1_442/Y GND 0.20fF
C67647 PAND2X1_443/Y GND 0.25fF
C67648 PAND2X1_444/CTRL2 GND 0.02fF
C67649 POR2X1_832/A GND 0.41fF
C67650 PAND2X1_433/O GND 0.02fF
C67651 PAND2X1_445/Y GND -0.14fF
C67652 PAND2X1_455/m4_208_n4# GND 0.00fF
C67653 PAND2X1_403/B GND 0.11fF
C67654 POR2X1_393/Y GND -0.09fF
C67655 POR2X1_394/Y GND 0.18fF
C67656 PAND2X1_400/CTRL GND 0.02fF
C67657 PAND2X1_93/B GND -6.07fF
C67658 PAND2X1_422/m4_208_n4# GND 0.00fF
C67659 POR2X1_410/Y GND -0.13fF
C67660 PAND2X1_411/m4_208_n4# GND 0.00fF
C67661 POR2X1_481/Y GND 0.21fF
C67662 POR2X1_477/B GND 0.30fF
C67663 POR2X1_467/Y GND -0.99fF
C67664 POR2X1_466/Y GND 0.13fF
C67665 POR2X1_470/m4_208_n4# GND -0.00fF
C67666 POR2X1_470/O GND 0.02fF
C67667 PAND2X1_659/B GND 0.50fF
C67668 PAND2X1_669/m4_208_n4# GND -0.00fF
C67669 PAND2X1_656/B GND 0.21fF
C67670 PAND2X1_400/m4_208_n4# GND -0.00fF
C67671 PAND2X1_647/CTRL GND 0.02fF
C67672 POR2X1_631/A GND -0.02fF
C67673 PAND2X1_625/m4_208_n4# GND 0.00fF
C67674 PAND2X1_625/CTRL GND 0.02fF
C67675 PAND2X1_639/B GND 0.20fF
C67676 PAND2X1_614/m4_208_n4# GND 0.00fF
C67677 PAND2X1_614/CTRL2 GND 0.02fF
C67678 POR2X1_605/B GND 0.20fF
C67679 PAND2X1_603/O GND 0.02fF
C67680 POR2X1_695/Y GND 0.18fF
C67681 POR2X1_48/A GND 1.53fF
C67682 POR2X1_23/Y GND 1.48fF
C67683 POR2X1_695/m4_208_n4# GND 0.00fF
C67684 POR2X1_684/m4_208_n4# GND 0.00fF
C67685 POR2X1_673/m4_208_n4# GND 0.00fF
C67686 POR2X1_661/Y GND 0.00fF
C67687 POR2X1_660/Y GND 0.13fF
C67688 POR2X1_662/m4_208_n4# GND 0.00fF
C67689 POR2X1_639/Y GND 0.32fF
C67690 POR2X1_638/Y GND 0.09fF
C67691 POR2X1_633/Y GND -0.34fF
C67692 POR2X1_79/O GND 0.02fF
C67693 POR2X1_57/CTRL2 GND 0.02fF
C67694 POR2X1_46/CTRL GND 0.02fF
C67695 POR2X1_68/m4_208_n4# GND 0.00fF
C67696 POR2X1_68/CTRL2 GND 0.02fF
C67697 PAND2X1_82/CTRL2 GND 0.02fF
C67698 POR2X1_98/B GND 0.38fF
C67699 PAND2X1_93/m4_208_n4# GND 0.00fF
C67700 POR2X1_13/Y GND 0.36fF
C67701 POR2X1_13/CTRL GND 0.02fF
C67702 POR2X1_24/CTRL GND 0.02fF
C67703 POR2X1_34/Y GND 0.15fF
C67704 PAND2X1_60/m4_208_n4# GND 0.00fF
C67705 POR2X1_137/Y GND -0.65fF
C67706 POR2X1_140/B GND 0.51fF
C67707 POR2X1_128/m4_208_n4# GND 0.00fF
C67708 POR2X1_251/A GND 0.18fF
C67709 POR2X1_106/m4_208_n4# GND 0.00fF
C67710 PAND2X1_852/B GND 0.30fF
C67711 PAND2X1_835/Y GND 0.20fF
C67712 PAND2X1_839/CTRL GND 0.02fF
C67713 POR2X1_829/A GND 0.53fF
C67714 PAND2X1_828/CTRL GND 0.02fF
C67715 POR2X1_847/B GND 0.18fF
C67716 PAND2X1_807/B GND 0.27fF
C67717 PAND2X1_362/A GND -0.13fF
C67718 POR2X1_866/A GND 0.83fF
C67719 POR2X1_862/Y GND 0.13fF
C67720 POR2X1_865/m4_208_n4# GND 0.00fF
C67721 POR2X1_832/m4_208_n4# GND 0.00fF
C67722 POR2X1_832/CTRL GND 0.01fF
C67723 POR2X1_850/A GND 0.14fF
C67724 POR2X1_287/B GND 0.23fF
C67725 POR2X1_343/A GND 0.43fF
C67726 POR2X1_843/m4_208_n4# GND -0.00fF
C67727 POR2X1_856/B GND 1.76fF
C67728 POR2X1_567/B GND 2.42fF
C67729 POR2X1_854/m4_208_n4# GND 0.00fF
C67730 POR2X1_812/B GND 0.21fF
C67731 POR2X1_809/Y GND 0.14fF
C67732 POR2X1_821/CTRL GND 0.02fF
C67733 POR2X1_309/m4_208_n4# GND 0.00fF
C67734 POR2X1_346/A GND 0.27fF
C67735 POR2X1_294/Y GND 0.75fF
C67736 PAND2X1_295/m4_208_n4# GND 0.00fF
C67737 PAND2X1_284/CTRL2 GND 0.02fF
C67738 PAND2X1_243/B GND 0.36fF
C67739 POR2X1_234/Y GND 0.16fF
C67740 PAND2X1_240/m4_208_n4# GND 0.00fF
C67741 POR2X1_786/A GND -0.54fF
C67742 PAND2X1_262/m4_208_n4# GND 0.00fF
C67743 PAND2X1_262/O GND 0.01fF
C67744 PAND2X1_471/B GND 0.15fF
C67745 PAND2X1_455/Y GND -0.10fF
C67746 PAND2X1_465/m4_208_n4# GND 0.00fF
C67747 PAND2X1_465/CTRL GND 0.02fF
C67748 POR2X1_489/B GND -0.09fF
C67749 PAND2X1_479/B GND 0.20fF
C67750 PAND2X1_473/Y GND 0.20fF
C67751 PAND2X1_475/m4_208_n4# GND -0.01fF
C67752 PAND2X1_443/m4_208_n4# GND -0.00fF
C67753 PAND2X1_443/CTRL GND 0.02fF
C67754 PAND2X1_466/B GND 0.11fF
C67755 PAND2X1_446/Y GND -0.05fF
C67756 POR2X1_130/A GND 0.82fF
C67757 POR2X1_596/A GND 0.33fF
C67758 PAND2X1_421/m4_208_n4# GND 0.00fF
C67759 POR2X1_491/CTRL GND 0.02fF
C67760 D_GATE_479 GND 0.07fF
C67761 POR2X1_478/Y GND 0.13fF
C67762 POR2X1_480/m4_208_n4# GND 0.00fF
C67763 POR2X1_669/A GND 0.16fF
C67764 PAND2X1_668/m4_208_n4# GND 0.00fF
C67765 POR2X1_728/B GND 0.23fF
C67766 POR2X1_676/Y GND 0.16fF
C67767 PAND2X1_659/A GND 0.28fF
C67768 PAND2X1_217/B GND 0.82fF
C67769 PAND2X1_647/B GND 0.15fF
C67770 POR2X1_609/Y GND 0.52fF
C67771 PAND2X1_646/m4_208_n4# GND 0.00fF
C67772 POR2X1_428/Y GND 0.35fF
C67773 POR2X1_582/Y GND 0.14fF
C67774 PAND2X1_635/m4_208_n4# GND -0.00fF
C67775 PAND2X1_658/A GND -0.84fF
C67776 PAND2X1_623/Y GND -0.23fF
C67777 POR2X1_601/Y GND 0.20fF
C67778 PAND2X1_602/m4_208_n4# GND 0.00fF
C67779 POR2X1_620/A GND 0.20fF
C67780 POR2X1_694/Y GND 0.17fF
C67781 POR2X1_257/A GND 1.81fF
C67782 POR2X1_694/m4_208_n4# GND 0.00fF
C67783 POR2X1_683/Y GND 0.07fF
C67784 POR2X1_683/m4_208_n4# GND 0.00fF
C67785 POR2X1_661/m4_208_n4# GND 0.00fF
C67786 POR2X1_654/B GND -0.79fF
C67787 POR2X1_640/Y GND 0.09fF
C67788 POR2X1_89/Y GND 0.15fF
C67789 POR2X1_89/m4_208_n4# GND 0.00fF
C67790 POR2X1_672/Y GND 0.16fF
C67791 POR2X1_672/m4_208_n4# GND -0.00fF
C67792 POR2X1_45/Y GND 0.29fF
C67793 POR2X1_45/m4_208_n4# GND 0.00fF
C67794 POR2X1_78/m4_208_n4# GND 0.00fF
C67795 PAND2X1_92/CTRL GND 0.02fF
C67796 POR2X1_13/A GND 1.76fF
C67797 POR2X1_34/A GND 0.15fF
C67798 POR2X1_34/B GND 0.30fF
C67799 POR2X1_34/CTRL2 GND 0.02fF
C67800 POR2X1_84/B GND 0.29fF
C67801 PAND2X1_95/B GND -1.36fF
C67802 PAND2X1_70/m4_208_n4# GND 0.00fF
C67803 POR2X1_127/Y GND 0.21fF
C67804 POR2X1_127/CTRL GND 0.02fF
C67805 POR2X1_149/m4_208_n4# GND -0.01fF
C67806 POR2X1_139/A GND 0.19fF
C67807 POR2X1_114/Y GND 0.30fF
C67808 POR2X1_116/m4_208_n4# GND 0.00fF
C67809 POR2X1_105/Y GND 0.20fF
C67810 POR2X1_814/B GND 2.22fF
C67811 PAND2X1_859/B GND 0.35fF
C67812 PAND2X1_844/Y GND 0.26fF
C67813 POR2X1_838/B GND 0.45fF
C67814 PAND2X1_827/m4_208_n4# GND 0.00fF
C67815 PAND2X1_852/A GND 0.26fF
C67816 POR2X1_827/Y GND 0.19fF
C67817 PAND2X1_195/m4_208_n4# GND -0.00fF
C67818 PAND2X1_838/CTRL GND 0.02fF
C67819 PAND2X1_793/Y GND 0.48fF
C67820 POR2X1_866/B GND 0.18fF
C67821 POR2X1_774/Y GND 0.28fF
C67822 POR2X1_864/m4_208_n4# GND 0.00fF
C67823 POR2X1_864/CTRL GND 0.01fF
C67824 POR2X1_850/B GND 0.27fF
C67825 POR2X1_830/Y GND 0.23fF
C67826 POR2X1_842/m4_208_n4# GND 0.00fF
C67827 POR2X1_841/B GND 0.20fF
C67828 POR2X1_301/A GND 0.34fF
C67829 POR2X1_274/A GND 0.52fF
C67830 POR2X1_831/m4_208_n4# GND 0.00fF
C67831 POR2X1_857/A GND 0.14fF
C67832 POR2X1_820/Y GND 0.23fF
C67833 POR2X1_820/B GND -0.02fF
C67834 POR2X1_820/CTRL GND 0.02fF
C67835 POR2X1_317/Y GND 0.26fF
C67836 POR2X1_367/m4_208_n4# GND -0.01fF
C67837 POR2X1_307/Y GND 0.22fF
C67838 POR2X1_308/m4_208_n4# GND 0.00fF
C67839 PAND2X1_337/m4_208_n4# GND -0.01fF
C67840 POR2X1_286/B GND 0.24fF
C67841 PAND2X1_283/m4_208_n4# GND 0.00fF
C67842 POR2X1_260/Y GND 0.20fF
C67843 PAND2X1_261/CTRL GND 0.02fF
C67844 PAND2X1_250/m4_208_n4# GND -0.00fF
C67845 PAND2X1_272/m4_208_n4# GND 0.00fF
C67846 PAND2X1_272/CTRL GND 0.02fF
C67847 POR2X1_484/Y GND 0.03fF
C67848 POR2X1_485/Y GND 0.22fF
C67849 PAND2X1_486/CTRL GND 0.02fF
C67850 PAND2X1_479/A GND 0.21fF
C67851 POR2X1_406/Y GND 0.45fF
C67852 PAND2X1_474/Y GND 0.27fF
C67853 PAND2X1_79/m4_208_n4# GND -0.00fF
C67854 PAND2X1_497/CTRL GND 0.02fF
C67855 PAND2X1_457/Y GND 0.14fF
C67856 PAND2X1_464/O GND 0.02fF
C67857 PAND2X1_466/A GND 0.47fF
C67858 PAND2X1_449/Y GND 0.22fF
C67859 PAND2X1_442/m4_208_n4# GND 0.00fF
C67860 PAND2X1_420/m4_208_n4# GND 0.00fF
C67861 PAND2X1_431/m4_208_n4# GND 0.00fF
C67862 POR2X1_490/Y GND 0.31fF
C67863 POR2X1_490/CTRL GND 0.02fF
C67864 PAND2X1_689/m4_208_n4# GND 0.00fF
C67865 PAND2X1_678/O GND 0.02fF
C67866 POR2X1_720/B GND 0.19fF
C67867 POR2X1_264/Y GND 0.18fF
C67868 PAND2X1_667/m4_208_n4# GND 0.00fF
C67869 PAND2X1_660/B GND 0.38fF
C67870 POR2X1_394/m4_208_n4# GND -0.01fF
C67871 PAND2X1_656/CTRL GND 0.02fF
C67872 PAND2X1_640/B GND 0.17fF
C67873 PAND2X1_602/Y GND 0.54fF
C67874 PAND2X1_645/m4_208_n4# GND 0.00fF
C67875 PAND2X1_620/Y GND 0.19fF
C67876 PAND2X1_623/m4_208_n4# GND 0.00fF
C67877 PAND2X1_601/m4_208_n4# GND -0.00fF
C67878 POR2X1_647/B GND 0.09fF
C67879 POR2X1_610/Y GND 0.12fF
C67880 POR2X1_693/Y GND 0.33fF
C67881 POR2X1_682/Y GND 0.15fF
C67882 POR2X1_655/Y GND 0.19fF
C67883 POR2X1_660/m4_208_n4# GND -0.00fF
C67884 POR2X1_88/m4_208_n4# GND -0.00fF
C67885 POR2X1_88/CTRL GND 0.02fF
C67886 POR2X1_99/Y GND 0.24fF
C67887 POR2X1_99/CTRL2 GND 0.02fF
C67888 POR2X1_672/A GND 0.16fF
C67889 D_INPUT_2 GND -1.33fF
C67890 POR2X1_671/m4_208_n4# GND -0.00fF
C67891 POR2X1_55/CTRL2 GND 0.02fF
C67892 POR2X1_66/Y GND 0.00fF
C67893 POR2X1_66/m4_208_n4# GND 0.00fF
C67894 POR2X1_43/B GND 0.97fF
C67895 POR2X1_44/m4_208_n4# GND 0.00fF
C67896 POR2X1_35/B GND 0.37fF
C67897 POR2X1_33/B GND 0.20fF
C67898 POR2X1_33/m4_208_n4# GND 0.00fF
C67899 POR2X1_97/A GND -1.21fF
C67900 PAND2X1_91/O GND 0.02fF
C67901 POR2X1_12/A GND 0.87fF
C67902 D_INPUT_5 GND 0.33fF
C67903 POR2X1_11/m4_208_n4# GND 0.00fF
C67904 PAND2X1_81/B GND 0.26fF
C67905 PAND2X1_80/m4_208_n4# GND 0.00fF
C67906 POR2X1_149/A GND 0.30fF
C67907 POR2X1_137/B GND 0.13fF
C67908 POR2X1_113/m4_208_n4# GND -0.01fF
C67909 POR2X1_159/CTRL GND 0.02fF
C67910 POR2X1_126/m4_208_n4# GND 0.00fF
C67911 POR2X1_116/A GND -0.27fF
C67912 POR2X1_554/B GND 0.15fF
C67913 PAND2X1_862/B GND 0.18fF
C67914 PAND2X1_859/A GND 0.37fF
C67915 PAND2X1_848/m4_208_n4# GND 0.00fF
C67916 PAND2X1_826/m4_208_n4# GND 0.00fF
C67917 PAND2X1_838/B GND 0.39fF
C67918 POR2X1_826/Y GND 0.18fF
C67919 PAND2X1_837/m4_208_n4# GND 0.00fF
C67920 PAND2X1_837/CTRL2 GND 0.02fF
C67921 POR2X1_846/B GND 0.16fF
C67922 PAND2X1_808/B GND 0.07fF
C67923 PAND2X1_804/CTRL2 GND 0.02fF
C67924 POR2X1_851/A GND 0.21fF
C67925 POR2X1_832/Y GND 0.17fF
C67926 POR2X1_841/m4_208_n4# GND 0.00fF
C67927 POR2X1_864/A GND 0.60fF
C67928 POR2X1_863/m4_208_n4# GND 0.00fF
C67929 POR2X1_857/B GND 0.43fF
C67930 POR2X1_852/m4_208_n4# GND -0.00fF
C67931 POR2X1_852/CTRL GND 0.02fF
C67932 POR2X1_319/A GND 0.24fF
C67933 POR2X1_445/A GND 0.36fF
C67934 POR2X1_318/m4_208_n4# GND 0.00fF
C67935 POR2X1_329/Y GND 0.12fF
C67936 POR2X1_760/A GND 0.47fF
C67937 POR2X1_329/CTRL GND 0.02fF
C67938 POR2X1_307/B GND 0.10fF
C67939 POR2X1_307/m4_208_n4# GND 0.00fF
C67940 PAND2X1_293/m4_208_n4# GND 0.00fF
C67941 POR2X1_261/A GND 0.16fF
C67942 PAND2X1_260/m4_208_n4# GND 0.00fF
C67943 PAND2X1_282/m4_208_n4# GND 0.00fF
C67944 POR2X1_270/Y GND 0.33fF
C67945 PAND2X1_485/m4_208_n4# GND 0.00fF
C67946 PAND2X1_404/Y GND -0.95fF
C67947 POR2X1_499/A GND 0.70fF
C67948 PAND2X1_472/B GND 0.57fF
C67949 PAND2X1_459/Y GND 0.15fF
C67950 PAND2X1_460/Y GND -0.34fF
C67951 PAND2X1_463/CTRL GND 0.02fF
C67952 PAND2X1_467/B GND -0.39fF
C67953 POR2X1_443/A GND 0.33fF
C67954 PAND2X1_441/CTRL GND 0.02fF
C67955 PAND2X1_429/Y GND 0.10fF
C67956 PAND2X1_430/m4_208_n4# GND 0.00fF
C67957 PAND2X1_9/CTRL GND 0.02fF
C67958 POR2X1_709/A GND 0.23fF
C67959 PAND2X1_699/m4_208_n4# GND 0.00fF
C67960 POR2X1_689/A GND 0.25fF
C67961 PAND2X1_677/CTRL2 GND 0.02fF
C67962 POR2X1_719/A GND -0.33fF
C67963 PAND2X1_20/A GND 1.94fF
C67964 PAND2X1_666/O GND 0.02fF
C67965 PAND2X1_648/Y GND 0.19fF
C67966 POR2X1_597/Y GND 0.29fF
C67967 PAND2X1_644/m4_208_n4# GND 0.00fF
C67968 PAND2X1_633/m4_208_n4# GND 0.00fF
C67969 POR2X1_602/B GND 0.26fF
C67970 POR2X1_719/m4_208_n4# GND -0.01fF
C67971 PAND2X1_612/B GND 0.27fF
C67972 POR2X1_54/Y GND 1.63fF
C67973 PAND2X1_611/m4_208_n4# GND 0.00fF
C67974 PAND2X1_624/A GND 0.17fF
C67975 PAND2X1_621/Y GND 0.14fF
C67976 POR2X1_692/m4_208_n4# GND 0.00fF
C67977 POR2X1_681/Y GND 0.30fF
C67978 POR2X1_681/m4_208_n4# GND 0.00fF
C67979 POR2X1_670/m4_208_n4# GND 0.00fF
C67980 POR2X1_99/A GND 0.26fF
C67981 POR2X1_76/m4_208_n4# GND -0.01fF
C67982 POR2X1_65/Y GND 0.20fF
C67983 POR2X1_63/Y GND 0.58fF
C67984 POR2X1_65/CTRL GND 0.02fF
C67985 POR2X1_87/B GND 0.33fF
C67986 POR2X1_87/m4_208_n4# GND 0.00fF
C67987 POR2X1_54/m4_208_n4# GND 0.00fF
C67988 POR2X1_21/CTRL2 GND 0.02fF
C67989 POR2X1_32/Y GND 0.21fF
C67990 POR2X1_29/Y GND 0.12fF
C67991 POR2X1_32/CTRL GND 0.02fF
C67992 POR2X1_43/Y GND 0.25fF
C67993 POR2X1_43/m4_208_n4# GND 0.00fF
C67994 POR2X1_43/CTRL GND 0.02fF
C67995 PAND2X1_90/m4_208_n4# GND 0.00fF
C67996 POR2X1_169/B GND 0.14fF
C67997 POR2X1_169/m4_208_n4# GND 0.00fF
C67998 POR2X1_136/Y GND 0.18fF
C67999 POR2X1_136/m4_208_n4# GND 0.00fF
C68000 POR2X1_149/B GND 0.22fF
C68001 POR2X1_147/A GND -0.08fF
C68002 POR2X1_147/CTRL2 GND 0.02fF
C68003 POR2X1_158/Y GND 0.43fF
C68004 POR2X1_416/B GND 2.64fF
C68005 POR2X1_158/m4_208_n4# GND 0.00fF
C68006 POR2X1_125/Y GND 0.17fF
C68007 POR2X1_125/m4_208_n4# GND 0.00fF
C68008 POR2X1_113/Y GND -0.87fF
C68009 POR2X1_114/O GND 0.02fF
C68010 PAND2X1_850/Y GND 0.36fF
C68011 PAND2X1_858/m4_208_n4# GND 0.00fF
C68012 PAND2X1_825/m4_208_n4# GND 0.00fF
C68013 PAND2X1_839/B GND 0.23fF
C68014 POR2X1_823/Y GND 0.23fF
C68015 POR2X1_824/Y GND 0.19fF
C68016 PAND2X1_836/m4_208_n4# GND 0.00fF
C68017 PAND2X1_836/CTRL2 GND 0.02fF
C68018 PAND2X1_848/B GND -0.27fF
C68019 POR2X1_817/Y GND 0.01fF
C68020 PAND2X1_797/Y GND 0.37fF
C68021 PAND2X1_803/O GND 0.02fF
C68022 PAND2X1_814/m4_208_n4# GND 0.00fF
C68023 POR2X1_862/m4_208_n4# GND 0.00fF
C68024 POR2X1_858/A GND 0.17fF
C68025 POR2X1_840/Y GND 0.15fF
C68026 POR2X1_851/m4_208_n4# GND -0.00fF
C68027 POR2X1_834/Y GND 0.82fF
C68028 POR2X1_840/m4_208_n4# GND 0.00fF
C68029 POR2X1_328/m4_208_n4# GND -0.00fF
C68030 POR2X1_332/Y GND -0.21fF
C68031 POR2X1_339/CTRL GND 0.02fF
C68032 POR2X1_306/CTRL GND 0.02fF
C68033 POR2X1_510/A GND -0.18fF
C68034 POR2X1_509/A GND 0.15fF
C68035 POR2X1_509/m4_208_n4# GND -0.00fF
C68036 POR2X1_509/O GND 0.02fF
C68037 PAND2X1_292/m4_208_n4# GND 0.00fF
C68038 POR2X1_285/B GND 0.30fF
C68039 POR2X1_271/A GND 0.38fF
C68040 POR2X1_486/B GND 0.09fF
C68041 PAND2X1_484/m4_208_n4# GND 0.00fF
C68042 POR2X1_833/A GND 0.50fF
C68043 PAND2X1_495/m4_208_n4# GND 0.00fF
C68044 PAND2X1_472/A GND 0.16fF
C68045 POR2X1_416/Y GND 0.36fF
C68046 PAND2X1_462/m4_208_n4# GND 0.00fF
C68047 PAND2X1_452/B GND 0.22fF
C68048 PAND2X1_216/B GND 0.31fF
C68049 POR2X1_437/Y GND 0.14fF
C68050 PAND2X1_675/A GND 0.40fF
C68051 PAND2X1_440/CTRL2 GND 0.02fF
C68052 INPUT_2 GND 0.19fF
C68053 PAND2X1_8/m4_208_n4# GND 0.00fF
C68054 PAND2X1_687/O GND 0.02fF
C68055 PAND2X1_698/m4_208_n4# GND 0.00fF
C68056 POR2X1_679/B GND 0.20fF
C68057 PAND2X1_676/O GND 0.02fF
C68058 PAND2X1_661/B GND 0.25fF
C68059 PAND2X1_651/Y GND 1.57fF
C68060 PAND2X1_654/m4_208_n4# GND 0.00fF
C68061 PAND2X1_665/m4_208_n4# GND 0.00fF
C68062 POR2X1_616/Y GND 0.19fF
C68063 POR2X1_617/Y GND 0.12fF
C68064 PAND2X1_621/CTRL GND 0.02fF
C68065 POR2X1_855/B GND 0.30fF
C68066 POR2X1_691/B GND 0.17fF
C68067 POR2X1_691/m4_208_n4# GND 0.00fF
C68068 POR2X1_680/Y GND 0.18fF
C68069 POR2X1_680/CTRL GND 0.02fF
C68070 POR2X1_99/B GND 0.59fF
C68071 POR2X1_97/B GND -0.05fF
C68072 POR2X1_97/m4_208_n4# GND 0.00fF
C68073 POR2X1_75/CTRL GND 0.02fF
C68074 POR2X1_22/A GND 0.08fF
C68075 POR2X1_64/m4_208_n4# GND -0.00fF
C68076 POR2X1_64/O GND 0.02fF
C68077 POR2X1_86/Y GND 0.17fF
C68078 POR2X1_85/Y GND -0.33fF
C68079 POR2X1_86/m4_208_n4# GND -0.01fF
C68080 POR2X1_53/m4_208_n4# GND 0.00fF
C68081 POR2X1_31/m4_208_n4# GND 0.00fF
C68082 POR2X1_42/m4_208_n4# GND 0.00fF
C68083 POR2X1_20/Y GND 0.21fF
C68084 POR2X1_20/m4_208_n4# GND 0.00fF
C68085 POR2X1_775/A GND -0.45fF
C68086 PAND2X1_109/m4_208_n4# GND 0.00fF
C68087 POR2X1_179/Y GND 0.19fF
C68088 POR2X1_311/m4_208_n4# GND -0.01fF
C68089 POR2X1_146/Y GND 0.20fF
C68090 POR2X1_146/m4_208_n4# GND -0.00fF
C68091 POR2X1_36/B GND 0.70fF
C68092 POR2X1_3/A GND 0.63fF
C68093 POR2X1_157/m4_208_n4# GND 0.00fF
C68094 POR2X1_170/B GND 0.23fF
C68095 POR2X1_168/A GND 0.19fF
C68096 POR2X1_113/A GND 0.11fF
C68097 POR2X1_123/Y GND -0.14fF
C68098 POR2X1_124/B GND 0.31fF
C68099 POR2X1_124/m4_208_n4# GND 0.00fF
C68100 POR2X1_124/CTRL GND 0.01fF
C68101 PAND2X1_863/B GND 0.44fF
C68102 PAND2X1_857/CTRL2 GND 0.02fF
C68103 POR2X1_821/Y GND -0.24fF
C68104 POR2X1_822/Y GND 0.18fF
C68105 PAND2X1_835/CTRL GND 0.02fF
C68106 PAND2X1_848/A GND 0.19fF
C68107 PAND2X1_809/B GND 0.17fF
C68108 PAND2X1_798/Y GND 0.61fF
C68109 POR2X1_845/A GND 0.13fF
C68110 POR2X1_62/Y GND 0.84fF
C68111 POR2X1_266/A GND 0.61fF
C68112 PAND2X1_813/CTRL GND 0.02fF
C68113 POR2X1_858/B GND 0.25fF
C68114 POR2X1_865/B GND 0.32fF
C68115 POR2X1_861/m4_208_n4# GND 0.00fF
C68116 PAND2X1_63/Y GND 0.77fF
C68117 POR2X1_327/m4_208_n4# GND -0.00fF
C68118 POR2X1_327/CTRL GND 0.01fF
C68119 POR2X1_343/Y GND 1.46fF
C68120 POR2X1_342/Y GND 0.13fF
C68121 POR2X1_349/m4_208_n4# GND -0.01fF
C68122 POR2X1_351/B GND 0.21fF
C68123 POR2X1_334/Y GND 0.84fF
C68124 POR2X1_333/Y GND -0.34fF
C68125 POR2X1_338/m4_208_n4# GND 0.00fF
C68126 POR2X1_305/Y GND 0.33fF
C68127 POR2X1_316/Y GND 0.36fF
C68128 POR2X1_81/A GND 0.74fF
C68129 POR2X1_316/CTRL GND 0.02fF
C68130 POR2X1_519/m4_208_n4# GND 0.00fF
C68131 POR2X1_519/CTRL GND 0.02fF
C68132 POR2X1_510/B GND 0.17fF
C68133 POR2X1_508/m4_208_n4# GND 0.00fF
C68134 POR2X1_334/A GND 0.32fF
C68135 PAND2X1_824/B GND 0.37fF
C68136 POR2X1_542/B GND 0.40fF
C68137 PAND2X1_631/A GND 0.72fF
C68138 POR2X1_252/Y GND -0.18fF
C68139 PAND2X1_483/m4_208_n4# GND 0.00fF
C68140 PAND2X1_462/B GND 0.22fF
C68141 POR2X1_411/Y GND -0.05fF
C68142 POR2X1_413/Y GND 0.12fF
C68143 PAND2X1_461/m4_208_n4# GND 0.00fF
C68144 PAND2X1_476/A GND 0.46fF
C68145 PAND2X1_452/A GND 0.03fF
C68146 PAND2X1_450/m4_208_n4# GND 0.00fF
C68147 PAND2X1_7/O GND 0.02fF
C68148 PAND2X1_687/B GND 0.30fF
C68149 POR2X1_684/Y GND 0.11fF
C68150 PAND2X1_686/m4_208_n4# GND 0.00fF
C68151 POR2X1_383/A GND 1.61fF
C68152 PAND2X1_736/A GND 0.45fF
C68153 PAND2X1_649/A GND 0.37fF
C68154 PAND2X1_642/m4_208_n4# GND 0.00fF
C68155 PAND2X1_642/CTRL2 GND 0.02fF
C68156 PAND2X1_664/m4_208_n4# GND 0.00fF
C68157 POR2X1_594/Y GND 0.05fF
C68158 PAND2X1_652/Y GND 0.04fF
C68159 POR2X1_613/Y GND 0.08fF
C68160 PAND2X1_620/m4_208_n4# GND 0.00fF
C68161 PAND2X1_632/B GND 0.28fF
C68162 PAND2X1_631/m4_208_n4# GND 0.00fF
C68163 POR2X1_690/Y GND 0.17fF
C68164 POR2X1_413/A GND 0.61fF
C68165 POR2X1_74/Y GND 0.19fF
C68166 POR2X1_85/m4_208_n4# GND -0.01fF
C68167 POR2X1_96/Y GND 0.35fF
C68168 POR2X1_51/B GND 0.74fF
C68169 POR2X1_30/m4_208_n4# GND 0.00fF
C68170 POR2X1_41/Y GND 0.21fF
C68171 POR2X1_41/m4_208_n4# GND 0.00fF
C68172 POR2X1_41/CTRL2 GND 0.02fF
C68173 INPUT_1 GND -6.56fF
C68174 PAND2X1_94/A GND 1.68fF
C68175 PAND2X1_119/m4_208_n4# GND 0.00fF
C68176 POR2X1_114/B GND 0.29fF
C68177 PAND2X1_108/m4_208_n4# GND 0.00fF
C68178 POR2X1_178/Y GND 0.37fF
C68179 POR2X1_178/CTRL GND 0.02fF
C68180 POR2X1_189/Y GND 0.31fF
C68181 POR2X1_189/m4_208_n4# GND 0.00fF
C68182 POR2X1_167/CTRL GND 0.02fF
C68183 POR2X1_145/Y GND 0.33fF
C68184 POR2X1_145/m4_208_n4# GND -0.00fF
C68185 POR2X1_145/CTRL GND 0.02fF
C68186 POR2X1_155/Y GND 0.13fF
C68187 POR2X1_134/CTRL GND 0.02fF
C68188 POR2X1_123/m4_208_n4# GND 0.00fF
C68189 POR2X1_123/CTRL GND 0.01fF
C68190 POR2X1_332/B GND -0.47fF
C68191 PAND2X1_863/A GND 0.27fF
C68192 PAND2X1_854/Y GND 0.18fF
C68193 PAND2X1_849/B GND 0.31fF
C68194 POR2X1_813/Y GND 0.20fF
C68195 PAND2X1_845/CTRL GND 0.02fF
C68196 PAND2X1_840/B GND 0.18fF
C68197 PAND2X1_834/m4_208_n4# GND 0.00fF
C68198 PAND2X1_823/CTRL GND 0.02fF
C68199 GATE_811 GND 0.17fF
C68200 PAND2X1_811/Y GND 0.24fF
C68201 PAND2X1_811/m4_208_n4# GND -0.01fF
C68202 PAND2X1_809/A GND 0.26fF
C68203 POR2X1_861/A GND 0.60fF
C68204 POR2X1_860/m4_208_n4# GND 0.00fF
C68205 POR2X1_335/Y GND -0.24fF
C68206 POR2X1_337/m4_208_n4# GND -0.00fF
C68207 POR2X1_337/CTRL2 GND 0.02fF
C68208 POR2X1_349/Y GND -0.25fF
C68209 POR2X1_359/B GND 0.05fF
C68210 POR2X1_344/Y GND 0.12fF
C68211 POR2X1_348/CTRL GND 0.02fF
C68212 POR2X1_56/B GND 0.54fF
C68213 POR2X1_304/CTRL2 GND 0.02fF
C68214 POR2X1_324/Y GND 0.30fF
C68215 POR2X1_324/m4_208_n4# GND -0.01fF
C68216 POR2X1_326/CTRL GND 0.02fF
C68217 POR2X1_315/Y GND 0.58fF
C68218 POR2X1_315/m4_208_n4# GND 0.00fF
C68219 POR2X1_529/Y GND 0.34fF
C68220 D_INPUT_3 GND 0.59fF
C68221 POR2X1_529/m4_208_n4# GND 0.00fF
C68222 POR2X1_518/m4_208_n4# GND 0.00fF
C68223 POR2X1_508/A GND 0.10fF
C68224 POR2X1_507/B GND 0.17fF
C68225 POR2X1_507/O GND 0.02fF
C68226 POR2X1_334/B GND 2.03fF
C68227 PAND2X1_290/m4_208_n4# GND 0.00fF
C68228 POR2X1_491/Y GND 0.23fF
C68229 POR2X1_492/Y GND 0.18fF
C68230 PAND2X1_493/CTRL2 GND 0.02fF
C68231 POR2X1_409/Y GND 0.11fF
C68232 PAND2X1_460/m4_208_n4# GND 0.00fF
C68233 PAND2X1_477/B GND 0.30fF
C68234 PAND2X1_464/Y GND -0.08fF
C68235 POR2X1_237/m4_208_n4# GND -0.01fF
C68236 POR2X1_483/A GND 0.29fF
C68237 PAND2X1_482/m4_208_n4# GND 0.00fF
C68238 PAND2X1_687/A GND 0.17fF
C68239 POR2X1_708/B GND 0.21fF
C68240 POR2X1_502/A GND 1.72fF
C68241 GATE_662 GND 0.04fF
C68242 PAND2X1_659/Y GND 0.82fF
C68243 PAND2X1_662/Y GND 0.16fF
C68244 PAND2X1_663/m4_208_n4# GND 0.00fF
C68245 PAND2X1_674/CTRL2 GND 0.01fF
C68246 POR2X1_594/m4_208_n4# GND -0.01fF
C68247 PAND2X1_341/B GND 0.51fF
C68248 POR2X1_265/Y GND 0.40fF
C68249 PAND2X1_632/A GND 0.25fF
C68250 PAND2X1_630/m4_208_n4# GND 0.00fF
C68251 POR2X1_96/A GND 1.01fF
C68252 POR2X1_51/A GND 0.13fF
C68253 POR2X1_95/CTRL GND 0.02fF
C68254 POR2X1_73/m4_208_n4# GND 0.00fF
C68255 POR2X1_73/CTRL2 GND 0.02fF
C68256 POR2X1_84/m4_208_n4# GND 0.00fF
C68257 POR2X1_84/CTRL GND 0.02fF
C68258 POR2X1_51/m4_208_n4# GND 0.00fF
C68259 POR2X1_25/Y GND 0.48fF
C68260 POR2X1_40/m4_208_n4# GND 0.00fF
C68261 POR2X1_62/CTRL2 GND 0.02fF
C68262 PAND2X1_90/A GND 1.17fF
C68263 PAND2X1_129/m4_208_n4# GND 0.00fF
C68264 POR2X1_123/A GND -0.49fF
C68265 POR2X1_733/m4_208_n4# GND -0.01fF
C68266 POR2X1_207/B GND 0.19fF
C68267 POR2X1_196/Y GND 0.22fF
C68268 POR2X1_199/CTRL GND 0.02fF
C68269 POR2X1_177/Y GND 0.27fF
C68270 POR2X1_16/A GND 0.87fF
C68271 POR2X1_166/CTRL2 GND 0.02fF
C68272 POR2X1_407/A GND 0.73fF
C68273 POR2X1_68/A GND 1.71fF
C68274 POR2X1_144/Y GND 0.19fF
C68275 POR2X1_144/CTRL GND 0.02fF
C68276 POR2X1_111/Y GND 0.27fF
C68277 POR2X1_111/CTRL GND 0.02fF
C68278 POR2X1_133/m4_208_n4# GND 0.00fF
C68279 POR2X1_122/Y GND 0.19fF
C68280 POR2X1_122/A GND 0.13fF
C68281 POR2X1_122/m4_208_n4# GND -0.00fF
C68282 POR2X1_101/A GND 0.23fF
C68283 PAND2X1_86/Y GND 0.17fF
C68284 GATE_865 GND 0.17fF
C68285 PAND2X1_865/Y GND 0.84fF
C68286 PAND2X1_856/B GND 0.35fF
C68287 PAND2X1_691/Y GND 0.68fF
C68288 PAND2X1_840/A GND 0.33fF
C68289 POR2X1_495/Y GND -0.18fF
C68290 PAND2X1_351/m4_208_n4# GND -0.00fF
C68291 PAND2X1_808/Y GND 0.24fF
C68292 PAND2X1_801/B GND 0.20fF
C68293 POR2X1_760/Y GND 0.29fF
C68294 POR2X1_760/m4_208_n4# GND -0.01fF
C68295 POR2X1_369/Y GND 0.10fF
C68296 POR2X1_119/Y GND 1.51fF
C68297 POR2X1_369/m4_208_n4# GND 0.00fF
C68298 POR2X1_337/A GND 0.22fF
C68299 POR2X1_538/A GND 0.10fF
C68300 POR2X1_336/m4_208_n4# GND -0.00fF
C68301 POR2X1_364/A GND 0.35fF
C68302 POR2X1_351/Y GND 0.26fF
C68303 POR2X1_350/Y GND 0.14fF
C68304 POR2X1_333/m4_208_n4# GND -0.01fF
C68305 POR2X1_360/A GND 0.41fF
C68306 POR2X1_347/B GND -1.18fF
C68307 POR2X1_347/m4_208_n4# GND 0.00fF
C68308 POR2X1_326/A GND -1.05fF
C68309 POR2X1_325/m4_208_n4# GND 0.00fF
C68310 POR2X1_566/A GND 2.10fF
C68311 POR2X1_302/Y GND 0.58fF
C68312 POR2X1_303/m4_208_n4# GND 0.00fF
C68313 POR2X1_567/A GND 0.40fF
C68314 POR2X1_537/Y GND -0.87fF
C68315 POR2X1_528/Y GND 0.41fF
C68316 POR2X1_528/O GND 0.02fF
C68317 POR2X1_517/Y GND 0.18fF
C68318 POR2X1_517/m4_208_n4# GND 0.00fF
C68319 POR2X1_508/B GND 0.53fF
C68320 POR2X1_447/B GND 0.90fF
C68321 POR2X1_506/m4_208_n4# GND 0.00fF
C68322 POR2X1_711/B GND -0.17fF
C68323 POR2X1_709/B GND 0.25fF
C68324 POR2X1_709/m4_208_n4# GND 0.00fF
C68325 POR2X1_555/A GND -0.99fF
C68326 PAND2X1_477/A GND 0.20fF
C68327 PAND2X1_467/Y GND 0.25fF
C68328 PAND2X1_470/CTRL2 GND 0.02fF
C68329 PAND2X1_5/m4_208_n4# GND -0.00fF
C68330 PAND2X1_23/Y GND 2.37fF
C68331 PAND2X1_48/B GND 1.67fF
C68332 POR2X1_686/A GND 0.43fF
C68333 PAND2X1_684/O GND 0.02fF
C68334 PAND2X1_660/Y GND 0.16fF
C68335 PAND2X1_661/Y GND 0.49fF
C68336 PAND2X1_662/m4_208_n4# GND 0.00fF
C68337 POR2X1_670/Y GND 0.15fF
C68338 PAND2X1_639/Y GND -0.27fF
C68339 PAND2X1_651/m4_208_n4# GND 0.00fF
C68340 PAND2X1_651/O GND 0.02fF
C68341 PAND2X1_650/A GND 0.26fF
C68342 PAND2X1_633/Y GND -0.10fF
C68343 PAND2X1_640/m4_208_n4# GND 0.00fF
C68344 POR2X1_72/Y GND 0.28fF
C68345 POR2X1_71/Y GND 0.44fF
C68346 POR2X1_83/Y GND -0.66fF
C68347 POR2X1_83/m4_208_n4# GND 0.00fF
C68348 POR2X1_96/B GND 0.20fF
C68349 POR2X1_50/m4_208_n4# GND 0.00fF
C68350 POR2X1_61/A GND 0.16fF
C68351 POR2X1_61/m4_208_n4# GND 0.00fF
C68352 PAND2X1_140/A GND 0.15fF
C68353 PAND2X1_128/m4_208_n4# GND 0.00fF
C68354 PAND2X1_137/Y GND 0.42fF
C68355 PAND2X1_106/m4_208_n4# GND 0.00fF
C68356 POR2X1_123/B GND 0.19fF
C68357 PAND2X1_117/m4_208_n4# GND 0.00fF
C68358 PAND2X1_117/CTRL GND 0.01fF
C68359 POR2X1_187/Y GND 0.21fF
C68360 POR2X1_208/A GND 0.46fF
C68361 POR2X1_197/Y GND 0.25fF
C68362 POR2X1_176/m4_208_n4# GND 0.00fF
C68363 POR2X1_165/Y GND 0.17fF
C68364 POR2X1_156/B GND -0.26fF
C68365 PAND2X1_6/Y GND 1.77fF
C68366 POR2X1_121/m4_208_n4# GND -0.00fF
C68367 POR2X1_143/m4_208_n4# GND 0.00fF
C68368 POR2X1_110/m4_208_n4# GND 0.00fF
C68369 PAND2X1_535/Y GND 0.31fF
C68370 POR2X1_251/Y GND 0.29fF
C68371 POR2X1_278/Y GND 0.98fF
C68372 PAND2X1_843/m4_208_n4# GND 0.00fF
C68373 PAND2X1_862/Y GND 0.08fF
C68374 PAND2X1_821/m4_208_n4# GND 0.00fF
C68375 PAND2X1_841/B GND 0.18fF
C68376 PAND2X1_832/O GND 0.02fF
C68377 PAND2X1_812/A GND 0.37fF
C68378 POR2X1_335/B GND -0.13fF
C68379 PAND2X1_309/m4_208_n4# GND 0.00fF
C68380 POR2X1_379/Y GND 0.19fF
C68381 POR2X1_379/m4_208_n4# GND 0.00fF
C68382 POR2X1_368/Y GND 0.11fF
C68383 POR2X1_368/m4_208_n4# GND 0.00fF
C68384 POR2X1_353/Y GND 0.27fF
C68385 POR2X1_357/CTRL GND 0.02fF
C68386 POR2X1_347/A GND 0.48fF
C68387 POR2X1_346/B GND 0.42fF
C68388 POR2X1_346/m4_208_n4# GND 0.00fF
C68389 POR2X1_346/CTRL GND 0.02fF
C68390 POR2X1_302/A GND 0.13fF
C68391 POR2X1_302/m4_208_n4# GND 0.00fF
C68392 POR2X1_302/CTRL GND 0.01fF
C68393 POR2X1_324/A GND 0.19fF
C68394 POR2X1_324/B GND 0.15fF
C68395 POR2X1_324/CTRL GND 0.02fF
C68396 POR2X1_313/Y GND -0.00fF
C68397 POR2X1_335/A GND -0.12fF
C68398 POR2X1_335/m4_208_n4# GND 0.00fF
C68399 POR2X1_110/Y GND 0.55fF
C68400 POR2X1_527/m4_208_n4# GND 0.00fF
C68401 POR2X1_539/A GND 0.31fF
C68402 POR2X1_538/m4_208_n4# GND 0.00fF
C68403 POR2X1_565/B GND -0.43fF
C68404 POR2X1_549/m4_208_n4# GND 0.00fF
C68405 POR2X1_505/Y GND 0.22fF
C68406 POR2X1_516/A GND 0.13fF
C68407 POR2X1_722/A GND 0.32fF
C68408 POR2X1_719/B GND -0.19fF
C68409 POR2X1_712/A GND -0.05fF
C68410 POR2X1_779/A GND 0.39fF
C68411 POR2X1_708/CTRL2 GND 0.02fF
C68412 GATE_479 GND 0.12fF
C68413 PAND2X1_478/Y GND 0.20fF
C68414 PAND2X1_776/m4_208_n4# GND -0.01fF
C68415 POR2X1_493/B GND -0.24fF
C68416 PAND2X1_4/m4_208_n4# GND -0.00fF
C68417 POR2X1_614/A GND -10.13fF
C68418 PAND2X1_694/m4_208_n4# GND 0.00fF
C68419 POR2X1_673/A GND 0.21fF
C68420 PAND2X1_671/Y GND -0.19fF
C68421 PAND2X1_672/CTRL GND 0.02fF
C68422 PAND2X1_654/A GND 0.20fF
C68423 PAND2X1_641/Y GND -0.16fF
C68424 PAND2X1_650/m4_208_n4# GND 0.00fF
C68425 PAND2X1_653/Y GND 0.04fF
C68426 PAND2X1_661/m4_208_n4# GND 0.00fF
C68427 POR2X1_686/B GND 0.08fF
C68428 POR2X1_78/B GND 2.00fF
C68429 PAND2X1_683/CTRL GND 0.02fF
C68430 POR2X1_93/O GND 0.02fF
C68431 POR2X1_83/A GND -0.44fF
C68432 POR2X1_82/m4_208_n4# GND 0.00fF
C68433 POR2X1_71/m4_208_n4# GND -0.01fF
C68434 PAND2X1_209/A GND -0.30fF
C68435 PAND2X1_148/Y GND 0.03fF
C68436 PAND2X1_149/m4_208_n4# GND 0.00fF
C68437 PAND2X1_139/B GND 0.43fF
C68438 POR2X1_135/Y GND 0.28fF
C68439 PAND2X1_114/Y GND 0.20fF
C68440 PAND2X1_115/Y GND 0.23fF
C68441 PAND2X1_116/m4_208_n4# GND 0.00fF
C68442 POR2X1_128/A GND 0.30fF
C68443 PAND2X1_127/O GND 0.02fF
C68444 PAND2X1_56/Y GND 2.18fF
C68445 POR2X1_197/CTRL GND 0.02fF
C68446 POR2X1_188/A GND 0.36fF
C68447 POR2X1_186/m4_208_n4# GND 0.00fF
C68448 POR2X1_164/Y GND 0.47fF
C68449 POR2X1_853/A GND 0.61fF
C68450 POR2X1_175/m4_208_n4# GND 0.00fF
C68451 POR2X1_153/CTRL GND 0.02fF
C68452 POR2X1_131/Y GND 0.20fF
C68453 POR2X1_131/m4_208_n4# GND -0.01fF
C68454 POR2X1_121/A GND -0.77fF
C68455 POR2X1_120/m4_208_n4# GND 0.00fF
C68456 POR2X1_65/A GND 1.80fF
C68457 POR2X1_49/Y GND 1.47fF
C68458 POR2X1_142/CTRL GND 0.02fF
C68459 PAND2X1_830/Y GND 0.16fF
C68460 PAND2X1_842/CTRL GND 0.02fF
C68461 PAND2X1_866/A GND 0.19fF
C68462 PAND2X1_810/A GND 0.05fF
C68463 PAND2X1_857/B GND 0.21fF
C68464 PAND2X1_853/CTRL2 GND 0.02fF
C68465 POR2X1_847/A GND 0.21fF
C68466 PAND2X1_820/CTRL2 GND 0.02fF
C68467 PAND2X1_317/Y GND 0.56fF
C68468 PAND2X1_319/m4_208_n4# GND -0.00fF
C68469 POR2X1_306/Y GND 0.40fF
C68470 PAND2X1_308/CTRL GND 0.02fF
C68471 POR2X1_389/A GND -0.49fF
C68472 POR2X1_389/m4_208_n4# GND 0.00fF
C68473 POR2X1_378/Y GND 0.18fF
C68474 POR2X1_378/m4_208_n4# GND 0.00fF
C68475 D_GATE_366 GND 0.26fF
C68476 POR2X1_366/Y GND 0.45fF
C68477 POR2X1_365/Y GND 0.20fF
C68478 POR2X1_348/A GND 0.24fF
C68479 POR2X1_345/A GND 0.17fF
C68480 POR2X1_345/CTRL GND 0.02fF
C68481 POR2X1_312/m4_208_n4# GND -0.00fF
C68482 POR2X1_323/Y GND 0.19fF
C68483 POR2X1_164/m4_208_n4# GND -0.01fF
C68484 POR2X1_537/m4_208_n4# GND 0.00fF
C68485 POR2X1_559/B GND 0.18fF
C68486 POR2X1_549/A GND 0.17fF
C68487 POR2X1_548/B GND 0.08fF
C68488 POR2X1_504/Y GND -0.03fF
C68489 POR2X1_504/m4_208_n4# GND 0.00fF
C68490 POR2X1_526/m4_208_n4# GND -0.01fF
C68491 POR2X1_526/CTRL GND 0.02fF
C68492 POR2X1_514/Y GND 0.21fF
C68493 POR2X1_687/Y GND 0.30fF
C68494 POR2X1_729/m4_208_n4# GND 0.00fF
C68495 POR2X1_729/CTRL GND 0.01fF
C68496 POR2X1_722/B GND 0.22fF
C68497 POR2X1_718/m4_208_n4# GND 0.00fF
C68498 POR2X1_707/A GND 0.06fF
C68499 POR2X1_707/B GND 0.17fF
C68500 POR2X1_557/A GND 0.53fF
C68501 PAND2X1_63/m4_208_n4# GND -0.01fF
C68502 POR2X1_66/B GND 1.33fF
C68503 PAND2X1_3/CTRL2 GND 0.02fF
C68504 PAND2X1_693/m4_208_n4# GND 0.00fF
C68505 PAND2X1_655/Y GND 0.24fF
C68506 PAND2X1_671/CTRL GND 0.02fF
C68507 POR2X1_685/A GND 0.38fF
C68508 PAND2X1_682/m4_208_n4# GND 0.00fF
C68509 POR2X1_81/m4_208_n4# GND 0.00fF
C68510 POR2X1_8/Y GND -0.40fF
C68511 POR2X1_92/m4_208_n4# GND -0.00fF
C68512 POR2X1_70/m4_208_n4# GND 0.00fF
C68513 PAND2X1_159/O GND 0.02fF
C68514 POR2X1_132/Y GND 0.17fF
C68515 POR2X1_134/Y GND 0.41fF
C68516 PAND2X1_104/m4_208_n4# GND 0.00fF
C68517 PAND2X1_104/CTRL2 GND 0.02fF
C68518 PAND2X1_126/CTRL GND 0.02fF
C68519 PAND2X1_115/m4_208_n4# GND 0.00fF
C68520 PAND2X1_48/Y GND 0.06fF
C68521 POR2X1_702/B GND 0.10fF
C68522 POR2X1_196/CTRL GND 0.02fF
C68523 POR2X1_163/A GND 0.35fF
C68524 POR2X1_52/A GND 1.19fF
C68525 POR2X1_175/A GND 0.17fF
C68526 POR2X1_174/m4_208_n4# GND 0.00fF
C68527 POR2X1_174/CTRL GND 0.02fF
C68528 POR2X1_152/m4_208_n4# GND -0.00fF
C68529 POR2X1_139/Y GND 0.13fF
C68530 POR2X1_141/m4_208_n4# GND -0.01fF
C68531 PAND2X1_857/A GND 0.55fF
C68532 POR2X1_821/m4_208_n4# GND -0.00fF
C68533 PAND2X1_852/CTRL GND 0.02fF
C68534 PAND2X1_864/B GND 0.47fF
C68535 PAND2X1_863/O GND 0.02fF
C68536 PAND2X1_830/O GND 0.02fF
C68537 PAND2X1_831/Y GND -0.11fF
C68538 PAND2X1_841/m4_208_n4# GND 0.00fF
C68539 POR2X1_327/Y GND 0.72fF
C68540 PAND2X1_319/B GND 0.65fF
C68541 PAND2X1_318/m4_208_n4# GND 0.00fF
C68542 PAND2X1_308/B GND 0.21fF
C68543 POR2X1_304/Y GND 0.23fF
C68544 PAND2X1_307/CTRL2 GND 0.02fF
C68545 POR2X1_390/B GND 0.49fF
C68546 POR2X1_180/B GND 0.51fF
C68547 POR2X1_388/m4_208_n4# GND 0.00fF
C68548 POR2X1_399/A GND 0.16fF
C68549 POR2X1_362/Y GND 0.22fF
C68550 POR2X1_378/A GND 0.19fF
C68551 POR2X1_377/m4_208_n4# GND 0.00fF
C68552 POR2X1_356/A GND 2.93fF
C68553 POR2X1_355/B GND 0.43fF
C68554 POR2X1_355/m4_208_n4# GND 0.00fF
C68555 POR2X1_311/Y GND 0.43fF
C68556 POR2X1_322/Y GND 0.22fF
C68557 POR2X1_57/A GND 0.79fF
C68558 POR2X1_322/CTRL GND 0.02fF
C68559 POR2X1_344/A GND 0.21fF
C68560 POR2X1_254/Y GND 0.26fF
C68561 POR2X1_333/A GND 1.10fF
C68562 POR2X1_174/B GND 0.40fF
C68563 POR2X1_558/A GND 0.17fF
C68564 POR2X1_564/Y GND 0.27fF
C68565 POR2X1_536/Y GND -0.19fF
C68566 POR2X1_536/CTRL GND 0.02fF
C68567 POR2X1_550/A GND 0.42fF
C68568 POR2X1_547/m4_208_n4# GND 0.00fF
C68569 POR2X1_547/CTRL GND 0.02fF
C68570 POR2X1_525/Y GND -0.01fF
C68571 POR2X1_41/B GND 1.96fF
C68572 POR2X1_740/A GND 0.16fF
C68573 POR2X1_730/Y GND 0.34fF
C68574 POR2X1_739/m4_208_n4# GND 0.00fF
C68575 POR2X1_730/B GND -0.51fF
C68576 POR2X1_728/m4_208_n4# GND 0.00fF
C68577 POR2X1_728/O GND 0.02fF
C68578 POR2X1_713/A GND 0.15fF
C68579 POR2X1_706/A GND 0.14fF
C68580 POR2X1_706/B GND 0.28fF
C68581 POR2X1_706/m4_208_n4# GND 0.00fF
C68582 POR2X1_717/m4_208_n4# GND 0.00fF
.ends

