*** TEST 045 : compensed AND2 structure ***
*
* ngSPICE test for PLS experiments
*
* NAND PLS test - gate area exported directly from Magic VLSI layout
*
* Author: Jan Belohoubek, 09/2020
* jan.belohoubek@fit.cvut.cz
*
* https://users.fit.cvut.cz/~belohja4/
*
*
* **************************************

.include ../models.lib
.include ../tsmc180nmcmos.lib
.include magic/PAND2X1.spice

* **************************************
* --- Test ---
* **************************************

* --- Settings
.param showPlots = 1
.param writeFile = 1
* redefine ...
.include test04X_settings.inc
.csparam showPlots = {showPlots}
.csparam writeFile = {writeFile}
.global showPlots writeFile
* --- End of Settins

Vtrig LaserTrig 0 0 PWL(0ns 0V 40ns 0V 42ns SUPP 62ns SUPP 64ns 0V 100ns 0V)

.param beamDistanceTop = 0
.param beamDistanceBot = 0

.global LaserTrig beamDistanceTop beamDistanceBot

* --- inputs
*Vvin0 A 0 0 PWL(0ns 0V 30ns 0V 31ns SUPP)

* --- outputs
C1 VSS O 10fF

* --- circuit layout model
Xgate VDD VSS B A Y PAND2X1

*Ra Xgate.A A 0.001
*Rb Xgate.B B 0.001
Ro Xgate.O O 0.001
*Ry Xgate.Y Y 0.001
*Rsupply Xgate.VDD VDD 0.001
*Rground Xgate.GND VSS 0.001
Rctrl Xgate.CTRL CTRL 0.001
Rctrl2 Xgate.CTRL2 CTRL2 0.001

* **************************************
* --- Simulation Settings ---
* **************************************

.tran 0.1ns 100ns
.param SIMSTEP = '100ns/0.1ns'
.csparam SIMSTEP = {SIMSTEP}

* **************************************
* --- Simulation Control ---
* **************************************

.control
    let INHIGH_NEW = 'SUPP-0.3V'
    let INLOW_NEW = '0V - 0.3V'
    
    alterparam INHIGH = $&INHIGH_NEW
    alterparam INLOW = $&INLOW_NEW
    reset
    
    run
    
    if ('showPlots' > 0)   
        plot i(vvdd) i(vvss)
        
        plot v(A)
        plot v(O) 
    end
    
    let timeIndex = 0
    while time[timeIndex] < 55ns
      let timeIndex= timeIndex + 1
    end
    
    print i(VVDD)[$&timeIndex]
    print v(O)[$&timeIndex]
    print v(Y)[$&timeIndex]
    print v(CTRL)[$&timeIndex]
    print v(CTRL2)[$&timeIndex]
    print time[$&timeIndex]
    
    if ('writeFile' > 0)   
      wrdata ivdd.out i(vvdd)
      wrdata ivss.out i(vvss)
    end
    
    if ('showPlots' < 1)
        quit
    end
    
.endc

.end
