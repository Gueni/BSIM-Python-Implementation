*** NAND2 gate symetric elements + serial R ***
*
* ngSPICE compensed NAND gate
*
*
* Author: Jan Belohoubek, 01/2020
* jan.belohoubek@fit.cvut.cz
*
* https://users.fit.cvut.cz/~belohja4/
*
*
* **************************************

.subckt NAND2 A B O VSS VDD

*** block P ***
Xpmos1 Y A VDD_TOP VDD_TOP VSS LaserTrig SUBCKT_PMOS beamDistance = beamDistanceTop ch_w=2u ch_l=0.2u mos_ad=0.6p mos_pd=2.6u mos_as=1p mos_ps=5u
Xpmos2 Y B VDD_TOP VDD_TOP VSS LaserTrig SUBCKT_PMOS beamDistance = beamDistanceTop ch_w=2u ch_l=0.2u mos_ad=0.6p mos_pd=2.6u mos_as=1p mos_ps=5u

*** block N ***
Xnmos1 MIDDLE A VSS_BOT VSS psubIn LaserTrig SUBCKT_NMOS beamDistance = beamDistanceBot ch_w=1u ch_l=0.2u mos_ad=0.15p mos_pd=1.7u mos_as=0.5p  mos_ps=2.5u commonDrain = 1 commonSource = 0
Xnmos2 Y B MIDDLE       VSS psubIn LaserTrig SUBCKT_NMOS beamDistance = beamDistanceBot ch_w=1u ch_l=0.2u mos_ad=0.5p  mos_pd=2.5u mos_as=0.15p mos_ps=1.2u commonDrain = 0 commonSource = 1

Xnmos1c MIDDLE2 B VSS_BOT VSS psubIn LaserTrig SUBCKT_NMOS beamDistance = beamDistanceBot ch_w=1u ch_l=0.2u mos_ad=0.15p mos_pd=1.7u mos_as=0.5p  mos_ps=2.5u commonDrain = 1 commonSource = 0
Xnmos2c Y A MIDDLE2       VSS psubIn LaserTrig SUBCKT_NMOS beamDistance = beamDistanceBot ch_w=1u ch_l=0.2u mos_ad=0.5p  mos_pd=2.5u mos_as=0.15p mos_ps=1.2u commonDrain = 0 commonSource = 1

*** Compensation Serial PMOS - TOP ***
XpmosTOP VDD_TOP VSS VDD VDD VSS LaserTrig SUBCKT_PMOS beamDistance = beamDistanceTop ch_w=2u ch_l=0.2u mos_ad=1.1p mos_pd=5u mos_as=1.1p mos_ps=5u

*** Compensation Serial NMOS - BOT ***
Rbot VSS_BOT VSS 0.001

*** Output ***
R1 Y O 1

*** common NMOS substarte virtual node ***
XpsubIn psubIn VSS PSUB_IN

.ends
