* SPICE3 file created from PAND2X1.ext - technology: scmos

*.subckt PAND2X1 VDD GND B A Y a_36_28# O m4_240_n4# a_48_308# a_8_28# CTRL2 CTRL a_88_28#
.subckt PAND2X1 VDD GND B A Y
X0 CTRL GND VDD VDD PMOS_MAGIC ad=0.2p pd=1.8u as=4.78p ps=22.2u w=0.4u l=0.2u
**devattr s=S d=D
X1 O B a_48_308# VDD PMOS_MAGIC ad=1.16p pd=6.2u as=1.76p ps=8.6u w=1.6u l=0.2u
**devattr s=S d=D
X2 CTRL2 CTRL VDD VDD PMOS_MAGIC ad=1.95p pd=8.8u as=0p ps=0u w=3.9u l=0.2u
**devattr s=S d=D
X3 Y O GND GND NMOS_MAGIC ad=0.8p pd=4.2u as=2.83p ps=13.6u w=1.6u l=0.2u
**devattr s=S d=D
X4 O CTRL4 GND GND NMOS_MAGIC ad=0.84p pd=5.4u as=0p ps=0u w=1.2u l=0.2u
**devattr s=S d=D
X5 CTRL2 CTRL GND GND NMOS_MAGIC ad=0.2p pd=1.8u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X6 CTRL GND GND GND NMOS_MAGIC ad=1.75p pd=8u as=0p ps=0u w=3.5u l=0.2u
**devattr s=S d=D
X7 a_48_308# CTRL4 VDD VDD PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=1.6u l=0.2u
**devattr s=S d=D
X8 a_36_28# B a_8_28# GND NMOS_MAGIC ad=0.12p pd=1.4u as=0.84p ps=5.4u w=0.4u l=0.2u
**devattr s=S d=D
X9 a_88_28# A a_8_28# GND NMOS_MAGIC ad=0.12p pd=1.4u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X10 O B a_88_28# GND NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X11 O A a_36_28# GND NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X12 Y O VDD VDD PMOS_MAGIC ad=1.95p pd=8.8u as=0p ps=0u w=3.9u l=0.2u
**devattr s=S d=D
X13 a_8_28# CTRL3 GND GND NMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=1.2u l=0.2u
**devattr s=S d=D
X14 O CTRL3 VDD VDD PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=0.4u l=0.2u
**devattr s=S d=D
X15 O A a_48_308# VDD PMOS_MAGIC ad=0p pd=0u as=0p ps=0u w=1.6u l=0.2u

X22 CTRL4 CTRL3 VDD VDD PMOS_MAGIC ad=1.95p pd=8.8u as=0p ps=0u w=3.9u l=0.2u
X55 CTRL4 CTRL3 GND GND NMOS_MAGIC ad=0.2p pd=1.8u as=0p ps=0u w=0.4u l=0.2u

X00 CTRL3 CTRL2 VDD VDD PMOS_MAGIC ad=0.2p pd=1.8u as=4.78p ps=22.2u w=0.4u l=0.2u
X66 CTRL3 CTRL2 GND GND NMOS_MAGIC ad=1.75p pd=8u as=0p ps=0u w=3.5u l=0.2u


**devattr s=S d=D
C0 CTRL2 VDD 0.73fF
C1 CTRL2 CTRL 0.34fF
C2 CTRL VDD 1.51fF
C3 CTRL2 O 0.90fF
C4 VDD B 0.36fF
C5 a_8_28# a_36_28# 0.00fF
C6 CTRL2 A 0.06fF
C7 O VDD 0.71fF
C8 CTRL O 0.21fF
C9 VDD A 0.22fF
C10 a_8_28# a_88_28# 0.00fF
C11 a_48_308# VDD 0.29fF
C12 CTRL A 0.13fF
C13 O B 0.04fF
C14 VDD Y 0.54fF
C15 B A 0.82fF
C16 O A 0.12fF
C17 a_48_308# B 0.01fF
C18 O a_48_308# 0.41fF
C19 O Y 0.05fF
C20 a_48_308# A 0.01fF
C21 a_8_28# B 0.01fF
C22 O a_8_28# 0.08fF
C23 a_8_28# A 0.01fF
C24 Y GND 0.50fF
C25 A GND 0.60fF
C26 B GND 0.55fF
C27 VDD GND 4.94fF
C28 GND GND -0.17fF

*C29 m4_240_n4# GND 0.01fF
Rcorr m4_240_n4# GND 0.001

C30 a_8_28# GND 0.26fF
C31 a_48_308# GND 0.00fF
C32 O GND 0.49fF
C33 CTRL GND 0.65fF
C34 CTRL2 GND 0.44fF
.ends
