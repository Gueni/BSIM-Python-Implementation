magic
tech scmos
magscale 1 2
timestamp 1598358390
<< error_s >>
rect 188 3956 196 3964
rect 140 3876 148 3884
rect 5324 3876 5332 3884
rect 5388 3876 5396 3884
rect 252 3836 256 3844
rect 5340 3776 5348 3784
rect 5452 3756 5460 3764
rect 5516 3756 5524 3764
rect 5312 3696 5316 3704
rect 5388 3696 5396 3704
rect 5436 3696 5444 3704
rect 5516 3696 5524 3704
rect 5452 3536 5460 3544
rect 5324 3516 5332 3524
rect 5388 3516 5396 3524
rect 5532 3516 5540 3524
rect 5436 3496 5444 3504
rect 28 3476 36 3484
rect 204 3476 212 3484
rect 5324 3476 5332 3484
rect 252 3456 256 3464
rect 124 3356 132 3364
rect 252 3356 256 3364
rect 5388 3336 5396 3344
rect 5324 3316 5332 3324
rect 60 3296 68 3304
rect 5532 3296 5540 3304
rect 76 3196 84 3204
rect 5312 3156 5316 3164
rect 5564 3156 5572 3164
rect 5532 3116 5540 3124
rect 252 3076 256 3084
rect 188 3056 196 3064
rect 204 3056 212 3064
rect 5372 2996 5380 3004
rect 5372 2976 5380 2984
rect 12 2896 20 2904
rect 28 2896 36 2904
rect 76 2896 84 2904
rect 156 2716 164 2724
rect 5452 2716 5460 2724
rect 5516 2716 5524 2724
rect 5372 2696 5380 2704
rect 5484 2696 5492 2704
rect 92 2676 100 2684
rect 60 2556 68 2564
rect 124 2536 132 2544
rect 172 2536 180 2544
rect 5388 2536 5396 2544
rect 5452 2536 5460 2544
rect 5516 2536 5524 2544
rect 5372 2496 5380 2504
rect 252 2396 260 2404
rect 5324 2316 5332 2324
rect 5468 2316 5476 2324
rect 140 2276 148 2284
rect 204 2276 212 2284
rect 76 2256 84 2264
rect 5564 2176 5572 2184
rect 108 2136 116 2144
rect 172 2136 180 2144
rect 5372 2136 5380 2144
rect 5452 2136 5460 2144
rect 5484 2136 5492 2144
rect 5516 2136 5524 2144
rect 12 2096 20 2104
rect 236 2096 244 2104
rect 5516 2096 5524 2104
rect 5372 1916 5380 1924
rect 5468 1916 5476 1924
rect 140 1896 148 1904
rect 172 1876 180 1884
rect 204 1876 212 1884
rect 5404 1876 5412 1884
rect 140 1776 148 1784
rect 5500 1756 5508 1764
rect 124 1736 132 1744
rect 204 1716 212 1724
rect 5324 1516 5332 1524
rect 5372 1516 5380 1524
rect 5452 1516 5460 1524
rect 172 1476 180 1484
rect 188 1476 196 1484
rect 60 1456 68 1464
rect 188 1456 196 1464
rect 5312 1436 5316 1444
rect 5356 1376 5364 1384
rect 5372 1376 5380 1384
rect 5452 1376 5460 1384
rect 220 1336 228 1344
rect 5500 1336 5508 1344
rect 5484 1296 5492 1304
rect 252 1156 260 1164
rect 5312 1136 5316 1144
rect 5436 1096 5444 1104
rect 28 1076 36 1084
rect 5468 1076 5476 1084
rect 60 1036 68 1044
rect 5388 976 5396 984
rect 5452 976 5460 984
rect 252 956 260 964
rect 5500 936 5508 944
rect 5312 896 5316 904
rect 5356 896 5364 904
rect 5484 896 5492 904
rect 5500 736 5508 744
rect 188 716 196 724
rect 204 696 212 704
rect 5388 696 5396 704
rect 5452 696 5460 704
rect 188 676 196 684
rect 252 676 260 684
rect 5312 676 5316 684
rect 124 656 132 664
rect 124 536 132 544
rect 5404 536 5412 544
rect 5324 516 5332 524
rect 5452 516 5460 524
rect 12 496 20 504
rect 108 496 116 504
rect 236 496 244 504
rect 5452 496 5460 504
rect 5436 436 5444 444
rect 5372 356 5380 364
rect 5388 336 5396 344
rect 28 316 36 324
rect 140 316 148 324
rect 220 276 228 284
rect 5324 276 5332 284
rect 124 236 132 244
rect 5312 176 5316 184
rect 5580 176 5588 184
rect 5324 156 5332 164
rect 44 136 52 144
rect 220 136 228 144
rect 140 116 148 124
rect 5404 96 5412 104
<< metal1 >>
rect -412 4016 -312 4020
rect -412 4004 10 4016
rect -412 3616 -312 4004
rect 1860 3937 1875 3943
rect 125 3917 163 3923
rect 1837 3917 1852 3923
rect 1924 3917 1939 3923
rect 2164 3917 2211 3923
rect 3325 3917 3363 3923
rect 3581 3917 3596 3923
rect 4029 3917 4044 3923
rect 4605 3917 4620 3923
rect 4797 3917 4835 3923
rect 5012 3917 5027 3923
rect 5181 3917 5196 3923
rect 5373 3917 5411 3923
rect 1900 3904 1908 3916
rect 3548 3904 3556 3916
rect 4764 3904 4772 3916
rect 3517 3897 3540 3903
rect 3340 3892 3348 3896
rect 3532 3892 3540 3897
rect 3836 3897 3859 3903
rect 4029 3897 4052 3903
rect 3836 3892 3844 3897
rect 4044 3892 4052 3897
rect 4236 3892 4244 3896
rect 4412 3897 4435 3903
rect 4412 3892 4420 3897
rect 5340 3904 5348 3916
rect 4989 3897 5012 3903
rect 5004 3892 5012 3897
rect 62 3877 83 3883
rect 77 3857 83 3877
rect 317 3877 338 3883
rect 317 3857 323 3877
rect 446 3877 483 3883
rect 557 3877 594 3883
rect 637 3877 658 3883
rect 637 3857 643 3877
rect 708 3877 722 3883
rect 1085 3877 1106 3883
rect 1085 3857 1091 3877
rect 1261 3877 1298 3883
rect 1348 3877 1362 3883
rect 1389 3877 1404 3883
rect 2301 3877 2332 3883
rect 2580 3877 2588 3883
rect 2622 3877 2643 3883
rect 2637 3857 2643 3877
rect 2942 3877 2956 3883
rect 3892 3877 3939 3883
rect 956 3844 964 3848
rect 1164 3844 1172 3848
rect 1468 3844 1476 3848
rect 1548 3844 1556 3848
rect 1676 3844 1684 3848
rect 2044 3844 2052 3848
rect 2060 3844 2068 3848
rect 2124 3844 2132 3848
rect 2236 3844 2244 3848
rect 2252 3844 2260 3848
rect 4092 3844 4100 3848
rect 4220 3844 4228 3848
rect 4284 3844 4292 3848
rect 4364 3844 4372 3848
rect 4668 3844 4676 3848
rect 4860 3844 4868 3848
rect 5052 3844 5060 3848
rect 5244 3844 5252 3848
rect 5260 3844 5268 3848
rect 5436 3844 5444 3848
rect 5500 3843 5508 3848
rect 5500 3837 5516 3843
rect 5894 3816 5994 4018
rect 5552 3804 5994 3816
rect 780 3772 788 3776
rect 844 3772 852 3776
rect 1036 3772 1044 3776
rect 1100 3772 1108 3776
rect 1228 3772 1236 3776
rect 1292 3772 1300 3776
rect 1356 3772 1364 3776
rect 1484 3772 1492 3776
rect 1724 3772 1732 3776
rect 1788 3772 1796 3776
rect 1804 3772 1812 3776
rect 2316 3772 2324 3776
rect 3468 3772 3476 3776
rect 4156 3772 4164 3776
rect 4412 3772 4420 3776
rect 4476 3772 4484 3776
rect 4668 3772 4676 3776
rect 4876 3772 4884 3776
rect 5132 3772 5140 3776
rect 84 3737 99 3743
rect 148 3737 163 3743
rect 237 3737 252 3743
rect 429 3737 466 3743
rect 685 3737 722 3743
rect 1933 3743 1939 3763
rect 2884 3757 2899 3763
rect 4733 3744 4739 3763
rect 1918 3737 1939 3743
rect 2052 3737 2067 3743
rect 4052 3737 4067 3743
rect 4180 3737 4195 3743
rect 4756 3737 4764 3743
rect 5460 3737 5475 3743
rect 316 3724 324 3728
rect 2492 3724 2500 3728
rect 2500 3717 2515 3723
rect 3516 3723 3524 3728
rect 3916 3724 3924 3728
rect 3516 3717 3539 3723
rect 4108 3723 4116 3728
rect 4364 3723 4372 3728
rect 4556 3723 4564 3728
rect 4093 3717 4116 3723
rect 4349 3717 4372 3723
rect 4541 3717 4564 3723
rect 4620 3724 4628 3728
rect 4860 3724 4868 3728
rect 4924 3724 4932 3728
rect 5004 3723 5012 3728
rect 4989 3717 5012 3723
rect 5388 3723 5396 3728
rect 5516 3723 5524 3728
rect 5373 3717 5396 3723
rect 5501 3717 5524 3723
rect 4908 3704 4916 3716
rect 5164 3704 5172 3716
rect 1156 3697 1171 3703
rect 1684 3697 1699 3703
rect 2157 3697 2172 3703
rect 2413 3697 2428 3703
rect 3309 3697 3324 3703
rect 3501 3697 3516 3703
rect 3901 3697 3939 3703
rect 4564 3697 4579 3703
rect 5396 3697 5411 3703
rect 5524 3697 5539 3703
rect 2237 3677 2252 3683
rect 2436 3677 2451 3683
rect 4349 3677 4364 3683
rect 5565 3637 5580 3643
rect -412 3604 16 3616
rect -412 3216 -312 3604
rect 4221 3537 4236 3543
rect 365 3517 380 3523
rect 429 3517 460 3523
rect 1325 3517 1356 3523
rect 2388 3517 2403 3523
rect 3284 3517 3299 3523
rect 3453 3517 3491 3523
rect 3517 3517 3532 3523
rect 3668 3517 3683 3523
rect 3901 3517 3939 3523
rect 4093 3517 4124 3523
rect 4308 3517 4323 3523
rect 4612 3517 4643 3523
rect 4740 3517 4771 3523
rect 5012 3517 5027 3523
rect 5053 3517 5068 3523
rect 5268 3517 5283 3523
rect 5309 3517 5324 3523
rect 5396 3517 5411 3523
rect 5460 3517 5475 3523
rect 3148 3492 3156 3496
rect 3468 3492 3476 3496
rect 3660 3492 3668 3496
rect 3916 3492 3924 3496
rect 4108 3492 4116 3496
rect 5245 3497 5268 3503
rect 4748 3492 4756 3496
rect 5260 3492 5268 3497
rect 173 3477 188 3483
rect 237 3477 252 3483
rect 638 3477 659 3483
rect 653 3457 659 3477
rect 877 3477 914 3483
rect 2052 3477 2067 3483
rect 2558 3477 2579 3483
rect 2573 3457 2579 3477
rect 2813 3477 2828 3483
rect 4733 3477 4755 3483
rect 4868 3477 4882 3483
rect 4990 3477 5011 3483
rect 332 3444 340 3448
rect 396 3444 404 3448
rect 508 3444 516 3448
rect 1020 3444 1028 3448
rect 1084 3444 1092 3448
rect 1164 3444 1172 3448
rect 1228 3444 1236 3448
rect 1292 3444 1300 3448
rect 1404 3444 1412 3448
rect 1532 3444 1540 3448
rect 1724 3444 1732 3448
rect 1740 3444 1748 3448
rect 1852 3444 1860 3448
rect 1916 3444 1924 3448
rect 1932 3444 1940 3448
rect 1996 3444 2004 3448
rect 2108 3444 2116 3448
rect 2124 3444 2132 3448
rect 2236 3444 2244 3448
rect 2252 3444 2260 3448
rect 2428 3444 2436 3448
rect 2492 3444 2500 3448
rect 2684 3444 2692 3448
rect 3196 3444 3204 3448
rect 3324 3444 3332 3448
rect 3580 3444 3588 3448
rect 3644 3444 3652 3448
rect 3708 3444 3716 3448
rect 3788 3444 3796 3448
rect 4156 3444 4164 3448
rect 4284 3444 4292 3448
rect 4348 3444 4356 3448
rect 4668 3444 4676 3448
rect 4684 3444 4692 3448
rect 4796 3444 4804 3448
rect 5116 3444 5124 3448
rect 5372 3444 5380 3448
rect 5500 3444 5508 3448
rect 5564 3444 5572 3448
rect 5894 3416 5994 3804
rect 5552 3404 5994 3416
rect 12 3372 20 3376
rect 588 3372 596 3376
rect 780 3372 788 3376
rect 844 3372 852 3376
rect 908 3372 916 3376
rect 972 3372 980 3376
rect 1484 3372 1492 3376
rect 1548 3372 1556 3376
rect 1932 3372 1940 3376
rect 2060 3372 2068 3376
rect 2188 3372 2196 3376
rect 2252 3372 2260 3376
rect 2444 3372 2452 3376
rect 2636 3372 2644 3376
rect 2828 3372 2836 3376
rect 3148 3372 3156 3376
rect 3532 3372 3540 3376
rect 3836 3372 3844 3376
rect 4236 3372 4244 3376
rect 4300 3372 4308 3376
rect 4540 3372 4548 3376
rect 4556 3372 4564 3376
rect 4748 3372 4756 3376
rect 4876 3372 4884 3376
rect 4940 3372 4948 3376
rect 5244 3372 5252 3376
rect 5308 3372 5316 3376
rect 5452 3372 5460 3376
rect 109 3337 146 3343
rect 237 3337 252 3343
rect 381 3343 387 3363
rect 381 3337 396 3343
rect 701 3343 707 3363
rect 701 3337 722 3343
rect 1165 3343 1171 3363
rect 1140 3337 1171 3343
rect 1229 3343 1235 3363
rect 1214 3337 1235 3343
rect 1389 3337 1404 3343
rect 1869 3343 1875 3363
rect 2941 3357 2956 3363
rect 1812 3337 1827 3343
rect 1854 3337 1875 3343
rect 2605 3337 2620 3343
rect 2964 3337 2979 3343
rect 3972 3337 3987 3343
rect 4109 3343 4115 3363
rect 4084 3337 4115 3343
rect 4158 3337 4172 3343
rect 4349 3337 4370 3343
rect 5373 3337 5388 3343
rect 1724 3324 1732 3328
rect 2236 3323 2244 3328
rect 2684 3324 2692 3328
rect 2876 3324 2884 3328
rect 3404 3324 3412 3328
rect 2236 3317 2259 3323
rect 3788 3323 3796 3328
rect 3773 3317 3796 3323
rect 4604 3323 4612 3328
rect 4796 3324 4804 3328
rect 4604 3317 4627 3323
rect 5260 3324 5268 3328
rect 45 3297 60 3303
rect 556 3303 564 3316
rect 3804 3304 3812 3316
rect 3996 3304 4004 3316
rect 556 3300 572 3303
rect 557 3297 572 3300
rect 3181 3297 3196 3303
rect 3389 3297 3427 3303
rect 3629 3297 3667 3303
rect 4781 3297 4819 3303
rect 5181 3297 5196 3303
rect 5565 3237 5580 3243
rect -412 3204 16 3216
rect -412 2816 -312 3204
rect 1796 3137 1811 3143
rect 1917 3117 1955 3123
rect 2196 3117 2211 3123
rect 2260 3117 2275 3123
rect 2900 3117 2915 3123
rect 3005 3117 3020 3123
rect 3140 3117 3155 3123
rect 3204 3117 3219 3123
rect 3245 3117 3283 3123
rect 3581 3117 3619 3123
rect 3773 3117 3811 3123
rect 4029 3117 4044 3123
rect 4180 3117 4195 3123
rect 4333 3117 4364 3123
rect 5204 3117 5219 3123
rect 5437 3117 5452 3123
rect 4252 3104 4260 3116
rect 4524 3104 4532 3116
rect 1212 3092 1220 3096
rect 1276 3092 1284 3096
rect 2877 3097 2900 3103
rect 2444 3092 2452 3096
rect 2892 3092 2900 3097
rect 3965 3097 3988 3103
rect 3260 3092 3268 3096
rect 3980 3092 3988 3097
rect 4172 3092 4180 3096
rect 4236 3092 4244 3096
rect 4348 3092 4356 3096
rect 4540 3092 4548 3096
rect 4988 3092 4996 3096
rect 5196 3092 5204 3096
rect 45 3077 82 3083
rect 109 3077 146 3083
rect 180 3077 188 3083
rect 365 3077 380 3083
rect 621 3077 636 3083
rect 749 3077 786 3083
rect 829 3077 850 3083
rect 829 3057 835 3077
rect 941 3077 956 3083
rect 1405 3077 1426 3083
rect 1405 3057 1411 3077
rect 3908 3077 3939 3083
rect 204 3044 212 3048
rect 1020 3044 1028 3048
rect 1084 3044 1092 3048
rect 1164 3044 1172 3048
rect 1228 3044 1236 3048
rect 1484 3044 1492 3048
rect 1548 3044 1556 3048
rect 1660 3044 1668 3048
rect 1740 3044 1748 3048
rect 1980 3044 1988 3048
rect 2236 3044 2244 3048
rect 2300 3044 2308 3048
rect 2428 3044 2436 3048
rect 2492 3044 2500 3048
rect 2508 3044 2516 3048
rect 2636 3044 2644 3048
rect 3084 3044 3092 3048
rect 3836 3044 3844 3048
rect 4092 3044 4100 3048
rect 4156 3044 4164 3048
rect 4220 3044 4228 3048
rect 4300 3044 4308 3048
rect 4412 3044 4420 3048
rect 4492 3044 4500 3048
rect 4556 3044 4564 3048
rect 4732 3044 4740 3048
rect 4940 3044 4948 3048
rect 5068 3044 5076 3048
rect 5244 3044 5252 3048
rect 5372 3044 5380 3048
rect 5500 3044 5508 3048
rect 5894 3016 5994 3404
rect 5552 3004 5994 3016
rect 188 2972 196 2976
rect 316 2972 324 2976
rect 380 2972 388 2976
rect 700 2972 708 2976
rect 780 2972 788 2976
rect 908 2972 916 2976
rect 972 2972 980 2976
rect 1084 2972 1092 2976
rect 1404 2972 1412 2976
rect 1852 2972 1860 2976
rect 1868 2972 1876 2976
rect 1980 2972 1988 2976
rect 2188 2972 2196 2976
rect 2428 2972 2436 2976
rect 2684 2972 2692 2976
rect 2764 2972 2772 2976
rect 3084 2972 3092 2976
rect 3276 2972 3284 2976
rect 3980 2972 3988 2976
rect 4092 2972 4100 2976
rect 4364 2972 4372 2976
rect 4492 2972 4500 2976
rect 4556 2972 4564 2976
rect 4684 2972 4692 2976
rect 5116 2972 5124 2976
rect 5180 2972 5188 2976
rect 5308 2972 5316 2976
rect 5564 2972 5572 2976
rect 1485 2943 1491 2963
rect 1470 2937 1491 2943
rect 1709 2937 1724 2943
rect 2372 2937 2387 2943
rect 2573 2943 2579 2963
rect 2516 2937 2531 2943
rect 2558 2937 2579 2943
rect 3325 2937 3340 2943
rect 5374 2937 5395 2943
rect 2812 2924 2820 2928
rect 3132 2924 3140 2928
rect 3596 2924 3604 2928
rect 3900 2923 3908 2928
rect 3900 2917 3923 2923
rect 4172 2923 4180 2928
rect 4876 2924 4884 2928
rect 5068 2924 5076 2928
rect 4164 2917 4180 2923
rect 5132 2924 5140 2928
rect 5452 2923 5460 2928
rect 5437 2917 5460 2923
rect 1948 2904 1956 2916
rect 4892 2904 4900 2916
rect 253 2897 268 2903
rect 493 2897 508 2903
rect 637 2897 675 2903
rect 1005 2897 1020 2903
rect 1812 2897 1827 2903
rect 4589 2897 4627 2903
rect 5460 2897 5475 2903
rect 1341 2877 1356 2883
rect -412 2804 18 2816
rect -412 2416 -312 2804
rect 788 2717 803 2723
rect 3012 2717 3027 2723
rect 3348 2717 3363 2723
rect 3837 2717 3875 2723
rect 3924 2717 3939 2723
rect 4077 2717 4092 2723
rect 4692 2717 4707 2723
rect 4932 2717 4963 2723
rect 4989 2717 5004 2723
rect 5437 2717 5452 2723
rect 5524 2717 5539 2723
rect 2813 2697 2836 2703
rect 2828 2692 2836 2697
rect 3197 2697 3220 2703
rect 2940 2692 2948 2696
rect 3212 2692 3220 2697
rect 3708 2692 3716 2696
rect 5181 2697 5204 2703
rect 3852 2692 3860 2696
rect 5196 2692 5204 2697
rect 62 2677 83 2683
rect 77 2657 83 2677
rect 660 2677 675 2683
rect 1156 2677 1187 2683
rect 2388 2677 2403 2683
rect 2516 2677 2531 2683
rect 2580 2677 2595 2683
rect 2749 2677 2780 2683
rect 2749 2657 2755 2677
rect 3524 2677 3539 2683
rect 4477 2677 4492 2683
rect 4798 2677 4819 2683
rect 188 2644 196 2648
rect 268 2644 276 2648
rect 460 2644 468 2648
rect 828 2644 836 2648
rect 972 2644 980 2648
rect 1036 2644 1044 2648
rect 1468 2644 1476 2648
rect 1532 2644 1540 2648
rect 1596 2644 1604 2648
rect 1852 2644 1860 2648
rect 1868 2644 1876 2648
rect 2044 2644 2052 2648
rect 2364 2644 2372 2648
rect 2684 2644 2692 2648
rect 2876 2644 2884 2648
rect 2956 2644 2964 2648
rect 3132 2644 3140 2648
rect 3260 2644 3268 2648
rect 3388 2644 3396 2648
rect 3580 2644 3588 2648
rect 3660 2644 3668 2648
rect 3900 2644 3908 2648
rect 4028 2644 4036 2648
rect 4044 2644 4052 2648
rect 4172 2644 4180 2648
rect 4284 2644 4292 2648
rect 4364 2644 4372 2648
rect 4540 2644 4548 2648
rect 4732 2644 4740 2648
rect 5052 2644 5060 2648
rect 5308 2644 5316 2648
rect 5500 2644 5508 2648
rect 5564 2643 5572 2648
rect 5564 2637 5580 2643
rect 5894 2616 5994 3004
rect 5552 2604 5994 2616
rect 204 2572 212 2576
rect 316 2572 324 2576
rect 1356 2572 1364 2576
rect 2108 2572 2116 2576
rect 2316 2572 2324 2576
rect 2492 2572 2500 2576
rect 2556 2572 2564 2576
rect 2940 2572 2948 2576
rect 3324 2572 3332 2576
rect 3580 2572 3588 2576
rect 3596 2572 3604 2576
rect 3772 2572 3780 2576
rect 3836 2572 3844 2576
rect 4108 2572 4116 2576
rect 4300 2572 4308 2576
rect 4492 2572 4500 2576
rect 4860 2572 4868 2576
rect 4876 2572 4884 2576
rect 5052 2572 5060 2576
rect 5116 2572 5124 2576
rect 5180 2572 5188 2576
rect 5308 2572 5316 2576
rect 5436 2572 5444 2576
rect 5564 2572 5572 2576
rect 365 2537 380 2543
rect 429 2537 460 2543
rect 621 2537 668 2543
rect 772 2537 786 2543
rect 829 2543 835 2563
rect 829 2537 850 2543
rect 1214 2537 1228 2543
rect 1709 2537 1746 2543
rect 1773 2537 1788 2543
rect 1981 2543 1987 2563
rect 1981 2537 2002 2543
rect 2173 2543 2179 2563
rect 2173 2537 2194 2543
rect 2221 2537 2252 2543
rect 2605 2537 2642 2543
rect 4212 2537 4259 2543
rect 4948 2537 4963 2543
rect 2764 2523 2772 2528
rect 2828 2523 2836 2528
rect 2892 2523 2900 2528
rect 2749 2517 2772 2523
rect 2813 2517 2836 2523
rect 2877 2517 2900 2523
rect 3452 2523 3460 2528
rect 3452 2517 3475 2523
rect 4156 2523 4164 2528
rect 4732 2524 4740 2528
rect 4156 2517 4172 2523
rect 4812 2523 4820 2528
rect 4797 2517 4820 2523
rect 5004 2524 5012 2528
rect 2349 2497 2387 2503
rect 2900 2497 2915 2503
rect 3348 2497 3363 2503
rect 3732 2497 3747 2503
rect 4909 2497 4924 2503
rect 5396 2497 5411 2503
rect 5245 2477 5260 2483
rect -412 2404 26 2416
rect -412 2016 -312 2404
rect 109 2317 124 2323
rect 2196 2317 2211 2323
rect 2621 2317 2659 2323
rect 3604 2317 3619 2323
rect 4084 2317 4115 2323
rect 4740 2317 4755 2323
rect 3372 2304 3380 2316
rect 3676 2304 3684 2316
rect 4268 2304 4276 2316
rect 2956 2292 2964 2296
rect 3516 2292 3524 2296
rect 3724 2292 3732 2296
rect 3916 2292 3924 2296
rect 4092 2292 4100 2296
rect 4284 2292 4292 2296
rect 4940 2292 4948 2296
rect 125 2277 140 2283
rect 276 2277 291 2283
rect 852 2277 867 2283
rect 980 2277 995 2283
rect 1213 2277 1234 2283
rect 1213 2257 1219 2277
rect 1364 2277 1379 2283
rect 1645 2277 1660 2283
rect 2365 2277 2386 2283
rect 2413 2277 2428 2283
rect 2365 2257 2371 2277
rect 4484 2277 4499 2283
rect 4564 2277 4579 2283
rect 4606 2277 4627 2283
rect 76 2244 84 2248
rect 188 2244 196 2248
rect 652 2244 660 2248
rect 908 2244 916 2248
rect 1100 2244 1108 2248
rect 1292 2244 1300 2248
rect 1532 2244 1540 2248
rect 1740 2244 1748 2248
rect 1996 2244 2004 2248
rect 2236 2244 2244 2248
rect 2684 2244 2692 2248
rect 2748 2244 2756 2248
rect 2812 2244 2820 2248
rect 2876 2244 2884 2248
rect 3004 2244 3012 2248
rect 3148 2244 3156 2248
rect 3324 2244 3332 2248
rect 3468 2244 3476 2248
rect 3708 2244 3716 2248
rect 3772 2244 3780 2248
rect 3836 2244 3844 2248
rect 3964 2244 3972 2248
rect 4044 2244 4052 2248
rect 4220 2244 4228 2248
rect 4540 2244 4548 2248
rect 4668 2244 4676 2248
rect 4684 2244 4692 2248
rect 4988 2244 4996 2248
rect 5052 2244 5060 2248
rect 5180 2244 5188 2248
rect 5436 2244 5444 2248
rect 5894 2216 5994 2604
rect 5552 2204 5994 2216
rect 204 2172 212 2176
rect 572 2172 580 2176
rect 716 2172 724 2176
rect 1036 2172 1044 2176
rect 1100 2172 1108 2176
rect 1276 2172 1284 2176
rect 1292 2172 1300 2176
rect 1420 2172 1428 2176
rect 1740 2172 1748 2176
rect 1868 2172 1876 2176
rect 1980 2172 1988 2176
rect 2108 2172 2116 2176
rect 2172 2172 2180 2176
rect 2364 2172 2372 2176
rect 2380 2172 2388 2176
rect 2492 2172 2500 2176
rect 2876 2172 2884 2176
rect 2892 2172 2900 2176
rect 2956 2172 2964 2176
rect 3260 2172 3268 2176
rect 3276 2172 3284 2176
rect 3452 2172 3460 2176
rect 3580 2172 3588 2176
rect 3772 2172 3780 2176
rect 3788 2172 3796 2176
rect 3900 2172 3908 2176
rect 3916 2172 3924 2176
rect 4156 2172 4164 2176
rect 4220 2172 4228 2176
rect 4236 2172 4244 2176
rect 4364 2172 4372 2176
rect 4620 2172 4628 2176
rect 4940 2172 4948 2176
rect 5324 2172 5332 2176
rect 5500 2172 5508 2176
rect 5564 2172 5572 2176
rect 125 2143 131 2163
rect 125 2137 146 2143
rect 381 2143 387 2163
rect 381 2137 402 2143
rect 660 2137 675 2143
rect 829 2143 835 2163
rect 829 2137 860 2143
rect 1604 2137 1618 2143
rect 2765 2143 2771 2163
rect 3069 2157 3084 2163
rect 2708 2137 2723 2143
rect 2750 2137 2771 2143
rect 3524 2137 3539 2143
rect 3710 2137 3731 2143
rect 3988 2137 4003 2143
rect 4077 2137 4092 2143
rect 4493 2143 4499 2163
rect 4468 2137 4499 2143
rect 4557 2143 4563 2163
rect 4542 2137 4563 2143
rect 2940 2124 2948 2128
rect 3148 2123 3156 2128
rect 3133 2117 3156 2123
rect 3212 2124 3220 2128
rect 4172 2124 4180 2128
rect 4284 2124 4292 2128
rect 4684 2124 4692 2128
rect 4812 2123 4820 2128
rect 5068 2124 5076 2128
rect 4797 2117 4820 2123
rect 924 2103 932 2116
rect 4396 2104 4404 2116
rect 916 2100 932 2103
rect 916 2097 931 2100
rect 1796 2097 1811 2103
rect 1901 2097 1932 2103
rect 3156 2097 3171 2103
rect 3309 2097 3340 2103
rect 4676 2097 4707 2103
rect 4733 2097 4771 2103
rect 5524 2097 5539 2103
rect 5437 2077 5452 2083
rect -412 2004 26 2016
rect -412 1616 -312 2004
rect 1684 1917 1699 1923
rect 3133 1917 3171 1923
rect 3325 1917 3340 1923
rect 3476 1917 3491 1923
rect 4868 1917 4883 1923
rect 5309 1917 5324 1923
rect 3612 1904 3620 1916
rect 4076 1904 4084 1916
rect 4908 1904 4916 1916
rect 3453 1897 3476 1903
rect 3148 1892 3156 1896
rect 3468 1892 3476 1897
rect 3901 1897 3924 1903
rect 3916 1892 3924 1897
rect 5245 1897 5268 1903
rect 4748 1892 4756 1896
rect 5068 1892 5076 1896
rect 5260 1892 5268 1897
rect 61 1877 82 1883
rect 61 1857 67 1877
rect 637 1877 652 1883
rect 893 1877 908 1883
rect 893 1857 899 1877
rect 1389 1877 1426 1883
rect 1533 1877 1554 1883
rect 1213 1857 1219 1876
rect 1533 1857 1539 1877
rect 1917 1877 1938 1883
rect 1917 1857 1923 1877
rect 1988 1877 2019 1883
rect 2110 1877 2131 1883
rect 2125 1857 2131 1877
rect 2477 1877 2514 1883
rect 2797 1877 2828 1883
rect 3540 1877 3555 1883
rect 3860 1877 3875 1883
rect 4093 1877 4108 1883
rect 5181 1877 5196 1883
rect 4548 1857 4563 1863
rect 252 1844 260 1848
rect 380 1844 388 1848
rect 460 1844 468 1848
rect 588 1844 596 1848
rect 972 1844 980 1848
rect 1036 1844 1044 1848
rect 2300 1844 2308 1848
rect 2380 1844 2388 1848
rect 2700 1844 2708 1848
rect 3644 1844 3652 1848
rect 3772 1844 3780 1848
rect 3964 1844 3972 1848
rect 3980 1844 3988 1848
rect 4172 1844 4180 1848
rect 4412 1844 4420 1848
rect 4796 1844 4804 1848
rect 5116 1844 5124 1848
rect 5500 1844 5508 1848
rect 5564 1844 5572 1848
rect 5894 1816 5994 2204
rect 5552 1804 5994 1816
rect 140 1772 148 1776
rect 828 1772 836 1776
rect 844 1772 852 1776
rect 1036 1772 1044 1776
rect 1276 1772 1284 1776
rect 1356 1772 1364 1776
rect 1548 1772 1556 1776
rect 1612 1772 1620 1776
rect 1916 1772 1924 1776
rect 2188 1772 2196 1776
rect 2252 1772 2260 1776
rect 2492 1772 2500 1776
rect 2572 1772 2580 1776
rect 2684 1772 2692 1776
rect 2748 1772 2756 1776
rect 2876 1772 2884 1776
rect 2956 1772 2964 1776
rect 3212 1772 3220 1776
rect 3324 1772 3332 1776
rect 3404 1772 3412 1776
rect 3516 1772 3524 1776
rect 3596 1772 3604 1776
rect 3772 1772 3780 1776
rect 3964 1772 3972 1776
rect 4028 1772 4036 1776
rect 4092 1772 4100 1776
rect 4108 1772 4116 1776
rect 4364 1772 4372 1776
rect 4860 1772 4868 1776
rect 4988 1772 4996 1776
rect 5244 1772 5252 1776
rect 5260 1772 5268 1776
rect 5372 1772 5380 1776
rect 5436 1772 5444 1776
rect 5564 1772 5572 1776
rect 45 1737 60 1743
rect 237 1737 274 1743
rect 429 1737 444 1743
rect 1476 1737 1507 1743
rect 1709 1737 1724 1743
rect 1773 1737 1788 1743
rect 2324 1737 2339 1743
rect 4285 1737 4300 1743
rect 4541 1737 4562 1743
rect 4717 1737 4732 1743
rect 5012 1737 5027 1743
rect 2300 1724 2308 1728
rect 3004 1724 3012 1728
rect 3452 1724 3460 1728
rect 3724 1723 3732 1728
rect 3916 1723 3924 1728
rect 3709 1717 3732 1723
rect 3901 1717 3924 1723
rect 4044 1724 4052 1728
rect 4156 1723 4164 1728
rect 4220 1723 4228 1728
rect 4412 1724 4420 1728
rect 4156 1717 4179 1723
rect 4220 1717 4243 1723
rect 4748 1724 4756 1728
rect 4940 1723 4948 1728
rect 4925 1717 4948 1723
rect 5196 1724 5204 1728
rect 173 1697 188 1703
rect 765 1697 803 1703
rect 1213 1697 1251 1703
rect 2221 1697 2236 1703
rect 2285 1697 2300 1703
rect 2452 1697 2467 1703
rect 2836 1697 2851 1703
rect 3092 1697 3107 1703
rect 3629 1697 3644 1703
rect 4397 1697 4435 1703
rect 5181 1697 5219 1703
rect 5300 1697 5347 1703
rect -412 1604 28 1616
rect -412 1216 -312 1604
rect 2244 1537 2259 1543
rect 3076 1537 3091 1543
rect 813 1517 828 1523
rect 3284 1517 3299 1523
rect 3885 1517 3900 1523
rect 3988 1517 4003 1523
rect 4180 1517 4195 1523
rect 4397 1517 4435 1523
rect 4884 1517 4899 1523
rect 5140 1517 5155 1523
rect 5332 1517 5347 1523
rect 5460 1517 5475 1523
rect 5501 1517 5516 1523
rect 1884 1504 1892 1516
rect 3068 1492 3076 1496
rect 3580 1497 3603 1503
rect 3340 1492 3348 1496
rect 3580 1492 3588 1497
rect 4412 1492 4420 1496
rect 4684 1492 4692 1496
rect 5116 1492 5124 1496
rect 5436 1492 5444 1496
rect 237 1477 274 1483
rect 301 1477 338 1483
rect 509 1477 530 1483
rect 557 1477 594 1483
rect 621 1477 636 1483
rect 509 1457 515 1477
rect 660 1477 675 1483
rect 749 1477 764 1483
rect 893 1477 914 1483
rect 893 1457 899 1477
rect 2477 1477 2492 1483
rect 2925 1477 2956 1483
rect 3245 1477 3260 1483
rect 3901 1477 3916 1483
rect 4084 1477 4092 1483
rect 4996 1477 5011 1483
rect 5204 1477 5219 1483
rect 5246 1477 5267 1483
rect 444 1444 452 1448
rect 780 1444 788 1448
rect 972 1444 980 1448
rect 2188 1444 2196 1448
rect 2364 1444 2372 1448
rect 2636 1444 2644 1448
rect 3020 1444 3028 1448
rect 3388 1444 3396 1448
rect 3532 1444 3540 1448
rect 3836 1444 3844 1448
rect 4108 1444 4116 1448
rect 4220 1444 4228 1448
rect 4300 1444 4308 1448
rect 4492 1444 4500 1448
rect 4668 1444 4676 1448
rect 4924 1444 4932 1448
rect 5052 1444 5060 1448
rect 5068 1444 5076 1448
rect 5308 1444 5316 1448
rect 5388 1444 5396 1448
rect 5564 1444 5572 1448
rect 5894 1416 5994 1804
rect 5552 1404 5994 1416
rect 140 1372 148 1376
rect 316 1372 324 1376
rect 572 1372 580 1376
rect 716 1372 724 1376
rect 780 1372 788 1376
rect 1660 1372 1668 1376
rect 1804 1372 1812 1376
rect 1996 1372 2004 1376
rect 2300 1372 2308 1376
rect 2684 1372 2692 1376
rect 2812 1372 2820 1376
rect 3084 1372 3092 1376
rect 3276 1372 3284 1376
rect 3468 1372 3476 1376
rect 3532 1372 3540 1376
rect 3644 1372 3652 1376
rect 3916 1372 3924 1376
rect 4028 1372 4036 1376
rect 4044 1372 4052 1376
rect 4108 1372 4116 1376
rect 4540 1372 4548 1376
rect 4620 1372 4628 1376
rect 4860 1372 4868 1376
rect 4924 1372 4932 1376
rect 5116 1372 5124 1376
rect 5132 1372 5140 1376
rect 5244 1372 5252 1376
rect 5372 1372 5380 1376
rect 5436 1372 5444 1376
rect 5452 1372 5460 1376
rect 365 1337 380 1343
rect 877 1337 892 1343
rect 1492 1337 1500 1343
rect 1556 1337 1571 1343
rect 2196 1337 2211 1343
rect 2429 1337 2444 1343
rect 3725 1343 3731 1363
rect 3716 1337 3731 1343
rect 2572 1323 2580 1328
rect 2557 1317 2580 1323
rect 2892 1323 2900 1328
rect 2877 1317 2900 1323
rect 3004 1323 3012 1328
rect 3004 1317 3027 1323
rect 4668 1323 4676 1328
rect 4668 1317 4691 1323
rect 2029 1297 2044 1303
rect 2836 1297 2851 1303
rect 2989 1297 3004 1303
rect 3972 1297 4003 1303
rect 4077 1297 4092 1303
rect 4244 1297 4259 1303
rect 4413 1297 4451 1303
rect 4477 1297 4492 1303
rect 4653 1297 4668 1303
rect 4989 1297 5027 1303
rect 5165 1297 5180 1303
rect 5204 1297 5219 1303
rect 3837 1277 3852 1283
rect 4221 1277 4236 1283
rect 4349 1277 4364 1283
rect -412 1204 26 1216
rect -412 816 -312 1204
rect 4164 1137 4179 1143
rect 429 1117 476 1123
rect 813 1117 828 1123
rect 980 1117 995 1123
rect 1405 1123 1411 1136
rect 1405 1117 1443 1123
rect 2116 1117 2147 1123
rect 3437 1117 3452 1123
rect 3796 1117 3811 1123
rect 4461 1117 4476 1123
rect 4733 1117 4748 1123
rect 2860 1104 2868 1116
rect 4396 1104 4404 1116
rect 4764 1104 4772 1116
rect 572 1097 595 1103
rect 572 1092 580 1097
rect 3324 1097 3347 1103
rect 3773 1097 3796 1103
rect 2876 1092 2884 1096
rect 3324 1092 3332 1097
rect 3788 1092 3796 1097
rect 4044 1092 4052 1096
rect 4156 1092 4164 1096
rect 4348 1092 4356 1096
rect 4620 1092 4628 1096
rect 5004 1092 5012 1096
rect 5436 1092 5444 1096
rect 1534 1077 1555 1083
rect 1549 1057 1555 1077
rect 2989 1077 3004 1083
rect 3508 1077 3539 1083
rect 3533 1057 3539 1077
rect 4477 1077 4492 1083
rect 396 1044 404 1048
rect 508 1044 516 1048
rect 716 1044 724 1048
rect 892 1044 900 1048
rect 1020 1044 1028 1048
rect 1036 1044 1044 1048
rect 1148 1044 1156 1048
rect 1164 1044 1172 1048
rect 1228 1044 1236 1048
rect 1356 1044 1364 1048
rect 1468 1044 1476 1048
rect 1788 1044 1796 1048
rect 1980 1044 1988 1048
rect 2060 1044 2068 1048
rect 2172 1044 2180 1048
rect 2188 1044 2196 1048
rect 2572 1044 2580 1048
rect 2764 1044 2772 1048
rect 3404 1044 3412 1048
rect 3836 1044 3844 1048
rect 4300 1044 4308 1048
rect 4364 1044 4372 1048
rect 4556 1044 4564 1048
rect 4668 1044 4676 1048
rect 4796 1044 4804 1048
rect 4940 1044 4948 1048
rect 5052 1044 5060 1048
rect 5116 1044 5124 1048
rect 5244 1044 5252 1048
rect 5372 1044 5380 1048
rect 5501 1037 5516 1043
rect 5894 1016 5994 1404
rect 5552 1004 5994 1016
rect 140 972 148 976
rect 332 972 340 976
rect 652 972 660 976
rect 1548 972 1556 976
rect 1996 972 2004 976
rect 2108 972 2116 976
rect 2252 972 2260 976
rect 2572 972 2580 976
rect 2700 972 2708 976
rect 2812 972 2820 976
rect 2828 972 2836 976
rect 2940 972 2948 976
rect 3260 972 3268 976
rect 3324 972 3332 976
rect 3340 972 3348 976
rect 3532 972 3540 976
rect 3852 972 3860 976
rect 3964 972 3972 976
rect 3980 972 3988 976
rect 4092 972 4100 976
rect 4364 972 4372 976
rect 4604 972 4612 976
rect 4860 972 4868 976
rect 4876 972 4884 976
rect 4988 972 4996 976
rect 5244 972 5252 976
rect 5436 972 5444 976
rect 5452 972 5460 976
rect 61 943 67 963
rect 61 937 82 943
rect 244 937 274 943
rect 916 937 931 943
rect 1037 943 1043 963
rect 1028 937 1043 943
rect 1156 937 1170 943
rect 1197 937 1212 943
rect 1277 943 1283 963
rect 1277 937 1298 943
rect 1453 937 1484 943
rect 1726 937 1763 943
rect 1965 937 1980 943
rect 2045 937 2060 943
rect 3149 943 3155 963
rect 3134 937 3155 943
rect 3636 937 3683 943
rect 3757 937 3772 943
rect 2508 924 2516 928
rect 596 897 611 903
rect 2484 897 2531 903
rect 2765 883 2771 928
rect 3212 923 3220 928
rect 3197 917 3220 923
rect 3580 923 3588 928
rect 4220 924 4228 928
rect 3580 917 3603 923
rect 4492 923 4500 928
rect 4812 924 4820 928
rect 4477 917 4500 923
rect 5196 924 5204 928
rect 4012 904 4020 916
rect 4508 904 4516 916
rect 2861 897 2876 903
rect 2989 897 3020 903
rect 4205 897 4220 903
rect 4541 897 4579 903
rect 2756 877 2771 883
rect -412 804 22 816
rect -412 416 -312 804
rect 445 737 460 743
rect 173 717 188 723
rect 237 717 252 723
rect 445 692 451 737
rect 685 717 700 723
rect 724 717 739 723
rect 1389 720 1404 723
rect 1388 717 1404 720
rect 1388 704 1396 717
rect 1661 717 1699 723
rect 2477 717 2492 723
rect 3476 717 3491 723
rect 3565 717 3603 723
rect 4269 717 4300 723
rect 4925 717 4963 723
rect 5165 717 5180 723
rect 5204 717 5219 723
rect 2908 704 2916 716
rect 3868 704 3876 716
rect 5292 704 5300 716
rect 3453 697 3476 703
rect 3468 692 3476 697
rect 3580 692 3588 696
rect 3852 692 3860 696
rect 4940 692 4948 696
rect 5452 692 5460 696
rect 45 677 82 683
rect 941 677 978 683
rect 1021 677 1042 683
rect 1021 657 1027 677
rect 1517 677 1532 683
rect 1790 677 1811 683
rect 1805 657 1811 677
rect 2685 677 2700 683
rect 3326 677 3347 683
rect 3341 664 3347 677
rect 3629 677 3644 683
rect 140 644 148 648
rect 204 644 212 648
rect 316 644 324 648
rect 396 644 404 648
rect 508 644 516 648
rect 572 644 580 648
rect 652 644 660 648
rect 764 644 772 648
rect 828 644 836 648
rect 1212 644 1220 648
rect 1356 644 1364 648
rect 1468 644 1476 648
rect 1724 644 1732 648
rect 1916 644 1924 648
rect 2300 644 2308 648
rect 2316 644 2324 648
rect 2380 644 2388 648
rect 2444 644 2452 648
rect 2508 644 2516 648
rect 2748 644 2756 648
rect 3532 644 3540 648
rect 4236 644 4244 648
rect 4348 644 4356 648
rect 4428 644 4436 648
rect 4540 644 4548 648
rect 4604 644 4612 648
rect 4988 644 4996 648
rect 5004 644 5012 648
rect 5436 644 5444 648
rect 5894 616 5994 1004
rect 5552 604 5994 616
rect 204 572 212 576
rect 316 572 324 576
rect 460 572 468 576
rect 764 572 772 576
rect 908 572 916 576
rect 1228 572 1236 576
rect 2172 572 2180 576
rect 2380 572 2388 576
rect 2492 572 2500 576
rect 2556 572 2564 576
rect 2956 572 2964 576
rect 3084 572 3092 576
rect 3148 572 3156 576
rect 3276 572 3284 576
rect 3468 572 3476 576
rect 3772 572 3780 576
rect 3964 572 3972 576
rect 4092 572 4100 576
rect 4236 572 4244 576
rect 4348 572 4356 576
rect 4364 572 4372 576
rect 4556 572 4564 576
rect 4796 572 4804 576
rect 4876 572 4884 576
rect 5132 572 5140 576
rect 5500 572 5508 576
rect 589 543 595 563
rect 574 537 595 543
rect 653 543 659 563
rect 638 537 659 543
rect 1022 537 1059 543
rect 1620 537 1635 543
rect 1901 537 1916 543
rect 2237 543 2243 563
rect 2237 537 2258 543
rect 2285 537 2300 543
rect 2733 537 2748 543
rect 4740 537 4755 543
rect 4996 537 5010 543
rect 3580 523 3588 528
rect 3724 523 3732 528
rect 3916 523 3924 528
rect 4044 523 4052 528
rect 4284 524 4292 528
rect 5452 524 5460 528
rect 3580 517 3603 523
rect 3709 517 3732 523
rect 3901 517 3924 523
rect 4029 517 4052 523
rect 3564 504 3572 516
rect 4060 504 4068 516
rect 877 497 915 503
rect 1149 497 1187 503
rect 2132 497 2147 503
rect 2797 497 2835 503
rect 3501 497 3539 503
rect 3732 497 3747 503
rect 3924 497 3939 503
rect 4397 497 4435 503
rect -412 404 24 416
rect -412 16 -312 404
rect 580 337 595 343
rect 1220 317 1235 323
rect 1837 317 1875 323
rect 2093 317 2124 323
rect 2733 317 2748 323
rect 2772 317 2780 323
rect 2964 317 2979 323
rect 4973 317 4988 323
rect 4012 304 4020 316
rect 4572 304 4580 316
rect 4780 304 4788 316
rect 2941 297 2964 303
rect 2956 292 2964 297
rect 4541 297 4564 303
rect 4476 292 4484 296
rect 4556 292 4564 297
rect 4988 297 5011 303
rect 4620 292 4628 296
rect 4796 292 4804 296
rect 4988 292 4996 297
rect 637 277 658 283
rect 685 277 700 283
rect 637 257 643 277
rect 772 277 786 283
rect 958 277 995 283
rect 2324 277 2339 283
rect 2756 277 2771 283
rect 3092 277 3100 283
rect 4029 277 4044 283
rect 4158 277 4179 283
rect 4173 257 4179 277
rect 4292 277 4323 283
rect 5460 277 5475 283
rect 60 244 68 248
rect 268 244 276 248
rect 332 244 340 248
rect 524 244 532 248
rect 1740 244 1748 248
rect 1804 244 1812 248
rect 1980 244 1988 248
rect 1996 244 2004 248
rect 2060 244 2068 248
rect 2172 244 2180 248
rect 2300 244 2308 248
rect 2380 244 2388 248
rect 3980 244 3988 248
rect 4428 244 4436 248
rect 4604 244 4612 248
rect 4668 244 4676 248
rect 4748 244 4756 248
rect 4940 244 4948 248
rect 5068 244 5076 248
rect 5196 244 5204 248
rect 5894 216 5994 604
rect 5552 204 5994 216
rect 956 172 964 176
rect 1036 172 1044 176
rect 2188 172 2196 176
rect 2700 172 2708 176
rect 2764 172 2772 176
rect 2876 172 2884 176
rect 3148 172 3156 176
rect 3660 172 3668 176
rect 4044 172 4052 176
rect 4156 172 4164 176
rect 4796 172 4804 176
rect 5052 172 5060 176
rect 5068 172 5076 176
rect 5132 172 5140 176
rect 5244 172 5252 176
rect 5308 172 5316 176
rect 5436 172 5444 176
rect 5500 177 5580 183
rect 5500 172 5508 177
rect 333 143 339 163
rect 318 137 339 143
rect 382 137 419 143
rect 781 143 787 163
rect 766 137 787 143
rect 1165 143 1171 163
rect 1150 137 1171 143
rect 1389 137 1420 143
rect 1485 143 1491 163
rect 1470 137 1491 143
rect 1581 137 1612 143
rect 1997 143 2003 163
rect 1988 137 2003 143
rect 2093 137 2108 143
rect 2301 143 2307 163
rect 2301 137 2322 143
rect 2349 137 2364 143
rect 2413 137 2428 143
rect 3373 137 3404 143
rect 3476 137 3491 143
rect 4093 137 4108 143
rect 3260 124 3268 128
rect 173 97 211 103
rect 893 97 924 103
rect 980 97 995 103
rect 2157 97 2172 103
rect 2484 97 2515 103
rect 2733 97 2748 103
rect 2796 103 2804 116
rect 3708 123 3716 128
rect 3900 123 3908 128
rect 4364 124 4372 128
rect 3708 117 3731 123
rect 3900 117 3923 123
rect 4492 123 4500 128
rect 4748 124 4756 128
rect 4477 117 4500 123
rect 4860 123 4868 128
rect 4860 117 4883 123
rect 2796 100 2812 103
rect 2797 97 2812 100
rect 2844 103 2852 116
rect 4076 104 4084 116
rect 4844 104 4852 116
rect 5020 104 5028 116
rect 5388 123 5396 128
rect 5373 117 5396 123
rect 5164 104 5172 116
rect 2820 100 2852 103
rect 2820 97 2851 100
rect 3181 97 3219 103
rect 3245 97 3283 103
rect 4100 97 4131 103
rect 4372 97 4387 103
rect -412 4 30 16
rect -412 0 -312 4
rect 5894 -2 5994 204
<< m2contact >>
rect 508 3976 516 3984
rect 1612 3976 1620 3984
rect 1740 3976 1748 3984
rect 188 3956 196 3964
rect 1804 3956 1812 3964
rect 2684 3956 2692 3964
rect 1852 3936 1860 3944
rect 3388 3936 3396 3944
rect 3644 3936 3652 3944
rect 3964 3936 3972 3944
rect 4156 3936 4164 3944
rect 4348 3936 4356 3944
rect 5068 3936 5076 3944
rect 268 3916 276 3924
rect 860 3916 868 3924
rect 924 3916 932 3924
rect 1036 3916 1044 3924
rect 1196 3916 1204 3924
rect 1436 3916 1444 3924
rect 1484 3916 1492 3924
rect 1516 3916 1524 3924
rect 1580 3916 1588 3924
rect 1644 3916 1652 3924
rect 1708 3916 1716 3924
rect 1772 3916 1780 3924
rect 1852 3916 1860 3924
rect 1916 3916 1924 3924
rect 1964 3916 1972 3924
rect 2012 3916 2020 3924
rect 2092 3916 2100 3924
rect 2156 3916 2164 3924
rect 2284 3916 2292 3924
rect 2428 3916 2436 3924
rect 2556 3916 2564 3924
rect 3132 3916 3140 3924
rect 3180 3916 3188 3924
rect 3596 3916 3604 3924
rect 3612 3916 3620 3924
rect 3820 3916 3828 3924
rect 4044 3916 4052 3924
rect 4060 3916 4068 3924
rect 4188 3916 4196 3924
rect 4252 3916 4260 3924
rect 4396 3916 4404 3924
rect 4524 3916 4532 3924
rect 4572 3916 4580 3924
rect 4620 3916 4628 3924
rect 4636 3916 4644 3924
rect 4684 3916 4692 3924
rect 4716 3916 4724 3924
rect 4924 3916 4932 3924
rect 5004 3916 5012 3924
rect 5100 3916 5108 3924
rect 5148 3916 5156 3924
rect 5196 3916 5204 3924
rect 5212 3916 5220 3924
rect 5292 3916 5300 3924
rect 5468 3916 5476 3924
rect 892 3896 900 3904
rect 1228 3896 1236 3904
rect 1900 3896 1908 3904
rect 2364 3896 2372 3904
rect 3004 3896 3012 3904
rect 3148 3896 3156 3904
rect 3260 3896 3268 3904
rect 3340 3896 3348 3904
rect 3452 3896 3460 3904
rect 3548 3896 3556 3904
rect 3724 3896 3732 3904
rect 3788 3896 3796 3904
rect 4236 3896 4244 3904
rect 4492 3896 4500 3904
rect 4764 3896 4772 3904
rect 5340 3896 5348 3904
rect 28 3876 36 3884
rect 12 3856 20 3864
rect 92 3876 100 3884
rect 140 3876 148 3884
rect 220 3876 228 3884
rect 300 3876 308 3884
rect 204 3856 212 3864
rect 364 3876 372 3884
rect 412 3876 420 3884
rect 522 3876 530 3884
rect 620 3876 628 3884
rect 380 3856 388 3864
rect 396 3856 404 3864
rect 460 3856 468 3864
rect 572 3856 580 3864
rect 684 3876 692 3884
rect 700 3876 708 3884
rect 748 3876 756 3884
rect 812 3876 820 3884
rect 844 3876 852 3884
rect 908 3876 916 3884
rect 988 3876 996 3884
rect 1022 3876 1030 3884
rect 1068 3876 1076 3884
rect 700 3856 708 3864
rect 764 3856 772 3864
rect 828 3856 836 3864
rect 972 3856 980 3864
rect 1132 3876 1140 3884
rect 1212 3876 1220 3884
rect 1324 3876 1332 3884
rect 1340 3876 1348 3884
rect 1404 3876 1412 3884
rect 1420 3876 1428 3884
rect 1532 3876 1540 3884
rect 1596 3876 1604 3884
rect 1660 3876 1668 3884
rect 1724 3876 1732 3884
rect 1788 3876 1796 3884
rect 1852 3876 1860 3884
rect 1916 3876 1924 3884
rect 1980 3876 1988 3884
rect 1996 3876 2004 3884
rect 2108 3876 2116 3884
rect 2172 3876 2180 3884
rect 2188 3876 2196 3884
rect 2332 3876 2340 3884
rect 2396 3876 2404 3884
rect 2460 3876 2468 3884
rect 2524 3876 2532 3884
rect 2572 3876 2580 3884
rect 2588 3876 2596 3884
rect 1148 3856 1156 3864
rect 1276 3856 1284 3864
rect 1340 3856 1348 3864
rect 1404 3856 1412 3864
rect 2316 3856 2324 3864
rect 2380 3856 2388 3864
rect 2444 3856 2452 3864
rect 2508 3856 2516 3864
rect 2572 3856 2580 3864
rect 2652 3876 2660 3884
rect 2716 3876 2724 3884
rect 2762 3876 2770 3884
rect 2796 3876 2804 3884
rect 2844 3876 2852 3884
rect 2908 3876 2916 3884
rect 2956 3876 2964 3884
rect 2972 3876 2980 3884
rect 3036 3876 3044 3884
rect 3070 3876 3078 3884
rect 3100 3876 3108 3884
rect 3196 3876 3204 3884
rect 3228 3876 3236 3884
rect 3292 3876 3300 3884
rect 3420 3876 3428 3884
rect 3484 3876 3492 3884
rect 3596 3876 3604 3884
rect 3692 3876 3700 3884
rect 3756 3876 3764 3884
rect 3884 3876 3892 3884
rect 3996 3876 4004 3884
rect 4124 3876 4132 3884
rect 4172 3876 4180 3884
rect 4316 3876 4324 3884
rect 4460 3876 4468 3884
rect 4540 3876 4548 3884
rect 4556 3876 4564 3884
rect 4620 3876 4628 3884
rect 4732 3876 4740 3884
rect 4748 3876 4756 3884
rect 4812 3876 4820 3884
rect 4892 3876 4900 3884
rect 4956 3876 4964 3884
rect 5116 3876 5124 3884
rect 5132 3876 5140 3884
rect 5196 3876 5204 3884
rect 5308 3876 5316 3884
rect 5324 3876 5332 3884
rect 5388 3876 5396 3884
rect 5452 3876 5460 3884
rect 2700 3856 2708 3864
rect 2812 3856 2820 3864
rect 2828 3856 2836 3864
rect 2892 3856 2900 3864
rect 2956 3856 2964 3864
rect 3020 3856 3028 3864
rect 3084 3856 3092 3864
rect 3212 3856 3220 3864
rect 3276 3856 3284 3864
rect 3404 3856 3412 3864
rect 3468 3856 3476 3864
rect 3708 3856 3716 3864
rect 3772 3856 3780 3864
rect 3900 3856 3908 3864
rect 3916 3856 3924 3864
rect 3980 3856 3988 3864
rect 4108 3856 4116 3864
rect 4300 3856 4308 3864
rect 4476 3856 4484 3864
rect 4876 3856 4884 3864
rect 4940 3856 4948 3864
rect 252 3836 260 3844
rect 780 3836 788 3844
rect 956 3836 964 3844
rect 1164 3836 1172 3844
rect 1468 3836 1476 3844
rect 1548 3836 1556 3844
rect 1676 3836 1684 3844
rect 2044 3836 2052 3844
rect 2060 3836 2068 3844
rect 2124 3836 2132 3844
rect 2236 3836 2244 3844
rect 2252 3836 2260 3844
rect 2492 3836 2500 3844
rect 2620 3836 2628 3844
rect 2748 3836 2756 3844
rect 2876 3836 2884 3844
rect 3660 3836 3668 3844
rect 4092 3836 4100 3844
rect 4220 3836 4228 3844
rect 4284 3836 4292 3844
rect 4364 3836 4372 3844
rect 4668 3836 4676 3844
rect 4860 3836 4868 3844
rect 5052 3836 5060 3844
rect 5244 3836 5252 3844
rect 5260 3836 5268 3844
rect 5436 3836 5444 3844
rect 5516 3836 5524 3844
rect 124 3776 132 3784
rect 188 3776 196 3784
rect 524 3776 532 3784
rect 780 3776 788 3784
rect 844 3776 852 3784
rect 1036 3776 1044 3784
rect 1100 3776 1108 3784
rect 1228 3776 1236 3784
rect 1292 3776 1300 3784
rect 1356 3776 1364 3784
rect 1484 3776 1492 3784
rect 1660 3776 1668 3784
rect 1724 3776 1732 3784
rect 1788 3776 1796 3784
rect 1804 3776 1812 3784
rect 2316 3776 2324 3784
rect 3468 3776 3476 3784
rect 4156 3776 4164 3784
rect 4412 3776 4420 3784
rect 4476 3776 4484 3784
rect 4668 3776 4676 3784
rect 4876 3776 4884 3784
rect 5132 3776 5140 3784
rect 76 3756 84 3764
rect 140 3756 148 3764
rect 252 3756 260 3764
rect 380 3756 388 3764
rect 444 3756 452 3764
rect 508 3756 516 3764
rect 572 3756 580 3764
rect 588 3756 596 3764
rect 700 3756 708 3764
rect 764 3756 772 3764
rect 1020 3756 1028 3764
rect 1212 3756 1220 3764
rect 1596 3756 1604 3764
rect 1612 3756 1620 3764
rect 1868 3756 1876 3764
rect 12 3736 20 3744
rect 76 3736 84 3744
rect 140 3736 148 3744
rect 252 3736 260 3744
rect 330 3736 338 3744
rect 364 3736 372 3744
rect 492 3736 500 3744
rect 556 3736 564 3744
rect 604 3736 612 3744
rect 748 3736 756 3744
rect 828 3736 836 3744
rect 892 3736 900 3744
rect 956 3736 964 3744
rect 1004 3736 1012 3744
rect 1084 3736 1092 3744
rect 1148 3736 1156 3744
rect 1196 3736 1204 3744
rect 1276 3736 1284 3744
rect 1340 3736 1348 3744
rect 1404 3736 1412 3744
rect 1468 3736 1476 3744
rect 1532 3736 1540 3744
rect 1580 3736 1588 3744
rect 1628 3736 1636 3744
rect 1676 3736 1684 3744
rect 1740 3736 1748 3744
rect 1852 3736 1860 3744
rect 1884 3736 1892 3744
rect 2572 3756 2580 3764
rect 2636 3756 2644 3764
rect 2700 3756 2708 3764
rect 2764 3756 2772 3764
rect 2876 3756 2884 3764
rect 2956 3756 2964 3764
rect 3020 3756 3028 3764
rect 3084 3756 3092 3764
rect 3148 3756 3156 3764
rect 3260 3756 3268 3764
rect 3388 3756 3396 3764
rect 3452 3756 3460 3764
rect 3580 3756 3588 3764
rect 3644 3756 3652 3764
rect 3772 3756 3780 3764
rect 3788 3756 3796 3764
rect 3852 3756 3860 3764
rect 4044 3756 4052 3764
rect 4172 3756 4180 3764
rect 4236 3756 4244 3764
rect 4300 3756 4308 3764
rect 4748 3756 4756 3764
rect 4940 3756 4948 3764
rect 5116 3756 5124 3764
rect 5260 3756 5268 3764
rect 5324 3756 5332 3764
rect 5452 3756 5460 3764
rect 1948 3736 1956 3744
rect 2044 3736 2052 3744
rect 2172 3736 2180 3744
rect 2188 3736 2196 3744
rect 2252 3736 2260 3744
rect 2364 3736 2372 3744
rect 2428 3736 2436 3744
rect 2556 3736 2564 3744
rect 2588 3736 2596 3744
rect 2652 3736 2660 3744
rect 2716 3736 2724 3744
rect 2780 3736 2788 3744
rect 2860 3736 2868 3744
rect 2908 3736 2916 3744
rect 2942 3736 2950 3744
rect 2972 3736 2980 3744
rect 3036 3736 3044 3744
rect 3100 3736 3108 3744
rect 3164 3736 3172 3744
rect 3244 3736 3252 3744
rect 3324 3736 3332 3744
rect 3372 3736 3380 3744
rect 3436 3736 3444 3744
rect 3564 3736 3572 3744
rect 3628 3736 3636 3744
rect 3660 3736 3668 3744
rect 3756 3736 3764 3744
rect 3804 3736 3812 3744
rect 3868 3736 3876 3744
rect 4028 3736 4036 3744
rect 4044 3736 4052 3744
rect 4172 3736 4180 3744
rect 4252 3736 4260 3744
rect 4316 3736 4324 3744
rect 4428 3736 4436 3744
rect 4492 3736 4500 3744
rect 4716 3736 4724 3744
rect 4732 3736 4740 3744
rect 4748 3736 4756 3744
rect 4764 3736 4772 3744
rect 4956 3736 4964 3744
rect 5100 3736 5108 3744
rect 5180 3736 5188 3744
rect 5244 3736 5252 3744
rect 5276 3736 5284 3744
rect 5340 3736 5348 3744
rect 5452 3736 5460 3744
rect 60 3716 68 3724
rect 268 3716 276 3724
rect 316 3716 324 3724
rect 908 3716 916 3724
rect 1420 3716 1428 3724
rect 2300 3716 2308 3724
rect 2492 3716 2500 3724
rect 2620 3716 2628 3724
rect 3836 3716 3844 3724
rect 3916 3716 3924 3724
rect 4620 3716 4628 3724
rect 4812 3716 4820 3724
rect 4860 3716 4868 3724
rect 4908 3716 4916 3724
rect 4924 3716 4932 3724
rect 5164 3716 5172 3724
rect 5196 3716 5204 3724
rect 28 3696 36 3704
rect 300 3696 308 3704
rect 396 3696 404 3704
rect 652 3696 660 3704
rect 812 3696 820 3704
rect 876 3696 884 3704
rect 940 3696 948 3704
rect 1068 3696 1076 3704
rect 1132 3696 1140 3704
rect 1148 3696 1156 3704
rect 1260 3696 1268 3704
rect 1324 3696 1332 3704
rect 1388 3696 1396 3704
rect 1452 3696 1460 3704
rect 1516 3696 1524 3704
rect 1676 3696 1684 3704
rect 1756 3696 1764 3704
rect 1836 3696 1844 3704
rect 2028 3696 2036 3704
rect 2076 3696 2084 3704
rect 2172 3696 2180 3704
rect 2204 3696 2212 3704
rect 2268 3696 2276 3704
rect 2348 3696 2356 3704
rect 2428 3696 2436 3704
rect 2476 3696 2484 3704
rect 2540 3696 2548 3704
rect 3068 3696 3076 3704
rect 3324 3696 3332 3704
rect 3516 3696 3524 3704
rect 3596 3696 3604 3704
rect 3676 3696 3684 3704
rect 3724 3696 3732 3704
rect 4012 3696 4020 3704
rect 4124 3696 4132 3704
rect 4220 3696 4228 3704
rect 4284 3696 4292 3704
rect 4380 3696 4388 3704
rect 4444 3696 4452 3704
rect 4508 3696 4516 3704
rect 4556 3696 4564 3704
rect 4636 3696 4644 3704
rect 4684 3696 4692 3704
rect 4796 3696 4804 3704
rect 4844 3696 4852 3704
rect 5020 3696 5028 3704
rect 5228 3696 5236 3704
rect 5308 3696 5316 3704
rect 5388 3696 5396 3704
rect 5436 3696 5444 3704
rect 5516 3696 5524 3704
rect 2252 3676 2260 3684
rect 2428 3676 2436 3684
rect 3964 3676 3972 3684
rect 4364 3676 4372 3684
rect 5068 3676 5076 3684
rect 204 3636 212 3644
rect 636 3636 644 3644
rect 972 3636 980 3644
rect 1548 3636 1556 3644
rect 1980 3636 1988 3644
rect 1996 3636 2004 3644
rect 2108 3636 2116 3644
rect 2124 3636 2132 3644
rect 2380 3636 2388 3644
rect 2684 3636 2692 3644
rect 2748 3636 2756 3644
rect 2812 3636 2820 3644
rect 2828 3636 2836 3644
rect 3004 3636 3012 3644
rect 3132 3636 3140 3644
rect 3196 3636 3204 3644
rect 3212 3636 3220 3644
rect 3276 3636 3284 3644
rect 3340 3636 3348 3644
rect 3404 3636 3412 3644
rect 3708 3636 3716 3644
rect 3980 3636 3988 3644
rect 4604 3636 4612 3644
rect 5052 3636 5060 3644
rect 5580 3636 5588 3644
rect 60 3576 68 3584
rect 140 3576 148 3584
rect 716 3576 724 3584
rect 2764 3576 2772 3584
rect 4492 3576 4500 3584
rect 4556 3576 4564 3584
rect 2556 3556 2564 3564
rect 4428 3556 4436 3564
rect 524 3536 532 3544
rect 780 3536 788 3544
rect 3084 3536 3092 3544
rect 3260 3536 3268 3544
rect 3388 3536 3396 3544
rect 3964 3536 3972 3544
rect 4236 3536 4244 3544
rect 4412 3536 4420 3544
rect 108 3516 116 3524
rect 300 3516 308 3524
rect 380 3516 388 3524
rect 460 3516 468 3524
rect 476 3516 484 3524
rect 556 3516 564 3524
rect 844 3516 852 3524
rect 988 3516 996 3524
rect 1052 3516 1060 3524
rect 1196 3516 1204 3524
rect 1260 3516 1268 3524
rect 1356 3516 1364 3524
rect 1372 3516 1380 3524
rect 1500 3516 1508 3524
rect 1692 3516 1700 3524
rect 1772 3516 1780 3524
rect 1820 3516 1828 3524
rect 1884 3516 1892 3524
rect 1964 3516 1972 3524
rect 2028 3516 2036 3524
rect 2076 3516 2084 3524
rect 2156 3516 2164 3524
rect 2204 3516 2212 3524
rect 2284 3516 2292 3524
rect 2348 3516 2356 3524
rect 2380 3516 2388 3524
rect 2460 3516 2468 3524
rect 2652 3516 2660 3524
rect 2748 3516 2756 3524
rect 2796 3516 2804 3524
rect 3068 3516 3076 3524
rect 3116 3516 3124 3524
rect 3164 3516 3172 3524
rect 3276 3516 3284 3524
rect 3532 3516 3540 3524
rect 3548 3516 3556 3524
rect 3612 3516 3620 3524
rect 3660 3516 3668 3524
rect 3820 3516 3828 3524
rect 4028 3516 4036 3524
rect 4124 3516 4132 3524
rect 4252 3516 4260 3524
rect 4300 3516 4308 3524
rect 4380 3516 4388 3524
rect 4524 3516 4532 3524
rect 4588 3516 4596 3524
rect 4604 3516 4612 3524
rect 4716 3516 4724 3524
rect 4732 3516 4740 3524
rect 4812 3516 4820 3524
rect 5004 3516 5012 3524
rect 5068 3516 5076 3524
rect 5084 3516 5092 3524
rect 5180 3516 5188 3524
rect 5260 3516 5268 3524
rect 5324 3516 5332 3524
rect 5340 3516 5348 3524
rect 5388 3516 5396 3524
rect 5452 3516 5460 3524
rect 5532 3516 5540 3524
rect 76 3496 84 3504
rect 268 3496 276 3504
rect 1612 3496 1620 3504
rect 2316 3496 2324 3504
rect 3148 3496 3156 3504
rect 3468 3496 3476 3504
rect 3660 3496 3668 3504
rect 3772 3496 3780 3504
rect 3916 3496 3924 3504
rect 4108 3496 4116 3504
rect 4748 3496 4756 3504
rect 5436 3496 5444 3504
rect 28 3476 36 3484
rect 124 3476 132 3484
rect 188 3476 196 3484
rect 252 3476 260 3484
rect 316 3476 324 3484
rect 380 3476 388 3484
rect 444 3476 452 3484
rect 460 3476 468 3484
rect 572 3476 580 3484
rect 604 3476 612 3484
rect 12 3456 20 3464
rect 188 3456 196 3464
rect 252 3456 260 3464
rect 588 3456 596 3464
rect 668 3476 676 3484
rect 748 3476 756 3484
rect 812 3476 820 3484
rect 940 3476 948 3484
rect 972 3476 980 3484
rect 1036 3476 1044 3484
rect 1116 3476 1124 3484
rect 1212 3476 1220 3484
rect 1276 3476 1284 3484
rect 1340 3476 1348 3484
rect 1356 3476 1364 3484
rect 1436 3476 1444 3484
rect 1484 3476 1492 3484
rect 1564 3476 1572 3484
rect 1644 3476 1652 3484
rect 1676 3476 1684 3484
rect 1788 3476 1796 3484
rect 1804 3476 1812 3484
rect 1868 3476 1876 3484
rect 1980 3476 1988 3484
rect 2044 3476 2052 3484
rect 2172 3476 2180 3484
rect 2188 3476 2196 3484
rect 2300 3476 2308 3484
rect 2364 3476 2372 3484
rect 2380 3476 2388 3484
rect 2444 3476 2452 3484
rect 2524 3476 2532 3484
rect 764 3456 772 3464
rect 828 3456 836 3464
rect 892 3456 900 3464
rect 956 3456 964 3464
rect 1100 3456 1108 3464
rect 1420 3456 1428 3464
rect 1548 3456 1556 3464
rect 1660 3456 1668 3464
rect 2508 3456 2516 3464
rect 2588 3476 2596 3484
rect 2636 3476 2644 3484
rect 2716 3476 2724 3484
rect 2828 3476 2836 3484
rect 2844 3476 2852 3484
rect 2890 3476 2898 3484
rect 2924 3476 2932 3484
rect 2972 3476 2980 3484
rect 3006 3476 3014 3484
rect 3036 3476 3044 3484
rect 3132 3476 3140 3484
rect 3228 3476 3236 3484
rect 3276 3476 3284 3484
rect 3356 3476 3364 3484
rect 3420 3476 3428 3484
rect 3532 3476 3540 3484
rect 3596 3476 3604 3484
rect 3740 3476 3748 3484
rect 3836 3476 3844 3484
rect 3868 3476 3876 3484
rect 3996 3476 4004 3484
rect 4060 3476 4068 3484
rect 4188 3476 4196 3484
rect 4236 3476 4244 3484
rect 4300 3476 4308 3484
rect 4364 3476 4372 3484
rect 4460 3476 4468 3484
rect 4540 3476 4548 3484
rect 4604 3476 4612 3484
rect 4620 3476 4628 3484
rect 4844 3476 4852 3484
rect 4860 3476 4868 3484
rect 4908 3476 4916 3484
rect 4956 3476 4964 3484
rect 5068 3476 5076 3484
rect 5148 3476 5156 3484
rect 5212 3476 5220 3484
rect 5324 3476 5332 3484
rect 5388 3476 5396 3484
rect 5452 3476 5460 3484
rect 5516 3476 5524 3484
rect 2700 3456 2708 3464
rect 2828 3456 2836 3464
rect 2940 3456 2948 3464
rect 2956 3456 2964 3464
rect 3020 3456 3028 3464
rect 3212 3456 3220 3464
rect 3340 3456 3348 3464
rect 3404 3456 3412 3464
rect 3724 3456 3732 3464
rect 3852 3456 3860 3464
rect 3980 3456 3988 3464
rect 4044 3456 4052 3464
rect 4172 3456 4180 3464
rect 4476 3456 4484 3464
rect 4860 3456 4868 3464
rect 4924 3456 4932 3464
rect 4940 3456 4948 3464
rect 5132 3456 5140 3464
rect 5196 3456 5204 3464
rect 140 3436 148 3444
rect 204 3436 212 3444
rect 332 3436 340 3444
rect 396 3436 404 3444
rect 508 3436 516 3444
rect 700 3436 708 3444
rect 1020 3436 1028 3444
rect 1084 3436 1092 3444
rect 1148 3436 1156 3444
rect 1164 3436 1172 3444
rect 1228 3436 1236 3444
rect 1292 3436 1300 3444
rect 1404 3436 1412 3444
rect 1468 3436 1476 3444
rect 1532 3436 1540 3444
rect 1596 3436 1604 3444
rect 1724 3436 1732 3444
rect 1740 3436 1748 3444
rect 1852 3436 1860 3444
rect 1916 3436 1924 3444
rect 1932 3436 1940 3444
rect 1996 3436 2004 3444
rect 2108 3436 2116 3444
rect 2124 3436 2132 3444
rect 2236 3436 2244 3444
rect 2252 3436 2260 3444
rect 2428 3436 2436 3444
rect 2492 3436 2500 3444
rect 2620 3436 2628 3444
rect 2684 3436 2692 3444
rect 2876 3436 2884 3444
rect 3196 3436 3204 3444
rect 3324 3436 3332 3444
rect 3580 3436 3588 3444
rect 3644 3436 3652 3444
rect 3708 3436 3716 3444
rect 3788 3436 3796 3444
rect 4156 3436 4164 3444
rect 4284 3436 4292 3444
rect 4348 3436 4356 3444
rect 4668 3436 4676 3444
rect 4684 3436 4692 3444
rect 4796 3436 4804 3444
rect 4988 3436 4996 3444
rect 5116 3436 5124 3444
rect 5372 3436 5380 3444
rect 5500 3436 5508 3444
rect 5564 3436 5572 3444
rect 12 3376 20 3384
rect 332 3376 340 3384
rect 588 3376 596 3384
rect 780 3376 788 3384
rect 844 3376 852 3384
rect 908 3376 916 3384
rect 972 3376 980 3384
rect 1484 3376 1492 3384
rect 1548 3376 1556 3384
rect 1932 3376 1940 3384
rect 2060 3376 2068 3384
rect 2188 3376 2196 3384
rect 2252 3376 2260 3384
rect 2444 3376 2452 3384
rect 2636 3376 2644 3384
rect 2828 3376 2836 3384
rect 3148 3376 3156 3384
rect 3468 3376 3476 3384
rect 3532 3376 3540 3384
rect 3836 3376 3844 3384
rect 4236 3376 4244 3384
rect 4300 3376 4308 3384
rect 4540 3376 4548 3384
rect 4556 3376 4564 3384
rect 4748 3376 4756 3384
rect 4876 3376 4884 3384
rect 4940 3376 4948 3384
rect 5244 3376 5252 3384
rect 5308 3376 5316 3384
rect 5452 3376 5460 3384
rect 124 3356 132 3364
rect 188 3356 196 3364
rect 252 3356 260 3364
rect 60 3336 68 3344
rect 172 3336 180 3344
rect 252 3336 260 3344
rect 316 3336 324 3344
rect 364 3336 372 3344
rect 396 3356 404 3364
rect 508 3356 516 3364
rect 396 3336 404 3344
rect 412 3336 420 3344
rect 446 3336 454 3344
rect 492 3336 500 3344
rect 572 3336 580 3344
rect 636 3336 644 3344
rect 684 3336 692 3344
rect 764 3356 772 3364
rect 1036 3356 1044 3364
rect 1148 3356 1156 3364
rect 748 3336 756 3344
rect 828 3336 836 3344
rect 892 3336 900 3344
rect 956 3336 964 3344
rect 1020 3336 1028 3344
rect 1052 3336 1060 3344
rect 1132 3336 1140 3344
rect 1180 3336 1188 3344
rect 1292 3356 1300 3364
rect 1404 3356 1412 3364
rect 1612 3356 1620 3364
rect 1788 3356 1796 3364
rect 1804 3356 1812 3364
rect 1244 3336 1252 3344
rect 1308 3336 1316 3344
rect 1404 3336 1412 3344
rect 1468 3336 1476 3344
rect 1532 3336 1540 3344
rect 1596 3336 1604 3344
rect 1628 3336 1636 3344
rect 1738 3336 1746 3344
rect 1772 3336 1780 3344
rect 1804 3336 1812 3344
rect 2044 3356 2052 3364
rect 2172 3356 2180 3364
rect 2316 3356 2324 3364
rect 2428 3356 2436 3364
rect 2556 3356 2564 3364
rect 2620 3356 2628 3364
rect 2700 3356 2708 3364
rect 2812 3356 2820 3364
rect 2956 3356 2964 3364
rect 3020 3356 3028 3364
rect 3084 3356 3092 3364
rect 3212 3356 3220 3364
rect 3276 3356 3284 3364
rect 3340 3356 3348 3364
rect 3516 3356 3524 3364
rect 3708 3356 3716 3364
rect 3724 3356 3732 3364
rect 3900 3356 3908 3364
rect 4092 3356 4100 3364
rect 1884 3336 1892 3344
rect 1980 3336 1988 3344
rect 2028 3336 2036 3344
rect 2108 3336 2116 3344
rect 2156 3336 2164 3344
rect 2300 3336 2308 3344
rect 2332 3336 2340 3344
rect 2378 3336 2386 3344
rect 2412 3336 2420 3344
rect 2492 3336 2500 3344
rect 2540 3336 2548 3344
rect 2620 3336 2628 3344
rect 2716 3336 2724 3344
rect 2750 3336 2758 3344
rect 2796 3336 2804 3344
rect 2924 3336 2932 3344
rect 2956 3336 2964 3344
rect 3036 3336 3044 3344
rect 3100 3336 3108 3344
rect 3134 3336 3142 3344
rect 3196 3336 3204 3344
rect 3228 3336 3236 3344
rect 3292 3336 3300 3344
rect 3356 3336 3364 3344
rect 3500 3336 3508 3344
rect 3580 3336 3588 3344
rect 3644 3336 3652 3344
rect 3692 3336 3700 3344
rect 3740 3336 3748 3344
rect 3884 3336 3892 3344
rect 3964 3336 3972 3344
rect 4042 3336 4050 3344
rect 4076 3336 4084 3344
rect 4172 3356 4180 3364
rect 4412 3356 4420 3364
rect 4428 3356 4436 3364
rect 4668 3356 4676 3364
rect 4732 3356 4740 3364
rect 4860 3356 4868 3364
rect 5004 3356 5012 3364
rect 5068 3356 5076 3364
rect 5132 3356 5140 3364
rect 5388 3356 5396 3364
rect 4124 3336 4132 3344
rect 4172 3336 4180 3344
rect 4188 3336 4196 3344
rect 4284 3336 4292 3344
rect 4396 3336 4404 3344
rect 4444 3336 4452 3344
rect 4492 3336 4500 3344
rect 4652 3336 4660 3344
rect 4716 3336 4724 3344
rect 4844 3336 4852 3344
rect 4924 3336 4932 3344
rect 4988 3336 4996 3344
rect 5020 3336 5028 3344
rect 5084 3336 5092 3344
rect 5148 3336 5156 3344
rect 5196 3336 5204 3344
rect 5388 3336 5396 3344
rect 5404 3336 5412 3344
rect 5438 3336 5446 3344
rect 5500 3336 5508 3344
rect 5516 3336 5524 3344
rect 268 3316 276 3324
rect 524 3316 532 3324
rect 556 3316 564 3324
rect 1356 3316 1364 3324
rect 1420 3316 1428 3324
rect 1676 3316 1684 3324
rect 1724 3316 1732 3324
rect 2684 3316 2692 3324
rect 2764 3316 2772 3324
rect 2876 3316 2884 3324
rect 3324 3316 3332 3324
rect 3404 3316 3412 3324
rect 3804 3316 3812 3324
rect 3852 3316 3860 3324
rect 3996 3316 4004 3324
rect 4796 3316 4804 3324
rect 5260 3316 5268 3324
rect 5324 3316 5332 3324
rect 60 3296 68 3304
rect 300 3296 308 3304
rect 572 3296 580 3304
rect 620 3296 628 3304
rect 812 3296 820 3304
rect 876 3296 884 3304
rect 940 3296 948 3304
rect 1004 3296 1012 3304
rect 1452 3296 1460 3304
rect 1516 3296 1524 3304
rect 1580 3296 1588 3304
rect 1708 3296 1716 3304
rect 1964 3296 1972 3304
rect 2092 3296 2100 3304
rect 2220 3296 2228 3304
rect 2284 3296 2292 3304
rect 2476 3296 2484 3304
rect 2572 3296 2580 3304
rect 2668 3296 2676 3304
rect 2860 3296 2868 3304
rect 3196 3296 3204 3304
rect 3260 3296 3268 3304
rect 3564 3296 3572 3304
rect 3916 3296 3924 3304
rect 3948 3296 3956 3304
rect 4268 3296 4276 3304
rect 4332 3296 4340 3304
rect 4476 3296 4484 3304
rect 4508 3296 4516 3304
rect 4588 3296 4596 3304
rect 4684 3296 4692 3304
rect 4908 3296 4916 3304
rect 4972 3296 4980 3304
rect 5052 3296 5060 3304
rect 5196 3296 5204 3304
rect 5212 3296 5220 3304
rect 5276 3296 5284 3304
rect 5356 3296 5364 3304
rect 5484 3296 5492 3304
rect 5532 3296 5540 3304
rect 1340 3256 1348 3264
rect 76 3236 84 3244
rect 204 3236 212 3244
rect 460 3236 468 3244
rect 652 3236 660 3244
rect 1084 3236 1092 3244
rect 1100 3236 1108 3244
rect 1276 3236 1284 3244
rect 1660 3236 1668 3244
rect 1916 3236 1924 3244
rect 1996 3236 2004 3244
rect 2124 3236 2132 3244
rect 2364 3236 2372 3244
rect 2508 3236 2516 3244
rect 2892 3236 2900 3244
rect 3004 3236 3012 3244
rect 3068 3236 3076 3244
rect 3452 3236 3460 3244
rect 3596 3236 3604 3244
rect 4028 3236 4036 3244
rect 4220 3236 4228 3244
rect 4364 3236 4372 3244
rect 4556 3236 4564 3244
rect 5116 3236 5124 3244
rect 5580 3236 5588 3244
rect 396 3176 404 3184
rect 700 3176 708 3184
rect 1724 3176 1732 3184
rect 2364 3176 2372 3184
rect 4284 3176 4292 3184
rect 5180 3176 5188 3184
rect 1996 3156 2004 3164
rect 2940 3156 2948 3164
rect 3644 3156 3652 3164
rect 5308 3156 5316 3164
rect 5564 3156 5572 3164
rect 1020 3136 1028 3144
rect 1356 3136 1364 3144
rect 1788 3136 1796 3144
rect 2124 3136 2132 3144
rect 2812 3136 2820 3144
rect 3468 3136 3476 3144
rect 3852 3136 3860 3144
rect 236 3116 244 3124
rect 332 3116 340 3124
rect 476 3116 484 3124
rect 524 3116 532 3124
rect 588 3116 596 3124
rect 668 3116 676 3124
rect 716 3116 724 3124
rect 908 3116 916 3124
rect 988 3116 996 3124
rect 1052 3116 1060 3124
rect 1196 3116 1204 3124
rect 1260 3116 1268 3124
rect 1516 3116 1524 3124
rect 1580 3116 1588 3124
rect 1628 3116 1636 3124
rect 1772 3116 1780 3124
rect 1836 3116 1844 3124
rect 2108 3116 2116 3124
rect 2188 3116 2196 3124
rect 2252 3116 2260 3124
rect 2396 3116 2404 3124
rect 2460 3116 2468 3124
rect 2540 3116 2548 3124
rect 2668 3116 2676 3124
rect 2732 3116 2740 3124
rect 2892 3116 2900 3124
rect 2972 3116 2980 3124
rect 3020 3116 3028 3124
rect 3036 3116 3044 3124
rect 3116 3116 3124 3124
rect 3132 3116 3140 3124
rect 3180 3116 3188 3124
rect 3196 3116 3204 3124
rect 3340 3116 3348 3124
rect 3452 3116 3460 3124
rect 3548 3116 3556 3124
rect 3884 3116 3892 3124
rect 3996 3116 4004 3124
rect 4044 3116 4052 3124
rect 4060 3116 4068 3124
rect 4124 3116 4132 3124
rect 4172 3116 4180 3124
rect 4364 3116 4372 3124
rect 4380 3116 4388 3124
rect 4588 3116 4596 3124
rect 4700 3116 4708 3124
rect 4892 3116 4900 3124
rect 4924 3116 4932 3124
rect 4972 3116 4980 3124
rect 5052 3116 5060 3124
rect 5100 3116 5108 3124
rect 5196 3116 5204 3124
rect 5340 3116 5348 3124
rect 5404 3116 5412 3124
rect 5452 3116 5460 3124
rect 5468 3116 5476 3124
rect 5532 3116 5540 3124
rect 508 3096 516 3104
rect 1100 3096 1108 3104
rect 1212 3096 1220 3104
rect 1276 3096 1284 3104
rect 2444 3096 2452 3104
rect 2700 3096 2708 3104
rect 3068 3096 3076 3104
rect 3260 3096 3268 3104
rect 4172 3096 4180 3104
rect 4236 3096 4244 3104
rect 4252 3096 4260 3104
rect 4348 3096 4356 3104
rect 4476 3096 4484 3104
rect 4524 3096 4532 3104
rect 4540 3096 4548 3104
rect 4748 3096 4756 3104
rect 4860 3096 4868 3104
rect 4988 3096 4996 3104
rect 5196 3096 5204 3104
rect 172 3076 180 3084
rect 188 3076 196 3084
rect 252 3076 260 3084
rect 300 3076 308 3084
rect 380 3076 388 3084
rect 428 3076 436 3084
rect 460 3076 468 3084
rect 556 3076 564 3084
rect 636 3076 644 3084
rect 652 3076 660 3084
rect 812 3076 820 3084
rect 60 3056 68 3064
rect 124 3056 132 3064
rect 188 3056 196 3064
rect 316 3056 324 3064
rect 380 3056 388 3064
rect 444 3056 452 3064
rect 572 3056 580 3064
rect 636 3056 644 3064
rect 764 3056 772 3064
rect 876 3076 884 3084
rect 956 3076 964 3084
rect 972 3076 980 3084
rect 1036 3076 1044 3084
rect 1132 3076 1140 3084
rect 1324 3076 1332 3084
rect 1388 3076 1396 3084
rect 892 3056 900 3064
rect 956 3056 964 3064
rect 1148 3056 1156 3064
rect 1340 3056 1348 3064
rect 1452 3076 1460 3084
rect 1532 3076 1540 3084
rect 1596 3076 1604 3084
rect 1612 3076 1620 3084
rect 1692 3076 1700 3084
rect 1788 3076 1796 3084
rect 1852 3076 1860 3084
rect 1884 3076 1892 3084
rect 1932 3076 1940 3084
rect 2028 3076 2036 3084
rect 2076 3076 2084 3084
rect 2156 3076 2164 3084
rect 2188 3076 2196 3084
rect 2252 3076 2260 3084
rect 2332 3076 2340 3084
rect 2380 3076 2388 3084
rect 2556 3076 2564 3084
rect 2604 3076 2612 3084
rect 2684 3076 2692 3084
rect 2748 3076 2756 3084
rect 2780 3076 2788 3084
rect 2844 3076 2852 3084
rect 2956 3076 2964 3084
rect 3020 3076 3028 3084
rect 3132 3076 3140 3084
rect 3196 3076 3204 3084
rect 3308 3076 3316 3084
rect 3372 3076 3380 3084
rect 3420 3076 3428 3084
rect 3500 3076 3508 3084
rect 3532 3076 3540 3084
rect 3596 3076 3604 3084
rect 3676 3076 3684 3084
rect 3740 3076 3748 3084
rect 3788 3076 3796 3084
rect 3900 3076 3908 3084
rect 4044 3076 4052 3084
rect 4108 3076 4116 3084
rect 4364 3076 4372 3084
rect 4444 3076 4452 3084
rect 4604 3076 4612 3084
rect 4636 3076 4644 3084
rect 4684 3076 4692 3084
rect 4780 3076 4788 3084
rect 4828 3076 4836 3084
rect 4876 3076 4884 3084
rect 5020 3076 5028 3084
rect 5116 3076 5124 3084
rect 5148 3076 5156 3084
rect 5276 3076 5284 3084
rect 5324 3076 5332 3084
rect 5388 3076 5396 3084
rect 5452 3076 5460 3084
rect 5516 3076 5524 3084
rect 1468 3056 1476 3064
rect 1676 3056 1684 3064
rect 1868 3056 1876 3064
rect 2044 3056 2052 3064
rect 2060 3056 2068 3064
rect 2172 3056 2180 3064
rect 2316 3056 2324 3064
rect 2620 3056 2628 3064
rect 2764 3056 2772 3064
rect 2828 3056 2836 3064
rect 3324 3056 3332 3064
rect 3388 3056 3396 3064
rect 3404 3056 3412 3064
rect 3516 3056 3524 3064
rect 3660 3056 3668 3064
rect 3724 3056 3732 3064
rect 3916 3056 3924 3064
rect 4428 3056 4436 3064
rect 4620 3056 4628 3064
rect 4796 3056 4804 3064
rect 4812 3056 4820 3064
rect 5004 3056 5012 3064
rect 5132 3056 5140 3064
rect 5260 3056 5268 3064
rect 12 3036 20 3044
rect 204 3036 212 3044
rect 268 3036 276 3044
rect 1020 3036 1028 3044
rect 1084 3036 1092 3044
rect 1164 3036 1172 3044
rect 1228 3036 1236 3044
rect 1292 3036 1300 3044
rect 1484 3036 1492 3044
rect 1548 3036 1556 3044
rect 1660 3036 1668 3044
rect 1740 3036 1748 3044
rect 1980 3036 1988 3044
rect 2236 3036 2244 3044
rect 2300 3036 2308 3044
rect 2428 3036 2436 3044
rect 2492 3036 2500 3044
rect 2508 3036 2516 3044
rect 2572 3036 2580 3044
rect 2636 3036 2644 3044
rect 3084 3036 3092 3044
rect 3708 3036 3716 3044
rect 3836 3036 3844 3044
rect 4092 3036 4100 3044
rect 4156 3036 4164 3044
rect 4220 3036 4228 3044
rect 4300 3036 4308 3044
rect 4412 3036 4420 3044
rect 4492 3036 4500 3044
rect 4556 3036 4564 3044
rect 4668 3036 4676 3044
rect 4732 3036 4740 3044
rect 4940 3036 4948 3044
rect 5068 3036 5076 3044
rect 5244 3036 5252 3044
rect 5372 3036 5380 3044
rect 5500 3036 5508 3044
rect 188 2976 196 2984
rect 316 2976 324 2984
rect 380 2976 388 2984
rect 700 2976 708 2984
rect 780 2976 788 2984
rect 908 2976 916 2984
rect 972 2976 980 2984
rect 1084 2976 1092 2984
rect 1228 2976 1236 2984
rect 1404 2976 1412 2984
rect 1852 2976 1860 2984
rect 1868 2976 1876 2984
rect 1980 2976 1988 2984
rect 2188 2976 2196 2984
rect 2252 2976 2260 2984
rect 2428 2976 2436 2984
rect 2684 2976 2692 2984
rect 2764 2976 2772 2984
rect 2956 2976 2964 2984
rect 3084 2976 3092 2984
rect 3260 2976 3268 2984
rect 3276 2976 3284 2984
rect 3980 2976 3988 2984
rect 4092 2976 4100 2984
rect 4364 2976 4372 2984
rect 4492 2976 4500 2984
rect 4556 2976 4564 2984
rect 4684 2976 4692 2984
rect 4940 2976 4948 2984
rect 5116 2976 5124 2984
rect 5180 2976 5188 2984
rect 5308 2976 5316 2984
rect 5372 2976 5380 2984
rect 5564 2976 5572 2984
rect 124 2956 132 2964
rect 204 2956 212 2964
rect 396 2956 404 2964
rect 524 2956 532 2964
rect 588 2956 596 2964
rect 716 2956 724 2964
rect 892 2956 900 2964
rect 1100 2956 1108 2964
rect 1212 2956 1220 2964
rect 1276 2956 1284 2964
rect 1292 2956 1300 2964
rect 1420 2956 1428 2964
rect 12 2936 20 2944
rect 108 2936 116 2944
rect 140 2936 148 2944
rect 220 2936 228 2944
rect 268 2936 276 2944
rect 332 2936 340 2944
rect 412 2936 420 2944
rect 508 2936 516 2944
rect 540 2936 548 2944
rect 604 2936 612 2944
rect 652 2936 660 2944
rect 732 2936 740 2944
rect 828 2936 836 2944
rect 876 2936 884 2944
rect 956 2936 964 2944
rect 1020 2936 1028 2944
rect 1036 2936 1044 2944
rect 1116 2936 1124 2944
rect 1196 2936 1204 2944
rect 1260 2936 1268 2944
rect 1308 2936 1316 2944
rect 1356 2936 1364 2944
rect 1436 2936 1444 2944
rect 1548 2956 1556 2964
rect 1612 2956 1620 2964
rect 1724 2956 1732 2964
rect 1996 2956 2004 2964
rect 2060 2956 2068 2964
rect 2172 2956 2180 2964
rect 2300 2956 2308 2964
rect 2364 2956 2372 2964
rect 2508 2956 2516 2964
rect 1500 2936 1508 2944
rect 1564 2936 1572 2944
rect 1628 2936 1636 2944
rect 1674 2936 1682 2944
rect 1724 2936 1732 2944
rect 1788 2936 1796 2944
rect 1804 2936 1812 2944
rect 1916 2936 1924 2944
rect 1932 2936 1940 2944
rect 2012 2936 2020 2944
rect 2076 2936 2084 2944
rect 2156 2936 2164 2944
rect 2236 2936 2244 2944
rect 2284 2936 2292 2944
rect 2348 2936 2356 2944
rect 2364 2936 2372 2944
rect 2444 2936 2452 2944
rect 2508 2936 2516 2944
rect 2748 2956 2756 2964
rect 2876 2956 2884 2964
rect 2940 2956 2948 2964
rect 3004 2956 3012 2964
rect 3068 2956 3076 2964
rect 3148 2956 3156 2964
rect 3212 2956 3220 2964
rect 3340 2956 3348 2964
rect 3452 2956 3460 2964
rect 3580 2956 3588 2964
rect 3708 2956 3716 2964
rect 4796 2956 4804 2964
rect 4988 2956 4996 2964
rect 5004 2956 5012 2964
rect 5324 2956 5332 2964
rect 2588 2936 2596 2944
rect 2636 2936 2644 2944
rect 2732 2936 2740 2944
rect 2860 2936 2868 2944
rect 2924 2936 2932 2944
rect 2988 2936 2996 2944
rect 3052 2936 3060 2944
rect 3164 2936 3172 2944
rect 3228 2936 3236 2944
rect 3340 2936 3348 2944
rect 3356 2936 3364 2944
rect 3436 2936 3444 2944
rect 3468 2936 3476 2944
rect 3564 2936 3572 2944
rect 3692 2936 3700 2944
rect 3724 2936 3732 2944
rect 3836 2936 3844 2944
rect 3964 2936 3972 2944
rect 4028 2936 4036 2944
rect 4044 2936 4052 2944
rect 4108 2936 4116 2944
rect 4284 2936 4292 2944
rect 4300 2936 4308 2944
rect 4412 2936 4420 2944
rect 4428 2936 4436 2944
rect 4540 2936 4548 2944
rect 4604 2936 4612 2944
rect 4668 2936 4676 2944
rect 4732 2936 4740 2944
rect 4780 2936 4788 2944
rect 4860 2936 4868 2944
rect 4972 2936 4980 2944
rect 5020 2936 5028 2944
rect 5054 2936 5062 2944
rect 5196 2936 5204 2944
rect 5260 2936 5268 2944
rect 5340 2936 5348 2944
rect 5516 2936 5524 2944
rect 60 2916 68 2924
rect 460 2916 468 2924
rect 1340 2916 1348 2924
rect 1740 2916 1748 2924
rect 1948 2916 1956 2924
rect 2492 2916 2500 2924
rect 2812 2916 2820 2924
rect 3132 2916 3140 2924
rect 3596 2916 3604 2924
rect 3644 2916 3652 2924
rect 4156 2916 4164 2924
rect 4220 2916 4228 2924
rect 4348 2916 4356 2924
rect 4476 2916 4484 2924
rect 4748 2916 4756 2924
rect 4876 2916 4884 2924
rect 4892 2916 4900 2924
rect 5068 2916 5076 2924
rect 5132 2916 5140 2924
rect 5244 2916 5252 2924
rect 5500 2916 5508 2924
rect 28 2896 36 2904
rect 76 2896 84 2904
rect 156 2896 164 2904
rect 268 2896 276 2904
rect 284 2896 292 2904
rect 348 2896 356 2904
rect 508 2896 516 2904
rect 812 2896 820 2904
rect 940 2896 948 2904
rect 1020 2896 1028 2904
rect 1052 2896 1060 2904
rect 1372 2896 1380 2904
rect 1772 2896 1780 2904
rect 1804 2896 1812 2904
rect 1900 2896 1908 2904
rect 2108 2896 2116 2904
rect 2220 2896 2228 2904
rect 2396 2896 2404 2904
rect 2460 2896 2468 2904
rect 2652 2896 2660 2904
rect 2796 2896 2804 2904
rect 2892 2896 2900 2904
rect 3020 2896 3028 2904
rect 3116 2896 3124 2904
rect 3196 2896 3204 2904
rect 3308 2896 3316 2904
rect 3388 2896 3396 2904
rect 3484 2896 3492 2904
rect 3532 2896 3540 2904
rect 3612 2896 3620 2904
rect 3660 2896 3668 2904
rect 3740 2896 3748 2904
rect 3820 2896 3828 2904
rect 3884 2896 3892 2904
rect 3948 2896 3956 2904
rect 4012 2896 4020 2904
rect 4060 2896 4068 2904
rect 4124 2896 4132 2904
rect 4188 2896 4196 2904
rect 4268 2896 4276 2904
rect 4316 2896 4324 2904
rect 4396 2896 4404 2904
rect 4444 2896 4452 2904
rect 4524 2896 4532 2904
rect 4652 2896 4660 2904
rect 4716 2896 4724 2904
rect 4844 2896 4852 2904
rect 5084 2896 5092 2904
rect 5148 2896 5156 2904
rect 5212 2896 5220 2904
rect 5276 2896 5284 2904
rect 5404 2896 5412 2904
rect 5452 2896 5460 2904
rect 5532 2896 5540 2904
rect 1148 2876 1156 2884
rect 1356 2876 1364 2884
rect 2700 2876 2708 2884
rect 3404 2856 3412 2864
rect 3772 2856 3780 2864
rect 444 2836 452 2844
rect 572 2836 580 2844
rect 764 2836 772 2844
rect 844 2836 852 2844
rect 1164 2836 1172 2844
rect 1532 2836 1540 2844
rect 1596 2836 1604 2844
rect 1660 2836 1668 2844
rect 2044 2836 2052 2844
rect 2124 2836 2132 2844
rect 2316 2836 2324 2844
rect 2620 2836 2628 2844
rect 2828 2836 2836 2844
rect 2956 2836 2964 2844
rect 3516 2836 3524 2844
rect 3788 2836 3796 2844
rect 3852 2836 3860 2844
rect 4236 2836 4244 2844
rect 4812 2836 4820 2844
rect 4924 2836 4932 2844
rect 1212 2776 1220 2784
rect 1740 2776 1748 2784
rect 2044 2776 2052 2784
rect 2252 2776 2260 2784
rect 844 2756 852 2764
rect 1612 2756 1620 2764
rect 3452 2756 3460 2764
rect 4156 2756 4164 2764
rect 4428 2756 4436 2764
rect 156 2716 164 2724
rect 300 2716 308 2724
rect 364 2716 372 2724
rect 492 2716 500 2724
rect 540 2716 548 2724
rect 604 2716 612 2724
rect 780 2716 788 2724
rect 1004 2716 1012 2724
rect 1068 2716 1076 2724
rect 1436 2716 1444 2724
rect 1500 2716 1508 2724
rect 1564 2716 1572 2724
rect 1644 2716 1652 2724
rect 1772 2716 1780 2724
rect 1820 2716 1828 2724
rect 1900 2716 1908 2724
rect 2012 2716 2020 2724
rect 2204 2716 2212 2724
rect 2236 2716 2244 2724
rect 2332 2716 2340 2724
rect 2428 2716 2436 2724
rect 2476 2716 2484 2724
rect 2652 2716 2660 2724
rect 2844 2716 2852 2724
rect 2892 2716 2900 2724
rect 2924 2716 2932 2724
rect 2988 2716 2996 2724
rect 3004 2716 3012 2724
rect 3100 2716 3108 2724
rect 3228 2716 3236 2724
rect 3276 2716 3284 2724
rect 3340 2716 3348 2724
rect 3420 2716 3428 2724
rect 3548 2716 3556 2724
rect 3596 2716 3604 2724
rect 3692 2716 3700 2724
rect 3772 2716 3780 2724
rect 3916 2716 3924 2724
rect 3996 2716 4004 2724
rect 4092 2716 4100 2724
rect 4124 2716 4132 2724
rect 4204 2716 4212 2724
rect 4252 2716 4260 2724
rect 4316 2716 4324 2724
rect 4396 2716 4404 2724
rect 4460 2716 4468 2724
rect 4508 2716 4516 2724
rect 4588 2716 4596 2724
rect 4684 2716 4692 2724
rect 4796 2716 4804 2724
rect 4828 2716 4836 2724
rect 4876 2716 4884 2724
rect 4908 2716 4916 2724
rect 4924 2716 4932 2724
rect 5004 2716 5012 2724
rect 5020 2716 5028 2724
rect 5212 2716 5220 2724
rect 5276 2716 5284 2724
rect 5340 2716 5348 2724
rect 5404 2716 5412 2724
rect 5452 2716 5460 2724
rect 5468 2716 5476 2724
rect 5516 2716 5524 2724
rect 332 2696 340 2704
rect 572 2696 580 2704
rect 636 2696 644 2704
rect 1100 2696 1108 2704
rect 1932 2696 1940 2704
rect 2444 2696 2452 2704
rect 2940 2696 2948 2704
rect 3468 2696 3476 2704
rect 3708 2696 3716 2704
rect 3852 2696 3860 2704
rect 3964 2696 3972 2704
rect 4348 2696 4356 2704
rect 4556 2696 4564 2704
rect 4620 2696 4628 2704
rect 4860 2696 4868 2704
rect 5244 2696 5252 2704
rect 5372 2696 5380 2704
rect 28 2676 36 2684
rect 12 2656 20 2664
rect 92 2676 100 2684
rect 140 2676 148 2684
rect 220 2676 228 2684
rect 316 2676 324 2684
rect 380 2676 388 2684
rect 412 2676 420 2684
rect 508 2676 516 2684
rect 524 2676 532 2684
rect 588 2676 596 2684
rect 652 2676 660 2684
rect 732 2676 740 2684
rect 780 2676 788 2684
rect 876 2676 884 2684
rect 940 2676 948 2684
rect 1020 2676 1028 2684
rect 1084 2676 1092 2684
rect 1132 2676 1140 2684
rect 1148 2676 1156 2684
rect 1226 2676 1234 2684
rect 1260 2676 1268 2684
rect 1324 2676 1332 2684
rect 1372 2676 1380 2684
rect 1420 2676 1428 2684
rect 1484 2676 1492 2684
rect 1548 2676 1556 2684
rect 1660 2676 1668 2684
rect 1692 2676 1700 2684
rect 1788 2676 1796 2684
rect 1804 2676 1812 2684
rect 1916 2676 1924 2684
rect 1964 2676 1972 2684
rect 1996 2676 2004 2684
rect 2092 2676 2100 2684
rect 2140 2676 2148 2684
rect 2188 2676 2196 2684
rect 2284 2676 2292 2684
rect 2316 2676 2324 2684
rect 2380 2676 2388 2684
rect 2492 2676 2500 2684
rect 2508 2676 2516 2684
rect 2572 2676 2580 2684
rect 2636 2676 2644 2684
rect 2732 2676 2740 2684
rect 204 2656 212 2664
rect 396 2656 404 2664
rect 652 2656 660 2664
rect 716 2656 724 2664
rect 892 2656 900 2664
rect 956 2656 964 2664
rect 1148 2656 1156 2664
rect 1164 2656 1172 2664
rect 1276 2656 1284 2664
rect 1340 2656 1348 2664
rect 1356 2656 1364 2664
rect 1676 2656 1684 2664
rect 1980 2656 1988 2664
rect 2108 2656 2116 2664
rect 2124 2656 2132 2664
rect 2300 2656 2308 2664
rect 2380 2656 2388 2664
rect 2508 2656 2516 2664
rect 2572 2656 2580 2664
rect 2780 2676 2788 2684
rect 3004 2676 3012 2684
rect 3052 2676 3060 2684
rect 3084 2676 3092 2684
rect 3164 2676 3172 2684
rect 3308 2676 3316 2684
rect 3340 2676 3348 2684
rect 3404 2676 3412 2684
rect 3500 2676 3508 2684
rect 3516 2676 3524 2684
rect 3628 2676 3636 2684
rect 3740 2676 3748 2684
rect 3804 2676 3812 2684
rect 3916 2676 3924 2684
rect 3980 2676 3988 2684
rect 4092 2676 4100 2684
rect 4108 2676 4116 2684
rect 4220 2676 4228 2684
rect 4236 2676 4244 2684
rect 4300 2676 4308 2684
rect 4412 2676 4420 2684
rect 4492 2676 4500 2684
rect 4604 2676 4612 2684
rect 4652 2676 4660 2684
rect 4684 2676 4692 2684
rect 4764 2676 4772 2684
rect 4924 2676 4932 2684
rect 4940 2676 4948 2684
rect 5004 2676 5012 2684
rect 5100 2676 5108 2684
rect 5148 2676 5156 2684
rect 5260 2676 5268 2684
rect 5324 2676 5332 2684
rect 5388 2676 5396 2684
rect 5452 2676 5460 2684
rect 5516 2676 5524 2684
rect 2764 2656 2772 2664
rect 3068 2656 3076 2664
rect 3148 2656 3156 2664
rect 3324 2656 3332 2664
rect 3516 2656 3524 2664
rect 3644 2656 3652 2664
rect 3724 2656 3732 2664
rect 3788 2656 3796 2664
rect 4668 2656 4676 2664
rect 4748 2656 4756 2664
rect 5116 2656 5124 2664
rect 5132 2656 5140 2664
rect 124 2636 132 2644
rect 188 2636 196 2644
rect 252 2636 260 2644
rect 268 2636 276 2644
rect 444 2636 452 2644
rect 460 2636 468 2644
rect 700 2636 708 2644
rect 764 2636 772 2644
rect 828 2636 836 2644
rect 908 2636 916 2644
rect 972 2636 980 2644
rect 1036 2636 1044 2644
rect 1292 2636 1300 2644
rect 1404 2636 1412 2644
rect 1468 2636 1476 2644
rect 1532 2636 1540 2644
rect 1596 2636 1604 2644
rect 1724 2636 1732 2644
rect 1852 2636 1860 2644
rect 1868 2636 1876 2644
rect 2044 2636 2052 2644
rect 2060 2636 2068 2644
rect 2172 2636 2180 2644
rect 2364 2636 2372 2644
rect 2556 2636 2564 2644
rect 2620 2636 2628 2644
rect 2684 2636 2692 2644
rect 2700 2636 2708 2644
rect 2876 2636 2884 2644
rect 2956 2636 2964 2644
rect 3132 2636 3140 2644
rect 3260 2636 3268 2644
rect 3388 2636 3396 2644
rect 3580 2636 3588 2644
rect 3660 2636 3668 2644
rect 3900 2636 3908 2644
rect 4028 2636 4036 2644
rect 4044 2636 4052 2644
rect 4172 2636 4180 2644
rect 4284 2636 4292 2644
rect 4364 2636 4372 2644
rect 4540 2636 4548 2644
rect 4732 2636 4740 2644
rect 5052 2636 5060 2644
rect 5068 2636 5076 2644
rect 5308 2636 5316 2644
rect 5500 2636 5508 2644
rect 5580 2636 5588 2644
rect 140 2576 148 2584
rect 204 2576 212 2584
rect 316 2576 324 2584
rect 1276 2576 1284 2584
rect 1356 2576 1364 2584
rect 1596 2576 1604 2584
rect 2108 2576 2116 2584
rect 2316 2576 2324 2584
rect 2492 2576 2500 2584
rect 2556 2576 2564 2584
rect 2940 2576 2948 2584
rect 3324 2576 3332 2584
rect 3580 2576 3588 2584
rect 3596 2576 3604 2584
rect 3772 2576 3780 2584
rect 3836 2576 3844 2584
rect 4108 2576 4116 2584
rect 4300 2576 4308 2584
rect 4492 2576 4500 2584
rect 4860 2576 4868 2584
rect 4876 2576 4884 2584
rect 5052 2576 5060 2584
rect 5116 2576 5124 2584
rect 5180 2576 5188 2584
rect 5308 2576 5316 2584
rect 5436 2576 5444 2584
rect 5564 2576 5572 2584
rect 60 2556 68 2564
rect 124 2556 132 2564
rect 188 2556 196 2564
rect 380 2556 388 2564
rect 444 2556 452 2564
rect 460 2556 468 2564
rect 572 2556 580 2564
rect 636 2556 644 2564
rect 652 2556 660 2564
rect 764 2556 772 2564
rect 44 2536 52 2544
rect 108 2536 116 2544
rect 172 2536 180 2544
rect 252 2536 260 2544
rect 268 2536 276 2544
rect 380 2536 388 2544
rect 460 2536 468 2544
rect 476 2536 484 2544
rect 510 2536 518 2544
rect 556 2536 564 2544
rect 668 2536 676 2544
rect 702 2536 710 2544
rect 748 2536 756 2544
rect 764 2536 772 2544
rect 812 2536 820 2544
rect 892 2556 900 2564
rect 972 2556 980 2564
rect 1084 2556 1092 2564
rect 1100 2556 1108 2564
rect 1164 2556 1172 2564
rect 1228 2556 1236 2564
rect 1292 2556 1300 2564
rect 1468 2556 1476 2564
rect 1532 2556 1540 2564
rect 1548 2556 1556 2564
rect 1612 2556 1620 2564
rect 1724 2556 1732 2564
rect 1788 2556 1796 2564
rect 1916 2556 1924 2564
rect 876 2536 884 2544
rect 956 2536 964 2544
rect 988 2536 996 2544
rect 1022 2536 1030 2544
rect 1068 2536 1076 2544
rect 1116 2536 1124 2544
rect 1180 2536 1188 2544
rect 1228 2536 1236 2544
rect 1244 2536 1252 2544
rect 1308 2536 1316 2544
rect 1342 2536 1350 2544
rect 1404 2536 1412 2544
rect 1452 2536 1460 2544
rect 1516 2536 1524 2544
rect 1564 2536 1572 2544
rect 1628 2536 1636 2544
rect 1788 2536 1796 2544
rect 1852 2536 1860 2544
rect 1900 2536 1908 2544
rect 1964 2536 1972 2544
rect 2044 2556 2052 2564
rect 2028 2536 2036 2544
rect 2060 2536 2068 2544
rect 2156 2536 2164 2544
rect 2236 2556 2244 2564
rect 2252 2556 2260 2564
rect 2428 2556 2436 2564
rect 2620 2556 2628 2564
rect 2684 2556 2692 2564
rect 2700 2556 2708 2564
rect 3004 2556 3012 2564
rect 3084 2556 3092 2564
rect 3516 2556 3524 2564
rect 3708 2556 3716 2564
rect 3916 2556 3924 2564
rect 4044 2556 4052 2564
rect 4220 2556 4228 2564
rect 4236 2556 4244 2564
rect 4476 2556 4484 2564
rect 4620 2556 4628 2564
rect 4940 2556 4948 2564
rect 5324 2556 5332 2564
rect 2252 2536 2260 2544
rect 2268 2536 2276 2544
rect 2302 2536 2310 2544
rect 2364 2536 2372 2544
rect 2412 2536 2420 2544
rect 2444 2536 2452 2544
rect 2508 2536 2516 2544
rect 2668 2536 2676 2544
rect 2716 2536 2724 2544
rect 2892 2536 2900 2544
rect 2988 2536 2996 2544
rect 3020 2536 3028 2544
rect 3100 2536 3108 2544
rect 3196 2536 3204 2544
rect 3212 2536 3220 2544
rect 3276 2536 3284 2544
rect 3340 2536 3348 2544
rect 3500 2536 3508 2544
rect 3532 2536 3540 2544
rect 3644 2536 3652 2544
rect 3692 2536 3700 2544
rect 3724 2536 3732 2544
rect 3788 2536 3796 2544
rect 3900 2536 3908 2544
rect 3932 2536 3940 2544
rect 4028 2536 4036 2544
rect 4060 2536 4068 2544
rect 4204 2536 4212 2544
rect 4348 2536 4356 2544
rect 4364 2536 4372 2544
rect 4460 2536 4468 2544
rect 4540 2536 4548 2544
rect 4604 2536 4612 2544
rect 4636 2536 4644 2544
rect 4748 2536 4756 2544
rect 4924 2536 4932 2544
rect 4940 2536 4948 2544
rect 4990 2536 4998 2544
rect 5068 2536 5076 2544
rect 5132 2536 5140 2544
rect 5196 2536 5204 2544
rect 5260 2536 5268 2544
rect 5340 2536 5348 2544
rect 5388 2536 5396 2544
rect 5452 2536 5460 2544
rect 5516 2536 5524 2544
rect 332 2516 340 2524
rect 908 2516 916 2524
rect 1036 2516 1044 2524
rect 1804 2516 1812 2524
rect 2572 2516 2580 2524
rect 3260 2516 3268 2524
rect 3852 2516 3860 2524
rect 4172 2516 4180 2524
rect 4684 2516 4692 2524
rect 4732 2516 4740 2524
rect 5004 2516 5012 2524
rect 5500 2516 5508 2524
rect 236 2496 244 2504
rect 284 2496 292 2504
rect 588 2496 596 2504
rect 940 2496 948 2504
rect 1388 2496 1396 2504
rect 1484 2496 1492 2504
rect 1676 2496 1684 2504
rect 1836 2496 1844 2504
rect 2076 2496 2084 2504
rect 2460 2496 2468 2504
rect 2524 2496 2532 2504
rect 2780 2496 2788 2504
rect 2844 2496 2852 2504
rect 2892 2496 2900 2504
rect 2956 2496 2964 2504
rect 3036 2496 3044 2504
rect 3132 2496 3140 2504
rect 3180 2496 3188 2504
rect 3228 2496 3236 2504
rect 3292 2496 3300 2504
rect 3340 2496 3348 2504
rect 3436 2496 3444 2504
rect 3548 2496 3556 2504
rect 3628 2496 3636 2504
rect 3660 2496 3668 2504
rect 3724 2496 3732 2504
rect 3804 2496 3812 2504
rect 3884 2496 3892 2504
rect 3980 2496 3988 2504
rect 4012 2496 4020 2504
rect 4092 2496 4100 2504
rect 4140 2496 4148 2504
rect 4284 2496 4292 2504
rect 4332 2496 4340 2504
rect 4380 2496 4388 2504
rect 4524 2496 4532 2504
rect 4556 2496 4564 2504
rect 4588 2496 4596 2504
rect 4668 2496 4676 2504
rect 4716 2496 4724 2504
rect 4764 2496 4772 2504
rect 4828 2496 4836 2504
rect 4924 2496 4932 2504
rect 5020 2496 5028 2504
rect 5084 2496 5092 2504
rect 5148 2496 5156 2504
rect 5212 2496 5220 2504
rect 5276 2496 5284 2504
rect 5372 2496 5380 2504
rect 5388 2496 5396 2504
rect 5468 2496 5476 2504
rect 5532 2496 5540 2504
rect 1148 2476 1156 2484
rect 3388 2476 3396 2484
rect 3404 2476 3412 2484
rect 4412 2476 4420 2484
rect 5260 2476 5268 2484
rect 3068 2456 3076 2464
rect 12 2436 20 2444
rect 76 2436 84 2444
rect 396 2436 404 2444
rect 524 2436 532 2444
rect 716 2436 724 2444
rect 1420 2436 1428 2444
rect 1660 2436 1668 2444
rect 1740 2436 1748 2444
rect 1868 2436 1876 2444
rect 1932 2436 1940 2444
rect 2124 2436 2132 2444
rect 3148 2436 3156 2444
rect 3964 2436 3972 2444
rect 4428 2436 4436 2444
rect 316 2376 324 2384
rect 380 2376 388 2384
rect 716 2376 724 2384
rect 892 2376 900 2384
rect 1596 2376 1604 2384
rect 2316 2376 2324 2384
rect 3212 2376 3220 2384
rect 3644 2376 3652 2384
rect 4044 2376 4052 2384
rect 4236 2376 4244 2384
rect 4860 2376 4868 2384
rect 5180 2376 5188 2384
rect 5244 2376 5252 2384
rect 5500 2376 5508 2384
rect 908 2356 916 2364
rect 1916 2356 1924 2364
rect 2124 2356 2132 2364
rect 3900 2356 3908 2364
rect 4348 2356 4356 2364
rect 5260 2356 5268 2364
rect 1980 2336 1988 2344
rect 2892 2336 2900 2344
rect 4876 2336 4884 2344
rect 124 2316 132 2324
rect 156 2316 164 2324
rect 220 2316 228 2324
rect 588 2316 596 2324
rect 684 2316 692 2324
rect 748 2316 756 2324
rect 796 2316 804 2324
rect 940 2316 948 2324
rect 1132 2316 1140 2324
rect 1324 2316 1332 2324
rect 1500 2316 1508 2324
rect 1772 2316 1780 2324
rect 1884 2316 1892 2324
rect 2028 2316 2036 2324
rect 2188 2316 2196 2324
rect 2476 2316 2484 2324
rect 2716 2316 2724 2324
rect 2780 2316 2788 2324
rect 2844 2316 2852 2324
rect 2972 2316 2980 2324
rect 3020 2316 3028 2324
rect 3180 2316 3188 2324
rect 3292 2316 3300 2324
rect 3420 2316 3428 2324
rect 3500 2316 3508 2324
rect 3596 2316 3604 2324
rect 3740 2316 3748 2324
rect 3804 2316 3812 2324
rect 3868 2316 3876 2324
rect 3932 2316 3940 2324
rect 4076 2316 4084 2324
rect 4188 2316 4196 2324
rect 4380 2316 4388 2324
rect 4412 2316 4420 2324
rect 4508 2316 4516 2324
rect 4604 2316 4612 2324
rect 4636 2316 4644 2324
rect 4716 2316 4724 2324
rect 4732 2316 4740 2324
rect 4780 2316 4788 2324
rect 4956 2316 4964 2324
rect 5020 2316 5028 2324
rect 5116 2316 5124 2324
rect 5148 2316 5156 2324
rect 5212 2316 5220 2324
rect 5324 2316 5332 2324
rect 5404 2316 5412 2324
rect 5468 2316 5476 2324
rect 5516 2316 5524 2324
rect 252 2296 260 2304
rect 572 2296 580 2304
rect 828 2296 836 2304
rect 1036 2296 1044 2304
rect 1676 2296 1684 2304
rect 2444 2296 2452 2304
rect 2956 2296 2964 2304
rect 3084 2296 3092 2304
rect 3340 2296 3348 2304
rect 3372 2296 3380 2304
rect 3452 2296 3460 2304
rect 3516 2296 3524 2304
rect 3676 2296 3684 2304
rect 3724 2296 3732 2304
rect 3916 2296 3924 2304
rect 3980 2296 3988 2304
rect 4092 2296 4100 2304
rect 4268 2296 4276 2304
rect 4284 2296 4292 2304
rect 4428 2296 4436 2304
rect 4940 2296 4948 2304
rect 28 2276 36 2284
rect 140 2276 148 2284
rect 204 2276 212 2284
rect 268 2276 276 2284
rect 348 2276 356 2284
rect 412 2276 420 2284
rect 492 2276 500 2284
rect 540 2276 548 2284
rect 620 2276 628 2284
rect 700 2276 708 2284
rect 764 2276 772 2284
rect 780 2276 788 2284
rect 844 2276 852 2284
rect 956 2276 964 2284
rect 972 2276 980 2284
rect 1068 2276 1076 2284
rect 1148 2276 1156 2284
rect 1196 2276 1204 2284
rect 12 2256 20 2264
rect 268 2256 276 2264
rect 332 2256 340 2264
rect 396 2256 404 2264
rect 508 2256 516 2264
rect 524 2256 532 2264
rect 636 2256 644 2264
rect 844 2256 852 2264
rect 972 2256 980 2264
rect 1084 2256 1092 2264
rect 1260 2276 1268 2284
rect 1340 2276 1348 2284
rect 1356 2276 1364 2284
rect 1436 2276 1444 2284
rect 1484 2276 1492 2284
rect 1564 2276 1572 2284
rect 1610 2276 1618 2284
rect 1660 2276 1668 2284
rect 1708 2276 1716 2284
rect 1788 2276 1796 2284
rect 1820 2276 1828 2284
rect 1868 2276 1876 2284
rect 1948 2276 1956 2284
rect 2044 2276 2052 2284
rect 2076 2276 2084 2284
rect 2156 2276 2164 2284
rect 2188 2276 2196 2284
rect 2268 2276 2276 2284
rect 2348 2276 2356 2284
rect 1276 2256 1284 2264
rect 1356 2256 1364 2264
rect 1420 2256 1428 2264
rect 1548 2256 1556 2264
rect 1660 2256 1668 2264
rect 1724 2256 1732 2264
rect 1804 2256 1812 2264
rect 1932 2256 1940 2264
rect 2060 2256 2068 2264
rect 2172 2256 2180 2264
rect 2252 2256 2260 2264
rect 2428 2276 2436 2284
rect 2492 2276 2500 2284
rect 2540 2276 2548 2284
rect 2588 2276 2596 2284
rect 2636 2276 2644 2284
rect 2700 2276 2708 2284
rect 2764 2276 2772 2284
rect 2828 2276 2836 2284
rect 2924 2276 2932 2284
rect 3052 2276 3060 2284
rect 3116 2276 3124 2284
rect 3196 2276 3204 2284
rect 3244 2276 3252 2284
rect 3276 2276 3284 2284
rect 3388 2276 3396 2284
rect 3404 2276 3412 2284
rect 3530 2276 3538 2284
rect 3564 2276 3572 2284
rect 3596 2276 3604 2284
rect 3660 2276 3668 2284
rect 3788 2276 3796 2284
rect 3852 2276 3860 2284
rect 4012 2276 4020 2284
rect 4140 2276 4148 2284
rect 4172 2276 4180 2284
rect 4316 2276 4324 2284
rect 4364 2276 4372 2284
rect 4460 2276 4468 2284
rect 4476 2276 4484 2284
rect 4556 2276 4564 2284
rect 4732 2276 4740 2284
rect 4796 2276 4804 2284
rect 4828 2276 4836 2284
rect 4908 2276 4916 2284
rect 5004 2276 5012 2284
rect 5084 2276 5092 2284
rect 5132 2276 5140 2284
rect 5196 2276 5204 2284
rect 5292 2276 5300 2284
rect 5356 2276 5364 2284
rect 5388 2276 5396 2284
rect 5452 2276 5460 2284
rect 5548 2276 5556 2284
rect 2428 2256 2436 2264
rect 2556 2256 2564 2264
rect 2572 2256 2580 2264
rect 2940 2256 2948 2264
rect 3068 2256 3076 2264
rect 3132 2256 3140 2264
rect 3260 2256 3268 2264
rect 3580 2256 3588 2264
rect 4028 2256 4036 2264
rect 4156 2256 4164 2264
rect 4300 2256 4308 2264
rect 4476 2256 4484 2264
rect 4556 2256 4564 2264
rect 4812 2256 4820 2264
rect 4924 2256 4932 2264
rect 5068 2256 5076 2264
rect 5308 2256 5316 2264
rect 5372 2256 5380 2264
rect 5564 2256 5572 2264
rect 60 2236 68 2244
rect 76 2236 84 2244
rect 188 2236 196 2244
rect 444 2236 452 2244
rect 460 2236 468 2244
rect 652 2236 660 2244
rect 908 2236 916 2244
rect 1020 2236 1028 2244
rect 1100 2236 1108 2244
rect 1164 2236 1172 2244
rect 1292 2236 1300 2244
rect 1404 2236 1412 2244
rect 1468 2236 1476 2244
rect 1532 2236 1540 2244
rect 1740 2236 1748 2244
rect 1852 2236 1860 2244
rect 1996 2236 2004 2244
rect 2108 2236 2116 2244
rect 2236 2236 2244 2244
rect 2300 2236 2308 2244
rect 2508 2236 2516 2244
rect 2684 2236 2692 2244
rect 2748 2236 2756 2244
rect 2812 2236 2820 2244
rect 2876 2236 2884 2244
rect 3004 2236 3012 2244
rect 3148 2236 3156 2244
rect 3324 2236 3332 2244
rect 3468 2236 3476 2244
rect 3708 2236 3716 2244
rect 3772 2236 3780 2244
rect 3836 2236 3844 2244
rect 3964 2236 3972 2244
rect 4044 2236 4052 2244
rect 4220 2236 4228 2244
rect 4540 2236 4548 2244
rect 4668 2236 4676 2244
rect 4684 2236 4692 2244
rect 4988 2236 4996 2244
rect 5052 2236 5060 2244
rect 5180 2236 5188 2244
rect 5436 2236 5444 2244
rect 204 2176 212 2184
rect 268 2176 276 2184
rect 572 2176 580 2184
rect 636 2176 644 2184
rect 716 2176 724 2184
rect 892 2176 900 2184
rect 972 2176 980 2184
rect 1036 2176 1044 2184
rect 1100 2176 1108 2184
rect 1276 2176 1284 2184
rect 1292 2176 1300 2184
rect 1420 2176 1428 2184
rect 1740 2176 1748 2184
rect 1804 2176 1812 2184
rect 1868 2176 1876 2184
rect 1980 2176 1988 2184
rect 2108 2176 2116 2184
rect 2172 2176 2180 2184
rect 2252 2176 2260 2184
rect 2364 2176 2372 2184
rect 2380 2176 2388 2184
rect 2492 2176 2500 2184
rect 2876 2176 2884 2184
rect 2892 2176 2900 2184
rect 2956 2176 2964 2184
rect 3020 2176 3028 2184
rect 3260 2176 3268 2184
rect 3276 2176 3284 2184
rect 3452 2176 3460 2184
rect 3580 2176 3588 2184
rect 3772 2176 3780 2184
rect 3788 2176 3796 2184
rect 3900 2176 3908 2184
rect 3916 2176 3924 2184
rect 4028 2176 4036 2184
rect 4156 2176 4164 2184
rect 4220 2176 4228 2184
rect 4236 2176 4244 2184
rect 4364 2176 4372 2184
rect 4620 2176 4628 2184
rect 4940 2176 4948 2184
rect 5324 2176 5332 2184
rect 5500 2176 5508 2184
rect 5564 2176 5572 2184
rect 60 2156 68 2164
rect 44 2136 52 2144
rect 108 2136 116 2144
rect 188 2156 196 2164
rect 316 2156 324 2164
rect 172 2136 180 2144
rect 252 2136 260 2144
rect 300 2136 308 2144
rect 364 2136 372 2144
rect 444 2156 452 2164
rect 508 2156 516 2164
rect 588 2156 596 2164
rect 652 2156 660 2164
rect 428 2136 436 2144
rect 492 2136 500 2144
rect 524 2136 532 2144
rect 604 2136 612 2144
rect 652 2136 660 2144
rect 702 2136 710 2144
rect 764 2136 772 2144
rect 812 2136 820 2144
rect 844 2156 852 2164
rect 1020 2156 1028 2164
rect 1212 2156 1220 2164
rect 1404 2156 1412 2164
rect 1532 2156 1540 2164
rect 1596 2156 1604 2164
rect 1660 2156 1668 2164
rect 1724 2156 1732 2164
rect 1852 2156 1860 2164
rect 1996 2156 2004 2164
rect 2236 2156 2244 2164
rect 2300 2156 2308 2164
rect 2508 2156 2516 2164
rect 2572 2156 2580 2164
rect 2700 2156 2708 2164
rect 860 2136 868 2144
rect 908 2136 916 2144
rect 1004 2136 1012 2144
rect 1084 2136 1092 2144
rect 1148 2136 1156 2144
rect 1196 2136 1204 2144
rect 1228 2136 1236 2144
rect 1340 2136 1348 2144
rect 1388 2136 1396 2144
rect 1468 2136 1476 2144
rect 1516 2136 1524 2144
rect 1580 2136 1588 2144
rect 1596 2136 1604 2144
rect 1644 2136 1652 2144
rect 1708 2136 1716 2144
rect 1788 2136 1796 2144
rect 1836 2136 1844 2144
rect 1916 2136 1924 2144
rect 1932 2136 1940 2144
rect 2012 2136 2020 2144
rect 2060 2136 2068 2144
rect 2124 2136 2132 2144
rect 2220 2136 2228 2144
rect 2284 2136 2292 2144
rect 2316 2136 2324 2144
rect 2428 2136 2436 2144
rect 2444 2136 2452 2144
rect 2524 2136 2532 2144
rect 2588 2136 2596 2144
rect 2636 2136 2644 2144
rect 2700 2136 2708 2144
rect 3084 2156 3092 2164
rect 3516 2156 3524 2164
rect 3596 2156 3604 2164
rect 3660 2156 3668 2164
rect 3980 2156 3988 2164
rect 4092 2156 4100 2164
rect 4348 2156 4356 2164
rect 4476 2156 4484 2164
rect 2780 2136 2788 2144
rect 2828 2136 2836 2144
rect 3004 2136 3012 2144
rect 3052 2136 3060 2144
rect 3100 2136 3108 2144
rect 3148 2136 3156 2144
rect 3324 2136 3332 2144
rect 3340 2136 3348 2144
rect 3404 2136 3412 2144
rect 3500 2136 3508 2144
rect 3516 2136 3524 2144
rect 3612 2136 3620 2144
rect 3676 2136 3684 2144
rect 3836 2136 3844 2144
rect 3852 2136 3860 2144
rect 3964 2136 3972 2144
rect 3980 2136 3988 2144
rect 4092 2136 4100 2144
rect 4108 2136 4116 2144
rect 4332 2136 4340 2144
rect 4412 2136 4420 2144
rect 4460 2136 4468 2144
rect 4508 2136 4516 2144
rect 4876 2156 4884 2164
rect 5196 2156 5204 2164
rect 5308 2156 5316 2164
rect 4572 2136 4580 2144
rect 4668 2136 4676 2144
rect 4748 2136 4756 2144
rect 4892 2136 4900 2144
rect 4988 2136 4996 2144
rect 5004 2136 5012 2144
rect 5132 2136 5140 2144
rect 5212 2136 5220 2144
rect 5258 2136 5266 2144
rect 5292 2136 5300 2144
rect 5372 2136 5380 2144
rect 5388 2136 5396 2144
rect 5452 2136 5460 2144
rect 5516 2136 5524 2144
rect 332 2116 340 2124
rect 924 2116 932 2124
rect 956 2116 964 2124
rect 1484 2116 1492 2124
rect 2684 2116 2692 2124
rect 2812 2116 2820 2124
rect 2940 2116 2948 2124
rect 3212 2116 3220 2124
rect 4172 2116 4180 2124
rect 4284 2116 4292 2124
rect 4396 2116 4404 2124
rect 4428 2116 4436 2124
rect 4540 2116 4548 2124
rect 4604 2116 4612 2124
rect 4684 2116 4692 2124
rect 4860 2116 4868 2124
rect 5052 2116 5060 2124
rect 5068 2116 5076 2124
rect 5116 2116 5124 2124
rect 5180 2116 5188 2124
rect 12 2096 20 2104
rect 236 2096 244 2104
rect 460 2096 468 2104
rect 540 2096 548 2104
rect 748 2096 756 2104
rect 908 2096 916 2104
rect 1068 2096 1076 2104
rect 1132 2096 1140 2104
rect 1244 2096 1252 2104
rect 1324 2096 1332 2104
rect 1452 2096 1460 2104
rect 1772 2096 1780 2104
rect 1788 2096 1796 2104
rect 1932 2096 1940 2104
rect 1948 2096 1956 2104
rect 2076 2096 2084 2104
rect 2140 2096 2148 2104
rect 2332 2096 2340 2104
rect 2412 2096 2420 2104
rect 2460 2096 2468 2104
rect 2652 2096 2660 2104
rect 2844 2096 2852 2104
rect 2924 2096 2932 2104
rect 2988 2096 2996 2104
rect 3148 2096 3156 2104
rect 3228 2096 3236 2104
rect 3340 2096 3348 2104
rect 3356 2096 3364 2104
rect 3420 2096 3428 2104
rect 3548 2096 3556 2104
rect 3644 2096 3652 2104
rect 3740 2096 3748 2104
rect 3820 2096 3828 2104
rect 3868 2096 3876 2104
rect 3948 2096 3956 2104
rect 4044 2096 4052 2104
rect 4124 2096 4132 2104
rect 4188 2096 4196 2104
rect 4268 2096 4276 2104
rect 4652 2096 4660 2104
rect 4668 2096 4676 2104
rect 4828 2096 4836 2104
rect 4924 2096 4932 2104
rect 4972 2096 4980 2104
rect 5020 2096 5028 2104
rect 5084 2096 5092 2104
rect 5148 2096 5156 2104
rect 5244 2096 5252 2104
rect 5356 2096 5364 2104
rect 5404 2096 5412 2104
rect 5468 2096 5476 2104
rect 5516 2096 5524 2104
rect 3388 2076 3396 2084
rect 5452 2076 5460 2084
rect 2620 2056 2628 2064
rect 76 2036 84 2044
rect 716 2036 724 2044
rect 780 2036 788 2044
rect 1100 2036 1108 2044
rect 1164 2036 1172 2044
rect 1356 2036 1364 2044
rect 1548 2036 1556 2044
rect 1676 2036 1684 2044
rect 2044 2036 2052 2044
rect 2188 2036 2196 2044
rect 2556 2036 2564 2044
rect 2956 2036 2964 2044
rect 3196 2036 3204 2044
rect 3468 2036 3476 2044
rect 3708 2036 3716 2044
rect 4300 2036 4308 2044
rect 12 1976 20 1984
rect 316 1976 324 1984
rect 524 1976 532 1984
rect 828 1976 836 1984
rect 844 1976 852 1984
rect 1292 1976 1300 1984
rect 1612 1976 1620 1984
rect 1868 1976 1876 1984
rect 2764 1976 2772 1984
rect 2956 1976 2964 1984
rect 3020 1976 3028 1984
rect 3196 1976 3204 1984
rect 3212 1976 3220 1984
rect 3660 1976 3668 1984
rect 4988 1976 4996 1984
rect 5436 1976 5444 1984
rect 700 1956 708 1964
rect 1484 1956 1492 1964
rect 1724 1956 1732 1964
rect 2444 1956 2452 1964
rect 4044 1956 4052 1964
rect 4284 1956 4292 1964
rect 4668 1956 4676 1964
rect 5132 1956 5140 1964
rect 2684 1936 2692 1944
rect 2892 1936 2900 1944
rect 3388 1936 3396 1944
rect 4732 1936 4740 1944
rect 5052 1936 5060 1944
rect 220 1916 228 1924
rect 348 1916 356 1924
rect 444 1916 452 1924
rect 492 1916 500 1924
rect 620 1916 628 1924
rect 1004 1916 1012 1924
rect 1068 1916 1076 1924
rect 1356 1916 1364 1924
rect 1676 1916 1684 1924
rect 1852 1916 1860 1924
rect 2268 1916 2276 1924
rect 2412 1916 2420 1924
rect 2588 1916 2596 1924
rect 2652 1916 2660 1924
rect 2732 1916 2740 1924
rect 2876 1916 2884 1924
rect 3244 1916 3252 1924
rect 3292 1916 3300 1924
rect 3340 1916 3348 1924
rect 3356 1916 3364 1924
rect 3468 1916 3476 1924
rect 3516 1916 3524 1924
rect 3580 1916 3588 1924
rect 3740 1916 3748 1924
rect 3932 1916 3940 1924
rect 4012 1916 4020 1924
rect 4204 1916 4212 1924
rect 4252 1916 4260 1924
rect 4300 1916 4308 1924
rect 4380 1916 4388 1924
rect 4428 1916 4436 1924
rect 4460 1916 4468 1924
rect 4604 1916 4612 1924
rect 4764 1916 4772 1924
rect 4844 1916 4852 1924
rect 4860 1916 4868 1924
rect 4956 1916 4964 1924
rect 5084 1916 5092 1924
rect 5164 1916 5172 1924
rect 5276 1916 5284 1924
rect 5324 1916 5332 1924
rect 5340 1916 5348 1924
rect 5372 1916 5380 1924
rect 5468 1916 5476 1924
rect 5532 1916 5540 1924
rect 140 1896 148 1904
rect 2188 1896 2196 1904
rect 2620 1896 2628 1904
rect 3148 1896 3156 1904
rect 3612 1896 3620 1904
rect 3836 1896 3844 1904
rect 4076 1896 4084 1904
rect 4492 1896 4500 1904
rect 4748 1896 4756 1904
rect 4812 1896 4820 1904
rect 4908 1896 4916 1904
rect 5068 1896 5076 1904
rect 44 1876 52 1884
rect 108 1876 116 1884
rect 172 1876 180 1884
rect 204 1876 212 1884
rect 284 1876 292 1884
rect 332 1876 340 1884
rect 412 1876 420 1884
rect 508 1876 516 1884
rect 556 1876 564 1884
rect 652 1876 660 1884
rect 668 1876 676 1884
rect 748 1876 756 1884
rect 796 1876 804 1884
rect 876 1876 884 1884
rect 124 1856 132 1864
rect 188 1856 196 1864
rect 268 1856 276 1864
rect 396 1856 404 1864
rect 572 1856 580 1864
rect 652 1856 660 1864
rect 764 1856 772 1864
rect 780 1856 788 1864
rect 908 1876 916 1884
rect 924 1876 932 1884
rect 1020 1876 1028 1884
rect 1084 1876 1092 1884
rect 1116 1876 1124 1884
rect 1196 1876 1204 1884
rect 1212 1876 1220 1884
rect 1244 1876 1252 1884
rect 1324 1876 1332 1884
rect 1452 1876 1460 1884
rect 1516 1876 1524 1884
rect 908 1856 916 1864
rect 1100 1856 1108 1864
rect 1228 1856 1236 1864
rect 1340 1856 1348 1864
rect 1404 1856 1412 1864
rect 1468 1856 1476 1864
rect 1580 1876 1588 1884
rect 1644 1876 1652 1884
rect 1676 1876 1684 1884
rect 1756 1876 1764 1884
rect 1820 1876 1828 1884
rect 1900 1876 1908 1884
rect 1596 1856 1604 1864
rect 1660 1856 1668 1864
rect 1740 1856 1748 1864
rect 1804 1856 1812 1864
rect 1964 1876 1972 1884
rect 1980 1876 1988 1884
rect 2076 1876 2084 1884
rect 1980 1856 1988 1864
rect 1996 1856 2004 1864
rect 2060 1856 2068 1864
rect 2140 1876 2148 1884
rect 2220 1876 2228 1884
rect 2252 1876 2260 1884
rect 2348 1876 2356 1884
rect 2428 1876 2436 1884
rect 2540 1876 2548 1884
rect 2572 1876 2580 1884
rect 2636 1876 2644 1884
rect 2748 1876 2756 1884
rect 2828 1876 2836 1884
rect 2844 1876 2852 1884
rect 2924 1876 2932 1884
rect 2988 1876 2996 1884
rect 3052 1876 3060 1884
rect 3100 1876 3108 1884
rect 3260 1876 3268 1884
rect 3276 1876 3284 1884
rect 3340 1876 3348 1884
rect 3420 1876 3428 1884
rect 3532 1876 3540 1884
rect 3596 1876 3604 1884
rect 3692 1876 3700 1884
rect 3724 1876 3732 1884
rect 3804 1876 3812 1884
rect 3852 1876 3860 1884
rect 4028 1876 4036 1884
rect 4108 1876 4116 1884
rect 4124 1876 4132 1884
rect 4158 1876 4166 1884
rect 4220 1876 4228 1884
rect 4236 1876 4244 1884
rect 4332 1876 4340 1884
rect 4364 1876 4372 1884
rect 4476 1876 4484 1884
rect 4524 1876 4532 1884
rect 4572 1876 4580 1884
rect 4636 1876 4644 1884
rect 4700 1876 4708 1884
rect 4860 1876 4868 1884
rect 4924 1876 4932 1884
rect 4940 1876 4948 1884
rect 5020 1876 5028 1884
rect 5196 1876 5204 1884
rect 5212 1876 5220 1884
rect 5324 1876 5332 1884
rect 5404 1876 5412 1884
rect 5452 1876 5460 1884
rect 5516 1876 5524 1884
rect 2236 1856 2244 1864
rect 2364 1856 2372 1864
rect 2492 1856 2500 1864
rect 2556 1856 2564 1864
rect 2812 1856 2820 1864
rect 2828 1856 2836 1864
rect 2940 1856 2948 1864
rect 3004 1856 3012 1864
rect 3068 1856 3076 1864
rect 3084 1856 3092 1864
rect 3404 1856 3412 1864
rect 3532 1856 3540 1864
rect 3708 1856 3716 1864
rect 3788 1856 3796 1864
rect 3852 1856 3860 1864
rect 4108 1856 4116 1864
rect 4348 1856 4356 1864
rect 4540 1856 4548 1864
rect 4620 1856 4628 1864
rect 4684 1856 4692 1864
rect 5004 1856 5012 1864
rect 5196 1856 5204 1864
rect 5388 1856 5396 1864
rect 252 1836 260 1844
rect 380 1836 388 1844
rect 460 1836 468 1844
rect 588 1836 596 1844
rect 700 1836 708 1844
rect 716 1836 724 1844
rect 956 1836 964 1844
rect 972 1836 980 1844
rect 1036 1836 1044 1844
rect 1148 1836 1156 1844
rect 1164 1836 1172 1844
rect 1276 1836 1284 1844
rect 1788 1836 1796 1844
rect 2044 1836 2052 1844
rect 2172 1836 2180 1844
rect 2300 1836 2308 1844
rect 2316 1836 2324 1844
rect 2380 1836 2388 1844
rect 2700 1836 2708 1844
rect 3644 1836 3652 1844
rect 3772 1836 3780 1844
rect 3964 1836 3972 1844
rect 3980 1836 3988 1844
rect 4172 1836 4180 1844
rect 4412 1836 4420 1844
rect 4796 1836 4804 1844
rect 5116 1836 5124 1844
rect 5500 1836 5508 1844
rect 5564 1836 5572 1844
rect 140 1776 148 1784
rect 396 1776 404 1784
rect 828 1776 836 1784
rect 844 1776 852 1784
rect 908 1776 916 1784
rect 1036 1776 1044 1784
rect 1276 1776 1284 1784
rect 1340 1776 1348 1784
rect 1356 1776 1364 1784
rect 1532 1776 1540 1784
rect 1548 1776 1556 1784
rect 1612 1776 1620 1784
rect 1676 1776 1684 1784
rect 1740 1776 1748 1784
rect 1916 1776 1924 1784
rect 2188 1776 2196 1784
rect 2252 1776 2260 1784
rect 2492 1776 2500 1784
rect 2572 1776 2580 1784
rect 2684 1776 2692 1784
rect 2748 1776 2756 1784
rect 2876 1776 2884 1784
rect 2956 1776 2964 1784
rect 3212 1776 3220 1784
rect 3324 1776 3332 1784
rect 3404 1776 3412 1784
rect 3516 1776 3524 1784
rect 3596 1776 3604 1784
rect 3772 1776 3780 1784
rect 3964 1776 3972 1784
rect 4028 1776 4036 1784
rect 4092 1776 4100 1784
rect 4108 1776 4116 1784
rect 4364 1776 4372 1784
rect 4860 1776 4868 1784
rect 4988 1776 4996 1784
rect 5244 1776 5252 1784
rect 5260 1776 5268 1784
rect 5372 1776 5380 1784
rect 5436 1776 5444 1784
rect 5564 1776 5572 1784
rect 60 1756 68 1764
rect 252 1756 260 1764
rect 316 1756 324 1764
rect 332 1756 340 1764
rect 444 1756 452 1764
rect 636 1756 644 1764
rect 700 1756 708 1764
rect 716 1756 724 1764
rect 956 1756 964 1764
rect 1020 1756 1028 1764
rect 1164 1756 1172 1764
rect 1292 1756 1300 1764
rect 1468 1756 1476 1764
rect 1484 1756 1492 1764
rect 1724 1756 1732 1764
rect 1788 1756 1796 1764
rect 1932 1756 1940 1764
rect 2060 1756 2068 1764
rect 2172 1756 2180 1764
rect 2316 1756 2324 1764
rect 2556 1756 2564 1764
rect 2892 1756 2900 1764
rect 3068 1756 3076 1764
rect 3196 1756 3204 1764
rect 3388 1756 3396 1764
rect 3580 1756 3588 1764
rect 3660 1756 3668 1764
rect 3788 1756 3796 1764
rect 4300 1756 4308 1764
rect 4476 1756 4484 1764
rect 4604 1756 4612 1764
rect 4620 1756 4628 1764
rect 4732 1756 4740 1764
rect 4876 1756 4884 1764
rect 5004 1756 5012 1764
rect 5132 1756 5140 1764
rect 5500 1756 5508 1764
rect 60 1736 68 1744
rect 124 1736 132 1744
rect 188 1736 196 1744
rect 300 1736 308 1744
rect 348 1736 356 1744
rect 444 1736 452 1744
rect 508 1736 516 1744
rect 524 1736 532 1744
rect 620 1736 628 1744
rect 684 1736 692 1744
rect 732 1736 740 1744
rect 780 1736 788 1744
rect 892 1736 900 1744
rect 940 1736 948 1744
rect 1004 1736 1012 1744
rect 1084 1736 1092 1744
rect 1100 1736 1108 1744
rect 1180 1736 1188 1744
rect 1228 1736 1236 1744
rect 1308 1736 1316 1744
rect 1404 1736 1412 1744
rect 1452 1736 1460 1744
rect 1468 1736 1476 1744
rect 1596 1736 1604 1744
rect 1660 1736 1668 1744
rect 1724 1736 1732 1744
rect 1788 1736 1796 1744
rect 1852 1736 1860 1744
rect 1868 1736 1876 1744
rect 1948 1736 1956 1744
rect 1996 1736 2004 1744
rect 2076 1736 2084 1744
rect 2156 1736 2164 1744
rect 2236 1736 2244 1744
rect 2316 1736 2324 1744
rect 2380 1736 2388 1744
rect 2444 1736 2452 1744
rect 2540 1736 2548 1744
rect 2620 1736 2628 1744
rect 2636 1736 2644 1744
rect 2700 1736 2708 1744
rect 2764 1736 2772 1744
rect 2828 1736 2836 1744
rect 2908 1736 2916 1744
rect 3018 1736 3026 1744
rect 3052 1736 3060 1744
rect 3084 1736 3092 1744
rect 3180 1736 3188 1744
rect 3260 1736 3268 1744
rect 3276 1736 3284 1744
rect 3372 1736 3380 1744
rect 3468 1736 3476 1744
rect 3564 1736 3572 1744
rect 3644 1736 3652 1744
rect 3676 1736 3684 1744
rect 3804 1736 3812 1744
rect 3852 1736 3860 1744
rect 3980 1736 3988 1744
rect 4156 1736 4164 1744
rect 4300 1736 4308 1744
rect 4316 1736 4324 1744
rect 4460 1736 4468 1744
rect 4588 1736 4596 1744
rect 4636 1736 4644 1744
rect 4732 1736 4740 1744
rect 4812 1736 4820 1744
rect 4892 1736 4900 1744
rect 5004 1736 5012 1744
rect 5068 1736 5076 1744
rect 5148 1736 5156 1744
rect 5308 1736 5316 1744
rect 5324 1736 5332 1744
rect 5388 1736 5396 1744
rect 5484 1736 5492 1744
rect 5516 1736 5524 1744
rect 204 1716 212 1724
rect 460 1716 468 1724
rect 572 1716 580 1724
rect 1420 1716 1428 1724
rect 1804 1716 1812 1724
rect 2044 1716 2052 1724
rect 2124 1716 2132 1724
rect 2300 1716 2308 1724
rect 2428 1716 2436 1724
rect 2812 1716 2820 1724
rect 3004 1716 3012 1724
rect 3132 1716 3140 1724
rect 3452 1716 3460 1724
rect 4044 1716 4052 1724
rect 4412 1716 4420 1724
rect 4748 1716 4756 1724
rect 5196 1716 5204 1724
rect 108 1696 116 1704
rect 188 1696 196 1704
rect 380 1696 388 1704
rect 492 1696 500 1704
rect 540 1696 548 1704
rect 876 1696 884 1704
rect 1068 1696 1076 1704
rect 1116 1696 1124 1704
rect 1388 1696 1396 1704
rect 1580 1696 1588 1704
rect 1644 1696 1652 1704
rect 1836 1696 1844 1704
rect 1884 1696 1892 1704
rect 2012 1696 2020 1704
rect 2236 1696 2244 1704
rect 2300 1696 2308 1704
rect 2396 1696 2404 1704
rect 2444 1696 2452 1704
rect 2604 1696 2612 1704
rect 2652 1696 2660 1704
rect 2716 1696 2724 1704
rect 2780 1696 2788 1704
rect 2828 1696 2836 1704
rect 2940 1696 2948 1704
rect 2988 1696 2996 1704
rect 3084 1696 3092 1704
rect 3244 1696 3252 1704
rect 3292 1696 3300 1704
rect 3436 1696 3444 1704
rect 3484 1696 3492 1704
rect 3532 1696 3540 1704
rect 3644 1696 3652 1704
rect 3740 1696 3748 1704
rect 3868 1696 3876 1704
rect 3932 1696 3940 1704
rect 3996 1696 4004 1704
rect 4060 1696 4068 1704
rect 4140 1696 4148 1704
rect 4204 1696 4212 1704
rect 4268 1696 4276 1704
rect 4524 1696 4532 1704
rect 4764 1696 4772 1704
rect 4828 1696 4836 1704
rect 4956 1696 4964 1704
rect 5052 1696 5060 1704
rect 5084 1696 5092 1704
rect 5292 1696 5300 1704
rect 5404 1696 5412 1704
rect 5532 1696 5540 1704
rect 3340 1676 3348 1684
rect 3836 1676 3844 1684
rect 4348 1676 4356 1684
rect 4556 1676 4564 1684
rect 4684 1676 4692 1684
rect 12 1636 20 1644
rect 76 1636 84 1644
rect 396 1636 404 1644
rect 588 1636 596 1644
rect 652 1636 660 1644
rect 972 1636 980 1644
rect 1148 1636 1156 1644
rect 1980 1636 1988 1644
rect 2108 1636 2116 1644
rect 2364 1636 2372 1644
rect 2508 1636 2516 1644
rect 3148 1636 3156 1644
rect 4492 1636 4500 1644
rect 4668 1636 4676 1644
rect 4796 1636 4804 1644
rect 5116 1636 5124 1644
rect 5452 1636 5460 1644
rect 140 1576 148 1584
rect 204 1576 212 1584
rect 1404 1576 1412 1584
rect 1548 1576 1556 1584
rect 1676 1576 1684 1584
rect 1916 1576 1924 1584
rect 1932 1576 1940 1584
rect 2700 1576 2708 1584
rect 2828 1576 2836 1584
rect 3004 1576 3012 1584
rect 3324 1576 3332 1584
rect 3708 1576 3716 1584
rect 3724 1576 3732 1584
rect 4284 1576 4292 1584
rect 4364 1576 4372 1584
rect 4860 1576 4868 1584
rect 1036 1556 1044 1564
rect 1660 1556 1668 1564
rect 2060 1556 2068 1564
rect 4732 1556 4740 1564
rect 4860 1556 4868 1564
rect 1164 1536 1172 1544
rect 1420 1536 1428 1544
rect 2236 1536 2244 1544
rect 3068 1536 3076 1544
rect 3468 1536 3476 1544
rect 3596 1536 3604 1544
rect 4028 1536 4036 1544
rect 4860 1536 4868 1544
rect 4940 1536 4948 1544
rect 5180 1536 5188 1544
rect 412 1516 420 1524
rect 828 1516 836 1524
rect 1004 1516 1012 1524
rect 1068 1516 1076 1524
rect 1196 1516 1204 1524
rect 1244 1516 1252 1524
rect 1452 1516 1460 1524
rect 1740 1516 1748 1524
rect 1804 1516 1812 1524
rect 2092 1516 2100 1524
rect 2172 1516 2180 1524
rect 2220 1516 2228 1524
rect 2332 1516 2340 1524
rect 2428 1516 2436 1524
rect 2524 1516 2532 1524
rect 2572 1516 2580 1524
rect 2668 1516 2676 1524
rect 2732 1516 2740 1524
rect 2892 1516 2900 1524
rect 3052 1516 3060 1524
rect 3148 1516 3156 1524
rect 3212 1516 3220 1524
rect 3276 1516 3284 1524
rect 3356 1516 3364 1524
rect 3564 1516 3572 1524
rect 3756 1516 3764 1524
rect 3804 1516 3812 1524
rect 3900 1516 3908 1524
rect 3964 1516 3972 1524
rect 3980 1516 3988 1524
rect 4044 1516 4052 1524
rect 4140 1516 4148 1524
rect 4172 1516 4180 1524
rect 4332 1516 4340 1524
rect 4524 1516 4532 1524
rect 4556 1516 4564 1524
rect 4636 1516 4644 1524
rect 4700 1516 4708 1524
rect 4748 1516 4756 1524
rect 4876 1516 4884 1524
rect 5020 1516 5028 1524
rect 5100 1516 5108 1524
rect 5132 1516 5140 1524
rect 5276 1516 5284 1524
rect 5324 1516 5332 1524
rect 5372 1516 5380 1524
rect 5420 1516 5428 1524
rect 5452 1516 5460 1524
rect 5516 1516 5524 1524
rect 5532 1516 5540 1524
rect 460 1496 468 1504
rect 700 1496 708 1504
rect 1276 1496 1284 1504
rect 1484 1496 1492 1504
rect 1884 1496 1892 1504
rect 2444 1496 2452 1504
rect 2556 1496 2564 1504
rect 3068 1496 3076 1504
rect 3340 1496 3348 1504
rect 3452 1496 3460 1504
rect 3852 1496 3860 1504
rect 4412 1496 4420 1504
rect 4684 1496 4692 1504
rect 5116 1496 5124 1504
rect 5244 1496 5252 1504
rect 5436 1496 5444 1504
rect 44 1476 52 1484
rect 108 1476 116 1484
rect 172 1476 180 1484
rect 364 1476 372 1484
rect 396 1476 404 1484
rect 492 1476 500 1484
rect 60 1456 68 1464
rect 124 1456 132 1464
rect 188 1456 196 1464
rect 252 1456 260 1464
rect 316 1456 324 1464
rect 380 1456 388 1464
rect 636 1476 644 1484
rect 652 1476 660 1484
rect 714 1476 722 1484
rect 764 1476 772 1484
rect 828 1476 836 1484
rect 876 1476 884 1484
rect 572 1456 580 1464
rect 636 1456 644 1464
rect 652 1456 660 1464
rect 764 1456 772 1464
rect 940 1476 948 1484
rect 1020 1476 1028 1484
rect 1084 1476 1092 1484
rect 1116 1476 1124 1484
rect 1150 1476 1158 1484
rect 1212 1476 1220 1484
rect 1228 1476 1236 1484
rect 1324 1476 1332 1484
rect 1372 1476 1380 1484
rect 1468 1476 1476 1484
rect 1516 1476 1524 1484
rect 1580 1476 1588 1484
rect 1628 1476 1636 1484
rect 1708 1476 1716 1484
rect 1772 1476 1780 1484
rect 1836 1476 1844 1484
rect 1868 1476 1876 1484
rect 1964 1476 1972 1484
rect 2028 1476 2036 1484
rect 2108 1476 2116 1484
rect 2140 1476 2148 1484
rect 2236 1476 2244 1484
rect 2284 1476 2292 1484
rect 2316 1476 2324 1484
rect 2396 1476 2404 1484
rect 2492 1476 2500 1484
rect 2508 1476 2516 1484
rect 2604 1476 2612 1484
rect 2684 1476 2692 1484
rect 2748 1476 2756 1484
rect 2780 1476 2788 1484
rect 2860 1476 2868 1484
rect 2956 1476 2964 1484
rect 2972 1476 2980 1484
rect 3116 1476 3124 1484
rect 3180 1476 3188 1484
rect 3260 1476 3268 1484
rect 3276 1476 3284 1484
rect 3420 1476 3428 1484
rect 3500 1476 3508 1484
rect 3628 1476 3636 1484
rect 3676 1476 3684 1484
rect 3772 1476 3780 1484
rect 3788 1476 3796 1484
rect 3916 1476 3924 1484
rect 3932 1476 3940 1484
rect 3980 1476 3988 1484
rect 4076 1476 4084 1484
rect 4092 1476 4100 1484
rect 4156 1476 4164 1484
rect 4172 1476 4180 1484
rect 4252 1476 4260 1484
rect 4348 1476 4356 1484
rect 4460 1476 4468 1484
rect 4540 1476 4548 1484
rect 4588 1476 4596 1484
rect 4620 1476 4628 1484
rect 4780 1476 4788 1484
rect 4828 1476 4836 1484
rect 4876 1476 4884 1484
rect 4972 1476 4980 1484
rect 4988 1476 4996 1484
rect 5132 1476 5140 1484
rect 5196 1476 5204 1484
rect 5324 1476 5332 1484
rect 5452 1476 5460 1484
rect 5516 1476 5524 1484
rect 956 1456 964 1464
rect 1100 1456 1108 1464
rect 1340 1456 1348 1464
rect 1356 1456 1364 1464
rect 1532 1456 1540 1464
rect 1596 1456 1604 1464
rect 1612 1456 1620 1464
rect 1724 1456 1732 1464
rect 1788 1456 1796 1464
rect 1852 1456 1860 1464
rect 1980 1456 1988 1464
rect 2044 1456 2052 1464
rect 2124 1456 2132 1464
rect 2300 1456 2308 1464
rect 2380 1456 2388 1464
rect 2492 1456 2500 1464
rect 2620 1456 2628 1464
rect 2764 1456 2772 1464
rect 2876 1456 2884 1464
rect 2940 1456 2948 1464
rect 2956 1456 2964 1464
rect 3132 1456 3140 1464
rect 3196 1456 3204 1464
rect 3260 1456 3268 1464
rect 3404 1456 3412 1464
rect 3516 1456 3524 1464
rect 3644 1456 3652 1464
rect 3660 1456 3668 1464
rect 3916 1456 3924 1464
rect 4092 1456 4100 1464
rect 4236 1456 4244 1464
rect 4476 1456 4484 1464
rect 4604 1456 4612 1464
rect 4796 1456 4804 1464
rect 4812 1456 4820 1464
rect 4988 1456 4996 1464
rect 5196 1456 5204 1464
rect 12 1436 20 1444
rect 76 1436 84 1444
rect 444 1436 452 1444
rect 780 1436 788 1444
rect 844 1436 852 1444
rect 972 1436 980 1444
rect 1292 1436 1300 1444
rect 1996 1436 2004 1444
rect 2188 1436 2196 1444
rect 2364 1436 2372 1444
rect 2636 1436 2644 1444
rect 2812 1436 2820 1444
rect 3020 1436 3028 1444
rect 3388 1436 3396 1444
rect 3532 1436 3540 1444
rect 3708 1436 3716 1444
rect 3836 1436 3844 1444
rect 4108 1436 4116 1444
rect 4220 1436 4228 1444
rect 4300 1436 4308 1444
rect 4492 1436 4500 1444
rect 4668 1436 4676 1444
rect 4860 1436 4868 1444
rect 4924 1436 4932 1444
rect 5052 1436 5060 1444
rect 5068 1436 5076 1444
rect 5308 1436 5316 1444
rect 5388 1436 5396 1444
rect 5564 1436 5572 1444
rect 140 1376 148 1384
rect 252 1376 260 1384
rect 316 1376 324 1384
rect 396 1376 404 1384
rect 572 1376 580 1384
rect 652 1376 660 1384
rect 716 1376 724 1384
rect 780 1376 788 1384
rect 844 1376 852 1384
rect 972 1376 980 1384
rect 1660 1376 1668 1384
rect 1804 1376 1812 1384
rect 1996 1376 2004 1384
rect 2300 1376 2308 1384
rect 2316 1376 2324 1384
rect 2684 1376 2692 1384
rect 2748 1376 2756 1384
rect 2812 1376 2820 1384
rect 3084 1376 3092 1384
rect 3276 1376 3284 1384
rect 3388 1376 3396 1384
rect 3468 1376 3476 1384
rect 3532 1376 3540 1384
rect 3644 1376 3652 1384
rect 3916 1376 3924 1384
rect 4028 1376 4036 1384
rect 4044 1376 4052 1384
rect 4108 1376 4116 1384
rect 4540 1376 4548 1384
rect 4620 1376 4628 1384
rect 4860 1376 4868 1384
rect 4924 1376 4932 1384
rect 5116 1376 5124 1384
rect 5132 1376 5140 1384
rect 5244 1376 5252 1384
rect 5308 1376 5316 1384
rect 5372 1376 5380 1384
rect 5436 1376 5444 1384
rect 5452 1376 5460 1384
rect 12 1356 20 1364
rect 124 1356 132 1364
rect 204 1356 212 1364
rect 380 1356 388 1364
rect 444 1356 452 1364
rect 508 1356 516 1364
rect 636 1356 644 1364
rect 700 1356 708 1364
rect 892 1356 900 1364
rect 1020 1356 1028 1364
rect 1084 1356 1092 1364
rect 1100 1356 1108 1364
rect 1212 1356 1220 1364
rect 1228 1356 1236 1364
rect 1356 1356 1364 1364
rect 1420 1356 1428 1364
rect 1484 1356 1492 1364
rect 1548 1356 1556 1364
rect 1724 1356 1732 1364
rect 1788 1356 1796 1364
rect 1980 1356 1988 1364
rect 2060 1356 2068 1364
rect 2124 1356 2132 1364
rect 2188 1356 2196 1364
rect 2364 1356 2372 1364
rect 2444 1356 2452 1364
rect 2508 1356 2516 1364
rect 2700 1356 2708 1364
rect 3068 1356 3076 1364
rect 3196 1356 3204 1364
rect 3260 1356 3268 1364
rect 3340 1356 3348 1364
rect 3404 1356 3412 1364
rect 3708 1356 3716 1364
rect 28 1336 36 1344
rect 108 1336 116 1344
rect 188 1336 196 1344
rect 220 1336 228 1344
rect 268 1336 276 1344
rect 330 1336 338 1344
rect 380 1336 388 1344
rect 428 1336 436 1344
rect 492 1336 500 1344
rect 524 1336 532 1344
rect 620 1336 628 1344
rect 684 1336 692 1344
rect 764 1336 772 1344
rect 828 1336 836 1344
rect 892 1336 900 1344
rect 956 1336 964 1344
rect 1004 1336 1012 1344
rect 1068 1336 1076 1344
rect 1116 1336 1124 1344
rect 1162 1336 1170 1344
rect 1196 1336 1204 1344
rect 1244 1336 1252 1344
rect 1292 1336 1300 1344
rect 1372 1336 1380 1344
rect 1436 1336 1444 1344
rect 1484 1336 1492 1344
rect 1500 1336 1508 1344
rect 1548 1336 1556 1344
rect 1612 1336 1620 1344
rect 1674 1336 1682 1344
rect 1708 1336 1716 1344
rect 1772 1336 1780 1344
rect 1852 1336 1860 1344
rect 1916 1336 1924 1344
rect 1964 1336 1972 1344
rect 2044 1336 2052 1344
rect 2076 1336 2084 1344
rect 2140 1336 2148 1344
rect 2188 1336 2196 1344
rect 2252 1336 2260 1344
rect 2348 1336 2356 1344
rect 2444 1336 2452 1344
rect 2460 1336 2468 1344
rect 2524 1336 2532 1344
rect 2636 1336 2644 1344
rect 2716 1336 2724 1344
rect 2764 1336 2772 1344
rect 2828 1336 2836 1344
rect 3052 1336 3060 1344
rect 3132 1336 3140 1344
rect 3180 1336 3188 1344
rect 3244 1336 3252 1344
rect 3324 1336 3332 1344
rect 3356 1336 3364 1344
rect 3420 1336 3428 1344
rect 3516 1336 3524 1344
rect 3580 1336 3588 1344
rect 3596 1336 3604 1344
rect 3692 1336 3700 1344
rect 3708 1336 3716 1344
rect 4732 1356 4740 1364
rect 4796 1356 4804 1364
rect 4940 1356 4948 1364
rect 5260 1356 5268 1364
rect 3740 1336 3748 1344
rect 3788 1336 3796 1344
rect 3852 1336 3860 1344
rect 3964 1336 3972 1344
rect 3980 1336 3988 1344
rect 4092 1336 4100 1344
rect 4156 1336 4164 1344
rect 4172 1336 4180 1344
rect 4236 1336 4244 1344
rect 4300 1336 4308 1344
rect 4364 1336 4372 1344
rect 4428 1336 4436 1344
rect 4492 1336 4500 1344
rect 4604 1336 4612 1344
rect 4716 1336 4724 1344
rect 4780 1336 4788 1344
rect 4812 1336 4820 1344
rect 4876 1336 4884 1344
rect 4956 1336 4964 1344
rect 5004 1336 5012 1344
rect 5068 1336 5076 1344
rect 5180 1336 5188 1344
rect 5196 1336 5204 1344
rect 5276 1336 5284 1344
rect 5324 1336 5332 1344
rect 5388 1336 5396 1344
rect 5500 1336 5508 1344
rect 908 1316 916 1324
rect 1468 1316 1476 1324
rect 2620 1316 2628 1324
rect 4284 1316 4292 1324
rect 4556 1316 4564 1324
rect 172 1296 180 1304
rect 284 1296 292 1304
rect 540 1296 548 1304
rect 748 1296 756 1304
rect 812 1296 820 1304
rect 940 1296 948 1304
rect 1308 1296 1316 1304
rect 1628 1296 1636 1304
rect 1836 1296 1844 1304
rect 1868 1296 1876 1304
rect 1900 1296 1908 1304
rect 2044 1296 2052 1304
rect 2108 1296 2116 1304
rect 2172 1296 2180 1304
rect 2268 1296 2276 1304
rect 2412 1296 2420 1304
rect 2588 1296 2596 1304
rect 2652 1296 2660 1304
rect 2780 1296 2788 1304
rect 2828 1296 2836 1304
rect 2908 1296 2916 1304
rect 2956 1296 2964 1304
rect 3004 1296 3012 1304
rect 3116 1296 3124 1304
rect 3148 1296 3156 1304
rect 3308 1296 3316 1304
rect 3500 1296 3508 1304
rect 3564 1296 3572 1304
rect 3612 1296 3620 1304
rect 3804 1296 3812 1304
rect 3868 1296 3876 1304
rect 3948 1296 3956 1304
rect 3964 1296 3972 1304
rect 4092 1296 4100 1304
rect 4140 1296 4148 1304
rect 4188 1296 4196 1304
rect 4236 1296 4244 1304
rect 4316 1296 4324 1304
rect 4380 1296 4388 1304
rect 4492 1296 4500 1304
rect 4508 1296 4516 1304
rect 4588 1296 4596 1304
rect 4668 1296 4676 1304
rect 4748 1296 4756 1304
rect 4828 1296 4836 1304
rect 4892 1296 4900 1304
rect 5052 1296 5060 1304
rect 5084 1296 5092 1304
rect 5180 1296 5188 1304
rect 5196 1296 5204 1304
rect 5340 1296 5348 1304
rect 5404 1296 5412 1304
rect 5484 1296 5492 1304
rect 460 1276 468 1284
rect 1340 1276 1348 1284
rect 1932 1276 1940 1284
rect 2236 1276 2244 1284
rect 2492 1276 2500 1284
rect 2940 1276 2948 1284
rect 3772 1276 3780 1284
rect 3852 1276 3860 1284
rect 3900 1276 3908 1284
rect 4236 1276 4244 1284
rect 4364 1276 4372 1284
rect 1036 1256 1044 1264
rect 1596 1256 1604 1264
rect 3212 1256 3220 1264
rect 60 1236 68 1244
rect 76 1236 84 1244
rect 588 1236 596 1244
rect 972 1236 980 1244
rect 1148 1236 1156 1244
rect 1276 1236 1284 1244
rect 1404 1236 1412 1244
rect 1532 1236 1540 1244
rect 1740 1236 1748 1244
rect 2380 1236 2388 1244
rect 3452 1236 3460 1244
rect 3660 1236 3668 1244
rect 76 1176 84 1184
rect 140 1176 148 1184
rect 780 1176 788 1184
rect 908 1176 916 1184
rect 1148 1176 1156 1184
rect 1340 1176 1348 1184
rect 1596 1176 1604 1184
rect 1676 1176 1684 1184
rect 2252 1176 2260 1184
rect 2380 1176 2388 1184
rect 2444 1176 2452 1184
rect 2508 1176 2516 1184
rect 2828 1176 2836 1184
rect 3132 1176 3140 1184
rect 3196 1176 3204 1184
rect 3468 1176 3476 1184
rect 3596 1176 3604 1184
rect 3660 1176 3668 1184
rect 3900 1176 3908 1184
rect 4108 1176 4116 1184
rect 5388 1176 5396 1184
rect 252 1156 260 1164
rect 1612 1156 1620 1164
rect 2364 1156 2372 1164
rect 4428 1156 4436 1164
rect 4876 1156 4884 1164
rect 524 1136 532 1144
rect 1404 1136 1412 1144
rect 2892 1136 2900 1144
rect 3980 1136 3988 1144
rect 4156 1136 4164 1144
rect 5052 1136 5060 1144
rect 5308 1136 5316 1144
rect 268 1116 276 1124
rect 476 1116 484 1124
rect 556 1116 564 1124
rect 748 1116 756 1124
rect 828 1116 836 1124
rect 860 1116 868 1124
rect 972 1116 980 1124
rect 1068 1116 1076 1124
rect 1116 1116 1124 1124
rect 1196 1116 1204 1124
rect 1260 1116 1268 1124
rect 1388 1116 1396 1124
rect 1756 1116 1764 1124
rect 1804 1116 1812 1124
rect 1948 1116 1956 1124
rect 2044 1116 2052 1124
rect 2092 1116 2100 1124
rect 2108 1116 2116 1124
rect 2220 1116 2228 1124
rect 2332 1116 2340 1124
rect 2412 1116 2420 1124
rect 2540 1116 2548 1124
rect 2604 1116 2612 1124
rect 2796 1116 2804 1124
rect 3020 1116 3028 1124
rect 3260 1116 3268 1124
rect 3308 1116 3316 1124
rect 3452 1116 3460 1124
rect 3580 1116 3588 1124
rect 3788 1116 3796 1124
rect 3964 1116 3972 1124
rect 4060 1116 4068 1124
rect 4092 1116 4100 1124
rect 4140 1116 4148 1124
rect 4332 1116 4340 1124
rect 4476 1116 4484 1124
rect 4588 1116 4596 1124
rect 4636 1116 4644 1124
rect 4700 1116 4708 1124
rect 4748 1116 4756 1124
rect 4812 1116 4820 1124
rect 4908 1116 4916 1124
rect 4972 1116 4980 1124
rect 5020 1116 5028 1124
rect 5084 1116 5092 1124
rect 5212 1116 5220 1124
rect 5340 1116 5348 1124
rect 5420 1116 5428 1124
rect 2860 1096 2868 1104
rect 2876 1096 2884 1104
rect 3276 1096 3284 1104
rect 4044 1096 4052 1104
rect 4156 1096 4164 1104
rect 4236 1096 4244 1104
rect 4348 1096 4356 1104
rect 4396 1096 4404 1104
rect 4620 1096 4628 1104
rect 4764 1096 4772 1104
rect 5004 1096 5012 1104
rect 5180 1096 5188 1104
rect 5436 1096 5444 1104
rect 28 1076 36 1084
rect 108 1076 116 1084
rect 172 1076 180 1084
rect 220 1076 228 1084
rect 300 1076 308 1084
rect 348 1076 356 1084
rect 444 1076 452 1084
rect 460 1076 468 1084
rect 620 1076 628 1084
rect 668 1076 676 1084
rect 764 1076 772 1084
rect 828 1076 836 1084
rect 844 1076 852 1084
rect 940 1076 948 1084
rect 972 1076 980 1084
rect 1084 1076 1092 1084
rect 1100 1076 1108 1084
rect 1212 1076 1220 1084
rect 1276 1076 1284 1084
rect 1308 1076 1316 1084
rect 1342 1076 1350 1084
rect 1404 1076 1412 1084
rect 1420 1076 1428 1084
rect 1500 1076 1508 1084
rect 12 1056 20 1064
rect 124 1056 132 1064
rect 188 1056 196 1064
rect 204 1056 212 1064
rect 316 1056 324 1064
rect 332 1056 340 1064
rect 636 1056 644 1064
rect 652 1056 660 1064
rect 956 1056 964 1064
rect 1292 1056 1300 1064
rect 1484 1056 1492 1064
rect 1564 1076 1572 1084
rect 1644 1076 1652 1084
rect 1708 1076 1716 1084
rect 1740 1076 1748 1084
rect 1836 1076 1844 1084
rect 1900 1076 1908 1084
rect 1932 1076 1940 1084
rect 2012 1076 2020 1084
rect 2108 1076 2116 1084
rect 2124 1076 2132 1084
rect 2236 1076 2244 1084
rect 2284 1076 2292 1084
rect 2316 1076 2324 1084
rect 2428 1076 2436 1084
rect 2476 1076 2484 1084
rect 2556 1076 2564 1084
rect 2620 1076 2628 1084
rect 2668 1076 2676 1084
rect 2732 1076 2740 1084
rect 2812 1076 2820 1084
rect 2924 1076 2932 1084
rect 2954 1076 2962 1084
rect 3004 1076 3012 1084
rect 3052 1076 3060 1084
rect 3100 1076 3108 1084
rect 3164 1076 3172 1084
rect 3228 1076 3236 1084
rect 3372 1076 3380 1084
rect 3452 1076 3460 1084
rect 3500 1076 3508 1084
rect 1660 1056 1668 1064
rect 1724 1056 1732 1064
rect 1852 1056 1860 1064
rect 1916 1056 1924 1064
rect 1996 1056 2004 1064
rect 2300 1056 2308 1064
rect 2492 1056 2500 1064
rect 2684 1056 2692 1064
rect 2748 1056 2756 1064
rect 2940 1056 2948 1064
rect 3004 1056 3012 1064
rect 3068 1056 3076 1064
rect 3084 1056 3092 1064
rect 3148 1056 3156 1064
rect 3212 1056 3220 1064
rect 3388 1056 3396 1064
rect 3516 1056 3524 1064
rect 3548 1076 3556 1084
rect 3628 1076 3636 1084
rect 3692 1076 3700 1084
rect 3740 1076 3748 1084
rect 3868 1076 3876 1084
rect 3932 1076 3940 1084
rect 4012 1076 4020 1084
rect 4204 1076 4212 1084
rect 4268 1076 4276 1084
rect 4412 1076 4420 1084
rect 4492 1076 4500 1084
rect 4508 1076 4516 1084
rect 4542 1076 4550 1084
rect 4604 1076 4612 1084
rect 4684 1076 4692 1084
rect 4748 1076 4756 1084
rect 4844 1076 4852 1084
rect 4924 1076 4932 1084
rect 4988 1076 4996 1084
rect 5068 1076 5076 1084
rect 5148 1076 5156 1084
rect 5196 1076 5204 1084
rect 5276 1076 5284 1084
rect 5324 1076 5332 1084
rect 5468 1076 5476 1084
rect 3644 1056 3652 1064
rect 3708 1056 3716 1064
rect 3724 1056 3732 1064
rect 3852 1056 3860 1064
rect 3916 1056 3924 1064
rect 4028 1056 4036 1064
rect 4220 1056 4228 1064
rect 4284 1056 4292 1064
rect 4492 1056 4500 1064
rect 4860 1056 4868 1064
rect 5132 1056 5140 1064
rect 5260 1056 5268 1064
rect 5452 1056 5460 1064
rect 60 1036 68 1044
rect 380 1036 388 1044
rect 396 1036 404 1044
rect 508 1036 516 1044
rect 700 1036 708 1044
rect 716 1036 724 1044
rect 892 1036 900 1044
rect 1020 1036 1028 1044
rect 1036 1036 1044 1044
rect 1148 1036 1156 1044
rect 1164 1036 1172 1044
rect 1228 1036 1236 1044
rect 1356 1036 1364 1044
rect 1468 1036 1476 1044
rect 1788 1036 1796 1044
rect 1868 1036 1876 1044
rect 1980 1036 1988 1044
rect 2060 1036 2068 1044
rect 2172 1036 2180 1044
rect 2188 1036 2196 1044
rect 2572 1036 2580 1044
rect 2636 1036 2644 1044
rect 2700 1036 2708 1044
rect 2764 1036 2772 1044
rect 3404 1036 3412 1044
rect 3660 1036 3668 1044
rect 3836 1036 3844 1044
rect 4300 1036 4308 1044
rect 4364 1036 4372 1044
rect 4556 1036 4564 1044
rect 4668 1036 4676 1044
rect 4796 1036 4804 1044
rect 4940 1036 4948 1044
rect 5052 1036 5060 1044
rect 5116 1036 5124 1044
rect 5244 1036 5252 1044
rect 5372 1036 5380 1044
rect 5516 1036 5524 1044
rect 12 976 20 984
rect 140 976 148 984
rect 332 976 340 984
rect 652 976 660 984
rect 1548 976 1556 984
rect 1724 976 1732 984
rect 1996 976 2004 984
rect 2108 976 2116 984
rect 2252 976 2260 984
rect 2316 976 2324 984
rect 2572 976 2580 984
rect 2684 976 2692 984
rect 2700 976 2708 984
rect 2812 976 2820 984
rect 2828 976 2836 984
rect 2940 976 2948 984
rect 3260 976 3268 984
rect 3324 976 3332 984
rect 3340 976 3348 984
rect 3404 976 3412 984
rect 3532 976 3540 984
rect 3788 976 3796 984
rect 3852 976 3860 984
rect 3964 976 3972 984
rect 3980 976 3988 984
rect 4092 976 4100 984
rect 4364 976 4372 984
rect 4604 976 4612 984
rect 4732 976 4740 984
rect 4860 976 4868 984
rect 4876 976 4884 984
rect 4988 976 4996 984
rect 5244 976 5252 984
rect 5436 976 5444 984
rect 5452 976 5460 984
rect 44 936 52 944
rect 124 956 132 964
rect 252 956 260 964
rect 316 956 324 964
rect 444 956 452 964
rect 508 956 516 964
rect 572 956 580 964
rect 764 956 772 964
rect 828 956 836 964
rect 908 956 916 964
rect 1020 956 1028 964
rect 108 936 116 944
rect 188 936 196 944
rect 236 936 244 944
rect 300 936 308 944
rect 380 936 388 944
rect 428 936 436 944
rect 492 936 500 944
rect 556 936 564 944
rect 588 936 596 944
rect 700 936 708 944
rect 748 936 756 944
rect 812 936 820 944
rect 844 936 852 944
rect 908 936 916 944
rect 958 936 966 944
rect 1004 936 1012 944
rect 1020 936 1028 944
rect 1148 956 1156 964
rect 1212 956 1220 964
rect 1052 936 1060 944
rect 1132 936 1140 944
rect 1148 936 1156 944
rect 1212 936 1220 944
rect 1260 936 1268 944
rect 1340 956 1348 964
rect 1404 956 1412 964
rect 1468 956 1476 964
rect 1484 956 1492 964
rect 1660 956 1668 964
rect 1676 956 1684 964
rect 1740 956 1748 964
rect 1804 956 1812 964
rect 1916 956 1924 964
rect 1980 956 1988 964
rect 2172 956 2180 964
rect 2236 956 2244 964
rect 2364 956 2372 964
rect 2428 956 2436 964
rect 2636 956 2644 964
rect 3084 956 3092 964
rect 1324 936 1332 944
rect 1388 936 1396 944
rect 1484 936 1492 944
rect 1500 936 1508 944
rect 1534 936 1542 944
rect 1596 936 1604 944
rect 1644 936 1652 944
rect 1692 936 1700 944
rect 1820 936 1828 944
rect 1900 936 1908 944
rect 1980 936 1988 944
rect 2060 936 2068 944
rect 2156 936 2164 944
rect 2220 936 2228 944
rect 2300 936 2308 944
rect 2348 936 2356 944
rect 2412 936 2420 944
rect 2492 936 2500 944
rect 2620 936 2628 944
rect 2652 936 2660 944
rect 2748 936 2756 944
rect 2876 936 2884 944
rect 2892 936 2900 944
rect 3004 936 3012 944
rect 3020 936 3028 944
rect 3100 936 3108 944
rect 3452 956 3460 964
rect 3468 956 3476 964
rect 3644 956 3652 964
rect 3660 956 3668 964
rect 3772 956 3780 964
rect 3836 956 3844 964
rect 4108 956 4116 964
rect 4236 956 4244 964
rect 4348 956 4356 964
rect 4428 956 4436 964
rect 4684 956 4692 964
rect 5052 956 5060 964
rect 5068 956 5076 964
rect 5132 956 5140 964
rect 3164 936 3172 944
rect 3276 936 3284 944
rect 3388 936 3396 944
rect 3436 936 3444 944
rect 3484 936 3492 944
rect 3628 936 3636 944
rect 3772 936 3780 944
rect 3820 936 3828 944
rect 3900 936 3908 944
rect 3916 936 3924 944
rect 4028 936 4036 944
rect 4044 936 4052 944
rect 4124 936 4132 944
rect 4252 936 4260 944
rect 4332 936 4340 944
rect 4412 936 4420 944
rect 4444 936 4452 944
rect 4556 936 4564 944
rect 4620 936 4628 944
rect 4700 936 4708 944
rect 4748 936 4756 944
rect 4924 936 4932 944
rect 4940 936 4948 944
rect 5036 936 5044 944
rect 5084 936 5092 944
rect 5148 936 5156 944
rect 5260 936 5268 944
rect 5372 936 5380 944
rect 5388 936 5396 944
rect 5500 936 5508 944
rect 636 916 644 924
rect 1868 916 1876 924
rect 2188 916 2196 924
rect 2444 916 2452 924
rect 2508 916 2516 924
rect 172 896 180 904
rect 364 896 372 904
rect 588 896 596 904
rect 684 896 692 904
rect 860 896 868 904
rect 1580 896 1588 904
rect 1932 896 1940 904
rect 2028 896 2036 904
rect 2076 896 2084 904
rect 2124 896 2132 904
rect 2284 896 2292 904
rect 2476 896 2484 904
rect 2556 896 2564 904
rect 2604 896 2612 904
rect 2732 896 2740 904
rect 460 876 468 884
rect 524 876 532 884
rect 892 876 900 884
rect 2748 876 2756 884
rect 3068 916 3076 924
rect 3708 916 3716 924
rect 4012 916 4020 924
rect 4220 916 4228 924
rect 4508 916 4516 924
rect 4668 916 4676 924
rect 4812 916 4820 924
rect 5196 916 5204 924
rect 2780 896 2788 904
rect 2876 896 2884 904
rect 2908 896 2916 904
rect 2956 896 2964 904
rect 3020 896 3028 904
rect 3036 896 3044 904
rect 3228 896 3236 904
rect 3292 896 3300 904
rect 3372 896 3380 904
rect 3564 896 3572 904
rect 3884 896 3892 904
rect 3932 896 3940 904
rect 4060 896 4068 904
rect 4220 896 4228 904
rect 4396 896 4404 904
rect 4636 896 4644 904
rect 4764 896 4772 904
rect 4828 896 4836 904
rect 4908 896 4916 904
rect 4956 896 4964 904
rect 5004 896 5012 904
rect 5116 896 5124 904
rect 5212 896 5220 904
rect 5276 896 5284 904
rect 5308 896 5316 904
rect 5356 896 5364 904
rect 5404 896 5412 904
rect 5484 896 5492 904
rect 3516 876 3524 884
rect 3724 856 3732 864
rect 4284 856 4292 864
rect 4300 856 4308 864
rect 4796 856 4804 864
rect 204 836 212 844
rect 396 836 404 844
rect 716 836 724 844
rect 780 836 788 844
rect 972 836 980 844
rect 1084 836 1092 844
rect 1100 836 1108 844
rect 1228 836 1236 844
rect 1356 836 1364 844
rect 1420 836 1428 844
rect 1612 836 1620 844
rect 1788 836 1796 844
rect 1852 836 1860 844
rect 2380 836 2388 844
rect 4156 836 4164 844
rect 4172 836 4180 844
rect 5180 836 5188 844
rect 5324 836 5332 844
rect 12 776 20 784
rect 396 776 404 784
rect 892 776 900 784
rect 1100 776 1108 784
rect 1340 776 1348 784
rect 1980 776 1988 784
rect 2172 776 2180 784
rect 2188 776 2196 784
rect 2444 776 2452 784
rect 2636 776 2644 784
rect 2764 776 2772 784
rect 2940 776 2948 784
rect 2956 776 2964 784
rect 3084 776 3092 784
rect 3196 776 3204 784
rect 3212 776 3220 784
rect 3516 776 3524 784
rect 4156 776 4164 784
rect 4412 776 4420 784
rect 5324 776 5332 784
rect 1228 756 1236 764
rect 1852 756 1860 764
rect 1996 756 2004 764
rect 3660 756 3668 764
rect 3900 756 3908 764
rect 4028 756 4036 764
rect 4620 756 4628 764
rect 4732 756 4740 764
rect 5260 756 5268 764
rect 188 716 196 724
rect 252 716 260 724
rect 284 716 292 724
rect 428 716 436 724
rect 460 736 468 744
rect 2876 736 2884 744
rect 3388 736 3396 744
rect 4172 736 4180 744
rect 4796 736 4804 744
rect 5244 736 5252 744
rect 5500 736 5508 744
rect 476 716 484 724
rect 540 716 548 724
rect 588 716 596 724
rect 700 716 708 724
rect 716 716 724 724
rect 796 716 804 724
rect 1132 716 1140 724
rect 1180 716 1188 724
rect 1260 716 1268 724
rect 1404 716 1412 724
rect 1436 716 1444 724
rect 1580 716 1588 724
rect 1884 716 1892 724
rect 2028 716 2036 724
rect 2140 716 2148 724
rect 2220 716 2228 724
rect 2268 716 2276 724
rect 2348 716 2356 724
rect 2412 716 2420 724
rect 2492 716 2500 724
rect 2540 716 2548 724
rect 2668 716 2676 724
rect 2716 716 2724 724
rect 2796 716 2804 724
rect 2844 716 2852 724
rect 2988 716 2996 724
rect 3020 716 3028 724
rect 3468 716 3476 724
rect 3772 716 3780 724
rect 3836 716 3844 724
rect 4124 716 4132 724
rect 4300 716 4308 724
rect 4316 716 4324 724
rect 4460 716 4468 724
rect 4508 716 4516 724
rect 4572 716 4580 724
rect 4652 716 4660 724
rect 4700 716 4708 724
rect 5036 716 5044 724
rect 5116 716 5124 724
rect 5180 716 5188 724
rect 5196 716 5204 724
rect 5356 716 5364 724
rect 5404 716 5412 724
rect 5468 716 5476 724
rect 1388 696 1396 704
rect 1548 696 1556 704
rect 2572 696 2580 704
rect 2908 696 2916 704
rect 3580 696 3588 704
rect 3852 696 3860 704
rect 3868 696 3876 704
rect 4860 696 4868 704
rect 4940 696 4948 704
rect 5132 696 5140 704
rect 5292 696 5300 704
rect 5452 696 5460 704
rect 108 676 116 684
rect 188 676 196 684
rect 252 676 260 684
rect 268 676 276 684
rect 348 676 356 684
rect 460 676 468 684
rect 524 676 532 684
rect 620 676 628 684
rect 700 676 708 684
rect 716 676 724 684
rect 780 676 788 684
rect 860 676 868 684
rect 906 676 914 684
rect 1004 676 1012 684
rect 60 656 68 664
rect 124 656 132 664
rect 332 656 340 664
rect 636 656 644 664
rect 844 656 852 664
rect 956 656 964 664
rect 1068 676 1076 684
rect 1148 676 1156 684
rect 1164 676 1172 684
rect 1276 676 1284 684
rect 1308 676 1316 684
rect 1404 676 1412 684
rect 1420 676 1428 684
rect 1532 676 1540 684
rect 1596 676 1604 684
rect 1628 676 1636 684
rect 1676 676 1684 684
rect 1756 676 1764 684
rect 1084 656 1092 664
rect 1292 656 1300 664
rect 1532 656 1540 664
rect 1612 656 1620 664
rect 1740 656 1748 664
rect 1820 676 1828 684
rect 1868 676 1876 684
rect 1948 676 1956 684
rect 2044 676 2052 684
rect 2092 676 2100 684
rect 2124 676 2132 684
rect 2236 676 2244 684
rect 2252 676 2260 684
rect 2364 676 2372 684
rect 2428 676 2436 684
rect 2492 676 2500 684
rect 2556 676 2564 684
rect 2604 676 2612 684
rect 2700 676 2708 684
rect 2812 676 2820 684
rect 2828 676 2836 684
rect 2892 676 2900 684
rect 3004 676 3012 684
rect 3052 676 3060 684
rect 3116 676 3124 684
rect 3164 676 3172 684
rect 3244 676 3252 684
rect 3292 676 3300 684
rect 3356 676 3364 684
rect 3420 676 3428 684
rect 3644 676 3652 684
rect 3692 676 3700 684
rect 3740 676 3748 684
rect 3804 676 3812 684
rect 3932 676 3940 684
rect 3966 676 3974 684
rect 3996 676 4004 684
rect 4060 676 4068 684
rect 4108 676 4116 684
rect 4204 676 4212 684
rect 4284 676 4292 684
rect 4300 676 4308 684
rect 4380 676 4388 684
rect 4476 676 4484 684
rect 4492 676 4500 684
rect 4556 676 4564 684
rect 4668 676 4676 684
rect 4684 676 4692 684
rect 4764 676 4772 684
rect 4828 676 4836 684
rect 4892 676 4900 684
rect 5052 676 5060 684
rect 5084 676 5092 684
rect 5180 676 5188 684
rect 5196 676 5204 684
rect 5308 676 5316 684
rect 5372 676 5380 684
rect 5388 676 5396 684
rect 1932 656 1940 664
rect 2108 656 2116 664
rect 2620 656 2628 664
rect 3068 656 3076 664
rect 3132 656 3140 664
rect 3148 656 3156 664
rect 3260 656 3268 664
rect 3276 656 3284 664
rect 3340 656 3348 664
rect 3404 656 3412 664
rect 3644 656 3652 664
rect 3708 656 3716 664
rect 3724 656 3732 664
rect 3788 656 3796 664
rect 3916 656 3924 664
rect 3980 656 3988 664
rect 4044 656 4052 664
rect 4220 656 4228 664
rect 4364 656 4372 664
rect 4748 656 4756 664
rect 4812 656 4820 664
rect 4876 656 4884 664
rect 5068 656 5076 664
rect 140 636 148 644
rect 204 636 212 644
rect 316 636 324 644
rect 380 636 388 644
rect 396 636 404 644
rect 508 636 516 644
rect 572 636 580 644
rect 652 636 660 644
rect 764 636 772 644
rect 828 636 836 644
rect 972 636 980 644
rect 1212 636 1220 644
rect 1356 636 1364 644
rect 1468 636 1476 644
rect 1484 636 1492 644
rect 1724 636 1732 644
rect 1916 636 1924 644
rect 2060 636 2068 644
rect 2300 636 2308 644
rect 2316 636 2324 644
rect 2380 636 2388 644
rect 2444 636 2452 644
rect 2508 636 2516 644
rect 2748 636 2756 644
rect 3532 636 3540 644
rect 4092 636 4100 644
rect 4236 636 4244 644
rect 4348 636 4356 644
rect 4428 636 4436 644
rect 4540 636 4548 644
rect 4604 636 4612 644
rect 4988 636 4996 644
rect 5004 636 5012 644
rect 5436 636 5444 644
rect 140 576 148 584
rect 204 576 212 584
rect 316 576 324 584
rect 460 576 468 584
rect 764 576 772 584
rect 908 576 916 584
rect 1228 576 1236 584
rect 1292 576 1300 584
rect 1532 576 1540 584
rect 2060 576 2068 584
rect 2172 576 2180 584
rect 2380 576 2388 584
rect 2492 576 2500 584
rect 2556 576 2564 584
rect 2956 576 2964 584
rect 3084 576 3092 584
rect 3148 576 3156 584
rect 3276 576 3284 584
rect 3388 576 3396 584
rect 3468 576 3476 584
rect 3772 576 3780 584
rect 3836 576 3844 584
rect 3964 576 3972 584
rect 4092 576 4100 584
rect 4220 576 4228 584
rect 4236 576 4244 584
rect 4348 576 4356 584
rect 4364 576 4372 584
rect 4556 576 4564 584
rect 4796 576 4804 584
rect 4876 576 4884 584
rect 5132 576 5140 584
rect 5500 576 5508 584
rect 60 556 68 564
rect 188 556 196 564
rect 332 556 340 564
rect 396 556 404 564
rect 524 556 532 564
rect 44 536 52 544
rect 124 536 132 544
rect 172 536 180 544
rect 252 536 260 544
rect 268 536 276 544
rect 348 536 356 544
rect 412 536 420 544
rect 508 536 516 544
rect 540 536 548 544
rect 604 536 612 544
rect 780 556 788 564
rect 972 556 980 564
rect 1036 556 1044 564
rect 1100 556 1108 564
rect 1340 556 1348 564
rect 1356 556 1364 564
rect 1420 556 1428 564
rect 1484 556 1492 564
rect 1596 556 1604 564
rect 1612 556 1620 564
rect 1676 556 1684 564
rect 1740 556 1748 564
rect 1852 556 1860 564
rect 1916 556 1924 564
rect 2108 556 2116 564
rect 668 536 676 544
rect 716 536 724 544
rect 796 536 804 544
rect 892 536 900 544
rect 956 536 964 544
rect 988 536 996 544
rect 1116 536 1124 544
rect 1164 536 1172 544
rect 1276 536 1284 544
rect 1324 536 1332 544
rect 1372 536 1380 544
rect 1436 536 1444 544
rect 1500 536 1508 544
rect 1580 536 1588 544
rect 1612 536 1620 544
rect 1692 536 1700 544
rect 1756 536 1764 544
rect 1790 536 1798 544
rect 1836 536 1844 544
rect 1916 536 1924 544
rect 1980 536 1988 544
rect 1996 536 2004 544
rect 2092 536 2100 544
rect 2124 536 2132 544
rect 2220 536 2228 544
rect 2300 556 2308 564
rect 2636 556 2644 564
rect 2748 556 2756 564
rect 3020 556 3028 564
rect 3212 556 3220 564
rect 3340 556 3348 564
rect 3452 556 3460 564
rect 3644 556 3652 564
rect 3660 556 3668 564
rect 3788 556 3796 564
rect 3852 556 3860 564
rect 3980 556 3988 564
rect 4156 556 4164 564
rect 4172 556 4180 564
rect 4540 556 4548 564
rect 4668 556 4676 564
rect 4732 556 4740 564
rect 4860 556 4868 564
rect 4988 556 4996 564
rect 5052 556 5060 564
rect 5068 556 5076 564
rect 5196 556 5204 564
rect 5308 556 5316 564
rect 5372 556 5380 564
rect 5388 556 5396 564
rect 2300 536 2308 544
rect 2364 536 2372 544
rect 2428 536 2436 544
rect 2444 536 2452 544
rect 2508 536 2516 544
rect 2620 536 2628 544
rect 2652 536 2660 544
rect 2686 536 2694 544
rect 2748 536 2756 544
rect 2812 536 2820 544
rect 2876 536 2884 544
rect 2892 536 2900 544
rect 3004 536 3012 544
rect 3036 536 3044 544
rect 3132 536 3140 544
rect 3196 536 3204 544
rect 3228 536 3236 544
rect 3262 536 3270 544
rect 3324 536 3332 544
rect 3356 536 3364 544
rect 3436 536 3444 544
rect 3516 536 3524 544
rect 3628 536 3636 544
rect 3676 536 3684 544
rect 3804 536 3812 544
rect 3868 536 3876 544
rect 3996 536 4004 544
rect 4140 536 4148 544
rect 4188 536 4196 544
rect 4300 536 4308 544
rect 4412 536 4420 544
rect 4476 536 4484 544
rect 4524 536 4532 544
rect 4604 536 4612 544
rect 4652 536 4660 544
rect 4682 536 4690 544
rect 4716 536 4724 544
rect 4732 536 4740 544
rect 4844 536 4852 544
rect 4924 536 4932 544
rect 4972 536 4980 544
rect 4988 536 4996 544
rect 5036 536 5044 544
rect 5084 536 5092 544
rect 5180 536 5188 544
rect 5212 536 5220 544
rect 5292 536 5300 544
rect 5356 536 5364 544
rect 5404 536 5412 544
rect 844 516 852 524
rect 1660 516 1668 524
rect 1932 516 1940 524
rect 2316 516 2324 524
rect 2572 516 2580 524
rect 2700 516 2708 524
rect 2764 516 2772 524
rect 3068 516 3076 524
rect 3404 516 3412 524
rect 3564 516 3572 524
rect 4060 516 4068 524
rect 4108 516 4116 524
rect 4284 516 4292 524
rect 5260 516 5268 524
rect 5324 516 5332 524
rect 5452 516 5460 524
rect 12 496 20 504
rect 108 496 116 504
rect 236 496 244 504
rect 284 496 292 504
rect 492 496 500 504
rect 732 496 740 504
rect 940 496 948 504
rect 1260 496 1268 504
rect 1964 496 1972 504
rect 2012 496 2020 504
rect 2124 496 2132 504
rect 2188 496 2196 504
rect 2348 496 2356 504
rect 2412 496 2420 504
rect 2460 496 2468 504
rect 2524 496 2532 504
rect 2604 496 2612 504
rect 2860 496 2868 504
rect 2908 496 2916 504
rect 2988 496 2996 504
rect 3116 496 3124 504
rect 3180 496 3188 504
rect 3308 496 3316 504
rect 3724 496 3732 504
rect 3916 496 3924 504
rect 4268 496 4276 504
rect 4316 496 4324 504
rect 4460 496 4468 504
rect 4492 496 4500 504
rect 4588 496 4596 504
rect 4764 496 4772 504
rect 4812 496 4820 504
rect 4908 496 4916 504
rect 5116 496 5124 504
rect 5164 496 5172 504
rect 5468 496 5476 504
rect 1212 476 1220 484
rect 5244 476 5252 484
rect 1404 456 1412 464
rect 76 436 84 444
rect 380 436 388 444
rect 444 436 452 444
rect 700 436 708 444
rect 828 436 836 444
rect 1084 436 1092 444
rect 1148 436 1156 444
rect 1468 436 1476 444
rect 1548 436 1556 444
rect 1724 436 1732 444
rect 1804 436 1812 444
rect 1868 436 1876 444
rect 2044 436 2052 444
rect 2940 436 2948 444
rect 4620 436 4628 444
rect 4940 436 4948 444
rect 5436 436 5444 444
rect 1612 376 1620 384
rect 2444 376 2452 384
rect 2700 376 2708 384
rect 2828 376 2836 384
rect 3004 376 3012 384
rect 3068 376 3076 384
rect 3132 376 3140 384
rect 3196 376 3204 384
rect 3404 376 3412 384
rect 3516 376 3524 384
rect 3580 376 3588 384
rect 3644 376 3652 384
rect 3708 376 3716 384
rect 3772 376 3780 384
rect 3900 376 3908 384
rect 4220 376 4228 384
rect 4348 376 4356 384
rect 4412 376 4420 384
rect 5132 376 5140 384
rect 5260 376 5268 384
rect 2508 356 2516 364
rect 2812 356 2820 364
rect 4236 356 4244 364
rect 5372 356 5380 364
rect 460 336 468 344
rect 572 336 580 344
rect 716 336 724 344
rect 2684 336 2692 344
rect 5388 336 5396 344
rect 28 316 36 324
rect 140 316 148 324
rect 300 316 308 324
rect 364 316 372 324
rect 492 316 500 324
rect 556 316 564 324
rect 1196 316 1204 324
rect 1212 316 1220 324
rect 1260 316 1268 324
rect 1356 316 1364 324
rect 1772 316 1780 324
rect 1948 316 1956 324
rect 2028 316 2036 324
rect 2124 316 2132 324
rect 2140 316 2148 324
rect 2204 316 2212 324
rect 2268 316 2276 324
rect 2412 316 2420 324
rect 2476 316 2484 324
rect 2620 316 2628 324
rect 2652 316 2660 324
rect 2748 316 2756 324
rect 2764 316 2772 324
rect 2780 316 2788 324
rect 2860 316 2868 324
rect 2956 316 2964 324
rect 3964 316 3972 324
rect 4268 316 4276 324
rect 4460 316 4468 324
rect 4636 316 4644 324
rect 4684 316 4692 324
rect 4892 316 4900 324
rect 4988 316 4996 324
rect 5100 316 5108 324
rect 5228 316 5236 324
rect 5292 316 5300 324
rect 5340 316 5348 324
rect 5420 316 5428 324
rect 1036 296 1044 304
rect 1100 296 1108 304
rect 1164 296 1172 304
rect 2236 296 2244 304
rect 3836 296 3844 304
rect 4012 296 4020 304
rect 4156 296 4164 304
rect 4476 296 4484 304
rect 4572 296 4580 304
rect 4620 296 4628 304
rect 4780 296 4788 304
rect 4796 296 4804 304
rect 4812 296 4820 304
rect 4924 296 4932 304
rect 12 276 20 284
rect 92 276 100 284
rect 172 276 180 284
rect 220 276 228 284
rect 254 276 262 284
rect 316 276 324 284
rect 380 276 388 284
rect 428 276 436 284
rect 508 276 516 284
rect 572 276 580 284
rect 620 276 628 284
rect 76 256 84 264
rect 188 256 196 264
rect 204 256 212 264
rect 444 256 452 264
rect 700 276 708 284
rect 748 276 756 284
rect 764 276 772 284
rect 812 276 820 284
rect 876 276 884 284
rect 924 276 932 284
rect 1068 276 1076 284
rect 1132 276 1140 284
rect 1212 276 1220 284
rect 1276 276 1284 284
rect 1324 276 1332 284
rect 1388 276 1396 284
rect 1436 276 1444 284
rect 1516 276 1524 284
rect 1564 276 1572 284
rect 1644 276 1652 284
rect 1692 276 1700 284
rect 1788 276 1796 284
rect 1852 276 1860 284
rect 1900 276 1908 284
rect 1932 276 1940 284
rect 2044 276 2052 284
rect 2108 276 2116 284
rect 2124 276 2132 284
rect 2188 276 2196 284
rect 2252 276 2260 284
rect 2316 276 2324 284
rect 2428 276 2436 284
rect 2492 276 2500 284
rect 2540 276 2548 284
rect 2588 276 2596 284
rect 2636 276 2644 284
rect 2748 276 2756 284
rect 2876 276 2884 284
rect 2908 276 2916 284
rect 3036 276 3044 284
rect 3084 276 3092 284
rect 3100 276 3108 284
rect 3164 276 3172 284
rect 3244 276 3252 284
rect 3292 276 3300 284
rect 3356 276 3364 284
rect 3436 276 3444 284
rect 3484 276 3492 284
rect 3548 276 3556 284
rect 3612 276 3620 284
rect 3676 276 3684 284
rect 3740 276 3748 284
rect 3804 276 3812 284
rect 3868 276 3876 284
rect 3932 276 3940 284
rect 4044 276 4052 284
rect 4060 276 4068 284
rect 4124 276 4132 284
rect 700 256 708 264
rect 764 256 772 264
rect 828 256 836 264
rect 892 256 900 264
rect 908 256 916 264
rect 972 256 980 264
rect 1084 256 1092 264
rect 1148 256 1156 264
rect 1340 256 1348 264
rect 1404 256 1412 264
rect 1420 256 1428 264
rect 1532 256 1540 264
rect 1548 256 1556 264
rect 1660 256 1668 264
rect 1676 256 1684 264
rect 1916 256 1924 264
rect 2316 256 2324 264
rect 2556 256 2564 264
rect 2572 256 2580 264
rect 2892 256 2900 264
rect 3020 256 3028 264
rect 3084 256 3092 264
rect 3148 256 3156 264
rect 3260 256 3268 264
rect 3276 256 3284 264
rect 3340 256 3348 264
rect 3452 256 3460 264
rect 3468 256 3476 264
rect 3532 256 3540 264
rect 3596 256 3604 264
rect 3660 256 3668 264
rect 3724 256 3732 264
rect 3788 256 3796 264
rect 3852 256 3860 264
rect 3916 256 3924 264
rect 4044 256 4052 264
rect 4108 256 4116 264
rect 4188 276 4196 284
rect 4284 276 4292 284
rect 4380 276 4388 284
rect 4508 276 4516 284
rect 4716 276 4724 284
rect 4844 276 4852 284
rect 4876 276 4884 284
rect 5036 276 5044 284
rect 5116 276 5124 284
rect 5164 276 5172 284
rect 5244 276 5252 284
rect 5308 276 5316 284
rect 5324 276 5332 284
rect 5436 276 5444 284
rect 5452 276 5460 284
rect 4300 256 4308 264
rect 4364 256 4372 264
rect 4492 256 4500 264
rect 4732 256 4740 264
rect 4860 256 4868 264
rect 5052 256 5060 264
rect 5180 256 5188 264
rect 5452 256 5460 264
rect 60 236 68 244
rect 124 236 132 244
rect 268 236 276 244
rect 332 236 340 244
rect 396 236 404 244
rect 524 236 532 244
rect 844 236 852 244
rect 1020 236 1028 244
rect 1292 236 1300 244
rect 1468 236 1476 244
rect 1484 236 1492 244
rect 1596 236 1604 244
rect 1612 236 1620 244
rect 1724 236 1732 244
rect 1740 236 1748 244
rect 1804 236 1812 244
rect 1980 236 1988 244
rect 1996 236 2004 244
rect 2060 236 2068 244
rect 2172 236 2180 244
rect 2300 236 2308 244
rect 2364 236 2372 244
rect 2380 236 2388 244
rect 3212 236 3220 244
rect 3324 236 3332 244
rect 3388 236 3396 244
rect 3580 236 3588 244
rect 3980 236 3988 244
rect 4092 236 4100 244
rect 4428 236 4436 244
rect 4604 236 4612 244
rect 4668 236 4676 244
rect 4748 236 4756 244
rect 4940 236 4948 244
rect 5068 236 5076 244
rect 5196 236 5204 244
rect 5500 236 5508 244
rect 12 176 20 184
rect 956 176 964 184
rect 1036 176 1044 184
rect 1212 176 1220 184
rect 1276 176 1284 184
rect 1660 176 1668 184
rect 2188 176 2196 184
rect 2572 176 2580 184
rect 2700 176 2708 184
rect 2764 176 2772 184
rect 2876 176 2884 184
rect 3068 176 3076 184
rect 3148 176 3156 184
rect 3516 176 3524 184
rect 3660 176 3668 184
rect 4044 176 4052 184
rect 4156 176 4164 184
rect 4796 176 4804 184
rect 5052 176 5060 184
rect 5068 176 5076 184
rect 5132 176 5140 184
rect 5244 176 5252 184
rect 5308 176 5316 184
rect 5436 176 5444 184
rect 5580 176 5588 184
rect 60 156 68 164
rect 76 156 84 164
rect 252 156 260 164
rect 268 156 276 164
rect 44 136 52 144
rect 92 136 100 144
rect 126 136 134 144
rect 188 136 196 144
rect 236 136 244 144
rect 284 136 292 144
rect 396 156 404 164
rect 508 156 516 164
rect 572 156 580 164
rect 588 156 596 164
rect 700 156 708 164
rect 716 156 724 164
rect 348 136 356 144
rect 492 136 500 144
rect 556 136 564 144
rect 604 136 612 144
rect 684 136 692 144
rect 732 136 740 144
rect 844 156 852 164
rect 1100 156 1108 164
rect 796 136 804 144
rect 860 136 868 144
rect 908 136 916 144
rect 972 136 980 144
rect 1084 136 1092 144
rect 1116 136 1124 144
rect 1228 156 1236 164
rect 1340 156 1348 164
rect 1404 156 1412 164
rect 1420 156 1428 164
rect 1180 136 1188 144
rect 1244 136 1252 144
rect 1324 136 1332 144
rect 1420 136 1428 144
rect 1436 136 1444 144
rect 1596 156 1604 164
rect 1612 156 1620 164
rect 1724 156 1732 164
rect 1788 156 1796 164
rect 1852 156 1860 164
rect 1868 156 1876 164
rect 1980 156 1988 164
rect 1500 136 1508 144
rect 1612 136 1620 144
rect 1628 136 1636 144
rect 1708 136 1716 144
rect 1772 136 1780 144
rect 1836 136 1844 144
rect 1884 136 1892 144
rect 1930 136 1938 144
rect 1964 136 1972 144
rect 1980 136 1988 144
rect 2108 156 2116 164
rect 2012 136 2020 144
rect 2046 136 2054 144
rect 2108 136 2116 144
rect 2172 136 2180 144
rect 2236 136 2244 144
rect 2284 136 2292 144
rect 2364 156 2372 164
rect 2428 156 2436 164
rect 2620 156 2628 164
rect 2892 156 2900 164
rect 2956 156 2964 164
rect 3020 156 3028 164
rect 3084 156 3092 164
rect 3324 156 3332 164
rect 3388 156 3396 164
rect 3404 156 3412 164
rect 3468 156 3476 164
rect 3596 156 3604 164
rect 3772 156 3780 164
rect 3788 156 3796 164
rect 3964 156 3972 164
rect 3980 156 3988 164
rect 4220 156 4228 164
rect 4236 156 4244 164
rect 4348 156 4356 164
rect 4428 156 4436 164
rect 4732 156 4740 164
rect 4924 156 4932 164
rect 4988 156 4996 164
rect 5324 156 5332 164
rect 2364 136 2372 144
rect 2428 136 2436 144
rect 2492 136 2500 144
rect 2556 136 2564 144
rect 2604 136 2612 144
rect 2684 136 2692 144
rect 2748 136 2756 144
rect 2812 136 2820 144
rect 2828 136 2836 144
rect 2908 136 2916 144
rect 2972 136 2980 144
rect 3006 136 3014 144
rect 3036 136 3044 144
rect 3100 136 3108 144
rect 3196 136 3204 144
rect 3308 136 3316 144
rect 3404 136 3412 144
rect 3420 136 3428 144
rect 3468 136 3476 144
rect 3580 136 3588 144
rect 3612 136 3620 144
rect 3756 136 3764 144
rect 3804 136 3812 144
rect 3948 136 3956 144
rect 3996 136 4004 144
rect 4108 136 4116 144
rect 4204 136 4212 144
rect 4252 136 4260 144
rect 4332 136 4340 144
rect 4444 136 4452 144
rect 4604 136 4612 144
rect 4668 136 4676 144
rect 4716 136 4724 144
rect 4908 136 4916 144
rect 4972 136 4980 144
rect 5004 136 5012 144
rect 5116 136 5124 144
rect 5180 136 5188 144
rect 5196 136 5204 144
rect 5260 136 5268 144
rect 5340 136 5348 144
rect 5452 136 5460 144
rect 140 116 148 124
rect 444 116 452 124
rect 652 116 660 124
rect 1020 116 1028 124
rect 2124 116 2132 124
rect 2444 116 2452 124
rect 2636 116 2644 124
rect 2796 116 2804 124
rect 524 96 532 104
rect 636 96 644 104
rect 924 96 932 104
rect 972 96 980 104
rect 1068 96 1076 104
rect 1292 96 1300 104
rect 1356 96 1364 104
rect 1548 96 1556 104
rect 1676 96 1684 104
rect 2060 96 2068 104
rect 2172 96 2180 104
rect 2220 96 2228 104
rect 2380 96 2388 104
rect 2476 96 2484 104
rect 2540 96 2548 104
rect 2668 96 2676 104
rect 2748 96 2756 104
rect 2844 116 2852 124
rect 2940 116 2948 124
rect 3260 116 3268 124
rect 3340 116 3348 124
rect 3532 116 3540 124
rect 4076 116 4084 124
rect 4364 116 4372 124
rect 4540 116 4548 124
rect 4684 116 4692 124
rect 4748 116 4756 124
rect 4812 116 4820 124
rect 4844 116 4852 124
rect 4940 116 4948 124
rect 5020 116 5028 124
rect 2812 96 2820 104
rect 5164 116 5172 124
rect 3132 96 3140 104
rect 3564 96 3572 104
rect 3692 96 3700 104
rect 3884 96 3892 104
rect 4028 96 4036 104
rect 4092 96 4100 104
rect 4172 96 4180 104
rect 4284 96 4292 104
rect 4300 96 4308 104
rect 4364 96 4372 104
rect 4412 96 4420 104
rect 4508 96 4516 104
rect 4588 96 4596 104
rect 4652 96 4660 104
rect 4764 96 4772 104
rect 5100 96 5108 104
rect 5212 96 5220 104
rect 5276 96 5284 104
rect 5404 96 5412 104
rect 5468 96 5476 104
rect 1804 76 1812 84
rect 1916 76 1924 84
rect 3452 76 3460 84
rect 3644 76 3652 84
rect 3836 76 3844 84
rect 1740 56 1748 64
rect 2252 56 2260 64
rect 3852 56 3860 64
rect 4620 56 4628 64
rect 460 36 468 44
rect 828 36 836 44
rect 1532 36 1540 44
rect 4556 36 4564 44
<< metal2 >>
rect 605 3984 611 4083
rect 861 3924 867 3956
rect 925 3924 931 3956
rect 1197 3924 1203 3996
rect 1517 3924 1523 3936
rect 221 3884 227 3916
rect 365 3884 371 3896
rect 29 3864 35 3876
rect 13 3844 19 3856
rect 68 3757 76 3763
rect 93 3744 99 3876
rect 212 3857 227 3863
rect 61 3737 76 3743
rect 13 3724 19 3736
rect 61 3724 67 3737
rect 29 3684 35 3696
rect 61 3584 67 3696
rect 109 3544 115 3836
rect 189 3784 195 3796
rect 125 3763 131 3776
rect 125 3757 140 3763
rect 141 3584 147 3736
rect 109 3524 115 3536
rect 77 3484 83 3496
rect 205 3484 211 3636
rect 180 3477 188 3483
rect 13 3384 19 3456
rect 125 3384 131 3476
rect 196 3457 211 3463
rect 205 3444 211 3457
rect 141 3404 147 3436
rect 173 3344 179 3396
rect 61 3324 67 3336
rect 77 3204 83 3236
rect 189 3084 195 3356
rect 221 3324 227 3857
rect 253 3764 259 3776
rect 260 3737 275 3743
rect 269 3724 275 3737
rect 269 3483 275 3496
rect 260 3477 275 3483
rect 285 3483 291 3876
rect 381 3864 387 3916
rect 685 3884 691 3896
rect 893 3884 899 3896
rect 1533 3884 1539 4083
rect 1741 3984 1747 3996
rect 1597 3884 1603 3936
rect 1709 3924 1715 3936
rect 820 3877 828 3883
rect 852 3877 860 3883
rect 1396 3877 1404 3883
rect 397 3844 403 3856
rect 413 3844 419 3876
rect 573 3864 579 3876
rect 461 3844 467 3856
rect 532 3777 540 3783
rect 573 3764 579 3776
rect 589 3764 595 3796
rect 365 3724 371 3736
rect 317 3704 323 3716
rect 301 3684 307 3696
rect 381 3524 387 3756
rect 445 3744 451 3756
rect 509 3704 515 3756
rect 557 3724 563 3736
rect 605 3704 611 3736
rect 621 3724 627 3876
rect 909 3864 915 3876
rect 836 3857 851 3863
rect 701 3844 707 3856
rect 765 3844 771 3856
rect 781 3823 787 3836
rect 765 3817 787 3823
rect 765 3764 771 3817
rect 781 3784 787 3796
rect 845 3784 851 3857
rect 980 3857 988 3863
rect 909 3784 915 3856
rect 957 3804 963 3836
rect 1133 3824 1139 3876
rect 1213 3864 1219 3876
rect 1277 3864 1283 3876
rect 1156 3857 1171 3863
rect 1165 3844 1171 3857
rect 1325 3804 1331 3876
rect 1341 3823 1347 3856
rect 1341 3817 1363 3823
rect 1101 3784 1107 3796
rect 1293 3784 1299 3796
rect 1357 3784 1363 3817
rect 1037 3763 1043 3776
rect 1028 3757 1043 3763
rect 701 3724 707 3756
rect 461 3524 467 3536
rect 381 3504 387 3516
rect 461 3484 467 3496
rect 285 3477 316 3483
rect 260 3337 275 3343
rect 269 3324 275 3337
rect 157 3077 172 3083
rect 61 3064 67 3076
rect 125 3064 131 3076
rect 13 2964 19 3036
rect 125 2964 131 2976
rect 141 2944 147 2956
rect 157 2944 163 3077
rect 205 3064 211 3236
rect 237 3104 243 3116
rect 269 3044 275 3056
rect 205 2983 211 3036
rect 285 2984 291 3316
rect 301 3304 307 3477
rect 333 3444 339 3456
rect 381 3384 387 3476
rect 397 3364 403 3436
rect 445 3344 451 3356
rect 349 3337 364 3343
rect 301 3284 307 3296
rect 317 3084 323 3336
rect 301 3064 307 3076
rect 317 2984 323 3036
rect 205 2977 227 2983
rect 189 2963 195 2976
rect 189 2957 204 2963
rect 221 2944 227 2977
rect 13 2904 19 2936
rect 61 2924 67 2936
rect 13 2664 19 2876
rect 109 2724 115 2936
rect 157 2904 163 2916
rect 148 2677 156 2683
rect 13 2264 19 2436
rect 29 2284 35 2676
rect 189 2657 204 2663
rect 189 2644 195 2657
rect 221 2643 227 2676
rect 205 2637 227 2643
rect 109 2544 115 2596
rect 125 2584 131 2636
rect 205 2584 211 2637
rect 141 2563 147 2576
rect 132 2557 147 2563
rect 205 2563 211 2576
rect 196 2557 211 2563
rect 45 2524 51 2536
rect 29 2023 35 2276
rect 77 2264 83 2436
rect 125 2324 131 2536
rect 237 2504 243 2956
rect 333 2944 339 3076
rect 349 3044 355 3337
rect 445 3337 446 3344
rect 413 3324 419 3336
rect 477 3324 483 3516
rect 493 3344 499 3376
rect 509 3364 515 3436
rect 525 3324 531 3336
rect 557 3324 563 3516
rect 605 3484 611 3536
rect 573 3464 579 3476
rect 589 3444 595 3456
rect 637 3384 643 3636
rect 669 3484 675 3596
rect 749 3584 755 3736
rect 829 3724 835 3736
rect 877 3704 883 3756
rect 893 3724 899 3736
rect 909 3724 915 3756
rect 957 3744 963 3756
rect 1092 3737 1100 3743
rect 1005 3724 1011 3736
rect 1133 3704 1139 3776
rect 1229 3763 1235 3776
rect 1220 3757 1235 3763
rect 1405 3763 1411 3856
rect 1421 3784 1427 3876
rect 1533 3864 1539 3876
rect 1469 3804 1475 3836
rect 1549 3804 1555 3836
rect 1485 3784 1491 3796
rect 1629 3784 1635 3816
rect 1597 3764 1603 3776
rect 1613 3764 1619 3776
rect 1405 3757 1427 3763
rect 1284 3737 1292 3743
rect 1149 3724 1155 3736
rect 813 3684 819 3696
rect 941 3684 947 3696
rect 973 3624 979 3636
rect 1069 3524 1075 3696
rect 989 3504 995 3516
rect 925 3477 940 3483
rect 701 3383 707 3436
rect 749 3424 755 3476
rect 765 3444 771 3456
rect 765 3423 771 3436
rect 765 3417 787 3423
rect 781 3384 787 3417
rect 813 3384 819 3476
rect 829 3423 835 3456
rect 893 3444 899 3456
rect 829 3417 851 3423
rect 845 3384 851 3417
rect 685 3377 707 3383
rect 685 3344 691 3377
rect 772 3357 780 3363
rect 749 3344 755 3356
rect 893 3344 899 3356
rect 813 3304 819 3316
rect 829 3304 835 3336
rect 884 3297 892 3303
rect 573 3264 579 3296
rect 397 3184 403 3256
rect 381 3084 387 3116
rect 461 3104 467 3236
rect 477 3124 483 3136
rect 397 3063 403 3096
rect 429 3064 435 3076
rect 461 3064 467 3076
rect 388 3057 403 3063
rect 381 2963 387 2976
rect 381 2957 396 2963
rect 260 2897 268 2903
rect 285 2684 291 2896
rect 445 2884 451 3056
rect 477 2944 483 3116
rect 516 3097 547 3103
rect 541 3083 547 3097
rect 541 3077 556 3083
rect 509 2944 515 3076
rect 573 3044 579 3056
rect 589 2964 595 2976
rect 605 2964 611 3276
rect 621 3144 627 3296
rect 813 3284 819 3296
rect 653 3164 659 3236
rect 669 3124 675 3136
rect 813 3124 819 3276
rect 637 3084 643 3116
rect 829 3103 835 3176
rect 829 3097 883 3103
rect 877 3084 883 3097
rect 797 3077 812 3083
rect 637 3044 643 3056
rect 653 2984 659 3076
rect 765 3044 771 3056
rect 701 2963 707 2976
rect 701 2957 716 2963
rect 525 2944 531 2956
rect 589 2944 595 2956
rect 605 2944 611 2956
rect 733 2944 739 2976
rect 461 2924 467 2936
rect 541 2924 547 2936
rect 653 2924 659 2936
rect 541 2904 547 2916
rect 509 2884 515 2896
rect 333 2844 339 2876
rect 301 2724 307 2776
rect 365 2724 371 2876
rect 445 2704 451 2836
rect 493 2724 499 2736
rect 541 2724 547 2776
rect 573 2724 579 2836
rect 653 2764 659 2916
rect 765 2804 771 2836
rect 797 2764 803 3077
rect 813 2904 819 2976
rect 877 2944 883 3076
rect 893 3044 899 3056
rect 909 2963 915 2976
rect 900 2957 915 2963
rect 845 2804 851 2836
rect 644 2717 780 2723
rect 413 2684 419 2696
rect 253 2644 259 2656
rect 269 2544 275 2616
rect 253 2404 259 2536
rect 285 2504 291 2676
rect 381 2624 387 2676
rect 397 2644 403 2656
rect 445 2583 451 2636
rect 445 2577 467 2583
rect 461 2564 467 2577
rect 493 2564 499 2716
rect 605 2704 611 2716
rect 925 2704 931 3477
rect 957 3423 963 3456
rect 973 3444 979 3476
rect 957 3417 979 3423
rect 973 3404 979 3417
rect 973 3384 979 3396
rect 957 3324 963 3336
rect 989 3324 995 3496
rect 1037 3464 1043 3476
rect 1021 3423 1027 3436
rect 1021 3417 1043 3423
rect 1037 3404 1043 3417
rect 1021 3344 1027 3396
rect 1037 3364 1043 3396
rect 1053 3384 1059 3516
rect 1133 3504 1139 3696
rect 1197 3624 1203 3736
rect 1261 3684 1267 3696
rect 1325 3664 1331 3696
rect 1405 3604 1411 3736
rect 1421 3724 1427 3757
rect 1629 3744 1635 3776
rect 1469 3704 1475 3736
rect 1533 3704 1539 3736
rect 1444 3697 1452 3703
rect 1357 3524 1363 3556
rect 1197 3504 1203 3516
rect 1124 3477 1139 3483
rect 1133 3463 1139 3477
rect 1133 3457 1171 3463
rect 1101 3444 1107 3456
rect 1165 3444 1171 3457
rect 1085 3424 1091 3436
rect 1133 3344 1139 3416
rect 1149 3364 1155 3436
rect 1053 3324 1059 3336
rect 941 3164 947 3296
rect 1005 3264 1011 3296
rect 1085 3224 1091 3236
rect 1101 3204 1107 3236
rect 957 3084 963 3136
rect 964 3057 979 3063
rect 941 2904 947 3056
rect 973 2984 979 3057
rect 941 2704 947 2896
rect 957 2884 963 2916
rect 573 2684 579 2696
rect 589 2684 595 2696
rect 637 2683 643 2696
rect 637 2677 652 2683
rect 724 2677 732 2683
rect 509 2604 515 2676
rect 525 2664 531 2676
rect 669 2663 675 2676
rect 781 2664 787 2676
rect 660 2657 675 2663
rect 701 2657 716 2663
rect 701 2644 707 2657
rect 797 2643 803 2656
rect 772 2637 803 2643
rect 317 2384 323 2556
rect 381 2384 387 2536
rect 477 2524 483 2536
rect 157 2324 163 2336
rect 61 2183 67 2236
rect 77 2203 83 2236
rect 77 2197 99 2203
rect 45 2177 67 2183
rect 45 2144 51 2177
rect 13 2017 35 2023
rect 13 1984 19 2017
rect 61 1944 67 2156
rect 45 1784 51 1876
rect 52 1757 60 1763
rect 77 1743 83 2036
rect 93 1883 99 2197
rect 93 1877 108 1883
rect 125 1763 131 1856
rect 125 1757 147 1763
rect 68 1737 83 1743
rect 109 1684 115 1696
rect 13 1603 19 1636
rect 77 1624 83 1636
rect 13 1597 35 1603
rect 13 1364 19 1436
rect 29 1344 35 1597
rect 109 1484 115 1616
rect 141 1584 147 1757
rect 45 1204 51 1476
rect 125 1464 131 1476
rect 77 1364 83 1436
rect 125 1423 131 1456
rect 125 1417 147 1423
rect 141 1384 147 1417
rect 132 1357 140 1363
rect 109 1344 115 1356
rect 157 1303 163 2276
rect 189 2184 195 2236
rect 173 2177 188 2183
rect 173 2144 179 2177
rect 205 2163 211 2176
rect 196 2157 211 2163
rect 221 2084 227 2316
rect 253 2283 259 2296
rect 349 2284 355 2316
rect 253 2277 268 2283
rect 269 2184 275 2256
rect 317 2164 323 2176
rect 301 2144 307 2156
rect 333 2143 339 2256
rect 365 2144 371 2356
rect 381 2304 387 2376
rect 397 2264 403 2436
rect 493 2284 499 2296
rect 413 2264 419 2276
rect 509 2264 515 2296
rect 525 2264 531 2436
rect 541 2364 547 2596
rect 557 2544 563 2616
rect 829 2584 835 2636
rect 877 2584 883 2676
rect 893 2644 899 2656
rect 941 2644 947 2676
rect 957 2664 963 2736
rect 989 2644 995 3116
rect 1037 3084 1043 3096
rect 1053 3064 1059 3116
rect 1108 3097 1116 3103
rect 1133 3064 1139 3076
rect 1156 3057 1164 3063
rect 1021 2984 1027 3036
rect 1085 3004 1091 3036
rect 1085 2963 1091 2976
rect 1085 2957 1100 2963
rect 1037 2944 1043 2956
rect 1165 2944 1171 3036
rect 1021 2924 1027 2936
rect 1021 2724 1027 2896
rect 1053 2884 1059 2896
rect 909 2604 915 2636
rect 573 2564 579 2576
rect 893 2564 899 2576
rect 973 2564 979 2636
rect 653 2544 659 2556
rect 701 2544 707 2556
rect 749 2544 755 2556
rect 893 2544 899 2556
rect 989 2544 995 2556
rect 701 2537 702 2544
rect 717 2404 723 2436
rect 621 2284 627 2356
rect 461 2244 467 2256
rect 445 2183 451 2236
rect 429 2177 451 2183
rect 429 2144 435 2177
rect 509 2164 515 2176
rect 445 2144 451 2156
rect 317 2137 339 2143
rect 253 2124 259 2136
rect 221 1924 227 2076
rect 317 1984 323 2137
rect 349 2123 355 2136
rect 541 2123 547 2276
rect 637 2264 643 2376
rect 692 2317 700 2323
rect 740 2317 748 2323
rect 701 2284 707 2296
rect 765 2284 771 2336
rect 797 2324 803 2336
rect 813 2324 819 2536
rect 877 2524 883 2536
rect 957 2524 963 2536
rect 893 2384 899 2396
rect 829 2283 835 2296
rect 829 2277 844 2283
rect 781 2264 787 2276
rect 573 2163 579 2176
rect 573 2157 588 2163
rect 605 2144 611 2196
rect 621 2183 627 2216
rect 637 2204 643 2256
rect 653 2184 659 2236
rect 621 2177 636 2183
rect 653 2164 659 2176
rect 717 2164 723 2176
rect 660 2137 668 2143
rect 340 2117 355 2123
rect 525 2117 547 2123
rect 525 1984 531 2117
rect 173 1857 188 1863
rect 173 1504 179 1857
rect 189 1744 195 1756
rect 189 1484 195 1696
rect 205 1584 211 1616
rect 221 1463 227 1916
rect 349 1904 355 1916
rect 621 1904 627 1916
rect 653 1884 659 2096
rect 733 1964 739 2176
rect 765 2144 771 2156
rect 813 2144 819 2236
rect 845 2224 851 2256
rect 845 2164 851 2176
rect 925 2124 931 2316
rect 941 2284 947 2316
rect 957 2284 963 2296
rect 973 2284 979 2536
rect 1005 2264 1011 2716
rect 1021 2644 1027 2676
rect 1037 2584 1043 2636
rect 1053 2604 1059 2876
rect 1149 2864 1155 2876
rect 1069 2664 1075 2716
rect 1181 2704 1187 3336
rect 1197 3284 1203 3496
rect 1213 3404 1219 3476
rect 1229 3383 1235 3436
rect 1229 3377 1251 3383
rect 1245 3344 1251 3377
rect 1245 3324 1251 3336
rect 1261 3284 1267 3516
rect 1485 3484 1491 3596
rect 1501 3524 1507 3556
rect 1341 3464 1347 3476
rect 1405 3457 1420 3463
rect 1405 3444 1411 3457
rect 1293 3424 1299 3436
rect 1293 3364 1299 3376
rect 1405 3364 1411 3396
rect 1437 3384 1443 3476
rect 1309 3344 1315 3356
rect 1412 3337 1427 3343
rect 1421 3324 1427 3337
rect 1453 3304 1459 3476
rect 1517 3464 1523 3696
rect 1549 3564 1555 3636
rect 1581 3544 1587 3736
rect 1645 3664 1651 3916
rect 1661 3884 1667 3896
rect 1661 3784 1667 3796
rect 1677 3764 1683 3836
rect 1725 3804 1731 3876
rect 1677 3544 1683 3696
rect 1741 3544 1747 3736
rect 1757 3684 1763 3696
rect 1661 3537 1676 3543
rect 1661 3504 1667 3537
rect 1757 3523 1763 3656
rect 1773 3543 1779 3916
rect 1789 3884 1795 3976
rect 1853 3944 1859 3956
rect 1965 3924 1971 4083
rect 1981 4077 2003 4083
rect 1981 3884 1987 4077
rect 2013 3944 2019 3976
rect 2093 3964 2099 4083
rect 2013 3924 2019 3936
rect 1853 3804 1859 3876
rect 1805 3764 1811 3776
rect 1869 3764 1875 3776
rect 1885 3744 1891 3756
rect 1828 3697 1836 3703
rect 1773 3537 1795 3543
rect 1757 3517 1772 3523
rect 1565 3497 1612 3503
rect 1565 3484 1571 3497
rect 1549 3444 1555 3456
rect 1533 3384 1539 3436
rect 1549 3384 1555 3396
rect 1469 3324 1475 3336
rect 1453 3284 1459 3296
rect 1197 3124 1203 3236
rect 1213 3104 1219 3136
rect 1261 3124 1267 3136
rect 1277 3104 1283 3236
rect 1533 3204 1539 3336
rect 1581 3304 1587 3476
rect 1597 3404 1603 3436
rect 1645 3384 1651 3476
rect 1677 3464 1683 3476
rect 1661 3424 1667 3456
rect 1693 3444 1699 3516
rect 1789 3484 1795 3537
rect 1821 3524 1827 3536
rect 1821 3504 1827 3516
rect 1805 3484 1811 3496
rect 1725 3424 1731 3436
rect 1741 3404 1747 3436
rect 1613 3364 1619 3376
rect 1773 3344 1779 3416
rect 1805 3364 1811 3396
rect 1581 3224 1587 3296
rect 1364 3137 1372 3143
rect 1325 3084 1331 3136
rect 1389 3084 1395 3096
rect 1453 3084 1459 3096
rect 1533 3084 1539 3096
rect 1597 3084 1603 3336
rect 1677 3324 1683 3336
rect 1700 3297 1708 3303
rect 1661 3124 1667 3236
rect 1725 3204 1731 3316
rect 1789 3184 1795 3356
rect 1837 3344 1843 3696
rect 1885 3524 1891 3656
rect 1869 3484 1875 3496
rect 1853 3424 1859 3436
rect 1885 3324 1891 3336
rect 1732 3177 1740 3183
rect 1284 3057 1299 3063
rect 1293 3044 1299 3057
rect 1476 3057 1491 3063
rect 1229 3004 1235 3036
rect 1229 2963 1235 2976
rect 1220 2957 1235 2963
rect 1261 2944 1267 2976
rect 1204 2937 1212 2943
rect 1277 2864 1283 2956
rect 1309 2944 1315 3056
rect 1341 3044 1347 3056
rect 1485 3044 1491 3057
rect 1485 3004 1491 3036
rect 1549 3024 1555 3036
rect 1405 2963 1411 2976
rect 1405 2957 1420 2963
rect 1437 2944 1443 2956
rect 1501 2944 1507 2976
rect 1549 2964 1555 2996
rect 1565 2944 1571 3036
rect 1597 3024 1603 3076
rect 1629 3044 1635 3116
rect 1700 3077 1715 3083
rect 1661 3057 1676 3063
rect 1661 3044 1667 3057
rect 1709 3063 1715 3077
rect 1709 3057 1747 3063
rect 1741 3044 1747 3057
rect 1613 2964 1619 2976
rect 1213 2784 1219 2796
rect 1108 2697 1116 2703
rect 1085 2684 1091 2696
rect 1261 2684 1267 2756
rect 1325 2684 1331 2696
rect 1085 2664 1091 2676
rect 1149 2664 1155 2676
rect 1149 2644 1155 2656
rect 1165 2584 1171 2656
rect 1229 2644 1235 2676
rect 1357 2664 1363 2876
rect 1501 2764 1507 2776
rect 1501 2724 1507 2756
rect 1373 2684 1379 2696
rect 1533 2684 1539 2836
rect 1565 2804 1571 2936
rect 1549 2684 1555 2716
rect 1565 2684 1571 2716
rect 1597 2684 1603 2836
rect 1277 2644 1283 2656
rect 1341 2644 1347 2656
rect 1357 2644 1363 2656
rect 1053 2523 1059 2556
rect 1069 2544 1075 2576
rect 1085 2544 1091 2556
rect 1044 2517 1059 2523
rect 1101 2404 1107 2556
rect 1117 2444 1123 2536
rect 1165 2444 1171 2556
rect 1181 2544 1187 2636
rect 1405 2604 1411 2636
rect 1236 2557 1244 2563
rect 1277 2563 1283 2576
rect 1421 2564 1427 2676
rect 1469 2624 1475 2636
rect 1277 2557 1292 2563
rect 1437 2557 1468 2563
rect 1229 2523 1235 2536
rect 1261 2523 1267 2556
rect 1309 2544 1315 2556
rect 1341 2544 1347 2556
rect 1341 2537 1342 2544
rect 1229 2517 1267 2523
rect 1389 2523 1395 2556
rect 1437 2523 1443 2557
rect 1469 2523 1475 2536
rect 1389 2517 1443 2523
rect 1453 2517 1475 2523
rect 1421 2424 1427 2436
rect 1133 2304 1139 2316
rect 1181 2277 1196 2283
rect 973 2244 979 2256
rect 1021 2184 1027 2236
rect 1069 2204 1075 2276
rect 1092 2257 1107 2263
rect 1101 2244 1107 2257
rect 1101 2184 1107 2196
rect 980 2177 988 2183
rect 1037 2163 1043 2176
rect 1028 2157 1043 2163
rect 1085 2144 1091 2176
rect 1149 2164 1155 2276
rect 1165 2224 1171 2236
rect 989 2137 1004 2143
rect 989 2123 995 2137
rect 964 2117 995 2123
rect 1069 2104 1075 2116
rect 749 2064 755 2096
rect 909 2084 915 2096
rect 1133 2084 1139 2096
rect 1149 2084 1155 2136
rect 285 1864 291 1876
rect 253 1857 268 1863
rect 253 1844 259 1857
rect 413 1843 419 1876
rect 397 1837 419 1843
rect 381 1824 387 1836
rect 317 1764 323 1776
rect 333 1764 339 1776
rect 253 1704 259 1756
rect 349 1744 355 1816
rect 397 1784 403 1837
rect 461 1803 467 1836
rect 445 1797 467 1803
rect 301 1724 307 1736
rect 397 1543 403 1636
rect 381 1537 403 1543
rect 317 1464 323 1476
rect 221 1457 243 1463
rect 189 1324 195 1336
rect 157 1297 172 1303
rect 61 1224 67 1236
rect 77 1223 83 1236
rect 77 1217 99 1223
rect 77 1184 83 1196
rect 13 984 19 1056
rect 93 943 99 1217
rect 141 1184 147 1196
rect 173 1104 179 1296
rect 205 1204 211 1356
rect 237 1164 243 1457
rect 253 1384 259 1456
rect 365 1384 371 1476
rect 381 1464 387 1537
rect 413 1524 419 1796
rect 445 1784 451 1797
rect 445 1764 451 1776
rect 461 1743 467 1776
rect 509 1744 515 1876
rect 557 1784 563 1876
rect 573 1764 579 1856
rect 589 1844 595 1856
rect 653 1823 659 1856
rect 669 1844 675 1876
rect 749 1864 755 1876
rect 781 1864 787 2036
rect 1101 2024 1107 2036
rect 1165 2004 1171 2036
rect 845 1984 851 1996
rect 1181 1964 1187 2277
rect 1261 2264 1267 2276
rect 1284 2257 1299 2263
rect 1197 2144 1203 2256
rect 1293 2244 1299 2257
rect 1213 2164 1219 2176
rect 1229 2144 1235 2156
rect 1229 2104 1235 2136
rect 1245 2084 1251 2096
rect 797 1884 803 1956
rect 1069 1924 1075 1936
rect 909 1917 963 1923
rect 765 1844 771 1856
rect 685 1823 691 1836
rect 653 1817 691 1823
rect 701 1764 707 1836
rect 829 1764 835 1776
rect 644 1757 668 1763
rect 685 1744 691 1756
rect 452 1737 467 1743
rect 461 1724 467 1737
rect 621 1724 627 1736
rect 500 1697 508 1703
rect 397 1484 403 1516
rect 397 1363 403 1376
rect 388 1357 403 1363
rect 269 1324 275 1336
rect 285 1164 291 1296
rect 381 1284 387 1336
rect 221 1084 227 1096
rect 349 1084 355 1116
rect 109 1004 115 1076
rect 173 1064 179 1076
rect 205 1064 211 1076
rect 132 1057 140 1063
rect 189 1024 195 1056
rect 141 984 147 996
rect 132 957 140 963
rect 93 937 108 943
rect 180 937 188 943
rect 45 804 51 936
rect 173 884 179 896
rect 13 784 19 796
rect 61 664 67 816
rect 205 704 211 836
rect 221 684 227 1076
rect 301 1064 307 1076
rect 317 1044 323 1056
rect 333 1024 339 1056
rect 237 944 243 1016
rect 381 984 387 1036
rect 333 963 339 976
rect 397 964 403 1036
rect 413 964 419 1516
rect 589 1504 595 1636
rect 493 1464 499 1476
rect 580 1457 588 1463
rect 445 1383 451 1436
rect 445 1377 467 1383
rect 461 1363 467 1377
rect 573 1364 579 1376
rect 461 1357 499 1363
rect 493 1344 499 1357
rect 621 1344 627 1536
rect 637 1484 643 1496
rect 653 1484 659 1636
rect 717 1604 723 1756
rect 733 1724 739 1736
rect 781 1724 787 1736
rect 765 1484 771 1556
rect 829 1524 835 1536
rect 829 1484 835 1496
rect 637 1364 643 1436
rect 653 1384 659 1456
rect 845 1424 851 1436
rect 701 1364 707 1376
rect 717 1364 723 1376
rect 845 1364 851 1376
rect 532 1337 540 1343
rect 477 1124 483 1316
rect 541 1304 547 1316
rect 445 1084 451 1116
rect 461 1064 467 1076
rect 445 964 451 976
rect 509 964 515 1036
rect 324 957 339 963
rect 301 944 307 956
rect 381 924 387 936
rect 253 724 259 776
rect 285 724 291 896
rect 413 884 419 956
rect 429 884 435 936
rect 397 784 403 796
rect 429 724 435 736
rect 445 723 451 936
rect 461 744 467 756
rect 477 724 483 736
rect 445 717 467 723
rect 269 684 275 696
rect 45 544 51 656
rect 109 604 115 676
rect 333 664 339 716
rect 461 684 467 717
rect 205 644 211 656
rect 141 623 147 636
rect 141 617 163 623
rect 61 564 67 576
rect 13 264 19 276
rect 45 264 51 536
rect 77 284 83 436
rect 93 284 99 596
rect 141 584 147 596
rect 157 543 163 617
rect 205 563 211 576
rect 196 557 211 563
rect 253 544 259 556
rect 269 544 275 656
rect 349 644 355 676
rect 317 584 323 616
rect 317 563 323 576
rect 317 557 332 563
rect 381 563 387 636
rect 397 583 403 636
rect 461 584 467 636
rect 397 577 419 583
rect 381 557 396 563
rect 413 544 419 577
rect 157 537 172 543
rect 493 504 499 836
rect 541 743 547 1296
rect 589 1203 595 1236
rect 589 1197 611 1203
rect 557 1124 563 1156
rect 573 964 579 976
rect 557 944 563 956
rect 589 944 595 956
rect 589 884 595 896
rect 525 737 547 743
rect 525 684 531 737
rect 557 723 563 776
rect 548 717 563 723
rect 605 683 611 1197
rect 621 1084 627 1136
rect 637 1083 643 1276
rect 637 1077 659 1083
rect 653 1064 659 1077
rect 637 1024 643 1056
rect 669 1043 675 1076
rect 653 1037 675 1043
rect 653 984 659 1037
rect 685 944 691 1336
rect 813 1264 819 1296
rect 749 1124 755 1136
rect 829 1124 835 1276
rect 861 1124 867 1896
rect 877 1884 883 1896
rect 909 1884 915 1917
rect 957 1904 963 1917
rect 1053 1917 1068 1923
rect 925 1884 931 1896
rect 1021 1884 1027 1896
rect 973 1844 979 1856
rect 957 1784 963 1836
rect 1053 1823 1059 1917
rect 1197 1903 1203 1996
rect 1197 1897 1219 1903
rect 1213 1884 1219 1897
rect 1181 1877 1196 1883
rect 1085 1864 1091 1876
rect 1069 1843 1075 1856
rect 1101 1843 1107 1856
rect 1117 1844 1123 1876
rect 1181 1863 1187 1877
rect 1245 1864 1251 1876
rect 1149 1857 1187 1863
rect 1197 1857 1228 1863
rect 1149 1844 1155 1857
rect 1069 1837 1107 1843
rect 1037 1817 1059 1823
rect 1037 1784 1043 1817
rect 893 1744 899 1756
rect 925 1737 940 1743
rect 893 1364 899 1436
rect 900 1337 915 1343
rect 909 1324 915 1337
rect 909 1284 915 1316
rect 925 1203 931 1737
rect 957 1704 963 1756
rect 1005 1744 1011 1776
rect 1021 1764 1027 1776
rect 1165 1764 1171 1776
rect 1181 1744 1187 1756
rect 973 1483 979 1636
rect 1069 1623 1075 1696
rect 1053 1617 1075 1623
rect 1005 1524 1011 1536
rect 1021 1484 1027 1516
rect 973 1477 995 1483
rect 941 1464 947 1476
rect 964 1457 972 1463
rect 973 1384 979 1396
rect 957 1344 963 1356
rect 957 1204 963 1336
rect 909 1197 931 1203
rect 909 1184 915 1197
rect 973 1124 979 1236
rect 868 1117 883 1123
rect 701 1024 707 1036
rect 717 1024 723 1036
rect 749 944 755 1056
rect 829 1044 835 1076
rect 845 1024 851 1076
rect 765 964 771 996
rect 637 924 643 936
rect 685 764 691 896
rect 701 724 707 816
rect 717 724 723 836
rect 781 784 787 836
rect 797 743 803 956
rect 813 944 819 996
rect 829 964 835 1016
rect 845 944 851 996
rect 861 904 867 1076
rect 877 784 883 1117
rect 973 1084 979 1096
rect 941 1064 947 1076
rect 893 943 899 1036
rect 957 1024 963 1056
rect 989 1004 995 1477
rect 1005 1344 1011 1376
rect 1021 1364 1027 1396
rect 1053 1364 1059 1617
rect 1069 1524 1075 1536
rect 1085 1484 1091 1736
rect 1101 1664 1107 1736
rect 1124 1697 1132 1703
rect 1133 1684 1139 1696
rect 1117 1484 1123 1536
rect 1181 1504 1187 1736
rect 1197 1644 1203 1857
rect 1229 1744 1235 1836
rect 1229 1544 1235 1736
rect 1197 1524 1203 1536
rect 1245 1524 1251 1596
rect 1213 1484 1219 1496
rect 1229 1484 1235 1516
rect 1085 1364 1091 1376
rect 1101 1364 1107 1416
rect 1069 1344 1075 1356
rect 1037 1264 1043 1276
rect 1085 1224 1091 1356
rect 1117 1344 1123 1436
rect 1069 1124 1075 1136
rect 1005 963 1011 1116
rect 1085 1084 1091 1196
rect 1101 1084 1107 1336
rect 1133 1223 1139 1456
rect 1213 1364 1219 1376
rect 1156 1336 1162 1344
rect 1170 1337 1171 1343
rect 1188 1337 1196 1343
rect 1229 1284 1235 1356
rect 1245 1344 1251 1436
rect 1261 1384 1267 2196
rect 1277 2184 1283 2216
rect 1293 2184 1299 2196
rect 1325 2104 1331 2316
rect 1357 2284 1363 2396
rect 1341 2264 1347 2276
rect 1428 2257 1443 2263
rect 1357 2244 1363 2256
rect 1405 2204 1411 2236
rect 1421 2184 1427 2236
rect 1437 2224 1443 2257
rect 1453 2244 1459 2517
rect 1485 2484 1491 2496
rect 1501 2324 1507 2596
rect 1533 2564 1539 2636
rect 1597 2603 1603 2636
rect 1581 2597 1603 2603
rect 1533 2544 1539 2556
rect 1485 2284 1491 2316
rect 1549 2284 1555 2556
rect 1581 2543 1587 2597
rect 1629 2563 1635 2796
rect 1645 2724 1651 3016
rect 1725 2964 1731 2976
rect 1732 2937 1747 2943
rect 1741 2924 1747 2937
rect 1661 2764 1667 2836
rect 1741 2784 1747 2796
rect 1645 2684 1651 2716
rect 1757 2684 1763 3176
rect 1789 3144 1795 3176
rect 1837 3124 1843 3136
rect 1773 3044 1779 3116
rect 1789 3104 1795 3116
rect 1789 3084 1795 3096
rect 1773 2904 1779 2996
rect 1789 2963 1795 3076
rect 1789 2957 1811 2963
rect 1805 2944 1811 2957
rect 1837 2944 1843 3116
rect 1869 3064 1875 3156
rect 1901 3083 1907 3756
rect 1949 3744 1955 3776
rect 1965 3563 1971 3876
rect 1997 3864 2003 3876
rect 2029 3763 2035 3956
rect 2093 3944 2099 3956
rect 2157 3944 2163 4083
rect 2093 3924 2099 3936
rect 2157 3924 2163 3936
rect 2285 3924 2291 4083
rect 2285 3904 2291 3916
rect 2173 3864 2179 3876
rect 2285 3864 2291 3896
rect 2317 3864 2323 3916
rect 2333 3844 2339 3876
rect 2381 3864 2387 3956
rect 2461 3904 2467 4083
rect 2557 4063 2563 4083
rect 2557 4057 2579 4063
rect 2397 3884 2403 3896
rect 2045 3824 2051 3836
rect 2061 3763 2067 3836
rect 2029 3757 2051 3763
rect 2061 3757 2083 3763
rect 2045 3744 2051 3757
rect 2077 3704 2083 3757
rect 2125 3724 2131 3836
rect 2237 3804 2243 3836
rect 2173 3744 2179 3796
rect 2237 3743 2243 3796
rect 2237 3737 2252 3743
rect 2189 3723 2195 3736
rect 2157 3717 2195 3723
rect 2029 3644 2035 3696
rect 1981 3584 1987 3636
rect 1997 3604 2003 3636
rect 1965 3557 1987 3563
rect 1965 3524 1971 3536
rect 1981 3504 1987 3557
rect 2029 3524 2035 3636
rect 1981 3484 1987 3496
rect 2045 3484 2051 3696
rect 2077 3544 2083 3696
rect 2077 3524 2083 3536
rect 1933 3404 1939 3436
rect 1997 3404 2003 3436
rect 2029 3344 2035 3416
rect 2061 3363 2067 3376
rect 2052 3357 2067 3363
rect 1965 3304 1971 3316
rect 1933 3084 1939 3196
rect 1965 3084 1971 3296
rect 1981 3204 1987 3336
rect 2061 3324 2067 3357
rect 2093 3304 2099 3676
rect 2109 3644 2115 3716
rect 2125 3664 2131 3716
rect 2109 3604 2115 3636
rect 2125 3464 2131 3636
rect 2157 3564 2163 3717
rect 2260 3697 2268 3703
rect 2157 3524 2163 3556
rect 2173 3484 2179 3696
rect 2189 3683 2195 3696
rect 2189 3677 2211 3683
rect 2189 3484 2195 3656
rect 2205 3524 2211 3677
rect 2253 3524 2259 3676
rect 2285 3563 2291 3836
rect 2381 3824 2387 3856
rect 2397 3804 2403 3876
rect 2317 3764 2323 3776
rect 2429 3764 2435 3816
rect 2429 3744 2435 3756
rect 2301 3724 2307 3736
rect 2349 3704 2355 3736
rect 2365 3724 2371 3736
rect 2285 3557 2307 3563
rect 2285 3524 2291 3536
rect 2301 3524 2307 3557
rect 2173 3464 2179 3476
rect 2109 3384 2115 3436
rect 2125 3404 2131 3436
rect 2189 3363 2195 3376
rect 2180 3357 2195 3363
rect 2157 3324 2163 3336
rect 1997 3204 2003 3236
rect 1988 3157 1996 3163
rect 2077 3084 2083 3096
rect 1892 3077 1907 3083
rect 1869 2984 1875 2996
rect 1805 2924 1811 2936
rect 1805 2804 1811 2896
rect 1837 2764 1843 2936
rect 1773 2724 1779 2736
rect 1805 2684 1811 2756
rect 1821 2724 1827 2736
rect 1821 2704 1827 2716
rect 1661 2664 1667 2676
rect 1677 2644 1683 2656
rect 1725 2564 1731 2636
rect 1853 2604 1859 2636
rect 1869 2604 1875 2636
rect 1789 2564 1795 2596
rect 1620 2557 1635 2563
rect 1853 2544 1859 2556
rect 1572 2537 1587 2543
rect 1796 2537 1804 2543
rect 1805 2524 1811 2536
rect 1597 2384 1603 2436
rect 1661 2364 1667 2436
rect 1741 2403 1747 2436
rect 1741 2397 1763 2403
rect 1645 2297 1676 2303
rect 1645 2284 1651 2297
rect 1709 2284 1715 2376
rect 1572 2277 1610 2283
rect 1618 2277 1619 2283
rect 1725 2264 1731 2276
rect 1549 2244 1555 2256
rect 1661 2244 1667 2256
rect 1533 2183 1539 2236
rect 1725 2223 1731 2256
rect 1725 2217 1747 2223
rect 1517 2177 1539 2183
rect 1421 2163 1427 2176
rect 1412 2157 1427 2163
rect 1469 2144 1475 2156
rect 1517 2144 1523 2177
rect 1540 2157 1548 2163
rect 1581 2144 1587 2196
rect 1597 2164 1603 2216
rect 1661 2164 1667 2196
rect 1741 2184 1747 2217
rect 1725 2164 1731 2176
rect 1716 2137 1724 2143
rect 1341 2104 1347 2136
rect 1293 1984 1299 2096
rect 1325 2084 1331 2096
rect 1389 2064 1395 2136
rect 1613 2123 1619 2136
rect 1492 2117 1619 2123
rect 1389 2044 1395 2056
rect 1357 2003 1363 2036
rect 1549 2004 1555 2036
rect 1357 1997 1379 2003
rect 1277 1844 1283 1856
rect 1325 1824 1331 1876
rect 1373 1864 1379 1997
rect 1581 1884 1587 2096
rect 1645 2024 1651 2136
rect 1677 1924 1683 2036
rect 1629 1877 1644 1883
rect 1453 1864 1459 1876
rect 1476 1857 1484 1863
rect 1341 1823 1347 1856
rect 1405 1824 1411 1856
rect 1341 1817 1363 1823
rect 1341 1784 1347 1796
rect 1357 1784 1363 1817
rect 1469 1777 1484 1783
rect 1277 1763 1283 1776
rect 1277 1757 1292 1763
rect 1453 1744 1459 1776
rect 1469 1764 1475 1777
rect 1501 1763 1507 1796
rect 1492 1757 1507 1763
rect 1309 1464 1315 1736
rect 1469 1723 1475 1736
rect 1428 1717 1475 1723
rect 1325 1484 1331 1496
rect 1373 1464 1379 1476
rect 1293 1444 1299 1456
rect 1357 1443 1363 1456
rect 1341 1437 1363 1443
rect 1341 1343 1347 1437
rect 1389 1424 1395 1696
rect 1405 1584 1411 1636
rect 1453 1524 1459 1676
rect 1517 1604 1523 1876
rect 1533 1784 1539 1796
rect 1565 1644 1571 1856
rect 1597 1763 1603 1796
rect 1613 1784 1619 1796
rect 1597 1757 1619 1763
rect 1581 1704 1587 1716
rect 1549 1584 1555 1596
rect 1581 1564 1587 1696
rect 1453 1504 1459 1516
rect 1581 1484 1587 1536
rect 1597 1484 1603 1736
rect 1613 1724 1619 1757
rect 1629 1524 1635 1877
rect 1661 1864 1667 1916
rect 1757 1884 1763 2397
rect 1773 2324 1779 2356
rect 1789 2284 1795 2356
rect 1837 2304 1843 2496
rect 1885 2344 1891 3056
rect 1901 2984 1907 3077
rect 1965 3064 1971 3076
rect 2029 3064 2035 3076
rect 2077 3064 2083 3076
rect 1933 2944 1939 2956
rect 1917 2904 1923 2936
rect 1949 2924 1955 2996
rect 1981 2963 1987 2976
rect 1981 2957 1996 2963
rect 1901 2884 1907 2896
rect 1981 2884 1987 2957
rect 2013 2944 2019 3036
rect 2045 3004 2051 3056
rect 2061 3044 2067 3056
rect 2061 2964 2067 2976
rect 2045 2804 2051 2836
rect 1901 2724 1907 2756
rect 2013 2704 2019 2716
rect 2093 2704 2099 3296
rect 2125 3163 2131 3236
rect 2125 3157 2147 3163
rect 1917 2644 1923 2676
rect 1917 2564 1923 2596
rect 1949 2543 1955 2696
rect 1965 2664 1971 2676
rect 1997 2664 2003 2676
rect 1981 2644 1987 2656
rect 2093 2643 2099 2676
rect 2109 2664 2115 2756
rect 2125 2664 2131 2836
rect 2141 2764 2147 3157
rect 2189 3124 2195 3136
rect 2157 3084 2163 3116
rect 2189 3084 2195 3096
rect 2221 3064 2227 3296
rect 2237 3203 2243 3436
rect 2253 3404 2259 3436
rect 2285 3304 2291 3516
rect 2301 3484 2307 3516
rect 2317 3484 2323 3496
rect 2365 3484 2371 3716
rect 2429 3704 2435 3716
rect 2381 3524 2387 3636
rect 2381 3484 2387 3496
rect 2445 3484 2451 3796
rect 2461 3684 2467 3876
rect 2509 3864 2515 3936
rect 2573 3884 2579 4057
rect 2685 3964 2691 3976
rect 2653 3884 2659 3936
rect 2493 3804 2499 3836
rect 2525 3784 2531 3876
rect 2589 3844 2595 3876
rect 2637 3843 2643 3876
rect 2701 3864 2707 3936
rect 2717 3884 2723 3896
rect 2797 3864 2803 3876
rect 2829 3864 2835 3916
rect 2973 3884 2979 3896
rect 3069 3876 3070 3883
rect 2637 3837 2659 3843
rect 2557 3744 2563 3836
rect 2589 3824 2595 3836
rect 2621 3804 2627 3836
rect 2653 3804 2659 3837
rect 2589 3744 2595 3776
rect 2493 3724 2499 3736
rect 2301 3344 2307 3456
rect 2317 3364 2323 3396
rect 2429 3383 2435 3436
rect 2413 3377 2435 3383
rect 2349 3357 2387 3363
rect 2349 3343 2355 3357
rect 2381 3344 2387 3357
rect 2413 3344 2419 3377
rect 2340 3337 2355 3343
rect 2386 3337 2387 3344
rect 2301 3324 2307 3336
rect 2365 3224 2371 3236
rect 2237 3197 2259 3203
rect 2253 3124 2259 3197
rect 2429 3184 2435 3356
rect 2477 3304 2483 3696
rect 2493 3603 2499 3696
rect 2493 3597 2515 3603
rect 2509 3464 2515 3597
rect 2525 3484 2531 3676
rect 2589 3484 2595 3736
rect 2637 3564 2643 3756
rect 2653 3744 2659 3796
rect 2701 3783 2707 3856
rect 2749 3844 2755 3856
rect 2813 3804 2819 3856
rect 2701 3777 2723 3783
rect 2717 3744 2723 3777
rect 2845 3764 2851 3876
rect 2861 3744 2867 3796
rect 2877 3784 2883 3836
rect 2893 3804 2899 3856
rect 2909 3764 2915 3876
rect 2957 3844 2963 3856
rect 2973 3804 2979 3876
rect 3037 3844 3043 3876
rect 3069 3864 3075 3876
rect 3085 3864 3091 3896
rect 3197 3884 3203 3896
rect 3101 3844 3107 3876
rect 2964 3757 2972 3763
rect 2989 3743 2995 3756
rect 2980 3737 2995 3743
rect 2781 3724 2787 3736
rect 2813 3644 2819 3716
rect 3021 3704 3027 3756
rect 3037 3744 3043 3836
rect 3085 3764 3091 3836
rect 3213 3764 3219 3856
rect 3101 3744 3107 3756
rect 2692 3637 2700 3643
rect 2653 3524 2659 3596
rect 2749 3543 2755 3636
rect 2765 3584 2771 3596
rect 2749 3537 2771 3543
rect 2493 3424 2499 3436
rect 2509 3403 2515 3456
rect 2493 3397 2515 3403
rect 2493 3344 2499 3397
rect 2637 3384 2643 3476
rect 2701 3444 2707 3456
rect 2621 3364 2627 3376
rect 2685 3344 2691 3436
rect 2717 3404 2723 3476
rect 2765 3464 2771 3537
rect 2813 3524 2819 3636
rect 2829 3504 2835 3636
rect 2829 3363 2835 3376
rect 2820 3357 2835 3363
rect 2701 3344 2707 3356
rect 2845 3344 2851 3476
rect 2925 3444 2931 3476
rect 2941 3464 2947 3536
rect 2973 3484 2979 3556
rect 3005 3524 3011 3636
rect 3037 3484 3043 3556
rect 3028 3457 3036 3463
rect 2877 3424 2883 3436
rect 2973 3384 2979 3456
rect 2973 3363 2979 3376
rect 2964 3357 2979 3363
rect 2925 3344 2931 3356
rect 2804 3337 2812 3343
rect 2621 3324 2627 3336
rect 2516 3237 2531 3243
rect 2525 3143 2531 3237
rect 2525 3137 2547 3143
rect 2541 3124 2547 3137
rect 2260 3077 2275 3083
rect 2173 3004 2179 3056
rect 2189 2984 2195 3036
rect 2237 2984 2243 3036
rect 2253 2984 2259 2996
rect 2173 2964 2179 2976
rect 2269 2944 2275 3077
rect 2317 3044 2323 3056
rect 2301 2984 2307 3036
rect 2333 2984 2339 3076
rect 2365 2964 2371 2996
rect 2397 2964 2403 3116
rect 2445 3104 2451 3116
rect 2557 3084 2563 3096
rect 2605 3064 2611 3076
rect 2621 3064 2627 3096
rect 2685 3064 2691 3076
rect 2509 3044 2515 3056
rect 2429 3004 2435 3036
rect 2493 2963 2499 3036
rect 2573 2983 2579 3036
rect 2637 3024 2643 3036
rect 2573 2977 2595 2983
rect 2493 2957 2508 2963
rect 2276 2937 2284 2943
rect 2157 2884 2163 2936
rect 2157 2864 2163 2876
rect 2205 2724 2211 2936
rect 2301 2904 2307 2956
rect 2349 2944 2355 2956
rect 2445 2944 2451 2956
rect 2589 2944 2595 2977
rect 2372 2937 2380 2943
rect 2493 2937 2508 2943
rect 2404 2897 2419 2903
rect 2221 2703 2227 2896
rect 2253 2784 2259 2876
rect 2333 2724 2339 2736
rect 2205 2697 2227 2703
rect 2141 2644 2147 2676
rect 2189 2664 2195 2676
rect 2093 2637 2115 2643
rect 2045 2584 2051 2636
rect 2061 2563 2067 2636
rect 2109 2584 2115 2637
rect 2173 2583 2179 2636
rect 2157 2577 2179 2583
rect 2052 2557 2067 2563
rect 2157 2544 2163 2577
rect 1949 2537 1964 2543
rect 2068 2537 2076 2543
rect 2029 2444 2035 2536
rect 2077 2504 2083 2516
rect 1917 2364 1923 2376
rect 1933 2344 1939 2436
rect 2125 2404 2131 2436
rect 1885 2324 1891 2336
rect 1789 2144 1795 2276
rect 1805 2264 1811 2276
rect 1821 2243 1827 2276
rect 1805 2237 1827 2243
rect 1805 2184 1811 2237
rect 1837 2144 1843 2176
rect 1869 2163 1875 2176
rect 1860 2157 1875 2163
rect 1789 2124 1795 2136
rect 1773 2084 1779 2096
rect 1869 1984 1875 2016
rect 1821 1884 1827 1936
rect 1805 1864 1811 1876
rect 1677 1784 1683 1856
rect 1789 1824 1795 1836
rect 1741 1784 1747 1796
rect 1661 1744 1667 1776
rect 1789 1764 1795 1776
rect 1709 1757 1724 1763
rect 1709 1724 1715 1757
rect 1796 1737 1811 1743
rect 1725 1724 1731 1736
rect 1805 1724 1811 1737
rect 1837 1704 1843 1956
rect 1885 1864 1891 2316
rect 1949 2284 1955 2336
rect 1933 2244 1939 2256
rect 1917 2144 1923 2156
rect 1949 2143 1955 2256
rect 1940 2137 1955 2143
rect 1853 1744 1859 1776
rect 1869 1724 1875 1736
rect 1837 1684 1843 1696
rect 1677 1584 1683 1596
rect 1629 1484 1635 1496
rect 1620 1457 1635 1463
rect 1533 1424 1539 1456
rect 1597 1424 1603 1456
rect 1629 1424 1635 1457
rect 1725 1424 1731 1456
rect 1357 1364 1363 1396
rect 1421 1364 1427 1376
rect 1485 1364 1491 1376
rect 1341 1337 1363 1343
rect 1133 1217 1155 1223
rect 1149 1184 1155 1217
rect 1277 1144 1283 1236
rect 1309 1164 1315 1296
rect 1341 1264 1347 1276
rect 1357 1223 1363 1337
rect 1380 1337 1388 1343
rect 1444 1337 1484 1343
rect 1517 1343 1523 1376
rect 1549 1364 1555 1396
rect 1613 1344 1619 1356
rect 1508 1337 1523 1343
rect 1533 1337 1548 1343
rect 1533 1323 1539 1337
rect 1629 1323 1635 1416
rect 1789 1404 1795 1456
rect 1805 1424 1811 1516
rect 1837 1484 1843 1636
rect 1869 1524 1875 1716
rect 1885 1704 1891 1716
rect 1885 1664 1891 1696
rect 1901 1604 1907 1876
rect 1949 1784 1955 2096
rect 1965 1924 1971 2376
rect 2125 2364 2131 2376
rect 2029 2244 2035 2316
rect 2077 2284 2083 2356
rect 2189 2324 2195 2336
rect 2052 2277 2060 2283
rect 2141 2277 2156 2283
rect 2141 2263 2147 2277
rect 2189 2264 2195 2276
rect 2109 2257 2147 2263
rect 2157 2257 2172 2263
rect 2061 2244 2067 2256
rect 2109 2244 2115 2257
rect 2157 2244 2163 2257
rect 1988 2237 1996 2243
rect 1997 2124 2003 2156
rect 2013 2124 2019 2136
rect 1965 1884 1971 1916
rect 1981 1864 1987 1876
rect 1981 1804 1987 1856
rect 1917 1763 1923 1776
rect 1917 1757 1932 1763
rect 1997 1704 2003 1736
rect 2029 1724 2035 2236
rect 2173 2184 2179 2236
rect 2061 2144 2067 2156
rect 2045 1964 2051 2036
rect 2077 1924 2083 2096
rect 2141 1964 2147 2096
rect 2189 1964 2195 2036
rect 2093 1897 2188 1903
rect 2093 1883 2099 1897
rect 2084 1877 2099 1883
rect 2045 1844 2051 1856
rect 2061 1824 2067 1856
rect 2141 1824 2147 1876
rect 2061 1764 2067 1796
rect 2173 1783 2179 1836
rect 2205 1823 2211 2697
rect 2285 2604 2291 2676
rect 2365 2657 2380 2663
rect 2301 2584 2307 2656
rect 2365 2644 2371 2657
rect 2317 2584 2323 2596
rect 2413 2583 2419 2897
rect 2445 2804 2451 2936
rect 2493 2924 2499 2937
rect 2637 2924 2643 2936
rect 2717 2924 2723 3336
rect 3037 3324 3043 3336
rect 2733 3104 2739 3116
rect 2845 3084 2851 3276
rect 2861 3264 2867 3296
rect 2877 3284 2883 3316
rect 2893 3164 2899 3236
rect 3005 3203 3011 3236
rect 2989 3197 3011 3203
rect 2893 3124 2899 3136
rect 2973 3124 2979 3136
rect 2733 3077 2748 3083
rect 2733 3044 2739 3077
rect 2749 2964 2755 3056
rect 2749 2904 2755 2956
rect 2461 2884 2467 2896
rect 2621 2804 2627 2836
rect 2653 2764 2659 2896
rect 2653 2724 2659 2736
rect 2468 2717 2476 2723
rect 2781 2704 2787 3076
rect 2829 3024 2835 3056
rect 2813 2904 2819 2916
rect 2797 2884 2803 2896
rect 2829 2744 2835 2836
rect 2845 2804 2851 3076
rect 2861 2944 2867 3016
rect 2957 2984 2963 3076
rect 2884 2957 2892 2963
rect 2925 2924 2931 2936
rect 2941 2764 2947 2956
rect 2957 2824 2963 2836
rect 2925 2724 2931 2736
rect 2941 2704 2947 2716
rect 2445 2684 2451 2696
rect 2493 2684 2499 2696
rect 2788 2677 2803 2683
rect 2733 2664 2739 2676
rect 2765 2664 2771 2676
rect 2797 2664 2803 2677
rect 2557 2657 2572 2663
rect 2509 2604 2515 2656
rect 2557 2644 2563 2657
rect 2557 2584 2563 2596
rect 2413 2577 2435 2583
rect 2253 2564 2259 2576
rect 2429 2564 2435 2577
rect 2621 2564 2627 2636
rect 2685 2583 2691 2636
rect 2669 2577 2691 2583
rect 2237 2544 2243 2556
rect 2253 2504 2259 2536
rect 2269 2444 2275 2536
rect 2317 2384 2323 2436
rect 2237 2257 2252 2263
rect 2237 2244 2243 2257
rect 2269 2244 2275 2276
rect 2253 2163 2259 2176
rect 2301 2164 2307 2176
rect 2244 2157 2259 2163
rect 2228 2137 2236 2143
rect 2276 2137 2284 2143
rect 2317 2124 2323 2136
rect 2333 2104 2339 2556
rect 2349 2244 2355 2276
rect 2365 2184 2371 2196
rect 2397 2103 2403 2536
rect 2413 2524 2419 2536
rect 2429 2524 2435 2556
rect 2445 2283 2451 2296
rect 2436 2277 2451 2283
rect 2429 2184 2435 2256
rect 2461 2164 2467 2496
rect 2477 2324 2483 2556
rect 2509 2544 2515 2556
rect 2669 2544 2675 2577
rect 2701 2564 2707 2636
rect 2717 2524 2723 2536
rect 2589 2284 2595 2296
rect 2637 2284 2643 2296
rect 2493 2244 2499 2276
rect 2516 2237 2524 2243
rect 2493 2184 2499 2216
rect 2541 2204 2547 2276
rect 2573 2264 2579 2276
rect 2557 2224 2563 2256
rect 2525 2144 2531 2196
rect 2573 2144 2579 2156
rect 2429 2124 2435 2136
rect 2589 2124 2595 2136
rect 2605 2124 2611 2156
rect 2397 2097 2412 2103
rect 2221 1884 2227 1976
rect 2253 1884 2259 1996
rect 2269 1844 2275 1916
rect 2317 1844 2323 1856
rect 2292 1837 2300 1843
rect 2189 1817 2211 1823
rect 2189 1784 2195 1817
rect 2253 1784 2259 1796
rect 2157 1777 2179 1783
rect 2157 1744 2163 1777
rect 2189 1764 2195 1776
rect 2045 1724 2051 1736
rect 2077 1724 2083 1736
rect 2013 1684 2019 1696
rect 1917 1584 1923 1616
rect 1933 1584 1939 1596
rect 1853 1503 1859 1516
rect 1853 1497 1884 1503
rect 1876 1477 1884 1483
rect 1773 1383 1779 1396
rect 1773 1377 1795 1383
rect 1789 1364 1795 1377
rect 1805 1364 1811 1376
rect 1677 1344 1683 1356
rect 1709 1344 1715 1356
rect 1682 1337 1683 1344
rect 1476 1317 1539 1323
rect 1613 1317 1635 1323
rect 1341 1217 1363 1223
rect 1341 1184 1347 1217
rect 1405 1144 1411 1236
rect 1261 1124 1267 1136
rect 1396 1117 1404 1123
rect 1421 1103 1427 1156
rect 1405 1097 1427 1103
rect 1405 1084 1411 1097
rect 1284 1077 1292 1083
rect 1316 1077 1324 1083
rect 1101 1044 1107 1076
rect 1421 1064 1427 1076
rect 1293 1044 1299 1056
rect 1021 1004 1027 1036
rect 1037 983 1043 1036
rect 1037 977 1059 983
rect 916 957 931 963
rect 1005 957 1020 963
rect 925 944 931 957
rect 1053 944 1059 977
rect 1133 944 1139 1016
rect 1149 964 1155 1036
rect 1165 1024 1171 1036
rect 1357 1003 1363 1036
rect 1341 997 1363 1003
rect 1341 964 1347 997
rect 1197 957 1212 963
rect 893 937 908 943
rect 989 923 995 936
rect 1021 923 1027 936
rect 989 917 1027 923
rect 900 877 908 883
rect 1197 864 1203 957
rect 1389 944 1395 1016
rect 1405 964 1411 996
rect 893 784 899 856
rect 973 824 979 836
rect 1085 824 1091 836
rect 1101 803 1107 836
rect 1085 797 1107 803
rect 781 737 803 743
rect 605 677 620 683
rect 509 604 515 636
rect 525 583 531 676
rect 573 603 579 636
rect 605 604 611 677
rect 637 664 643 716
rect 701 684 707 696
rect 781 684 787 737
rect 804 717 812 723
rect 717 664 723 676
rect 829 657 844 663
rect 829 644 835 657
rect 772 637 787 643
rect 653 604 659 636
rect 509 577 531 583
rect 557 597 579 603
rect 509 544 515 577
rect 557 563 563 597
rect 532 557 563 563
rect 669 544 675 596
rect 765 584 771 616
rect 781 564 787 637
rect 861 624 867 676
rect 877 584 883 776
rect 957 664 963 676
rect 893 544 899 616
rect 909 584 915 616
rect 973 564 979 636
rect 957 544 963 556
rect 989 544 995 576
rect 1037 564 1043 716
rect 1069 624 1075 676
rect 1085 664 1091 797
rect 1133 724 1139 836
rect 1213 804 1219 936
rect 1261 924 1267 936
rect 1325 884 1331 936
rect 1229 824 1235 836
rect 1181 724 1187 756
rect 1261 724 1267 796
rect 1341 784 1347 876
rect 1357 824 1363 836
rect 1405 724 1411 936
rect 1421 724 1427 836
rect 1140 677 1148 683
rect 1172 677 1180 683
rect 1213 624 1219 636
rect 1229 584 1235 716
rect 1277 684 1283 716
rect 1101 564 1107 576
rect 1165 544 1171 556
rect 1277 544 1283 656
rect 1293 584 1299 656
rect 1309 644 1315 676
rect 1357 603 1363 636
rect 1341 597 1363 603
rect 1341 564 1347 597
rect 1357 564 1363 576
rect 1373 544 1379 616
rect 1124 537 1132 543
rect 173 284 179 296
rect 189 264 195 496
rect 285 484 291 496
rect 301 324 307 496
rect 365 324 371 476
rect 381 364 387 436
rect 61 257 76 263
rect 61 244 67 257
rect 205 244 211 256
rect 20 177 28 183
rect 61 164 67 176
rect 77 164 83 176
rect 253 164 259 176
rect 269 164 275 236
rect 333 204 339 236
rect 237 144 243 156
rect 285 144 291 156
rect 349 144 355 196
rect 365 164 371 316
rect 381 284 387 316
rect 429 284 435 396
rect 445 283 451 436
rect 493 343 499 496
rect 477 337 499 343
rect 477 284 483 337
rect 509 284 515 536
rect 541 524 547 536
rect 605 524 611 536
rect 797 524 803 536
rect 941 504 947 516
rect 1325 504 1331 536
rect 580 337 588 343
rect 701 303 707 436
rect 717 344 723 356
rect 685 297 707 303
rect 445 277 467 283
rect 445 244 451 256
rect 461 244 467 277
rect 685 263 691 297
rect 733 264 739 496
rect 685 257 700 263
rect 397 164 403 236
rect 525 204 531 236
rect 509 164 515 176
rect 429 157 483 163
rect 93 124 99 136
rect 189 124 195 136
rect 365 124 371 156
rect 429 124 435 157
rect 477 143 483 157
rect 557 144 563 196
rect 573 164 579 176
rect 701 164 707 216
rect 749 204 755 276
rect 781 263 787 356
rect 829 284 835 436
rect 1085 424 1091 436
rect 909 297 1036 303
rect 804 277 812 283
rect 893 264 899 276
rect 909 264 915 297
rect 1069 284 1075 316
rect 772 257 787 263
rect 836 257 851 263
rect 845 244 851 257
rect 925 244 931 276
rect 1085 264 1091 396
rect 1149 344 1155 436
rect 1197 324 1203 336
rect 1261 324 1267 496
rect 1101 284 1107 296
rect 1149 264 1155 316
rect 1165 284 1171 296
rect 1325 284 1331 336
rect 1220 277 1228 283
rect 1373 283 1379 316
rect 1389 284 1395 696
rect 1421 664 1427 676
rect 1453 644 1459 1196
rect 1501 1044 1507 1076
rect 1469 1023 1475 1036
rect 1469 1017 1491 1023
rect 1469 964 1475 996
rect 1485 964 1491 1017
rect 1533 1004 1539 1236
rect 1613 1223 1619 1317
rect 1725 1304 1731 1356
rect 1837 1343 1843 1476
rect 1853 1364 1859 1456
rect 1837 1337 1852 1343
rect 1629 1284 1635 1296
rect 1773 1264 1779 1336
rect 1853 1324 1859 1336
rect 1885 1324 1891 1476
rect 1901 1464 1907 1516
rect 1981 1464 1987 1636
rect 2029 1484 2035 1556
rect 2093 1543 2099 1696
rect 2173 1544 2179 1756
rect 2237 1744 2243 1756
rect 2285 1743 2291 1796
rect 2301 1764 2307 1776
rect 2308 1757 2316 1763
rect 2333 1763 2339 2096
rect 2349 1864 2355 1876
rect 2372 1857 2387 1863
rect 2381 1844 2387 1857
rect 2413 1764 2419 1916
rect 2429 1784 2435 1876
rect 2493 1844 2499 1856
rect 2333 1757 2355 1763
rect 2285 1737 2316 1743
rect 2093 1537 2115 1543
rect 2045 1464 2051 1536
rect 1901 1343 1907 1456
rect 1981 1383 1987 1456
rect 1997 1404 2003 1436
rect 2093 1424 2099 1516
rect 2109 1484 2115 1537
rect 2221 1524 2227 1616
rect 2173 1497 2211 1503
rect 2173 1483 2179 1497
rect 2205 1484 2211 1497
rect 2237 1484 2243 1496
rect 2285 1484 2291 1516
rect 2301 1484 2307 1696
rect 2349 1484 2355 1757
rect 2381 1744 2387 1756
rect 2445 1724 2451 1736
rect 2420 1717 2428 1723
rect 2397 1704 2403 1716
rect 2365 1624 2371 1636
rect 2397 1503 2403 1696
rect 2445 1684 2451 1696
rect 2445 1604 2451 1676
rect 2397 1497 2419 1503
rect 2148 1477 2179 1483
rect 2125 1424 2131 1456
rect 2189 1444 2195 1476
rect 2317 1464 2323 1476
rect 2301 1443 2307 1456
rect 2381 1444 2387 1456
rect 2301 1437 2323 1443
rect 1965 1377 1987 1383
rect 1965 1344 1971 1377
rect 1997 1363 2003 1376
rect 2061 1364 2067 1376
rect 2125 1364 2131 1396
rect 2189 1364 2195 1436
rect 1988 1357 2003 1363
rect 2077 1344 2083 1356
rect 2141 1344 2147 1356
rect 2253 1344 2259 1416
rect 2301 1384 2307 1396
rect 2317 1384 2323 1437
rect 2365 1383 2371 1436
rect 2365 1377 2387 1383
rect 1901 1337 1916 1343
rect 1597 1217 1619 1223
rect 1597 1184 1603 1217
rect 1741 1124 1747 1236
rect 1837 1144 1843 1296
rect 1853 1204 1859 1316
rect 1892 1297 1900 1303
rect 1949 1143 1955 1336
rect 1933 1137 1955 1143
rect 1764 1117 1772 1123
rect 1821 1097 1859 1103
rect 1549 984 1555 1036
rect 1533 944 1539 956
rect 1533 937 1534 944
rect 1485 924 1491 936
rect 1501 864 1507 936
rect 1565 884 1571 1076
rect 1581 804 1587 896
rect 1613 764 1619 836
rect 1581 724 1587 756
rect 1549 683 1555 696
rect 1629 684 1635 1056
rect 1709 1044 1715 1076
rect 1741 1064 1747 1076
rect 1821 1063 1827 1097
rect 1853 1083 1859 1097
rect 1933 1084 1939 1137
rect 1853 1077 1875 1083
rect 1789 1057 1827 1063
rect 1725 984 1731 1056
rect 1789 1044 1795 1057
rect 1748 957 1756 963
rect 1645 904 1651 936
rect 1661 904 1667 956
rect 1693 904 1699 936
rect 1805 924 1811 956
rect 1821 944 1827 1036
rect 1837 1024 1843 1076
rect 1869 1064 1875 1077
rect 1981 1083 1987 1116
rect 1949 1077 1987 1083
rect 1901 1064 1907 1076
rect 1853 1024 1859 1056
rect 1917 1044 1923 1056
rect 1949 1044 1955 1077
rect 1997 1064 2003 1156
rect 2077 1124 2083 1336
rect 2093 1104 2099 1116
rect 2109 1084 2115 1116
rect 2125 1084 2131 1316
rect 2020 1077 2035 1083
rect 2029 1063 2035 1077
rect 2109 1064 2115 1076
rect 2189 1064 2195 1336
rect 2221 1124 2227 1236
rect 2253 1203 2259 1336
rect 2349 1304 2355 1336
rect 2365 1284 2371 1356
rect 2381 1304 2387 1377
rect 2237 1197 2259 1203
rect 2237 1084 2243 1197
rect 2381 1184 2387 1196
rect 2397 1104 2403 1476
rect 2413 1304 2419 1497
rect 2477 1463 2483 1516
rect 2509 1503 2515 1636
rect 2525 1524 2531 1936
rect 2541 1864 2547 1876
rect 2557 1864 2563 2036
rect 2573 1884 2579 1896
rect 2557 1764 2563 1796
rect 2541 1724 2547 1736
rect 2589 1644 2595 1916
rect 2605 1784 2611 2116
rect 2653 2104 2659 2116
rect 2621 1877 2636 1883
rect 2621 1864 2627 1877
rect 2621 1744 2627 1856
rect 2637 1764 2643 1816
rect 2637 1744 2643 1756
rect 2605 1684 2611 1696
rect 2621 1504 2627 1736
rect 2493 1497 2515 1503
rect 2493 1484 2499 1497
rect 2605 1484 2611 1496
rect 2477 1457 2492 1463
rect 2628 1457 2643 1463
rect 2637 1444 2643 1457
rect 2445 1364 2451 1396
rect 2509 1344 2515 1356
rect 2445 1204 2451 1336
rect 2461 1304 2467 1336
rect 2525 1324 2531 1336
rect 2509 1184 2515 1296
rect 2541 1204 2547 1336
rect 2589 1304 2595 1356
rect 2653 1323 2659 1696
rect 2669 1524 2675 2316
rect 2717 2304 2723 2316
rect 2685 2143 2691 2236
rect 2685 2137 2700 2143
rect 2685 2104 2691 2116
rect 2733 2024 2739 2656
rect 2765 2264 2771 2276
rect 2749 2204 2755 2236
rect 2765 2224 2771 2256
rect 2765 1984 2771 2036
rect 2781 1984 2787 2136
rect 2685 1784 2691 1916
rect 2701 1804 2707 1836
rect 2701 1704 2707 1736
rect 2717 1704 2723 1736
rect 2797 1724 2803 2656
rect 2877 2503 2883 2636
rect 2941 2584 2947 2596
rect 2957 2564 2963 2636
rect 2893 2544 2899 2556
rect 2973 2523 2979 3056
rect 2989 3024 2995 3197
rect 3021 3084 3027 3116
rect 3037 3104 3043 3116
rect 3053 2963 3059 3736
rect 3133 3624 3139 3636
rect 3149 3584 3155 3756
rect 3165 3744 3171 3756
rect 3229 3724 3235 3876
rect 3277 3864 3283 3916
rect 3293 3884 3299 3956
rect 3613 3924 3619 3936
rect 4061 3924 4067 3936
rect 4253 3924 4259 3936
rect 3828 3917 3836 3923
rect 3469 3884 3475 3916
rect 3597 3884 3603 3916
rect 3732 3897 3740 3903
rect 3421 3864 3427 3876
rect 3469 3864 3475 3876
rect 3405 3844 3411 3856
rect 3261 3764 3267 3796
rect 3357 3743 3363 3756
rect 3373 3744 3379 3816
rect 3332 3737 3363 3743
rect 3197 3623 3203 3636
rect 3197 3617 3219 3623
rect 3117 3484 3123 3516
rect 3149 3504 3155 3536
rect 3117 3364 3123 3476
rect 3165 3463 3171 3516
rect 3213 3484 3219 3617
rect 3245 3584 3251 3736
rect 3325 3684 3331 3696
rect 3229 3484 3235 3536
rect 3277 3524 3283 3636
rect 3341 3584 3347 3636
rect 3389 3604 3395 3756
rect 3437 3744 3443 3816
rect 3453 3764 3459 3796
rect 3469 3764 3475 3776
rect 3405 3483 3411 3636
rect 3421 3484 3427 3696
rect 3485 3544 3491 3876
rect 3645 3764 3651 3776
rect 3629 3744 3635 3756
rect 3661 3744 3667 3836
rect 3565 3724 3571 3736
rect 3469 3504 3475 3536
rect 3549 3524 3555 3596
rect 3661 3524 3667 3576
rect 3533 3484 3539 3516
rect 3389 3477 3411 3483
rect 3149 3457 3171 3463
rect 3149 3384 3155 3457
rect 3197 3424 3203 3436
rect 3213 3403 3219 3456
rect 3277 3424 3283 3476
rect 3213 3397 3235 3403
rect 3213 3364 3219 3376
rect 3229 3344 3235 3397
rect 3133 3337 3134 3343
rect 3142 3337 3196 3343
rect 3229 3324 3235 3336
rect 3277 3264 3283 3356
rect 3293 3344 3299 3356
rect 3325 3344 3331 3436
rect 3341 3424 3347 3456
rect 3357 3424 3363 3476
rect 3389 3384 3395 3477
rect 3405 3444 3411 3456
rect 3341 3364 3347 3376
rect 3421 3364 3427 3476
rect 3469 3364 3475 3376
rect 3501 3344 3507 3396
rect 3533 3384 3539 3416
rect 3517 3364 3523 3376
rect 3581 3364 3587 3436
rect 3597 3424 3603 3476
rect 3613 3404 3619 3516
rect 3693 3484 3699 3876
rect 3709 3864 3715 3896
rect 3757 3884 3763 3896
rect 3789 3884 3795 3896
rect 4173 3884 4179 3916
rect 4237 3904 4243 3916
rect 3876 3877 3884 3883
rect 3997 3864 4003 3876
rect 4109 3864 4115 3876
rect 3773 3804 3779 3856
rect 3789 3764 3795 3816
rect 3757 3744 3763 3756
rect 3709 3604 3715 3636
rect 3757 3524 3763 3736
rect 3773 3704 3779 3756
rect 3805 3744 3811 3836
rect 3901 3824 3907 3856
rect 3917 3764 3923 3856
rect 3853 3744 3859 3756
rect 3981 3744 3987 3856
rect 3844 3717 3916 3723
rect 3997 3683 4003 3856
rect 4093 3804 4099 3836
rect 4029 3744 4035 3796
rect 4109 3784 4115 3856
rect 4125 3824 4131 3876
rect 4301 3864 4307 3956
rect 4397 3924 4403 3936
rect 4708 3917 4716 3923
rect 4461 3884 4467 3896
rect 4317 3864 4323 3876
rect 4157 3784 4163 3796
rect 4173 3764 4179 3816
rect 4221 3804 4227 3836
rect 4052 3757 4147 3763
rect 4045 3724 4051 3736
rect 3997 3677 4019 3683
rect 3965 3664 3971 3676
rect 3821 3524 3827 3596
rect 3645 3364 3651 3436
rect 3693 3344 3699 3476
rect 3725 3464 3731 3476
rect 3741 3464 3747 3476
rect 3709 3383 3715 3436
rect 3709 3377 3731 3383
rect 3725 3364 3731 3377
rect 3757 3344 3763 3516
rect 3780 3497 3916 3503
rect 3981 3483 3987 3636
rect 3965 3477 3987 3483
rect 3069 3204 3075 3236
rect 3117 3104 3123 3116
rect 3133 3084 3139 3116
rect 3085 3023 3091 3036
rect 3085 3017 3107 3023
rect 3085 2984 3091 2996
rect 3053 2957 3068 2963
rect 2989 2924 2995 2936
rect 3053 2884 3059 2936
rect 2989 2604 2995 2716
rect 3021 2683 3027 2736
rect 3012 2677 3027 2683
rect 3053 2644 3059 2676
rect 3069 2664 3075 2776
rect 3101 2744 3107 3017
rect 3181 3004 3187 3116
rect 3197 3084 3203 3116
rect 3261 3104 3267 3116
rect 3293 3104 3299 3336
rect 3309 3124 3315 3336
rect 3501 3324 3507 3336
rect 3581 3324 3587 3336
rect 3309 3084 3315 3116
rect 3325 3083 3331 3176
rect 3421 3084 3427 3096
rect 3325 3077 3347 3083
rect 3149 2964 3155 2976
rect 3213 2964 3219 2996
rect 3261 2984 3267 2996
rect 3277 2984 3283 3056
rect 3325 3044 3331 3056
rect 3341 3023 3347 3077
rect 3357 3077 3372 3083
rect 3357 3064 3363 3077
rect 3380 3057 3388 3063
rect 3325 3017 3347 3023
rect 3165 2924 3171 2936
rect 3229 2904 3235 2936
rect 3204 2897 3212 2903
rect 3309 2864 3315 2896
rect 3325 2824 3331 3017
rect 3341 2964 3347 2996
rect 3357 2944 3363 3016
rect 3405 2984 3411 3056
rect 3341 2904 3347 2936
rect 3085 2684 3091 2696
rect 3165 2684 3171 2696
rect 3325 2684 3331 2796
rect 3341 2724 3347 2896
rect 3405 2844 3411 2856
rect 3421 2824 3427 3076
rect 3437 2944 3443 3316
rect 3453 3184 3459 3236
rect 3565 3204 3571 3296
rect 3501 3084 3507 3096
rect 3533 3084 3539 3136
rect 3597 3084 3603 3236
rect 3677 3084 3683 3096
rect 3517 3044 3523 3056
rect 3597 3004 3603 3076
rect 3661 3024 3667 3056
rect 3693 3044 3699 3336
rect 3741 3184 3747 3336
rect 3757 3083 3763 3336
rect 3789 3224 3795 3436
rect 3837 3384 3843 3476
rect 3789 3084 3795 3136
rect 3748 3077 3763 3083
rect 3709 3004 3715 3036
rect 3453 2964 3459 2976
rect 3437 2924 3443 2936
rect 3469 2904 3475 2936
rect 3501 2924 3507 2976
rect 3581 2964 3587 2976
rect 3716 2957 3724 2963
rect 3565 2944 3571 2956
rect 3693 2924 3699 2936
rect 3725 2924 3731 2936
rect 3540 2897 3548 2903
rect 3517 2784 3523 2836
rect 3661 2824 3667 2896
rect 3741 2864 3747 2896
rect 3693 2724 3699 2816
rect 3476 2697 3523 2703
rect 3517 2684 3523 2697
rect 3300 2677 3308 2683
rect 3325 2664 3331 2676
rect 3005 2564 3011 2576
rect 2989 2544 2995 2556
rect 3021 2544 3027 2556
rect 2973 2517 2995 2523
rect 2852 2497 2867 2503
rect 2877 2497 2892 2503
rect 2845 2324 2851 2336
rect 2813 2244 2819 2256
rect 2829 2164 2835 2276
rect 2861 2203 2867 2497
rect 2989 2264 2995 2517
rect 3037 2484 3043 2496
rect 3069 2483 3075 2656
rect 3133 2624 3139 2636
rect 3101 2544 3107 2576
rect 3149 2544 3155 2656
rect 3261 2603 3267 2636
rect 3261 2597 3283 2603
rect 3069 2477 3091 2483
rect 3085 2324 3091 2477
rect 3181 2464 3187 2496
rect 3140 2437 3148 2443
rect 3197 2364 3203 2536
rect 3213 2464 3219 2536
rect 3229 2504 3235 2576
rect 3277 2544 3283 2597
rect 3341 2584 3347 2676
rect 3405 2644 3411 2676
rect 3517 2644 3523 2656
rect 3357 2543 3363 2616
rect 3389 2603 3395 2636
rect 3581 2624 3587 2636
rect 3389 2597 3411 2603
rect 3348 2537 3363 2543
rect 3261 2524 3267 2536
rect 3277 2504 3283 2536
rect 3405 2504 3411 2597
rect 3517 2564 3523 2576
rect 3533 2544 3539 2616
rect 3581 2584 3587 2596
rect 3597 2584 3603 2596
rect 3293 2464 3299 2496
rect 3373 2477 3388 2483
rect 3213 2384 3219 2396
rect 3373 2344 3379 2477
rect 3197 2284 3203 2296
rect 3117 2264 3123 2276
rect 3140 2257 3155 2263
rect 2877 2224 2883 2236
rect 2861 2197 2883 2203
rect 2877 2184 2883 2197
rect 2893 2164 2899 2176
rect 2925 2104 2931 2116
rect 2845 1944 2851 2096
rect 2941 2044 2947 2116
rect 2973 2104 2979 2256
rect 3149 2244 3155 2257
rect 3005 2184 3011 2236
rect 3021 2164 3027 2176
rect 3085 2144 3091 2156
rect 3156 2137 3171 2143
rect 3005 2124 3011 2136
rect 3165 2104 3171 2137
rect 3245 2124 3251 2276
rect 3261 2244 3267 2256
rect 3293 2204 3299 2316
rect 3389 2304 3395 2456
rect 3613 2344 3619 2696
rect 3757 2684 3763 3077
rect 3837 3024 3843 3036
rect 3837 2944 3843 2996
rect 3853 2824 3859 2836
rect 3869 2804 3875 3476
rect 3885 3464 3891 3476
rect 3885 3344 3891 3456
rect 3901 3364 3907 3396
rect 3965 3344 3971 3477
rect 3997 3464 4003 3476
rect 4013 3464 4019 3677
rect 4029 3524 4035 3536
rect 4045 3504 4051 3716
rect 4061 3524 4067 3757
rect 4141 3684 4147 3757
rect 4109 3504 4115 3516
rect 4173 3484 4179 3736
rect 4237 3584 4243 3756
rect 4285 3743 4291 3836
rect 4301 3824 4307 3856
rect 4285 3737 4307 3743
rect 4301 3723 4307 3737
rect 4333 3723 4339 3756
rect 4301 3717 4339 3723
rect 4365 3704 4371 3836
rect 4413 3784 4419 3816
rect 4461 3764 4467 3876
rect 4477 3844 4483 3856
rect 4525 3824 4531 3916
rect 4557 3884 4563 3896
rect 4541 3863 4547 3876
rect 4541 3857 4563 3863
rect 4477 3784 4483 3796
rect 4557 3783 4563 3857
rect 4573 3804 4579 3916
rect 4621 3884 4627 3916
rect 4733 3884 4739 3916
rect 4765 3904 4771 3956
rect 4765 3883 4771 3896
rect 4957 3884 4963 3936
rect 4765 3877 4787 3883
rect 4749 3864 4755 3876
rect 4669 3804 4675 3836
rect 4557 3777 4595 3783
rect 4589 3763 4595 3777
rect 4669 3763 4675 3776
rect 4749 3764 4755 3776
rect 4541 3757 4579 3763
rect 4589 3757 4675 3763
rect 4429 3744 4435 3756
rect 4445 3743 4451 3756
rect 4445 3737 4492 3743
rect 4541 3743 4547 3757
rect 4525 3737 4547 3743
rect 4573 3743 4579 3757
rect 4717 3744 4723 3756
rect 4733 3744 4739 3756
rect 4765 3744 4771 3856
rect 4573 3737 4707 3743
rect 4292 3697 4300 3703
rect 4525 3703 4531 3737
rect 4621 3704 4627 3716
rect 4701 3704 4707 3737
rect 4749 3724 4755 3736
rect 4516 3697 4531 3703
rect 4365 3484 4371 3676
rect 4381 3564 4387 3696
rect 4381 3524 4387 3536
rect 4061 3464 4067 3476
rect 4189 3464 4195 3476
rect 4237 3464 4243 3476
rect 3981 3424 3987 3456
rect 4045 3424 4051 3456
rect 3997 3337 4042 3343
rect 3885 3264 3891 3336
rect 3997 3324 4003 3337
rect 4050 3337 4051 3343
rect 3949 3184 3955 3296
rect 4029 3203 4035 3236
rect 4013 3197 4035 3203
rect 4013 3123 4019 3197
rect 4061 3144 4067 3456
rect 4093 3304 4099 3356
rect 4109 3124 4115 3396
rect 4125 3264 4131 3336
rect 4157 3204 4163 3436
rect 4173 3364 4179 3396
rect 4237 3384 4243 3416
rect 4285 3344 4291 3396
rect 4301 3384 4307 3476
rect 4365 3464 4371 3476
rect 4349 3404 4355 3436
rect 4397 3344 4403 3456
rect 4445 3384 4451 3696
rect 4493 3584 4499 3596
rect 4525 3524 4531 3636
rect 4557 3584 4563 3696
rect 4781 3664 4787 3877
rect 4813 3784 4819 3876
rect 4861 3857 4876 3863
rect 4861 3844 4867 3857
rect 4813 3724 4819 3756
rect 4605 3524 4611 3636
rect 4717 3524 4723 3536
rect 4541 3517 4588 3523
rect 4461 3484 4467 3516
rect 4509 3503 4515 3516
rect 4541 3503 4547 3517
rect 4749 3504 4755 3516
rect 4509 3497 4547 3503
rect 4477 3444 4483 3456
rect 4541 3423 4547 3476
rect 4541 3417 4563 3423
rect 4541 3384 4547 3396
rect 4557 3384 4563 3417
rect 4429 3364 4435 3376
rect 4125 3124 4131 3176
rect 4173 3124 4179 3336
rect 4189 3304 4195 3336
rect 4269 3284 4275 3296
rect 4228 3237 4243 3243
rect 4004 3117 4019 3123
rect 3885 3004 3891 3116
rect 4045 3084 4051 3116
rect 3917 3044 3923 3056
rect 3885 2904 3891 2916
rect 3949 2904 3955 3016
rect 3981 2984 3987 2996
rect 3965 2924 3971 2936
rect 4029 2924 4035 2936
rect 4061 2924 4067 3116
rect 4077 2964 4083 3116
rect 4237 3104 4243 3237
rect 4109 3023 4115 3076
rect 4093 3017 4115 3023
rect 4093 2984 4099 3017
rect 4157 2964 4163 3036
rect 4221 3003 4227 3036
rect 4205 2997 4227 3003
rect 4109 2944 4115 2956
rect 4157 2924 4163 2936
rect 3965 2904 3971 2916
rect 4189 2904 4195 2996
rect 4132 2897 4147 2903
rect 3780 2717 3788 2723
rect 3805 2684 3811 2696
rect 3741 2664 3747 2676
rect 3789 2664 3795 2676
rect 3716 2657 3724 2663
rect 3661 2603 3667 2636
rect 3773 2617 3788 2623
rect 3661 2597 3683 2603
rect 3677 2484 3683 2597
rect 3709 2564 3715 2576
rect 3732 2537 3740 2543
rect 3693 2464 3699 2536
rect 3725 2384 3731 2496
rect 3501 2324 3507 2336
rect 3341 2284 3347 2296
rect 3373 2284 3379 2296
rect 3389 2284 3395 2296
rect 3405 2264 3411 2276
rect 3325 2244 3331 2256
rect 3421 2204 3427 2316
rect 3565 2284 3571 2316
rect 3597 2304 3603 2316
rect 3661 2284 3667 2336
rect 3741 2324 3747 2476
rect 3469 2244 3475 2256
rect 3261 2184 3267 2196
rect 3309 2183 3315 2196
rect 3453 2184 3459 2196
rect 3581 2184 3587 2216
rect 3284 2177 3315 2183
rect 3341 2144 3347 2176
rect 3213 2104 3219 2116
rect 2957 2004 2963 2036
rect 2973 1983 2979 2096
rect 2989 2084 2995 2096
rect 3021 1984 3027 2056
rect 3197 2024 3203 2036
rect 3213 1984 3219 2076
rect 2964 1977 2979 1983
rect 2829 1884 2835 1896
rect 2845 1884 2851 1896
rect 3053 1884 3059 1896
rect 3101 1884 3107 1956
rect 3149 1904 3155 1916
rect 3229 1904 3235 2096
rect 3325 2083 3331 2136
rect 3309 2077 3331 2083
rect 2916 1877 2924 1883
rect 2941 1864 2947 1876
rect 2813 1784 2819 1856
rect 2829 1844 2835 1856
rect 2989 1844 2995 1876
rect 3012 1857 3020 1863
rect 2829 1763 2835 1796
rect 2813 1757 2835 1763
rect 2813 1724 2819 1757
rect 2893 1744 2899 1756
rect 2909 1744 2915 1756
rect 2836 1737 2844 1743
rect 2701 1683 2707 1696
rect 2701 1677 2723 1683
rect 2701 1584 2707 1596
rect 2717 1543 2723 1677
rect 2781 1563 2787 1696
rect 2829 1584 2835 1696
rect 2781 1557 2803 1563
rect 2717 1537 2739 1543
rect 2733 1524 2739 1537
rect 2685 1484 2691 1516
rect 2685 1364 2691 1376
rect 2701 1364 2707 1416
rect 2653 1317 2675 1323
rect 2317 1084 2323 1096
rect 2413 1084 2419 1116
rect 2477 1084 2483 1156
rect 2541 1124 2547 1196
rect 2605 1144 2611 1276
rect 2605 1124 2611 1136
rect 2669 1124 2675 1317
rect 2701 1203 2707 1276
rect 2733 1264 2739 1516
rect 2797 1504 2803 1557
rect 2749 1484 2755 1496
rect 2749 1464 2755 1476
rect 2765 1444 2771 1456
rect 2797 1423 2803 1496
rect 2909 1484 2915 1736
rect 2797 1417 2819 1423
rect 2813 1384 2819 1417
rect 2749 1364 2755 1376
rect 2829 1344 2835 1356
rect 2765 1324 2771 1336
rect 2685 1197 2707 1203
rect 2237 1064 2243 1076
rect 2029 1057 2067 1063
rect 2061 1044 2067 1057
rect 1789 803 1795 836
rect 1853 824 1859 836
rect 1773 797 1795 803
rect 1677 684 1683 776
rect 1757 684 1763 776
rect 1540 677 1555 683
rect 1597 664 1603 676
rect 1613 664 1619 676
rect 1533 644 1539 656
rect 1421 564 1427 636
rect 1485 624 1491 636
rect 1437 584 1443 616
rect 1565 584 1571 596
rect 1540 577 1548 583
rect 1437 544 1443 576
rect 1485 564 1491 576
rect 1501 444 1507 536
rect 1469 403 1475 436
rect 1453 397 1475 403
rect 1357 277 1379 283
rect 1357 263 1363 277
rect 1405 264 1411 316
rect 1453 283 1459 397
rect 1444 277 1459 283
rect 1517 264 1523 276
rect 1533 264 1539 376
rect 1549 364 1555 436
rect 1565 284 1571 576
rect 1597 564 1603 596
rect 1613 564 1619 616
rect 1629 564 1635 676
rect 1725 657 1740 663
rect 1725 644 1731 657
rect 1668 557 1676 563
rect 1732 557 1740 563
rect 1773 543 1779 797
rect 1821 684 1827 696
rect 1869 684 1875 736
rect 1885 724 1891 976
rect 1901 944 1907 996
rect 1965 963 1971 1016
rect 1981 1004 1987 1036
rect 2109 984 2115 1056
rect 2173 983 2179 1036
rect 2189 1004 2195 1036
rect 2157 977 2179 983
rect 1997 964 2003 976
rect 1924 957 1939 963
rect 1965 957 1980 963
rect 1933 923 1939 957
rect 2061 944 2067 956
rect 2157 944 2163 977
rect 1933 917 1955 923
rect 1949 904 1955 917
rect 1981 784 1987 936
rect 2029 844 2035 896
rect 1949 684 1955 756
rect 1869 664 1875 676
rect 1917 657 1932 663
rect 1917 644 1923 657
rect 1917 564 1923 636
rect 1764 537 1779 543
rect 1789 544 1795 556
rect 1837 544 1843 556
rect 1789 537 1790 544
rect 1924 537 1939 543
rect 1581 464 1587 536
rect 1613 384 1619 536
rect 1693 524 1699 536
rect 1933 524 1939 537
rect 1933 504 1939 516
rect 1693 424 1699 436
rect 1725 424 1731 436
rect 1693 284 1699 416
rect 1773 324 1779 336
rect 1645 264 1651 276
rect 1348 257 1363 263
rect 1805 263 1811 436
rect 1853 284 1859 356
rect 1853 264 1859 276
rect 1805 257 1827 263
rect 973 244 979 256
rect 1421 244 1427 256
rect 1469 244 1475 256
rect 1613 244 1619 256
rect 1492 237 1500 243
rect 957 184 963 196
rect 717 164 723 176
rect 845 164 851 176
rect 1021 164 1027 236
rect 1037 184 1043 216
rect 1213 184 1219 236
rect 1293 224 1299 236
rect 1277 184 1283 196
rect 1661 184 1667 256
rect 1677 244 1683 256
rect 1725 244 1731 256
rect 1805 224 1811 236
rect 1309 177 1507 183
rect 1213 157 1228 163
rect 477 137 492 143
rect 557 124 563 136
rect 589 124 595 156
rect 861 144 867 156
rect 605 124 611 136
rect 685 124 691 136
rect 733 124 739 136
rect 797 124 803 136
rect 1021 124 1027 136
rect 1069 123 1075 156
rect 1085 144 1091 156
rect 1101 144 1107 156
rect 1213 144 1219 157
rect 1309 144 1315 177
rect 1501 163 1507 177
rect 1565 177 1619 183
rect 1565 163 1571 177
rect 1613 164 1619 177
rect 1709 177 1747 183
rect 1428 157 1459 163
rect 1501 157 1571 163
rect 1124 137 1132 143
rect 1188 137 1196 143
rect 1236 137 1244 143
rect 1149 123 1155 136
rect 1069 117 1155 123
rect 1341 104 1347 156
rect 1405 104 1411 156
rect 1421 104 1427 136
rect 1364 97 1372 103
rect 637 84 643 96
rect 1437 84 1443 136
rect 1453 84 1459 157
rect 1709 163 1715 177
rect 1645 157 1715 163
rect 1508 137 1523 143
rect 1517 123 1523 137
rect 1517 117 1571 123
rect 1565 104 1571 117
rect 1597 104 1603 156
rect 1645 143 1651 157
rect 1636 137 1651 143
rect 1613 104 1619 136
rect 1709 84 1715 136
rect 1725 64 1731 156
rect 1741 144 1747 177
rect 1757 84 1763 216
rect 1789 164 1795 196
rect 1805 64 1811 76
rect 1741 44 1747 56
rect 461 -37 467 36
rect 445 -43 467 -37
rect 829 -43 835 36
rect 1533 -43 1539 36
rect 1821 -37 1827 257
rect 1853 164 1859 196
rect 1869 164 1875 436
rect 1949 324 1955 656
rect 1965 524 1971 716
rect 1981 544 1987 656
rect 2013 543 2019 836
rect 2077 804 2083 896
rect 2029 724 2035 736
rect 2045 684 2051 756
rect 2093 684 2099 696
rect 2125 684 2131 736
rect 2141 724 2147 936
rect 2173 784 2179 956
rect 2157 663 2163 776
rect 2173 744 2179 776
rect 2141 657 2163 663
rect 2109 644 2115 656
rect 2141 644 2147 657
rect 2045 583 2051 616
rect 2061 604 2067 636
rect 2173 584 2179 596
rect 2045 577 2060 583
rect 2004 537 2019 543
rect 1965 504 1971 516
rect 2093 504 2099 536
rect 2109 523 2115 556
rect 2125 544 2131 556
rect 2109 517 2147 523
rect 2141 504 2147 517
rect 2020 497 2028 503
rect 2045 344 2051 436
rect 2125 364 2131 496
rect 2125 324 2131 356
rect 2157 323 2163 536
rect 2205 363 2211 1056
rect 2285 1004 2291 1076
rect 2429 1064 2435 1076
rect 2301 1044 2307 1056
rect 2493 1044 2499 1056
rect 2237 964 2243 996
rect 2285 984 2291 996
rect 2429 964 2435 996
rect 2301 944 2307 956
rect 2221 924 2227 936
rect 2285 904 2291 916
rect 2221 724 2227 736
rect 2237 684 2243 856
rect 2253 684 2259 816
rect 2269 724 2275 776
rect 2349 724 2355 736
rect 2365 703 2371 956
rect 2493 944 2499 956
rect 2541 944 2547 1116
rect 2621 1084 2627 1116
rect 2653 1077 2668 1083
rect 2404 937 2412 943
rect 2445 924 2451 936
rect 2557 924 2563 1076
rect 2653 1063 2659 1077
rect 2685 1064 2691 1197
rect 2573 1057 2659 1063
rect 2573 1044 2579 1057
rect 2381 784 2387 836
rect 2429 744 2435 916
rect 2461 897 2476 903
rect 2461 803 2467 897
rect 2445 797 2467 803
rect 2445 784 2451 797
rect 2349 697 2371 703
rect 2301 584 2307 636
rect 2221 544 2227 576
rect 2317 563 2323 636
rect 2349 584 2355 697
rect 2429 684 2435 736
rect 2365 664 2371 676
rect 2381 604 2387 636
rect 2445 624 2451 636
rect 2365 597 2380 603
rect 2308 557 2323 563
rect 2365 544 2371 597
rect 2429 544 2435 576
rect 2445 544 2451 576
rect 2308 537 2323 543
rect 2317 524 2323 537
rect 2340 497 2348 503
rect 2413 384 2419 496
rect 2461 484 2467 496
rect 2445 384 2451 416
rect 2148 317 2163 323
rect 2189 357 2211 363
rect 1901 284 1907 316
rect 2029 304 2035 316
rect 2045 284 2051 296
rect 2125 284 2131 296
rect 2189 284 2195 357
rect 2477 343 2483 876
rect 2493 724 2499 876
rect 2509 864 2515 916
rect 2589 903 2595 976
rect 2637 964 2643 1036
rect 2733 1004 2739 1076
rect 2756 1057 2771 1063
rect 2765 1044 2771 1057
rect 2701 984 2707 996
rect 2781 984 2787 1276
rect 2829 1184 2835 1296
rect 2861 1283 2867 1476
rect 2877 1324 2883 1456
rect 2845 1277 2867 1283
rect 2797 1104 2803 1116
rect 2813 984 2819 996
rect 2653 944 2659 976
rect 2621 924 2627 936
rect 2749 904 2755 936
rect 2564 897 2595 903
rect 2724 897 2732 903
rect 2605 884 2611 896
rect 2749 844 2755 876
rect 2765 784 2771 896
rect 2781 884 2787 896
rect 2845 883 2851 1277
rect 2877 1104 2883 1116
rect 2925 1104 2931 1736
rect 2941 1704 2947 1836
rect 3005 1584 3011 1596
rect 2957 1484 2963 1496
rect 2957 1444 2963 1456
rect 3021 1404 3027 1436
rect 3037 1343 3043 1856
rect 3053 1744 3059 1856
rect 3069 1764 3075 1856
rect 3213 1784 3219 1796
rect 3197 1764 3203 1776
rect 3069 1544 3075 1756
rect 3181 1744 3187 1756
rect 3085 1604 3091 1696
rect 3069 1504 3075 1516
rect 3117 1484 3123 1716
rect 3156 1637 3171 1643
rect 3165 1544 3171 1637
rect 3181 1484 3187 1516
rect 3133 1477 3171 1483
rect 3085 1363 3091 1376
rect 3117 1364 3123 1476
rect 3133 1464 3139 1477
rect 3165 1464 3171 1477
rect 3076 1357 3091 1363
rect 3133 1344 3139 1436
rect 3037 1337 3052 1343
rect 3149 1304 3155 1456
rect 3197 1364 3203 1376
rect 3181 1324 3187 1336
rect 3012 1297 3020 1303
rect 2861 1084 2867 1096
rect 2925 1084 2931 1096
rect 3005 1084 3011 1096
rect 3108 1077 3123 1083
rect 2941 984 2947 1056
rect 3069 1044 3075 1056
rect 3085 1024 3091 1056
rect 3005 944 3011 956
rect 3101 944 3107 996
rect 2877 924 2883 936
rect 2845 877 2867 883
rect 2541 724 2547 776
rect 2493 684 2499 696
rect 2557 684 2563 776
rect 2765 764 2771 776
rect 2589 677 2604 683
rect 2493 603 2499 676
rect 2509 623 2515 636
rect 2509 617 2531 623
rect 2493 597 2515 603
rect 2509 544 2515 597
rect 2525 504 2531 617
rect 2564 577 2572 583
rect 2589 563 2595 677
rect 2621 664 2627 736
rect 2669 704 2675 716
rect 2701 584 2707 676
rect 2717 664 2723 716
rect 2749 624 2755 636
rect 2781 584 2787 876
rect 2813 724 2819 776
rect 2845 724 2851 816
rect 2861 724 2867 877
rect 2877 864 2883 896
rect 2893 884 2899 936
rect 3021 904 3027 936
rect 3069 924 3075 936
rect 2893 744 2899 876
rect 2957 784 2963 816
rect 2989 724 2995 896
rect 3021 804 3027 896
rect 3037 884 3043 896
rect 2797 704 2803 716
rect 2637 564 2643 576
rect 2573 557 2595 563
rect 2573 524 2579 557
rect 2797 563 2803 696
rect 2813 684 2819 716
rect 2909 704 2915 716
rect 2781 557 2803 563
rect 2621 544 2627 556
rect 2653 544 2659 556
rect 2685 544 2691 556
rect 2685 537 2686 544
rect 2756 537 2771 543
rect 2765 524 2771 537
rect 2525 484 2531 496
rect 2477 337 2499 343
rect 2413 324 2419 336
rect 2212 317 2220 323
rect 2276 317 2284 323
rect 2468 317 2476 323
rect 2317 284 2323 296
rect 2493 284 2499 337
rect 2541 284 2547 336
rect 1924 277 1932 283
rect 2436 277 2444 283
rect 2109 264 2115 276
rect 2557 264 2563 356
rect 2589 284 2595 336
rect 2653 324 2659 376
rect 2749 324 2755 336
rect 2781 324 2787 557
rect 2813 544 2819 556
rect 2893 544 2899 656
rect 2909 544 2915 696
rect 3053 684 3059 796
rect 3076 777 3084 783
rect 2829 384 2835 396
rect 2637 264 2643 276
rect 1917 244 1923 256
rect 2317 244 2323 256
rect 2573 244 2579 256
rect 1981 183 1987 236
rect 1965 177 1987 183
rect 1965 144 1971 177
rect 1997 163 2003 236
rect 2061 163 2067 236
rect 1988 157 2003 163
rect 2029 157 2067 163
rect 2077 157 2108 163
rect 2029 143 2035 157
rect 2020 137 2035 143
rect 2045 137 2046 143
rect 2077 143 2083 157
rect 2285 144 2291 196
rect 2301 184 2307 236
rect 2365 164 2371 176
rect 2054 137 2083 143
rect 2381 143 2387 236
rect 2701 184 2707 276
rect 2765 184 2771 316
rect 2564 177 2572 183
rect 2429 164 2435 176
rect 2621 164 2627 176
rect 2493 144 2499 156
rect 2605 144 2611 156
rect 2372 137 2387 143
rect 2436 137 2451 143
rect 1837 104 1843 136
rect 1981 123 1987 136
rect 1949 117 1987 123
rect 1949 84 1955 117
rect 2109 104 2115 136
rect 2125 124 2131 136
rect 2221 104 2227 136
rect 2445 124 2451 137
rect 2173 84 2179 96
rect 2477 84 2483 96
rect 2253 44 2259 56
rect 1821 -43 1859 -37
rect 2493 -43 2499 136
rect 2557 124 2563 136
rect 2637 124 2643 136
rect 2541 104 2547 116
rect 2669 104 2675 116
rect 2669 -43 2675 96
rect 2685 44 2691 136
rect 2717 -43 2723 36
rect 2749 -43 2755 96
rect 2781 -43 2787 136
rect 2797 124 2803 176
rect 2829 144 2835 156
rect 2845 144 2851 516
rect 2989 504 2995 556
rect 3005 544 3011 676
rect 3021 564 3027 616
rect 3005 504 3011 536
rect 2861 344 2867 496
rect 2909 484 2915 496
rect 2877 284 2883 456
rect 2941 403 2947 436
rect 2989 404 2995 496
rect 2941 397 2963 403
rect 2957 324 2963 397
rect 3005 384 3011 416
rect 3021 283 3027 556
rect 3037 524 3043 536
rect 3053 504 3059 676
rect 3085 584 3091 676
rect 3101 664 3107 936
rect 3117 744 3123 1077
rect 3149 1044 3155 1056
rect 3165 1024 3171 1076
rect 3181 1024 3187 1316
rect 3197 1184 3203 1316
rect 3213 1244 3219 1256
rect 3197 1104 3203 1176
rect 3229 1084 3235 1856
rect 3245 1804 3251 1916
rect 3261 1884 3267 1936
rect 3277 1804 3283 1876
rect 3261 1744 3267 1776
rect 3245 1604 3251 1696
rect 3293 1684 3299 1696
rect 3277 1524 3283 1536
rect 3261 1484 3267 1496
rect 3261 1444 3267 1456
rect 3245 1384 3251 1436
rect 3277 1404 3283 1476
rect 3309 1384 3315 2077
rect 3341 2024 3347 2096
rect 3357 2084 3363 2096
rect 3405 2084 3411 2136
rect 3421 2104 3427 2176
rect 3597 2164 3603 2176
rect 3661 2164 3667 2216
rect 3677 2164 3683 2296
rect 3613 2144 3619 2156
rect 3709 2144 3715 2236
rect 3741 2184 3747 2256
rect 3501 2104 3507 2136
rect 3501 2084 3507 2096
rect 3389 2064 3395 2076
rect 3517 2064 3523 2136
rect 3373 2024 3379 2056
rect 3469 2044 3475 2056
rect 3469 1924 3475 2036
rect 3517 1924 3523 1936
rect 3341 1884 3347 1916
rect 3357 1804 3363 1916
rect 3421 1884 3427 1896
rect 3405 1824 3411 1856
rect 3405 1784 3411 1796
rect 3389 1744 3395 1756
rect 3325 1584 3331 1596
rect 3357 1524 3363 1696
rect 3373 1404 3379 1736
rect 3469 1724 3475 1736
rect 3437 1704 3443 1716
rect 3453 1704 3459 1716
rect 3485 1504 3491 1696
rect 3501 1504 3507 1796
rect 3517 1784 3523 1896
rect 3533 1884 3539 2096
rect 3540 1857 3555 1863
rect 3549 1844 3555 1857
rect 3501 1484 3507 1496
rect 3421 1464 3427 1476
rect 3389 1424 3395 1436
rect 3405 1404 3411 1456
rect 3517 1424 3523 1456
rect 3549 1444 3555 1836
rect 3597 1803 3603 1876
rect 3629 1823 3635 2136
rect 3661 1984 3667 2136
rect 3677 2124 3683 2136
rect 3629 1817 3651 1823
rect 3597 1797 3619 1803
rect 3565 1744 3571 1776
rect 3597 1763 3603 1776
rect 3588 1757 3603 1763
rect 3613 1684 3619 1797
rect 3645 1744 3651 1817
rect 3661 1764 3667 1776
rect 3677 1764 3683 2116
rect 3693 2037 3708 2043
rect 3693 1904 3699 2037
rect 3604 1537 3612 1543
rect 3565 1524 3571 1536
rect 3693 1484 3699 1876
rect 3725 1864 3731 1876
rect 3709 1844 3715 1856
rect 3741 1804 3747 1896
rect 3741 1664 3747 1696
rect 3725 1584 3731 1596
rect 3629 1464 3635 1476
rect 3725 1464 3731 1536
rect 3757 1524 3763 2616
rect 3773 2584 3779 2617
rect 3837 2584 3843 2736
rect 3885 2704 3891 2816
rect 3917 2724 3923 2756
rect 3997 2724 4003 2836
rect 4013 2784 4019 2896
rect 4093 2724 4099 2756
rect 4125 2724 4131 2736
rect 3860 2697 3868 2703
rect 3917 2684 3923 2696
rect 4093 2684 4099 2696
rect 4141 2683 4147 2897
rect 4189 2723 4195 2756
rect 4205 2744 4211 2997
rect 4189 2717 4204 2723
rect 4221 2684 4227 2756
rect 4237 2744 4243 2836
rect 4253 2764 4259 2976
rect 4269 2944 4275 3156
rect 4333 3124 4339 3296
rect 4413 3264 4419 3356
rect 4429 3344 4435 3356
rect 4605 3344 4611 3476
rect 4621 3404 4627 3476
rect 4484 3337 4492 3343
rect 4445 3244 4451 3336
rect 4509 3284 4515 3296
rect 4365 3124 4371 3236
rect 4381 3124 4387 3156
rect 4349 3077 4364 3083
rect 4349 3064 4355 3077
rect 4285 2944 4291 3016
rect 4301 2964 4307 3036
rect 4365 2984 4371 3056
rect 4269 2904 4275 2936
rect 4301 2924 4307 2936
rect 4333 2903 4339 2956
rect 4397 2943 4403 3116
rect 4445 3084 4451 3236
rect 4557 3224 4563 3236
rect 4589 3124 4595 3156
rect 4525 3064 4531 3096
rect 4605 3084 4611 3116
rect 4637 3084 4643 3376
rect 4653 3344 4659 3496
rect 4669 3424 4675 3436
rect 4685 3404 4691 3436
rect 4669 3344 4675 3356
rect 4717 3344 4723 3476
rect 4781 3384 4787 3656
rect 4845 3624 4851 3696
rect 4861 3484 4867 3716
rect 4893 3644 4899 3876
rect 4941 3784 4947 3856
rect 5053 3804 5059 3836
rect 5101 3804 5107 3916
rect 5149 3904 5155 3916
rect 5117 3864 5123 3876
rect 5197 3824 5203 3876
rect 5133 3784 5139 3796
rect 4909 3724 4915 3756
rect 4941 3724 4947 3756
rect 4941 3684 4947 3716
rect 5021 3684 5027 3696
rect 5005 3524 5011 3616
rect 5053 3524 5059 3636
rect 4957 3484 4963 3496
rect 5069 3484 5075 3516
rect 4845 3464 4851 3476
rect 4909 3464 4915 3476
rect 4756 3377 4764 3383
rect 4733 3364 4739 3376
rect 4781 3264 4787 3376
rect 4797 3344 4803 3436
rect 4861 3423 4867 3456
rect 4941 3424 4947 3456
rect 4861 3417 4883 3423
rect 4877 3384 4883 3417
rect 4941 3384 4947 3396
rect 4845 3324 4851 3336
rect 4797 3304 4803 3316
rect 4708 3117 4716 3123
rect 4429 3044 4435 3056
rect 4621 3044 4627 3056
rect 4413 3004 4419 3036
rect 4493 3024 4499 3036
rect 4557 3024 4563 3036
rect 4493 2964 4499 2976
rect 4397 2937 4412 2943
rect 4324 2897 4339 2903
rect 4397 2884 4403 2896
rect 4429 2864 4435 2936
rect 4445 2904 4451 2916
rect 4525 2904 4531 2916
rect 4317 2724 4323 2756
rect 4397 2704 4403 2716
rect 4301 2684 4307 2696
rect 4349 2684 4355 2696
rect 4413 2684 4419 2856
rect 4125 2677 4147 2683
rect 3901 2544 3907 2636
rect 3981 2624 3987 2676
rect 3981 2604 3987 2616
rect 4029 2603 4035 2636
rect 4013 2597 4035 2603
rect 3917 2544 3923 2556
rect 3933 2544 3939 2576
rect 3853 2524 3859 2536
rect 4013 2504 4019 2597
rect 4045 2583 4051 2636
rect 4029 2577 4051 2583
rect 4029 2544 4035 2577
rect 4061 2524 4067 2536
rect 4077 2524 4083 2596
rect 4109 2584 4115 2676
rect 3805 2484 3811 2496
rect 3885 2404 3891 2496
rect 3981 2484 3987 2496
rect 3965 2344 3971 2436
rect 4045 2384 4051 2496
rect 3933 2324 3939 2336
rect 3805 2263 3811 2316
rect 3869 2304 3875 2316
rect 3853 2264 3859 2276
rect 3997 2264 4003 2336
rect 4013 2284 4019 2296
rect 3789 2257 3811 2263
rect 3773 2204 3779 2236
rect 3789 2184 3795 2257
rect 4036 2257 4044 2263
rect 3837 2184 3843 2236
rect 3885 2184 3891 2236
rect 3917 2184 3923 2236
rect 3901 2164 3907 2176
rect 3965 2164 3971 2236
rect 4029 2184 4035 2236
rect 4045 2224 4051 2236
rect 3981 2164 3987 2176
rect 3837 2144 3843 2156
rect 3805 1884 3811 2136
rect 3828 2097 3836 2103
rect 3853 2044 3859 2136
rect 3933 2104 3939 2156
rect 4061 2144 4067 2516
rect 4077 2324 4083 2336
rect 4093 2304 4099 2336
rect 3933 1924 3939 2096
rect 3965 2083 3971 2136
rect 3949 2077 3971 2083
rect 3789 1824 3795 1856
rect 3773 1784 3779 1796
rect 3780 1757 3788 1763
rect 3805 1744 3811 1856
rect 3853 1844 3859 1856
rect 3949 1823 3955 2077
rect 4013 1924 4019 1976
rect 4077 1943 4083 2216
rect 4125 2184 4131 2677
rect 4244 2677 4252 2683
rect 4173 2544 4179 2636
rect 4205 2544 4211 2656
rect 4237 2564 4243 2576
rect 4221 2544 4227 2556
rect 4285 2544 4291 2636
rect 4301 2584 4307 2676
rect 4349 2544 4355 2596
rect 4365 2584 4371 2636
rect 4461 2584 4467 2716
rect 4493 2684 4499 2696
rect 4509 2624 4515 2716
rect 4525 2623 4531 2876
rect 4589 2724 4595 2736
rect 4573 2683 4579 2696
rect 4557 2677 4579 2683
rect 4557 2623 4563 2677
rect 4525 2617 4563 2623
rect 4493 2584 4499 2596
rect 4477 2564 4483 2576
rect 4541 2544 4547 2617
rect 4605 2604 4611 2676
rect 4605 2544 4611 2576
rect 4621 2564 4627 2576
rect 4637 2544 4643 3016
rect 4653 2924 4659 3116
rect 4685 3084 4691 3096
rect 4781 3084 4787 3096
rect 4669 3044 4675 3056
rect 4685 2984 4691 3056
rect 4733 2984 4739 3036
rect 4733 2944 4739 2956
rect 4781 2944 4787 3076
rect 4813 3064 4819 3116
rect 4845 3104 4851 3316
rect 4909 3304 4915 3356
rect 4957 3344 4963 3476
rect 5101 3464 5107 3736
rect 5117 3603 5123 3756
rect 5172 3737 5180 3743
rect 5197 3724 5203 3736
rect 5213 3683 5219 3916
rect 5469 3904 5475 3916
rect 5309 3864 5315 3876
rect 5245 3804 5251 3836
rect 5261 3824 5267 3836
rect 5341 3784 5347 3896
rect 5437 3804 5443 3836
rect 5453 3784 5459 3876
rect 5261 3764 5267 3776
rect 5517 3764 5523 3836
rect 5236 3737 5244 3743
rect 5213 3677 5235 3683
rect 5117 3597 5139 3603
rect 5133 3464 5139 3597
rect 5165 3464 5171 3636
rect 5213 3464 5219 3476
rect 4989 3404 4995 3436
rect 5021 3344 5027 3456
rect 5117 3404 5123 3436
rect 5133 3384 5139 3456
rect 5069 3364 5075 3376
rect 5124 3357 5132 3363
rect 4925 3324 4931 3336
rect 4989 3304 4995 3336
rect 5149 3324 5155 3336
rect 4893 3124 4899 3136
rect 4861 3084 4867 3096
rect 4836 3077 4844 3083
rect 4877 3064 4883 3076
rect 4877 3024 4883 3056
rect 4797 2964 4803 2976
rect 4861 2944 4867 2996
rect 4909 2964 4915 3296
rect 4941 3003 4947 3036
rect 4925 2997 4947 3003
rect 4781 2924 4787 2936
rect 4740 2917 4748 2923
rect 4653 2904 4659 2916
rect 4845 2884 4851 2896
rect 4925 2863 4931 2997
rect 4941 2964 4947 2976
rect 4957 2924 4963 3296
rect 4973 3244 4979 3296
rect 4973 3124 4979 3136
rect 5053 3124 5059 3136
rect 5101 3124 5107 3156
rect 4989 3104 4995 3116
rect 5021 3084 5027 3096
rect 5117 3084 5123 3096
rect 5021 3004 5027 3076
rect 5149 3064 5155 3076
rect 5165 3064 5171 3456
rect 5197 3444 5203 3456
rect 5197 3384 5203 3436
rect 5197 3344 5203 3356
rect 5229 3324 5235 3677
rect 5277 3624 5283 3736
rect 5325 3664 5331 3756
rect 5341 3724 5347 3736
rect 5453 3544 5459 3736
rect 5437 3523 5443 3536
rect 5581 3524 5587 3636
rect 5437 3517 5452 3523
rect 5341 3424 5347 3516
rect 5517 3484 5523 3496
rect 5309 3384 5315 3396
rect 5373 3364 5379 3436
rect 5389 3404 5395 3476
rect 5453 3384 5459 3476
rect 5501 3384 5507 3436
rect 5389 3364 5395 3376
rect 5517 3363 5523 3476
rect 5501 3357 5523 3363
rect 5405 3344 5411 3356
rect 5501 3344 5507 3357
rect 5517 3324 5523 3336
rect 5181 3184 5187 3216
rect 5197 3124 5203 3236
rect 5213 3164 5219 3296
rect 5261 3104 5267 3316
rect 5341 3124 5347 3236
rect 5357 3224 5363 3296
rect 5485 3284 5491 3296
rect 5396 3117 5404 3123
rect 5268 3057 5276 3063
rect 5133 3044 5139 3056
rect 4973 2944 4979 2996
rect 5117 2984 5123 3016
rect 5245 3004 5251 3036
rect 5325 3024 5331 3076
rect 5373 3004 5379 3036
rect 5309 2984 5315 2996
rect 4989 2964 4995 2976
rect 5325 2964 5331 2976
rect 5005 2944 5011 2956
rect 5021 2944 5027 2956
rect 5261 2944 5267 2956
rect 5341 2944 5347 2956
rect 5389 2944 5395 3076
rect 5421 2984 5427 3276
rect 5565 3244 5571 3436
rect 5469 3124 5475 3156
rect 5581 3124 5587 3236
rect 5453 3084 5459 3116
rect 5508 3077 5516 3083
rect 5501 2963 5507 3036
rect 5517 2984 5523 3016
rect 5565 2984 5571 2996
rect 5501 2957 5523 2963
rect 5517 2944 5523 2957
rect 4925 2857 4947 2863
rect 4813 2744 4819 2836
rect 4685 2724 4691 2736
rect 4925 2724 4931 2836
rect 4861 2684 4867 2696
rect 4909 2683 4915 2716
rect 4941 2704 4947 2857
rect 5028 2717 5036 2723
rect 4925 2684 4931 2696
rect 5005 2684 5011 2716
rect 4893 2677 4915 2683
rect 4653 2544 4659 2676
rect 4685 2664 4691 2676
rect 4733 2544 4739 2636
rect 4877 2584 4883 2616
rect 4365 2524 4371 2536
rect 4461 2524 4467 2536
rect 4637 2524 4643 2536
rect 4685 2524 4691 2536
rect 4237 2384 4243 2396
rect 4189 2324 4195 2376
rect 4260 2297 4268 2303
rect 4285 2284 4291 2296
rect 4317 2284 4323 2296
rect 4141 2264 4147 2276
rect 4157 2244 4163 2256
rect 4157 2224 4163 2236
rect 4100 2157 4108 2163
rect 4141 2143 4147 2196
rect 4157 2184 4163 2196
rect 4116 2137 4147 2143
rect 4093 2124 4099 2136
rect 4173 2124 4179 2236
rect 4221 2204 4227 2236
rect 4301 2224 4307 2256
rect 4333 2244 4339 2496
rect 4381 2324 4387 2496
rect 4429 2404 4435 2436
rect 4509 2324 4515 2476
rect 4525 2364 4531 2496
rect 4845 2383 4851 2516
rect 4893 2444 4899 2677
rect 4948 2677 4963 2683
rect 4941 2564 4947 2656
rect 4925 2524 4931 2536
rect 4941 2524 4947 2536
rect 4916 2497 4924 2503
rect 4845 2377 4860 2383
rect 4557 2337 4659 2343
rect 4557 2324 4563 2337
rect 4653 2323 4659 2337
rect 4781 2324 4787 2336
rect 4653 2317 4716 2323
rect 4436 2297 4483 2303
rect 4477 2284 4483 2297
rect 4452 2277 4460 2283
rect 4365 2244 4371 2276
rect 4484 2257 4499 2263
rect 4301 2204 4307 2216
rect 4221 2164 4227 2176
rect 4260 2157 4323 2163
rect 4317 2143 4323 2157
rect 4365 2163 4371 2176
rect 4356 2157 4371 2163
rect 4413 2144 4419 2156
rect 4461 2144 4467 2256
rect 4477 2164 4483 2236
rect 4493 2184 4499 2257
rect 4317 2137 4332 2143
rect 4077 1937 4099 1943
rect 4093 1924 4099 1937
rect 4109 1884 4115 1996
rect 4125 1984 4131 2096
rect 4173 2003 4179 2116
rect 4285 2104 4291 2116
rect 4269 2024 4275 2096
rect 4301 2004 4307 2036
rect 4173 1997 4195 2003
rect 4125 1884 4131 1896
rect 3965 1844 3971 1856
rect 3949 1817 3971 1823
rect 3965 1784 3971 1817
rect 3981 1784 3987 1836
rect 4029 1784 4035 1876
rect 4109 1844 4115 1856
rect 4109 1764 4115 1776
rect 3981 1744 3987 1756
rect 3853 1704 3859 1736
rect 3869 1704 3875 1736
rect 3924 1697 3932 1703
rect 3805 1524 3811 1536
rect 3789 1484 3795 1496
rect 3773 1464 3779 1476
rect 3668 1457 3683 1463
rect 3677 1444 3683 1457
rect 3533 1424 3539 1436
rect 3460 1377 3468 1383
rect 3245 1344 3251 1376
rect 3277 1084 3283 1096
rect 3165 944 3171 976
rect 3213 964 3219 1056
rect 3261 984 3267 996
rect 3277 944 3283 1016
rect 3277 924 3283 936
rect 3293 904 3299 1356
rect 3309 1264 3315 1296
rect 3325 1244 3331 1336
rect 3357 1104 3363 1336
rect 3437 1124 3443 1376
rect 3453 1224 3459 1236
rect 3485 1183 3491 1396
rect 3501 1304 3507 1376
rect 3581 1344 3587 1416
rect 3645 1364 3651 1376
rect 3597 1344 3603 1356
rect 3517 1224 3523 1336
rect 3581 1324 3587 1336
rect 3565 1284 3571 1296
rect 3597 1184 3603 1256
rect 3613 1204 3619 1296
rect 3661 1184 3667 1196
rect 3476 1177 3491 1183
rect 3444 1117 3452 1123
rect 3549 1084 3555 1096
rect 3613 1077 3628 1083
rect 3453 1064 3459 1076
rect 3396 1057 3411 1063
rect 3405 1044 3411 1057
rect 3341 964 3347 976
rect 3405 964 3411 976
rect 3437 944 3443 996
rect 3469 964 3475 976
rect 3453 944 3459 956
rect 3293 884 3299 896
rect 3245 844 3251 856
rect 3197 784 3203 816
rect 3220 777 3228 783
rect 3165 684 3171 756
rect 3245 684 3251 836
rect 3357 684 3363 876
rect 3421 684 3427 936
rect 3117 643 3123 676
rect 3133 644 3139 656
rect 3101 637 3123 643
rect 3101 584 3107 637
rect 3037 284 3043 496
rect 3101 464 3107 576
rect 3117 504 3123 616
rect 3133 544 3139 576
rect 3117 484 3123 496
rect 3133 484 3139 536
rect 3181 504 3187 576
rect 3213 564 3219 676
rect 3245 624 3251 676
rect 3261 664 3267 676
rect 3277 644 3283 656
rect 3293 624 3299 676
rect 3357 664 3363 676
rect 3412 657 3427 663
rect 3341 644 3347 656
rect 3277 584 3283 616
rect 3197 483 3203 536
rect 3181 477 3203 483
rect 3133 384 3139 456
rect 3060 377 3068 383
rect 3133 324 3139 376
rect 3165 284 3171 296
rect 3005 277 3027 283
rect 2893 264 2899 276
rect 2909 264 2915 276
rect 2877 184 2883 236
rect 2893 164 2899 176
rect 2957 164 2963 196
rect 3005 164 3011 277
rect 3044 277 3084 283
rect 3101 263 3107 276
rect 3101 257 3123 263
rect 3021 244 3027 256
rect 3069 184 3075 236
rect 3021 164 3027 176
rect 2845 124 2851 136
rect 2893 104 2899 156
rect 3005 144 3011 156
rect 3101 144 3107 176
rect 3005 137 3006 144
rect 2813 -43 2819 96
rect 2909 44 2915 136
rect 2973 44 2979 136
rect 3037 44 3043 136
rect 2941 -43 2947 16
rect 3117 -37 3123 257
rect 3149 244 3155 256
rect 3181 204 3187 477
rect 3213 403 3219 556
rect 3229 544 3235 556
rect 3261 544 3267 556
rect 3325 544 3331 616
rect 3373 584 3379 636
rect 3389 584 3395 616
rect 3357 544 3363 556
rect 3261 537 3262 544
rect 3396 517 3404 523
rect 3197 397 3219 403
rect 3197 384 3203 397
rect 3197 264 3203 376
rect 3245 284 3251 336
rect 3293 284 3299 496
rect 3197 237 3212 243
rect 3149 184 3155 196
rect 3197 144 3203 237
rect 3277 224 3283 256
rect 3293 244 3299 276
rect 3341 264 3347 456
rect 3405 384 3411 416
rect 3357 284 3363 316
rect 3421 264 3427 657
rect 3437 564 3443 936
rect 3485 844 3491 936
rect 3469 724 3475 736
rect 3501 644 3507 1076
rect 3517 1044 3523 1056
rect 3549 804 3555 1076
rect 3565 784 3571 896
rect 3581 704 3587 756
rect 3501 604 3507 636
rect 3533 603 3539 636
rect 3517 597 3539 603
rect 3453 564 3459 576
rect 3469 564 3475 576
rect 3517 544 3523 597
rect 3613 584 3619 1077
rect 3645 1044 3651 1056
rect 3645 964 3651 996
rect 3661 964 3667 1036
rect 3677 984 3683 1436
rect 3693 1384 3699 1456
rect 3709 1403 3715 1436
rect 3709 1397 3731 1403
rect 3709 1364 3715 1376
rect 3693 1344 3699 1356
rect 3709 1324 3715 1336
rect 3725 1184 3731 1397
rect 3821 1364 3827 1696
rect 3981 1524 3987 1696
rect 3997 1664 4003 1696
rect 3917 1517 3964 1523
rect 3917 1484 3923 1517
rect 3933 1484 3939 1496
rect 3837 1403 3843 1436
rect 3837 1397 3859 1403
rect 3741 1324 3747 1336
rect 3693 1084 3699 1096
rect 3741 1064 3747 1076
rect 3757 1064 3763 1356
rect 3789 1344 3795 1356
rect 3789 1124 3795 1216
rect 3805 1164 3811 1296
rect 3709 984 3715 1056
rect 3725 1044 3731 1056
rect 3725 1004 3731 1036
rect 3629 824 3635 936
rect 3645 684 3651 936
rect 3661 764 3667 776
rect 3437 524 3443 536
rect 3437 284 3443 296
rect 3485 284 3491 536
rect 3508 377 3516 383
rect 3325 224 3331 236
rect 3389 224 3395 236
rect 3325 164 3331 176
rect 3389 164 3395 216
rect 3309 144 3315 156
rect 3437 143 3443 276
rect 3533 264 3539 296
rect 3549 284 3555 576
rect 3661 564 3667 656
rect 3629 544 3635 556
rect 3645 544 3651 556
rect 3677 544 3683 916
rect 3565 524 3571 536
rect 3693 484 3699 676
rect 3709 664 3715 716
rect 3725 664 3731 836
rect 3741 684 3747 976
rect 3757 963 3763 1056
rect 3789 984 3795 1036
rect 3821 1024 3827 1356
rect 3853 1344 3859 1397
rect 3917 1384 3923 1436
rect 3933 1404 3939 1416
rect 3869 1304 3875 1356
rect 3885 1284 3891 1336
rect 3860 1277 3875 1283
rect 3869 1263 3875 1277
rect 3917 1263 3923 1356
rect 3869 1257 3923 1263
rect 3869 1084 3875 1096
rect 3933 1084 3939 1396
rect 3981 1364 3987 1476
rect 3949 1323 3955 1336
rect 3949 1317 3971 1323
rect 3965 1304 3971 1317
rect 3949 1284 3955 1296
rect 3981 1284 3987 1336
rect 3853 1044 3859 1056
rect 3837 1004 3843 1036
rect 3853 984 3859 1016
rect 3981 984 3987 996
rect 3956 977 3964 983
rect 3837 964 3843 976
rect 3757 957 3772 963
rect 3821 944 3827 956
rect 3773 924 3779 936
rect 3853 924 3859 956
rect 3901 944 3907 976
rect 3917 944 3923 956
rect 3645 384 3651 416
rect 3588 377 3596 383
rect 3725 383 3731 496
rect 3716 377 3731 383
rect 3597 264 3603 276
rect 3453 164 3459 256
rect 3469 244 3475 256
rect 3469 164 3475 196
rect 3517 184 3523 196
rect 3453 144 3459 156
rect 3581 144 3587 236
rect 3597 184 3603 256
rect 3613 224 3619 276
rect 3677 264 3683 276
rect 3725 264 3731 296
rect 3741 284 3747 476
rect 3757 383 3763 896
rect 3789 703 3795 796
rect 3837 724 3843 916
rect 3885 904 3891 916
rect 3940 897 3955 903
rect 3773 697 3795 703
rect 3821 697 3852 703
rect 3773 584 3779 697
rect 3821 684 3827 697
rect 3876 697 3891 703
rect 3885 684 3891 697
rect 3789 664 3795 676
rect 3805 644 3811 676
rect 3837 623 3843 676
rect 3837 617 3859 623
rect 3789 564 3795 576
rect 3805 544 3811 596
rect 3837 584 3843 596
rect 3853 564 3859 617
rect 3869 544 3875 676
rect 3917 624 3923 656
rect 3933 644 3939 676
rect 3949 603 3955 897
rect 3997 684 4003 1096
rect 4013 1084 4019 1696
rect 4045 1604 4051 1716
rect 4141 1704 4147 1956
rect 4189 1844 4195 1997
rect 4365 1884 4371 1936
rect 4397 1884 4403 2116
rect 4461 1924 4467 2116
rect 4477 1884 4483 1916
rect 4525 1884 4531 2296
rect 4733 2284 4739 2316
rect 4781 2277 4796 2283
rect 4573 2263 4579 2276
rect 4564 2257 4579 2263
rect 4541 2163 4547 2236
rect 4541 2157 4595 2163
rect 4589 2144 4595 2157
rect 4669 2144 4675 2236
rect 4685 2184 4691 2236
rect 4781 2224 4787 2277
rect 4813 2224 4819 2256
rect 4829 2164 4835 2276
rect 4845 2144 4851 2377
rect 4877 2164 4883 2196
rect 4893 2144 4899 2376
rect 4941 2304 4947 2496
rect 4957 2484 4963 2677
rect 5053 2623 5059 2636
rect 5069 2624 5075 2636
rect 5037 2617 5059 2623
rect 4980 2537 4990 2543
rect 5037 2524 5043 2617
rect 5085 2604 5091 2896
rect 5101 2684 5107 2696
rect 5133 2684 5139 2916
rect 5149 2884 5155 2896
rect 5197 2844 5203 2936
rect 5284 2897 5299 2903
rect 5213 2824 5219 2896
rect 5117 2664 5123 2676
rect 5133 2644 5139 2656
rect 5053 2584 5059 2596
rect 5117 2584 5123 2616
rect 5149 2564 5155 2676
rect 5213 2604 5219 2716
rect 5245 2704 5251 2816
rect 5261 2684 5267 2776
rect 5181 2584 5187 2596
rect 5261 2564 5267 2656
rect 5277 2644 5283 2716
rect 5293 2664 5299 2897
rect 5341 2803 5347 2936
rect 5501 2924 5507 2936
rect 5453 2904 5459 2916
rect 5405 2884 5411 2896
rect 5341 2797 5363 2803
rect 5341 2724 5347 2736
rect 5325 2684 5331 2696
rect 5309 2604 5315 2636
rect 5069 2524 5075 2536
rect 5229 2524 5235 2556
rect 5245 2537 5260 2543
rect 5021 2384 5027 2496
rect 5021 2324 5027 2336
rect 4909 2264 4915 2276
rect 4932 2257 4940 2263
rect 4564 2137 4572 2143
rect 4548 2117 4556 2123
rect 4669 2104 4675 2136
rect 4893 2124 4899 2136
rect 4324 1877 4332 1883
rect 4509 1877 4524 1883
rect 4061 1684 4067 1696
rect 4141 1544 4147 1696
rect 4173 1684 4179 1836
rect 4221 1804 4227 1876
rect 4333 1857 4348 1863
rect 4333 1784 4339 1857
rect 4413 1804 4419 1836
rect 4365 1784 4371 1796
rect 4301 1764 4307 1776
rect 4461 1744 4467 1876
rect 4477 1744 4483 1756
rect 4301 1703 4307 1736
rect 4317 1724 4323 1736
rect 4301 1697 4323 1703
rect 4205 1684 4211 1696
rect 4269 1604 4275 1696
rect 4317 1684 4323 1697
rect 4413 1684 4419 1716
rect 4285 1584 4291 1656
rect 4365 1584 4371 1596
rect 4493 1584 4499 1636
rect 4260 1537 4323 1543
rect 4173 1524 4179 1536
rect 4317 1523 4323 1537
rect 4317 1517 4332 1523
rect 4093 1484 4099 1496
rect 4157 1484 4163 1516
rect 4349 1484 4355 1576
rect 4413 1504 4419 1516
rect 4260 1477 4275 1483
rect 4077 1464 4083 1476
rect 4173 1464 4179 1476
rect 4237 1464 4243 1476
rect 4109 1423 4115 1436
rect 4109 1417 4131 1423
rect 4045 1384 4051 1396
rect 4109 1384 4115 1396
rect 4029 1364 4035 1376
rect 4125 1363 4131 1417
rect 4109 1357 4131 1363
rect 4093 1344 4099 1356
rect 4109 1303 4115 1357
rect 4157 1344 4163 1356
rect 4125 1324 4131 1336
rect 4100 1297 4115 1303
rect 4061 1124 4067 1236
rect 4052 1097 4060 1103
rect 4013 1064 4019 1076
rect 4029 1044 4035 1056
rect 4045 944 4051 956
rect 4029 804 4035 936
rect 4061 884 4067 896
rect 4036 757 4044 763
rect 3965 664 3971 676
rect 4061 664 4067 676
rect 3988 657 3996 663
rect 4045 604 4051 656
rect 4077 623 4083 1276
rect 4125 1223 4131 1316
rect 4141 1284 4147 1296
rect 4109 1217 4131 1223
rect 4109 1184 4115 1217
rect 4157 1144 4163 1336
rect 4173 1324 4179 1336
rect 4189 1304 4195 1456
rect 4205 1084 4211 1456
rect 4237 1444 4243 1456
rect 4221 1404 4227 1436
rect 4237 1344 4243 1356
rect 4253 1283 4259 1296
rect 4269 1284 4275 1477
rect 4301 1344 4307 1436
rect 4365 1324 4371 1336
rect 4381 1304 4387 1336
rect 4308 1297 4316 1303
rect 4244 1277 4259 1283
rect 4333 1124 4339 1136
rect 4349 1104 4355 1116
rect 4397 1104 4403 1436
rect 4429 1324 4435 1336
rect 4461 1143 4467 1476
rect 4477 1464 4483 1496
rect 4509 1464 4515 1877
rect 4573 1864 4579 1876
rect 4621 1864 4627 2096
rect 4637 1904 4643 2076
rect 4637 1884 4643 1896
rect 4541 1844 4547 1856
rect 4621 1844 4627 1856
rect 4525 1664 4531 1696
rect 4525 1524 4531 1576
rect 4541 1484 4547 1576
rect 4477 1384 4483 1456
rect 4493 1363 4499 1436
rect 4477 1357 4499 1363
rect 4477 1324 4483 1357
rect 4493 1304 4499 1336
rect 4557 1324 4563 1336
rect 4445 1137 4467 1143
rect 4269 1084 4275 1096
rect 4189 1077 4204 1083
rect 4093 984 4099 1016
rect 4109 744 4115 956
rect 4125 944 4131 1036
rect 4125 724 4131 736
rect 4109 664 4115 676
rect 4093 644 4099 656
rect 4077 617 4099 623
rect 3949 597 3971 603
rect 3965 584 3971 597
rect 3981 564 3987 596
rect 3997 544 4003 596
rect 3869 524 3875 536
rect 3917 424 3923 496
rect 3757 377 3772 383
rect 3908 377 3916 383
rect 3805 284 3811 296
rect 3853 264 3859 316
rect 3869 284 3875 316
rect 3661 224 3667 256
rect 3789 244 3795 256
rect 3597 144 3603 156
rect 3757 144 3763 176
rect 3773 164 3779 196
rect 3901 184 3907 356
rect 3917 264 3923 336
rect 3933 284 3939 316
rect 3997 284 4003 536
rect 4013 304 4019 596
rect 4093 584 4099 617
rect 4141 544 4147 1076
rect 4157 784 4163 816
rect 4173 784 4179 836
rect 4173 744 4179 756
rect 4189 704 4195 1077
rect 4292 1057 4307 1063
rect 4221 1004 4227 1056
rect 4301 1044 4307 1057
rect 4237 964 4243 996
rect 4365 984 4371 996
rect 4397 964 4403 1096
rect 4356 957 4364 963
rect 4253 924 4259 936
rect 4228 917 4236 923
rect 4221 884 4227 896
rect 4253 864 4259 916
rect 4276 857 4284 863
rect 4301 844 4307 856
rect 4205 684 4211 696
rect 4205 664 4211 676
rect 4228 657 4243 663
rect 4237 644 4243 657
rect 4157 564 4163 616
rect 4237 584 4243 596
rect 4173 564 4179 576
rect 4141 524 4147 536
rect 4013 264 4019 296
rect 4061 284 4067 296
rect 4125 284 4131 436
rect 4141 284 4147 516
rect 4173 304 4179 556
rect 4189 544 4195 576
rect 4253 504 4259 736
rect 4317 724 4323 956
rect 4413 944 4419 1056
rect 4429 964 4435 976
rect 4445 944 4451 1137
rect 4477 1124 4483 1216
rect 4484 1057 4492 1063
rect 4509 984 4515 1076
rect 4509 924 4515 936
rect 4397 884 4403 896
rect 4413 784 4419 816
rect 4301 704 4307 716
rect 4285 684 4291 696
rect 4301 684 4307 696
rect 4381 684 4387 696
rect 4301 544 4307 616
rect 4349 603 4355 636
rect 4365 604 4371 656
rect 4333 597 4355 603
rect 4253 323 4259 496
rect 4285 384 4291 516
rect 4308 497 4316 503
rect 4333 404 4339 597
rect 4365 564 4371 576
rect 4397 564 4403 776
rect 4461 724 4467 756
rect 4477 684 4483 836
rect 4509 724 4515 736
rect 4493 684 4499 716
rect 4429 624 4435 636
rect 4525 623 4531 1056
rect 4557 1004 4563 1036
rect 4573 943 4579 1836
rect 4621 1764 4627 1796
rect 4637 1744 4643 1756
rect 4589 1704 4595 1736
rect 4637 1524 4643 1576
rect 4621 1484 4627 1516
rect 4589 1464 4595 1476
rect 4621 1364 4627 1376
rect 4605 1324 4611 1336
rect 4589 1164 4595 1296
rect 4605 1084 4611 1156
rect 4637 1124 4643 1416
rect 4621 1104 4627 1116
rect 4605 984 4611 1036
rect 4621 944 4627 956
rect 4573 937 4595 943
rect 4557 804 4563 936
rect 4557 684 4563 756
rect 4573 724 4579 756
rect 4541 624 4547 636
rect 4509 617 4531 623
rect 4413 544 4419 556
rect 4477 544 4483 556
rect 4413 384 4419 476
rect 4461 384 4467 496
rect 4253 317 4268 323
rect 4285 284 4291 296
rect 4109 264 4115 276
rect 4189 244 4195 276
rect 3789 164 3795 176
rect 3805 144 3811 176
rect 3965 164 3971 176
rect 3981 164 3987 236
rect 4093 204 4099 236
rect 4045 164 4051 176
rect 3949 144 3955 156
rect 3997 144 4003 156
rect 4109 144 4115 216
rect 4164 177 4172 183
rect 4205 144 4211 276
rect 4221 164 4227 176
rect 4237 164 4243 276
rect 4301 264 4307 276
rect 4349 164 4355 276
rect 4365 264 4371 356
rect 4381 284 4387 296
rect 4413 284 4419 376
rect 4461 324 4467 336
rect 4493 264 4499 296
rect 4509 284 4515 617
rect 4557 584 4563 596
rect 4557 563 4563 576
rect 4589 564 4595 937
rect 4637 904 4643 1076
rect 4653 1044 4659 2036
rect 4765 1924 4771 1956
rect 4749 1904 4755 1916
rect 4701 1744 4707 1876
rect 4685 1664 4691 1676
rect 4676 1637 4691 1643
rect 4685 1504 4691 1637
rect 4669 1323 4675 1436
rect 4717 1344 4723 1896
rect 4829 1883 4835 2096
rect 4909 1943 4915 2256
rect 4941 2184 4947 2196
rect 4957 2104 4963 2316
rect 5005 2284 5011 2316
rect 5085 2303 5091 2496
rect 5213 2484 5219 2496
rect 5181 2384 5187 2396
rect 5108 2317 5116 2323
rect 5085 2297 5107 2303
rect 4989 2204 4995 2236
rect 5037 2123 5043 2196
rect 5053 2144 5059 2236
rect 5101 2224 5107 2297
rect 5133 2284 5139 2356
rect 5149 2324 5155 2336
rect 5213 2324 5219 2336
rect 5197 2284 5203 2316
rect 5085 2124 5091 2196
rect 5181 2143 5187 2236
rect 5197 2164 5203 2176
rect 5213 2144 5219 2156
rect 5181 2137 5203 2143
rect 5117 2124 5123 2136
rect 5133 2124 5139 2136
rect 5037 2117 5052 2123
rect 5172 2117 5180 2123
rect 4893 1937 4915 1943
rect 4861 1884 4867 1916
rect 4829 1877 4851 1883
rect 4733 1764 4739 1856
rect 4733 1644 4739 1736
rect 4749 1684 4755 1716
rect 4765 1604 4771 1696
rect 4781 1484 4787 1816
rect 4797 1664 4803 1836
rect 4829 1743 4835 1816
rect 4845 1803 4851 1877
rect 4845 1797 4867 1803
rect 4861 1784 4867 1797
rect 4877 1784 4883 1816
rect 4877 1764 4883 1776
rect 4893 1764 4899 1937
rect 4909 1904 4915 1916
rect 4925 1884 4931 1976
rect 4973 1964 4979 2096
rect 4957 1924 4963 1936
rect 5005 1884 5011 2096
rect 5085 1924 5091 2096
rect 5149 2064 5155 2096
rect 5165 1924 5171 1936
rect 5069 1904 5075 1916
rect 5197 1884 5203 2137
rect 5028 1877 5036 1883
rect 5229 1883 5235 2516
rect 5245 2444 5251 2537
rect 5277 2504 5283 2596
rect 5245 2384 5251 2416
rect 5277 1944 5283 2436
rect 5293 2284 5299 2576
rect 5309 2564 5315 2576
rect 5325 2564 5331 2576
rect 5341 2524 5347 2536
rect 5357 2304 5363 2797
rect 5405 2724 5411 2736
rect 5469 2704 5475 2716
rect 5453 2684 5459 2696
rect 5517 2684 5523 2696
rect 5380 2677 5388 2683
rect 5437 2584 5443 2596
rect 5501 2544 5507 2636
rect 5533 2604 5539 2896
rect 5565 2584 5571 2616
rect 5581 2544 5587 2636
rect 5501 2504 5507 2516
rect 5389 2484 5395 2496
rect 5469 2404 5475 2496
rect 5533 2464 5539 2496
rect 5501 2384 5507 2396
rect 5508 2317 5516 2323
rect 5341 2277 5356 2283
rect 5309 2244 5315 2256
rect 5325 2184 5331 2196
rect 5309 2164 5315 2176
rect 5220 1877 5235 1883
rect 4941 1763 4947 1876
rect 5005 1864 5011 1876
rect 4989 1784 4995 1796
rect 4925 1757 4947 1763
rect 4893 1744 4899 1756
rect 4820 1737 4835 1743
rect 4925 1704 4931 1757
rect 4996 1757 5004 1763
rect 5069 1744 5075 1756
rect 5005 1724 5011 1736
rect 4836 1697 4851 1703
rect 4797 1584 4803 1636
rect 4733 1364 4739 1436
rect 4781 1364 4787 1476
rect 4797 1464 4803 1516
rect 4813 1464 4819 1676
rect 4797 1364 4803 1456
rect 4813 1444 4819 1456
rect 4829 1424 4835 1476
rect 4845 1384 4851 1697
rect 4861 1584 4867 1596
rect 4861 1564 4867 1576
rect 4861 1544 4867 1556
rect 4877 1524 4883 1536
rect 4877 1484 4883 1496
rect 4925 1483 4931 1596
rect 4948 1537 4956 1543
rect 4973 1484 4979 1496
rect 4989 1484 4995 1576
rect 4909 1477 4931 1483
rect 4861 1403 4867 1436
rect 4861 1397 4883 1403
rect 4861 1364 4867 1376
rect 4797 1344 4803 1356
rect 4877 1344 4883 1397
rect 4909 1364 4915 1477
rect 4925 1403 4931 1436
rect 4989 1424 4995 1456
rect 4925 1397 4947 1403
rect 4941 1364 4947 1397
rect 4957 1344 4963 1356
rect 5005 1344 5011 1556
rect 5021 1524 5027 1556
rect 4669 1317 4691 1323
rect 4685 1143 4691 1317
rect 4669 1137 4691 1143
rect 4669 1063 4675 1137
rect 4692 1117 4700 1123
rect 4717 1103 4723 1196
rect 4740 1117 4748 1123
rect 4765 1104 4771 1116
rect 4685 1097 4723 1103
rect 4685 1084 4691 1097
rect 4781 1084 4787 1336
rect 4813 1244 4819 1336
rect 4829 1284 4835 1296
rect 4820 1117 4828 1123
rect 4845 1104 4851 1336
rect 4845 1084 4851 1096
rect 4701 1077 4748 1083
rect 4701 1063 4707 1077
rect 4861 1064 4867 1096
rect 4669 1057 4707 1063
rect 4877 1043 4883 1116
rect 4861 1037 4883 1043
rect 4653 923 4659 996
rect 4669 943 4675 1036
rect 4685 964 4691 996
rect 4701 944 4707 996
rect 4733 984 4739 996
rect 4749 944 4755 1016
rect 4797 1003 4803 1036
rect 4781 997 4803 1003
rect 4669 937 4691 943
rect 4653 917 4668 923
rect 4685 923 4691 937
rect 4685 917 4723 923
rect 4717 903 4723 917
rect 4717 897 4755 903
rect 4605 604 4611 636
rect 4637 584 4643 896
rect 4749 883 4755 897
rect 4781 903 4787 997
rect 4861 984 4867 1037
rect 4877 984 4883 996
rect 4813 904 4819 916
rect 4772 897 4787 903
rect 4829 883 4835 896
rect 4749 877 4835 883
rect 4804 857 4812 863
rect 4893 844 4899 1296
rect 4909 1077 4924 1083
rect 4909 1004 4915 1077
rect 4925 944 4931 996
rect 4957 943 4963 1336
rect 5037 1283 5043 1716
rect 5085 1704 5091 1876
rect 5229 1864 5235 1877
rect 5197 1844 5203 1856
rect 5117 1743 5123 1836
rect 5133 1764 5139 1776
rect 5117 1737 5139 1743
rect 5117 1564 5123 1636
rect 5101 1524 5107 1536
rect 5133 1524 5139 1737
rect 5181 1563 5187 1836
rect 5197 1624 5203 1716
rect 5181 1557 5203 1563
rect 5085 1483 5091 1496
rect 5197 1484 5203 1557
rect 5085 1477 5132 1483
rect 5053 1364 5059 1436
rect 5069 1364 5075 1436
rect 5117 1384 5123 1396
rect 5133 1364 5139 1376
rect 5021 1277 5043 1283
rect 5021 1124 5027 1277
rect 5069 1184 5075 1336
rect 5085 1284 5091 1296
rect 5085 1124 5091 1176
rect 4973 1063 4979 1116
rect 4989 1084 4995 1116
rect 5149 1084 5155 1096
rect 4973 1057 4995 1063
rect 4989 984 4995 1057
rect 5069 1044 5075 1076
rect 5133 1064 5139 1076
rect 5053 983 5059 1036
rect 5053 977 5075 983
rect 5069 964 5075 977
rect 5037 944 5043 956
rect 5053 944 5059 956
rect 5085 944 5091 1056
rect 5117 964 5123 1036
rect 5133 964 5139 976
rect 4957 937 4979 943
rect 4653 724 4659 776
rect 4788 737 4796 743
rect 4669 684 4675 736
rect 4685 684 4691 696
rect 4749 664 4755 736
rect 4765 684 4771 736
rect 4813 664 4819 756
rect 4829 684 4835 816
rect 4845 684 4851 776
rect 4861 684 4867 696
rect 4548 557 4563 563
rect 4589 504 4595 556
rect 4605 544 4611 576
rect 4669 564 4675 596
rect 4797 584 4803 596
rect 4589 484 4595 496
rect 4621 304 4627 436
rect 4653 284 4659 536
rect 4429 164 4435 236
rect 4605 224 4611 236
rect 4669 184 4675 236
rect 4253 144 4259 156
rect 3428 137 3443 143
rect 3476 137 3484 143
rect 3405 124 3411 136
rect 3533 124 3539 136
rect 4333 124 4339 136
rect 3268 117 3292 123
rect 4084 117 4115 123
rect 4109 104 4115 117
rect 4372 117 4380 123
rect 4509 104 4515 176
rect 4701 143 4707 556
rect 4845 544 4851 676
rect 4877 664 4883 756
rect 4893 684 4899 696
rect 4909 604 4915 896
rect 4941 884 4947 936
rect 4941 684 4947 696
rect 4884 577 4892 583
rect 4861 564 4867 576
rect 4717 524 4723 536
rect 4717 284 4723 316
rect 4717 164 4723 276
rect 4733 264 4739 396
rect 4733 164 4739 216
rect 4749 184 4755 236
rect 4765 224 4771 356
rect 4797 304 4803 376
rect 4781 204 4787 296
rect 4845 284 4851 296
rect 4861 264 4867 556
rect 4973 544 4979 937
rect 5037 724 5043 736
rect 5085 664 5091 676
rect 5069 644 5075 656
rect 4989 604 4995 636
rect 5005 604 5011 636
rect 4989 564 4995 576
rect 5037 544 5043 576
rect 5053 564 5059 596
rect 5069 564 5075 596
rect 4925 464 4931 536
rect 4941 384 4947 436
rect 4893 324 4899 336
rect 4989 324 4995 536
rect 5037 304 5043 516
rect 5101 324 5107 956
rect 5149 944 5155 1036
rect 5124 717 5132 723
rect 5149 704 5155 936
rect 5165 884 5171 1476
rect 5181 1344 5187 1436
rect 5197 1344 5203 1356
rect 5181 1204 5187 1296
rect 5213 1124 5219 1136
rect 5229 1084 5235 1856
rect 5277 1804 5283 1916
rect 5293 1904 5299 2136
rect 5341 2084 5347 2277
rect 5389 2264 5395 2276
rect 5373 2244 5379 2256
rect 5405 2184 5411 2316
rect 5549 2284 5555 2296
rect 5437 2203 5443 2236
rect 5453 2204 5459 2276
rect 5565 2264 5571 2276
rect 5421 2197 5443 2203
rect 5389 2144 5395 2156
rect 5357 2044 5363 2096
rect 5405 2084 5411 2096
rect 5421 1944 5427 2197
rect 5469 2084 5475 2096
rect 5437 1984 5443 1996
rect 5341 1924 5347 1936
rect 5293 1884 5299 1896
rect 5325 1884 5331 1916
rect 5453 1884 5459 2076
rect 5389 1823 5395 1856
rect 5373 1817 5395 1823
rect 5245 1784 5251 1796
rect 5373 1784 5379 1817
rect 5437 1784 5443 1796
rect 5261 1764 5267 1776
rect 5277 1543 5283 1776
rect 5373 1764 5379 1776
rect 5485 1744 5491 2236
rect 5501 2184 5507 2196
rect 5508 1877 5516 1883
rect 5501 1783 5507 1836
rect 5533 1804 5539 1916
rect 5565 1824 5571 1836
rect 5565 1784 5571 1796
rect 5501 1777 5523 1783
rect 5517 1744 5523 1777
rect 5300 1737 5308 1743
rect 5325 1724 5331 1736
rect 5389 1584 5395 1736
rect 5277 1537 5299 1543
rect 5293 1383 5299 1537
rect 5325 1384 5331 1476
rect 5293 1377 5308 1383
rect 5261 1344 5267 1356
rect 5277 1324 5283 1336
rect 5261 1064 5267 1096
rect 5277 1064 5283 1076
rect 5245 1023 5251 1036
rect 5245 1017 5267 1023
rect 5245 984 5251 996
rect 5261 944 5267 1017
rect 5133 684 5139 696
rect 5133 584 5139 616
rect 5149 544 5155 696
rect 5165 604 5171 876
rect 5181 844 5187 936
rect 5197 844 5203 916
rect 5277 884 5283 896
rect 5181 724 5187 836
rect 5197 724 5203 736
rect 5293 724 5299 1377
rect 5309 1304 5315 1356
rect 5325 1324 5331 1336
rect 5341 1304 5347 1376
rect 5357 1223 5363 1576
rect 5389 1363 5395 1436
rect 5405 1384 5411 1696
rect 5453 1623 5459 1636
rect 5437 1617 5459 1623
rect 5421 1524 5427 1536
rect 5437 1504 5443 1617
rect 5533 1604 5539 1696
rect 5517 1484 5523 1516
rect 5533 1504 5539 1516
rect 5437 1477 5452 1483
rect 5437 1384 5443 1477
rect 5389 1357 5411 1363
rect 5405 1344 5411 1357
rect 5389 1284 5395 1336
rect 5405 1304 5411 1336
rect 5341 1217 5363 1223
rect 5325 1084 5331 1156
rect 5341 1124 5347 1217
rect 5389 1184 5395 1196
rect 5421 1124 5427 1136
rect 5453 1044 5459 1056
rect 5309 837 5324 843
rect 5309 703 5315 837
rect 5341 823 5347 1016
rect 5357 943 5363 976
rect 5373 964 5379 1036
rect 5437 984 5443 996
rect 5357 937 5372 943
rect 5389 924 5395 936
rect 5405 904 5411 916
rect 5325 817 5347 823
rect 5325 784 5331 817
rect 5357 724 5363 736
rect 5309 697 5331 703
rect 5165 584 5171 596
rect 5181 544 5187 676
rect 5300 557 5308 563
rect 5284 537 5292 543
rect 5325 543 5331 697
rect 5373 684 5379 736
rect 5357 544 5363 676
rect 5389 664 5395 676
rect 5405 644 5411 716
rect 5373 564 5379 576
rect 5389 564 5395 596
rect 5309 537 5331 543
rect 5341 537 5356 543
rect 5181 524 5187 536
rect 5117 303 5123 456
rect 5261 384 5267 496
rect 5101 297 5123 303
rect 5037 284 5043 296
rect 4877 264 4883 276
rect 5060 257 5075 263
rect 4797 184 4803 216
rect 4925 164 4931 256
rect 5069 244 5075 257
rect 4941 224 4947 236
rect 5053 184 5059 196
rect 5069 184 5075 216
rect 4909 144 4915 156
rect 4701 137 4716 143
rect 4605 124 4611 136
rect 4669 124 4675 136
rect 4692 117 4700 123
rect 4541 104 4547 116
rect 4589 104 4595 116
rect 4765 104 4771 116
rect 5101 104 5107 297
rect 5165 284 5171 296
rect 5117 244 5123 276
rect 5188 257 5203 263
rect 5197 244 5203 257
rect 5117 144 5123 216
rect 5165 124 5171 156
rect 5181 144 5187 196
rect 5197 144 5203 216
rect 5213 104 5219 376
rect 5309 324 5315 537
rect 5341 324 5347 537
rect 5421 324 5427 556
rect 5437 464 5443 636
rect 5469 604 5475 716
rect 5501 584 5507 596
rect 5245 284 5251 296
rect 5309 284 5315 296
rect 5245 184 5251 216
rect 5261 144 5267 176
rect 5341 144 5347 276
rect 5357 184 5363 316
rect 5453 284 5459 496
rect 5469 484 5475 496
rect 5437 244 5443 276
rect 5453 244 5459 256
rect 5501 244 5507 256
rect 5437 184 5443 196
rect 5444 137 5452 143
rect 5517 124 5523 1036
rect 5565 384 5571 1436
rect 4308 97 4316 103
rect 3565 84 3571 96
rect 3693 84 3699 96
rect 3885 84 3891 96
rect 5277 84 5283 96
rect 5469 84 5475 96
rect 3853 44 3859 56
rect 3117 -43 3139 -37
rect 4701 -43 4707 16
<< m3contact >>
rect 1196 3996 1204 4004
rect 508 3976 516 3984
rect 604 3976 612 3984
rect 188 3956 196 3964
rect 860 3956 868 3964
rect 924 3956 932 3964
rect 1516 3936 1524 3944
rect 220 3916 228 3924
rect 268 3916 276 3924
rect 380 3916 388 3924
rect 1036 3916 1044 3924
rect 1436 3916 1444 3924
rect 1484 3916 1492 3924
rect 364 3896 372 3904
rect 140 3876 148 3884
rect 284 3876 292 3884
rect 300 3876 308 3884
rect 28 3856 36 3864
rect 12 3836 20 3844
rect 60 3756 68 3764
rect 108 3836 116 3844
rect 92 3736 100 3744
rect 12 3716 20 3724
rect 60 3696 68 3704
rect 28 3676 36 3684
rect 188 3796 196 3804
rect 108 3536 116 3544
rect 28 3476 36 3484
rect 76 3476 84 3484
rect 172 3476 180 3484
rect 204 3476 212 3484
rect 140 3396 148 3404
rect 172 3396 180 3404
rect 124 3376 132 3384
rect 124 3356 132 3364
rect 60 3316 68 3324
rect 60 3296 68 3304
rect 76 3196 84 3204
rect 252 3836 260 3844
rect 252 3776 260 3784
rect 684 3896 692 3904
rect 1228 3896 1236 3904
rect 1740 3996 1748 4004
rect 1612 3976 1620 3984
rect 1788 3976 1796 3984
rect 1596 3936 1604 3944
rect 1708 3936 1716 3944
rect 1580 3916 1588 3924
rect 1644 3916 1652 3924
rect 1772 3916 1780 3924
rect 524 3876 530 3884
rect 530 3876 532 3884
rect 572 3876 580 3884
rect 700 3876 708 3884
rect 748 3876 756 3884
rect 828 3876 836 3884
rect 860 3876 868 3884
rect 892 3876 900 3884
rect 988 3876 996 3884
rect 1020 3876 1022 3884
rect 1022 3876 1028 3884
rect 1068 3876 1076 3884
rect 1276 3876 1284 3884
rect 1340 3876 1348 3884
rect 1388 3876 1396 3884
rect 396 3836 404 3844
rect 412 3836 420 3844
rect 460 3836 468 3844
rect 588 3796 596 3804
rect 540 3776 548 3784
rect 572 3776 580 3784
rect 380 3756 388 3764
rect 332 3736 338 3744
rect 338 3736 340 3744
rect 364 3716 372 3724
rect 316 3696 324 3704
rect 300 3676 308 3684
rect 444 3736 452 3744
rect 492 3736 500 3744
rect 556 3716 564 3724
rect 700 3836 708 3844
rect 764 3836 772 3844
rect 780 3796 788 3804
rect 908 3856 916 3864
rect 988 3856 996 3864
rect 1212 3856 1220 3864
rect 1132 3816 1140 3824
rect 956 3796 964 3804
rect 1100 3796 1108 3804
rect 1292 3796 1300 3804
rect 1324 3796 1332 3804
rect 908 3776 916 3784
rect 1132 3776 1140 3784
rect 876 3756 884 3764
rect 908 3756 916 3764
rect 956 3756 964 3764
rect 620 3716 628 3724
rect 700 3716 708 3724
rect 396 3696 404 3704
rect 508 3696 516 3704
rect 604 3696 612 3704
rect 652 3696 660 3704
rect 460 3536 468 3544
rect 524 3536 532 3544
rect 604 3536 612 3544
rect 300 3516 308 3524
rect 380 3496 388 3504
rect 460 3496 468 3504
rect 252 3456 260 3464
rect 252 3356 260 3364
rect 220 3316 228 3324
rect 284 3316 292 3324
rect 60 3076 68 3084
rect 124 3076 132 3084
rect 124 2976 132 2984
rect 12 2956 20 2964
rect 140 2956 148 2964
rect 236 3096 244 3104
rect 252 3076 260 3084
rect 188 3056 196 3064
rect 204 3056 212 3064
rect 268 3056 276 3064
rect 188 2976 196 2984
rect 444 3476 452 3484
rect 332 3456 340 3464
rect 332 3376 340 3384
rect 380 3376 388 3384
rect 396 3356 404 3364
rect 444 3356 452 3364
rect 316 3336 324 3344
rect 300 3276 308 3284
rect 332 3116 340 3124
rect 316 3076 324 3084
rect 332 3076 340 3084
rect 300 3056 308 3064
rect 316 3056 324 3064
rect 316 3036 324 3044
rect 284 2976 292 2984
rect 236 2956 244 2964
rect 60 2936 68 2944
rect 156 2936 164 2944
rect 12 2896 20 2904
rect 28 2896 36 2904
rect 76 2896 84 2904
rect 12 2876 20 2884
rect 156 2916 164 2924
rect 108 2716 116 2724
rect 156 2716 164 2724
rect 92 2676 100 2684
rect 156 2676 164 2684
rect 108 2596 116 2604
rect 60 2556 68 2564
rect 124 2576 132 2584
rect 124 2536 132 2544
rect 172 2536 180 2544
rect 44 2516 52 2524
rect 12 2096 20 2104
rect 396 3336 404 3344
rect 492 3376 500 3384
rect 524 3336 532 3344
rect 572 3456 580 3464
rect 588 3436 596 3444
rect 668 3596 676 3604
rect 828 3716 836 3724
rect 1100 3736 1108 3744
rect 892 3716 900 3724
rect 1004 3716 1012 3724
rect 1532 3856 1540 3864
rect 1628 3816 1636 3824
rect 1468 3796 1476 3804
rect 1484 3796 1492 3804
rect 1548 3796 1556 3804
rect 1420 3776 1428 3784
rect 1596 3776 1604 3784
rect 1612 3776 1620 3784
rect 1628 3776 1636 3784
rect 1292 3736 1300 3744
rect 1340 3736 1348 3744
rect 1148 3716 1156 3724
rect 1148 3696 1156 3704
rect 812 3676 820 3684
rect 940 3676 948 3684
rect 972 3616 980 3624
rect 716 3576 724 3584
rect 748 3576 756 3584
rect 780 3536 788 3544
rect 844 3516 852 3524
rect 1068 3516 1076 3524
rect 988 3496 996 3504
rect 588 3376 596 3384
rect 636 3376 644 3384
rect 764 3436 772 3444
rect 748 3416 756 3424
rect 892 3436 900 3444
rect 812 3376 820 3384
rect 908 3376 916 3384
rect 748 3356 756 3364
rect 780 3356 788 3364
rect 892 3356 900 3364
rect 572 3336 580 3344
rect 636 3336 644 3344
rect 828 3336 836 3344
rect 412 3316 420 3324
rect 476 3316 484 3324
rect 812 3316 820 3324
rect 828 3296 836 3304
rect 892 3296 900 3304
rect 604 3276 612 3284
rect 396 3256 404 3264
rect 572 3256 580 3264
rect 380 3116 388 3124
rect 476 3136 484 3144
rect 524 3116 532 3124
rect 588 3116 596 3124
rect 396 3096 404 3104
rect 460 3096 468 3104
rect 428 3056 436 3064
rect 460 3056 468 3064
rect 348 3036 356 3044
rect 268 2936 276 2944
rect 412 2936 420 2944
rect 252 2896 260 2904
rect 284 2896 292 2904
rect 348 2896 356 2904
rect 508 3076 516 3084
rect 572 3036 580 3044
rect 588 2976 596 2984
rect 812 3276 820 3284
rect 700 3176 708 3184
rect 652 3156 660 3164
rect 620 3136 628 3144
rect 668 3136 676 3144
rect 828 3176 836 3184
rect 636 3116 644 3124
rect 716 3116 724 3124
rect 812 3116 820 3124
rect 908 3116 916 3124
rect 636 3036 644 3044
rect 764 3036 772 3044
rect 652 2976 660 2984
rect 732 2976 740 2984
rect 780 2976 788 2984
rect 604 2956 612 2964
rect 460 2936 468 2944
rect 476 2936 484 2944
rect 524 2936 532 2944
rect 588 2936 596 2944
rect 540 2916 548 2924
rect 652 2916 660 2924
rect 540 2896 548 2904
rect 332 2876 340 2884
rect 364 2876 372 2884
rect 444 2876 452 2884
rect 508 2876 516 2884
rect 332 2836 340 2844
rect 300 2776 308 2784
rect 364 2716 372 2724
rect 540 2776 548 2784
rect 492 2736 500 2744
rect 764 2796 772 2804
rect 812 2976 820 2984
rect 892 3036 900 3044
rect 828 2936 836 2944
rect 844 2796 852 2804
rect 652 2756 660 2764
rect 796 2756 804 2764
rect 844 2756 852 2764
rect 572 2716 580 2724
rect 636 2716 644 2724
rect 332 2696 340 2704
rect 412 2696 420 2704
rect 444 2696 452 2704
rect 284 2676 292 2684
rect 316 2676 324 2684
rect 252 2656 260 2664
rect 268 2636 276 2644
rect 268 2616 276 2624
rect 396 2636 404 2644
rect 460 2636 468 2644
rect 380 2616 388 2624
rect 316 2576 324 2584
rect 972 3436 980 3444
rect 972 3396 980 3404
rect 1036 3456 1044 3464
rect 1020 3396 1028 3404
rect 1036 3396 1044 3404
rect 1388 3696 1396 3704
rect 1260 3676 1268 3684
rect 1324 3656 1332 3664
rect 1196 3616 1204 3624
rect 1436 3696 1444 3704
rect 1468 3696 1476 3704
rect 1532 3696 1540 3704
rect 1404 3596 1412 3604
rect 1484 3596 1492 3604
rect 1356 3556 1364 3564
rect 1372 3516 1380 3524
rect 1132 3496 1140 3504
rect 1196 3496 1204 3504
rect 1100 3436 1108 3444
rect 1084 3416 1092 3424
rect 1132 3416 1140 3424
rect 1052 3376 1060 3384
rect 956 3316 964 3324
rect 988 3316 996 3324
rect 1052 3316 1060 3324
rect 1004 3256 1012 3264
rect 1084 3216 1092 3224
rect 1100 3196 1108 3204
rect 940 3156 948 3164
rect 956 3136 964 3144
rect 1020 3136 1028 3144
rect 988 3116 996 3124
rect 972 3076 980 3084
rect 940 3056 948 3064
rect 956 2936 964 2944
rect 956 2916 964 2924
rect 956 2876 964 2884
rect 956 2736 964 2744
rect 588 2696 596 2704
rect 604 2696 612 2704
rect 924 2696 932 2704
rect 940 2696 948 2704
rect 572 2676 580 2684
rect 652 2676 660 2684
rect 668 2676 676 2684
rect 716 2676 724 2684
rect 780 2676 788 2684
rect 524 2656 532 2664
rect 780 2656 788 2664
rect 796 2656 804 2664
rect 556 2616 564 2624
rect 508 2596 516 2604
rect 540 2596 548 2604
rect 316 2556 324 2564
rect 380 2556 388 2564
rect 444 2556 452 2564
rect 492 2556 500 2564
rect 252 2396 260 2404
rect 460 2536 468 2544
rect 508 2536 510 2544
rect 510 2536 516 2544
rect 332 2516 340 2524
rect 476 2516 484 2524
rect 364 2356 372 2364
rect 156 2336 164 2344
rect 348 2316 356 2324
rect 140 2276 148 2284
rect 156 2276 164 2284
rect 204 2276 212 2284
rect 76 2256 84 2264
rect 60 1936 68 1944
rect 44 1776 52 1784
rect 44 1756 52 1764
rect 108 2136 116 2144
rect 140 1896 148 1904
rect 140 1776 148 1784
rect 124 1736 132 1744
rect 108 1676 116 1684
rect 76 1616 84 1624
rect 108 1616 116 1624
rect 124 1476 132 1484
rect 60 1456 68 1464
rect 76 1356 84 1364
rect 108 1356 116 1364
rect 140 1356 148 1364
rect 188 2176 196 2184
rect 316 2176 324 2184
rect 300 2156 308 2164
rect 380 2296 388 2304
rect 492 2296 500 2304
rect 508 2296 516 2304
rect 1036 3096 1044 3104
rect 1116 3096 1124 3104
rect 1052 3056 1060 3064
rect 1132 3056 1140 3064
rect 1164 3056 1172 3064
rect 1084 2996 1092 3004
rect 1020 2976 1028 2984
rect 1036 2956 1044 2964
rect 1116 2936 1124 2944
rect 1164 2936 1172 2944
rect 1020 2916 1028 2924
rect 1020 2896 1028 2904
rect 1052 2876 1060 2884
rect 1004 2716 1012 2724
rect 1020 2716 1028 2724
rect 892 2636 900 2644
rect 940 2636 948 2644
rect 988 2636 996 2644
rect 908 2596 916 2604
rect 572 2576 580 2584
rect 828 2576 836 2584
rect 876 2576 884 2584
rect 892 2576 900 2584
rect 636 2556 644 2564
rect 700 2556 708 2564
rect 748 2556 756 2564
rect 764 2556 772 2564
rect 988 2556 996 2564
rect 652 2536 660 2544
rect 668 2536 676 2544
rect 764 2536 772 2544
rect 892 2536 900 2544
rect 972 2536 980 2544
rect 588 2496 596 2504
rect 716 2396 724 2404
rect 636 2376 644 2384
rect 716 2376 724 2384
rect 540 2356 548 2364
rect 620 2356 628 2364
rect 588 2316 596 2324
rect 572 2296 580 2304
rect 412 2256 420 2264
rect 460 2256 468 2264
rect 508 2176 516 2184
rect 252 2116 260 2124
rect 236 2096 244 2104
rect 220 2076 228 2084
rect 348 2136 356 2144
rect 444 2136 452 2144
rect 492 2136 500 2144
rect 524 2136 532 2144
rect 764 2336 772 2344
rect 796 2336 804 2344
rect 700 2316 708 2324
rect 732 2316 740 2324
rect 700 2296 708 2304
rect 876 2516 884 2524
rect 908 2516 916 2524
rect 956 2516 964 2524
rect 940 2496 948 2504
rect 892 2396 900 2404
rect 908 2356 916 2364
rect 812 2316 820 2324
rect 924 2316 932 2324
rect 780 2256 788 2264
rect 620 2216 628 2224
rect 604 2196 612 2204
rect 572 2176 580 2184
rect 812 2236 820 2244
rect 636 2196 644 2204
rect 652 2176 660 2184
rect 732 2176 740 2184
rect 716 2156 724 2164
rect 668 2136 676 2144
rect 700 2136 702 2144
rect 702 2136 708 2144
rect 460 2096 468 2104
rect 540 2096 548 2104
rect 652 2096 660 2104
rect 444 1916 452 1924
rect 492 1916 500 1924
rect 172 1876 180 1884
rect 204 1876 212 1884
rect 188 1756 196 1764
rect 204 1716 212 1724
rect 172 1496 180 1504
rect 204 1616 212 1624
rect 172 1476 180 1484
rect 188 1476 196 1484
rect 188 1456 196 1464
rect 348 1896 356 1904
rect 620 1896 628 1904
rect 716 2036 724 2044
rect 764 2156 772 2164
rect 908 2236 916 2244
rect 844 2216 852 2224
rect 844 2176 852 2184
rect 892 2176 900 2184
rect 860 2136 868 2144
rect 908 2136 916 2144
rect 956 2296 964 2304
rect 940 2276 948 2284
rect 956 2276 964 2284
rect 1020 2636 1028 2644
rect 1148 2856 1156 2864
rect 1164 2836 1172 2844
rect 1212 3396 1220 3404
rect 1244 3316 1252 3324
rect 1500 3556 1508 3564
rect 1276 3476 1284 3484
rect 1356 3476 1364 3484
rect 1452 3476 1460 3484
rect 1484 3476 1492 3484
rect 1340 3456 1348 3464
rect 1292 3416 1300 3424
rect 1404 3396 1412 3404
rect 1292 3376 1300 3384
rect 1436 3376 1444 3384
rect 1308 3356 1316 3364
rect 1356 3316 1364 3324
rect 1548 3556 1556 3564
rect 1660 3896 1668 3904
rect 1660 3796 1668 3804
rect 1724 3796 1732 3804
rect 1724 3776 1732 3784
rect 1676 3756 1684 3764
rect 1676 3736 1684 3744
rect 1644 3656 1652 3664
rect 1756 3676 1764 3684
rect 1756 3656 1764 3664
rect 1580 3536 1588 3544
rect 1676 3536 1684 3544
rect 1740 3536 1748 3544
rect 1804 3956 1812 3964
rect 1852 3956 1860 3964
rect 1852 3936 1860 3944
rect 1852 3916 1860 3924
rect 1916 3916 1924 3924
rect 1964 3916 1972 3924
rect 1900 3896 1908 3904
rect 2012 3976 2020 3984
rect 2028 3956 2036 3964
rect 2092 3956 2100 3964
rect 2012 3936 2020 3944
rect 1916 3876 1924 3884
rect 1964 3876 1972 3884
rect 1980 3876 1988 3884
rect 1852 3796 1860 3804
rect 1788 3776 1796 3784
rect 1868 3776 1876 3784
rect 1948 3776 1956 3784
rect 1804 3756 1812 3764
rect 1884 3756 1892 3764
rect 1900 3756 1908 3764
rect 1852 3736 1860 3744
rect 1820 3696 1828 3704
rect 1660 3496 1668 3504
rect 1580 3476 1588 3484
rect 1516 3456 1524 3464
rect 1468 3436 1476 3444
rect 1548 3436 1556 3444
rect 1548 3396 1556 3404
rect 1484 3376 1492 3384
rect 1532 3376 1540 3384
rect 1468 3316 1476 3324
rect 1516 3296 1524 3304
rect 1196 3276 1204 3284
rect 1260 3276 1268 3284
rect 1452 3276 1460 3284
rect 1340 3256 1348 3264
rect 1196 3236 1204 3244
rect 1212 3136 1220 3144
rect 1260 3136 1268 3144
rect 1596 3396 1604 3404
rect 1676 3456 1684 3464
rect 1820 3536 1828 3544
rect 1804 3496 1812 3504
rect 1820 3496 1828 3504
rect 1692 3436 1700 3444
rect 1660 3416 1668 3424
rect 1724 3416 1732 3424
rect 1772 3416 1780 3424
rect 1740 3396 1748 3404
rect 1612 3376 1620 3384
rect 1644 3376 1652 3384
rect 1804 3396 1812 3404
rect 1628 3336 1636 3344
rect 1676 3336 1684 3344
rect 1740 3336 1746 3344
rect 1746 3336 1748 3344
rect 1580 3216 1588 3224
rect 1532 3196 1540 3204
rect 1324 3136 1332 3144
rect 1372 3136 1380 3144
rect 1516 3116 1524 3124
rect 1580 3116 1588 3124
rect 1388 3096 1396 3104
rect 1452 3096 1460 3104
rect 1532 3096 1540 3104
rect 1692 3296 1700 3304
rect 1724 3196 1732 3204
rect 1884 3656 1892 3664
rect 1868 3496 1876 3504
rect 1852 3416 1860 3424
rect 1804 3336 1812 3344
rect 1836 3336 1844 3344
rect 1884 3316 1892 3324
rect 1740 3176 1748 3184
rect 1756 3176 1764 3184
rect 1788 3176 1796 3184
rect 1660 3116 1668 3124
rect 1612 3076 1620 3084
rect 1276 3056 1284 3064
rect 1308 3056 1316 3064
rect 1228 2996 1236 3004
rect 1260 2976 1268 2984
rect 1292 2956 1300 2964
rect 1212 2936 1220 2944
rect 1340 3036 1348 3044
rect 1564 3036 1572 3044
rect 1548 3016 1556 3024
rect 1484 2996 1492 3004
rect 1548 2996 1556 3004
rect 1500 2976 1508 2984
rect 1436 2956 1444 2964
rect 1628 3036 1636 3044
rect 1596 3016 1604 3024
rect 1644 3016 1652 3024
rect 1612 2976 1620 2984
rect 1356 2936 1364 2944
rect 1628 2936 1636 2944
rect 1340 2916 1348 2924
rect 1372 2896 1380 2904
rect 1276 2856 1284 2864
rect 1212 2796 1220 2804
rect 1260 2756 1268 2764
rect 1084 2696 1092 2704
rect 1116 2696 1124 2704
rect 1180 2696 1188 2704
rect 1324 2696 1332 2704
rect 1132 2676 1140 2684
rect 1228 2676 1234 2684
rect 1234 2676 1236 2684
rect 1068 2656 1076 2664
rect 1084 2656 1092 2664
rect 1148 2636 1156 2644
rect 1052 2596 1060 2604
rect 1500 2776 1508 2784
rect 1500 2756 1508 2764
rect 1436 2716 1444 2724
rect 1372 2696 1380 2704
rect 1564 2796 1572 2804
rect 1548 2716 1556 2724
rect 1628 2796 1636 2804
rect 1612 2756 1620 2764
rect 1484 2676 1492 2684
rect 1532 2676 1540 2684
rect 1564 2676 1572 2684
rect 1596 2676 1604 2684
rect 1180 2636 1188 2644
rect 1228 2636 1236 2644
rect 1276 2636 1284 2644
rect 1292 2636 1300 2644
rect 1340 2636 1348 2644
rect 1356 2636 1364 2644
rect 1036 2576 1044 2584
rect 1068 2576 1076 2584
rect 1164 2576 1172 2584
rect 1052 2556 1060 2564
rect 1020 2536 1022 2544
rect 1022 2536 1028 2544
rect 1068 2536 1076 2544
rect 1084 2536 1092 2544
rect 1148 2476 1156 2484
rect 1404 2596 1412 2604
rect 1356 2576 1364 2584
rect 1244 2556 1252 2564
rect 1260 2556 1268 2564
rect 1468 2636 1476 2644
rect 1468 2616 1476 2624
rect 1500 2596 1508 2604
rect 1308 2556 1316 2564
rect 1340 2556 1348 2564
rect 1388 2556 1396 2564
rect 1420 2556 1428 2564
rect 1244 2536 1252 2544
rect 1404 2536 1412 2544
rect 1452 2536 1460 2544
rect 1468 2536 1476 2544
rect 1388 2496 1396 2504
rect 1116 2436 1124 2444
rect 1164 2436 1172 2444
rect 1420 2416 1428 2424
rect 1100 2396 1108 2404
rect 1356 2396 1364 2404
rect 1036 2296 1044 2304
rect 1132 2296 1140 2304
rect 1004 2256 1012 2264
rect 972 2236 980 2244
rect 1068 2196 1076 2204
rect 1100 2196 1108 2204
rect 988 2176 996 2184
rect 1020 2176 1028 2184
rect 1084 2176 1092 2184
rect 1164 2216 1172 2224
rect 1148 2156 1156 2164
rect 1068 2116 1076 2124
rect 908 2076 916 2084
rect 1132 2076 1140 2084
rect 1148 2076 1156 2084
rect 748 2056 756 2064
rect 700 1956 708 1964
rect 732 1956 740 1964
rect 332 1876 340 1884
rect 508 1876 516 1884
rect 284 1856 292 1864
rect 396 1856 404 1864
rect 348 1816 356 1824
rect 380 1816 388 1824
rect 316 1776 324 1784
rect 332 1776 340 1784
rect 412 1796 420 1804
rect 300 1716 308 1724
rect 252 1696 260 1704
rect 380 1696 388 1704
rect 316 1476 324 1484
rect 188 1316 196 1324
rect 60 1216 68 1224
rect 44 1196 52 1204
rect 76 1196 84 1204
rect 28 1076 36 1084
rect 60 1036 68 1044
rect 140 1196 148 1204
rect 220 1336 228 1344
rect 204 1196 212 1204
rect 444 1776 452 1784
rect 460 1776 468 1784
rect 588 1856 596 1864
rect 556 1776 564 1784
rect 1100 2016 1108 2024
rect 844 1996 852 2004
rect 1164 1996 1172 2004
rect 828 1976 836 1984
rect 1196 2256 1204 2264
rect 1260 2256 1268 2264
rect 1276 2216 1284 2224
rect 1260 2196 1268 2204
rect 1212 2176 1220 2184
rect 1228 2156 1236 2164
rect 1228 2096 1236 2104
rect 1244 2076 1252 2084
rect 1196 1996 1204 2004
rect 796 1956 804 1964
rect 1180 1956 1188 1964
rect 1068 1936 1076 1944
rect 860 1896 868 1904
rect 876 1896 884 1904
rect 748 1856 756 1864
rect 668 1836 676 1844
rect 684 1836 692 1844
rect 716 1836 724 1844
rect 764 1836 772 1844
rect 844 1776 852 1784
rect 572 1756 580 1764
rect 668 1756 676 1764
rect 684 1756 692 1764
rect 828 1756 836 1764
rect 524 1736 532 1744
rect 572 1716 580 1724
rect 620 1716 628 1724
rect 508 1696 516 1704
rect 540 1696 548 1704
rect 396 1516 404 1524
rect 316 1376 324 1384
rect 364 1376 372 1384
rect 332 1336 338 1344
rect 338 1336 340 1344
rect 268 1316 276 1324
rect 380 1276 388 1284
rect 236 1156 244 1164
rect 252 1156 260 1164
rect 284 1156 292 1164
rect 268 1116 276 1124
rect 348 1116 356 1124
rect 172 1096 180 1104
rect 220 1096 228 1104
rect 204 1076 212 1084
rect 140 1056 148 1064
rect 172 1056 180 1064
rect 188 1016 196 1024
rect 108 996 116 1004
rect 140 996 148 1004
rect 140 956 148 964
rect 172 936 180 944
rect 172 876 180 884
rect 60 816 68 824
rect 12 796 20 804
rect 44 796 52 804
rect 188 716 196 724
rect 204 696 212 704
rect 300 1056 308 1064
rect 316 1036 324 1044
rect 236 1016 244 1024
rect 332 1016 340 1024
rect 380 976 388 984
rect 252 956 260 964
rect 300 956 308 964
rect 620 1536 628 1544
rect 460 1496 468 1504
rect 588 1496 596 1504
rect 492 1456 500 1464
rect 588 1456 596 1464
rect 444 1356 452 1364
rect 508 1356 516 1364
rect 572 1356 580 1364
rect 636 1496 644 1504
rect 732 1716 740 1724
rect 780 1716 788 1724
rect 716 1596 724 1604
rect 764 1556 772 1564
rect 700 1496 708 1504
rect 828 1536 836 1544
rect 828 1496 836 1504
rect 716 1476 722 1484
rect 722 1476 724 1484
rect 636 1456 644 1464
rect 764 1456 772 1464
rect 636 1436 644 1444
rect 780 1436 788 1444
rect 844 1416 852 1424
rect 700 1376 708 1384
rect 780 1376 788 1384
rect 716 1356 724 1364
rect 844 1356 852 1364
rect 428 1336 436 1344
rect 540 1336 548 1344
rect 764 1336 772 1344
rect 828 1336 836 1344
rect 476 1316 484 1324
rect 540 1316 548 1324
rect 460 1276 468 1284
rect 524 1136 532 1144
rect 444 1116 452 1124
rect 460 1056 468 1064
rect 508 1036 516 1044
rect 444 976 452 984
rect 396 956 404 964
rect 412 956 420 964
rect 380 916 388 924
rect 284 896 292 904
rect 364 896 372 904
rect 252 776 260 784
rect 444 936 452 944
rect 492 936 500 944
rect 412 876 420 884
rect 428 876 436 884
rect 396 836 404 844
rect 396 796 404 804
rect 428 736 436 744
rect 284 716 292 724
rect 332 716 340 724
rect 460 876 468 884
rect 524 876 532 884
rect 492 836 500 844
rect 460 756 468 764
rect 476 736 484 744
rect 268 696 276 704
rect 188 676 196 684
rect 220 676 228 684
rect 252 676 260 684
rect 44 656 52 664
rect 124 656 132 664
rect 204 656 212 664
rect 268 656 276 664
rect 92 596 100 604
rect 108 596 116 604
rect 140 596 148 604
rect 60 576 68 584
rect 12 496 20 504
rect 28 316 36 324
rect 124 536 132 544
rect 252 556 260 564
rect 316 636 324 644
rect 348 636 356 644
rect 460 636 468 644
rect 316 616 324 624
rect 348 536 356 544
rect 636 1276 644 1284
rect 556 1156 564 1164
rect 572 976 580 984
rect 556 956 564 964
rect 588 956 596 964
rect 588 876 596 884
rect 556 776 564 784
rect 588 716 596 724
rect 620 1136 628 1144
rect 636 1016 644 1024
rect 748 1296 756 1304
rect 828 1276 836 1284
rect 812 1256 820 1264
rect 780 1176 788 1184
rect 748 1136 756 1144
rect 1004 1916 1012 1924
rect 924 1896 932 1904
rect 956 1896 964 1904
rect 1020 1896 1028 1904
rect 908 1856 916 1864
rect 972 1856 980 1864
rect 972 1836 980 1844
rect 1036 1836 1044 1844
rect 1068 1856 1076 1864
rect 1084 1856 1092 1864
rect 1116 1836 1124 1844
rect 1164 1836 1172 1844
rect 908 1776 916 1784
rect 956 1776 964 1784
rect 1004 1776 1012 1784
rect 1020 1776 1028 1784
rect 1164 1776 1172 1784
rect 892 1756 900 1764
rect 876 1696 884 1704
rect 876 1476 884 1484
rect 892 1436 900 1444
rect 908 1276 916 1284
rect 1180 1756 1188 1764
rect 956 1696 964 1704
rect 1036 1556 1044 1564
rect 1004 1536 1012 1544
rect 1020 1516 1028 1524
rect 940 1456 948 1464
rect 972 1456 980 1464
rect 972 1436 980 1444
rect 972 1396 980 1404
rect 956 1356 964 1364
rect 940 1296 948 1304
rect 956 1196 964 1204
rect 764 1076 772 1084
rect 860 1076 868 1084
rect 748 1056 756 1064
rect 700 1016 708 1024
rect 716 1016 724 1024
rect 828 1036 836 1044
rect 828 1016 836 1024
rect 844 1016 852 1024
rect 764 996 772 1004
rect 812 996 820 1004
rect 796 956 804 964
rect 636 936 644 944
rect 684 936 692 944
rect 700 936 708 944
rect 700 816 708 824
rect 684 756 692 764
rect 780 776 788 784
rect 844 996 852 1004
rect 972 1096 980 1104
rect 940 1056 948 1064
rect 956 1016 964 1024
rect 1020 1396 1028 1404
rect 1004 1376 1012 1384
rect 1068 1536 1076 1544
rect 1132 1696 1140 1704
rect 1132 1676 1140 1684
rect 1100 1656 1108 1664
rect 1148 1636 1156 1644
rect 1116 1536 1124 1544
rect 1164 1536 1172 1544
rect 1244 1856 1252 1864
rect 1228 1836 1236 1844
rect 1196 1636 1204 1644
rect 1244 1596 1252 1604
rect 1196 1536 1204 1544
rect 1228 1536 1236 1544
rect 1228 1516 1236 1524
rect 1244 1516 1252 1524
rect 1180 1496 1188 1504
rect 1212 1496 1220 1504
rect 1084 1476 1092 1484
rect 1148 1476 1150 1484
rect 1150 1476 1156 1484
rect 1100 1456 1108 1464
rect 1132 1456 1140 1464
rect 1116 1436 1124 1444
rect 1100 1416 1108 1424
rect 1084 1376 1092 1384
rect 1052 1356 1060 1364
rect 1068 1356 1076 1364
rect 1036 1276 1044 1284
rect 1036 1256 1044 1264
rect 1100 1336 1108 1344
rect 1084 1216 1092 1224
rect 1084 1196 1092 1204
rect 1068 1136 1076 1144
rect 1004 1116 1012 1124
rect 988 996 996 1004
rect 1244 1436 1252 1444
rect 1212 1376 1220 1384
rect 1148 1336 1156 1344
rect 1180 1336 1188 1344
rect 1292 2196 1300 2204
rect 1276 2176 1284 2184
rect 1436 2276 1444 2284
rect 1340 2256 1348 2264
rect 1356 2236 1364 2244
rect 1420 2236 1428 2244
rect 1404 2196 1412 2204
rect 1484 2476 1492 2484
rect 1516 2536 1524 2544
rect 1532 2536 1540 2544
rect 1484 2316 1492 2324
rect 1596 2576 1604 2584
rect 1724 2976 1732 2984
rect 1676 2936 1682 2944
rect 1682 2936 1684 2944
rect 1740 2796 1748 2804
rect 1660 2756 1668 2764
rect 1868 3156 1876 3164
rect 1836 3136 1844 3144
rect 1788 3116 1796 3124
rect 1788 3096 1796 3104
rect 1772 3036 1780 3044
rect 1772 2996 1780 3004
rect 1852 3076 1860 3084
rect 1996 3856 2004 3864
rect 2092 3936 2100 3944
rect 2156 3936 2164 3944
rect 2380 3956 2388 3964
rect 2316 3916 2324 3924
rect 2284 3896 2292 3904
rect 2108 3876 2116 3884
rect 2188 3876 2196 3884
rect 2364 3896 2372 3904
rect 2172 3856 2180 3864
rect 2284 3856 2292 3864
rect 2428 3916 2436 3924
rect 2508 3936 2516 3944
rect 2396 3896 2404 3904
rect 2460 3896 2468 3904
rect 2396 3876 2404 3884
rect 2460 3876 2468 3884
rect 2252 3836 2260 3844
rect 2284 3836 2292 3844
rect 2332 3836 2340 3844
rect 2044 3816 2052 3824
rect 2172 3796 2180 3804
rect 2236 3796 2244 3804
rect 2108 3716 2116 3724
rect 2124 3716 2132 3724
rect 2044 3696 2052 3704
rect 2028 3636 2036 3644
rect 1996 3596 2004 3604
rect 1980 3576 1988 3584
rect 1964 3536 1972 3544
rect 1980 3496 1988 3504
rect 2092 3676 2100 3684
rect 2076 3536 2084 3544
rect 1916 3436 1924 3444
rect 2028 3416 2036 3424
rect 1932 3396 1940 3404
rect 1996 3396 2004 3404
rect 1932 3376 1940 3384
rect 1964 3316 1972 3324
rect 1916 3236 1924 3244
rect 1932 3196 1940 3204
rect 2060 3316 2068 3324
rect 2124 3656 2132 3664
rect 2108 3596 2116 3604
rect 2188 3696 2196 3704
rect 2204 3696 2212 3704
rect 2252 3696 2260 3704
rect 2156 3556 2164 3564
rect 2188 3656 2196 3664
rect 2380 3816 2388 3824
rect 2444 3856 2452 3864
rect 2428 3816 2436 3824
rect 2396 3796 2404 3804
rect 2444 3796 2452 3804
rect 2316 3756 2324 3764
rect 2428 3756 2436 3764
rect 2300 3736 2308 3744
rect 2348 3736 2356 3744
rect 2364 3716 2372 3724
rect 2428 3716 2436 3724
rect 2284 3536 2292 3544
rect 2252 3516 2260 3524
rect 2300 3516 2308 3524
rect 2348 3516 2356 3524
rect 2124 3456 2132 3464
rect 2172 3456 2180 3464
rect 2124 3396 2132 3404
rect 2108 3376 2116 3384
rect 2108 3336 2116 3344
rect 2156 3316 2164 3324
rect 1980 3196 1988 3204
rect 1996 3196 2004 3204
rect 1980 3156 1988 3164
rect 2076 3096 2084 3104
rect 1884 3056 1892 3064
rect 1868 2996 1876 3004
rect 1852 2976 1860 2984
rect 1788 2936 1796 2944
rect 1836 2936 1844 2944
rect 1804 2916 1812 2924
rect 1804 2796 1812 2804
rect 1804 2756 1812 2764
rect 1836 2756 1844 2764
rect 1772 2736 1780 2744
rect 1820 2736 1828 2744
rect 1820 2696 1828 2704
rect 1644 2676 1652 2684
rect 1692 2676 1700 2684
rect 1756 2676 1764 2684
rect 1788 2676 1796 2684
rect 1660 2656 1668 2664
rect 1676 2636 1684 2644
rect 1788 2596 1796 2604
rect 1852 2596 1860 2604
rect 1868 2596 1876 2604
rect 1852 2556 1860 2564
rect 1628 2536 1636 2544
rect 1804 2536 1812 2544
rect 1676 2496 1684 2504
rect 1596 2436 1604 2444
rect 1708 2376 1716 2384
rect 1660 2356 1668 2364
rect 1548 2276 1556 2284
rect 1644 2276 1652 2284
rect 1660 2276 1668 2284
rect 1724 2276 1732 2284
rect 1452 2236 1460 2244
rect 1468 2236 1476 2244
rect 1548 2236 1556 2244
rect 1660 2236 1668 2244
rect 1436 2216 1444 2224
rect 1596 2216 1604 2224
rect 1740 2236 1748 2244
rect 1580 2196 1588 2204
rect 1468 2156 1476 2164
rect 1548 2156 1556 2164
rect 1660 2196 1668 2204
rect 1724 2176 1732 2184
rect 1596 2136 1604 2144
rect 1612 2136 1620 2144
rect 1724 2136 1732 2144
rect 1292 2096 1300 2104
rect 1340 2096 1348 2104
rect 1324 2076 1332 2084
rect 1452 2096 1460 2104
rect 1580 2096 1588 2104
rect 1388 2056 1396 2064
rect 1388 2036 1396 2044
rect 1356 1916 1364 1924
rect 1276 1856 1284 1864
rect 1548 1996 1556 2004
rect 1484 1956 1492 1964
rect 1644 2016 1652 2024
rect 1612 1976 1620 1984
rect 1724 1956 1732 1964
rect 1660 1916 1668 1924
rect 1372 1856 1380 1864
rect 1452 1856 1460 1864
rect 1484 1856 1492 1864
rect 1324 1816 1332 1824
rect 1340 1796 1348 1804
rect 1404 1816 1412 1824
rect 1500 1796 1508 1804
rect 1452 1776 1460 1784
rect 1484 1776 1492 1784
rect 1404 1736 1412 1744
rect 1276 1496 1284 1504
rect 1324 1496 1332 1504
rect 1292 1456 1300 1464
rect 1308 1456 1316 1464
rect 1340 1456 1348 1464
rect 1372 1456 1380 1464
rect 1260 1376 1268 1384
rect 1292 1336 1300 1344
rect 1452 1676 1460 1684
rect 1404 1636 1412 1644
rect 1420 1536 1428 1544
rect 1564 1856 1572 1864
rect 1596 1856 1604 1864
rect 1532 1796 1540 1804
rect 1548 1776 1556 1784
rect 1596 1796 1604 1804
rect 1612 1796 1620 1804
rect 1580 1716 1588 1724
rect 1564 1636 1572 1644
rect 1516 1596 1524 1604
rect 1548 1596 1556 1604
rect 1580 1556 1588 1564
rect 1580 1536 1588 1544
rect 1452 1496 1460 1504
rect 1484 1496 1492 1504
rect 1612 1716 1620 1724
rect 1772 2356 1780 2364
rect 1788 2356 1796 2364
rect 1868 2436 1876 2444
rect 1932 3076 1940 3084
rect 1964 3076 1972 3084
rect 1964 3056 1972 3064
rect 2028 3056 2036 3064
rect 2076 3056 2084 3064
rect 1980 3036 1988 3044
rect 2012 3036 2020 3044
rect 1948 2996 1956 3004
rect 1900 2976 1908 2984
rect 1932 2956 1940 2964
rect 1916 2896 1924 2904
rect 2060 3036 2068 3044
rect 2044 2996 2052 3004
rect 2060 2976 2068 2984
rect 2076 2936 2084 2944
rect 1900 2876 1908 2884
rect 1980 2876 1988 2884
rect 2044 2796 2052 2804
rect 2044 2776 2052 2784
rect 1900 2756 1908 2764
rect 2124 3136 2132 3144
rect 2108 3116 2116 3124
rect 2108 2896 2116 2904
rect 2108 2756 2116 2764
rect 1932 2696 1940 2704
rect 1948 2696 1956 2704
rect 2012 2696 2020 2704
rect 2092 2696 2100 2704
rect 1916 2636 1924 2644
rect 1916 2596 1924 2604
rect 1900 2536 1908 2544
rect 1964 2656 1972 2664
rect 1996 2656 2004 2664
rect 1980 2636 1988 2644
rect 2188 3136 2196 3144
rect 2156 3116 2164 3124
rect 2188 3096 2196 3104
rect 2252 3396 2260 3404
rect 2252 3376 2260 3384
rect 2428 3676 2436 3684
rect 2380 3496 2388 3504
rect 2556 3916 2564 3924
rect 2684 3976 2692 3984
rect 3292 3956 3300 3964
rect 4300 3956 4308 3964
rect 4764 3956 4772 3964
rect 2652 3936 2660 3944
rect 2700 3936 2708 3944
rect 2636 3876 2644 3884
rect 2492 3796 2500 3804
rect 2572 3856 2580 3864
rect 2556 3836 2564 3844
rect 2588 3836 2596 3844
rect 2828 3916 2836 3924
rect 3132 3916 3140 3924
rect 3180 3916 3188 3924
rect 3276 3916 3284 3924
rect 2716 3896 2724 3904
rect 2764 3876 2770 3884
rect 2770 3876 2772 3884
rect 2972 3896 2980 3904
rect 3004 3896 3012 3904
rect 3084 3896 3092 3904
rect 3148 3896 3156 3904
rect 3196 3896 3204 3904
rect 3260 3896 3268 3904
rect 2956 3876 2964 3884
rect 2748 3856 2756 3864
rect 2796 3856 2804 3864
rect 2828 3856 2836 3864
rect 2524 3776 2532 3784
rect 2588 3816 2596 3824
rect 2620 3796 2628 3804
rect 2652 3796 2660 3804
rect 2588 3776 2596 3784
rect 2572 3756 2580 3764
rect 2492 3736 2500 3744
rect 2492 3716 2500 3724
rect 2492 3696 2500 3704
rect 2540 3696 2548 3704
rect 2460 3676 2468 3684
rect 2460 3516 2468 3524
rect 2316 3476 2324 3484
rect 2300 3456 2308 3464
rect 2316 3396 2324 3404
rect 2444 3376 2452 3384
rect 2300 3316 2308 3324
rect 2284 3296 2292 3304
rect 2364 3216 2372 3224
rect 2524 3676 2532 3684
rect 2556 3556 2564 3564
rect 2620 3716 2628 3724
rect 2812 3796 2820 3804
rect 2700 3756 2708 3764
rect 2860 3796 2868 3804
rect 2764 3756 2772 3764
rect 2844 3756 2852 3764
rect 2892 3796 2900 3804
rect 2876 3776 2884 3784
rect 2956 3836 2964 3844
rect 3020 3856 3028 3864
rect 3068 3856 3076 3864
rect 3036 3836 3044 3844
rect 3084 3836 3092 3844
rect 3100 3836 3108 3844
rect 2972 3796 2980 3804
rect 2876 3756 2884 3764
rect 2908 3756 2916 3764
rect 2972 3756 2980 3764
rect 2988 3756 2996 3764
rect 2908 3736 2916 3744
rect 2940 3736 2942 3744
rect 2942 3736 2948 3744
rect 2780 3716 2788 3724
rect 2812 3716 2820 3724
rect 3100 3756 3108 3764
rect 3164 3756 3172 3764
rect 3212 3756 3220 3764
rect 3052 3736 3060 3744
rect 3020 3696 3028 3704
rect 2700 3636 2708 3644
rect 2652 3596 2660 3604
rect 2636 3556 2644 3564
rect 2764 3596 2772 3604
rect 2748 3516 2756 3524
rect 2492 3416 2500 3424
rect 2620 3436 2628 3444
rect 2700 3436 2708 3444
rect 2620 3376 2628 3384
rect 2556 3356 2564 3364
rect 2796 3516 2804 3524
rect 2812 3516 2820 3524
rect 2972 3556 2980 3564
rect 2940 3536 2948 3544
rect 2828 3496 2836 3504
rect 2828 3476 2836 3484
rect 2892 3476 2898 3484
rect 2898 3476 2900 3484
rect 2764 3456 2772 3464
rect 2828 3456 2836 3464
rect 2716 3396 2724 3404
rect 3036 3556 3044 3564
rect 3004 3516 3012 3524
rect 3004 3476 3006 3484
rect 3006 3476 3012 3484
rect 2956 3456 2964 3464
rect 2972 3456 2980 3464
rect 3036 3456 3044 3464
rect 2924 3436 2932 3444
rect 2876 3416 2884 3424
rect 2972 3376 2980 3384
rect 2924 3356 2932 3364
rect 3020 3356 3028 3364
rect 2540 3336 2548 3344
rect 2684 3336 2692 3344
rect 2700 3336 2708 3344
rect 2748 3336 2750 3344
rect 2750 3336 2756 3344
rect 2812 3336 2820 3344
rect 2844 3336 2852 3344
rect 2956 3336 2964 3344
rect 2620 3316 2628 3324
rect 2684 3316 2692 3324
rect 2476 3296 2484 3304
rect 2572 3296 2580 3304
rect 2668 3296 2676 3304
rect 2364 3176 2372 3184
rect 2428 3176 2436 3184
rect 2444 3116 2452 3124
rect 2460 3116 2468 3124
rect 2668 3116 2676 3124
rect 2220 3056 2228 3064
rect 2188 3036 2196 3044
rect 2172 2996 2180 3004
rect 2252 2996 2260 3004
rect 2172 2976 2180 2984
rect 2236 2976 2244 2984
rect 2380 3076 2388 3084
rect 2316 3036 2324 3044
rect 2364 2996 2372 3004
rect 2300 2976 2308 2984
rect 2332 2976 2340 2984
rect 2556 3096 2564 3104
rect 2620 3096 2628 3104
rect 2700 3096 2708 3104
rect 2508 3056 2516 3064
rect 2604 3056 2612 3064
rect 2684 3056 2692 3064
rect 2428 2996 2436 3004
rect 2428 2976 2436 2984
rect 2348 2956 2356 2964
rect 2396 2956 2404 2964
rect 2444 2956 2452 2964
rect 2636 3016 2644 3024
rect 2204 2936 2212 2944
rect 2236 2936 2244 2944
rect 2268 2936 2276 2944
rect 2156 2876 2164 2884
rect 2156 2856 2164 2864
rect 2140 2756 2148 2764
rect 2684 2976 2692 2984
rect 2380 2936 2388 2944
rect 2300 2896 2308 2904
rect 2396 2896 2404 2904
rect 2204 2716 2212 2724
rect 2252 2876 2260 2884
rect 2316 2836 2324 2844
rect 2332 2736 2340 2744
rect 2236 2716 2244 2724
rect 2188 2656 2196 2664
rect 2044 2576 2052 2584
rect 2140 2636 2148 2644
rect 2076 2536 2084 2544
rect 2076 2516 2084 2524
rect 2028 2436 2036 2444
rect 1916 2376 1924 2384
rect 1916 2356 1924 2364
rect 2124 2396 2132 2404
rect 1964 2376 1972 2384
rect 2124 2376 2132 2384
rect 1884 2336 1892 2344
rect 1932 2336 1940 2344
rect 1948 2336 1956 2344
rect 1836 2296 1844 2304
rect 1804 2276 1812 2284
rect 1868 2276 1876 2284
rect 1852 2236 1860 2244
rect 1836 2176 1844 2184
rect 1788 2116 1796 2124
rect 1788 2096 1796 2104
rect 1772 2076 1780 2084
rect 1868 2016 1876 2024
rect 1836 1956 1844 1964
rect 1820 1936 1828 1944
rect 1676 1876 1684 1884
rect 1804 1876 1812 1884
rect 1676 1856 1684 1864
rect 1740 1856 1748 1864
rect 1788 1816 1796 1824
rect 1740 1796 1748 1804
rect 1660 1776 1668 1784
rect 1788 1776 1796 1784
rect 1708 1716 1716 1724
rect 1724 1716 1732 1724
rect 1852 1916 1860 1924
rect 1948 2256 1956 2264
rect 1932 2236 1940 2244
rect 1916 2156 1924 2164
rect 1932 2096 1940 2104
rect 1884 1856 1892 1864
rect 1852 1776 1860 1784
rect 1852 1736 1860 1744
rect 1868 1716 1876 1724
rect 1884 1716 1892 1724
rect 1644 1696 1652 1704
rect 1836 1676 1844 1684
rect 1836 1636 1844 1644
rect 1676 1596 1684 1604
rect 1660 1556 1668 1564
rect 1628 1516 1636 1524
rect 1740 1516 1748 1524
rect 1804 1516 1812 1524
rect 1628 1496 1636 1504
rect 1468 1476 1476 1484
rect 1516 1476 1524 1484
rect 1580 1476 1588 1484
rect 1596 1476 1604 1484
rect 1708 1476 1716 1484
rect 1772 1476 1780 1484
rect 1388 1416 1396 1424
rect 1532 1416 1540 1424
rect 1596 1416 1604 1424
rect 1628 1416 1636 1424
rect 1724 1416 1732 1424
rect 1356 1396 1364 1404
rect 1548 1396 1556 1404
rect 1420 1376 1428 1384
rect 1484 1376 1492 1384
rect 1516 1376 1524 1384
rect 1228 1276 1236 1284
rect 1148 1236 1156 1244
rect 1340 1256 1348 1264
rect 1388 1336 1396 1344
rect 1612 1356 1620 1364
rect 1884 1656 1892 1664
rect 2076 2356 2084 2364
rect 1980 2336 1988 2344
rect 2188 2336 2196 2344
rect 2060 2276 2068 2284
rect 2188 2256 2196 2264
rect 1980 2236 1988 2244
rect 2028 2236 2036 2244
rect 2060 2236 2068 2244
rect 2156 2236 2164 2244
rect 2172 2236 2180 2244
rect 1980 2176 1988 2184
rect 1996 2116 2004 2124
rect 2012 2116 2020 2124
rect 1964 1916 1972 1924
rect 1996 1856 2004 1864
rect 1980 1796 1988 1804
rect 1948 1776 1956 1784
rect 1948 1736 1956 1744
rect 2108 2176 2116 2184
rect 2060 2156 2068 2164
rect 2124 2136 2132 2144
rect 2044 1956 2052 1964
rect 2140 1956 2148 1964
rect 2188 1956 2196 1964
rect 2076 1916 2084 1924
rect 2044 1856 2052 1864
rect 2060 1816 2068 1824
rect 2140 1816 2148 1824
rect 2060 1796 2068 1804
rect 2316 2676 2324 2684
rect 2380 2676 2388 2684
rect 2284 2596 2292 2604
rect 2316 2596 2324 2604
rect 2252 2576 2260 2584
rect 2300 2576 2308 2584
rect 2764 3316 2772 3324
rect 3036 3316 3044 3324
rect 2844 3276 2852 3284
rect 2812 3136 2820 3144
rect 2732 3096 2740 3104
rect 2876 3276 2884 3284
rect 2860 3256 2868 3264
rect 2892 3156 2900 3164
rect 2940 3156 2948 3164
rect 2892 3136 2900 3144
rect 2972 3136 2980 3144
rect 2780 3076 2788 3084
rect 2748 3056 2756 3064
rect 2764 3056 2772 3064
rect 2732 3036 2740 3044
rect 2764 2976 2772 2984
rect 2732 2936 2740 2944
rect 2636 2916 2644 2924
rect 2716 2916 2724 2924
rect 2748 2896 2756 2904
rect 2460 2876 2468 2884
rect 2444 2796 2452 2804
rect 2620 2796 2628 2804
rect 2700 2876 2708 2884
rect 2652 2756 2660 2764
rect 2652 2736 2660 2744
rect 2428 2716 2436 2724
rect 2460 2716 2468 2724
rect 2828 3016 2836 3024
rect 2812 2896 2820 2904
rect 2796 2876 2804 2884
rect 2860 3016 2868 3024
rect 2972 3056 2980 3064
rect 2892 2956 2900 2964
rect 2924 2916 2932 2924
rect 2892 2896 2900 2904
rect 2844 2796 2852 2804
rect 2956 2816 2964 2824
rect 2940 2756 2948 2764
rect 2828 2736 2836 2744
rect 2924 2736 2932 2744
rect 2844 2716 2852 2724
rect 2892 2716 2900 2724
rect 2940 2716 2948 2724
rect 2492 2696 2500 2704
rect 2780 2696 2788 2704
rect 2444 2676 2452 2684
rect 2508 2676 2516 2684
rect 2572 2676 2580 2684
rect 2636 2676 2644 2684
rect 2764 2676 2772 2684
rect 2732 2656 2740 2664
rect 2796 2656 2804 2664
rect 2508 2596 2516 2604
rect 2556 2596 2564 2604
rect 2492 2576 2500 2584
rect 2332 2556 2340 2564
rect 2476 2556 2484 2564
rect 2508 2556 2516 2564
rect 2236 2536 2244 2544
rect 2300 2536 2302 2544
rect 2302 2536 2308 2544
rect 2252 2496 2260 2504
rect 2268 2436 2276 2444
rect 2316 2436 2324 2444
rect 2268 2236 2276 2244
rect 2300 2236 2308 2244
rect 2300 2176 2308 2184
rect 2236 2136 2244 2144
rect 2268 2136 2276 2144
rect 2316 2116 2324 2124
rect 2364 2536 2372 2544
rect 2396 2536 2404 2544
rect 2348 2236 2356 2244
rect 2364 2196 2372 2204
rect 2380 2176 2388 2184
rect 2444 2536 2452 2544
rect 2412 2516 2420 2524
rect 2428 2516 2436 2524
rect 2428 2176 2436 2184
rect 2684 2556 2692 2564
rect 2572 2516 2580 2524
rect 2716 2516 2724 2524
rect 2524 2496 2532 2504
rect 2668 2316 2676 2324
rect 2588 2296 2596 2304
rect 2636 2296 2644 2304
rect 2572 2276 2580 2284
rect 2492 2236 2500 2244
rect 2524 2236 2532 2244
rect 2492 2216 2500 2224
rect 2556 2216 2564 2224
rect 2524 2196 2532 2204
rect 2540 2196 2548 2204
rect 2460 2156 2468 2164
rect 2508 2156 2516 2164
rect 2604 2156 2612 2164
rect 2444 2136 2452 2144
rect 2572 2136 2580 2144
rect 2636 2136 2644 2144
rect 2428 2116 2436 2124
rect 2588 2116 2596 2124
rect 2604 2116 2612 2124
rect 2652 2116 2660 2124
rect 2460 2096 2468 2104
rect 2252 1996 2260 2004
rect 2220 1976 2228 1984
rect 2236 1856 2244 1864
rect 2316 1856 2324 1864
rect 2268 1836 2276 1844
rect 2284 1836 2292 1844
rect 2252 1796 2260 1804
rect 2284 1796 2292 1804
rect 2188 1756 2196 1764
rect 2236 1756 2244 1764
rect 2044 1736 2052 1744
rect 2028 1716 2036 1724
rect 2076 1716 2084 1724
rect 2124 1716 2132 1724
rect 1996 1696 2004 1704
rect 2092 1696 2100 1704
rect 2012 1676 2020 1684
rect 1916 1616 1924 1624
rect 1900 1596 1908 1604
rect 1932 1596 1940 1604
rect 1852 1516 1860 1524
rect 1868 1516 1876 1524
rect 1900 1516 1908 1524
rect 1884 1476 1892 1484
rect 1804 1416 1812 1424
rect 1772 1396 1780 1404
rect 1788 1396 1796 1404
rect 1660 1376 1668 1384
rect 1676 1356 1684 1364
rect 1708 1356 1716 1364
rect 1804 1356 1812 1364
rect 1596 1256 1604 1264
rect 1308 1156 1316 1164
rect 1452 1196 1460 1204
rect 1420 1156 1428 1164
rect 1260 1136 1268 1144
rect 1276 1136 1284 1144
rect 1116 1116 1124 1124
rect 1196 1116 1204 1124
rect 1404 1116 1412 1124
rect 1212 1076 1220 1084
rect 1292 1076 1300 1084
rect 1324 1076 1332 1084
rect 1340 1076 1342 1084
rect 1342 1076 1348 1084
rect 1420 1076 1428 1084
rect 1420 1056 1428 1064
rect 1100 1036 1108 1044
rect 1228 1036 1236 1044
rect 1292 1036 1300 1044
rect 1020 996 1028 1004
rect 1132 1016 1140 1024
rect 1164 1016 1172 1024
rect 1388 1016 1396 1024
rect 924 936 932 944
rect 956 936 958 944
rect 958 936 964 944
rect 988 936 996 944
rect 1004 936 1012 944
rect 1148 936 1156 944
rect 908 876 916 884
rect 1404 996 1412 1004
rect 1212 936 1220 944
rect 1404 936 1412 944
rect 892 856 900 864
rect 1196 856 1204 864
rect 1132 836 1140 844
rect 972 816 980 824
rect 1084 816 1092 824
rect 876 776 884 784
rect 636 716 644 724
rect 508 596 516 604
rect 700 696 708 704
rect 812 716 820 724
rect 780 676 788 684
rect 716 656 724 664
rect 764 616 772 624
rect 604 596 612 604
rect 652 596 660 604
rect 668 596 676 604
rect 860 616 868 624
rect 1036 716 1044 724
rect 908 676 914 684
rect 914 676 916 684
rect 956 676 964 684
rect 1004 676 1012 684
rect 892 616 900 624
rect 908 616 916 624
rect 876 576 884 584
rect 988 576 996 584
rect 956 556 964 564
rect 1100 776 1108 784
rect 1260 916 1268 924
rect 1324 876 1332 884
rect 1340 876 1348 884
rect 1228 816 1236 824
rect 1212 796 1220 804
rect 1260 796 1268 804
rect 1180 756 1188 764
rect 1228 756 1236 764
rect 1356 816 1364 824
rect 1228 716 1236 724
rect 1276 716 1284 724
rect 1420 716 1428 724
rect 1436 716 1444 724
rect 1132 676 1140 684
rect 1180 676 1188 684
rect 1068 616 1076 624
rect 1212 616 1220 624
rect 1276 656 1284 664
rect 1100 576 1108 584
rect 1164 556 1172 564
rect 1308 636 1316 644
rect 1372 616 1380 624
rect 1356 576 1364 584
rect 716 536 724 544
rect 1132 536 1140 544
rect 1276 536 1284 544
rect 108 496 116 504
rect 188 496 196 504
rect 236 496 244 504
rect 300 496 308 504
rect 140 316 148 324
rect 172 296 180 304
rect 76 276 84 284
rect 284 476 292 484
rect 364 476 372 484
rect 428 396 436 404
rect 380 356 388 364
rect 380 316 388 324
rect 220 276 228 284
rect 252 276 254 284
rect 254 276 260 284
rect 316 276 324 284
rect 12 256 20 264
rect 44 256 52 264
rect 124 236 132 244
rect 204 236 212 244
rect 28 176 36 184
rect 60 176 68 184
rect 76 176 84 184
rect 252 176 260 184
rect 332 196 340 204
rect 348 196 356 204
rect 236 156 244 164
rect 284 156 292 164
rect 460 336 468 344
rect 492 316 500 324
rect 540 516 548 524
rect 604 516 612 524
rect 796 516 804 524
rect 844 516 852 524
rect 940 516 948 524
rect 1324 496 1332 504
rect 588 336 596 344
rect 556 316 564 324
rect 716 356 724 364
rect 476 276 484 284
rect 572 276 580 284
rect 620 276 628 284
rect 700 276 708 284
rect 1212 476 1220 484
rect 780 356 788 364
rect 764 276 772 284
rect 732 256 740 264
rect 444 236 452 244
rect 460 236 468 244
rect 700 216 708 224
rect 524 196 532 204
rect 556 196 564 204
rect 508 176 516 184
rect 364 156 372 164
rect 44 136 52 144
rect 124 136 126 144
rect 126 136 132 144
rect 572 176 580 184
rect 1084 416 1092 424
rect 1084 396 1092 404
rect 1068 316 1076 324
rect 796 276 804 284
rect 828 276 836 284
rect 876 276 884 284
rect 892 276 900 284
rect 1148 336 1156 344
rect 1196 336 1204 344
rect 1324 336 1332 344
rect 1148 316 1156 324
rect 1212 316 1220 324
rect 1260 316 1268 324
rect 1100 276 1108 284
rect 1132 276 1140 284
rect 1356 316 1364 324
rect 1372 316 1380 324
rect 1164 276 1172 284
rect 1228 276 1236 284
rect 1276 276 1284 284
rect 1404 676 1412 684
rect 1420 656 1428 664
rect 1484 1056 1492 1064
rect 1500 1036 1508 1044
rect 1468 996 1476 1004
rect 1852 1456 1860 1464
rect 1852 1356 1860 1364
rect 1724 1296 1732 1304
rect 1628 1276 1636 1284
rect 1964 1476 1972 1484
rect 2028 1556 2036 1564
rect 2060 1556 2068 1564
rect 2044 1536 2052 1544
rect 2108 1636 2116 1644
rect 2300 1776 2308 1784
rect 2300 1756 2308 1764
rect 2444 1956 2452 1964
rect 2524 1936 2532 1944
rect 2348 1856 2356 1864
rect 2428 1876 2436 1884
rect 2492 1836 2500 1844
rect 2428 1776 2436 1784
rect 2492 1776 2500 1784
rect 2300 1716 2308 1724
rect 2236 1696 2244 1704
rect 2220 1616 2228 1624
rect 1900 1456 1908 1464
rect 2172 1536 2180 1544
rect 2236 1536 2244 1544
rect 2172 1516 2180 1524
rect 2284 1516 2292 1524
rect 2236 1496 2244 1504
rect 2332 1516 2340 1524
rect 2380 1756 2388 1764
rect 2412 1756 2420 1764
rect 2396 1716 2404 1724
rect 2412 1716 2420 1724
rect 2444 1716 2452 1724
rect 2364 1616 2372 1624
rect 2444 1676 2452 1684
rect 2444 1596 2452 1604
rect 2428 1516 2436 1524
rect 2476 1516 2484 1524
rect 2188 1476 2196 1484
rect 2204 1476 2212 1484
rect 2300 1476 2308 1484
rect 2348 1476 2356 1484
rect 2316 1456 2324 1464
rect 2380 1456 2388 1464
rect 2092 1416 2100 1424
rect 2124 1416 2132 1424
rect 1996 1396 2004 1404
rect 2124 1396 2132 1404
rect 2060 1376 2068 1384
rect 2252 1416 2260 1424
rect 2076 1356 2084 1364
rect 2140 1356 2148 1364
rect 2300 1396 2308 1404
rect 2380 1436 2388 1444
rect 1948 1336 1956 1344
rect 2044 1336 2052 1344
rect 1852 1316 1860 1324
rect 1884 1316 1892 1324
rect 1772 1256 1780 1264
rect 1676 1176 1684 1184
rect 1612 1156 1620 1164
rect 1868 1296 1876 1304
rect 1884 1296 1892 1304
rect 1932 1276 1940 1284
rect 1852 1196 1860 1204
rect 1836 1136 1844 1144
rect 2044 1296 2052 1304
rect 1996 1156 2004 1164
rect 1740 1116 1748 1124
rect 1772 1116 1780 1124
rect 1804 1116 1812 1124
rect 1644 1076 1652 1084
rect 1548 1036 1556 1044
rect 1532 996 1540 1004
rect 1532 956 1540 964
rect 1484 916 1492 924
rect 1628 1056 1636 1064
rect 1660 1056 1668 1064
rect 1596 936 1604 944
rect 1564 876 1572 884
rect 1500 856 1508 864
rect 1580 796 1588 804
rect 1580 756 1588 764
rect 1612 756 1620 764
rect 1740 1056 1748 1064
rect 1948 1116 1956 1124
rect 1980 1116 1988 1124
rect 1708 1036 1716 1044
rect 1820 1036 1828 1044
rect 1676 956 1684 964
rect 1756 956 1764 964
rect 1868 1056 1876 1064
rect 1900 1056 1908 1064
rect 2124 1316 2132 1324
rect 2108 1296 2116 1304
rect 2044 1116 2052 1124
rect 2076 1116 2084 1124
rect 2092 1096 2100 1104
rect 2172 1296 2180 1304
rect 2236 1276 2244 1284
rect 2220 1236 2228 1244
rect 2268 1296 2276 1304
rect 2348 1296 2356 1304
rect 2380 1296 2388 1304
rect 2364 1276 2372 1284
rect 2380 1236 2388 1244
rect 2380 1196 2388 1204
rect 2252 1176 2260 1184
rect 2364 1156 2372 1164
rect 2332 1116 2340 1124
rect 2444 1496 2452 1504
rect 2572 1896 2580 1904
rect 2540 1856 2548 1864
rect 2556 1796 2564 1804
rect 2572 1776 2580 1784
rect 2540 1716 2548 1724
rect 2620 2056 2628 2064
rect 2652 1916 2660 1924
rect 2620 1896 2628 1904
rect 2620 1856 2628 1864
rect 2604 1776 2612 1784
rect 2636 1816 2644 1824
rect 2636 1756 2644 1764
rect 2604 1676 2612 1684
rect 2588 1636 2596 1644
rect 2572 1516 2580 1524
rect 2556 1496 2564 1504
rect 2604 1496 2612 1504
rect 2620 1496 2628 1504
rect 2508 1476 2516 1484
rect 2444 1396 2452 1404
rect 2588 1356 2596 1364
rect 2444 1336 2452 1344
rect 2508 1336 2516 1344
rect 2540 1336 2548 1344
rect 2524 1316 2532 1324
rect 2460 1296 2468 1304
rect 2508 1296 2516 1304
rect 2492 1276 2500 1284
rect 2444 1196 2452 1204
rect 2636 1336 2644 1344
rect 2620 1316 2628 1324
rect 2716 2296 2724 2304
rect 2700 2276 2708 2284
rect 2700 2156 2708 2164
rect 2684 2096 2692 2104
rect 2780 2496 2788 2504
rect 2780 2316 2788 2324
rect 2764 2256 2772 2264
rect 2764 2216 2772 2224
rect 2748 2196 2756 2204
rect 2764 2036 2772 2044
rect 2732 2016 2740 2024
rect 2780 1976 2788 1984
rect 2684 1936 2692 1944
rect 2684 1916 2692 1924
rect 2732 1916 2740 1924
rect 2748 1876 2756 1884
rect 2700 1796 2708 1804
rect 2748 1776 2756 1784
rect 2716 1736 2724 1744
rect 2764 1736 2772 1744
rect 2940 2596 2948 2604
rect 2892 2556 2900 2564
rect 2956 2556 2964 2564
rect 3036 3096 3044 3104
rect 2988 3016 2996 3024
rect 3004 2956 3012 2964
rect 3068 3696 3076 3704
rect 3132 3616 3140 3624
rect 3388 3936 3396 3944
rect 3612 3936 3620 3944
rect 3644 3936 3652 3944
rect 3964 3936 3972 3944
rect 4060 3936 4068 3944
rect 4156 3936 4164 3944
rect 4252 3936 4260 3944
rect 3468 3916 3476 3924
rect 3836 3916 3844 3924
rect 4044 3916 4052 3924
rect 4172 3916 4180 3924
rect 4188 3916 4196 3924
rect 4236 3916 4244 3924
rect 3340 3896 3348 3904
rect 3452 3896 3460 3904
rect 3548 3896 3556 3904
rect 3708 3896 3716 3904
rect 3740 3896 3748 3904
rect 3756 3896 3764 3904
rect 3468 3876 3476 3884
rect 3692 3876 3700 3884
rect 3420 3856 3428 3864
rect 3404 3836 3412 3844
rect 3372 3816 3380 3824
rect 3436 3816 3444 3824
rect 3260 3796 3268 3804
rect 3356 3756 3364 3764
rect 3228 3716 3236 3724
rect 3212 3636 3220 3644
rect 3148 3576 3156 3584
rect 3084 3536 3092 3544
rect 3148 3536 3156 3544
rect 3068 3516 3076 3524
rect 3116 3476 3124 3484
rect 3132 3476 3140 3484
rect 3324 3676 3332 3684
rect 3244 3576 3252 3584
rect 3228 3536 3236 3544
rect 3260 3536 3268 3544
rect 3452 3796 3460 3804
rect 3468 3756 3476 3764
rect 3420 3696 3428 3704
rect 3388 3596 3396 3604
rect 3340 3576 3348 3584
rect 3388 3536 3396 3544
rect 3212 3476 3220 3484
rect 3644 3776 3652 3784
rect 3580 3756 3588 3764
rect 3628 3756 3636 3764
rect 3564 3716 3572 3724
rect 3516 3696 3524 3704
rect 3596 3696 3604 3704
rect 3676 3696 3684 3704
rect 3548 3596 3556 3604
rect 3468 3536 3476 3544
rect 3484 3536 3492 3544
rect 3660 3576 3668 3584
rect 3212 3456 3220 3464
rect 3196 3416 3204 3424
rect 3276 3416 3284 3424
rect 3212 3376 3220 3384
rect 3084 3356 3092 3364
rect 3116 3356 3124 3364
rect 3292 3356 3300 3364
rect 3100 3336 3108 3344
rect 3228 3316 3236 3324
rect 3196 3296 3204 3304
rect 3260 3296 3268 3304
rect 3340 3416 3348 3424
rect 3356 3416 3364 3424
rect 3404 3436 3412 3444
rect 3340 3376 3348 3384
rect 3388 3376 3396 3384
rect 3532 3416 3540 3424
rect 3500 3396 3508 3404
rect 3420 3356 3428 3364
rect 3468 3356 3476 3364
rect 3516 3376 3524 3384
rect 3596 3416 3604 3424
rect 3660 3496 3668 3504
rect 3756 3876 3764 3884
rect 3788 3876 3796 3884
rect 3868 3876 3876 3884
rect 4108 3876 4116 3884
rect 3996 3856 4004 3864
rect 3804 3836 3812 3844
rect 3788 3816 3796 3824
rect 3772 3796 3780 3804
rect 3756 3756 3764 3764
rect 3724 3696 3732 3704
rect 3708 3596 3716 3604
rect 3900 3816 3908 3824
rect 3916 3756 3924 3764
rect 3852 3736 3860 3744
rect 3868 3736 3876 3744
rect 3980 3736 3988 3744
rect 3772 3696 3780 3704
rect 4028 3796 4036 3804
rect 4092 3796 4100 3804
rect 4348 3936 4356 3944
rect 4396 3936 4404 3944
rect 4636 3916 4644 3924
rect 4684 3916 4692 3924
rect 4700 3916 4708 3924
rect 4732 3916 4740 3924
rect 4460 3896 4468 3904
rect 4492 3896 4500 3904
rect 4316 3856 4324 3864
rect 4124 3816 4132 3824
rect 4172 3816 4180 3824
rect 4156 3796 4164 3804
rect 4108 3776 4116 3784
rect 4220 3796 4228 3804
rect 4044 3716 4052 3724
rect 4012 3696 4020 3704
rect 3964 3656 3972 3664
rect 3820 3596 3828 3604
rect 3964 3536 3972 3544
rect 3756 3516 3764 3524
rect 3692 3476 3700 3484
rect 3724 3476 3732 3484
rect 3612 3396 3620 3404
rect 3580 3356 3588 3364
rect 3644 3356 3652 3364
rect 3740 3456 3748 3464
rect 3708 3356 3716 3364
rect 3884 3476 3892 3484
rect 3308 3336 3316 3344
rect 3324 3336 3332 3344
rect 3356 3336 3364 3344
rect 3644 3336 3652 3344
rect 3756 3336 3764 3344
rect 3276 3256 3284 3264
rect 3068 3196 3076 3204
rect 3260 3116 3268 3124
rect 3068 3096 3076 3104
rect 3116 3096 3124 3104
rect 3084 2996 3092 3004
rect 2988 2916 2996 2924
rect 3020 2896 3028 2904
rect 3052 2876 3060 2884
rect 3068 2776 3076 2784
rect 3020 2736 3028 2744
rect 3004 2716 3012 2724
rect 3324 3316 3332 3324
rect 3404 3316 3412 3324
rect 3436 3316 3444 3324
rect 3500 3316 3508 3324
rect 3580 3316 3588 3324
rect 3324 3176 3332 3184
rect 3308 3116 3316 3124
rect 3292 3096 3300 3104
rect 3340 3116 3348 3124
rect 3420 3096 3428 3104
rect 3276 3056 3284 3064
rect 3180 2996 3188 3004
rect 3212 2996 3220 3004
rect 3260 2996 3268 3004
rect 3148 2976 3156 2984
rect 3324 3036 3332 3044
rect 3356 3056 3364 3064
rect 3372 3056 3380 3064
rect 3404 3056 3412 3064
rect 3132 2916 3140 2924
rect 3164 2916 3172 2924
rect 3116 2896 3124 2904
rect 3212 2896 3220 2904
rect 3228 2896 3236 2904
rect 3308 2856 3316 2864
rect 3356 3016 3364 3024
rect 3340 2996 3348 3004
rect 3404 2976 3412 2984
rect 3340 2896 3348 2904
rect 3388 2896 3396 2904
rect 3324 2816 3332 2824
rect 3324 2796 3332 2804
rect 3100 2736 3108 2744
rect 3100 2716 3108 2724
rect 3228 2716 3236 2724
rect 3276 2716 3284 2724
rect 3084 2696 3092 2704
rect 3164 2696 3172 2704
rect 3404 2836 3412 2844
rect 3564 3196 3572 3204
rect 3452 3176 3460 3184
rect 3468 3136 3476 3144
rect 3532 3136 3540 3144
rect 3452 3116 3460 3124
rect 3500 3096 3508 3104
rect 3548 3116 3556 3124
rect 3644 3156 3652 3164
rect 3676 3096 3684 3104
rect 3516 3036 3524 3044
rect 3740 3176 3748 3184
rect 3852 3456 3860 3464
rect 3804 3316 3812 3324
rect 3852 3316 3860 3324
rect 3788 3216 3796 3224
rect 3788 3136 3796 3144
rect 3852 3136 3860 3144
rect 3724 3056 3732 3064
rect 3692 3036 3700 3044
rect 3660 3016 3668 3024
rect 3596 2996 3604 3004
rect 3708 2996 3716 3004
rect 3452 2976 3460 2984
rect 3500 2976 3508 2984
rect 3580 2976 3588 2984
rect 3436 2916 3444 2924
rect 3564 2956 3572 2964
rect 3724 2956 3732 2964
rect 3500 2916 3508 2924
rect 3596 2916 3604 2924
rect 3644 2916 3652 2924
rect 3692 2916 3700 2924
rect 3724 2916 3732 2924
rect 3468 2896 3476 2904
rect 3484 2896 3492 2904
rect 3548 2896 3556 2904
rect 3612 2896 3620 2904
rect 3660 2896 3668 2904
rect 3420 2816 3428 2824
rect 3740 2856 3748 2864
rect 3660 2816 3668 2824
rect 3692 2816 3700 2824
rect 3516 2776 3524 2784
rect 3452 2756 3460 2764
rect 3420 2716 3428 2724
rect 3548 2716 3556 2724
rect 3596 2716 3604 2724
rect 3612 2696 3620 2704
rect 3708 2696 3716 2704
rect 3292 2676 3300 2684
rect 3324 2676 3332 2684
rect 3500 2676 3508 2684
rect 3052 2636 3060 2644
rect 2988 2596 2996 2604
rect 3004 2576 3012 2584
rect 2988 2556 2996 2564
rect 3020 2556 3028 2564
rect 2844 2336 2852 2344
rect 2812 2256 2820 2264
rect 2956 2496 2964 2504
rect 2892 2336 2900 2344
rect 2972 2316 2980 2324
rect 2956 2296 2964 2304
rect 2924 2276 2932 2284
rect 3036 2476 3044 2484
rect 3132 2616 3140 2624
rect 3100 2576 3108 2584
rect 3084 2556 3092 2564
rect 3228 2576 3236 2584
rect 3100 2536 3108 2544
rect 3148 2536 3156 2544
rect 3132 2496 3140 2504
rect 3068 2456 3076 2464
rect 3180 2456 3188 2464
rect 3132 2436 3140 2444
rect 3404 2636 3412 2644
rect 3516 2636 3524 2644
rect 3356 2616 3364 2624
rect 3324 2576 3332 2584
rect 3340 2576 3348 2584
rect 3260 2536 3268 2544
rect 3532 2616 3540 2624
rect 3580 2616 3588 2624
rect 3516 2576 3524 2584
rect 3580 2596 3588 2604
rect 3596 2596 3604 2604
rect 3500 2536 3508 2544
rect 3276 2496 3284 2504
rect 3340 2496 3348 2504
rect 3404 2496 3412 2504
rect 3436 2496 3444 2504
rect 3548 2496 3556 2504
rect 3212 2456 3220 2464
rect 3292 2456 3300 2464
rect 3212 2396 3220 2404
rect 3196 2356 3204 2364
rect 3404 2476 3412 2484
rect 3388 2456 3396 2464
rect 3372 2336 3380 2344
rect 3020 2316 3028 2324
rect 3084 2316 3092 2324
rect 3180 2316 3188 2324
rect 3084 2296 3092 2304
rect 3196 2296 3204 2304
rect 3052 2276 3060 2284
rect 3276 2276 3284 2284
rect 2940 2256 2948 2264
rect 2972 2256 2980 2264
rect 2988 2256 2996 2264
rect 3068 2256 3076 2264
rect 3116 2256 3124 2264
rect 2876 2216 2884 2224
rect 2956 2176 2964 2184
rect 2828 2156 2836 2164
rect 2892 2156 2900 2164
rect 2828 2136 2836 2144
rect 2812 2116 2820 2124
rect 2924 2116 2932 2124
rect 3004 2176 3012 2184
rect 3020 2156 3028 2164
rect 3052 2136 3060 2144
rect 3084 2136 3092 2144
rect 3100 2136 3108 2144
rect 3004 2116 3012 2124
rect 3260 2236 3268 2244
rect 3836 3016 3844 3024
rect 3836 2996 3844 3004
rect 3820 2896 3828 2904
rect 3772 2856 3780 2864
rect 3788 2836 3796 2844
rect 3852 2816 3860 2824
rect 3884 3456 3892 3464
rect 3900 3396 3908 3404
rect 4028 3536 4036 3544
rect 4124 3696 4132 3704
rect 4140 3676 4148 3684
rect 4060 3516 4068 3524
rect 4108 3516 4116 3524
rect 4124 3516 4132 3524
rect 4044 3496 4052 3504
rect 4220 3696 4228 3704
rect 4252 3736 4260 3744
rect 4300 3816 4308 3824
rect 4300 3756 4308 3764
rect 4332 3756 4340 3764
rect 4316 3736 4324 3744
rect 4412 3816 4420 3824
rect 4476 3836 4484 3844
rect 4556 3896 4564 3904
rect 4524 3816 4532 3824
rect 4476 3796 4484 3804
rect 4956 3936 4964 3944
rect 5068 3936 5076 3944
rect 4924 3916 4932 3924
rect 5004 3916 5012 3924
rect 5196 3916 5204 3924
rect 5292 3916 5300 3924
rect 4748 3856 4756 3864
rect 4764 3856 4772 3864
rect 4572 3796 4580 3804
rect 4668 3796 4676 3804
rect 4428 3756 4436 3764
rect 4444 3756 4452 3764
rect 4460 3756 4468 3764
rect 4748 3776 4756 3784
rect 4716 3756 4724 3764
rect 4732 3756 4740 3764
rect 4300 3696 4308 3704
rect 4364 3696 4372 3704
rect 4748 3716 4756 3724
rect 4620 3696 4628 3704
rect 4636 3696 4644 3704
rect 4684 3696 4692 3704
rect 4700 3696 4708 3704
rect 4236 3576 4244 3584
rect 4236 3536 4244 3544
rect 4252 3516 4260 3524
rect 4300 3516 4308 3524
rect 4380 3556 4388 3564
rect 4428 3556 4436 3564
rect 4380 3536 4388 3544
rect 4412 3536 4420 3544
rect 4172 3476 4180 3484
rect 3996 3456 4004 3464
rect 4012 3456 4020 3464
rect 4060 3456 4068 3464
rect 4172 3456 4180 3464
rect 4188 3456 4196 3464
rect 4236 3456 4244 3464
rect 3980 3416 3988 3424
rect 4044 3416 4052 3424
rect 3916 3296 3924 3304
rect 3884 3256 3892 3264
rect 3948 3176 3956 3184
rect 4284 3436 4292 3444
rect 4108 3396 4116 3404
rect 4076 3336 4084 3344
rect 4092 3296 4100 3304
rect 4060 3136 4068 3144
rect 4124 3256 4132 3264
rect 4236 3416 4244 3424
rect 4172 3396 4180 3404
rect 4284 3396 4292 3404
rect 4364 3456 4372 3464
rect 4396 3456 4404 3464
rect 4348 3396 4356 3404
rect 4524 3636 4532 3644
rect 4492 3596 4500 3604
rect 4892 3876 4900 3884
rect 4812 3776 4820 3784
rect 4876 3776 4884 3784
rect 4812 3756 4820 3764
rect 4796 3696 4804 3704
rect 4844 3696 4852 3704
rect 4780 3656 4788 3664
rect 4716 3536 4724 3544
rect 4460 3516 4468 3524
rect 4508 3516 4516 3524
rect 4524 3516 4532 3524
rect 4732 3516 4740 3524
rect 4748 3516 4756 3524
rect 4652 3496 4660 3504
rect 4476 3436 4484 3444
rect 4540 3396 4548 3404
rect 4428 3376 4436 3384
rect 4444 3376 4452 3384
rect 4396 3336 4404 3344
rect 4156 3196 4164 3204
rect 4124 3176 4132 3184
rect 4188 3296 4196 3304
rect 4268 3276 4276 3284
rect 4076 3116 4084 3124
rect 4108 3116 4116 3124
rect 4172 3116 4180 3124
rect 3900 3076 3908 3084
rect 3916 3036 3924 3044
rect 3948 3016 3956 3024
rect 3884 2996 3892 3004
rect 3884 2916 3892 2924
rect 3980 2996 3988 3004
rect 4044 2936 4052 2944
rect 4284 3176 4292 3184
rect 4268 3156 4276 3164
rect 4172 3096 4180 3104
rect 4252 3096 4260 3104
rect 4092 3036 4100 3044
rect 4188 2996 4196 3004
rect 4076 2956 4084 2964
rect 4108 2956 4116 2964
rect 4156 2956 4164 2964
rect 4156 2936 4164 2944
rect 3964 2916 3972 2924
rect 4028 2916 4036 2924
rect 4060 2916 4068 2924
rect 3964 2896 3972 2904
rect 4060 2896 4068 2904
rect 3996 2836 4004 2844
rect 3884 2816 3892 2824
rect 3868 2796 3876 2804
rect 3836 2736 3844 2744
rect 3788 2716 3796 2724
rect 3804 2696 3812 2704
rect 3628 2676 3636 2684
rect 3756 2676 3764 2684
rect 3788 2676 3796 2684
rect 3644 2656 3652 2664
rect 3708 2656 3716 2664
rect 3740 2656 3748 2664
rect 3756 2616 3764 2624
rect 3644 2536 3652 2544
rect 3628 2496 3636 2504
rect 3660 2496 3668 2504
rect 3708 2576 3716 2584
rect 3740 2536 3748 2544
rect 3676 2476 3684 2484
rect 3692 2456 3700 2464
rect 3740 2476 3748 2484
rect 3644 2376 3652 2384
rect 3724 2376 3732 2384
rect 3500 2336 3508 2344
rect 3612 2336 3620 2344
rect 3660 2336 3668 2344
rect 3564 2316 3572 2324
rect 3388 2296 3396 2304
rect 3340 2276 3348 2284
rect 3372 2276 3380 2284
rect 3324 2256 3332 2264
rect 3404 2256 3412 2264
rect 3452 2296 3460 2304
rect 3516 2296 3524 2304
rect 3596 2296 3604 2304
rect 3724 2296 3732 2304
rect 3532 2276 3538 2284
rect 3538 2276 3540 2284
rect 3596 2276 3604 2284
rect 3468 2256 3476 2264
rect 3580 2256 3588 2264
rect 3580 2216 3588 2224
rect 3660 2216 3668 2224
rect 3260 2196 3268 2204
rect 3292 2196 3300 2204
rect 3308 2196 3316 2204
rect 3420 2196 3428 2204
rect 3452 2196 3460 2204
rect 3340 2176 3348 2184
rect 3420 2176 3428 2184
rect 3596 2176 3604 2184
rect 3244 2116 3252 2124
rect 2972 2096 2980 2104
rect 3148 2096 3156 2104
rect 3164 2096 3172 2104
rect 3212 2096 3220 2104
rect 2940 2036 2948 2044
rect 2956 1996 2964 2004
rect 2988 2076 2996 2084
rect 3212 2076 3220 2084
rect 3020 2056 3028 2064
rect 3196 2016 3204 2024
rect 3196 1976 3204 1984
rect 3100 1956 3108 1964
rect 2844 1936 2852 1944
rect 2892 1936 2900 1944
rect 2876 1916 2884 1924
rect 2828 1896 2836 1904
rect 2844 1896 2852 1904
rect 3052 1896 3060 1904
rect 3148 1916 3156 1924
rect 3260 1936 3268 1944
rect 3228 1896 3236 1904
rect 2908 1876 2916 1884
rect 2940 1876 2948 1884
rect 3020 1856 3028 1864
rect 3036 1856 3044 1864
rect 3052 1856 3060 1864
rect 3084 1856 3092 1864
rect 3228 1856 3236 1864
rect 2828 1836 2836 1844
rect 2940 1836 2948 1844
rect 2988 1836 2996 1844
rect 2828 1796 2836 1804
rect 2812 1776 2820 1784
rect 2876 1776 2884 1784
rect 2908 1756 2916 1764
rect 2844 1736 2852 1744
rect 2892 1736 2900 1744
rect 2924 1736 2932 1744
rect 2796 1716 2804 1724
rect 2700 1696 2708 1704
rect 2700 1596 2708 1604
rect 2684 1516 2692 1524
rect 2700 1416 2708 1424
rect 2684 1356 2692 1364
rect 2716 1336 2724 1344
rect 2652 1296 2660 1304
rect 2604 1276 2612 1284
rect 2540 1196 2548 1204
rect 2444 1176 2452 1184
rect 2476 1156 2484 1164
rect 2316 1096 2324 1104
rect 2396 1096 2404 1104
rect 2604 1136 2612 1144
rect 2700 1276 2708 1284
rect 2892 1516 2900 1524
rect 2748 1496 2756 1504
rect 2796 1496 2804 1504
rect 2780 1476 2788 1484
rect 2748 1456 2756 1464
rect 2764 1436 2772 1444
rect 2908 1476 2916 1484
rect 2812 1436 2820 1444
rect 2748 1356 2756 1364
rect 2828 1356 2836 1364
rect 2764 1316 2772 1324
rect 2780 1296 2788 1304
rect 2780 1276 2788 1284
rect 2732 1256 2740 1264
rect 2620 1116 2628 1124
rect 2668 1116 2676 1124
rect 2412 1076 2420 1084
rect 2108 1056 2116 1064
rect 2188 1056 2196 1064
rect 2204 1056 2212 1064
rect 2236 1056 2244 1064
rect 1868 1036 1876 1044
rect 1916 1036 1924 1044
rect 1948 1036 1956 1044
rect 1836 1016 1844 1024
rect 1852 1016 1860 1024
rect 1964 1016 1972 1024
rect 1900 996 1908 1004
rect 1884 976 1892 984
rect 1804 916 1812 924
rect 1868 916 1876 924
rect 1644 896 1652 904
rect 1660 896 1668 904
rect 1692 896 1700 904
rect 1852 816 1860 824
rect 1676 776 1684 784
rect 1756 776 1764 784
rect 1612 676 1620 684
rect 1628 676 1636 684
rect 1596 656 1604 664
rect 1420 636 1428 644
rect 1452 636 1460 644
rect 1468 636 1476 644
rect 1532 636 1540 644
rect 1436 616 1444 624
rect 1484 616 1492 624
rect 1612 616 1620 624
rect 1564 596 1572 604
rect 1596 596 1604 604
rect 1436 576 1444 584
rect 1484 576 1492 584
rect 1548 576 1556 584
rect 1564 576 1572 584
rect 1404 456 1412 464
rect 1500 436 1508 444
rect 1404 316 1412 324
rect 1532 376 1540 384
rect 1548 356 1556 364
rect 1628 556 1636 564
rect 1660 556 1668 564
rect 1724 556 1732 564
rect 1852 756 1860 764
rect 1868 736 1876 744
rect 1820 696 1828 704
rect 1980 996 1988 1004
rect 2172 1036 2180 1044
rect 2188 996 2196 1004
rect 1996 956 2004 964
rect 2060 956 2068 964
rect 2140 936 2148 944
rect 1932 896 1940 904
rect 1948 896 1956 904
rect 2124 896 2132 904
rect 2012 836 2020 844
rect 2028 836 2036 844
rect 1948 756 1956 764
rect 1996 756 2004 764
rect 1964 716 1972 724
rect 1868 656 1876 664
rect 1948 656 1956 664
rect 1788 556 1796 564
rect 1836 556 1844 564
rect 1852 556 1860 564
rect 1580 456 1588 464
rect 1660 516 1668 524
rect 1692 516 1700 524
rect 1932 496 1940 504
rect 1692 436 1700 444
rect 1692 416 1700 424
rect 1724 416 1732 424
rect 1772 336 1780 344
rect 1788 276 1796 284
rect 1404 256 1412 264
rect 1468 256 1476 264
rect 1516 256 1524 264
rect 1548 256 1556 264
rect 1612 256 1620 264
rect 1644 256 1652 264
rect 1724 256 1732 264
rect 1852 356 1860 364
rect 924 236 932 244
rect 972 236 980 244
rect 1212 236 1220 244
rect 1420 236 1428 244
rect 1500 236 1508 244
rect 1596 236 1604 244
rect 748 196 756 204
rect 956 196 964 204
rect 716 176 724 184
rect 844 176 852 184
rect 1036 216 1044 224
rect 1292 216 1300 224
rect 1276 196 1284 204
rect 1676 236 1684 244
rect 1740 236 1748 244
rect 1756 216 1764 224
rect 1804 216 1812 224
rect 844 156 852 164
rect 860 156 868 164
rect 1020 156 1028 164
rect 1068 156 1076 164
rect 1084 156 1092 164
rect 908 136 916 144
rect 972 136 980 144
rect 1020 136 1028 144
rect 92 116 100 124
rect 140 116 148 124
rect 188 116 196 124
rect 364 116 372 124
rect 428 116 436 124
rect 444 116 452 124
rect 556 116 564 124
rect 588 116 596 124
rect 604 116 612 124
rect 652 116 660 124
rect 684 116 692 124
rect 732 116 740 124
rect 796 116 804 124
rect 1100 136 1108 144
rect 1132 136 1140 144
rect 1148 136 1156 144
rect 1196 136 1204 144
rect 1212 136 1220 144
rect 1228 136 1236 144
rect 1308 136 1316 144
rect 1324 136 1332 144
rect 524 96 532 104
rect 924 96 932 104
rect 972 96 980 104
rect 1068 96 1076 104
rect 1292 96 1300 104
rect 1340 96 1348 104
rect 1372 96 1380 104
rect 1404 96 1412 104
rect 1420 96 1428 104
rect 1548 96 1556 104
rect 1564 96 1572 104
rect 1596 96 1604 104
rect 1612 96 1620 104
rect 1676 96 1684 104
rect 636 76 644 84
rect 1436 76 1444 84
rect 1452 76 1460 84
rect 1708 76 1716 84
rect 1740 136 1748 144
rect 1788 196 1796 204
rect 1772 136 1780 144
rect 1756 76 1764 84
rect 1724 56 1732 64
rect 1804 56 1812 64
rect 1740 36 1748 44
rect 1852 256 1860 264
rect 1852 196 1860 204
rect 1980 656 1988 664
rect 1980 536 1988 544
rect 2076 796 2084 804
rect 2044 756 2052 764
rect 2028 736 2036 744
rect 2124 736 2132 744
rect 2092 696 2100 704
rect 2188 916 2196 924
rect 2156 776 2164 784
rect 2188 776 2196 784
rect 2140 716 2148 724
rect 2172 736 2180 744
rect 2108 636 2116 644
rect 2140 636 2148 644
rect 2044 616 2052 624
rect 2060 596 2068 604
rect 2172 596 2180 604
rect 2124 556 2132 564
rect 1964 516 1972 524
rect 2156 536 2164 544
rect 2028 496 2036 504
rect 2092 496 2100 504
rect 2140 496 2148 504
rect 2124 356 2132 364
rect 2044 336 2052 344
rect 1900 316 1908 324
rect 2188 496 2196 504
rect 2428 1056 2436 1064
rect 2300 1036 2308 1044
rect 2492 1036 2500 1044
rect 2236 996 2244 1004
rect 2284 996 2292 1004
rect 2428 996 2436 1004
rect 2252 976 2260 984
rect 2284 976 2292 984
rect 2316 976 2324 984
rect 2300 956 2308 964
rect 2492 956 2500 964
rect 2348 936 2356 944
rect 2220 916 2228 924
rect 2284 916 2292 924
rect 2236 856 2244 864
rect 2220 736 2228 744
rect 2252 816 2260 824
rect 2268 776 2276 784
rect 2348 736 2356 744
rect 2396 936 2404 944
rect 2444 936 2452 944
rect 2540 936 2548 944
rect 2700 1036 2708 1044
rect 2572 976 2580 984
rect 2588 976 2596 984
rect 2428 916 2436 924
rect 2556 916 2564 924
rect 2380 776 2388 784
rect 2476 876 2484 884
rect 2492 876 2500 884
rect 2428 736 2436 744
rect 2412 716 2420 724
rect 2220 576 2228 584
rect 2300 576 2308 584
rect 2364 656 2372 664
rect 2444 616 2452 624
rect 2348 576 2356 584
rect 2380 596 2388 604
rect 2380 576 2388 584
rect 2428 576 2436 584
rect 2444 576 2452 584
rect 2332 496 2340 504
rect 2460 476 2468 484
rect 2444 416 2452 424
rect 2412 376 2420 384
rect 2028 296 2036 304
rect 2044 296 2052 304
rect 2124 296 2132 304
rect 2412 336 2420 344
rect 2700 996 2708 1004
rect 2732 996 2740 1004
rect 2876 1316 2884 1324
rect 2908 1296 2916 1304
rect 2796 1096 2804 1104
rect 2812 1076 2820 1084
rect 2812 996 2820 1004
rect 2652 976 2660 984
rect 2684 976 2692 984
rect 2780 976 2788 984
rect 2828 976 2836 984
rect 2620 916 2628 924
rect 2716 896 2724 904
rect 2748 896 2756 904
rect 2764 896 2772 904
rect 2604 876 2612 884
rect 2508 856 2516 864
rect 2748 836 2756 844
rect 2780 876 2788 884
rect 2892 1136 2900 1144
rect 2876 1116 2884 1124
rect 2956 1776 2964 1784
rect 3020 1736 3026 1744
rect 3026 1736 3028 1744
rect 3004 1716 3012 1724
rect 2940 1696 2948 1704
rect 2988 1696 2996 1704
rect 3004 1596 3012 1604
rect 2956 1496 2964 1504
rect 2972 1476 2980 1484
rect 2940 1456 2948 1464
rect 2956 1436 2964 1444
rect 3020 1396 3028 1404
rect 3212 1796 3220 1804
rect 3196 1776 3204 1784
rect 3180 1756 3188 1764
rect 3084 1736 3092 1744
rect 3116 1716 3124 1724
rect 3132 1716 3140 1724
rect 3084 1596 3092 1604
rect 3052 1516 3060 1524
rect 3068 1516 3076 1524
rect 3164 1536 3172 1544
rect 3148 1516 3156 1524
rect 3180 1516 3188 1524
rect 3212 1516 3220 1524
rect 3148 1456 3156 1464
rect 3164 1456 3172 1464
rect 3196 1456 3204 1464
rect 3132 1436 3140 1444
rect 3116 1356 3124 1364
rect 3196 1376 3204 1384
rect 3180 1316 3188 1324
rect 3196 1316 3204 1324
rect 2956 1296 2964 1304
rect 3020 1296 3028 1304
rect 3116 1296 3124 1304
rect 3148 1296 3156 1304
rect 2940 1276 2948 1284
rect 3132 1176 3140 1184
rect 3020 1116 3028 1124
rect 2924 1096 2932 1104
rect 3004 1096 3012 1104
rect 2860 1076 2868 1084
rect 2956 1076 2962 1084
rect 2962 1076 2964 1084
rect 3052 1076 3060 1084
rect 3004 1056 3012 1064
rect 3068 1036 3076 1044
rect 3084 1016 3092 1024
rect 3100 996 3108 1004
rect 3004 956 3012 964
rect 3084 956 3092 964
rect 3068 936 3076 944
rect 2876 916 2884 924
rect 2540 776 2548 784
rect 2556 776 2564 784
rect 2636 776 2644 784
rect 2492 716 2500 724
rect 2540 716 2548 724
rect 2492 696 2500 704
rect 2764 756 2772 764
rect 2620 736 2628 744
rect 2572 696 2580 704
rect 2492 576 2500 584
rect 2572 576 2580 584
rect 2668 696 2676 704
rect 2716 656 2724 664
rect 2748 616 2756 624
rect 2844 816 2852 824
rect 2812 776 2820 784
rect 2908 896 2916 904
rect 2956 896 2964 904
rect 2988 896 2996 904
rect 2892 876 2900 884
rect 2876 856 2884 864
rect 2956 816 2964 824
rect 2940 776 2948 784
rect 2876 736 2884 744
rect 2892 736 2900 744
rect 3036 876 3044 884
rect 3020 796 3028 804
rect 3052 796 3060 804
rect 2812 716 2820 724
rect 2860 716 2868 724
rect 2908 716 2916 724
rect 3020 716 3028 724
rect 2796 696 2804 704
rect 2636 576 2644 584
rect 2700 576 2708 584
rect 2780 576 2788 584
rect 2620 556 2628 564
rect 2652 556 2660 564
rect 2684 556 2692 564
rect 2748 556 2756 564
rect 2828 676 2836 684
rect 2892 676 2900 684
rect 2892 656 2900 664
rect 2700 516 2708 524
rect 2604 496 2612 504
rect 2524 476 2532 484
rect 2652 376 2660 384
rect 2700 376 2708 384
rect 2508 356 2516 364
rect 2556 356 2564 364
rect 2220 316 2228 324
rect 2284 316 2292 324
rect 2460 316 2468 324
rect 2236 296 2244 304
rect 2316 296 2324 304
rect 2540 336 2548 344
rect 1916 276 1924 284
rect 2252 276 2260 284
rect 2444 276 2452 284
rect 2492 276 2500 284
rect 2588 336 2596 344
rect 2684 336 2692 344
rect 2748 336 2756 344
rect 2812 556 2820 564
rect 3068 776 3076 784
rect 3004 676 3012 684
rect 3084 676 3092 684
rect 2956 576 2964 584
rect 2988 556 2996 564
rect 2876 536 2884 544
rect 2908 536 2916 544
rect 2844 516 2852 524
rect 2828 396 2836 404
rect 2812 356 2820 364
rect 2620 316 2628 324
rect 2700 276 2708 284
rect 2748 276 2756 284
rect 2108 256 2116 264
rect 2636 256 2644 264
rect 1916 236 1924 244
rect 2172 236 2180 244
rect 2316 236 2324 244
rect 2364 236 2372 244
rect 2572 236 2580 244
rect 2284 196 2292 204
rect 2188 176 2196 184
rect 1884 136 1892 144
rect 1932 136 1938 144
rect 1938 136 1940 144
rect 2300 176 2308 184
rect 2364 176 2372 184
rect 2124 136 2132 144
rect 2172 136 2180 144
rect 2220 136 2228 144
rect 2236 136 2244 144
rect 2428 176 2436 184
rect 2556 176 2564 184
rect 2620 176 2628 184
rect 2796 176 2804 184
rect 2492 156 2500 164
rect 2604 156 2612 164
rect 1836 96 1844 104
rect 2636 136 2644 144
rect 2684 136 2692 144
rect 2748 136 2756 144
rect 2780 136 2788 144
rect 2060 96 2068 104
rect 2108 96 2116 104
rect 2220 96 2228 104
rect 2380 96 2388 104
rect 1916 76 1924 84
rect 1948 76 1956 84
rect 2172 76 2180 84
rect 2476 76 2484 84
rect 2252 36 2260 44
rect 2540 116 2548 124
rect 2556 116 2564 124
rect 2668 116 2676 124
rect 2748 96 2756 104
rect 2684 36 2692 44
rect 2716 36 2724 44
rect 2828 156 2836 164
rect 3020 616 3028 624
rect 2860 496 2868 504
rect 3004 496 3012 504
rect 2908 476 2916 484
rect 2876 456 2884 464
rect 2860 336 2868 344
rect 2860 316 2868 324
rect 3004 416 3012 424
rect 2988 396 2996 404
rect 2892 276 2900 284
rect 3036 516 3044 524
rect 3068 656 3076 664
rect 3148 1036 3156 1044
rect 3212 1236 3220 1244
rect 3196 1096 3204 1104
rect 3292 1916 3300 1924
rect 3244 1796 3252 1804
rect 3276 1796 3284 1804
rect 3260 1776 3268 1784
rect 3276 1736 3284 1744
rect 3292 1676 3300 1684
rect 3244 1596 3252 1604
rect 3276 1536 3284 1544
rect 3260 1496 3268 1504
rect 3244 1436 3252 1444
rect 3260 1436 3268 1444
rect 3276 1396 3284 1404
rect 3740 2256 3748 2264
rect 3516 2156 3524 2164
rect 3612 2156 3620 2164
rect 3676 2156 3684 2164
rect 3740 2176 3748 2184
rect 3628 2136 3636 2144
rect 3660 2136 3668 2144
rect 3708 2136 3716 2144
rect 3500 2096 3508 2104
rect 3356 2076 3364 2084
rect 3404 2076 3412 2084
rect 3500 2076 3508 2084
rect 3532 2096 3540 2104
rect 3548 2096 3556 2104
rect 3372 2056 3380 2064
rect 3388 2056 3396 2064
rect 3468 2056 3476 2064
rect 3516 2056 3524 2064
rect 3340 2016 3348 2024
rect 3372 2016 3380 2024
rect 3388 1936 3396 1944
rect 3516 1936 3524 1944
rect 3516 1916 3524 1924
rect 3420 1896 3428 1904
rect 3516 1896 3524 1904
rect 3404 1816 3412 1824
rect 3356 1796 3364 1804
rect 3404 1796 3412 1804
rect 3500 1796 3508 1804
rect 3324 1776 3332 1784
rect 3388 1736 3396 1744
rect 3356 1696 3364 1704
rect 3340 1676 3348 1684
rect 3324 1596 3332 1604
rect 3340 1496 3348 1504
rect 3436 1716 3444 1724
rect 3468 1716 3476 1724
rect 3452 1696 3460 1704
rect 3468 1536 3476 1544
rect 3580 1916 3588 1924
rect 3612 1896 3620 1904
rect 3548 1836 3556 1844
rect 3532 1696 3540 1704
rect 3452 1496 3460 1504
rect 3484 1496 3492 1504
rect 3500 1496 3508 1504
rect 3420 1456 3428 1464
rect 3388 1416 3396 1424
rect 3644 2096 3652 2104
rect 3676 2116 3684 2124
rect 3644 1836 3652 1844
rect 3564 1776 3572 1784
rect 3596 1776 3604 1784
rect 3660 1776 3668 1784
rect 3740 2096 3748 2104
rect 3740 1916 3748 1924
rect 3692 1896 3700 1904
rect 3740 1896 3748 1904
rect 3676 1756 3684 1764
rect 3676 1736 3684 1744
rect 3644 1696 3652 1704
rect 3612 1676 3620 1684
rect 3564 1536 3572 1544
rect 3612 1536 3620 1544
rect 3724 1856 3732 1864
rect 3708 1836 3716 1844
rect 3740 1796 3748 1804
rect 3740 1656 3748 1664
rect 3724 1596 3732 1604
rect 3708 1576 3716 1584
rect 3724 1536 3732 1544
rect 3676 1476 3684 1484
rect 3692 1476 3700 1484
rect 3788 2616 3796 2624
rect 3916 2756 3924 2764
rect 4012 2776 4020 2784
rect 4092 2756 4100 2764
rect 4124 2736 4132 2744
rect 3868 2696 3876 2704
rect 3884 2696 3892 2704
rect 3916 2696 3924 2704
rect 3964 2696 3972 2704
rect 4092 2696 4100 2704
rect 4156 2756 4164 2764
rect 4188 2756 4196 2764
rect 4252 2976 4260 2984
rect 4220 2916 4228 2924
rect 4220 2756 4228 2764
rect 4204 2736 4212 2744
rect 4620 3396 4628 3404
rect 4636 3376 4644 3384
rect 4428 3336 4436 3344
rect 4476 3336 4484 3344
rect 4604 3336 4612 3344
rect 4412 3256 4420 3264
rect 4476 3296 4484 3304
rect 4588 3296 4596 3304
rect 4508 3276 4516 3284
rect 4444 3236 4452 3244
rect 4380 3156 4388 3164
rect 4332 3116 4340 3124
rect 4364 3116 4372 3124
rect 4396 3116 4404 3124
rect 4348 3096 4356 3104
rect 4348 3056 4356 3064
rect 4364 3056 4372 3064
rect 4284 3016 4292 3024
rect 4300 2956 4308 2964
rect 4332 2956 4340 2964
rect 4268 2936 4276 2944
rect 4300 2916 4308 2924
rect 4556 3216 4564 3224
rect 4588 3156 4596 3164
rect 4604 3116 4612 3124
rect 4476 3096 4484 3104
rect 4540 3096 4548 3104
rect 4716 3476 4724 3484
rect 4668 3416 4676 3424
rect 4684 3396 4692 3404
rect 4844 3616 4852 3624
rect 4812 3516 4820 3524
rect 4940 3856 4948 3864
rect 5148 3896 5156 3904
rect 5132 3876 5140 3884
rect 5116 3856 5124 3864
rect 5196 3816 5204 3824
rect 5052 3796 5060 3804
rect 5100 3796 5108 3804
rect 5132 3796 5140 3804
rect 4940 3776 4948 3784
rect 4908 3756 4916 3764
rect 5116 3756 5124 3764
rect 4956 3736 4964 3744
rect 4924 3716 4932 3724
rect 4940 3716 4948 3724
rect 4940 3676 4948 3684
rect 5020 3676 5028 3684
rect 5068 3676 5076 3684
rect 4892 3636 4900 3644
rect 5004 3616 5012 3624
rect 5052 3516 5060 3524
rect 5084 3516 5092 3524
rect 4956 3496 4964 3504
rect 4844 3456 4852 3464
rect 4908 3456 4916 3464
rect 4924 3456 4932 3464
rect 4732 3376 4740 3384
rect 4764 3376 4772 3384
rect 4780 3376 4788 3384
rect 4668 3336 4676 3344
rect 4684 3296 4692 3304
rect 4940 3416 4948 3424
rect 4940 3396 4948 3404
rect 4860 3356 4868 3364
rect 4908 3356 4916 3364
rect 4796 3336 4804 3344
rect 4844 3316 4852 3324
rect 4796 3296 4804 3304
rect 4780 3256 4788 3264
rect 4652 3116 4660 3124
rect 4716 3116 4724 3124
rect 4812 3116 4820 3124
rect 4636 3076 4644 3084
rect 4524 3056 4532 3064
rect 4428 3036 4436 3044
rect 4620 3036 4628 3044
rect 4492 3016 4500 3024
rect 4556 3016 4564 3024
rect 4636 3016 4644 3024
rect 4412 2996 4420 3004
rect 4556 2976 4564 2984
rect 4492 2956 4500 2964
rect 4540 2936 4548 2944
rect 4604 2936 4612 2944
rect 4348 2916 4356 2924
rect 4396 2876 4404 2884
rect 4444 2916 4452 2924
rect 4476 2916 4484 2924
rect 4524 2916 4532 2924
rect 4524 2876 4532 2884
rect 4412 2856 4420 2864
rect 4428 2856 4436 2864
rect 4252 2756 4260 2764
rect 4316 2756 4324 2764
rect 4236 2736 4244 2744
rect 4252 2716 4260 2724
rect 4300 2696 4308 2704
rect 4396 2696 4404 2704
rect 4428 2756 4436 2764
rect 3980 2616 3988 2624
rect 3980 2596 3988 2604
rect 3932 2576 3940 2584
rect 3788 2536 3796 2544
rect 3852 2536 3860 2544
rect 3916 2536 3924 2544
rect 4076 2596 4084 2604
rect 4044 2556 4052 2564
rect 4060 2516 4068 2524
rect 4076 2516 4084 2524
rect 3804 2496 3812 2504
rect 4044 2496 4052 2504
rect 3804 2476 3812 2484
rect 3980 2476 3988 2484
rect 3884 2396 3892 2404
rect 3900 2356 3908 2364
rect 3932 2336 3940 2344
rect 3964 2336 3972 2344
rect 3996 2336 4004 2344
rect 3788 2276 3796 2284
rect 3868 2296 3876 2304
rect 3916 2296 3924 2304
rect 3980 2296 3988 2304
rect 4012 2296 4020 2304
rect 3772 2196 3780 2204
rect 3852 2256 3860 2264
rect 3996 2256 4004 2264
rect 4044 2256 4052 2264
rect 3884 2236 3892 2244
rect 3916 2236 3924 2244
rect 4028 2236 4036 2244
rect 3772 2176 3780 2184
rect 3836 2176 3844 2184
rect 3884 2176 3892 2184
rect 4044 2216 4052 2224
rect 3980 2176 3988 2184
rect 3836 2156 3844 2164
rect 3900 2156 3908 2164
rect 3932 2156 3940 2164
rect 3964 2156 3972 2164
rect 3804 2136 3812 2144
rect 3836 2096 3844 2104
rect 4092 2496 4100 2504
rect 4076 2336 4084 2344
rect 4092 2336 4100 2344
rect 4076 2216 4084 2224
rect 3980 2136 3988 2144
rect 4060 2136 4068 2144
rect 3868 2096 3876 2104
rect 3932 2096 3940 2104
rect 3948 2096 3956 2104
rect 3852 2036 3860 2044
rect 4044 2096 4052 2104
rect 3836 1896 3844 1904
rect 3852 1876 3860 1884
rect 3804 1856 3812 1864
rect 3772 1836 3780 1844
rect 3788 1816 3796 1824
rect 3772 1796 3780 1804
rect 3772 1756 3780 1764
rect 3852 1836 3860 1844
rect 4012 1976 4020 1984
rect 4044 1956 4052 1964
rect 4252 2676 4260 2684
rect 4348 2676 4356 2684
rect 4204 2656 4212 2664
rect 4236 2576 4244 2584
rect 4348 2596 4356 2604
rect 4492 2696 4500 2704
rect 4508 2616 4516 2624
rect 4588 2736 4596 2744
rect 4556 2696 4564 2704
rect 4572 2696 4580 2704
rect 4620 2696 4628 2704
rect 4540 2636 4548 2644
rect 4492 2596 4500 2604
rect 4364 2576 4372 2584
rect 4460 2576 4468 2584
rect 4476 2576 4484 2584
rect 4604 2596 4612 2604
rect 4604 2576 4612 2584
rect 4620 2576 4628 2584
rect 4684 3096 4692 3104
rect 4748 3096 4756 3104
rect 4780 3096 4788 3104
rect 4668 3056 4676 3064
rect 4684 3056 4692 3064
rect 4732 2976 4740 2984
rect 4732 2956 4740 2964
rect 5164 3736 5172 3744
rect 5196 3736 5204 3744
rect 5164 3716 5172 3724
rect 5468 3896 5476 3904
rect 5324 3876 5332 3884
rect 5308 3856 5316 3864
rect 5260 3816 5268 3824
rect 5244 3796 5252 3804
rect 5388 3876 5396 3884
rect 5436 3796 5444 3804
rect 5260 3776 5268 3784
rect 5340 3776 5348 3784
rect 5452 3776 5460 3784
rect 5452 3756 5460 3764
rect 5516 3756 5524 3764
rect 5228 3736 5236 3744
rect 5228 3696 5236 3704
rect 5164 3636 5172 3644
rect 5148 3476 5156 3484
rect 5180 3516 5188 3524
rect 5020 3456 5028 3464
rect 5100 3456 5108 3464
rect 5164 3456 5172 3464
rect 5212 3456 5220 3464
rect 4988 3396 4996 3404
rect 5004 3356 5012 3364
rect 5116 3396 5124 3404
rect 5068 3376 5076 3384
rect 5132 3376 5140 3384
rect 5116 3356 5124 3364
rect 4956 3336 4964 3344
rect 5084 3336 5092 3344
rect 4924 3316 4932 3324
rect 5148 3316 5156 3324
rect 4956 3296 4964 3304
rect 4988 3296 4996 3304
rect 5052 3296 5060 3304
rect 4892 3136 4900 3144
rect 4844 3096 4852 3104
rect 4844 3076 4852 3084
rect 4860 3076 4868 3084
rect 4796 3056 4804 3064
rect 4876 3056 4884 3064
rect 4876 3016 4884 3024
rect 4860 2996 4868 3004
rect 4796 2976 4804 2984
rect 4924 3116 4932 3124
rect 4908 2956 4916 2964
rect 4668 2936 4676 2944
rect 4652 2916 4660 2924
rect 4732 2916 4740 2924
rect 4780 2916 4788 2924
rect 4876 2916 4884 2924
rect 4892 2916 4900 2924
rect 4716 2896 4724 2904
rect 4844 2876 4852 2884
rect 4940 2956 4948 2964
rect 4972 3236 4980 3244
rect 5116 3236 5124 3244
rect 5100 3156 5108 3164
rect 4972 3136 4980 3144
rect 5052 3136 5060 3144
rect 4988 3116 4996 3124
rect 5020 3096 5028 3104
rect 5116 3096 5124 3104
rect 5004 3056 5012 3064
rect 5196 3436 5204 3444
rect 5196 3376 5204 3384
rect 5196 3356 5204 3364
rect 5308 3696 5316 3704
rect 5340 3716 5348 3724
rect 5388 3696 5396 3704
rect 5436 3696 5444 3704
rect 5324 3656 5332 3664
rect 5276 3616 5284 3624
rect 5516 3696 5524 3704
rect 5436 3536 5444 3544
rect 5452 3536 5460 3544
rect 5260 3516 5268 3524
rect 5324 3516 5332 3524
rect 5388 3516 5396 3524
rect 5532 3516 5540 3524
rect 5580 3516 5588 3524
rect 5324 3476 5332 3484
rect 5436 3496 5444 3504
rect 5516 3496 5524 3504
rect 5340 3416 5348 3424
rect 5308 3396 5316 3404
rect 5244 3376 5252 3384
rect 5388 3396 5396 3404
rect 5388 3376 5396 3384
rect 5500 3376 5508 3384
rect 5372 3356 5380 3364
rect 5404 3356 5412 3364
rect 5388 3336 5396 3344
rect 5436 3336 5438 3344
rect 5438 3336 5444 3344
rect 5228 3316 5236 3324
rect 5324 3316 5332 3324
rect 5516 3316 5524 3324
rect 5196 3296 5204 3304
rect 5196 3236 5204 3244
rect 5180 3216 5188 3224
rect 5212 3156 5220 3164
rect 5276 3296 5284 3304
rect 5532 3296 5540 3304
rect 5340 3236 5348 3244
rect 5308 3156 5316 3164
rect 5420 3276 5428 3284
rect 5484 3276 5492 3284
rect 5356 3216 5364 3224
rect 5388 3116 5396 3124
rect 5196 3096 5204 3104
rect 5260 3096 5268 3104
rect 5276 3076 5284 3084
rect 5148 3056 5156 3064
rect 5164 3056 5172 3064
rect 5276 3056 5284 3064
rect 5068 3036 5076 3044
rect 5132 3036 5140 3044
rect 5116 3016 5124 3024
rect 4972 2996 4980 3004
rect 5020 2996 5028 3004
rect 5324 3016 5332 3024
rect 5244 2996 5252 3004
rect 5308 2996 5316 3004
rect 5372 2996 5380 3004
rect 4988 2976 4996 2984
rect 5180 2976 5188 2984
rect 5324 2976 5332 2984
rect 5372 2976 5380 2984
rect 5020 2956 5028 2964
rect 5260 2956 5268 2964
rect 5340 2956 5348 2964
rect 5564 3236 5572 3244
rect 5468 3156 5476 3164
rect 5564 3156 5572 3164
rect 5532 3116 5540 3124
rect 5580 3116 5588 3124
rect 5500 3076 5508 3084
rect 5420 2976 5428 2984
rect 5516 3016 5524 3024
rect 5564 2996 5572 3004
rect 5516 2976 5524 2984
rect 5004 2936 5012 2944
rect 5052 2936 5054 2944
rect 5054 2936 5060 2944
rect 5388 2936 5396 2944
rect 5500 2936 5508 2944
rect 4956 2916 4964 2924
rect 5068 2916 5076 2924
rect 4684 2736 4692 2744
rect 4812 2736 4820 2744
rect 4796 2716 4804 2724
rect 4828 2716 4836 2724
rect 4876 2716 4884 2724
rect 4924 2716 4932 2724
rect 4764 2676 4772 2684
rect 4860 2676 4868 2684
rect 5036 2716 5044 2724
rect 4924 2696 4932 2704
rect 4940 2696 4948 2704
rect 4668 2656 4676 2664
rect 4684 2656 4692 2664
rect 4748 2656 4756 2664
rect 4876 2616 4884 2624
rect 4860 2576 4868 2584
rect 4172 2536 4180 2544
rect 4220 2536 4228 2544
rect 4284 2536 4292 2544
rect 4652 2536 4660 2544
rect 4684 2536 4692 2544
rect 4732 2536 4740 2544
rect 4748 2536 4756 2544
rect 4172 2516 4180 2524
rect 4364 2516 4372 2524
rect 4460 2516 4468 2524
rect 4636 2516 4644 2524
rect 4732 2516 4740 2524
rect 4844 2516 4852 2524
rect 4140 2496 4148 2504
rect 4284 2496 4292 2504
rect 4380 2496 4388 2504
rect 4556 2496 4564 2504
rect 4588 2496 4596 2504
rect 4668 2496 4676 2504
rect 4716 2496 4724 2504
rect 4764 2496 4772 2504
rect 4828 2496 4836 2504
rect 4236 2396 4244 2404
rect 4188 2376 4196 2384
rect 4252 2296 4260 2304
rect 4316 2296 4324 2304
rect 4140 2276 4148 2284
rect 4172 2276 4180 2284
rect 4284 2276 4292 2284
rect 4140 2256 4148 2264
rect 4156 2236 4164 2244
rect 4172 2236 4180 2244
rect 4156 2216 4164 2224
rect 4140 2196 4148 2204
rect 4156 2196 4164 2204
rect 4124 2176 4132 2184
rect 4108 2156 4116 2164
rect 4348 2356 4356 2364
rect 4412 2476 4420 2484
rect 4508 2476 4516 2484
rect 4428 2396 4436 2404
rect 4940 2656 4948 2664
rect 4924 2516 4932 2524
rect 4940 2516 4948 2524
rect 4908 2496 4916 2504
rect 4940 2496 4948 2504
rect 4892 2436 4900 2444
rect 4524 2356 4532 2364
rect 4412 2316 4420 2324
rect 4556 2316 4564 2324
rect 4604 2316 4612 2324
rect 4636 2316 4644 2324
rect 4780 2336 4788 2344
rect 4524 2296 4532 2304
rect 4444 2276 4452 2284
rect 4460 2256 4468 2264
rect 4332 2236 4340 2244
rect 4364 2236 4372 2244
rect 4300 2216 4308 2224
rect 4220 2196 4228 2204
rect 4300 2196 4308 2204
rect 4236 2176 4244 2184
rect 4364 2176 4372 2184
rect 4220 2156 4228 2164
rect 4252 2156 4260 2164
rect 4412 2156 4420 2164
rect 4476 2236 4484 2244
rect 4492 2176 4500 2184
rect 4508 2136 4516 2144
rect 4092 2116 4100 2124
rect 4396 2116 4404 2124
rect 4428 2116 4436 2124
rect 4460 2116 4468 2124
rect 4108 1996 4116 2004
rect 4092 1916 4100 1924
rect 4076 1896 4084 1904
rect 4188 2096 4196 2104
rect 4284 2096 4292 2104
rect 4268 2016 4276 2024
rect 4124 1976 4132 1984
rect 4140 1956 4148 1964
rect 4124 1896 4132 1904
rect 3964 1856 3972 1864
rect 4108 1836 4116 1844
rect 3980 1776 3988 1784
rect 4092 1776 4100 1784
rect 3980 1756 3988 1764
rect 4108 1756 4116 1764
rect 3868 1736 3876 1744
rect 3820 1696 3828 1704
rect 3852 1696 3860 1704
rect 3916 1696 3924 1704
rect 3980 1696 3988 1704
rect 4012 1696 4020 1704
rect 3804 1536 3812 1544
rect 3756 1516 3764 1524
rect 3788 1496 3796 1504
rect 3628 1456 3636 1464
rect 3644 1456 3652 1464
rect 3692 1456 3700 1464
rect 3724 1456 3732 1464
rect 3772 1456 3780 1464
rect 3548 1436 3556 1444
rect 3676 1436 3684 1444
rect 3516 1416 3524 1424
rect 3532 1416 3540 1424
rect 3580 1416 3588 1424
rect 3372 1396 3380 1404
rect 3404 1396 3412 1404
rect 3484 1396 3492 1404
rect 3244 1376 3252 1384
rect 3276 1376 3284 1384
rect 3308 1376 3316 1384
rect 3388 1376 3396 1384
rect 3436 1376 3444 1384
rect 3452 1376 3460 1384
rect 3260 1356 3268 1364
rect 3292 1356 3300 1364
rect 3340 1356 3348 1364
rect 3404 1356 3412 1364
rect 3260 1116 3268 1124
rect 3228 1076 3236 1084
rect 3276 1076 3284 1084
rect 3164 1016 3172 1024
rect 3180 1016 3188 1024
rect 3164 976 3172 984
rect 3276 1016 3284 1024
rect 3260 996 3268 1004
rect 3212 956 3220 964
rect 3276 916 3284 924
rect 3420 1336 3428 1344
rect 3308 1256 3316 1264
rect 3324 1236 3332 1244
rect 3308 1116 3316 1124
rect 3452 1216 3460 1224
rect 3500 1376 3508 1384
rect 3532 1376 3540 1384
rect 3596 1356 3604 1364
rect 3644 1356 3652 1364
rect 3580 1316 3588 1324
rect 3564 1276 3572 1284
rect 3596 1256 3604 1264
rect 3516 1216 3524 1224
rect 3660 1236 3668 1244
rect 3612 1196 3620 1204
rect 3660 1196 3668 1204
rect 3436 1116 3444 1124
rect 3580 1116 3588 1124
rect 3356 1096 3364 1104
rect 3548 1096 3556 1104
rect 3372 1076 3380 1084
rect 3452 1056 3460 1064
rect 3436 996 3444 1004
rect 3324 976 3332 984
rect 3340 956 3348 964
rect 3404 956 3412 964
rect 3468 976 3476 984
rect 3388 936 3396 944
rect 3420 936 3428 944
rect 3452 936 3460 944
rect 3228 896 3236 904
rect 3372 896 3380 904
rect 3292 876 3300 884
rect 3356 876 3364 884
rect 3244 856 3252 864
rect 3244 836 3252 844
rect 3196 816 3204 824
rect 3228 776 3236 784
rect 3164 756 3172 764
rect 3116 736 3124 744
rect 3388 736 3396 744
rect 3164 676 3172 684
rect 3212 676 3220 684
rect 3260 676 3268 684
rect 3100 656 3108 664
rect 3148 656 3156 664
rect 3132 636 3140 644
rect 3116 616 3124 624
rect 3100 576 3108 584
rect 3068 516 3076 524
rect 3036 496 3044 504
rect 3052 496 3060 504
rect 3132 576 3140 584
rect 3148 576 3156 584
rect 3180 576 3188 584
rect 3276 636 3284 644
rect 3356 656 3364 664
rect 3340 636 3348 644
rect 3372 636 3380 644
rect 3244 616 3252 624
rect 3276 616 3284 624
rect 3292 616 3300 624
rect 3324 616 3332 624
rect 3228 556 3236 564
rect 3260 556 3268 564
rect 3116 476 3124 484
rect 3132 476 3140 484
rect 3100 456 3108 464
rect 3132 456 3140 464
rect 3052 376 3060 384
rect 3132 316 3140 324
rect 3164 296 3172 304
rect 2908 256 2916 264
rect 2876 236 2884 244
rect 2956 196 2964 204
rect 2892 176 2900 184
rect 3084 256 3092 264
rect 3020 236 3028 244
rect 3068 236 3076 244
rect 3020 176 3028 184
rect 3100 176 3108 184
rect 3004 156 3012 164
rect 3084 156 3092 164
rect 2812 136 2820 144
rect 2844 136 2852 144
rect 2892 96 2900 104
rect 2940 116 2948 124
rect 2908 36 2916 44
rect 2972 36 2980 44
rect 3036 36 3044 44
rect 2940 16 2948 24
rect 3148 236 3156 244
rect 3388 616 3396 624
rect 3372 576 3380 584
rect 3340 556 3348 564
rect 3356 556 3364 564
rect 3324 536 3332 544
rect 3388 516 3396 524
rect 3292 496 3300 504
rect 3308 496 3316 504
rect 3244 336 3252 344
rect 3340 456 3348 464
rect 3196 256 3204 264
rect 3260 256 3268 264
rect 3148 196 3156 204
rect 3180 196 3188 204
rect 3404 416 3412 424
rect 3356 316 3364 324
rect 3484 836 3492 844
rect 3468 736 3476 744
rect 3516 1036 3524 1044
rect 3532 976 3540 984
rect 3516 876 3524 884
rect 3548 796 3556 804
rect 3516 776 3524 784
rect 3564 776 3572 784
rect 3580 756 3588 764
rect 3500 636 3508 644
rect 3500 596 3508 604
rect 3452 576 3460 584
rect 3436 556 3444 564
rect 3468 556 3476 564
rect 3644 1036 3652 1044
rect 3644 996 3652 1004
rect 3692 1376 3700 1384
rect 3708 1376 3716 1384
rect 3692 1356 3700 1364
rect 3708 1316 3716 1324
rect 3836 1676 3844 1684
rect 3996 1656 4004 1664
rect 3900 1516 3908 1524
rect 3852 1496 3860 1504
rect 3932 1496 3940 1504
rect 3916 1456 3924 1464
rect 3916 1436 3924 1444
rect 3756 1356 3764 1364
rect 3788 1356 3796 1364
rect 3820 1356 3828 1364
rect 3740 1316 3748 1324
rect 3724 1176 3732 1184
rect 3692 1096 3700 1104
rect 3772 1276 3780 1284
rect 3788 1216 3796 1224
rect 3804 1156 3812 1164
rect 3740 1056 3748 1064
rect 3756 1056 3764 1064
rect 3724 1036 3732 1044
rect 3724 996 3732 1004
rect 3676 976 3684 984
rect 3708 976 3716 984
rect 3740 976 3748 984
rect 3644 936 3652 944
rect 3628 816 3636 824
rect 3676 916 3684 924
rect 3708 916 3716 924
rect 3660 776 3668 784
rect 3644 656 3652 664
rect 3660 656 3668 664
rect 3548 576 3556 584
rect 3612 576 3620 584
rect 3484 536 3492 544
rect 3436 516 3444 524
rect 3436 296 3444 304
rect 3500 376 3508 384
rect 3532 296 3540 304
rect 3420 256 3428 264
rect 3292 236 3300 244
rect 3276 216 3284 224
rect 3324 216 3332 224
rect 3388 216 3396 224
rect 3324 176 3332 184
rect 3308 156 3316 164
rect 3404 156 3412 164
rect 3628 556 3636 564
rect 3724 856 3732 864
rect 3724 836 3732 844
rect 3708 716 3716 724
rect 3564 536 3572 544
rect 3644 536 3652 544
rect 3676 536 3684 544
rect 3788 1036 3796 1044
rect 3932 1416 3940 1424
rect 3932 1396 3940 1404
rect 3868 1356 3876 1364
rect 3916 1356 3924 1364
rect 3884 1336 3892 1344
rect 3884 1276 3892 1284
rect 3900 1276 3908 1284
rect 3900 1176 3908 1184
rect 3868 1096 3876 1104
rect 3980 1356 3988 1364
rect 3948 1336 3956 1344
rect 3964 1336 3972 1344
rect 3948 1276 3956 1284
rect 3980 1276 3988 1284
rect 3980 1136 3988 1144
rect 3964 1116 3972 1124
rect 3996 1096 4004 1104
rect 3916 1056 3924 1064
rect 3852 1036 3860 1044
rect 3820 1016 3828 1024
rect 3852 1016 3860 1024
rect 3836 996 3844 1004
rect 3980 996 3988 1004
rect 3836 976 3844 984
rect 3900 976 3908 984
rect 3948 976 3956 984
rect 3820 956 3828 964
rect 3852 956 3860 964
rect 3916 956 3924 964
rect 3772 916 3780 924
rect 3836 916 3844 924
rect 3852 916 3860 924
rect 3884 916 3892 924
rect 3756 896 3764 904
rect 3740 676 3748 684
rect 3692 476 3700 484
rect 3644 416 3652 424
rect 3596 376 3604 384
rect 3740 476 3748 484
rect 3724 296 3732 304
rect 3548 276 3556 284
rect 3596 276 3604 284
rect 3468 236 3476 244
rect 3468 196 3476 204
rect 3516 196 3524 204
rect 3452 156 3460 164
rect 3788 796 3796 804
rect 3772 716 3780 724
rect 3900 756 3908 764
rect 3836 716 3844 724
rect 3788 676 3796 684
rect 3820 676 3828 684
rect 3836 676 3844 684
rect 3868 676 3876 684
rect 3884 676 3892 684
rect 3804 636 3812 644
rect 3804 596 3812 604
rect 3836 596 3844 604
rect 3788 576 3796 584
rect 3932 636 3940 644
rect 3916 616 3924 624
rect 4156 1876 4158 1884
rect 4158 1876 4164 1884
rect 4300 1996 4308 2004
rect 4284 1956 4292 1964
rect 4364 1936 4372 1944
rect 4204 1916 4212 1924
rect 4252 1916 4260 1924
rect 4300 1916 4308 1924
rect 4380 1916 4388 1924
rect 4428 1916 4436 1924
rect 4476 1916 4484 1924
rect 4492 1896 4500 1904
rect 4556 2276 4564 2284
rect 4572 2276 4580 2284
rect 4620 2176 4628 2184
rect 4780 2216 4788 2224
rect 4812 2216 4820 2224
rect 4684 2176 4692 2184
rect 4828 2156 4836 2164
rect 4892 2376 4900 2384
rect 4876 2336 4884 2344
rect 4876 2196 4884 2204
rect 4972 2536 4980 2544
rect 5068 2616 5076 2624
rect 5100 2696 5108 2704
rect 5148 2876 5156 2884
rect 5244 2916 5252 2924
rect 5196 2836 5204 2844
rect 5212 2816 5220 2824
rect 5244 2816 5252 2824
rect 5116 2676 5124 2684
rect 5132 2676 5140 2684
rect 5132 2636 5140 2644
rect 5116 2616 5124 2624
rect 5052 2596 5060 2604
rect 5084 2596 5092 2604
rect 5260 2776 5268 2784
rect 5244 2696 5252 2704
rect 5260 2656 5268 2664
rect 5180 2596 5188 2604
rect 5212 2596 5220 2604
rect 5452 2916 5460 2924
rect 5404 2876 5412 2884
rect 5340 2736 5348 2744
rect 5324 2696 5332 2704
rect 5292 2656 5300 2664
rect 5276 2636 5284 2644
rect 5276 2596 5284 2604
rect 5308 2596 5316 2604
rect 5148 2556 5156 2564
rect 5228 2556 5236 2564
rect 5260 2556 5268 2564
rect 5132 2536 5140 2544
rect 5196 2536 5204 2544
rect 5004 2516 5012 2524
rect 5036 2516 5044 2524
rect 5068 2516 5076 2524
rect 5228 2516 5236 2524
rect 5148 2496 5156 2504
rect 4956 2476 4964 2484
rect 5020 2376 5028 2384
rect 5020 2336 5028 2344
rect 5004 2316 5012 2324
rect 4908 2256 4916 2264
rect 4940 2256 4948 2264
rect 4556 2136 4564 2144
rect 4588 2136 4596 2144
rect 4748 2136 4756 2144
rect 4844 2136 4852 2144
rect 4556 2116 4564 2124
rect 4604 2116 4612 2124
rect 4684 2116 4692 2124
rect 4860 2116 4868 2124
rect 4892 2116 4900 2124
rect 4620 2096 4628 2104
rect 4652 2096 4660 2104
rect 4604 1916 4612 1924
rect 4236 1876 4244 1884
rect 4316 1876 4324 1884
rect 4396 1876 4404 1884
rect 4460 1876 4468 1884
rect 4188 1836 4196 1844
rect 4156 1736 4164 1744
rect 4060 1676 4068 1684
rect 4044 1596 4052 1604
rect 4220 1796 4228 1804
rect 4364 1796 4372 1804
rect 4412 1796 4420 1804
rect 4300 1776 4308 1784
rect 4332 1776 4340 1784
rect 4476 1736 4484 1744
rect 4316 1716 4324 1724
rect 4172 1676 4180 1684
rect 4204 1676 4212 1684
rect 4316 1676 4324 1684
rect 4348 1676 4356 1684
rect 4412 1676 4420 1684
rect 4284 1656 4292 1664
rect 4268 1596 4276 1604
rect 4364 1596 4372 1604
rect 4348 1576 4356 1584
rect 4492 1576 4500 1584
rect 4028 1536 4036 1544
rect 4140 1536 4148 1544
rect 4172 1536 4180 1544
rect 4252 1536 4260 1544
rect 4044 1516 4052 1524
rect 4140 1516 4148 1524
rect 4156 1516 4164 1524
rect 4092 1496 4100 1504
rect 4412 1516 4420 1524
rect 4476 1496 4484 1504
rect 4236 1476 4244 1484
rect 4076 1456 4084 1464
rect 4092 1456 4100 1464
rect 4172 1456 4180 1464
rect 4188 1456 4196 1464
rect 4204 1456 4212 1464
rect 4044 1396 4052 1404
rect 4108 1396 4116 1404
rect 4028 1356 4036 1364
rect 4092 1356 4100 1364
rect 4156 1356 4164 1364
rect 4124 1336 4132 1344
rect 4124 1316 4132 1324
rect 4076 1276 4084 1284
rect 4060 1236 4068 1244
rect 4060 1096 4068 1104
rect 4012 1056 4020 1064
rect 4028 1036 4036 1044
rect 4044 956 4052 964
rect 4012 916 4020 924
rect 4060 876 4068 884
rect 4028 796 4036 804
rect 4044 756 4052 764
rect 3964 676 3966 684
rect 3966 676 3972 684
rect 3964 656 3972 664
rect 3996 656 4004 664
rect 4060 656 4068 664
rect 4140 1276 4148 1284
rect 4172 1316 4180 1324
rect 4092 1116 4100 1124
rect 4140 1116 4148 1124
rect 4156 1096 4164 1104
rect 4236 1436 4244 1444
rect 4220 1396 4228 1404
rect 4236 1356 4244 1364
rect 4236 1336 4244 1344
rect 4236 1296 4244 1304
rect 4252 1296 4260 1304
rect 4460 1476 4468 1484
rect 4396 1436 4404 1444
rect 4380 1336 4388 1344
rect 4284 1316 4292 1324
rect 4364 1316 4372 1324
rect 4300 1296 4308 1304
rect 4268 1276 4276 1284
rect 4364 1276 4372 1284
rect 4332 1136 4340 1144
rect 4348 1116 4356 1124
rect 4428 1316 4436 1324
rect 4428 1156 4436 1164
rect 4636 2076 4644 2084
rect 4652 2036 4660 2044
rect 4636 1896 4644 1904
rect 4572 1856 4580 1864
rect 4540 1836 4548 1844
rect 4572 1836 4580 1844
rect 4620 1836 4628 1844
rect 4556 1676 4564 1684
rect 4524 1656 4532 1664
rect 4524 1576 4532 1584
rect 4540 1576 4548 1584
rect 4556 1516 4564 1524
rect 4508 1456 4516 1464
rect 4476 1376 4484 1384
rect 4540 1376 4548 1384
rect 4556 1336 4564 1344
rect 4476 1316 4484 1324
rect 4508 1296 4516 1304
rect 4476 1216 4484 1224
rect 4236 1096 4244 1104
rect 4268 1096 4276 1104
rect 4140 1076 4148 1084
rect 4124 1036 4132 1044
rect 4092 1016 4100 1024
rect 4108 956 4116 964
rect 4108 736 4116 744
rect 4124 736 4132 744
rect 4092 656 4100 664
rect 4108 656 4116 664
rect 3980 596 3988 604
rect 3996 596 4004 604
rect 4012 596 4020 604
rect 4044 596 4052 604
rect 3868 516 3876 524
rect 3916 416 3924 424
rect 3916 376 3924 384
rect 3900 356 3908 364
rect 3852 316 3860 324
rect 3868 316 3876 324
rect 3804 296 3812 304
rect 3836 296 3844 304
rect 3676 256 3684 264
rect 3788 236 3796 244
rect 3612 216 3620 224
rect 3660 216 3668 224
rect 3772 196 3780 204
rect 3596 176 3604 184
rect 3660 176 3668 184
rect 3756 176 3764 184
rect 3916 336 3924 344
rect 3932 316 3940 324
rect 3964 316 3972 324
rect 4156 836 4164 844
rect 4156 816 4164 824
rect 4172 776 4180 784
rect 4172 756 4180 764
rect 4364 1036 4372 1044
rect 4220 996 4228 1004
rect 4236 996 4244 1004
rect 4364 996 4372 1004
rect 4412 1076 4420 1084
rect 4412 1056 4420 1064
rect 4316 956 4324 964
rect 4364 956 4372 964
rect 4396 956 4404 964
rect 4236 916 4244 924
rect 4252 916 4260 924
rect 4220 876 4228 884
rect 4252 856 4260 864
rect 4268 856 4276 864
rect 4300 836 4308 844
rect 4252 736 4260 744
rect 4188 696 4196 704
rect 4204 696 4212 704
rect 4204 656 4212 664
rect 4156 616 4164 624
rect 4236 596 4244 604
rect 4172 576 4180 584
rect 4188 576 4196 584
rect 4220 576 4228 584
rect 4060 516 4068 524
rect 4108 516 4116 524
rect 4140 516 4148 524
rect 4124 436 4132 444
rect 4060 296 4068 304
rect 3996 276 4004 284
rect 4428 976 4436 984
rect 4492 1076 4500 1084
rect 4540 1076 4542 1084
rect 4542 1076 4548 1084
rect 4476 1056 4484 1064
rect 4524 1056 4532 1064
rect 4508 976 4516 984
rect 4332 936 4340 944
rect 4444 936 4452 944
rect 4508 936 4516 944
rect 4396 876 4404 884
rect 4476 836 4484 844
rect 4412 816 4420 824
rect 4396 776 4404 784
rect 4300 716 4308 724
rect 4284 696 4292 704
rect 4300 696 4308 704
rect 4380 696 4388 704
rect 4300 616 4308 624
rect 4252 496 4260 504
rect 4268 496 4276 504
rect 4220 376 4228 384
rect 4236 356 4244 364
rect 4300 496 4308 504
rect 4364 596 4372 604
rect 4348 576 4356 584
rect 4460 756 4468 764
rect 4508 736 4516 744
rect 4492 716 4500 724
rect 4428 616 4436 624
rect 4556 996 4564 1004
rect 4620 1796 4628 1804
rect 4604 1756 4612 1764
rect 4636 1756 4644 1764
rect 4588 1696 4596 1704
rect 4636 1576 4644 1584
rect 4620 1516 4628 1524
rect 4588 1456 4596 1464
rect 4604 1456 4612 1464
rect 4636 1416 4644 1424
rect 4620 1356 4628 1364
rect 4604 1316 4612 1324
rect 4588 1156 4596 1164
rect 4604 1156 4612 1164
rect 4588 1116 4596 1124
rect 4620 1116 4628 1124
rect 4636 1076 4644 1084
rect 4604 1036 4612 1044
rect 4620 956 4628 964
rect 4556 796 4564 804
rect 4556 756 4564 764
rect 4572 756 4580 764
rect 4364 556 4372 564
rect 4396 556 4404 564
rect 4412 556 4420 564
rect 4476 556 4484 564
rect 4492 496 4500 504
rect 4412 476 4420 484
rect 4332 396 4340 404
rect 4284 376 4292 384
rect 4348 376 4356 384
rect 4460 376 4468 384
rect 4364 356 4372 364
rect 4156 296 4164 304
rect 4172 296 4180 304
rect 4284 296 4292 304
rect 4044 276 4052 284
rect 4108 276 4116 284
rect 4140 276 4148 284
rect 4204 276 4212 284
rect 4236 276 4244 284
rect 4300 276 4308 284
rect 4348 276 4356 284
rect 4012 256 4020 264
rect 4044 256 4052 264
rect 4188 236 4196 244
rect 3788 176 3796 184
rect 3804 176 3812 184
rect 3900 176 3908 184
rect 3964 176 3972 184
rect 4108 216 4116 224
rect 4092 196 4100 204
rect 3948 156 3956 164
rect 3996 156 4004 164
rect 4044 156 4052 164
rect 4172 176 4180 184
rect 4220 176 4228 184
rect 4380 296 4388 304
rect 4460 336 4468 344
rect 4476 296 4484 304
rect 4492 296 4500 304
rect 4412 276 4420 284
rect 4540 616 4548 624
rect 4556 596 4564 604
rect 4668 1956 4676 1964
rect 4764 1956 4772 1964
rect 4732 1936 4740 1944
rect 4748 1916 4756 1924
rect 4716 1896 4724 1904
rect 4812 1896 4820 1904
rect 4700 1876 4708 1884
rect 4684 1856 4692 1864
rect 4700 1736 4708 1744
rect 4684 1676 4692 1684
rect 4684 1656 4692 1664
rect 4700 1516 4708 1524
rect 4940 2196 4948 2204
rect 5212 2476 5220 2484
rect 5180 2396 5188 2404
rect 5132 2356 5140 2364
rect 5100 2316 5108 2324
rect 5084 2276 5092 2284
rect 5068 2256 5076 2264
rect 4988 2196 4996 2204
rect 5036 2196 5044 2204
rect 4988 2136 4996 2144
rect 5004 2136 5012 2144
rect 5148 2336 5156 2344
rect 5212 2336 5220 2344
rect 5196 2316 5204 2324
rect 5212 2316 5220 2324
rect 5100 2216 5108 2224
rect 5084 2196 5092 2204
rect 5052 2136 5060 2144
rect 5116 2136 5124 2144
rect 5196 2176 5204 2184
rect 5212 2156 5220 2164
rect 5068 2116 5076 2124
rect 5084 2116 5092 2124
rect 5132 2116 5140 2124
rect 5164 2116 5172 2124
rect 4924 2096 4932 2104
rect 4956 2096 4964 2104
rect 5004 2096 5012 2104
rect 5020 2096 5028 2104
rect 5084 2096 5092 2104
rect 4924 1976 4932 1984
rect 4844 1916 4852 1924
rect 4732 1856 4740 1864
rect 4780 1816 4788 1824
rect 4748 1676 4756 1684
rect 4732 1636 4740 1644
rect 4764 1596 4772 1604
rect 4732 1556 4740 1564
rect 4748 1516 4756 1524
rect 4828 1816 4836 1824
rect 4876 1816 4884 1824
rect 4876 1776 4884 1784
rect 4908 1916 4916 1924
rect 4988 1976 4996 1984
rect 4972 1956 4980 1964
rect 4956 1936 4964 1944
rect 4956 1916 4964 1924
rect 5052 1936 5060 1944
rect 5148 2056 5156 2064
rect 5132 1956 5140 1964
rect 5164 1936 5172 1944
rect 5068 1916 5076 1924
rect 5004 1876 5012 1884
rect 5036 1876 5044 1884
rect 5084 1876 5092 1884
rect 5292 2576 5300 2584
rect 5324 2576 5332 2584
rect 5260 2476 5268 2484
rect 5244 2436 5252 2444
rect 5276 2436 5284 2444
rect 5244 2416 5252 2424
rect 5260 2356 5268 2364
rect 5260 2136 5266 2144
rect 5266 2136 5268 2144
rect 5244 2096 5252 2104
rect 5308 2556 5316 2564
rect 5340 2516 5348 2524
rect 5324 2316 5332 2324
rect 5404 2736 5412 2744
rect 5452 2716 5460 2724
rect 5516 2716 5524 2724
rect 5372 2696 5380 2704
rect 5452 2696 5460 2704
rect 5468 2696 5476 2704
rect 5516 2696 5524 2704
rect 5372 2676 5380 2684
rect 5436 2596 5444 2604
rect 5564 2616 5572 2624
rect 5532 2596 5540 2604
rect 5388 2536 5396 2544
rect 5452 2536 5460 2544
rect 5500 2536 5508 2544
rect 5516 2536 5524 2544
rect 5580 2536 5588 2544
rect 5372 2496 5380 2504
rect 5500 2496 5508 2504
rect 5388 2476 5396 2484
rect 5532 2456 5540 2464
rect 5468 2396 5476 2404
rect 5500 2396 5508 2404
rect 5468 2316 5476 2324
rect 5500 2316 5508 2324
rect 5356 2296 5364 2304
rect 5308 2236 5316 2244
rect 5324 2196 5332 2204
rect 5308 2176 5316 2184
rect 5276 1936 5284 1944
rect 4892 1756 4900 1764
rect 4988 1796 4996 1804
rect 4988 1756 4996 1764
rect 5068 1756 5076 1764
rect 5004 1716 5012 1724
rect 5036 1716 5044 1724
rect 4812 1676 4820 1684
rect 4796 1656 4804 1664
rect 4796 1576 4804 1584
rect 4796 1516 4804 1524
rect 4732 1436 4740 1444
rect 4812 1436 4820 1444
rect 4828 1416 4836 1424
rect 4924 1696 4932 1704
rect 4956 1696 4964 1704
rect 4860 1596 4868 1604
rect 4924 1596 4932 1604
rect 4860 1576 4868 1584
rect 4876 1536 4884 1544
rect 4876 1496 4884 1504
rect 4988 1576 4996 1584
rect 4956 1536 4964 1544
rect 4972 1496 4980 1504
rect 5004 1556 5012 1564
rect 5020 1556 5028 1564
rect 4844 1376 4852 1384
rect 4780 1356 4788 1364
rect 4860 1356 4868 1364
rect 4988 1416 4996 1424
rect 4924 1376 4932 1384
rect 4908 1356 4916 1364
rect 4956 1356 4964 1364
rect 4796 1336 4804 1344
rect 4844 1336 4852 1344
rect 4668 1296 4676 1304
rect 4748 1296 4756 1304
rect 4716 1196 4724 1204
rect 4684 1116 4692 1124
rect 4732 1116 4740 1124
rect 4764 1116 4772 1124
rect 4828 1276 4836 1284
rect 4812 1236 4820 1244
rect 4828 1116 4836 1124
rect 4876 1156 4884 1164
rect 4876 1116 4884 1124
rect 4844 1096 4852 1104
rect 4860 1096 4868 1104
rect 4780 1076 4788 1084
rect 4652 1036 4660 1044
rect 4652 996 4660 1004
rect 4748 1016 4756 1024
rect 4684 996 4692 1004
rect 4700 996 4708 1004
rect 4732 996 4740 1004
rect 4620 756 4628 764
rect 4604 596 4612 604
rect 4876 996 4884 1004
rect 4812 896 4820 904
rect 4812 856 4820 864
rect 4908 1116 4916 1124
rect 4940 1036 4948 1044
rect 4908 996 4916 1004
rect 4924 996 4932 1004
rect 5228 1856 5236 1864
rect 5180 1836 5188 1844
rect 5196 1836 5204 1844
rect 5132 1776 5140 1784
rect 5052 1696 5060 1704
rect 5116 1556 5124 1564
rect 5100 1536 5108 1544
rect 5148 1736 5156 1744
rect 5196 1616 5204 1624
rect 5180 1536 5188 1544
rect 5084 1496 5092 1504
rect 5116 1496 5124 1504
rect 5164 1476 5172 1484
rect 5196 1476 5204 1484
rect 5116 1396 5124 1404
rect 5052 1356 5060 1364
rect 5068 1356 5076 1364
rect 5132 1356 5140 1364
rect 5052 1296 5060 1304
rect 5084 1276 5092 1284
rect 5068 1176 5076 1184
rect 5084 1176 5092 1184
rect 5052 1136 5060 1144
rect 4988 1116 4996 1124
rect 5020 1116 5028 1124
rect 5004 1096 5012 1104
rect 5148 1096 5156 1104
rect 5132 1076 5140 1084
rect 5084 1056 5092 1064
rect 5068 1036 5076 1044
rect 5036 956 5044 964
rect 5052 956 5060 964
rect 5148 1036 5156 1044
rect 5132 976 5140 984
rect 5100 956 5108 964
rect 5116 956 5124 964
rect 4892 836 4900 844
rect 4828 816 4836 824
rect 4652 776 4660 784
rect 4732 756 4740 764
rect 4812 756 4820 764
rect 4668 736 4676 744
rect 4748 736 4756 744
rect 4764 736 4772 744
rect 4780 736 4788 744
rect 4700 716 4708 724
rect 4684 696 4692 704
rect 4844 776 4852 784
rect 4876 756 4884 764
rect 4844 676 4852 684
rect 4860 676 4868 684
rect 4668 596 4676 604
rect 4796 596 4804 604
rect 4604 576 4612 584
rect 4636 576 4644 584
rect 4588 556 4596 564
rect 4524 536 4532 544
rect 4700 556 4708 564
rect 4732 556 4740 564
rect 4652 536 4660 544
rect 4684 536 4690 544
rect 4690 536 4692 544
rect 4588 476 4596 484
rect 4636 316 4644 324
rect 4572 296 4580 304
rect 4684 316 4692 324
rect 4652 276 4660 284
rect 4604 216 4612 224
rect 4508 176 4516 184
rect 4668 176 4676 184
rect 4252 156 4260 164
rect 3452 136 3460 144
rect 3484 136 3492 144
rect 3532 136 3540 144
rect 3596 136 3604 144
rect 3612 136 3620 144
rect 4204 136 4212 144
rect 4332 136 4340 144
rect 4444 136 4452 144
rect 3292 116 3300 124
rect 3340 116 3348 124
rect 3404 116 3412 124
rect 4332 116 4340 124
rect 4380 116 4388 124
rect 4892 696 4900 704
rect 4956 896 4964 904
rect 4940 876 4948 884
rect 4940 676 4948 684
rect 4908 596 4916 604
rect 4860 576 4868 584
rect 4892 576 4900 584
rect 4732 536 4740 544
rect 4716 516 4724 524
rect 4764 496 4772 504
rect 4812 496 4820 504
rect 4732 396 4740 404
rect 4716 316 4724 324
rect 4796 376 4804 384
rect 4764 356 4772 364
rect 4732 216 4740 224
rect 4812 296 4820 304
rect 4844 296 4852 304
rect 4764 216 4772 224
rect 5052 936 5060 944
rect 5004 896 5012 904
rect 5036 736 5044 744
rect 5052 676 5060 684
rect 5084 656 5092 664
rect 5068 636 5076 644
rect 4988 596 4996 604
rect 5004 596 5012 604
rect 5052 596 5060 604
rect 5068 596 5076 604
rect 4988 576 4996 584
rect 5036 576 5044 584
rect 4972 536 4980 544
rect 5084 536 5092 544
rect 4908 496 4916 504
rect 4924 456 4932 464
rect 4940 376 4948 384
rect 4892 336 4900 344
rect 5036 516 5044 524
rect 5116 896 5124 904
rect 5132 716 5140 724
rect 5196 1456 5204 1464
rect 5180 1436 5188 1444
rect 5196 1356 5204 1364
rect 5196 1296 5204 1304
rect 5180 1196 5188 1204
rect 5212 1136 5220 1144
rect 5180 1096 5188 1104
rect 5388 2256 5396 2264
rect 5372 2236 5380 2244
rect 5548 2296 5556 2304
rect 5564 2276 5572 2284
rect 5484 2236 5492 2244
rect 5404 2176 5412 2184
rect 5388 2156 5396 2164
rect 5372 2136 5380 2144
rect 5340 2076 5348 2084
rect 5404 2076 5412 2084
rect 5356 2036 5364 2044
rect 5452 2196 5460 2204
rect 5452 2136 5460 2144
rect 5468 2076 5476 2084
rect 5436 1996 5444 2004
rect 5340 1936 5348 1944
rect 5420 1936 5428 1944
rect 5372 1916 5380 1924
rect 5292 1896 5300 1904
rect 5468 1916 5476 1924
rect 5292 1876 5300 1884
rect 5404 1876 5412 1884
rect 5244 1796 5252 1804
rect 5276 1796 5284 1804
rect 5436 1796 5444 1804
rect 5276 1776 5284 1784
rect 5260 1756 5268 1764
rect 5372 1756 5380 1764
rect 5500 2196 5508 2204
rect 5564 2176 5572 2184
rect 5516 2136 5524 2144
rect 5516 2096 5524 2104
rect 5500 1876 5508 1884
rect 5564 1816 5572 1824
rect 5532 1796 5540 1804
rect 5564 1796 5572 1804
rect 5500 1756 5508 1764
rect 5292 1736 5300 1744
rect 5388 1736 5396 1744
rect 5324 1716 5332 1724
rect 5292 1696 5300 1704
rect 5356 1576 5364 1584
rect 5388 1576 5396 1584
rect 5276 1516 5284 1524
rect 5244 1496 5252 1504
rect 5244 1376 5252 1384
rect 5324 1516 5332 1524
rect 5308 1436 5316 1444
rect 5260 1336 5268 1344
rect 5276 1316 5284 1324
rect 5260 1096 5268 1104
rect 5196 1076 5204 1084
rect 5228 1076 5236 1084
rect 5276 1056 5284 1064
rect 5244 996 5252 1004
rect 5180 936 5188 944
rect 5164 876 5172 884
rect 5148 696 5156 704
rect 5132 676 5140 684
rect 5132 616 5140 624
rect 5212 896 5220 904
rect 5276 876 5284 884
rect 5196 836 5204 844
rect 5260 756 5268 764
rect 5196 736 5204 744
rect 5244 736 5252 744
rect 5324 1376 5332 1384
rect 5340 1376 5348 1384
rect 5308 1356 5316 1364
rect 5324 1316 5332 1324
rect 5308 1296 5316 1304
rect 5372 1516 5380 1524
rect 5372 1376 5380 1384
rect 5420 1536 5428 1544
rect 5532 1596 5540 1604
rect 5452 1516 5460 1524
rect 5532 1496 5540 1504
rect 5404 1376 5412 1384
rect 5452 1376 5460 1384
rect 5404 1336 5412 1344
rect 5500 1336 5508 1344
rect 5484 1296 5492 1304
rect 5388 1276 5396 1284
rect 5324 1156 5332 1164
rect 5308 1136 5316 1144
rect 5388 1196 5396 1204
rect 5420 1136 5428 1144
rect 5436 1096 5444 1104
rect 5468 1076 5476 1084
rect 5452 1036 5460 1044
rect 5340 1016 5348 1024
rect 5308 896 5316 904
rect 5292 716 5300 724
rect 5292 696 5300 704
rect 5356 976 5364 984
rect 5436 996 5444 1004
rect 5452 976 5460 984
rect 5372 956 5380 964
rect 5500 936 5508 944
rect 5388 916 5396 924
rect 5404 916 5412 924
rect 5356 896 5364 904
rect 5484 896 5492 904
rect 5356 736 5364 744
rect 5372 736 5380 744
rect 5500 736 5508 744
rect 5196 676 5204 684
rect 5308 676 5316 684
rect 5164 596 5172 604
rect 5164 576 5172 584
rect 5196 556 5204 564
rect 5292 556 5300 564
rect 5148 536 5156 544
rect 5212 536 5220 544
rect 5276 536 5284 544
rect 5356 676 5364 684
rect 5388 656 5396 664
rect 5452 696 5460 704
rect 5404 636 5412 644
rect 5388 596 5396 604
rect 5372 576 5380 584
rect 5420 556 5428 564
rect 5180 516 5188 524
rect 5260 516 5268 524
rect 5116 496 5124 504
rect 5164 496 5172 504
rect 5260 496 5268 504
rect 5244 476 5252 484
rect 5116 456 5124 464
rect 4924 296 4932 304
rect 5036 296 5044 304
rect 5132 376 5140 384
rect 5212 376 5220 384
rect 4860 256 4868 264
rect 4876 256 4884 264
rect 4924 256 4932 264
rect 4796 216 4804 224
rect 4780 196 4788 204
rect 4748 176 4756 184
rect 4940 216 4948 224
rect 5068 216 5076 224
rect 5052 196 5060 204
rect 4716 156 4724 164
rect 4908 156 4916 164
rect 4988 156 4996 164
rect 4972 136 4980 144
rect 5004 136 5012 144
rect 4588 116 4596 124
rect 4604 116 4612 124
rect 4668 116 4676 124
rect 4700 116 4708 124
rect 4748 116 4756 124
rect 4764 116 4772 124
rect 4812 116 4820 124
rect 4844 116 4852 124
rect 4940 116 4948 124
rect 5020 116 5028 124
rect 5164 296 5172 304
rect 5180 256 5188 264
rect 5116 236 5124 244
rect 5116 216 5124 224
rect 5196 216 5204 224
rect 5180 196 5188 204
rect 5132 176 5140 184
rect 5164 156 5172 164
rect 5324 516 5332 524
rect 5404 536 5412 544
rect 5372 356 5380 364
rect 5388 336 5396 344
rect 5468 596 5476 604
rect 5500 596 5508 604
rect 5452 516 5460 524
rect 5452 496 5460 504
rect 5436 456 5444 464
rect 5436 436 5444 444
rect 5228 316 5236 324
rect 5292 316 5300 324
rect 5308 316 5316 324
rect 5356 316 5364 324
rect 5244 296 5252 304
rect 5308 296 5316 304
rect 5324 276 5332 284
rect 5340 276 5348 284
rect 5244 216 5252 224
rect 5260 176 5268 184
rect 5308 176 5316 184
rect 5324 156 5332 164
rect 5468 476 5476 484
rect 5500 256 5508 264
rect 5436 236 5444 244
rect 5452 236 5460 244
rect 5436 196 5444 204
rect 5356 176 5364 184
rect 5436 136 5444 144
rect 5564 376 5572 384
rect 5580 176 5588 184
rect 5516 116 5524 124
rect 3132 96 3140 104
rect 4028 96 4036 104
rect 4092 96 4100 104
rect 4108 96 4116 104
rect 4172 96 4180 104
rect 4284 96 4292 104
rect 4316 96 4324 104
rect 4364 96 4372 104
rect 4412 96 4420 104
rect 4540 96 4548 104
rect 4652 96 4660 104
rect 5404 96 5412 104
rect 3452 76 3460 84
rect 3564 76 3572 84
rect 3644 76 3652 84
rect 3692 76 3700 84
rect 3836 76 3844 84
rect 3884 76 3892 84
rect 5276 76 5284 84
rect 5468 76 5476 84
rect 4620 56 4628 64
rect 3852 36 3860 44
rect 4556 36 4564 44
rect 4700 16 4708 24
<< metal3 >>
rect 1204 3997 1740 4003
rect 516 3977 604 3983
rect 1117 3977 1612 3983
rect 196 3957 252 3963
rect 868 3957 924 3963
rect 1117 3963 1123 3977
rect 1796 3977 2012 3983
rect 2685 3964 2691 3976
rect 932 3957 1123 3963
rect 1492 3957 1804 3963
rect 1860 3957 2028 3963
rect 2100 3957 2380 3963
rect 3300 3957 4300 3963
rect 4308 3957 4764 3963
rect 1524 3937 1596 3943
rect 1604 3937 1708 3943
rect 1716 3937 1852 3943
rect 2020 3937 2092 3943
rect 2164 3937 2508 3943
rect 2516 3937 2652 3943
rect 2660 3937 2700 3943
rect 3396 3937 3612 3943
rect 3652 3937 3948 3943
rect 3972 3937 4060 3943
rect 4164 3937 4252 3943
rect 4356 3937 4396 3943
rect 4964 3937 5068 3943
rect 228 3917 268 3923
rect 388 3917 1036 3923
rect 1444 3917 1484 3923
rect 1588 3917 1644 3923
rect 1780 3917 1852 3923
rect 1860 3917 1916 3923
rect 1972 3917 2316 3923
rect 2324 3917 2332 3923
rect 2436 3917 2492 3923
rect 2564 3917 2828 3923
rect 3140 3917 3180 3923
rect 3268 3917 3276 3923
rect 3476 3917 3788 3923
rect 3828 3917 3836 3923
rect 4052 3917 4172 3923
rect 4196 3917 4236 3923
rect 4244 3917 4524 3923
rect 4644 3917 4684 3923
rect 4708 3917 4723 3923
rect 4740 3917 4924 3923
rect 4932 3917 5004 3923
rect 5204 3917 5292 3923
rect 5469 3904 5475 3916
rect 260 3897 364 3903
rect 692 3897 1068 3903
rect 1236 3897 1308 3903
rect 1668 3897 1900 3903
rect 1908 3897 2284 3903
rect 2372 3897 2380 3903
rect 2404 3897 2460 3903
rect 2468 3897 2716 3903
rect 2724 3897 2972 3903
rect 3012 3897 3084 3903
rect 3156 3897 3164 3903
rect 3204 3897 3260 3903
rect 3268 3897 3340 3903
rect 3460 3897 3548 3903
rect 3652 3897 3708 3903
rect 3725 3897 3740 3903
rect 3764 3897 4460 3903
rect 4500 3897 4556 3903
rect 5156 3897 5324 3903
rect 148 3877 284 3883
rect 308 3877 524 3883
rect 580 3877 700 3883
rect 756 3877 764 3883
rect 820 3877 828 3883
rect 852 3877 860 3883
rect 900 3877 988 3883
rect 1028 3877 1068 3883
rect 1284 3877 1340 3883
rect 1396 3877 1404 3883
rect 1924 3877 1964 3883
rect 1972 3877 1980 3883
rect 1988 3877 2092 3883
rect 2116 3877 2188 3883
rect 2196 3877 2396 3883
rect 2420 3877 2460 3883
rect 2500 3877 2636 3883
rect 2772 3877 2860 3883
rect 2964 3877 3468 3883
rect 3700 3877 3756 3883
rect 3796 3877 3804 3883
rect 3876 3877 3891 3883
rect 4116 3877 4892 3883
rect 5140 3877 5212 3883
rect 5300 3877 5324 3883
rect 5364 3877 5388 3883
rect 1213 3864 1219 3876
rect 36 3857 908 3863
rect 980 3857 988 3863
rect 1540 3857 1996 3863
rect 2004 3857 2172 3863
rect 2180 3857 2188 3863
rect 2292 3857 2300 3863
rect 2308 3857 2444 3863
rect 2452 3857 2572 3863
rect 2836 3857 3020 3863
rect 3076 3857 3420 3863
rect 3428 3857 3500 3863
rect 3508 3857 3996 3863
rect 4004 3857 4316 3863
rect 4333 3857 4748 3863
rect 20 3837 108 3843
rect 260 3837 396 3843
rect 436 3837 460 3843
rect 756 3837 764 3843
rect 2260 3837 2284 3843
rect 2340 3837 2556 3843
rect 2564 3837 2588 3843
rect 2804 3837 2956 3843
rect 2964 3837 3036 3843
rect 3044 3837 3084 3843
rect 3108 3837 3404 3843
rect 3412 3837 3564 3843
rect 3572 3837 3804 3843
rect 4333 3843 4339 3857
rect 4772 3857 4940 3863
rect 5124 3857 5132 3863
rect 5309 3844 5315 3856
rect 3812 3837 4339 3843
rect 1140 3817 1628 3823
rect 2036 3817 2044 3823
rect 2388 3817 2428 3823
rect 2596 3817 3372 3823
rect 3380 3817 3436 3823
rect 4180 3817 4300 3823
rect 4420 3817 4524 3823
rect 4548 3817 5196 3823
rect 5252 3817 5260 3823
rect 196 3797 588 3803
rect 1092 3797 1100 3803
rect 1300 3797 1324 3803
rect 1492 3797 1500 3803
rect 1556 3797 1564 3803
rect 1732 3797 1852 3803
rect 1860 3797 2172 3803
rect 2180 3797 2236 3803
rect 2404 3797 2444 3803
rect 2500 3797 2588 3803
rect 2660 3797 2812 3803
rect 2820 3797 2860 3803
rect 2868 3797 2892 3803
rect 2900 3797 2956 3803
rect 2980 3797 3212 3803
rect 3252 3797 3260 3803
rect 3268 3797 3452 3803
rect 3780 3797 3788 3803
rect 4036 3797 4044 3803
rect 4084 3797 4092 3803
rect 4116 3797 4156 3803
rect 4228 3797 4236 3803
rect 4484 3797 4572 3803
rect 4676 3797 4684 3803
rect 5060 3797 5068 3803
rect 5108 3797 5132 3803
rect 5252 3797 5308 3803
rect 5428 3797 5436 3803
rect 1613 3784 1619 3796
rect 532 3777 540 3783
rect 580 3777 828 3783
rect 916 3777 1132 3783
rect 1140 3777 1420 3783
rect 1428 3777 1596 3783
rect 1636 3777 1724 3783
rect 1796 3777 1868 3783
rect 1940 3777 1948 3783
rect 2196 3777 2524 3783
rect 2532 3777 2588 3783
rect 2884 3777 3068 3783
rect 3076 3777 3644 3783
rect 3652 3777 4108 3783
rect 4180 3777 4748 3783
rect 4820 3777 4876 3783
rect 4948 3777 5260 3783
rect 5444 3777 5452 3783
rect 253 3764 259 3776
rect 68 3757 76 3763
rect 388 3757 876 3763
rect 900 3757 908 3763
rect 964 3757 1020 3763
rect 1028 3757 1676 3763
rect 1812 3757 1884 3763
rect 1908 3757 2316 3763
rect 2436 3757 2572 3763
rect 2596 3757 2700 3763
rect 2708 3757 2764 3763
rect 2772 3757 2844 3763
rect 2852 3757 2876 3763
rect 2964 3757 2972 3763
rect 2996 3757 3036 3763
rect 3044 3757 3100 3763
rect 3108 3757 3164 3763
rect 3220 3757 3340 3763
rect 3396 3757 3468 3763
rect 3588 3757 3596 3763
rect 3636 3757 3740 3763
rect 3764 3757 3916 3763
rect 3924 3757 4300 3763
rect 4340 3757 4428 3763
rect 4468 3757 4716 3763
rect 4772 3757 4812 3763
rect 4916 3757 5116 3763
rect 5188 3757 5452 3763
rect 100 3737 332 3743
rect 452 3737 476 3743
rect 500 3737 508 3743
rect 525 3737 1084 3743
rect 13 3724 19 3736
rect 525 3723 531 3737
rect 1092 3737 1100 3743
rect 1277 3737 1292 3743
rect 1348 3737 1676 3743
rect 1684 3737 1852 3743
rect 1860 3737 2300 3743
rect 2308 3737 2316 3743
rect 2356 3737 2492 3743
rect 2916 3737 2924 3743
rect 2948 3737 3052 3743
rect 3060 3737 3852 3743
rect 3876 3737 3932 3743
rect 3956 3737 3980 3743
rect 3988 3737 4252 3743
rect 4308 3737 4316 3743
rect 4340 3737 4956 3743
rect 5172 3737 5180 3743
rect 5236 3737 5244 3743
rect 5197 3724 5203 3736
rect 5341 3724 5347 3736
rect 372 3717 531 3723
rect 548 3717 556 3723
rect 628 3717 636 3723
rect 708 3717 716 3723
rect 836 3717 892 3723
rect 900 3717 908 3723
rect 964 3717 1004 3723
rect 1156 3717 2108 3723
rect 2132 3717 2364 3723
rect 2436 3717 2492 3723
rect 2628 3717 2780 3723
rect 2788 3717 2796 3723
rect 2820 3717 3228 3723
rect 3236 3717 3564 3723
rect 3572 3717 4044 3723
rect 4148 3717 4748 3723
rect 4820 3717 4924 3723
rect 4948 3717 5164 3723
rect 68 3697 76 3703
rect 324 3697 396 3703
rect 516 3697 524 3703
rect 612 3697 652 3703
rect 868 3697 1148 3703
rect 1220 3697 1372 3703
rect 1380 3697 1388 3703
rect 1444 3697 1452 3703
rect 1476 3697 1484 3703
rect 1524 3697 1532 3703
rect 1828 3697 1836 3703
rect 1924 3697 2044 3703
rect 2052 3697 2188 3703
rect 2212 3697 2252 3703
rect 2260 3697 2284 3703
rect 2340 3697 2492 3703
rect 2500 3697 2540 3703
rect 2548 3697 2908 3703
rect 3012 3697 3020 3703
rect 3076 3697 3420 3703
rect 3524 3697 3596 3703
rect 3684 3697 3724 3703
rect 3812 3697 4012 3703
rect 4132 3697 4220 3703
rect 4276 3697 4300 3703
rect 4388 3697 4620 3703
rect 4644 3697 4684 3703
rect 4708 3697 4764 3703
rect 4804 3697 4844 3703
rect 4932 3697 5228 3703
rect 5316 3697 5388 3703
rect 5444 3697 5516 3703
rect 301 3684 307 3696
rect 813 3684 819 3696
rect 36 3677 284 3683
rect 836 3677 940 3683
rect 948 3677 1180 3683
rect 1252 3677 1260 3683
rect 1268 3677 1756 3683
rect 1764 3677 2092 3683
rect 2100 3677 2428 3683
rect 2468 3677 2524 3683
rect 4148 3677 4940 3683
rect 5028 3677 5068 3683
rect 3965 3664 3971 3676
rect 1652 3657 1756 3663
rect 1764 3657 1884 3663
rect 1892 3657 2124 3663
rect 4788 3657 5324 3663
rect 2692 3637 2700 3643
rect 3220 3637 3228 3643
rect 4372 3637 4524 3643
rect 4900 3637 5164 3643
rect 3133 3624 3139 3636
rect 717 3617 972 3623
rect 717 3603 723 3617
rect 4852 3617 5004 3623
rect 676 3597 723 3603
rect 1412 3597 1484 3603
rect 1972 3597 1996 3603
rect 2116 3597 2124 3603
rect 2660 3597 2764 3603
rect 3028 3597 3388 3603
rect 3556 3597 3708 3603
rect 3828 3597 4492 3603
rect 724 3577 748 3583
rect 2628 3577 3148 3583
rect 3156 3577 3196 3583
rect 3204 3577 3244 3583
rect 3348 3577 3660 3583
rect 3668 3577 4156 3583
rect 4164 3577 4236 3583
rect 1364 3557 1500 3563
rect 1508 3557 1548 3563
rect 2564 3557 2636 3563
rect 2644 3557 2956 3563
rect 2964 3557 2972 3563
rect 2980 3557 3036 3563
rect 4388 3557 4428 3563
rect 116 3537 460 3543
rect 468 3537 476 3543
rect 532 3537 604 3543
rect 772 3537 780 3543
rect 820 3537 1580 3543
rect 1684 3537 1692 3543
rect 1748 3537 1820 3543
rect 1972 3537 2076 3543
rect 2084 3537 2284 3543
rect 2948 3537 3084 3543
rect 3108 3537 3148 3543
rect 3220 3537 3228 3543
rect 3268 3537 3292 3543
rect 3396 3537 3468 3543
rect 3972 3537 4012 3543
rect 4244 3537 4380 3543
rect 4420 3537 4716 3543
rect 5076 3537 5436 3543
rect 308 3517 812 3523
rect 836 3517 844 3523
rect 1076 3517 1372 3523
rect 1380 3517 1388 3523
rect 1396 3517 2252 3523
rect 2276 3517 2300 3523
rect 2308 3517 2348 3523
rect 2356 3517 2460 3523
rect 2756 3517 2796 3523
rect 2820 3517 2844 3523
rect 3076 3517 3756 3523
rect 4029 3523 4035 3536
rect 4020 3517 4035 3523
rect 4052 3517 4060 3523
rect 4100 3517 4108 3523
rect 4132 3517 4252 3523
rect 4292 3517 4300 3523
rect 4532 3517 4732 3523
rect 4756 3517 4812 3523
rect 5060 3517 5084 3523
rect 5188 3517 5260 3523
rect 5332 3517 5388 3523
rect 5540 3517 5580 3523
rect 388 3497 396 3503
rect 468 3497 588 3503
rect 596 3497 908 3503
rect 996 3497 1132 3503
rect 1204 3497 1660 3503
rect 1684 3497 1788 3503
rect 1796 3497 1804 3503
rect 1876 3497 1980 3503
rect 2084 3497 2380 3503
rect 2836 3497 3212 3503
rect 3220 3497 3660 3503
rect 3668 3497 4028 3503
rect 4052 3497 4652 3503
rect 4660 3497 4956 3503
rect 5444 3497 5516 3503
rect 36 3477 76 3483
rect 180 3477 188 3483
rect 452 3477 1276 3483
rect 1284 3477 1340 3483
rect 1364 3477 1452 3483
rect 1492 3477 1580 3483
rect 1588 3477 2316 3483
rect 2836 3477 2892 3483
rect 3012 3477 3116 3483
rect 3140 3477 3212 3483
rect 3220 3477 3692 3483
rect 3732 3477 3820 3483
rect 3892 3477 4172 3483
rect 4180 3477 4716 3483
rect 4724 3477 4988 3483
rect 4996 3477 5148 3483
rect 5172 3477 5260 3483
rect 5268 3477 5324 3483
rect 260 3457 332 3463
rect 580 3457 956 3463
rect 1044 3457 1340 3463
rect 1348 3457 1516 3463
rect 1524 3457 1676 3463
rect 1684 3457 2124 3463
rect 2132 3457 2140 3463
rect 2180 3457 2268 3463
rect 2772 3457 2828 3463
rect 2932 3457 2940 3463
rect 2948 3457 2956 3463
rect 2980 3457 3020 3463
rect 3028 3457 3036 3463
rect 3204 3457 3212 3463
rect 3236 3457 3740 3463
rect 3748 3457 3836 3463
rect 3860 3457 3884 3463
rect 3924 3457 3996 3463
rect 4020 3457 4060 3463
rect 4100 3457 4172 3463
rect 4244 3457 4364 3463
rect 4404 3457 4844 3463
rect 4932 3457 4940 3463
rect 5028 3457 5100 3463
rect 5172 3457 5212 3463
rect 596 3437 764 3443
rect 884 3437 892 3443
rect 964 3437 972 3443
rect 1012 3437 1100 3443
rect 1476 3437 1548 3443
rect 1700 3437 1708 3443
rect 1924 3437 1932 3443
rect 2628 3437 2700 3443
rect 2932 3437 3404 3443
rect 3412 3437 4268 3443
rect 4292 3437 4316 3443
rect 4484 3437 5196 3443
rect 756 3417 1036 3423
rect 1092 3417 1132 3423
rect 1284 3417 1292 3423
rect 1668 3417 1724 3423
rect 1780 3417 1852 3423
rect 1860 3417 2028 3423
rect 2484 3417 2492 3423
rect 2884 3417 3100 3423
rect 3204 3417 3276 3423
rect 3300 3417 3340 3423
rect 3373 3417 3532 3423
rect 148 3397 172 3403
rect 980 3397 1004 3403
rect 1044 3397 1155 3403
rect 132 3377 140 3383
rect 324 3377 332 3383
rect 372 3377 380 3383
rect 500 3377 588 3383
rect 820 3377 908 3383
rect 1149 3383 1155 3397
rect 1220 3397 1292 3403
rect 1412 3397 1548 3403
rect 1604 3397 1612 3403
rect 1924 3397 1932 3403
rect 1988 3397 1996 3403
rect 2116 3397 2124 3403
rect 2244 3397 2252 3403
rect 2276 3397 2316 3403
rect 3373 3403 3379 3417
rect 3540 3417 3596 3423
rect 4061 3417 4236 3423
rect 2724 3397 3379 3403
rect 3620 3397 3900 3403
rect 4061 3403 4067 3417
rect 4244 3417 4652 3423
rect 4948 3417 4956 3423
rect 5092 3417 5340 3423
rect 3908 3397 4067 3403
rect 4084 3397 4108 3403
rect 4164 3397 4172 3403
rect 4356 3397 4364 3403
rect 4548 3397 4620 3403
rect 4676 3397 4684 3403
rect 4788 3397 4940 3403
rect 4996 3397 5020 3403
rect 5124 3397 5132 3403
rect 5316 3397 5388 3403
rect 4445 3384 4451 3396
rect 1149 3377 1292 3383
rect 1428 3377 1436 3383
rect 1444 3377 1484 3383
rect 1540 3377 1612 3383
rect 1652 3377 1932 3383
rect 2100 3377 2108 3383
rect 2164 3377 2252 3383
rect 2276 3377 2444 3383
rect 2628 3377 2636 3383
rect 2980 3377 3212 3383
rect 3348 3377 3388 3383
rect 3524 3377 3724 3383
rect 3860 3377 4428 3383
rect 4644 3377 4732 3383
rect 4749 3377 4764 3383
rect 4788 3377 5068 3383
rect 5124 3377 5132 3383
rect 5188 3377 5196 3383
rect 5252 3377 5388 3383
rect 5492 3377 5500 3383
rect 3469 3364 3475 3376
rect 132 3357 204 3363
rect 260 3357 396 3363
rect 452 3357 748 3363
rect 772 3357 780 3363
rect 900 3357 1308 3363
rect 1316 3357 1484 3363
rect 1572 3357 2556 3363
rect 2564 3357 2572 3363
rect 2612 3357 2924 3363
rect 2948 3357 3020 3363
rect 3092 3357 3100 3363
rect 3124 3357 3292 3363
rect 3396 3357 3420 3363
rect 3652 3357 3660 3363
rect 3700 3357 3708 3363
rect 3716 3357 4860 3363
rect 4868 3357 4908 3363
rect 4916 3357 5004 3363
rect 5124 3357 5132 3363
rect 5380 3357 5404 3363
rect 5197 3344 5203 3356
rect 324 3337 380 3343
rect 404 3337 524 3343
rect 580 3337 636 3343
rect 644 3337 652 3343
rect 836 3337 1564 3343
rect 1636 3337 1676 3343
rect 1748 3337 1804 3343
rect 1844 3337 2108 3343
rect 2324 3337 2540 3343
rect 2676 3337 2684 3343
rect 2724 3337 2748 3343
rect 2797 3337 2812 3343
rect 2820 3337 2844 3343
rect 2916 3337 2956 3343
rect 3012 3337 3100 3343
rect 3108 3337 3308 3343
rect 3364 3337 3500 3343
rect 3620 3337 3644 3343
rect 3764 3337 4076 3343
rect 4084 3337 4396 3343
rect 4436 3337 4444 3343
rect 4484 3337 4492 3343
rect 4612 3337 4636 3343
rect 4676 3337 4684 3343
rect 61 3324 67 3336
rect 2621 3324 2627 3336
rect 3581 3324 3587 3336
rect 4925 3324 4931 3343
rect 4964 3337 5084 3343
rect 5396 3337 5436 3343
rect 196 3317 220 3323
rect 292 3317 412 3323
rect 484 3317 812 3323
rect 948 3317 956 3323
rect 996 3317 1020 3323
rect 1044 3317 1052 3323
rect 1060 3317 1244 3323
rect 1268 3317 1356 3323
rect 1476 3317 1740 3323
rect 1764 3317 1884 3323
rect 2068 3317 2156 3323
rect 2308 3317 2604 3323
rect 2692 3317 2764 3323
rect 3044 3317 3228 3323
rect 3332 3317 3404 3323
rect 3412 3317 3420 3323
rect 3444 3317 3500 3323
rect 3812 3317 3852 3323
rect 3901 3317 4844 3323
rect 68 3297 300 3303
rect 308 3297 828 3303
rect 884 3297 892 3303
rect 916 3297 1516 3303
rect 1524 3297 1532 3303
rect 1700 3297 1724 3303
rect 2292 3297 2476 3303
rect 2580 3297 2668 3303
rect 3204 3297 3244 3303
rect 3901 3303 3907 3317
rect 4948 3317 5148 3323
rect 5204 3317 5228 3323
rect 5332 3317 5516 3323
rect 3268 3297 3907 3303
rect 3924 3297 4060 3303
rect 4084 3297 4092 3303
rect 4196 3297 4204 3303
rect 4484 3297 4588 3303
rect 4692 3297 4796 3303
rect 4804 3297 4892 3303
rect 4964 3297 4988 3303
rect 4996 3297 5052 3303
rect 5204 3297 5276 3303
rect 5405 3297 5532 3303
rect 308 3277 604 3283
rect 820 3277 1196 3283
rect 1268 3277 1452 3283
rect 1460 3277 1884 3283
rect 2852 3277 2876 3283
rect 3444 3277 4268 3283
rect 4500 3277 4508 3283
rect 5405 3283 5411 3297
rect 4868 3277 5411 3283
rect 5428 3277 5484 3283
rect 404 3257 412 3263
rect 580 3257 604 3263
rect 948 3257 1004 3263
rect 1245 3257 1340 3263
rect 1245 3243 1251 3257
rect 2852 3257 2860 3263
rect 4420 3257 4732 3263
rect 4740 3257 4780 3263
rect 1204 3237 1251 3243
rect 1924 3237 1948 3243
rect 3652 3237 4444 3243
rect 4980 3237 5116 3243
rect 5124 3237 5196 3243
rect 5348 3237 5564 3243
rect 1085 3224 1091 3236
rect 1588 3217 1596 3223
rect 2340 3217 2364 3223
rect 3796 3217 3804 3223
rect 4564 3217 4572 3223
rect 5188 3217 5356 3223
rect 1092 3197 1100 3203
rect 1540 3197 1548 3203
rect 1716 3197 1724 3203
rect 1940 3197 1980 3203
rect 2004 3197 2012 3203
rect 3076 3197 3084 3203
rect 3572 3197 3676 3203
rect 3684 3197 4044 3203
rect 708 3177 828 3183
rect 1732 3177 1740 3183
rect 1764 3177 1788 3183
rect 2372 3177 2428 3183
rect 3460 3177 3468 3183
rect 3748 3177 3756 3183
rect 3812 3177 3948 3183
rect 4132 3177 4284 3183
rect 644 3157 652 3163
rect 836 3157 940 3163
rect 948 3157 1868 3163
rect 1876 3157 1916 3163
rect 1997 3163 2003 3176
rect 1988 3157 2003 3163
rect 2900 3157 2908 3163
rect 2948 3157 3612 3163
rect 3652 3157 4268 3163
rect 4292 3157 4316 3163
rect 4372 3157 4380 3163
rect 5108 3157 5212 3163
rect 5220 3157 5308 3163
rect 5476 3157 5564 3163
rect 404 3137 476 3143
rect 628 3137 668 3143
rect 676 3137 940 3143
rect 964 3137 1020 3143
rect 1220 3137 1228 3143
rect 1364 3137 1372 3143
rect 1492 3137 1836 3143
rect 2132 3137 2188 3143
rect 2820 3137 2892 3143
rect 2980 3137 3468 3143
rect 3476 3137 3532 3143
rect 3796 3137 3804 3143
rect 3860 3137 4044 3143
rect 4068 3137 4892 3143
rect 4973 3124 4979 3136
rect 5053 3124 5059 3136
rect 180 3117 332 3123
rect 388 3117 524 3123
rect 548 3117 588 3123
rect 644 3117 716 3123
rect 804 3117 812 3123
rect 868 3117 908 3123
rect 996 3117 1452 3123
rect 1460 3117 1516 3123
rect 1572 3117 1580 3123
rect 1652 3117 1660 3123
rect 2116 3117 2156 3123
rect 2164 3117 2444 3123
rect 2468 3117 2476 3123
rect 2676 3117 3100 3123
rect 3316 3117 3324 3123
rect 3348 3117 3356 3123
rect 3460 3117 3548 3123
rect 3556 3117 3923 3123
rect 3261 3104 3267 3116
rect 244 3097 364 3103
rect 404 3097 460 3103
rect 516 3097 1036 3103
rect 1101 3097 1116 3103
rect 1204 3097 1212 3103
rect 1220 3097 1388 3103
rect 1460 3097 1468 3103
rect 1540 3097 1660 3103
rect 1668 3097 1788 3103
rect 1860 3097 2076 3103
rect 2196 3097 2236 3103
rect 2388 3097 2556 3103
rect 2628 3097 2700 3103
rect 2820 3097 3036 3103
rect 3076 3097 3116 3103
rect 3300 3097 3420 3103
rect 3556 3097 3676 3103
rect 3684 3097 3900 3103
rect 3917 3103 3923 3117
rect 4084 3117 4108 3123
rect 4180 3117 4332 3123
rect 4340 3117 4348 3123
rect 4372 3117 4396 3123
rect 4420 3117 4604 3123
rect 4660 3117 4668 3123
rect 4701 3117 4716 3123
rect 4820 3117 4924 3123
rect 4996 3117 5020 3123
rect 5028 3117 5043 3123
rect 3917 3097 4172 3103
rect 4260 3097 4332 3103
rect 4356 3097 4476 3103
rect 4548 3097 4684 3103
rect 4692 3097 4748 3103
rect 4788 3097 4844 3103
rect 4861 3097 4876 3103
rect 125 3084 131 3096
rect 68 3077 92 3083
rect 260 3077 316 3083
rect 324 3077 332 3083
rect 365 3083 371 3096
rect 4861 3084 4867 3097
rect 4932 3097 5020 3103
rect 5037 3103 5043 3117
rect 5396 3117 5411 3123
rect 5540 3117 5580 3123
rect 5629 3117 5660 3123
rect 5037 3097 5116 3103
rect 5140 3097 5196 3103
rect 5252 3097 5260 3103
rect 365 3077 508 3083
rect 516 3077 972 3083
rect 980 3077 1596 3083
rect 1604 3077 1612 3083
rect 1636 3077 1820 3083
rect 1844 3077 1852 3083
rect 1860 3077 1932 3083
rect 1972 3077 2380 3083
rect 2404 3077 2780 3083
rect 2788 3077 3900 3083
rect 4157 3077 4636 3083
rect 180 3057 188 3063
rect 260 3057 268 3063
rect 324 3057 348 3063
rect 356 3057 428 3063
rect 452 3057 460 3063
rect 468 3057 940 3063
rect 948 3057 1052 3063
rect 1140 3057 1148 3063
rect 1172 3057 1276 3063
rect 1300 3057 1308 3063
rect 1316 3057 1852 3063
rect 1892 3057 1964 3063
rect 2084 3057 2220 3063
rect 2516 3057 2604 3063
rect 2692 3057 2748 3063
rect 2772 3057 2972 3063
rect 3284 3057 3308 3063
rect 3380 3057 3388 3063
rect 3412 3057 3692 3063
rect 3716 3057 3724 3063
rect 4157 3063 4163 3077
rect 4836 3077 4844 3083
rect 4916 3077 5100 3083
rect 5108 3077 5276 3083
rect 5508 3077 5516 3083
rect 3796 3057 4163 3063
rect 4324 3057 4348 3063
rect 4372 3057 4412 3063
rect 4532 3057 4668 3063
rect 4692 3057 4796 3063
rect 4884 3057 5004 3063
rect 5012 3057 5148 3063
rect 5156 3057 5164 3063
rect 5268 3057 5276 3063
rect 2061 3044 2067 3056
rect 4429 3044 4435 3056
rect 324 3037 332 3043
rect 340 3037 348 3043
rect 900 3037 1212 3043
rect 1348 3037 1564 3043
rect 1588 3037 1628 3043
rect 1988 3037 2012 3043
rect 2196 3037 2316 3043
rect 2740 3037 3324 3043
rect 3332 3037 3356 3043
rect 3524 3037 3692 3043
rect 3860 3037 3916 3043
rect 4068 3037 4092 3043
rect 4628 3037 4940 3043
rect 5060 3037 5068 3043
rect 5092 3037 5132 3043
rect 573 3024 579 3036
rect 1172 3017 1548 3023
rect 1556 3017 1587 3023
rect 1044 2997 1068 3003
rect 1076 2997 1084 3003
rect 1492 2997 1548 3003
rect 1581 3003 1587 3017
rect 1604 3017 1644 3023
rect 2644 3017 2828 3023
rect 2868 3017 2988 3023
rect 2996 3017 3356 3023
rect 3844 3017 3852 3023
rect 3956 3017 4284 3023
rect 4292 3017 4492 3023
rect 4644 3017 4876 3023
rect 5124 3017 5324 3023
rect 5357 3017 5516 3023
rect 1581 2997 1772 3003
rect 1956 2997 2044 3003
rect 2052 2997 2172 3003
rect 2180 2997 2252 3003
rect 2372 2997 2428 3003
rect 3092 2997 3180 3003
rect 3252 2997 3260 3003
rect 3604 2997 3612 3003
rect 3716 2997 3836 3003
rect 3844 2997 3884 3003
rect 4196 2997 4412 3003
rect 4420 2997 4860 3003
rect 4980 2997 5020 3003
rect 5236 2997 5244 3003
rect 5357 3003 5363 3017
rect 5316 2997 5363 3003
rect 5572 2997 5660 3003
rect 116 2977 124 2983
rect 196 2977 284 2983
rect 596 2977 652 2983
rect 740 2977 780 2983
rect 820 2977 828 2983
rect 1028 2977 1116 2983
rect 1268 2977 1308 2983
rect 1508 2977 1516 2983
rect 1620 2977 1644 2983
rect 1732 2977 1852 2983
rect 1869 2977 1875 2996
rect 2068 2977 2108 2983
rect 2180 2977 2236 2983
rect 2308 2977 2323 2983
rect 20 2957 28 2963
rect 148 2957 236 2963
rect 244 2957 588 2963
rect 612 2957 764 2963
rect 772 2957 1036 2963
rect 1044 2957 1244 2963
rect 1284 2957 1292 2963
rect 1316 2957 1436 2963
rect 1604 2957 1932 2963
rect 1940 2957 2300 2963
rect 2317 2963 2323 2977
rect 2340 2977 2428 2983
rect 2692 2977 2732 2983
rect 2772 2977 2812 2983
rect 3156 2977 3404 2983
rect 3460 2977 3468 2983
rect 3492 2977 3500 2983
rect 3572 2977 3580 2983
rect 4260 2977 4556 2983
rect 4804 2977 4828 2983
rect 5188 2977 5324 2983
rect 5380 2977 5420 2983
rect 5524 2977 5635 2983
rect 4989 2964 4995 2976
rect 2317 2957 2348 2963
rect 2404 2957 2444 2963
rect 2877 2957 2892 2963
rect 3012 2957 3020 2963
rect 3092 2957 3548 2963
rect 3556 2957 3564 2963
rect 3716 2957 3724 2963
rect 3732 2957 3772 2963
rect 4084 2957 4108 2963
rect 4308 2957 4316 2963
rect 4340 2957 4492 2963
rect 4740 2957 4876 2963
rect 4884 2957 4908 2963
rect 4932 2957 4940 2963
rect 5012 2957 5020 2963
rect 5172 2957 5260 2963
rect 5348 2957 5452 2963
rect 68 2937 156 2943
rect 276 2937 284 2943
rect 420 2937 460 2943
rect 484 2937 524 2943
rect 532 2937 540 2943
rect 596 2937 748 2943
rect 836 2937 924 2943
rect 964 2937 972 2943
rect 1124 2937 1164 2943
rect 1204 2937 1212 2943
rect 1252 2937 1356 2943
rect 1636 2937 1676 2943
rect 1796 2937 1804 2943
rect 1844 2937 2076 2943
rect 2132 2937 2204 2943
rect 2212 2937 2236 2943
rect 2276 2937 2284 2943
rect 2356 2937 2380 2943
rect 2692 2937 2732 2943
rect 2740 2937 3884 2943
rect 4052 2937 4156 2943
rect 4276 2937 4540 2943
rect 4612 2937 4636 2943
rect 4676 2937 4780 2943
rect 4852 2937 5004 2943
rect 5060 2937 5068 2943
rect 5076 2937 5244 2943
rect 5396 2937 5500 2943
rect 4029 2924 4035 2936
rect 164 2917 540 2923
rect 660 2917 956 2923
rect 1012 2917 1020 2923
rect 1028 2917 1308 2923
rect 1348 2917 1708 2923
rect 1812 2917 2636 2923
rect 2724 2917 2924 2923
rect 2932 2917 2988 2923
rect 2996 2917 3004 2923
rect 3140 2917 3148 2923
rect 3172 2917 3436 2923
rect 3444 2917 3484 2923
rect 3508 2917 3596 2923
rect 3652 2917 3683 2923
rect 36 2897 76 2903
rect 260 2897 275 2903
rect 292 2897 348 2903
rect 356 2897 444 2903
rect 548 2897 1020 2903
rect 1092 2897 1292 2903
rect 1300 2897 1372 2903
rect 1924 2897 1932 2903
rect 2116 2897 2275 2903
rect 20 2877 332 2883
rect 372 2877 380 2883
rect 516 2877 620 2883
rect 964 2877 1052 2883
rect 1908 2877 1980 2883
rect 2164 2877 2252 2883
rect 2269 2883 2275 2897
rect 2308 2897 2396 2903
rect 2820 2897 2892 2903
rect 3028 2897 3116 2903
rect 3188 2897 3212 2903
rect 3236 2897 3244 2903
rect 3316 2897 3340 2903
rect 3396 2897 3436 2903
rect 3460 2897 3468 2903
rect 3492 2897 3532 2903
rect 3540 2897 3548 2903
rect 3620 2897 3660 2903
rect 3677 2903 3683 2917
rect 3732 2917 3740 2923
rect 3860 2917 3884 2923
rect 3940 2917 3964 2923
rect 4068 2917 4204 2923
rect 4228 2917 4300 2923
rect 4340 2917 4348 2923
rect 4420 2917 4444 2923
rect 4484 2917 4508 2923
rect 4532 2917 4652 2923
rect 4740 2917 4748 2923
rect 4788 2917 4828 2923
rect 4868 2917 4876 2923
rect 4900 2917 4956 2923
rect 5060 2917 5068 2923
rect 5252 2917 5452 2923
rect 3677 2897 3820 2903
rect 3972 2897 4060 2903
rect 4260 2897 4268 2903
rect 4276 2897 4716 2903
rect 4724 2897 5116 2903
rect 5405 2884 5411 2896
rect 2269 2877 2460 2883
rect 2708 2877 2796 2883
rect 3060 2877 3196 2883
rect 3204 2877 3372 2883
rect 3380 2877 3916 2883
rect 4404 2877 4524 2883
rect 4788 2877 4844 2883
rect 4852 2877 4860 2883
rect 4932 2877 5148 2883
rect 1149 2864 1155 2876
rect 1284 2857 2156 2863
rect 3316 2857 3340 2863
rect 3780 2857 4412 2863
rect 4420 2857 4428 2863
rect 3405 2844 3411 2856
rect 3741 2844 3747 2856
rect 340 2837 1164 2843
rect 2292 2837 2316 2843
rect 3796 2837 3996 2843
rect 4004 2837 5196 2843
rect 2964 2817 3004 2823
rect 3332 2817 3340 2823
rect 3412 2817 3420 2823
rect 3668 2817 3692 2823
rect 3860 2817 3884 2823
rect 5220 2817 5244 2823
rect 772 2797 780 2803
rect 852 2797 860 2803
rect 1204 2797 1212 2803
rect 1572 2797 1628 2803
rect 1636 2797 1740 2803
rect 2388 2797 2444 2803
rect 2612 2797 2620 2803
rect 2852 2797 3324 2803
rect 308 2777 540 2783
rect 548 2777 1500 2783
rect 1556 2777 2044 2783
rect 3524 2777 4012 2783
rect 5268 2777 5372 2783
rect 644 2757 652 2763
rect 804 2757 844 2763
rect 1204 2757 1260 2763
rect 1508 2757 1612 2763
rect 1636 2757 1660 2763
rect 1812 2757 1836 2763
rect 1844 2757 1852 2763
rect 1908 2757 1916 2763
rect 2116 2757 2140 2763
rect 2660 2757 2668 2763
rect 2948 2757 3132 2763
rect 3460 2757 3468 2763
rect 3821 2757 3916 2763
rect 500 2737 844 2743
rect 932 2737 956 2743
rect 1028 2737 1772 2743
rect 1780 2737 1788 2743
rect 1828 2737 2332 2743
rect 2580 2737 2652 2743
rect 2836 2737 2924 2743
rect 3028 2737 3100 2743
rect 3821 2743 3827 2757
rect 4100 2757 4156 2763
rect 4196 2757 4204 2763
rect 4228 2757 4252 2763
rect 4324 2757 4428 2763
rect 3156 2737 3827 2743
rect 3844 2737 4060 2743
rect 4132 2737 4204 2743
rect 4244 2737 4284 2743
rect 4324 2737 4588 2743
rect 4676 2737 4684 2743
rect 4820 2737 5340 2743
rect 5412 2737 5484 2743
rect 116 2717 156 2723
rect 164 2717 268 2723
rect 276 2717 364 2723
rect 580 2717 636 2723
rect 660 2717 1004 2723
rect 1028 2717 1436 2723
rect 1444 2717 1452 2723
rect 1556 2717 1788 2723
rect 1796 2717 2204 2723
rect 2244 2717 2252 2723
rect 2436 2717 2444 2723
rect 2468 2717 2483 2723
rect 2852 2717 2892 2723
rect 2948 2717 3004 2723
rect 3012 2717 3100 2723
rect 3236 2717 3276 2723
rect 3348 2717 3420 2723
rect 3556 2717 3596 2723
rect 3780 2717 3788 2723
rect 3812 2717 4252 2723
rect 4532 2717 4796 2723
rect 4820 2717 4828 2723
rect 4884 2717 4908 2723
rect 4932 2717 4972 2723
rect 5028 2717 5036 2723
rect 5460 2717 5516 2723
rect 340 2697 412 2703
rect 452 2697 556 2703
rect 612 2697 780 2703
rect 916 2697 924 2703
rect 948 2697 1084 2703
rect 1108 2697 1116 2703
rect 1188 2697 1260 2703
rect 1380 2697 1404 2703
rect 1460 2697 1820 2703
rect 1924 2697 1932 2703
rect 2020 2697 2028 2703
rect 2052 2697 2092 2703
rect 2100 2697 2492 2703
rect 3012 2697 3084 2703
rect 3172 2697 3196 2703
rect 3204 2697 3516 2703
rect 3716 2697 3740 2703
rect 3764 2697 3804 2703
rect 3844 2697 3868 2703
rect 3892 2697 3916 2703
rect 3972 2697 4060 2703
rect 4100 2697 4300 2703
rect 4388 2697 4396 2703
rect 4500 2697 4556 2703
rect 4580 2697 4620 2703
rect 4660 2697 4924 2703
rect 4948 2697 5100 2703
rect 5252 2697 5324 2703
rect 5380 2697 5452 2703
rect 5476 2697 5484 2703
rect 573 2684 579 2696
rect 589 2684 595 2696
rect 1325 2684 1331 2696
rect 5517 2684 5523 2696
rect 36 2677 92 2683
rect 148 2677 156 2683
rect 292 2677 316 2683
rect 676 2677 684 2683
rect 724 2677 732 2683
rect 788 2677 1004 2683
rect 1140 2677 1228 2683
rect 1348 2677 1468 2683
rect 1476 2677 1484 2683
rect 1524 2677 1532 2683
rect 1556 2677 1564 2683
rect 1700 2677 1756 2683
rect 1796 2677 1980 2683
rect 2180 2677 2195 2683
rect 2189 2664 2195 2677
rect 2244 2677 2316 2683
rect 2372 2677 2380 2683
rect 2452 2677 2508 2683
rect 2564 2677 2572 2683
rect 2628 2677 2636 2683
rect 2644 2677 2652 2683
rect 2772 2677 3004 2683
rect 3012 2677 3212 2683
rect 3300 2677 3315 2683
rect 3332 2677 3420 2683
rect 3428 2677 3500 2683
rect 3524 2677 3628 2683
rect 3636 2677 3740 2683
rect 3764 2677 3788 2683
rect 3796 2677 4220 2683
rect 4237 2677 4252 2683
rect 4237 2664 4243 2677
rect 4356 2677 4412 2683
rect 4452 2677 4748 2683
rect 4756 2677 4764 2683
rect 4868 2677 5116 2683
rect 5140 2677 5148 2683
rect 5380 2677 5395 2683
rect 260 2657 508 2663
rect 532 2657 780 2663
rect 804 2657 844 2663
rect 868 2657 1068 2663
rect 1092 2657 1244 2663
rect 1268 2657 1660 2663
rect 1668 2657 1932 2663
rect 1956 2657 1964 2663
rect 2004 2657 2124 2663
rect 2212 2657 2732 2663
rect 2804 2657 3612 2663
rect 3652 2657 3660 2663
rect 3716 2657 3731 2663
rect 3748 2657 3884 2663
rect 3892 2657 4044 2663
rect 4196 2657 4204 2663
rect 4484 2657 4668 2663
rect 4692 2657 4700 2663
rect 4756 2657 4764 2663
rect 4932 2657 4940 2663
rect 5268 2657 5292 2663
rect 260 2637 268 2643
rect 404 2637 460 2643
rect 548 2637 892 2643
rect 932 2637 940 2643
rect 996 2637 1004 2643
rect 1012 2637 1020 2643
rect 1060 2637 1148 2643
rect 1188 2637 1228 2643
rect 1268 2637 1276 2643
rect 1300 2637 1324 2643
rect 1364 2637 1436 2643
rect 1476 2637 1676 2643
rect 1972 2637 1980 2643
rect 2132 2637 2140 2643
rect 3300 2637 3404 2643
rect 3524 2637 3580 2643
rect 3588 2637 4124 2643
rect 4532 2637 4540 2643
rect 4692 2637 5132 2643
rect 5165 2637 5276 2643
rect 564 2617 1468 2623
rect 3140 2617 3356 2623
rect 3364 2617 3532 2623
rect 3588 2617 3596 2623
rect 3764 2617 3772 2623
rect 3796 2617 3804 2623
rect 3988 2617 4508 2623
rect 4868 2617 4876 2623
rect 5060 2617 5068 2623
rect 5165 2623 5171 2637
rect 5124 2617 5171 2623
rect 5572 2617 5635 2623
rect 116 2597 204 2603
rect 548 2597 908 2603
rect 1060 2597 1404 2603
rect 1412 2597 1500 2603
rect 1796 2597 1852 2603
rect 1876 2597 1916 2603
rect 2292 2597 2316 2603
rect 2516 2597 2556 2603
rect 2948 2597 2988 2603
rect 3604 2597 3980 2603
rect 4356 2597 4492 2603
rect 4612 2597 4620 2603
rect 5060 2597 5084 2603
rect 5188 2597 5212 2603
rect 5284 2597 5308 2603
rect 5444 2597 5532 2603
rect 3581 2584 3587 2596
rect 116 2577 124 2583
rect 324 2577 540 2583
rect 548 2577 572 2583
rect 836 2577 867 2583
rect 68 2557 76 2563
rect 324 2557 348 2563
rect 388 2557 396 2563
rect 452 2557 460 2563
rect 644 2557 668 2563
rect 708 2557 748 2563
rect 772 2557 780 2563
rect 861 2563 867 2577
rect 884 2577 892 2583
rect 900 2577 1036 2583
rect 1076 2577 1164 2583
rect 1220 2577 1356 2583
rect 1380 2577 1596 2583
rect 1604 2577 2012 2583
rect 2036 2577 2044 2583
rect 2260 2577 2268 2583
rect 2308 2577 2492 2583
rect 3012 2577 3100 2583
rect 3236 2577 3324 2583
rect 3716 2577 3788 2583
rect 3924 2577 3932 2583
rect 4084 2577 4236 2583
rect 4372 2577 4380 2583
rect 4452 2577 4460 2583
rect 4628 2577 4668 2583
rect 4868 2577 4988 2583
rect 5012 2577 5292 2583
rect 5300 2577 5324 2583
rect 5508 2577 5635 2583
rect 861 2557 988 2563
rect 1236 2557 1244 2563
rect 1268 2557 1308 2563
rect 1348 2557 1388 2563
rect 1412 2557 1420 2563
rect 1428 2557 1852 2563
rect 1860 2557 2108 2563
rect 2116 2557 2332 2563
rect 2340 2557 2476 2563
rect 2484 2557 2508 2563
rect 2692 2557 2716 2563
rect 2900 2557 2908 2563
rect 2980 2557 2988 2563
rect 3028 2557 3036 2563
rect 3092 2557 3388 2563
rect 3396 2557 4044 2563
rect 4052 2557 4428 2563
rect 4436 2557 5148 2563
rect 5156 2557 5228 2563
rect 5268 2557 5308 2563
rect 180 2537 252 2543
rect 468 2537 508 2543
rect 516 2537 652 2543
rect 676 2537 764 2543
rect 900 2537 972 2543
rect 1028 2537 1068 2543
rect 1092 2537 1244 2543
rect 1252 2537 1324 2543
rect 1396 2537 1404 2543
rect 1428 2537 1452 2543
rect 1476 2537 1516 2543
rect 1540 2537 1628 2543
rect 1812 2537 1900 2543
rect 2068 2537 2076 2543
rect 2244 2537 2300 2543
rect 2324 2537 2364 2543
rect 2372 2537 2396 2543
rect 2413 2524 2419 2543
rect 2436 2537 2444 2543
rect 2452 2537 3068 2543
rect 3108 2537 3148 2543
rect 3156 2537 3244 2543
rect 3268 2537 3292 2543
rect 3492 2537 3500 2543
rect 3572 2537 3644 2543
rect 3716 2537 3740 2543
rect 3780 2537 3788 2543
rect 3860 2537 3884 2543
rect 3924 2537 4140 2543
rect 4180 2537 4188 2543
rect 4228 2537 4236 2543
rect 4644 2537 4652 2543
rect 4676 2537 4684 2543
rect 4756 2537 4796 2543
rect 4925 2524 4931 2543
rect 4980 2537 5004 2543
rect 5044 2537 5132 2543
rect 5172 2537 5196 2543
rect 5380 2537 5388 2543
rect 5460 2537 5500 2543
rect 5524 2537 5580 2543
rect 4941 2524 4947 2536
rect 52 2517 332 2523
rect 484 2517 716 2523
rect 884 2517 908 2523
rect 964 2517 972 2523
rect 980 2517 1084 2523
rect 1092 2517 1772 2523
rect 1908 2517 2076 2523
rect 2436 2517 2444 2523
rect 2461 2517 2572 2523
rect 404 2497 588 2503
rect 932 2497 940 2503
rect 948 2497 1164 2503
rect 1396 2497 1420 2503
rect 1508 2497 1676 2503
rect 2461 2503 2467 2517
rect 2724 2517 3228 2523
rect 3236 2517 3580 2523
rect 3620 2517 4060 2523
rect 4180 2517 4364 2523
rect 4468 2517 4620 2523
rect 4628 2517 4636 2523
rect 4740 2517 4844 2523
rect 5012 2517 5020 2523
rect 5044 2517 5068 2523
rect 5236 2517 5340 2523
rect 5501 2504 5507 2516
rect 2260 2497 2467 2503
rect 2532 2497 2620 2503
rect 2788 2497 2956 2503
rect 3140 2497 3260 2503
rect 3284 2497 3340 2503
rect 3412 2497 3436 2503
rect 3556 2497 3564 2503
rect 3604 2497 3628 2503
rect 3668 2497 3804 2503
rect 4036 2497 4044 2503
rect 4100 2497 4140 2503
rect 4292 2497 4380 2503
rect 4564 2497 4572 2503
rect 4596 2497 4604 2503
rect 4676 2497 4716 2503
rect 4772 2497 4780 2503
rect 4820 2497 4828 2503
rect 4916 2497 4931 2503
rect 4948 2497 4956 2503
rect 5156 2497 5292 2503
rect 5300 2497 5372 2503
rect 1485 2484 1491 2496
rect 3981 2484 3987 2496
rect 452 2477 1148 2483
rect 3044 2477 3404 2483
rect 3412 2477 3628 2483
rect 3684 2477 3724 2483
rect 3748 2477 3804 2483
rect 4420 2477 4508 2483
rect 4516 2477 4956 2483
rect 5220 2477 5244 2483
rect 5268 2477 5388 2483
rect 3076 2457 3180 2463
rect 3220 2457 3228 2463
rect 3348 2457 3388 2463
rect 4004 2457 5532 2463
rect 1124 2437 1164 2443
rect 1172 2437 1596 2443
rect 1716 2437 1868 2443
rect 2036 2437 2268 2443
rect 2276 2437 2316 2443
rect 3140 2437 3148 2443
rect 4900 2437 4908 2443
rect 5252 2437 5276 2443
rect 1380 2417 1420 2423
rect 5252 2417 5356 2423
rect 420 2397 716 2403
rect 900 2397 1100 2403
rect 1108 2397 1356 2403
rect 2116 2397 2124 2403
rect 3892 2397 4236 2403
rect 5124 2397 5180 2403
rect 5476 2397 5500 2403
rect 3213 2384 3219 2396
rect 644 2377 716 2383
rect 1716 2377 1916 2383
rect 1972 2377 1996 2383
rect 3652 2377 3724 2383
rect 4196 2377 4268 2383
rect 4852 2377 4892 2383
rect 5028 2377 5036 2383
rect 2125 2364 2131 2376
rect 372 2357 540 2363
rect 628 2357 908 2363
rect 1668 2357 1676 2363
rect 1764 2357 1772 2363
rect 1924 2357 2076 2363
rect 3204 2357 3212 2363
rect 3524 2357 3900 2363
rect 4340 2357 4348 2363
rect 4532 2357 5132 2363
rect 5140 2357 5260 2363
rect 164 2337 284 2343
rect 292 2337 556 2343
rect 564 2337 764 2343
rect 804 2337 988 2343
rect 1172 2337 1884 2343
rect 1908 2337 1932 2343
rect 1988 2337 1996 2343
rect 2036 2337 2188 2343
rect 2692 2337 2844 2343
rect 2884 2337 2892 2343
rect 3380 2337 3500 2343
rect 3620 2337 3660 2343
rect 3940 2337 3964 2343
rect 4004 2337 4076 2343
rect 4100 2337 4332 2343
rect 4356 2337 4780 2343
rect 4868 2337 4876 2343
rect 4884 2337 5020 2343
rect 5156 2337 5212 2343
rect 356 2317 588 2323
rect 692 2317 700 2323
rect 740 2317 748 2323
rect 820 2317 892 2323
rect 932 2317 1299 2323
rect 388 2297 492 2303
rect 516 2297 572 2303
rect 708 2297 956 2303
rect 980 2297 1036 2303
rect 1140 2297 1276 2303
rect 1293 2303 1299 2317
rect 1316 2317 1484 2323
rect 1492 2317 1500 2323
rect 1508 2317 2092 2323
rect 2100 2317 2668 2323
rect 2676 2317 2780 2323
rect 2980 2317 3020 2323
rect 3092 2317 3180 2323
rect 3188 2317 3564 2323
rect 4420 2317 4556 2323
rect 4580 2317 4604 2323
rect 4644 2317 4956 2323
rect 5108 2317 5132 2323
rect 5140 2317 5196 2323
rect 5220 2317 5324 2323
rect 5460 2317 5468 2323
rect 5508 2317 5523 2323
rect 1293 2297 1804 2303
rect 1812 2297 1836 2303
rect 1860 2297 2588 2303
rect 2708 2297 2716 2303
rect 2964 2297 3084 2303
rect 3268 2297 3388 2303
rect 3460 2297 3500 2303
rect 3524 2297 3532 2303
rect 3604 2297 3612 2303
rect 3716 2297 3724 2303
rect 3732 2297 3868 2303
rect 3924 2297 3980 2303
rect 4020 2297 4220 2303
rect 4260 2297 4275 2303
rect 2637 2284 2643 2296
rect 3197 2284 3203 2296
rect 4269 2284 4275 2297
rect 4324 2297 4476 2303
rect 4532 2297 4748 2303
rect 4756 2297 5356 2303
rect 5364 2297 5548 2303
rect 4285 2284 4291 2296
rect 148 2277 156 2283
rect 164 2277 204 2283
rect 212 2277 924 2283
rect 964 2277 1404 2283
rect 1428 2277 1436 2283
rect 1556 2277 1644 2283
rect 1668 2277 1724 2283
rect 1796 2277 1804 2283
rect 1876 2277 2028 2283
rect 2052 2277 2060 2283
rect 2068 2277 2572 2283
rect 2708 2277 2780 2283
rect 2916 2277 2924 2283
rect 3060 2277 3068 2283
rect 3284 2277 3340 2283
rect 3380 2277 3532 2283
rect 3565 2277 3596 2283
rect 3117 2264 3123 2276
rect 420 2257 460 2263
rect 788 2257 988 2263
rect 996 2257 1004 2263
rect 1044 2257 1196 2263
rect 1204 2257 1260 2263
rect 1348 2257 1420 2263
rect 1428 2257 1948 2263
rect 1956 2257 2140 2263
rect 2148 2257 2188 2263
rect 2228 2257 2764 2263
rect 2820 2257 2940 2263
rect 2980 2257 2988 2263
rect 2996 2257 3068 2263
rect 3124 2257 3276 2263
rect 3332 2257 3404 2263
rect 3565 2263 3571 2277
rect 3796 2277 3804 2283
rect 3892 2277 4140 2283
rect 4180 2277 4204 2283
rect 4308 2277 4444 2283
rect 4468 2277 4556 2283
rect 4580 2277 4588 2283
rect 4644 2277 5084 2283
rect 5092 2277 5100 2283
rect 5268 2277 5564 2283
rect 3476 2257 3571 2263
rect 3588 2257 3708 2263
rect 3748 2257 3836 2263
rect 3860 2257 3996 2263
rect 4020 2257 4044 2263
rect 4148 2257 4460 2263
rect 4468 2257 4908 2263
rect 4932 2257 4940 2263
rect 4948 2257 5068 2263
rect 5076 2257 5180 2263
rect 5236 2257 5388 2263
rect 820 2237 828 2243
rect 916 2237 972 2243
rect 1236 2237 1356 2243
rect 1428 2237 1452 2243
rect 1476 2237 1548 2243
rect 1668 2237 1676 2243
rect 1732 2237 1740 2243
rect 1860 2237 1932 2243
rect 1988 2237 2003 2243
rect 1165 2224 1171 2236
rect 1997 2224 2003 2237
rect 2020 2237 2028 2243
rect 2052 2237 2060 2243
rect 2180 2237 2268 2243
rect 2308 2237 2348 2243
rect 2516 2237 2524 2243
rect 2676 2237 3260 2243
rect 3268 2237 3868 2243
rect 3876 2237 3884 2243
rect 3924 2237 3996 2243
rect 4036 2237 4156 2243
rect 4340 2237 4348 2243
rect 4484 2237 4796 2243
rect 4900 2237 5020 2243
rect 5028 2237 5308 2243
rect 5316 2237 5372 2243
rect 5380 2237 5484 2243
rect 628 2217 636 2223
rect 644 2217 844 2223
rect 1284 2217 1436 2223
rect 1604 2217 1708 2223
rect 2500 2217 2556 2223
rect 3572 2217 3580 2223
rect 3668 2217 3676 2223
rect 4052 2217 4076 2223
rect 4164 2217 4300 2223
rect 4804 2217 4812 2223
rect 3309 2204 3315 2216
rect 612 2197 636 2203
rect 1076 2197 1100 2203
rect 1124 2197 1260 2203
rect 1300 2197 1308 2203
rect 1412 2197 1532 2203
rect 1572 2197 1580 2203
rect 1668 2197 1692 2203
rect 1972 2197 2003 2203
rect 196 2177 316 2183
rect 516 2177 572 2183
rect 628 2177 652 2183
rect 740 2177 844 2183
rect 900 2177 956 2183
rect 980 2177 988 2183
rect 1028 2177 1036 2183
rect 1220 2177 1276 2183
rect 1300 2177 1692 2183
rect 1700 2177 1724 2183
rect 1844 2177 1980 2183
rect 1997 2183 2003 2197
rect 2372 2197 2524 2203
rect 2532 2197 2540 2203
rect 2724 2197 2748 2203
rect 3268 2197 3292 2203
rect 3428 2197 3452 2203
rect 3780 2197 3804 2203
rect 4116 2197 4140 2203
rect 4228 2197 4236 2203
rect 4308 2197 4876 2203
rect 4948 2197 4956 2203
rect 4996 2197 5004 2203
rect 5044 2197 5084 2203
rect 5252 2197 5324 2203
rect 5460 2197 5500 2203
rect 1997 2177 2108 2183
rect 2308 2177 2332 2183
rect 2388 2177 2428 2183
rect 2452 2177 2956 2183
rect 2996 2177 3004 2183
rect 3236 2177 3340 2183
rect 3428 2177 3516 2183
rect 3604 2177 3660 2183
rect 3668 2177 3708 2183
rect 3748 2177 3772 2183
rect 3844 2177 3852 2183
rect 3892 2177 3980 2183
rect 4132 2177 4236 2183
rect 4372 2177 4492 2183
rect 4612 2177 4620 2183
rect 4676 2177 4684 2183
rect 4708 2177 5148 2183
rect 5156 2177 5196 2183
rect 5236 2177 5308 2183
rect 5412 2177 5564 2183
rect 308 2157 716 2163
rect 772 2157 1116 2163
rect 1124 2157 1148 2163
rect 1236 2157 1404 2163
rect 1540 2157 1548 2163
rect 1588 2157 1916 2163
rect 1940 2157 2060 2163
rect 2068 2157 2428 2163
rect 2468 2157 2508 2163
rect 2516 2157 2604 2163
rect 2692 2157 2700 2163
rect 2836 2157 2892 2163
rect 3005 2157 3020 2163
rect 765 2144 771 2156
rect 1469 2144 1475 2156
rect 116 2137 172 2143
rect 484 2137 492 2143
rect 532 2137 540 2143
rect 660 2137 668 2143
rect 708 2137 732 2143
rect 868 2137 892 2143
rect 916 2137 1196 2143
rect 1204 2137 1468 2143
rect 1524 2137 1596 2143
rect 1709 2137 1724 2143
rect 1748 2137 2124 2143
rect 2228 2137 2236 2143
rect 2276 2137 2284 2143
rect 2308 2137 2444 2143
rect 2564 2137 2572 2143
rect 2644 2137 2780 2143
rect 3005 2143 3011 2157
rect 3092 2157 3404 2163
rect 3524 2157 3548 2163
rect 3556 2157 3612 2163
rect 3661 2157 3676 2163
rect 3085 2144 3091 2156
rect 3661 2144 3667 2157
rect 3844 2157 3900 2163
rect 3940 2157 3964 2163
rect 4093 2157 4108 2163
rect 4228 2157 4252 2163
rect 4276 2157 4412 2163
rect 4420 2157 4812 2163
rect 4820 2157 4828 2163
rect 4836 2157 5212 2163
rect 5396 2157 5420 2163
rect 2836 2137 3011 2143
rect 3028 2137 3052 2143
rect 3108 2137 3132 2143
rect 3140 2137 3628 2143
rect 3636 2137 3644 2143
rect 3716 2137 3724 2143
rect 3812 2137 3900 2143
rect 3908 2137 3980 2143
rect 4068 2137 4508 2143
rect 4564 2137 4579 2143
rect 4596 2137 4748 2143
rect 4852 2137 4988 2143
rect 5012 2137 5052 2143
rect 5108 2137 5116 2143
rect 5268 2137 5372 2143
rect 5380 2137 5452 2143
rect 5492 2137 5516 2143
rect 2589 2124 2595 2136
rect -51 2103 -45 2123
rect 20 2117 252 2123
rect 260 2117 1068 2123
rect 1076 2117 1084 2123
rect 1092 2117 1388 2123
rect 1412 2117 1788 2123
rect 1956 2117 1996 2123
rect 2036 2117 2316 2123
rect 2612 2117 2652 2123
rect 2740 2117 2812 2123
rect 2996 2117 3004 2123
rect 3012 2117 3244 2123
rect 3252 2117 3660 2123
rect 2685 2104 2691 2116
rect 2925 2104 2931 2116
rect 3533 2104 3539 2117
rect 3684 2117 4044 2123
rect 4052 2117 4092 2123
rect 4100 2117 4396 2123
rect 4420 2117 4428 2123
rect 4436 2117 4460 2123
rect 4541 2117 4556 2123
rect 4612 2117 4684 2123
rect 4852 2117 4860 2123
rect 4900 2117 4956 2123
rect 4996 2117 5068 2123
rect 5092 2117 5132 2123
rect 5172 2117 5180 2123
rect -51 2097 12 2103
rect 244 2097 348 2103
rect 404 2097 460 2103
rect 548 2097 652 2103
rect 660 2097 748 2103
rect 756 2097 828 2103
rect 836 2097 1228 2103
rect 1268 2097 1292 2103
rect 1460 2097 1484 2103
rect 1588 2097 1676 2103
rect 1716 2097 1788 2103
rect 1940 2097 1980 2103
rect 2468 2097 2620 2103
rect 2980 2097 3148 2103
rect 3172 2097 3212 2103
rect 3252 2097 3500 2103
rect 3556 2097 3644 2103
rect 3652 2097 3740 2103
rect 3828 2097 3836 2103
rect 3876 2097 3932 2103
rect 3956 2097 3964 2103
rect 4052 2097 4188 2103
rect 4660 2097 4716 2103
rect 4916 2097 4924 2103
rect 4964 2097 5004 2103
rect 5028 2097 5036 2103
rect 5092 2097 5244 2103
rect 5300 2097 5516 2103
rect 1325 2084 1331 2096
rect 228 2077 908 2083
rect 1188 2077 1244 2083
rect 1460 2077 1772 2083
rect 2068 2077 2636 2083
rect 2644 2077 2988 2083
rect 3220 2077 3356 2083
rect 3389 2064 3395 2083
rect 3508 2077 3564 2083
rect 3572 2077 4636 2083
rect 4644 2077 5260 2083
rect 5268 2077 5340 2083
rect 5396 2077 5404 2083
rect 5460 2077 5468 2083
rect 1396 2057 2556 2063
rect 2612 2057 2620 2063
rect 3028 2057 3372 2063
rect 3476 2057 3516 2063
rect 4100 2057 4188 2063
rect 724 2037 1388 2043
rect 1684 2037 1820 2043
rect 1828 2037 2492 2043
rect 2772 2037 2940 2043
rect 2948 2037 3852 2043
rect 4660 2037 5356 2043
rect 1108 2017 1132 2023
rect 1652 2017 1868 2023
rect 3204 2017 3340 2023
rect 3380 2017 4268 2023
rect 845 2004 851 2016
rect 1172 1997 1196 2003
rect 1556 1997 1564 2003
rect 2004 1997 2108 2003
rect 2244 1997 2252 2003
rect 2948 1997 2956 2003
rect 4116 1997 4300 2003
rect 5437 1984 5443 1996
rect 820 1977 828 1983
rect 852 1977 1612 1983
rect 2228 1977 2684 1983
rect 2692 1977 2780 1983
rect 3204 1977 3260 1983
rect 3268 1977 3308 1983
rect 4020 1977 4092 1983
rect 4116 1977 4124 1983
rect 4932 1977 4988 1983
rect 708 1957 732 1963
rect 772 1957 796 1963
rect 820 1957 1180 1963
rect 1220 1957 1484 1963
rect 1620 1957 1724 1963
rect 1844 1957 1868 1963
rect 2052 1957 2092 1963
rect 2148 1957 2156 1963
rect 2452 1957 2460 1963
rect 2756 1957 3100 1963
rect 3108 1957 3180 1963
rect 3188 1957 3372 1963
rect 4052 1957 4140 1963
rect 4292 1957 4492 1963
rect 4676 1957 4764 1963
rect 4772 1957 4972 1963
rect 5140 1957 5244 1963
rect 68 1937 844 1943
rect 1076 1937 1180 1943
rect 1828 1937 1900 1943
rect 1924 1937 2524 1943
rect 2532 1937 2684 1943
rect 2852 1937 2892 1943
rect 3268 1937 3388 1943
rect 3524 1937 4364 1943
rect 4740 1937 4956 1943
rect 5060 1937 5164 1943
rect 5252 1937 5276 1943
rect 5348 1937 5420 1943
rect 452 1917 460 1923
rect 500 1917 1004 1923
rect 1012 1917 1260 1923
rect 1300 1917 1356 1923
rect 1668 1917 1852 1923
rect 1956 1917 1964 1923
rect 2084 1917 2476 1923
rect 2484 1917 2652 1923
rect 2724 1917 2732 1923
rect 2884 1917 3148 1923
rect 3300 1917 3516 1923
rect 3588 1917 3676 1923
rect 3732 1917 3740 1923
rect 4100 1917 4204 1923
rect 4260 1917 4300 1923
rect 4388 1917 4428 1923
rect 4484 1917 4604 1923
rect 4612 1917 4748 1923
rect 4788 1917 4844 1923
rect 4900 1917 4908 1923
rect 4964 1917 5068 1923
rect 5380 1917 5468 1923
rect 349 1904 355 1916
rect -51 1897 140 1903
rect 628 1897 860 1903
rect 884 1897 892 1903
rect 932 1897 940 1903
rect 996 1897 1020 1903
rect 1028 1897 1212 1903
rect 1220 1897 1980 1903
rect 1988 1897 2252 1903
rect 2260 1897 2572 1903
rect 2596 1897 2620 1903
rect 2852 1897 2972 1903
rect 3060 1897 3196 1903
rect 3620 1897 3692 1903
rect 3716 1897 3740 1903
rect 3844 1897 4076 1903
rect 4116 1897 4124 1903
rect 4132 1897 4268 1903
rect 4500 1897 4620 1903
rect 4644 1897 4716 1903
rect 4788 1897 4812 1903
rect 4836 1897 5292 1903
rect 116 1877 172 1883
rect 212 1877 236 1883
rect 340 1877 380 1883
rect 516 1877 1420 1883
rect 1508 1877 1676 1883
rect 1725 1877 1804 1883
rect 148 1857 284 1863
rect 372 1857 396 1863
rect 628 1857 748 1863
rect 772 1857 908 1863
rect 980 1857 1068 1863
rect 1092 1857 1203 1863
rect 589 1843 595 1856
rect 580 1837 595 1843
rect 612 1837 668 1843
rect 692 1837 700 1843
rect 724 1837 748 1843
rect 772 1837 972 1843
rect 1044 1837 1068 1843
rect 1076 1837 1116 1843
rect 1156 1837 1164 1843
rect 1197 1843 1203 1857
rect 1236 1857 1244 1863
rect 1284 1857 1324 1863
rect 1380 1857 1452 1863
rect 1469 1863 1475 1876
rect 1469 1857 1484 1863
rect 1572 1857 1596 1863
rect 1725 1863 1731 1877
rect 1892 1877 2428 1883
rect 2516 1877 2748 1883
rect 2829 1883 2835 1896
rect 3421 1884 3427 1896
rect 2829 1877 2844 1883
rect 2916 1877 2924 1883
rect 2948 1877 3420 1883
rect 3428 1877 3852 1883
rect 3805 1864 3811 1877
rect 3860 1877 3884 1883
rect 4164 1877 4236 1883
rect 4324 1877 4332 1883
rect 4404 1877 4460 1883
rect 4468 1877 4700 1883
rect 4916 1877 5004 1883
rect 5028 1877 5036 1883
rect 5076 1877 5084 1883
rect 5300 1877 5388 1883
rect 5396 1877 5404 1883
rect 5508 1877 5523 1883
rect 1684 1857 1731 1863
rect 1748 1857 1772 1863
rect 1876 1857 1884 1863
rect 1956 1857 1996 1863
rect 2052 1857 2124 1863
rect 2180 1857 2236 1863
rect 2244 1857 2316 1863
rect 2340 1857 2348 1863
rect 2628 1857 2988 1863
rect 3012 1857 3020 1863
rect 3028 1857 3036 1863
rect 3060 1857 3084 1863
rect 3092 1857 3228 1863
rect 3236 1857 3548 1863
rect 3732 1857 3756 1863
rect 3972 1857 3980 1863
rect 4420 1857 4572 1863
rect 4580 1857 4636 1863
rect 4692 1857 4700 1863
rect 4740 1857 5228 1863
rect 3709 1844 3715 1856
rect 1197 1837 1228 1843
rect 1284 1837 2108 1843
rect 2116 1837 2268 1843
rect 2292 1837 2300 1843
rect 2468 1837 2492 1843
rect 2836 1837 2940 1843
rect 2996 1837 3548 1843
rect 3652 1837 3699 1843
rect 356 1817 380 1823
rect 388 1817 460 1823
rect 468 1817 1324 1823
rect 1396 1817 1404 1823
rect 1796 1817 2060 1823
rect 2100 1817 2140 1823
rect 2580 1817 2636 1823
rect 3693 1823 3699 1837
rect 3780 1837 3852 1843
rect 3860 1837 3964 1843
rect 4100 1837 4108 1843
rect 4196 1837 4540 1843
rect 4548 1837 4572 1843
rect 4628 1837 5180 1843
rect 5204 1837 5276 1843
rect 3693 1817 3788 1823
rect 4788 1817 4812 1823
rect 4836 1817 4844 1823
rect 5236 1817 5564 1823
rect 68 1797 412 1803
rect 420 1797 1276 1803
rect 1348 1797 1500 1803
rect 1540 1797 1596 1803
rect 1620 1797 1731 1803
rect 52 1777 140 1783
rect 340 1777 444 1783
rect 468 1777 556 1783
rect 653 1777 844 1783
rect 52 1757 60 1763
rect 196 1757 428 1763
rect 436 1757 524 1763
rect 653 1763 659 1777
rect 900 1777 908 1783
rect 948 1777 956 1783
rect 980 1777 1004 1783
rect 1028 1777 1036 1783
rect 1156 1777 1164 1783
rect 1172 1777 1324 1783
rect 1460 1777 1468 1783
rect 1492 1777 1548 1783
rect 1668 1777 1676 1783
rect 1725 1783 1731 1797
rect 1748 1797 1980 1803
rect 2068 1797 2124 1803
rect 2260 1797 2268 1803
rect 2292 1797 2428 1803
rect 2708 1797 2716 1803
rect 2836 1797 2908 1803
rect 3220 1797 3244 1803
rect 3284 1797 3292 1803
rect 3364 1797 3404 1803
rect 3492 1797 3500 1803
rect 3748 1797 3772 1803
rect 4196 1797 4220 1803
rect 4356 1797 4364 1803
rect 4420 1797 4428 1803
rect 4724 1797 4748 1803
rect 4756 1797 4988 1803
rect 5252 1797 5276 1803
rect 5380 1797 5436 1803
rect 5540 1797 5564 1803
rect 1725 1777 1788 1783
rect 1892 1777 1948 1783
rect 1956 1777 2300 1783
rect 2436 1777 2492 1783
rect 2532 1777 2572 1783
rect 2612 1777 2748 1783
rect 2820 1777 2876 1783
rect 2964 1777 3196 1783
rect 3268 1777 3324 1783
rect 3572 1777 3580 1783
rect 3604 1777 3660 1783
rect 3988 1777 3996 1783
rect 4084 1777 4092 1783
rect 4100 1777 4284 1783
rect 4308 1777 4332 1783
rect 4340 1777 4876 1783
rect 4884 1777 5132 1783
rect 5284 1777 5292 1783
rect 580 1757 659 1763
rect 692 1757 812 1763
rect 820 1757 828 1763
rect 900 1757 1180 1763
rect 1188 1757 2060 1763
rect 2100 1757 2188 1763
rect 2244 1757 2284 1763
rect 2308 1757 2316 1763
rect 2388 1757 2396 1763
rect 2420 1757 2604 1763
rect 2612 1757 2636 1763
rect 2676 1757 2908 1763
rect 3188 1757 3436 1763
rect 3444 1757 3676 1763
rect 3780 1757 3788 1763
rect 3860 1757 3980 1763
rect 4100 1757 4108 1763
rect 4148 1757 4604 1763
rect 4612 1757 4620 1763
rect 4644 1757 4892 1763
rect 4996 1757 5004 1763
rect 5060 1757 5068 1763
rect 5092 1757 5260 1763
rect 5268 1757 5340 1763
rect 5380 1757 5500 1763
rect 132 1737 268 1743
rect 276 1737 444 1743
rect 516 1737 524 1743
rect 532 1737 1404 1743
rect 1412 1737 1436 1743
rect 1444 1737 1852 1743
rect 1956 1737 2044 1743
rect 2084 1737 2268 1743
rect 2276 1737 2716 1743
rect 2724 1737 2764 1743
rect 2836 1737 2844 1743
rect 2884 1737 2892 1743
rect 2932 1737 2940 1743
rect 3028 1737 3084 1743
rect 3268 1737 3276 1743
rect 3396 1737 3644 1743
rect 3684 1737 3692 1743
rect 3700 1737 3836 1743
rect 3876 1737 4156 1743
rect 4260 1737 4476 1743
rect 4484 1737 4684 1743
rect 4708 1737 4892 1743
rect 4900 1737 5148 1743
rect 5300 1737 5315 1743
rect 5380 1737 5388 1743
rect 68 1717 204 1723
rect 308 1717 316 1723
rect 580 1717 604 1723
rect 628 1717 652 1723
rect 740 1717 764 1723
rect 788 1717 1244 1723
rect 1252 1717 1580 1723
rect 1620 1717 1708 1723
rect 1748 1717 1868 1723
rect 1892 1717 2028 1723
rect 2084 1717 2124 1723
rect 2292 1717 2300 1723
rect 2340 1717 2396 1723
rect 2420 1717 2428 1723
rect 2452 1717 2460 1723
rect 2548 1717 2572 1723
rect 2804 1717 3004 1723
rect 3012 1717 3116 1723
rect 3140 1717 3436 1723
rect 3444 1717 3468 1723
rect 3556 1717 4316 1723
rect 4324 1717 4940 1723
rect 4948 1717 5004 1723
rect 5044 1717 5324 1723
rect 260 1697 380 1703
rect 500 1697 508 1703
rect 548 1697 556 1703
rect 564 1697 796 1703
rect 884 1697 924 1703
rect 1124 1697 1132 1703
rect 1204 1697 1644 1703
rect 1652 1697 1996 1703
rect 2004 1697 2092 1703
rect 2244 1697 2700 1703
rect 2948 1697 2988 1703
rect 2996 1697 3052 1703
rect 3060 1697 3356 1703
rect 3364 1697 3372 1703
rect 3460 1697 3532 1703
rect 3652 1697 3708 1703
rect 3716 1697 3724 1703
rect 3828 1697 3852 1703
rect 3924 1697 3932 1703
rect 3949 1697 3980 1703
rect 116 1677 220 1683
rect 228 1677 924 1683
rect 1140 1677 1404 1683
rect 1460 1677 1676 1683
rect 1844 1677 1900 1683
rect 1924 1677 2012 1683
rect 2020 1677 2364 1683
rect 2452 1677 2604 1683
rect 3300 1677 3340 1683
rect 3620 1677 3836 1683
rect 3949 1683 3955 1697
rect 4020 1697 4124 1703
rect 4132 1697 4588 1703
rect 4596 1697 4700 1703
rect 4932 1697 4940 1703
rect 4964 1697 5052 1703
rect 5124 1697 5292 1703
rect 3844 1677 3955 1683
rect 3972 1677 4060 1683
rect 4180 1677 4204 1683
rect 4324 1677 4348 1683
rect 4420 1677 4556 1683
rect 4692 1677 4748 1683
rect 4820 1677 4828 1683
rect 1108 1657 1132 1663
rect 3732 1657 3740 1663
rect 3924 1657 3996 1663
rect 4292 1657 4508 1663
rect 4532 1657 4684 1663
rect 4804 1657 4812 1663
rect 1156 1637 1180 1643
rect 1188 1637 1196 1643
rect 1412 1637 1564 1643
rect 1988 1637 2108 1643
rect 2548 1637 2588 1643
rect 84 1617 108 1623
rect 116 1617 140 1623
rect 196 1617 204 1623
rect 1924 1617 1948 1623
rect 2228 1617 2364 1623
rect 4516 1617 5196 1623
rect 3725 1604 3731 1616
rect 500 1597 716 1603
rect 724 1597 1244 1603
rect 1524 1597 1548 1603
rect 1908 1597 1932 1603
rect 2436 1597 2444 1603
rect 2660 1597 2700 1603
rect 3012 1597 3084 1603
rect 3252 1597 3324 1603
rect 4276 1597 4364 1603
rect 4772 1597 4860 1603
rect 4932 1597 5532 1603
rect 1677 1584 1683 1596
rect 3716 1577 3724 1583
rect 4356 1577 4492 1583
rect 4644 1577 4652 1583
rect 4788 1577 4796 1583
rect 4868 1577 4988 1583
rect 5364 1577 5388 1583
rect 772 1557 1036 1563
rect 1588 1557 1596 1563
rect 1652 1557 1660 1563
rect 2036 1557 2060 1563
rect 3508 1557 4732 1563
rect 4740 1557 5004 1563
rect 5028 1557 5116 1563
rect 628 1537 636 1543
rect 836 1537 860 1543
rect 1012 1537 1020 1543
rect 1076 1537 1116 1543
rect 1124 1537 1164 1543
rect 1396 1537 1420 1543
rect 1588 1537 1612 1543
rect 2180 1537 2236 1543
rect 3172 1537 3276 1543
rect 3460 1537 3468 1543
rect 3572 1537 3580 1543
rect 3604 1537 3612 1543
rect 3700 1537 3724 1543
rect 4036 1537 4124 1543
rect 4148 1537 4172 1543
rect 4228 1537 4252 1543
rect 4276 1537 4796 1543
rect 4804 1537 4876 1543
rect 4948 1537 4956 1543
rect 4980 1537 5100 1543
rect 5188 1537 5420 1543
rect 1197 1524 1203 1536
rect 3805 1524 3811 1536
rect 388 1517 396 1523
rect 404 1517 1020 1523
rect 1028 1517 1196 1523
rect 1204 1517 1228 1523
rect 1252 1517 1452 1523
rect 1636 1517 1740 1523
rect 1812 1517 1852 1523
rect 1876 1517 1900 1523
rect 2036 1517 2172 1523
rect 2180 1517 2284 1523
rect 2340 1517 2428 1523
rect 2484 1517 2572 1523
rect 2900 1517 3052 1523
rect 3076 1517 3148 1523
rect 3220 1517 3756 1523
rect 3908 1517 4044 1523
rect 4052 1517 4140 1523
rect 4164 1517 4412 1523
rect 4420 1517 4556 1523
rect 4628 1517 4652 1523
rect 4708 1517 4748 1523
rect 4772 1517 4796 1523
rect 4916 1517 5276 1523
rect 5300 1517 5324 1523
rect 5380 1517 5452 1523
rect 2797 1504 2803 1516
rect 5533 1504 5539 1516
rect 180 1497 460 1503
rect 596 1497 604 1503
rect 644 1497 700 1503
rect 1156 1497 1180 1503
rect 1188 1497 1212 1503
rect 1284 1497 1324 1503
rect 1364 1497 1452 1503
rect 1492 1497 1500 1503
rect 1636 1497 1644 1503
rect 1668 1497 2236 1503
rect 2253 1497 2444 1503
rect 829 1484 835 1496
rect 132 1477 172 1483
rect 324 1477 716 1483
rect 884 1477 940 1483
rect 1092 1477 1100 1483
rect 1124 1477 1148 1483
rect 1220 1477 1468 1483
rect 1524 1477 1580 1483
rect 1604 1477 1708 1483
rect 1716 1477 1740 1483
rect 1764 1477 1772 1483
rect 1876 1477 1884 1483
rect 1972 1477 2188 1483
rect 2253 1483 2259 1497
rect 2564 1497 2604 1503
rect 2628 1497 2748 1503
rect 2964 1497 3244 1503
rect 3268 1497 3276 1503
rect 3300 1497 3340 1503
rect 3460 1497 3484 1503
rect 3508 1497 3692 1503
rect 3796 1497 3852 1503
rect 3908 1497 3932 1503
rect 3940 1497 3948 1503
rect 4100 1497 4428 1503
rect 4484 1497 4876 1503
rect 4884 1497 4924 1503
rect 5044 1497 5084 1503
rect 5124 1497 5244 1503
rect 2212 1477 2259 1483
rect 2356 1477 2508 1483
rect 2516 1477 2732 1483
rect 2788 1477 2908 1483
rect 2916 1477 2956 1483
rect 2980 1477 3084 1483
rect 3092 1477 3676 1483
rect 3684 1477 3692 1483
rect 3700 1477 3868 1483
rect 3876 1477 4236 1483
rect 4468 1477 4956 1483
rect 4973 1477 4979 1496
rect 5172 1477 5196 1483
rect 68 1457 76 1463
rect 180 1457 188 1463
rect 484 1457 492 1463
rect 580 1457 588 1463
rect 644 1457 652 1463
rect 772 1457 780 1463
rect 788 1457 940 1463
rect 957 1457 972 1463
rect 1108 1457 1132 1463
rect 1172 1457 1292 1463
rect 1332 1457 1340 1463
rect 1380 1457 1388 1463
rect 1492 1457 1500 1463
rect 1508 1457 1852 1463
rect 1908 1457 2124 1463
rect 2132 1457 2316 1463
rect 2388 1457 2396 1463
rect 2948 1457 3148 1463
rect 3204 1457 3260 1463
rect 3268 1457 3420 1463
rect 3428 1457 3628 1463
rect 3652 1457 3660 1463
rect 3700 1457 3724 1463
rect 3780 1457 3852 1463
rect 3924 1457 3996 1463
rect 4004 1457 4076 1463
rect 4100 1457 4156 1463
rect 4180 1457 4188 1463
rect 4212 1457 4508 1463
rect 4516 1457 4588 1463
rect 4612 1457 4844 1463
rect 4852 1457 5132 1463
rect 5140 1457 5196 1463
rect 644 1437 780 1443
rect 900 1437 972 1443
rect 980 1437 1116 1443
rect 1252 1437 1260 1443
rect 1268 1437 2380 1443
rect 2692 1437 2764 1443
rect 2781 1437 2812 1443
rect 660 1417 844 1423
rect 1076 1417 1100 1423
rect 1524 1417 1532 1423
rect 1588 1417 1596 1423
rect 1620 1417 1628 1423
rect 1732 1417 1804 1423
rect 1812 1417 1964 1423
rect 1972 1417 2092 1423
rect 2132 1417 2156 1423
rect 2781 1423 2787 1437
rect 2820 1437 2956 1443
rect 3092 1437 3132 1443
rect 3252 1437 3260 1443
rect 3268 1437 3548 1443
rect 3556 1437 3676 1443
rect 3924 1437 3932 1443
rect 4244 1437 4396 1443
rect 4404 1437 4412 1443
rect 4436 1437 4732 1443
rect 4740 1437 4812 1443
rect 5188 1437 5308 1443
rect 2708 1417 2787 1423
rect 3540 1417 3548 1423
rect 3572 1417 3580 1423
rect 3940 1417 4044 1423
rect 4820 1417 4828 1423
rect 4836 1417 4988 1423
rect 196 1397 972 1403
rect 1028 1397 1036 1403
rect 1348 1397 1356 1403
rect 1540 1397 1548 1403
rect 1764 1397 1772 1403
rect 1844 1397 1996 1403
rect 2116 1397 2124 1403
rect 2308 1397 2444 1403
rect 3012 1397 3020 1403
rect 3380 1397 3404 1403
rect 3412 1397 3484 1403
rect 3492 1397 3932 1403
rect 3956 1397 4044 1403
rect 4116 1397 4124 1403
rect 5124 1397 5452 1403
rect 324 1377 364 1383
rect 708 1377 780 1383
rect 996 1377 1004 1383
rect 1012 1377 1084 1383
rect 1188 1377 1212 1383
rect 1268 1377 1420 1383
rect 1524 1377 1660 1383
rect 1700 1377 2060 1383
rect 2068 1377 2908 1383
rect 3204 1377 3244 1383
rect 3284 1377 3308 1383
rect 3396 1377 3436 1383
rect 3460 1377 3468 1383
rect 3540 1377 3660 1383
rect 3668 1377 3692 1383
rect 3716 1377 4476 1383
rect 4484 1377 4492 1383
rect 4548 1377 4572 1383
rect 4852 1377 4924 1383
rect 5252 1377 5324 1383
rect 5332 1377 5340 1383
rect 5364 1377 5372 1383
rect 5412 1377 5452 1383
rect 1677 1364 1683 1376
rect 84 1357 108 1363
rect 132 1357 140 1363
rect 452 1357 460 1363
rect 516 1357 572 1363
rect 580 1357 620 1363
rect 644 1357 716 1363
rect 740 1357 844 1363
rect 964 1357 1052 1363
rect 1076 1357 1340 1363
rect 1412 1357 1612 1363
rect 1716 1357 1804 1363
rect 1860 1357 2076 1363
rect 2100 1357 2140 1363
rect 2148 1357 2412 1363
rect 2596 1357 2684 1363
rect 2756 1357 2828 1363
rect 3108 1357 3116 1363
rect 3252 1357 3260 1363
rect 3268 1357 3292 1363
rect 3332 1357 3340 1363
rect 3396 1357 3404 1363
rect 3492 1357 3596 1363
rect 3620 1357 3644 1363
rect 3700 1357 3756 1363
rect 3796 1357 3820 1363
rect 3876 1357 3884 1363
rect 4020 1357 4028 1363
rect 4100 1357 4147 1363
rect 2509 1344 2515 1356
rect 228 1337 332 1343
rect 436 1337 460 1343
rect 532 1337 540 1343
rect 596 1337 764 1343
rect 820 1337 828 1343
rect 836 1337 1100 1343
rect 1156 1337 1164 1343
rect 1204 1337 1292 1343
rect 1380 1337 1388 1343
rect 1428 1337 1596 1343
rect 1604 1337 1948 1343
rect 1956 1337 2044 1343
rect 2052 1337 2236 1343
rect 2308 1337 2444 1343
rect 2548 1337 2636 1343
rect 2724 1337 3420 1343
rect 3428 1337 3836 1343
rect 3892 1337 3948 1343
rect 3972 1337 4124 1343
rect 4141 1343 4147 1357
rect 4164 1357 4188 1363
rect 4244 1357 4620 1363
rect 4788 1357 4796 1363
rect 4868 1357 4908 1363
rect 5044 1357 5052 1363
rect 5140 1357 5196 1363
rect 5316 1357 5324 1363
rect 4141 1337 4236 1343
rect 4388 1337 4556 1343
rect 4580 1337 4796 1343
rect 4852 1337 5260 1343
rect 5316 1337 5331 1343
rect 5325 1324 5331 1337
rect 5412 1337 5500 1343
rect 196 1317 252 1323
rect 260 1317 268 1323
rect 276 1317 460 1323
rect 484 1317 540 1323
rect 548 1317 1212 1323
rect 1348 1317 1852 1323
rect 1892 1317 2124 1323
rect 2132 1317 2348 1323
rect 2356 1317 2524 1323
rect 2564 1317 2620 1323
rect 2708 1317 2764 1323
rect 2884 1317 3180 1323
rect 3204 1317 3580 1323
rect 3748 1317 4108 1323
rect 4132 1317 4172 1323
rect 4292 1317 4364 1323
rect 4436 1317 4476 1323
rect 4596 1317 4604 1323
rect 4740 1317 5148 1323
rect 5156 1317 5276 1323
rect 628 1297 748 1303
rect 756 1297 844 1303
rect 932 1297 940 1303
rect 948 1297 1612 1303
rect 1732 1297 1868 1303
rect 1892 1297 1900 1303
rect 1908 1297 1932 1303
rect 2052 1297 2108 1303
rect 2180 1297 2268 1303
rect 2340 1297 2348 1303
rect 2388 1297 2460 1303
rect 2500 1297 2508 1303
rect 2660 1297 2780 1303
rect 2788 1297 2796 1303
rect 2916 1297 2956 1303
rect 3012 1297 3020 1303
rect 3044 1297 3116 1303
rect 3156 1297 4156 1303
rect 4212 1297 4236 1303
rect 4260 1297 4291 1303
rect 388 1277 460 1283
rect 468 1277 636 1283
rect 836 1277 908 1283
rect 1044 1277 1228 1283
rect 1460 1277 1628 1283
rect 1812 1277 1932 1283
rect 2164 1277 2236 1283
rect 2372 1277 2492 1283
rect 2708 1277 2716 1283
rect 2772 1277 2780 1283
rect 2948 1277 3164 1283
rect 3188 1277 3564 1283
rect 3780 1277 3884 1283
rect 3908 1277 3948 1283
rect 3988 1277 4076 1283
rect 4084 1277 4140 1283
rect 4244 1277 4268 1283
rect 4285 1283 4291 1297
rect 4308 1297 4316 1303
rect 4333 1297 4508 1303
rect 4333 1283 4339 1297
rect 4676 1297 4748 1303
rect 5060 1297 5196 1303
rect 5316 1297 5484 1303
rect 4285 1277 4339 1283
rect 4372 1277 4828 1283
rect 4980 1277 5084 1283
rect 5092 1277 5388 1283
rect 1341 1264 1347 1276
rect 820 1257 1036 1263
rect 1604 1257 1772 1263
rect 2724 1257 2732 1263
rect 3300 1257 3308 1263
rect 3316 1257 3340 1263
rect 3524 1257 3596 1263
rect 3604 1257 4812 1263
rect 3213 1244 3219 1256
rect 1156 1237 1164 1243
rect 1396 1237 2220 1243
rect 2228 1237 2380 1243
rect 3332 1237 3660 1243
rect 3668 1237 4060 1243
rect 4813 1224 4819 1236
rect 52 1217 60 1223
rect 1092 1217 1116 1223
rect 3460 1217 3516 1223
rect 3524 1217 3788 1223
rect 52 1197 76 1203
rect 148 1197 204 1203
rect 1460 1197 1836 1203
rect 2324 1197 2380 1203
rect 2452 1197 2540 1203
rect 3620 1197 3660 1203
rect 4724 1197 5068 1203
rect 5188 1197 5388 1203
rect 276 1177 780 1183
rect 1684 1177 1788 1183
rect 1812 1177 2252 1183
rect 2452 1177 2524 1183
rect 3140 1177 3148 1183
rect 3716 1177 3724 1183
rect 3908 1177 3948 1183
rect 4100 1177 5068 1183
rect 5076 1177 5084 1183
rect 68 1157 236 1163
rect 260 1157 284 1163
rect 292 1157 556 1163
rect 1316 1157 1420 1163
rect 1428 1157 1612 1163
rect 2004 1157 2364 1163
rect 2372 1157 2476 1163
rect 3300 1157 3804 1163
rect 3940 1157 4428 1163
rect 4612 1157 4876 1163
rect 4884 1157 5324 1163
rect 532 1137 540 1143
rect 756 1137 1052 1143
rect 1060 1137 1068 1143
rect 1172 1137 1260 1143
rect 1284 1137 1292 1143
rect 1396 1137 1596 1143
rect 1620 1137 1836 1143
rect 1844 1137 2044 1143
rect 2052 1137 2604 1143
rect 2861 1137 2892 1143
rect -51 1117 268 1123
rect -51 1097 -45 1117
rect 356 1117 412 1123
rect 452 1117 1004 1123
rect 1012 1117 1116 1123
rect 1124 1117 1196 1123
rect 1396 1117 1404 1123
rect 1764 1117 1772 1123
rect 1796 1117 1804 1123
rect 1956 1117 1964 1123
rect 1988 1117 2044 1123
rect 2084 1117 2332 1123
rect 2340 1117 2540 1123
rect 2861 1123 2867 1137
rect 3796 1137 3980 1143
rect 4340 1137 5052 1143
rect 5172 1137 5212 1143
rect 5316 1137 5420 1143
rect 2676 1117 2867 1123
rect 2884 1117 3020 1123
rect 3268 1117 3308 1123
rect 3444 1117 3452 1123
rect 3588 1117 3804 1123
rect 3956 1117 3964 1123
rect 4100 1117 4140 1123
rect 4340 1117 4348 1123
rect 4372 1117 4588 1123
rect 4628 1117 4652 1123
rect 4692 1117 4700 1123
rect 4740 1117 4748 1123
rect 4820 1117 4828 1123
rect 4884 1117 4908 1123
rect 4980 1117 4988 1123
rect 5028 1117 5324 1123
rect 180 1097 188 1103
rect 228 1097 812 1103
rect 836 1097 972 1103
rect 980 1097 2092 1103
rect 2100 1097 2316 1103
rect 2404 1097 2764 1103
rect 2772 1097 2796 1103
rect 2820 1097 2924 1103
rect 3012 1097 3196 1103
rect 3364 1097 3548 1103
rect 3684 1097 3692 1103
rect 3812 1097 3868 1103
rect 3876 1097 3996 1103
rect 4052 1097 4060 1103
rect 4164 1097 4236 1103
rect 4276 1097 4460 1103
rect 4468 1097 4844 1103
rect 4884 1097 5004 1103
rect 5012 1097 5148 1103
rect 5188 1097 5244 1103
rect 5300 1097 5436 1103
rect 36 1077 44 1083
rect 212 1077 764 1083
rect 772 1077 860 1083
rect 868 1077 1212 1083
rect 1220 1077 1228 1083
rect 1277 1077 1292 1083
rect 1316 1077 1324 1083
rect 1348 1077 1372 1083
rect 1428 1077 1436 1083
rect 1492 1077 1644 1083
rect 1652 1077 1660 1083
rect 1668 1077 1836 1083
rect 1853 1077 2268 1083
rect 173 1064 179 1076
rect 205 1064 211 1076
rect 132 1057 140 1063
rect 292 1057 300 1063
rect 468 1057 748 1063
rect 756 1057 860 1063
rect 996 1057 1420 1063
rect 1476 1057 1484 1063
rect 1636 1057 1660 1063
rect 1732 1057 1740 1063
rect 1853 1063 1859 1077
rect 2404 1077 2412 1083
rect 2452 1077 2812 1083
rect 2868 1077 2956 1083
rect 3060 1077 3228 1083
rect 3380 1077 3820 1083
rect 3844 1077 4140 1083
rect 4148 1077 4412 1083
rect 4500 1077 4540 1083
rect 4628 1077 4636 1083
rect 4644 1077 4780 1083
rect 4788 1077 5132 1083
rect 5172 1077 5196 1083
rect 5236 1077 5356 1083
rect 5364 1077 5468 1083
rect 1748 1057 1859 1063
rect 1876 1057 1900 1063
rect 1956 1057 2108 1063
rect 2212 1057 2236 1063
rect 2436 1057 2700 1063
rect 3012 1057 3436 1063
rect 3460 1057 3628 1063
rect 3732 1057 3740 1063
rect 3764 1057 3916 1063
rect 4020 1057 4364 1063
rect 4420 1057 4476 1063
rect 4484 1057 4492 1063
rect 4532 1057 4796 1063
rect 4804 1057 5084 1063
rect 5092 1057 5276 1063
rect 5284 1057 5452 1063
rect 68 1037 275 1043
rect 196 1017 236 1023
rect 269 1023 275 1037
rect 292 1037 316 1043
rect 516 1037 780 1043
rect 836 1037 844 1043
rect 1108 1037 1116 1043
rect 1236 1037 1292 1043
rect 1332 1037 1500 1043
rect 1716 1037 1820 1043
rect 1828 1037 1868 1043
rect 1924 1037 1948 1043
rect 2180 1037 2300 1043
rect 2532 1037 2700 1043
rect 3076 1037 3116 1043
rect 3156 1037 3324 1043
rect 3524 1037 3644 1043
rect 3732 1037 3788 1043
rect 3796 1037 3852 1043
rect 4036 1037 4124 1043
rect 4132 1037 4364 1043
rect 4612 1037 4652 1043
rect 4948 1037 4956 1043
rect 5300 1037 5452 1043
rect 2493 1024 2499 1036
rect 269 1017 332 1023
rect 692 1017 700 1023
rect 820 1017 828 1023
rect 964 1017 1132 1023
rect 1140 1017 1164 1023
rect 1396 1017 1740 1023
rect 1828 1017 1836 1023
rect 1860 1017 1884 1023
rect 1956 1017 1964 1023
rect 3076 1017 3084 1023
rect 3172 1017 3180 1023
rect 3268 1017 3276 1023
rect 3828 1017 3852 1023
rect 4660 1017 4748 1023
rect 5316 1017 5340 1023
rect 116 997 140 1003
rect 772 997 796 1003
rect 804 997 812 1003
rect 852 997 860 1003
rect 980 997 988 1003
rect 1028 997 1036 1003
rect 1380 997 1404 1003
rect 1972 997 1980 1003
rect 2196 997 2204 1003
rect 2244 997 2284 1003
rect 2436 997 2444 1003
rect 2708 997 2732 1003
rect 2820 997 2828 1003
rect 3268 997 3292 1003
rect 3652 997 3724 1003
rect 3988 997 4012 1003
rect 4228 997 4236 1003
rect 4244 997 4364 1003
rect 4660 997 4684 1003
rect 4708 997 4716 1003
rect 4884 997 4908 1003
rect 4932 997 4972 1003
rect 5044 997 5244 1003
rect 5373 997 5436 1003
rect 404 977 444 983
rect 564 977 572 983
rect 580 977 1500 983
rect 1524 977 1884 983
rect 1892 977 2252 983
rect 2292 977 2316 983
rect 2372 977 2572 983
rect 2596 977 2652 983
rect 2676 977 2684 983
rect 2788 977 2828 983
rect 3172 977 3324 983
rect 3348 977 3468 983
rect 3540 977 3564 983
rect 3684 977 3708 983
rect 3716 977 3740 983
rect 3748 977 3836 983
rect 3908 977 3948 983
rect 3972 977 4428 983
rect 4516 977 4716 983
rect 4724 977 5004 983
rect 5012 977 5132 983
rect 5140 977 5308 983
rect 5373 983 5379 997
rect 5364 977 5379 983
rect 5396 977 5452 983
rect 132 957 140 963
rect 260 957 268 963
rect 308 957 396 963
rect 420 957 556 963
rect 596 957 796 963
rect 804 957 1484 963
rect 1540 957 1676 963
rect 1748 957 1756 963
rect 1860 957 1996 963
rect 2068 957 2300 963
rect 2308 957 2476 963
rect 2500 957 2780 963
rect 2788 957 2828 963
rect 2836 957 3004 963
rect 3060 957 3084 963
rect 3220 957 3340 963
rect 3396 957 3404 963
rect 3844 957 3852 963
rect 3924 957 3932 963
rect 4052 957 4060 963
rect 4116 957 4316 963
rect 4356 957 4364 963
rect 4404 957 4620 963
rect 4628 957 5036 963
rect 5060 957 5100 963
rect 5124 957 5132 963
rect 5380 957 5388 963
rect 3453 944 3459 956
rect 180 937 188 943
rect 196 937 236 943
rect 244 937 444 943
rect 468 937 492 943
rect 644 937 684 943
rect 708 937 828 943
rect 900 937 924 943
rect 964 937 988 943
rect 1012 937 1020 943
rect 1060 937 1148 943
rect 1220 937 1324 943
rect 1412 937 1500 943
rect 1588 937 1596 943
rect 1604 937 2140 943
rect 2340 937 2348 943
rect 2404 937 2412 943
rect 2436 937 2444 943
rect 2548 937 2876 943
rect 2916 937 3068 943
rect 3092 937 3388 943
rect 3396 937 3420 943
rect 3652 937 4332 943
rect 4340 937 4444 943
rect 4516 937 4540 943
rect 4580 937 5052 943
rect 5108 937 5180 943
rect 5444 937 5500 943
rect 2221 924 2227 936
rect 2877 924 2883 936
rect 5405 924 5411 936
rect 388 917 1212 923
rect 1252 917 1260 923
rect 1492 917 1804 923
rect 1812 917 1868 923
rect 1892 917 2188 923
rect 2292 917 2396 923
rect 2404 917 2428 923
rect 2564 917 2620 923
rect 2628 917 2787 923
rect 292 897 348 903
rect 356 897 364 903
rect 372 897 1004 903
rect 1540 897 1644 903
rect 1668 897 1676 903
rect 1700 897 1932 903
rect 1956 897 2124 903
rect 2436 897 2716 903
rect 2724 897 2732 903
rect 2781 903 2787 917
rect 3284 917 3676 923
rect 3716 917 3740 923
rect 3764 917 3772 923
rect 3780 917 3836 923
rect 3860 917 3884 923
rect 3924 917 4012 923
rect 4212 917 4236 923
rect 4260 917 4956 923
rect 5092 917 5212 923
rect 5220 917 5388 923
rect 2781 897 2908 903
rect 2916 897 2956 903
rect 2964 897 2988 903
rect 3236 897 3276 903
rect 3380 897 3404 903
rect 3412 897 3756 903
rect 3853 897 4812 903
rect 180 877 412 883
rect 436 877 460 883
rect 516 877 524 883
rect 532 877 588 883
rect 900 877 908 883
rect 948 877 1324 883
rect 1348 877 1564 883
rect 2292 877 2476 883
rect 2500 877 2604 883
rect 2612 877 2716 883
rect 2724 877 2780 883
rect 2868 877 2892 883
rect 2948 877 3036 883
rect 3300 877 3356 883
rect 3853 883 3859 897
rect 4820 897 4956 903
rect 4980 897 5004 903
rect 5124 897 5212 903
rect 5316 897 5356 903
rect 5396 897 5484 903
rect 3524 877 3859 883
rect 4068 877 4076 883
rect 4212 877 4220 883
rect 4260 877 4396 883
rect 4452 877 4940 883
rect 4964 877 5164 883
rect 5268 877 5276 883
rect 900 857 1196 863
rect 1204 857 1500 863
rect 2244 857 2508 863
rect 2516 857 2780 863
rect 2868 857 2876 863
rect 3005 857 3244 863
rect 93 837 396 843
rect 93 823 99 837
rect 900 837 1132 843
rect 1140 837 2012 843
rect 2020 837 2028 843
rect 2036 837 2748 843
rect 3005 843 3011 857
rect 3668 857 3724 863
rect 4020 857 4252 863
rect 4276 857 4284 863
rect 4804 857 4812 863
rect 4301 844 4307 856
rect 2756 837 3011 843
rect 3108 837 3164 843
rect 3252 837 3484 843
rect 3524 837 3724 843
rect 4164 837 4172 843
rect 4484 837 4892 843
rect 4900 837 5132 843
rect 5172 837 5196 843
rect 68 817 99 823
rect 708 817 972 823
rect 1076 817 1084 823
rect 1236 817 1244 823
rect 1268 817 1356 823
rect 1556 817 1852 823
rect 2260 817 2268 823
rect 2852 817 2956 823
rect 3188 817 3196 823
rect 3396 817 3628 823
rect 4164 817 4188 823
rect 4420 817 4588 823
rect 20 797 44 803
rect 308 797 396 803
rect 1220 797 1228 803
rect 1268 797 1580 803
rect 1588 797 2076 803
rect 2084 797 2156 803
rect 2468 797 2492 803
rect 2500 797 3020 803
rect 3028 797 3052 803
rect 3060 797 3548 803
rect 3796 797 4028 803
rect 4036 797 4556 803
rect 260 777 556 783
rect 564 777 780 783
rect 884 777 1100 783
rect 1108 777 1676 783
rect 1764 777 1964 783
rect 2164 777 2188 783
rect 2276 777 2380 783
rect 2484 777 2540 783
rect 2573 777 2636 783
rect 468 757 684 763
rect 692 757 1180 763
rect 1188 757 1228 763
rect 1572 757 1580 763
rect 1620 757 1628 763
rect 1716 757 1852 763
rect 1956 757 1996 763
rect 2052 757 2268 763
rect 2573 763 2579 777
rect 2820 777 2940 783
rect 3076 777 3084 783
rect 3220 777 3228 783
rect 3524 777 3564 783
rect 4157 777 4172 783
rect 3661 764 3667 776
rect 2276 757 2579 763
rect 2628 757 2764 763
rect 2900 757 3164 763
rect 3588 757 3644 763
rect 3908 757 3932 763
rect 4029 757 4044 763
rect 484 737 828 743
rect 852 737 1868 743
rect 1876 737 2028 743
rect 2132 737 2140 743
rect 2180 737 2220 743
rect 2356 737 2364 743
rect 2436 737 2444 743
rect 2628 737 2876 743
rect 3092 737 3116 743
rect 3396 737 3468 743
rect 3661 737 4108 743
rect 429 724 435 736
rect 196 717 284 723
rect 484 717 588 723
rect 644 717 780 723
rect 797 717 812 723
rect 1044 717 1164 723
rect 1300 717 1420 723
rect 1444 717 1452 723
rect 1460 717 1964 723
rect 2148 717 2412 723
rect 2420 717 2492 723
rect 2548 717 2812 723
rect 2868 717 2908 723
rect 3028 717 3036 723
rect 3661 723 3667 737
rect 4157 743 4163 777
rect 4404 777 4652 783
rect 4196 757 4460 763
rect 4548 757 4556 763
rect 4580 757 4620 763
rect 4740 757 4812 763
rect 4820 757 4876 763
rect 5060 757 5116 763
rect 5124 757 5260 763
rect 4132 737 4163 743
rect 4173 743 4179 756
rect 5037 744 5043 756
rect 4173 737 4188 743
rect 4260 737 4268 743
rect 4292 737 4508 743
rect 4564 737 4668 743
rect 4788 737 4796 743
rect 5076 737 5196 743
rect 5252 737 5356 743
rect 5380 737 5500 743
rect 3044 717 3667 723
rect 3780 717 3820 723
rect 3844 717 4300 723
rect 4388 717 4492 723
rect 4516 717 4700 723
rect 4708 717 4860 723
rect 4868 717 5068 723
rect 5124 717 5132 723
rect 5268 717 5292 723
rect 260 697 268 703
rect 276 697 700 703
rect 708 697 1724 703
rect 1828 697 2092 703
rect 2100 697 2108 703
rect 2132 697 2492 703
rect 2532 697 2572 703
rect 2676 697 2796 703
rect 2804 697 2860 703
rect 3476 697 4188 703
rect 4196 697 4204 703
rect 4276 697 4284 703
rect 4308 697 4316 703
rect 4356 697 4380 703
rect 4500 697 4684 703
rect 4692 697 4844 703
rect 5044 697 5148 703
rect 5252 697 5276 703
rect 5284 697 5292 703
rect 5396 697 5452 703
rect 4861 684 4867 696
rect 4893 684 4899 696
rect 4941 684 4947 696
rect 196 677 220 683
rect 260 677 380 683
rect 388 677 780 683
rect 804 677 908 683
rect 964 677 972 683
rect 1012 677 1036 683
rect 1140 677 1148 683
rect 1172 677 1180 683
rect 1220 677 1404 683
rect 1412 677 1420 683
rect 1597 664 1603 683
rect 1636 677 2428 683
rect 2612 677 2828 683
rect 2900 677 3004 683
rect 3076 677 3084 683
rect 3172 677 3212 683
rect 3252 677 3260 683
rect 3284 677 3724 683
rect 3732 677 3740 683
rect 3812 677 3820 683
rect 3892 677 3948 683
rect 3972 677 4844 683
rect 5060 677 5132 683
rect 5140 677 5196 683
rect 5300 677 5308 683
rect 5364 677 5372 683
rect 1613 664 1619 676
rect 52 657 60 663
rect 132 657 204 663
rect 276 657 716 663
rect 724 657 1084 663
rect 1092 657 1276 663
rect 1428 657 1564 663
rect 1876 657 1948 663
rect 1988 657 2364 663
rect 2372 657 2508 663
rect 2516 657 2716 663
rect 2724 657 2892 663
rect 3076 657 3100 663
rect 3156 657 3276 663
rect 3364 657 3468 663
rect 3636 657 3644 663
rect 3652 657 3660 663
rect 3668 657 3964 663
rect 3988 657 3996 663
rect 4052 657 4060 663
rect 4116 657 4140 663
rect 4212 657 5084 663
rect 5108 657 5388 663
rect 4093 644 4099 656
rect 324 637 332 643
rect 356 637 460 643
rect 468 637 1308 643
rect 1428 637 1452 643
rect 1476 637 1532 643
rect 2116 637 2140 643
rect 3140 637 3276 643
rect 3284 637 3324 643
rect 3348 637 3372 643
rect 3508 637 3804 643
rect 3812 637 3932 643
rect 4132 637 5068 643
rect 5156 637 5404 643
rect 772 617 860 623
rect 1076 617 1212 623
rect 1220 617 1372 623
rect 1444 617 1484 623
rect 1508 617 1612 623
rect 1620 617 2044 623
rect 2452 617 2476 623
rect 2724 617 2748 623
rect 3028 617 3084 623
rect 3124 617 3148 623
rect 3252 617 3276 623
rect 3300 617 3324 623
rect 3364 617 3388 623
rect 3524 617 3836 623
rect 3844 617 3916 623
rect 4308 617 4428 623
rect 4452 617 4540 623
rect 100 597 108 603
rect 116 597 140 603
rect 516 597 524 603
rect 644 597 652 603
rect 676 597 1564 603
rect 1604 597 2060 603
rect 2180 597 2220 603
rect 3092 597 3500 603
rect 3764 597 3804 603
rect 3844 597 3852 603
rect 4020 597 4044 603
rect 4228 597 4236 603
rect 4372 597 4556 603
rect 4612 597 4620 603
rect 4804 597 4908 603
rect 4980 597 4988 603
rect 5172 597 5388 603
rect 5476 597 5500 603
rect 68 577 876 583
rect 996 577 1004 583
rect 1108 577 1116 583
rect 1364 577 1436 583
rect 1540 577 1548 583
rect 1572 577 1628 583
rect 2228 577 2300 583
rect 2356 577 2380 583
rect 2500 577 2524 583
rect 2564 577 2572 583
rect 2644 577 2652 583
rect 2708 577 2780 583
rect 2788 577 2956 583
rect 3108 577 3132 583
rect 3156 577 3164 583
rect 3188 577 3308 583
rect 3380 577 3452 583
rect 3556 577 3612 583
rect 3620 577 3788 583
rect 3796 577 4172 583
rect 4212 577 4220 583
rect 4356 577 4380 583
rect 4596 577 4604 583
rect 4644 577 4860 583
rect 4877 577 4892 583
rect 4877 564 4883 577
rect 5044 577 5164 583
rect 260 557 556 563
rect 596 557 956 563
rect 964 557 1164 563
rect 1172 557 1628 563
rect 1668 557 1676 563
rect 1732 557 1740 563
rect 1796 557 1836 563
rect 1860 557 1980 563
rect 2356 557 2620 563
rect 2644 557 2652 563
rect 2692 557 2748 563
rect 2900 557 2988 563
rect 2996 557 3228 563
rect 3268 557 3340 563
rect 3364 557 3436 563
rect 3460 557 3468 563
rect 3636 557 4012 563
rect 4372 557 4396 563
rect 4420 557 4444 563
rect 4596 557 4700 563
rect 4708 557 4732 563
rect 4900 557 5196 563
rect 5300 557 5308 563
rect 5373 563 5379 576
rect 5373 557 5388 563
rect 5396 557 5420 563
rect 2125 544 2131 556
rect 2813 544 2819 556
rect 132 537 252 543
rect 340 537 348 543
rect 436 537 716 543
rect 724 537 844 543
rect 1117 537 1132 543
rect 1284 537 1980 543
rect 2164 537 2812 543
rect 2884 537 2892 543
rect 2900 537 2908 543
rect 2964 537 3324 543
rect 3332 537 3484 543
rect 3508 537 3564 543
rect 3652 537 3660 543
rect 3684 537 4524 543
rect 4532 537 4652 543
rect 4692 537 4732 543
rect 4980 537 5084 543
rect 5156 537 5212 543
rect 5284 537 5299 543
rect 5332 537 5404 543
rect 532 517 540 523
rect 612 517 636 523
rect 804 517 844 523
rect 948 517 956 523
rect 964 517 1580 523
rect 1636 517 1660 523
rect 1700 517 1948 523
rect 1972 517 2620 523
rect 2644 517 2700 523
rect 2852 517 3036 523
rect 3076 517 3331 523
rect 20 497 108 503
rect 196 497 220 503
rect 228 497 236 503
rect 244 497 300 503
rect 1332 497 1932 503
rect 2013 497 2028 503
rect 2100 497 2124 503
rect 2148 497 2188 503
rect 2340 497 2348 503
rect 2612 497 2620 503
rect 2692 497 2860 503
rect 3012 497 3036 503
rect 3060 497 3292 503
rect 3300 497 3308 503
rect 3325 503 3331 517
rect 3396 517 3420 523
rect 3444 517 3868 523
rect 4068 517 4108 523
rect 4148 517 4716 523
rect 4724 517 5036 523
rect 5188 517 5260 523
rect 5332 517 5452 523
rect 3325 497 4252 503
rect 4276 497 4284 503
rect 4308 497 4316 503
rect 4340 497 4492 503
rect 4772 497 4812 503
rect 4916 497 5004 503
rect 5124 497 5164 503
rect 5268 497 5436 503
rect 292 477 364 483
rect 1220 477 1772 483
rect 1812 477 2460 483
rect 2516 477 2524 483
rect 2916 477 3116 483
rect 3140 477 3404 483
rect 3412 477 3532 483
rect 3540 477 3692 483
rect 3700 477 3740 483
rect 3748 477 3788 483
rect 4228 477 4412 483
rect 4420 477 4588 483
rect 5252 477 5468 483
rect 1412 457 1580 463
rect 2884 457 3100 463
rect 3268 457 3340 463
rect 3348 457 3452 463
rect 4148 457 4924 463
rect 5124 457 5436 463
rect 1508 437 1692 443
rect 2900 437 4124 443
rect 4132 437 4268 443
rect 5316 437 5436 443
rect 1700 417 1724 423
rect 1828 417 2444 423
rect 2468 417 3004 423
rect 3652 417 3916 423
rect 436 397 1084 403
rect 1092 397 2828 403
rect 2980 397 2988 403
rect 4228 397 4332 403
rect 4340 397 4732 403
rect 1540 377 1548 383
rect 2420 377 2652 383
rect 2660 377 2700 383
rect 3060 377 3068 383
rect 3508 377 3516 383
rect 3581 377 3596 383
rect 3908 377 3916 383
rect 4228 377 4284 383
rect 4356 377 4364 383
rect 4468 377 4476 383
rect 4804 377 4940 383
rect 5140 377 5164 383
rect 5220 377 5564 383
rect 388 357 396 363
rect 788 357 1292 363
rect 1540 357 1548 363
rect 1844 357 1852 363
rect 2132 357 2508 363
rect 2548 357 2556 363
rect 2564 357 2812 363
rect 3908 357 4236 363
rect 4356 357 4364 363
rect 4772 357 5372 363
rect 100 337 460 343
rect 573 343 579 356
rect 717 344 723 356
rect 573 337 588 343
rect 1156 337 1196 343
rect 1492 337 1772 343
rect 2052 337 2412 343
rect 2420 337 2540 343
rect 2596 337 2684 343
rect 3252 337 3260 343
rect 4372 337 4460 343
rect 4900 337 4972 343
rect 5044 337 5388 343
rect 2749 324 2755 336
rect 36 317 140 323
rect 500 317 508 323
rect 564 317 1020 323
rect 1076 317 1148 323
rect 1156 317 1212 323
rect 1268 317 1356 323
rect 1380 317 1388 323
rect 1412 317 1900 323
rect 1908 317 2204 323
rect 2212 317 2220 323
rect 2276 317 2284 323
rect 2468 317 2476 323
rect 2516 317 2620 323
rect 2852 317 2860 323
rect 3140 317 3356 323
rect 3364 317 3788 323
rect 3844 317 3852 323
rect 3924 317 3932 323
rect 3972 317 4492 323
rect 4644 317 4684 323
rect 4852 317 5228 323
rect 5284 317 5292 323
rect 5316 317 5324 323
rect 5364 317 5635 323
rect 180 297 988 303
rect 1028 297 1916 303
rect 1924 297 2028 303
rect 2244 297 2316 303
rect 2836 297 3164 303
rect 3172 297 3436 303
rect 3844 297 3964 303
rect 4100 297 4156 303
rect 4180 297 4284 303
rect 4292 297 4380 303
rect 4404 297 4476 303
rect 4500 297 4508 303
rect 4580 297 4812 303
rect 4932 297 5020 303
rect 5044 297 5164 303
rect 5300 297 5308 303
rect 2045 284 2051 296
rect 68 277 76 283
rect 212 277 220 283
rect 260 277 300 283
rect 324 277 476 283
rect 580 277 588 283
rect 628 277 684 283
rect 708 277 764 283
rect 804 277 819 283
rect 836 277 876 283
rect 900 277 1100 283
rect 1140 277 1164 283
rect 1220 277 1228 283
rect 1284 277 1404 283
rect 1412 277 1788 283
rect 1796 277 1804 283
rect 1924 277 1932 283
rect 2125 283 2131 296
rect 2116 277 2131 283
rect 2244 277 2252 283
rect 2436 277 2444 283
rect 2500 277 2572 283
rect 2708 277 2748 283
rect 2900 277 2908 283
rect 3076 277 3548 283
rect 3604 277 3996 283
rect 4052 277 4108 283
rect 4148 277 4204 283
rect 4276 277 4300 283
rect 4356 277 4412 283
rect 4660 277 5324 283
rect 5332 277 5340 283
rect 5348 277 5356 283
rect 20 257 44 263
rect 52 257 732 263
rect 740 257 1404 263
rect 1476 257 1516 263
rect 1556 257 1612 263
rect 1636 257 1644 263
rect 1860 257 2108 263
rect 2116 257 2636 263
rect 2660 257 2876 263
rect 2884 257 2908 263
rect 2980 257 3084 263
rect 3204 257 3244 263
rect 3268 257 3420 263
rect 3428 257 3676 263
rect 3684 257 4012 263
rect 4020 257 4044 263
rect 4052 257 4860 263
rect 4932 257 5180 263
rect 5252 257 5500 263
rect 132 237 204 243
rect 404 237 444 243
rect 468 237 924 243
rect 964 237 972 243
rect 1220 237 1420 243
rect 1492 237 1500 243
rect 1604 237 1676 243
rect 1716 237 1740 243
rect 2180 237 2316 243
rect 2372 237 2572 243
rect 2868 237 2876 243
rect 2900 237 3020 243
rect 3076 237 3132 243
rect 3156 237 3292 243
rect 3300 237 3468 243
rect 3572 237 3788 243
rect 3796 237 4188 243
rect 4196 237 4236 243
rect 4260 237 5116 243
rect 5124 237 5436 243
rect 5444 237 5452 243
rect 708 217 748 223
rect 1028 217 1036 223
rect 1060 217 1292 223
rect 1764 217 1804 223
rect 3396 217 3612 223
rect 3636 217 3660 223
rect 4116 217 4604 223
rect 4740 217 4764 223
rect 4804 217 4828 223
rect 4932 217 4940 223
rect 5076 217 5084 223
rect 5124 217 5180 223
rect 5204 217 5228 223
rect 5252 217 5635 223
rect 324 197 332 203
rect 356 197 524 203
rect 564 197 748 203
rect 1284 197 1452 203
rect 1796 197 1820 203
rect 1860 197 1980 203
rect 2292 197 2300 203
rect 2964 197 2972 203
rect 3156 197 3180 203
rect 3460 197 3468 203
rect 3780 197 4092 203
rect 4100 197 4780 203
rect 5060 197 5148 203
rect 5188 197 5244 203
rect 5444 197 5468 203
rect 13 177 28 183
rect 260 177 428 183
rect 580 177 604 183
rect 708 177 716 183
rect 852 177 2188 183
rect 2308 177 2364 183
rect 2436 177 2460 183
rect 2564 177 2572 183
rect 2628 177 2796 183
rect 2948 177 3020 183
rect 3028 177 3100 183
rect 3332 177 3596 183
rect 3668 177 3692 183
rect 3780 177 3788 183
rect 3812 177 3900 183
rect 3972 177 4092 183
rect 4164 177 4172 183
rect 4516 177 4668 183
rect 4692 177 4748 183
rect 5140 177 5196 183
rect 5252 177 5260 183
rect 5316 177 5356 183
rect 5588 177 5635 183
rect 61 164 67 176
rect 77 164 83 176
rect 4221 164 4227 176
rect 292 157 316 163
rect 372 157 844 163
rect 868 157 876 163
rect 1028 157 1068 163
rect 1092 157 1100 163
rect 1108 157 2492 163
rect 2612 157 2828 163
rect 2836 157 2956 163
rect 3012 157 3084 163
rect 3092 157 3244 163
rect 3332 157 3404 163
rect 3460 157 3948 163
rect 3988 157 3996 163
rect 4052 157 4140 163
rect 4260 157 4716 163
rect 4724 157 4908 163
rect 4996 157 5036 163
rect 5172 157 5292 163
rect 5332 157 5340 163
rect 237 144 243 156
rect 52 137 92 143
rect 132 137 220 143
rect 244 137 908 143
rect 980 137 988 143
rect 1028 137 1100 143
rect 1117 137 1132 143
rect 1156 137 1164 143
rect 1188 137 1196 143
rect 1236 137 1251 143
rect 1332 137 1724 143
rect 1748 137 1756 143
rect 1780 137 1884 143
rect 1892 137 1932 143
rect 1956 137 2124 143
rect 2180 137 2220 143
rect 2244 137 2636 143
rect 2644 137 2652 143
rect 2692 137 2748 143
rect 2788 137 2812 143
rect 2820 137 2828 143
rect 2852 137 3452 143
rect 3476 137 3484 143
rect 3540 137 3596 143
rect 3620 137 4204 143
rect 4340 137 4444 143
rect 4452 137 4460 143
rect 4468 137 4972 143
rect 5012 137 5260 143
rect 5444 137 5459 143
rect 100 117 140 123
rect 196 117 364 123
rect 420 117 428 123
rect 452 117 556 123
rect 580 117 588 123
rect 612 117 652 123
rect 708 117 732 123
rect 804 117 812 123
rect 996 117 2428 123
rect 2436 117 2540 123
rect 2564 117 2668 123
rect 2676 117 2876 123
rect 2948 117 3276 123
rect 3300 117 3340 123
rect 3412 117 4332 123
rect 4365 117 4380 123
rect 4676 117 4684 123
rect 4708 117 4748 123
rect 4772 117 4812 123
rect 4852 117 4940 123
rect 5028 117 5516 123
rect 4541 104 4547 116
rect 532 97 556 103
rect 932 97 972 103
rect 1076 97 1148 103
rect 1172 97 1292 103
rect 1348 97 1356 103
rect 1428 97 1548 103
rect 1588 97 1596 103
rect 1620 97 1676 103
rect 1732 97 1836 103
rect 1844 97 2060 103
rect 2116 97 2124 103
rect 2228 97 2332 103
rect 2356 97 2380 103
rect 2756 97 2892 103
rect 3124 97 3132 103
rect 3140 97 3980 103
rect 4036 97 4092 103
rect 4116 97 4172 103
rect 4292 97 4300 103
rect 4324 97 4364 103
rect 4420 97 4524 103
rect 4564 97 4652 103
rect 4788 97 5404 103
rect 637 84 643 96
rect 1716 77 1756 83
rect 1924 77 1948 83
rect 2180 77 2476 83
rect 3460 77 3564 83
rect 3652 77 3692 83
rect 3844 77 3884 83
rect 4004 77 5276 83
rect 5332 77 5468 83
rect 1805 64 1811 76
rect 1716 57 1724 63
rect 4628 57 5420 63
rect 1741 44 1747 56
rect 2253 44 2259 56
rect 3853 44 3859 56
rect 2692 37 2716 43
rect 2724 37 2908 43
rect 2916 37 2972 43
rect 2980 37 3036 43
rect 4564 37 4652 43
rect 2948 17 2956 23
rect 4692 17 4700 23
<< m4contact >>
rect 252 3956 260 3964
rect 1484 3956 1492 3964
rect 2684 3956 2692 3964
rect 3948 3936 3956 3944
rect 1916 3916 1924 3924
rect 2332 3916 2340 3924
rect 2492 3916 2500 3924
rect 3260 3916 3268 3924
rect 3788 3916 3796 3924
rect 3820 3916 3828 3924
rect 4524 3916 4532 3924
rect 4700 3916 4708 3924
rect 5468 3916 5476 3924
rect 252 3896 260 3904
rect 1068 3896 1076 3904
rect 1308 3896 1316 3904
rect 2380 3896 2388 3904
rect 3164 3896 3172 3904
rect 3644 3896 3652 3904
rect 3740 3896 3748 3904
rect 5324 3896 5332 3904
rect 764 3876 772 3884
rect 812 3876 820 3884
rect 844 3876 852 3884
rect 1212 3876 1220 3884
rect 1404 3876 1412 3884
rect 2092 3876 2100 3884
rect 2412 3876 2420 3884
rect 2492 3876 2500 3884
rect 2860 3876 2868 3884
rect 3804 3876 3812 3884
rect 3868 3876 3876 3884
rect 5212 3876 5220 3884
rect 5292 3876 5300 3884
rect 5356 3876 5364 3884
rect 972 3856 980 3864
rect 2188 3856 2196 3864
rect 2300 3856 2308 3864
rect 2748 3856 2756 3864
rect 2796 3856 2804 3864
rect 3020 3856 3028 3864
rect 3500 3856 3508 3864
rect 412 3836 420 3844
rect 428 3836 436 3844
rect 700 3836 708 3844
rect 748 3836 756 3844
rect 2796 3836 2804 3844
rect 3564 3836 3572 3844
rect 4748 3856 4756 3864
rect 5132 3856 5140 3864
rect 4476 3836 4484 3844
rect 5308 3836 5316 3844
rect 2028 3816 2036 3824
rect 3788 3816 3796 3824
rect 3900 3816 3908 3824
rect 4124 3816 4132 3824
rect 4540 3816 4548 3824
rect 5244 3816 5252 3824
rect 780 3796 788 3804
rect 956 3796 964 3804
rect 1084 3796 1092 3804
rect 1468 3796 1476 3804
rect 1500 3796 1508 3804
rect 1564 3796 1572 3804
rect 1612 3796 1620 3804
rect 1660 3796 1668 3804
rect 2588 3796 2596 3804
rect 2620 3796 2628 3804
rect 2956 3796 2964 3804
rect 3212 3796 3220 3804
rect 3244 3796 3252 3804
rect 3788 3796 3796 3804
rect 4044 3796 4052 3804
rect 4076 3796 4084 3804
rect 4108 3796 4116 3804
rect 4236 3796 4244 3804
rect 4684 3796 4692 3804
rect 5068 3796 5076 3804
rect 5308 3796 5316 3804
rect 5420 3796 5428 3804
rect 524 3776 532 3784
rect 828 3776 836 3784
rect 1932 3776 1940 3784
rect 2188 3776 2196 3784
rect 3068 3776 3076 3784
rect 4172 3776 4180 3784
rect 5340 3776 5348 3784
rect 5436 3776 5444 3784
rect 76 3756 84 3764
rect 252 3756 260 3764
rect 892 3756 900 3764
rect 1020 3756 1028 3764
rect 1676 3756 1684 3764
rect 2588 3756 2596 3764
rect 2908 3756 2916 3764
rect 2956 3756 2964 3764
rect 3036 3756 3044 3764
rect 3340 3756 3348 3764
rect 3356 3756 3364 3764
rect 3388 3756 3396 3764
rect 3596 3756 3604 3764
rect 3628 3756 3636 3764
rect 3740 3756 3748 3764
rect 4444 3756 4452 3764
rect 4716 3756 4724 3764
rect 4732 3756 4740 3764
rect 4764 3756 4772 3764
rect 5180 3756 5188 3764
rect 5516 3756 5524 3764
rect 12 3736 20 3744
rect 476 3736 484 3744
rect 508 3736 516 3744
rect 1084 3736 1092 3744
rect 1292 3736 1300 3744
rect 1340 3736 1348 3744
rect 2316 3736 2324 3744
rect 2348 3736 2356 3744
rect 2924 3736 2932 3744
rect 3852 3736 3860 3744
rect 3868 3736 3876 3744
rect 3932 3736 3940 3744
rect 3948 3736 3956 3744
rect 4300 3736 4308 3744
rect 4332 3736 4340 3744
rect 5180 3736 5188 3744
rect 5244 3736 5252 3744
rect 5340 3736 5348 3744
rect 540 3716 548 3724
rect 636 3716 644 3724
rect 716 3716 724 3724
rect 908 3716 916 3724
rect 956 3716 964 3724
rect 2796 3716 2804 3724
rect 4140 3716 4148 3724
rect 4812 3716 4820 3724
rect 5196 3716 5204 3724
rect 76 3696 84 3704
rect 300 3696 308 3704
rect 524 3696 532 3704
rect 812 3696 820 3704
rect 860 3696 868 3704
rect 1212 3696 1220 3704
rect 1372 3696 1380 3704
rect 1452 3696 1460 3704
rect 1484 3696 1492 3704
rect 1516 3696 1524 3704
rect 1836 3696 1844 3704
rect 1916 3696 1924 3704
rect 2284 3696 2292 3704
rect 2332 3696 2340 3704
rect 2908 3696 2916 3704
rect 3004 3696 3012 3704
rect 3772 3696 3780 3704
rect 3804 3696 3812 3704
rect 4268 3696 4276 3704
rect 4364 3696 4372 3704
rect 4380 3696 4388 3704
rect 4764 3696 4772 3704
rect 4924 3696 4932 3704
rect 284 3676 292 3684
rect 828 3676 836 3684
rect 1180 3676 1188 3684
rect 1244 3676 1252 3684
rect 3324 3676 3332 3684
rect 3964 3676 3972 3684
rect 1324 3656 1332 3664
rect 2188 3656 2196 3664
rect 2028 3636 2036 3644
rect 2684 3636 2692 3644
rect 3132 3636 3140 3644
rect 3228 3636 3236 3644
rect 4364 3636 4372 3644
rect 1196 3616 1204 3624
rect 5276 3616 5284 3624
rect 1964 3596 1972 3604
rect 2124 3596 2132 3604
rect 3020 3596 3028 3604
rect 1980 3576 1988 3584
rect 2620 3576 2628 3584
rect 3196 3576 3204 3584
rect 4156 3576 4164 3584
rect 2156 3556 2164 3564
rect 2956 3556 2964 3564
rect 476 3536 484 3544
rect 764 3536 772 3544
rect 812 3536 820 3544
rect 1692 3536 1700 3544
rect 3100 3536 3108 3544
rect 3212 3536 3220 3544
rect 3292 3536 3300 3544
rect 3484 3536 3492 3544
rect 4012 3536 4020 3544
rect 5068 3536 5076 3544
rect 5452 3536 5460 3544
rect 812 3516 820 3524
rect 828 3516 836 3524
rect 1388 3516 1396 3524
rect 2268 3516 2276 3524
rect 2844 3516 2852 3524
rect 3004 3516 3012 3524
rect 4012 3516 4020 3524
rect 4044 3516 4052 3524
rect 4092 3516 4100 3524
rect 4284 3516 4292 3524
rect 4460 3516 4468 3524
rect 4508 3516 4516 3524
rect 396 3496 404 3504
rect 588 3496 596 3504
rect 908 3496 916 3504
rect 1676 3496 1684 3504
rect 1788 3496 1796 3504
rect 1820 3496 1828 3504
rect 2076 3496 2084 3504
rect 2380 3496 2388 3504
rect 3212 3496 3220 3504
rect 4028 3496 4036 3504
rect 188 3476 196 3484
rect 204 3476 212 3484
rect 1340 3476 1348 3484
rect 3820 3476 3828 3484
rect 4988 3476 4996 3484
rect 5164 3476 5172 3484
rect 5260 3476 5268 3484
rect 956 3456 964 3464
rect 2140 3456 2148 3464
rect 2268 3456 2276 3464
rect 2300 3456 2308 3464
rect 2924 3456 2932 3464
rect 2940 3456 2948 3464
rect 3020 3456 3028 3464
rect 3196 3456 3204 3464
rect 3228 3456 3236 3464
rect 3836 3456 3844 3464
rect 3916 3456 3924 3464
rect 4092 3456 4100 3464
rect 4188 3456 4196 3464
rect 4844 3456 4852 3464
rect 4908 3456 4916 3464
rect 4940 3456 4948 3464
rect 5020 3456 5028 3464
rect 876 3436 884 3444
rect 956 3436 964 3444
rect 1004 3436 1012 3444
rect 1708 3436 1716 3444
rect 1932 3436 1940 3444
rect 4268 3436 4276 3444
rect 4316 3436 4324 3444
rect 1036 3416 1044 3424
rect 1276 3416 1284 3424
rect 2476 3416 2484 3424
rect 3100 3416 3108 3424
rect 3292 3416 3300 3424
rect 3356 3416 3364 3424
rect 1004 3396 1012 3404
rect 1020 3396 1028 3404
rect 140 3376 148 3384
rect 316 3376 324 3384
rect 364 3376 372 3384
rect 636 3376 644 3384
rect 1052 3376 1060 3384
rect 1292 3396 1300 3404
rect 1612 3396 1620 3404
rect 1740 3396 1748 3404
rect 1804 3396 1812 3404
rect 1916 3396 1924 3404
rect 1980 3396 1988 3404
rect 2108 3396 2116 3404
rect 2236 3396 2244 3404
rect 2268 3396 2276 3404
rect 3980 3416 3988 3424
rect 4044 3416 4052 3424
rect 3500 3396 3508 3404
rect 4652 3416 4660 3424
rect 4668 3416 4676 3424
rect 4956 3416 4964 3424
rect 5084 3416 5092 3424
rect 4076 3396 4084 3404
rect 4156 3396 4164 3404
rect 4284 3396 4292 3404
rect 4364 3396 4372 3404
rect 4444 3396 4452 3404
rect 4668 3396 4676 3404
rect 4780 3396 4788 3404
rect 5020 3396 5028 3404
rect 5132 3396 5140 3404
rect 1420 3376 1428 3384
rect 2092 3376 2100 3384
rect 2156 3376 2164 3384
rect 2268 3376 2276 3384
rect 2636 3376 2644 3384
rect 3468 3376 3476 3384
rect 3724 3376 3732 3384
rect 3852 3376 3860 3384
rect 4764 3376 4772 3384
rect 5116 3376 5124 3384
rect 5180 3376 5188 3384
rect 5484 3376 5492 3384
rect 204 3356 212 3364
rect 764 3356 772 3364
rect 1484 3356 1492 3364
rect 1564 3356 1572 3364
rect 2572 3356 2580 3364
rect 2604 3356 2612 3364
rect 2940 3356 2948 3364
rect 3100 3356 3108 3364
rect 3388 3356 3396 3364
rect 3580 3356 3588 3364
rect 3660 3356 3668 3364
rect 3692 3356 3700 3364
rect 5132 3356 5140 3364
rect 60 3336 68 3344
rect 380 3336 388 3344
rect 652 3336 660 3344
rect 1564 3336 1572 3344
rect 2316 3336 2324 3344
rect 2620 3336 2628 3344
rect 2668 3336 2676 3344
rect 2700 3336 2708 3344
rect 2716 3336 2724 3344
rect 2812 3336 2820 3344
rect 2908 3336 2916 3344
rect 3004 3336 3012 3344
rect 3324 3336 3332 3344
rect 3500 3336 3508 3344
rect 3580 3336 3588 3344
rect 3612 3336 3620 3344
rect 4444 3336 4452 3344
rect 4492 3336 4500 3344
rect 4636 3336 4644 3344
rect 4684 3336 4692 3344
rect 4796 3336 4804 3344
rect 5196 3336 5204 3344
rect 188 3316 196 3324
rect 940 3316 948 3324
rect 1020 3316 1028 3324
rect 1036 3316 1044 3324
rect 1260 3316 1268 3324
rect 1740 3316 1748 3324
rect 1756 3316 1764 3324
rect 1964 3316 1972 3324
rect 2604 3316 2612 3324
rect 3420 3316 3428 3324
rect 3852 3316 3860 3324
rect 300 3296 308 3304
rect 876 3296 884 3304
rect 908 3296 916 3304
rect 1532 3296 1540 3304
rect 1724 3296 1732 3304
rect 3244 3296 3252 3304
rect 4924 3316 4932 3324
rect 4940 3316 4948 3324
rect 5196 3316 5204 3324
rect 4060 3296 4068 3304
rect 4076 3296 4084 3304
rect 4204 3296 4212 3304
rect 4892 3296 4900 3304
rect 1884 3276 1892 3284
rect 2844 3276 2852 3284
rect 3436 3276 3444 3284
rect 4492 3276 4500 3284
rect 4860 3276 4868 3284
rect 412 3256 420 3264
rect 604 3256 612 3264
rect 940 3256 948 3264
rect 1084 3236 1092 3244
rect 2844 3256 2852 3264
rect 2860 3256 2868 3264
rect 3276 3256 3284 3264
rect 3884 3256 3892 3264
rect 4124 3256 4132 3264
rect 4732 3256 4740 3264
rect 1948 3236 1956 3244
rect 3644 3236 3652 3244
rect 1596 3216 1604 3224
rect 2332 3216 2340 3224
rect 3804 3216 3812 3224
rect 4572 3216 4580 3224
rect 76 3196 84 3204
rect 1084 3196 1092 3204
rect 1548 3196 1556 3204
rect 1708 3196 1716 3204
rect 2012 3196 2020 3204
rect 3084 3196 3092 3204
rect 3676 3196 3684 3204
rect 4044 3196 4052 3204
rect 4156 3196 4164 3204
rect 1724 3176 1732 3184
rect 1996 3176 2004 3184
rect 3324 3176 3332 3184
rect 3468 3176 3476 3184
rect 3756 3176 3764 3184
rect 3804 3176 3812 3184
rect 636 3156 644 3164
rect 828 3156 836 3164
rect 1916 3156 1924 3164
rect 2908 3156 2916 3164
rect 3612 3156 3620 3164
rect 4284 3156 4292 3164
rect 4316 3156 4324 3164
rect 4364 3156 4372 3164
rect 4588 3156 4596 3164
rect 396 3136 404 3144
rect 620 3136 628 3144
rect 940 3136 948 3144
rect 1228 3136 1236 3144
rect 1260 3136 1268 3144
rect 1324 3136 1332 3144
rect 1356 3136 1364 3144
rect 1484 3136 1492 3144
rect 3804 3136 3812 3144
rect 4044 3136 4052 3144
rect 4892 3136 4900 3144
rect 172 3116 180 3124
rect 540 3116 548 3124
rect 796 3116 804 3124
rect 860 3116 868 3124
rect 1452 3116 1460 3124
rect 1564 3116 1572 3124
rect 1644 3116 1652 3124
rect 1788 3116 1796 3124
rect 2476 3116 2484 3124
rect 3100 3116 3108 3124
rect 3324 3116 3332 3124
rect 3356 3116 3364 3124
rect 124 3096 132 3104
rect 236 3096 244 3104
rect 364 3096 372 3104
rect 508 3096 516 3104
rect 1036 3096 1044 3104
rect 1116 3096 1124 3104
rect 1196 3096 1204 3104
rect 1212 3096 1220 3104
rect 1468 3096 1476 3104
rect 1660 3096 1668 3104
rect 1852 3096 1860 3104
rect 2236 3096 2244 3104
rect 2380 3096 2388 3104
rect 2732 3096 2740 3104
rect 2812 3096 2820 3104
rect 3260 3096 3268 3104
rect 3500 3096 3508 3104
rect 3548 3096 3556 3104
rect 3900 3096 3908 3104
rect 4348 3116 4356 3124
rect 4412 3116 4420 3124
rect 4668 3116 4676 3124
rect 4716 3116 4724 3124
rect 4972 3116 4980 3124
rect 5020 3116 5028 3124
rect 4332 3096 4340 3104
rect 92 3076 100 3084
rect 4876 3096 4884 3104
rect 4924 3096 4932 3104
rect 5052 3116 5060 3124
rect 5388 3116 5396 3124
rect 5660 3116 5668 3124
rect 5132 3096 5140 3104
rect 5244 3096 5252 3104
rect 1596 3076 1604 3084
rect 1628 3076 1636 3084
rect 1820 3076 1828 3084
rect 1836 3076 1844 3084
rect 2396 3076 2404 3084
rect 3900 3076 3908 3084
rect 172 3056 180 3064
rect 204 3056 212 3064
rect 252 3056 260 3064
rect 300 3056 308 3064
rect 348 3056 356 3064
rect 444 3056 452 3064
rect 1148 3056 1156 3064
rect 1292 3056 1300 3064
rect 1852 3056 1860 3064
rect 2028 3056 2036 3064
rect 2060 3056 2068 3064
rect 2220 3056 2228 3064
rect 3308 3056 3316 3064
rect 3356 3056 3364 3064
rect 3388 3056 3396 3064
rect 3692 3056 3700 3064
rect 3708 3056 3716 3064
rect 3788 3056 3796 3064
rect 4828 3076 4836 3084
rect 4908 3076 4916 3084
rect 5100 3076 5108 3084
rect 5516 3076 5524 3084
rect 4316 3056 4324 3064
rect 4412 3056 4420 3064
rect 4428 3056 4436 3064
rect 5260 3056 5268 3064
rect 332 3036 340 3044
rect 636 3036 644 3044
rect 764 3036 772 3044
rect 1212 3036 1220 3044
rect 1580 3036 1588 3044
rect 1772 3036 1780 3044
rect 3356 3036 3364 3044
rect 3516 3036 3524 3044
rect 3852 3036 3860 3044
rect 4060 3036 4068 3044
rect 4940 3036 4948 3044
rect 5052 3036 5060 3044
rect 5084 3036 5092 3044
rect 572 3016 580 3024
rect 1164 3016 1172 3024
rect 1036 2996 1044 3004
rect 1068 2996 1076 3004
rect 1228 2996 1236 3004
rect 3660 3016 3668 3024
rect 3852 3016 3860 3024
rect 4556 3016 4564 3024
rect 1868 2996 1876 3004
rect 3212 2996 3220 3004
rect 3244 2996 3252 3004
rect 3340 2996 3348 3004
rect 3612 2996 3620 3004
rect 3980 2996 3988 3004
rect 5228 2996 5236 3004
rect 5372 2996 5380 3004
rect 5660 2996 5668 3004
rect 108 2976 116 2984
rect 828 2976 836 2984
rect 1116 2976 1124 2984
rect 1308 2976 1316 2984
rect 1516 2976 1524 2984
rect 1644 2976 1652 2984
rect 1900 2976 1908 2984
rect 2108 2976 2116 2984
rect 28 2956 36 2964
rect 588 2956 596 2964
rect 764 2956 772 2964
rect 1244 2956 1252 2964
rect 1276 2956 1284 2964
rect 1308 2956 1316 2964
rect 1596 2956 1604 2964
rect 2300 2956 2308 2964
rect 2732 2976 2740 2984
rect 2812 2976 2820 2984
rect 3468 2976 3476 2984
rect 3484 2976 3492 2984
rect 3564 2976 3572 2984
rect 4732 2976 4740 2984
rect 4828 2976 4836 2984
rect 2892 2956 2900 2964
rect 3020 2956 3028 2964
rect 3084 2956 3092 2964
rect 3548 2956 3556 2964
rect 3708 2956 3716 2964
rect 3772 2956 3780 2964
rect 4156 2956 4164 2964
rect 4316 2956 4324 2964
rect 4876 2956 4884 2964
rect 4924 2956 4932 2964
rect 4988 2956 4996 2964
rect 5004 2956 5012 2964
rect 5164 2956 5172 2964
rect 5452 2956 5460 2964
rect 284 2936 292 2944
rect 540 2936 548 2944
rect 748 2936 756 2944
rect 924 2936 932 2944
rect 972 2936 980 2944
rect 1196 2936 1204 2944
rect 1244 2936 1252 2944
rect 1804 2936 1812 2944
rect 2124 2936 2132 2944
rect 2284 2936 2292 2944
rect 2348 2936 2356 2944
rect 2684 2936 2692 2944
rect 3884 2936 3892 2944
rect 4028 2936 4036 2944
rect 4636 2936 4644 2944
rect 4780 2936 4788 2944
rect 4844 2936 4852 2944
rect 5068 2936 5076 2944
rect 5244 2936 5252 2944
rect 1004 2916 1012 2924
rect 1308 2916 1316 2924
rect 1708 2916 1716 2924
rect 3004 2916 3012 2924
rect 3148 2916 3156 2924
rect 3484 2916 3492 2924
rect 12 2896 20 2904
rect 252 2896 260 2904
rect 444 2896 452 2904
rect 1084 2896 1092 2904
rect 1292 2896 1300 2904
rect 1932 2896 1940 2904
rect 380 2876 388 2884
rect 444 2876 452 2884
rect 620 2876 628 2884
rect 1148 2876 1156 2884
rect 2748 2896 2756 2904
rect 3180 2896 3188 2904
rect 3244 2896 3252 2904
rect 3308 2896 3316 2904
rect 3436 2896 3444 2904
rect 3452 2896 3460 2904
rect 3532 2896 3540 2904
rect 3692 2916 3700 2924
rect 3740 2916 3748 2924
rect 3852 2916 3860 2924
rect 3932 2916 3940 2924
rect 4204 2916 4212 2924
rect 4332 2916 4340 2924
rect 4412 2916 4420 2924
rect 4508 2916 4516 2924
rect 4748 2916 4756 2924
rect 4828 2916 4836 2924
rect 4860 2916 4868 2924
rect 5052 2916 5060 2924
rect 4252 2896 4260 2904
rect 4268 2896 4276 2904
rect 5116 2896 5124 2904
rect 5404 2896 5412 2904
rect 3196 2876 3204 2884
rect 3372 2876 3380 2884
rect 3916 2876 3924 2884
rect 4780 2876 4788 2884
rect 4860 2876 4868 2884
rect 4924 2876 4932 2884
rect 3340 2856 3348 2864
rect 3404 2856 3412 2864
rect 2284 2836 2292 2844
rect 3740 2836 3748 2844
rect 3004 2816 3012 2824
rect 3340 2816 3348 2824
rect 3404 2816 3412 2824
rect 780 2796 788 2804
rect 860 2796 868 2804
rect 1196 2796 1204 2804
rect 1804 2796 1812 2804
rect 2044 2796 2052 2804
rect 2380 2796 2388 2804
rect 2604 2796 2612 2804
rect 3868 2796 3876 2804
rect 1548 2776 1556 2784
rect 3068 2776 3076 2784
rect 5372 2776 5380 2784
rect 636 2756 644 2764
rect 1196 2756 1204 2764
rect 1628 2756 1636 2764
rect 1852 2756 1860 2764
rect 1916 2756 1924 2764
rect 2668 2756 2676 2764
rect 3132 2756 3140 2764
rect 3468 2756 3476 2764
rect 844 2736 852 2744
rect 924 2736 932 2744
rect 1020 2736 1028 2744
rect 1788 2736 1796 2744
rect 2572 2736 2580 2744
rect 3148 2736 3156 2744
rect 4204 2756 4212 2764
rect 4060 2736 4068 2744
rect 4284 2736 4292 2744
rect 4316 2736 4324 2744
rect 4668 2736 4676 2744
rect 5484 2736 5492 2744
rect 268 2716 276 2724
rect 652 2716 660 2724
rect 1452 2716 1460 2724
rect 1788 2716 1796 2724
rect 2252 2716 2260 2724
rect 2444 2716 2452 2724
rect 2460 2716 2468 2724
rect 3340 2716 3348 2724
rect 3772 2716 3780 2724
rect 3804 2716 3812 2724
rect 4524 2716 4532 2724
rect 4812 2716 4820 2724
rect 4908 2716 4916 2724
rect 4972 2716 4980 2724
rect 5020 2716 5028 2724
rect 556 2696 564 2704
rect 572 2696 580 2704
rect 604 2696 612 2704
rect 780 2696 788 2704
rect 908 2696 916 2704
rect 1100 2696 1108 2704
rect 1260 2696 1268 2704
rect 1404 2696 1412 2704
rect 1452 2696 1460 2704
rect 1916 2696 1924 2704
rect 1948 2696 1956 2704
rect 2028 2696 2036 2704
rect 2044 2696 2052 2704
rect 2780 2696 2788 2704
rect 3004 2696 3012 2704
rect 3196 2696 3204 2704
rect 3516 2696 3524 2704
rect 3612 2696 3620 2704
rect 3740 2696 3748 2704
rect 3756 2696 3764 2704
rect 3836 2696 3844 2704
rect 4060 2696 4068 2704
rect 4380 2696 4388 2704
rect 4652 2696 4660 2704
rect 5484 2696 5492 2704
rect 28 2676 36 2684
rect 140 2676 148 2684
rect 588 2676 596 2684
rect 652 2676 660 2684
rect 684 2676 692 2684
rect 732 2676 740 2684
rect 1004 2676 1012 2684
rect 1324 2676 1332 2684
rect 1340 2676 1348 2684
rect 1468 2676 1476 2684
rect 1516 2676 1524 2684
rect 1548 2676 1556 2684
rect 1596 2676 1604 2684
rect 1644 2676 1652 2684
rect 1980 2676 1988 2684
rect 2172 2676 2180 2684
rect 2236 2676 2244 2684
rect 2364 2676 2372 2684
rect 2556 2676 2564 2684
rect 2620 2676 2628 2684
rect 2652 2676 2660 2684
rect 3004 2676 3012 2684
rect 3212 2676 3220 2684
rect 3292 2676 3300 2684
rect 3420 2676 3428 2684
rect 3516 2676 3524 2684
rect 3740 2676 3748 2684
rect 4220 2676 4228 2684
rect 4412 2676 4420 2684
rect 4444 2676 4452 2684
rect 4748 2676 4756 2684
rect 5148 2676 5156 2684
rect 5372 2676 5380 2684
rect 5516 2676 5524 2684
rect 508 2656 516 2664
rect 524 2656 532 2664
rect 844 2656 852 2664
rect 860 2656 868 2664
rect 1068 2656 1076 2664
rect 1244 2656 1252 2664
rect 1260 2656 1268 2664
rect 1932 2656 1940 2664
rect 1948 2656 1956 2664
rect 1996 2656 2004 2664
rect 2124 2656 2132 2664
rect 2204 2656 2212 2664
rect 3612 2656 3620 2664
rect 3660 2656 3668 2664
rect 3708 2656 3716 2664
rect 3884 2656 3892 2664
rect 4044 2656 4052 2664
rect 4188 2656 4196 2664
rect 4236 2656 4244 2664
rect 4476 2656 4484 2664
rect 4700 2656 4708 2664
rect 4764 2656 4772 2664
rect 4924 2656 4932 2664
rect 252 2636 260 2644
rect 540 2636 548 2644
rect 924 2636 932 2644
rect 1004 2636 1012 2644
rect 1052 2636 1060 2644
rect 1260 2636 1268 2644
rect 1324 2636 1332 2644
rect 1340 2636 1348 2644
rect 1436 2636 1444 2644
rect 1916 2636 1924 2644
rect 1964 2636 1972 2644
rect 2124 2636 2132 2644
rect 3052 2636 3060 2644
rect 3292 2636 3300 2644
rect 3580 2636 3588 2644
rect 4124 2636 4132 2644
rect 4524 2636 4532 2644
rect 4684 2636 4692 2644
rect 268 2616 276 2624
rect 380 2616 388 2624
rect 3596 2616 3604 2624
rect 3772 2616 3780 2624
rect 3804 2616 3812 2624
rect 4860 2616 4868 2624
rect 5052 2616 5060 2624
rect 204 2596 212 2604
rect 508 2596 516 2604
rect 4076 2596 4084 2604
rect 4620 2596 4628 2604
rect 108 2576 116 2584
rect 316 2576 324 2584
rect 540 2576 548 2584
rect 828 2576 836 2584
rect 76 2556 84 2564
rect 348 2556 356 2564
rect 396 2556 404 2564
rect 460 2556 468 2564
rect 492 2556 500 2564
rect 668 2556 676 2564
rect 780 2556 788 2564
rect 1212 2576 1220 2584
rect 1372 2576 1380 2584
rect 2012 2576 2020 2584
rect 2028 2576 2036 2584
rect 2268 2576 2276 2584
rect 3340 2576 3348 2584
rect 3516 2576 3524 2584
rect 3580 2576 3588 2584
rect 3788 2576 3796 2584
rect 3916 2576 3924 2584
rect 4076 2576 4084 2584
rect 4380 2576 4388 2584
rect 4444 2576 4452 2584
rect 4476 2576 4484 2584
rect 4604 2576 4612 2584
rect 4668 2576 4676 2584
rect 4988 2576 4996 2584
rect 5004 2576 5012 2584
rect 5500 2576 5508 2584
rect 1052 2556 1060 2564
rect 1228 2556 1236 2564
rect 1404 2556 1412 2564
rect 2108 2556 2116 2564
rect 2716 2556 2724 2564
rect 2908 2556 2916 2564
rect 2956 2556 2964 2564
rect 2972 2556 2980 2564
rect 3036 2556 3044 2564
rect 3388 2556 3396 2564
rect 4428 2556 4436 2564
rect 124 2536 132 2544
rect 252 2536 260 2544
rect 1324 2536 1332 2544
rect 1388 2536 1396 2544
rect 1420 2536 1428 2544
rect 2060 2536 2068 2544
rect 2316 2536 2324 2544
rect 2428 2536 2436 2544
rect 3068 2536 3076 2544
rect 3244 2536 3252 2544
rect 3292 2536 3300 2544
rect 3484 2536 3492 2544
rect 3564 2536 3572 2544
rect 3708 2536 3716 2544
rect 3772 2536 3780 2544
rect 3884 2536 3892 2544
rect 4140 2536 4148 2544
rect 4188 2536 4196 2544
rect 4236 2536 4244 2544
rect 4284 2536 4292 2544
rect 4636 2536 4644 2544
rect 4668 2536 4676 2544
rect 4732 2536 4740 2544
rect 4796 2536 4804 2544
rect 4940 2536 4948 2544
rect 5004 2536 5012 2544
rect 5036 2536 5044 2544
rect 5164 2536 5172 2544
rect 5372 2536 5380 2544
rect 716 2516 724 2524
rect 972 2516 980 2524
rect 1084 2516 1092 2524
rect 1772 2516 1780 2524
rect 1900 2516 1908 2524
rect 2076 2516 2084 2524
rect 2412 2516 2420 2524
rect 2444 2516 2452 2524
rect 396 2496 404 2504
rect 924 2496 932 2504
rect 1164 2496 1172 2504
rect 1420 2496 1428 2504
rect 1484 2496 1492 2504
rect 1500 2496 1508 2504
rect 3228 2516 3236 2524
rect 3580 2516 3588 2524
rect 3612 2516 3620 2524
rect 4076 2516 4084 2524
rect 4620 2516 4628 2524
rect 4924 2516 4932 2524
rect 5020 2516 5028 2524
rect 5340 2516 5348 2524
rect 5500 2516 5508 2524
rect 2620 2496 2628 2504
rect 3260 2496 3268 2504
rect 3564 2496 3572 2504
rect 3596 2496 3604 2504
rect 3980 2496 3988 2504
rect 4028 2496 4036 2504
rect 4572 2496 4580 2504
rect 4604 2496 4612 2504
rect 4780 2496 4788 2504
rect 4812 2496 4820 2504
rect 4908 2496 4916 2504
rect 4956 2496 4964 2504
rect 5292 2496 5300 2504
rect 444 2476 452 2484
rect 3628 2476 3636 2484
rect 3724 2476 3732 2484
rect 5244 2476 5252 2484
rect 3228 2456 3236 2464
rect 3292 2456 3300 2464
rect 3340 2456 3348 2464
rect 3692 2456 3700 2464
rect 3996 2456 4004 2464
rect 1708 2436 1716 2444
rect 3148 2436 3156 2444
rect 4908 2436 4916 2444
rect 1372 2416 1380 2424
rect 5356 2416 5364 2424
rect 252 2396 260 2404
rect 412 2396 420 2404
rect 2108 2396 2116 2404
rect 4428 2396 4436 2404
rect 5116 2396 5124 2404
rect 1996 2376 2004 2384
rect 3212 2376 3220 2384
rect 4268 2376 4276 2384
rect 4844 2376 4852 2384
rect 5036 2376 5044 2384
rect 1676 2356 1684 2364
rect 1756 2356 1764 2364
rect 1788 2356 1796 2364
rect 2124 2356 2132 2364
rect 3212 2356 3220 2364
rect 3516 2356 3524 2364
rect 4332 2356 4340 2364
rect 284 2336 292 2344
rect 556 2336 564 2344
rect 988 2336 996 2344
rect 1164 2336 1172 2344
rect 1900 2336 1908 2344
rect 1948 2336 1956 2344
rect 1996 2336 2004 2344
rect 2028 2336 2036 2344
rect 2684 2336 2692 2344
rect 2876 2336 2884 2344
rect 4332 2336 4340 2344
rect 4348 2336 4356 2344
rect 4860 2336 4868 2344
rect 684 2316 692 2324
rect 748 2316 756 2324
rect 892 2316 900 2324
rect 956 2296 964 2304
rect 972 2296 980 2304
rect 1276 2296 1284 2304
rect 1308 2316 1316 2324
rect 1500 2316 1508 2324
rect 2092 2316 2100 2324
rect 4572 2316 4580 2324
rect 4956 2316 4964 2324
rect 5004 2316 5012 2324
rect 5132 2316 5140 2324
rect 5452 2316 5460 2324
rect 5500 2316 5508 2324
rect 1804 2296 1812 2304
rect 1852 2296 1860 2304
rect 2700 2296 2708 2304
rect 3260 2296 3268 2304
rect 3500 2296 3508 2304
rect 3532 2296 3540 2304
rect 3612 2296 3620 2304
rect 3708 2296 3716 2304
rect 4220 2296 4228 2304
rect 4284 2296 4292 2304
rect 4476 2296 4484 2304
rect 4748 2296 4756 2304
rect 140 2276 148 2284
rect 924 2276 932 2284
rect 940 2276 948 2284
rect 1404 2276 1412 2284
rect 1420 2276 1428 2284
rect 1788 2276 1796 2284
rect 1868 2276 1876 2284
rect 2028 2276 2036 2284
rect 2044 2276 2052 2284
rect 2636 2276 2644 2284
rect 2780 2276 2788 2284
rect 2908 2276 2916 2284
rect 3068 2276 3076 2284
rect 3116 2276 3124 2284
rect 3196 2276 3204 2284
rect 76 2256 84 2264
rect 988 2256 996 2264
rect 1036 2256 1044 2264
rect 1420 2256 1428 2264
rect 2140 2256 2148 2264
rect 2220 2256 2228 2264
rect 3276 2256 3284 2264
rect 3804 2276 3812 2284
rect 3884 2276 3892 2284
rect 4204 2276 4212 2284
rect 4268 2276 4276 2284
rect 4300 2276 4308 2284
rect 4460 2276 4468 2284
rect 4588 2276 4596 2284
rect 4636 2276 4644 2284
rect 5100 2276 5108 2284
rect 5260 2276 5268 2284
rect 3708 2256 3716 2264
rect 3836 2256 3844 2264
rect 4012 2256 4020 2264
rect 4924 2256 4932 2264
rect 5180 2256 5188 2264
rect 5228 2256 5236 2264
rect 828 2236 836 2244
rect 1164 2236 1172 2244
rect 1228 2236 1236 2244
rect 1676 2236 1684 2244
rect 1724 2236 1732 2244
rect 2012 2236 2020 2244
rect 2044 2236 2052 2244
rect 2156 2236 2164 2244
rect 2492 2236 2500 2244
rect 2508 2236 2516 2244
rect 2668 2236 2676 2244
rect 3868 2236 3876 2244
rect 3996 2236 4004 2244
rect 4172 2236 4180 2244
rect 4348 2236 4356 2244
rect 4364 2236 4372 2244
rect 4796 2236 4804 2244
rect 4892 2236 4900 2244
rect 5020 2236 5028 2244
rect 636 2216 644 2224
rect 1708 2216 1716 2224
rect 1996 2216 2004 2224
rect 2764 2216 2772 2224
rect 2876 2216 2884 2224
rect 3308 2216 3316 2224
rect 3564 2216 3572 2224
rect 3676 2216 3684 2224
rect 4780 2216 4788 2224
rect 4796 2216 4804 2224
rect 4812 2216 4820 2224
rect 5100 2216 5108 2224
rect 1116 2196 1124 2204
rect 1308 2196 1316 2204
rect 1532 2196 1540 2204
rect 1564 2196 1572 2204
rect 1692 2196 1700 2204
rect 1964 2196 1972 2204
rect 620 2176 628 2184
rect 956 2176 964 2184
rect 972 2176 980 2184
rect 1036 2176 1044 2184
rect 1084 2176 1092 2184
rect 1292 2176 1300 2184
rect 1692 2176 1700 2184
rect 2716 2196 2724 2204
rect 3804 2196 3812 2204
rect 4108 2196 4116 2204
rect 4156 2196 4164 2204
rect 4236 2196 4244 2204
rect 4956 2196 4964 2204
rect 5004 2196 5012 2204
rect 5244 2196 5252 2204
rect 2332 2176 2340 2184
rect 2444 2176 2452 2184
rect 2988 2176 2996 2184
rect 3228 2176 3236 2184
rect 3516 2176 3524 2184
rect 3660 2176 3668 2184
rect 3708 2176 3716 2184
rect 3852 2176 3860 2184
rect 4604 2176 4612 2184
rect 4668 2176 4676 2184
rect 4700 2176 4708 2184
rect 5148 2176 5156 2184
rect 5228 2176 5236 2184
rect 1116 2156 1124 2164
rect 1404 2156 1412 2164
rect 1532 2156 1540 2164
rect 1580 2156 1588 2164
rect 1932 2156 1940 2164
rect 2428 2156 2436 2164
rect 2684 2156 2692 2164
rect 172 2136 180 2144
rect 348 2136 356 2144
rect 444 2136 452 2144
rect 476 2136 484 2144
rect 540 2136 548 2144
rect 652 2136 660 2144
rect 732 2136 740 2144
rect 764 2136 772 2144
rect 892 2136 900 2144
rect 1196 2136 1204 2144
rect 1468 2136 1476 2144
rect 1516 2136 1524 2144
rect 1612 2136 1620 2144
rect 1724 2136 1732 2144
rect 1740 2136 1748 2144
rect 2220 2136 2228 2144
rect 2284 2136 2292 2144
rect 2300 2136 2308 2144
rect 2444 2136 2452 2144
rect 2556 2136 2564 2144
rect 2588 2136 2596 2144
rect 2780 2136 2788 2144
rect 3084 2156 3092 2164
rect 3404 2156 3412 2164
rect 3548 2156 3556 2164
rect 4108 2156 4116 2164
rect 4268 2156 4276 2164
rect 4812 2156 4820 2164
rect 5420 2156 5428 2164
rect 3020 2136 3028 2144
rect 3132 2136 3140 2144
rect 3644 2136 3652 2144
rect 3724 2136 3732 2144
rect 3900 2136 3908 2144
rect 4556 2136 4564 2144
rect 5100 2136 5108 2144
rect 5484 2136 5492 2144
rect 12 2116 20 2124
rect 1084 2116 1092 2124
rect 1388 2116 1396 2124
rect 1404 2116 1412 2124
rect 1948 2116 1956 2124
rect 2012 2116 2020 2124
rect 2028 2116 2036 2124
rect 2428 2116 2436 2124
rect 2684 2116 2692 2124
rect 2732 2116 2740 2124
rect 2988 2116 2996 2124
rect 3660 2116 3668 2124
rect 4044 2116 4052 2124
rect 4412 2116 4420 2124
rect 4556 2116 4564 2124
rect 4844 2116 4852 2124
rect 4956 2116 4964 2124
rect 4988 2116 4996 2124
rect 5180 2116 5188 2124
rect 348 2096 356 2104
rect 396 2096 404 2104
rect 748 2096 756 2104
rect 828 2096 836 2104
rect 1260 2096 1268 2104
rect 1324 2096 1332 2104
rect 1340 2096 1348 2104
rect 1484 2096 1492 2104
rect 1676 2096 1684 2104
rect 1708 2096 1716 2104
rect 1980 2096 1988 2104
rect 2620 2096 2628 2104
rect 2924 2096 2932 2104
rect 3244 2096 3252 2104
rect 3820 2096 3828 2104
rect 3964 2096 3972 2104
rect 4284 2096 4292 2104
rect 4620 2096 4628 2104
rect 4716 2096 4724 2104
rect 4908 2096 4916 2104
rect 5036 2096 5044 2104
rect 5292 2096 5300 2104
rect 1132 2076 1140 2084
rect 1148 2076 1156 2084
rect 1180 2076 1188 2084
rect 1452 2076 1460 2084
rect 2060 2076 2068 2084
rect 2636 2076 2644 2084
rect 3404 2076 3412 2084
rect 3564 2076 3572 2084
rect 5260 2076 5268 2084
rect 5388 2076 5396 2084
rect 5452 2076 5460 2084
rect 748 2056 756 2064
rect 2556 2056 2564 2064
rect 2604 2056 2612 2064
rect 3388 2056 3396 2064
rect 4092 2056 4100 2064
rect 4188 2056 4196 2064
rect 5148 2056 5156 2064
rect 1676 2036 1684 2044
rect 1820 2036 1828 2044
rect 2492 2036 2500 2044
rect 844 2016 852 2024
rect 1132 2016 1140 2024
rect 2732 2016 2740 2024
rect 1564 1996 1572 2004
rect 1996 1996 2004 2004
rect 2108 1996 2116 2004
rect 2236 1996 2244 2004
rect 2940 1996 2948 2004
rect 812 1976 820 1984
rect 844 1976 852 1984
rect 2684 1976 2692 1984
rect 3260 1976 3268 1984
rect 3308 1976 3316 1984
rect 4092 1976 4100 1984
rect 4108 1976 4116 1984
rect 5436 1976 5444 1984
rect 764 1956 772 1964
rect 812 1956 820 1964
rect 1212 1956 1220 1964
rect 1612 1956 1620 1964
rect 1868 1956 1876 1964
rect 2092 1956 2100 1964
rect 2156 1956 2164 1964
rect 2188 1956 2196 1964
rect 2460 1956 2468 1964
rect 2748 1956 2756 1964
rect 3180 1956 3188 1964
rect 3372 1956 3380 1964
rect 4492 1956 4500 1964
rect 5244 1956 5252 1964
rect 844 1936 852 1944
rect 1180 1936 1188 1944
rect 1900 1936 1908 1944
rect 1916 1936 1924 1944
rect 5244 1936 5252 1944
rect 348 1916 356 1924
rect 460 1916 468 1924
rect 492 1916 500 1924
rect 1260 1916 1268 1924
rect 1292 1916 1300 1924
rect 1948 1916 1956 1924
rect 2476 1916 2484 1924
rect 2684 1916 2692 1924
rect 2716 1916 2724 1924
rect 3676 1916 3684 1924
rect 3724 1916 3732 1924
rect 4780 1916 4788 1924
rect 4892 1916 4900 1924
rect 860 1896 868 1904
rect 892 1896 900 1904
rect 940 1896 948 1904
rect 956 1896 964 1904
rect 988 1896 996 1904
rect 1212 1896 1220 1904
rect 1980 1896 1988 1904
rect 2252 1896 2260 1904
rect 2588 1896 2596 1904
rect 2972 1896 2980 1904
rect 3196 1896 3204 1904
rect 3228 1896 3236 1904
rect 3516 1896 3524 1904
rect 3708 1896 3716 1904
rect 4108 1896 4116 1904
rect 4268 1896 4276 1904
rect 4620 1896 4628 1904
rect 4780 1896 4788 1904
rect 4828 1896 4836 1904
rect 108 1876 116 1884
rect 204 1876 212 1884
rect 236 1876 244 1884
rect 380 1876 388 1884
rect 1420 1876 1428 1884
rect 1468 1876 1476 1884
rect 1500 1876 1508 1884
rect 140 1856 148 1864
rect 364 1856 372 1864
rect 396 1856 404 1864
rect 620 1856 628 1864
rect 764 1856 772 1864
rect 572 1836 580 1844
rect 604 1836 612 1844
rect 700 1836 708 1844
rect 716 1836 724 1844
rect 748 1836 756 1844
rect 1068 1836 1076 1844
rect 1148 1836 1156 1844
rect 1228 1856 1236 1864
rect 1324 1856 1332 1864
rect 1884 1876 1892 1884
rect 2508 1876 2516 1884
rect 2844 1876 2852 1884
rect 2924 1876 2932 1884
rect 3420 1876 3428 1884
rect 3884 1876 3892 1884
rect 4332 1876 4340 1884
rect 4908 1876 4916 1884
rect 5020 1876 5028 1884
rect 5068 1876 5076 1884
rect 5388 1876 5396 1884
rect 5500 1876 5508 1884
rect 1772 1856 1780 1864
rect 1868 1856 1876 1864
rect 1948 1856 1956 1864
rect 2124 1856 2132 1864
rect 2172 1856 2180 1864
rect 2332 1856 2340 1864
rect 2540 1856 2548 1864
rect 2988 1856 2996 1864
rect 3004 1856 3012 1864
rect 3548 1856 3556 1864
rect 3708 1856 3716 1864
rect 3756 1856 3764 1864
rect 3980 1856 3988 1864
rect 4412 1856 4420 1864
rect 4636 1856 4644 1864
rect 4700 1856 4708 1864
rect 1276 1836 1284 1844
rect 2108 1836 2116 1844
rect 2300 1836 2308 1844
rect 2460 1836 2468 1844
rect 460 1816 468 1824
rect 1388 1816 1396 1824
rect 2092 1816 2100 1824
rect 2572 1816 2580 1824
rect 3404 1816 3412 1824
rect 3964 1836 3972 1844
rect 4092 1836 4100 1844
rect 5276 1836 5284 1844
rect 4812 1816 4820 1824
rect 4844 1816 4852 1824
rect 4876 1816 4884 1824
rect 5228 1816 5236 1824
rect 60 1796 68 1804
rect 1276 1796 1284 1804
rect 316 1776 324 1784
rect 60 1756 68 1764
rect 428 1756 436 1764
rect 524 1756 532 1764
rect 892 1776 900 1784
rect 940 1776 948 1784
rect 972 1776 980 1784
rect 1036 1776 1044 1784
rect 1148 1776 1156 1784
rect 1324 1776 1332 1784
rect 1468 1776 1476 1784
rect 1676 1776 1684 1784
rect 2124 1796 2132 1804
rect 2268 1796 2276 1804
rect 2428 1796 2436 1804
rect 2556 1796 2564 1804
rect 2716 1796 2724 1804
rect 2908 1796 2916 1804
rect 3292 1796 3300 1804
rect 3484 1796 3492 1804
rect 4188 1796 4196 1804
rect 4348 1796 4356 1804
rect 4428 1796 4436 1804
rect 4620 1796 4628 1804
rect 4716 1796 4724 1804
rect 4748 1796 4756 1804
rect 5372 1796 5380 1804
rect 1852 1776 1860 1784
rect 1884 1776 1892 1784
rect 2524 1776 2532 1784
rect 3580 1776 3588 1784
rect 3996 1776 4004 1784
rect 4076 1776 4084 1784
rect 4284 1776 4292 1784
rect 5132 1776 5140 1784
rect 5292 1776 5300 1784
rect 668 1756 676 1764
rect 812 1756 820 1764
rect 2060 1756 2068 1764
rect 2092 1756 2100 1764
rect 2284 1756 2292 1764
rect 2316 1756 2324 1764
rect 2396 1756 2404 1764
rect 2604 1756 2612 1764
rect 2668 1756 2676 1764
rect 3436 1756 3444 1764
rect 3788 1756 3796 1764
rect 3852 1756 3860 1764
rect 4092 1756 4100 1764
rect 4140 1756 4148 1764
rect 4620 1756 4628 1764
rect 4988 1756 4996 1764
rect 5004 1756 5012 1764
rect 5052 1756 5060 1764
rect 5084 1756 5092 1764
rect 5340 1756 5348 1764
rect 268 1736 276 1744
rect 444 1736 452 1744
rect 508 1736 516 1744
rect 1436 1736 1444 1744
rect 2076 1736 2084 1744
rect 2268 1736 2276 1744
rect 2828 1736 2836 1744
rect 2876 1736 2884 1744
rect 2940 1736 2948 1744
rect 3260 1736 3268 1744
rect 3644 1736 3652 1744
rect 3692 1736 3700 1744
rect 3836 1736 3844 1744
rect 4252 1736 4260 1744
rect 4684 1736 4692 1744
rect 4892 1736 4900 1744
rect 5292 1736 5300 1744
rect 5372 1736 5380 1744
rect 60 1716 68 1724
rect 316 1716 324 1724
rect 604 1716 612 1724
rect 652 1716 660 1724
rect 764 1716 772 1724
rect 1244 1716 1252 1724
rect 1724 1716 1732 1724
rect 1740 1716 1748 1724
rect 2284 1716 2292 1724
rect 2332 1716 2340 1724
rect 2428 1716 2436 1724
rect 2460 1716 2468 1724
rect 2572 1716 2580 1724
rect 3548 1716 3556 1724
rect 4940 1716 4948 1724
rect 5004 1716 5012 1724
rect 5036 1716 5044 1724
rect 492 1696 500 1704
rect 556 1696 564 1704
rect 796 1696 804 1704
rect 924 1696 932 1704
rect 956 1696 964 1704
rect 1116 1696 1124 1704
rect 1196 1696 1204 1704
rect 3052 1696 3060 1704
rect 3372 1696 3380 1704
rect 3708 1696 3716 1704
rect 3724 1696 3732 1704
rect 3932 1696 3940 1704
rect 220 1676 228 1684
rect 924 1676 932 1684
rect 1404 1676 1412 1684
rect 1676 1676 1684 1684
rect 1900 1676 1908 1684
rect 1916 1676 1924 1684
rect 2364 1676 2372 1684
rect 4124 1696 4132 1704
rect 4700 1696 4708 1704
rect 4940 1696 4948 1704
rect 5116 1696 5124 1704
rect 3964 1676 3972 1684
rect 4348 1676 4356 1684
rect 4828 1676 4836 1684
rect 1132 1656 1140 1664
rect 1884 1656 1892 1664
rect 3724 1656 3732 1664
rect 3916 1656 3924 1664
rect 4508 1656 4516 1664
rect 4812 1656 4820 1664
rect 1180 1636 1188 1644
rect 1836 1636 1844 1644
rect 1980 1636 1988 1644
rect 2540 1636 2548 1644
rect 4732 1636 4740 1644
rect 140 1616 148 1624
rect 188 1616 196 1624
rect 1916 1616 1924 1624
rect 1948 1616 1956 1624
rect 3724 1616 3732 1624
rect 4508 1616 4516 1624
rect 492 1596 500 1604
rect 2428 1596 2436 1604
rect 2652 1596 2660 1604
rect 4044 1596 4052 1604
rect 1676 1576 1684 1584
rect 3724 1576 3732 1584
rect 4524 1576 4532 1584
rect 4540 1576 4548 1584
rect 4652 1576 4660 1584
rect 4780 1576 4788 1584
rect 1596 1556 1604 1564
rect 1644 1556 1652 1564
rect 3500 1556 3508 1564
rect 636 1536 644 1544
rect 860 1536 868 1544
rect 1004 1536 1012 1544
rect 1020 1536 1028 1544
rect 1228 1536 1236 1544
rect 1388 1536 1396 1544
rect 1612 1536 1620 1544
rect 2044 1536 2052 1544
rect 3452 1536 3460 1544
rect 3580 1536 3588 1544
rect 3596 1536 3604 1544
rect 3692 1536 3700 1544
rect 4124 1536 4132 1544
rect 4220 1536 4228 1544
rect 4268 1536 4276 1544
rect 4796 1536 4804 1544
rect 4940 1536 4948 1544
rect 4972 1536 4980 1544
rect 380 1516 388 1524
rect 1196 1516 1204 1524
rect 1452 1516 1460 1524
rect 2028 1516 2036 1524
rect 2684 1516 2692 1524
rect 2796 1516 2804 1524
rect 3180 1516 3188 1524
rect 3804 1516 3812 1524
rect 4652 1516 4660 1524
rect 4764 1516 4772 1524
rect 4908 1516 4916 1524
rect 5292 1516 5300 1524
rect 5532 1516 5540 1524
rect 604 1496 612 1504
rect 1148 1496 1156 1504
rect 1356 1496 1364 1504
rect 1500 1496 1508 1504
rect 1644 1496 1652 1504
rect 1660 1496 1668 1504
rect 188 1476 196 1484
rect 828 1476 836 1484
rect 940 1476 948 1484
rect 1100 1476 1108 1484
rect 1116 1476 1124 1484
rect 1212 1476 1220 1484
rect 1740 1476 1748 1484
rect 1756 1476 1764 1484
rect 1868 1476 1876 1484
rect 3244 1496 3252 1504
rect 3276 1496 3284 1504
rect 3292 1496 3300 1504
rect 3484 1496 3492 1504
rect 3692 1496 3700 1504
rect 3900 1496 3908 1504
rect 3948 1496 3956 1504
rect 4428 1496 4436 1504
rect 4924 1496 4932 1504
rect 4972 1496 4980 1504
rect 5036 1496 5044 1504
rect 2300 1476 2308 1484
rect 2732 1476 2740 1484
rect 2956 1476 2964 1484
rect 3084 1476 3092 1484
rect 3868 1476 3876 1484
rect 4956 1476 4964 1484
rect 76 1456 84 1464
rect 172 1456 180 1464
rect 476 1456 484 1464
rect 572 1456 580 1464
rect 652 1456 660 1464
rect 780 1456 788 1464
rect 972 1456 980 1464
rect 1164 1456 1172 1464
rect 1308 1456 1316 1464
rect 1324 1456 1332 1464
rect 1388 1456 1396 1464
rect 1484 1456 1492 1464
rect 1500 1456 1508 1464
rect 2124 1456 2132 1464
rect 2396 1456 2404 1464
rect 2748 1456 2756 1464
rect 3164 1456 3172 1464
rect 3260 1456 3268 1464
rect 3660 1456 3668 1464
rect 3852 1456 3860 1464
rect 3996 1456 4004 1464
rect 4156 1456 4164 1464
rect 4172 1456 4180 1464
rect 4844 1456 4852 1464
rect 5132 1456 5140 1464
rect 1260 1436 1268 1444
rect 2684 1436 2692 1444
rect 652 1416 660 1424
rect 1068 1416 1076 1424
rect 1388 1416 1396 1424
rect 1516 1416 1524 1424
rect 1580 1416 1588 1424
rect 1612 1416 1620 1424
rect 1964 1416 1972 1424
rect 2156 1416 2164 1424
rect 2252 1416 2260 1424
rect 3084 1436 3092 1444
rect 3132 1436 3140 1444
rect 3932 1436 3940 1444
rect 4412 1436 4420 1444
rect 4428 1436 4436 1444
rect 3388 1416 3396 1424
rect 3516 1416 3524 1424
rect 3548 1416 3556 1424
rect 3564 1416 3572 1424
rect 4044 1416 4052 1424
rect 4636 1416 4644 1424
rect 4812 1416 4820 1424
rect 188 1396 196 1404
rect 1036 1396 1044 1404
rect 1340 1396 1348 1404
rect 1532 1396 1540 1404
rect 1756 1396 1764 1404
rect 1788 1396 1796 1404
rect 1836 1396 1844 1404
rect 2108 1396 2116 1404
rect 3004 1396 3012 1404
rect 3276 1396 3284 1404
rect 3948 1396 3956 1404
rect 4124 1396 4132 1404
rect 4220 1396 4228 1404
rect 5452 1396 5460 1404
rect 988 1376 996 1384
rect 1180 1376 1188 1384
rect 1484 1376 1492 1384
rect 1676 1376 1684 1384
rect 1692 1376 1700 1384
rect 2908 1376 2916 1384
rect 3468 1376 3476 1384
rect 3500 1376 3508 1384
rect 3660 1376 3668 1384
rect 3708 1376 3716 1384
rect 4492 1376 4500 1384
rect 4572 1376 4580 1384
rect 5356 1376 5364 1384
rect 124 1356 132 1364
rect 460 1356 468 1364
rect 620 1356 628 1364
rect 636 1356 644 1364
rect 732 1356 740 1364
rect 1068 1356 1076 1364
rect 1340 1356 1348 1364
rect 1404 1356 1412 1364
rect 2092 1356 2100 1364
rect 2412 1356 2420 1364
rect 2508 1356 2516 1364
rect 3100 1356 3108 1364
rect 3244 1356 3252 1364
rect 3324 1356 3332 1364
rect 3388 1356 3396 1364
rect 3484 1356 3492 1364
rect 3612 1356 3620 1364
rect 3692 1356 3700 1364
rect 3884 1356 3892 1364
rect 3916 1356 3924 1364
rect 3980 1356 3988 1364
rect 4012 1356 4020 1364
rect 460 1336 468 1344
rect 524 1336 532 1344
rect 540 1336 548 1344
rect 588 1336 596 1344
rect 812 1336 820 1344
rect 1164 1336 1172 1344
rect 1180 1336 1188 1344
rect 1196 1336 1204 1344
rect 1372 1336 1380 1344
rect 1420 1336 1428 1344
rect 1596 1336 1604 1344
rect 2236 1336 2244 1344
rect 2300 1336 2308 1344
rect 2636 1336 2644 1344
rect 3836 1336 3844 1344
rect 4188 1356 4196 1364
rect 4796 1356 4804 1364
rect 4956 1356 4964 1364
rect 5036 1356 5044 1364
rect 5068 1356 5076 1364
rect 5324 1356 5332 1364
rect 4572 1336 4580 1344
rect 5308 1336 5316 1344
rect 252 1316 260 1324
rect 460 1316 468 1324
rect 1212 1316 1220 1324
rect 1340 1316 1348 1324
rect 2348 1316 2356 1324
rect 2556 1316 2564 1324
rect 2700 1316 2708 1324
rect 3708 1316 3716 1324
rect 3740 1316 3748 1324
rect 4108 1316 4116 1324
rect 4588 1316 4596 1324
rect 4732 1316 4740 1324
rect 5148 1316 5156 1324
rect 620 1296 628 1304
rect 844 1296 852 1304
rect 924 1296 932 1304
rect 1612 1296 1620 1304
rect 1900 1296 1908 1304
rect 1932 1296 1940 1304
rect 2332 1296 2340 1304
rect 2492 1296 2500 1304
rect 2796 1296 2804 1304
rect 3004 1296 3012 1304
rect 3036 1296 3044 1304
rect 4156 1296 4164 1304
rect 4204 1296 4212 1304
rect 1340 1276 1348 1284
rect 1452 1276 1460 1284
rect 1804 1276 1812 1284
rect 2156 1276 2164 1284
rect 2604 1276 2612 1284
rect 2716 1276 2724 1284
rect 2764 1276 2772 1284
rect 3164 1276 3172 1284
rect 3180 1276 3188 1284
rect 3948 1276 3956 1284
rect 4236 1276 4244 1284
rect 4316 1296 4324 1304
rect 5308 1296 5316 1304
rect 4972 1276 4980 1284
rect 2716 1256 2724 1264
rect 3212 1256 3220 1264
rect 3292 1256 3300 1264
rect 3340 1256 3348 1264
rect 3516 1256 3524 1264
rect 4812 1256 4820 1264
rect 1164 1236 1172 1244
rect 1388 1236 1396 1244
rect 44 1216 52 1224
rect 1116 1216 1124 1224
rect 4476 1216 4484 1224
rect 4812 1216 4820 1224
rect 956 1196 964 1204
rect 1084 1196 1092 1204
rect 1836 1196 1844 1204
rect 1852 1196 1860 1204
rect 2316 1196 2324 1204
rect 5068 1196 5076 1204
rect 268 1176 276 1184
rect 1788 1176 1796 1184
rect 1804 1176 1812 1184
rect 2524 1176 2532 1184
rect 3148 1176 3156 1184
rect 3708 1176 3716 1184
rect 3948 1176 3956 1184
rect 4092 1176 4100 1184
rect 60 1156 68 1164
rect 3292 1156 3300 1164
rect 3932 1156 3940 1164
rect 4588 1156 4596 1164
rect 540 1136 548 1144
rect 620 1136 628 1144
rect 1052 1136 1060 1144
rect 1164 1136 1172 1144
rect 1292 1136 1300 1144
rect 1388 1136 1396 1144
rect 1596 1136 1604 1144
rect 1612 1136 1620 1144
rect 2044 1136 2052 1144
rect 412 1116 420 1124
rect 444 1116 452 1124
rect 1196 1116 1204 1124
rect 1388 1116 1396 1124
rect 1740 1116 1748 1124
rect 1756 1116 1764 1124
rect 1788 1116 1796 1124
rect 1964 1116 1972 1124
rect 2540 1116 2548 1124
rect 2620 1116 2628 1124
rect 3788 1136 3796 1144
rect 5164 1136 5172 1144
rect 3452 1116 3460 1124
rect 3804 1116 3812 1124
rect 3948 1116 3956 1124
rect 4332 1116 4340 1124
rect 4364 1116 4372 1124
rect 4652 1116 4660 1124
rect 4700 1116 4708 1124
rect 4748 1116 4756 1124
rect 4764 1116 4772 1124
rect 4812 1116 4820 1124
rect 4972 1116 4980 1124
rect 5324 1116 5332 1124
rect 188 1096 196 1104
rect 812 1096 820 1104
rect 828 1096 836 1104
rect 2764 1096 2772 1104
rect 2812 1096 2820 1104
rect 3676 1096 3684 1104
rect 3804 1096 3812 1104
rect 4044 1096 4052 1104
rect 4460 1096 4468 1104
rect 4860 1096 4868 1104
rect 4876 1096 4884 1104
rect 5244 1096 5252 1104
rect 5260 1096 5268 1104
rect 5292 1096 5300 1104
rect 44 1076 52 1084
rect 172 1076 180 1084
rect 1228 1076 1236 1084
rect 1292 1076 1300 1084
rect 1308 1076 1316 1084
rect 1372 1076 1380 1084
rect 1436 1076 1444 1084
rect 1484 1076 1492 1084
rect 1660 1076 1668 1084
rect 1836 1076 1844 1084
rect 124 1056 132 1064
rect 204 1056 212 1064
rect 284 1056 292 1064
rect 460 1056 468 1064
rect 860 1056 868 1064
rect 940 1056 948 1064
rect 988 1056 996 1064
rect 1468 1056 1476 1064
rect 1724 1056 1732 1064
rect 2268 1076 2276 1084
rect 2396 1076 2404 1084
rect 2444 1076 2452 1084
rect 2812 1076 2820 1084
rect 3276 1076 3284 1084
rect 3820 1076 3828 1084
rect 3836 1076 3844 1084
rect 4620 1076 4628 1084
rect 5164 1076 5172 1084
rect 5356 1076 5364 1084
rect 1948 1056 1956 1064
rect 2188 1056 2196 1064
rect 2428 1056 2436 1064
rect 2700 1056 2708 1064
rect 3436 1056 3444 1064
rect 3628 1056 3636 1064
rect 3724 1056 3732 1064
rect 4364 1056 4372 1064
rect 4492 1056 4500 1064
rect 4796 1056 4804 1064
rect 5452 1056 5460 1064
rect 284 1036 292 1044
rect 780 1036 788 1044
rect 844 1036 852 1044
rect 1116 1036 1124 1044
rect 1324 1036 1332 1044
rect 1548 1036 1556 1044
rect 2524 1036 2532 1044
rect 3116 1036 3124 1044
rect 3324 1036 3332 1044
rect 3516 1036 3524 1044
rect 4956 1036 4964 1044
rect 5068 1036 5076 1044
rect 5148 1036 5156 1044
rect 5292 1036 5300 1044
rect 636 1016 644 1024
rect 684 1016 692 1024
rect 716 1016 724 1024
rect 812 1016 820 1024
rect 844 1016 852 1024
rect 1740 1016 1748 1024
rect 1820 1016 1828 1024
rect 1884 1016 1892 1024
rect 1948 1016 1956 1024
rect 2492 1016 2500 1024
rect 3068 1016 3076 1024
rect 3164 1016 3172 1024
rect 3260 1016 3268 1024
rect 4092 1016 4100 1024
rect 4652 1016 4660 1024
rect 5308 1016 5316 1024
rect 796 996 804 1004
rect 860 996 868 1004
rect 972 996 980 1004
rect 1036 996 1044 1004
rect 1372 996 1380 1004
rect 1468 996 1476 1004
rect 1532 996 1540 1004
rect 1900 996 1908 1004
rect 1964 996 1972 1004
rect 2204 996 2212 1004
rect 2444 996 2452 1004
rect 2828 996 2836 1004
rect 3100 996 3108 1004
rect 3292 996 3300 1004
rect 3436 996 3444 1004
rect 3836 996 3844 1004
rect 4012 996 4020 1004
rect 4556 996 4564 1004
rect 4716 996 4724 1004
rect 4732 996 4740 1004
rect 4972 996 4980 1004
rect 5036 996 5044 1004
rect 380 976 388 984
rect 396 976 404 984
rect 556 976 564 984
rect 1500 976 1508 984
rect 1516 976 1524 984
rect 2364 976 2372 984
rect 2668 976 2676 984
rect 3340 976 3348 984
rect 3564 976 3572 984
rect 3964 976 3972 984
rect 4716 976 4724 984
rect 5004 976 5012 984
rect 5308 976 5316 984
rect 5388 976 5396 984
rect 124 956 132 964
rect 268 956 276 964
rect 396 956 404 964
rect 1484 956 1492 964
rect 1740 956 1748 964
rect 1852 956 1860 964
rect 2476 956 2484 964
rect 2780 956 2788 964
rect 2828 956 2836 964
rect 3052 956 3060 964
rect 3388 956 3396 964
rect 3452 956 3460 964
rect 3820 956 3828 964
rect 3836 956 3844 964
rect 3932 956 3940 964
rect 4060 956 4068 964
rect 4348 956 4356 964
rect 5132 956 5140 964
rect 5388 956 5396 964
rect 188 936 196 944
rect 236 936 244 944
rect 460 936 468 944
rect 828 936 836 944
rect 892 936 900 944
rect 1020 936 1028 944
rect 1052 936 1060 944
rect 1324 936 1332 944
rect 1500 936 1508 944
rect 1580 936 1588 944
rect 2220 936 2228 944
rect 2332 936 2340 944
rect 2412 936 2420 944
rect 2428 936 2436 944
rect 2876 936 2884 944
rect 2908 936 2916 944
rect 3084 936 3092 944
rect 3644 936 3652 944
rect 4540 936 4548 944
rect 4572 936 4580 944
rect 5100 936 5108 944
rect 5404 936 5412 944
rect 5436 936 5444 944
rect 1212 916 1220 924
rect 1244 916 1252 924
rect 1884 916 1892 924
rect 2396 916 2404 924
rect 2556 916 2564 924
rect 348 896 356 904
rect 1004 896 1012 904
rect 1532 896 1540 904
rect 1676 896 1684 904
rect 2428 896 2436 904
rect 2732 896 2740 904
rect 2748 896 2756 904
rect 2764 896 2772 904
rect 3740 916 3748 924
rect 3756 916 3764 924
rect 3916 916 3924 924
rect 4204 916 4212 924
rect 4956 916 4964 924
rect 5084 916 5092 924
rect 5212 916 5220 924
rect 2988 896 2996 904
rect 3276 896 3284 904
rect 3404 896 3412 904
rect 460 876 468 884
rect 508 876 516 884
rect 892 876 900 884
rect 940 876 948 884
rect 2284 876 2292 884
rect 2716 876 2724 884
rect 2860 876 2868 884
rect 2940 876 2948 884
rect 4972 896 4980 904
rect 5388 896 5396 904
rect 4076 876 4084 884
rect 4204 876 4212 884
rect 4252 876 4260 884
rect 4444 876 4452 884
rect 4956 876 4964 884
rect 5260 876 5268 884
rect 2780 856 2788 864
rect 2860 856 2868 864
rect 492 836 500 844
rect 892 836 900 844
rect 3660 856 3668 864
rect 4012 856 4020 864
rect 4284 856 4292 864
rect 4300 856 4308 864
rect 4796 856 4804 864
rect 3100 836 3108 844
rect 3164 836 3172 844
rect 3516 836 3524 844
rect 4172 836 4180 844
rect 5132 836 5140 844
rect 5164 836 5172 844
rect 1068 816 1076 824
rect 1244 816 1252 824
rect 1260 816 1268 824
rect 1548 816 1556 824
rect 2268 816 2276 824
rect 3180 816 3188 824
rect 3388 816 3396 824
rect 4188 816 4196 824
rect 4588 816 4596 824
rect 4828 816 4836 824
rect 300 796 308 804
rect 1228 796 1236 804
rect 2156 796 2164 804
rect 2460 796 2468 804
rect 2492 796 2500 804
rect 1964 776 1972 784
rect 2476 776 2484 784
rect 2556 776 2564 784
rect 1564 756 1572 764
rect 1628 756 1636 764
rect 1708 756 1716 764
rect 2268 756 2276 764
rect 2940 776 2948 784
rect 3084 776 3092 784
rect 3212 776 3220 784
rect 2620 756 2628 764
rect 2892 756 2900 764
rect 3644 756 3652 764
rect 3660 756 3668 764
rect 3932 756 3940 764
rect 4044 756 4052 764
rect 828 736 836 744
rect 844 736 852 744
rect 2140 736 2148 744
rect 2364 736 2372 744
rect 2444 736 2452 744
rect 2892 736 2900 744
rect 3084 736 3092 744
rect 332 716 340 724
rect 428 716 436 724
rect 476 716 484 724
rect 780 716 788 724
rect 812 716 820 724
rect 1164 716 1172 724
rect 1228 716 1236 724
rect 1276 716 1284 724
rect 1292 716 1300 724
rect 1452 716 1460 724
rect 3036 716 3044 724
rect 4844 776 4852 784
rect 4188 756 4196 764
rect 4540 756 4548 764
rect 5036 756 5044 764
rect 5052 756 5060 764
rect 5116 756 5124 764
rect 4188 736 4196 744
rect 4268 736 4276 744
rect 4284 736 4292 744
rect 4556 736 4564 744
rect 4748 736 4756 744
rect 4764 736 4772 744
rect 4796 736 4804 744
rect 5068 736 5076 744
rect 3708 716 3716 724
rect 3820 716 3828 724
rect 4380 716 4388 724
rect 4508 716 4516 724
rect 4860 716 4868 724
rect 5068 716 5076 724
rect 5116 716 5124 724
rect 5260 716 5268 724
rect 204 696 212 704
rect 252 696 260 704
rect 1724 696 1732 704
rect 2108 696 2116 704
rect 2124 696 2132 704
rect 2524 696 2532 704
rect 2860 696 2868 704
rect 3468 696 3476 704
rect 4268 696 4276 704
rect 4316 696 4324 704
rect 4348 696 4356 704
rect 4492 696 4500 704
rect 4844 696 4852 704
rect 4860 696 4868 704
rect 4940 696 4948 704
rect 5036 696 5044 704
rect 5244 696 5252 704
rect 5276 696 5284 704
rect 5388 696 5396 704
rect 380 676 388 684
rect 796 676 804 684
rect 972 676 980 684
rect 1036 676 1044 684
rect 1148 676 1156 684
rect 1164 676 1172 684
rect 1212 676 1220 684
rect 1420 676 1428 684
rect 2428 676 2436 684
rect 2604 676 2612 684
rect 3068 676 3076 684
rect 3244 676 3252 684
rect 3276 676 3284 684
rect 3724 676 3732 684
rect 3788 676 3796 684
rect 3804 676 3812 684
rect 3836 676 3844 684
rect 3868 676 3876 684
rect 3948 676 3956 684
rect 4892 676 4900 684
rect 5292 676 5300 684
rect 5372 676 5380 684
rect 60 656 68 664
rect 1084 656 1092 664
rect 1564 656 1572 664
rect 1596 656 1604 664
rect 1612 656 1620 664
rect 2508 656 2516 664
rect 3068 656 3076 664
rect 3276 656 3284 664
rect 3468 656 3476 664
rect 3628 656 3636 664
rect 3980 656 3988 664
rect 4044 656 4052 664
rect 4140 656 4148 664
rect 5100 656 5108 664
rect 332 636 340 644
rect 3132 636 3140 644
rect 3324 636 3332 644
rect 3804 636 3812 644
rect 4092 636 4100 644
rect 4124 636 4132 644
rect 5148 636 5156 644
rect 316 616 324 624
rect 892 616 900 624
rect 908 616 916 624
rect 1500 616 1508 624
rect 2476 616 2484 624
rect 2716 616 2724 624
rect 3084 616 3092 624
rect 3148 616 3156 624
rect 3356 616 3364 624
rect 3516 616 3524 624
rect 3836 616 3844 624
rect 3916 616 3924 624
rect 4156 616 4164 624
rect 4444 616 4452 624
rect 5132 616 5140 624
rect 524 596 532 604
rect 604 596 612 604
rect 636 596 644 604
rect 2220 596 2228 604
rect 2380 596 2388 604
rect 3084 596 3092 604
rect 3756 596 3764 604
rect 3852 596 3860 604
rect 3980 596 3988 604
rect 3996 596 4004 604
rect 4220 596 4228 604
rect 4620 596 4628 604
rect 4668 596 4676 604
rect 4972 596 4980 604
rect 5004 596 5012 604
rect 5052 596 5060 604
rect 5068 596 5076 604
rect 1004 576 1012 584
rect 1116 576 1124 584
rect 1484 576 1492 584
rect 1532 576 1540 584
rect 1628 576 1636 584
rect 2428 576 2436 584
rect 2444 576 2452 584
rect 2524 576 2532 584
rect 2556 576 2564 584
rect 2652 576 2660 584
rect 3164 576 3172 584
rect 3308 576 3316 584
rect 3452 576 3460 584
rect 4188 576 4196 584
rect 4204 576 4212 584
rect 4380 576 4388 584
rect 4588 576 4596 584
rect 4988 576 4996 584
rect 556 556 564 564
rect 588 556 596 564
rect 1676 556 1684 564
rect 1740 556 1748 564
rect 1980 556 1988 564
rect 2348 556 2356 564
rect 2636 556 2644 564
rect 2892 556 2900 564
rect 3452 556 3460 564
rect 4012 556 4020 564
rect 4444 556 4452 564
rect 4476 556 4484 564
rect 4876 556 4884 564
rect 4892 556 4900 564
rect 5308 556 5316 564
rect 5388 556 5396 564
rect 252 536 260 544
rect 332 536 340 544
rect 428 536 436 544
rect 844 536 852 544
rect 1132 536 1140 544
rect 2124 536 2132 544
rect 2812 536 2820 544
rect 2892 536 2900 544
rect 2956 536 2964 544
rect 3484 536 3492 544
rect 3500 536 3508 544
rect 3660 536 3668 544
rect 5276 536 5284 544
rect 5324 536 5332 544
rect 524 516 532 524
rect 636 516 644 524
rect 956 516 964 524
rect 1580 516 1588 524
rect 1628 516 1636 524
rect 1948 516 1956 524
rect 2620 516 2628 524
rect 2636 516 2644 524
rect 2844 516 2852 524
rect 220 496 228 504
rect 2028 496 2036 504
rect 2124 496 2132 504
rect 2348 496 2356 504
rect 2620 496 2628 504
rect 2684 496 2692 504
rect 3420 516 3428 524
rect 4284 496 4292 504
rect 4316 496 4324 504
rect 4332 496 4340 504
rect 5004 496 5012 504
rect 5436 496 5444 504
rect 5452 496 5460 504
rect 364 476 372 484
rect 1772 476 1780 484
rect 1804 476 1812 484
rect 2508 476 2516 484
rect 3404 476 3412 484
rect 3532 476 3540 484
rect 3788 476 3796 484
rect 4220 476 4228 484
rect 3132 456 3140 464
rect 3260 456 3268 464
rect 3452 456 3460 464
rect 4140 456 4148 464
rect 2892 436 2900 444
rect 4268 436 4276 444
rect 5308 436 5316 444
rect 1084 416 1092 424
rect 1820 416 1828 424
rect 2460 416 2468 424
rect 3404 416 3412 424
rect 2972 396 2980 404
rect 4220 396 4228 404
rect 1548 376 1556 384
rect 3068 376 3076 384
rect 3516 376 3524 384
rect 3596 376 3604 384
rect 3900 376 3908 384
rect 4364 376 4372 384
rect 4476 376 4484 384
rect 5164 376 5172 384
rect 396 356 404 364
rect 572 356 580 364
rect 1292 356 1300 364
rect 1532 356 1540 364
rect 1836 356 1844 364
rect 2540 356 2548 364
rect 4348 356 4356 364
rect 92 336 100 344
rect 716 336 724 344
rect 1324 336 1332 344
rect 1484 336 1492 344
rect 2412 336 2420 344
rect 2860 336 2868 344
rect 3260 336 3268 344
rect 3916 336 3924 344
rect 4364 336 4372 344
rect 4972 336 4980 344
rect 5036 336 5044 344
rect 380 316 388 324
rect 508 316 516 324
rect 1020 316 1028 324
rect 1388 316 1396 324
rect 2204 316 2212 324
rect 2268 316 2276 324
rect 2476 316 2484 324
rect 2508 316 2516 324
rect 2748 316 2756 324
rect 2844 316 2852 324
rect 3788 316 3796 324
rect 3836 316 3844 324
rect 3868 316 3876 324
rect 3916 316 3924 324
rect 4492 316 4500 324
rect 4716 316 4724 324
rect 4844 316 4852 324
rect 5276 316 5284 324
rect 5324 316 5332 324
rect 988 296 996 304
rect 1020 296 1028 304
rect 1916 296 1924 304
rect 2828 296 2836 304
rect 3532 296 3540 304
rect 3724 296 3732 304
rect 3804 296 3812 304
rect 3964 296 3972 304
rect 4060 296 4068 304
rect 4092 296 4100 304
rect 4396 296 4404 304
rect 4508 296 4516 304
rect 4844 296 4852 304
rect 5020 296 5028 304
rect 5244 296 5252 304
rect 5292 296 5300 304
rect 60 276 68 284
rect 204 276 212 284
rect 300 276 308 284
rect 588 276 596 284
rect 684 276 692 284
rect 796 276 804 284
rect 1212 276 1220 284
rect 1404 276 1412 284
rect 1804 276 1812 284
rect 1932 276 1940 284
rect 2044 276 2052 284
rect 2108 276 2116 284
rect 2236 276 2244 284
rect 2428 276 2436 284
rect 2572 276 2580 284
rect 2700 276 2708 284
rect 2908 276 2916 284
rect 3068 276 3076 284
rect 4108 276 4116 284
rect 4236 276 4244 284
rect 4268 276 4276 284
rect 5356 276 5364 284
rect 1628 256 1636 264
rect 1724 256 1732 264
rect 2652 256 2660 264
rect 2876 256 2884 264
rect 2972 256 2980 264
rect 3244 256 3252 264
rect 4876 256 4884 264
rect 5244 256 5252 264
rect 396 236 404 244
rect 956 236 964 244
rect 1484 236 1492 244
rect 1708 236 1716 244
rect 1916 236 1924 244
rect 2860 236 2868 244
rect 2892 236 2900 244
rect 3132 236 3140 244
rect 3564 236 3572 244
rect 4236 236 4244 244
rect 4252 236 4260 244
rect 748 216 756 224
rect 1020 216 1028 224
rect 1052 216 1060 224
rect 3276 216 3284 224
rect 3324 216 3332 224
rect 3628 216 3636 224
rect 4828 216 4836 224
rect 4924 216 4932 224
rect 5084 216 5092 224
rect 5180 216 5188 224
rect 5228 216 5236 224
rect 316 196 324 204
rect 956 196 964 204
rect 1452 196 1460 204
rect 1820 196 1828 204
rect 1980 196 1988 204
rect 2300 196 2308 204
rect 2972 196 2980 204
rect 3452 196 3460 204
rect 3516 196 3524 204
rect 5148 196 5156 204
rect 5244 196 5252 204
rect 5468 196 5476 204
rect 28 176 36 184
rect 428 176 436 184
rect 508 176 516 184
rect 604 176 612 184
rect 700 176 708 184
rect 2460 176 2468 184
rect 2572 176 2580 184
rect 2892 176 2900 184
rect 2940 176 2948 184
rect 3100 176 3108 184
rect 3692 176 3700 184
rect 3756 176 3764 184
rect 3772 176 3780 184
rect 4092 176 4100 184
rect 4156 176 4164 184
rect 4684 176 4692 184
rect 5196 176 5204 184
rect 5244 176 5252 184
rect 60 156 68 164
rect 76 156 84 164
rect 316 156 324 164
rect 876 156 884 164
rect 1100 156 1108 164
rect 2492 156 2500 164
rect 2956 156 2964 164
rect 3244 156 3252 164
rect 3308 156 3316 164
rect 3324 156 3332 164
rect 3948 156 3956 164
rect 3980 156 3988 164
rect 4140 156 4148 164
rect 4220 156 4228 164
rect 5036 156 5044 164
rect 5292 156 5300 164
rect 5340 156 5348 164
rect 92 136 100 144
rect 220 136 228 144
rect 236 136 244 144
rect 988 136 996 144
rect 1132 136 1140 144
rect 1164 136 1172 144
rect 1180 136 1188 144
rect 1212 136 1220 144
rect 1228 136 1236 144
rect 1308 136 1316 144
rect 1724 136 1732 144
rect 1756 136 1764 144
rect 1948 136 1956 144
rect 2652 136 2660 144
rect 2828 136 2836 144
rect 3468 136 3476 144
rect 4460 136 4468 144
rect 5260 136 5268 144
rect 5436 136 5444 144
rect 412 116 420 124
rect 572 116 580 124
rect 684 116 692 124
rect 700 116 708 124
rect 812 116 820 124
rect 988 116 996 124
rect 2428 116 2436 124
rect 2876 116 2884 124
rect 3276 116 3284 124
rect 4380 116 4388 124
rect 4540 116 4548 124
rect 4588 116 4596 124
rect 4604 116 4612 124
rect 4684 116 4692 124
rect 556 96 564 104
rect 636 96 644 104
rect 1148 96 1156 104
rect 1164 96 1172 104
rect 1356 96 1364 104
rect 1372 96 1380 104
rect 1404 96 1412 104
rect 1564 96 1572 104
rect 1580 96 1588 104
rect 1724 96 1732 104
rect 2124 96 2132 104
rect 2332 96 2340 104
rect 2348 96 2356 104
rect 3116 96 3124 104
rect 3980 96 3988 104
rect 4300 96 4308 104
rect 4524 96 4532 104
rect 4556 96 4564 104
rect 4780 96 4788 104
rect 1436 76 1444 84
rect 1452 76 1460 84
rect 1804 76 1812 84
rect 3996 76 4004 84
rect 5324 76 5332 84
rect 1708 56 1716 64
rect 1740 56 1748 64
rect 2252 56 2260 64
rect 3852 56 3860 64
rect 5420 56 5428 64
rect 4652 36 4660 44
rect 2956 16 2964 24
rect 4684 16 4692 24
<< metal4 >>
rect 253 3904 259 3956
rect 253 3764 259 3896
rect 13 2904 19 3736
rect 77 3704 83 3756
rect 285 3684 291 3716
rect 13 2124 19 2896
rect 29 2684 35 2956
rect 61 1804 67 3336
rect 77 2564 83 3196
rect 93 3084 99 3096
rect 125 3084 131 3096
rect 116 2977 124 2983
rect 141 2684 147 3376
rect 189 3344 195 3476
rect 205 3364 211 3476
rect 173 3064 179 3116
rect 61 1724 67 1756
rect 77 1464 83 2256
rect 109 1884 115 2576
rect 125 2544 131 2556
rect 141 2284 147 2676
rect 141 1624 147 1856
rect 189 1624 195 3316
rect 205 2604 211 3056
rect 237 1884 243 3096
rect 253 3064 259 3076
rect 285 2944 291 3676
rect 301 3304 307 3696
rect 317 3344 323 3376
rect 365 3104 371 3376
rect 397 3144 403 3496
rect 413 3264 419 3836
rect 301 3024 307 3056
rect 260 2897 268 2903
rect 253 2544 259 2636
rect 269 2624 275 2716
rect 125 1304 131 1356
rect 45 1084 51 1216
rect 61 664 67 1156
rect 125 1064 131 1116
rect 173 1084 179 1456
rect 189 1404 195 1476
rect 173 1064 179 1076
rect 125 924 131 956
rect 189 944 195 1096
rect 205 1064 211 1876
rect 20 177 28 183
rect 61 164 67 276
rect 77 164 83 176
rect 93 144 99 336
rect 205 284 211 696
rect 221 504 227 1676
rect 253 1324 259 2396
rect 269 1744 275 2616
rect 285 2344 291 2936
rect 317 1784 323 2576
rect 269 964 275 1176
rect 285 1064 291 1076
rect 237 144 243 936
rect 253 544 259 696
rect 285 344 291 1036
rect 301 804 307 1056
rect 317 624 323 1716
rect 333 724 339 3036
rect 349 2564 355 3056
rect 349 2124 355 2136
rect 349 1924 355 2096
rect 349 904 355 1916
rect 365 1864 371 2896
rect 381 2884 387 2956
rect 381 1884 387 2616
rect 397 2504 403 2556
rect 397 2104 403 2136
rect 381 1524 387 1876
rect 333 544 339 636
rect 365 484 371 1076
rect 397 984 403 1856
rect 413 1124 419 2396
rect 429 1964 435 3836
rect 701 3784 707 3836
rect 525 3744 531 3776
rect 468 3537 476 3543
rect 509 3104 515 3736
rect 548 3717 556 3723
rect 525 3124 531 3696
rect 637 3524 643 3716
rect 717 3504 723 3716
rect 541 3104 547 3116
rect 445 2904 451 3056
rect 573 3024 579 3036
rect 445 2484 451 2876
rect 461 2564 467 3016
rect 589 2964 595 3496
rect 532 2937 540 2943
rect 573 2684 579 2696
rect 589 2684 595 2956
rect 605 2704 611 3256
rect 637 3184 643 3376
rect 621 2884 627 3136
rect 637 3044 643 3156
rect 509 2624 515 2656
rect 445 2124 451 2136
rect 493 1924 499 2556
rect 381 704 387 976
rect 397 944 403 956
rect 429 724 435 1756
rect 445 1124 451 1736
rect 461 1364 467 1816
rect 509 1744 515 2596
rect 525 1764 531 2656
rect 541 2584 547 2636
rect 637 2564 643 2756
rect 653 2724 659 3336
rect 749 3104 755 3836
rect 765 3744 771 3876
rect 781 3784 787 3796
rect 813 3764 819 3876
rect 813 3544 819 3696
rect 829 3684 835 3776
rect 765 3524 771 3536
rect 813 3524 819 3536
rect 765 3324 771 3356
rect 765 3044 771 3076
rect 733 2684 739 2696
rect 676 2677 684 2683
rect 493 1684 499 1696
rect 461 1064 467 1316
rect 477 724 483 1456
rect 493 844 499 1596
rect 541 1344 547 2136
rect 557 1704 563 2336
rect 621 2144 627 2176
rect 580 1837 588 1843
rect 605 1724 611 1836
rect 573 1464 579 1496
rect 525 1324 531 1336
rect 541 1104 547 1136
rect 381 324 387 676
rect 429 544 435 716
rect 397 244 403 356
rect 317 164 323 196
rect 429 184 435 536
rect 509 324 515 876
rect 525 524 531 596
rect 557 564 563 976
rect 589 564 595 1336
rect 605 624 611 1496
rect 621 1364 627 1856
rect 637 1544 643 2216
rect 653 2144 659 2676
rect 685 2304 691 2316
rect 669 1764 675 1856
rect 717 1844 723 2516
rect 749 2324 755 2936
rect 733 2124 739 2136
rect 749 2104 755 2316
rect 765 2144 771 2956
rect 781 2544 787 2556
rect 749 2064 755 2076
rect 765 1924 771 1956
rect 749 1857 764 1863
rect 749 1844 755 1857
rect 692 1837 700 1843
rect 653 1424 659 1456
rect 637 1344 643 1356
rect 733 1304 739 1356
rect 621 1144 627 1296
rect 621 1084 627 1136
rect 637 1024 643 1056
rect 717 1024 723 1056
rect 692 1017 700 1023
rect 573 344 579 356
rect 589 284 595 556
rect 509 184 515 256
rect 605 184 611 596
rect 637 524 643 596
rect 717 304 723 336
rect 685 284 691 296
rect 749 224 755 1536
rect 781 1464 787 2116
rect 797 1764 803 3116
rect 813 2304 819 3516
rect 829 3504 835 3516
rect 829 2984 835 3156
rect 845 2744 851 3876
rect 861 3704 867 3736
rect 957 3724 963 3796
rect 973 3784 979 3856
rect 909 3504 915 3716
rect 884 3437 899 3443
rect 893 3424 899 3437
rect 909 3304 915 3496
rect 957 3444 963 3456
rect 861 3104 867 3116
rect 861 2684 867 2796
rect 829 2244 835 2576
rect 813 1764 819 1956
rect 829 1484 835 2096
rect 845 2004 851 2016
rect 845 1944 851 1976
rect 861 1904 867 2656
rect 877 1944 883 3296
rect 941 3264 947 3316
rect 941 3144 947 3256
rect 925 2924 931 2936
rect 925 2744 931 2756
rect 893 2144 899 2156
rect 884 1897 892 1903
rect 797 1004 803 1356
rect 813 1104 819 1336
rect 829 1104 835 1476
rect 845 1304 851 1756
rect 861 1524 867 1536
rect 813 964 819 1016
rect 829 944 835 1096
rect 861 1064 867 1336
rect 845 1044 851 1056
rect 845 744 851 1016
rect 861 1004 867 1056
rect 893 884 899 936
rect 804 717 812 723
rect 781 703 787 716
rect 781 697 803 703
rect 797 684 803 697
rect 845 544 851 736
rect 893 624 899 836
rect 909 624 915 2696
rect 925 2644 931 2716
rect 925 2284 931 2496
rect 941 2284 947 3136
rect 957 2304 963 3436
rect 1005 3404 1011 3436
rect 1021 3404 1027 3756
rect 1037 3324 1043 3416
rect 1053 3384 1059 3496
rect 973 2524 979 2936
rect 989 2684 995 2976
rect 1005 2684 1011 2916
rect 1021 2744 1027 3316
rect 1037 3084 1043 3096
rect 989 2344 995 2676
rect 973 2304 979 2316
rect 925 1704 931 2276
rect 941 2084 947 2276
rect 973 2164 979 2176
rect 957 1904 963 1916
rect 989 1904 995 2256
rect 925 1304 931 1676
rect 941 1484 947 1776
rect 957 1704 963 1796
rect 989 1724 995 1736
rect 964 1457 972 1463
rect 989 1384 995 1716
rect 1005 1544 1011 2636
rect 1021 2104 1027 2736
rect 1037 2264 1043 2996
rect 1053 2704 1059 3376
rect 1069 3004 1075 3896
rect 1085 3784 1091 3796
rect 1085 3364 1091 3736
rect 1213 3704 1219 3876
rect 1284 3737 1292 3743
rect 1085 3217 1091 3236
rect 1085 3024 1091 3196
rect 1108 3097 1116 3103
rect 1140 3057 1148 3063
rect 1181 3044 1187 3676
rect 1197 3104 1203 3616
rect 1213 3544 1219 3696
rect 1229 3144 1235 3156
rect 1213 3044 1219 3096
rect 1165 3024 1171 3036
rect 1085 2904 1091 2916
rect 1101 2704 1107 2716
rect 1053 2644 1059 2656
rect 1053 2544 1059 2556
rect 1085 2184 1091 2516
rect 1117 2204 1123 2976
rect 1149 2884 1155 2916
rect 1037 2164 1043 2176
rect 1037 1784 1043 1836
rect 941 1044 947 1056
rect 957 524 963 1196
rect 973 804 979 996
rect 973 684 979 776
rect 989 304 995 1056
rect 1005 904 1011 976
rect 1021 944 1027 1536
rect 1037 1384 1043 1396
rect 1053 1144 1059 1936
rect 1069 1424 1075 1836
rect 1085 1204 1091 2116
rect 1117 1704 1123 2156
rect 1133 2104 1139 2696
rect 1165 2344 1171 2496
rect 1165 2244 1171 2276
rect 1133 2084 1139 2096
rect 1149 2084 1155 2116
rect 1181 2084 1187 3036
rect 1197 2924 1203 2936
rect 1197 2784 1203 2796
rect 1213 2584 1219 3036
rect 1229 2584 1235 2996
rect 1245 2964 1251 3676
rect 1261 3104 1267 3136
rect 1277 2984 1283 3416
rect 1293 3384 1299 3396
rect 1293 2964 1299 3056
rect 1309 2984 1315 3896
rect 1405 3764 1411 3876
rect 1469 3784 1475 3796
rect 1325 3664 1331 3676
rect 1341 3484 1347 3736
rect 1485 3704 1491 3956
rect 2685 3924 2691 3956
rect 3949 3924 3955 3936
rect 3268 3917 3276 3923
rect 4708 3917 4716 3923
rect 1501 3764 1507 3796
rect 1517 3704 1523 3736
rect 1325 3104 1331 3136
rect 1309 2964 1315 2976
rect 1245 2664 1251 2936
rect 1261 2664 1267 2696
rect 1229 2284 1235 2556
rect 1229 2244 1235 2276
rect 1133 1864 1139 2016
rect 1181 1944 1187 2076
rect 1149 1704 1155 1776
rect 1197 1704 1203 2136
rect 1037 684 1043 996
rect 1053 924 1059 936
rect 1085 664 1091 1196
rect 1005 584 1011 616
rect 1021 304 1027 316
rect 804 277 812 283
rect 964 237 972 243
rect 957 184 963 196
rect 708 177 716 183
rect 868 157 876 163
rect 989 144 995 296
rect 1021 224 1027 296
rect 1085 284 1091 416
rect 1053 224 1059 256
rect 1101 164 1107 1476
rect 1133 1324 1139 1656
rect 1117 1204 1123 1216
rect 1117 684 1123 1036
rect 1117 564 1123 576
rect 1133 544 1139 1316
rect 1149 704 1155 1496
rect 1181 1384 1187 1636
rect 1197 1524 1203 1696
rect 1213 1484 1219 1896
rect 1245 1724 1251 2656
rect 1261 2104 1267 2636
rect 1277 2304 1283 2956
rect 1181 1344 1187 1356
rect 1165 1324 1171 1336
rect 1165 1144 1171 1236
rect 1197 1124 1203 1336
rect 1213 1324 1219 1476
rect 1229 1084 1235 1536
rect 1261 1444 1267 1916
rect 1277 1844 1283 2296
rect 1293 2184 1299 2896
rect 1309 2324 1315 2916
rect 1325 2684 1331 2696
rect 1341 2684 1347 3476
rect 1325 2584 1331 2636
rect 1341 2624 1347 2636
rect 1325 2504 1331 2536
rect 1309 2204 1315 2276
rect 1341 2104 1347 2116
rect 1325 2084 1331 2096
rect 1277 1804 1283 1836
rect 1325 1464 1331 1476
rect 1309 1364 1315 1456
rect 1341 1404 1347 2076
rect 1357 1504 1363 2936
rect 1373 2664 1379 3696
rect 1453 3544 1459 3696
rect 1373 2564 1379 2576
rect 1389 2544 1395 3516
rect 1421 3104 1427 3376
rect 1453 3124 1459 3536
rect 1485 3364 1491 3696
rect 1485 3144 1491 3356
rect 1517 3144 1523 3696
rect 1565 3364 1571 3796
rect 1613 3784 1619 3796
rect 1661 3784 1667 3796
rect 1677 3504 1683 3756
rect 1837 3704 1843 3716
rect 1917 3704 1923 3916
rect 1940 3777 1948 3783
rect 2029 3644 2035 3816
rect 2189 3784 2195 3856
rect 2189 3664 2195 3776
rect 2276 3697 2284 3703
rect 1460 3097 1468 3103
rect 1533 3064 1539 3296
rect 1549 3204 1555 3356
rect 1565 3344 1571 3356
rect 1549 2784 1555 3196
rect 1565 3124 1571 3336
rect 1613 3324 1619 3396
rect 1581 3044 1587 3116
rect 1597 3084 1603 3216
rect 1453 2704 1459 2716
rect 1405 2684 1411 2696
rect 1373 1743 1379 2416
rect 1389 2124 1395 2536
rect 1405 2284 1411 2556
rect 1421 2544 1427 2596
rect 1421 2344 1427 2496
rect 1405 2124 1411 2156
rect 1421 1884 1427 2256
rect 1396 1817 1411 1823
rect 1437 1763 1443 2636
rect 1453 2084 1459 2696
rect 1549 2684 1555 2696
rect 1469 2144 1475 2676
rect 1517 2604 1523 2676
rect 1485 2504 1491 2536
rect 1485 2104 1491 2296
rect 1421 1757 1443 1763
rect 1373 1737 1395 1743
rect 1341 1324 1347 1356
rect 1341 1284 1347 1296
rect 1284 1137 1292 1143
rect 1309 1084 1315 1096
rect 1284 1077 1292 1083
rect 1325 944 1331 1036
rect 1252 917 1260 923
rect 1165 724 1171 816
rect 1149 684 1155 696
rect 1213 684 1219 916
rect 1229 724 1235 796
rect 1245 784 1251 816
rect 1357 724 1363 1496
rect 1373 1344 1379 1716
rect 1389 1564 1395 1737
rect 1389 1484 1395 1536
rect 1389 1244 1395 1416
rect 1405 1364 1411 1676
rect 1421 1384 1427 1757
rect 1389 1144 1395 1216
rect 1389 1104 1395 1116
rect 1373 1044 1379 1076
rect 1389 964 1395 1096
rect 1277 704 1283 716
rect 1124 537 1132 543
rect 1124 137 1132 143
rect 685 124 691 136
rect 989 124 995 136
rect 420 117 428 123
rect 557 117 572 123
rect 557 104 563 117
rect 804 117 812 123
rect 637 104 643 116
rect 1149 104 1155 676
rect 1165 664 1171 676
rect 1213 284 1219 676
rect 1293 364 1299 716
rect 1325 284 1331 336
rect 1380 317 1388 323
rect 1405 284 1411 1356
rect 1421 684 1427 1336
rect 1437 1084 1443 1736
rect 1453 1524 1459 2076
rect 1469 1864 1475 1876
rect 1469 1764 1475 1776
rect 1453 1284 1459 1516
rect 1453 724 1459 1276
rect 1469 1064 1475 1656
rect 1485 1464 1491 2096
rect 1501 1884 1507 2316
rect 1533 2164 1539 2196
rect 1485 1324 1491 1376
rect 1469 964 1475 996
rect 1485 964 1491 1076
rect 1501 984 1507 1456
rect 1524 1417 1539 1423
rect 1533 1364 1539 1396
rect 1549 1044 1555 2676
rect 1581 2544 1587 3036
rect 1597 2964 1603 3076
rect 1645 2984 1651 3116
rect 1565 2164 1571 2196
rect 1581 2164 1587 2536
rect 1565 1804 1571 1996
rect 1501 944 1507 976
rect 1533 904 1539 996
rect 1549 944 1555 1036
rect 1485 584 1491 776
rect 1533 584 1539 596
rect 1549 384 1555 816
rect 1565 764 1571 1776
rect 1581 1744 1587 2156
rect 1597 1584 1603 2676
rect 1613 2144 1619 2156
rect 1581 964 1587 1416
rect 1597 1344 1603 1556
rect 1613 1544 1619 1956
rect 1629 1544 1635 2756
rect 1645 2684 1651 2696
rect 1661 1504 1667 3096
rect 1693 2724 1699 3536
rect 1709 3444 1715 3536
rect 1709 3364 1715 3436
rect 1741 3324 1747 3396
rect 1716 3297 1724 3303
rect 1709 2924 1715 3196
rect 1725 3184 1731 3196
rect 1677 2284 1683 2356
rect 1677 2244 1683 2256
rect 1693 2204 1699 2316
rect 1709 2224 1715 2436
rect 1725 2244 1731 2256
rect 1693 2144 1699 2176
rect 1741 2144 1747 3316
rect 1773 3044 1779 3136
rect 1789 3124 1795 3496
rect 1805 3184 1811 3396
rect 1821 3084 1827 3496
rect 1837 3084 1843 3336
rect 1757 2364 1763 2716
rect 1773 2524 1779 3036
rect 1789 2744 1795 3076
rect 1805 2764 1811 2796
rect 1716 2137 1724 2143
rect 1741 2124 1747 2136
rect 1773 2124 1779 2516
rect 1789 2364 1795 2716
rect 1796 2277 1804 2283
rect 1677 2084 1683 2096
rect 1677 1784 1683 2036
rect 1677 1724 1683 1776
rect 1677 1584 1683 1656
rect 1677 1524 1683 1576
rect 1636 1497 1644 1503
rect 1613 1424 1619 1456
rect 1597 1144 1603 1156
rect 1613 1144 1619 1296
rect 1581 524 1587 936
rect 1597 664 1603 676
rect 1613 664 1619 1136
rect 1661 1084 1667 1496
rect 1693 1384 1699 2096
rect 1709 1744 1715 2096
rect 1741 1724 1747 2116
rect 1821 2044 1827 3076
rect 1837 2684 1843 3076
rect 1853 3064 1859 3096
rect 1869 2984 1875 2996
rect 1885 2924 1891 3276
rect 1917 3164 1923 3396
rect 1901 2984 1907 3056
rect 1677 1364 1683 1376
rect 1725 1124 1731 1716
rect 1757 1464 1763 1476
rect 1757 1124 1763 1136
rect 1668 897 1676 903
rect 1629 584 1635 756
rect 1709 724 1715 756
rect 1725 704 1731 1056
rect 1741 1024 1747 1116
rect 1741 964 1747 1016
rect 1677 564 1683 576
rect 1741 564 1747 596
rect 1629 504 1635 516
rect 1773 484 1779 1856
rect 1837 1644 1843 2676
rect 1853 2304 1859 2756
rect 1853 1784 1859 2296
rect 1869 1964 1875 2276
rect 1885 2144 1891 2916
rect 1901 2524 1907 2976
rect 1933 2923 1939 3436
rect 1965 3324 1971 3596
rect 1981 3424 1987 3576
rect 2029 3544 2035 3636
rect 1917 2917 1939 2923
rect 1917 2764 1923 2917
rect 1917 2704 1923 2736
rect 1933 2664 1939 2896
rect 1949 2704 1955 3236
rect 1981 2684 1987 3396
rect 1997 3164 2003 3176
rect 1956 2657 1964 2663
rect 1885 1884 1891 2136
rect 1901 1944 1907 2336
rect 1917 1944 1923 2636
rect 1933 2164 1939 2656
rect 1949 2324 1955 2336
rect 1965 2204 1971 2636
rect 1949 2124 1955 2176
rect 1981 2104 1987 2676
rect 1997 2664 2003 2936
rect 2013 2603 2019 3196
rect 2029 3064 2035 3076
rect 2061 3044 2067 3056
rect 2045 2744 2051 2796
rect 1997 2597 2019 2603
rect 1997 2384 2003 2597
rect 2029 2344 2035 2576
rect 1997 2284 2003 2336
rect 2013 2244 2019 2336
rect 2029 2284 2035 2336
rect 2045 2284 2051 2696
rect 1997 2224 2003 2236
rect 2013 2124 2019 2136
rect 1949 1904 1955 1916
rect 1981 1904 1987 2096
rect 2061 2084 2067 2536
rect 1869 1484 1875 1856
rect 1789 1184 1795 1396
rect 1805 1284 1811 1396
rect 1837 1204 1843 1396
rect 1805 1164 1811 1176
rect 1805 1044 1811 1116
rect 1309 144 1315 176
rect 1236 137 1244 143
rect 1181 124 1187 136
rect 1165 104 1171 116
rect 1213 104 1219 136
rect 1261 104 1267 136
rect 1373 104 1379 136
rect 1405 104 1411 256
rect 1485 244 1491 316
rect 1533 264 1539 356
rect 1805 284 1811 476
rect 1636 257 1644 263
rect 1725 244 1731 256
rect 1348 97 1356 103
rect 1437 84 1443 236
rect 1453 84 1459 196
rect 1565 104 1571 136
rect 1588 97 1596 103
rect 1709 64 1715 236
rect 1821 204 1827 416
rect 1837 364 1843 1076
rect 1853 964 1859 1196
rect 1885 1144 1891 1656
rect 1901 1304 1907 1676
rect 1949 1624 1955 1856
rect 1917 1163 1923 1616
rect 1901 1157 1923 1163
rect 1885 924 1891 1016
rect 1901 1004 1907 1157
rect 1917 304 1923 1136
rect 1933 544 1939 1296
rect 1949 1064 1955 1476
rect 1965 1124 1971 1416
rect 1949 984 1955 1016
rect 1965 784 1971 996
rect 1981 564 1987 1636
rect 1917 244 1923 296
rect 1933 284 1939 536
rect 1949 524 1955 536
rect 1997 323 2003 1996
rect 2061 1764 2067 2076
rect 2077 1744 2083 2516
rect 2093 2324 2099 3376
rect 2109 2984 2115 3396
rect 2109 2564 2115 2976
rect 2125 2944 2131 3596
rect 2157 3544 2163 3556
rect 2269 3464 2275 3516
rect 2301 3464 2307 3856
rect 2141 2944 2147 3456
rect 2237 3104 2243 3396
rect 2269 3344 2275 3376
rect 2317 3344 2323 3736
rect 2333 3704 2339 3916
rect 2493 3884 2499 3916
rect 3732 3897 3740 3903
rect 2749 3864 2755 3876
rect 2797 3864 2803 3896
rect 2797 3844 2803 3856
rect 2589 3764 2595 3796
rect 2349 3704 2355 3736
rect 2621 3584 2627 3796
rect 2797 3724 2803 3756
rect 2109 2004 2115 2396
rect 2125 2324 2131 2356
rect 2141 2264 2147 2936
rect 2180 2677 2188 2683
rect 2093 1824 2099 1956
rect 2125 1844 2131 1856
rect 2029 1504 2035 1516
rect 2045 1484 2051 1536
rect 2109 1404 2115 1836
rect 2125 1804 2131 1816
rect 2020 497 2028 503
rect 1981 317 2003 323
rect 1981 204 1987 317
rect 2045 284 2051 1136
rect 2109 984 2115 1396
rect 2125 704 2131 1456
rect 2141 744 2147 2256
rect 2157 2244 2163 2276
rect 2221 2264 2227 3056
rect 2237 2684 2243 3096
rect 2285 2924 2291 2936
rect 2253 2684 2259 2716
rect 2221 2144 2227 2156
rect 2237 2004 2243 2676
rect 2260 2577 2268 2583
rect 2285 2164 2291 2836
rect 2301 2144 2307 2956
rect 2317 2544 2323 3336
rect 2333 2184 2339 3216
rect 2381 3104 2387 3496
rect 2477 3124 2483 3416
rect 2397 3084 2403 3096
rect 2356 2937 2364 2943
rect 2381 2403 2387 2796
rect 2573 2744 2579 3356
rect 2605 3324 2611 3356
rect 2621 3344 2627 3356
rect 2637 3344 2643 3376
rect 2468 2717 2476 2723
rect 2445 2684 2451 2716
rect 2413 2524 2419 2536
rect 2365 2397 2387 2403
rect 2157 1784 2163 1956
rect 2173 1484 2179 1856
rect 2189 1824 2195 1956
rect 2157 1284 2163 1416
rect 2237 1344 2243 1996
rect 2285 1924 2291 2136
rect 2253 1424 2259 1896
rect 2340 1857 2348 1863
rect 2301 1844 2307 1856
rect 2269 1784 2275 1796
rect 2285 1744 2291 1756
rect 2189 944 2195 1056
rect 2205 964 2211 996
rect 2100 697 2108 703
rect 2125 684 2131 696
rect 2125 544 2131 676
rect 2141 664 2147 736
rect 2221 604 2227 936
rect 2125 324 2131 496
rect 2205 324 2211 476
rect 2237 284 2243 1336
rect 2269 1084 2275 1736
rect 2269 824 2275 1076
rect 2285 1064 2291 1716
rect 2301 1344 2307 1476
rect 2317 1204 2323 1756
rect 2333 1724 2339 1736
rect 2365 1684 2371 2397
rect 2429 2164 2435 2536
rect 2445 2184 2451 2516
rect 2509 2244 2515 2276
rect 2429 1804 2435 2116
rect 2388 1757 2396 1763
rect 2413 1743 2419 1776
rect 2397 1737 2419 1743
rect 2333 1304 2339 1316
rect 2285 884 2291 1056
rect 2269 324 2275 756
rect 2269 304 2275 316
rect 2116 277 2124 283
rect 2301 204 2307 1136
rect 2333 944 2339 956
rect 2349 564 2355 1316
rect 2365 984 2371 1676
rect 2397 1464 2403 1737
rect 2429 1724 2435 1796
rect 2413 1104 2419 1356
rect 2365 744 2371 976
rect 2397 924 2403 1076
rect 2413 944 2419 1096
rect 2429 1064 2435 1596
rect 2445 1084 2451 2136
rect 2493 2044 2499 2236
rect 2461 1924 2467 1956
rect 2477 1764 2483 1916
rect 2445 1004 2451 1056
rect 2381 564 2387 596
rect 2349 504 2355 556
rect 2413 344 2419 936
rect 2429 684 2435 896
rect 2461 804 2467 1716
rect 2477 964 2483 1756
rect 2493 1304 2499 2036
rect 2509 1364 2515 1876
rect 2541 1763 2547 1856
rect 2557 1804 2563 2056
rect 2573 1824 2579 2736
rect 2605 2144 2611 2796
rect 2621 2684 2627 3336
rect 2669 2783 2675 3336
rect 2685 2944 2691 3636
rect 2804 3337 2812 3343
rect 2669 2777 2691 2783
rect 2589 2124 2595 2136
rect 2621 2104 2627 2496
rect 2637 2284 2643 2296
rect 2605 2064 2611 2076
rect 2621 1944 2627 2096
rect 2525 1757 2547 1763
rect 2493 1024 2499 1036
rect 2477 784 2483 956
rect 2429 584 2435 676
rect 2445 664 2451 736
rect 2445 564 2451 576
rect 1748 137 1756 143
rect 1725 104 1731 136
rect 1741 64 1747 116
rect 1805 84 1811 156
rect 2333 104 2339 136
rect 2429 124 2435 276
rect 2461 184 2467 416
rect 2477 324 2483 616
rect 2493 164 2499 796
rect 2509 664 2515 1356
rect 2525 1184 2531 1757
rect 2589 1743 2595 1896
rect 2573 1737 2595 1743
rect 2573 1724 2579 1737
rect 2541 1124 2547 1636
rect 2605 1284 2611 1756
rect 2637 1344 2643 2076
rect 2653 1604 2659 2676
rect 2669 2244 2675 2756
rect 2685 2344 2691 2777
rect 2701 2704 2707 3336
rect 2845 3284 2851 3516
rect 2861 3264 2867 3876
rect 2909 3704 2915 3756
rect 2925 3744 2931 3876
rect 2909 3344 2915 3696
rect 2925 3464 2931 3736
rect 2957 3564 2963 3756
rect 3005 3704 3011 3736
rect 3021 3604 3027 3856
rect 3165 3784 3171 3896
rect 3645 3884 3651 3896
rect 3252 3797 3260 3803
rect 2941 3364 2947 3456
rect 3005 3344 3011 3516
rect 3021 3464 3027 3596
rect 2733 2984 2739 3096
rect 2813 2984 2819 3096
rect 2701 2304 2707 2696
rect 2717 2344 2723 2556
rect 2669 1764 2675 2236
rect 2685 2124 2691 2156
rect 2685 1924 2691 1976
rect 2685 1504 2691 1516
rect 2525 1044 2531 1116
rect 2541 364 2547 1116
rect 2557 784 2563 916
rect 2605 684 2611 1276
rect 2621 1104 2627 1116
rect 2637 1064 2643 1096
rect 2685 1064 2691 1436
rect 2701 1324 2707 2296
rect 2717 1944 2723 2196
rect 2717 1924 2723 1936
rect 2701 1064 2707 1316
rect 2717 1284 2723 1796
rect 2733 1564 2739 2016
rect 2749 1964 2755 2896
rect 2781 2284 2787 2696
rect 2669 904 2675 976
rect 2557 564 2563 576
rect 2621 524 2627 756
rect 2685 664 2691 1056
rect 2644 577 2652 583
rect 2637 524 2643 536
rect 2621 504 2627 516
rect 2685 504 2691 656
rect 2701 504 2707 1056
rect 2717 884 2723 1256
rect 2733 904 2739 1476
rect 2749 1044 2755 1456
rect 2765 1284 2771 2216
rect 2781 2144 2787 2276
rect 2749 904 2755 916
rect 2765 904 2771 1096
rect 2781 964 2787 2136
rect 2845 1884 2851 3256
rect 2909 3004 2915 3156
rect 2884 2957 2892 2963
rect 2996 2917 3004 2923
rect 3005 2704 3011 2816
rect 3021 2684 3027 2956
rect 3069 2784 3075 3776
rect 3133 3644 3139 3736
rect 3101 3424 3107 3536
rect 3085 2964 3091 3196
rect 3101 3124 3107 3356
rect 2980 2557 2988 2563
rect 2909 2544 2915 2556
rect 2877 2184 2883 2216
rect 2836 1877 2844 1883
rect 2909 1804 2915 2276
rect 2957 2164 2963 2556
rect 2925 2104 2931 2136
rect 2925 1864 2931 1876
rect 2941 1744 2947 1996
rect 2973 1904 2979 2556
rect 2989 2144 2995 2176
rect 2989 1864 2995 2116
rect 3005 1864 3011 2676
rect 3021 2144 3027 2676
rect 3053 2644 3059 2656
rect 3037 2544 3043 2556
rect 2884 1737 2892 1743
rect 2829 1724 2835 1736
rect 2797 1504 2803 1516
rect 2717 624 2723 856
rect 2781 844 2787 856
rect 2701 284 2707 496
rect 2717 344 2723 616
rect 2749 324 2755 756
rect 2797 624 2803 1296
rect 2813 544 2819 1076
rect 2829 984 2835 996
rect 2829 304 2835 956
rect 2845 524 2851 1036
rect 2861 884 2867 916
rect 2861 704 2867 856
rect 2845 324 2851 336
rect 2573 184 2579 276
rect 2653 144 2659 256
rect 2829 144 2835 296
rect 2861 244 2867 336
rect 2877 264 2883 936
rect 2893 764 2899 1736
rect 2909 944 2915 1376
rect 2989 1084 2995 1556
rect 3005 1304 3011 1396
rect 3037 1304 3043 1716
rect 3053 1704 3059 2636
rect 3069 2524 3075 2536
rect 3069 2284 3075 2516
rect 2893 564 2899 736
rect 2893 444 2899 536
rect 2893 244 2899 436
rect 2909 284 2915 936
rect 2941 784 2947 876
rect 2957 544 2963 1076
rect 2989 904 2995 1076
rect 3037 724 3043 1296
rect 3069 1064 3075 1496
rect 3085 1484 3091 2156
rect 3101 1724 3107 3116
rect 3133 2924 3139 3636
rect 3197 3464 3203 3576
rect 3213 3544 3219 3796
rect 3357 3764 3363 3776
rect 3325 3684 3331 3756
rect 3213 3004 3219 3496
rect 3229 3464 3235 3636
rect 3149 2924 3155 2936
rect 3188 2897 3196 2903
rect 3069 1024 3075 1056
rect 3053 884 3059 956
rect 3085 944 3091 1436
rect 3101 1004 3107 1356
rect 3117 1044 3123 2276
rect 3133 2144 3139 2756
rect 3149 2444 3155 2736
rect 3197 2724 3203 2876
rect 3197 2284 3203 2696
rect 3213 2684 3219 2996
rect 3213 2384 3219 2576
rect 3229 2524 3235 3456
rect 3293 3424 3299 3536
rect 3245 3304 3251 3316
rect 3261 3104 3267 3116
rect 3252 2997 3267 3003
rect 3261 2984 3267 2997
rect 3245 2904 3251 2936
rect 3245 2544 3251 2896
rect 3133 1444 3139 2136
rect 3149 1464 3155 1856
rect 3181 1524 3187 1956
rect 3197 1904 3203 2276
rect 3213 1883 3219 2356
rect 3229 2204 3235 2456
rect 3229 2164 3235 2176
rect 3245 2104 3251 2536
rect 3261 2304 3267 2496
rect 3277 2264 3283 3256
rect 3325 3184 3331 3336
rect 3325 3104 3331 3116
rect 3300 2677 3308 2683
rect 3293 2544 3299 2636
rect 3325 2564 3331 3096
rect 3341 3004 3347 3756
rect 3357 3424 3363 3436
rect 3357 3064 3363 3076
rect 3341 2984 3347 2996
rect 3373 2884 3379 3436
rect 3389 3064 3395 3356
rect 3421 3304 3427 3316
rect 3437 3284 3443 3356
rect 3469 3324 3475 3376
rect 3469 3144 3475 3176
rect 3485 3063 3491 3536
rect 3501 3404 3507 3856
rect 3501 3324 3507 3336
rect 3501 3084 3507 3096
rect 3485 3057 3507 3063
rect 3341 2864 3347 2876
rect 3341 2724 3347 2816
rect 3293 2464 3299 2476
rect 3341 2464 3347 2576
rect 3309 2204 3315 2216
rect 3309 1984 3315 2116
rect 3197 1877 3219 1883
rect 3165 1464 3171 1496
rect 3149 1184 3155 1456
rect 3181 1284 3187 1516
rect 3069 684 3075 796
rect 3085 784 3091 936
rect 2861 144 2867 236
rect 2893 184 2899 236
rect 2957 164 2963 536
rect 2973 264 2979 396
rect 3069 384 3075 656
rect 3085 624 3091 736
rect 3085 604 3091 616
rect 3069 284 3075 376
rect 2973 204 2979 256
rect 2877 124 2883 136
rect 2349 104 2355 116
rect 2116 97 2124 103
rect 2253 64 2259 96
rect 2957 24 2963 156
rect 2973 144 2979 196
rect 3101 184 3107 836
rect 3101 164 3107 176
rect 3117 104 3123 1036
rect 3165 844 3171 1016
rect 3181 824 3187 1276
rect 3133 464 3139 636
rect 3197 604 3203 1877
rect 3213 1264 3219 1296
rect 3229 944 3235 1896
rect 3261 1744 3267 1976
rect 3293 1524 3299 1796
rect 3268 1497 3276 1503
rect 3245 1364 3251 1496
rect 3293 1464 3299 1496
rect 3261 1024 3267 1456
rect 3277 1124 3283 1396
rect 3325 1364 3331 1476
rect 3293 1264 3299 1296
rect 3277 904 3283 1076
rect 3293 1004 3299 1156
rect 3325 1044 3331 1356
rect 3213 784 3219 836
rect 3252 677 3260 683
rect 3165 584 3171 596
rect 3261 464 3267 676
rect 3277 664 3283 676
rect 3133 244 3139 276
rect 3261 264 3267 336
rect 3245 244 3251 256
rect 3277 224 3283 656
rect 3325 644 3331 1036
rect 3341 984 3347 1256
rect 3357 624 3363 2776
rect 3389 2564 3395 3056
rect 3460 2977 3468 2983
rect 3485 2963 3491 2976
rect 3437 2957 3491 2963
rect 3437 2904 3443 2957
rect 3460 2897 3468 2903
rect 3405 2864 3411 2876
rect 3405 2164 3411 2816
rect 3405 2084 3411 2116
rect 3389 2064 3395 2076
rect 3373 1964 3379 1996
rect 3421 1884 3427 2676
rect 3485 2544 3491 2916
rect 3501 2644 3507 3057
rect 3517 2704 3523 3036
rect 3565 2984 3571 3836
rect 3597 3764 3603 3776
rect 3581 3364 3587 3376
rect 3581 2964 3587 3336
rect 3533 2884 3539 2896
rect 3517 2684 3523 2696
rect 3517 2564 3523 2576
rect 3373 1704 3379 1836
rect 3405 1824 3411 1856
rect 3389 1364 3395 1416
rect 3389 944 3395 956
rect 3405 904 3411 1816
rect 3437 1064 3443 1756
rect 3453 1524 3459 1536
rect 3469 1524 3475 2476
rect 3485 1804 3491 2536
rect 3517 2184 3523 2356
rect 3517 1904 3523 2036
rect 3469 1384 3475 1396
rect 3485 1364 3491 1496
rect 3501 1384 3507 1556
rect 3517 1264 3523 1416
rect 3533 1404 3539 2296
rect 3549 2164 3555 2956
rect 3581 2644 3587 2956
rect 3597 2664 3603 3756
rect 3613 3304 3619 3336
rect 3613 2704 3619 2996
rect 3629 2684 3635 3756
rect 3645 3244 3651 3876
rect 3789 3824 3795 3916
rect 3821 3904 3827 3916
rect 3876 3877 3884 3883
rect 3773 3704 3779 3716
rect 3581 2584 3587 2596
rect 3565 2504 3571 2536
rect 3565 2224 3571 2496
rect 3549 1864 3555 2156
rect 3549 1724 3555 1856
rect 3565 1424 3571 2076
rect 3581 1784 3587 2516
rect 3597 2504 3603 2616
rect 3613 2524 3619 2656
rect 3629 2484 3635 2496
rect 3604 2297 3612 2303
rect 3645 2144 3651 3236
rect 3661 3064 3667 3336
rect 3661 3024 3667 3056
rect 3661 2644 3667 2656
rect 3661 2184 3667 2636
rect 3677 2224 3683 3196
rect 3693 3064 3699 3356
rect 3709 3024 3715 3056
rect 3693 2464 3699 2916
rect 3709 2664 3715 2956
rect 3725 2684 3731 3376
rect 3757 3084 3763 3176
rect 3741 2924 3747 2956
rect 3741 2844 3747 2856
rect 3757 2704 3763 3076
rect 3773 2964 3779 3696
rect 3789 3064 3795 3796
rect 3805 3704 3811 3876
rect 4125 3824 4131 3876
rect 3821 3444 3827 3476
rect 3853 3384 3859 3736
rect 3805 3204 3811 3216
rect 3805 3164 3811 3176
rect 3805 3144 3811 3156
rect 3789 3044 3795 3056
rect 3853 3044 3859 3316
rect 3773 2704 3779 2716
rect 3716 2657 3724 2663
rect 3716 2537 3724 2543
rect 3661 2124 3667 2136
rect 3677 1924 3683 2216
rect 3581 1764 3587 1776
rect 3581 1384 3587 1536
rect 3597 1524 3603 1536
rect 3613 1364 3619 1376
rect 3453 1104 3459 1116
rect 3437 1004 3443 1056
rect 3389 804 3395 816
rect 3453 584 3459 956
rect 3469 664 3475 696
rect 3309 564 3315 576
rect 3412 517 3420 523
rect 3405 424 3411 476
rect 3245 144 3251 156
rect 3277 124 3283 216
rect 3309 164 3315 276
rect 3325 224 3331 256
rect 3453 204 3459 456
rect 3325 144 3331 156
rect 3469 144 3475 656
rect 3485 544 3491 1056
rect 3517 844 3523 1036
rect 3565 984 3571 1136
rect 3629 664 3635 1056
rect 3645 944 3651 1736
rect 3661 1384 3667 1396
rect 3677 1104 3683 1896
rect 3693 1744 3699 2456
rect 3709 2304 3715 2336
rect 3709 2244 3715 2256
rect 3709 2104 3715 2176
rect 3725 2124 3731 2136
rect 3709 1904 3715 2056
rect 3709 1723 3715 1856
rect 3693 1717 3715 1723
rect 3693 1544 3699 1717
rect 3725 1704 3731 1916
rect 3693 1364 3699 1496
rect 3709 1384 3715 1696
rect 3725 1604 3731 1616
rect 3709 1324 3715 1356
rect 3661 783 3667 856
rect 3645 777 3667 783
rect 3645 764 3651 777
rect 3661 684 3667 756
rect 3709 724 3715 1176
rect 3725 1064 3731 1496
rect 3741 1324 3747 2676
rect 3757 1864 3763 2696
rect 3773 2624 3779 2676
rect 3789 2584 3795 3036
rect 3853 2924 3859 3016
rect 3869 2944 3875 3736
rect 3901 3484 3907 3816
rect 4036 3797 4044 3803
rect 3917 3757 3955 3763
rect 3917 3724 3923 3757
rect 3949 3744 3955 3757
rect 3933 3724 3939 3736
rect 3965 3684 3971 3696
rect 4020 3517 4028 3523
rect 3885 2944 3891 3256
rect 3901 3104 3907 3476
rect 3981 3424 3987 3456
rect 4045 3424 4051 3516
rect 3981 3384 3987 3416
rect 4045 3204 4051 3416
rect 4077 3404 4083 3796
rect 4077 3304 4083 3336
rect 4045 3124 4051 3136
rect 3805 2624 3811 2716
rect 3844 2697 3852 2703
rect 3773 2524 3779 2536
rect 3732 1057 3740 1063
rect 3757 924 3763 1856
rect 3773 1504 3779 2516
rect 3789 1764 3795 2576
rect 3805 2284 3811 2296
rect 3837 2264 3843 2296
rect 3869 2244 3875 2796
rect 3885 2664 3891 2936
rect 3789 1483 3795 1756
rect 3805 1524 3811 2196
rect 3821 2104 3827 2116
rect 3853 1764 3859 2176
rect 3885 1884 3891 2276
rect 3901 2144 3907 3076
rect 3981 3004 3987 3016
rect 4061 2944 4067 3036
rect 3917 2584 3923 2876
rect 3933 2544 3939 2916
rect 3965 2263 3971 2656
rect 3981 2504 3987 2516
rect 4029 2504 4035 2936
rect 4061 2724 4067 2736
rect 3949 2257 3971 2263
rect 3773 1477 3795 1483
rect 3725 664 3731 676
rect 3501 524 3507 536
rect 3517 384 3523 616
rect 3652 537 3660 543
rect 3533 304 3539 476
rect 3588 377 3596 383
rect 3725 304 3731 656
rect 3517 184 3523 196
rect 3693 184 3699 236
rect 3757 184 3763 596
rect 3773 264 3779 1477
rect 3789 1124 3795 1136
rect 3805 1084 3811 1096
rect 3821 1084 3827 1756
rect 3837 1344 3843 1736
rect 3837 1084 3843 1336
rect 3821 964 3827 1076
rect 3837 964 3843 996
rect 3837 684 3843 756
rect 3853 704 3859 1456
rect 3789 484 3795 676
rect 3805 304 3811 636
rect 3837 324 3843 616
rect 3853 604 3859 696
rect 3869 684 3875 1476
rect 3901 524 3907 1496
rect 3917 1364 3923 1656
rect 3933 1444 3939 1696
rect 3949 1504 3955 2257
rect 3997 2244 4003 2456
rect 4020 2257 4028 2263
rect 3965 2084 3971 2096
rect 4013 1864 4019 2256
rect 4045 2124 4051 2656
rect 3965 1684 3971 1836
rect 3965 1464 3971 1676
rect 3981 1524 3987 1856
rect 3997 1484 4003 1776
rect 3949 1384 3955 1396
rect 3949 1284 3955 1336
rect 3949 1184 3955 1256
rect 3933 964 3939 1156
rect 3949 1084 3955 1116
rect 3965 984 3971 1456
rect 3933 644 3939 756
rect 3901 384 3907 516
rect 3917 344 3923 616
rect 3924 317 3932 323
rect 3837 244 3843 316
rect 3869 304 3875 316
rect 3885 264 3891 296
rect 3933 264 3939 316
rect 3780 177 3788 183
rect 3757 164 3763 176
rect 3949 164 3955 556
rect 3965 344 3971 736
rect 3981 684 3987 1356
rect 3981 664 3987 676
rect 3997 604 4003 1456
rect 4045 1424 4051 1596
rect 4013 1004 4019 1156
rect 4045 1084 4051 1096
rect 4061 964 4067 2636
rect 4077 2604 4083 3296
rect 4077 1784 4083 2516
rect 4093 2163 4099 3316
rect 4109 3064 4115 3456
rect 4109 2284 4115 3056
rect 4125 2644 4131 3256
rect 4109 2184 4115 2196
rect 4093 2157 4108 2163
rect 4093 1984 4099 2056
rect 4093 1764 4099 1776
rect 4109 1764 4115 1896
rect 4125 1704 4131 2636
rect 4141 2544 4147 3716
rect 4157 3404 4163 3576
rect 4157 3164 4163 3196
rect 4173 2984 4179 3776
rect 4237 3524 4243 3796
rect 4477 3784 4483 3836
rect 4301 3744 4307 3756
rect 4276 3697 4284 3703
rect 4189 3464 4195 3476
rect 4157 2684 4163 2956
rect 4141 1884 4147 2536
rect 4157 2204 4163 2356
rect 4173 2244 4179 2976
rect 4189 2664 4195 3456
rect 4205 3304 4211 3336
rect 4269 2904 4275 3436
rect 4285 3404 4291 3436
rect 4189 2064 4195 2536
rect 4221 2304 4227 2676
rect 4237 2664 4243 2676
rect 4205 2284 4211 2296
rect 4237 2244 4243 2536
rect 4237 1944 4243 2196
rect 4141 1764 4147 1876
rect 4173 1424 4179 1456
rect 4125 1324 4131 1396
rect 4189 1364 4195 1796
rect 4253 1784 4259 2896
rect 4285 2763 4291 3156
rect 4269 2757 4291 2763
rect 4269 2384 4275 2757
rect 4285 2344 4291 2536
rect 4285 2304 4291 2316
rect 4269 2284 4275 2296
rect 4301 2284 4307 3736
rect 4445 3704 4451 3756
rect 4365 3644 4371 3696
rect 4509 3524 4515 3536
rect 4461 3504 4467 3516
rect 4317 3164 4323 3436
rect 4365 3364 4371 3396
rect 4445 3384 4451 3396
rect 4372 3157 4380 3163
rect 4317 3064 4323 3096
rect 4317 2744 4323 2956
rect 4317 2283 4323 2356
rect 4349 2344 4355 3116
rect 4413 3064 4419 3116
rect 4413 2924 4419 2936
rect 4388 2697 4396 2703
rect 4317 2277 4339 2283
rect 4269 1904 4275 2156
rect 4285 2104 4291 2116
rect 4093 1024 4099 1176
rect 3981 584 3987 596
rect 3981 164 3987 576
rect 4013 564 4019 856
rect 4036 757 4044 763
rect 4052 657 4060 663
rect 4077 624 4083 876
rect 4093 644 4099 676
rect 4109 664 4115 1316
rect 3981 104 3987 156
rect 3997 84 4003 336
rect 4061 264 4067 296
rect 4093 184 4099 296
rect 4109 284 4115 656
rect 4125 644 4131 1116
rect 4141 644 4147 656
rect 4157 624 4163 1296
rect 4205 1264 4211 1296
rect 4221 1124 4227 1396
rect 4237 1304 4243 1776
rect 4285 1764 4291 1776
rect 4212 917 4220 923
rect 4212 877 4220 883
rect 4189 784 4195 816
rect 4180 737 4188 743
rect 4205 684 4211 756
rect 4237 684 4243 1276
rect 4253 884 4259 1736
rect 4301 1724 4307 2276
rect 4333 2224 4339 2277
rect 4333 1884 4339 1896
rect 4228 597 4236 603
rect 4253 584 4259 876
rect 4269 744 4275 1536
rect 4333 1484 4339 1876
rect 4349 1804 4355 2236
rect 4365 2124 4371 2236
rect 4349 1684 4355 1736
rect 4317 1304 4323 1316
rect 4333 1104 4339 1116
rect 4285 864 4291 876
rect 4301 864 4307 916
rect 4317 704 4323 1056
rect 4349 964 4355 1396
rect 4276 697 4284 703
rect 4189 564 4195 576
rect 4205 504 4211 576
rect 4221 484 4227 536
rect 4237 524 4243 556
rect 4141 164 4147 456
rect 4157 184 4163 216
rect 4221 164 4227 396
rect 4237 284 4243 516
rect 4237 244 4243 256
rect 4253 244 4259 576
rect 4269 444 4275 676
rect 4349 664 4355 696
rect 4365 544 4371 1056
rect 4381 744 4387 2576
rect 4429 2564 4435 3056
rect 4445 2684 4451 3336
rect 4429 2404 4435 2516
rect 4445 2504 4451 2576
rect 4429 2124 4435 2396
rect 4461 2284 4467 3496
rect 4493 3344 4499 3356
rect 4500 3277 4508 3283
rect 4509 2924 4515 2956
rect 4525 2724 4531 3916
rect 4541 2784 4547 3816
rect 4669 3424 4675 3476
rect 4573 3124 4579 3216
rect 4589 3144 4595 3156
rect 4605 3123 4611 3136
rect 4589 3117 4611 3123
rect 4557 3103 4563 3116
rect 4589 3103 4595 3117
rect 4557 3097 4595 3103
rect 4477 2584 4483 2656
rect 4541 2643 4547 2656
rect 4557 2644 4563 3016
rect 4653 2704 4659 3356
rect 4669 3124 4675 3396
rect 4685 3364 4691 3796
rect 4717 3364 4723 3756
rect 4733 3744 4739 3756
rect 4749 3484 4755 3856
rect 4765 3704 4771 3756
rect 4756 3377 4764 3383
rect 4781 3344 4787 3396
rect 4685 2644 4691 3336
rect 4708 3117 4716 3123
rect 4733 3004 4739 3256
rect 4733 2744 4739 2976
rect 4749 2924 4755 2936
rect 4781 2884 4787 2936
rect 4532 2637 4547 2643
rect 4557 2484 4563 2616
rect 4605 2584 4611 2596
rect 4621 2583 4627 2596
rect 4621 2577 4659 2583
rect 4653 2563 4659 2577
rect 4653 2557 4675 2563
rect 4669 2544 4675 2557
rect 4573 2484 4579 2496
rect 4413 1444 4419 1856
rect 4429 1704 4435 1796
rect 4445 1764 4451 1836
rect 4429 1444 4435 1496
rect 4461 1104 4467 2276
rect 4477 2164 4483 2296
rect 4580 2277 4588 2283
rect 4605 2184 4611 2496
rect 4564 2137 4572 2143
rect 4548 2117 4556 2123
rect 4477 1224 4483 2116
rect 4621 2104 4627 2516
rect 4637 2284 4643 2536
rect 4493 1544 4499 1956
rect 4621 1904 4627 1916
rect 4621 1843 4627 1896
rect 4637 1864 4643 2276
rect 4653 1924 4659 2256
rect 4669 2084 4675 2176
rect 4621 1837 4643 1843
rect 4621 1784 4627 1796
rect 4509 1624 4515 1656
rect 4525 1524 4531 1576
rect 4541 1544 4547 1576
rect 4381 584 4387 716
rect 4445 564 4451 616
rect 4285 504 4291 516
rect 4333 504 4339 516
rect 4269 244 4275 276
rect 4317 224 4323 496
rect 4365 384 4371 536
rect 4349 264 4355 356
rect 4365 344 4371 376
rect 4365 284 4371 336
rect 4397 304 4403 316
rect 4461 144 4467 1096
rect 4493 1064 4499 1376
rect 4477 564 4483 876
rect 4493 704 4499 1056
rect 4509 724 4515 1456
rect 4573 1384 4579 1496
rect 4477 184 4483 376
rect 4493 324 4499 696
rect 4509 304 4515 716
rect 4541 684 4547 756
rect 4557 744 4563 996
rect 4573 944 4579 1336
rect 4596 1317 4604 1323
rect 4573 504 4579 936
rect 4589 824 4595 1156
rect 4621 1084 4627 1756
rect 4637 1424 4643 1837
rect 4685 1744 4691 2636
rect 4701 1864 4707 2176
rect 4653 1544 4659 1576
rect 4589 564 4595 576
rect 4541 124 4547 176
rect 4605 124 4611 256
rect 4372 117 4380 123
rect 4301 104 4307 116
rect 4589 84 4595 116
rect 3853 64 3859 76
rect 4621 -17 4627 596
rect 4653 44 4659 1016
rect 4669 604 4675 1736
rect 4701 1704 4707 1856
rect 4717 1804 4723 2096
rect 4733 1884 4739 2536
rect 4749 2304 4755 2676
rect 4765 2544 4771 2656
rect 4797 2544 4803 3336
rect 4829 3064 4835 3076
rect 4829 2984 4835 3056
rect 4845 2944 4851 3456
rect 4884 3297 4892 3303
rect 4861 3284 4867 3296
rect 4868 3097 4876 3103
rect 4733 1644 4739 1716
rect 4733 1324 4739 1636
rect 4749 1324 4755 1796
rect 4765 1524 4771 2536
rect 4813 2484 4819 2496
rect 4781 2224 4787 2256
rect 4813 2224 4819 2276
rect 4781 1924 4787 1936
rect 4781 1604 4787 1896
rect 4701 1124 4707 1136
rect 4765 1124 4771 1156
rect 4749 1104 4755 1116
rect 4708 997 4716 1003
rect 4669 584 4675 596
rect 4717 324 4723 976
rect 4733 944 4739 996
rect 4749 884 4755 1096
rect 4749 744 4755 796
rect 4765 684 4771 736
rect 4685 124 4691 176
rect 4781 104 4787 1576
rect 4797 1544 4803 2216
rect 4829 2164 4835 2916
rect 4845 2384 4851 2936
rect 4861 2924 4867 2936
rect 4861 2624 4867 2876
rect 4813 1824 4819 2156
rect 4829 1904 4835 2156
rect 4845 2124 4851 2196
rect 4829 1684 4835 1896
rect 4845 1704 4851 1816
rect 4813 1544 4819 1656
rect 4797 1064 4803 1356
rect 4813 1264 4819 1416
rect 4813 1224 4819 1236
rect 4797 864 4803 876
rect 4829 824 4835 1476
rect 4845 784 4851 1456
rect 4861 1104 4867 2236
rect 4877 1824 4883 2956
rect 4893 2244 4899 3136
rect 4909 3084 4915 3456
rect 4925 3324 4931 3696
rect 4941 3384 4947 3456
rect 4957 3424 4963 3436
rect 4925 3084 4931 3096
rect 4941 3044 4947 3316
rect 4925 2944 4931 2956
rect 4909 2704 4915 2716
rect 4925 2664 4931 2876
rect 4925 2564 4931 2656
rect 4941 2544 4947 3036
rect 4925 2524 4931 2536
rect 4916 2497 4924 2503
rect 4909 2204 4915 2436
rect 4909 2104 4915 2136
rect 4900 1917 4908 1923
rect 4909 1844 4915 1876
rect 4797 724 4803 736
rect 4861 724 4867 1096
rect 4877 1064 4883 1096
rect 4845 324 4851 696
rect 4861 664 4867 696
rect 4893 684 4899 1736
rect 4909 1524 4915 1596
rect 4925 1504 4931 2256
rect 4941 1724 4947 2536
rect 4957 2504 4963 3416
rect 4973 3124 4979 3136
rect 4989 2964 4995 3476
rect 5005 2964 5011 3776
rect 5069 3544 5075 3796
rect 5133 3744 5139 3856
rect 5181 3764 5187 3776
rect 5181 3744 5187 3756
rect 5197 3724 5203 3736
rect 5021 3464 5027 3496
rect 5117 3397 5132 3403
rect 5021 3124 5027 3396
rect 5053 3104 5059 3116
rect 5085 3044 5091 3056
rect 4957 2164 4963 2196
rect 4941 1524 4947 1536
rect 4957 1484 4963 2116
rect 4973 1664 4979 2716
rect 5005 2584 5011 2956
rect 5021 2724 5027 2736
rect 4989 2564 4995 2576
rect 4996 2537 5004 2543
rect 5021 2524 5027 2616
rect 5037 2524 5043 2536
rect 5005 2324 5011 2516
rect 5005 2184 5011 2196
rect 5021 1884 5027 2236
rect 5037 2164 5043 2376
rect 5005 1764 5011 1776
rect 4973 1484 4979 1496
rect 4957 1364 4963 1476
rect 4957 1044 4963 1056
rect 4957 884 4963 916
rect 4973 904 4979 996
rect 4941 704 4947 716
rect 4877 564 4883 576
rect 4893 564 4899 676
rect 4973 344 4979 596
rect 4989 584 4995 1756
rect 5037 1724 5043 1996
rect 5053 1863 5059 2616
rect 5069 1884 5075 2936
rect 5053 1857 5075 1863
rect 5005 984 5011 1716
rect 5069 1544 5075 1857
rect 5085 1764 5091 3036
rect 5101 2284 5107 3076
rect 5117 2904 5123 3376
rect 5133 3364 5139 3376
rect 5124 2317 5132 2323
rect 5101 2183 5107 2216
rect 5149 2184 5155 2676
rect 5165 2544 5171 2556
rect 5181 2264 5187 3376
rect 5197 3344 5203 3356
rect 5101 2177 5123 2183
rect 5117 2164 5123 2177
rect 5101 2144 5107 2156
rect 5181 2124 5187 2156
rect 5149 2044 5155 2056
rect 5037 1504 5043 1516
rect 5037 1124 5043 1356
rect 5069 1204 5075 1356
rect 5069 1044 5075 1096
rect 5037 984 5043 996
rect 5101 944 5107 1856
rect 5037 744 5043 756
rect 5053 684 5059 756
rect 5069 744 5075 756
rect 5053 604 5059 676
rect 5069 604 5075 716
rect 5005 504 5011 596
rect 4845 304 4851 316
rect 5021 304 5027 316
rect 4829 224 4835 296
rect 4877 204 4883 256
rect 4925 224 4931 256
rect 5037 164 5043 336
rect 5085 224 5091 916
rect 5117 764 5123 1696
rect 5133 1464 5139 1776
rect 5149 1044 5155 1316
rect 5165 1144 5171 1156
rect 5165 1064 5171 1076
rect 5133 924 5139 956
rect 5117 704 5123 716
rect 5133 624 5139 836
rect 5149 204 5155 636
rect 5165 384 5171 836
rect 5181 224 5187 1776
rect 5197 184 5203 3316
rect 5213 924 5219 3876
rect 5245 3784 5251 3816
rect 5245 3744 5251 3756
rect 5229 2264 5235 2996
rect 5245 2944 5251 3096
rect 5261 3064 5267 3476
rect 5245 2204 5251 2476
rect 5261 2284 5267 3056
rect 5277 2584 5283 3616
rect 5261 2244 5267 2276
rect 5229 224 5235 1816
rect 5245 1724 5251 1936
rect 5261 1104 5267 2076
rect 5277 1844 5283 2576
rect 5293 2504 5299 3876
rect 5309 3844 5315 3863
rect 5245 304 5251 696
rect 5245 204 5251 256
rect 5245 164 5251 176
rect 5261 144 5267 716
rect 5277 704 5283 1836
rect 5293 1784 5299 2096
rect 5309 1784 5315 3796
rect 5300 1737 5308 1743
rect 5293 1524 5299 1536
rect 5325 1364 5331 3896
rect 5341 3764 5347 3776
rect 5341 2524 5347 3736
rect 5357 2424 5363 3876
rect 5396 3117 5404 3123
rect 5373 2784 5379 2996
rect 5380 2677 5388 2683
rect 5373 1804 5379 2536
rect 5405 2143 5411 2896
rect 5421 2164 5427 3796
rect 5405 2137 5427 2143
rect 5396 2077 5404 2083
rect 5316 1337 5324 1343
rect 5293 684 5299 1036
rect 5309 1024 5315 1296
rect 5293 544 5299 676
rect 5309 564 5315 976
rect 5325 544 5331 1116
rect 5284 537 5292 543
rect 5309 263 5315 436
rect 5293 257 5315 263
rect 5293 164 5299 257
rect 5325 84 5331 316
rect 5341 164 5347 1756
rect 5373 1744 5379 1756
rect 5389 1683 5395 1876
rect 5373 1677 5395 1683
rect 5357 284 5363 1076
rect 5373 684 5379 1677
rect 5389 904 5395 956
rect 5405 924 5411 936
rect 5380 557 5388 563
rect 5421 64 5427 2137
rect 5437 1984 5443 3776
rect 5453 2964 5459 3536
rect 5453 2224 5459 2316
rect 5453 1404 5459 2076
rect 5437 504 5443 936
rect 5453 504 5459 1056
rect 5469 204 5475 3916
rect 5485 2744 5491 3376
rect 5517 3084 5523 3756
rect 5517 2684 5523 3076
rect 5661 3004 5667 3116
rect 5501 2524 5507 2576
rect 5508 2317 5516 2323
rect 5508 1877 5516 1883
rect 5533 1504 5539 1516
rect 5444 137 5452 143
rect 4685 -17 4691 16
rect 4621 -23 4691 -17
<< m5contact >>
rect 284 3716 292 3724
rect 92 3096 100 3104
rect 124 3076 132 3084
rect 124 2976 132 2984
rect 188 3336 196 3344
rect 124 2556 132 2564
rect 172 2136 180 2144
rect 252 3076 260 3084
rect 316 3336 324 3344
rect 380 3336 388 3344
rect 300 3016 308 3024
rect 268 2896 276 2904
rect 124 1296 132 1304
rect 124 1116 132 1124
rect 172 1056 180 1064
rect 124 916 132 924
rect 12 176 20 184
rect 76 176 84 184
rect 284 1076 292 1084
rect 300 1056 308 1064
rect 380 2956 388 2964
rect 364 2896 372 2904
rect 348 2116 356 2124
rect 348 2096 356 2104
rect 396 2136 404 2144
rect 364 1076 372 1084
rect 700 3776 708 3784
rect 476 3736 484 3744
rect 524 3736 532 3744
rect 460 3536 468 3544
rect 556 3716 564 3724
rect 636 3516 644 3524
rect 716 3496 724 3504
rect 524 3116 532 3124
rect 540 3096 548 3104
rect 572 3036 580 3044
rect 460 3016 468 3024
rect 524 2936 532 2944
rect 556 2696 564 2704
rect 636 3176 644 3184
rect 572 2676 580 2684
rect 508 2616 516 2624
rect 476 2136 484 2144
rect 444 2116 452 2124
rect 428 1956 436 1964
rect 460 1916 468 1924
rect 396 936 404 944
rect 780 3776 788 3784
rect 812 3756 820 3764
rect 764 3736 772 3744
rect 764 3516 772 3524
rect 764 3316 772 3324
rect 748 3096 756 3104
rect 764 3076 772 3084
rect 732 2696 740 2704
rect 668 2676 676 2684
rect 636 2556 644 2564
rect 492 1676 500 1684
rect 460 1336 468 1344
rect 460 936 468 944
rect 460 876 468 884
rect 620 2136 628 2144
rect 588 1836 596 1844
rect 572 1496 580 1504
rect 524 1316 532 1324
rect 540 1096 548 1104
rect 380 696 388 704
rect 284 336 292 344
rect 300 276 308 284
rect 668 2556 676 2564
rect 684 2296 692 2304
rect 668 1856 676 1864
rect 732 2116 740 2124
rect 780 2796 788 2804
rect 780 2696 788 2704
rect 780 2536 788 2544
rect 780 2116 788 2124
rect 748 2076 756 2084
rect 764 1916 772 1924
rect 684 1836 692 1844
rect 652 1716 660 1724
rect 764 1716 772 1724
rect 748 1536 756 1544
rect 636 1336 644 1344
rect 732 1296 740 1304
rect 620 1076 628 1084
rect 636 1056 644 1064
rect 716 1056 724 1064
rect 700 1016 708 1024
rect 604 616 612 624
rect 572 336 580 344
rect 508 256 516 264
rect 684 296 692 304
rect 716 296 724 304
rect 828 3496 836 3504
rect 892 3756 900 3764
rect 860 3736 868 3744
rect 972 3776 980 3784
rect 892 3416 900 3424
rect 860 3096 868 3104
rect 860 2676 868 2684
rect 844 2656 852 2664
rect 812 2296 820 2304
rect 812 1976 820 1984
rect 796 1756 804 1764
rect 796 1696 804 1704
rect 844 1996 852 2004
rect 924 2916 932 2924
rect 924 2756 932 2764
rect 924 2716 932 2724
rect 892 2316 900 2324
rect 892 2156 900 2164
rect 876 1936 884 1944
rect 876 1896 884 1904
rect 892 1776 900 1784
rect 844 1756 852 1764
rect 796 1356 804 1364
rect 780 1036 788 1044
rect 860 1516 868 1524
rect 860 1336 868 1344
rect 812 956 820 964
rect 844 1056 852 1064
rect 828 736 836 744
rect 796 716 804 724
rect 1052 3496 1060 3504
rect 988 2976 996 2984
rect 1036 3076 1044 3084
rect 988 2676 996 2684
rect 972 2316 980 2324
rect 956 2176 964 2184
rect 972 2156 980 2164
rect 940 2076 948 2084
rect 956 1916 964 1924
rect 940 1896 948 1904
rect 956 1796 964 1804
rect 972 1776 980 1784
rect 988 1736 996 1744
rect 988 1716 996 1724
rect 956 1456 964 1464
rect 1084 3776 1092 3784
rect 1276 3736 1284 3744
rect 1180 3676 1188 3684
rect 1084 3356 1092 3364
rect 1084 3236 1092 3244
rect 1100 3096 1108 3104
rect 1132 3056 1140 3064
rect 1212 3536 1220 3544
rect 1228 3156 1236 3164
rect 1164 3036 1172 3044
rect 1180 3036 1188 3044
rect 1084 3016 1092 3024
rect 1084 2916 1092 2924
rect 1100 2716 1108 2724
rect 1052 2696 1060 2704
rect 1052 2656 1060 2664
rect 1068 2656 1076 2664
rect 1052 2536 1060 2544
rect 1148 2916 1156 2924
rect 1132 2696 1140 2704
rect 1036 2156 1044 2164
rect 1020 2096 1028 2104
rect 1052 1936 1060 1944
rect 1036 1836 1044 1844
rect 940 1036 948 1044
rect 940 876 948 884
rect 972 796 980 804
rect 972 776 980 784
rect 1004 976 1012 984
rect 1036 1376 1044 1384
rect 1068 1356 1076 1364
rect 1164 2276 1172 2284
rect 1148 2116 1156 2124
rect 1132 2096 1140 2104
rect 1196 2916 1204 2924
rect 1196 2776 1204 2784
rect 1196 2756 1204 2764
rect 1260 3316 1268 3324
rect 1260 3096 1268 3104
rect 1292 3376 1300 3384
rect 1276 2976 1284 2984
rect 1468 3776 1476 3784
rect 1404 3756 1412 3764
rect 1324 3676 1332 3684
rect 2684 3916 2692 3924
rect 3276 3916 3284 3924
rect 3948 3916 3956 3924
rect 4716 3916 4724 3924
rect 1500 3756 1508 3764
rect 1516 3736 1524 3744
rect 1324 3096 1332 3104
rect 1292 2956 1300 2964
rect 1228 2576 1236 2584
rect 1228 2276 1236 2284
rect 1132 1856 1140 1864
rect 1148 1836 1156 1844
rect 1212 1956 1220 1964
rect 1148 1696 1156 1704
rect 1116 1476 1124 1484
rect 1052 916 1060 924
rect 1068 816 1076 824
rect 1004 616 1012 624
rect 812 276 820 284
rect 972 236 980 244
rect 716 176 724 184
rect 956 176 964 184
rect 860 156 868 164
rect 1084 276 1092 284
rect 1052 256 1060 264
rect 1132 1316 1140 1324
rect 1116 1196 1124 1204
rect 1116 676 1124 684
rect 1116 556 1124 564
rect 1164 1456 1172 1464
rect 1228 1856 1236 1864
rect 1180 1356 1188 1364
rect 1164 1316 1172 1324
rect 1324 2696 1332 2704
rect 1356 3136 1364 3144
rect 1356 2936 1364 2944
rect 1340 2616 1348 2624
rect 1324 2576 1332 2584
rect 1324 2496 1332 2504
rect 1308 2276 1316 2284
rect 1340 2116 1348 2124
rect 1324 2076 1332 2084
rect 1340 2076 1348 2084
rect 1292 1916 1300 1924
rect 1324 1856 1332 1864
rect 1324 1776 1332 1784
rect 1324 1476 1332 1484
rect 1452 3536 1460 3544
rect 1372 2656 1380 2664
rect 1372 2556 1380 2564
rect 1612 3776 1620 3784
rect 1660 3776 1668 3784
rect 1836 3716 1844 3724
rect 2092 3876 2100 3884
rect 1948 3776 1956 3784
rect 2268 3696 2276 3704
rect 1708 3536 1716 3544
rect 1548 3356 1556 3364
rect 1516 3136 1524 3144
rect 1420 3096 1428 3104
rect 1452 3096 1460 3104
rect 1532 3056 1540 3064
rect 1516 2976 1524 2984
rect 1612 3316 1620 3324
rect 1580 3116 1588 3124
rect 1628 3076 1636 3084
rect 1404 2696 1412 2704
rect 1548 2696 1556 2704
rect 1404 2676 1412 2684
rect 1420 2596 1428 2604
rect 1420 2336 1428 2344
rect 1420 2276 1428 2284
rect 1388 1816 1396 1824
rect 1516 2596 1524 2604
rect 1484 2536 1492 2544
rect 1500 2496 1508 2504
rect 1484 2296 1492 2304
rect 1372 1716 1380 1724
rect 1308 1356 1316 1364
rect 1340 1296 1348 1304
rect 1276 1136 1284 1144
rect 1308 1096 1316 1104
rect 1276 1076 1284 1084
rect 1260 916 1268 924
rect 1164 816 1172 824
rect 1148 696 1156 704
rect 1260 816 1268 824
rect 1244 776 1252 784
rect 1388 1556 1396 1564
rect 1388 1476 1396 1484
rect 1388 1456 1396 1464
rect 1372 1336 1380 1344
rect 1420 1376 1428 1384
rect 1388 1216 1396 1224
rect 1388 1096 1396 1104
rect 1372 1036 1380 1044
rect 1372 996 1380 1004
rect 1388 956 1396 964
rect 1356 716 1364 724
rect 1276 696 1284 704
rect 1116 536 1124 544
rect 220 136 228 144
rect 684 136 692 144
rect 1116 136 1124 144
rect 428 116 436 124
rect 636 116 644 124
rect 700 116 708 124
rect 796 116 804 124
rect 1164 656 1172 664
rect 1372 316 1380 324
rect 1468 1856 1476 1864
rect 1468 1756 1476 1764
rect 1468 1656 1476 1664
rect 1516 2136 1524 2144
rect 1500 1496 1508 1504
rect 1484 1316 1492 1324
rect 1516 1416 1524 1424
rect 1532 1356 1540 1364
rect 1580 2536 1588 2544
rect 1564 2156 1572 2164
rect 1564 1796 1572 1804
rect 1564 1776 1572 1784
rect 1516 976 1524 984
rect 1468 956 1476 964
rect 1548 936 1556 944
rect 1484 776 1492 784
rect 1500 616 1508 624
rect 1532 596 1540 604
rect 1580 1736 1588 1744
rect 1612 2156 1620 2164
rect 1596 1576 1604 1584
rect 1644 2696 1652 2704
rect 1644 1556 1652 1564
rect 1628 1536 1636 1544
rect 1708 3356 1716 3364
rect 1756 3316 1764 3324
rect 1708 3296 1716 3304
rect 1724 3196 1732 3204
rect 1692 2716 1700 2724
rect 1692 2316 1700 2324
rect 1676 2276 1684 2284
rect 1676 2256 1684 2264
rect 1724 2256 1732 2264
rect 1772 3136 1780 3144
rect 1804 3176 1812 3184
rect 1836 3336 1844 3344
rect 1788 3076 1796 3084
rect 1756 2716 1764 2724
rect 1804 2936 1812 2944
rect 1804 2756 1812 2764
rect 1692 2136 1700 2144
rect 1708 2136 1716 2144
rect 1804 2296 1812 2304
rect 1804 2276 1812 2284
rect 1740 2116 1748 2124
rect 1772 2116 1780 2124
rect 1692 2096 1700 2104
rect 1676 2076 1684 2084
rect 1676 1716 1684 1724
rect 1676 1676 1684 1684
rect 1676 1656 1684 1664
rect 1676 1516 1684 1524
rect 1628 1496 1636 1504
rect 1612 1456 1620 1464
rect 1596 1156 1604 1164
rect 1580 956 1588 964
rect 1564 656 1572 664
rect 1596 676 1604 684
rect 1708 1736 1716 1744
rect 1868 2976 1876 2984
rect 1900 3056 1908 3064
rect 1884 2916 1892 2924
rect 1836 2676 1844 2684
rect 1676 1356 1684 1364
rect 1740 1476 1748 1484
rect 1756 1456 1764 1464
rect 1756 1396 1764 1404
rect 1756 1136 1764 1144
rect 1724 1116 1732 1124
rect 1660 896 1668 904
rect 1708 716 1716 724
rect 1740 596 1748 604
rect 1676 576 1684 584
rect 1628 496 1636 504
rect 2028 3536 2036 3544
rect 2076 3496 2084 3504
rect 1980 3416 1988 3424
rect 1916 2736 1924 2744
rect 1996 3156 2004 3164
rect 1996 2936 2004 2944
rect 1964 2656 1972 2664
rect 1884 2136 1892 2144
rect 1948 2316 1956 2324
rect 1948 2176 1956 2184
rect 2028 3076 2036 3084
rect 2060 3036 2068 3044
rect 2044 2736 2052 2744
rect 2028 2696 2036 2704
rect 2012 2576 2020 2584
rect 2012 2336 2020 2344
rect 1996 2276 2004 2284
rect 1996 2236 2004 2244
rect 2044 2236 2052 2244
rect 2012 2136 2020 2144
rect 2028 2116 2036 2124
rect 1916 1936 1924 1944
rect 1948 1896 1956 1904
rect 1884 1776 1892 1784
rect 1916 1676 1924 1684
rect 1804 1396 1812 1404
rect 1804 1156 1812 1164
rect 1788 1116 1796 1124
rect 1804 1116 1812 1124
rect 1804 1036 1812 1044
rect 1820 1016 1828 1024
rect 1484 336 1492 344
rect 1484 316 1492 324
rect 1324 276 1332 284
rect 1404 256 1412 264
rect 1308 176 1316 184
rect 1164 136 1172 144
rect 1244 136 1252 144
rect 1260 136 1268 144
rect 1372 136 1380 144
rect 1164 116 1172 124
rect 1180 116 1188 124
rect 1532 256 1540 264
rect 1644 256 1652 264
rect 1436 236 1444 244
rect 1724 236 1732 244
rect 1212 96 1220 104
rect 1260 96 1268 104
rect 1340 96 1348 104
rect 1564 136 1572 144
rect 1596 96 1604 104
rect 1948 1476 1956 1484
rect 1884 1136 1892 1144
rect 1916 1136 1924 1144
rect 1948 976 1956 984
rect 1932 536 1940 544
rect 1948 536 1956 544
rect 2156 3536 2164 3544
rect 2268 3396 2276 3404
rect 2156 3376 2164 3384
rect 2380 3896 2388 3904
rect 2796 3896 2804 3904
rect 3724 3896 3732 3904
rect 2412 3876 2420 3884
rect 2748 3876 2756 3884
rect 2924 3876 2932 3884
rect 2348 3696 2356 3704
rect 2796 3756 2804 3764
rect 2268 3336 2276 3344
rect 2140 2936 2148 2944
rect 2124 2656 2132 2664
rect 2124 2636 2132 2644
rect 2124 2316 2132 2324
rect 2188 2676 2196 2684
rect 2204 2656 2212 2664
rect 2156 2276 2164 2284
rect 2124 1836 2132 1844
rect 2092 1756 2100 1764
rect 2028 1496 2036 1504
rect 2044 1476 2052 1484
rect 2124 1816 2132 1824
rect 2092 1356 2100 1364
rect 2012 496 2020 504
rect 1932 276 1940 284
rect 2108 976 2116 984
rect 2284 2916 2292 2924
rect 2252 2676 2260 2684
rect 2220 2156 2228 2164
rect 2252 2576 2260 2584
rect 2284 2156 2292 2164
rect 2620 3356 2628 3364
rect 2396 3096 2404 3104
rect 2364 2936 2372 2944
rect 2364 2676 2372 2684
rect 2636 3336 2644 3344
rect 2476 2716 2484 2724
rect 2444 2676 2452 2684
rect 2556 2676 2564 2684
rect 2412 2536 2420 2544
rect 2156 1776 2164 1784
rect 2188 1816 2196 1824
rect 2172 1476 2180 1484
rect 2284 1916 2292 1924
rect 2300 1856 2308 1864
rect 2348 1856 2356 1864
rect 2268 1776 2276 1784
rect 2284 1736 2292 1744
rect 2204 956 2212 964
rect 2188 936 2196 944
rect 2156 796 2164 804
rect 2092 696 2100 704
rect 2124 676 2132 684
rect 2140 656 2148 664
rect 2204 476 2212 484
rect 2124 316 2132 324
rect 2332 1736 2340 1744
rect 2508 2276 2516 2284
rect 2412 1776 2420 1784
rect 2380 1756 2388 1764
rect 2332 1316 2340 1324
rect 2300 1136 2308 1144
rect 2284 1056 2292 1064
rect 2268 296 2276 304
rect 2124 276 2132 284
rect 2332 956 2340 964
rect 2412 1096 2420 1104
rect 2556 2136 2564 2144
rect 2460 1916 2468 1924
rect 2460 1836 2468 1844
rect 2476 1756 2484 1764
rect 2444 1056 2452 1064
rect 2428 936 2436 944
rect 2380 556 2388 564
rect 2524 1776 2532 1784
rect 2716 3336 2724 3344
rect 2796 3336 2804 3344
rect 2604 2136 2612 2144
rect 2588 2116 2596 2124
rect 2636 2296 2644 2304
rect 2604 2076 2612 2084
rect 2620 1936 2628 1944
rect 2492 1036 2500 1044
rect 2444 656 2452 664
rect 2444 556 2452 564
rect 1804 156 1812 164
rect 1740 136 1748 144
rect 1740 116 1748 124
rect 1948 136 1956 144
rect 2332 136 2340 144
rect 2556 1316 2564 1324
rect 2956 3796 2964 3804
rect 2924 3736 2932 3744
rect 3004 3736 3012 3744
rect 3644 3876 3652 3884
rect 3260 3796 3268 3804
rect 3164 3776 3172 3784
rect 3036 3756 3044 3764
rect 2700 2696 2708 2704
rect 2716 2336 2724 2344
rect 2684 1496 2692 1504
rect 2524 1116 2532 1124
rect 2524 696 2532 704
rect 2524 576 2532 584
rect 2508 476 2516 484
rect 2620 1096 2628 1104
rect 2636 1096 2644 1104
rect 2732 2116 2740 2124
rect 2716 1936 2724 1944
rect 2732 1556 2740 1564
rect 2636 1056 2644 1064
rect 2684 1056 2692 1064
rect 2668 896 2676 904
rect 2556 556 2564 564
rect 2684 656 2692 664
rect 2636 576 2644 584
rect 2636 556 2644 564
rect 2636 536 2644 544
rect 2748 1036 2756 1044
rect 2748 916 2756 924
rect 2908 2996 2916 3004
rect 2876 2956 2884 2964
rect 2988 2916 2996 2924
rect 3132 3736 3140 3744
rect 3100 3356 3108 3364
rect 3020 2676 3028 2684
rect 2988 2556 2996 2564
rect 2908 2536 2916 2544
rect 2876 2336 2884 2344
rect 2876 2176 2884 2184
rect 2828 1876 2836 1884
rect 2956 2156 2964 2164
rect 2924 2136 2932 2144
rect 2924 1856 2932 1864
rect 2988 2136 2996 2144
rect 2972 1896 2980 1904
rect 3052 2656 3060 2664
rect 3036 2536 3044 2544
rect 2892 1736 2900 1744
rect 2828 1716 2836 1724
rect 2796 1496 2804 1504
rect 2716 856 2724 864
rect 2780 836 2788 844
rect 2748 756 2756 764
rect 2700 496 2708 504
rect 2508 316 2516 324
rect 2716 336 2724 344
rect 2812 1096 2820 1104
rect 2796 616 2804 624
rect 2844 1036 2852 1044
rect 2828 976 2836 984
rect 2860 916 2868 924
rect 2860 856 2868 864
rect 2844 336 2852 344
rect 2572 176 2580 184
rect 3036 1716 3044 1724
rect 2988 1556 2996 1564
rect 2956 1476 2964 1484
rect 3068 2516 3076 2524
rect 3068 1496 3076 1504
rect 2956 1076 2964 1084
rect 2988 1076 2996 1084
rect 2892 756 2900 764
rect 3356 3776 3364 3784
rect 3324 3756 3332 3764
rect 3388 3756 3396 3764
rect 3148 2936 3156 2944
rect 3132 2916 3140 2924
rect 3196 2896 3204 2904
rect 3100 1716 3108 1724
rect 3068 1056 3076 1064
rect 3196 2716 3204 2724
rect 3212 2576 3220 2584
rect 3244 3316 3252 3324
rect 3260 3116 3268 3124
rect 3260 2976 3268 2984
rect 3244 2936 3252 2944
rect 3148 1856 3156 1864
rect 3228 2196 3236 2204
rect 3228 2156 3236 2164
rect 3324 3096 3332 3104
rect 3308 3056 3316 3064
rect 3308 2896 3316 2904
rect 3308 2676 3316 2684
rect 3356 3436 3364 3444
rect 3372 3436 3380 3444
rect 3356 3116 3364 3124
rect 3356 3076 3364 3084
rect 3356 3036 3364 3044
rect 3340 2976 3348 2984
rect 3436 3356 3444 3364
rect 3420 3296 3428 3304
rect 3468 3316 3476 3324
rect 3468 3136 3476 3144
rect 3500 3316 3508 3324
rect 3548 3096 3556 3104
rect 3500 3076 3508 3084
rect 3340 2876 3348 2884
rect 3356 2776 3364 2784
rect 3324 2556 3332 2564
rect 3292 2476 3300 2484
rect 3308 2196 3316 2204
rect 3308 2116 3316 2124
rect 3164 1496 3172 1504
rect 3148 1456 3156 1464
rect 3164 1276 3172 1284
rect 3052 876 3060 884
rect 3068 796 3076 804
rect 2940 176 2948 184
rect 2860 136 2868 144
rect 2876 136 2884 144
rect 2348 116 2356 124
rect 2108 96 2116 104
rect 2252 96 2260 104
rect 3100 156 3108 164
rect 2972 136 2980 144
rect 3148 616 3156 624
rect 3212 1296 3220 1304
rect 3292 1516 3300 1524
rect 3260 1496 3268 1504
rect 3324 1476 3332 1484
rect 3292 1456 3300 1464
rect 3292 1296 3300 1304
rect 3276 1116 3284 1124
rect 3228 936 3236 944
rect 3212 836 3220 844
rect 3260 676 3268 684
rect 3164 596 3172 604
rect 3196 596 3204 604
rect 3132 276 3140 284
rect 3260 256 3268 264
rect 3244 236 3252 244
rect 3452 2976 3460 2984
rect 3468 2896 3476 2904
rect 3404 2876 3412 2884
rect 3468 2756 3476 2764
rect 3404 2116 3412 2124
rect 3388 2076 3396 2084
rect 3372 1996 3380 2004
rect 3596 3776 3604 3784
rect 3580 3376 3588 3384
rect 3580 2956 3588 2964
rect 3532 2876 3540 2884
rect 3500 2636 3508 2644
rect 3516 2556 3524 2564
rect 3468 2476 3476 2484
rect 3404 1856 3412 1864
rect 3372 1836 3380 1844
rect 3388 936 3396 944
rect 3500 2296 3508 2304
rect 3516 2036 3524 2044
rect 3452 1516 3460 1524
rect 3468 1516 3476 1524
rect 3468 1396 3476 1404
rect 3612 3296 3620 3304
rect 3612 3156 3620 3164
rect 3820 3896 3828 3904
rect 3884 3876 3892 3884
rect 4124 3876 4132 3884
rect 3740 3756 3748 3764
rect 3772 3716 3780 3724
rect 3724 3376 3732 3384
rect 3660 3356 3668 3364
rect 3660 3336 3668 3344
rect 3628 2676 3636 2684
rect 3596 2656 3604 2664
rect 3580 2596 3588 2604
rect 3628 2496 3636 2504
rect 3596 2296 3604 2304
rect 3660 3056 3668 3064
rect 3660 2636 3668 2644
rect 3708 3016 3716 3024
rect 3692 2916 3700 2924
rect 3756 3076 3764 3084
rect 3740 2956 3748 2964
rect 3740 2856 3748 2864
rect 3836 3456 3844 3464
rect 3820 3436 3828 3444
rect 3804 3196 3812 3204
rect 3804 3156 3812 3164
rect 3788 3036 3796 3044
rect 3740 2696 3748 2704
rect 3772 2696 3780 2704
rect 3724 2676 3732 2684
rect 3724 2656 3732 2664
rect 3724 2536 3732 2544
rect 3724 2476 3732 2484
rect 3660 2136 3668 2144
rect 3676 1896 3684 1904
rect 3580 1756 3588 1764
rect 3548 1416 3556 1424
rect 3532 1396 3540 1404
rect 3596 1516 3604 1524
rect 3580 1376 3588 1384
rect 3612 1376 3620 1384
rect 3564 1136 3572 1144
rect 3452 1096 3460 1104
rect 3484 1056 3492 1064
rect 3388 796 3396 804
rect 3308 556 3316 564
rect 3452 556 3460 564
rect 3404 516 3412 524
rect 3308 276 3316 284
rect 3244 136 3252 144
rect 3324 256 3332 264
rect 3516 836 3524 844
rect 3660 1456 3668 1464
rect 3660 1396 3668 1404
rect 3708 2336 3716 2344
rect 3708 2236 3716 2244
rect 3724 2116 3732 2124
rect 3708 2096 3716 2104
rect 3708 2056 3716 2064
rect 3724 1656 3732 1664
rect 3724 1596 3732 1604
rect 3724 1576 3732 1584
rect 3724 1496 3732 1504
rect 3708 1356 3716 1364
rect 3772 2676 3780 2684
rect 4028 3796 4036 3804
rect 4108 3796 4116 3804
rect 3916 3716 3924 3724
rect 3932 3716 3940 3724
rect 3964 3696 3972 3704
rect 4012 3536 4020 3544
rect 4028 3516 4036 3524
rect 4028 3496 4036 3504
rect 3900 3476 3908 3484
rect 3916 3456 3924 3464
rect 3980 3456 3988 3464
rect 3980 3376 3988 3384
rect 4092 3516 4100 3524
rect 4092 3456 4100 3464
rect 4108 3456 4116 3464
rect 4076 3336 4084 3344
rect 4092 3316 4100 3324
rect 4060 3296 4068 3304
rect 4044 3116 4052 3124
rect 3868 2936 3876 2944
rect 3852 2696 3860 2704
rect 3772 2516 3780 2524
rect 3740 1056 3748 1064
rect 3804 2296 3812 2304
rect 3836 2296 3844 2304
rect 3884 2536 3892 2544
rect 3772 1496 3780 1504
rect 3820 2116 3828 2124
rect 3980 3016 3988 3024
rect 4060 2936 4068 2944
rect 3964 2656 3972 2664
rect 3932 2536 3940 2544
rect 3980 2516 3988 2524
rect 4060 2716 4068 2724
rect 4060 2696 4068 2704
rect 3820 1756 3828 1764
rect 3740 916 3748 924
rect 3660 676 3668 684
rect 3724 656 3732 664
rect 3516 616 3524 624
rect 3500 516 3508 524
rect 3644 536 3652 544
rect 3580 376 3588 384
rect 3724 296 3732 304
rect 3564 236 3572 244
rect 3692 236 3700 244
rect 3628 216 3636 224
rect 3788 1116 3796 1124
rect 3804 1116 3812 1124
rect 3804 1076 3812 1084
rect 3836 756 3844 764
rect 3820 716 3828 724
rect 3852 696 3860 704
rect 3804 676 3812 684
rect 3788 316 3796 324
rect 3884 1356 3892 1364
rect 4028 2256 4036 2264
rect 3964 2076 3972 2084
rect 4060 2636 4068 2644
rect 4012 1856 4020 1864
rect 3980 1516 3988 1524
rect 3996 1476 4004 1484
rect 3964 1456 3972 1464
rect 3948 1376 3956 1384
rect 3948 1336 3956 1344
rect 3948 1256 3956 1264
rect 3948 1076 3956 1084
rect 3916 916 3924 924
rect 3964 736 3972 744
rect 3948 676 3956 684
rect 3932 636 3940 644
rect 3900 516 3908 524
rect 3948 556 3956 564
rect 3932 316 3940 324
rect 3772 256 3780 264
rect 3868 296 3876 304
rect 3884 296 3892 304
rect 3884 256 3892 264
rect 3932 256 3940 264
rect 3836 236 3844 244
rect 3516 176 3524 184
rect 3788 176 3796 184
rect 3980 676 3988 684
rect 4012 1356 4020 1364
rect 4012 1156 4020 1164
rect 4044 1076 4052 1084
rect 4076 2576 4084 2584
rect 4108 3056 4116 3064
rect 4108 2276 4116 2284
rect 4108 2176 4116 2184
rect 4108 2156 4116 2164
rect 4108 1976 4116 1984
rect 4092 1836 4100 1844
rect 4092 1776 4100 1784
rect 4108 1756 4116 1764
rect 4156 3156 4164 3164
rect 4476 3776 4484 3784
rect 4300 3756 4308 3764
rect 4332 3736 4340 3744
rect 4284 3696 4292 3704
rect 4236 3516 4244 3524
rect 4284 3516 4292 3524
rect 4188 3476 4196 3484
rect 4172 2976 4180 2984
rect 4156 2676 4164 2684
rect 4156 2356 4164 2364
rect 4284 3436 4292 3444
rect 4204 3336 4212 3344
rect 4204 2916 4212 2924
rect 4204 2756 4212 2764
rect 4236 2676 4244 2684
rect 4236 2536 4244 2544
rect 4204 2296 4212 2304
rect 4236 2236 4244 2244
rect 4236 1936 4244 1944
rect 4140 1876 4148 1884
rect 4124 1536 4132 1544
rect 4156 1456 4164 1464
rect 4172 1416 4180 1424
rect 4284 2736 4292 2744
rect 4284 2336 4292 2344
rect 4284 2316 4292 2324
rect 4268 2296 4276 2304
rect 4380 3696 4388 3704
rect 4444 3696 4452 3704
rect 4508 3536 4516 3544
rect 4460 3496 4468 3504
rect 4444 3376 4452 3384
rect 4364 3356 4372 3364
rect 4380 3156 4388 3164
rect 4316 3096 4324 3104
rect 4332 3096 4340 3104
rect 4332 2916 4340 2924
rect 4316 2356 4324 2364
rect 4332 2356 4340 2364
rect 4412 2936 4420 2944
rect 4396 2696 4404 2704
rect 4412 2676 4420 2684
rect 4332 2336 4340 2344
rect 4284 2116 4292 2124
rect 4236 1776 4244 1784
rect 4252 1776 4260 1784
rect 4220 1536 4228 1544
rect 4124 1316 4132 1324
rect 3980 576 3988 584
rect 3964 336 3972 344
rect 3964 296 3972 304
rect 4028 756 4036 764
rect 4060 656 4068 664
rect 4092 676 4100 684
rect 4156 1296 4164 1304
rect 4124 1116 4132 1124
rect 4108 656 4116 664
rect 4076 616 4084 624
rect 3996 336 4004 344
rect 3756 156 3764 164
rect 3324 136 3332 144
rect 4060 256 4068 264
rect 4140 636 4148 644
rect 4204 1256 4212 1264
rect 4284 1756 4292 1764
rect 4236 1296 4244 1304
rect 4220 1116 4228 1124
rect 4220 916 4228 924
rect 4220 876 4228 884
rect 4172 836 4180 844
rect 4188 776 4196 784
rect 4188 756 4196 764
rect 4204 756 4212 764
rect 4172 736 4180 744
rect 4332 2216 4340 2224
rect 4332 1896 4340 1904
rect 4300 1716 4308 1724
rect 4204 676 4212 684
rect 4236 676 4244 684
rect 4236 596 4244 604
rect 4364 2116 4372 2124
rect 4348 1736 4356 1744
rect 4332 1476 4340 1484
rect 4348 1396 4356 1404
rect 4316 1316 4324 1324
rect 4332 1096 4340 1104
rect 4316 1056 4324 1064
rect 4300 916 4308 924
rect 4284 876 4292 884
rect 4284 736 4292 744
rect 4364 1116 4372 1124
rect 4284 696 4292 704
rect 4268 676 4276 684
rect 4252 576 4260 584
rect 4188 556 4196 564
rect 4236 556 4244 564
rect 4220 536 4228 544
rect 4204 496 4212 504
rect 4236 516 4244 524
rect 4156 216 4164 224
rect 4236 256 4244 264
rect 4348 656 4356 664
rect 4428 2516 4436 2524
rect 4444 2496 4452 2504
rect 4492 3356 4500 3364
rect 4508 3276 4516 3284
rect 4508 2956 4516 2964
rect 4668 3476 4676 3484
rect 4652 3416 4660 3424
rect 4652 3356 4660 3364
rect 4636 3336 4644 3344
rect 4588 3136 4596 3144
rect 4604 3136 4612 3144
rect 4556 3116 4564 3124
rect 4572 3116 4580 3124
rect 4540 2776 4548 2784
rect 4476 2656 4484 2664
rect 4540 2656 4548 2664
rect 4636 2936 4644 2944
rect 4732 3736 4740 3744
rect 5004 3776 5012 3784
rect 4812 3716 4820 3724
rect 4748 3476 4756 3484
rect 4748 3376 4756 3384
rect 4684 3356 4692 3364
rect 4716 3356 4724 3364
rect 4780 3336 4788 3344
rect 4668 2736 4676 2744
rect 4700 3116 4708 3124
rect 4732 2996 4740 3004
rect 4748 2936 4756 2944
rect 4732 2736 4740 2744
rect 4700 2656 4708 2664
rect 4556 2636 4564 2644
rect 4556 2616 4564 2624
rect 4604 2596 4612 2604
rect 4668 2576 4676 2584
rect 4556 2476 4564 2484
rect 4572 2476 4580 2484
rect 4572 2316 4580 2324
rect 4412 2116 4420 2124
rect 4428 2116 4436 2124
rect 4444 1836 4452 1844
rect 4444 1756 4452 1764
rect 4428 1696 4436 1704
rect 4572 2276 4580 2284
rect 4476 2156 4484 2164
rect 4572 2136 4580 2144
rect 4476 2116 4484 2124
rect 4540 2116 4548 2124
rect 4620 1916 4628 1924
rect 4652 2256 4660 2264
rect 4668 2076 4676 2084
rect 4652 1916 4660 1924
rect 4620 1776 4628 1784
rect 4492 1536 4500 1544
rect 4540 1536 4548 1544
rect 4524 1516 4532 1524
rect 4572 1496 4580 1504
rect 4508 1456 4516 1464
rect 4444 876 4452 884
rect 4380 736 4388 744
rect 4364 536 4372 544
rect 4284 516 4292 524
rect 4332 516 4340 524
rect 4268 236 4276 244
rect 4396 316 4404 324
rect 4364 276 4372 284
rect 4348 256 4356 264
rect 4316 216 4324 224
rect 4476 876 4484 884
rect 4540 936 4548 944
rect 4604 1316 4612 1324
rect 4540 676 4548 684
rect 4668 1736 4676 1744
rect 4652 1536 4660 1544
rect 4652 1516 4660 1524
rect 4652 1116 4660 1124
rect 4588 556 4596 564
rect 4572 496 4580 504
rect 4508 296 4516 304
rect 4604 256 4612 264
rect 4476 176 4484 184
rect 4540 176 4548 184
rect 4300 116 4308 124
rect 4364 116 4372 124
rect 4524 96 4532 104
rect 4556 96 4564 104
rect 3852 76 3860 84
rect 4588 76 4596 84
rect 4828 3056 4836 3064
rect 4860 3296 4868 3304
rect 4876 3296 4884 3304
rect 4860 3096 4868 3104
rect 4860 2936 4868 2944
rect 4812 2716 4820 2724
rect 4764 2536 4772 2544
rect 4732 1876 4740 1884
rect 4732 1716 4740 1724
rect 4780 2496 4788 2504
rect 4812 2476 4820 2484
rect 4812 2276 4820 2284
rect 4780 2256 4788 2264
rect 4796 2236 4804 2244
rect 4780 1936 4788 1944
rect 4780 1596 4788 1604
rect 4748 1316 4756 1324
rect 4764 1156 4772 1164
rect 4700 1136 4708 1144
rect 4748 1096 4756 1104
rect 4700 996 4708 1004
rect 4668 576 4676 584
rect 4732 936 4740 944
rect 4748 876 4756 884
rect 4748 796 4756 804
rect 4764 676 4772 684
rect 4860 2336 4868 2344
rect 4860 2236 4868 2244
rect 4844 2196 4852 2204
rect 4828 2156 4836 2164
rect 4844 1696 4852 1704
rect 4812 1536 4820 1544
rect 4828 1476 4836 1484
rect 4812 1236 4820 1244
rect 4812 1116 4820 1124
rect 4796 876 4804 884
rect 4940 3456 4948 3464
rect 4956 3436 4964 3444
rect 4940 3376 4948 3384
rect 4924 3316 4932 3324
rect 4924 3076 4932 3084
rect 4924 2936 4932 2944
rect 4908 2696 4916 2704
rect 4924 2556 4932 2564
rect 4924 2536 4932 2544
rect 4924 2496 4932 2504
rect 4908 2196 4916 2204
rect 4908 2136 4916 2144
rect 4908 1916 4916 1924
rect 4908 1836 4916 1844
rect 4876 1056 4884 1064
rect 4796 716 4804 724
rect 4908 1596 4916 1604
rect 4972 3136 4980 3144
rect 5180 3776 5188 3784
rect 5132 3736 5140 3744
rect 5196 3736 5204 3744
rect 5020 3496 5028 3504
rect 5164 3476 5172 3484
rect 5084 3416 5092 3424
rect 5132 3396 5140 3404
rect 5132 3376 5140 3384
rect 5052 3096 5060 3104
rect 5084 3056 5092 3064
rect 5052 3036 5060 3044
rect 4956 2316 4964 2324
rect 4956 2156 4964 2164
rect 4940 1696 4948 1704
rect 4940 1516 4948 1524
rect 5052 2916 5060 2924
rect 5020 2736 5028 2744
rect 5020 2616 5028 2624
rect 4988 2556 4996 2564
rect 4988 2536 4996 2544
rect 5004 2516 5012 2524
rect 5036 2516 5044 2524
rect 5004 2176 5012 2184
rect 4988 2116 4996 2124
rect 5036 2156 5044 2164
rect 5036 2096 5044 2104
rect 5036 1996 5044 2004
rect 5004 1776 5012 1784
rect 4972 1656 4980 1664
rect 4972 1536 4980 1544
rect 4972 1476 4980 1484
rect 4972 1276 4980 1284
rect 4972 1116 4980 1124
rect 4956 1056 4964 1064
rect 4940 716 4948 724
rect 4860 656 4868 664
rect 4876 576 4884 584
rect 5052 1756 5060 1764
rect 5132 3096 5140 3104
rect 5164 2956 5172 2964
rect 5116 2396 5124 2404
rect 5116 2316 5124 2324
rect 5164 2556 5172 2564
rect 5196 3356 5204 3364
rect 5100 2156 5108 2164
rect 5116 2156 5124 2164
rect 5180 2156 5188 2164
rect 5148 2036 5156 2044
rect 5100 1856 5108 1864
rect 5068 1536 5076 1544
rect 5036 1516 5044 1524
rect 5036 1116 5044 1124
rect 5068 1096 5076 1104
rect 5036 976 5044 984
rect 5180 1776 5188 1784
rect 5068 756 5076 764
rect 5036 736 5044 744
rect 5036 696 5044 704
rect 5052 676 5060 684
rect 5020 316 5028 324
rect 4828 296 4836 304
rect 4924 256 4932 264
rect 4876 196 4884 204
rect 5164 1156 5172 1164
rect 5164 1056 5172 1064
rect 5132 916 5140 924
rect 5116 696 5124 704
rect 5100 656 5108 664
rect 5244 3776 5252 3784
rect 5244 3756 5252 3764
rect 5276 2576 5284 2584
rect 5260 2236 5268 2244
rect 5228 2176 5236 2184
rect 5244 1956 5252 1964
rect 5244 1716 5252 1724
rect 5308 3836 5316 3844
rect 5244 1096 5252 1104
rect 5260 876 5268 884
rect 5244 156 5252 164
rect 5308 1776 5316 1784
rect 5308 1736 5316 1744
rect 5292 1536 5300 1544
rect 5340 3756 5348 3764
rect 5404 3116 5412 3124
rect 5388 2676 5396 2684
rect 5404 2076 5412 2084
rect 5372 1756 5380 1764
rect 5324 1336 5332 1344
rect 5292 1096 5300 1104
rect 5292 536 5300 544
rect 5276 316 5284 324
rect 5292 296 5300 304
rect 5356 1376 5364 1384
rect 5388 976 5396 984
rect 5404 916 5412 924
rect 5388 696 5396 704
rect 5372 556 5380 564
rect 5452 2216 5460 2224
rect 5484 2696 5492 2704
rect 5516 2316 5524 2324
rect 5484 2136 5492 2144
rect 5516 1876 5524 1884
rect 5532 1496 5540 1504
rect 5452 136 5460 144
<< metal5 >>
rect 2692 3917 3276 3923
rect 3956 3917 4716 3923
rect 2388 3897 2796 3903
rect 3732 3897 3820 3903
rect 2100 3877 2412 3883
rect 2756 3877 2924 3883
rect 3652 3877 3884 3883
rect 3892 3877 4124 3883
rect 5309 3844 5315 3855
rect 2964 3797 3260 3803
rect 4036 3797 4108 3803
rect 708 3777 780 3783
rect 980 3777 1084 3783
rect 1476 3777 1612 3783
rect 1668 3777 1948 3783
rect 3172 3777 3356 3783
rect 3604 3777 4476 3783
rect 4484 3777 5004 3783
rect 5012 3777 5180 3783
rect 820 3757 892 3763
rect 1412 3757 1500 3763
rect 2804 3757 3036 3763
rect 3332 3757 3388 3763
rect 3748 3757 4300 3763
rect 4308 3757 5244 3763
rect 484 3737 524 3743
rect 772 3737 860 3743
rect 1284 3737 1516 3743
rect 2932 3737 3004 3743
rect 3140 3737 4332 3743
rect 4357 3737 4732 3743
rect 5140 3737 5196 3743
rect 292 3717 556 3723
rect 564 3717 1836 3723
rect 3780 3717 3916 3723
rect 3940 3717 4812 3723
rect 2276 3697 2348 3703
rect 3972 3697 4267 3703
rect 4292 3697 4380 3703
rect 4405 3697 4444 3703
rect 1188 3677 1324 3683
rect 468 3537 1212 3543
rect 1460 3537 1708 3543
rect 2036 3537 2156 3543
rect 4020 3537 4508 3543
rect 644 3517 764 3523
rect 4036 3517 4092 3523
rect 4244 3517 4284 3523
rect 724 3497 828 3503
rect 1060 3497 2076 3503
rect 4036 3497 4460 3503
rect 4468 3497 5020 3503
rect 3908 3477 4188 3483
rect 4756 3477 5164 3483
rect 3844 3457 3916 3463
rect 3988 3457 4092 3463
rect 4116 3457 4940 3463
rect 3364 3437 3372 3443
rect 3380 3437 3820 3443
rect 3828 3437 4284 3443
rect 4292 3437 4956 3443
rect 893 3424 899 3435
rect 4660 3417 5084 3423
rect 2181 3397 2268 3403
rect 5125 3397 5132 3403
rect 1300 3377 2156 3383
rect 3732 3377 3980 3383
rect 4452 3377 4748 3383
rect 4948 3377 5132 3383
rect 3581 3365 3587 3376
rect 1092 3357 1548 3363
rect 1716 3357 2620 3363
rect 3108 3357 3436 3363
rect 3668 3357 3675 3363
rect 4372 3357 4492 3363
rect 4660 3357 4684 3363
rect 4724 3357 5196 3363
rect 196 3337 316 3343
rect 388 3337 1836 3343
rect 1861 3337 2268 3343
rect 2644 3337 2716 3343
rect 2804 3337 3660 3343
rect 4084 3337 4204 3343
rect 4644 3337 4780 3343
rect 772 3317 1260 3323
rect 1620 3317 1756 3323
rect 3252 3317 3468 3323
rect 3508 3317 4092 3323
rect 4100 3317 4123 3323
rect 4925 3324 4931 3335
rect 1716 3297 1723 3303
rect 3428 3297 3612 3303
rect 4068 3297 4860 3303
rect 4884 3297 4891 3303
rect 4101 3277 4508 3283
rect 1085 3225 1091 3236
rect 1725 3183 1731 3196
rect 1725 3177 1804 3183
rect 1236 3157 1996 3163
rect 3620 3157 3804 3163
rect 4164 3157 4380 3163
rect 1349 3137 1356 3143
rect 1524 3137 1772 3143
rect 3476 3137 4588 3143
rect 4612 3137 4972 3143
rect 532 3117 1580 3123
rect 3268 3117 3356 3123
rect 4052 3117 4556 3123
rect 4580 3117 4700 3123
rect 4741 3117 5404 3123
rect 100 3097 540 3103
rect 756 3097 860 3103
rect 877 3097 1100 3103
rect 132 3077 252 3083
rect 877 3083 883 3097
rect 1268 3097 1307 3103
rect 1332 3097 1420 3103
rect 1460 3097 2396 3103
rect 3332 3097 3548 3103
rect 3653 3097 4316 3103
rect 4340 3097 4860 3103
rect 5060 3097 5132 3103
rect 772 3077 883 3083
rect 1044 3077 1628 3083
rect 1796 3077 2028 3083
rect 3364 3077 3500 3083
rect 3508 3077 3756 3083
rect 3764 3077 4924 3083
rect 1140 3057 1339 3063
rect 1540 3057 1900 3063
rect 3316 3057 3643 3063
rect 3668 3057 4108 3063
rect 4836 3057 5084 3063
rect 580 3037 1164 3043
rect 1188 3037 2060 3043
rect 3364 3037 3788 3043
rect 4997 3037 5052 3043
rect 308 3017 460 3023
rect 468 3017 1084 3023
rect 3685 3017 3708 3023
rect 3988 3017 4091 3023
rect 2916 2997 2939 3003
rect 132 2977 988 2983
rect 1284 2977 1307 2983
rect 3261 2984 3267 2995
rect 1524 2977 1868 2983
rect 3268 2977 3323 2983
rect 3348 2977 3452 2983
rect 3460 2977 4172 2983
rect 388 2957 1292 2963
rect 2884 2957 3580 2963
rect 3621 2957 3740 2963
rect 4516 2957 5164 2963
rect 532 2937 1356 2943
rect 1812 2937 1996 2943
rect 2148 2937 2364 2943
rect 3156 2937 3227 2943
rect 3252 2937 3868 2943
rect 4068 2937 4412 2943
rect 4644 2937 4748 2943
rect 4868 2937 4924 2943
rect 932 2917 1084 2923
rect 1156 2917 1196 2923
rect 1892 2917 2284 2923
rect 2996 2917 3132 2923
rect 3140 2917 3692 2923
rect 4212 2917 4332 2923
rect 5060 2917 5115 2923
rect 276 2897 364 2903
rect 3204 2897 3308 2903
rect 3333 2897 3468 2903
rect 3348 2877 3404 2883
rect 3540 2877 3643 2883
rect 3748 2857 3771 2863
rect 788 2797 795 2803
rect 1204 2777 1211 2783
rect 3364 2777 4540 2783
rect 925 2745 931 2756
rect 1029 2757 1196 2763
rect 1812 2757 1819 2763
rect 3476 2757 4204 2763
rect 4292 2737 4668 2743
rect 4740 2737 5020 2743
rect 932 2717 1100 2723
rect 1700 2717 1756 2723
rect 1764 2717 2476 2723
rect 4068 2717 4812 2723
rect 564 2697 732 2703
rect 788 2697 1052 2703
rect 1060 2697 1132 2703
rect 1317 2697 1324 2703
rect 1412 2697 1548 2703
rect 1652 2697 2028 2703
rect 2036 2697 2700 2703
rect 3685 2697 3740 2703
rect 3780 2697 3852 2703
rect 4068 2697 4396 2703
rect 4916 2697 5484 2703
rect 580 2677 668 2683
rect 868 2677 955 2683
rect 996 2677 1404 2683
rect 1844 2677 2188 2683
rect 2260 2677 2364 2683
rect 2452 2677 2556 2683
rect 3028 2677 3308 2683
rect 3316 2677 3628 2683
rect 3732 2677 3772 2683
rect 4164 2677 4236 2683
rect 4420 2677 5388 2683
rect 852 2657 1052 2663
rect 1076 2657 1372 2663
rect 1380 2657 1964 2663
rect 2132 2657 2204 2663
rect 3060 2657 3596 2663
rect 3732 2657 3964 2663
rect 3972 2657 4476 2663
rect 4548 2657 4700 2663
rect 805 2637 923 2643
rect 1221 2637 2124 2643
rect 3508 2637 3660 2643
rect 3668 2637 3739 2643
rect 4068 2637 4556 2643
rect 516 2617 1340 2623
rect 4564 2617 5020 2623
rect 1428 2597 1516 2603
rect 3588 2597 4604 2603
rect 1236 2577 1243 2583
rect 1332 2577 1627 2583
rect 2020 2577 2252 2583
rect 3205 2577 3212 2583
rect 3749 2577 4076 2583
rect 4453 2577 4668 2583
rect 4676 2577 5276 2583
rect 132 2557 636 2563
rect 676 2557 1372 2563
rect 2996 2557 3324 2563
rect 3524 2557 4571 2563
rect 4581 2557 4924 2563
rect 4996 2557 5164 2563
rect 788 2537 1052 2543
rect 1349 2537 1467 2543
rect 1477 2537 1484 2543
rect 1588 2537 2412 2543
rect 2916 2537 3036 2543
rect 3732 2537 3867 2543
rect 3892 2537 3932 2543
rect 4244 2537 4764 2543
rect 4932 2537 4988 2543
rect 3076 2517 3772 2523
rect 3909 2517 3980 2523
rect 4436 2517 5004 2523
rect 5012 2517 5036 2523
rect 1332 2497 1500 2503
rect 3636 2497 4444 2503
rect 4773 2497 4780 2503
rect 4932 2497 5083 2503
rect 3300 2477 3468 2483
rect 3732 2477 4556 2483
rect 4580 2477 4812 2483
rect 5093 2397 5116 2403
rect 4164 2357 4316 2363
rect 4340 2357 4347 2363
rect 1381 2337 1420 2343
rect 1428 2337 2012 2343
rect 2724 2337 2876 2343
rect 3653 2337 3708 2343
rect 4340 2337 4860 2343
rect 900 2317 972 2323
rect 1700 2317 1851 2323
rect 1956 2317 2124 2323
rect 4292 2317 4572 2323
rect 4964 2317 5116 2323
rect 5349 2317 5516 2323
rect 692 2297 812 2303
rect 820 2297 1484 2303
rect 1812 2297 2636 2303
rect 3508 2297 3596 2303
rect 3844 2297 4204 2303
rect 4276 2297 4347 2303
rect 3805 2285 3811 2296
rect 1172 2277 1228 2283
rect 1316 2277 1420 2283
rect 1684 2277 1804 2283
rect 1861 2277 1996 2283
rect 2164 2277 2508 2283
rect 4116 2277 4572 2283
rect 4580 2277 4812 2283
rect 1684 2257 1724 2263
rect 4036 2257 4443 2263
rect 4660 2257 4780 2263
rect 2004 2237 2044 2243
rect 3716 2237 4236 2243
rect 4804 2237 4860 2243
rect 4868 2237 5260 2243
rect 4340 2217 5452 2223
rect 3236 2197 3308 2203
rect 4852 2197 4908 2203
rect 964 2177 1948 2183
rect 2884 2177 4108 2183
rect 5012 2177 5228 2183
rect 900 2157 972 2163
rect 1044 2157 1564 2163
rect 1620 2157 2220 2163
rect 2292 2157 2299 2163
rect 2964 2157 3228 2163
rect 4101 2157 4108 2163
rect 4484 2157 4828 2163
rect 5044 2157 5100 2163
rect 5124 2157 5180 2163
rect 180 2137 396 2143
rect 484 2137 620 2143
rect 637 2137 1516 2143
rect 325 2117 348 2123
rect 637 2123 643 2137
rect 1716 2137 1884 2143
rect 2020 2137 2043 2143
rect 2564 2137 2604 2143
rect 2932 2137 2988 2143
rect 3668 2137 4572 2143
rect 4916 2137 5484 2143
rect 452 2117 643 2123
rect 740 2117 780 2123
rect 1156 2117 1340 2123
rect 1348 2117 1740 2123
rect 1780 2117 1851 2123
rect 1861 2117 2028 2123
rect 2596 2117 2732 2123
rect 3316 2117 3404 2123
rect 3732 2117 3820 2123
rect 4292 2117 4364 2123
rect 4372 2117 4412 2123
rect 4436 2117 4476 2123
rect 4548 2117 4988 2123
rect 356 2097 1020 2103
rect 1140 2097 1692 2103
rect 4965 2097 5036 2103
rect 756 2077 940 2083
rect 948 2077 1211 2083
rect 1332 2077 1340 2083
rect 1348 2077 1659 2083
rect 1684 2077 2604 2083
rect 3396 2077 3964 2083
rect 4676 2077 5404 2083
rect 3716 2057 3771 2063
rect 3524 2037 5148 2043
rect 852 1997 859 2003
rect 3380 1997 4923 2003
rect 4933 1997 5036 2003
rect 820 1977 827 1983
rect 4116 1977 4123 1983
rect 436 1957 1212 1963
rect 5252 1957 5275 1963
rect 884 1937 1052 1943
rect 1060 1937 1916 1943
rect 2628 1937 2716 1943
rect 4244 1937 4780 1943
rect 468 1917 764 1923
rect 964 1917 1292 1923
rect 2292 1917 2460 1923
rect 4628 1917 4652 1923
rect 4916 1917 4987 1923
rect 837 1897 876 1903
rect 948 1897 1948 1903
rect 2980 1897 3676 1903
rect 3684 1897 4332 1903
rect 2836 1877 4140 1883
rect 4740 1877 5516 1883
rect 676 1857 859 1863
rect 1140 1857 1228 1863
rect 1332 1857 1468 1863
rect 2308 1857 2348 1863
rect 2932 1857 3148 1863
rect 3412 1857 4012 1863
rect 4965 1857 5100 1863
rect 596 1837 684 1843
rect 1044 1837 1148 1843
rect 2132 1837 2460 1843
rect 3380 1837 4092 1843
rect 4452 1837 4908 1843
rect 1396 1817 1403 1823
rect 2132 1817 2188 1823
rect 964 1797 1083 1803
rect 900 1777 972 1783
rect 1332 1777 1564 1783
rect 1572 1777 1884 1783
rect 2164 1777 2268 1783
rect 2420 1777 2524 1783
rect 4100 1777 4123 1783
rect 4244 1777 4252 1783
rect 4260 1777 4620 1783
rect 4628 1777 5004 1783
rect 5188 1777 5308 1783
rect 804 1757 844 1763
rect 1476 1757 1651 1763
rect 996 1737 1580 1743
rect 1645 1743 1651 1757
rect 1669 1757 2092 1763
rect 2388 1757 2476 1763
rect 3588 1757 3820 1763
rect 3828 1757 4108 1763
rect 4292 1757 4444 1763
rect 4557 1757 5052 1763
rect 1645 1737 1708 1743
rect 2292 1737 2332 1743
rect 2340 1737 2892 1743
rect 4557 1743 4563 1757
rect 5285 1757 5372 1763
rect 4356 1737 4563 1743
rect 4581 1737 4668 1743
rect 4676 1737 5308 1743
rect 645 1717 652 1723
rect 772 1717 988 1723
rect 1380 1717 1676 1723
rect 2836 1717 3036 1723
rect 3044 1717 3100 1723
rect 4308 1717 4732 1723
rect 5252 1717 5275 1723
rect 804 1697 1148 1703
rect 4436 1697 4844 1703
rect 4948 1697 4955 1703
rect 500 1677 1371 1683
rect 1684 1677 1916 1683
rect 1684 1657 1691 1663
rect 3732 1657 3771 1663
rect 4980 1657 4987 1663
rect 3732 1597 3739 1603
rect 4788 1597 4795 1603
rect 4901 1597 4908 1603
rect 3685 1577 3724 1583
rect 1381 1557 1388 1563
rect 1652 1557 1659 1563
rect 2740 1557 2988 1563
rect 756 1537 1628 1543
rect 4132 1537 4220 1543
rect 4500 1537 4540 1543
rect 4548 1537 4652 1543
rect 4820 1537 4972 1543
rect 5076 1537 5292 1543
rect 868 1517 1676 1523
rect 3300 1517 3452 1523
rect 3476 1517 3596 1523
rect 3988 1517 4524 1523
rect 4660 1517 4940 1523
rect 4948 1517 5036 1523
rect 580 1497 1500 1503
rect 1636 1497 2028 1503
rect 2692 1497 2796 1503
rect 3076 1497 3164 1503
rect 3172 1497 3260 1503
rect 3732 1497 3772 1503
rect 4580 1497 5532 1503
rect 901 1477 1116 1483
rect 1332 1477 1388 1483
rect 1748 1477 1948 1483
rect 2052 1477 2172 1483
rect 2964 1477 3324 1483
rect 3973 1477 3996 1483
rect 4340 1477 4828 1483
rect 4836 1477 4972 1483
rect 964 1457 1147 1463
rect 1157 1457 1164 1463
rect 1396 1457 1612 1463
rect 1669 1457 1756 1463
rect 3156 1457 3292 1463
rect 3668 1457 3964 1463
rect 4164 1457 4508 1463
rect 1524 1417 1531 1423
rect 3556 1417 4172 1423
rect 1764 1397 1804 1403
rect 3476 1397 3532 1403
rect 3668 1397 4348 1403
rect 1044 1377 1420 1383
rect 1428 1377 1435 1383
rect 3588 1377 3612 1383
rect 3781 1377 3948 1383
rect 5317 1377 5356 1383
rect 804 1357 1068 1363
rect 1093 1357 1180 1363
rect 1316 1357 1339 1363
rect 1540 1357 1676 1363
rect 1861 1357 2092 1363
rect 3716 1357 3739 1363
rect 3892 1357 4012 1363
rect 468 1337 636 1343
rect 644 1337 843 1343
rect 868 1337 1372 1343
rect 3956 1337 5324 1343
rect 532 1317 1132 1323
rect 1172 1317 1484 1323
rect 2340 1317 2556 1323
rect 4132 1317 4316 1323
rect 4612 1317 4748 1323
rect 132 1297 732 1303
rect 3220 1297 3292 1303
rect 4164 1297 4236 1303
rect 3172 1277 4972 1283
rect 3956 1257 4204 1263
rect 4820 1237 4827 1243
rect 1396 1217 1403 1223
rect 1117 1204 1123 1215
rect 1604 1157 1804 1163
rect 4020 1157 4764 1163
rect 4805 1157 5164 1163
rect 1284 1137 1756 1143
rect 1892 1137 1916 1143
rect 3572 1137 4700 1143
rect 132 1117 1467 1123
rect 1732 1117 1788 1123
rect 1812 1117 2524 1123
rect 3284 1117 3788 1123
rect 3812 1117 3835 1123
rect 3845 1117 4091 1123
rect 4101 1117 4124 1123
rect 4228 1117 4364 1123
rect 4660 1117 4812 1123
rect 4980 1117 5036 1123
rect 548 1097 1308 1103
rect 1396 1097 2299 1103
rect 2420 1097 2620 1103
rect 2644 1097 2812 1103
rect 3460 1097 3707 1103
rect 3717 1097 4332 1103
rect 4756 1097 5068 1103
rect 5252 1097 5292 1103
rect 292 1077 315 1083
rect 372 1077 620 1083
rect 1284 1077 2956 1083
rect 2996 1077 3804 1083
rect 3956 1077 4044 1083
rect 180 1057 300 1063
rect 644 1057 716 1063
rect 852 1057 2284 1063
rect 2309 1057 2444 1063
rect 2452 1057 2636 1063
rect 2692 1057 3068 1063
rect 3492 1057 3740 1063
rect 4324 1057 4876 1063
rect 4964 1057 5164 1063
rect 788 1037 940 1043
rect 1380 1037 1403 1043
rect 1477 1037 1804 1043
rect 2500 1037 2683 1043
rect 2756 1037 2844 1043
rect 708 1017 1820 1023
rect 1253 997 1372 1003
rect 4708 997 4731 1003
rect 1012 977 1516 983
rect 1605 977 1948 983
rect 2116 977 2828 983
rect 4773 977 5036 983
rect 5285 977 5388 983
rect 820 957 1388 963
rect 1413 957 1468 963
rect 1588 957 1595 963
rect 2212 957 2332 963
rect 404 937 460 943
rect 997 937 1548 943
rect 2196 937 2428 943
rect 3236 937 3388 943
rect 4548 937 4732 943
rect 132 917 1052 923
rect 1093 917 1260 923
rect 2756 917 2860 923
rect 3748 917 3916 923
rect 4228 917 4300 923
rect 5140 917 5404 923
rect 1668 897 2668 903
rect 468 877 940 883
rect 2877 877 3052 883
rect 2693 857 2716 863
rect 2877 863 2883 877
rect 3060 877 3099 883
rect 4228 877 4284 883
rect 4292 877 4444 883
rect 4484 877 4748 883
rect 4804 877 5260 883
rect 2868 857 2883 863
rect 2788 837 3212 843
rect 3220 837 3516 843
rect 4165 837 4172 843
rect 1076 817 1083 823
rect 1172 817 1260 823
rect 965 797 972 803
rect 2164 797 3068 803
rect 3076 797 3388 803
rect 3813 797 4748 803
rect 980 777 1244 783
rect 1252 777 1484 783
rect 2756 757 2892 763
rect 4036 757 4188 763
rect 4212 757 5068 763
rect 836 737 987 743
rect 4069 737 4172 743
rect 4197 737 4284 743
rect 4997 737 5036 743
rect 804 717 1356 723
rect 1541 717 1708 723
rect 2949 717 3803 723
rect 3828 717 4539 723
rect 4804 717 4940 723
rect 1156 697 1276 703
rect 2100 697 2524 703
rect 3860 697 4284 703
rect 4292 697 5036 703
rect 5124 697 5388 703
rect 1124 677 1596 683
rect 1604 677 2124 683
rect 3109 677 3260 683
rect 3668 677 3804 683
rect 3956 677 3963 683
rect 3988 677 4092 683
rect 4165 677 4204 683
rect 4244 677 4268 683
rect 4293 677 4540 683
rect 4772 677 5052 683
rect 1172 657 1564 663
rect 1572 657 2140 663
rect 2452 657 2684 663
rect 3732 657 4060 663
rect 4116 657 4348 663
rect 4868 657 5100 663
rect 3940 637 4140 643
rect 1012 617 1500 623
rect 2804 617 3148 623
rect 3156 617 3516 623
rect 4069 617 4076 623
rect 1540 597 1740 603
rect 3172 597 3196 603
rect 4229 597 4236 603
rect 1637 577 1676 583
rect 2532 577 2636 583
rect 3988 577 4252 583
rect 4549 577 4668 583
rect 4837 577 4876 583
rect 1125 557 2380 563
rect 2388 557 2444 563
rect 2564 557 2636 563
rect 3316 557 3452 563
rect 3956 557 4188 563
rect 4244 557 4588 563
rect 4741 557 5372 563
rect 1124 537 1932 543
rect 1956 537 2636 543
rect 3652 537 4220 543
rect 4372 537 5292 543
rect 3412 517 3500 523
rect 3908 517 4236 523
rect 4292 517 4332 523
rect 1605 497 1628 503
rect 2020 497 2700 503
rect 4212 497 4572 503
rect 2212 477 2508 483
rect 3588 377 4731 383
rect 292 337 572 343
rect 1445 337 1484 343
rect 2724 337 2844 343
rect 3972 337 3996 343
rect 1380 317 1484 323
rect 2132 317 2508 323
rect 3796 317 3932 323
rect 3949 317 4396 323
rect 692 297 716 303
rect 1221 297 2268 303
rect 3732 297 3868 303
rect 3949 303 3955 317
rect 5028 317 5276 323
rect 3892 297 3955 303
rect 3972 297 4508 303
rect 4836 297 5292 303
rect 308 277 812 283
rect 1092 277 1324 283
rect 1940 277 2124 283
rect 3140 277 3291 283
rect 3316 277 4364 283
rect 516 257 1052 263
rect 1412 257 1532 263
rect 1573 257 1644 263
rect 3268 257 3324 263
rect 3332 257 3772 263
rect 3780 257 3884 263
rect 3940 257 4060 263
rect 4244 257 4348 263
rect 4612 257 4924 263
rect 965 237 972 243
rect 1444 237 1724 243
rect 3252 237 3564 243
rect 3700 237 3803 243
rect 3844 237 4268 243
rect 3301 217 3628 223
rect 4164 217 4316 223
rect 3845 197 4876 203
rect 20 177 76 183
rect 613 177 716 183
rect 964 177 1308 183
rect 2580 177 2940 183
rect 3524 177 3788 183
rect 4484 177 4540 183
rect 868 157 1211 163
rect 5245 164 5251 175
rect 1677 157 1804 163
rect 228 137 684 143
rect 1124 137 1147 143
rect 1172 137 1244 143
rect 1268 137 1372 143
rect 1677 143 1683 157
rect 3108 157 3756 163
rect 1572 137 1683 143
rect 1748 137 1948 143
rect 2340 137 2860 143
rect 2884 137 2972 143
rect 3252 137 3324 143
rect 4389 137 5452 143
rect 389 117 428 123
rect 644 117 700 123
rect 804 117 1164 123
rect 1188 117 1740 123
rect 1757 117 2348 123
rect 1220 97 1260 103
rect 1348 97 1371 103
rect 1757 103 1763 117
rect 4308 117 4364 123
rect 1604 97 1763 103
rect 2116 97 2252 103
rect 4532 97 4556 103
rect 3860 77 4588 83
<< m6contact >>
rect 5307 3855 5317 3865
rect 5243 3784 5253 3785
rect 5243 3776 5244 3784
rect 5244 3776 5252 3784
rect 5252 3776 5253 3784
rect 5243 3775 5253 3776
rect 5339 3764 5349 3765
rect 5339 3756 5340 3764
rect 5340 3756 5348 3764
rect 5348 3756 5349 3764
rect 5339 3755 5349 3756
rect 4347 3735 4357 3745
rect 4267 3695 4277 3705
rect 4395 3695 4405 3705
rect 4667 3484 4677 3485
rect 4667 3476 4668 3484
rect 4668 3476 4676 3484
rect 4676 3476 4677 3484
rect 4667 3475 4677 3476
rect 891 3435 901 3445
rect 1979 3424 1989 3425
rect 1979 3416 1980 3424
rect 1980 3416 1988 3424
rect 1988 3416 1989 3424
rect 1979 3415 1989 3416
rect 2171 3395 2181 3405
rect 5115 3395 5125 3405
rect 3579 3355 3589 3365
rect 3675 3355 3685 3365
rect 1851 3335 1861 3345
rect 4923 3335 4933 3345
rect 4123 3315 4133 3325
rect 1723 3295 1733 3305
rect 4891 3295 4901 3305
rect 4091 3275 4101 3285
rect 1083 3215 1093 3225
rect 3803 3204 3813 3205
rect 3803 3196 3804 3204
rect 3804 3196 3812 3204
rect 3812 3196 3813 3204
rect 635 3184 645 3185
rect 635 3176 636 3184
rect 636 3176 644 3184
rect 644 3176 645 3184
rect 3803 3195 3813 3196
rect 635 3175 645 3176
rect 1339 3135 1349 3145
rect 4731 3115 4741 3125
rect 1307 3095 1317 3105
rect 3643 3095 3653 3105
rect 1339 3055 1349 3065
rect 3643 3055 3653 3065
rect 4987 3035 4997 3045
rect 3675 3015 3685 3025
rect 4091 3015 4101 3025
rect 2939 2995 2949 3005
rect 3259 2995 3269 3005
rect 4731 3004 4741 3005
rect 4731 2996 4732 3004
rect 4732 2996 4740 3004
rect 4740 2996 4741 3004
rect 4731 2995 4741 2996
rect 1307 2975 1317 2985
rect 3323 2975 3333 2985
rect 3611 2955 3621 2965
rect 3227 2935 3237 2945
rect 5115 2915 5125 2925
rect 3323 2895 3333 2905
rect 3643 2875 3653 2885
rect 3771 2855 3781 2865
rect 795 2795 805 2805
rect 1211 2775 1221 2785
rect 1019 2755 1029 2765
rect 1819 2755 1829 2765
rect 923 2735 933 2745
rect 1915 2744 1925 2745
rect 1915 2736 1916 2744
rect 1916 2736 1924 2744
rect 1924 2736 1925 2744
rect 1915 2735 1925 2736
rect 2043 2744 2053 2745
rect 2043 2736 2044 2744
rect 2044 2736 2052 2744
rect 2052 2736 2053 2744
rect 2043 2735 2053 2736
rect 3195 2724 3205 2725
rect 3195 2716 3196 2724
rect 3196 2716 3204 2724
rect 3204 2716 3205 2724
rect 3195 2715 3205 2716
rect 1307 2695 1317 2705
rect 3675 2695 3685 2705
rect 955 2675 965 2685
rect 795 2635 805 2645
rect 923 2635 933 2645
rect 1211 2635 1221 2645
rect 3739 2635 3749 2645
rect 1243 2575 1253 2585
rect 1627 2575 1637 2585
rect 3195 2575 3205 2585
rect 3739 2575 3749 2585
rect 4443 2575 4453 2585
rect 4571 2555 4581 2565
rect 1339 2535 1349 2545
rect 1467 2535 1477 2545
rect 3867 2535 3877 2545
rect 3899 2515 3909 2525
rect 4763 2495 4773 2505
rect 5083 2495 5093 2505
rect 5083 2395 5093 2405
rect 4347 2355 4357 2365
rect 1371 2335 1381 2345
rect 3643 2335 3653 2345
rect 4283 2344 4293 2345
rect 4283 2336 4284 2344
rect 4284 2336 4292 2344
rect 4292 2336 4293 2344
rect 4283 2335 4293 2336
rect 1851 2315 1861 2325
rect 5339 2315 5349 2325
rect 4347 2295 4357 2305
rect 1851 2275 1861 2285
rect 3803 2275 3813 2285
rect 4443 2255 4453 2265
rect 2299 2155 2309 2165
rect 4091 2155 4101 2165
rect 4955 2164 4965 2165
rect 4955 2156 4956 2164
rect 4956 2156 4964 2164
rect 4964 2156 4965 2164
rect 4955 2155 4965 2156
rect 1691 2144 1701 2145
rect 315 2115 325 2125
rect 1691 2136 1692 2144
rect 1692 2136 1700 2144
rect 1700 2136 1701 2144
rect 1691 2135 1701 2136
rect 2043 2135 2053 2145
rect 1851 2115 1861 2125
rect 3707 2104 3717 2105
rect 3707 2096 3708 2104
rect 3708 2096 3716 2104
rect 3716 2096 3717 2104
rect 3707 2095 3717 2096
rect 4955 2095 4965 2105
rect 1211 2075 1221 2085
rect 1659 2075 1669 2085
rect 3771 2055 3781 2065
rect 859 1995 869 2005
rect 4923 1995 4933 2005
rect 827 1975 837 1985
rect 4123 1975 4133 1985
rect 5275 1955 5285 1965
rect 4987 1915 4997 1925
rect 827 1895 837 1905
rect 859 1855 869 1865
rect 4955 1855 4965 1865
rect 1403 1815 1413 1825
rect 1083 1795 1093 1805
rect 1563 1804 1573 1805
rect 1563 1796 1564 1804
rect 1564 1796 1572 1804
rect 1572 1796 1573 1804
rect 1563 1795 1573 1796
rect 4123 1775 4133 1785
rect 1659 1755 1669 1765
rect 5275 1755 5285 1765
rect 4571 1735 4581 1745
rect 635 1715 645 1725
rect 5275 1715 5285 1725
rect 4955 1695 4965 1705
rect 1371 1675 1381 1685
rect 1467 1664 1477 1665
rect 1467 1656 1468 1664
rect 1468 1656 1476 1664
rect 1476 1656 1477 1664
rect 1467 1655 1477 1656
rect 1691 1655 1701 1665
rect 3771 1655 3781 1665
rect 4987 1655 4997 1665
rect 3739 1595 3749 1605
rect 4795 1595 4805 1605
rect 4891 1595 4901 1605
rect 1595 1584 1605 1585
rect 1595 1576 1596 1584
rect 1596 1576 1604 1584
rect 1604 1576 1605 1584
rect 1595 1575 1605 1576
rect 3675 1575 3685 1585
rect 1371 1555 1381 1565
rect 1659 1555 1669 1565
rect 891 1475 901 1485
rect 3963 1475 3973 1485
rect 1147 1455 1157 1465
rect 1659 1455 1669 1465
rect 1531 1415 1541 1425
rect 1435 1375 1445 1385
rect 3771 1375 3781 1385
rect 5307 1375 5317 1385
rect 1083 1355 1093 1365
rect 1339 1355 1349 1365
rect 1851 1355 1861 1365
rect 3739 1355 3749 1365
rect 843 1335 853 1345
rect 1339 1304 1349 1305
rect 1339 1296 1340 1304
rect 1340 1296 1348 1304
rect 1348 1296 1349 1304
rect 1339 1295 1349 1296
rect 4827 1235 4837 1245
rect 1115 1215 1125 1225
rect 1403 1215 1413 1225
rect 4795 1155 4805 1165
rect 2299 1144 2309 1145
rect 2299 1136 2300 1144
rect 2300 1136 2308 1144
rect 2308 1136 2309 1144
rect 2299 1135 2309 1136
rect 1467 1115 1477 1125
rect 3835 1115 3845 1125
rect 4091 1115 4101 1125
rect 2299 1095 2309 1105
rect 3707 1095 3717 1105
rect 315 1075 325 1085
rect 2299 1055 2309 1065
rect 1403 1035 1413 1045
rect 1467 1035 1477 1045
rect 2683 1035 2693 1045
rect 1243 995 1253 1005
rect 4731 995 4741 1005
rect 1595 975 1605 985
rect 4763 975 4773 985
rect 5275 975 5285 985
rect 1403 955 1413 965
rect 1595 955 1605 965
rect 987 935 997 945
rect 1083 915 1093 925
rect 2683 855 2693 865
rect 3099 875 3109 885
rect 4155 835 4165 845
rect 1083 815 1093 825
rect 955 795 965 805
rect 3803 795 3813 805
rect 4187 784 4197 785
rect 4187 776 4188 784
rect 4188 776 4196 784
rect 4196 776 4197 784
rect 4187 775 4197 776
rect 3835 764 3845 765
rect 3835 756 3836 764
rect 3836 756 3844 764
rect 3844 756 3845 764
rect 3835 755 3845 756
rect 987 735 997 745
rect 3963 744 3973 745
rect 3963 736 3964 744
rect 3964 736 3972 744
rect 3972 736 3973 744
rect 3963 735 3973 736
rect 4059 735 4069 745
rect 4187 735 4197 745
rect 4379 744 4389 745
rect 4379 736 4380 744
rect 4380 736 4388 744
rect 4388 736 4389 744
rect 4379 735 4389 736
rect 4987 735 4997 745
rect 1531 715 1541 725
rect 2939 715 2949 725
rect 3803 715 3813 725
rect 4539 715 4549 725
rect 379 704 389 705
rect 379 696 380 704
rect 380 696 388 704
rect 388 696 389 704
rect 379 695 389 696
rect 3099 675 3109 685
rect 3963 675 3973 685
rect 4155 675 4165 685
rect 4283 675 4293 685
rect 603 624 613 625
rect 603 616 604 624
rect 604 616 612 624
rect 612 616 613 624
rect 603 615 613 616
rect 4059 615 4069 625
rect 4219 595 4229 605
rect 1627 575 1637 585
rect 4539 575 4549 585
rect 4827 575 4837 585
rect 1115 564 1125 565
rect 1115 556 1116 564
rect 1116 556 1124 564
rect 1124 556 1125 564
rect 1115 555 1125 556
rect 4731 555 4741 565
rect 1595 495 1605 505
rect 4731 375 4741 385
rect 1435 335 1445 345
rect 1211 295 1221 305
rect 3291 275 3301 285
rect 1563 255 1573 265
rect 955 235 965 245
rect 3803 235 3813 245
rect 3291 215 3301 225
rect 3835 195 3845 205
rect 603 175 613 185
rect 5243 175 5253 185
rect 1211 155 1221 165
rect 1147 135 1157 145
rect 4379 135 4389 145
rect 379 115 389 125
rect 1371 95 1381 105
<< metal6 >>
rect 4123 3735 4347 3745
rect 315 1085 325 2115
rect 635 1725 645 3175
rect 795 2645 805 2795
rect 827 1905 837 1975
rect 859 1865 869 1995
rect 891 1485 901 3435
rect 1979 3385 1989 3415
rect 2171 3385 2181 3395
rect 1979 3375 2181 3385
rect 1723 3335 1851 3345
rect 1723 3305 1733 3335
rect 923 2645 933 2735
rect 1019 2705 1029 2755
rect 955 2695 1029 2705
rect 955 2685 965 2695
rect 1083 1805 1093 3215
rect 1339 3105 1349 3135
rect 1317 3095 1349 3105
rect 1211 2645 1221 2775
rect 1307 2705 1317 2975
rect 1083 1345 1093 1355
rect 853 1335 1093 1345
rect 379 125 389 695
rect 603 185 613 615
rect 955 245 965 795
rect 987 745 997 935
rect 1083 825 1093 915
rect 1115 565 1125 1215
rect 1147 145 1157 1455
rect 1211 305 1221 2075
rect 1243 1005 1253 2575
rect 1339 2545 1349 3055
rect 1819 2705 1829 2755
rect 1915 2705 1925 2735
rect 1819 2695 1925 2705
rect 1371 1685 1381 2335
rect 1339 1305 1349 1355
rect 1211 165 1221 295
rect 1371 105 1381 1555
rect 1403 1225 1413 1815
rect 1467 1665 1477 2535
rect 1403 965 1413 1035
rect 1435 345 1445 1375
rect 1467 1045 1477 1115
rect 1531 725 1541 1415
rect 1563 265 1573 1795
rect 1595 985 1605 1575
rect 1595 505 1605 955
rect 1627 585 1637 2575
rect 1851 2285 1861 2315
rect 2043 2145 2053 2735
rect 1659 1765 1669 2075
rect 1691 1665 1701 2135
rect 1659 1465 1669 1555
rect 1851 1365 1861 2115
rect 2299 1145 2309 2155
rect 2299 1065 2309 1095
rect 2683 865 2693 1035
rect 2939 725 2949 2995
rect 3259 2945 3269 2995
rect 3237 2935 3269 2945
rect 3323 2905 3333 2975
rect 3579 2945 3589 3355
rect 3643 3065 3653 3095
rect 3675 3025 3685 3355
rect 4123 3325 4133 3735
rect 4277 3695 4395 3705
rect 3611 2945 3621 2955
rect 3579 2935 3621 2945
rect 3195 2585 3205 2715
rect 3643 2345 3653 2875
rect 3675 1585 3685 2695
rect 3739 2585 3749 2635
rect 3707 1105 3717 2095
rect 3771 2065 3781 2855
rect 3803 2285 3813 3195
rect 4091 3025 4101 3275
rect 4667 3145 4677 3475
rect 4667 3135 4741 3145
rect 4731 3125 4741 3135
rect 3877 2535 3909 2545
rect 3899 2525 3909 2535
rect 3739 1365 3749 1595
rect 3771 1385 3781 1655
rect 3099 685 3109 875
rect 3803 725 3813 795
rect 3835 765 3845 1115
rect 3963 745 3973 1475
rect 4091 1125 4101 2155
rect 4123 1785 4133 1975
rect 4059 705 4069 735
rect 3963 695 4069 705
rect 3963 685 3973 695
rect 4155 685 4165 835
rect 4187 745 4197 775
rect 4283 685 4293 2335
rect 4347 2305 4357 2355
rect 4443 2265 4453 2575
rect 4571 1745 4581 2555
rect 4731 1005 4741 2995
rect 4059 585 4069 615
rect 4219 585 4229 595
rect 4059 575 4229 585
rect 3291 225 3301 275
rect 3803 255 3845 265
rect 3803 245 3813 255
rect 3835 205 3845 255
rect 4379 145 4389 735
rect 4539 585 4549 715
rect 4731 565 4741 995
rect 4763 985 4773 2495
rect 4891 1605 4901 3295
rect 4923 2005 4933 3335
rect 4955 2105 4965 2155
rect 4987 1925 4997 3035
rect 5115 2925 5125 3395
rect 5083 2405 5093 2495
rect 4955 1705 4965 1855
rect 4795 1165 4805 1595
rect 4827 585 4837 1235
rect 4987 745 4997 1655
rect 4731 385 4741 555
rect 5243 185 5253 3775
rect 5275 1765 5285 1955
rect 5275 985 5285 1715
rect 5307 1385 5317 3855
rect 5339 2325 5349 3755
use FILL  FILL_20_4
timestamp 1598358358
transform 1 0 5560 0 1 3810
box -16 -6 32 210
use AND2X1  AND2X1_192
timestamp 1598358358
transform 1 0 5448 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_551
timestamp 1598358358
transform 1 0 5384 0 1 3810
box -16 -6 80 210
use FILL  FILL_20_3
timestamp 1598358358
transform 1 0 5544 0 1 3810
box -16 -6 32 210
use FILL  FILL_20_2
timestamp 1598358358
transform 1 0 5528 0 1 3810
box -16 -6 32 210
use FILL  FILL_20_1
timestamp 1598358358
transform 1 0 5512 0 1 3810
box -16 -6 32 210
use AND2X1  AND2X1_545
timestamp 1598358358
transform 1 0 5320 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_659
timestamp 1598358358
transform -1 0 5320 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_622
timestamp 1598358358
transform 1 0 5192 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_658
timestamp 1598358358
transform 1 0 5128 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_158
timestamp 1598358358
transform 1 0 4936 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_156
timestamp 1598358358
transform -1 0 5128 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_210
timestamp 1598358358
transform 1 0 5000 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_163
timestamp 1598358358
transform 1 0 4872 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_162
timestamp 1598358358
transform 1 0 4808 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_161
timestamp 1598358358
transform 1 0 4744 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_467
timestamp 1598358358
transform -1 0 4744 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_603
timestamp 1598358358
transform -1 0 4488 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_470
timestamp 1598358358
transform 1 0 4616 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_466
timestamp 1598358358
transform 1 0 4552 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_453
timestamp 1598358358
transform -1 0 4552 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_604
timestamp 1598358358
transform 1 0 4296 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_605
timestamp 1598358358
transform -1 0 4424 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_446
timestamp 1598358358
transform 1 0 4232 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_418
timestamp 1598358358
transform 1 0 4104 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_313
timestamp 1598358358
transform 1 0 3976 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_704
timestamp 1598358358
transform 1 0 4168 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_317
timestamp 1598358358
transform 1 0 4040 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_314
timestamp 1598358358
transform 1 0 3912 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_683
timestamp 1598358358
transform -1 0 3912 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_686
timestamp 1598358358
transform -1 0 3848 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_684
timestamp 1598358358
transform -1 0 3784 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_765
timestamp 1598358358
transform -1 0 3720 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_452
timestamp 1598358358
transform 1 0 3592 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_450
timestamp 1598358358
transform 1 0 3528 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_426
timestamp 1598358358
transform 1 0 3464 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_427
timestamp 1598358358
transform 1 0 3400 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_451
timestamp 1598358358
transform 1 0 3336 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_430
timestamp 1598358358
transform 1 0 3272 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_428
timestamp 1598358358
transform 1 0 3208 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_582
timestamp 1598358358
transform 1 0 3080 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_635
timestamp 1598358358
transform -1 0 3208 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_70
timestamp 1598358358
transform 1 0 3016 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_581
timestamp 1598358358
transform 1 0 2952 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_425
timestamp 1598358358
transform 1 0 2888 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_51
timestamp 1598358358
transform 1 0 2824 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_157
timestamp 1598358358
transform -1 0 2824 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_25
timestamp 1598358358
transform 1 0 2696 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_429
timestamp 1598358358
transform 1 0 2632 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_11
timestamp 1598358358
transform 1 0 2568 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_50
timestamp 1598358358
transform 1 0 2504 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_30
timestamp 1598358358
transform 1 0 2440 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_17
timestamp 1598358358
transform 1 0 2376 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_2
timestamp 1598358358
transform 1 0 2312 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_21
timestamp 1598358358
transform -1 0 2312 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_1
timestamp 1598358358
transform 1 0 2184 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_17
timestamp 1598358358
transform -1 0 2184 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_50
timestamp 1598358358
transform -1 0 2120 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_25
timestamp 1598358358
transform 1 0 1992 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_11
timestamp 1598358358
transform -1 0 1992 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_2
timestamp 1598358358
transform -1 0 1928 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_12
timestamp 1598358358
transform -1 0 1864 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_429
timestamp 1598358358
transform -1 0 1800 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_3
timestamp 1598358358
transform -1 0 1736 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_425
timestamp 1598358358
transform -1 0 1672 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_157
timestamp 1598358358
transform -1 0 1608 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_686
timestamp 1598358358
transform -1 0 1416 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_685
timestamp 1598358358
transform -1 0 1352 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_581
timestamp 1598358358
transform -1 0 1544 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_582
timestamp 1598358358
transform 1 0 1416 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_687
timestamp 1598358358
transform -1 0 1288 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_451
timestamp 1598358358
transform -1 0 1160 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_430
timestamp 1598358358
transform -1 0 1224 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_452
timestamp 1598358358
transform -1 0 1096 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_450
timestamp 1598358358
transform 1 0 968 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_694
timestamp 1598358358
transform 1 0 904 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_426
timestamp 1598358358
transform 1 0 840 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_780
timestamp 1598358358
transform -1 0 840 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_454
timestamp 1598358358
transform -1 0 776 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_449
timestamp 1598358358
transform -1 0 712 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_453
timestamp 1598358358
transform -1 0 648 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_466
timestamp 1598358358
transform -1 0 584 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_480
timestamp 1598358358
transform 1 0 456 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_478
timestamp 1598358358
transform 1 0 392 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_467
timestamp 1598358358
transform -1 0 392 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_470
timestamp 1598358358
transform -1 0 328 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_477
timestamp 1598358358
transform 1 0 200 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_162
timestamp 1598358358
transform 1 0 72 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_161
timestamp 1598358358
transform 1 0 8 0 1 3810
box -16 -6 80 210
use AND2X1  AND2X1_163
timestamp 1598358358
transform 1 0 136 0 1 3810
box -16 -6 80 210
use OR2X1  OR2X1_747
timestamp 1598358358
transform 1 0 5448 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_782
timestamp 1598358358
transform 1 0 5512 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_797
timestamp 1598358358
transform 1 0 5512 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_213
timestamp 1598358358
transform 1 0 5448 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_781
timestamp 1598358358
transform 1 0 5384 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_149
timestamp 1598358358
transform 1 0 5384 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_745
timestamp 1598358358
transform 1 0 5320 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_746
timestamp 1598358358
transform 1 0 5256 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_145
timestamp 1598358358
transform 1 0 5192 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_146
timestamp 1598358358
transform 1 0 5128 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_676
timestamp 1598358358
transform 1 0 5320 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_148
timestamp 1598358358
transform 1 0 5256 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_154
timestamp 1598358358
transform -1 0 5256 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_155
timestamp 1598358358
transform -1 0 5192 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_744
timestamp 1598358358
transform -1 0 5128 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_743
timestamp 1598358358
transform 1 0 4936 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_511
timestamp 1598358358
transform 1 0 4936 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_783
timestamp 1598358358
transform 1 0 5064 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_780
timestamp 1598358358
transform 1 0 5000 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_779
timestamp 1598358358
transform 1 0 5000 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_696
timestamp 1598358358
transform -1 0 4936 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_591
timestamp 1598358358
transform -1 0 4872 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_697
timestamp 1598358358
transform 1 0 4744 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_422
timestamp 1598358358
transform -1 0 4744 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_160
timestamp 1598358358
transform -1 0 4936 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_708
timestamp 1598358358
transform -1 0 4872 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_718
timestamp 1598358358
transform 1 0 4744 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_593
timestamp 1598358358
transform -1 0 4744 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_424
timestamp 1598358358
transform -1 0 4488 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_448
timestamp 1598358358
transform 1 0 4616 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_732
timestamp 1598358358
transform 1 0 4616 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_725
timestamp 1598358358
transform 1 0 4552 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_713
timestamp 1598358358
transform -1 0 4616 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_712
timestamp 1598358358
transform 1 0 4488 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_645
timestamp 1598358358
transform -1 0 4552 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_454
timestamp 1598358358
transform 1 0 4424 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_423
timestamp 1598358358
transform 1 0 4296 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_421
timestamp 1598358358
transform 1 0 4232 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_449
timestamp 1598358358
transform 1 0 4360 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_592
timestamp 1598358358
transform 1 0 4360 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_714
timestamp 1598358358
transform 1 0 4296 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_832
timestamp 1598358358
transform 1 0 4232 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_682
timestamp 1598358358
transform 1 0 4168 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_589
timestamp 1598358358
transform 1 0 4168 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_681
timestamp 1598358358
transform 1 0 4040 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_433
timestamp 1598358358
transform 1 0 4040 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_432
timestamp 1598358358
transform 1 0 3976 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_685
timestamp 1598358358
transform 1 0 4104 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_435
timestamp 1598358358
transform 1 0 4104 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_687
timestamp 1598358358
transform -1 0 4040 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_695
timestamp 1598358358
transform 1 0 3848 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_694
timestamp 1598358358
transform 1 0 3784 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_693
timestamp 1598358358
transform 1 0 3848 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_707
timestamp 1598358358
transform 1 0 3912 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_706
timestamp 1598358358
transform 1 0 3912 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_648
timestamp 1598358358
transform -1 0 3848 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_766
timestamp 1598358358
transform -1 0 3784 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_692
timestamp 1598358358
transform 1 0 3720 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_584
timestamp 1598358358
transform -1 0 3656 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_583
timestamp 1598358358
transform -1 0 3592 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_770
timestamp 1598358358
transform 1 0 3656 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_596
timestamp 1598358358
transform 1 0 3656 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_828
timestamp 1598358358
transform 1 0 3592 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_771
timestamp 1598358358
transform 1 0 3528 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_386
timestamp 1598358358
transform -1 0 3464 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_764
timestamp 1598358358
transform 1 0 3400 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_328
timestamp 1598358358
transform -1 0 3400 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_763
timestamp 1598358358
transform 1 0 3336 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_636
timestamp 1598358358
transform -1 0 3528 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_769
timestamp 1598358358
transform 1 0 3464 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_18
timestamp 1598358358
transform -1 0 3272 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_762
timestamp 1598358358
transform 1 0 3208 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_12
timestamp 1598358358
transform 1 0 3144 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_3
timestamp 1598358358
transform 1 0 3080 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_639
timestamp 1598358358
transform -1 0 3336 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_651
timestamp 1598358358
transform 1 0 3272 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_638
timestamp 1598358358
transform 1 0 3144 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_379
timestamp 1598358358
transform -1 0 3144 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_40
timestamp 1598358358
transform 1 0 3016 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_64
timestamp 1598358358
transform 1 0 3016 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_22
timestamp 1598358358
transform 1 0 2952 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_26
timestamp 1598358358
transform 1 0 2952 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_47
timestamp 1598358358
transform 1 0 2888 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_380
timestamp 1598358358
transform -1 0 2952 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_44
timestamp 1598358358
transform -1 0 2888 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_588
timestamp 1598358358
transform 1 0 2824 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_31
timestamp 1598358358
transform 1 0 2760 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_587
timestamp 1598358358
transform 1 0 2696 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_409
timestamp 1598358358
transform 1 0 2696 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_36
timestamp 1598358358
transform 1 0 2632 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_460
timestamp 1598358358
transform -1 0 2824 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_463
timestamp 1598358358
transform 1 0 2632 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_1
timestamp 1598358358
transform 1 0 2568 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_408
timestamp 1598358358
transform 1 0 2568 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_21
timestamp 1598358358
transform 1 0 2504 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_30
timestamp 1598358358
transform -1 0 2568 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_51
timestamp 1598358358
transform -1 0 2504 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_408
timestamp 1598358358
transform 1 0 2440 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_587
timestamp 1598358358
transform -1 0 2440 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_588
timestamp 1598358358
transform 1 0 2376 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_44
timestamp 1598358358
transform -1 0 2376 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_36
timestamp 1598358358
transform -1 0 2376 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_31
timestamp 1598358358
transform 1 0 2248 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_47
timestamp 1598358358
transform 1 0 2184 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_64
timestamp 1598358358
transform -1 0 2312 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_762
timestamp 1598358358
transform 1 0 2184 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_22
timestamp 1598358358
transform -1 0 2184 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_26
timestamp 1598358358
transform -1 0 2184 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_70
timestamp 1598358358
transform 1 0 2056 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_95
timestamp 1598358358
transform 1 0 2056 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_40
timestamp 1598358358
transform -1 0 2056 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_59
timestamp 1598358358
transform -1 0 2056 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_639
timestamp 1598358358
transform 1 0 1928 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_636
timestamp 1598358358
transform 1 0 1864 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_328
timestamp 1598358358
transform -1 0 1992 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_386
timestamp 1598358358
transform 1 0 1864 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_583
timestamp 1598358358
transform -1 0 1864 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_7
timestamp 1598358358
transform 1 0 1800 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_584
timestamp 1598358358
transform 1 0 1736 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_18
timestamp 1598358358
transform -1 0 1800 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_635
timestamp 1598358358
transform 1 0 1608 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_195
timestamp 1598358358
transform -1 0 1672 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_614
timestamp 1598358358
transform -1 0 1608 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_199
timestamp 1598358358
transform 1 0 1544 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_428
timestamp 1598358358
transform 1 0 1672 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_43
timestamp 1598358358
transform 1 0 1672 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_196
timestamp 1598358358
transform 1 0 1416 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_683
timestamp 1598358358
transform -1 0 1544 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_754
timestamp 1598358358
transform 1 0 1480 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_684
timestamp 1598358358
transform -1 0 1480 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_682
timestamp 1598358358
transform -1 0 1416 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_48
timestamp 1598358358
transform 1 0 1352 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_681
timestamp 1598358358
transform -1 0 1352 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_615
timestamp 1598358358
transform -1 0 1352 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_446
timestamp 1598358358
transform -1 0 1224 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_307
timestamp 1598358358
transform 1 0 1096 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_418
timestamp 1598358358
transform -1 0 1288 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_511
timestamp 1598358358
transform -1 0 1288 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_427
timestamp 1598358358
transform -1 0 1160 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_304
timestamp 1598358358
transform -1 0 1224 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_707
timestamp 1598358358
transform -1 0 1032 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_777
timestamp 1598358358
transform -1 0 968 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_784
timestamp 1598358358
transform -1 0 904 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_695
timestamp 1598358358
transform -1 0 1096 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_306
timestamp 1598358358
transform 1 0 1032 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_677
timestamp 1598358358
transform 1 0 968 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_743
timestamp 1598358358
transform -1 0 968 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_744
timestamp 1598358358
transform -1 0 904 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_448
timestamp 1598358358
transform -1 0 840 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_783
timestamp 1598358358
transform -1 0 776 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_779
timestamp 1598358358
transform -1 0 776 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_796
timestamp 1598358358
transform -1 0 712 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_712
timestamp 1598358358
transform 1 0 648 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_424
timestamp 1598358358
transform -1 0 840 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_803
timestamp 1598358358
transform 1 0 584 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_155
timestamp 1598358358
transform -1 0 584 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_708
timestamp 1598358358
transform 1 0 584 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_154
timestamp 1598358358
transform -1 0 520 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_156
timestamp 1598358358
transform -1 0 456 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_696
timestamp 1598358358
transform -1 0 584 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_701
timestamp 1598358358
transform 1 0 456 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_526
timestamp 1598358358
transform -1 0 456 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_160
timestamp 1598358358
transform -1 0 392 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_210
timestamp 1598358358
transform -1 0 264 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_148
timestamp 1598358358
transform -1 0 264 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_146
timestamp 1598358358
transform -1 0 392 0 1 3410
box -16 -6 80 210
use AND2X1  AND2X1_158
timestamp 1598358358
transform -1 0 328 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_145
timestamp 1598358358
transform -1 0 328 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_781
timestamp 1598358358
transform 1 0 8 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_797
timestamp 1598358358
transform 1 0 136 0 -1 3810
box -16 -6 80 210
use OR2X1  OR2X1_149
timestamp 1598358358
transform -1 0 200 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_782
timestamp 1598358358
transform 1 0 72 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_747
timestamp 1598358358
transform 1 0 8 0 -1 3810
box -16 -6 80 210
use AND2X1  AND2X1_745
timestamp 1598358358
transform -1 0 136 0 1 3410
box -16 -6 80 210
use OR2X1  OR2X1_679
timestamp 1598358358
transform 1 0 5384 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_730
timestamp 1598358358
transform 1 0 5512 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_209
timestamp 1598358358
transform -1 0 5512 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_144
timestamp 1598358358
transform 1 0 5128 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_728
timestamp 1598358358
transform -1 0 5384 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_147
timestamp 1598358358
transform 1 0 5256 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_678
timestamp 1598358358
transform 1 0 5192 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_526
timestamp 1598358358
transform 1 0 5064 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_485
timestamp 1598358358
transform 1 0 5000 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_705
timestamp 1598358358
transform -1 0 5000 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_420
timestamp 1598358358
transform -1 0 4872 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_419
timestamp 1598358358
transform -1 0 4744 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_590
timestamp 1598358358
transform -1 0 4936 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_447
timestamp 1598358358
transform -1 0 4808 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_600
timestamp 1598358358
transform -1 0 4680 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_601
timestamp 1598358358
transform 1 0 4424 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_602
timestamp 1598358358
transform -1 0 4616 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_724
timestamp 1598358358
transform 1 0 4488 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_167
timestamp 1598358358
transform -1 0 4424 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_703
timestamp 1598358358
transform -1 0 4360 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_598
timestamp 1598358358
transform -1 0 4296 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_329
timestamp 1598358358
transform 1 0 4168 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_312
timestamp 1598358358
transform 1 0 4104 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_760
timestamp 1598358358
transform -1 0 4104 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_800
timestamp 1598358358
transform 1 0 3976 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_599
timestamp 1598358358
transform -1 0 3912 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_729
timestamp 1598358358
transform -1 0 3976 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_644
timestamp 1598358358
transform 1 0 3784 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_597
timestamp 1598358358
transform 1 0 3720 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_536
timestamp 1598358358
transform -1 0 3720 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_537
timestamp 1598358358
transform -1 0 3656 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_407
timestamp 1598358358
transform -1 0 3592 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_586
timestamp 1598358358
transform -1 0 3528 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_387
timestamp 1598358358
transform 1 0 3336 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_389
timestamp 1598358358
transform 1 0 3400 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_385
timestamp 1598358358
transform 1 0 3272 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_95
timestamp 1598358358
transform 1 0 3208 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_585
timestamp 1598358358
transform 1 0 3080 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_637
timestamp 1598358358
transform -1 0 3208 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_59
timestamp 1598358358
transform 1 0 3016 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_53
timestamp 1598358358
transform 1 0 2952 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_752
timestamp 1598358358
transform -1 0 2952 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_376
timestamp 1598358358
transform -1 0 2824 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_377
timestamp 1598358358
transform 1 0 2696 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_375
timestamp 1598358358
transform -1 0 2888 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_459
timestamp 1598358358
transform -1 0 2696 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_378
timestamp 1598358358
transform -1 0 2632 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_375
timestamp 1598358358
transform -1 0 2568 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_752
timestamp 1598358358
transform -1 0 2504 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_638
timestamp 1598358358
transform -1 0 2440 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_651
timestamp 1598358358
transform 1 0 2312 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_53
timestamp 1598358358
transform -1 0 2312 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_56
timestamp 1598358358
transform -1 0 2248 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_197
timestamp 1598358358
transform -1 0 2184 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_228
timestamp 1598358358
transform -1 0 2056 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_52
timestamp 1598358358
transform -1 0 2120 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_207
timestamp 1598358358
transform 1 0 1864 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_200
timestamp 1598358358
transform 1 0 1800 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_193
timestamp 1598358358
transform -1 0 1800 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_41
timestamp 1598358358
transform -1 0 1992 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_790
timestamp 1598358358
transform 1 0 1608 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_753
timestamp 1598358358
transform -1 0 1736 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_693
timestamp 1598358358
transform -1 0 1608 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_706
timestamp 1598358358
transform -1 0 1416 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_678
timestamp 1598358358
transform 1 0 1288 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_45
timestamp 1598358358
transform -1 0 1544 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_692
timestamp 1598358358
transform -1 0 1480 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_513
timestamp 1598358358
transform 1 0 1224 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_512
timestamp 1598358358
transform 1 0 1160 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_308
timestamp 1598358358
transform -1 0 1160 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_834
timestamp 1598358358
transform 1 0 1032 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_305
timestamp 1598358358
transform -1 0 1032 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_421
timestamp 1598358358
transform -1 0 968 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_422
timestamp 1598358358
transform -1 0 904 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_713
timestamp 1598358358
transform -1 0 776 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_725
timestamp 1598358358
transform -1 0 712 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_697
timestamp 1598358358
transform -1 0 840 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_710
timestamp 1598358358
transform -1 0 520 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_705
timestamp 1598358358
transform 1 0 392 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_700
timestamp 1598358358
transform -1 0 648 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_144
timestamp 1598358358
transform -1 0 584 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_147
timestamp 1598358358
transform -1 0 392 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_546
timestamp 1598358358
transform -1 0 264 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_525
timestamp 1598358358
transform -1 0 328 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_209
timestamp 1598358358
transform -1 0 200 0 -1 3410
box -16 -6 80 210
use OR2X1  OR2X1_213
timestamp 1598358358
transform -1 0 136 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_746
timestamp 1598358358
transform -1 0 72 0 -1 3410
box -16 -6 80 210
use AND2X1  AND2X1_739
timestamp 1598358358
transform 1 0 5512 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_740
timestamp 1598358358
transform 1 0 5448 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_738
timestamp 1598358358
transform 1 0 5384 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_677
timestamp 1598358358
transform 1 0 5256 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_680
timestamp 1598358358
transform 1 0 5128 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_803
timestamp 1598358358
transform 1 0 5320 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_546
timestamp 1598358358
transform 1 0 5192 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_525
timestamp 1598358358
transform 1 0 5000 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_834
timestamp 1598358358
transform -1 0 5128 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_513
timestamp 1598358358
transform -1 0 5000 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_331
timestamp 1598358358
transform 1 0 4808 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_533
timestamp 1598358358
transform -1 0 4808 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_330
timestamp 1598358358
transform 1 0 4872 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_788
timestamp 1598358358
transform 1 0 4680 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_534
timestamp 1598358358
transform 1 0 4616 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_166
timestamp 1598358358
transform 1 0 4424 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_390
timestamp 1598358358
transform -1 0 4616 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_535
timestamp 1598358358
transform -1 0 4552 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_436
timestamp 1598358358
transform 1 0 4360 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_169
timestamp 1598358358
transform -1 0 4360 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_355
timestamp 1598358358
transform 1 0 4232 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_336
timestamp 1598358358
transform 1 0 4168 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_356
timestamp 1598358358
transform 1 0 4104 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_809
timestamp 1598358358
transform 1 0 4040 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_801
timestamp 1598358358
transform 1 0 3976 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_761
timestamp 1598358358
transform 1 0 3912 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_512
timestamp 1598358358
transform -1 0 3912 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_855
timestamp 1598358358
transform 1 0 3784 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_829
timestamp 1598358358
transform 1 0 3720 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_306
timestamp 1598358358
transform 1 0 3656 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_539
timestamp 1598358358
transform 1 0 3592 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_538
timestamp 1598358358
transform 1 0 3528 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_13
timestamp 1598358358
transform -1 0 3528 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_311
timestamp 1598358358
transform 1 0 3400 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_41
timestamp 1598358358
transform -1 0 3400 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_43
timestamp 1598358358
transform -1 0 3336 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_195
timestamp 1598358358
transform -1 0 3272 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_199
timestamp 1598358358
transform -1 0 3208 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_207
timestamp 1598358358
transform -1 0 3144 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_200
timestamp 1598358358
transform 1 0 3016 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_193
timestamp 1598358358
transform 1 0 2952 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_691
timestamp 1598358358
transform 1 0 2888 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_689
timestamp 1598358358
transform 1 0 2824 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_690
timestamp 1598358358
transform 1 0 2760 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_378
timestamp 1598358358
transform -1 0 2760 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_688
timestamp 1598358358
transform -1 0 2696 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_459
timestamp 1598358358
transform -1 0 2632 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_376
timestamp 1598358358
transform -1 0 2568 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_409
timestamp 1598358358
transform 1 0 2440 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_637
timestamp 1598358358
transform 1 0 2312 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_764
timestamp 1598358358
transform 1 0 2376 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_763
timestamp 1598358358
transform 1 0 2248 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_829
timestamp 1598358358
transform 1 0 2184 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_828
timestamp 1598358358
transform -1 0 2184 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_407
timestamp 1598358358
transform 1 0 2056 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_676
timestamp 1598358358
transform -1 0 2056 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_596
timestamp 1598358358
transform 1 0 1864 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_597
timestamp 1598358358
transform 1 0 1928 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_13
timestamp 1598358358
transform -1 0 1864 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_16
timestamp 1598358358
transform -1 0 1800 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_194
timestamp 1598358358
transform 1 0 1672 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_39
timestamp 1598358358
transform 1 0 1608 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_699
timestamp 1598358358
transform -1 0 1608 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_514
timestamp 1598358358
transform -1 0 1480 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_515
timestamp 1598358358
transform -1 0 1416 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_702
timestamp 1598358358
transform -1 0 1352 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_136
timestamp 1598358358
transform -1 0 1544 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_715
timestamp 1598358358
transform -1 0 1160 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_516
timestamp 1598358358
transform -1 0 1288 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_679
timestamp 1598358358
transform -1 0 1224 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_447
timestamp 1598358358
transform -1 0 968 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_704
timestamp 1598358358
transform -1 0 904 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_423
timestamp 1598358358
transform 1 0 1032 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_419
timestamp 1598358358
transform 1 0 968 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_714
timestamp 1598358358
transform -1 0 840 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_724
timestamp 1598358358
transform -1 0 776 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_313
timestamp 1598358358
transform 1 0 648 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_732
timestamp 1598358358
transform -1 0 648 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_709
timestamp 1598358358
transform -1 0 584 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_469
timestamp 1598358358
transform -1 0 456 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_698
timestamp 1598358358
transform 1 0 456 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_711
timestamp 1598358358
transform -1 0 392 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_727
timestamp 1598358358
transform -1 0 328 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_484
timestamp 1598358358
transform -1 0 264 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_738
timestamp 1598358358
transform -1 0 72 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_726
timestamp 1598358358
transform -1 0 200 0 1 3010
box -16 -6 80 210
use OR2X1  OR2X1_731
timestamp 1598358358
transform -1 0 136 0 1 3010
box -16 -6 80 210
use AND2X1  AND2X1_742
timestamp 1598358358
transform 1 0 5512 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_731
timestamp 1598358358
transform 1 0 5448 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_726
timestamp 1598358358
transform 1 0 5384 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_152
timestamp 1598358358
transform 1 0 5320 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_812
timestamp 1598358358
transform 1 0 5256 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_727
timestamp 1598358358
transform 1 0 5192 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_151
timestamp 1598358358
transform 1 0 5128 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_142
timestamp 1598358358
transform 1 0 5000 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_484
timestamp 1598358358
transform -1 0 5000 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_796
timestamp 1598358358
transform 1 0 5064 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_594
timestamp 1598358358
transform -1 0 4808 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_486
timestamp 1598358358
transform 1 0 4872 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_468
timestamp 1598358358
transform -1 0 4872 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_532
timestamp 1598358358
transform -1 0 4744 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_652
timestamp 1598358358
transform -1 0 4680 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_653
timestamp 1598358358
transform -1 0 4616 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_799
timestamp 1598358358
transform -1 0 4552 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_810
timestamp 1598358358
transform 1 0 4424 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_388
timestamp 1598358358
transform -1 0 4424 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_802
timestamp 1598358358
transform 1 0 4296 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_567
timestamp 1598358358
transform -1 0 4296 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_798
timestamp 1598358358
transform 1 0 4168 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_319
timestamp 1598358358
transform 1 0 4104 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_354
timestamp 1598358358
transform 1 0 4040 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_715
timestamp 1598358358
transform -1 0 4040 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_854
timestamp 1598358358
transform -1 0 3976 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_856
timestamp 1598358358
transform -1 0 3912 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_308
timestamp 1598358358
transform -1 0 3848 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_305
timestamp 1598358358
transform -1 0 3720 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_135
timestamp 1598358358
transform -1 0 3592 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_774
timestamp 1598358358
transform 1 0 3720 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_307
timestamp 1598358358
transform 1 0 3592 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_431
timestamp 1598358358
transform -1 0 3464 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_304
timestamp 1598358358
transform 1 0 3336 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_702
timestamp 1598358358
transform 1 0 3464 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_45
timestamp 1598358358
transform 1 0 3208 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_172
timestamp 1598358358
transform 1 0 3144 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_434
timestamp 1598358358
transform -1 0 3336 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_196
timestamp 1598358358
transform -1 0 3144 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_48
timestamp 1598358358
transform -1 0 3080 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_7
timestamp 1598358358
transform -1 0 3016 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_16
timestamp 1598358358
transform -1 0 2952 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_56
timestamp 1598358358
transform -1 0 2888 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_39
timestamp 1598358358
transform -1 0 2760 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_194
timestamp 1598358358
transform -1 0 2824 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_377
timestamp 1598358358
transform 1 0 2632 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_463
timestamp 1598358358
transform 1 0 2568 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_460
timestamp 1598358358
transform 1 0 2504 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_380
timestamp 1598358358
transform 1 0 2440 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_769
timestamp 1598358358
transform -1 0 2376 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_598
timestamp 1598358358
transform -1 0 2312 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_585
timestamp 1598358358
transform 1 0 2376 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_586
timestamp 1598358358
transform -1 0 2248 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_855
timestamp 1598358358
transform -1 0 2184 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_379
timestamp 1598358358
transform 1 0 2056 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_644
timestamp 1598358358
transform 1 0 1992 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_599
timestamp 1598358358
transform 1 0 1928 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_761
timestamp 1598358358
transform -1 0 1928 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_751
timestamp 1598358358
transform 1 0 1800 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_748
timestamp 1598358358
transform -1 0 1800 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_789
timestamp 1598358358
transform -1 0 1736 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_793
timestamp 1598358358
transform 1 0 1608 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_138
timestamp 1598358358
transform 1 0 1544 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_801
timestamp 1598358358
transform 1 0 1480 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_800
timestamp 1598358358
transform 1 0 1416 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_185
timestamp 1598358358
transform 1 0 1288 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_760
timestamp 1598358358
transform 1 0 1352 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_729
timestamp 1598358358
transform -1 0 1288 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_730
timestamp 1598358358
transform -1 0 1224 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_728
timestamp 1598358358
transform 1 0 1096 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_317
timestamp 1598358358
transform -1 0 904 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_680
timestamp 1598358358
transform 1 0 1032 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_420
timestamp 1598358358
transform -1 0 1032 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_314
timestamp 1598358358
transform -1 0 968 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_355
timestamp 1598358358
transform 1 0 712 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_329
timestamp 1598358358
transform -1 0 840 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_331
timestamp 1598358358
transform 1 0 648 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_330
timestamp 1598358358
transform 1 0 584 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_532
timestamp 1598358358
transform 1 0 520 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_324
timestamp 1598358358
transform 1 0 392 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_320
timestamp 1598358358
transform -1 0 520 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_486
timestamp 1598358358
transform 1 0 200 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_321
timestamp 1598358358
transform 1 0 328 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_142
timestamp 1598358358
transform 1 0 264 0 -1 3010
box -16 -6 80 210
use OR2X1  OR2X1_151
timestamp 1598358358
transform -1 0 136 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_485
timestamp 1598358358
transform 1 0 136 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_152
timestamp 1598358358
transform 1 0 8 0 -1 3010
box -16 -6 80 210
use AND2X1  AND2X1_221
timestamp 1598358358
transform 1 0 5512 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_478
timestamp 1598358358
transform 1 0 5448 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_220
timestamp 1598358358
transform 1 0 5384 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_442
timestamp 1598358358
transform 1 0 5128 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_469
timestamp 1598358358
transform 1 0 5320 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_808
timestamp 1598358358
transform 1 0 5256 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_444
timestamp 1598358358
transform 1 0 5192 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_516
timestamp 1598358358
transform -1 0 5128 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_794
timestamp 1598358358
transform 1 0 5000 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_787
timestamp 1598358358
transform 1 0 4936 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_417
timestamp 1598358358
transform 1 0 4744 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_477
timestamp 1598358358
transform -1 0 4936 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_515
timestamp 1598358358
transform 1 0 4808 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_568
timestamp 1598358358
transform 1 0 4680 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_176
timestamp 1598358358
transform -1 0 4680 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_170
timestamp 1598358358
transform -1 0 4616 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_566
timestamp 1598358358
transform 1 0 4488 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_211
timestamp 1598358358
transform -1 0 4488 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_864
timestamp 1598358358
transform -1 0 4424 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_212
timestamp 1598358358
transform 1 0 4296 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_365
timestamp 1598358358
transform 1 0 4232 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_661
timestamp 1598358358
transform -1 0 4232 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_337
timestamp 1598358358
transform 1 0 4104 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_352
timestamp 1598358358
transform -1 0 4104 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_353
timestamp 1598358358
transform 1 0 3976 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_321
timestamp 1598358358
transform 1 0 3784 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_863
timestamp 1598358358
transform 1 0 3912 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_324
timestamp 1598358358
transform 1 0 3848 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_320
timestamp 1598358358
transform 1 0 3720 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_299
timestamp 1598358358
transform -1 0 3656 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_777
timestamp 1598358358
transform -1 0 3720 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_302
timestamp 1598358358
transform 1 0 3528 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_298
timestamp 1598358358
transform -1 0 3528 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_654
timestamp 1598358358
transform 1 0 3400 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_174
timestamp 1598358358
transform 1 0 3336 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_230
timestamp 1598358358
transform -1 0 3336 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_229
timestamp 1598358358
transform 1 0 3144 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_231
timestamp 1598358358
transform 1 0 3208 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_228
timestamp 1598358358
transform 1 0 3080 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_52
timestamp 1598358358
transform -1 0 3080 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_214
timestamp 1598358358
transform -1 0 3016 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_197
timestamp 1598358358
transform -1 0 2952 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_57
timestamp 1598358358
transform 1 0 2760 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_19
timestamp 1598358358
transform -1 0 2760 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_198
timestamp 1598358358
transform 1 0 2824 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_827
timestamp 1598358358
transform 1 0 2632 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_839
timestamp 1598358358
transform 1 0 2568 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_836
timestamp 1598358358
transform 1 0 2504 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_823
timestamp 1598358358
transform -1 0 2504 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_835
timestamp 1598358358
transform 1 0 2376 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_691
timestamp 1598358358
transform -1 0 2312 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_822
timestamp 1598358358
transform 1 0 2312 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_821
timestamp 1598358358
transform 1 0 2184 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_856
timestamp 1598358358
transform 1 0 2120 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_198
timestamp 1598358358
transform -1 0 2120 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_23
timestamp 1598358358
transform 1 0 1992 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_750
timestamp 1598358358
transform -1 0 1992 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_387
timestamp 1598358358
transform -1 0 1928 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_536
timestamp 1598358358
transform 1 0 1800 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_135
timestamp 1598358358
transform -1 0 1800 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_538
timestamp 1598358358
transform 1 0 1672 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_110
timestamp 1598358358
transform -1 0 1672 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_173
timestamp 1598358358
transform 1 0 1544 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_186
timestamp 1598358358
transform 1 0 1352 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_623
timestamp 1598358358
transform -1 0 1352 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_111
timestamp 1598358358
transform 1 0 1480 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_311
timestamp 1598358358
transform 1 0 1416 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_319
timestamp 1598358358
transform -1 0 1288 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_854
timestamp 1598358358
transform 1 0 1160 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_354
timestamp 1598358358
transform -1 0 1160 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_356
timestamp 1598358358
transform -1 0 968 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_703
timestamp 1598358358
transform -1 0 904 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_167
timestamp 1598358358
transform -1 0 1096 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_534
timestamp 1598358358
transform -1 0 1032 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_326
timestamp 1598358358
transform 1 0 712 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_325
timestamp 1598358358
transform 1 0 648 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_533
timestamp 1598358358
transform 1 0 776 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_302
timestamp 1598358358
transform 1 0 392 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_322
timestamp 1598358358
transform 1 0 584 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_323
timestamp 1598358358
transform 1 0 520 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_299
timestamp 1598358358
transform -1 0 520 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_620
timestamp 1598358358
transform 1 0 200 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_298
timestamp 1598358358
transform -1 0 392 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_527
timestamp 1598358358
transform -1 0 328 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_739
timestamp 1598358358
transform 1 0 8 0 1 2610
box -16 -6 80 210
use OR2X1  OR2X1_740
timestamp 1598358358
transform 1 0 72 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_613
timestamp 1598358358
transform 1 0 136 0 1 2610
box -16 -6 80 210
use AND2X1  AND2X1_223
timestamp 1598358358
transform 1 0 5512 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_480
timestamp 1598358358
transform 1 0 5448 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_741
timestamp 1598358358
transform 1 0 5384 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_441
timestamp 1598358358
transform 1 0 5320 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_811
timestamp 1598358358
transform 1 0 5256 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_737
timestamp 1598358358
transform 1 0 5192 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_443
timestamp 1598358358
transform 1 0 5128 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_437
timestamp 1598358358
transform 1 0 4936 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_804
timestamp 1598358358
transform 1 0 5064 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_784
timestamp 1598358358
transform 1 0 5000 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_440
timestamp 1598358358
transform -1 0 4936 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_733
timestamp 1598358358
transform 1 0 4808 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_722
timestamp 1598358358
transform 1 0 4744 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_168
timestamp 1598358358
transform -1 0 4744 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_165
timestamp 1598358358
transform 1 0 4616 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_91
timestamp 1598358358
transform -1 0 4488 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_723
timestamp 1598358358
transform -1 0 4616 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_180
timestamp 1598358358
transform -1 0 4552 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_369
timestamp 1598358358
transform 1 0 4232 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_370
timestamp 1598358358
transform 1 0 4360 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_182
timestamp 1598358358
transform -1 0 4360 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_309
timestamp 1598358358
transform -1 0 4232 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_310
timestamp 1598358358
transform 1 0 4040 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_335
timestamp 1598358358
transform -1 0 4168 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_357
timestamp 1598358358
transform -1 0 4040 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_519
timestamp 1598358358
transform 1 0 3912 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_326
timestamp 1598358358
transform -1 0 3912 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_514
timestamp 1598358358
transform 1 0 3784 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_136
timestamp 1598358358
transform -1 0 3720 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_364
timestamp 1598358358
transform 1 0 3720 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_303
timestamp 1598358358
transform -1 0 3656 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_716
timestamp 1598358358
transform 1 0 3528 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_173
timestamp 1598358358
transform -1 0 3528 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_175
timestamp 1598358358
transform -1 0 3464 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_341
timestamp 1598358358
transform 1 0 3336 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_171
timestamp 1598358358
transform 1 0 3080 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_641
timestamp 1598358358
transform 1 0 3272 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_650
timestamp 1598358358
transform 1 0 3208 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_857
timestamp 1598358358
transform -1 0 3208 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_24
timestamp 1598358358
transform -1 0 3016 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_853
timestamp 1598358358
transform 1 0 3016 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_208
timestamp 1598358358
transform 1 0 2888 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_20
timestamp 1598358358
transform 1 0 2696 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_838
timestamp 1598358358
transform -1 0 2696 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_35
timestamp 1598358358
transform 1 0 2824 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_33
timestamp 1598358358
transform 1 0 2760 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_852
timestamp 1598358358
transform -1 0 2632 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_824
timestamp 1598358358
transform 1 0 2504 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_690
timestamp 1598358358
transform 1 0 2440 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_688
timestamp 1598358358
transform -1 0 2440 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_853
timestamp 1598358358
transform 1 0 2248 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_857
timestamp 1598358358
transform -1 0 2248 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_689
timestamp 1598358358
transform -1 0 2376 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_863
timestamp 1598358358
transform -1 0 2184 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_208
timestamp 1598358358
transform -1 0 2056 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_57
timestamp 1598358358
transform 1 0 2056 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_214
timestamp 1598358358
transform -1 0 1992 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_389
timestamp 1598358358
transform -1 0 1928 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_537
timestamp 1598358358
transform -1 0 1800 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_385
timestamp 1598358358
transform -1 0 1864 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_539
timestamp 1598358358
transform -1 0 1736 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_332
timestamp 1598358358
transform 1 0 1608 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_175
timestamp 1598358358
transform 1 0 1544 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_112
timestamp 1598358358
transform -1 0 1544 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_809
timestamp 1598358358
transform -1 0 1480 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_802
timestamp 1598358358
transform 1 0 1288 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_417
timestamp 1598358358
transform -1 0 1416 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_799
timestamp 1598358358
transform 1 0 1224 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_798
timestamp 1598358358
transform 1 0 1160 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_468
timestamp 1598358358
transform 1 0 1096 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_567
timestamp 1598358358
transform -1 0 1096 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_535
timestamp 1598358358
transform 1 0 968 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_169
timestamp 1598358358
transform -1 0 904 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_166
timestamp 1598358358
transform -1 0 968 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_170
timestamp 1598358358
transform -1 0 840 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_568
timestamp 1598358358
transform -1 0 776 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_566
timestamp 1598358358
transform 1 0 648 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_211
timestamp 1598358358
transform -1 0 648 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_336
timestamp 1598358358
transform -1 0 584 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_303
timestamp 1598358358
transform 1 0 456 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_353
timestamp 1598358358
transform -1 0 456 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_212
timestamp 1598358358
transform -1 0 392 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_312
timestamp 1598358358
transform 1 0 264 0 -1 2610
box -16 -6 80 210
use AND2X1  AND2X1_528
timestamp 1598358358
transform -1 0 264 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_220
timestamp 1598358358
transform -1 0 72 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_547
timestamp 1598358358
transform -1 0 200 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_550
timestamp 1598358358
transform -1 0 136 0 -1 2610
box -16 -6 80 210
use OR2X1  OR2X1_524
timestamp 1598358358
transform -1 0 5576 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_479
timestamp 1598358358
transform 1 0 5448 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_550
timestamp 1598358358
transform 1 0 5384 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_438
timestamp 1598358358
transform -1 0 5384 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_177
timestamp 1598358358
transform -1 0 5320 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_544
timestamp 1598358358
transform 1 0 5192 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_439
timestamp 1598358358
transform 1 0 5128 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_373
timestamp 1598358358
transform 1 0 5064 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_775
timestamp 1598358358
transform 1 0 5000 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_405
timestamp 1598358358
transform 1 0 4936 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_109
timestamp 1598358358
transform -1 0 4936 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_164
timestamp 1598358358
transform 1 0 4808 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_542
timestamp 1598358358
transform -1 0 4808 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_552
timestamp 1598358358
transform -1 0 4744 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_322
timestamp 1598358358
transform 1 0 4552 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_368
timestamp 1598358358
transform -1 0 4488 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_374
timestamp 1598358358
transform 1 0 4616 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_457
timestamp 1598358358
transform 1 0 4488 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_323
timestamp 1598358358
transform 1 0 4296 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_543
timestamp 1598358358
transform 1 0 4360 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_325
timestamp 1598358358
transform -1 0 4296 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_111
timestamp 1598358358
transform -1 0 4168 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_518
timestamp 1598358358
transform -1 0 4040 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_841
timestamp 1598358358
transform 1 0 4168 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_112
timestamp 1598358358
transform -1 0 4104 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_520
timestamp 1598358358
transform 1 0 3912 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_332
timestamp 1598358358
transform 1 0 3848 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_655
timestamp 1598358358
transform 1 0 3784 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_289
timestamp 1598358358
transform -1 0 3592 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_138
timestamp 1598358358
transform 1 0 3720 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_643
timestamp 1598358358
transform 1 0 3656 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_358
timestamp 1598358358
transform 1 0 3592 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_350
timestamp 1598358358
transform -1 0 3528 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_351
timestamp 1598358358
transform 1 0 3400 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_333
timestamp 1598358358
transform -1 0 3400 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_46
timestamp 1598358358
transform -1 0 3272 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_411
timestamp 1598358358
transform -1 0 3144 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_338
timestamp 1598358358
transform 1 0 3272 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_410
timestamp 1598358358
transform -1 0 3208 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_413
timestamp 1598358358
transform -1 0 3080 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_837
timestamp 1598358358
transform -1 0 2952 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_461
timestamp 1598358358
transform 1 0 2952 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_472
timestamp 1598358358
transform 1 0 2824 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_826
timestamp 1598358358
transform 1 0 2760 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_233
timestamp 1598358358
transform 1 0 2696 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_411
timestamp 1598358358
transform 1 0 2632 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_410
timestamp 1598358358
transform 1 0 2568 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_334
timestamp 1598358358
transform -1 0 2568 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_27
timestamp 1598358358
transform -1 0 2504 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_34
timestamp 1598358358
transform -1 0 2440 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_35
timestamp 1598358358
transform -1 0 2376 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_33
timestamp 1598358358
transform 1 0 2248 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_24
timestamp 1598358358
transform 1 0 2184 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_338
timestamp 1598358358
transform -1 0 2184 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_333
timestamp 1598358358
transform 1 0 2056 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_289
timestamp 1598358358
transform -1 0 2056 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_351
timestamp 1598358358
transform 1 0 1928 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_339
timestamp 1598358358
transform 1 0 1800 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_171
timestamp 1598358358
transform 1 0 1864 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_431
timestamp 1598358358
transform -1 0 1800 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_174
timestamp 1598358358
transform -1 0 1736 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_434
timestamp 1598358358
transform -1 0 1672 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_436
timestamp 1598358358
transform 1 0 1544 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_435
timestamp 1598358358
transform 1 0 1416 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_652
timestamp 1598358358
transform 1 0 1352 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_594
timestamp 1598358358
transform 1 0 1480 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_589
timestamp 1598358358
transform -1 0 1352 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_592
timestamp 1598358358
transform -1 0 1288 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_593
timestamp 1598358358
transform -1 0 1224 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_165
timestamp 1598358358
transform -1 0 1160 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_168
timestamp 1598358358
transform -1 0 1096 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_388
timestamp 1598358358
transform 1 0 968 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_440
timestamp 1598358358
transform 1 0 840 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_176
timestamp 1598358358
transform -1 0 968 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_437
timestamp 1598358358
transform 1 0 776 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_177
timestamp 1598358358
transform -1 0 776 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_373
timestamp 1598358358
transform -1 0 712 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_180
timestamp 1598358358
transform -1 0 648 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_337
timestamp 1598358358
transform 1 0 520 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_352
timestamp 1598358358
transform -1 0 520 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_357
timestamp 1598358358
transform 1 0 392 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_182
timestamp 1598358358
transform 1 0 328 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_444
timestamp 1598358358
transform 1 0 264 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_442
timestamp 1598358358
transform 1 0 200 0 1 2210
box -16 -6 80 210
use OR2X1  OR2X1_221
timestamp 1598358358
transform 1 0 8 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_441
timestamp 1598358358
transform 1 0 136 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_187
timestamp 1598358358
transform -1 0 136 0 1 2210
box -16 -6 80 210
use AND2X1  AND2X1_547
timestamp 1598358358
transform 1 0 5512 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_475
timestamp 1598358358
transform 1 0 5448 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_564
timestamp 1598358358
transform 1 0 5384 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_406
timestamp 1598358358
transform -1 0 5320 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_496
timestamp 1598358358
transform 1 0 5192 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_734
timestamp 1598358358
transform -1 0 5384 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_795
timestamp 1598358358
transform 1 0 5128 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_778
timestamp 1598358358
transform 1 0 5064 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_785
timestamp 1598358358
transform 1 0 5000 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_776
timestamp 1598358358
transform -1 0 5000 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_527
timestamp 1598358358
transform 1 0 4872 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_471
timestamp 1598358358
transform 1 0 4808 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_464
timestamp 1598358358
transform 1 0 4744 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_458
timestamp 1598358358
transform 1 0 4680 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_372
timestamp 1598358358
transform 1 0 4552 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_371
timestamp 1598358358
transform 1 0 4488 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_315
timestamp 1598358358
transform -1 0 4488 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_717
timestamp 1598358358
transform -1 0 4680 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_271
timestamp 1598358358
transform -1 0 4360 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_270
timestamp 1598358358
transform -1 0 4424 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_318
timestamp 1598358358
transform -1 0 4296 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_268
timestamp 1598358358
transform -1 0 4104 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_110
timestamp 1598358358
transform 1 0 3976 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_269
timestamp 1598358358
transform 1 0 4168 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_476
timestamp 1598358358
transform 1 0 4104 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_222
timestamp 1598358358
transform -1 0 3976 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_642
timestamp 1598358358
transform 1 0 3848 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_649
timestamp 1598358358
transform -1 0 3848 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_273
timestamp 1598358358
transform 1 0 3656 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_300
timestamp 1598358358
transform 1 0 3592 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_831
timestamp 1598358358
transform 1 0 3720 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_301
timestamp 1598358358
transform 1 0 3528 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_75
timestamp 1598358358
transform -1 0 3528 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_339
timestamp 1598358358
transform 1 0 3400 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_219
timestamp 1598358358
transform 1 0 3336 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_290
timestamp 1598358358
transform 1 0 3080 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_640
timestamp 1598358358
transform -1 0 3336 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_334
timestamp 1598358358
transform 1 0 3208 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_634
timestamp 1598358358
transform 1 0 3144 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_27
timestamp 1598358358
transform -1 0 3080 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_293
timestamp 1598358358
transform -1 0 3016 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_462
timestamp 1598358358
transform -1 0 2952 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_462
timestamp 1598358358
transform 1 0 2760 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_461
timestamp 1598358358
transform 1 0 2696 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_34
timestamp 1598358358
transform 1 0 2824 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_413
timestamp 1598358358
transform 1 0 2632 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_472
timestamp 1598358358
transform 1 0 2568 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_634
timestamp 1598358358
transform 1 0 2504 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_291
timestamp 1598358358
transform 1 0 2440 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_654
timestamp 1598358358
transform -1 0 2312 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_661
timestamp 1598358358
transform -1 0 2248 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_32
timestamp 1598358358
transform -1 0 2440 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_290
timestamp 1598358358
transform 1 0 2312 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_648
timestamp 1598358358
transform 1 0 1992 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_20
timestamp 1598358358
transform 1 0 2120 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_749
timestamp 1598358358
transform 1 0 2056 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_61
timestamp 1598358358
transform -1 0 1864 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_58
timestamp 1598358358
transform 1 0 1928 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_60
timestamp 1598358358
transform -1 0 1928 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_172
timestamp 1598358358
transform -1 0 1800 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_405
timestamp 1598358358
transform -1 0 1736 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_358
timestamp 1598358358
transform -1 0 1672 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_390
timestamp 1598358358
transform -1 0 1608 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_653
timestamp 1598358358
transform -1 0 1544 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_775
timestamp 1598358358
transform -1 0 1416 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_109
timestamp 1598358358
transform -1 0 1480 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_432
timestamp 1598358358
transform -1 0 1352 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_832
timestamp 1598358358
transform -1 0 1224 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_433
timestamp 1598358358
transform 1 0 1224 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_164
timestamp 1598358358
transform -1 0 1160 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_602
timestamp 1598358358
transform -1 0 1032 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_645
timestamp 1598358358
transform 1 0 840 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_601
timestamp 1598358358
transform -1 0 1096 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_600
timestamp 1598358358
transform 1 0 904 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_788
timestamp 1598358358
transform -1 0 840 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_374
timestamp 1598358358
transform 1 0 648 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_91
timestamp 1598358358
transform -1 0 776 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_439
timestamp 1598358358
transform 1 0 584 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_544
timestamp 1598358358
transform -1 0 520 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_364
timestamp 1598358358
transform -1 0 456 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_438
timestamp 1598358358
transform 1 0 520 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_365
timestamp 1598358358
transform -1 0 392 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_443
timestamp 1598358358
transform -1 0 328 0 -1 2210
box -16 -6 80 210
use AND2X1  AND2X1_524
timestamp 1598358358
transform -1 0 264 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_223
timestamp 1598358358
transform -1 0 72 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_545
timestamp 1598358358
transform -1 0 200 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_551
timestamp 1598358358
transform -1 0 136 0 -1 2210
box -16 -6 80 210
use OR2X1  OR2X1_189
timestamp 1598358358
transform 1 0 5384 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_498
timestamp 1598358358
transform -1 0 5512 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_578
timestamp 1598358358
transform 1 0 5512 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_569
timestamp 1598358358
transform 1 0 5448 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_577
timestamp 1598358358
transform 1 0 5512 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_736
timestamp 1598358358
transform 1 0 5384 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_531
timestamp 1598358358
transform 1 0 5192 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_530
timestamp 1598358358
transform 1 0 5128 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_565
timestamp 1598358358
transform 1 0 5320 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_549
timestamp 1598358358
transform 1 0 5256 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_675
timestamp 1598358358
transform -1 0 5192 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_188
timestamp 1598358358
transform 1 0 5320 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_186
timestamp 1598358358
transform -1 0 5320 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_548
timestamp 1598358358
transform 1 0 5192 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_674
timestamp 1598358358
transform 1 0 5000 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_492
timestamp 1598358358
transform 1 0 5000 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_499
timestamp 1598358358
transform 1 0 5064 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_833
timestamp 1598358358
transform 1 0 4936 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_830
timestamp 1598358358
transform 1 0 5064 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_493
timestamp 1598358358
transform 1 0 4936 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_495
timestamp 1598358358
transform 1 0 4680 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_491
timestamp 1598358358
transform 1 0 4872 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_183
timestamp 1598358358
transform -1 0 4744 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_840
timestamp 1598358358
transform -1 0 4936 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_851
timestamp 1598358358
transform -1 0 4872 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_241
timestamp 1598358358
transform 1 0 4744 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_465
timestamp 1598358358
transform 1 0 4808 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_190
timestamp 1598358358
transform 1 0 4744 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_238
timestamp 1598358358
transform 1 0 4616 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_237
timestamp 1598358358
transform 1 0 4552 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_280
timestamp 1598358358
transform -1 0 4552 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_224
timestamp 1598358358
transform 1 0 4616 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_178
timestamp 1598358358
transform -1 0 4616 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_179
timestamp 1598358358
transform -1 0 4488 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_445
timestamp 1598358358
transform -1 0 4488 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_540
timestamp 1598358358
transform -1 0 4552 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_522
timestamp 1598358358
transform -1 0 4360 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_108
timestamp 1598358358
transform 1 0 4296 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_455
timestamp 1598358358
transform 1 0 4360 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_523
timestamp 1598358358
transform 1 0 4232 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_181
timestamp 1598358358
transform -1 0 4424 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_114
timestamp 1598358358
transform -1 0 4296 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_521
timestamp 1598358358
transform 1 0 4104 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_115
timestamp 1598358358
transform -1 0 4232 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_276
timestamp 1598358358
transform -1 0 4104 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_662
timestamp 1598358358
transform -1 0 4040 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_116
timestamp 1598358358
transform -1 0 4232 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_473
timestamp 1598358358
transform -1 0 4168 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_327
timestamp 1598358358
transform 1 0 4040 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_660
timestamp 1598358358
transform 1 0 3976 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_517
timestamp 1598358358
transform 1 0 3848 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_275
timestamp 1598358358
transform 1 0 3784 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_272
timestamp 1598358358
transform 1 0 3784 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_559
timestamp 1598358358
transform 1 0 3912 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_218
timestamp 1598358358
transform 1 0 3912 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_216
timestamp 1598358358
transform 1 0 3848 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_595
timestamp 1598358358
transform -1 0 3720 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_153
timestamp 1598358358
transform 1 0 3528 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_767
timestamp 1598358358
transform 1 0 3656 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_79
timestamp 1598358358
transform -1 0 3592 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_264
timestamp 1598358358
transform 1 0 3720 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_274
timestamp 1598358358
transform 1 0 3592 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_773
timestamp 1598358358
transform 1 0 3720 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_78
timestamp 1598358358
transform -1 0 3656 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_74
timestamp 1598358358
transform 1 0 3400 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_65
timestamp 1598358358
transform -1 0 3400 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_76
timestamp 1598358358
transform 1 0 3464 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_205
timestamp 1598358358
transform 1 0 3336 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_786
timestamp 1598358358
transform 1 0 3464 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_204
timestamp 1598358358
transform -1 0 3464 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_60
timestamp 1598358358
transform 1 0 3080 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_69
timestamp 1598358358
transform -1 0 3208 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_203
timestamp 1598358358
transform 1 0 3272 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_215
timestamp 1598358358
transform -1 0 3272 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_61
timestamp 1598358358
transform 1 0 3144 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_201
timestamp 1598358358
transform 1 0 3272 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_206
timestamp 1598358358
transform -1 0 3272 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_84
timestamp 1598358358
transform 1 0 3080 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_316
timestamp 1598358358
transform -1 0 3080 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_412
timestamp 1598358358
transform -1 0 3016 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_32
timestamp 1598358358
transform -1 0 2952 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_81
timestamp 1598358358
transform -1 0 3080 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_49
timestamp 1598358358
transform 1 0 2888 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_68
timestamp 1598358358
transform -1 0 3016 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_58
timestamp 1598358358
transform 1 0 2824 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_416
timestamp 1598358358
transform -1 0 2824 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_234
timestamp 1598358358
transform -1 0 2760 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_92
timestamp 1598358358
transform 1 0 2632 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_415
timestamp 1598358358
transform 1 0 2824 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_825
timestamp 1598358358
transform 1 0 2760 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_412
timestamp 1598358358
transform 1 0 2696 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_416
timestamp 1598358358
transform 1 0 2632 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_640
timestamp 1598358358
transform -1 0 2568 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_650
timestamp 1598358358
transform -1 0 2504 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_97
timestamp 1598358358
transform -1 0 2568 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_89
timestamp 1598358358
transform 1 0 2568 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_119
timestamp 1598358358
transform -1 0 2632 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_46
timestamp 1598358358
transform 1 0 2440 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_520
timestamp 1598358358
transform -1 0 2376 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_642
timestamp 1598358358
transform -1 0 2248 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_87
timestamp 1598358358
transform 1 0 2312 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_519
timestamp 1598358358
transform -1 0 2440 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_518
timestamp 1598358358
transform 1 0 2248 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_29
timestamp 1598358358
transform 1 0 2376 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_19
timestamp 1598358358
transform -1 0 2312 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_129
timestamp 1598358358
transform -1 0 2248 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_655
timestamp 1598358358
transform 1 0 2120 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_649
timestamp 1598358358
transform 1 0 2056 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_641
timestamp 1598358358
transform 1 0 1992 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_660
timestamp 1598358358
transform -1 0 2184 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_662
timestamp 1598358358
transform 1 0 2056 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_224
timestamp 1598358358
transform 1 0 1992 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_341
timestamp 1598358358
transform -1 0 1992 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_350
timestamp 1598358358
transform -1 0 1928 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_219
timestamp 1598358358
transform 1 0 1800 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_643
timestamp 1598358358
transform 1 0 1736 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_227
timestamp 1598358358
transform 1 0 1928 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_231
timestamp 1598358358
transform -1 0 1800 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_226
timestamp 1598358358
transform 1 0 1864 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_229
timestamp 1598358358
transform -1 0 1864 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_222
timestamp 1598358358
transform -1 0 1672 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_476
timestamp 1598358358
transform -1 0 1608 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_215
timestamp 1598358358
transform -1 0 1736 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_406
timestamp 1598358358
transform 1 0 1672 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_230
timestamp 1598358358
transform -1 0 1672 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_65
timestamp 1598358358
transform -1 0 1608 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_479
timestamp 1598358358
transform -1 0 1544 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_785
timestamp 1598358358
transform -1 0 1480 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_795
timestamp 1598358358
transform -1 0 1416 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_318
timestamp 1598358358
transform -1 0 1352 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_206
timestamp 1598358358
transform 1 0 1480 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_201
timestamp 1598358358
transform -1 0 1480 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_202
timestamp 1598358358
transform 1 0 1288 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_316
timestamp 1598358358
transform -1 0 1416 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_776
timestamp 1598358358
transform 1 0 1224 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_841
timestamp 1598358358
transform -1 0 1224 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_831
timestamp 1598358358
transform 1 0 1096 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_68
timestamp 1598358358
transform 1 0 1160 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_69
timestamp 1598358358
transform 1 0 1224 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_238
timestamp 1598358358
transform 1 0 1096 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_716
timestamp 1598358358
transform 1 0 904 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_804
timestamp 1598358358
transform -1 0 904 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_851
timestamp 1598358358
transform -1 0 1032 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_840
timestamp 1598358358
transform -1 0 968 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_273
timestamp 1598358358
transform -1 0 1096 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_300
timestamp 1598358358
transform -1 0 1032 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_153
timestamp 1598358358
transform -1 0 1096 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_310
timestamp 1598358358
transform -1 0 904 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_794
timestamp 1598358358
transform 1 0 776 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_301
timestamp 1598358358
transform -1 0 776 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_605
timestamp 1598358358
transform 1 0 648 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_590
timestamp 1598358358
transform 1 0 712 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_718
timestamp 1598358358
transform -1 0 712 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_591
timestamp 1598358358
transform 1 0 776 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_335
timestamp 1598358358
transform -1 0 584 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_787
timestamp 1598358358
transform 1 0 392 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_808
timestamp 1598358358
transform -1 0 648 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_370
timestamp 1598358358
transform -1 0 456 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_604
timestamp 1598358358
transform -1 0 648 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_369
timestamp 1598358358
transform -1 0 520 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_603
timestamp 1598358358
transform 1 0 520 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_309
timestamp 1598358358
transform -1 0 520 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_181
timestamp 1598358358
transform 1 0 264 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_543
timestamp 1598358358
transform 1 0 328 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_542
timestamp 1598358358
transform -1 0 328 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_552
timestamp 1598358358
transform -1 0 264 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_315
timestamp 1598358358
transform 1 0 328 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_179
timestamp 1598358358
transform 1 0 200 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_192
timestamp 1598358358
transform -1 0 72 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_564
timestamp 1598358358
transform -1 0 72 0 -1 1810
box -16 -6 80 210
use OR2X1  OR2X1_742
timestamp 1598358358
transform -1 0 200 0 1 1810
box -16 -6 80 210
use OR2X1  OR2X1_191
timestamp 1598358358
transform -1 0 136 0 1 1810
box -16 -6 80 210
use AND2X1  AND2X1_189
timestamp 1598358358
transform -1 0 200 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_178
timestamp 1598358358
transform -1 0 136 0 -1 1810
box -16 -6 80 210
use AND2X1  AND2X1_579
timestamp 1598358358
transform 1 0 5512 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_575
timestamp 1598358358
transform 1 0 5448 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_501
timestamp 1598358358
transform -1 0 5448 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_239
timestamp 1598358358
transform 1 0 5192 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_574
timestamp 1598358358
transform 1 0 5320 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_506
timestamp 1598358358
transform 1 0 5256 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_500
timestamp 1598358358
transform 1 0 5128 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_497
timestamp 1598358358
transform -1 0 5000 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_242
timestamp 1598358358
transform -1 0 5128 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_842
timestamp 1598358358
transform 1 0 5000 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_184
timestamp 1598358358
transform 1 0 4808 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_226
timestamp 1598358358
transform -1 0 4808 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_502
timestamp 1598358358
transform 1 0 4872 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_227
timestamp 1598358358
transform 1 0 4680 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_103
timestamp 1598358358
transform -1 0 4616 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_107
timestamp 1598358358
transform -1 0 4488 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_844
timestamp 1598358358
transform 1 0 4616 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_560
timestamp 1598358358
transform -1 0 4552 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_529
timestamp 1598358358
transform 1 0 4232 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_113
timestamp 1598358358
transform -1 0 4424 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_553
timestamp 1598358358
transform -1 0 4360 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_134
timestamp 1598358358
transform -1 0 4104 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_361
timestamp 1598358358
transform 1 0 4168 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_768
timestamp 1598358358
transform -1 0 4168 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_541
timestamp 1598358358
transform 1 0 3976 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_132
timestamp 1598358358
transform 1 0 3912 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_137
timestamp 1598358358
transform -1 0 3912 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_139
timestamp 1598358358
transform 1 0 3784 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_245
timestamp 1598358358
transform 1 0 3656 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_265
timestamp 1598358358
transform -1 0 3656 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_130
timestamp 1598358358
transform -1 0 3784 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_267
timestamp 1598358358
transform -1 0 3592 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_72
timestamp 1598358358
transform -1 0 3528 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_262
timestamp 1598358358
transform 1 0 3400 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_87
timestamp 1598358358
transform 1 0 3336 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_129
timestamp 1598358358
transform -1 0 3272 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_393
timestamp 1598358358
transform -1 0 3208 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_80
timestamp 1598358358
transform -1 0 3144 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_202
timestamp 1598358358
transform 1 0 3272 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_83
timestamp 1598358358
transform 1 0 2952 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_394
timestamp 1598358358
transform -1 0 2952 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_400
timestamp 1598358358
transform -1 0 3080 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_414
timestamp 1598358358
transform -1 0 2888 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_82
timestamp 1598358358
transform 1 0 2760 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_42
timestamp 1598358358
transform -1 0 2760 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_96
timestamp 1598358358
transform -1 0 2696 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_98
timestamp 1598358358
transform -1 0 2632 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_99
timestamp 1598358358
transform -1 0 2504 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_93
timestamp 1598358358
transform 1 0 2504 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_606
timestamp 1598358358
transform 1 0 2376 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_656
timestamp 1598358358
transform -1 0 2312 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_607
timestamp 1598358358
transform 1 0 2312 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_88
timestamp 1598358358
transform -1 0 2248 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_101
timestamp 1598358358
transform 1 0 2120 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_559
timestamp 1598358358
transform -1 0 2056 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_517
timestamp 1598358358
transform -1 0 2120 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_340
timestamp 1598358358
transform -1 0 1992 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_264
timestamp 1598358358
transform -1 0 1864 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_218
timestamp 1598358358
transform -1 0 1800 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_265
timestamp 1598358358
transform 1 0 1864 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_327
timestamp 1598358358
transform -1 0 1736 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_216
timestamp 1598358358
transform 1 0 1608 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_475
timestamp 1598358358
transform -1 0 1608 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_734
timestamp 1598358358
transform -1 0 1544 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_473
timestamp 1598358358
transform 1 0 1352 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_493
timestamp 1598358358
transform -1 0 1352 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_492
timestamp 1598358358
transform -1 0 1480 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_778
timestamp 1598358358
transform 1 0 1096 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_491
timestamp 1598358358
transform 1 0 1224 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_371
timestamp 1598358358
transform -1 0 1224 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_717
timestamp 1598358358
transform -1 0 968 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_723
timestamp 1598358358
transform -1 0 904 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_372
timestamp 1598358358
transform -1 0 1096 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_272
timestamp 1598358358
transform -1 0 1032 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_458
timestamp 1598358358
transform -1 0 776 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_722
timestamp 1598358358
transform 1 0 648 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_674
timestamp 1598358358
transform -1 0 840 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_733
timestamp 1598358358
transform -1 0 648 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_737
timestamp 1598358358
transform -1 0 584 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_741
timestamp 1598358358
transform -1 0 520 0 1 1410
box -16 -6 80 210
use AND2X1  AND2X1_74
timestamp 1598358358
transform 1 0 392 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_457
timestamp 1598358358
transform -1 0 392 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_464
timestamp 1598358358
transform -1 0 328 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_471
timestamp 1598358358
transform -1 0 264 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_565
timestamp 1598358358
transform -1 0 72 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_190
timestamp 1598358358
transform -1 0 200 0 1 1410
box -16 -6 80 210
use OR2X1  OR2X1_540
timestamp 1598358358
transform -1 0 136 0 1 1410
box -16 -6 80 210
use FILL  FILL_7_4
timestamp 1598358358
transform -1 0 5576 0 -1 1410
box -16 -6 32 210
use AND2X1  AND2X1_735
timestamp 1598358358
transform -1 0 5512 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_573
timestamp 1598358358
transform 1 0 5384 0 -1 1410
box -16 -6 80 210
use FILL  FILL_7_3
timestamp 1598358358
transform -1 0 5560 0 -1 1410
box -16 -6 32 210
use FILL  FILL_7_2
timestamp 1598358358
transform -1 0 5544 0 -1 1410
box -16 -6 32 210
use FILL  FILL_7_1
timestamp 1598358358
transform -1 0 5528 0 -1 1410
box -16 -6 32 210
use OR2X1  OR2X1_528
timestamp 1598358358
transform 1 0 5256 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_657
timestamp 1598358358
transform 1 0 5320 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_510
timestamp 1598358358
transform 1 0 5192 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_508
timestamp 1598358358
transform -1 0 5192 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_503
timestamp 1598358358
transform 1 0 4936 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_474
timestamp 1598358358
transform 1 0 5064 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_509
timestamp 1598358358
transform 1 0 5000 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_488
timestamp 1598358358
transform -1 0 4808 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_487
timestamp 1598358358
transform -1 0 4744 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_456
timestamp 1598358358
transform 1 0 4872 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_570
timestamp 1598358358
transform 1 0 4808 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_489
timestamp 1598358358
transform -1 0 4680 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_558
timestamp 1598358358
transform -1 0 4616 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_576
timestamp 1598358358
transform 1 0 4488 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_571
timestamp 1598358358
transform 1 0 4424 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_561
timestamp 1598358358
transform 1 0 4360 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_563
timestamp 1598358358
transform 1 0 4296 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_557
timestamp 1598358358
transform 1 0 4232 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_572
timestamp 1598358358
transform 1 0 4168 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_554
timestamp 1598358358
transform -1 0 4168 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_772
timestamp 1598358358
transform -1 0 4104 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_140
timestamp 1598358358
transform 1 0 3976 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_217
timestamp 1598358358
transform -1 0 3976 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_141
timestamp 1598358358
transform 1 0 3848 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_656
timestamp 1598358358
transform 1 0 3784 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_131
timestamp 1598358358
transform 1 0 3720 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_118
timestamp 1598358358
transform -1 0 3720 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_266
timestamp 1598358358
transform 1 0 3592 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_249
timestamp 1598358358
transform -1 0 3592 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_88
timestamp 1598358358
transform 1 0 3400 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_119
timestamp 1598358358
transform 1 0 3336 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_340
timestamp 1598358358
transform -1 0 3528 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_277
timestamp 1598358358
transform -1 0 3272 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_126
timestamp 1598358358
transform -1 0 3208 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_633
timestamp 1598358358
transform -1 0 3336 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_398
timestamp 1598358358
transform -1 0 3144 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_399
timestamp 1598358358
transform -1 0 3080 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_403
timestamp 1598358358
transform -1 0 3016 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_404
timestamp 1598358358
transform 1 0 2888 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_397
timestamp 1598358358
transform 1 0 2696 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_402
timestamp 1598358358
transform 1 0 2824 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_94
timestamp 1598358358
transform 1 0 2760 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_611
timestamp 1598358358
transform 1 0 2632 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_610
timestamp 1598358358
transform 1 0 2504 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_646
timestamp 1598358358
transform 1 0 2440 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_612
timestamp 1598358358
transform 1 0 2568 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_647
timestamp 1598358358
transform -1 0 2376 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_100
timestamp 1598358358
transform 1 0 2184 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_80
timestamp 1598358358
transform -1 0 2440 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_609
timestamp 1598358358
transform 1 0 2248 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_608
timestamp 1598358358
transform 1 0 2120 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_502
timestamp 1598358358
transform 1 0 2056 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_503
timestamp 1598358358
transform -1 0 2056 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_509
timestamp 1598358358
transform -1 0 1992 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_510
timestamp 1598358358
transform -1 0 1800 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_505
timestamp 1598358358
transform -1 0 1928 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_504
timestamp 1598358358
transform -1 0 1864 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_507
timestamp 1598358358
transform -1 0 1736 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_508
timestamp 1598358358
transform 1 0 1544 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_239
timestamp 1598358358
transform 1 0 1608 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_242
timestamp 1598358358
transform 1 0 1480 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_506
timestamp 1598358358
transform 1 0 1416 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_130
timestamp 1598358358
transform 1 0 1352 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_67
timestamp 1598358358
transform 1 0 1288 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_121
timestamp 1598358358
transform 1 0 1224 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_241
timestamp 1598358358
transform -1 0 1224 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_274
timestamp 1598358358
transform 1 0 1096 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_120
timestamp 1598358358
transform -1 0 1096 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_188
timestamp 1598358358
transform -1 0 1032 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_541
timestamp 1598358358
transform -1 0 904 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_255
timestamp 1598358358
transform -1 0 968 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_719
timestamp 1598358358
transform -1 0 712 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_666
timestamp 1598358358
transform -1 0 840 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_237
timestamp 1598358358
transform -1 0 776 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_675
timestamp 1598358358
transform -1 0 648 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_76
timestamp 1598358358
transform -1 0 520 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_445
timestamp 1598358358
transform -1 0 456 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_75
timestamp 1598358358
transform 1 0 520 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_455
timestamp 1598358358
transform -1 0 392 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_465
timestamp 1598358358
transform 1 0 200 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_368
timestamp 1598358358
transform 1 0 264 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_569
timestamp 1598358358
transform 1 0 8 0 -1 1410
box -16 -6 80 210
use OR2X1  OR2X1_553
timestamp 1598358358
transform -1 0 136 0 -1 1410
box -16 -6 80 210
use AND2X1  AND2X1_183
timestamp 1598358358
transform -1 0 200 0 -1 1410
box -16 -6 80 210
use FILL  FILL_6_4
timestamp 1598358358
transform 1 0 5560 0 1 1010
box -16 -6 32 210
use OR2X1  OR2X1_613
timestamp 1598358358
transform 1 0 5448 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_507
timestamp 1598358358
transform -1 0 5448 0 1 1010
box -16 -6 80 210
use FILL  FILL_6_3
timestamp 1598358358
transform 1 0 5544 0 1 1010
box -16 -6 32 210
use FILL  FILL_6_2
timestamp 1598358358
transform 1 0 5528 0 1 1010
box -16 -6 32 210
use FILL  FILL_6_1
timestamp 1598358358
transform 1 0 5512 0 1 1010
box -16 -6 32 210
use OR2X1  OR2X1_505
timestamp 1598358358
transform 1 0 5256 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_504
timestamp 1598358358
transform 1 0 5128 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_806
timestamp 1598358358
transform 1 0 5320 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_858
timestamp 1598358358
transform 1 0 5192 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_860
timestamp 1598358358
transform 1 0 5064 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_120
timestamp 1598358358
transform 1 0 5000 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_850
timestamp 1598358358
transform -1 0 5000 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_279
timestamp 1598358358
transform -1 0 4872 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_288
timestamp 1598358358
transform -1 0 4936 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_849
timestamp 1598358358
transform 1 0 4744 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_244
timestamp 1598358358
transform 1 0 4680 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_89
timestamp 1598358358
transform 1 0 4488 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_284
timestamp 1598358358
transform 1 0 4616 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_362
timestamp 1598358358
transform -1 0 4616 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_97
timestamp 1598358358
transform -1 0 4488 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_122
timestamp 1598358358
transform -1 0 4296 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_66
timestamp 1598358358
transform -1 0 4424 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_121
timestamp 1598358358
transform -1 0 4360 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_106
timestamp 1598358358
transform -1 0 4232 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_67
timestamp 1598358358
transform -1 0 4040 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_124
timestamp 1598358358
transform -1 0 4168 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_123
timestamp 1598358358
transform 1 0 4040 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_117
timestamp 1598358358
transform 1 0 3912 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_490
timestamp 1598358358
transform 1 0 3848 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_100
timestamp 1598358358
transform 1 0 3784 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_86
timestamp 1598358358
transform 1 0 3720 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_263
timestamp 1598358358
transform -1 0 3720 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_71
timestamp 1598358358
transform -1 0 3656 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_92
timestamp 1598358358
transform 1 0 3528 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_63
timestamp 1598358358
transform -1 0 3528 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_607
timestamp 1598358358
transform -1 0 3400 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_606
timestamp 1598358358
transform -1 0 3464 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_609
timestamp 1598358358
transform 1 0 3208 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_23
timestamp 1598358358
transform 1 0 3144 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_29
timestamp 1598358358
transform 1 0 3080 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_646
timestamp 1598358358
transform -1 0 3336 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_395
timestamp 1598358358
transform -1 0 3080 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_396
timestamp 1598358358
transform -1 0 3016 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_415
timestamp 1598358358
transform -1 0 2952 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_548
timestamp 1598358358
transform -1 0 2760 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_240
timestamp 1598358358
transform -1 0 2696 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_401
timestamp 1598358358
transform -1 0 2888 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_530
timestamp 1598358358
transform -1 0 2824 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_633
timestamp 1598358358
transform -1 0 2504 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_232
timestamp 1598358358
transform -1 0 2632 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_6
timestamp 1598358358
transform -1 0 2568 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_786
timestamp 1598358358
transform -1 0 2312 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_49
timestamp 1598358358
transform -1 0 2440 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_118
timestamp 1598358358
transform 1 0 2312 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_81
timestamp 1598358358
transform -1 0 2248 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_123
timestamp 1598358358
transform 1 0 1992 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_262
timestamp 1598358358
transform 1 0 2120 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_117
timestamp 1598358358
transform -1 0 2120 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_124
timestamp 1598358358
transform -1 0 1928 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_205
timestamp 1598358358
transform -1 0 1864 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_667
timestamp 1598358358
transform 1 0 1928 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_122
timestamp 1598358358
transform 1 0 1736 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_217
timestamp 1598358358
transform -1 0 1736 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_66
timestamp 1598358358
transform -1 0 1672 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_116
timestamp 1598358358
transform 1 0 1544 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_115
timestamp 1598358358
transform 1 0 1480 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_276
timestamp 1598358358
transform 1 0 1288 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_131
timestamp 1598358358
transform 1 0 1416 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_625
timestamp 1598358358
transform -1 0 1416 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_275
timestamp 1598358358
transform -1 0 1288 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_495
timestamp 1598358358
transform -1 0 1224 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_496
timestamp 1598358358
transform 1 0 1096 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_833
timestamp 1598358358
transform -1 0 968 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_628
timestamp 1598358358
transform -1 0 1096 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_498
timestamp 1598358358
transform 1 0 968 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_626
timestamp 1598358358
transform 1 0 840 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_203
timestamp 1598358358
transform 1 0 648 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_256
timestamp 1598358358
transform -1 0 840 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_268
timestamp 1598358358
transform -1 0 776 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_269
timestamp 1598358358
transform -1 0 648 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_271
timestamp 1598358358
transform -1 0 584 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_482
timestamp 1598358358
transform 1 0 456 0 1 1010
box -16 -6 80 210
use AND2X1  AND2X1_252
timestamp 1598358358
transform -1 0 456 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_578
timestamp 1598358358
transform 1 0 328 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_367
timestamp 1598358358
transform -1 0 328 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_270
timestamp 1598358358
transform 1 0 200 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_577
timestamp 1598358358
transform 1 0 8 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_456
timestamp 1598358358
transform -1 0 200 0 1 1010
box -16 -6 80 210
use OR2X1  OR2X1_549
timestamp 1598358358
transform -1 0 136 0 1 1010
box -16 -6 80 210
use FILL  FILL_5_4
timestamp 1598358358
transform -1 0 5576 0 -1 1010
box -16 -6 32 210
use AND2X1  AND2X1_807
timestamp 1598358358
transform -1 0 5512 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_861
timestamp 1598358358
transform 1 0 5384 0 -1 1010
box -16 -6 80 210
use FILL  FILL_5_3
timestamp 1598358358
transform -1 0 5560 0 -1 1010
box -16 -6 32 210
use FILL  FILL_5_2
timestamp 1598358358
transform -1 0 5544 0 -1 1010
box -16 -6 32 210
use FILL  FILL_5_1
timestamp 1598358358
transform -1 0 5528 0 -1 1010
box -16 -6 32 210
use OR2X1  OR2X1_482
timestamp 1598358358
transform 1 0 5128 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_865
timestamp 1598358358
transform -1 0 5384 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_862
timestamp 1598358358
transform 1 0 5256 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_719
timestamp 1598358358
transform 1 0 5192 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_666
timestamp 1598358358
transform 1 0 5064 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_283
timestamp 1598358358
transform -1 0 5064 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_843
timestamp 1598358358
transform 1 0 4936 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_669
timestamp 1598358358
transform 1 0 4680 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_286
timestamp 1598358358
transform -1 0 4936 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_287
timestamp 1598358358
transform 1 0 4808 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_859
timestamp 1598358358
transform 1 0 4744 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_667
timestamp 1598358358
transform 1 0 4424 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_668
timestamp 1598358358
transform 1 0 4616 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_721
timestamp 1598358358
transform 1 0 4552 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_720
timestamp 1598358358
transform 1 0 4488 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_250
timestamp 1598358358
transform -1 0 4360 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_251
timestamp 1598358358
transform 1 0 4232 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_105
timestamp 1598358358
transform -1 0 4424 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_625
timestamp 1598358358
transform 1 0 4104 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_343
timestamp 1598358358
transform -1 0 4232 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_392
timestamp 1598358358
transform 1 0 4040 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_845
timestamp 1598358358
transform -1 0 4040 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_85
timestamp 1598358358
transform -1 0 3848 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_99
timestamp 1598358358
transform 1 0 3912 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_101
timestamp 1598358358
transform -1 0 3912 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_821
timestamp 1598358358
transform -1 0 3784 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_813
timestamp 1598358358
transform 1 0 3656 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_235
timestamp 1598358358
transform -1 0 3656 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_243
timestamp 1598358358
transform -1 0 3592 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_278
timestamp 1598358358
transform 1 0 3464 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_291
timestamp 1598358358
transform -1 0 3464 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_608
timestamp 1598358358
transform -1 0 3400 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_612
timestamp 1598358358
transform 1 0 3144 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_611
timestamp 1598358358
transform 1 0 3080 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_610
timestamp 1598358358
transform 1 0 3272 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_647
timestamp 1598358358
transform 1 0 3208 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_143
timestamp 1598358358
transform 1 0 3016 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_4
timestamp 1598358358
transform -1 0 3016 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_414
timestamp 1598358358
transform 1 0 2888 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_243
timestamp 1598358358
transform 1 0 2632 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_55
timestamp 1598358358
transform -1 0 2888 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_73
timestamp 1598358358
transform 1 0 2760 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_529
timestamp 1598358358
transform -1 0 2760 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_126
timestamp 1598358358
transform -1 0 2632 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_235
timestamp 1598358358
transform 1 0 2504 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_86
timestamp 1598358358
transform -1 0 2504 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_398
timestamp 1598358358
transform -1 0 2440 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_84
timestamp 1598358358
transform -1 0 2376 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_204
timestamp 1598358358
transform -1 0 2248 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_133
timestamp 1598358358
transform -1 0 2312 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_266
timestamp 1598358358
transform -1 0 2184 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_63
timestamp 1598358358
transform 1 0 2056 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_10
timestamp 1598358358
transform -1 0 2056 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_139
timestamp 1598358358
transform -1 0 1992 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_267
timestamp 1598358358
transform -1 0 1928 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_572
timestamp 1598358358
transform 1 0 1800 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_657
timestamp 1598358358
transform 1 0 1736 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_141
timestamp 1598358358
transform 1 0 1672 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_244
timestamp 1598358358
transform -1 0 1672 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_150
timestamp 1598358358
transform -1 0 1608 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_140
timestamp 1598358358
transform 1 0 1480 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_361
timestamp 1598358358
transform -1 0 1480 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_574
timestamp 1598358358
transform -1 0 1416 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_631
timestamp 1598358358
transform -1 0 1352 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_632
timestamp 1598358358
transform -1 0 1288 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_554
timestamp 1598358358
transform -1 0 1224 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_499
timestamp 1598358358
transform -1 0 1160 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_630
timestamp 1598358358
transform 1 0 1032 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_296
timestamp 1598358358
transform -1 0 1032 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_629
timestamp 1598358358
transform 1 0 904 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_627
timestamp 1598358358
transform 1 0 840 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_294
timestamp 1598358358
transform -1 0 840 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_247
timestamp 1598358358
transform -1 0 776 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_72
timestamp 1598358358
transform -1 0 712 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_664
timestamp 1598358358
transform -1 0 584 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_483
timestamp 1598358358
transform -1 0 520 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_556
timestamp 1598358358
transform -1 0 456 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_665
timestamp 1598358358
transform 1 0 584 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_254
timestamp 1598358358
transform -1 0 328 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_344
timestamp 1598358358
transform -1 0 264 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_253
timestamp 1598358358
transform -1 0 392 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_570
timestamp 1598358358
transform -1 0 72 0 -1 1010
box -16 -6 80 210
use OR2X1  OR2X1_563
timestamp 1598358358
transform -1 0 136 0 -1 1010
box -16 -6 80 210
use AND2X1  AND2X1_531
timestamp 1598358358
transform -1 0 200 0 -1 1010
box -16 -6 80 210
use FILL  FILL_4_4
timestamp 1598358358
transform 1 0 5560 0 1 610
box -16 -6 32 210
use AND2X1  AND2X1_630
timestamp 1598358358
transform 1 0 5448 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_623
timestamp 1598358358
transform 1 0 5384 0 1 610
box -16 -6 80 210
use FILL  FILL_4_3
timestamp 1598358358
transform 1 0 5544 0 1 610
box -16 -6 32 210
use FILL  FILL_4_2
timestamp 1598358358
transform 1 0 5528 0 1 610
box -16 -6 32 210
use FILL  FILL_4_1
timestamp 1598358358
transform 1 0 5512 0 1 610
box -16 -6 32 210
use AND2X1  AND2X1_632
timestamp 1598358358
transform -1 0 5384 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_185
timestamp 1598358358
transform -1 0 5320 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_631
timestamp 1598358358
transform 1 0 5192 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_483
timestamp 1598358358
transform -1 0 5192 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_628
timestamp 1598358358
transform 1 0 5064 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_556
timestamp 1598358358
transform -1 0 5064 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_790
timestamp 1598358358
transform 1 0 4936 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_754
timestamp 1598358358
transform 1 0 4872 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_615
timestamp 1598358358
transform 1 0 4808 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_753
timestamp 1598358358
transform 1 0 4744 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_614
timestamp 1598358358
transform 1 0 4680 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_366
timestamp 1598358358
transform -1 0 4680 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_367
timestamp 1598358358
transform 1 0 4552 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_359
timestamp 1598358358
transform 1 0 4488 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_344
timestamp 1598358358
transform -1 0 4488 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_494
timestamp 1598358358
transform 1 0 4360 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_294
timestamp 1598358358
transform 1 0 4296 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_247
timestamp 1598358358
transform -1 0 4296 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_248
timestamp 1598358358
transform -1 0 4232 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_255
timestamp 1598358358
transform 1 0 4040 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_256
timestamp 1598358358
transform 1 0 3976 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_349
timestamp 1598358358
transform 1 0 4104 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_102
timestamp 1598358358
transform 1 0 3912 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_10
timestamp 1598358358
transform 1 0 3784 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_342
timestamp 1598358358
transform 1 0 3848 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_150
timestamp 1598358358
transform 1 0 3720 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_246
timestamp 1598358358
transform -1 0 3720 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_822
timestamp 1598358358
transform -1 0 3656 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_835
timestamp 1598358358
transform -1 0 3592 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_232
timestamp 1598358358
transform 1 0 3400 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_234
timestamp 1598358358
transform 1 0 3336 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_240
timestamp 1598358358
transform 1 0 3464 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_233
timestamp 1598358358
transform 1 0 3272 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_62
timestamp 1598358358
transform -1 0 3272 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_38
timestamp 1598358358
transform 1 0 3144 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_15
timestamp 1598358358
transform -1 0 3144 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_293
timestamp 1598358358
transform -1 0 3080 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_671
timestamp 1598358358
transform -1 0 3016 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_8
timestamp 1598358358
transform 1 0 2888 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_672
timestamp 1598358358
transform 1 0 2824 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_102
timestamp 1598358358
transform -1 0 2824 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_277
timestamp 1598358358
transform 1 0 2696 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_90
timestamp 1598358358
transform -1 0 2696 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_673
timestamp 1598358358
transform -1 0 2632 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_104
timestamp 1598358358
transform -1 0 2568 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_85
timestamp 1598358358
transform -1 0 2504 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_38
timestamp 1598358358
transform -1 0 2440 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_394
timestamp 1598358358
transform -1 0 2376 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_399
timestamp 1598358358
transform 1 0 2248 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_813
timestamp 1598358358
transform -1 0 2248 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_845
timestamp 1598358358
transform -1 0 2120 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_263
timestamp 1598358358
transform 1 0 2120 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_132
timestamp 1598358358
transform -1 0 2056 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_137
timestamp 1598358358
transform 1 0 1928 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_721
timestamp 1598358358
transform 1 0 1800 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_720
timestamp 1598358358
transform 1 0 1736 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_134
timestamp 1598358358
transform 1 0 1864 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_668
timestamp 1598358358
transform 1 0 1608 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_669
timestamp 1598358358
transform 1 0 1672 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_521
timestamp 1598358358
transform -1 0 1608 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_523
timestamp 1598358358
transform -1 0 1544 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_114
timestamp 1598358358
transform 1 0 1288 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_522
timestamp 1598358358
transform 1 0 1416 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_107
timestamp 1598358358
transform -1 0 1416 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_71
timestamp 1598358358
transform -1 0 1288 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_497
timestamp 1598358358
transform 1 0 1160 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_159
timestamp 1598358358
transform -1 0 1160 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_500
timestamp 1598358358
transform -1 0 1096 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_501
timestamp 1598358358
transform -1 0 1032 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_735
timestamp 1598358358
transform -1 0 968 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_128
timestamp 1598358358
transform 1 0 840 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_127
timestamp 1598358358
transform 1 0 776 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_248
timestamp 1598358358
transform 1 0 712 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_297
timestamp 1598358358
transform -1 0 712 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_736
timestamp 1598358358
transform -1 0 648 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_295
timestamp 1598358358
transform 1 0 520 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_292
timestamp 1598358358
transform 1 0 456 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_184
timestamp 1598358358
transform -1 0 456 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_830
timestamp 1598358358
transform 1 0 328 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_279
timestamp 1598358358
transform 1 0 264 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_481
timestamp 1598358358
transform -1 0 264 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_562
timestamp 1598358358
transform -1 0 72 0 1 610
box -16 -6 80 210
use OR2X1  OR2X1_555
timestamp 1598358358
transform -1 0 136 0 1 610
box -16 -6 80 210
use AND2X1  AND2X1_257
timestamp 1598358358
transform -1 0 200 0 1 610
box -16 -6 80 210
use FILL  FILL_3_4
timestamp 1598358358
transform -1 0 5576 0 -1 610
box -16 -6 32 210
use OR2X1  OR2X1_617
timestamp 1598358358
transform 1 0 5384 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_629
timestamp 1598358358
transform 1 0 5448 0 -1 610
box -16 -6 80 210
use FILL  FILL_3_3
timestamp 1598358358
transform -1 0 5560 0 -1 610
box -16 -6 32 210
use FILL  FILL_3_2
timestamp 1598358358
transform -1 0 5544 0 -1 610
box -16 -6 32 210
use FILL  FILL_3_1
timestamp 1598358358
transform -1 0 5528 0 -1 610
box -16 -6 32 210
use OR2X1  OR2X1_626
timestamp 1598358358
transform -1 0 5384 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_252
timestamp 1598358358
transform -1 0 5320 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_627
timestamp 1598358358
transform 1 0 5192 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_254
timestamp 1598358358
transform -1 0 5192 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_253
timestamp 1598358358
transform 1 0 5064 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_816
timestamp 1598358358
transform -1 0 5064 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_698
timestamp 1598358358
transform -1 0 5000 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_282
timestamp 1598358358
transform -1 0 4872 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_281
timestamp 1598358358
transform -1 0 4744 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_562
timestamp 1598358358
transform -1 0 4936 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_285
timestamp 1598358358
transform 1 0 4744 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_292
timestamp 1598358358
transform -1 0 4680 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_384
timestamp 1598358358
transform -1 0 4552 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_383
timestamp 1598358358
transform -1 0 4616 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_360
timestamp 1598358358
transform -1 0 4488 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_363
timestamp 1598358358
transform -1 0 4424 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_348
timestamp 1598358358
transform 1 0 4296 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_391
timestamp 1598358358
transform -1 0 4296 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_225
timestamp 1598358358
transform 1 0 4168 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_127
timestamp 1598358358
transform -1 0 4168 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_125
timestamp 1598358358
transform 1 0 3976 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_128
timestamp 1598358358
transform 1 0 4040 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_93
timestamp 1598358358
transform 1 0 3848 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_6
timestamp 1598358358
transform 1 0 3784 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_98
timestamp 1598358358
transform 1 0 3912 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_670
timestamp 1598358358
transform 1 0 3656 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_823
timestamp 1598358358
transform -1 0 3656 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_673
timestamp 1598358358
transform 1 0 3720 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_836
timestamp 1598358358
transform -1 0 3592 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_824
timestamp 1598358358
transform -1 0 3464 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_619
timestamp 1598358358
transform 1 0 3336 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_839
timestamp 1598358358
transform -1 0 3528 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_618
timestamp 1598358358
transform 1 0 3208 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_9
timestamp 1598358358
transform -1 0 3336 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_852
timestamp 1598358358
transform -1 0 3208 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_62
timestamp 1598358358
transform -1 0 3144 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_143
timestamp 1598358358
transform 1 0 3016 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_37
timestamp 1598358358
transform -1 0 3016 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_819
timestamp 1598358358
transform 1 0 2888 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_622
timestamp 1598358358
transform -1 0 2760 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_621
timestamp 1598358358
transform 1 0 2632 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_618
timestamp 1598358358
transform -1 0 2888 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_619
timestamp 1598358358
transform -1 0 2824 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_670
timestamp 1598358358
transform -1 0 2632 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_616
timestamp 1598358358
transform 1 0 2504 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_617
timestamp 1598358358
transform 1 0 2440 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_400
timestamp 1598358358
transform -1 0 2312 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_403
timestamp 1598358358
transform -1 0 2248 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_83
timestamp 1598358358
transform -1 0 2440 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_393
timestamp 1598358358
transform -1 0 2376 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_404
timestamp 1598358358
transform -1 0 2120 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_79
timestamp 1598358358
transform 1 0 2120 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_15
timestamp 1598358358
transform 1 0 1992 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_768
timestamp 1598358358
transform -1 0 1928 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_663
timestamp 1598358358
transform -1 0 1864 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_659
timestamp 1598358358
transform 1 0 1736 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_103
timestamp 1598358358
transform -1 0 1992 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_624
timestamp 1598358358
transform 1 0 1672 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_474
timestamp 1598358358
transform 1 0 1608 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_849
timestamp 1598358358
transform -1 0 1608 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_658
timestamp 1598358358
transform 1 0 1480 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_560
timestamp 1598358358
transform 1 0 1416 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_844
timestamp 1598358358
transform 1 0 1352 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_113
timestamp 1598358358
transform -1 0 1352 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_249
timestamp 1598358358
transform 1 0 1096 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_106
timestamp 1598358358
transform -1 0 1288 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_595
timestamp 1598358358
transform 1 0 1160 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_575
timestamp 1598358358
transform 1 0 1032 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_573
timestamp 1598358358
transform 1 0 968 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_245
timestamp 1598358358
transform -1 0 968 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_246
timestamp 1598358358
transform -1 0 904 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_342
timestamp 1598358358
transform 1 0 776 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_360
timestamp 1598358358
transform 1 0 648 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_125
timestamp 1598358358
transform 1 0 712 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_347
timestamp 1598358358
transform 1 0 584 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_346
timestamp 1598358358
transform 1 0 520 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_842
timestamp 1598358358
transform 1 0 392 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_108
timestamp 1598358358
transform -1 0 520 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_284
timestamp 1598358358
transform 1 0 328 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_280
timestamp 1598358358
transform 1 0 264 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_258
timestamp 1598358358
transform -1 0 264 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_756
timestamp 1598358358
transform -1 0 72 0 -1 610
box -16 -6 80 210
use OR2X1  OR2X1_259
timestamp 1598358358
transform -1 0 200 0 -1 610
box -16 -6 80 210
use AND2X1  AND2X1_757
timestamp 1598358358
transform -1 0 136 0 -1 610
box -16 -6 80 210
use FILL  FILL_2_4
timestamp 1598358358
transform 1 0 5560 0 1 210
box -16 -6 32 210
use OR2X1  OR2X1_616
timestamp 1598358358
transform 1 0 5448 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_756
timestamp 1598358358
transform -1 0 5448 0 1 210
box -16 -6 80 210
use FILL  FILL_2_3
timestamp 1598358358
transform 1 0 5544 0 1 210
box -16 -6 32 210
use FILL  FILL_2_2
timestamp 1598358358
transform 1 0 5528 0 1 210
box -16 -6 32 210
use FILL  FILL_2_1
timestamp 1598358358
transform 1 0 5512 0 1 210
box -16 -6 32 210
use OR2X1  OR2X1_665
timestamp 1598358358
transform -1 0 5192 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_758
timestamp 1598358358
transform 1 0 5320 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_805
timestamp 1598358358
transform -1 0 5320 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_664
timestamp 1598358358
transform -1 0 5256 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_815
timestamp 1598358358
transform -1 0 5064 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_814
timestamp 1598358358
transform -1 0 5128 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_846
timestamp 1598358358
transform -1 0 5000 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_258
timestamp 1598358358
transform -1 0 4872 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_295
timestamp 1598358358
transform -1 0 4744 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_793
timestamp 1598358358
transform 1 0 4872 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_709
timestamp 1598358358
transform -1 0 4808 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_257
timestamp 1598358358
transform 1 0 4488 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_346
timestamp 1598358358
transform 1 0 4616 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_259
timestamp 1598358358
transform 1 0 4552 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_296
timestamp 1598358358
transform -1 0 4488 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_236
timestamp 1598358358
transform 1 0 4360 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_55
timestamp 1598358358
transform 1 0 4296 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_818
timestamp 1598358358
transform -1 0 4296 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_382
timestamp 1598358358
transform 1 0 4168 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_381
timestamp 1598358358
transform 1 0 4104 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_699
timestamp 1598358358
transform 1 0 4040 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_260
timestamp 1598358358
transform -1 0 4040 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_77
timestamp 1598358358
transform 1 0 3912 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_90
timestamp 1598358358
transform 1 0 3848 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_133
timestamp 1598358358
transform 1 0 3784 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_73
timestamp 1598358358
transform 1 0 3720 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_672
timestamp 1598358358
transform 1 0 3656 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_96
timestamp 1598358358
transform 1 0 3592 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_159
timestamp 1598358358
transform 1 0 3528 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_54
timestamp 1598358358
transform 1 0 3464 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_9
timestamp 1598358358
transform -1 0 3464 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_94
timestamp 1598358358
transform 1 0 3336 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_42
timestamp 1598358358
transform 1 0 3272 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_827
timestamp 1598358358
transform -1 0 3272 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_28
timestamp 1598358358
transform 1 0 3144 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_14
timestamp 1598358358
transform 1 0 3080 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_5
timestamp 1598358358
transform 1 0 3016 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_818
timestamp 1598358358
transform 1 0 2888 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_820
timestamp 1598358358
transform 1 0 2952 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_278
timestamp 1598358358
transform -1 0 2888 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_77
timestamp 1598358358
transform 1 0 2760 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_82
timestamp 1598358358
transform -1 0 2760 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_397
timestamp 1598358358
transform 1 0 2632 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_402
timestamp 1598358358
transform 1 0 2568 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_78
timestamp 1598358358
transform -1 0 2568 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_490
timestamp 1598358358
transform -1 0 2504 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_401
timestamp 1598358358
transform 1 0 2312 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_765
timestamp 1598358358
transform -1 0 2440 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_766
timestamp 1598358358
transform 1 0 2248 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_395
timestamp 1598358358
transform 1 0 2184 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_396
timestamp 1598358358
transform 1 0 2120 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_767
timestamp 1598358358
transform -1 0 2120 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_488
timestamp 1598358358
transform -1 0 2056 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_814
timestamp 1598358358
transform -1 0 1928 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_487
timestamp 1598358358
transform 1 0 1928 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_815
timestamp 1598358358
transform -1 0 1864 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_816
timestamp 1598358358
transform -1 0 1800 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_861
timestamp 1598358358
transform 1 0 1672 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_392
timestamp 1598358358
transform -1 0 1672 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_860
timestamp 1598358358
transform 1 0 1544 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_576
timestamp 1598358358
transform -1 0 1544 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_571
timestamp 1598358358
transform 1 0 1416 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_105
timestamp 1598358358
transform -1 0 1416 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_579
timestamp 1598358358
transform -1 0 1352 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_343
timestamp 1598358358
transform -1 0 1160 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_251
timestamp 1598358358
transform -1 0 1288 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_250
timestamp 1598358358
transform -1 0 1224 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_843
timestamp 1598358358
transform -1 0 1096 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_858
timestamp 1598358358
transform 1 0 968 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_850
timestamp 1598358358
transform 1 0 904 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_349
timestamp 1598358358
transform -1 0 904 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_359
timestamp 1598358358
transform -1 0 840 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_362
timestamp 1598358358
transform -1 0 776 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_363
timestamp 1598358358
transform -1 0 712 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_366
timestamp 1598358358
transform -1 0 648 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_287
timestamp 1598358358
transform -1 0 456 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_283
timestamp 1598358358
transform -1 0 584 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_755
timestamp 1598358358
transform -1 0 520 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_348
timestamp 1598358358
transform 1 0 200 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_281
timestamp 1598358358
transform -1 0 392 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_282
timestamp 1598358358
transform -1 0 328 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_260
timestamp 1598358358
transform -1 0 200 0 1 210
box -16 -6 80 210
use OR2X1  OR2X1_345
timestamp 1598358358
transform 1 0 72 0 1 210
box -16 -6 80 210
use AND2X1  AND2X1_261
timestamp 1598358358
transform 1 0 8 0 1 210
box -16 -6 80 210
use FILL  FILL_1_4
timestamp 1598358358
transform -1 0 5576 0 -1 210
box -16 -6 32 210
use AND2X1  AND2X1_866
timestamp 1598358358
transform 1 0 5448 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_191
timestamp 1598358358
transform 1 0 5384 0 -1 210
box -16 -6 80 210
use FILL  FILL_1_3
timestamp 1598358358
transform -1 0 5560 0 -1 210
box -16 -6 32 210
use FILL  FILL_1_2
timestamp 1598358358
transform -1 0 5544 0 -1 210
box -16 -6 32 210
use FILL  FILL_1_1
timestamp 1598358358
transform -1 0 5528 0 -1 210
box -16 -6 32 210
use OR2X1  OR2X1_187
timestamp 1598358358
transform 1 0 5320 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_663
timestamp 1598358358
transform 1 0 5256 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_580
timestamp 1598358358
transform 1 0 5192 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_621
timestamp 1598358358
transform -1 0 5192 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_757
timestamp 1598358358
transform -1 0 5000 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_624
timestamp 1598358358
transform -1 0 5128 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_620
timestamp 1598358358
transform 1 0 5000 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_755
timestamp 1598358358
transform -1 0 4936 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_759
timestamp 1598358358
transform -1 0 4744 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_791
timestamp 1598358358
transform -1 0 4872 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_792
timestamp 1598358358
transform 1 0 4744 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_297
timestamp 1598358358
transform 1 0 4424 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_711
timestamp 1598358358
transform -1 0 4680 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_848
timestamp 1598358358
transform -1 0 4616 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_347
timestamp 1598358358
transform 1 0 4488 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_701
timestamp 1598358358
transform -1 0 4360 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_700
timestamp 1598358358
transform 1 0 4232 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_710
timestamp 1598358358
transform 1 0 4360 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_481
timestamp 1598358358
transform -1 0 4232 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_261
timestamp 1598358358
transform 1 0 3976 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_345
timestamp 1598358358
transform 1 0 4104 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_555
timestamp 1598358358
transform -1 0 4104 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_817
timestamp 1598358358
transform -1 0 3976 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_820
timestamp 1598358358
transform 1 0 3784 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_847
timestamp 1598358358
transform -1 0 3912 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_748
timestamp 1598358358
transform -1 0 3784 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_751
timestamp 1598358358
transform 1 0 3592 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_789
timestamp 1598358358
transform -1 0 3720 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_750
timestamp 1598358358
transform -1 0 3592 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_819
timestamp 1598358358
transform 1 0 3464 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_749
timestamp 1598358358
transform 1 0 3400 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_825
timestamp 1598358358
transform -1 0 3400 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_826
timestamp 1598358358
transform -1 0 3336 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_104
timestamp 1598358358
transform 1 0 3080 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_837
timestamp 1598358358
transform -1 0 3272 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_838
timestamp 1598358358
transform -1 0 3208 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_671
timestamp 1598358358
transform 1 0 3016 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_8
timestamp 1598358358
transform 1 0 2952 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_37
timestamp 1598358358
transform 1 0 2888 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_28
timestamp 1598358358
transform 1 0 2824 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_54
timestamp 1598358358
transform -1 0 2824 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_14
timestamp 1598358358
transform -1 0 2760 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_5
timestamp 1598358358
transform -1 0 2696 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_4
timestamp 1598358358
transform -1 0 2632 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_381
timestamp 1598358358
transform -1 0 2568 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_817
timestamp 1598358358
transform -1 0 2504 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_847
timestamp 1598358358
transform -1 0 2440 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_770
timestamp 1598358358
transform -1 0 2376 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_771
timestamp 1598358358
transform -1 0 2312 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_236
timestamp 1598358358
transform -1 0 2248 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_774
timestamp 1598358358
transform -1 0 2120 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_773
timestamp 1598358358
transform 1 0 1992 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_382
timestamp 1598358358
transform -1 0 2184 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_489
timestamp 1598358358
transform -1 0 1992 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_772
timestamp 1598358358
transform 1 0 1864 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_864
timestamp 1598358358
transform -1 0 1864 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_557
timestamp 1598358358
transform -1 0 1800 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_846
timestamp 1598358358
transform -1 0 1736 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_391
timestamp 1598358358
transform 1 0 1608 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_848
timestamp 1598358358
transform -1 0 1608 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_866
timestamp 1598358358
transform 1 0 1480 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_865
timestamp 1598358358
transform 1 0 1416 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_859
timestamp 1598358358
transform -1 0 1416 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_810
timestamp 1598358358
transform -1 0 1352 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_862
timestamp 1598358358
transform 1 0 1224 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_561
timestamp 1598358358
transform 1 0 1160 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_558
timestamp 1598358358
transform 1 0 1096 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_383
timestamp 1598358358
transform 1 0 840 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_225
timestamp 1598358358
transform -1 0 1096 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_494
timestamp 1598358358
transform 1 0 968 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_384
timestamp 1598358358
transform 1 0 904 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_812
timestamp 1598358358
transform 1 0 776 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_811
timestamp 1598358358
transform 1 0 712 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_805
timestamp 1598358358
transform -1 0 712 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_807
timestamp 1598358358
transform 1 0 584 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_806
timestamp 1598358358
transform -1 0 584 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_580
timestamp 1598358358
transform -1 0 520 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_288
timestamp 1598358358
transform 1 0 392 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_286
timestamp 1598358358
transform 1 0 328 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_285
timestamp 1598358358
transform 1 0 264 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_758
timestamp 1598358358
transform -1 0 264 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_792
timestamp 1598358358
transform 1 0 72 0 -1 210
box -16 -6 80 210
use OR2X1  OR2X1_791
timestamp 1598358358
transform -1 0 72 0 -1 210
box -16 -6 80 210
use AND2X1  AND2X1_759
timestamp 1598358358
transform -1 0 200 0 -1 210
box -16 -6 80 210
<< labels >>
rlabel metal2 s 2784 -40 2784 -40 8 INPUT_0
port 0 nsew
rlabel metal2 s 2944 -40 2944 -40 8 D_INPUT_0
port 1 nsew
rlabel metal2 s 2816 -40 2816 -40 8 INPUT_1
port 2 nsew
rlabel metal2 s 2496 -40 2496 -40 8 D_INPUT_1
port 3 nsew
rlabel metal2 s 3136 -40 3136 -40 8 INPUT_2
port 4 nsew
rlabel metal2 s 2720 -40 2720 -40 8 D_INPUT_2
port 5 nsew
rlabel metal2 s 2672 -40 2672 -40 8 INPUT_3
port 6 nsew
rlabel metal2 s 2752 -40 2752 -40 8 D_INPUT_3
port 7 nsew
rlabel metal2 s 2560 4080 2560 4080 6 INPUT_4
port 8 nsew
rlabel metal2 s 2000 4080 2000 4080 6 D_INPUT_4
port 9 nsew
rlabel metal2 s 1968 4080 1968 4080 6 INPUT_5
port 10 nsew
rlabel metal2 s 2288 4080 2288 4080 6 D_INPUT_5
port 11 nsew
rlabel metal2 s 1536 4080 1536 4080 6 INPUT_6
port 12 nsew
rlabel metal2 s 2464 4080 2464 4080 6 D_INPUT_6
port 13 nsew
rlabel metal2 s 2160 4080 2160 4080 6 INPUT_7
port 14 nsew
rlabel metal2 s 2096 4080 2096 4080 6 D_INPUT_7
port 15 nsew
rlabel metal3 s -48 2120 -48 2120 4 D_GATE_222
port 16 nsew
rlabel metal3 s -48 1100 -48 1100 4 D_GATE_366
port 17 nsew
rlabel metal2 s 608 4080 608 4080 6 D_GATE_479
port 18 nsew
rlabel metal2 s 448 -40 448 -40 8 D_GATE_579
port 19 nsew
rlabel metal2 s 1856 -40 1856 -40 8 D_GATE_662
port 20 nsew
rlabel metal3 s -48 1900 -48 1900 4 D_GATE_741
port 21 nsew
rlabel metal2 s 832 -40 832 -40 8 D_GATE_811
port 22 nsew
rlabel metal2 s 1536 -40 1536 -40 8 D_GATE_865
port 23 nsew
rlabel metal3 s 5632 2620 5632 2620 6 GATE_222
port 24 nsew
rlabel metal2 s 4704 -40 4704 -40 8 GATE_366
port 25 nsew
rlabel metal3 s 5632 2580 5632 2580 6 GATE_479
port 26 nsew
rlabel metal3 s 5632 220 5632 220 6 GATE_579
port 27 nsew
rlabel metal3 s 5632 320 5632 320 6 GATE_662
port 28 nsew
rlabel metal3 s 5632 3120 5632 3120 6 GATE_741
port 29 nsew
rlabel metal3 s 5632 2980 5632 2980 6 GATE_811
port 30 nsew
rlabel metal3 s 5632 180 5632 180 6 GATE_865
port 31 nsew
rlabel metal2 s 3696 -40 3696 -40 8 gate
port 32 nsew
rlabel metal3 s 5632 3880 5632 3880 6 type:
port 33 nsew
rlabel metal2 s 4992 4080 4992 4080 6 AND;
port 34 nsew
rlabel metal2 s 4560 4080 4560 4080 6 name:
port 35 nsew
rlabel metal2 s 928 -40 928 -40 8 GATE_0_I0
port 36 nsew
rlabel space -412 -43 5994 4083 1 vdd
rlabel space -412 -43 5994 4083 1 gnd
<< end >>
