*** TEST 009 ***
*
* ngSPICE test for PLS experiments
*
* dynamic NAND (positive) gate (not a standard cell (!!!) - it's a pseudo cell) under PLS
*
* Author: Jan Belohoubek, 04/2019
* jan.belohoubek@fit.cvut.cz
*
* https://users.fit.cvut.cz/~belohja4/
*
*
* **************************************

.include ../models.lib
.include ../tsmc180nmcmos.lib

* **************************************
* --- Test ---
* **************************************

* --- Settings
.param showPlots = 1
* redefine ...
.include test00X_settings.inc
.csparam showPlots = {showPlots}
.global showPlots
* --- End of Settins

Vtrig LaserTrig 0 0 PWL(0ns 0V 40ns 0V 42ns SUPP 62ns SUPP 64ns 0V 100ns 0V)
*Vtrig LaserTrig 0 0V

.global LaserTrig 

* --- outputs
*R1 VSS out 1000000
C1 VSS out 1pF


*
* 2-input NOR Gate
*
.subckt dynamicNANDp Y VSS A B CLK VDD beamDistanceTop = 0 beamDistanceBot = 0

Xpmos1 Y A VDD VDD VSS LaserTrig SUBCKT_PMOS beamDistance = beamDistanceTop ch_w=2u ch_l=0.2u mos_ad=1.2p mos_pd=5.2u mos_as=2p mos_ps=10u
Xpmos2 VDD B Y VDD VSS LaserTrig SUBCKT_PMOS beamDistance = beamDistanceTop ch_w=2u ch_l=0.2u mos_ad=0p mos_pd=0u mos_as=0p mos_ps=0u

Xnmos1 Y CLK VSS VSS LaserTrig SUBCKT_NMOS beamDistance = beamDistanceBot ch_w=1u ch_l=0.2u mos_ad=0.6p mos_pd=3.2u mos_as=1.32p mos_ps=9.2u

C1 VSS Y 0.09fF
C2 Y B 0.10fF
C3 VSS A 0.05fF
C4 Y A 0.08fF
C5 Y VDD 0.57fF
C6 B A 0.22fF
C7 B VDD 0.27fF
C8 A VDD 0.20fF
C9 VSS VSS 0.17fF
C10 Y VSS 0.11fF
C11 B VSS 0.19fF
C12 A VSS 0.25fF
C13 VDD VSS 1.73fF

.ends


* --- circuit layout model
xNOR out VSS A B CLK VDD dynamicNANDp


* **************************************
* --- Simulation Settings ---
* **************************************

* --- inputs
*Vvin0 A 0 0 PWL(0ns 0V 20ns SUPP 22ns SUPP)
*Vvin1 B 0 0 PWL(0ns 0V 21ns SUPP 23ns SUPP)

* precharge to 0
VvCK CLK 0 0 PWL(0ns SUPP 15ns SUPP 17ns 0V)
* open pull-down transistor
*VvCK CLK 0 0 PWL(0ns SUPP 15ns SUPP 17ns SUPP)

.tran 0.1ns 100ns
.param SIMSTEP = '100ns/0.1ns'
.csparam SIMSTEP = {SIMSTEP}

* **************************************
* --- Simulation Control ---
* **************************************

.control
    run
    
    if ('showPlots' > 0)
      plot i(vvdd) i(vvss)
      plot v(vss) v(vdd) v(LaserTrig)
      plot v(A) v(B) v(CLK) v(out)
    end
    
    print '(i(vvdd)[length(i(vvdd)) - 1] + i(vvdd)[length(i(vvdd)) - 2])/2'
    print '(i(vvss)[length(i(vvss)) - 1] + i(vvss)[length(i(vvss)) - 2])/2'
    
    print i(vvdd)[length(i(vvdd))/2]
    print i(vvss)[length(i(vvss))/2]
    
    print v(out)[length(v(out))/2]
    
    if ('showPlots' < 1)
        quit
    end
    
.endc

.end
